// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18;

output N25612,N25598,N25616,N25591,N25601,N25613,N25617,N25610,N25607,N25618;

not NOT1 (N19, N2);
nand NAND3 (N20, N11, N15, N4);
nand NAND4 (N21, N15, N8, N8, N12);
xor XOR2 (N22, N2, N13);
nor NOR2 (N23, N13, N6);
or OR4 (N24, N21, N21, N16, N11);
xor XOR2 (N25, N15, N12);
and AND4 (N26, N1, N12, N8, N19);
buf BUF1 (N27, N12);
not NOT1 (N28, N13);
not NOT1 (N29, N18);
nand NAND4 (N30, N9, N10, N24, N17);
not NOT1 (N31, N30);
and AND4 (N32, N8, N20, N27, N14);
nor NOR4 (N33, N6, N31, N4, N27);
and AND3 (N34, N32, N11, N14);
buf BUF1 (N35, N22);
and AND4 (N36, N25, N22, N9, N29);
nor NOR3 (N37, N12, N22, N15);
nor NOR2 (N38, N36, N29);
xor XOR2 (N39, N4, N9);
not NOT1 (N40, N18);
nor NOR3 (N41, N23, N11, N12);
nand NAND2 (N42, N28, N34);
and AND4 (N43, N22, N26, N12, N12);
nor NOR3 (N44, N27, N23, N11);
and AND3 (N45, N40, N18, N30);
or OR3 (N46, N42, N37, N24);
buf BUF1 (N47, N2);
or OR2 (N48, N46, N25);
nor NOR2 (N49, N41, N31);
xor XOR2 (N50, N39, N40);
buf BUF1 (N51, N47);
or OR3 (N52, N35, N9, N2);
not NOT1 (N53, N48);
or OR3 (N54, N44, N11, N7);
or OR4 (N55, N51, N20, N38, N43);
or OR2 (N56, N2, N44);
or OR4 (N57, N17, N56, N14, N49);
or OR3 (N58, N16, N8, N9);
nor NOR3 (N59, N40, N29, N10);
not NOT1 (N60, N59);
and AND3 (N61, N60, N54, N12);
xor XOR2 (N62, N7, N61);
nor NOR2 (N63, N23, N60);
xor XOR2 (N64, N62, N26);
nand NAND4 (N65, N33, N8, N59, N44);
nor NOR4 (N66, N63, N2, N47, N33);
or OR4 (N67, N64, N50, N48, N41);
not NOT1 (N68, N17);
nand NAND2 (N69, N55, N53);
nor NOR3 (N70, N13, N45, N36);
xor XOR2 (N71, N9, N59);
or OR3 (N72, N70, N40, N14);
and AND4 (N73, N52, N11, N66, N67);
buf BUF1 (N74, N60);
nand NAND3 (N75, N68, N57, N26);
and AND3 (N76, N73, N48, N43);
or OR3 (N77, N74, N17, N27);
nor NOR2 (N78, N49, N34);
or OR3 (N79, N17, N12, N20);
nand NAND4 (N80, N58, N16, N50, N45);
buf BUF1 (N81, N71);
nor NOR3 (N82, N80, N6, N36);
buf BUF1 (N83, N75);
buf BUF1 (N84, N77);
nand NAND2 (N85, N78, N30);
nor NOR2 (N86, N69, N64);
xor XOR2 (N87, N82, N73);
and AND4 (N88, N72, N78, N5, N73);
not NOT1 (N89, N88);
buf BUF1 (N90, N89);
nor NOR4 (N91, N76, N31, N50, N69);
and AND2 (N92, N84, N65);
buf BUF1 (N93, N20);
xor XOR2 (N94, N92, N63);
nor NOR2 (N95, N90, N38);
not NOT1 (N96, N91);
or OR2 (N97, N85, N16);
xor XOR2 (N98, N83, N22);
buf BUF1 (N99, N95);
not NOT1 (N100, N96);
or OR4 (N101, N86, N83, N83, N53);
xor XOR2 (N102, N101, N65);
xor XOR2 (N103, N102, N46);
buf BUF1 (N104, N81);
and AND2 (N105, N99, N45);
not NOT1 (N106, N79);
nor NOR4 (N107, N100, N71, N85, N90);
and AND4 (N108, N107, N102, N31, N11);
or OR4 (N109, N87, N25, N46, N22);
and AND3 (N110, N103, N70, N33);
or OR4 (N111, N109, N22, N100, N64);
and AND3 (N112, N98, N15, N3);
and AND4 (N113, N106, N43, N7, N55);
buf BUF1 (N114, N108);
buf BUF1 (N115, N97);
xor XOR2 (N116, N113, N39);
or OR3 (N117, N110, N115, N18);
and AND4 (N118, N90, N99, N18, N82);
not NOT1 (N119, N94);
xor XOR2 (N120, N93, N107);
nor NOR4 (N121, N112, N18, N22, N59);
not NOT1 (N122, N104);
nand NAND2 (N123, N111, N104);
xor XOR2 (N124, N114, N88);
or OR3 (N125, N116, N110, N13);
or OR4 (N126, N122, N67, N119, N108);
buf BUF1 (N127, N74);
nor NOR2 (N128, N125, N114);
buf BUF1 (N129, N118);
and AND4 (N130, N120, N35, N2, N84);
nand NAND4 (N131, N121, N24, N86, N71);
or OR3 (N132, N124, N91, N90);
xor XOR2 (N133, N123, N110);
nor NOR2 (N134, N127, N86);
buf BUF1 (N135, N133);
and AND4 (N136, N130, N128, N132, N89);
xor XOR2 (N137, N37, N131);
or OR3 (N138, N101, N119, N20);
nand NAND2 (N139, N14, N40);
not NOT1 (N140, N105);
or OR4 (N141, N138, N115, N9, N46);
nand NAND4 (N142, N140, N106, N123, N70);
not NOT1 (N143, N117);
and AND4 (N144, N136, N112, N87, N113);
not NOT1 (N145, N134);
nor NOR3 (N146, N126, N75, N134);
xor XOR2 (N147, N145, N126);
nor NOR3 (N148, N135, N75, N123);
xor XOR2 (N149, N129, N64);
xor XOR2 (N150, N143, N140);
xor XOR2 (N151, N142, N42);
xor XOR2 (N152, N150, N40);
or OR2 (N153, N148, N135);
nor NOR3 (N154, N152, N81, N8);
or OR3 (N155, N153, N94, N39);
buf BUF1 (N156, N155);
nor NOR3 (N157, N154, N149, N131);
not NOT1 (N158, N113);
xor XOR2 (N159, N137, N69);
xor XOR2 (N160, N147, N135);
buf BUF1 (N161, N141);
buf BUF1 (N162, N151);
not NOT1 (N163, N158);
nand NAND2 (N164, N163, N43);
nor NOR4 (N165, N156, N56, N157, N4);
and AND4 (N166, N85, N24, N88, N161);
buf BUF1 (N167, N11);
xor XOR2 (N168, N162, N166);
buf BUF1 (N169, N77);
or OR3 (N170, N167, N4, N18);
buf BUF1 (N171, N164);
xor XOR2 (N172, N159, N112);
xor XOR2 (N173, N160, N34);
not NOT1 (N174, N165);
nor NOR4 (N175, N174, N106, N69, N98);
nand NAND3 (N176, N144, N146, N2);
nor NOR4 (N177, N133, N59, N85, N72);
nor NOR3 (N178, N139, N12, N97);
or OR4 (N179, N170, N100, N72, N89);
nor NOR2 (N180, N176, N175);
buf BUF1 (N181, N113);
or OR2 (N182, N177, N57);
nand NAND4 (N183, N168, N156, N79, N52);
or OR2 (N184, N180, N139);
xor XOR2 (N185, N181, N138);
not NOT1 (N186, N172);
or OR3 (N187, N171, N12, N111);
and AND3 (N188, N169, N68, N89);
nand NAND2 (N189, N182, N176);
and AND4 (N190, N184, N169, N130, N94);
xor XOR2 (N191, N190, N13);
xor XOR2 (N192, N187, N131);
or OR3 (N193, N186, N35, N75);
or OR2 (N194, N178, N13);
not NOT1 (N195, N183);
xor XOR2 (N196, N192, N169);
nand NAND4 (N197, N179, N76, N13, N77);
or OR3 (N198, N188, N91, N76);
and AND2 (N199, N173, N54);
buf BUF1 (N200, N199);
buf BUF1 (N201, N196);
nand NAND4 (N202, N198, N26, N126, N11);
xor XOR2 (N203, N193, N158);
buf BUF1 (N204, N194);
nor NOR4 (N205, N195, N187, N138, N22);
buf BUF1 (N206, N201);
xor XOR2 (N207, N185, N188);
not NOT1 (N208, N200);
not NOT1 (N209, N202);
or OR2 (N210, N207, N206);
or OR4 (N211, N13, N139, N144, N39);
buf BUF1 (N212, N209);
buf BUF1 (N213, N189);
xor XOR2 (N214, N210, N104);
nand NAND2 (N215, N205, N31);
buf BUF1 (N216, N212);
and AND2 (N217, N213, N153);
and AND3 (N218, N204, N102, N47);
buf BUF1 (N219, N208);
and AND3 (N220, N215, N215, N192);
xor XOR2 (N221, N211, N105);
not NOT1 (N222, N218);
nor NOR4 (N223, N219, N150, N221, N152);
or OR3 (N224, N213, N106, N164);
xor XOR2 (N225, N223, N197);
or OR2 (N226, N216, N138);
nor NOR2 (N227, N69, N58);
nor NOR2 (N228, N191, N126);
nand NAND2 (N229, N225, N93);
not NOT1 (N230, N203);
nand NAND3 (N231, N228, N163, N5);
nor NOR2 (N232, N222, N157);
nand NAND4 (N233, N227, N182, N131, N6);
or OR2 (N234, N214, N227);
nand NAND4 (N235, N231, N158, N152, N190);
not NOT1 (N236, N226);
or OR3 (N237, N230, N228, N127);
nor NOR4 (N238, N235, N115, N17, N78);
nor NOR3 (N239, N232, N87, N186);
and AND2 (N240, N233, N175);
not NOT1 (N241, N238);
nor NOR2 (N242, N220, N210);
xor XOR2 (N243, N224, N85);
xor XOR2 (N244, N234, N67);
nand NAND3 (N245, N229, N66, N104);
not NOT1 (N246, N244);
or OR4 (N247, N217, N183, N105, N104);
xor XOR2 (N248, N240, N170);
not NOT1 (N249, N246);
buf BUF1 (N250, N241);
nand NAND4 (N251, N249, N111, N18, N79);
not NOT1 (N252, N251);
buf BUF1 (N253, N247);
xor XOR2 (N254, N252, N101);
and AND4 (N255, N243, N122, N42, N18);
buf BUF1 (N256, N253);
nand NAND2 (N257, N248, N248);
nor NOR3 (N258, N239, N42, N131);
buf BUF1 (N259, N257);
and AND3 (N260, N245, N5, N90);
not NOT1 (N261, N237);
nor NOR2 (N262, N250, N11);
buf BUF1 (N263, N258);
or OR4 (N264, N263, N14, N93, N100);
or OR2 (N265, N255, N35);
nor NOR2 (N266, N254, N221);
not NOT1 (N267, N236);
xor XOR2 (N268, N267, N80);
not NOT1 (N269, N259);
nand NAND2 (N270, N261, N150);
and AND2 (N271, N242, N52);
or OR4 (N272, N256, N26, N35, N240);
or OR3 (N273, N271, N72, N219);
nor NOR4 (N274, N262, N168, N32, N71);
and AND4 (N275, N270, N268, N149, N190);
buf BUF1 (N276, N18);
nand NAND3 (N277, N266, N151, N157);
nand NAND2 (N278, N276, N120);
buf BUF1 (N279, N273);
nand NAND3 (N280, N278, N207, N262);
xor XOR2 (N281, N269, N38);
xor XOR2 (N282, N272, N191);
or OR3 (N283, N260, N60, N114);
or OR2 (N284, N282, N2);
not NOT1 (N285, N284);
or OR3 (N286, N275, N185, N164);
or OR3 (N287, N283, N5, N235);
and AND4 (N288, N280, N69, N101, N64);
nand NAND2 (N289, N285, N82);
nand NAND2 (N290, N264, N234);
buf BUF1 (N291, N289);
nor NOR4 (N292, N265, N119, N39, N234);
xor XOR2 (N293, N286, N2);
xor XOR2 (N294, N281, N197);
xor XOR2 (N295, N294, N92);
and AND2 (N296, N279, N234);
xor XOR2 (N297, N287, N157);
buf BUF1 (N298, N293);
xor XOR2 (N299, N290, N30);
nand NAND3 (N300, N298, N145, N189);
buf BUF1 (N301, N296);
nor NOR3 (N302, N301, N201, N180);
buf BUF1 (N303, N292);
xor XOR2 (N304, N299, N117);
nand NAND2 (N305, N303, N263);
or OR2 (N306, N304, N211);
nor NOR2 (N307, N295, N297);
nor NOR2 (N308, N20, N223);
nor NOR4 (N309, N300, N12, N146, N99);
buf BUF1 (N310, N274);
nand NAND4 (N311, N291, N291, N42, N232);
and AND4 (N312, N308, N168, N222, N55);
xor XOR2 (N313, N309, N296);
xor XOR2 (N314, N313, N118);
xor XOR2 (N315, N305, N105);
buf BUF1 (N316, N315);
nand NAND2 (N317, N306, N55);
nand NAND2 (N318, N312, N171);
not NOT1 (N319, N277);
or OR2 (N320, N319, N92);
xor XOR2 (N321, N302, N84);
xor XOR2 (N322, N320, N67);
nand NAND3 (N323, N317, N253, N301);
or OR3 (N324, N310, N21, N263);
nand NAND3 (N325, N323, N73, N323);
nand NAND2 (N326, N316, N234);
nor NOR4 (N327, N324, N203, N259, N157);
and AND2 (N328, N307, N174);
nand NAND4 (N329, N325, N55, N210, N70);
and AND3 (N330, N314, N88, N256);
nor NOR3 (N331, N288, N232, N233);
not NOT1 (N332, N327);
buf BUF1 (N333, N326);
or OR3 (N334, N328, N246, N107);
nor NOR2 (N335, N330, N6);
xor XOR2 (N336, N311, N166);
nor NOR2 (N337, N332, N284);
not NOT1 (N338, N329);
buf BUF1 (N339, N322);
xor XOR2 (N340, N336, N280);
buf BUF1 (N341, N335);
nor NOR3 (N342, N321, N232, N92);
not NOT1 (N343, N342);
nor NOR3 (N344, N333, N329, N204);
or OR3 (N345, N339, N314, N104);
not NOT1 (N346, N334);
nand NAND2 (N347, N340, N100);
and AND2 (N348, N346, N81);
buf BUF1 (N349, N331);
xor XOR2 (N350, N343, N68);
nand NAND3 (N351, N318, N334, N325);
nor NOR3 (N352, N350, N156, N114);
not NOT1 (N353, N351);
and AND3 (N354, N348, N219, N297);
and AND2 (N355, N353, N107);
buf BUF1 (N356, N341);
nor NOR2 (N357, N345, N356);
nor NOR3 (N358, N150, N179, N357);
or OR2 (N359, N167, N230);
not NOT1 (N360, N337);
buf BUF1 (N361, N355);
nor NOR3 (N362, N359, N71, N137);
nor NOR4 (N363, N338, N292, N48, N181);
and AND2 (N364, N358, N248);
buf BUF1 (N365, N352);
buf BUF1 (N366, N361);
not NOT1 (N367, N347);
or OR4 (N368, N367, N278, N298, N267);
and AND3 (N369, N362, N356, N72);
buf BUF1 (N370, N369);
nand NAND3 (N371, N366, N61, N160);
nor NOR4 (N372, N349, N367, N4, N33);
nand NAND3 (N373, N360, N122, N298);
not NOT1 (N374, N365);
and AND4 (N375, N371, N222, N278, N176);
or OR4 (N376, N363, N252, N135, N259);
or OR4 (N377, N344, N231, N311, N36);
nand NAND3 (N378, N373, N221, N14);
or OR4 (N379, N364, N78, N80, N310);
not NOT1 (N380, N378);
not NOT1 (N381, N377);
buf BUF1 (N382, N375);
and AND3 (N383, N382, N38, N249);
and AND2 (N384, N376, N28);
not NOT1 (N385, N374);
not NOT1 (N386, N379);
nor NOR2 (N387, N354, N54);
not NOT1 (N388, N384);
nor NOR2 (N389, N386, N175);
and AND2 (N390, N368, N42);
and AND2 (N391, N388, N231);
or OR2 (N392, N372, N170);
xor XOR2 (N393, N381, N30);
or OR2 (N394, N393, N365);
not NOT1 (N395, N387);
and AND3 (N396, N390, N167, N345);
or OR3 (N397, N395, N29, N79);
nor NOR2 (N398, N385, N161);
or OR3 (N399, N391, N104, N135);
not NOT1 (N400, N399);
nand NAND4 (N401, N383, N341, N355, N210);
and AND4 (N402, N380, N235, N350, N282);
and AND3 (N403, N398, N396, N175);
buf BUF1 (N404, N315);
not NOT1 (N405, N401);
and AND2 (N406, N392, N12);
xor XOR2 (N407, N406, N200);
xor XOR2 (N408, N394, N185);
and AND3 (N409, N408, N115, N45);
buf BUF1 (N410, N370);
not NOT1 (N411, N402);
nand NAND2 (N412, N407, N36);
xor XOR2 (N413, N410, N332);
nand NAND4 (N414, N397, N225, N126, N230);
buf BUF1 (N415, N403);
and AND3 (N416, N411, N293, N66);
buf BUF1 (N417, N389);
not NOT1 (N418, N400);
or OR3 (N419, N413, N87, N110);
buf BUF1 (N420, N414);
and AND2 (N421, N409, N72);
nor NOR2 (N422, N416, N330);
not NOT1 (N423, N405);
and AND2 (N424, N420, N115);
nor NOR3 (N425, N417, N93, N368);
or OR3 (N426, N421, N181, N76);
and AND4 (N427, N424, N46, N325, N115);
buf BUF1 (N428, N422);
and AND4 (N429, N418, N230, N221, N232);
nor NOR2 (N430, N427, N342);
buf BUF1 (N431, N415);
not NOT1 (N432, N429);
and AND3 (N433, N432, N409, N290);
buf BUF1 (N434, N430);
buf BUF1 (N435, N425);
buf BUF1 (N436, N426);
or OR2 (N437, N436, N272);
nor NOR4 (N438, N412, N396, N329, N337);
and AND3 (N439, N434, N94, N60);
nand NAND2 (N440, N435, N197);
nor NOR4 (N441, N440, N77, N235, N261);
or OR3 (N442, N404, N439, N333);
nand NAND3 (N443, N424, N310, N260);
buf BUF1 (N444, N423);
and AND4 (N445, N437, N346, N383, N346);
xor XOR2 (N446, N444, N370);
nor NOR3 (N447, N438, N360, N162);
not NOT1 (N448, N447);
nor NOR4 (N449, N433, N218, N294, N10);
nor NOR2 (N450, N428, N272);
nand NAND2 (N451, N419, N300);
nor NOR2 (N452, N431, N31);
not NOT1 (N453, N451);
or OR4 (N454, N452, N284, N87, N103);
or OR2 (N455, N448, N330);
nand NAND3 (N456, N450, N69, N209);
or OR4 (N457, N446, N305, N71, N179);
xor XOR2 (N458, N445, N121);
xor XOR2 (N459, N454, N236);
buf BUF1 (N460, N441);
or OR3 (N461, N456, N178, N364);
nor NOR4 (N462, N455, N239, N282, N443);
nand NAND3 (N463, N432, N71, N405);
and AND3 (N464, N453, N24, N216);
xor XOR2 (N465, N461, N131);
and AND2 (N466, N462, N276);
xor XOR2 (N467, N459, N272);
or OR4 (N468, N463, N315, N246, N300);
not NOT1 (N469, N468);
nor NOR2 (N470, N460, N415);
nor NOR2 (N471, N457, N398);
not NOT1 (N472, N471);
xor XOR2 (N473, N464, N184);
nor NOR3 (N474, N458, N9, N126);
or OR4 (N475, N473, N408, N412, N94);
nor NOR2 (N476, N475, N353);
or OR2 (N477, N465, N104);
and AND2 (N478, N472, N372);
not NOT1 (N479, N470);
xor XOR2 (N480, N469, N250);
xor XOR2 (N481, N476, N403);
nor NOR2 (N482, N466, N441);
or OR3 (N483, N467, N180, N412);
not NOT1 (N484, N478);
buf BUF1 (N485, N484);
buf BUF1 (N486, N474);
and AND2 (N487, N449, N120);
nand NAND3 (N488, N485, N420, N446);
and AND3 (N489, N480, N164, N270);
nand NAND2 (N490, N481, N2);
nor NOR4 (N491, N483, N339, N124, N286);
and AND2 (N492, N491, N151);
or OR2 (N493, N477, N87);
nand NAND4 (N494, N489, N311, N28, N45);
and AND4 (N495, N493, N348, N188, N73);
not NOT1 (N496, N488);
and AND2 (N497, N442, N238);
xor XOR2 (N498, N487, N378);
not NOT1 (N499, N492);
nor NOR3 (N500, N494, N162, N5);
buf BUF1 (N501, N497);
xor XOR2 (N502, N499, N201);
xor XOR2 (N503, N490, N20);
buf BUF1 (N504, N500);
buf BUF1 (N505, N498);
nor NOR3 (N506, N504, N281, N18);
and AND2 (N507, N495, N289);
nand NAND3 (N508, N486, N11, N155);
nor NOR2 (N509, N479, N287);
xor XOR2 (N510, N509, N350);
and AND3 (N511, N501, N333, N444);
or OR2 (N512, N510, N267);
xor XOR2 (N513, N505, N32);
xor XOR2 (N514, N512, N390);
not NOT1 (N515, N513);
buf BUF1 (N516, N503);
nand NAND3 (N517, N511, N345, N122);
xor XOR2 (N518, N506, N7);
nand NAND4 (N519, N482, N417, N231, N515);
xor XOR2 (N520, N116, N44);
buf BUF1 (N521, N514);
and AND4 (N522, N517, N498, N5, N379);
nor NOR3 (N523, N522, N294, N315);
and AND4 (N524, N502, N450, N353, N256);
nor NOR3 (N525, N523, N377, N126);
buf BUF1 (N526, N521);
not NOT1 (N527, N496);
nand NAND4 (N528, N508, N517, N197, N297);
or OR3 (N529, N524, N301, N99);
buf BUF1 (N530, N526);
buf BUF1 (N531, N525);
xor XOR2 (N532, N529, N301);
buf BUF1 (N533, N507);
and AND3 (N534, N532, N86, N449);
nand NAND3 (N535, N516, N175, N141);
xor XOR2 (N536, N531, N188);
or OR2 (N537, N519, N340);
nor NOR2 (N538, N528, N226);
or OR4 (N539, N533, N118, N169, N193);
and AND2 (N540, N536, N455);
or OR3 (N541, N518, N342, N342);
nor NOR4 (N542, N520, N243, N397, N526);
or OR3 (N543, N535, N413, N123);
nor NOR3 (N544, N540, N283, N258);
nor NOR4 (N545, N530, N325, N111, N207);
nor NOR4 (N546, N544, N259, N510, N318);
or OR4 (N547, N534, N99, N90, N248);
nor NOR4 (N548, N545, N86, N374, N31);
nor NOR2 (N549, N538, N400);
and AND2 (N550, N546, N483);
or OR2 (N551, N550, N437);
xor XOR2 (N552, N548, N15);
not NOT1 (N553, N552);
nand NAND3 (N554, N542, N390, N282);
nand NAND3 (N555, N537, N22, N388);
or OR3 (N556, N554, N296, N2);
and AND4 (N557, N551, N177, N300, N455);
or OR4 (N558, N553, N147, N105, N524);
xor XOR2 (N559, N527, N513);
or OR3 (N560, N547, N72, N493);
or OR2 (N561, N555, N359);
and AND2 (N562, N539, N386);
buf BUF1 (N563, N543);
not NOT1 (N564, N562);
nor NOR2 (N565, N559, N282);
or OR2 (N566, N558, N427);
or OR3 (N567, N549, N250, N358);
nor NOR4 (N568, N561, N140, N216, N260);
not NOT1 (N569, N566);
or OR4 (N570, N557, N243, N440, N508);
nand NAND2 (N571, N570, N272);
buf BUF1 (N572, N567);
or OR2 (N573, N556, N490);
or OR4 (N574, N565, N107, N260, N287);
and AND4 (N575, N571, N390, N421, N246);
nor NOR4 (N576, N563, N419, N321, N473);
or OR4 (N577, N564, N421, N18, N48);
or OR3 (N578, N575, N394, N2);
or OR2 (N579, N569, N303);
buf BUF1 (N580, N573);
nand NAND3 (N581, N579, N212, N580);
nand NAND2 (N582, N462, N206);
buf BUF1 (N583, N574);
nor NOR2 (N584, N577, N41);
or OR4 (N585, N541, N290, N223, N105);
not NOT1 (N586, N568);
nor NOR2 (N587, N582, N568);
and AND2 (N588, N585, N209);
buf BUF1 (N589, N572);
or OR4 (N590, N587, N99, N504, N300);
buf BUF1 (N591, N578);
or OR3 (N592, N581, N321, N215);
nor NOR4 (N593, N560, N157, N184, N182);
nor NOR3 (N594, N586, N5, N218);
xor XOR2 (N595, N592, N79);
buf BUF1 (N596, N589);
nand NAND4 (N597, N576, N336, N473, N430);
buf BUF1 (N598, N597);
and AND2 (N599, N584, N236);
not NOT1 (N600, N596);
not NOT1 (N601, N600);
nor NOR3 (N602, N595, N172, N41);
nor NOR4 (N603, N588, N408, N187, N53);
buf BUF1 (N604, N593);
and AND3 (N605, N604, N498, N579);
nor NOR3 (N606, N591, N73, N27);
buf BUF1 (N607, N599);
nor NOR2 (N608, N590, N85);
buf BUF1 (N609, N605);
buf BUF1 (N610, N608);
not NOT1 (N611, N594);
xor XOR2 (N612, N607, N492);
or OR3 (N613, N583, N527, N429);
not NOT1 (N614, N606);
not NOT1 (N615, N601);
nand NAND2 (N616, N603, N200);
xor XOR2 (N617, N612, N10);
nand NAND3 (N618, N613, N613, N506);
xor XOR2 (N619, N598, N359);
nand NAND3 (N620, N619, N564, N329);
buf BUF1 (N621, N602);
buf BUF1 (N622, N616);
nor NOR4 (N623, N614, N184, N376, N166);
nor NOR3 (N624, N623, N584, N61);
buf BUF1 (N625, N609);
not NOT1 (N626, N624);
not NOT1 (N627, N625);
not NOT1 (N628, N620);
buf BUF1 (N629, N628);
not NOT1 (N630, N626);
or OR2 (N631, N622, N150);
or OR3 (N632, N631, N132, N271);
nand NAND3 (N633, N621, N367, N400);
buf BUF1 (N634, N633);
or OR2 (N635, N617, N29);
not NOT1 (N636, N618);
or OR3 (N637, N634, N588, N341);
not NOT1 (N638, N629);
nand NAND2 (N639, N615, N331);
xor XOR2 (N640, N611, N574);
nor NOR2 (N641, N639, N542);
nand NAND3 (N642, N640, N31, N584);
nand NAND2 (N643, N636, N375);
or OR2 (N644, N627, N125);
buf BUF1 (N645, N641);
and AND2 (N646, N635, N636);
xor XOR2 (N647, N644, N273);
nand NAND2 (N648, N645, N76);
nor NOR2 (N649, N638, N382);
buf BUF1 (N650, N632);
nor NOR3 (N651, N649, N330, N25);
buf BUF1 (N652, N610);
not NOT1 (N653, N650);
buf BUF1 (N654, N646);
nor NOR3 (N655, N651, N17, N634);
nor NOR2 (N656, N643, N311);
buf BUF1 (N657, N656);
nor NOR3 (N658, N647, N31, N243);
and AND2 (N659, N653, N108);
buf BUF1 (N660, N630);
and AND4 (N661, N648, N242, N5, N114);
not NOT1 (N662, N659);
and AND2 (N663, N658, N606);
xor XOR2 (N664, N662, N493);
and AND2 (N665, N664, N629);
and AND2 (N666, N655, N10);
buf BUF1 (N667, N637);
or OR3 (N668, N652, N438, N559);
or OR4 (N669, N668, N99, N283, N632);
not NOT1 (N670, N661);
nand NAND4 (N671, N667, N565, N276, N318);
xor XOR2 (N672, N642, N52);
not NOT1 (N673, N665);
or OR2 (N674, N672, N407);
and AND2 (N675, N654, N93);
not NOT1 (N676, N671);
xor XOR2 (N677, N663, N124);
not NOT1 (N678, N669);
buf BUF1 (N679, N660);
nand NAND2 (N680, N676, N656);
not NOT1 (N681, N678);
xor XOR2 (N682, N675, N542);
buf BUF1 (N683, N679);
not NOT1 (N684, N680);
buf BUF1 (N685, N681);
nor NOR3 (N686, N670, N547, N492);
nor NOR2 (N687, N684, N91);
xor XOR2 (N688, N685, N395);
not NOT1 (N689, N682);
nor NOR4 (N690, N677, N409, N120, N147);
not NOT1 (N691, N686);
nor NOR4 (N692, N683, N23, N45, N534);
nor NOR2 (N693, N666, N636);
and AND2 (N694, N673, N434);
xor XOR2 (N695, N694, N400);
nor NOR3 (N696, N657, N433, N339);
nand NAND2 (N697, N689, N659);
xor XOR2 (N698, N691, N337);
nand NAND4 (N699, N692, N121, N220, N677);
and AND4 (N700, N688, N540, N595, N647);
and AND3 (N701, N674, N539, N151);
xor XOR2 (N702, N687, N567);
and AND3 (N703, N695, N340, N429);
buf BUF1 (N704, N696);
not NOT1 (N705, N693);
or OR4 (N706, N702, N286, N363, N527);
and AND3 (N707, N701, N35, N483);
not NOT1 (N708, N706);
buf BUF1 (N709, N700);
nor NOR3 (N710, N705, N191, N691);
xor XOR2 (N711, N690, N200);
or OR2 (N712, N711, N611);
buf BUF1 (N713, N712);
nor NOR3 (N714, N710, N552, N589);
or OR3 (N715, N698, N618, N360);
or OR4 (N716, N697, N513, N712, N1);
not NOT1 (N717, N715);
buf BUF1 (N718, N717);
not NOT1 (N719, N718);
xor XOR2 (N720, N708, N203);
buf BUF1 (N721, N713);
buf BUF1 (N722, N721);
not NOT1 (N723, N707);
or OR2 (N724, N716, N378);
and AND2 (N725, N703, N475);
and AND3 (N726, N719, N323, N365);
nor NOR3 (N727, N714, N453, N353);
xor XOR2 (N728, N726, N217);
xor XOR2 (N729, N725, N280);
or OR2 (N730, N729, N34);
xor XOR2 (N731, N699, N678);
not NOT1 (N732, N727);
xor XOR2 (N733, N722, N8);
nor NOR2 (N734, N723, N730);
or OR2 (N735, N38, N410);
or OR4 (N736, N724, N259, N210, N268);
or OR2 (N737, N734, N538);
not NOT1 (N738, N737);
or OR4 (N739, N720, N410, N518, N516);
nand NAND2 (N740, N732, N546);
and AND3 (N741, N739, N266, N622);
and AND4 (N742, N731, N525, N730, N23);
xor XOR2 (N743, N728, N279);
nor NOR3 (N744, N738, N556, N8);
nor NOR3 (N745, N704, N5, N598);
nand NAND2 (N746, N744, N278);
and AND2 (N747, N742, N406);
nor NOR3 (N748, N747, N486, N141);
not NOT1 (N749, N745);
buf BUF1 (N750, N740);
nor NOR4 (N751, N709, N700, N748, N357);
xor XOR2 (N752, N33, N36);
or OR2 (N753, N733, N641);
xor XOR2 (N754, N743, N401);
buf BUF1 (N755, N754);
and AND3 (N756, N735, N285, N33);
xor XOR2 (N757, N750, N548);
nand NAND4 (N758, N752, N648, N542, N730);
nor NOR2 (N759, N758, N253);
nor NOR3 (N760, N757, N226, N426);
nand NAND2 (N761, N746, N475);
and AND4 (N762, N751, N655, N149, N442);
and AND4 (N763, N755, N197, N352, N262);
not NOT1 (N764, N759);
or OR2 (N765, N762, N366);
or OR3 (N766, N764, N232, N126);
and AND3 (N767, N756, N475, N485);
and AND2 (N768, N765, N240);
nor NOR3 (N769, N741, N40, N374);
not NOT1 (N770, N769);
nand NAND2 (N771, N749, N107);
nand NAND3 (N772, N753, N699, N400);
nor NOR4 (N773, N772, N403, N531, N744);
nor NOR3 (N774, N770, N89, N200);
not NOT1 (N775, N774);
or OR4 (N776, N773, N389, N532, N359);
nor NOR4 (N777, N760, N171, N334, N479);
not NOT1 (N778, N777);
nand NAND2 (N779, N767, N675);
or OR4 (N780, N768, N150, N732, N217);
nor NOR4 (N781, N780, N186, N767, N625);
nand NAND4 (N782, N763, N160, N216, N405);
and AND4 (N783, N779, N466, N745, N20);
or OR4 (N784, N776, N702, N257, N238);
not NOT1 (N785, N771);
or OR3 (N786, N781, N69, N618);
or OR2 (N787, N784, N38);
not NOT1 (N788, N761);
nand NAND2 (N789, N788, N641);
not NOT1 (N790, N775);
or OR3 (N791, N787, N599, N182);
not NOT1 (N792, N766);
nor NOR2 (N793, N792, N506);
or OR2 (N794, N793, N222);
not NOT1 (N795, N783);
nor NOR2 (N796, N785, N474);
not NOT1 (N797, N790);
and AND3 (N798, N796, N358, N730);
buf BUF1 (N799, N797);
nand NAND3 (N800, N789, N543, N76);
not NOT1 (N801, N778);
or OR2 (N802, N786, N39);
nand NAND2 (N803, N802, N757);
xor XOR2 (N804, N801, N294);
nand NAND2 (N805, N798, N327);
xor XOR2 (N806, N804, N177);
not NOT1 (N807, N782);
not NOT1 (N808, N803);
not NOT1 (N809, N791);
xor XOR2 (N810, N800, N23);
not NOT1 (N811, N808);
not NOT1 (N812, N805);
and AND2 (N813, N806, N463);
buf BUF1 (N814, N811);
buf BUF1 (N815, N809);
nand NAND4 (N816, N815, N742, N736, N332);
buf BUF1 (N817, N257);
not NOT1 (N818, N812);
and AND3 (N819, N807, N712, N768);
xor XOR2 (N820, N813, N476);
not NOT1 (N821, N814);
and AND2 (N822, N821, N324);
buf BUF1 (N823, N818);
and AND4 (N824, N817, N434, N645, N106);
xor XOR2 (N825, N816, N327);
not NOT1 (N826, N825);
xor XOR2 (N827, N794, N186);
and AND2 (N828, N822, N373);
buf BUF1 (N829, N828);
or OR3 (N830, N795, N474, N171);
and AND4 (N831, N820, N396, N740, N136);
nand NAND3 (N832, N799, N55, N395);
xor XOR2 (N833, N827, N780);
xor XOR2 (N834, N826, N364);
and AND3 (N835, N819, N622, N84);
and AND3 (N836, N829, N593, N565);
nand NAND3 (N837, N836, N382, N824);
nand NAND2 (N838, N568, N339);
or OR3 (N839, N823, N750, N743);
xor XOR2 (N840, N837, N534);
xor XOR2 (N841, N830, N626);
buf BUF1 (N842, N833);
nor NOR4 (N843, N834, N161, N325, N238);
or OR3 (N844, N832, N146, N625);
and AND2 (N845, N841, N353);
xor XOR2 (N846, N845, N220);
xor XOR2 (N847, N846, N349);
xor XOR2 (N848, N835, N537);
and AND3 (N849, N843, N223, N573);
not NOT1 (N850, N844);
and AND2 (N851, N850, N384);
nand NAND3 (N852, N839, N81, N545);
and AND2 (N853, N847, N578);
xor XOR2 (N854, N838, N230);
and AND2 (N855, N810, N549);
nand NAND3 (N856, N851, N826, N721);
not NOT1 (N857, N855);
not NOT1 (N858, N831);
nand NAND3 (N859, N858, N833, N263);
nor NOR4 (N860, N853, N32, N177, N834);
not NOT1 (N861, N848);
and AND4 (N862, N860, N519, N136, N101);
nor NOR4 (N863, N862, N588, N370, N823);
xor XOR2 (N864, N854, N66);
nand NAND3 (N865, N842, N659, N658);
or OR3 (N866, N856, N239, N210);
nor NOR4 (N867, N866, N504, N572, N406);
nor NOR2 (N868, N849, N256);
or OR3 (N869, N868, N772, N517);
or OR3 (N870, N869, N15, N632);
xor XOR2 (N871, N861, N244);
nand NAND4 (N872, N870, N304, N389, N854);
nand NAND3 (N873, N865, N338, N279);
and AND2 (N874, N872, N515);
nand NAND4 (N875, N840, N314, N245, N138);
or OR4 (N876, N875, N42, N480, N838);
buf BUF1 (N877, N857);
nand NAND3 (N878, N874, N756, N700);
or OR2 (N879, N876, N774);
not NOT1 (N880, N871);
and AND3 (N881, N877, N858, N63);
buf BUF1 (N882, N864);
nand NAND2 (N883, N859, N665);
or OR3 (N884, N863, N39, N828);
buf BUF1 (N885, N882);
and AND2 (N886, N883, N376);
or OR3 (N887, N884, N241, N745);
xor XOR2 (N888, N886, N531);
xor XOR2 (N889, N888, N527);
or OR3 (N890, N889, N432, N885);
and AND3 (N891, N887, N631, N260);
nor NOR3 (N892, N668, N787, N507);
xor XOR2 (N893, N891, N488);
not NOT1 (N894, N892);
or OR3 (N895, N867, N761, N393);
xor XOR2 (N896, N878, N158);
or OR3 (N897, N890, N590, N416);
not NOT1 (N898, N897);
and AND3 (N899, N873, N682, N89);
or OR2 (N900, N879, N852);
and AND2 (N901, N580, N545);
or OR3 (N902, N899, N315, N481);
xor XOR2 (N903, N901, N85);
and AND2 (N904, N903, N143);
and AND2 (N905, N895, N599);
not NOT1 (N906, N880);
xor XOR2 (N907, N898, N180);
xor XOR2 (N908, N894, N697);
and AND2 (N909, N893, N837);
buf BUF1 (N910, N896);
and AND3 (N911, N904, N48, N694);
xor XOR2 (N912, N911, N371);
not NOT1 (N913, N902);
buf BUF1 (N914, N906);
or OR2 (N915, N909, N500);
or OR4 (N916, N912, N775, N645, N280);
nor NOR3 (N917, N908, N701, N425);
not NOT1 (N918, N917);
buf BUF1 (N919, N907);
xor XOR2 (N920, N881, N245);
and AND2 (N921, N900, N806);
nand NAND2 (N922, N914, N437);
xor XOR2 (N923, N915, N820);
nor NOR4 (N924, N905, N296, N881, N696);
and AND4 (N925, N918, N331, N629, N214);
nand NAND3 (N926, N923, N712, N215);
buf BUF1 (N927, N916);
nor NOR2 (N928, N920, N558);
and AND3 (N929, N925, N926, N541);
nor NOR2 (N930, N744, N572);
not NOT1 (N931, N921);
nor NOR4 (N932, N930, N87, N496, N172);
or OR2 (N933, N928, N610);
or OR4 (N934, N913, N910, N764, N793);
and AND2 (N935, N876, N749);
nor NOR4 (N936, N929, N784, N109, N826);
xor XOR2 (N937, N924, N617);
buf BUF1 (N938, N933);
nand NAND4 (N939, N922, N417, N198, N349);
buf BUF1 (N940, N919);
buf BUF1 (N941, N927);
nor NOR4 (N942, N939, N124, N599, N872);
nand NAND4 (N943, N942, N914, N612, N446);
xor XOR2 (N944, N941, N792);
nand NAND3 (N945, N934, N843, N52);
xor XOR2 (N946, N935, N861);
xor XOR2 (N947, N944, N358);
and AND4 (N948, N932, N15, N285, N199);
or OR3 (N949, N946, N644, N484);
and AND2 (N950, N948, N398);
nor NOR3 (N951, N947, N319, N300);
not NOT1 (N952, N937);
or OR3 (N953, N943, N839, N204);
nor NOR4 (N954, N938, N86, N286, N554);
nor NOR4 (N955, N949, N100, N669, N308);
not NOT1 (N956, N945);
and AND4 (N957, N936, N313, N399, N765);
nand NAND2 (N958, N952, N592);
nand NAND3 (N959, N956, N773, N210);
xor XOR2 (N960, N931, N353);
not NOT1 (N961, N953);
buf BUF1 (N962, N950);
nor NOR4 (N963, N962, N111, N66, N846);
nor NOR4 (N964, N940, N922, N932, N303);
or OR4 (N965, N958, N575, N425, N787);
nand NAND4 (N966, N964, N335, N375, N66);
or OR3 (N967, N955, N573, N656);
or OR2 (N968, N959, N770);
and AND4 (N969, N951, N448, N518, N645);
not NOT1 (N970, N963);
or OR3 (N971, N961, N941, N799);
buf BUF1 (N972, N967);
or OR4 (N973, N968, N376, N508, N746);
or OR3 (N974, N960, N566, N825);
or OR2 (N975, N957, N284);
buf BUF1 (N976, N970);
and AND4 (N977, N954, N403, N566, N448);
and AND3 (N978, N969, N123, N309);
buf BUF1 (N979, N978);
buf BUF1 (N980, N971);
and AND4 (N981, N973, N749, N262, N779);
xor XOR2 (N982, N981, N934);
nor NOR4 (N983, N965, N293, N609, N114);
not NOT1 (N984, N976);
not NOT1 (N985, N983);
or OR2 (N986, N982, N654);
buf BUF1 (N987, N966);
and AND3 (N988, N974, N48, N733);
nand NAND3 (N989, N988, N287, N559);
nor NOR2 (N990, N989, N463);
buf BUF1 (N991, N979);
not NOT1 (N992, N985);
xor XOR2 (N993, N984, N395);
xor XOR2 (N994, N977, N951);
xor XOR2 (N995, N994, N888);
xor XOR2 (N996, N975, N449);
not NOT1 (N997, N992);
nand NAND2 (N998, N997, N915);
or OR2 (N999, N993, N782);
or OR3 (N1000, N991, N887, N819);
or OR4 (N1001, N980, N64, N802, N175);
nand NAND3 (N1002, N990, N198, N791);
or OR3 (N1003, N986, N891, N54);
not NOT1 (N1004, N972);
or OR3 (N1005, N1002, N634, N68);
nand NAND3 (N1006, N1003, N230, N910);
buf BUF1 (N1007, N1006);
nand NAND2 (N1008, N998, N320);
xor XOR2 (N1009, N1008, N997);
nor NOR3 (N1010, N1005, N123, N211);
not NOT1 (N1011, N1004);
nor NOR4 (N1012, N1009, N988, N393, N1);
and AND4 (N1013, N996, N372, N75, N357);
nor NOR4 (N1014, N995, N552, N240, N466);
not NOT1 (N1015, N987);
and AND4 (N1016, N1010, N411, N890, N38);
not NOT1 (N1017, N1016);
nor NOR2 (N1018, N1017, N333);
nor NOR2 (N1019, N1013, N502);
buf BUF1 (N1020, N1011);
or OR4 (N1021, N1018, N86, N950, N13);
buf BUF1 (N1022, N1012);
not NOT1 (N1023, N1015);
and AND3 (N1024, N1007, N737, N332);
buf BUF1 (N1025, N1020);
xor XOR2 (N1026, N1000, N460);
nand NAND4 (N1027, N1019, N434, N538, N703);
buf BUF1 (N1028, N1014);
xor XOR2 (N1029, N1021, N270);
buf BUF1 (N1030, N999);
and AND3 (N1031, N1025, N338, N746);
nand NAND2 (N1032, N1027, N75);
or OR2 (N1033, N1024, N178);
nand NAND3 (N1034, N1030, N488, N761);
nand NAND2 (N1035, N1026, N390);
and AND4 (N1036, N1035, N130, N611, N620);
nor NOR3 (N1037, N1028, N199, N855);
buf BUF1 (N1038, N1033);
nor NOR4 (N1039, N1023, N815, N613, N1023);
xor XOR2 (N1040, N1032, N116);
buf BUF1 (N1041, N1039);
buf BUF1 (N1042, N1040);
not NOT1 (N1043, N1022);
buf BUF1 (N1044, N1041);
and AND4 (N1045, N1036, N884, N637, N641);
nor NOR3 (N1046, N1029, N146, N639);
buf BUF1 (N1047, N1001);
xor XOR2 (N1048, N1044, N411);
nand NAND2 (N1049, N1042, N915);
and AND2 (N1050, N1034, N283);
nand NAND4 (N1051, N1050, N550, N100, N197);
nor NOR2 (N1052, N1045, N1036);
xor XOR2 (N1053, N1048, N1044);
nor NOR2 (N1054, N1038, N930);
nand NAND3 (N1055, N1049, N824, N968);
xor XOR2 (N1056, N1047, N58);
buf BUF1 (N1057, N1052);
and AND3 (N1058, N1053, N244, N620);
nor NOR2 (N1059, N1037, N9);
not NOT1 (N1060, N1059);
xor XOR2 (N1061, N1046, N359);
buf BUF1 (N1062, N1061);
and AND2 (N1063, N1055, N510);
nand NAND3 (N1064, N1057, N1029, N666);
xor XOR2 (N1065, N1054, N437);
nand NAND2 (N1066, N1031, N807);
nor NOR2 (N1067, N1062, N841);
nand NAND2 (N1068, N1056, N417);
and AND3 (N1069, N1051, N659, N3);
nand NAND3 (N1070, N1068, N137, N168);
xor XOR2 (N1071, N1043, N73);
xor XOR2 (N1072, N1069, N262);
nor NOR4 (N1073, N1070, N11, N820, N544);
and AND3 (N1074, N1072, N721, N153);
nor NOR4 (N1075, N1067, N300, N1017, N487);
and AND3 (N1076, N1063, N867, N521);
and AND4 (N1077, N1076, N1049, N599, N665);
or OR4 (N1078, N1071, N991, N1028, N590);
and AND2 (N1079, N1074, N412);
nor NOR2 (N1080, N1066, N596);
nand NAND2 (N1081, N1065, N1080);
nor NOR4 (N1082, N229, N396, N688, N1059);
xor XOR2 (N1083, N1079, N964);
buf BUF1 (N1084, N1081);
and AND4 (N1085, N1077, N694, N833, N998);
and AND3 (N1086, N1084, N17, N407);
buf BUF1 (N1087, N1085);
nand NAND2 (N1088, N1060, N668);
not NOT1 (N1089, N1082);
nand NAND2 (N1090, N1089, N986);
nand NAND3 (N1091, N1064, N668, N161);
or OR3 (N1092, N1073, N674, N649);
xor XOR2 (N1093, N1075, N421);
buf BUF1 (N1094, N1092);
nand NAND4 (N1095, N1091, N310, N474, N653);
buf BUF1 (N1096, N1095);
buf BUF1 (N1097, N1078);
xor XOR2 (N1098, N1058, N1019);
nand NAND4 (N1099, N1086, N991, N151, N571);
buf BUF1 (N1100, N1098);
nand NAND2 (N1101, N1083, N572);
buf BUF1 (N1102, N1093);
and AND4 (N1103, N1102, N202, N128, N608);
and AND4 (N1104, N1100, N956, N231, N760);
not NOT1 (N1105, N1104);
and AND2 (N1106, N1101, N728);
or OR2 (N1107, N1090, N671);
nand NAND3 (N1108, N1103, N174, N791);
or OR4 (N1109, N1099, N790, N936, N845);
nand NAND2 (N1110, N1106, N540);
xor XOR2 (N1111, N1105, N534);
not NOT1 (N1112, N1111);
not NOT1 (N1113, N1088);
and AND4 (N1114, N1113, N930, N494, N246);
and AND4 (N1115, N1087, N1031, N801, N128);
xor XOR2 (N1116, N1094, N36);
nor NOR3 (N1117, N1108, N752, N473);
and AND2 (N1118, N1116, N474);
nand NAND3 (N1119, N1096, N675, N145);
nand NAND3 (N1120, N1110, N363, N751);
xor XOR2 (N1121, N1115, N463);
nor NOR4 (N1122, N1119, N158, N606, N244);
xor XOR2 (N1123, N1121, N276);
xor XOR2 (N1124, N1120, N161);
buf BUF1 (N1125, N1118);
xor XOR2 (N1126, N1107, N421);
buf BUF1 (N1127, N1122);
or OR3 (N1128, N1117, N167, N652);
or OR4 (N1129, N1109, N212, N1054, N491);
xor XOR2 (N1130, N1128, N1021);
buf BUF1 (N1131, N1114);
and AND4 (N1132, N1126, N685, N164, N183);
not NOT1 (N1133, N1124);
not NOT1 (N1134, N1133);
xor XOR2 (N1135, N1131, N741);
not NOT1 (N1136, N1112);
or OR3 (N1137, N1136, N485, N712);
buf BUF1 (N1138, N1127);
and AND4 (N1139, N1137, N193, N630, N696);
buf BUF1 (N1140, N1123);
not NOT1 (N1141, N1097);
and AND3 (N1142, N1132, N979, N70);
buf BUF1 (N1143, N1142);
and AND3 (N1144, N1139, N704, N741);
nor NOR3 (N1145, N1138, N897, N365);
not NOT1 (N1146, N1140);
buf BUF1 (N1147, N1135);
xor XOR2 (N1148, N1129, N481);
or OR3 (N1149, N1144, N222, N284);
not NOT1 (N1150, N1134);
nor NOR3 (N1151, N1146, N493, N42);
and AND2 (N1152, N1130, N443);
buf BUF1 (N1153, N1149);
nor NOR3 (N1154, N1125, N255, N273);
or OR4 (N1155, N1143, N461, N698, N273);
xor XOR2 (N1156, N1150, N1011);
xor XOR2 (N1157, N1154, N641);
xor XOR2 (N1158, N1155, N97);
and AND2 (N1159, N1145, N426);
nand NAND2 (N1160, N1147, N594);
buf BUF1 (N1161, N1160);
xor XOR2 (N1162, N1161, N807);
not NOT1 (N1163, N1152);
or OR4 (N1164, N1163, N529, N543, N58);
or OR2 (N1165, N1164, N1125);
or OR4 (N1166, N1159, N283, N238, N406);
or OR2 (N1167, N1141, N54);
and AND4 (N1168, N1157, N443, N1056, N94);
and AND2 (N1169, N1158, N823);
or OR4 (N1170, N1169, N8, N610, N821);
or OR2 (N1171, N1151, N421);
nor NOR4 (N1172, N1156, N149, N383, N1097);
nor NOR2 (N1173, N1166, N823);
nor NOR3 (N1174, N1173, N285, N451);
nand NAND3 (N1175, N1174, N512, N116);
or OR3 (N1176, N1162, N666, N851);
or OR2 (N1177, N1168, N149);
and AND2 (N1178, N1167, N386);
nor NOR3 (N1179, N1165, N917, N268);
buf BUF1 (N1180, N1170);
and AND2 (N1181, N1172, N156);
or OR4 (N1182, N1181, N928, N430, N1168);
and AND4 (N1183, N1180, N281, N680, N364);
and AND2 (N1184, N1171, N232);
nor NOR2 (N1185, N1178, N626);
and AND2 (N1186, N1182, N57);
xor XOR2 (N1187, N1175, N1106);
or OR4 (N1188, N1184, N191, N1184, N819);
not NOT1 (N1189, N1187);
nor NOR4 (N1190, N1179, N1074, N1157, N826);
nor NOR2 (N1191, N1148, N192);
and AND3 (N1192, N1189, N808, N136);
nor NOR4 (N1193, N1176, N933, N798, N126);
not NOT1 (N1194, N1153);
nand NAND2 (N1195, N1193, N174);
or OR3 (N1196, N1177, N284, N579);
nor NOR3 (N1197, N1185, N709, N205);
nand NAND3 (N1198, N1195, N538, N1003);
nor NOR3 (N1199, N1191, N92, N901);
or OR3 (N1200, N1192, N614, N599);
and AND3 (N1201, N1183, N401, N1200);
nor NOR4 (N1202, N706, N729, N270, N763);
nor NOR3 (N1203, N1188, N499, N588);
not NOT1 (N1204, N1202);
nor NOR4 (N1205, N1194, N1012, N390, N195);
nor NOR4 (N1206, N1204, N429, N1034, N38);
buf BUF1 (N1207, N1190);
or OR2 (N1208, N1196, N939);
or OR2 (N1209, N1208, N875);
nand NAND3 (N1210, N1205, N444, N813);
nand NAND3 (N1211, N1206, N347, N1176);
nand NAND3 (N1212, N1207, N827, N208);
not NOT1 (N1213, N1186);
and AND2 (N1214, N1209, N322);
nor NOR3 (N1215, N1210, N1160, N45);
or OR2 (N1216, N1212, N198);
and AND3 (N1217, N1215, N1214, N472);
and AND3 (N1218, N803, N1184, N1217);
buf BUF1 (N1219, N225);
not NOT1 (N1220, N1201);
xor XOR2 (N1221, N1199, N698);
or OR2 (N1222, N1218, N319);
buf BUF1 (N1223, N1197);
xor XOR2 (N1224, N1219, N570);
buf BUF1 (N1225, N1211);
nand NAND3 (N1226, N1221, N107, N202);
not NOT1 (N1227, N1224);
and AND4 (N1228, N1198, N402, N1142, N153);
and AND3 (N1229, N1226, N938, N456);
and AND4 (N1230, N1228, N359, N905, N654);
not NOT1 (N1231, N1229);
buf BUF1 (N1232, N1223);
buf BUF1 (N1233, N1203);
not NOT1 (N1234, N1213);
and AND4 (N1235, N1230, N740, N701, N100);
nor NOR2 (N1236, N1225, N567);
or OR2 (N1237, N1235, N1081);
nand NAND4 (N1238, N1237, N76, N599, N700);
nand NAND4 (N1239, N1220, N149, N1031, N10);
nand NAND3 (N1240, N1227, N188, N752);
or OR3 (N1241, N1216, N519, N983);
nand NAND2 (N1242, N1231, N1116);
nand NAND4 (N1243, N1222, N229, N396, N1067);
buf BUF1 (N1244, N1243);
nor NOR2 (N1245, N1241, N208);
nand NAND4 (N1246, N1236, N336, N947, N632);
xor XOR2 (N1247, N1238, N794);
nand NAND3 (N1248, N1247, N408, N979);
buf BUF1 (N1249, N1246);
or OR3 (N1250, N1232, N327, N532);
or OR3 (N1251, N1239, N430, N743);
and AND4 (N1252, N1250, N1168, N442, N539);
xor XOR2 (N1253, N1240, N1150);
not NOT1 (N1254, N1245);
or OR3 (N1255, N1242, N248, N741);
or OR2 (N1256, N1249, N889);
nor NOR3 (N1257, N1252, N1090, N530);
or OR4 (N1258, N1233, N613, N1090, N376);
nand NAND4 (N1259, N1256, N1144, N542, N402);
buf BUF1 (N1260, N1257);
nand NAND2 (N1261, N1244, N93);
not NOT1 (N1262, N1260);
nand NAND3 (N1263, N1253, N711, N823);
not NOT1 (N1264, N1261);
xor XOR2 (N1265, N1254, N1142);
not NOT1 (N1266, N1259);
xor XOR2 (N1267, N1262, N31);
not NOT1 (N1268, N1251);
and AND3 (N1269, N1234, N699, N799);
nor NOR3 (N1270, N1268, N621, N547);
or OR3 (N1271, N1255, N706, N87);
nand NAND2 (N1272, N1270, N1034);
xor XOR2 (N1273, N1258, N884);
or OR2 (N1274, N1273, N752);
buf BUF1 (N1275, N1272);
xor XOR2 (N1276, N1265, N726);
nor NOR4 (N1277, N1267, N976, N1047, N980);
nor NOR4 (N1278, N1275, N529, N1181, N498);
xor XOR2 (N1279, N1271, N311);
and AND4 (N1280, N1278, N699, N877, N1097);
nor NOR2 (N1281, N1276, N565);
xor XOR2 (N1282, N1266, N318);
nor NOR2 (N1283, N1277, N555);
and AND2 (N1284, N1282, N1241);
or OR4 (N1285, N1274, N704, N44, N149);
buf BUF1 (N1286, N1248);
nor NOR3 (N1287, N1264, N703, N416);
nand NAND4 (N1288, N1280, N438, N944, N572);
buf BUF1 (N1289, N1283);
or OR3 (N1290, N1289, N353, N1060);
and AND3 (N1291, N1269, N582, N450);
buf BUF1 (N1292, N1287);
or OR3 (N1293, N1284, N1208, N1028);
nor NOR2 (N1294, N1279, N1125);
nor NOR4 (N1295, N1286, N340, N263, N406);
not NOT1 (N1296, N1281);
and AND2 (N1297, N1292, N675);
buf BUF1 (N1298, N1295);
nand NAND4 (N1299, N1263, N68, N980, N262);
buf BUF1 (N1300, N1290);
not NOT1 (N1301, N1293);
not NOT1 (N1302, N1298);
buf BUF1 (N1303, N1301);
nand NAND4 (N1304, N1299, N62, N675, N613);
not NOT1 (N1305, N1296);
nand NAND2 (N1306, N1294, N672);
nand NAND2 (N1307, N1305, N829);
and AND4 (N1308, N1288, N719, N1104, N406);
buf BUF1 (N1309, N1285);
nor NOR4 (N1310, N1300, N106, N1237, N1022);
buf BUF1 (N1311, N1308);
not NOT1 (N1312, N1311);
or OR2 (N1313, N1306, N529);
buf BUF1 (N1314, N1312);
nand NAND3 (N1315, N1297, N747, N1048);
xor XOR2 (N1316, N1307, N437);
and AND2 (N1317, N1291, N1130);
nand NAND4 (N1318, N1303, N1256, N970, N1204);
buf BUF1 (N1319, N1316);
not NOT1 (N1320, N1317);
not NOT1 (N1321, N1313);
or OR3 (N1322, N1318, N1303, N198);
xor XOR2 (N1323, N1319, N190);
xor XOR2 (N1324, N1323, N803);
and AND3 (N1325, N1310, N563, N273);
not NOT1 (N1326, N1302);
and AND2 (N1327, N1325, N272);
and AND3 (N1328, N1326, N684, N739);
not NOT1 (N1329, N1322);
buf BUF1 (N1330, N1320);
nor NOR3 (N1331, N1309, N823, N70);
buf BUF1 (N1332, N1324);
or OR3 (N1333, N1331, N1294, N1141);
nand NAND4 (N1334, N1333, N1299, N925, N389);
xor XOR2 (N1335, N1334, N109);
nand NAND2 (N1336, N1315, N401);
nand NAND4 (N1337, N1327, N486, N1072, N738);
or OR3 (N1338, N1314, N857, N1048);
or OR2 (N1339, N1336, N398);
nand NAND2 (N1340, N1321, N559);
xor XOR2 (N1341, N1338, N480);
nand NAND3 (N1342, N1330, N202, N1331);
and AND3 (N1343, N1340, N659, N568);
and AND3 (N1344, N1328, N546, N604);
not NOT1 (N1345, N1335);
nor NOR4 (N1346, N1337, N1108, N1107, N1336);
nand NAND2 (N1347, N1329, N171);
buf BUF1 (N1348, N1342);
nand NAND4 (N1349, N1344, N618, N1147, N1100);
and AND2 (N1350, N1332, N251);
and AND4 (N1351, N1348, N3, N143, N548);
not NOT1 (N1352, N1339);
or OR2 (N1353, N1349, N1230);
buf BUF1 (N1354, N1347);
or OR2 (N1355, N1352, N269);
nor NOR4 (N1356, N1350, N86, N1078, N695);
xor XOR2 (N1357, N1355, N193);
buf BUF1 (N1358, N1356);
nand NAND3 (N1359, N1358, N925, N180);
buf BUF1 (N1360, N1357);
nand NAND3 (N1361, N1359, N1149, N382);
nor NOR3 (N1362, N1346, N1256, N245);
and AND3 (N1363, N1361, N236, N655);
xor XOR2 (N1364, N1363, N365);
nand NAND4 (N1365, N1343, N733, N529, N826);
nand NAND4 (N1366, N1341, N613, N159, N1042);
or OR2 (N1367, N1364, N505);
nand NAND2 (N1368, N1360, N523);
not NOT1 (N1369, N1367);
xor XOR2 (N1370, N1368, N298);
nor NOR4 (N1371, N1369, N611, N339, N102);
or OR3 (N1372, N1345, N120, N313);
and AND3 (N1373, N1365, N817, N1013);
xor XOR2 (N1374, N1370, N287);
not NOT1 (N1375, N1372);
or OR3 (N1376, N1371, N1244, N349);
not NOT1 (N1377, N1375);
buf BUF1 (N1378, N1354);
xor XOR2 (N1379, N1351, N762);
not NOT1 (N1380, N1379);
or OR2 (N1381, N1304, N30);
buf BUF1 (N1382, N1378);
nor NOR3 (N1383, N1381, N1252, N1273);
and AND4 (N1384, N1373, N523, N134, N386);
nand NAND3 (N1385, N1384, N899, N209);
nand NAND2 (N1386, N1353, N1174);
and AND3 (N1387, N1377, N681, N902);
and AND3 (N1388, N1366, N599, N619);
not NOT1 (N1389, N1385);
xor XOR2 (N1390, N1380, N1193);
xor XOR2 (N1391, N1386, N266);
xor XOR2 (N1392, N1390, N453);
not NOT1 (N1393, N1376);
nor NOR3 (N1394, N1393, N264, N1211);
and AND4 (N1395, N1383, N1199, N262, N1173);
nor NOR3 (N1396, N1395, N603, N107);
buf BUF1 (N1397, N1382);
buf BUF1 (N1398, N1392);
xor XOR2 (N1399, N1397, N143);
not NOT1 (N1400, N1388);
not NOT1 (N1401, N1394);
nor NOR3 (N1402, N1391, N693, N880);
and AND2 (N1403, N1400, N1113);
xor XOR2 (N1404, N1374, N1387);
not NOT1 (N1405, N1094);
not NOT1 (N1406, N1389);
xor XOR2 (N1407, N1398, N1326);
not NOT1 (N1408, N1362);
nor NOR3 (N1409, N1408, N585, N1013);
or OR4 (N1410, N1404, N402, N639, N287);
nand NAND3 (N1411, N1406, N158, N746);
or OR4 (N1412, N1405, N328, N1389, N354);
nand NAND3 (N1413, N1411, N497, N729);
nand NAND4 (N1414, N1401, N95, N1174, N1298);
nor NOR3 (N1415, N1414, N239, N1180);
nand NAND4 (N1416, N1413, N910, N541, N955);
not NOT1 (N1417, N1412);
nor NOR3 (N1418, N1407, N278, N98);
xor XOR2 (N1419, N1416, N661);
or OR3 (N1420, N1410, N270, N1266);
not NOT1 (N1421, N1417);
or OR3 (N1422, N1396, N1115, N251);
buf BUF1 (N1423, N1421);
buf BUF1 (N1424, N1422);
and AND3 (N1425, N1403, N290, N602);
or OR2 (N1426, N1399, N1357);
or OR3 (N1427, N1420, N763, N1097);
nor NOR3 (N1428, N1419, N973, N729);
and AND4 (N1429, N1423, N55, N655, N1333);
xor XOR2 (N1430, N1428, N503);
xor XOR2 (N1431, N1409, N1083);
nor NOR4 (N1432, N1418, N1078, N378, N568);
nand NAND3 (N1433, N1429, N294, N525);
or OR4 (N1434, N1431, N1060, N293, N480);
and AND3 (N1435, N1402, N779, N1068);
nor NOR2 (N1436, N1424, N850);
and AND4 (N1437, N1433, N321, N1354, N10);
or OR3 (N1438, N1437, N1387, N1336);
xor XOR2 (N1439, N1425, N1256);
nor NOR2 (N1440, N1435, N1188);
or OR2 (N1441, N1440, N112);
or OR3 (N1442, N1438, N710, N1266);
nor NOR2 (N1443, N1434, N1248);
and AND4 (N1444, N1442, N307, N118, N411);
or OR3 (N1445, N1415, N624, N1103);
nor NOR3 (N1446, N1426, N862, N771);
nand NAND2 (N1447, N1430, N402);
and AND3 (N1448, N1441, N1338, N708);
buf BUF1 (N1449, N1447);
buf BUF1 (N1450, N1449);
nor NOR2 (N1451, N1439, N915);
not NOT1 (N1452, N1443);
and AND3 (N1453, N1427, N111, N752);
buf BUF1 (N1454, N1436);
nor NOR2 (N1455, N1453, N123);
or OR4 (N1456, N1444, N296, N1430, N409);
or OR2 (N1457, N1451, N1229);
xor XOR2 (N1458, N1456, N420);
xor XOR2 (N1459, N1457, N1046);
xor XOR2 (N1460, N1448, N1257);
xor XOR2 (N1461, N1455, N533);
nor NOR4 (N1462, N1454, N875, N1047, N791);
and AND2 (N1463, N1445, N1354);
nand NAND3 (N1464, N1459, N409, N1339);
and AND2 (N1465, N1458, N58);
nand NAND4 (N1466, N1432, N856, N707, N1271);
or OR3 (N1467, N1463, N1351, N1266);
nor NOR4 (N1468, N1462, N64, N844, N289);
nand NAND2 (N1469, N1450, N540);
xor XOR2 (N1470, N1464, N1043);
xor XOR2 (N1471, N1468, N1330);
nor NOR3 (N1472, N1471, N886, N729);
not NOT1 (N1473, N1466);
not NOT1 (N1474, N1465);
nand NAND2 (N1475, N1473, N70);
nor NOR2 (N1476, N1446, N425);
or OR4 (N1477, N1472, N1006, N351, N1150);
not NOT1 (N1478, N1477);
and AND3 (N1479, N1475, N1253, N1462);
nand NAND3 (N1480, N1461, N301, N1192);
nand NAND2 (N1481, N1467, N387);
nor NOR3 (N1482, N1470, N706, N1285);
not NOT1 (N1483, N1452);
or OR4 (N1484, N1479, N1400, N1045, N568);
and AND3 (N1485, N1481, N1469, N54);
nor NOR2 (N1486, N1411, N856);
not NOT1 (N1487, N1485);
not NOT1 (N1488, N1482);
nand NAND3 (N1489, N1484, N60, N1262);
and AND3 (N1490, N1487, N734, N721);
or OR4 (N1491, N1488, N427, N772, N1249);
or OR2 (N1492, N1476, N1203);
nand NAND4 (N1493, N1492, N350, N325, N191);
and AND2 (N1494, N1483, N400);
nor NOR3 (N1495, N1474, N220, N1212);
and AND2 (N1496, N1460, N893);
and AND4 (N1497, N1495, N638, N758, N349);
and AND4 (N1498, N1480, N1147, N93, N147);
nand NAND2 (N1499, N1496, N657);
or OR2 (N1500, N1499, N1237);
nand NAND2 (N1501, N1491, N1156);
nand NAND3 (N1502, N1489, N302, N437);
and AND4 (N1503, N1490, N1162, N572, N474);
nor NOR2 (N1504, N1497, N1035);
xor XOR2 (N1505, N1478, N563);
not NOT1 (N1506, N1503);
and AND3 (N1507, N1494, N412, N502);
nand NAND2 (N1508, N1505, N545);
buf BUF1 (N1509, N1498);
and AND2 (N1510, N1486, N914);
and AND4 (N1511, N1501, N436, N697, N142);
nor NOR4 (N1512, N1508, N723, N157, N657);
not NOT1 (N1513, N1510);
and AND4 (N1514, N1506, N1411, N180, N724);
nor NOR4 (N1515, N1493, N598, N1170, N571);
nand NAND4 (N1516, N1513, N616, N1277, N823);
or OR4 (N1517, N1509, N616, N1312, N286);
buf BUF1 (N1518, N1507);
buf BUF1 (N1519, N1515);
xor XOR2 (N1520, N1504, N996);
nor NOR4 (N1521, N1511, N319, N697, N1020);
nand NAND3 (N1522, N1516, N42, N345);
not NOT1 (N1523, N1521);
and AND2 (N1524, N1522, N201);
nor NOR2 (N1525, N1519, N774);
xor XOR2 (N1526, N1524, N51);
nand NAND3 (N1527, N1502, N474, N706);
or OR4 (N1528, N1520, N1483, N1125, N1283);
not NOT1 (N1529, N1518);
nand NAND4 (N1530, N1517, N1124, N723, N799);
nor NOR4 (N1531, N1512, N1390, N14, N1263);
nor NOR4 (N1532, N1525, N350, N359, N159);
xor XOR2 (N1533, N1523, N1115);
nor NOR3 (N1534, N1528, N1029, N115);
nand NAND3 (N1535, N1531, N1448, N26);
nor NOR2 (N1536, N1500, N497);
xor XOR2 (N1537, N1529, N1061);
nor NOR3 (N1538, N1526, N550, N1136);
xor XOR2 (N1539, N1527, N929);
nor NOR2 (N1540, N1538, N575);
buf BUF1 (N1541, N1537);
and AND3 (N1542, N1534, N484, N26);
buf BUF1 (N1543, N1530);
xor XOR2 (N1544, N1536, N1428);
or OR3 (N1545, N1543, N1405, N34);
xor XOR2 (N1546, N1535, N755);
buf BUF1 (N1547, N1533);
or OR4 (N1548, N1539, N15, N493, N849);
nor NOR4 (N1549, N1547, N1354, N303, N1376);
and AND3 (N1550, N1549, N908, N576);
and AND3 (N1551, N1541, N476, N847);
nor NOR3 (N1552, N1540, N1244, N686);
nand NAND2 (N1553, N1552, N1225);
not NOT1 (N1554, N1542);
and AND3 (N1555, N1551, N555, N701);
nor NOR4 (N1556, N1545, N531, N1336, N1203);
nor NOR2 (N1557, N1544, N1495);
buf BUF1 (N1558, N1548);
buf BUF1 (N1559, N1553);
not NOT1 (N1560, N1559);
and AND2 (N1561, N1555, N892);
nand NAND3 (N1562, N1532, N13, N329);
buf BUF1 (N1563, N1560);
buf BUF1 (N1564, N1562);
not NOT1 (N1565, N1563);
not NOT1 (N1566, N1546);
xor XOR2 (N1567, N1564, N985);
and AND2 (N1568, N1554, N139);
nand NAND3 (N1569, N1514, N1566, N222);
buf BUF1 (N1570, N1284);
xor XOR2 (N1571, N1558, N1021);
nand NAND2 (N1572, N1568, N293);
nand NAND2 (N1573, N1556, N712);
nor NOR4 (N1574, N1557, N143, N231, N393);
and AND3 (N1575, N1550, N389, N717);
and AND4 (N1576, N1567, N929, N596, N1169);
nor NOR3 (N1577, N1569, N1368, N1252);
not NOT1 (N1578, N1575);
not NOT1 (N1579, N1572);
or OR3 (N1580, N1570, N24, N1446);
not NOT1 (N1581, N1580);
nor NOR2 (N1582, N1565, N525);
and AND4 (N1583, N1574, N1185, N1015, N977);
nor NOR3 (N1584, N1561, N321, N1561);
and AND4 (N1585, N1581, N1360, N1534, N1210);
nor NOR3 (N1586, N1584, N660, N314);
xor XOR2 (N1587, N1573, N1530);
or OR2 (N1588, N1586, N1204);
or OR3 (N1589, N1583, N894, N1473);
xor XOR2 (N1590, N1587, N1012);
and AND2 (N1591, N1585, N1557);
nor NOR3 (N1592, N1578, N232, N329);
nand NAND2 (N1593, N1588, N328);
or OR4 (N1594, N1582, N145, N624, N1030);
nor NOR4 (N1595, N1576, N1364, N926, N988);
nand NAND3 (N1596, N1594, N1371, N715);
not NOT1 (N1597, N1591);
xor XOR2 (N1598, N1589, N1583);
or OR4 (N1599, N1593, N123, N466, N1556);
buf BUF1 (N1600, N1595);
not NOT1 (N1601, N1579);
nor NOR4 (N1602, N1601, N234, N263, N820);
nor NOR3 (N1603, N1600, N1103, N1393);
not NOT1 (N1604, N1603);
nor NOR4 (N1605, N1598, N1189, N1378, N990);
not NOT1 (N1606, N1592);
or OR4 (N1607, N1577, N1183, N1405, N1486);
or OR2 (N1608, N1597, N55);
not NOT1 (N1609, N1602);
nor NOR4 (N1610, N1596, N1399, N1259, N905);
nor NOR3 (N1611, N1590, N405, N280);
nand NAND2 (N1612, N1605, N1402);
and AND4 (N1613, N1599, N889, N1032, N1250);
xor XOR2 (N1614, N1613, N673);
xor XOR2 (N1615, N1614, N1099);
and AND4 (N1616, N1608, N1284, N638, N770);
xor XOR2 (N1617, N1606, N1507);
not NOT1 (N1618, N1610);
not NOT1 (N1619, N1615);
buf BUF1 (N1620, N1617);
and AND2 (N1621, N1604, N980);
and AND2 (N1622, N1616, N1470);
not NOT1 (N1623, N1611);
or OR4 (N1624, N1612, N640, N124, N1038);
buf BUF1 (N1625, N1622);
nor NOR2 (N1626, N1607, N1026);
and AND2 (N1627, N1618, N1136);
xor XOR2 (N1628, N1621, N470);
and AND3 (N1629, N1624, N1576, N1236);
nand NAND4 (N1630, N1623, N408, N1034, N238);
xor XOR2 (N1631, N1625, N1541);
buf BUF1 (N1632, N1628);
or OR4 (N1633, N1571, N357, N532, N199);
not NOT1 (N1634, N1631);
nand NAND3 (N1635, N1620, N1568, N773);
and AND3 (N1636, N1626, N878, N1050);
or OR4 (N1637, N1609, N999, N1493, N22);
nand NAND3 (N1638, N1634, N491, N1474);
nor NOR2 (N1639, N1638, N1262);
buf BUF1 (N1640, N1637);
buf BUF1 (N1641, N1629);
xor XOR2 (N1642, N1632, N1106);
not NOT1 (N1643, N1641);
not NOT1 (N1644, N1633);
and AND3 (N1645, N1635, N1388, N233);
xor XOR2 (N1646, N1643, N400);
xor XOR2 (N1647, N1619, N1124);
not NOT1 (N1648, N1640);
not NOT1 (N1649, N1639);
xor XOR2 (N1650, N1647, N20);
nor NOR2 (N1651, N1649, N1125);
not NOT1 (N1652, N1651);
xor XOR2 (N1653, N1636, N976);
nor NOR2 (N1654, N1646, N1629);
and AND4 (N1655, N1650, N180, N123, N715);
nand NAND4 (N1656, N1653, N1409, N752, N852);
and AND3 (N1657, N1645, N1265, N511);
or OR2 (N1658, N1654, N1364);
not NOT1 (N1659, N1658);
nand NAND3 (N1660, N1627, N577, N917);
nand NAND4 (N1661, N1655, N397, N1010, N412);
or OR2 (N1662, N1656, N1645);
xor XOR2 (N1663, N1657, N6);
not NOT1 (N1664, N1660);
buf BUF1 (N1665, N1644);
xor XOR2 (N1666, N1652, N597);
nor NOR3 (N1667, N1661, N321, N1352);
nand NAND2 (N1668, N1630, N619);
not NOT1 (N1669, N1664);
not NOT1 (N1670, N1663);
buf BUF1 (N1671, N1662);
buf BUF1 (N1672, N1642);
or OR3 (N1673, N1670, N402, N1158);
and AND3 (N1674, N1648, N643, N867);
nand NAND4 (N1675, N1666, N1673, N297, N618);
xor XOR2 (N1676, N972, N1448);
or OR4 (N1677, N1659, N1080, N1634, N1610);
nor NOR3 (N1678, N1667, N866, N915);
and AND4 (N1679, N1676, N1276, N932, N63);
nor NOR4 (N1680, N1679, N752, N1261, N102);
or OR2 (N1681, N1680, N1608);
and AND4 (N1682, N1675, N256, N267, N9);
not NOT1 (N1683, N1677);
and AND2 (N1684, N1681, N1348);
not NOT1 (N1685, N1683);
xor XOR2 (N1686, N1672, N918);
nor NOR4 (N1687, N1668, N1187, N1659, N981);
or OR2 (N1688, N1665, N740);
xor XOR2 (N1689, N1685, N1384);
xor XOR2 (N1690, N1688, N1662);
nand NAND4 (N1691, N1690, N1294, N1345, N303);
not NOT1 (N1692, N1671);
nor NOR2 (N1693, N1669, N930);
or OR3 (N1694, N1682, N1434, N761);
nor NOR4 (N1695, N1674, N827, N1619, N50);
nand NAND3 (N1696, N1692, N775, N193);
and AND2 (N1697, N1693, N1377);
and AND2 (N1698, N1691, N1618);
and AND2 (N1699, N1695, N479);
or OR4 (N1700, N1697, N1608, N1614, N1663);
nor NOR3 (N1701, N1686, N345, N1092);
or OR2 (N1702, N1684, N200);
and AND3 (N1703, N1701, N1627, N971);
or OR2 (N1704, N1703, N1438);
buf BUF1 (N1705, N1702);
or OR4 (N1706, N1687, N125, N1274, N1563);
and AND4 (N1707, N1696, N508, N193, N1031);
nand NAND4 (N1708, N1700, N69, N439, N738);
xor XOR2 (N1709, N1704, N894);
and AND2 (N1710, N1706, N91);
and AND4 (N1711, N1710, N478, N549, N888);
nand NAND4 (N1712, N1709, N1671, N749, N1483);
nor NOR4 (N1713, N1705, N1200, N556, N1104);
nor NOR2 (N1714, N1708, N489);
nor NOR4 (N1715, N1711, N133, N531, N354);
xor XOR2 (N1716, N1712, N98);
xor XOR2 (N1717, N1689, N782);
or OR4 (N1718, N1699, N304, N1006, N164);
nand NAND3 (N1719, N1717, N1682, N917);
nand NAND2 (N1720, N1678, N1124);
and AND2 (N1721, N1707, N648);
nand NAND3 (N1722, N1694, N606, N198);
and AND3 (N1723, N1722, N252, N463);
nor NOR3 (N1724, N1723, N976, N532);
buf BUF1 (N1725, N1719);
buf BUF1 (N1726, N1714);
not NOT1 (N1727, N1716);
nand NAND3 (N1728, N1715, N1495, N1002);
buf BUF1 (N1729, N1720);
xor XOR2 (N1730, N1721, N179);
and AND4 (N1731, N1724, N729, N390, N1668);
buf BUF1 (N1732, N1725);
nand NAND2 (N1733, N1718, N1702);
not NOT1 (N1734, N1698);
nor NOR4 (N1735, N1732, N454, N323, N1152);
nor NOR4 (N1736, N1735, N1519, N1714, N1050);
not NOT1 (N1737, N1734);
nand NAND4 (N1738, N1713, N1244, N558, N599);
buf BUF1 (N1739, N1736);
or OR3 (N1740, N1728, N596, N1007);
xor XOR2 (N1741, N1739, N1298);
xor XOR2 (N1742, N1741, N468);
nor NOR4 (N1743, N1727, N407, N242, N1016);
not NOT1 (N1744, N1729);
xor XOR2 (N1745, N1731, N364);
or OR2 (N1746, N1737, N1450);
and AND2 (N1747, N1746, N287);
or OR3 (N1748, N1740, N1309, N733);
xor XOR2 (N1749, N1748, N477);
not NOT1 (N1750, N1749);
nand NAND2 (N1751, N1747, N607);
not NOT1 (N1752, N1751);
or OR2 (N1753, N1752, N1627);
nand NAND2 (N1754, N1745, N903);
or OR2 (N1755, N1743, N1329);
buf BUF1 (N1756, N1730);
or OR3 (N1757, N1756, N666, N229);
xor XOR2 (N1758, N1733, N503);
buf BUF1 (N1759, N1742);
nand NAND3 (N1760, N1753, N566, N754);
xor XOR2 (N1761, N1758, N806);
or OR3 (N1762, N1755, N1420, N1615);
and AND3 (N1763, N1750, N1733, N398);
buf BUF1 (N1764, N1761);
not NOT1 (N1765, N1757);
buf BUF1 (N1766, N1754);
nand NAND4 (N1767, N1744, N465, N1251, N1758);
not NOT1 (N1768, N1767);
xor XOR2 (N1769, N1762, N396);
not NOT1 (N1770, N1759);
nand NAND3 (N1771, N1766, N1266, N83);
xor XOR2 (N1772, N1770, N1103);
and AND4 (N1773, N1769, N7, N143, N1378);
or OR2 (N1774, N1765, N1114);
nor NOR2 (N1775, N1772, N1454);
xor XOR2 (N1776, N1764, N1349);
and AND2 (N1777, N1768, N411);
or OR3 (N1778, N1774, N78, N967);
xor XOR2 (N1779, N1738, N880);
nand NAND4 (N1780, N1776, N1376, N299, N1719);
or OR2 (N1781, N1780, N1280);
buf BUF1 (N1782, N1777);
nand NAND4 (N1783, N1726, N1281, N1620, N115);
not NOT1 (N1784, N1779);
xor XOR2 (N1785, N1778, N1321);
nor NOR4 (N1786, N1775, N624, N454, N1424);
not NOT1 (N1787, N1763);
or OR3 (N1788, N1773, N620, N1392);
buf BUF1 (N1789, N1786);
and AND3 (N1790, N1789, N1001, N314);
buf BUF1 (N1791, N1787);
not NOT1 (N1792, N1781);
nand NAND3 (N1793, N1791, N1512, N805);
xor XOR2 (N1794, N1784, N1155);
buf BUF1 (N1795, N1790);
and AND3 (N1796, N1795, N992, N1007);
nand NAND2 (N1797, N1788, N311);
or OR2 (N1798, N1793, N1785);
buf BUF1 (N1799, N1410);
and AND4 (N1800, N1771, N805, N149, N1597);
xor XOR2 (N1801, N1792, N150);
buf BUF1 (N1802, N1783);
buf BUF1 (N1803, N1800);
nor NOR2 (N1804, N1798, N1444);
nand NAND2 (N1805, N1799, N217);
not NOT1 (N1806, N1796);
nand NAND3 (N1807, N1806, N1101, N231);
or OR4 (N1808, N1804, N1354, N528, N1524);
nand NAND3 (N1809, N1807, N394, N82);
nor NOR3 (N1810, N1797, N719, N1244);
or OR2 (N1811, N1808, N788);
and AND2 (N1812, N1782, N1380);
nor NOR4 (N1813, N1805, N430, N1598, N250);
or OR3 (N1814, N1803, N1166, N1353);
and AND3 (N1815, N1760, N407, N1432);
xor XOR2 (N1816, N1812, N1497);
nand NAND2 (N1817, N1810, N161);
buf BUF1 (N1818, N1816);
buf BUF1 (N1819, N1811);
and AND3 (N1820, N1809, N1312, N1205);
xor XOR2 (N1821, N1815, N1235);
not NOT1 (N1822, N1817);
not NOT1 (N1823, N1822);
nor NOR2 (N1824, N1820, N232);
nand NAND4 (N1825, N1823, N194, N1583, N1462);
or OR4 (N1826, N1802, N196, N656, N831);
nand NAND3 (N1827, N1814, N107, N1146);
buf BUF1 (N1828, N1824);
xor XOR2 (N1829, N1801, N871);
nand NAND3 (N1830, N1828, N697, N1396);
xor XOR2 (N1831, N1794, N1808);
nor NOR4 (N1832, N1829, N1250, N1514, N461);
xor XOR2 (N1833, N1832, N336);
not NOT1 (N1834, N1826);
nand NAND4 (N1835, N1833, N910, N76, N683);
and AND4 (N1836, N1819, N990, N1346, N540);
buf BUF1 (N1837, N1835);
or OR3 (N1838, N1827, N438, N698);
or OR2 (N1839, N1838, N1506);
buf BUF1 (N1840, N1831);
and AND4 (N1841, N1836, N571, N1264, N45);
buf BUF1 (N1842, N1813);
or OR4 (N1843, N1841, N826, N868, N910);
xor XOR2 (N1844, N1818, N1786);
xor XOR2 (N1845, N1837, N1049);
nor NOR4 (N1846, N1842, N1832, N1693, N945);
or OR2 (N1847, N1834, N1731);
nand NAND2 (N1848, N1845, N770);
or OR4 (N1849, N1844, N1809, N1595, N1656);
and AND3 (N1850, N1825, N789, N1831);
nand NAND2 (N1851, N1839, N405);
nand NAND4 (N1852, N1840, N1483, N150, N1589);
buf BUF1 (N1853, N1848);
or OR4 (N1854, N1852, N1146, N431, N1033);
not NOT1 (N1855, N1843);
buf BUF1 (N1856, N1849);
not NOT1 (N1857, N1856);
nor NOR2 (N1858, N1857, N1576);
and AND2 (N1859, N1851, N408);
and AND2 (N1860, N1854, N542);
buf BUF1 (N1861, N1846);
buf BUF1 (N1862, N1855);
nor NOR4 (N1863, N1861, N1775, N1031, N991);
not NOT1 (N1864, N1830);
or OR2 (N1865, N1847, N1579);
nand NAND2 (N1866, N1858, N1552);
and AND4 (N1867, N1864, N74, N1105, N1858);
nand NAND2 (N1868, N1862, N1610);
or OR2 (N1869, N1863, N1328);
buf BUF1 (N1870, N1865);
nand NAND4 (N1871, N1859, N1092, N395, N1778);
nor NOR2 (N1872, N1871, N942);
or OR4 (N1873, N1869, N1856, N1043, N1552);
not NOT1 (N1874, N1870);
not NOT1 (N1875, N1860);
and AND2 (N1876, N1853, N1767);
buf BUF1 (N1877, N1868);
nor NOR4 (N1878, N1867, N542, N231, N1383);
nand NAND2 (N1879, N1876, N130);
xor XOR2 (N1880, N1878, N381);
buf BUF1 (N1881, N1866);
nand NAND4 (N1882, N1873, N208, N545, N588);
nand NAND2 (N1883, N1875, N1799);
nand NAND4 (N1884, N1881, N1807, N1014, N104);
nor NOR2 (N1885, N1879, N341);
nand NAND4 (N1886, N1821, N1462, N1137, N777);
or OR2 (N1887, N1880, N188);
xor XOR2 (N1888, N1850, N380);
or OR2 (N1889, N1882, N1058);
or OR3 (N1890, N1887, N1715, N1029);
nor NOR2 (N1891, N1886, N1413);
nand NAND4 (N1892, N1891, N33, N1726, N177);
xor XOR2 (N1893, N1874, N921);
xor XOR2 (N1894, N1888, N389);
buf BUF1 (N1895, N1890);
not NOT1 (N1896, N1885);
nor NOR3 (N1897, N1884, N96, N1509);
nor NOR3 (N1898, N1895, N1544, N27);
buf BUF1 (N1899, N1897);
nor NOR2 (N1900, N1896, N148);
buf BUF1 (N1901, N1898);
nor NOR4 (N1902, N1889, N1683, N76, N850);
buf BUF1 (N1903, N1894);
nor NOR3 (N1904, N1900, N1785, N789);
xor XOR2 (N1905, N1901, N193);
xor XOR2 (N1906, N1905, N1824);
nor NOR3 (N1907, N1902, N691, N1638);
not NOT1 (N1908, N1907);
nor NOR3 (N1909, N1903, N750, N785);
and AND2 (N1910, N1904, N1406);
xor XOR2 (N1911, N1892, N280);
xor XOR2 (N1912, N1910, N1514);
nor NOR3 (N1913, N1911, N663, N980);
or OR4 (N1914, N1872, N1703, N222, N1652);
not NOT1 (N1915, N1908);
nand NAND4 (N1916, N1877, N479, N1639, N687);
buf BUF1 (N1917, N1914);
xor XOR2 (N1918, N1917, N1703);
not NOT1 (N1919, N1899);
and AND4 (N1920, N1918, N1583, N1532, N862);
nand NAND2 (N1921, N1883, N970);
nand NAND2 (N1922, N1912, N433);
xor XOR2 (N1923, N1920, N1735);
buf BUF1 (N1924, N1919);
buf BUF1 (N1925, N1921);
not NOT1 (N1926, N1923);
nor NOR2 (N1927, N1916, N1014);
nand NAND2 (N1928, N1906, N1429);
nand NAND2 (N1929, N1927, N1088);
and AND3 (N1930, N1926, N1144, N1629);
not NOT1 (N1931, N1928);
not NOT1 (N1932, N1915);
and AND4 (N1933, N1893, N847, N1410, N473);
nor NOR4 (N1934, N1929, N1128, N878, N1839);
nand NAND4 (N1935, N1931, N286, N238, N1795);
buf BUF1 (N1936, N1934);
and AND3 (N1937, N1936, N879, N427);
xor XOR2 (N1938, N1930, N922);
not NOT1 (N1939, N1909);
and AND4 (N1940, N1932, N1104, N164, N1806);
and AND3 (N1941, N1925, N172, N1134);
nand NAND3 (N1942, N1922, N1133, N451);
buf BUF1 (N1943, N1913);
nor NOR4 (N1944, N1938, N922, N207, N1406);
not NOT1 (N1945, N1933);
nand NAND2 (N1946, N1941, N487);
buf BUF1 (N1947, N1940);
buf BUF1 (N1948, N1946);
nor NOR4 (N1949, N1935, N916, N452, N581);
nor NOR3 (N1950, N1944, N696, N1622);
nor NOR2 (N1951, N1950, N445);
and AND2 (N1952, N1945, N1462);
not NOT1 (N1953, N1952);
not NOT1 (N1954, N1937);
buf BUF1 (N1955, N1947);
and AND2 (N1956, N1942, N902);
xor XOR2 (N1957, N1951, N1207);
not NOT1 (N1958, N1957);
nor NOR4 (N1959, N1956, N1134, N1941, N1801);
buf BUF1 (N1960, N1958);
not NOT1 (N1961, N1949);
buf BUF1 (N1962, N1954);
xor XOR2 (N1963, N1962, N980);
nand NAND2 (N1964, N1960, N216);
nor NOR4 (N1965, N1955, N729, N937, N1211);
and AND3 (N1966, N1943, N788, N375);
and AND3 (N1967, N1948, N289, N1604);
or OR4 (N1968, N1939, N1035, N872, N556);
nand NAND3 (N1969, N1967, N945, N1735);
nand NAND3 (N1970, N1966, N1194, N605);
or OR4 (N1971, N1924, N287, N213, N559);
nor NOR2 (N1972, N1965, N1912);
nand NAND4 (N1973, N1968, N251, N1018, N503);
and AND2 (N1974, N1969, N1009);
and AND4 (N1975, N1970, N1418, N1745, N1923);
xor XOR2 (N1976, N1963, N794);
buf BUF1 (N1977, N1971);
nor NOR2 (N1978, N1973, N1124);
xor XOR2 (N1979, N1975, N888);
not NOT1 (N1980, N1959);
or OR3 (N1981, N1979, N1224, N1829);
nand NAND3 (N1982, N1980, N1558, N406);
not NOT1 (N1983, N1982);
nor NOR2 (N1984, N1976, N79);
xor XOR2 (N1985, N1978, N355);
nand NAND3 (N1986, N1964, N1447, N1149);
and AND4 (N1987, N1985, N870, N37, N1699);
buf BUF1 (N1988, N1983);
xor XOR2 (N1989, N1953, N405);
nor NOR3 (N1990, N1981, N1714, N1538);
buf BUF1 (N1991, N1972);
xor XOR2 (N1992, N1991, N328);
nor NOR2 (N1993, N1974, N335);
not NOT1 (N1994, N1977);
not NOT1 (N1995, N1988);
and AND3 (N1996, N1993, N587, N861);
not NOT1 (N1997, N1990);
or OR4 (N1998, N1996, N137, N1010, N598);
not NOT1 (N1999, N1989);
buf BUF1 (N2000, N1998);
nor NOR3 (N2001, N1987, N1897, N1322);
xor XOR2 (N2002, N2000, N404);
or OR4 (N2003, N1961, N693, N662, N627);
buf BUF1 (N2004, N2001);
nor NOR3 (N2005, N2004, N52, N1280);
buf BUF1 (N2006, N1997);
buf BUF1 (N2007, N1986);
nand NAND3 (N2008, N2006, N731, N1708);
not NOT1 (N2009, N2008);
or OR2 (N2010, N1999, N96);
buf BUF1 (N2011, N1992);
nor NOR2 (N2012, N1994, N994);
or OR4 (N2013, N1995, N1291, N170, N1545);
or OR3 (N2014, N2011, N478, N1076);
xor XOR2 (N2015, N2005, N1957);
buf BUF1 (N2016, N2013);
buf BUF1 (N2017, N2009);
and AND4 (N2018, N2012, N706, N83, N413);
nand NAND4 (N2019, N2014, N400, N224, N762);
nor NOR2 (N2020, N2010, N1130);
nor NOR4 (N2021, N1984, N521, N1913, N1119);
or OR2 (N2022, N2018, N1105);
not NOT1 (N2023, N2002);
nand NAND4 (N2024, N2003, N326, N1199, N971);
not NOT1 (N2025, N2020);
xor XOR2 (N2026, N2017, N266);
and AND4 (N2027, N2026, N1953, N1947, N1840);
and AND4 (N2028, N2025, N911, N1397, N126);
xor XOR2 (N2029, N2028, N731);
xor XOR2 (N2030, N2022, N485);
nor NOR2 (N2031, N2007, N733);
not NOT1 (N2032, N2024);
and AND2 (N2033, N2030, N191);
xor XOR2 (N2034, N2015, N547);
nand NAND2 (N2035, N2033, N1740);
xor XOR2 (N2036, N2027, N1506);
and AND2 (N2037, N2016, N1392);
xor XOR2 (N2038, N2019, N1352);
not NOT1 (N2039, N2034);
or OR3 (N2040, N2021, N1528, N546);
or OR3 (N2041, N2040, N126, N860);
xor XOR2 (N2042, N2039, N1532);
or OR2 (N2043, N2035, N1522);
and AND3 (N2044, N2023, N317, N1301);
and AND4 (N2045, N2038, N1921, N403, N1911);
and AND3 (N2046, N2045, N1556, N337);
nor NOR4 (N2047, N2029, N662, N309, N528);
xor XOR2 (N2048, N2047, N1387);
not NOT1 (N2049, N2037);
and AND3 (N2050, N2042, N1616, N1977);
buf BUF1 (N2051, N2048);
not NOT1 (N2052, N2041);
nor NOR3 (N2053, N2052, N1270, N48);
not NOT1 (N2054, N2036);
xor XOR2 (N2055, N2050, N1259);
buf BUF1 (N2056, N2031);
not NOT1 (N2057, N2049);
and AND2 (N2058, N2032, N1454);
nand NAND2 (N2059, N2054, N2048);
not NOT1 (N2060, N2051);
and AND2 (N2061, N2053, N313);
and AND4 (N2062, N2058, N1829, N899, N1845);
xor XOR2 (N2063, N2044, N1304);
nor NOR3 (N2064, N2046, N1552, N811);
or OR3 (N2065, N2064, N45, N1129);
xor XOR2 (N2066, N2063, N2009);
xor XOR2 (N2067, N2062, N1737);
and AND4 (N2068, N2043, N915, N659, N985);
xor XOR2 (N2069, N2067, N1831);
or OR3 (N2070, N2057, N993, N766);
nor NOR3 (N2071, N2066, N1570, N1925);
and AND2 (N2072, N2061, N176);
or OR2 (N2073, N2069, N1521);
and AND2 (N2074, N2073, N1303);
not NOT1 (N2075, N2072);
xor XOR2 (N2076, N2071, N1171);
or OR2 (N2077, N2060, N601);
buf BUF1 (N2078, N2055);
buf BUF1 (N2079, N2065);
nand NAND3 (N2080, N2077, N1027, N1888);
buf BUF1 (N2081, N2075);
and AND2 (N2082, N2078, N1389);
not NOT1 (N2083, N2080);
nor NOR4 (N2084, N2070, N1352, N594, N1232);
nand NAND4 (N2085, N2059, N848, N922, N2030);
nand NAND3 (N2086, N2083, N313, N1744);
not NOT1 (N2087, N2082);
buf BUF1 (N2088, N2079);
nand NAND4 (N2089, N2085, N2072, N1872, N2031);
xor XOR2 (N2090, N2084, N585);
not NOT1 (N2091, N2076);
xor XOR2 (N2092, N2090, N643);
and AND4 (N2093, N2092, N1083, N1920, N175);
nor NOR4 (N2094, N2087, N960, N112, N1233);
buf BUF1 (N2095, N2074);
nor NOR4 (N2096, N2088, N2071, N905, N1664);
not NOT1 (N2097, N2091);
nand NAND2 (N2098, N2094, N1764);
and AND2 (N2099, N2068, N1850);
or OR2 (N2100, N2093, N778);
nand NAND4 (N2101, N2056, N1522, N719, N4);
nor NOR3 (N2102, N2081, N1739, N1328);
or OR4 (N2103, N2098, N1990, N815, N1889);
buf BUF1 (N2104, N2103);
and AND2 (N2105, N2096, N265);
buf BUF1 (N2106, N2100);
and AND3 (N2107, N2086, N1858, N376);
buf BUF1 (N2108, N2106);
buf BUF1 (N2109, N2101);
xor XOR2 (N2110, N2104, N58);
and AND2 (N2111, N2097, N1187);
nor NOR2 (N2112, N2111, N449);
not NOT1 (N2113, N2099);
or OR4 (N2114, N2108, N1144, N745, N945);
or OR4 (N2115, N2095, N1073, N505, N1848);
and AND4 (N2116, N2109, N344, N1431, N1122);
buf BUF1 (N2117, N2113);
xor XOR2 (N2118, N2107, N1644);
not NOT1 (N2119, N2117);
not NOT1 (N2120, N2110);
nand NAND2 (N2121, N2116, N2109);
not NOT1 (N2122, N2114);
nor NOR3 (N2123, N2105, N1186, N508);
xor XOR2 (N2124, N2118, N797);
and AND4 (N2125, N2089, N671, N1178, N642);
or OR2 (N2126, N2125, N1694);
or OR2 (N2127, N2102, N1532);
buf BUF1 (N2128, N2127);
or OR2 (N2129, N2115, N1460);
or OR3 (N2130, N2122, N1919, N1007);
xor XOR2 (N2131, N2130, N1970);
xor XOR2 (N2132, N2112, N537);
nand NAND4 (N2133, N2119, N1330, N1859, N803);
not NOT1 (N2134, N2120);
not NOT1 (N2135, N2123);
and AND4 (N2136, N2128, N1391, N1791, N1796);
xor XOR2 (N2137, N2131, N392);
nor NOR3 (N2138, N2136, N1204, N730);
xor XOR2 (N2139, N2121, N217);
and AND3 (N2140, N2129, N1556, N1331);
or OR4 (N2141, N2135, N431, N460, N12);
or OR3 (N2142, N2126, N1870, N2086);
buf BUF1 (N2143, N2133);
nor NOR2 (N2144, N2141, N1890);
and AND2 (N2145, N2144, N994);
buf BUF1 (N2146, N2124);
nand NAND4 (N2147, N2139, N174, N1705, N44);
nand NAND4 (N2148, N2142, N1906, N289, N1177);
xor XOR2 (N2149, N2145, N637);
nor NOR4 (N2150, N2132, N21, N1755, N463);
not NOT1 (N2151, N2148);
buf BUF1 (N2152, N2138);
nand NAND2 (N2153, N2146, N963);
buf BUF1 (N2154, N2140);
not NOT1 (N2155, N2147);
and AND4 (N2156, N2152, N123, N1600, N124);
and AND2 (N2157, N2137, N228);
buf BUF1 (N2158, N2150);
or OR2 (N2159, N2151, N821);
xor XOR2 (N2160, N2158, N448);
nand NAND4 (N2161, N2134, N898, N762, N816);
not NOT1 (N2162, N2161);
or OR4 (N2163, N2159, N1548, N1579, N245);
or OR3 (N2164, N2162, N1624, N470);
xor XOR2 (N2165, N2154, N1422);
or OR4 (N2166, N2157, N1623, N1545, N1189);
nand NAND2 (N2167, N2153, N1075);
or OR4 (N2168, N2155, N1360, N155, N1063);
not NOT1 (N2169, N2167);
or OR3 (N2170, N2166, N628, N376);
not NOT1 (N2171, N2160);
and AND4 (N2172, N2169, N571, N1810, N1491);
or OR2 (N2173, N2171, N440);
xor XOR2 (N2174, N2163, N1151);
buf BUF1 (N2175, N2143);
nor NOR2 (N2176, N2175, N265);
or OR2 (N2177, N2156, N67);
not NOT1 (N2178, N2164);
not NOT1 (N2179, N2172);
buf BUF1 (N2180, N2173);
not NOT1 (N2181, N2177);
xor XOR2 (N2182, N2180, N550);
or OR3 (N2183, N2170, N418, N716);
or OR3 (N2184, N2168, N304, N648);
nand NAND2 (N2185, N2178, N1714);
or OR4 (N2186, N2176, N252, N1720, N912);
or OR4 (N2187, N2183, N1617, N1508, N1747);
nor NOR4 (N2188, N2174, N1645, N1935, N281);
nor NOR4 (N2189, N2188, N856, N1774, N2029);
not NOT1 (N2190, N2185);
xor XOR2 (N2191, N2186, N471);
or OR4 (N2192, N2189, N1622, N2176, N1654);
and AND2 (N2193, N2187, N1747);
buf BUF1 (N2194, N2193);
nor NOR3 (N2195, N2184, N974, N1595);
buf BUF1 (N2196, N2191);
not NOT1 (N2197, N2196);
and AND4 (N2198, N2195, N1403, N1661, N466);
xor XOR2 (N2199, N2194, N496);
nor NOR3 (N2200, N2197, N312, N1406);
buf BUF1 (N2201, N2198);
or OR2 (N2202, N2179, N848);
not NOT1 (N2203, N2181);
buf BUF1 (N2204, N2200);
and AND4 (N2205, N2201, N219, N425, N1071);
nor NOR4 (N2206, N2149, N1026, N1458, N891);
nand NAND3 (N2207, N2199, N1645, N1823);
not NOT1 (N2208, N2203);
nor NOR4 (N2209, N2204, N1900, N1590, N1912);
xor XOR2 (N2210, N2209, N2050);
and AND2 (N2211, N2207, N345);
and AND4 (N2212, N2205, N1581, N392, N294);
not NOT1 (N2213, N2212);
nand NAND4 (N2214, N2210, N1215, N2043, N814);
and AND4 (N2215, N2206, N918, N1193, N832);
and AND3 (N2216, N2192, N1573, N2064);
or OR3 (N2217, N2213, N2069, N440);
and AND2 (N2218, N2208, N1024);
nor NOR3 (N2219, N2202, N2212, N1679);
not NOT1 (N2220, N2216);
xor XOR2 (N2221, N2215, N1633);
xor XOR2 (N2222, N2190, N813);
not NOT1 (N2223, N2222);
or OR2 (N2224, N2214, N1995);
nor NOR2 (N2225, N2220, N1473);
buf BUF1 (N2226, N2224);
xor XOR2 (N2227, N2211, N806);
xor XOR2 (N2228, N2225, N351);
nand NAND3 (N2229, N2218, N1579, N521);
not NOT1 (N2230, N2223);
nand NAND3 (N2231, N2227, N1501, N2115);
not NOT1 (N2232, N2226);
nor NOR2 (N2233, N2232, N333);
and AND3 (N2234, N2217, N2161, N1132);
buf BUF1 (N2235, N2228);
buf BUF1 (N2236, N2234);
or OR3 (N2237, N2236, N1242, N1694);
or OR4 (N2238, N2165, N2116, N1883, N1244);
not NOT1 (N2239, N2229);
and AND2 (N2240, N2239, N975);
not NOT1 (N2241, N2238);
buf BUF1 (N2242, N2241);
nand NAND4 (N2243, N2230, N1567, N949, N1510);
or OR4 (N2244, N2240, N1221, N412, N1766);
or OR2 (N2245, N2235, N2122);
xor XOR2 (N2246, N2243, N474);
buf BUF1 (N2247, N2242);
and AND3 (N2248, N2247, N1215, N1636);
xor XOR2 (N2249, N2237, N1932);
buf BUF1 (N2250, N2182);
nand NAND2 (N2251, N2245, N2087);
or OR2 (N2252, N2231, N465);
and AND3 (N2253, N2221, N1848, N2072);
or OR2 (N2254, N2249, N36);
and AND4 (N2255, N2251, N1155, N1961, N621);
and AND2 (N2256, N2246, N1915);
nor NOR3 (N2257, N2254, N1913, N233);
buf BUF1 (N2258, N2255);
nor NOR2 (N2259, N2233, N890);
xor XOR2 (N2260, N2258, N768);
and AND3 (N2261, N2256, N1345, N1349);
and AND2 (N2262, N2244, N62);
or OR4 (N2263, N2252, N1229, N244, N1189);
buf BUF1 (N2264, N2262);
and AND2 (N2265, N2263, N1365);
nor NOR2 (N2266, N2265, N702);
or OR4 (N2267, N2264, N395, N354, N97);
nor NOR3 (N2268, N2259, N1559, N253);
and AND2 (N2269, N2257, N10);
buf BUF1 (N2270, N2266);
nor NOR3 (N2271, N2253, N1868, N1342);
nand NAND4 (N2272, N2261, N1886, N1852, N583);
and AND3 (N2273, N2269, N127, N1149);
or OR4 (N2274, N2272, N1609, N1036, N422);
or OR2 (N2275, N2270, N369);
not NOT1 (N2276, N2267);
nand NAND2 (N2277, N2260, N446);
xor XOR2 (N2278, N2250, N1328);
nand NAND4 (N2279, N2275, N1058, N1650, N1263);
nand NAND3 (N2280, N2278, N2059, N441);
nand NAND4 (N2281, N2219, N1592, N565, N1725);
and AND2 (N2282, N2279, N1413);
buf BUF1 (N2283, N2282);
and AND4 (N2284, N2274, N425, N1433, N629);
nand NAND4 (N2285, N2277, N361, N2127, N183);
and AND2 (N2286, N2280, N684);
nand NAND4 (N2287, N2284, N317, N1923, N575);
and AND4 (N2288, N2285, N910, N1887, N1712);
nor NOR2 (N2289, N2286, N1092);
and AND4 (N2290, N2283, N1015, N641, N609);
not NOT1 (N2291, N2273);
and AND4 (N2292, N2289, N374, N544, N1393);
buf BUF1 (N2293, N2290);
nand NAND2 (N2294, N2271, N47);
nand NAND4 (N2295, N2292, N328, N285, N798);
buf BUF1 (N2296, N2268);
nor NOR3 (N2297, N2294, N804, N2230);
nor NOR4 (N2298, N2297, N97, N1211, N665);
or OR3 (N2299, N2293, N378, N321);
buf BUF1 (N2300, N2276);
xor XOR2 (N2301, N2299, N81);
or OR4 (N2302, N2287, N1623, N89, N306);
buf BUF1 (N2303, N2300);
or OR4 (N2304, N2281, N2101, N2184, N332);
not NOT1 (N2305, N2304);
buf BUF1 (N2306, N2305);
not NOT1 (N2307, N2301);
nand NAND3 (N2308, N2291, N2079, N2076);
or OR2 (N2309, N2308, N1003);
buf BUF1 (N2310, N2309);
or OR3 (N2311, N2310, N1081, N300);
buf BUF1 (N2312, N2306);
xor XOR2 (N2313, N2307, N2065);
xor XOR2 (N2314, N2298, N320);
nand NAND3 (N2315, N2302, N1407, N1141);
buf BUF1 (N2316, N2314);
nor NOR4 (N2317, N2316, N2115, N1343, N2112);
buf BUF1 (N2318, N2315);
buf BUF1 (N2319, N2311);
xor XOR2 (N2320, N2303, N1635);
not NOT1 (N2321, N2313);
nand NAND2 (N2322, N2296, N84);
or OR2 (N2323, N2320, N106);
xor XOR2 (N2324, N2318, N1137);
nor NOR2 (N2325, N2319, N7);
or OR4 (N2326, N2321, N1303, N1701, N1462);
and AND4 (N2327, N2322, N1791, N1387, N252);
or OR2 (N2328, N2317, N312);
nor NOR2 (N2329, N2327, N1567);
xor XOR2 (N2330, N2288, N1390);
buf BUF1 (N2331, N2328);
xor XOR2 (N2332, N2330, N1946);
buf BUF1 (N2333, N2248);
or OR3 (N2334, N2295, N2085, N1043);
buf BUF1 (N2335, N2325);
xor XOR2 (N2336, N2332, N262);
not NOT1 (N2337, N2329);
nor NOR2 (N2338, N2336, N1663);
not NOT1 (N2339, N2323);
not NOT1 (N2340, N2326);
not NOT1 (N2341, N2333);
buf BUF1 (N2342, N2338);
or OR2 (N2343, N2331, N271);
buf BUF1 (N2344, N2342);
nand NAND2 (N2345, N2343, N1578);
not NOT1 (N2346, N2337);
and AND3 (N2347, N2312, N1430, N365);
xor XOR2 (N2348, N2347, N2188);
or OR2 (N2349, N2345, N1034);
or OR2 (N2350, N2349, N197);
and AND3 (N2351, N2346, N2030, N1682);
or OR4 (N2352, N2335, N2206, N1168, N1278);
xor XOR2 (N2353, N2344, N1785);
nand NAND3 (N2354, N2352, N1884, N690);
nor NOR3 (N2355, N2324, N822, N2349);
nand NAND3 (N2356, N2355, N2259, N1719);
not NOT1 (N2357, N2339);
not NOT1 (N2358, N2353);
or OR2 (N2359, N2348, N1565);
nand NAND4 (N2360, N2340, N358, N1818, N1281);
nand NAND4 (N2361, N2358, N878, N1828, N2126);
nand NAND3 (N2362, N2360, N199, N75);
buf BUF1 (N2363, N2356);
nor NOR3 (N2364, N2359, N1297, N1414);
nand NAND3 (N2365, N2361, N894, N848);
and AND2 (N2366, N2357, N1885);
nand NAND3 (N2367, N2364, N1097, N104);
nor NOR2 (N2368, N2365, N2050);
nand NAND4 (N2369, N2350, N1284, N189, N1584);
or OR2 (N2370, N2351, N1899);
xor XOR2 (N2371, N2334, N181);
and AND3 (N2372, N2363, N1765, N1071);
xor XOR2 (N2373, N2366, N1139);
xor XOR2 (N2374, N2354, N2162);
nor NOR2 (N2375, N2367, N2133);
buf BUF1 (N2376, N2341);
or OR3 (N2377, N2368, N49, N1633);
and AND2 (N2378, N2370, N2195);
nor NOR4 (N2379, N2371, N1978, N388, N1979);
xor XOR2 (N2380, N2373, N658);
not NOT1 (N2381, N2378);
or OR2 (N2382, N2374, N1344);
or OR2 (N2383, N2379, N1580);
not NOT1 (N2384, N2380);
nor NOR4 (N2385, N2375, N2046, N1333, N2048);
nand NAND4 (N2386, N2383, N1813, N1845, N1885);
buf BUF1 (N2387, N2386);
nor NOR3 (N2388, N2382, N16, N657);
buf BUF1 (N2389, N2384);
not NOT1 (N2390, N2389);
nor NOR3 (N2391, N2362, N1077, N2376);
or OR3 (N2392, N660, N328, N2103);
nor NOR4 (N2393, N2387, N73, N786, N1235);
nand NAND4 (N2394, N2385, N1351, N2053, N122);
nor NOR2 (N2395, N2369, N1824);
xor XOR2 (N2396, N2372, N1669);
nand NAND4 (N2397, N2388, N1693, N1491, N77);
buf BUF1 (N2398, N2393);
or OR4 (N2399, N2390, N1162, N1409, N823);
xor XOR2 (N2400, N2399, N1832);
not NOT1 (N2401, N2397);
buf BUF1 (N2402, N2391);
nand NAND2 (N2403, N2398, N187);
not NOT1 (N2404, N2400);
and AND3 (N2405, N2404, N1753, N776);
or OR4 (N2406, N2403, N2216, N686, N890);
not NOT1 (N2407, N2402);
or OR2 (N2408, N2401, N2384);
nor NOR3 (N2409, N2395, N1057, N2401);
nand NAND4 (N2410, N2409, N1324, N1781, N2407);
buf BUF1 (N2411, N347);
not NOT1 (N2412, N2405);
buf BUF1 (N2413, N2381);
not NOT1 (N2414, N2410);
nor NOR2 (N2415, N2394, N1684);
nand NAND4 (N2416, N2414, N539, N1005, N589);
nor NOR4 (N2417, N2412, N1541, N983, N900);
or OR3 (N2418, N2413, N1644, N16);
and AND2 (N2419, N2408, N1173);
buf BUF1 (N2420, N2415);
buf BUF1 (N2421, N2417);
not NOT1 (N2422, N2392);
buf BUF1 (N2423, N2418);
xor XOR2 (N2424, N2377, N651);
not NOT1 (N2425, N2419);
nor NOR4 (N2426, N2396, N813, N156, N1804);
or OR4 (N2427, N2425, N505, N1282, N1714);
and AND2 (N2428, N2406, N363);
or OR2 (N2429, N2422, N121);
nand NAND2 (N2430, N2424, N1981);
xor XOR2 (N2431, N2427, N2049);
buf BUF1 (N2432, N2411);
nor NOR2 (N2433, N2428, N1033);
buf BUF1 (N2434, N2429);
not NOT1 (N2435, N2430);
not NOT1 (N2436, N2435);
and AND2 (N2437, N2433, N758);
buf BUF1 (N2438, N2436);
or OR2 (N2439, N2438, N2019);
or OR4 (N2440, N2420, N45, N932, N2413);
nor NOR2 (N2441, N2423, N801);
and AND3 (N2442, N2440, N1443, N1727);
not NOT1 (N2443, N2442);
not NOT1 (N2444, N2437);
and AND3 (N2445, N2434, N2168, N1296);
nor NOR3 (N2446, N2439, N2371, N1345);
and AND4 (N2447, N2443, N1101, N1026, N513);
not NOT1 (N2448, N2445);
and AND4 (N2449, N2447, N2017, N2196, N637);
or OR2 (N2450, N2449, N1425);
or OR3 (N2451, N2416, N567, N2218);
or OR2 (N2452, N2432, N21);
buf BUF1 (N2453, N2421);
not NOT1 (N2454, N2452);
not NOT1 (N2455, N2444);
and AND3 (N2456, N2455, N2389, N137);
or OR4 (N2457, N2431, N1083, N1880, N1983);
or OR4 (N2458, N2441, N1620, N197, N77);
nand NAND3 (N2459, N2450, N725, N2085);
buf BUF1 (N2460, N2448);
nor NOR3 (N2461, N2453, N1437, N850);
nand NAND4 (N2462, N2461, N315, N1558, N1604);
not NOT1 (N2463, N2456);
buf BUF1 (N2464, N2457);
xor XOR2 (N2465, N2459, N1254);
nand NAND2 (N2466, N2460, N153);
nand NAND3 (N2467, N2454, N684, N983);
nor NOR4 (N2468, N2462, N79, N1736, N2375);
nand NAND2 (N2469, N2446, N721);
and AND4 (N2470, N2467, N710, N627, N805);
and AND4 (N2471, N2466, N1473, N777, N2259);
not NOT1 (N2472, N2451);
or OR2 (N2473, N2472, N101);
or OR3 (N2474, N2468, N1746, N1955);
nand NAND4 (N2475, N2474, N2051, N1136, N211);
xor XOR2 (N2476, N2464, N453);
buf BUF1 (N2477, N2473);
nand NAND2 (N2478, N2458, N524);
or OR3 (N2479, N2471, N1428, N1152);
buf BUF1 (N2480, N2469);
and AND2 (N2481, N2475, N785);
nor NOR2 (N2482, N2465, N2050);
nor NOR2 (N2483, N2480, N757);
buf BUF1 (N2484, N2482);
or OR3 (N2485, N2470, N919, N185);
or OR4 (N2486, N2483, N1363, N1989, N867);
nor NOR3 (N2487, N2478, N515, N2113);
and AND3 (N2488, N2476, N1988, N1514);
xor XOR2 (N2489, N2488, N2075);
nor NOR3 (N2490, N2487, N2187, N2430);
nand NAND2 (N2491, N2486, N1099);
nand NAND3 (N2492, N2481, N102, N1427);
nand NAND2 (N2493, N2490, N33);
nor NOR4 (N2494, N2493, N2329, N473, N408);
nand NAND3 (N2495, N2492, N192, N2174);
not NOT1 (N2496, N2491);
and AND4 (N2497, N2494, N2166, N1017, N2299);
buf BUF1 (N2498, N2485);
or OR2 (N2499, N2426, N1980);
nand NAND3 (N2500, N2497, N1947, N1705);
buf BUF1 (N2501, N2498);
or OR3 (N2502, N2496, N2114, N1295);
or OR3 (N2503, N2495, N2268, N1361);
and AND2 (N2504, N2477, N116);
xor XOR2 (N2505, N2500, N984);
xor XOR2 (N2506, N2484, N793);
or OR2 (N2507, N2502, N779);
or OR3 (N2508, N2463, N1451, N2247);
buf BUF1 (N2509, N2501);
not NOT1 (N2510, N2507);
nand NAND2 (N2511, N2509, N2031);
and AND4 (N2512, N2504, N365, N1216, N2112);
or OR2 (N2513, N2506, N568);
nand NAND2 (N2514, N2505, N1896);
or OR2 (N2515, N2514, N496);
nor NOR4 (N2516, N2489, N1567, N1119, N2051);
nand NAND4 (N2517, N2499, N332, N217, N196);
or OR2 (N2518, N2515, N49);
nor NOR2 (N2519, N2512, N1589);
or OR2 (N2520, N2510, N111);
xor XOR2 (N2521, N2511, N1139);
nor NOR2 (N2522, N2520, N1964);
not NOT1 (N2523, N2513);
or OR3 (N2524, N2508, N1659, N1141);
nand NAND2 (N2525, N2479, N1758);
xor XOR2 (N2526, N2521, N747);
not NOT1 (N2527, N2523);
nand NAND3 (N2528, N2524, N452, N1706);
nor NOR2 (N2529, N2518, N2370);
or OR3 (N2530, N2525, N1878, N575);
not NOT1 (N2531, N2522);
not NOT1 (N2532, N2529);
not NOT1 (N2533, N2503);
nor NOR4 (N2534, N2531, N135, N128, N425);
buf BUF1 (N2535, N2516);
nand NAND3 (N2536, N2534, N180, N1720);
or OR4 (N2537, N2526, N289, N1158, N2198);
and AND2 (N2538, N2519, N2375);
not NOT1 (N2539, N2517);
or OR4 (N2540, N2533, N1751, N68, N273);
or OR2 (N2541, N2535, N1771);
nor NOR4 (N2542, N2538, N1191, N557, N2532);
buf BUF1 (N2543, N341);
or OR2 (N2544, N2541, N546);
or OR3 (N2545, N2537, N2195, N1569);
buf BUF1 (N2546, N2527);
buf BUF1 (N2547, N2543);
and AND4 (N2548, N2536, N1129, N2215, N801);
nand NAND2 (N2549, N2545, N2366);
nand NAND2 (N2550, N2540, N2510);
xor XOR2 (N2551, N2544, N884);
and AND4 (N2552, N2539, N586, N569, N1850);
buf BUF1 (N2553, N2530);
not NOT1 (N2554, N2550);
xor XOR2 (N2555, N2554, N2026);
and AND2 (N2556, N2549, N1005);
buf BUF1 (N2557, N2553);
buf BUF1 (N2558, N2557);
buf BUF1 (N2559, N2547);
not NOT1 (N2560, N2555);
and AND3 (N2561, N2556, N334, N1074);
not NOT1 (N2562, N2551);
nand NAND4 (N2563, N2560, N2067, N478, N98);
nor NOR4 (N2564, N2548, N1028, N1535, N169);
and AND4 (N2565, N2528, N1128, N2409, N1944);
not NOT1 (N2566, N2564);
nand NAND3 (N2567, N2561, N639, N1358);
xor XOR2 (N2568, N2552, N2449);
and AND3 (N2569, N2563, N2394, N301);
and AND2 (N2570, N2567, N2077);
nor NOR3 (N2571, N2562, N1049, N1096);
nor NOR4 (N2572, N2569, N1115, N1958, N2434);
or OR2 (N2573, N2559, N617);
nand NAND4 (N2574, N2566, N349, N2356, N1320);
not NOT1 (N2575, N2570);
xor XOR2 (N2576, N2575, N127);
and AND4 (N2577, N2571, N1241, N1543, N1312);
or OR2 (N2578, N2573, N480);
xor XOR2 (N2579, N2568, N1272);
and AND2 (N2580, N2576, N2527);
nand NAND4 (N2581, N2542, N808, N2489, N2115);
and AND2 (N2582, N2579, N324);
and AND3 (N2583, N2577, N1635, N333);
nor NOR3 (N2584, N2583, N1198, N2229);
or OR3 (N2585, N2580, N1440, N1483);
nor NOR3 (N2586, N2585, N195, N2519);
xor XOR2 (N2587, N2578, N446);
xor XOR2 (N2588, N2587, N27);
buf BUF1 (N2589, N2572);
xor XOR2 (N2590, N2558, N1083);
nor NOR2 (N2591, N2588, N796);
nand NAND4 (N2592, N2574, N1094, N1991, N1233);
buf BUF1 (N2593, N2546);
xor XOR2 (N2594, N2581, N723);
or OR4 (N2595, N2591, N2529, N255, N1007);
not NOT1 (N2596, N2586);
nand NAND3 (N2597, N2593, N121, N1691);
and AND3 (N2598, N2592, N1283, N2037);
not NOT1 (N2599, N2565);
nor NOR2 (N2600, N2589, N558);
and AND4 (N2601, N2595, N408, N2529, N436);
or OR2 (N2602, N2590, N465);
and AND4 (N2603, N2584, N2092, N93, N1213);
buf BUF1 (N2604, N2598);
nand NAND2 (N2605, N2600, N1252);
nand NAND3 (N2606, N2604, N637, N816);
buf BUF1 (N2607, N2599);
or OR2 (N2608, N2607, N592);
nand NAND2 (N2609, N2602, N2228);
not NOT1 (N2610, N2582);
buf BUF1 (N2611, N2605);
xor XOR2 (N2612, N2594, N39);
nand NAND3 (N2613, N2609, N1567, N1498);
buf BUF1 (N2614, N2611);
xor XOR2 (N2615, N2596, N2360);
buf BUF1 (N2616, N2610);
buf BUF1 (N2617, N2615);
buf BUF1 (N2618, N2612);
nor NOR3 (N2619, N2603, N2368, N2377);
nand NAND4 (N2620, N2597, N2161, N1151, N1646);
nor NOR2 (N2621, N2606, N367);
and AND3 (N2622, N2614, N699, N1910);
nor NOR4 (N2623, N2622, N1425, N1662, N2518);
nor NOR3 (N2624, N2619, N725, N1276);
not NOT1 (N2625, N2617);
not NOT1 (N2626, N2613);
nand NAND4 (N2627, N2620, N2287, N882, N2088);
xor XOR2 (N2628, N2608, N1562);
not NOT1 (N2629, N2621);
nor NOR4 (N2630, N2626, N1691, N998, N240);
and AND3 (N2631, N2630, N1615, N245);
buf BUF1 (N2632, N2624);
not NOT1 (N2633, N2625);
buf BUF1 (N2634, N2618);
or OR4 (N2635, N2631, N2125, N2213, N725);
nor NOR2 (N2636, N2623, N2156);
nor NOR3 (N2637, N2616, N432, N2203);
buf BUF1 (N2638, N2627);
not NOT1 (N2639, N2632);
xor XOR2 (N2640, N2628, N2305);
and AND2 (N2641, N2629, N2);
xor XOR2 (N2642, N2638, N193);
buf BUF1 (N2643, N2640);
not NOT1 (N2644, N2633);
not NOT1 (N2645, N2635);
not NOT1 (N2646, N2639);
not NOT1 (N2647, N2642);
nor NOR2 (N2648, N2641, N1603);
or OR2 (N2649, N2634, N860);
buf BUF1 (N2650, N2643);
xor XOR2 (N2651, N2645, N1300);
nand NAND2 (N2652, N2650, N812);
not NOT1 (N2653, N2644);
not NOT1 (N2654, N2649);
and AND4 (N2655, N2636, N2044, N2288, N479);
or OR3 (N2656, N2601, N2516, N1252);
buf BUF1 (N2657, N2653);
nor NOR3 (N2658, N2648, N2405, N48);
nor NOR2 (N2659, N2652, N2506);
nand NAND4 (N2660, N2656, N2538, N2322, N1700);
not NOT1 (N2661, N2651);
nor NOR4 (N2662, N2655, N2242, N2118, N1717);
xor XOR2 (N2663, N2659, N1723);
not NOT1 (N2664, N2663);
buf BUF1 (N2665, N2658);
nor NOR2 (N2666, N2646, N1740);
not NOT1 (N2667, N2665);
buf BUF1 (N2668, N2654);
and AND4 (N2669, N2668, N1174, N1333, N421);
xor XOR2 (N2670, N2657, N1593);
and AND4 (N2671, N2664, N1700, N1384, N2385);
buf BUF1 (N2672, N2670);
nor NOR4 (N2673, N2660, N1996, N1485, N525);
and AND2 (N2674, N2672, N874);
xor XOR2 (N2675, N2671, N1501);
or OR2 (N2676, N2637, N1313);
buf BUF1 (N2677, N2676);
nand NAND4 (N2678, N2647, N1389, N2554, N2041);
and AND3 (N2679, N2678, N24, N2647);
or OR2 (N2680, N2679, N332);
nand NAND3 (N2681, N2677, N2319, N1270);
not NOT1 (N2682, N2669);
and AND4 (N2683, N2667, N1910, N289, N999);
and AND3 (N2684, N2661, N942, N1581);
xor XOR2 (N2685, N2662, N2331);
nor NOR3 (N2686, N2684, N1548, N2380);
or OR4 (N2687, N2674, N1209, N322, N278);
buf BUF1 (N2688, N2687);
buf BUF1 (N2689, N2683);
xor XOR2 (N2690, N2680, N220);
not NOT1 (N2691, N2682);
nor NOR2 (N2692, N2675, N1456);
nand NAND3 (N2693, N2688, N364, N44);
not NOT1 (N2694, N2673);
or OR2 (N2695, N2689, N929);
nor NOR3 (N2696, N2685, N1827, N807);
buf BUF1 (N2697, N2691);
buf BUF1 (N2698, N2681);
or OR3 (N2699, N2690, N2569, N142);
nand NAND2 (N2700, N2699, N2041);
and AND3 (N2701, N2694, N2545, N1715);
nor NOR2 (N2702, N2693, N256);
buf BUF1 (N2703, N2692);
not NOT1 (N2704, N2696);
and AND3 (N2705, N2704, N156, N1648);
not NOT1 (N2706, N2703);
and AND4 (N2707, N2697, N924, N1964, N266);
or OR2 (N2708, N2695, N1254);
buf BUF1 (N2709, N2701);
nand NAND3 (N2710, N2709, N682, N1286);
nor NOR2 (N2711, N2702, N57);
and AND4 (N2712, N2698, N2270, N1822, N208);
nand NAND3 (N2713, N2705, N1391, N1350);
nand NAND2 (N2714, N2706, N2662);
xor XOR2 (N2715, N2686, N558);
and AND3 (N2716, N2714, N2465, N1416);
not NOT1 (N2717, N2710);
and AND4 (N2718, N2716, N1517, N413, N2449);
nand NAND3 (N2719, N2712, N2315, N166);
nand NAND2 (N2720, N2711, N205);
nor NOR4 (N2721, N2708, N1270, N1865, N1943);
nor NOR4 (N2722, N2721, N643, N1102, N2309);
and AND3 (N2723, N2666, N1896, N684);
nand NAND4 (N2724, N2720, N402, N1714, N1303);
buf BUF1 (N2725, N2724);
and AND2 (N2726, N2722, N2187);
or OR3 (N2727, N2700, N1368, N2166);
or OR3 (N2728, N2707, N518, N2508);
or OR3 (N2729, N2715, N2358, N2135);
not NOT1 (N2730, N2713);
and AND4 (N2731, N2729, N2446, N148, N1980);
and AND4 (N2732, N2719, N2211, N1986, N2020);
nand NAND2 (N2733, N2726, N820);
or OR3 (N2734, N2731, N362, N1979);
not NOT1 (N2735, N2728);
nand NAND3 (N2736, N2733, N2146, N1883);
nand NAND2 (N2737, N2734, N1120);
and AND4 (N2738, N2735, N2509, N777, N1714);
buf BUF1 (N2739, N2738);
nor NOR4 (N2740, N2732, N792, N755, N871);
not NOT1 (N2741, N2725);
nor NOR4 (N2742, N2737, N44, N2347, N509);
buf BUF1 (N2743, N2739);
and AND2 (N2744, N2727, N665);
xor XOR2 (N2745, N2742, N668);
not NOT1 (N2746, N2717);
or OR2 (N2747, N2730, N1102);
nand NAND3 (N2748, N2736, N1060, N853);
nor NOR3 (N2749, N2746, N1583, N2696);
nor NOR3 (N2750, N2749, N2131, N819);
not NOT1 (N2751, N2744);
or OR4 (N2752, N2748, N1834, N722, N177);
nor NOR2 (N2753, N2751, N1042);
not NOT1 (N2754, N2745);
buf BUF1 (N2755, N2743);
or OR3 (N2756, N2750, N2003, N2113);
or OR4 (N2757, N2723, N1141, N1565, N873);
nand NAND4 (N2758, N2757, N90, N1103, N2316);
buf BUF1 (N2759, N2753);
xor XOR2 (N2760, N2755, N76);
or OR4 (N2761, N2754, N2409, N2413, N741);
xor XOR2 (N2762, N2760, N696);
buf BUF1 (N2763, N2761);
nand NAND2 (N2764, N2763, N2524);
and AND2 (N2765, N2740, N1709);
not NOT1 (N2766, N2741);
xor XOR2 (N2767, N2718, N132);
nand NAND4 (N2768, N2756, N1915, N1025, N2377);
not NOT1 (N2769, N2766);
not NOT1 (N2770, N2752);
not NOT1 (N2771, N2770);
nor NOR3 (N2772, N2758, N564, N2210);
or OR2 (N2773, N2759, N968);
xor XOR2 (N2774, N2773, N2432);
or OR3 (N2775, N2768, N2066, N101);
nor NOR4 (N2776, N2772, N597, N221, N2593);
nand NAND2 (N2777, N2771, N169);
nor NOR3 (N2778, N2767, N2341, N1709);
xor XOR2 (N2779, N2775, N1963);
or OR2 (N2780, N2776, N1867);
and AND3 (N2781, N2764, N2666, N155);
nor NOR2 (N2782, N2778, N1909);
nand NAND4 (N2783, N2780, N1312, N1764, N2029);
nor NOR4 (N2784, N2782, N1850, N568, N966);
and AND2 (N2785, N2777, N499);
or OR3 (N2786, N2774, N1859, N2244);
buf BUF1 (N2787, N2762);
nor NOR3 (N2788, N2781, N1446, N474);
buf BUF1 (N2789, N2769);
nand NAND2 (N2790, N2779, N545);
not NOT1 (N2791, N2790);
nor NOR2 (N2792, N2786, N185);
and AND3 (N2793, N2789, N2272, N348);
and AND3 (N2794, N2788, N740, N1747);
or OR4 (N2795, N2783, N769, N622, N1898);
xor XOR2 (N2796, N2794, N460);
or OR4 (N2797, N2793, N617, N2486, N430);
or OR4 (N2798, N2797, N1129, N287, N2368);
and AND2 (N2799, N2792, N2113);
buf BUF1 (N2800, N2798);
xor XOR2 (N2801, N2791, N812);
and AND2 (N2802, N2787, N2105);
and AND4 (N2803, N2796, N1070, N946, N2657);
buf BUF1 (N2804, N2765);
nor NOR2 (N2805, N2800, N1316);
nor NOR2 (N2806, N2805, N2022);
not NOT1 (N2807, N2799);
buf BUF1 (N2808, N2803);
xor XOR2 (N2809, N2785, N201);
not NOT1 (N2810, N2804);
not NOT1 (N2811, N2801);
and AND3 (N2812, N2811, N487, N543);
nor NOR3 (N2813, N2808, N2143, N2401);
not NOT1 (N2814, N2809);
xor XOR2 (N2815, N2814, N97);
not NOT1 (N2816, N2813);
nor NOR4 (N2817, N2807, N771, N1133, N1471);
nor NOR4 (N2818, N2806, N1429, N2106, N2404);
or OR3 (N2819, N2818, N1824, N1403);
not NOT1 (N2820, N2810);
nor NOR4 (N2821, N2816, N2132, N618, N1887);
and AND2 (N2822, N2815, N2165);
nor NOR4 (N2823, N2822, N125, N1799, N451);
or OR2 (N2824, N2812, N924);
not NOT1 (N2825, N2823);
xor XOR2 (N2826, N2821, N1931);
or OR4 (N2827, N2825, N1224, N669, N36);
not NOT1 (N2828, N2826);
or OR3 (N2829, N2802, N432, N1076);
nand NAND3 (N2830, N2827, N566, N2746);
nor NOR2 (N2831, N2819, N1025);
xor XOR2 (N2832, N2747, N278);
nor NOR3 (N2833, N2831, N1403, N1958);
nand NAND2 (N2834, N2824, N1091);
nand NAND4 (N2835, N2784, N1290, N2386, N1918);
or OR3 (N2836, N2832, N2415, N67);
buf BUF1 (N2837, N2833);
nor NOR4 (N2838, N2834, N1964, N390, N475);
not NOT1 (N2839, N2835);
or OR4 (N2840, N2829, N2282, N12, N892);
xor XOR2 (N2841, N2820, N1366);
buf BUF1 (N2842, N2830);
or OR2 (N2843, N2795, N639);
nor NOR2 (N2844, N2817, N723);
buf BUF1 (N2845, N2843);
not NOT1 (N2846, N2840);
or OR4 (N2847, N2842, N1078, N1855, N2048);
xor XOR2 (N2848, N2844, N1947);
nor NOR4 (N2849, N2838, N2050, N1832, N1128);
nor NOR3 (N2850, N2845, N1531, N1600);
or OR2 (N2851, N2828, N2013);
buf BUF1 (N2852, N2851);
not NOT1 (N2853, N2837);
not NOT1 (N2854, N2841);
not NOT1 (N2855, N2847);
or OR4 (N2856, N2836, N388, N2282, N1496);
nor NOR2 (N2857, N2850, N53);
or OR4 (N2858, N2839, N1471, N1261, N1596);
buf BUF1 (N2859, N2854);
xor XOR2 (N2860, N2858, N1755);
xor XOR2 (N2861, N2856, N1601);
xor XOR2 (N2862, N2857, N1193);
and AND4 (N2863, N2853, N1816, N1834, N2647);
nand NAND2 (N2864, N2846, N2274);
not NOT1 (N2865, N2855);
or OR3 (N2866, N2862, N2225, N1556);
nand NAND2 (N2867, N2848, N1829);
nor NOR4 (N2868, N2852, N1982, N916, N811);
not NOT1 (N2869, N2863);
or OR2 (N2870, N2859, N1118);
nor NOR4 (N2871, N2864, N1409, N130, N899);
nand NAND3 (N2872, N2849, N2298, N479);
buf BUF1 (N2873, N2869);
xor XOR2 (N2874, N2860, N2170);
or OR3 (N2875, N2871, N979, N2172);
nand NAND3 (N2876, N2861, N896, N99);
buf BUF1 (N2877, N2865);
xor XOR2 (N2878, N2874, N1903);
nand NAND2 (N2879, N2866, N233);
not NOT1 (N2880, N2868);
and AND2 (N2881, N2878, N897);
xor XOR2 (N2882, N2877, N2052);
nand NAND3 (N2883, N2881, N643, N1812);
or OR2 (N2884, N2880, N2252);
or OR3 (N2885, N2884, N506, N103);
xor XOR2 (N2886, N2885, N1163);
nor NOR4 (N2887, N2870, N1654, N210, N622);
nor NOR3 (N2888, N2883, N1156, N503);
nor NOR2 (N2889, N2879, N2667);
nor NOR2 (N2890, N2873, N1862);
xor XOR2 (N2891, N2888, N2247);
nor NOR2 (N2892, N2890, N1770);
xor XOR2 (N2893, N2887, N51);
not NOT1 (N2894, N2876);
nor NOR4 (N2895, N2882, N2766, N1252, N433);
or OR2 (N2896, N2886, N2147);
and AND3 (N2897, N2894, N674, N2358);
and AND4 (N2898, N2895, N1056, N114, N2253);
buf BUF1 (N2899, N2892);
not NOT1 (N2900, N2867);
nand NAND4 (N2901, N2889, N2813, N635, N2748);
xor XOR2 (N2902, N2893, N2783);
buf BUF1 (N2903, N2872);
nor NOR2 (N2904, N2897, N2591);
and AND2 (N2905, N2896, N2626);
nand NAND3 (N2906, N2891, N2488, N1586);
or OR3 (N2907, N2899, N2714, N1326);
or OR4 (N2908, N2902, N2366, N2384, N1402);
xor XOR2 (N2909, N2875, N2746);
or OR3 (N2910, N2898, N845, N1164);
xor XOR2 (N2911, N2908, N1518);
or OR3 (N2912, N2904, N1318, N2191);
buf BUF1 (N2913, N2907);
buf BUF1 (N2914, N2913);
nor NOR4 (N2915, N2901, N817, N1664, N1089);
nor NOR3 (N2916, N2903, N444, N1220);
and AND2 (N2917, N2915, N1864);
not NOT1 (N2918, N2911);
or OR3 (N2919, N2916, N2294, N418);
or OR4 (N2920, N2905, N457, N1018, N2751);
xor XOR2 (N2921, N2919, N397);
not NOT1 (N2922, N2900);
buf BUF1 (N2923, N2910);
nand NAND3 (N2924, N2917, N2874, N1190);
nor NOR4 (N2925, N2921, N558, N1819, N1547);
xor XOR2 (N2926, N2920, N2569);
nor NOR4 (N2927, N2922, N2140, N636, N1638);
not NOT1 (N2928, N2909);
xor XOR2 (N2929, N2914, N2727);
buf BUF1 (N2930, N2927);
nand NAND4 (N2931, N2912, N1798, N2915, N2679);
nand NAND3 (N2932, N2931, N56, N1637);
not NOT1 (N2933, N2932);
nor NOR4 (N2934, N2923, N1149, N1102, N269);
or OR4 (N2935, N2925, N369, N211, N991);
not NOT1 (N2936, N2930);
nand NAND4 (N2937, N2918, N2725, N1176, N1853);
not NOT1 (N2938, N2928);
nor NOR2 (N2939, N2936, N1630);
nor NOR4 (N2940, N2924, N1573, N458, N2331);
xor XOR2 (N2941, N2933, N556);
and AND2 (N2942, N2926, N1196);
buf BUF1 (N2943, N2938);
and AND3 (N2944, N2906, N47, N2628);
xor XOR2 (N2945, N2929, N736);
nand NAND4 (N2946, N2937, N915, N1060, N921);
xor XOR2 (N2947, N2935, N64);
nor NOR4 (N2948, N2943, N2505, N1571, N839);
not NOT1 (N2949, N2947);
or OR3 (N2950, N2939, N722, N2129);
or OR3 (N2951, N2941, N1272, N2175);
nor NOR2 (N2952, N2948, N486);
and AND4 (N2953, N2946, N1063, N11, N1019);
buf BUF1 (N2954, N2944);
and AND3 (N2955, N2954, N516, N2860);
nor NOR2 (N2956, N2945, N665);
nand NAND2 (N2957, N2949, N452);
or OR3 (N2958, N2953, N1158, N1118);
nor NOR2 (N2959, N2934, N2467);
nor NOR2 (N2960, N2957, N2197);
not NOT1 (N2961, N2955);
not NOT1 (N2962, N2942);
nand NAND2 (N2963, N2940, N1470);
nand NAND3 (N2964, N2959, N2442, N1513);
xor XOR2 (N2965, N2961, N989);
buf BUF1 (N2966, N2962);
buf BUF1 (N2967, N2964);
nand NAND3 (N2968, N2952, N2101, N1514);
xor XOR2 (N2969, N2958, N1545);
or OR2 (N2970, N2969, N753);
not NOT1 (N2971, N2966);
and AND2 (N2972, N2956, N586);
xor XOR2 (N2973, N2950, N1221);
buf BUF1 (N2974, N2970);
or OR2 (N2975, N2963, N2298);
xor XOR2 (N2976, N2971, N1260);
or OR4 (N2977, N2976, N1355, N219, N2434);
nand NAND3 (N2978, N2977, N2671, N519);
xor XOR2 (N2979, N2978, N2337);
and AND3 (N2980, N2972, N2659, N2555);
nand NAND3 (N2981, N2965, N1126, N1463);
buf BUF1 (N2982, N2960);
nor NOR2 (N2983, N2980, N2887);
nor NOR3 (N2984, N2974, N2556, N2351);
or OR3 (N2985, N2975, N2024, N104);
nand NAND2 (N2986, N2968, N492);
xor XOR2 (N2987, N2967, N2701);
buf BUF1 (N2988, N2973);
and AND4 (N2989, N2985, N1928, N2300, N64);
nor NOR2 (N2990, N2982, N2498);
nand NAND4 (N2991, N2981, N1821, N1060, N1177);
not NOT1 (N2992, N2984);
nor NOR2 (N2993, N2951, N2503);
and AND4 (N2994, N2979, N1946, N2604, N923);
nand NAND4 (N2995, N2994, N2120, N2402, N1878);
buf BUF1 (N2996, N2993);
nor NOR4 (N2997, N2991, N645, N135, N2950);
or OR4 (N2998, N2987, N1509, N143, N843);
buf BUF1 (N2999, N2983);
not NOT1 (N3000, N2997);
and AND2 (N3001, N2990, N2069);
xor XOR2 (N3002, N2988, N394);
buf BUF1 (N3003, N2996);
not NOT1 (N3004, N3001);
xor XOR2 (N3005, N3003, N2822);
or OR3 (N3006, N3005, N1515, N2671);
not NOT1 (N3007, N2999);
nor NOR3 (N3008, N2995, N178, N2406);
and AND2 (N3009, N3008, N1844);
not NOT1 (N3010, N3004);
and AND2 (N3011, N2998, N1085);
not NOT1 (N3012, N2989);
and AND4 (N3013, N3007, N723, N931, N1888);
and AND2 (N3014, N3013, N2731);
and AND4 (N3015, N2992, N1194, N2612, N1065);
nand NAND3 (N3016, N3015, N1663, N512);
or OR3 (N3017, N3011, N1825, N1431);
and AND3 (N3018, N3010, N2564, N1497);
nor NOR4 (N3019, N2986, N2641, N337, N1020);
nand NAND3 (N3020, N3006, N889, N2434);
xor XOR2 (N3021, N3016, N1596);
xor XOR2 (N3022, N3020, N1722);
nor NOR2 (N3023, N3000, N2372);
buf BUF1 (N3024, N3017);
xor XOR2 (N3025, N3024, N997);
nor NOR3 (N3026, N3002, N1457, N672);
buf BUF1 (N3027, N3025);
nor NOR4 (N3028, N3012, N1938, N2337, N290);
nor NOR4 (N3029, N3014, N2796, N338, N765);
and AND4 (N3030, N3009, N2984, N2097, N2630);
nor NOR3 (N3031, N3029, N20, N2298);
not NOT1 (N3032, N3031);
buf BUF1 (N3033, N3032);
xor XOR2 (N3034, N3033, N1626);
nand NAND2 (N3035, N3027, N509);
and AND3 (N3036, N3034, N2865, N1931);
or OR3 (N3037, N3019, N2976, N174);
not NOT1 (N3038, N3028);
nand NAND2 (N3039, N3038, N3038);
not NOT1 (N3040, N3023);
nand NAND2 (N3041, N3035, N1283);
or OR3 (N3042, N3036, N2802, N2160);
nor NOR2 (N3043, N3041, N650);
not NOT1 (N3044, N3022);
nand NAND4 (N3045, N3044, N1920, N2208, N1077);
nor NOR3 (N3046, N3045, N1901, N2734);
not NOT1 (N3047, N3046);
xor XOR2 (N3048, N3026, N820);
not NOT1 (N3049, N3040);
buf BUF1 (N3050, N3049);
not NOT1 (N3051, N3030);
xor XOR2 (N3052, N3039, N727);
xor XOR2 (N3053, N3043, N1574);
xor XOR2 (N3054, N3042, N1982);
not NOT1 (N3055, N3047);
or OR3 (N3056, N3018, N907, N1235);
not NOT1 (N3057, N3054);
or OR3 (N3058, N3048, N1816, N2912);
nand NAND3 (N3059, N3037, N2438, N2294);
nor NOR3 (N3060, N3050, N1558, N67);
xor XOR2 (N3061, N3055, N872);
or OR4 (N3062, N3056, N1072, N1789, N1596);
xor XOR2 (N3063, N3058, N109);
xor XOR2 (N3064, N3057, N2983);
not NOT1 (N3065, N3064);
xor XOR2 (N3066, N3063, N2210);
xor XOR2 (N3067, N3021, N1499);
and AND3 (N3068, N3066, N1631, N1734);
and AND4 (N3069, N3065, N980, N1366, N939);
and AND4 (N3070, N3052, N2804, N391, N591);
nor NOR2 (N3071, N3053, N1871);
xor XOR2 (N3072, N3060, N2218);
or OR3 (N3073, N3069, N2744, N2217);
or OR3 (N3074, N3061, N1715, N1756);
xor XOR2 (N3075, N3074, N1249);
xor XOR2 (N3076, N3068, N2356);
or OR4 (N3077, N3070, N2377, N1163, N236);
nor NOR2 (N3078, N3071, N649);
and AND4 (N3079, N3076, N1547, N1384, N1739);
xor XOR2 (N3080, N3075, N1037);
and AND3 (N3081, N3077, N2579, N941);
xor XOR2 (N3082, N3078, N2021);
xor XOR2 (N3083, N3051, N1183);
or OR4 (N3084, N3080, N274, N2431, N2482);
and AND4 (N3085, N3081, N1744, N2546, N3082);
buf BUF1 (N3086, N223);
not NOT1 (N3087, N3073);
nand NAND4 (N3088, N3087, N1319, N107, N198);
and AND3 (N3089, N3079, N2335, N2864);
or OR2 (N3090, N3062, N590);
not NOT1 (N3091, N3067);
and AND3 (N3092, N3091, N533, N969);
nor NOR2 (N3093, N3092, N1450);
not NOT1 (N3094, N3083);
xor XOR2 (N3095, N3088, N3064);
or OR3 (N3096, N3084, N2952, N113);
xor XOR2 (N3097, N3093, N1593);
buf BUF1 (N3098, N3095);
not NOT1 (N3099, N3098);
buf BUF1 (N3100, N3090);
xor XOR2 (N3101, N3059, N511);
and AND2 (N3102, N3072, N1406);
nand NAND2 (N3103, N3094, N1784);
nor NOR4 (N3104, N3099, N1842, N2575, N3007);
not NOT1 (N3105, N3102);
or OR2 (N3106, N3101, N1328);
or OR4 (N3107, N3086, N801, N757, N2774);
nand NAND3 (N3108, N3089, N2485, N3062);
not NOT1 (N3109, N3108);
xor XOR2 (N3110, N3106, N992);
nor NOR3 (N3111, N3104, N2337, N1341);
and AND2 (N3112, N3100, N3075);
not NOT1 (N3113, N3111);
and AND4 (N3114, N3110, N412, N2469, N1502);
buf BUF1 (N3115, N3112);
not NOT1 (N3116, N3085);
not NOT1 (N3117, N3115);
nand NAND4 (N3118, N3114, N808, N2187, N3029);
xor XOR2 (N3119, N3103, N2967);
or OR4 (N3120, N3109, N1099, N2552, N2746);
and AND4 (N3121, N3119, N2991, N1519, N83);
buf BUF1 (N3122, N3107);
not NOT1 (N3123, N3116);
nand NAND4 (N3124, N3120, N2632, N1997, N145);
or OR3 (N3125, N3096, N44, N760);
nand NAND4 (N3126, N3124, N898, N2628, N453);
or OR4 (N3127, N3117, N1404, N250, N1372);
nand NAND3 (N3128, N3105, N2839, N1005);
not NOT1 (N3129, N3122);
and AND4 (N3130, N3121, N2480, N3028, N805);
and AND2 (N3131, N3118, N21);
not NOT1 (N3132, N3128);
xor XOR2 (N3133, N3126, N822);
and AND4 (N3134, N3125, N2952, N3014, N325);
nor NOR2 (N3135, N3132, N1992);
nor NOR3 (N3136, N3135, N2242, N1714);
nand NAND2 (N3137, N3129, N906);
buf BUF1 (N3138, N3130);
buf BUF1 (N3139, N3113);
nand NAND4 (N3140, N3134, N1152, N1543, N2670);
buf BUF1 (N3141, N3136);
or OR2 (N3142, N3127, N796);
xor XOR2 (N3143, N3140, N1250);
or OR4 (N3144, N3143, N2231, N775, N82);
xor XOR2 (N3145, N3139, N1844);
nor NOR3 (N3146, N3145, N195, N665);
buf BUF1 (N3147, N3131);
buf BUF1 (N3148, N3142);
nor NOR2 (N3149, N3123, N673);
buf BUF1 (N3150, N3147);
and AND4 (N3151, N3137, N748, N191, N2816);
xor XOR2 (N3152, N3141, N304);
buf BUF1 (N3153, N3151);
nor NOR3 (N3154, N3144, N2021, N1984);
buf BUF1 (N3155, N3133);
not NOT1 (N3156, N3149);
not NOT1 (N3157, N3153);
or OR3 (N3158, N3146, N1684, N2313);
buf BUF1 (N3159, N3158);
nand NAND2 (N3160, N3138, N2088);
buf BUF1 (N3161, N3152);
xor XOR2 (N3162, N3150, N2634);
and AND4 (N3163, N3161, N1924, N809, N1367);
buf BUF1 (N3164, N3160);
nand NAND3 (N3165, N3097, N1614, N1910);
xor XOR2 (N3166, N3163, N2542);
buf BUF1 (N3167, N3157);
or OR4 (N3168, N3164, N951, N2069, N2031);
nand NAND4 (N3169, N3154, N175, N1936, N2454);
not NOT1 (N3170, N3159);
not NOT1 (N3171, N3166);
nor NOR3 (N3172, N3148, N2616, N2774);
xor XOR2 (N3173, N3169, N2895);
nor NOR2 (N3174, N3155, N2182);
nor NOR4 (N3175, N3165, N1603, N1522, N679);
or OR4 (N3176, N3175, N1056, N1718, N1703);
nor NOR2 (N3177, N3162, N1262);
not NOT1 (N3178, N3177);
or OR3 (N3179, N3178, N1556, N587);
nor NOR4 (N3180, N3167, N596, N406, N932);
nand NAND4 (N3181, N3180, N2178, N1081, N2325);
and AND3 (N3182, N3156, N2968, N743);
nand NAND2 (N3183, N3173, N440);
xor XOR2 (N3184, N3183, N2575);
buf BUF1 (N3185, N3174);
or OR4 (N3186, N3185, N159, N2496, N1998);
and AND4 (N3187, N3170, N2831, N1100, N72);
and AND3 (N3188, N3181, N1436, N1526);
not NOT1 (N3189, N3186);
nand NAND3 (N3190, N3171, N1244, N2213);
and AND3 (N3191, N3179, N1530, N3162);
nand NAND2 (N3192, N3190, N2995);
not NOT1 (N3193, N3184);
xor XOR2 (N3194, N3191, N1039);
buf BUF1 (N3195, N3193);
and AND2 (N3196, N3188, N1770);
not NOT1 (N3197, N3194);
or OR4 (N3198, N3192, N3005, N2205, N1221);
or OR2 (N3199, N3187, N951);
nand NAND3 (N3200, N3172, N2572, N564);
and AND3 (N3201, N3200, N3115, N1849);
not NOT1 (N3202, N3189);
nor NOR4 (N3203, N3182, N1707, N2833, N368);
or OR4 (N3204, N3168, N2711, N3179, N1910);
and AND4 (N3205, N3201, N367, N867, N120);
buf BUF1 (N3206, N3198);
xor XOR2 (N3207, N3196, N1593);
nand NAND4 (N3208, N3203, N2730, N2921, N120);
and AND4 (N3209, N3202, N2893, N1543, N666);
nor NOR4 (N3210, N3206, N1095, N2982, N1075);
or OR4 (N3211, N3209, N2651, N2809, N1669);
nand NAND2 (N3212, N3205, N1176);
or OR2 (N3213, N3197, N2132);
and AND2 (N3214, N3210, N1567);
buf BUF1 (N3215, N3213);
not NOT1 (N3216, N3208);
or OR4 (N3217, N3215, N564, N390, N1511);
buf BUF1 (N3218, N3216);
xor XOR2 (N3219, N3204, N1497);
nor NOR2 (N3220, N3199, N1982);
not NOT1 (N3221, N3220);
nor NOR2 (N3222, N3176, N2830);
nand NAND2 (N3223, N3219, N2880);
and AND3 (N3224, N3214, N3093, N346);
buf BUF1 (N3225, N3223);
or OR4 (N3226, N3222, N899, N1763, N2539);
nor NOR3 (N3227, N3207, N994, N1162);
xor XOR2 (N3228, N3227, N1017);
xor XOR2 (N3229, N3211, N1543);
buf BUF1 (N3230, N3218);
not NOT1 (N3231, N3225);
and AND3 (N3232, N3212, N2230, N230);
not NOT1 (N3233, N3224);
xor XOR2 (N3234, N3232, N680);
nand NAND4 (N3235, N3234, N2247, N2419, N2825);
xor XOR2 (N3236, N3233, N685);
or OR3 (N3237, N3235, N526, N1242);
xor XOR2 (N3238, N3228, N1149);
and AND3 (N3239, N3238, N246, N2239);
buf BUF1 (N3240, N3239);
or OR3 (N3241, N3230, N3050, N2369);
not NOT1 (N3242, N3237);
buf BUF1 (N3243, N3226);
nand NAND2 (N3244, N3231, N2051);
and AND2 (N3245, N3242, N507);
xor XOR2 (N3246, N3229, N2059);
nor NOR3 (N3247, N3221, N1104, N2179);
or OR3 (N3248, N3195, N1438, N1460);
or OR2 (N3249, N3244, N3182);
nand NAND2 (N3250, N3243, N2720);
not NOT1 (N3251, N3245);
buf BUF1 (N3252, N3217);
xor XOR2 (N3253, N3241, N833);
buf BUF1 (N3254, N3246);
nand NAND3 (N3255, N3254, N3161, N1742);
buf BUF1 (N3256, N3247);
or OR3 (N3257, N3240, N2943, N1071);
nor NOR4 (N3258, N3251, N2296, N1617, N3100);
nor NOR2 (N3259, N3236, N1016);
xor XOR2 (N3260, N3257, N3097);
not NOT1 (N3261, N3255);
not NOT1 (N3262, N3250);
buf BUF1 (N3263, N3258);
or OR2 (N3264, N3261, N2987);
not NOT1 (N3265, N3263);
buf BUF1 (N3266, N3252);
nor NOR4 (N3267, N3248, N985, N1354, N858);
buf BUF1 (N3268, N3265);
buf BUF1 (N3269, N3267);
nand NAND3 (N3270, N3264, N2857, N391);
nand NAND2 (N3271, N3253, N643);
or OR4 (N3272, N3268, N1319, N675, N2555);
xor XOR2 (N3273, N3271, N2147);
and AND2 (N3274, N3273, N764);
nor NOR3 (N3275, N3270, N2342, N575);
nand NAND2 (N3276, N3260, N529);
and AND3 (N3277, N3272, N2071, N396);
nor NOR4 (N3278, N3269, N1038, N619, N2508);
buf BUF1 (N3279, N3266);
xor XOR2 (N3280, N3262, N657);
nand NAND2 (N3281, N3278, N2114);
nor NOR3 (N3282, N3281, N3163, N701);
not NOT1 (N3283, N3277);
buf BUF1 (N3284, N3274);
or OR2 (N3285, N3249, N1264);
and AND4 (N3286, N3280, N2178, N2690, N2609);
or OR2 (N3287, N3282, N1908);
and AND4 (N3288, N3259, N1694, N1548, N792);
or OR2 (N3289, N3287, N1820);
or OR3 (N3290, N3279, N1887, N2468);
or OR2 (N3291, N3286, N1762);
nand NAND4 (N3292, N3256, N656, N3075, N338);
not NOT1 (N3293, N3292);
xor XOR2 (N3294, N3283, N2961);
and AND2 (N3295, N3290, N2717);
xor XOR2 (N3296, N3276, N2331);
nor NOR2 (N3297, N3296, N1255);
buf BUF1 (N3298, N3275);
or OR2 (N3299, N3294, N3018);
or OR4 (N3300, N3285, N2649, N176, N1479);
xor XOR2 (N3301, N3299, N1055);
nor NOR2 (N3302, N3297, N736);
nor NOR2 (N3303, N3301, N2591);
nand NAND4 (N3304, N3298, N2697, N2910, N1659);
nor NOR2 (N3305, N3288, N278);
or OR3 (N3306, N3291, N1946, N3159);
and AND3 (N3307, N3300, N2301, N2043);
not NOT1 (N3308, N3289);
nand NAND3 (N3309, N3304, N2804, N2632);
nor NOR2 (N3310, N3302, N2247);
and AND4 (N3311, N3295, N2741, N1587, N1405);
not NOT1 (N3312, N3293);
and AND4 (N3313, N3311, N1743, N1224, N410);
not NOT1 (N3314, N3307);
nor NOR4 (N3315, N3308, N2834, N1996, N2187);
buf BUF1 (N3316, N3313);
not NOT1 (N3317, N3312);
xor XOR2 (N3318, N3310, N551);
or OR3 (N3319, N3303, N1031, N1182);
and AND3 (N3320, N3319, N1228, N3210);
not NOT1 (N3321, N3309);
nand NAND3 (N3322, N3318, N214, N1007);
nand NAND3 (N3323, N3284, N959, N122);
xor XOR2 (N3324, N3306, N1928);
nand NAND4 (N3325, N3321, N2641, N946, N1362);
nand NAND2 (N3326, N3325, N360);
not NOT1 (N3327, N3326);
and AND2 (N3328, N3327, N2865);
xor XOR2 (N3329, N3322, N664);
xor XOR2 (N3330, N3305, N1958);
nand NAND3 (N3331, N3330, N151, N97);
buf BUF1 (N3332, N3315);
nor NOR4 (N3333, N3317, N1083, N2215, N1410);
buf BUF1 (N3334, N3324);
xor XOR2 (N3335, N3320, N577);
and AND4 (N3336, N3323, N2163, N2737, N2182);
xor XOR2 (N3337, N3333, N827);
nor NOR2 (N3338, N3336, N2696);
or OR2 (N3339, N3338, N2650);
or OR3 (N3340, N3329, N1672, N961);
nor NOR3 (N3341, N3334, N3136, N1932);
buf BUF1 (N3342, N3328);
buf BUF1 (N3343, N3341);
buf BUF1 (N3344, N3331);
xor XOR2 (N3345, N3337, N2841);
not NOT1 (N3346, N3342);
nand NAND3 (N3347, N3314, N3133, N1204);
not NOT1 (N3348, N3346);
xor XOR2 (N3349, N3332, N276);
nor NOR4 (N3350, N3348, N1283, N1046, N1628);
not NOT1 (N3351, N3316);
or OR2 (N3352, N3351, N2451);
and AND3 (N3353, N3335, N1203, N2162);
buf BUF1 (N3354, N3349);
not NOT1 (N3355, N3350);
not NOT1 (N3356, N3343);
not NOT1 (N3357, N3354);
or OR3 (N3358, N3355, N566, N3307);
nand NAND4 (N3359, N3356, N3225, N343, N3127);
xor XOR2 (N3360, N3359, N888);
nor NOR3 (N3361, N3344, N2602, N1339);
not NOT1 (N3362, N3345);
nor NOR3 (N3363, N3347, N1762, N1531);
nor NOR3 (N3364, N3360, N294, N704);
not NOT1 (N3365, N3352);
nor NOR4 (N3366, N3358, N2352, N3094, N2535);
nand NAND3 (N3367, N3365, N1086, N2931);
or OR4 (N3368, N3367, N1118, N1369, N2805);
nand NAND4 (N3369, N3357, N149, N981, N816);
and AND4 (N3370, N3363, N1519, N1052, N2262);
and AND4 (N3371, N3369, N484, N1988, N52);
or OR4 (N3372, N3353, N2492, N2719, N1063);
buf BUF1 (N3373, N3364);
buf BUF1 (N3374, N3361);
buf BUF1 (N3375, N3374);
or OR3 (N3376, N3371, N3051, N2108);
and AND2 (N3377, N3339, N454);
and AND3 (N3378, N3340, N1140, N683);
or OR4 (N3379, N3372, N3065, N1300, N1791);
not NOT1 (N3380, N3377);
xor XOR2 (N3381, N3378, N1881);
nand NAND4 (N3382, N3380, N1197, N1408, N1582);
xor XOR2 (N3383, N3381, N1379);
nand NAND4 (N3384, N3375, N688, N2163, N2129);
nand NAND3 (N3385, N3370, N2887, N2240);
nor NOR4 (N3386, N3382, N2747, N941, N3103);
nand NAND2 (N3387, N3362, N1629);
or OR2 (N3388, N3385, N72);
and AND2 (N3389, N3387, N850);
nor NOR4 (N3390, N3386, N2050, N2680, N829);
buf BUF1 (N3391, N3366);
buf BUF1 (N3392, N3368);
buf BUF1 (N3393, N3383);
nand NAND3 (N3394, N3376, N770, N982);
xor XOR2 (N3395, N3391, N2616);
xor XOR2 (N3396, N3392, N249);
xor XOR2 (N3397, N3373, N1963);
nor NOR4 (N3398, N3394, N2616, N1509, N1283);
nand NAND3 (N3399, N3388, N2648, N515);
nor NOR2 (N3400, N3395, N2198);
not NOT1 (N3401, N3384);
buf BUF1 (N3402, N3393);
not NOT1 (N3403, N3397);
or OR2 (N3404, N3402, N2277);
and AND4 (N3405, N3404, N1143, N66, N3173);
or OR3 (N3406, N3403, N83, N1542);
not NOT1 (N3407, N3398);
or OR3 (N3408, N3400, N1945, N798);
xor XOR2 (N3409, N3407, N847);
buf BUF1 (N3410, N3399);
or OR3 (N3411, N3409, N565, N1714);
and AND2 (N3412, N3396, N1452);
and AND3 (N3413, N3412, N3159, N1796);
buf BUF1 (N3414, N3406);
xor XOR2 (N3415, N3379, N770);
not NOT1 (N3416, N3410);
not NOT1 (N3417, N3401);
or OR3 (N3418, N3389, N2551, N2432);
buf BUF1 (N3419, N3417);
nand NAND3 (N3420, N3408, N2011, N1916);
xor XOR2 (N3421, N3416, N1585);
or OR2 (N3422, N3414, N2043);
xor XOR2 (N3423, N3411, N2973);
nand NAND2 (N3424, N3405, N162);
not NOT1 (N3425, N3419);
or OR3 (N3426, N3413, N851, N712);
or OR2 (N3427, N3426, N2262);
and AND2 (N3428, N3418, N3007);
or OR4 (N3429, N3428, N2728, N2908, N501);
nor NOR3 (N3430, N3423, N2910, N235);
xor XOR2 (N3431, N3421, N279);
xor XOR2 (N3432, N3422, N859);
buf BUF1 (N3433, N3415);
nand NAND4 (N3434, N3430, N77, N2843, N1946);
buf BUF1 (N3435, N3390);
nor NOR2 (N3436, N3431, N1074);
nand NAND4 (N3437, N3433, N928, N136, N82);
and AND3 (N3438, N3424, N3372, N2547);
and AND2 (N3439, N3437, N1680);
nor NOR4 (N3440, N3438, N2477, N462, N974);
nor NOR4 (N3441, N3440, N3359, N1202, N1860);
xor XOR2 (N3442, N3427, N3358);
buf BUF1 (N3443, N3441);
xor XOR2 (N3444, N3420, N2586);
nand NAND4 (N3445, N3436, N17, N521, N185);
and AND4 (N3446, N3429, N2177, N682, N1691);
buf BUF1 (N3447, N3434);
and AND4 (N3448, N3446, N3010, N2838, N3035);
buf BUF1 (N3449, N3432);
or OR3 (N3450, N3442, N2316, N1905);
not NOT1 (N3451, N3448);
nand NAND3 (N3452, N3449, N2141, N2631);
nor NOR3 (N3453, N3425, N2136, N2121);
or OR3 (N3454, N3439, N1020, N1180);
nor NOR3 (N3455, N3450, N1676, N313);
buf BUF1 (N3456, N3435);
nor NOR2 (N3457, N3455, N3159);
nand NAND2 (N3458, N3453, N2236);
and AND4 (N3459, N3447, N874, N1302, N2241);
not NOT1 (N3460, N3457);
nor NOR4 (N3461, N3459, N387, N2608, N1926);
nand NAND4 (N3462, N3452, N2046, N801, N2256);
nand NAND4 (N3463, N3444, N2981, N2232, N812);
or OR3 (N3464, N3463, N1512, N819);
nand NAND4 (N3465, N3454, N1304, N2128, N394);
buf BUF1 (N3466, N3465);
nor NOR3 (N3467, N3443, N1229, N1200);
and AND2 (N3468, N3461, N2948);
nor NOR2 (N3469, N3445, N248);
and AND2 (N3470, N3458, N2001);
not NOT1 (N3471, N3470);
or OR2 (N3472, N3462, N2588);
xor XOR2 (N3473, N3471, N2876);
nand NAND3 (N3474, N3473, N2462, N1677);
or OR3 (N3475, N3467, N81, N1595);
not NOT1 (N3476, N3456);
not NOT1 (N3477, N3474);
nor NOR3 (N3478, N3460, N2736, N1331);
buf BUF1 (N3479, N3477);
nand NAND3 (N3480, N3478, N403, N376);
nor NOR3 (N3481, N3468, N673, N386);
buf BUF1 (N3482, N3480);
and AND4 (N3483, N3475, N1391, N2292, N1161);
or OR2 (N3484, N3469, N496);
and AND4 (N3485, N3481, N3215, N2851, N1445);
or OR3 (N3486, N3476, N2139, N3392);
xor XOR2 (N3487, N3472, N3133);
or OR3 (N3488, N3485, N450, N1667);
xor XOR2 (N3489, N3483, N1807);
and AND3 (N3490, N3488, N52, N589);
nor NOR4 (N3491, N3487, N771, N296, N758);
xor XOR2 (N3492, N3484, N3485);
nand NAND3 (N3493, N3486, N1254, N2532);
xor XOR2 (N3494, N3493, N2269);
nand NAND3 (N3495, N3466, N1688, N414);
nor NOR2 (N3496, N3479, N59);
nand NAND2 (N3497, N3491, N972);
xor XOR2 (N3498, N3494, N2742);
not NOT1 (N3499, N3497);
nor NOR4 (N3500, N3451, N952, N932, N354);
xor XOR2 (N3501, N3490, N1166);
and AND2 (N3502, N3496, N1735);
nand NAND3 (N3503, N3492, N2124, N1689);
nor NOR4 (N3504, N3498, N771, N2113, N1019);
and AND3 (N3505, N3501, N2755, N3126);
nor NOR2 (N3506, N3489, N3433);
and AND3 (N3507, N3506, N578, N2630);
nand NAND3 (N3508, N3505, N1261, N2251);
and AND3 (N3509, N3504, N1787, N3180);
and AND4 (N3510, N3464, N2942, N760, N1657);
nor NOR4 (N3511, N3499, N1372, N1835, N1931);
or OR2 (N3512, N3510, N3385);
or OR3 (N3513, N3503, N763, N1940);
or OR2 (N3514, N3509, N1395);
buf BUF1 (N3515, N3511);
nor NOR4 (N3516, N3513, N177, N592, N2967);
nand NAND4 (N3517, N3482, N2107, N2496, N1994);
not NOT1 (N3518, N3507);
and AND3 (N3519, N3495, N3071, N1174);
and AND2 (N3520, N3516, N588);
not NOT1 (N3521, N3508);
nor NOR4 (N3522, N3500, N3499, N3385, N334);
or OR3 (N3523, N3522, N1115, N2213);
and AND4 (N3524, N3518, N1175, N514, N2926);
and AND2 (N3525, N3502, N266);
or OR2 (N3526, N3521, N2417);
not NOT1 (N3527, N3519);
and AND2 (N3528, N3524, N2747);
not NOT1 (N3529, N3525);
buf BUF1 (N3530, N3523);
or OR4 (N3531, N3526, N1415, N525, N656);
xor XOR2 (N3532, N3528, N3477);
nor NOR3 (N3533, N3530, N233, N2136);
not NOT1 (N3534, N3532);
buf BUF1 (N3535, N3517);
and AND3 (N3536, N3535, N1252, N1672);
or OR3 (N3537, N3534, N1365, N563);
nor NOR4 (N3538, N3515, N3272, N1873, N1212);
or OR2 (N3539, N3520, N2215);
or OR4 (N3540, N3529, N3110, N3182, N2674);
buf BUF1 (N3541, N3537);
and AND4 (N3542, N3540, N3029, N2453, N2108);
buf BUF1 (N3543, N3527);
and AND4 (N3544, N3531, N1020, N1226, N1987);
nand NAND3 (N3545, N3541, N3324, N144);
nor NOR4 (N3546, N3542, N1701, N3430, N2691);
buf BUF1 (N3547, N3536);
nor NOR3 (N3548, N3543, N2306, N1263);
not NOT1 (N3549, N3546);
not NOT1 (N3550, N3548);
xor XOR2 (N3551, N3538, N1806);
and AND2 (N3552, N3550, N2091);
buf BUF1 (N3553, N3512);
or OR2 (N3554, N3549, N57);
not NOT1 (N3555, N3553);
not NOT1 (N3556, N3514);
nor NOR2 (N3557, N3551, N56);
and AND2 (N3558, N3539, N2441);
nand NAND2 (N3559, N3552, N3189);
nand NAND2 (N3560, N3559, N32);
and AND2 (N3561, N3554, N2339);
and AND3 (N3562, N3547, N1969, N2871);
nor NOR2 (N3563, N3533, N2674);
xor XOR2 (N3564, N3560, N1988);
not NOT1 (N3565, N3558);
not NOT1 (N3566, N3563);
and AND4 (N3567, N3561, N2054, N639, N1444);
buf BUF1 (N3568, N3564);
nor NOR4 (N3569, N3545, N2502, N2208, N1758);
nor NOR3 (N3570, N3555, N2353, N3267);
or OR2 (N3571, N3566, N29);
xor XOR2 (N3572, N3567, N3363);
nor NOR4 (N3573, N3544, N2177, N2704, N2791);
not NOT1 (N3574, N3570);
xor XOR2 (N3575, N3571, N3084);
xor XOR2 (N3576, N3572, N2264);
nand NAND3 (N3577, N3573, N1859, N767);
and AND3 (N3578, N3556, N814, N2687);
and AND4 (N3579, N3576, N1666, N2838, N3550);
not NOT1 (N3580, N3557);
not NOT1 (N3581, N3577);
not NOT1 (N3582, N3579);
buf BUF1 (N3583, N3582);
or OR4 (N3584, N3568, N1092, N374, N1595);
buf BUF1 (N3585, N3565);
and AND3 (N3586, N3583, N1783, N1902);
or OR4 (N3587, N3586, N2302, N2373, N2887);
xor XOR2 (N3588, N3581, N565);
nand NAND2 (N3589, N3588, N2402);
or OR4 (N3590, N3584, N2349, N2103, N2440);
or OR4 (N3591, N3578, N330, N1390, N426);
and AND3 (N3592, N3589, N89, N1078);
or OR3 (N3593, N3587, N3131, N2650);
nor NOR4 (N3594, N3592, N2710, N1763, N567);
nand NAND3 (N3595, N3593, N343, N2499);
not NOT1 (N3596, N3580);
nand NAND2 (N3597, N3585, N2206);
nand NAND4 (N3598, N3597, N888, N1113, N2726);
not NOT1 (N3599, N3590);
not NOT1 (N3600, N3596);
buf BUF1 (N3601, N3575);
and AND4 (N3602, N3598, N960, N1784, N1123);
buf BUF1 (N3603, N3600);
xor XOR2 (N3604, N3591, N1202);
or OR4 (N3605, N3562, N489, N3281, N360);
or OR3 (N3606, N3605, N1466, N1515);
nor NOR4 (N3607, N3594, N674, N756, N2257);
nor NOR4 (N3608, N3602, N3022, N3148, N2052);
buf BUF1 (N3609, N3607);
not NOT1 (N3610, N3603);
not NOT1 (N3611, N3604);
buf BUF1 (N3612, N3610);
nand NAND3 (N3613, N3611, N2302, N35);
nand NAND4 (N3614, N3599, N1728, N1221, N1547);
not NOT1 (N3615, N3612);
or OR4 (N3616, N3606, N918, N2692, N3492);
xor XOR2 (N3617, N3613, N664);
not NOT1 (N3618, N3595);
nand NAND3 (N3619, N3574, N838, N449);
xor XOR2 (N3620, N3601, N927);
and AND4 (N3621, N3616, N2668, N1222, N69);
nand NAND2 (N3622, N3614, N3447);
not NOT1 (N3623, N3569);
and AND3 (N3624, N3608, N1369, N2023);
nor NOR3 (N3625, N3617, N1314, N2618);
nor NOR4 (N3626, N3609, N976, N2425, N2202);
or OR2 (N3627, N3619, N3209);
xor XOR2 (N3628, N3627, N2968);
not NOT1 (N3629, N3628);
and AND3 (N3630, N3625, N1797, N139);
nor NOR3 (N3631, N3629, N1739, N1536);
nand NAND4 (N3632, N3624, N3112, N649, N2095);
xor XOR2 (N3633, N3615, N1743);
or OR2 (N3634, N3622, N3098);
and AND3 (N3635, N3620, N3582, N3172);
xor XOR2 (N3636, N3632, N2514);
nand NAND4 (N3637, N3636, N2740, N3345, N3545);
xor XOR2 (N3638, N3637, N796);
xor XOR2 (N3639, N3626, N113);
buf BUF1 (N3640, N3633);
xor XOR2 (N3641, N3635, N35);
xor XOR2 (N3642, N3623, N2181);
xor XOR2 (N3643, N3638, N2475);
not NOT1 (N3644, N3641);
nand NAND3 (N3645, N3630, N3442, N715);
not NOT1 (N3646, N3644);
not NOT1 (N3647, N3639);
buf BUF1 (N3648, N3645);
buf BUF1 (N3649, N3631);
or OR3 (N3650, N3634, N3589, N2361);
nand NAND3 (N3651, N3650, N3059, N3108);
or OR3 (N3652, N3640, N3221, N3579);
nor NOR4 (N3653, N3651, N1642, N1048, N3383);
xor XOR2 (N3654, N3643, N2458);
not NOT1 (N3655, N3654);
xor XOR2 (N3656, N3642, N1472);
and AND4 (N3657, N3618, N208, N111, N2329);
not NOT1 (N3658, N3656);
not NOT1 (N3659, N3655);
and AND2 (N3660, N3659, N366);
not NOT1 (N3661, N3652);
nor NOR3 (N3662, N3648, N849, N3017);
xor XOR2 (N3663, N3658, N3379);
not NOT1 (N3664, N3660);
xor XOR2 (N3665, N3646, N2240);
not NOT1 (N3666, N3662);
buf BUF1 (N3667, N3647);
not NOT1 (N3668, N3661);
nor NOR3 (N3669, N3664, N998, N3658);
and AND3 (N3670, N3649, N879, N2411);
or OR3 (N3671, N3669, N2839, N3413);
not NOT1 (N3672, N3621);
not NOT1 (N3673, N3665);
or OR3 (N3674, N3668, N40, N1265);
not NOT1 (N3675, N3663);
xor XOR2 (N3676, N3670, N1348);
or OR2 (N3677, N3653, N1661);
nand NAND3 (N3678, N3666, N3183, N1793);
not NOT1 (N3679, N3667);
and AND2 (N3680, N3677, N1191);
or OR4 (N3681, N3680, N2001, N1973, N3151);
nand NAND2 (N3682, N3673, N1246);
not NOT1 (N3683, N3672);
buf BUF1 (N3684, N3671);
nor NOR2 (N3685, N3682, N1893);
and AND4 (N3686, N3683, N560, N2258, N2405);
or OR4 (N3687, N3686, N1872, N3373, N3554);
xor XOR2 (N3688, N3679, N2806);
nand NAND2 (N3689, N3685, N3317);
not NOT1 (N3690, N3678);
buf BUF1 (N3691, N3684);
xor XOR2 (N3692, N3688, N618);
xor XOR2 (N3693, N3657, N2056);
nand NAND4 (N3694, N3689, N2004, N2355, N500);
buf BUF1 (N3695, N3690);
or OR4 (N3696, N3674, N2816, N3062, N471);
or OR3 (N3697, N3691, N110, N406);
xor XOR2 (N3698, N3696, N972);
and AND2 (N3699, N3676, N1230);
not NOT1 (N3700, N3687);
not NOT1 (N3701, N3699);
buf BUF1 (N3702, N3675);
and AND3 (N3703, N3695, N1730, N1719);
or OR3 (N3704, N3701, N2343, N719);
not NOT1 (N3705, N3704);
buf BUF1 (N3706, N3705);
and AND4 (N3707, N3692, N970, N3295, N3027);
nand NAND4 (N3708, N3693, N2230, N1481, N2283);
xor XOR2 (N3709, N3707, N3202);
or OR4 (N3710, N3700, N91, N490, N1476);
or OR3 (N3711, N3697, N1807, N1935);
nor NOR4 (N3712, N3706, N3022, N40, N3493);
nand NAND3 (N3713, N3708, N1688, N253);
not NOT1 (N3714, N3681);
buf BUF1 (N3715, N3711);
not NOT1 (N3716, N3712);
buf BUF1 (N3717, N3698);
xor XOR2 (N3718, N3709, N3610);
buf BUF1 (N3719, N3710);
not NOT1 (N3720, N3716);
nand NAND4 (N3721, N3694, N3252, N1947, N2784);
or OR4 (N3722, N3714, N1624, N2562, N2565);
or OR3 (N3723, N3713, N58, N1199);
and AND4 (N3724, N3715, N2576, N2378, N2857);
and AND2 (N3725, N3702, N1735);
not NOT1 (N3726, N3719);
and AND4 (N3727, N3721, N1791, N1097, N293);
or OR4 (N3728, N3723, N491, N3370, N1448);
nand NAND4 (N3729, N3727, N2282, N2156, N3226);
nand NAND2 (N3730, N3726, N2473);
nand NAND2 (N3731, N3722, N1848);
xor XOR2 (N3732, N3731, N1029);
or OR2 (N3733, N3717, N873);
buf BUF1 (N3734, N3725);
nor NOR3 (N3735, N3724, N1528, N1019);
not NOT1 (N3736, N3733);
nand NAND4 (N3737, N3718, N1947, N1452, N2929);
nand NAND3 (N3738, N3730, N275, N2096);
xor XOR2 (N3739, N3737, N1772);
buf BUF1 (N3740, N3720);
nor NOR3 (N3741, N3729, N1727, N2679);
nor NOR3 (N3742, N3740, N3455, N930);
buf BUF1 (N3743, N3734);
xor XOR2 (N3744, N3728, N117);
xor XOR2 (N3745, N3735, N136);
nor NOR4 (N3746, N3741, N3396, N1855, N837);
nand NAND2 (N3747, N3742, N2298);
nand NAND4 (N3748, N3746, N1311, N536, N1466);
nor NOR4 (N3749, N3747, N1221, N2974, N3437);
or OR4 (N3750, N3745, N3609, N842, N2006);
buf BUF1 (N3751, N3736);
and AND3 (N3752, N3750, N181, N3672);
nand NAND3 (N3753, N3732, N2770, N1541);
nor NOR4 (N3754, N3751, N285, N451, N2350);
or OR4 (N3755, N3743, N1746, N3467, N1517);
or OR2 (N3756, N3744, N176);
nor NOR4 (N3757, N3703, N3482, N2819, N1303);
xor XOR2 (N3758, N3753, N2439);
buf BUF1 (N3759, N3754);
nor NOR3 (N3760, N3755, N116, N2717);
nor NOR3 (N3761, N3759, N445, N1275);
not NOT1 (N3762, N3739);
xor XOR2 (N3763, N3748, N1580);
or OR3 (N3764, N3756, N1722, N1647);
and AND4 (N3765, N3760, N203, N301, N2876);
xor XOR2 (N3766, N3761, N2585);
not NOT1 (N3767, N3738);
or OR2 (N3768, N3764, N3486);
and AND3 (N3769, N3762, N1052, N1349);
nand NAND3 (N3770, N3757, N3561, N75);
and AND4 (N3771, N3767, N1561, N1618, N1782);
nand NAND2 (N3772, N3768, N3503);
or OR4 (N3773, N3749, N2766, N2917, N740);
not NOT1 (N3774, N3766);
not NOT1 (N3775, N3773);
nor NOR4 (N3776, N3765, N495, N1748, N2056);
nor NOR2 (N3777, N3758, N708);
nand NAND3 (N3778, N3777, N2846, N1116);
nand NAND2 (N3779, N3769, N3452);
xor XOR2 (N3780, N3774, N712);
or OR4 (N3781, N3770, N2190, N1627, N2569);
and AND4 (N3782, N3778, N2548, N784, N1925);
buf BUF1 (N3783, N3772);
buf BUF1 (N3784, N3783);
nor NOR3 (N3785, N3771, N3519, N1684);
and AND4 (N3786, N3782, N2371, N1133, N3475);
or OR2 (N3787, N3784, N592);
or OR3 (N3788, N3779, N2471, N1307);
or OR4 (N3789, N3780, N3367, N2550, N625);
nand NAND3 (N3790, N3776, N1918, N1408);
not NOT1 (N3791, N3763);
xor XOR2 (N3792, N3781, N1871);
not NOT1 (N3793, N3785);
and AND4 (N3794, N3790, N2961, N3050, N1765);
not NOT1 (N3795, N3786);
nor NOR3 (N3796, N3788, N2373, N1875);
nor NOR4 (N3797, N3787, N1093, N3238, N1112);
buf BUF1 (N3798, N3792);
not NOT1 (N3799, N3795);
buf BUF1 (N3800, N3752);
nor NOR4 (N3801, N3794, N2456, N2496, N676);
not NOT1 (N3802, N3798);
xor XOR2 (N3803, N3796, N855);
nor NOR3 (N3804, N3793, N636, N751);
nand NAND3 (N3805, N3791, N1380, N806);
or OR4 (N3806, N3805, N25, N561, N2762);
xor XOR2 (N3807, N3801, N3457);
and AND2 (N3808, N3800, N2693);
nor NOR4 (N3809, N3797, N1355, N48, N2888);
and AND3 (N3810, N3809, N3252, N1276);
nor NOR3 (N3811, N3810, N1195, N1036);
buf BUF1 (N3812, N3803);
or OR4 (N3813, N3775, N3129, N551, N1280);
nand NAND4 (N3814, N3802, N23, N3213, N845);
xor XOR2 (N3815, N3808, N1364);
and AND3 (N3816, N3804, N2404, N1851);
nand NAND3 (N3817, N3812, N232, N1640);
buf BUF1 (N3818, N3807);
nand NAND2 (N3819, N3789, N3035);
nand NAND3 (N3820, N3813, N1029, N2730);
buf BUF1 (N3821, N3811);
not NOT1 (N3822, N3816);
xor XOR2 (N3823, N3817, N2560);
buf BUF1 (N3824, N3823);
not NOT1 (N3825, N3822);
or OR4 (N3826, N3815, N1224, N846, N636);
and AND3 (N3827, N3825, N2283, N2560);
nand NAND2 (N3828, N3806, N53);
or OR3 (N3829, N3819, N2082, N680);
not NOT1 (N3830, N3824);
nand NAND4 (N3831, N3818, N2525, N825, N1962);
not NOT1 (N3832, N3820);
not NOT1 (N3833, N3828);
nand NAND4 (N3834, N3829, N672, N3468, N1892);
buf BUF1 (N3835, N3827);
and AND4 (N3836, N3821, N3036, N372, N3145);
buf BUF1 (N3837, N3826);
not NOT1 (N3838, N3799);
not NOT1 (N3839, N3814);
nor NOR3 (N3840, N3833, N895, N2410);
buf BUF1 (N3841, N3837);
buf BUF1 (N3842, N3836);
or OR2 (N3843, N3841, N3310);
xor XOR2 (N3844, N3840, N3713);
and AND3 (N3845, N3834, N2917, N3622);
nor NOR3 (N3846, N3832, N2385, N2079);
nand NAND2 (N3847, N3839, N3816);
nor NOR2 (N3848, N3846, N1443);
not NOT1 (N3849, N3848);
xor XOR2 (N3850, N3849, N1584);
xor XOR2 (N3851, N3842, N440);
nor NOR3 (N3852, N3850, N3831, N743);
xor XOR2 (N3853, N2536, N3444);
xor XOR2 (N3854, N3853, N2792);
nand NAND2 (N3855, N3843, N1444);
or OR3 (N3856, N3844, N368, N1593);
not NOT1 (N3857, N3845);
not NOT1 (N3858, N3854);
xor XOR2 (N3859, N3851, N1884);
xor XOR2 (N3860, N3855, N1779);
buf BUF1 (N3861, N3858);
not NOT1 (N3862, N3856);
buf BUF1 (N3863, N3862);
not NOT1 (N3864, N3835);
and AND4 (N3865, N3863, N3355, N295, N1911);
nand NAND2 (N3866, N3865, N332);
or OR2 (N3867, N3852, N2791);
nor NOR3 (N3868, N3861, N470, N1189);
nand NAND3 (N3869, N3867, N346, N555);
nand NAND4 (N3870, N3860, N2897, N2687, N2376);
buf BUF1 (N3871, N3857);
buf BUF1 (N3872, N3847);
not NOT1 (N3873, N3859);
and AND2 (N3874, N3873, N1734);
or OR2 (N3875, N3864, N1412);
nor NOR2 (N3876, N3872, N2646);
not NOT1 (N3877, N3868);
and AND2 (N3878, N3871, N1845);
nor NOR2 (N3879, N3878, N3249);
xor XOR2 (N3880, N3874, N910);
nand NAND4 (N3881, N3830, N433, N1362, N1166);
and AND4 (N3882, N3880, N2500, N3580, N2619);
and AND3 (N3883, N3882, N1727, N3408);
xor XOR2 (N3884, N3883, N1320);
nor NOR4 (N3885, N3876, N3779, N3529, N3045);
xor XOR2 (N3886, N3838, N2440);
buf BUF1 (N3887, N3866);
nor NOR2 (N3888, N3877, N3580);
and AND3 (N3889, N3875, N1689, N2522);
nor NOR3 (N3890, N3884, N1520, N1433);
and AND4 (N3891, N3869, N3068, N2241, N2930);
nor NOR2 (N3892, N3887, N756);
nand NAND4 (N3893, N3892, N1635, N3460, N3525);
xor XOR2 (N3894, N3891, N334);
nand NAND4 (N3895, N3885, N1217, N3578, N1664);
or OR3 (N3896, N3879, N3868, N2519);
buf BUF1 (N3897, N3895);
xor XOR2 (N3898, N3897, N1292);
xor XOR2 (N3899, N3893, N2498);
nand NAND4 (N3900, N3889, N3841, N3854, N3163);
or OR4 (N3901, N3881, N3521, N2539, N788);
and AND2 (N3902, N3900, N2424);
not NOT1 (N3903, N3898);
not NOT1 (N3904, N3903);
buf BUF1 (N3905, N3888);
nand NAND3 (N3906, N3902, N3198, N1392);
xor XOR2 (N3907, N3904, N3164);
not NOT1 (N3908, N3890);
or OR4 (N3909, N3908, N1107, N936, N2888);
xor XOR2 (N3910, N3906, N3827);
nand NAND2 (N3911, N3896, N2386);
buf BUF1 (N3912, N3899);
nor NOR4 (N3913, N3907, N2639, N2660, N1840);
nor NOR4 (N3914, N3870, N2019, N1465, N1216);
buf BUF1 (N3915, N3905);
and AND2 (N3916, N3912, N1356);
nor NOR3 (N3917, N3911, N385, N1329);
xor XOR2 (N3918, N3913, N1089);
xor XOR2 (N3919, N3909, N2253);
xor XOR2 (N3920, N3915, N1711);
or OR2 (N3921, N3901, N3318);
and AND4 (N3922, N3918, N2145, N3140, N2083);
nor NOR2 (N3923, N3886, N2618);
nor NOR4 (N3924, N3919, N1118, N2382, N2167);
nor NOR3 (N3925, N3914, N3149, N11);
not NOT1 (N3926, N3925);
and AND4 (N3927, N3910, N1145, N1750, N3266);
nand NAND4 (N3928, N3922, N1944, N3419, N1911);
or OR3 (N3929, N3920, N1137, N2370);
nand NAND4 (N3930, N3923, N2022, N2510, N2062);
nand NAND3 (N3931, N3921, N1031, N393);
nor NOR4 (N3932, N3924, N1318, N406, N1109);
xor XOR2 (N3933, N3929, N3890);
buf BUF1 (N3934, N3917);
nand NAND4 (N3935, N3930, N2734, N44, N854);
or OR2 (N3936, N3933, N3831);
buf BUF1 (N3937, N3927);
nor NOR4 (N3938, N3931, N260, N3456, N3554);
nor NOR3 (N3939, N3934, N1312, N271);
buf BUF1 (N3940, N3936);
and AND4 (N3941, N3938, N1610, N2788, N2125);
xor XOR2 (N3942, N3937, N3665);
nand NAND2 (N3943, N3926, N685);
buf BUF1 (N3944, N3939);
buf BUF1 (N3945, N3894);
nand NAND3 (N3946, N3928, N2560, N264);
not NOT1 (N3947, N3916);
nor NOR3 (N3948, N3944, N1527, N3482);
xor XOR2 (N3949, N3942, N1820);
nor NOR2 (N3950, N3945, N525);
xor XOR2 (N3951, N3949, N1471);
xor XOR2 (N3952, N3946, N2415);
not NOT1 (N3953, N3940);
and AND4 (N3954, N3932, N581, N3864, N1630);
buf BUF1 (N3955, N3947);
buf BUF1 (N3956, N3948);
and AND3 (N3957, N3953, N664, N3651);
or OR3 (N3958, N3957, N483, N2639);
xor XOR2 (N3959, N3951, N3142);
not NOT1 (N3960, N3950);
xor XOR2 (N3961, N3935, N1748);
buf BUF1 (N3962, N3952);
nor NOR4 (N3963, N3941, N1476, N241, N2067);
and AND3 (N3964, N3954, N480, N3702);
not NOT1 (N3965, N3956);
nand NAND4 (N3966, N3960, N151, N3563, N512);
xor XOR2 (N3967, N3966, N999);
xor XOR2 (N3968, N3955, N263);
not NOT1 (N3969, N3967);
buf BUF1 (N3970, N3962);
buf BUF1 (N3971, N3965);
not NOT1 (N3972, N3963);
nor NOR2 (N3973, N3943, N2196);
nor NOR3 (N3974, N3964, N825, N563);
nand NAND2 (N3975, N3972, N932);
or OR2 (N3976, N3970, N3427);
not NOT1 (N3977, N3959);
nand NAND4 (N3978, N3977, N1898, N2555, N3458);
buf BUF1 (N3979, N3971);
not NOT1 (N3980, N3975);
and AND4 (N3981, N3976, N2765, N1568, N2654);
buf BUF1 (N3982, N3979);
and AND4 (N3983, N3961, N928, N1732, N1249);
or OR2 (N3984, N3968, N1688);
nand NAND2 (N3985, N3981, N2340);
nor NOR3 (N3986, N3969, N1761, N3670);
xor XOR2 (N3987, N3982, N315);
not NOT1 (N3988, N3987);
not NOT1 (N3989, N3986);
or OR3 (N3990, N3978, N2620, N2981);
or OR2 (N3991, N3983, N1259);
xor XOR2 (N3992, N3991, N1911);
nand NAND2 (N3993, N3992, N145);
nand NAND4 (N3994, N3988, N1122, N2572, N1933);
nor NOR4 (N3995, N3974, N2604, N1412, N2951);
xor XOR2 (N3996, N3989, N1175);
xor XOR2 (N3997, N3996, N2456);
or OR3 (N3998, N3958, N1050, N857);
xor XOR2 (N3999, N3998, N796);
buf BUF1 (N4000, N3994);
not NOT1 (N4001, N3990);
buf BUF1 (N4002, N3980);
buf BUF1 (N4003, N3997);
or OR2 (N4004, N3995, N815);
and AND4 (N4005, N3999, N1164, N3398, N1557);
nand NAND4 (N4006, N3993, N2450, N1230, N2122);
xor XOR2 (N4007, N3973, N3646);
xor XOR2 (N4008, N4005, N707);
nor NOR2 (N4009, N4001, N3462);
xor XOR2 (N4010, N4008, N1470);
xor XOR2 (N4011, N4004, N2305);
nand NAND3 (N4012, N3985, N318, N2337);
nand NAND4 (N4013, N4003, N3500, N3906, N2665);
or OR2 (N4014, N4009, N1083);
or OR3 (N4015, N4012, N3328, N3949);
buf BUF1 (N4016, N4006);
and AND2 (N4017, N4015, N3800);
nor NOR4 (N4018, N4000, N328, N697, N260);
not NOT1 (N4019, N4018);
and AND2 (N4020, N4010, N1779);
and AND4 (N4021, N4014, N2531, N2097, N3506);
and AND3 (N4022, N4017, N3913, N2831);
buf BUF1 (N4023, N4021);
buf BUF1 (N4024, N4023);
xor XOR2 (N4025, N4024, N1613);
nand NAND4 (N4026, N4007, N2146, N3972, N3995);
not NOT1 (N4027, N4013);
xor XOR2 (N4028, N4016, N749);
xor XOR2 (N4029, N4026, N3314);
buf BUF1 (N4030, N4019);
not NOT1 (N4031, N4020);
nand NAND2 (N4032, N4011, N2403);
xor XOR2 (N4033, N4022, N177);
nand NAND4 (N4034, N4030, N3524, N2961, N1393);
or OR4 (N4035, N4002, N1914, N2956, N2469);
not NOT1 (N4036, N4027);
nand NAND4 (N4037, N4034, N90, N1456, N2235);
or OR4 (N4038, N4028, N754, N3202, N932);
nand NAND4 (N4039, N4031, N809, N1777, N194);
nand NAND4 (N4040, N4038, N3312, N2476, N3745);
nand NAND2 (N4041, N3984, N3570);
xor XOR2 (N4042, N4041, N1394);
xor XOR2 (N4043, N4029, N363);
not NOT1 (N4044, N4025);
buf BUF1 (N4045, N4039);
or OR3 (N4046, N4033, N3009, N2639);
and AND2 (N4047, N4044, N1052);
nor NOR2 (N4048, N4040, N2092);
buf BUF1 (N4049, N4048);
and AND4 (N4050, N4035, N2113, N2951, N1955);
or OR3 (N4051, N4032, N2994, N842);
or OR4 (N4052, N4043, N3448, N2172, N1008);
or OR4 (N4053, N4052, N1202, N1509, N2780);
nand NAND3 (N4054, N4046, N880, N3602);
not NOT1 (N4055, N4036);
or OR3 (N4056, N4053, N3684, N2557);
or OR3 (N4057, N4047, N1994, N2069);
and AND3 (N4058, N4057, N521, N264);
buf BUF1 (N4059, N4058);
and AND3 (N4060, N4037, N3789, N1724);
and AND4 (N4061, N4045, N266, N2919, N1198);
nor NOR3 (N4062, N4061, N516, N969);
nand NAND3 (N4063, N4049, N1122, N644);
not NOT1 (N4064, N4060);
xor XOR2 (N4065, N4056, N18);
or OR2 (N4066, N4050, N1163);
buf BUF1 (N4067, N4055);
and AND4 (N4068, N4051, N2585, N449, N608);
nor NOR3 (N4069, N4066, N1728, N2434);
not NOT1 (N4070, N4067);
and AND2 (N4071, N4070, N461);
and AND4 (N4072, N4054, N1451, N2069, N196);
buf BUF1 (N4073, N4071);
xor XOR2 (N4074, N4073, N2746);
xor XOR2 (N4075, N4064, N3202);
not NOT1 (N4076, N4059);
xor XOR2 (N4077, N4075, N4000);
nand NAND2 (N4078, N4076, N22);
xor XOR2 (N4079, N4062, N1624);
nand NAND4 (N4080, N4079, N1260, N2644, N1791);
nor NOR3 (N4081, N4077, N359, N432);
not NOT1 (N4082, N4069);
xor XOR2 (N4083, N4065, N2848);
nor NOR2 (N4084, N4042, N3535);
xor XOR2 (N4085, N4074, N2456);
nand NAND4 (N4086, N4072, N3790, N2173, N2079);
or OR3 (N4087, N4085, N1119, N1046);
not NOT1 (N4088, N4086);
nand NAND3 (N4089, N4081, N326, N1681);
xor XOR2 (N4090, N4082, N1252);
buf BUF1 (N4091, N4063);
nand NAND4 (N4092, N4080, N787, N2757, N1067);
not NOT1 (N4093, N4078);
nand NAND3 (N4094, N4089, N3167, N2851);
or OR3 (N4095, N4087, N2353, N117);
nor NOR3 (N4096, N4084, N914, N2843);
not NOT1 (N4097, N4068);
nand NAND4 (N4098, N4096, N765, N2307, N3987);
not NOT1 (N4099, N4088);
buf BUF1 (N4100, N4090);
not NOT1 (N4101, N4097);
nor NOR3 (N4102, N4091, N1851, N3621);
nand NAND4 (N4103, N4095, N3084, N3188, N605);
or OR3 (N4104, N4102, N3431, N2873);
not NOT1 (N4105, N4099);
xor XOR2 (N4106, N4093, N568);
nand NAND2 (N4107, N4105, N2689);
and AND4 (N4108, N4100, N2234, N1581, N1454);
buf BUF1 (N4109, N4103);
buf BUF1 (N4110, N4107);
xor XOR2 (N4111, N4108, N2748);
and AND2 (N4112, N4101, N2533);
and AND4 (N4113, N4094, N3259, N398, N92);
or OR3 (N4114, N4112, N2170, N2809);
xor XOR2 (N4115, N4104, N1118);
not NOT1 (N4116, N4111);
buf BUF1 (N4117, N4106);
buf BUF1 (N4118, N4110);
xor XOR2 (N4119, N4116, N83);
not NOT1 (N4120, N4109);
buf BUF1 (N4121, N4119);
nand NAND3 (N4122, N4098, N812, N2688);
buf BUF1 (N4123, N4118);
and AND4 (N4124, N4113, N1616, N258, N111);
nand NAND3 (N4125, N4117, N542, N381);
nand NAND4 (N4126, N4124, N2518, N2614, N1853);
xor XOR2 (N4127, N4115, N2034);
not NOT1 (N4128, N4083);
xor XOR2 (N4129, N4120, N1739);
xor XOR2 (N4130, N4126, N2060);
nor NOR3 (N4131, N4128, N2486, N3329);
nand NAND4 (N4132, N4122, N1999, N3690, N2968);
not NOT1 (N4133, N4114);
or OR3 (N4134, N4092, N2191, N626);
or OR2 (N4135, N4129, N3330);
and AND3 (N4136, N4127, N2019, N1443);
not NOT1 (N4137, N4125);
buf BUF1 (N4138, N4133);
or OR3 (N4139, N4132, N1870, N3377);
buf BUF1 (N4140, N4137);
nor NOR2 (N4141, N4139, N1031);
or OR3 (N4142, N4121, N3246, N476);
nand NAND4 (N4143, N4141, N3874, N2772, N1219);
buf BUF1 (N4144, N4136);
not NOT1 (N4145, N4123);
nor NOR2 (N4146, N4142, N770);
and AND3 (N4147, N4134, N1611, N3909);
nor NOR4 (N4148, N4145, N1335, N1210, N1867);
xor XOR2 (N4149, N4131, N2390);
not NOT1 (N4150, N4130);
or OR4 (N4151, N4143, N3063, N600, N166);
buf BUF1 (N4152, N4135);
nor NOR3 (N4153, N4147, N3493, N2554);
buf BUF1 (N4154, N4149);
nor NOR4 (N4155, N4153, N3654, N4137, N1845);
nor NOR2 (N4156, N4140, N3801);
and AND3 (N4157, N4151, N3842, N2695);
or OR2 (N4158, N4148, N751);
nor NOR3 (N4159, N4154, N1596, N1865);
nand NAND3 (N4160, N4159, N1015, N1540);
nand NAND2 (N4161, N4156, N379);
buf BUF1 (N4162, N4157);
buf BUF1 (N4163, N4160);
buf BUF1 (N4164, N4152);
nand NAND4 (N4165, N4138, N2229, N3822, N1515);
and AND4 (N4166, N4155, N3161, N844, N1699);
nor NOR4 (N4167, N4166, N605, N3385, N3491);
nor NOR2 (N4168, N4167, N3277);
nor NOR2 (N4169, N4161, N2811);
or OR2 (N4170, N4144, N690);
and AND2 (N4171, N4163, N638);
xor XOR2 (N4172, N4171, N3993);
not NOT1 (N4173, N4150);
xor XOR2 (N4174, N4173, N21);
nor NOR4 (N4175, N4168, N3509, N4060, N3044);
or OR3 (N4176, N4165, N4050, N119);
buf BUF1 (N4177, N4146);
and AND3 (N4178, N4172, N1508, N2158);
and AND4 (N4179, N4170, N2173, N3319, N2931);
not NOT1 (N4180, N4178);
buf BUF1 (N4181, N4158);
nand NAND2 (N4182, N4177, N1189);
nand NAND3 (N4183, N4181, N3605, N558);
buf BUF1 (N4184, N4162);
or OR3 (N4185, N4180, N2114, N1526);
xor XOR2 (N4186, N4185, N2474);
nand NAND2 (N4187, N4169, N1212);
xor XOR2 (N4188, N4174, N2099);
not NOT1 (N4189, N4184);
and AND3 (N4190, N4188, N2163, N912);
buf BUF1 (N4191, N4190);
buf BUF1 (N4192, N4191);
nor NOR2 (N4193, N4179, N1607);
and AND3 (N4194, N4175, N1146, N398);
not NOT1 (N4195, N4176);
nor NOR4 (N4196, N4164, N1635, N2085, N3265);
buf BUF1 (N4197, N4183);
nand NAND2 (N4198, N4195, N47);
buf BUF1 (N4199, N4186);
nor NOR2 (N4200, N4197, N3819);
nand NAND4 (N4201, N4192, N2028, N3829, N1764);
not NOT1 (N4202, N4198);
buf BUF1 (N4203, N4199);
nor NOR2 (N4204, N4196, N3596);
nor NOR2 (N4205, N4189, N1932);
or OR2 (N4206, N4205, N555);
buf BUF1 (N4207, N4202);
nor NOR3 (N4208, N4201, N3146, N1583);
and AND3 (N4209, N4194, N223, N5);
not NOT1 (N4210, N4209);
or OR2 (N4211, N4187, N4191);
xor XOR2 (N4212, N4200, N991);
nand NAND2 (N4213, N4206, N951);
and AND4 (N4214, N4212, N1173, N3107, N2654);
and AND4 (N4215, N4203, N1247, N3002, N3678);
or OR2 (N4216, N4215, N977);
or OR4 (N4217, N4211, N1408, N318, N3895);
xor XOR2 (N4218, N4208, N3835);
xor XOR2 (N4219, N4204, N3529);
nor NOR4 (N4220, N4193, N1304, N2502, N4097);
nor NOR4 (N4221, N4217, N478, N767, N2657);
or OR2 (N4222, N4216, N4022);
and AND3 (N4223, N4220, N1060, N1344);
or OR2 (N4224, N4223, N2325);
or OR4 (N4225, N4221, N743, N722, N659);
and AND3 (N4226, N4207, N2287, N3309);
xor XOR2 (N4227, N4218, N2429);
nor NOR2 (N4228, N4219, N711);
not NOT1 (N4229, N4225);
or OR4 (N4230, N4182, N2369, N1330, N4003);
not NOT1 (N4231, N4227);
nor NOR4 (N4232, N4228, N1334, N158, N1410);
not NOT1 (N4233, N4224);
xor XOR2 (N4234, N4232, N4177);
nand NAND4 (N4235, N4222, N1721, N237, N1165);
xor XOR2 (N4236, N4230, N718);
xor XOR2 (N4237, N4226, N422);
xor XOR2 (N4238, N4229, N2830);
buf BUF1 (N4239, N4233);
xor XOR2 (N4240, N4231, N2224);
nor NOR4 (N4241, N4235, N229, N3697, N331);
not NOT1 (N4242, N4238);
xor XOR2 (N4243, N4214, N4075);
nand NAND4 (N4244, N4239, N3459, N3965, N961);
or OR3 (N4245, N4234, N4232, N2082);
buf BUF1 (N4246, N4210);
and AND3 (N4247, N4213, N1593, N4182);
not NOT1 (N4248, N4236);
nor NOR3 (N4249, N4245, N1403, N2311);
buf BUF1 (N4250, N4243);
not NOT1 (N4251, N4247);
nand NAND3 (N4252, N4249, N510, N3935);
nor NOR2 (N4253, N4237, N3131);
buf BUF1 (N4254, N4253);
buf BUF1 (N4255, N4240);
not NOT1 (N4256, N4242);
nand NAND3 (N4257, N4246, N2899, N3922);
nand NAND4 (N4258, N4248, N355, N4197, N106);
nor NOR3 (N4259, N4241, N2657, N2850);
and AND3 (N4260, N4256, N2871, N2015);
or OR4 (N4261, N4244, N3469, N2327, N1001);
and AND3 (N4262, N4260, N868, N2277);
nand NAND4 (N4263, N4261, N1265, N3094, N3218);
or OR2 (N4264, N4258, N3250);
or OR3 (N4265, N4254, N3004, N707);
nand NAND3 (N4266, N4251, N2872, N3747);
not NOT1 (N4267, N4265);
nor NOR3 (N4268, N4250, N1602, N3178);
buf BUF1 (N4269, N4252);
or OR3 (N4270, N4268, N1642, N2597);
xor XOR2 (N4271, N4259, N600);
nand NAND2 (N4272, N4264, N4073);
or OR2 (N4273, N4262, N3505);
not NOT1 (N4274, N4263);
buf BUF1 (N4275, N4274);
xor XOR2 (N4276, N4257, N1414);
xor XOR2 (N4277, N4272, N1525);
xor XOR2 (N4278, N4277, N525);
or OR4 (N4279, N4270, N678, N1252, N2349);
nand NAND2 (N4280, N4278, N2267);
or OR4 (N4281, N4280, N1148, N4251, N1903);
and AND2 (N4282, N4255, N4045);
and AND3 (N4283, N4267, N1874, N4057);
buf BUF1 (N4284, N4266);
nand NAND3 (N4285, N4282, N4238, N244);
nand NAND4 (N4286, N4285, N3987, N4005, N892);
not NOT1 (N4287, N4281);
xor XOR2 (N4288, N4271, N1390);
and AND2 (N4289, N4283, N362);
and AND3 (N4290, N4276, N137, N478);
xor XOR2 (N4291, N4288, N2310);
not NOT1 (N4292, N4275);
nor NOR4 (N4293, N4269, N2580, N1822, N702);
xor XOR2 (N4294, N4286, N3664);
not NOT1 (N4295, N4289);
and AND3 (N4296, N4292, N2255, N1061);
xor XOR2 (N4297, N4296, N1881);
xor XOR2 (N4298, N4287, N1926);
xor XOR2 (N4299, N4290, N500);
nand NAND2 (N4300, N4279, N3763);
xor XOR2 (N4301, N4291, N4076);
not NOT1 (N4302, N4297);
buf BUF1 (N4303, N4301);
nor NOR3 (N4304, N4300, N1016, N1178);
or OR4 (N4305, N4298, N3867, N3076, N2704);
xor XOR2 (N4306, N4284, N3371);
not NOT1 (N4307, N4306);
nor NOR2 (N4308, N4307, N210);
xor XOR2 (N4309, N4308, N1961);
buf BUF1 (N4310, N4294);
not NOT1 (N4311, N4299);
nand NAND3 (N4312, N4303, N999, N1291);
not NOT1 (N4313, N4304);
or OR4 (N4314, N4302, N3838, N1135, N2469);
xor XOR2 (N4315, N4311, N2047);
or OR3 (N4316, N4309, N2663, N483);
or OR2 (N4317, N4310, N2402);
xor XOR2 (N4318, N4293, N482);
or OR3 (N4319, N4317, N2687, N3741);
and AND3 (N4320, N4316, N1376, N4091);
or OR4 (N4321, N4318, N3702, N4233, N3893);
nand NAND3 (N4322, N4313, N3083, N3853);
nor NOR3 (N4323, N4295, N3512, N3402);
buf BUF1 (N4324, N4322);
not NOT1 (N4325, N4324);
buf BUF1 (N4326, N4305);
nand NAND4 (N4327, N4273, N1360, N1970, N2439);
or OR2 (N4328, N4326, N3343);
nand NAND2 (N4329, N4320, N2367);
buf BUF1 (N4330, N4315);
not NOT1 (N4331, N4323);
nor NOR4 (N4332, N4312, N2972, N3625, N1136);
xor XOR2 (N4333, N4332, N4074);
nand NAND3 (N4334, N4330, N1268, N20);
nand NAND2 (N4335, N4331, N3982);
or OR3 (N4336, N4329, N1353, N3138);
nand NAND3 (N4337, N4314, N3539, N3319);
or OR4 (N4338, N4336, N1763, N3853, N1825);
and AND4 (N4339, N4338, N189, N448, N4265);
not NOT1 (N4340, N4328);
or OR3 (N4341, N4319, N799, N4297);
or OR3 (N4342, N4339, N2816, N2179);
nand NAND4 (N4343, N4334, N3906, N3384, N3196);
and AND3 (N4344, N4327, N2537, N3419);
nor NOR3 (N4345, N4335, N221, N1381);
not NOT1 (N4346, N4343);
and AND4 (N4347, N4342, N3661, N4145, N2558);
buf BUF1 (N4348, N4346);
nor NOR2 (N4349, N4325, N2654);
or OR2 (N4350, N4345, N4005);
nor NOR2 (N4351, N4340, N1653);
or OR2 (N4352, N4337, N3816);
or OR4 (N4353, N4352, N977, N84, N109);
and AND2 (N4354, N4351, N1458);
nand NAND3 (N4355, N4333, N2007, N405);
and AND2 (N4356, N4341, N1927);
nor NOR3 (N4357, N4353, N3943, N4186);
nand NAND3 (N4358, N4356, N3778, N104);
and AND2 (N4359, N4358, N3548);
buf BUF1 (N4360, N4349);
nor NOR2 (N4361, N4348, N3320);
buf BUF1 (N4362, N4361);
not NOT1 (N4363, N4360);
nor NOR3 (N4364, N4321, N892, N475);
nand NAND4 (N4365, N4362, N3223, N325, N969);
and AND2 (N4366, N4347, N1544);
nor NOR4 (N4367, N4366, N1969, N3004, N2876);
xor XOR2 (N4368, N4350, N1611);
nand NAND3 (N4369, N4357, N101, N4329);
xor XOR2 (N4370, N4363, N1948);
buf BUF1 (N4371, N4359);
buf BUF1 (N4372, N4367);
buf BUF1 (N4373, N4364);
not NOT1 (N4374, N4370);
or OR2 (N4375, N4365, N3421);
and AND3 (N4376, N4369, N1227, N374);
buf BUF1 (N4377, N4374);
buf BUF1 (N4378, N4371);
or OR2 (N4379, N4355, N2028);
buf BUF1 (N4380, N4377);
and AND3 (N4381, N4376, N199, N973);
nand NAND2 (N4382, N4381, N2871);
xor XOR2 (N4383, N4373, N215);
and AND3 (N4384, N4379, N3011, N1966);
or OR4 (N4385, N4354, N3244, N3901, N2942);
buf BUF1 (N4386, N4383);
xor XOR2 (N4387, N4385, N2083);
not NOT1 (N4388, N4368);
xor XOR2 (N4389, N4387, N236);
xor XOR2 (N4390, N4382, N2154);
nor NOR4 (N4391, N4386, N2547, N3318, N987);
xor XOR2 (N4392, N4390, N3651);
and AND2 (N4393, N4392, N2972);
or OR3 (N4394, N4393, N1012, N2504);
and AND4 (N4395, N4372, N791, N1230, N917);
or OR3 (N4396, N4378, N1712, N1385);
nor NOR2 (N4397, N4394, N1185);
not NOT1 (N4398, N4388);
nand NAND2 (N4399, N4391, N2131);
and AND3 (N4400, N4384, N2162, N2173);
or OR3 (N4401, N4397, N2463, N1176);
nor NOR3 (N4402, N4389, N844, N1848);
xor XOR2 (N4403, N4402, N3706);
or OR2 (N4404, N4399, N444);
nor NOR3 (N4405, N4401, N3568, N2559);
or OR3 (N4406, N4405, N821, N1576);
buf BUF1 (N4407, N4403);
and AND2 (N4408, N4375, N3144);
nand NAND3 (N4409, N4404, N1162, N3610);
xor XOR2 (N4410, N4407, N611);
not NOT1 (N4411, N4409);
nor NOR3 (N4412, N4380, N3949, N3219);
or OR3 (N4413, N4406, N1261, N423);
or OR2 (N4414, N4396, N3123);
and AND4 (N4415, N4412, N2751, N1264, N2058);
xor XOR2 (N4416, N4344, N2052);
nor NOR3 (N4417, N4411, N2512, N957);
xor XOR2 (N4418, N4410, N4403);
not NOT1 (N4419, N4400);
and AND3 (N4420, N4415, N710, N646);
and AND4 (N4421, N4413, N1996, N3458, N2514);
nor NOR3 (N4422, N4416, N1479, N440);
nand NAND3 (N4423, N4420, N2970, N1729);
nor NOR3 (N4424, N4398, N3759, N1184);
nor NOR2 (N4425, N4421, N3271);
not NOT1 (N4426, N4414);
and AND2 (N4427, N4423, N306);
not NOT1 (N4428, N4419);
nor NOR2 (N4429, N4424, N981);
and AND4 (N4430, N4418, N129, N2310, N4056);
and AND4 (N4431, N4425, N4261, N799, N2461);
or OR3 (N4432, N4429, N826, N384);
nor NOR4 (N4433, N4422, N2125, N1827, N3094);
nor NOR3 (N4434, N4432, N824, N3632);
and AND4 (N4435, N4434, N1362, N4198, N1655);
buf BUF1 (N4436, N4408);
nor NOR4 (N4437, N4395, N3440, N1537, N4132);
buf BUF1 (N4438, N4431);
and AND3 (N4439, N4438, N2294, N1353);
nand NAND4 (N4440, N4427, N3784, N3691, N4347);
buf BUF1 (N4441, N4436);
and AND2 (N4442, N4435, N1726);
not NOT1 (N4443, N4441);
nor NOR2 (N4444, N4439, N3070);
not NOT1 (N4445, N4417);
buf BUF1 (N4446, N4443);
nor NOR3 (N4447, N4444, N1971, N3173);
buf BUF1 (N4448, N4440);
and AND2 (N4449, N4437, N4389);
nand NAND2 (N4450, N4448, N4445);
nand NAND4 (N4451, N4355, N2743, N3152, N157);
and AND2 (N4452, N4447, N1370);
or OR3 (N4453, N4450, N315, N1291);
nand NAND4 (N4454, N4426, N1983, N4017, N3194);
not NOT1 (N4455, N4433);
nand NAND4 (N4456, N4430, N2751, N3889, N150);
not NOT1 (N4457, N4451);
not NOT1 (N4458, N4456);
xor XOR2 (N4459, N4454, N2478);
or OR4 (N4460, N4459, N4050, N2596, N4326);
or OR3 (N4461, N4458, N312, N1383);
or OR4 (N4462, N4460, N1859, N4391, N2774);
and AND3 (N4463, N4452, N2314, N3860);
not NOT1 (N4464, N4442);
buf BUF1 (N4465, N4449);
nor NOR4 (N4466, N4428, N3353, N3725, N2594);
not NOT1 (N4467, N4446);
buf BUF1 (N4468, N4455);
xor XOR2 (N4469, N4465, N2994);
and AND3 (N4470, N4453, N1355, N140);
and AND4 (N4471, N4470, N2627, N2642, N1143);
and AND2 (N4472, N4466, N2219);
xor XOR2 (N4473, N4468, N2283);
xor XOR2 (N4474, N4462, N2712);
and AND3 (N4475, N4461, N2966, N2388);
nand NAND3 (N4476, N4469, N2202, N3161);
buf BUF1 (N4477, N4457);
xor XOR2 (N4478, N4475, N3625);
or OR3 (N4479, N4477, N1842, N587);
and AND4 (N4480, N4476, N2267, N4412, N2244);
or OR2 (N4481, N4471, N1050);
not NOT1 (N4482, N4474);
nand NAND3 (N4483, N4480, N897, N978);
or OR4 (N4484, N4478, N2487, N542, N1330);
nor NOR4 (N4485, N4482, N3935, N513, N3971);
nor NOR3 (N4486, N4463, N23, N277);
xor XOR2 (N4487, N4485, N4133);
or OR3 (N4488, N4486, N76, N2226);
and AND2 (N4489, N4479, N2863);
nand NAND3 (N4490, N4487, N2913, N4284);
and AND3 (N4491, N4484, N4263, N592);
xor XOR2 (N4492, N4489, N1886);
nor NOR4 (N4493, N4473, N274, N3885, N3395);
buf BUF1 (N4494, N4490);
and AND3 (N4495, N4472, N819, N1640);
buf BUF1 (N4496, N4483);
and AND4 (N4497, N4488, N678, N3180, N2143);
xor XOR2 (N4498, N4492, N3509);
or OR4 (N4499, N4464, N166, N3526, N1695);
xor XOR2 (N4500, N4495, N4268);
nand NAND3 (N4501, N4481, N1746, N3900);
nand NAND4 (N4502, N4500, N154, N375, N4430);
nand NAND2 (N4503, N4496, N279);
and AND2 (N4504, N4502, N919);
or OR4 (N4505, N4499, N1885, N2229, N856);
xor XOR2 (N4506, N4504, N513);
nor NOR2 (N4507, N4505, N3492);
or OR3 (N4508, N4506, N3356, N3165);
or OR4 (N4509, N4467, N2390, N4231, N2484);
buf BUF1 (N4510, N4498);
nor NOR2 (N4511, N4507, N1740);
nor NOR3 (N4512, N4511, N3364, N346);
nand NAND2 (N4513, N4501, N2623);
and AND4 (N4514, N4503, N1586, N506, N1020);
xor XOR2 (N4515, N4491, N1379);
nand NAND3 (N4516, N4497, N4064, N4079);
buf BUF1 (N4517, N4515);
buf BUF1 (N4518, N4493);
and AND3 (N4519, N4517, N2915, N3251);
or OR3 (N4520, N4519, N269, N260);
nand NAND4 (N4521, N4516, N2404, N4498, N2922);
and AND2 (N4522, N4513, N1682);
or OR4 (N4523, N4509, N105, N2231, N4396);
xor XOR2 (N4524, N4494, N137);
xor XOR2 (N4525, N4523, N3181);
and AND2 (N4526, N4521, N1955);
nand NAND3 (N4527, N4514, N2093, N1789);
or OR2 (N4528, N4518, N2424);
buf BUF1 (N4529, N4510);
nor NOR3 (N4530, N4526, N2630, N104);
nor NOR2 (N4531, N4512, N2899);
nand NAND3 (N4532, N4520, N1525, N2583);
xor XOR2 (N4533, N4531, N1714);
nor NOR3 (N4534, N4525, N4108, N1992);
not NOT1 (N4535, N4508);
nor NOR4 (N4536, N4528, N3749, N1649, N1524);
buf BUF1 (N4537, N4524);
xor XOR2 (N4538, N4529, N1315);
buf BUF1 (N4539, N4535);
nand NAND2 (N4540, N4536, N3874);
not NOT1 (N4541, N4532);
nor NOR4 (N4542, N4540, N2317, N3551, N3910);
nor NOR4 (N4543, N4533, N2745, N1329, N3480);
buf BUF1 (N4544, N4543);
and AND2 (N4545, N4542, N4360);
or OR4 (N4546, N4522, N3198, N1529, N3868);
nor NOR3 (N4547, N4545, N1126, N2793);
and AND4 (N4548, N4544, N2394, N3005, N3200);
buf BUF1 (N4549, N4548);
not NOT1 (N4550, N4530);
nor NOR4 (N4551, N4550, N1337, N1902, N4076);
xor XOR2 (N4552, N4541, N3945);
nand NAND4 (N4553, N4549, N1559, N3858, N178);
nand NAND4 (N4554, N4537, N4324, N1810, N3088);
xor XOR2 (N4555, N4538, N299);
nand NAND2 (N4556, N4555, N2424);
not NOT1 (N4557, N4534);
buf BUF1 (N4558, N4527);
and AND2 (N4559, N4554, N4000);
nand NAND2 (N4560, N4552, N4357);
not NOT1 (N4561, N4551);
not NOT1 (N4562, N4547);
xor XOR2 (N4563, N4562, N3788);
buf BUF1 (N4564, N4539);
xor XOR2 (N4565, N4560, N4185);
not NOT1 (N4566, N4563);
xor XOR2 (N4567, N4561, N1996);
and AND2 (N4568, N4567, N997);
not NOT1 (N4569, N4558);
not NOT1 (N4570, N4569);
nor NOR4 (N4571, N4559, N2471, N3283, N856);
not NOT1 (N4572, N4570);
buf BUF1 (N4573, N4568);
buf BUF1 (N4574, N4573);
not NOT1 (N4575, N4557);
nor NOR3 (N4576, N4546, N4220, N3623);
not NOT1 (N4577, N4576);
nor NOR4 (N4578, N4577, N4344, N3432, N36);
xor XOR2 (N4579, N4564, N1331);
nor NOR4 (N4580, N4566, N1735, N2714, N1112);
or OR2 (N4581, N4574, N2202);
buf BUF1 (N4582, N4575);
xor XOR2 (N4583, N4571, N671);
and AND2 (N4584, N4556, N3583);
xor XOR2 (N4585, N4580, N2579);
or OR2 (N4586, N4579, N2390);
and AND4 (N4587, N4584, N99, N4418, N193);
buf BUF1 (N4588, N4583);
nor NOR4 (N4589, N4588, N3357, N1500, N1566);
buf BUF1 (N4590, N4587);
xor XOR2 (N4591, N4553, N94);
and AND4 (N4592, N4578, N2000, N3049, N2025);
and AND3 (N4593, N4585, N2554, N1287);
not NOT1 (N4594, N4586);
buf BUF1 (N4595, N4590);
or OR2 (N4596, N4592, N1581);
buf BUF1 (N4597, N4595);
nor NOR2 (N4598, N4589, N673);
not NOT1 (N4599, N4594);
buf BUF1 (N4600, N4596);
nand NAND4 (N4601, N4591, N3052, N3701, N3780);
or OR4 (N4602, N4593, N1837, N3584, N3005);
xor XOR2 (N4603, N4602, N181);
or OR3 (N4604, N4597, N644, N3134);
or OR3 (N4605, N4581, N3153, N2769);
buf BUF1 (N4606, N4582);
nor NOR4 (N4607, N4572, N933, N2626, N1856);
buf BUF1 (N4608, N4607);
buf BUF1 (N4609, N4604);
and AND2 (N4610, N4565, N1445);
nor NOR4 (N4611, N4603, N4113, N239, N2589);
nor NOR2 (N4612, N4605, N4220);
nand NAND4 (N4613, N4612, N3065, N4437, N3390);
buf BUF1 (N4614, N4600);
buf BUF1 (N4615, N4614);
or OR2 (N4616, N4615, N4154);
or OR2 (N4617, N4611, N2238);
nand NAND2 (N4618, N4613, N42);
xor XOR2 (N4619, N4617, N3003);
nor NOR4 (N4620, N4618, N3552, N4534, N1091);
or OR2 (N4621, N4619, N1848);
xor XOR2 (N4622, N4621, N96);
buf BUF1 (N4623, N4598);
nor NOR3 (N4624, N4623, N1207, N1453);
or OR4 (N4625, N4624, N3537, N2584, N2025);
and AND3 (N4626, N4625, N3317, N4443);
or OR2 (N4627, N4599, N4224);
xor XOR2 (N4628, N4610, N1611);
and AND3 (N4629, N4608, N1599, N2248);
nor NOR2 (N4630, N4616, N1283);
nor NOR2 (N4631, N4627, N1775);
xor XOR2 (N4632, N4631, N2001);
nor NOR3 (N4633, N4622, N3807, N1888);
or OR2 (N4634, N4630, N3194);
or OR4 (N4635, N4633, N483, N1126, N2644);
and AND2 (N4636, N4628, N484);
buf BUF1 (N4637, N4629);
nand NAND2 (N4638, N4609, N2638);
not NOT1 (N4639, N4606);
and AND4 (N4640, N4639, N3603, N346, N3896);
buf BUF1 (N4641, N4632);
and AND2 (N4642, N4641, N164);
xor XOR2 (N4643, N4637, N2196);
buf BUF1 (N4644, N4636);
xor XOR2 (N4645, N4642, N3260);
nor NOR4 (N4646, N4638, N3250, N1101, N1876);
not NOT1 (N4647, N4645);
not NOT1 (N4648, N4634);
and AND2 (N4649, N4648, N2473);
nor NOR3 (N4650, N4620, N1722, N2056);
xor XOR2 (N4651, N4635, N481);
nor NOR2 (N4652, N4649, N3278);
and AND3 (N4653, N4651, N1024, N2733);
or OR3 (N4654, N4646, N4591, N1156);
nor NOR2 (N4655, N4601, N3598);
or OR2 (N4656, N4652, N3354);
or OR3 (N4657, N4643, N1472, N2706);
xor XOR2 (N4658, N4654, N2150);
not NOT1 (N4659, N4644);
buf BUF1 (N4660, N4626);
or OR2 (N4661, N4658, N4553);
nand NAND4 (N4662, N4655, N1161, N3915, N2531);
or OR4 (N4663, N4647, N2304, N1506, N4556);
xor XOR2 (N4664, N4640, N2298);
xor XOR2 (N4665, N4659, N1785);
nand NAND3 (N4666, N4650, N1539, N2002);
or OR4 (N4667, N4666, N2818, N27, N1544);
not NOT1 (N4668, N4662);
not NOT1 (N4669, N4663);
and AND3 (N4670, N4660, N2800, N3161);
buf BUF1 (N4671, N4668);
buf BUF1 (N4672, N4664);
xor XOR2 (N4673, N4667, N3335);
not NOT1 (N4674, N4671);
and AND4 (N4675, N4665, N478, N1854, N1983);
not NOT1 (N4676, N4669);
nor NOR3 (N4677, N4653, N2445, N4572);
not NOT1 (N4678, N4672);
not NOT1 (N4679, N4677);
buf BUF1 (N4680, N4661);
xor XOR2 (N4681, N4656, N401);
and AND2 (N4682, N4670, N4355);
and AND4 (N4683, N4675, N1498, N950, N1055);
nand NAND4 (N4684, N4673, N253, N520, N1224);
buf BUF1 (N4685, N4679);
buf BUF1 (N4686, N4684);
and AND3 (N4687, N4683, N1867, N1895);
buf BUF1 (N4688, N4678);
nand NAND3 (N4689, N4687, N3123, N12);
and AND2 (N4690, N4686, N3240);
not NOT1 (N4691, N4681);
nand NAND4 (N4692, N4689, N4320, N2839, N3832);
not NOT1 (N4693, N4680);
buf BUF1 (N4694, N4690);
or OR4 (N4695, N4691, N784, N4618, N1071);
and AND2 (N4696, N4695, N108);
and AND2 (N4697, N4685, N3827);
and AND4 (N4698, N4694, N1203, N171, N1461);
xor XOR2 (N4699, N4692, N3177);
not NOT1 (N4700, N4698);
nand NAND3 (N4701, N4657, N2542, N3888);
and AND3 (N4702, N4676, N1835, N3835);
nand NAND4 (N4703, N4688, N2058, N778, N1280);
or OR4 (N4704, N4674, N2918, N4529, N1208);
xor XOR2 (N4705, N4700, N2426);
nor NOR3 (N4706, N4693, N4463, N1113);
nor NOR4 (N4707, N4702, N4450, N1099, N4105);
not NOT1 (N4708, N4703);
nand NAND4 (N4709, N4696, N1005, N4699, N3299);
nand NAND4 (N4710, N2253, N2058, N4180, N468);
nand NAND2 (N4711, N4710, N2709);
nand NAND4 (N4712, N4708, N3020, N1341, N1125);
not NOT1 (N4713, N4709);
and AND4 (N4714, N4705, N1133, N1985, N731);
nand NAND4 (N4715, N4714, N410, N1166, N2650);
nand NAND2 (N4716, N4711, N3685);
not NOT1 (N4717, N4682);
and AND3 (N4718, N4707, N4330, N2628);
nor NOR2 (N4719, N4701, N2294);
nor NOR2 (N4720, N4704, N2071);
nor NOR4 (N4721, N4719, N528, N574, N434);
or OR3 (N4722, N4720, N2650, N1989);
buf BUF1 (N4723, N4713);
nand NAND3 (N4724, N4716, N4535, N2065);
nor NOR3 (N4725, N4721, N2293, N2198);
and AND3 (N4726, N4725, N2346, N2775);
buf BUF1 (N4727, N4715);
nor NOR2 (N4728, N4722, N2652);
and AND3 (N4729, N4723, N3709, N2310);
not NOT1 (N4730, N4728);
nor NOR4 (N4731, N4727, N592, N7, N2842);
buf BUF1 (N4732, N4726);
xor XOR2 (N4733, N4732, N4357);
or OR3 (N4734, N4730, N1625, N1703);
xor XOR2 (N4735, N4712, N4713);
and AND4 (N4736, N4718, N3160, N1278, N3125);
nor NOR2 (N4737, N4736, N3629);
xor XOR2 (N4738, N4737, N508);
and AND3 (N4739, N4735, N3119, N3164);
buf BUF1 (N4740, N4706);
not NOT1 (N4741, N4724);
not NOT1 (N4742, N4733);
xor XOR2 (N4743, N4738, N1771);
or OR3 (N4744, N4742, N311, N1917);
and AND2 (N4745, N4731, N3314);
or OR3 (N4746, N4697, N2432, N2204);
xor XOR2 (N4747, N4739, N448);
buf BUF1 (N4748, N4743);
nor NOR3 (N4749, N4746, N2668, N1235);
buf BUF1 (N4750, N4749);
xor XOR2 (N4751, N4717, N24);
xor XOR2 (N4752, N4750, N1345);
buf BUF1 (N4753, N4745);
xor XOR2 (N4754, N4741, N977);
nor NOR3 (N4755, N4754, N3377, N3401);
or OR3 (N4756, N4744, N2047, N2651);
buf BUF1 (N4757, N4753);
xor XOR2 (N4758, N4752, N3328);
xor XOR2 (N4759, N4757, N1648);
buf BUF1 (N4760, N4748);
not NOT1 (N4761, N4760);
nand NAND3 (N4762, N4729, N3424, N1651);
nor NOR3 (N4763, N4756, N2242, N1547);
nor NOR2 (N4764, N4747, N1344);
not NOT1 (N4765, N4761);
nor NOR3 (N4766, N4755, N4653, N1444);
buf BUF1 (N4767, N4764);
buf BUF1 (N4768, N4758);
or OR4 (N4769, N4768, N119, N2776, N262);
buf BUF1 (N4770, N4765);
nor NOR3 (N4771, N4734, N252, N1);
nor NOR4 (N4772, N4740, N2788, N2184, N800);
buf BUF1 (N4773, N4767);
or OR4 (N4774, N4773, N3326, N959, N4109);
not NOT1 (N4775, N4772);
nand NAND3 (N4776, N4774, N522, N331);
buf BUF1 (N4777, N4762);
or OR2 (N4778, N4763, N2793);
not NOT1 (N4779, N4759);
buf BUF1 (N4780, N4770);
and AND4 (N4781, N4771, N1462, N727, N1923);
xor XOR2 (N4782, N4751, N3768);
nand NAND3 (N4783, N4769, N3741, N3209);
not NOT1 (N4784, N4777);
and AND4 (N4785, N4779, N220, N3953, N293);
buf BUF1 (N4786, N4782);
xor XOR2 (N4787, N4776, N462);
nand NAND3 (N4788, N4786, N2294, N769);
nand NAND3 (N4789, N4785, N662, N433);
xor XOR2 (N4790, N4775, N830);
and AND3 (N4791, N4781, N3135, N3083);
nand NAND3 (N4792, N4780, N2859, N3874);
and AND4 (N4793, N4778, N4617, N3031, N1089);
and AND3 (N4794, N4789, N4122, N2312);
xor XOR2 (N4795, N4792, N4304);
and AND4 (N4796, N4795, N1276, N4509, N3473);
nor NOR2 (N4797, N4766, N1718);
xor XOR2 (N4798, N4787, N4281);
and AND2 (N4799, N4798, N3438);
xor XOR2 (N4800, N4790, N2059);
buf BUF1 (N4801, N4796);
or OR2 (N4802, N4793, N4018);
nand NAND3 (N4803, N4788, N442, N3110);
not NOT1 (N4804, N4784);
buf BUF1 (N4805, N4783);
and AND4 (N4806, N4800, N3000, N697, N3942);
xor XOR2 (N4807, N4794, N4451);
or OR2 (N4808, N4802, N4462);
nor NOR3 (N4809, N4807, N1371, N4359);
buf BUF1 (N4810, N4801);
buf BUF1 (N4811, N4797);
buf BUF1 (N4812, N4791);
nand NAND3 (N4813, N4809, N1729, N2879);
or OR3 (N4814, N4806, N2463, N1231);
buf BUF1 (N4815, N4812);
nor NOR2 (N4816, N4813, N4325);
buf BUF1 (N4817, N4814);
or OR2 (N4818, N4815, N625);
buf BUF1 (N4819, N4799);
buf BUF1 (N4820, N4804);
buf BUF1 (N4821, N4803);
nand NAND2 (N4822, N4805, N4481);
not NOT1 (N4823, N4821);
nand NAND3 (N4824, N4822, N3399, N2499);
and AND2 (N4825, N4817, N3961);
nand NAND3 (N4826, N4819, N3323, N3914);
nand NAND2 (N4827, N4823, N2660);
buf BUF1 (N4828, N4825);
and AND3 (N4829, N4826, N1908, N3563);
nor NOR3 (N4830, N4811, N1899, N4019);
xor XOR2 (N4831, N4829, N4251);
nor NOR4 (N4832, N4828, N4757, N940, N124);
xor XOR2 (N4833, N4827, N2916);
or OR2 (N4834, N4816, N784);
or OR2 (N4835, N4833, N1531);
nor NOR4 (N4836, N4831, N1270, N4738, N2056);
not NOT1 (N4837, N4836);
nand NAND2 (N4838, N4810, N2335);
buf BUF1 (N4839, N4808);
and AND2 (N4840, N4832, N942);
nand NAND2 (N4841, N4837, N1976);
nor NOR3 (N4842, N4840, N4746, N504);
or OR4 (N4843, N4839, N1772, N1408, N3301);
nand NAND2 (N4844, N4843, N430);
not NOT1 (N4845, N4842);
buf BUF1 (N4846, N4844);
or OR2 (N4847, N4818, N1878);
buf BUF1 (N4848, N4835);
xor XOR2 (N4849, N4848, N1787);
nand NAND2 (N4850, N4824, N4474);
not NOT1 (N4851, N4838);
and AND4 (N4852, N4845, N3502, N3697, N673);
xor XOR2 (N4853, N4850, N1464);
xor XOR2 (N4854, N4846, N210);
buf BUF1 (N4855, N4852);
not NOT1 (N4856, N4834);
xor XOR2 (N4857, N4849, N475);
or OR2 (N4858, N4841, N3316);
xor XOR2 (N4859, N4830, N2429);
buf BUF1 (N4860, N4854);
buf BUF1 (N4861, N4859);
not NOT1 (N4862, N4851);
not NOT1 (N4863, N4857);
nand NAND2 (N4864, N4862, N3169);
and AND3 (N4865, N4856, N2682, N4589);
and AND4 (N4866, N4865, N2597, N140, N1304);
xor XOR2 (N4867, N4864, N3227);
and AND2 (N4868, N4861, N816);
and AND3 (N4869, N4853, N2405, N1206);
and AND3 (N4870, N4855, N2498, N1191);
not NOT1 (N4871, N4870);
nor NOR3 (N4872, N4863, N2535, N997);
nand NAND2 (N4873, N4866, N2455);
buf BUF1 (N4874, N4869);
xor XOR2 (N4875, N4871, N2559);
and AND3 (N4876, N4872, N2666, N476);
buf BUF1 (N4877, N4876);
not NOT1 (N4878, N4875);
and AND3 (N4879, N4858, N4845, N720);
xor XOR2 (N4880, N4868, N3114);
nor NOR4 (N4881, N4879, N4675, N4133, N3095);
and AND2 (N4882, N4878, N1490);
not NOT1 (N4883, N4877);
buf BUF1 (N4884, N4881);
buf BUF1 (N4885, N4883);
nand NAND4 (N4886, N4880, N740, N2171, N678);
xor XOR2 (N4887, N4867, N1186);
not NOT1 (N4888, N4847);
and AND4 (N4889, N4888, N3372, N561, N3911);
or OR2 (N4890, N4860, N4762);
and AND4 (N4891, N4873, N2302, N322, N1213);
and AND3 (N4892, N4874, N3419, N225);
nand NAND3 (N4893, N4882, N1887, N3273);
nor NOR4 (N4894, N4820, N1739, N211, N15);
xor XOR2 (N4895, N4887, N786);
nand NAND2 (N4896, N4891, N2877);
and AND4 (N4897, N4892, N679, N2062, N1861);
nor NOR2 (N4898, N4886, N1227);
and AND2 (N4899, N4895, N4136);
nand NAND3 (N4900, N4897, N4071, N3086);
buf BUF1 (N4901, N4899);
nand NAND2 (N4902, N4900, N4770);
or OR2 (N4903, N4889, N612);
nor NOR2 (N4904, N4890, N411);
and AND4 (N4905, N4904, N3333, N2260, N2825);
buf BUF1 (N4906, N4885);
xor XOR2 (N4907, N4903, N2897);
nand NAND3 (N4908, N4898, N4536, N4640);
buf BUF1 (N4909, N4901);
buf BUF1 (N4910, N4896);
xor XOR2 (N4911, N4910, N1808);
and AND4 (N4912, N4906, N4259, N1708, N329);
xor XOR2 (N4913, N4907, N947);
nand NAND4 (N4914, N4912, N2603, N2060, N676);
nand NAND4 (N4915, N4905, N4880, N3497, N4861);
xor XOR2 (N4916, N4909, N3453);
xor XOR2 (N4917, N4908, N1778);
nand NAND4 (N4918, N4884, N4057, N1759, N1022);
xor XOR2 (N4919, N4914, N4435);
xor XOR2 (N4920, N4918, N1913);
buf BUF1 (N4921, N4911);
not NOT1 (N4922, N4915);
not NOT1 (N4923, N4921);
or OR2 (N4924, N4894, N359);
and AND2 (N4925, N4919, N4314);
xor XOR2 (N4926, N4923, N2075);
xor XOR2 (N4927, N4893, N586);
or OR4 (N4928, N4925, N4059, N350, N3496);
not NOT1 (N4929, N4927);
or OR2 (N4930, N4917, N4141);
nand NAND2 (N4931, N4920, N2179);
nor NOR2 (N4932, N4922, N3759);
and AND2 (N4933, N4929, N808);
xor XOR2 (N4934, N4913, N2323);
not NOT1 (N4935, N4934);
and AND2 (N4936, N4933, N4574);
or OR3 (N4937, N4935, N687, N3948);
nor NOR2 (N4938, N4916, N3927);
not NOT1 (N4939, N4930);
xor XOR2 (N4940, N4939, N3889);
xor XOR2 (N4941, N4940, N4357);
and AND2 (N4942, N4938, N1736);
buf BUF1 (N4943, N4926);
nor NOR2 (N4944, N4928, N3976);
nand NAND2 (N4945, N4944, N162);
and AND3 (N4946, N4941, N545, N3963);
nor NOR2 (N4947, N4902, N3857);
nor NOR4 (N4948, N4932, N3076, N554, N3806);
nor NOR3 (N4949, N4943, N279, N2837);
not NOT1 (N4950, N4947);
not NOT1 (N4951, N4942);
and AND4 (N4952, N4945, N2361, N3943, N4369);
nor NOR2 (N4953, N4924, N1337);
or OR3 (N4954, N4936, N3632, N2117);
buf BUF1 (N4955, N4946);
nor NOR3 (N4956, N4953, N4691, N1545);
or OR4 (N4957, N4954, N463, N2896, N4361);
and AND4 (N4958, N4948, N476, N3207, N3925);
and AND2 (N4959, N4950, N169);
buf BUF1 (N4960, N4952);
nor NOR2 (N4961, N4951, N2221);
nand NAND4 (N4962, N4949, N4500, N3736, N4215);
nand NAND4 (N4963, N4931, N3907, N3381, N3115);
not NOT1 (N4964, N4963);
nand NAND4 (N4965, N4959, N2337, N3804, N3726);
nand NAND2 (N4966, N4937, N2753);
and AND2 (N4967, N4955, N375);
or OR4 (N4968, N4967, N188, N985, N2553);
xor XOR2 (N4969, N4965, N2126);
xor XOR2 (N4970, N4966, N577);
buf BUF1 (N4971, N4968);
not NOT1 (N4972, N4958);
and AND4 (N4973, N4960, N417, N918, N2425);
buf BUF1 (N4974, N4964);
buf BUF1 (N4975, N4961);
xor XOR2 (N4976, N4957, N1818);
buf BUF1 (N4977, N4975);
xor XOR2 (N4978, N4976, N4004);
and AND2 (N4979, N4970, N4358);
nor NOR3 (N4980, N4979, N2812, N3820);
xor XOR2 (N4981, N4972, N1233);
buf BUF1 (N4982, N4977);
buf BUF1 (N4983, N4971);
buf BUF1 (N4984, N4956);
nand NAND2 (N4985, N4982, N2987);
or OR2 (N4986, N4978, N356);
or OR4 (N4987, N4984, N487, N2753, N4621);
nor NOR4 (N4988, N4973, N4527, N1334, N3338);
and AND3 (N4989, N4981, N3336, N1927);
and AND2 (N4990, N4987, N276);
not NOT1 (N4991, N4980);
buf BUF1 (N4992, N4962);
xor XOR2 (N4993, N4974, N2036);
nand NAND2 (N4994, N4969, N4324);
and AND2 (N4995, N4993, N2903);
or OR3 (N4996, N4983, N1007, N729);
not NOT1 (N4997, N4990);
and AND2 (N4998, N4985, N3744);
nand NAND2 (N4999, N4986, N4090);
nor NOR3 (N5000, N4995, N1268, N1889);
not NOT1 (N5001, N4989);
and AND3 (N5002, N4996, N2525, N84);
xor XOR2 (N5003, N4991, N1813);
nand NAND4 (N5004, N5000, N3694, N781, N2425);
not NOT1 (N5005, N4994);
or OR3 (N5006, N5005, N4553, N1649);
not NOT1 (N5007, N4997);
xor XOR2 (N5008, N5007, N2568);
buf BUF1 (N5009, N5001);
nand NAND3 (N5010, N4992, N419, N3352);
not NOT1 (N5011, N5004);
nor NOR3 (N5012, N4998, N2491, N1625);
buf BUF1 (N5013, N5006);
nor NOR3 (N5014, N4988, N4175, N2878);
nand NAND4 (N5015, N4999, N3436, N2911, N1138);
nand NAND3 (N5016, N5002, N1196, N2058);
buf BUF1 (N5017, N5010);
nor NOR3 (N5018, N5013, N4339, N4351);
nand NAND2 (N5019, N5012, N472);
nand NAND4 (N5020, N5009, N3744, N550, N1097);
and AND3 (N5021, N5003, N4135, N1527);
nand NAND2 (N5022, N5011, N2826);
nand NAND4 (N5023, N5016, N4249, N1915, N1294);
not NOT1 (N5024, N5014);
nand NAND2 (N5025, N5015, N2355);
xor XOR2 (N5026, N5023, N2789);
buf BUF1 (N5027, N5020);
nand NAND4 (N5028, N5027, N3711, N4405, N4296);
nand NAND3 (N5029, N5022, N4128, N3442);
not NOT1 (N5030, N5028);
buf BUF1 (N5031, N5026);
nor NOR3 (N5032, N5031, N961, N1289);
nand NAND2 (N5033, N5024, N2240);
and AND4 (N5034, N5008, N1546, N3948, N3942);
not NOT1 (N5035, N5021);
or OR2 (N5036, N5025, N152);
buf BUF1 (N5037, N5032);
and AND2 (N5038, N5036, N2069);
and AND2 (N5039, N5017, N5003);
xor XOR2 (N5040, N5033, N3940);
nor NOR4 (N5041, N5037, N3344, N3814, N1272);
not NOT1 (N5042, N5034);
xor XOR2 (N5043, N5042, N452);
nor NOR4 (N5044, N5039, N3612, N2137, N3932);
or OR3 (N5045, N5019, N4416, N3265);
buf BUF1 (N5046, N5041);
and AND4 (N5047, N5043, N424, N3680, N2172);
buf BUF1 (N5048, N5044);
nor NOR4 (N5049, N5046, N4924, N1269, N4260);
xor XOR2 (N5050, N5035, N354);
nand NAND3 (N5051, N5018, N900, N381);
and AND3 (N5052, N5029, N3049, N3860);
buf BUF1 (N5053, N5045);
nor NOR4 (N5054, N5052, N3293, N4425, N3538);
nand NAND3 (N5055, N5047, N2536, N4546);
nand NAND3 (N5056, N5050, N4442, N3226);
and AND3 (N5057, N5054, N149, N557);
buf BUF1 (N5058, N5048);
not NOT1 (N5059, N5058);
nor NOR3 (N5060, N5030, N2799, N1043);
not NOT1 (N5061, N5049);
buf BUF1 (N5062, N5040);
and AND3 (N5063, N5053, N2288, N1026);
not NOT1 (N5064, N5063);
nor NOR4 (N5065, N5057, N3115, N1851, N4625);
nor NOR3 (N5066, N5056, N490, N2697);
buf BUF1 (N5067, N5038);
or OR4 (N5068, N5066, N2278, N229, N4127);
nor NOR3 (N5069, N5060, N42, N4798);
or OR3 (N5070, N5064, N2070, N2140);
nor NOR4 (N5071, N5070, N3751, N1219, N2571);
nand NAND3 (N5072, N5069, N1247, N373);
not NOT1 (N5073, N5065);
not NOT1 (N5074, N5068);
nand NAND2 (N5075, N5059, N3600);
xor XOR2 (N5076, N5071, N3098);
xor XOR2 (N5077, N5072, N764);
buf BUF1 (N5078, N5061);
and AND2 (N5079, N5055, N222);
xor XOR2 (N5080, N5079, N4267);
buf BUF1 (N5081, N5077);
buf BUF1 (N5082, N5076);
and AND3 (N5083, N5051, N4802, N2437);
nand NAND4 (N5084, N5062, N328, N3433, N114);
nor NOR4 (N5085, N5073, N4385, N3736, N2333);
and AND3 (N5086, N5078, N1739, N3984);
buf BUF1 (N5087, N5080);
nand NAND3 (N5088, N5087, N2190, N1659);
and AND3 (N5089, N5083, N1743, N2268);
and AND4 (N5090, N5084, N2422, N2578, N4970);
xor XOR2 (N5091, N5089, N3157);
buf BUF1 (N5092, N5075);
or OR4 (N5093, N5085, N4818, N728, N2404);
nand NAND4 (N5094, N5090, N1580, N808, N2562);
or OR4 (N5095, N5094, N4779, N1077, N177);
buf BUF1 (N5096, N5095);
xor XOR2 (N5097, N5096, N1040);
nor NOR2 (N5098, N5092, N2908);
nor NOR3 (N5099, N5093, N1854, N3884);
not NOT1 (N5100, N5097);
nand NAND2 (N5101, N5098, N4889);
nor NOR3 (N5102, N5086, N664, N2493);
buf BUF1 (N5103, N5101);
xor XOR2 (N5104, N5081, N2291);
or OR4 (N5105, N5100, N1774, N2915, N1977);
or OR2 (N5106, N5091, N3101);
xor XOR2 (N5107, N5067, N185);
xor XOR2 (N5108, N5099, N544);
or OR2 (N5109, N5074, N863);
nand NAND3 (N5110, N5108, N3560, N3416);
xor XOR2 (N5111, N5082, N4658);
not NOT1 (N5112, N5107);
nand NAND4 (N5113, N5111, N2963, N5044, N1939);
nand NAND2 (N5114, N5103, N3224);
xor XOR2 (N5115, N5109, N4691);
or OR3 (N5116, N5105, N361, N2876);
nand NAND3 (N5117, N5116, N1935, N821);
or OR3 (N5118, N5117, N4088, N2420);
xor XOR2 (N5119, N5114, N3341);
nand NAND4 (N5120, N5104, N212, N3367, N3988);
not NOT1 (N5121, N5088);
and AND2 (N5122, N5119, N2519);
not NOT1 (N5123, N5118);
or OR2 (N5124, N5112, N2793);
xor XOR2 (N5125, N5120, N526);
buf BUF1 (N5126, N5122);
not NOT1 (N5127, N5124);
not NOT1 (N5128, N5121);
or OR4 (N5129, N5128, N3949, N2438, N4445);
not NOT1 (N5130, N5106);
xor XOR2 (N5131, N5123, N4594);
nor NOR4 (N5132, N5131, N3580, N4258, N1821);
nand NAND3 (N5133, N5102, N1987, N2044);
buf BUF1 (N5134, N5133);
not NOT1 (N5135, N5134);
buf BUF1 (N5136, N5125);
or OR2 (N5137, N5130, N2277);
and AND2 (N5138, N5137, N755);
buf BUF1 (N5139, N5138);
not NOT1 (N5140, N5115);
not NOT1 (N5141, N5139);
buf BUF1 (N5142, N5136);
nand NAND4 (N5143, N5113, N767, N3571, N4831);
not NOT1 (N5144, N5140);
nand NAND4 (N5145, N5142, N497, N3594, N2966);
or OR2 (N5146, N5132, N2452);
nor NOR3 (N5147, N5127, N2170, N488);
nand NAND3 (N5148, N5146, N2687, N1893);
buf BUF1 (N5149, N5141);
and AND4 (N5150, N5149, N893, N3085, N3853);
buf BUF1 (N5151, N5144);
buf BUF1 (N5152, N5147);
and AND3 (N5153, N5150, N2070, N4774);
and AND4 (N5154, N5151, N5055, N4820, N416);
not NOT1 (N5155, N5129);
nand NAND2 (N5156, N5145, N713);
nor NOR4 (N5157, N5126, N3164, N3380, N4329);
xor XOR2 (N5158, N5153, N199);
xor XOR2 (N5159, N5156, N4226);
buf BUF1 (N5160, N5110);
nand NAND3 (N5161, N5135, N5150, N2084);
xor XOR2 (N5162, N5152, N739);
nand NAND3 (N5163, N5162, N948, N4488);
or OR4 (N5164, N5143, N4883, N252, N3578);
buf BUF1 (N5165, N5164);
buf BUF1 (N5166, N5154);
not NOT1 (N5167, N5166);
buf BUF1 (N5168, N5163);
not NOT1 (N5169, N5157);
buf BUF1 (N5170, N5158);
not NOT1 (N5171, N5160);
xor XOR2 (N5172, N5170, N3491);
buf BUF1 (N5173, N5161);
nor NOR3 (N5174, N5168, N2672, N1212);
not NOT1 (N5175, N5172);
and AND3 (N5176, N5171, N1631, N947);
xor XOR2 (N5177, N5169, N3481);
and AND2 (N5178, N5174, N4503);
not NOT1 (N5179, N5173);
nand NAND4 (N5180, N5165, N540, N3409, N3819);
nor NOR4 (N5181, N5155, N4641, N1249, N2160);
or OR2 (N5182, N5181, N4220);
or OR2 (N5183, N5159, N4703);
xor XOR2 (N5184, N5183, N4840);
nor NOR2 (N5185, N5179, N3627);
nand NAND4 (N5186, N5178, N3650, N3728, N1414);
and AND2 (N5187, N5186, N1192);
nand NAND3 (N5188, N5148, N784, N1286);
or OR2 (N5189, N5175, N2630);
nor NOR4 (N5190, N5182, N1472, N4643, N2156);
buf BUF1 (N5191, N5189);
nor NOR4 (N5192, N5167, N4498, N535, N564);
or OR3 (N5193, N5190, N4777, N108);
and AND2 (N5194, N5188, N3209);
buf BUF1 (N5195, N5180);
and AND2 (N5196, N5191, N2043);
buf BUF1 (N5197, N5185);
not NOT1 (N5198, N5176);
not NOT1 (N5199, N5184);
xor XOR2 (N5200, N5195, N3455);
or OR2 (N5201, N5194, N2121);
xor XOR2 (N5202, N5199, N3482);
or OR4 (N5203, N5177, N3712, N4364, N1708);
buf BUF1 (N5204, N5196);
xor XOR2 (N5205, N5201, N3539);
nor NOR2 (N5206, N5193, N4660);
not NOT1 (N5207, N5200);
and AND2 (N5208, N5207, N5020);
and AND4 (N5209, N5202, N529, N3369, N1885);
not NOT1 (N5210, N5204);
and AND4 (N5211, N5197, N570, N3705, N3127);
and AND2 (N5212, N5210, N2906);
or OR2 (N5213, N5205, N2168);
nand NAND3 (N5214, N5211, N812, N4464);
not NOT1 (N5215, N5192);
or OR2 (N5216, N5206, N357);
or OR4 (N5217, N5187, N467, N515, N179);
nand NAND4 (N5218, N5217, N4865, N787, N981);
not NOT1 (N5219, N5209);
xor XOR2 (N5220, N5203, N5107);
and AND3 (N5221, N5198, N5123, N4730);
and AND4 (N5222, N5219, N2779, N2092, N3574);
nor NOR3 (N5223, N5214, N4539, N3729);
not NOT1 (N5224, N5222);
nand NAND4 (N5225, N5220, N2916, N1286, N171);
nand NAND4 (N5226, N5225, N1629, N389, N4491);
nand NAND2 (N5227, N5208, N4996);
buf BUF1 (N5228, N5213);
nand NAND3 (N5229, N5212, N1561, N2290);
not NOT1 (N5230, N5228);
xor XOR2 (N5231, N5215, N2738);
not NOT1 (N5232, N5224);
nand NAND4 (N5233, N5227, N2742, N2511, N1568);
nand NAND2 (N5234, N5233, N138);
and AND4 (N5235, N5221, N720, N3799, N979);
nor NOR3 (N5236, N5229, N3478, N175);
and AND3 (N5237, N5226, N2879, N5091);
buf BUF1 (N5238, N5218);
xor XOR2 (N5239, N5216, N2307);
and AND3 (N5240, N5232, N158, N526);
not NOT1 (N5241, N5237);
xor XOR2 (N5242, N5238, N3487);
xor XOR2 (N5243, N5236, N3925);
buf BUF1 (N5244, N5234);
not NOT1 (N5245, N5241);
nor NOR3 (N5246, N5243, N3946, N2342);
not NOT1 (N5247, N5231);
nor NOR3 (N5248, N5230, N4689, N3352);
not NOT1 (N5249, N5246);
xor XOR2 (N5250, N5248, N485);
xor XOR2 (N5251, N5242, N987);
xor XOR2 (N5252, N5244, N2037);
and AND4 (N5253, N5251, N2278, N2253, N3727);
buf BUF1 (N5254, N5240);
and AND3 (N5255, N5245, N4816, N1386);
buf BUF1 (N5256, N5247);
and AND2 (N5257, N5252, N854);
or OR4 (N5258, N5249, N109, N4684, N1155);
xor XOR2 (N5259, N5253, N1567);
xor XOR2 (N5260, N5235, N3660);
and AND3 (N5261, N5250, N4365, N2498);
buf BUF1 (N5262, N5259);
and AND3 (N5263, N5262, N3396, N250);
or OR4 (N5264, N5258, N3286, N2543, N3232);
or OR3 (N5265, N5261, N1159, N1424);
nand NAND3 (N5266, N5239, N1026, N1968);
nor NOR3 (N5267, N5255, N3512, N848);
or OR4 (N5268, N5254, N3486, N791, N467);
nor NOR2 (N5269, N5264, N373);
or OR3 (N5270, N5266, N1577, N3508);
and AND3 (N5271, N5265, N406, N4818);
xor XOR2 (N5272, N5257, N1837);
or OR2 (N5273, N5263, N179);
nor NOR4 (N5274, N5271, N898, N3924, N181);
xor XOR2 (N5275, N5223, N4646);
xor XOR2 (N5276, N5267, N4826);
nor NOR3 (N5277, N5276, N1675, N870);
and AND4 (N5278, N5275, N2180, N2004, N4782);
and AND3 (N5279, N5272, N1809, N2582);
buf BUF1 (N5280, N5273);
buf BUF1 (N5281, N5270);
buf BUF1 (N5282, N5256);
not NOT1 (N5283, N5278);
buf BUF1 (N5284, N5283);
nor NOR4 (N5285, N5277, N304, N5045, N1414);
not NOT1 (N5286, N5269);
not NOT1 (N5287, N5284);
xor XOR2 (N5288, N5286, N3137);
and AND4 (N5289, N5287, N612, N2187, N2521);
not NOT1 (N5290, N5289);
nand NAND2 (N5291, N5280, N4179);
not NOT1 (N5292, N5260);
and AND4 (N5293, N5290, N955, N1976, N3899);
buf BUF1 (N5294, N5282);
not NOT1 (N5295, N5268);
not NOT1 (N5296, N5294);
or OR4 (N5297, N5279, N608, N1765, N508);
nand NAND4 (N5298, N5295, N795, N2158, N1782);
and AND3 (N5299, N5291, N4437, N3232);
and AND4 (N5300, N5296, N4895, N3835, N2280);
buf BUF1 (N5301, N5285);
buf BUF1 (N5302, N5298);
nand NAND4 (N5303, N5292, N3364, N4988, N2517);
nor NOR3 (N5304, N5301, N1682, N2986);
buf BUF1 (N5305, N5303);
not NOT1 (N5306, N5302);
or OR3 (N5307, N5288, N1045, N3679);
buf BUF1 (N5308, N5307);
nor NOR2 (N5309, N5274, N4476);
not NOT1 (N5310, N5297);
xor XOR2 (N5311, N5308, N941);
or OR4 (N5312, N5300, N389, N5246, N3222);
xor XOR2 (N5313, N5293, N4818);
nand NAND2 (N5314, N5305, N1275);
nor NOR2 (N5315, N5306, N1302);
or OR4 (N5316, N5304, N3690, N3814, N685);
not NOT1 (N5317, N5299);
or OR4 (N5318, N5316, N1103, N981, N2627);
not NOT1 (N5319, N5309);
nor NOR3 (N5320, N5314, N403, N4452);
buf BUF1 (N5321, N5311);
buf BUF1 (N5322, N5312);
buf BUF1 (N5323, N5281);
nand NAND4 (N5324, N5321, N2625, N4225, N2108);
nor NOR4 (N5325, N5319, N4954, N5268, N2697);
nor NOR2 (N5326, N5323, N139);
nor NOR3 (N5327, N5315, N373, N2196);
buf BUF1 (N5328, N5320);
buf BUF1 (N5329, N5325);
not NOT1 (N5330, N5317);
nor NOR4 (N5331, N5327, N3947, N1387, N4505);
and AND4 (N5332, N5326, N2001, N5005, N4056);
not NOT1 (N5333, N5328);
not NOT1 (N5334, N5322);
xor XOR2 (N5335, N5330, N4002);
not NOT1 (N5336, N5331);
and AND2 (N5337, N5332, N2534);
and AND2 (N5338, N5336, N1877);
buf BUF1 (N5339, N5337);
xor XOR2 (N5340, N5335, N5117);
or OR2 (N5341, N5313, N2757);
or OR2 (N5342, N5329, N4717);
buf BUF1 (N5343, N5339);
nand NAND2 (N5344, N5324, N1718);
nor NOR2 (N5345, N5344, N785);
and AND4 (N5346, N5343, N2595, N802, N865);
buf BUF1 (N5347, N5342);
xor XOR2 (N5348, N5340, N855);
nor NOR3 (N5349, N5345, N859, N2776);
or OR4 (N5350, N5338, N3435, N257, N2277);
buf BUF1 (N5351, N5346);
nor NOR4 (N5352, N5334, N3015, N3193, N1524);
nor NOR2 (N5353, N5352, N4103);
not NOT1 (N5354, N5310);
and AND4 (N5355, N5349, N1131, N1613, N994);
xor XOR2 (N5356, N5347, N4622);
nor NOR3 (N5357, N5354, N2620, N1597);
or OR2 (N5358, N5353, N3132);
and AND3 (N5359, N5341, N10, N4940);
or OR4 (N5360, N5333, N2709, N4630, N4023);
or OR3 (N5361, N5357, N1320, N1685);
and AND2 (N5362, N5359, N477);
and AND2 (N5363, N5355, N3373);
nand NAND4 (N5364, N5361, N3758, N2184, N2221);
not NOT1 (N5365, N5360);
nand NAND3 (N5366, N5364, N1071, N4553);
nor NOR3 (N5367, N5363, N3780, N3368);
or OR2 (N5368, N5362, N277);
xor XOR2 (N5369, N5348, N3816);
buf BUF1 (N5370, N5366);
buf BUF1 (N5371, N5318);
and AND4 (N5372, N5368, N3319, N2350, N2969);
buf BUF1 (N5373, N5358);
nand NAND3 (N5374, N5371, N1574, N568);
nand NAND4 (N5375, N5373, N654, N1857, N121);
or OR4 (N5376, N5367, N3304, N4106, N4325);
nand NAND3 (N5377, N5372, N4315, N4777);
and AND3 (N5378, N5374, N680, N5342);
nand NAND4 (N5379, N5370, N1271, N4815, N2588);
buf BUF1 (N5380, N5376);
nand NAND3 (N5381, N5378, N3602, N849);
nand NAND3 (N5382, N5377, N2882, N2350);
nand NAND4 (N5383, N5379, N5203, N1158, N321);
nor NOR4 (N5384, N5351, N4453, N146, N1489);
xor XOR2 (N5385, N5382, N3822);
xor XOR2 (N5386, N5384, N814);
nand NAND2 (N5387, N5380, N3758);
buf BUF1 (N5388, N5365);
nor NOR3 (N5389, N5375, N535, N2228);
xor XOR2 (N5390, N5369, N1199);
or OR2 (N5391, N5381, N3046);
nand NAND4 (N5392, N5350, N2472, N3868, N4390);
buf BUF1 (N5393, N5387);
and AND3 (N5394, N5383, N3349, N4153);
and AND3 (N5395, N5385, N1774, N2897);
nand NAND3 (N5396, N5389, N4317, N251);
nand NAND3 (N5397, N5395, N4926, N2636);
not NOT1 (N5398, N5397);
or OR2 (N5399, N5386, N3819);
or OR2 (N5400, N5391, N4355);
nor NOR4 (N5401, N5390, N4555, N71, N4131);
nor NOR4 (N5402, N5398, N482, N742, N903);
xor XOR2 (N5403, N5402, N1535);
xor XOR2 (N5404, N5394, N2828);
xor XOR2 (N5405, N5403, N4472);
nor NOR4 (N5406, N5393, N3188, N4955, N2542);
buf BUF1 (N5407, N5356);
not NOT1 (N5408, N5404);
buf BUF1 (N5409, N5399);
xor XOR2 (N5410, N5396, N1785);
nand NAND3 (N5411, N5405, N5113, N1483);
nor NOR4 (N5412, N5407, N4685, N2199, N2650);
and AND3 (N5413, N5400, N151, N1333);
not NOT1 (N5414, N5401);
not NOT1 (N5415, N5409);
nand NAND3 (N5416, N5413, N4685, N768);
or OR4 (N5417, N5392, N3006, N571, N3516);
buf BUF1 (N5418, N5415);
nor NOR2 (N5419, N5412, N4702);
xor XOR2 (N5420, N5406, N718);
not NOT1 (N5421, N5418);
or OR2 (N5422, N5419, N1761);
or OR3 (N5423, N5411, N908, N3654);
and AND3 (N5424, N5414, N2483, N5266);
or OR4 (N5425, N5408, N602, N2574, N1696);
nand NAND3 (N5426, N5420, N2272, N2401);
not NOT1 (N5427, N5422);
nor NOR2 (N5428, N5427, N924);
nand NAND2 (N5429, N5423, N278);
nand NAND2 (N5430, N5424, N4520);
and AND2 (N5431, N5426, N3962);
or OR2 (N5432, N5417, N3194);
xor XOR2 (N5433, N5410, N1169);
nor NOR4 (N5434, N5432, N2196, N1739, N2228);
not NOT1 (N5435, N5431);
nor NOR2 (N5436, N5421, N4421);
or OR4 (N5437, N5434, N1912, N5212, N785);
not NOT1 (N5438, N5437);
buf BUF1 (N5439, N5425);
and AND2 (N5440, N5430, N5234);
buf BUF1 (N5441, N5388);
xor XOR2 (N5442, N5438, N2647);
not NOT1 (N5443, N5416);
not NOT1 (N5444, N5433);
buf BUF1 (N5445, N5435);
and AND2 (N5446, N5439, N5316);
xor XOR2 (N5447, N5443, N3347);
or OR4 (N5448, N5436, N4974, N5412, N3121);
nand NAND4 (N5449, N5442, N216, N4822, N1471);
xor XOR2 (N5450, N5440, N2806);
xor XOR2 (N5451, N5449, N5331);
or OR3 (N5452, N5429, N2914, N4466);
nand NAND4 (N5453, N5441, N2705, N2393, N850);
not NOT1 (N5454, N5428);
and AND3 (N5455, N5453, N4847, N2321);
not NOT1 (N5456, N5451);
nand NAND3 (N5457, N5455, N2022, N585);
buf BUF1 (N5458, N5456);
not NOT1 (N5459, N5448);
and AND2 (N5460, N5458, N1912);
buf BUF1 (N5461, N5460);
nand NAND3 (N5462, N5444, N3412, N516);
nand NAND2 (N5463, N5450, N3814);
not NOT1 (N5464, N5452);
not NOT1 (N5465, N5447);
and AND4 (N5466, N5454, N3671, N1168, N2872);
buf BUF1 (N5467, N5465);
and AND2 (N5468, N5445, N3859);
xor XOR2 (N5469, N5457, N2721);
or OR4 (N5470, N5469, N5162, N2261, N4643);
buf BUF1 (N5471, N5467);
or OR4 (N5472, N5459, N4790, N4103, N4922);
buf BUF1 (N5473, N5461);
or OR4 (N5474, N5462, N5252, N2981, N4982);
or OR4 (N5475, N5471, N4236, N4248, N3708);
nand NAND4 (N5476, N5473, N4938, N2930, N5041);
nand NAND4 (N5477, N5468, N51, N1828, N610);
nand NAND4 (N5478, N5475, N3017, N2153, N1512);
not NOT1 (N5479, N5472);
nor NOR2 (N5480, N5476, N2035);
nor NOR4 (N5481, N5446, N3850, N1972, N560);
nor NOR3 (N5482, N5463, N5303, N783);
nand NAND4 (N5483, N5470, N1621, N935, N3765);
buf BUF1 (N5484, N5479);
xor XOR2 (N5485, N5482, N2355);
or OR3 (N5486, N5484, N4889, N2928);
nand NAND3 (N5487, N5474, N1038, N3304);
not NOT1 (N5488, N5478);
and AND4 (N5489, N5464, N5314, N1102, N4780);
xor XOR2 (N5490, N5477, N2777);
xor XOR2 (N5491, N5480, N3126);
xor XOR2 (N5492, N5488, N4164);
xor XOR2 (N5493, N5485, N1551);
buf BUF1 (N5494, N5490);
and AND2 (N5495, N5466, N3219);
or OR4 (N5496, N5493, N3260, N1500, N3671);
nor NOR2 (N5497, N5494, N1024);
not NOT1 (N5498, N5489);
or OR2 (N5499, N5491, N5287);
xor XOR2 (N5500, N5499, N290);
buf BUF1 (N5501, N5500);
not NOT1 (N5502, N5495);
xor XOR2 (N5503, N5492, N3701);
nor NOR2 (N5504, N5501, N3661);
not NOT1 (N5505, N5502);
or OR3 (N5506, N5497, N1222, N4719);
xor XOR2 (N5507, N5481, N4529);
buf BUF1 (N5508, N5498);
nor NOR3 (N5509, N5505, N4129, N2101);
xor XOR2 (N5510, N5486, N2844);
and AND2 (N5511, N5483, N1321);
and AND2 (N5512, N5506, N425);
xor XOR2 (N5513, N5487, N262);
nand NAND4 (N5514, N5508, N2213, N593, N4344);
or OR3 (N5515, N5507, N935, N174);
xor XOR2 (N5516, N5509, N3302);
buf BUF1 (N5517, N5504);
nor NOR2 (N5518, N5496, N5010);
or OR2 (N5519, N5516, N2402);
nand NAND4 (N5520, N5511, N586, N5333, N2849);
buf BUF1 (N5521, N5513);
nand NAND2 (N5522, N5515, N3118);
nor NOR4 (N5523, N5510, N4825, N852, N5048);
buf BUF1 (N5524, N5518);
and AND3 (N5525, N5522, N3306, N2476);
nand NAND4 (N5526, N5523, N761, N1238, N1360);
and AND3 (N5527, N5526, N3903, N3607);
nand NAND4 (N5528, N5512, N297, N4362, N4749);
or OR4 (N5529, N5519, N4937, N4954, N5302);
not NOT1 (N5530, N5528);
or OR4 (N5531, N5503, N1805, N3762, N4242);
or OR3 (N5532, N5529, N5490, N2172);
xor XOR2 (N5533, N5527, N15);
not NOT1 (N5534, N5533);
xor XOR2 (N5535, N5517, N4102);
nor NOR2 (N5536, N5521, N3919);
nand NAND3 (N5537, N5525, N3659, N826);
nand NAND3 (N5538, N5534, N3724, N961);
buf BUF1 (N5539, N5538);
not NOT1 (N5540, N5536);
buf BUF1 (N5541, N5540);
xor XOR2 (N5542, N5531, N1861);
xor XOR2 (N5543, N5532, N2549);
xor XOR2 (N5544, N5543, N5425);
and AND2 (N5545, N5537, N3907);
nor NOR4 (N5546, N5530, N3451, N3481, N4370);
and AND2 (N5547, N5545, N3277);
xor XOR2 (N5548, N5520, N2131);
buf BUF1 (N5549, N5541);
not NOT1 (N5550, N5535);
or OR2 (N5551, N5548, N872);
xor XOR2 (N5552, N5514, N5110);
nand NAND4 (N5553, N5542, N1745, N1724, N4245);
not NOT1 (N5554, N5553);
nor NOR4 (N5555, N5524, N714, N4637, N3449);
or OR2 (N5556, N5550, N4206);
or OR3 (N5557, N5552, N846, N2556);
or OR2 (N5558, N5539, N1030);
buf BUF1 (N5559, N5555);
buf BUF1 (N5560, N5557);
or OR2 (N5561, N5559, N1489);
nand NAND3 (N5562, N5544, N3466, N813);
and AND2 (N5563, N5551, N606);
or OR3 (N5564, N5554, N1661, N2880);
nand NAND3 (N5565, N5560, N3031, N2132);
and AND3 (N5566, N5564, N4162, N5190);
nor NOR3 (N5567, N5566, N3848, N2702);
or OR2 (N5568, N5563, N5069);
not NOT1 (N5569, N5568);
nor NOR2 (N5570, N5546, N2339);
buf BUF1 (N5571, N5565);
nand NAND2 (N5572, N5571, N100);
nor NOR3 (N5573, N5562, N2297, N2697);
nand NAND2 (N5574, N5547, N2377);
and AND3 (N5575, N5573, N3903, N3851);
or OR4 (N5576, N5570, N3929, N4040, N652);
buf BUF1 (N5577, N5576);
xor XOR2 (N5578, N5577, N2035);
xor XOR2 (N5579, N5569, N2162);
xor XOR2 (N5580, N5556, N1940);
buf BUF1 (N5581, N5575);
or OR4 (N5582, N5572, N2553, N54, N3138);
nand NAND3 (N5583, N5581, N2074, N5195);
or OR4 (N5584, N5561, N4990, N4697, N370);
and AND3 (N5585, N5567, N5332, N5396);
buf BUF1 (N5586, N5580);
xor XOR2 (N5587, N5585, N5072);
xor XOR2 (N5588, N5586, N2665);
not NOT1 (N5589, N5558);
nand NAND2 (N5590, N5587, N3498);
not NOT1 (N5591, N5588);
not NOT1 (N5592, N5574);
xor XOR2 (N5593, N5590, N2913);
not NOT1 (N5594, N5589);
or OR3 (N5595, N5592, N712, N674);
or OR2 (N5596, N5584, N5335);
nor NOR2 (N5597, N5594, N998);
nor NOR4 (N5598, N5595, N877, N2828, N1613);
nand NAND4 (N5599, N5597, N5141, N2000, N5030);
nor NOR3 (N5600, N5591, N885, N5348);
not NOT1 (N5601, N5596);
nand NAND2 (N5602, N5601, N1177);
nor NOR2 (N5603, N5582, N4641);
or OR3 (N5604, N5602, N2078, N2855);
and AND3 (N5605, N5593, N2684, N295);
nor NOR3 (N5606, N5599, N3388, N1791);
nand NAND4 (N5607, N5605, N1206, N2257, N4251);
not NOT1 (N5608, N5583);
not NOT1 (N5609, N5606);
buf BUF1 (N5610, N5604);
not NOT1 (N5611, N5578);
nand NAND4 (N5612, N5611, N3229, N791, N3907);
not NOT1 (N5613, N5609);
xor XOR2 (N5614, N5608, N4855);
or OR3 (N5615, N5610, N2663, N2652);
buf BUF1 (N5616, N5579);
buf BUF1 (N5617, N5613);
xor XOR2 (N5618, N5612, N2616);
or OR2 (N5619, N5614, N3433);
xor XOR2 (N5620, N5618, N3000);
xor XOR2 (N5621, N5615, N3908);
not NOT1 (N5622, N5619);
nor NOR4 (N5623, N5620, N3387, N4105, N250);
not NOT1 (N5624, N5616);
and AND4 (N5625, N5603, N679, N1804, N1476);
buf BUF1 (N5626, N5623);
buf BUF1 (N5627, N5624);
not NOT1 (N5628, N5600);
xor XOR2 (N5629, N5627, N4107);
nand NAND2 (N5630, N5629, N2860);
or OR2 (N5631, N5628, N360);
nor NOR3 (N5632, N5631, N645, N5329);
not NOT1 (N5633, N5625);
xor XOR2 (N5634, N5598, N3599);
xor XOR2 (N5635, N5634, N2388);
nor NOR4 (N5636, N5635, N2439, N3149, N1211);
nand NAND2 (N5637, N5549, N2694);
not NOT1 (N5638, N5622);
nand NAND4 (N5639, N5607, N905, N1594, N1940);
xor XOR2 (N5640, N5617, N361);
not NOT1 (N5641, N5636);
nand NAND4 (N5642, N5633, N1884, N4925, N4319);
buf BUF1 (N5643, N5638);
not NOT1 (N5644, N5637);
nor NOR2 (N5645, N5639, N5518);
nand NAND4 (N5646, N5643, N2801, N4036, N2034);
not NOT1 (N5647, N5621);
and AND3 (N5648, N5630, N2722, N2603);
or OR3 (N5649, N5626, N3182, N4003);
nor NOR3 (N5650, N5640, N5222, N850);
xor XOR2 (N5651, N5650, N3634);
nand NAND3 (N5652, N5645, N1458, N1497);
xor XOR2 (N5653, N5648, N5499);
or OR2 (N5654, N5651, N5404);
or OR3 (N5655, N5646, N2109, N3228);
buf BUF1 (N5656, N5641);
or OR4 (N5657, N5655, N1327, N5316, N3702);
nor NOR2 (N5658, N5647, N3777);
nor NOR3 (N5659, N5644, N591, N2825);
nand NAND2 (N5660, N5652, N72);
buf BUF1 (N5661, N5659);
and AND3 (N5662, N5656, N1326, N950);
buf BUF1 (N5663, N5657);
and AND2 (N5664, N5649, N4907);
nor NOR3 (N5665, N5654, N1314, N5579);
nand NAND3 (N5666, N5665, N3308, N5239);
nor NOR4 (N5667, N5660, N618, N2749, N1030);
buf BUF1 (N5668, N5632);
buf BUF1 (N5669, N5663);
or OR4 (N5670, N5668, N5565, N800, N2598);
nand NAND3 (N5671, N5669, N1335, N1902);
buf BUF1 (N5672, N5667);
xor XOR2 (N5673, N5670, N708);
not NOT1 (N5674, N5653);
and AND4 (N5675, N5674, N4351, N943, N1996);
not NOT1 (N5676, N5662);
nand NAND2 (N5677, N5672, N4325);
buf BUF1 (N5678, N5677);
nor NOR2 (N5679, N5642, N1592);
nor NOR2 (N5680, N5664, N2755);
xor XOR2 (N5681, N5673, N5180);
nand NAND4 (N5682, N5666, N4153, N3099, N3702);
or OR2 (N5683, N5679, N1387);
nand NAND3 (N5684, N5661, N1311, N4779);
and AND2 (N5685, N5684, N676);
nand NAND3 (N5686, N5678, N1318, N1128);
or OR2 (N5687, N5675, N2114);
not NOT1 (N5688, N5685);
or OR2 (N5689, N5682, N58);
nor NOR2 (N5690, N5681, N320);
or OR4 (N5691, N5683, N102, N5504, N1822);
buf BUF1 (N5692, N5658);
xor XOR2 (N5693, N5692, N26);
xor XOR2 (N5694, N5687, N3975);
not NOT1 (N5695, N5686);
or OR4 (N5696, N5680, N4172, N5225, N4421);
buf BUF1 (N5697, N5676);
not NOT1 (N5698, N5691);
not NOT1 (N5699, N5694);
not NOT1 (N5700, N5693);
not NOT1 (N5701, N5689);
buf BUF1 (N5702, N5695);
or OR4 (N5703, N5696, N5228, N3225, N234);
and AND2 (N5704, N5699, N5692);
not NOT1 (N5705, N5704);
and AND2 (N5706, N5698, N5313);
buf BUF1 (N5707, N5706);
xor XOR2 (N5708, N5705, N3407);
and AND4 (N5709, N5708, N1391, N5637, N4813);
nand NAND4 (N5710, N5702, N3494, N3258, N5315);
and AND3 (N5711, N5671, N2459, N2594);
buf BUF1 (N5712, N5701);
buf BUF1 (N5713, N5703);
or OR3 (N5714, N5711, N582, N4607);
buf BUF1 (N5715, N5713);
and AND3 (N5716, N5712, N297, N2130);
nor NOR4 (N5717, N5707, N5118, N5604, N2438);
xor XOR2 (N5718, N5709, N16);
or OR2 (N5719, N5700, N3755);
buf BUF1 (N5720, N5715);
nand NAND3 (N5721, N5720, N3765, N5166);
xor XOR2 (N5722, N5690, N1988);
nor NOR4 (N5723, N5688, N393, N887, N1512);
and AND4 (N5724, N5710, N68, N3778, N4400);
and AND3 (N5725, N5719, N1638, N2231);
buf BUF1 (N5726, N5724);
and AND3 (N5727, N5723, N3175, N101);
nand NAND2 (N5728, N5718, N539);
not NOT1 (N5729, N5721);
or OR3 (N5730, N5722, N3320, N4241);
xor XOR2 (N5731, N5730, N849);
not NOT1 (N5732, N5716);
or OR4 (N5733, N5725, N435, N4058, N43);
nor NOR4 (N5734, N5717, N4606, N104, N681);
nand NAND4 (N5735, N5732, N5314, N3583, N4988);
not NOT1 (N5736, N5714);
not NOT1 (N5737, N5734);
and AND3 (N5738, N5728, N2480, N4215);
buf BUF1 (N5739, N5737);
or OR3 (N5740, N5733, N505, N1295);
buf BUF1 (N5741, N5735);
nor NOR4 (N5742, N5697, N5612, N865, N4781);
nor NOR3 (N5743, N5727, N447, N3379);
xor XOR2 (N5744, N5743, N5464);
nor NOR3 (N5745, N5726, N476, N451);
nand NAND4 (N5746, N5736, N426, N4379, N2961);
buf BUF1 (N5747, N5741);
not NOT1 (N5748, N5738);
nor NOR3 (N5749, N5740, N4514, N1626);
or OR3 (N5750, N5731, N4857, N843);
and AND4 (N5751, N5747, N5336, N1923, N3975);
xor XOR2 (N5752, N5744, N4906);
and AND3 (N5753, N5739, N4391, N4404);
not NOT1 (N5754, N5750);
or OR2 (N5755, N5729, N2932);
nand NAND4 (N5756, N5754, N5709, N481, N5405);
nand NAND2 (N5757, N5753, N1294);
not NOT1 (N5758, N5752);
not NOT1 (N5759, N5758);
nand NAND4 (N5760, N5751, N2762, N3619, N1617);
xor XOR2 (N5761, N5756, N3582);
xor XOR2 (N5762, N5759, N5565);
buf BUF1 (N5763, N5745);
nor NOR4 (N5764, N5749, N5695, N2756, N3774);
xor XOR2 (N5765, N5746, N3216);
nor NOR3 (N5766, N5755, N1920, N5695);
nor NOR3 (N5767, N5757, N1208, N447);
xor XOR2 (N5768, N5762, N3423);
buf BUF1 (N5769, N5761);
nand NAND4 (N5770, N5760, N216, N747, N5221);
buf BUF1 (N5771, N5748);
not NOT1 (N5772, N5765);
and AND2 (N5773, N5763, N2795);
nor NOR4 (N5774, N5769, N192, N4827, N3157);
nor NOR2 (N5775, N5742, N2861);
xor XOR2 (N5776, N5775, N2475);
and AND2 (N5777, N5764, N2486);
not NOT1 (N5778, N5774);
xor XOR2 (N5779, N5773, N5608);
buf BUF1 (N5780, N5779);
xor XOR2 (N5781, N5776, N2759);
and AND3 (N5782, N5772, N1804, N3393);
and AND3 (N5783, N5771, N3896, N2836);
nor NOR4 (N5784, N5781, N1742, N770, N1935);
nor NOR4 (N5785, N5782, N3099, N220, N3029);
xor XOR2 (N5786, N5768, N1808);
not NOT1 (N5787, N5777);
nand NAND4 (N5788, N5766, N3562, N425, N191);
and AND4 (N5789, N5778, N738, N3064, N3962);
and AND4 (N5790, N5786, N5174, N1648, N5077);
nand NAND4 (N5791, N5770, N4988, N2193, N3994);
and AND4 (N5792, N5789, N3865, N3982, N4030);
not NOT1 (N5793, N5767);
buf BUF1 (N5794, N5791);
and AND4 (N5795, N5785, N5334, N1425, N4765);
xor XOR2 (N5796, N5787, N5683);
and AND3 (N5797, N5784, N5346, N1096);
xor XOR2 (N5798, N5793, N3627);
or OR3 (N5799, N5798, N1533, N2085);
and AND2 (N5800, N5795, N5649);
nor NOR3 (N5801, N5796, N5672, N4794);
not NOT1 (N5802, N5780);
xor XOR2 (N5803, N5797, N1626);
buf BUF1 (N5804, N5794);
xor XOR2 (N5805, N5799, N5652);
nand NAND4 (N5806, N5792, N3371, N2791, N4532);
buf BUF1 (N5807, N5804);
xor XOR2 (N5808, N5788, N4847);
buf BUF1 (N5809, N5783);
not NOT1 (N5810, N5803);
nand NAND4 (N5811, N5808, N2580, N1797, N5178);
nand NAND3 (N5812, N5810, N3645, N2991);
or OR4 (N5813, N5802, N1701, N3831, N326);
buf BUF1 (N5814, N5807);
xor XOR2 (N5815, N5813, N2296);
nor NOR4 (N5816, N5811, N1160, N1526, N1415);
or OR4 (N5817, N5814, N5733, N404, N4816);
xor XOR2 (N5818, N5806, N4564);
buf BUF1 (N5819, N5800);
not NOT1 (N5820, N5801);
nor NOR2 (N5821, N5816, N2683);
nor NOR4 (N5822, N5815, N1647, N644, N2834);
nand NAND3 (N5823, N5821, N3191, N725);
nor NOR4 (N5824, N5817, N2329, N2082, N1197);
or OR2 (N5825, N5809, N1906);
nor NOR2 (N5826, N5822, N3754);
nor NOR2 (N5827, N5819, N4738);
and AND4 (N5828, N5812, N1466, N3859, N547);
nand NAND3 (N5829, N5828, N4649, N2473);
buf BUF1 (N5830, N5818);
and AND2 (N5831, N5825, N4207);
xor XOR2 (N5832, N5826, N4108);
and AND3 (N5833, N5829, N342, N5526);
buf BUF1 (N5834, N5830);
and AND3 (N5835, N5820, N251, N2147);
nand NAND4 (N5836, N5834, N27, N4954, N1831);
and AND3 (N5837, N5831, N5490, N553);
or OR2 (N5838, N5837, N756);
and AND2 (N5839, N5790, N5831);
xor XOR2 (N5840, N5827, N1522);
buf BUF1 (N5841, N5836);
xor XOR2 (N5842, N5805, N2486);
not NOT1 (N5843, N5839);
not NOT1 (N5844, N5841);
and AND4 (N5845, N5832, N4176, N5369, N1430);
not NOT1 (N5846, N5833);
nand NAND4 (N5847, N5824, N1486, N1472, N808);
nand NAND4 (N5848, N5844, N1087, N4632, N445);
or OR4 (N5849, N5840, N1504, N5144, N5148);
not NOT1 (N5850, N5835);
or OR2 (N5851, N5823, N690);
xor XOR2 (N5852, N5850, N4785);
nor NOR3 (N5853, N5845, N419, N3814);
xor XOR2 (N5854, N5853, N895);
nor NOR3 (N5855, N5849, N5199, N1021);
buf BUF1 (N5856, N5854);
nor NOR2 (N5857, N5856, N219);
and AND4 (N5858, N5843, N3113, N509, N1320);
nand NAND4 (N5859, N5857, N3732, N3232, N5018);
buf BUF1 (N5860, N5842);
nor NOR3 (N5861, N5860, N5295, N4958);
nand NAND4 (N5862, N5858, N1160, N1294, N3752);
nand NAND4 (N5863, N5852, N122, N2015, N2808);
and AND4 (N5864, N5847, N4398, N1523, N4356);
not NOT1 (N5865, N5864);
not NOT1 (N5866, N5855);
xor XOR2 (N5867, N5861, N243);
and AND4 (N5868, N5862, N4401, N2754, N2047);
nand NAND4 (N5869, N5848, N3714, N4514, N4068);
and AND4 (N5870, N5865, N2893, N2470, N18);
or OR4 (N5871, N5851, N4967, N278, N5436);
nand NAND2 (N5872, N5846, N3893);
or OR4 (N5873, N5863, N232, N1721, N3685);
buf BUF1 (N5874, N5871);
buf BUF1 (N5875, N5870);
buf BUF1 (N5876, N5838);
or OR4 (N5877, N5872, N3545, N1004, N3544);
nand NAND3 (N5878, N5866, N2565, N4904);
nor NOR2 (N5879, N5868, N2962);
or OR2 (N5880, N5878, N5313);
not NOT1 (N5881, N5867);
and AND4 (N5882, N5876, N3829, N1947, N3904);
buf BUF1 (N5883, N5859);
buf BUF1 (N5884, N5881);
buf BUF1 (N5885, N5874);
nand NAND2 (N5886, N5869, N1784);
nand NAND2 (N5887, N5873, N5170);
xor XOR2 (N5888, N5883, N4562);
nor NOR2 (N5889, N5888, N428);
xor XOR2 (N5890, N5889, N2874);
xor XOR2 (N5891, N5882, N1186);
buf BUF1 (N5892, N5880);
not NOT1 (N5893, N5879);
not NOT1 (N5894, N5887);
nor NOR2 (N5895, N5893, N1094);
or OR4 (N5896, N5894, N992, N4696, N3550);
xor XOR2 (N5897, N5891, N5281);
buf BUF1 (N5898, N5892);
buf BUF1 (N5899, N5898);
not NOT1 (N5900, N5899);
xor XOR2 (N5901, N5877, N408);
and AND2 (N5902, N5875, N1885);
not NOT1 (N5903, N5895);
buf BUF1 (N5904, N5901);
and AND3 (N5905, N5900, N118, N5409);
xor XOR2 (N5906, N5903, N3133);
or OR3 (N5907, N5905, N3636, N4534);
nand NAND4 (N5908, N5885, N1015, N1946, N4959);
nand NAND4 (N5909, N5886, N5232, N1281, N2652);
xor XOR2 (N5910, N5897, N2362);
nand NAND2 (N5911, N5904, N3262);
nor NOR4 (N5912, N5911, N5295, N868, N1373);
not NOT1 (N5913, N5912);
nor NOR3 (N5914, N5907, N3761, N5697);
xor XOR2 (N5915, N5906, N4755);
not NOT1 (N5916, N5908);
nand NAND3 (N5917, N5896, N349, N5597);
xor XOR2 (N5918, N5909, N5502);
not NOT1 (N5919, N5915);
nor NOR4 (N5920, N5917, N3000, N380, N4932);
nor NOR4 (N5921, N5884, N3473, N1577, N5780);
and AND2 (N5922, N5890, N2119);
nand NAND2 (N5923, N5916, N5275);
or OR3 (N5924, N5920, N4452, N2227);
buf BUF1 (N5925, N5923);
buf BUF1 (N5926, N5914);
xor XOR2 (N5927, N5910, N3257);
xor XOR2 (N5928, N5919, N4119);
buf BUF1 (N5929, N5924);
not NOT1 (N5930, N5929);
xor XOR2 (N5931, N5913, N5746);
buf BUF1 (N5932, N5921);
nor NOR3 (N5933, N5931, N149, N5200);
buf BUF1 (N5934, N5902);
xor XOR2 (N5935, N5918, N3394);
and AND3 (N5936, N5932, N1349, N4897);
and AND4 (N5937, N5925, N5770, N3780, N1205);
buf BUF1 (N5938, N5936);
buf BUF1 (N5939, N5938);
not NOT1 (N5940, N5930);
nand NAND3 (N5941, N5939, N2270, N1703);
buf BUF1 (N5942, N5926);
nor NOR2 (N5943, N5933, N2532);
and AND2 (N5944, N5940, N2601);
and AND4 (N5945, N5944, N2512, N472, N3133);
not NOT1 (N5946, N5941);
nand NAND4 (N5947, N5937, N5157, N962, N5346);
and AND3 (N5948, N5942, N861, N1543);
nor NOR4 (N5949, N5947, N4608, N522, N837);
or OR3 (N5950, N5946, N3952, N2207);
buf BUF1 (N5951, N5934);
and AND2 (N5952, N5949, N1607);
nor NOR2 (N5953, N5948, N3958);
or OR2 (N5954, N5953, N2515);
and AND2 (N5955, N5922, N1360);
or OR4 (N5956, N5954, N4787, N1810, N993);
nor NOR2 (N5957, N5927, N3740);
or OR3 (N5958, N5951, N4335, N3855);
buf BUF1 (N5959, N5935);
and AND2 (N5960, N5956, N5668);
or OR2 (N5961, N5943, N2081);
nand NAND3 (N5962, N5945, N1193, N5927);
nand NAND2 (N5963, N5960, N4596);
and AND4 (N5964, N5950, N3824, N894, N1268);
buf BUF1 (N5965, N5961);
buf BUF1 (N5966, N5965);
not NOT1 (N5967, N5952);
nor NOR3 (N5968, N5959, N3710, N5855);
nor NOR2 (N5969, N5968, N2720);
nor NOR4 (N5970, N5969, N5856, N225, N3287);
not NOT1 (N5971, N5966);
nand NAND4 (N5972, N5964, N383, N5712, N4839);
nand NAND4 (N5973, N5971, N5757, N3882, N2108);
nand NAND2 (N5974, N5928, N5004);
and AND4 (N5975, N5955, N1885, N4705, N3305);
xor XOR2 (N5976, N5975, N3652);
xor XOR2 (N5977, N5957, N2383);
nand NAND4 (N5978, N5973, N527, N2261, N4546);
nor NOR3 (N5979, N5974, N5124, N635);
xor XOR2 (N5980, N5962, N2215);
and AND2 (N5981, N5967, N964);
not NOT1 (N5982, N5980);
xor XOR2 (N5983, N5976, N4157);
xor XOR2 (N5984, N5979, N4508);
nor NOR4 (N5985, N5972, N5347, N4163, N4095);
nor NOR4 (N5986, N5963, N3662, N5513, N4519);
not NOT1 (N5987, N5983);
not NOT1 (N5988, N5987);
buf BUF1 (N5989, N5985);
or OR3 (N5990, N5981, N1825, N4342);
nor NOR2 (N5991, N5984, N1539);
buf BUF1 (N5992, N5989);
nor NOR4 (N5993, N5977, N1844, N4068, N4151);
nand NAND3 (N5994, N5978, N3992, N1476);
nand NAND2 (N5995, N5986, N3282);
not NOT1 (N5996, N5958);
buf BUF1 (N5997, N5994);
xor XOR2 (N5998, N5997, N2400);
not NOT1 (N5999, N5970);
not NOT1 (N6000, N5993);
buf BUF1 (N6001, N5991);
buf BUF1 (N6002, N5999);
xor XOR2 (N6003, N5988, N4766);
not NOT1 (N6004, N5998);
buf BUF1 (N6005, N6003);
nand NAND3 (N6006, N5992, N4228, N1677);
and AND3 (N6007, N5996, N3484, N1191);
not NOT1 (N6008, N6004);
nor NOR4 (N6009, N6008, N3706, N2949, N3153);
or OR4 (N6010, N5995, N1024, N4923, N1570);
buf BUF1 (N6011, N6000);
buf BUF1 (N6012, N6006);
or OR4 (N6013, N6010, N4744, N4104, N5391);
buf BUF1 (N6014, N6009);
nor NOR2 (N6015, N5990, N4915);
not NOT1 (N6016, N6011);
nand NAND4 (N6017, N6014, N1165, N5822, N4515);
nor NOR4 (N6018, N6001, N5745, N3792, N3451);
nor NOR3 (N6019, N6007, N5004, N3752);
nor NOR4 (N6020, N5982, N3980, N5776, N100);
and AND3 (N6021, N6002, N5510, N3861);
not NOT1 (N6022, N6021);
xor XOR2 (N6023, N6018, N2500);
and AND3 (N6024, N6022, N2906, N2727);
not NOT1 (N6025, N6005);
not NOT1 (N6026, N6016);
nor NOR4 (N6027, N6025, N3702, N913, N23);
nor NOR3 (N6028, N6023, N2973, N3973);
xor XOR2 (N6029, N6015, N3064);
buf BUF1 (N6030, N6028);
or OR2 (N6031, N6012, N5825);
nor NOR2 (N6032, N6013, N1337);
and AND2 (N6033, N6031, N5902);
or OR3 (N6034, N6017, N3139, N3351);
nor NOR4 (N6035, N6033, N1620, N4883, N6024);
nand NAND2 (N6036, N4959, N4999);
buf BUF1 (N6037, N6036);
buf BUF1 (N6038, N6026);
not NOT1 (N6039, N6029);
nor NOR4 (N6040, N6039, N455, N516, N1750);
nand NAND4 (N6041, N6038, N5332, N3650, N4972);
and AND2 (N6042, N6034, N3668);
nor NOR4 (N6043, N6019, N159, N2823, N4257);
or OR4 (N6044, N6042, N5571, N110, N5040);
not NOT1 (N6045, N6020);
nor NOR4 (N6046, N6043, N397, N2372, N3065);
nand NAND2 (N6047, N6040, N5745);
not NOT1 (N6048, N6037);
nor NOR2 (N6049, N6032, N4200);
buf BUF1 (N6050, N6041);
nor NOR2 (N6051, N6035, N1106);
buf BUF1 (N6052, N6046);
nor NOR3 (N6053, N6048, N3979, N2081);
and AND4 (N6054, N6053, N4458, N3873, N4459);
nor NOR2 (N6055, N6052, N5027);
buf BUF1 (N6056, N6054);
buf BUF1 (N6057, N6049);
nor NOR2 (N6058, N6027, N5902);
nand NAND2 (N6059, N6044, N4227);
nor NOR3 (N6060, N6030, N5779, N5553);
nand NAND2 (N6061, N6059, N2233);
and AND4 (N6062, N6047, N2964, N4855, N2870);
not NOT1 (N6063, N6058);
and AND3 (N6064, N6057, N2050, N5791);
xor XOR2 (N6065, N6064, N2733);
xor XOR2 (N6066, N6065, N4557);
nand NAND4 (N6067, N6056, N4212, N5685, N474);
xor XOR2 (N6068, N6045, N2104);
not NOT1 (N6069, N6060);
not NOT1 (N6070, N6067);
nor NOR2 (N6071, N6069, N3972);
nor NOR2 (N6072, N6061, N757);
buf BUF1 (N6073, N6051);
and AND3 (N6074, N6073, N3159, N949);
nor NOR3 (N6075, N6055, N5076, N185);
or OR3 (N6076, N6068, N2934, N1602);
xor XOR2 (N6077, N6072, N2443);
or OR2 (N6078, N6050, N1077);
not NOT1 (N6079, N6070);
buf BUF1 (N6080, N6075);
or OR3 (N6081, N6080, N1468, N2812);
nand NAND4 (N6082, N6081, N2207, N5735, N2723);
and AND2 (N6083, N6079, N2738);
and AND4 (N6084, N6076, N3871, N1271, N2249);
xor XOR2 (N6085, N6063, N5807);
nand NAND2 (N6086, N6074, N4681);
nor NOR3 (N6087, N6082, N2140, N1121);
or OR3 (N6088, N6078, N125, N503);
xor XOR2 (N6089, N6086, N3954);
and AND3 (N6090, N6088, N2215, N2290);
nand NAND2 (N6091, N6087, N1152);
nor NOR3 (N6092, N6089, N4259, N3487);
nor NOR3 (N6093, N6085, N4442, N504);
or OR2 (N6094, N6071, N3945);
nor NOR4 (N6095, N6091, N5712, N337, N5592);
buf BUF1 (N6096, N6092);
or OR3 (N6097, N6094, N437, N1919);
nand NAND3 (N6098, N6090, N1523, N2945);
or OR3 (N6099, N6083, N4747, N2718);
or OR2 (N6100, N6084, N159);
nand NAND2 (N6101, N6095, N2497);
xor XOR2 (N6102, N6101, N1175);
nor NOR3 (N6103, N6097, N2830, N1229);
and AND4 (N6104, N6093, N1845, N2587, N1861);
xor XOR2 (N6105, N6102, N4365);
not NOT1 (N6106, N6099);
buf BUF1 (N6107, N6103);
buf BUF1 (N6108, N6062);
and AND3 (N6109, N6105, N5964, N5271);
or OR2 (N6110, N6098, N2768);
buf BUF1 (N6111, N6107);
xor XOR2 (N6112, N6111, N67);
buf BUF1 (N6113, N6112);
and AND4 (N6114, N6113, N813, N2727, N1038);
or OR3 (N6115, N6106, N3399, N4046);
and AND4 (N6116, N6096, N5778, N3056, N596);
nor NOR4 (N6117, N6115, N3227, N3776, N3599);
nor NOR2 (N6118, N6117, N3350);
nor NOR4 (N6119, N6116, N5281, N1215, N3982);
nor NOR4 (N6120, N6109, N1051, N664, N1158);
nand NAND2 (N6121, N6114, N335);
nand NAND4 (N6122, N6119, N3016, N4518, N3720);
nor NOR2 (N6123, N6104, N2387);
xor XOR2 (N6124, N6108, N5504);
buf BUF1 (N6125, N6100);
nand NAND4 (N6126, N6123, N3204, N2220, N309);
buf BUF1 (N6127, N6126);
and AND2 (N6128, N6121, N3342);
buf BUF1 (N6129, N6118);
or OR2 (N6130, N6124, N3560);
nor NOR4 (N6131, N6110, N450, N4796, N3095);
xor XOR2 (N6132, N6131, N3951);
or OR4 (N6133, N6127, N5719, N2446, N2042);
nor NOR4 (N6134, N6122, N817, N2685, N1462);
buf BUF1 (N6135, N6133);
buf BUF1 (N6136, N6128);
xor XOR2 (N6137, N6120, N4293);
not NOT1 (N6138, N6137);
nor NOR4 (N6139, N6129, N1293, N5936, N5705);
nand NAND3 (N6140, N6125, N1319, N1837);
not NOT1 (N6141, N6138);
nor NOR2 (N6142, N6135, N1419);
and AND2 (N6143, N6130, N1524);
nor NOR2 (N6144, N6139, N3647);
and AND4 (N6145, N6142, N1821, N5104, N3986);
nor NOR2 (N6146, N6134, N355);
or OR4 (N6147, N6146, N502, N173, N3145);
buf BUF1 (N6148, N6141);
not NOT1 (N6149, N6148);
and AND3 (N6150, N6145, N248, N6127);
nand NAND2 (N6151, N6066, N1373);
not NOT1 (N6152, N6144);
and AND4 (N6153, N6143, N4641, N4565, N1426);
nand NAND3 (N6154, N6152, N5065, N602);
nand NAND4 (N6155, N6077, N5028, N4812, N3384);
buf BUF1 (N6156, N6154);
nand NAND3 (N6157, N6136, N3036, N5486);
not NOT1 (N6158, N6157);
nand NAND3 (N6159, N6158, N1321, N1812);
buf BUF1 (N6160, N6156);
not NOT1 (N6161, N6140);
xor XOR2 (N6162, N6153, N2234);
buf BUF1 (N6163, N6149);
or OR4 (N6164, N6151, N3113, N957, N3740);
or OR2 (N6165, N6162, N3493);
not NOT1 (N6166, N6164);
or OR2 (N6167, N6166, N1748);
not NOT1 (N6168, N6159);
nand NAND4 (N6169, N6132, N5736, N5705, N2130);
or OR2 (N6170, N6161, N1490);
xor XOR2 (N6171, N6160, N2659);
and AND4 (N6172, N6167, N3240, N1328, N2819);
not NOT1 (N6173, N6168);
not NOT1 (N6174, N6169);
nor NOR2 (N6175, N6147, N1368);
not NOT1 (N6176, N6175);
nor NOR3 (N6177, N6165, N2624, N1111);
xor XOR2 (N6178, N6155, N32);
or OR3 (N6179, N6173, N4031, N1883);
and AND3 (N6180, N6179, N1081, N4326);
or OR4 (N6181, N6178, N3825, N1994, N1880);
not NOT1 (N6182, N6163);
or OR3 (N6183, N6172, N2832, N822);
and AND2 (N6184, N6176, N5204);
buf BUF1 (N6185, N6150);
nand NAND4 (N6186, N6170, N3308, N443, N494);
nand NAND3 (N6187, N6171, N618, N4113);
nor NOR4 (N6188, N6183, N1457, N3341, N3882);
buf BUF1 (N6189, N6180);
buf BUF1 (N6190, N6189);
or OR3 (N6191, N6181, N1718, N5911);
xor XOR2 (N6192, N6191, N2676);
not NOT1 (N6193, N6187);
or OR4 (N6194, N6177, N2482, N4918, N2671);
and AND2 (N6195, N6192, N5842);
and AND3 (N6196, N6174, N4932, N1946);
and AND2 (N6197, N6186, N1271);
xor XOR2 (N6198, N6194, N4846);
or OR2 (N6199, N6190, N2604);
nor NOR3 (N6200, N6184, N2324, N2105);
nand NAND3 (N6201, N6199, N2516, N1961);
nand NAND3 (N6202, N6185, N718, N4686);
or OR2 (N6203, N6196, N3262);
or OR4 (N6204, N6182, N3465, N5897, N3506);
nand NAND2 (N6205, N6203, N692);
and AND2 (N6206, N6198, N5127);
not NOT1 (N6207, N6195);
buf BUF1 (N6208, N6204);
or OR2 (N6209, N6206, N526);
or OR2 (N6210, N6205, N1018);
not NOT1 (N6211, N6200);
not NOT1 (N6212, N6193);
nor NOR4 (N6213, N6207, N1261, N4776, N5186);
and AND3 (N6214, N6213, N4096, N642);
not NOT1 (N6215, N6202);
nor NOR3 (N6216, N6197, N6062, N566);
nand NAND3 (N6217, N6214, N4569, N3801);
buf BUF1 (N6218, N6212);
and AND2 (N6219, N6211, N3338);
nor NOR2 (N6220, N6216, N1624);
xor XOR2 (N6221, N6201, N589);
not NOT1 (N6222, N6188);
or OR4 (N6223, N6219, N2521, N2027, N2896);
xor XOR2 (N6224, N6209, N5829);
xor XOR2 (N6225, N6218, N4720);
nor NOR4 (N6226, N6224, N4291, N2377, N4945);
buf BUF1 (N6227, N6220);
xor XOR2 (N6228, N6215, N1887);
nor NOR2 (N6229, N6227, N4352);
or OR2 (N6230, N6228, N1879);
and AND2 (N6231, N6217, N3056);
nor NOR4 (N6232, N6221, N1567, N4346, N2663);
nand NAND4 (N6233, N6223, N1508, N1896, N5149);
or OR3 (N6234, N6222, N4437, N5049);
nand NAND4 (N6235, N6234, N2195, N3279, N4776);
xor XOR2 (N6236, N6235, N5588);
xor XOR2 (N6237, N6226, N3940);
buf BUF1 (N6238, N6210);
or OR3 (N6239, N6230, N3385, N1257);
nor NOR2 (N6240, N6225, N4310);
and AND3 (N6241, N6232, N5307, N5224);
nand NAND4 (N6242, N6229, N5074, N1497, N503);
and AND2 (N6243, N6242, N4182);
or OR3 (N6244, N6231, N4978, N182);
not NOT1 (N6245, N6244);
nand NAND4 (N6246, N6233, N6015, N2495, N1795);
and AND4 (N6247, N6208, N3216, N676, N2242);
xor XOR2 (N6248, N6239, N5781);
buf BUF1 (N6249, N6243);
not NOT1 (N6250, N6237);
xor XOR2 (N6251, N6246, N5906);
or OR2 (N6252, N6236, N2171);
buf BUF1 (N6253, N6245);
and AND3 (N6254, N6238, N4663, N759);
buf BUF1 (N6255, N6252);
or OR2 (N6256, N6250, N4430);
or OR4 (N6257, N6255, N1504, N5443, N3358);
xor XOR2 (N6258, N6257, N5752);
or OR3 (N6259, N6254, N1366, N435);
and AND4 (N6260, N6251, N1835, N2259, N3697);
and AND3 (N6261, N6240, N2249, N2548);
buf BUF1 (N6262, N6260);
nand NAND4 (N6263, N6247, N841, N464, N4484);
nand NAND3 (N6264, N6263, N1868, N4857);
not NOT1 (N6265, N6241);
nand NAND4 (N6266, N6262, N9, N2339, N3487);
buf BUF1 (N6267, N6249);
and AND2 (N6268, N6261, N755);
nor NOR3 (N6269, N6258, N1604, N5097);
nor NOR4 (N6270, N6256, N505, N4168, N3305);
nor NOR2 (N6271, N6253, N4713);
buf BUF1 (N6272, N6266);
buf BUF1 (N6273, N6265);
or OR2 (N6274, N6264, N4540);
or OR3 (N6275, N6267, N3913, N3351);
nor NOR4 (N6276, N6273, N5652, N1627, N5397);
buf BUF1 (N6277, N6271);
nor NOR4 (N6278, N6269, N2983, N1811, N114);
or OR2 (N6279, N6276, N1470);
and AND4 (N6280, N6277, N6108, N104, N3351);
not NOT1 (N6281, N6259);
or OR4 (N6282, N6279, N3923, N5879, N2054);
nor NOR4 (N6283, N6282, N1322, N2257, N606);
xor XOR2 (N6284, N6274, N3036);
nor NOR4 (N6285, N6280, N2062, N3737, N1870);
buf BUF1 (N6286, N6275);
xor XOR2 (N6287, N6270, N952);
xor XOR2 (N6288, N6278, N2941);
and AND4 (N6289, N6281, N4627, N5142, N5752);
and AND3 (N6290, N6288, N3044, N795);
nand NAND4 (N6291, N6272, N486, N1194, N3626);
and AND3 (N6292, N6248, N5408, N958);
not NOT1 (N6293, N6268);
xor XOR2 (N6294, N6284, N4494);
not NOT1 (N6295, N6294);
nor NOR3 (N6296, N6289, N2798, N270);
or OR2 (N6297, N6287, N3502);
nand NAND4 (N6298, N6291, N5725, N1567, N3316);
xor XOR2 (N6299, N6285, N2284);
nor NOR3 (N6300, N6286, N6014, N4780);
nand NAND2 (N6301, N6299, N4864);
nor NOR3 (N6302, N6292, N5584, N2463);
nand NAND2 (N6303, N6301, N5144);
xor XOR2 (N6304, N6297, N469);
xor XOR2 (N6305, N6290, N4961);
nor NOR3 (N6306, N6305, N3768, N448);
or OR3 (N6307, N6296, N1926, N2788);
nor NOR3 (N6308, N6307, N4789, N767);
and AND2 (N6309, N6304, N2052);
xor XOR2 (N6310, N6300, N483);
not NOT1 (N6311, N6309);
nor NOR4 (N6312, N6310, N3790, N4165, N1709);
nor NOR3 (N6313, N6311, N5512, N5869);
not NOT1 (N6314, N6312);
or OR2 (N6315, N6308, N3868);
xor XOR2 (N6316, N6293, N5678);
nand NAND3 (N6317, N6303, N6096, N5061);
nand NAND4 (N6318, N6314, N26, N4006, N4594);
nand NAND3 (N6319, N6317, N5432, N1747);
nand NAND3 (N6320, N6315, N3537, N5571);
nor NOR4 (N6321, N6298, N883, N4473, N5541);
xor XOR2 (N6322, N6320, N3531);
not NOT1 (N6323, N6322);
nand NAND3 (N6324, N6319, N1129, N6089);
not NOT1 (N6325, N6323);
nand NAND2 (N6326, N6306, N3782);
or OR4 (N6327, N6326, N2112, N5092, N1964);
nand NAND3 (N6328, N6318, N1443, N3673);
nand NAND4 (N6329, N6313, N81, N4490, N1146);
buf BUF1 (N6330, N6295);
buf BUF1 (N6331, N6327);
not NOT1 (N6332, N6331);
xor XOR2 (N6333, N6283, N1368);
not NOT1 (N6334, N6316);
nand NAND4 (N6335, N6330, N830, N4688, N2539);
xor XOR2 (N6336, N6333, N2207);
xor XOR2 (N6337, N6321, N1711);
buf BUF1 (N6338, N6302);
nor NOR4 (N6339, N6332, N651, N6108, N5629);
buf BUF1 (N6340, N6329);
not NOT1 (N6341, N6337);
buf BUF1 (N6342, N6325);
xor XOR2 (N6343, N6334, N2759);
xor XOR2 (N6344, N6342, N564);
and AND3 (N6345, N6338, N4813, N1524);
buf BUF1 (N6346, N6336);
nand NAND4 (N6347, N6335, N6209, N2733, N2633);
nor NOR4 (N6348, N6324, N816, N3281, N423);
or OR2 (N6349, N6348, N4928);
buf BUF1 (N6350, N6349);
buf BUF1 (N6351, N6345);
or OR2 (N6352, N6344, N3919);
not NOT1 (N6353, N6350);
and AND2 (N6354, N6353, N82);
xor XOR2 (N6355, N6328, N1716);
and AND3 (N6356, N6352, N5418, N2960);
nand NAND2 (N6357, N6351, N1759);
and AND2 (N6358, N6356, N2440);
or OR4 (N6359, N6358, N2707, N2695, N3266);
and AND2 (N6360, N6340, N2249);
not NOT1 (N6361, N6343);
nor NOR3 (N6362, N6359, N1465, N1678);
buf BUF1 (N6363, N6354);
or OR3 (N6364, N6357, N226, N989);
or OR2 (N6365, N6360, N4877);
buf BUF1 (N6366, N6363);
nand NAND2 (N6367, N6364, N5164);
not NOT1 (N6368, N6355);
not NOT1 (N6369, N6365);
nor NOR4 (N6370, N6339, N3991, N5931, N3817);
and AND2 (N6371, N6347, N5194);
or OR3 (N6372, N6362, N5740, N5627);
not NOT1 (N6373, N6361);
and AND2 (N6374, N6372, N6285);
nor NOR4 (N6375, N6341, N5485, N5774, N2730);
not NOT1 (N6376, N6346);
or OR3 (N6377, N6366, N5637, N4150);
or OR2 (N6378, N6376, N2450);
or OR2 (N6379, N6367, N6191);
or OR3 (N6380, N6368, N4575, N622);
xor XOR2 (N6381, N6377, N3339);
nor NOR3 (N6382, N6378, N844, N205);
and AND3 (N6383, N6381, N877, N1506);
or OR4 (N6384, N6379, N3686, N5293, N1812);
or OR2 (N6385, N6383, N3441);
and AND4 (N6386, N6371, N246, N808, N5246);
and AND3 (N6387, N6375, N5080, N5101);
or OR2 (N6388, N6386, N1968);
buf BUF1 (N6389, N6382);
and AND3 (N6390, N6374, N125, N816);
and AND3 (N6391, N6369, N3713, N5842);
xor XOR2 (N6392, N6384, N3358);
not NOT1 (N6393, N6388);
nand NAND3 (N6394, N6373, N1288, N809);
or OR3 (N6395, N6391, N2305, N3605);
and AND2 (N6396, N6385, N5603);
buf BUF1 (N6397, N6393);
or OR3 (N6398, N6387, N297, N1096);
nand NAND2 (N6399, N6380, N3936);
nor NOR4 (N6400, N6394, N4478, N1400, N220);
or OR2 (N6401, N6398, N1804);
buf BUF1 (N6402, N6370);
nand NAND4 (N6403, N6401, N2371, N4801, N1681);
xor XOR2 (N6404, N6397, N4537);
xor XOR2 (N6405, N6392, N2790);
or OR3 (N6406, N6400, N5001, N5382);
and AND4 (N6407, N6406, N1885, N2926, N1092);
not NOT1 (N6408, N6389);
and AND4 (N6409, N6390, N6044, N981, N598);
nor NOR3 (N6410, N6408, N1356, N4906);
not NOT1 (N6411, N6403);
buf BUF1 (N6412, N6407);
buf BUF1 (N6413, N6411);
buf BUF1 (N6414, N6395);
xor XOR2 (N6415, N6414, N5968);
xor XOR2 (N6416, N6402, N3043);
not NOT1 (N6417, N6413);
not NOT1 (N6418, N6405);
or OR2 (N6419, N6416, N2389);
not NOT1 (N6420, N6418);
nor NOR4 (N6421, N6410, N3013, N5251, N790);
or OR2 (N6422, N6417, N11);
nor NOR3 (N6423, N6404, N6127, N6407);
not NOT1 (N6424, N6412);
not NOT1 (N6425, N6424);
not NOT1 (N6426, N6409);
nand NAND2 (N6427, N6415, N4560);
xor XOR2 (N6428, N6421, N1558);
nor NOR3 (N6429, N6422, N5786, N3961);
or OR3 (N6430, N6423, N4112, N1459);
and AND2 (N6431, N6430, N210);
and AND3 (N6432, N6425, N2848, N1628);
nand NAND3 (N6433, N6426, N3304, N4388);
or OR3 (N6434, N6432, N4026, N5554);
not NOT1 (N6435, N6429);
xor XOR2 (N6436, N6435, N2214);
nor NOR3 (N6437, N6431, N4702, N3530);
nor NOR4 (N6438, N6420, N2673, N5501, N3934);
nand NAND3 (N6439, N6438, N6415, N4031);
or OR3 (N6440, N6419, N4357, N302);
buf BUF1 (N6441, N6433);
xor XOR2 (N6442, N6396, N3732);
not NOT1 (N6443, N6441);
nand NAND2 (N6444, N6427, N3165);
buf BUF1 (N6445, N6437);
xor XOR2 (N6446, N6439, N1461);
xor XOR2 (N6447, N6445, N3418);
buf BUF1 (N6448, N6434);
nand NAND2 (N6449, N6399, N3816);
nor NOR4 (N6450, N6448, N1711, N5450, N2958);
xor XOR2 (N6451, N6442, N2757);
buf BUF1 (N6452, N6428);
or OR3 (N6453, N6449, N4322, N5920);
and AND2 (N6454, N6446, N3935);
or OR3 (N6455, N6443, N2446, N1028);
and AND3 (N6456, N6447, N1680, N6203);
or OR3 (N6457, N6440, N1424, N554);
or OR2 (N6458, N6456, N5939);
buf BUF1 (N6459, N6453);
xor XOR2 (N6460, N6451, N922);
nor NOR4 (N6461, N6452, N379, N5174, N4680);
not NOT1 (N6462, N6458);
not NOT1 (N6463, N6450);
nor NOR4 (N6464, N6444, N4522, N4102, N3816);
and AND2 (N6465, N6455, N3804);
nand NAND2 (N6466, N6460, N4838);
nand NAND3 (N6467, N6436, N5872, N5504);
buf BUF1 (N6468, N6464);
not NOT1 (N6469, N6463);
not NOT1 (N6470, N6466);
or OR3 (N6471, N6461, N2711, N688);
nand NAND2 (N6472, N6454, N4220);
not NOT1 (N6473, N6457);
not NOT1 (N6474, N6462);
xor XOR2 (N6475, N6472, N5819);
not NOT1 (N6476, N6471);
buf BUF1 (N6477, N6474);
nor NOR4 (N6478, N6475, N5165, N2595, N1771);
and AND3 (N6479, N6477, N1550, N731);
or OR3 (N6480, N6459, N4099, N2217);
xor XOR2 (N6481, N6470, N197);
buf BUF1 (N6482, N6481);
not NOT1 (N6483, N6468);
nand NAND2 (N6484, N6476, N4911);
buf BUF1 (N6485, N6478);
nor NOR3 (N6486, N6465, N5865, N3663);
nor NOR3 (N6487, N6482, N1777, N1393);
and AND3 (N6488, N6485, N3250, N5157);
or OR4 (N6489, N6469, N3454, N4236, N5323);
and AND2 (N6490, N6484, N2122);
buf BUF1 (N6491, N6490);
buf BUF1 (N6492, N6491);
not NOT1 (N6493, N6489);
nand NAND3 (N6494, N6467, N2805, N5436);
nor NOR4 (N6495, N6483, N1573, N255, N3796);
not NOT1 (N6496, N6495);
nor NOR4 (N6497, N6473, N6132, N575, N3278);
xor XOR2 (N6498, N6488, N5742);
and AND4 (N6499, N6486, N5138, N3176, N4001);
not NOT1 (N6500, N6493);
nand NAND2 (N6501, N6480, N3299);
nor NOR2 (N6502, N6497, N2597);
buf BUF1 (N6503, N6501);
not NOT1 (N6504, N6494);
or OR3 (N6505, N6500, N167, N1771);
nand NAND2 (N6506, N6479, N1624);
nand NAND2 (N6507, N6499, N2377);
and AND4 (N6508, N6503, N3723, N6284, N3708);
or OR4 (N6509, N6487, N830, N1545, N249);
not NOT1 (N6510, N6498);
or OR4 (N6511, N6502, N4929, N5497, N3821);
buf BUF1 (N6512, N6511);
xor XOR2 (N6513, N6510, N6108);
nor NOR3 (N6514, N6507, N587, N6436);
nand NAND3 (N6515, N6512, N5996, N3616);
nor NOR3 (N6516, N6513, N5397, N5040);
nand NAND3 (N6517, N6504, N1346, N2803);
or OR3 (N6518, N6514, N1880, N2896);
xor XOR2 (N6519, N6517, N433);
buf BUF1 (N6520, N6518);
xor XOR2 (N6521, N6519, N3625);
nor NOR4 (N6522, N6520, N5734, N3841, N5311);
buf BUF1 (N6523, N6492);
buf BUF1 (N6524, N6505);
or OR4 (N6525, N6523, N3406, N5756, N3655);
buf BUF1 (N6526, N6509);
not NOT1 (N6527, N6524);
nand NAND2 (N6528, N6515, N4567);
xor XOR2 (N6529, N6516, N4653);
nor NOR4 (N6530, N6496, N4179, N2329, N2602);
or OR4 (N6531, N6521, N3315, N335, N2086);
nor NOR3 (N6532, N6526, N671, N1648);
xor XOR2 (N6533, N6530, N4302);
nor NOR3 (N6534, N6533, N1332, N3685);
nor NOR2 (N6535, N6534, N3688);
not NOT1 (N6536, N6535);
buf BUF1 (N6537, N6525);
nand NAND2 (N6538, N6506, N757);
nand NAND2 (N6539, N6532, N3244);
xor XOR2 (N6540, N6531, N4191);
not NOT1 (N6541, N6540);
and AND3 (N6542, N6536, N3834, N4745);
nor NOR4 (N6543, N6542, N4649, N1002, N4629);
buf BUF1 (N6544, N6527);
or OR2 (N6545, N6537, N4209);
not NOT1 (N6546, N6508);
nand NAND4 (N6547, N6546, N1616, N3965, N4233);
nand NAND3 (N6548, N6528, N4116, N5065);
nand NAND4 (N6549, N6522, N2136, N2550, N5041);
nand NAND3 (N6550, N6538, N2946, N1853);
or OR2 (N6551, N6544, N2195);
nand NAND3 (N6552, N6549, N6535, N3705);
nand NAND3 (N6553, N6548, N2495, N6465);
xor XOR2 (N6554, N6547, N4495);
not NOT1 (N6555, N6552);
and AND2 (N6556, N6529, N1882);
and AND4 (N6557, N6541, N1199, N5063, N6252);
and AND4 (N6558, N6557, N3650, N2524, N2757);
nor NOR3 (N6559, N6554, N874, N1886);
or OR4 (N6560, N6545, N5735, N6044, N1877);
and AND2 (N6561, N6543, N583);
nand NAND4 (N6562, N6560, N5677, N1309, N1090);
xor XOR2 (N6563, N6551, N1043);
buf BUF1 (N6564, N6559);
nand NAND2 (N6565, N6555, N5431);
xor XOR2 (N6566, N6558, N1723);
not NOT1 (N6567, N6561);
buf BUF1 (N6568, N6563);
nor NOR3 (N6569, N6567, N1508, N50);
nand NAND2 (N6570, N6550, N3680);
or OR4 (N6571, N6564, N3146, N6271, N5725);
nand NAND4 (N6572, N6562, N3768, N1086, N4486);
or OR3 (N6573, N6556, N2515, N4117);
nor NOR2 (N6574, N6569, N4957);
not NOT1 (N6575, N6568);
nor NOR2 (N6576, N6570, N1158);
not NOT1 (N6577, N6571);
not NOT1 (N6578, N6576);
buf BUF1 (N6579, N6553);
buf BUF1 (N6580, N6565);
not NOT1 (N6581, N6579);
and AND2 (N6582, N6577, N1979);
buf BUF1 (N6583, N6539);
xor XOR2 (N6584, N6578, N4088);
xor XOR2 (N6585, N6566, N1726);
and AND2 (N6586, N6581, N3216);
and AND2 (N6587, N6572, N4063);
xor XOR2 (N6588, N6587, N6587);
buf BUF1 (N6589, N6583);
and AND4 (N6590, N6588, N391, N5098, N550);
or OR2 (N6591, N6590, N2819);
not NOT1 (N6592, N6575);
not NOT1 (N6593, N6584);
nor NOR3 (N6594, N6580, N2747, N4027);
and AND2 (N6595, N6594, N2143);
not NOT1 (N6596, N6593);
not NOT1 (N6597, N6574);
xor XOR2 (N6598, N6582, N3581);
nand NAND3 (N6599, N6592, N1697, N1544);
or OR3 (N6600, N6595, N1936, N4097);
not NOT1 (N6601, N6585);
xor XOR2 (N6602, N6601, N5124);
buf BUF1 (N6603, N6597);
or OR2 (N6604, N6596, N5578);
and AND2 (N6605, N6604, N4500);
nor NOR3 (N6606, N6598, N610, N499);
not NOT1 (N6607, N6605);
buf BUF1 (N6608, N6586);
not NOT1 (N6609, N6606);
buf BUF1 (N6610, N6600);
buf BUF1 (N6611, N6591);
or OR2 (N6612, N6573, N2686);
xor XOR2 (N6613, N6602, N2718);
buf BUF1 (N6614, N6607);
and AND2 (N6615, N6603, N5633);
nor NOR3 (N6616, N6615, N979, N5122);
and AND2 (N6617, N6608, N4428);
or OR4 (N6618, N6599, N3796, N5006, N6209);
or OR4 (N6619, N6613, N6321, N585, N2141);
nand NAND4 (N6620, N6589, N1091, N1465, N6414);
not NOT1 (N6621, N6614);
nand NAND4 (N6622, N6609, N712, N4505, N4401);
and AND3 (N6623, N6611, N3246, N1807);
and AND4 (N6624, N6616, N2993, N1420, N3885);
or OR3 (N6625, N6618, N1500, N717);
buf BUF1 (N6626, N6623);
or OR2 (N6627, N6612, N4073);
buf BUF1 (N6628, N6625);
or OR4 (N6629, N6620, N5477, N1510, N41);
buf BUF1 (N6630, N6626);
nor NOR2 (N6631, N6628, N1038);
not NOT1 (N6632, N6617);
or OR4 (N6633, N6621, N5921, N805, N2980);
xor XOR2 (N6634, N6622, N3620);
and AND2 (N6635, N6624, N2094);
xor XOR2 (N6636, N6629, N259);
nor NOR3 (N6637, N6630, N6264, N6375);
and AND3 (N6638, N6619, N2808, N4432);
or OR4 (N6639, N6633, N281, N784, N3155);
nor NOR4 (N6640, N6637, N1846, N5105, N6000);
not NOT1 (N6641, N6627);
nor NOR2 (N6642, N6610, N6365);
buf BUF1 (N6643, N6636);
not NOT1 (N6644, N6639);
nand NAND4 (N6645, N6642, N1724, N844, N1686);
nor NOR2 (N6646, N6641, N5550);
buf BUF1 (N6647, N6646);
nand NAND2 (N6648, N6632, N234);
buf BUF1 (N6649, N6645);
or OR4 (N6650, N6631, N5757, N62, N3581);
or OR4 (N6651, N6644, N4071, N374, N4068);
or OR3 (N6652, N6651, N2319, N363);
buf BUF1 (N6653, N6652);
nand NAND3 (N6654, N6653, N5131, N4419);
buf BUF1 (N6655, N6640);
buf BUF1 (N6656, N6635);
buf BUF1 (N6657, N6638);
or OR4 (N6658, N6656, N3083, N4452, N2927);
not NOT1 (N6659, N6650);
nor NOR4 (N6660, N6654, N310, N1721, N3291);
buf BUF1 (N6661, N6649);
buf BUF1 (N6662, N6643);
not NOT1 (N6663, N6661);
nand NAND4 (N6664, N6655, N6570, N4257, N6319);
nand NAND4 (N6665, N6659, N6418, N2787, N930);
nor NOR3 (N6666, N6660, N6371, N2606);
or OR2 (N6667, N6665, N6351);
nand NAND3 (N6668, N6658, N5346, N6612);
and AND4 (N6669, N6647, N6311, N3244, N4046);
and AND3 (N6670, N6648, N1851, N3274);
buf BUF1 (N6671, N6666);
nand NAND3 (N6672, N6657, N1815, N3035);
and AND2 (N6673, N6668, N3055);
not NOT1 (N6674, N6664);
nand NAND4 (N6675, N6662, N1939, N226, N3075);
xor XOR2 (N6676, N6634, N5818);
nor NOR4 (N6677, N6667, N4592, N6575, N612);
buf BUF1 (N6678, N6675);
buf BUF1 (N6679, N6676);
and AND3 (N6680, N6672, N18, N3844);
not NOT1 (N6681, N6674);
nand NAND4 (N6682, N6677, N3123, N3103, N2320);
and AND2 (N6683, N6679, N2790);
nand NAND2 (N6684, N6681, N528);
xor XOR2 (N6685, N6678, N3616);
or OR3 (N6686, N6680, N4147, N2299);
buf BUF1 (N6687, N6669);
nor NOR4 (N6688, N6670, N710, N1854, N1433);
or OR3 (N6689, N6683, N1313, N4355);
nor NOR2 (N6690, N6687, N4146);
nand NAND2 (N6691, N6686, N6489);
not NOT1 (N6692, N6684);
xor XOR2 (N6693, N6663, N2624);
buf BUF1 (N6694, N6692);
not NOT1 (N6695, N6689);
not NOT1 (N6696, N6682);
nor NOR3 (N6697, N6694, N1736, N6303);
xor XOR2 (N6698, N6690, N1226);
not NOT1 (N6699, N6685);
not NOT1 (N6700, N6671);
or OR4 (N6701, N6699, N4360, N426, N1389);
xor XOR2 (N6702, N6700, N2213);
nor NOR3 (N6703, N6701, N6245, N6590);
not NOT1 (N6704, N6691);
xor XOR2 (N6705, N6695, N2547);
not NOT1 (N6706, N6702);
nor NOR3 (N6707, N6704, N1850, N3806);
and AND3 (N6708, N6688, N2257, N3340);
nand NAND3 (N6709, N6673, N2740, N1099);
or OR3 (N6710, N6697, N1641, N1110);
xor XOR2 (N6711, N6703, N205);
nor NOR2 (N6712, N6705, N2943);
nor NOR4 (N6713, N6706, N791, N5824, N6619);
xor XOR2 (N6714, N6710, N880);
nand NAND3 (N6715, N6693, N4655, N1614);
xor XOR2 (N6716, N6712, N5244);
nor NOR4 (N6717, N6711, N3769, N5060, N4348);
nor NOR2 (N6718, N6707, N6638);
not NOT1 (N6719, N6698);
xor XOR2 (N6720, N6709, N6243);
buf BUF1 (N6721, N6713);
buf BUF1 (N6722, N6715);
and AND3 (N6723, N6708, N2321, N947);
or OR2 (N6724, N6723, N3394);
buf BUF1 (N6725, N6718);
xor XOR2 (N6726, N6720, N4392);
nor NOR4 (N6727, N6716, N1007, N3731, N1016);
nand NAND4 (N6728, N6714, N3937, N1239, N5422);
buf BUF1 (N6729, N6722);
nor NOR2 (N6730, N6727, N4543);
or OR4 (N6731, N6725, N958, N214, N4564);
or OR4 (N6732, N6717, N2551, N2899, N6430);
not NOT1 (N6733, N6732);
xor XOR2 (N6734, N6731, N2365);
buf BUF1 (N6735, N6728);
and AND4 (N6736, N6733, N3018, N2639, N4669);
or OR2 (N6737, N6696, N6263);
nand NAND3 (N6738, N6726, N1384, N893);
nor NOR2 (N6739, N6737, N5426);
nor NOR3 (N6740, N6719, N1543, N5588);
nor NOR2 (N6741, N6735, N4471);
and AND4 (N6742, N6734, N993, N1251, N1622);
not NOT1 (N6743, N6724);
or OR3 (N6744, N6740, N6392, N556);
and AND2 (N6745, N6743, N5537);
xor XOR2 (N6746, N6736, N4565);
and AND2 (N6747, N6730, N4046);
nor NOR4 (N6748, N6742, N1287, N5393, N2661);
xor XOR2 (N6749, N6746, N3983);
buf BUF1 (N6750, N6739);
buf BUF1 (N6751, N6750);
nand NAND3 (N6752, N6748, N2444, N5869);
xor XOR2 (N6753, N6721, N2904);
and AND4 (N6754, N6744, N6027, N1324, N1264);
nand NAND3 (N6755, N6754, N154, N5429);
nor NOR2 (N6756, N6729, N777);
xor XOR2 (N6757, N6755, N4116);
xor XOR2 (N6758, N6741, N1922);
or OR3 (N6759, N6751, N4338, N4631);
nor NOR2 (N6760, N6756, N3435);
buf BUF1 (N6761, N6758);
not NOT1 (N6762, N6757);
or OR2 (N6763, N6760, N6607);
or OR3 (N6764, N6747, N897, N6285);
and AND3 (N6765, N6764, N6069, N6356);
or OR3 (N6766, N6738, N846, N4337);
not NOT1 (N6767, N6759);
buf BUF1 (N6768, N6761);
buf BUF1 (N6769, N6753);
and AND2 (N6770, N6767, N1062);
and AND2 (N6771, N6745, N6313);
xor XOR2 (N6772, N6766, N539);
not NOT1 (N6773, N6772);
not NOT1 (N6774, N6771);
and AND4 (N6775, N6773, N4695, N4108, N783);
buf BUF1 (N6776, N6774);
and AND4 (N6777, N6752, N1049, N2643, N3180);
not NOT1 (N6778, N6769);
xor XOR2 (N6779, N6770, N2841);
or OR2 (N6780, N6775, N6460);
xor XOR2 (N6781, N6778, N3560);
not NOT1 (N6782, N6777);
nor NOR2 (N6783, N6765, N6324);
nand NAND4 (N6784, N6776, N1975, N532, N20);
not NOT1 (N6785, N6768);
nor NOR3 (N6786, N6782, N608, N2093);
or OR4 (N6787, N6780, N5113, N6292, N4330);
or OR3 (N6788, N6781, N2275, N2732);
and AND3 (N6789, N6762, N813, N2308);
not NOT1 (N6790, N6789);
not NOT1 (N6791, N6787);
nand NAND2 (N6792, N6786, N2000);
xor XOR2 (N6793, N6788, N4957);
or OR2 (N6794, N6791, N3212);
nor NOR4 (N6795, N6779, N1878, N933, N6160);
buf BUF1 (N6796, N6790);
nor NOR4 (N6797, N6785, N4900, N5864, N2602);
buf BUF1 (N6798, N6784);
nor NOR2 (N6799, N6792, N1829);
and AND3 (N6800, N6797, N2629, N609);
not NOT1 (N6801, N6794);
and AND2 (N6802, N6795, N4806);
or OR2 (N6803, N6793, N2122);
nand NAND3 (N6804, N6796, N1322, N1893);
xor XOR2 (N6805, N6763, N5902);
xor XOR2 (N6806, N6798, N1197);
xor XOR2 (N6807, N6804, N2041);
buf BUF1 (N6808, N6801);
or OR4 (N6809, N6803, N404, N3424, N3715);
xor XOR2 (N6810, N6809, N6450);
nand NAND2 (N6811, N6810, N906);
or OR3 (N6812, N6808, N4321, N1931);
buf BUF1 (N6813, N6802);
or OR2 (N6814, N6811, N5000);
xor XOR2 (N6815, N6814, N2682);
and AND2 (N6816, N6783, N2101);
nand NAND4 (N6817, N6800, N1767, N1407, N3629);
buf BUF1 (N6818, N6807);
nand NAND4 (N6819, N6817, N3631, N5828, N1925);
xor XOR2 (N6820, N6818, N5710);
or OR4 (N6821, N6812, N2095, N6177, N3859);
xor XOR2 (N6822, N6799, N3804);
nand NAND4 (N6823, N6815, N6604, N700, N3335);
not NOT1 (N6824, N6820);
xor XOR2 (N6825, N6816, N2032);
xor XOR2 (N6826, N6824, N1033);
not NOT1 (N6827, N6819);
or OR3 (N6828, N6827, N1458, N4384);
not NOT1 (N6829, N6826);
xor XOR2 (N6830, N6823, N763);
xor XOR2 (N6831, N6822, N4447);
not NOT1 (N6832, N6805);
nor NOR2 (N6833, N6832, N4142);
nand NAND2 (N6834, N6828, N2313);
xor XOR2 (N6835, N6806, N6024);
nand NAND2 (N6836, N6829, N2602);
and AND2 (N6837, N6835, N6309);
and AND2 (N6838, N6830, N5488);
not NOT1 (N6839, N6834);
and AND4 (N6840, N6837, N1069, N271, N3432);
not NOT1 (N6841, N6825);
buf BUF1 (N6842, N6821);
nand NAND3 (N6843, N6840, N541, N2945);
nor NOR3 (N6844, N6842, N2137, N1475);
or OR4 (N6845, N6833, N59, N1174, N3238);
xor XOR2 (N6846, N6838, N1571);
not NOT1 (N6847, N6749);
not NOT1 (N6848, N6844);
nand NAND3 (N6849, N6843, N6364, N3460);
xor XOR2 (N6850, N6841, N271);
not NOT1 (N6851, N6846);
nand NAND3 (N6852, N6847, N5478, N2005);
and AND3 (N6853, N6813, N3209, N5223);
buf BUF1 (N6854, N6850);
xor XOR2 (N6855, N6854, N5730);
not NOT1 (N6856, N6836);
buf BUF1 (N6857, N6856);
and AND4 (N6858, N6839, N1650, N17, N5211);
and AND4 (N6859, N6848, N4241, N3878, N3099);
xor XOR2 (N6860, N6857, N4075);
nand NAND2 (N6861, N6853, N4043);
not NOT1 (N6862, N6855);
nor NOR4 (N6863, N6859, N5688, N2063, N3638);
nand NAND4 (N6864, N6863, N5236, N5706, N6321);
buf BUF1 (N6865, N6862);
nand NAND4 (N6866, N6860, N5950, N6391, N2925);
or OR3 (N6867, N6845, N344, N1105);
and AND4 (N6868, N6851, N507, N479, N2917);
not NOT1 (N6869, N6866);
nand NAND4 (N6870, N6868, N1773, N5517, N5077);
not NOT1 (N6871, N6865);
and AND2 (N6872, N6870, N626);
and AND4 (N6873, N6867, N4957, N1654, N5435);
xor XOR2 (N6874, N6869, N6448);
and AND2 (N6875, N6871, N2901);
nand NAND3 (N6876, N6849, N3992, N2950);
nand NAND4 (N6877, N6864, N3926, N6817, N5885);
xor XOR2 (N6878, N6876, N734);
buf BUF1 (N6879, N6877);
and AND3 (N6880, N6858, N4328, N6582);
or OR2 (N6881, N6879, N4620);
and AND2 (N6882, N6831, N1912);
not NOT1 (N6883, N6882);
nor NOR2 (N6884, N6861, N6742);
not NOT1 (N6885, N6878);
nor NOR4 (N6886, N6875, N5575, N6229, N481);
xor XOR2 (N6887, N6881, N149);
not NOT1 (N6888, N6884);
xor XOR2 (N6889, N6885, N4188);
not NOT1 (N6890, N6874);
and AND3 (N6891, N6888, N3610, N1633);
not NOT1 (N6892, N6889);
xor XOR2 (N6893, N6891, N1735);
nand NAND3 (N6894, N6887, N5154, N4303);
nor NOR4 (N6895, N6894, N6112, N3187, N4859);
buf BUF1 (N6896, N6873);
nor NOR4 (N6897, N6893, N2676, N2050, N6167);
nor NOR4 (N6898, N6892, N4072, N1971, N4283);
or OR3 (N6899, N6886, N3281, N4568);
buf BUF1 (N6900, N6883);
or OR4 (N6901, N6899, N5260, N110, N6160);
nor NOR3 (N6902, N6852, N975, N1841);
nand NAND3 (N6903, N6890, N3604, N4833);
and AND4 (N6904, N6902, N3661, N4937, N3054);
nand NAND4 (N6905, N6872, N1137, N6102, N5075);
nand NAND3 (N6906, N6905, N6864, N2855);
xor XOR2 (N6907, N6901, N6504);
xor XOR2 (N6908, N6907, N1611);
not NOT1 (N6909, N6898);
not NOT1 (N6910, N6880);
buf BUF1 (N6911, N6904);
nand NAND2 (N6912, N6903, N927);
buf BUF1 (N6913, N6895);
nand NAND2 (N6914, N6911, N2719);
or OR2 (N6915, N6906, N3253);
not NOT1 (N6916, N6897);
xor XOR2 (N6917, N6914, N3696);
and AND4 (N6918, N6908, N5333, N5893, N417);
and AND3 (N6919, N6918, N2595, N86);
nor NOR3 (N6920, N6916, N5992, N1919);
buf BUF1 (N6921, N6910);
or OR4 (N6922, N6921, N3434, N5632, N1674);
not NOT1 (N6923, N6922);
not NOT1 (N6924, N6915);
not NOT1 (N6925, N6909);
nor NOR2 (N6926, N6913, N1334);
or OR4 (N6927, N6900, N3374, N598, N3361);
nand NAND2 (N6928, N6919, N6536);
buf BUF1 (N6929, N6927);
and AND2 (N6930, N6923, N2380);
not NOT1 (N6931, N6926);
nor NOR3 (N6932, N6924, N2939, N3367);
and AND2 (N6933, N6932, N802);
nor NOR4 (N6934, N6920, N1007, N6927, N4739);
nor NOR3 (N6935, N6931, N1132, N6639);
nor NOR4 (N6936, N6912, N2677, N6266, N1093);
and AND2 (N6937, N6896, N5375);
or OR3 (N6938, N6928, N2209, N1560);
not NOT1 (N6939, N6933);
not NOT1 (N6940, N6935);
and AND2 (N6941, N6936, N1988);
nor NOR4 (N6942, N6939, N593, N2101, N1659);
and AND3 (N6943, N6929, N2017, N4058);
xor XOR2 (N6944, N6937, N392);
nand NAND3 (N6945, N6941, N3430, N4696);
not NOT1 (N6946, N6943);
nor NOR3 (N6947, N6938, N5628, N6796);
not NOT1 (N6948, N6947);
nor NOR2 (N6949, N6944, N6406);
or OR2 (N6950, N6942, N1758);
nand NAND2 (N6951, N6930, N2941);
xor XOR2 (N6952, N6917, N2150);
nor NOR3 (N6953, N6950, N3206, N5489);
xor XOR2 (N6954, N6925, N1583);
not NOT1 (N6955, N6949);
and AND4 (N6956, N6953, N4425, N2455, N330);
not NOT1 (N6957, N6951);
nor NOR3 (N6958, N6940, N1368, N110);
buf BUF1 (N6959, N6934);
nor NOR4 (N6960, N6957, N3617, N6392, N5426);
or OR2 (N6961, N6958, N5641);
or OR3 (N6962, N6945, N862, N3206);
buf BUF1 (N6963, N6955);
nor NOR4 (N6964, N6946, N1906, N2618, N6454);
nand NAND3 (N6965, N6964, N5434, N5801);
xor XOR2 (N6966, N6961, N3253);
and AND2 (N6967, N6956, N4321);
nand NAND2 (N6968, N6954, N6696);
nand NAND2 (N6969, N6960, N6623);
nand NAND2 (N6970, N6968, N6749);
buf BUF1 (N6971, N6967);
not NOT1 (N6972, N6962);
nor NOR3 (N6973, N6948, N5561, N2390);
or OR3 (N6974, N6970, N6743, N3427);
buf BUF1 (N6975, N6965);
or OR2 (N6976, N6974, N2787);
xor XOR2 (N6977, N6972, N1289);
not NOT1 (N6978, N6969);
or OR2 (N6979, N6973, N742);
nor NOR2 (N6980, N6952, N2103);
nor NOR2 (N6981, N6966, N802);
not NOT1 (N6982, N6977);
buf BUF1 (N6983, N6978);
nand NAND3 (N6984, N6959, N1760, N6755);
nand NAND3 (N6985, N6982, N3024, N6513);
and AND4 (N6986, N6983, N1808, N5029, N6727);
not NOT1 (N6987, N6975);
or OR4 (N6988, N6963, N2192, N3821, N633);
nand NAND3 (N6989, N6985, N1207, N6923);
buf BUF1 (N6990, N6984);
nor NOR3 (N6991, N6981, N6390, N3757);
not NOT1 (N6992, N6988);
not NOT1 (N6993, N6991);
nor NOR3 (N6994, N6992, N6838, N3664);
nand NAND2 (N6995, N6989, N6504);
buf BUF1 (N6996, N6987);
not NOT1 (N6997, N6976);
xor XOR2 (N6998, N6995, N936);
and AND3 (N6999, N6996, N2632, N272);
xor XOR2 (N7000, N6971, N2956);
nand NAND2 (N7001, N6980, N645);
nand NAND2 (N7002, N7000, N4070);
nand NAND4 (N7003, N6979, N4460, N179, N685);
or OR2 (N7004, N6986, N2805);
or OR3 (N7005, N7002, N2763, N2089);
nand NAND4 (N7006, N6994, N2932, N4845, N1074);
buf BUF1 (N7007, N7004);
not NOT1 (N7008, N7007);
buf BUF1 (N7009, N7006);
and AND3 (N7010, N6998, N5197, N1861);
nor NOR4 (N7011, N7001, N639, N2654, N308);
nor NOR3 (N7012, N7003, N1608, N861);
or OR2 (N7013, N7009, N4149);
not NOT1 (N7014, N6997);
and AND2 (N7015, N7012, N3294);
xor XOR2 (N7016, N6993, N4335);
buf BUF1 (N7017, N6999);
nor NOR3 (N7018, N7011, N4664, N5562);
nand NAND3 (N7019, N7017, N2430, N3699);
and AND4 (N7020, N7005, N1574, N5401, N4627);
or OR2 (N7021, N6990, N4269);
nand NAND2 (N7022, N7010, N3257);
and AND4 (N7023, N7013, N3229, N1777, N1326);
buf BUF1 (N7024, N7014);
nor NOR3 (N7025, N7022, N2452, N5304);
xor XOR2 (N7026, N7019, N1870);
or OR3 (N7027, N7008, N2484, N6926);
nor NOR2 (N7028, N7015, N6309);
buf BUF1 (N7029, N7028);
and AND3 (N7030, N7016, N1834, N4514);
xor XOR2 (N7031, N7027, N1009);
buf BUF1 (N7032, N7021);
not NOT1 (N7033, N7026);
xor XOR2 (N7034, N7033, N3698);
or OR2 (N7035, N7024, N3018);
and AND4 (N7036, N7034, N961, N3660, N2251);
buf BUF1 (N7037, N7018);
and AND3 (N7038, N7029, N1336, N4272);
xor XOR2 (N7039, N7038, N3767);
nand NAND2 (N7040, N7035, N4166);
xor XOR2 (N7041, N7020, N5346);
nor NOR2 (N7042, N7023, N4733);
xor XOR2 (N7043, N7041, N5234);
and AND2 (N7044, N7030, N3342);
or OR2 (N7045, N7043, N1232);
xor XOR2 (N7046, N7042, N221);
nand NAND4 (N7047, N7031, N5780, N2415, N2591);
not NOT1 (N7048, N7046);
nand NAND4 (N7049, N7036, N5685, N5412, N1345);
and AND2 (N7050, N7047, N2996);
nor NOR3 (N7051, N7050, N187, N1347);
and AND4 (N7052, N7049, N2700, N3736, N1359);
not NOT1 (N7053, N7040);
xor XOR2 (N7054, N7048, N6649);
and AND4 (N7055, N7052, N4221, N3709, N6251);
and AND2 (N7056, N7032, N6251);
and AND2 (N7057, N7037, N3672);
and AND4 (N7058, N7054, N3220, N6803, N6615);
not NOT1 (N7059, N7045);
not NOT1 (N7060, N7058);
and AND3 (N7061, N7051, N5455, N927);
xor XOR2 (N7062, N7025, N5148);
and AND4 (N7063, N7057, N1362, N251, N255);
and AND3 (N7064, N7063, N2002, N6707);
nand NAND2 (N7065, N7056, N4272);
nor NOR4 (N7066, N7060, N277, N1085, N2720);
not NOT1 (N7067, N7066);
buf BUF1 (N7068, N7053);
or OR4 (N7069, N7044, N4249, N1299, N1586);
nand NAND2 (N7070, N7059, N3470);
nor NOR4 (N7071, N7068, N3690, N5989, N3426);
buf BUF1 (N7072, N7039);
or OR4 (N7073, N7062, N1063, N4077, N5956);
nor NOR3 (N7074, N7064, N1335, N744);
or OR4 (N7075, N7065, N3445, N3188, N434);
not NOT1 (N7076, N7072);
nor NOR3 (N7077, N7061, N257, N5638);
nand NAND2 (N7078, N7075, N4096);
and AND4 (N7079, N7077, N6290, N2192, N5603);
xor XOR2 (N7080, N7076, N2007);
nor NOR4 (N7081, N7070, N4584, N3515, N3169);
not NOT1 (N7082, N7067);
nor NOR4 (N7083, N7081, N2633, N2042, N38);
or OR3 (N7084, N7071, N5026, N6842);
nor NOR2 (N7085, N7069, N309);
buf BUF1 (N7086, N7055);
buf BUF1 (N7087, N7079);
buf BUF1 (N7088, N7080);
or OR4 (N7089, N7073, N6921, N4206, N1521);
buf BUF1 (N7090, N7086);
and AND2 (N7091, N7078, N5291);
nand NAND2 (N7092, N7074, N1959);
or OR2 (N7093, N7083, N4573);
and AND4 (N7094, N7082, N1409, N3141, N5504);
nor NOR2 (N7095, N7094, N3655);
nand NAND3 (N7096, N7087, N2447, N3276);
xor XOR2 (N7097, N7093, N4038);
xor XOR2 (N7098, N7091, N1689);
nor NOR3 (N7099, N7085, N1875, N1218);
not NOT1 (N7100, N7088);
nor NOR4 (N7101, N7100, N744, N2436, N4016);
xor XOR2 (N7102, N7089, N5938);
xor XOR2 (N7103, N7084, N2888);
or OR2 (N7104, N7098, N4466);
and AND2 (N7105, N7096, N2674);
or OR2 (N7106, N7097, N1037);
not NOT1 (N7107, N7105);
not NOT1 (N7108, N7095);
xor XOR2 (N7109, N7099, N1367);
not NOT1 (N7110, N7103);
nand NAND3 (N7111, N7102, N2211, N4608);
nor NOR4 (N7112, N7104, N1849, N3587, N1676);
buf BUF1 (N7113, N7090);
nor NOR2 (N7114, N7101, N6102);
nor NOR2 (N7115, N7107, N2714);
not NOT1 (N7116, N7114);
nor NOR4 (N7117, N7111, N5252, N3612, N4202);
nor NOR3 (N7118, N7106, N6792, N1209);
not NOT1 (N7119, N7116);
nor NOR3 (N7120, N7119, N2465, N4085);
and AND4 (N7121, N7108, N3149, N5837, N2807);
nand NAND4 (N7122, N7117, N718, N5122, N4575);
nor NOR3 (N7123, N7092, N6533, N1804);
xor XOR2 (N7124, N7112, N1214);
buf BUF1 (N7125, N7122);
buf BUF1 (N7126, N7115);
nand NAND4 (N7127, N7125, N4315, N4237, N2726);
nand NAND3 (N7128, N7110, N5500, N1980);
xor XOR2 (N7129, N7128, N1442);
buf BUF1 (N7130, N7124);
or OR2 (N7131, N7123, N4598);
not NOT1 (N7132, N7121);
not NOT1 (N7133, N7126);
and AND3 (N7134, N7120, N1940, N1495);
and AND3 (N7135, N7109, N5295, N1041);
and AND3 (N7136, N7135, N184, N6604);
not NOT1 (N7137, N7127);
xor XOR2 (N7138, N7137, N141);
xor XOR2 (N7139, N7133, N2273);
not NOT1 (N7140, N7113);
xor XOR2 (N7141, N7139, N5363);
nor NOR4 (N7142, N7131, N2696, N3326, N2524);
nor NOR2 (N7143, N7134, N2836);
or OR4 (N7144, N7129, N1430, N2798, N4236);
not NOT1 (N7145, N7140);
xor XOR2 (N7146, N7136, N1814);
nand NAND3 (N7147, N7132, N4953, N1367);
xor XOR2 (N7148, N7146, N3159);
or OR2 (N7149, N7118, N1021);
xor XOR2 (N7150, N7142, N896);
and AND3 (N7151, N7138, N5282, N6910);
xor XOR2 (N7152, N7143, N1298);
and AND2 (N7153, N7151, N2963);
or OR2 (N7154, N7141, N262);
or OR4 (N7155, N7145, N4865, N2089, N3754);
nand NAND2 (N7156, N7149, N6572);
and AND4 (N7157, N7144, N6132, N1787, N3902);
nor NOR3 (N7158, N7153, N5483, N3115);
nor NOR3 (N7159, N7152, N5045, N4214);
not NOT1 (N7160, N7154);
nor NOR3 (N7161, N7157, N5251, N5987);
not NOT1 (N7162, N7158);
nand NAND2 (N7163, N7148, N1451);
not NOT1 (N7164, N7147);
nor NOR2 (N7165, N7155, N323);
nor NOR4 (N7166, N7150, N1887, N374, N2734);
and AND2 (N7167, N7130, N6871);
nor NOR3 (N7168, N7156, N4637, N6133);
nand NAND4 (N7169, N7165, N639, N509, N5889);
or OR4 (N7170, N7167, N1060, N324, N7106);
or OR2 (N7171, N7164, N3048);
nand NAND2 (N7172, N7163, N1634);
xor XOR2 (N7173, N7171, N4371);
nor NOR2 (N7174, N7172, N106);
or OR4 (N7175, N7173, N5326, N6241, N5423);
and AND4 (N7176, N7175, N2054, N5007, N4299);
and AND4 (N7177, N7161, N6661, N5650, N5010);
nand NAND3 (N7178, N7166, N2555, N198);
and AND3 (N7179, N7170, N512, N1509);
or OR3 (N7180, N7179, N1672, N6290);
buf BUF1 (N7181, N7162);
nor NOR4 (N7182, N7169, N6835, N172, N2724);
xor XOR2 (N7183, N7182, N6066);
and AND4 (N7184, N7181, N3701, N3331, N432);
nor NOR3 (N7185, N7180, N1360, N372);
buf BUF1 (N7186, N7178);
not NOT1 (N7187, N7183);
nor NOR4 (N7188, N7168, N5103, N1468, N5643);
and AND4 (N7189, N7187, N1941, N2196, N1582);
and AND4 (N7190, N7176, N4603, N6837, N5352);
buf BUF1 (N7191, N7190);
nand NAND4 (N7192, N7177, N5855, N5703, N1601);
or OR2 (N7193, N7185, N282);
xor XOR2 (N7194, N7186, N4835);
not NOT1 (N7195, N7194);
nand NAND2 (N7196, N7189, N2897);
nor NOR2 (N7197, N7159, N5556);
not NOT1 (N7198, N7196);
xor XOR2 (N7199, N7193, N6705);
xor XOR2 (N7200, N7174, N2063);
and AND4 (N7201, N7199, N6797, N2979, N101);
nor NOR3 (N7202, N7198, N5161, N1206);
or OR4 (N7203, N7202, N5, N5837, N5773);
nor NOR2 (N7204, N7184, N6070);
not NOT1 (N7205, N7160);
not NOT1 (N7206, N7201);
buf BUF1 (N7207, N7195);
nand NAND3 (N7208, N7207, N3205, N952);
nor NOR2 (N7209, N7197, N4851);
and AND3 (N7210, N7203, N5860, N6883);
buf BUF1 (N7211, N7205);
nand NAND4 (N7212, N7200, N2779, N5255, N6558);
not NOT1 (N7213, N7191);
or OR3 (N7214, N7206, N2127, N5783);
nor NOR2 (N7215, N7213, N5957);
xor XOR2 (N7216, N7204, N3403);
and AND3 (N7217, N7215, N5392, N1420);
nor NOR2 (N7218, N7211, N3755);
buf BUF1 (N7219, N7212);
xor XOR2 (N7220, N7209, N3414);
not NOT1 (N7221, N7216);
xor XOR2 (N7222, N7217, N4504);
nor NOR2 (N7223, N7222, N3531);
xor XOR2 (N7224, N7220, N6893);
buf BUF1 (N7225, N7219);
nor NOR4 (N7226, N7214, N6127, N5185, N5995);
not NOT1 (N7227, N7221);
and AND2 (N7228, N7227, N5919);
nand NAND2 (N7229, N7225, N143);
buf BUF1 (N7230, N7229);
not NOT1 (N7231, N7226);
or OR4 (N7232, N7210, N3709, N4888, N4233);
buf BUF1 (N7233, N7231);
nor NOR4 (N7234, N7218, N2799, N3448, N4856);
xor XOR2 (N7235, N7223, N3738);
xor XOR2 (N7236, N7233, N4032);
and AND4 (N7237, N7188, N4354, N5495, N703);
or OR4 (N7238, N7192, N1618, N421, N6114);
nor NOR3 (N7239, N7208, N5050, N1167);
buf BUF1 (N7240, N7228);
or OR2 (N7241, N7240, N2226);
not NOT1 (N7242, N7238);
nor NOR3 (N7243, N7239, N5583, N5356);
or OR4 (N7244, N7243, N5664, N2462, N1320);
not NOT1 (N7245, N7235);
or OR4 (N7246, N7232, N1825, N3786, N1411);
nand NAND3 (N7247, N7246, N2232, N5109);
buf BUF1 (N7248, N7244);
or OR3 (N7249, N7248, N6554, N2582);
and AND4 (N7250, N7247, N3397, N89, N733);
buf BUF1 (N7251, N7241);
buf BUF1 (N7252, N7236);
and AND4 (N7253, N7252, N5938, N2427, N7156);
and AND4 (N7254, N7234, N3959, N6739, N6517);
or OR3 (N7255, N7254, N2934, N5675);
xor XOR2 (N7256, N7253, N1445);
not NOT1 (N7257, N7245);
or OR3 (N7258, N7242, N3151, N651);
not NOT1 (N7259, N7258);
nand NAND4 (N7260, N7249, N4433, N5278, N2729);
nor NOR2 (N7261, N7250, N6223);
and AND3 (N7262, N7230, N2782, N2491);
or OR4 (N7263, N7260, N4681, N2410, N4092);
not NOT1 (N7264, N7237);
not NOT1 (N7265, N7261);
or OR3 (N7266, N7257, N5565, N1883);
buf BUF1 (N7267, N7259);
and AND4 (N7268, N7267, N1280, N3323, N4948);
nand NAND3 (N7269, N7268, N4336, N3389);
or OR2 (N7270, N7256, N5763);
and AND2 (N7271, N7264, N1589);
not NOT1 (N7272, N7271);
buf BUF1 (N7273, N7251);
or OR2 (N7274, N7270, N3491);
xor XOR2 (N7275, N7266, N1479);
not NOT1 (N7276, N7224);
and AND3 (N7277, N7274, N143, N1925);
nor NOR4 (N7278, N7255, N2668, N140, N4248);
not NOT1 (N7279, N7273);
or OR4 (N7280, N7279, N727, N5282, N1933);
and AND3 (N7281, N7277, N4271, N184);
xor XOR2 (N7282, N7272, N3339);
xor XOR2 (N7283, N7280, N983);
not NOT1 (N7284, N7265);
or OR4 (N7285, N7262, N4396, N1797, N4012);
or OR2 (N7286, N7283, N7211);
not NOT1 (N7287, N7285);
buf BUF1 (N7288, N7278);
or OR4 (N7289, N7276, N5404, N4685, N7091);
not NOT1 (N7290, N7284);
or OR4 (N7291, N7286, N6005, N3809, N3802);
xor XOR2 (N7292, N7290, N1238);
and AND2 (N7293, N7282, N3008);
and AND3 (N7294, N7288, N6045, N5693);
nand NAND4 (N7295, N7292, N134, N4013, N2345);
buf BUF1 (N7296, N7281);
nand NAND4 (N7297, N7275, N5133, N4767, N29);
and AND3 (N7298, N7295, N3757, N1313);
or OR4 (N7299, N7289, N4564, N7246, N4011);
nand NAND4 (N7300, N7297, N2832, N2761, N3587);
nand NAND4 (N7301, N7263, N1970, N2843, N4922);
and AND2 (N7302, N7294, N5518);
and AND4 (N7303, N7298, N3436, N1856, N5778);
nor NOR4 (N7304, N7296, N4399, N6503, N6775);
nor NOR4 (N7305, N7287, N2210, N6188, N4454);
buf BUF1 (N7306, N7303);
not NOT1 (N7307, N7269);
and AND4 (N7308, N7301, N5974, N6920, N426);
xor XOR2 (N7309, N7299, N6439);
not NOT1 (N7310, N7300);
nand NAND2 (N7311, N7302, N3624);
buf BUF1 (N7312, N7305);
not NOT1 (N7313, N7308);
nand NAND2 (N7314, N7313, N6245);
xor XOR2 (N7315, N7291, N5412);
buf BUF1 (N7316, N7304);
xor XOR2 (N7317, N7311, N941);
and AND2 (N7318, N7315, N915);
nand NAND3 (N7319, N7318, N1691, N1181);
buf BUF1 (N7320, N7317);
nand NAND4 (N7321, N7312, N4189, N4149, N6120);
buf BUF1 (N7322, N7320);
nor NOR2 (N7323, N7316, N1564);
nor NOR4 (N7324, N7306, N4068, N2212, N655);
or OR4 (N7325, N7293, N1329, N5591, N5123);
nand NAND4 (N7326, N7309, N4207, N2773, N6165);
or OR3 (N7327, N7326, N6406, N3687);
not NOT1 (N7328, N7307);
not NOT1 (N7329, N7325);
nor NOR3 (N7330, N7324, N6789, N5606);
nor NOR4 (N7331, N7319, N5988, N2764, N5221);
nor NOR4 (N7332, N7329, N2933, N1311, N4500);
buf BUF1 (N7333, N7332);
or OR4 (N7334, N7322, N1857, N6945, N3007);
buf BUF1 (N7335, N7330);
nor NOR4 (N7336, N7333, N3001, N6319, N961);
or OR2 (N7337, N7334, N1985);
buf BUF1 (N7338, N7337);
or OR2 (N7339, N7321, N3268);
nand NAND3 (N7340, N7328, N3482, N3744);
nand NAND4 (N7341, N7310, N5058, N501, N862);
not NOT1 (N7342, N7340);
xor XOR2 (N7343, N7314, N1776);
or OR4 (N7344, N7323, N4723, N1536, N6713);
nor NOR3 (N7345, N7331, N3664, N4367);
or OR3 (N7346, N7338, N365, N3103);
buf BUF1 (N7347, N7327);
not NOT1 (N7348, N7346);
buf BUF1 (N7349, N7335);
xor XOR2 (N7350, N7345, N4256);
xor XOR2 (N7351, N7347, N7018);
not NOT1 (N7352, N7336);
buf BUF1 (N7353, N7351);
nor NOR3 (N7354, N7342, N1062, N5854);
nor NOR3 (N7355, N7354, N6283, N2196);
and AND3 (N7356, N7339, N5114, N1134);
or OR4 (N7357, N7344, N6401, N244, N2575);
or OR2 (N7358, N7343, N2241);
or OR2 (N7359, N7357, N1299);
or OR2 (N7360, N7358, N7167);
buf BUF1 (N7361, N7353);
or OR4 (N7362, N7348, N6580, N2407, N4723);
buf BUF1 (N7363, N7356);
buf BUF1 (N7364, N7355);
xor XOR2 (N7365, N7363, N5578);
buf BUF1 (N7366, N7365);
or OR3 (N7367, N7350, N3936, N5004);
and AND2 (N7368, N7349, N5863);
nor NOR2 (N7369, N7341, N6612);
xor XOR2 (N7370, N7359, N2005);
nor NOR4 (N7371, N7370, N4209, N2800, N3088);
buf BUF1 (N7372, N7364);
nor NOR3 (N7373, N7368, N419, N5378);
xor XOR2 (N7374, N7373, N4641);
and AND4 (N7375, N7361, N2895, N5522, N1428);
xor XOR2 (N7376, N7362, N3682);
or OR2 (N7377, N7352, N5497);
and AND3 (N7378, N7366, N4908, N5620);
xor XOR2 (N7379, N7371, N6709);
xor XOR2 (N7380, N7378, N3524);
buf BUF1 (N7381, N7380);
nand NAND4 (N7382, N7379, N1445, N898, N4528);
nand NAND4 (N7383, N7382, N6622, N350, N3486);
nand NAND2 (N7384, N7372, N3260);
xor XOR2 (N7385, N7376, N2913);
and AND2 (N7386, N7384, N6550);
buf BUF1 (N7387, N7367);
buf BUF1 (N7388, N7375);
not NOT1 (N7389, N7374);
xor XOR2 (N7390, N7387, N1675);
nor NOR2 (N7391, N7390, N7345);
not NOT1 (N7392, N7377);
buf BUF1 (N7393, N7385);
or OR2 (N7394, N7393, N4733);
nand NAND2 (N7395, N7381, N4857);
not NOT1 (N7396, N7391);
or OR2 (N7397, N7386, N3851);
not NOT1 (N7398, N7392);
buf BUF1 (N7399, N7369);
nand NAND4 (N7400, N7396, N4750, N5912, N3027);
nand NAND3 (N7401, N7389, N6754, N7051);
nor NOR4 (N7402, N7398, N6429, N1075, N2882);
not NOT1 (N7403, N7383);
buf BUF1 (N7404, N7403);
xor XOR2 (N7405, N7401, N1206);
buf BUF1 (N7406, N7397);
nor NOR4 (N7407, N7360, N5078, N2738, N3568);
or OR4 (N7408, N7402, N1160, N6232, N491);
or OR3 (N7409, N7404, N1488, N219);
nand NAND4 (N7410, N7400, N4344, N2978, N4862);
buf BUF1 (N7411, N7408);
nand NAND2 (N7412, N7405, N3033);
xor XOR2 (N7413, N7394, N401);
not NOT1 (N7414, N7411);
nor NOR2 (N7415, N7409, N349);
not NOT1 (N7416, N7399);
or OR4 (N7417, N7416, N5240, N2423, N2393);
nor NOR3 (N7418, N7413, N3123, N950);
not NOT1 (N7419, N7412);
buf BUF1 (N7420, N7418);
not NOT1 (N7421, N7414);
not NOT1 (N7422, N7406);
nor NOR2 (N7423, N7422, N2066);
nor NOR4 (N7424, N7420, N6285, N6566, N6401);
not NOT1 (N7425, N7423);
xor XOR2 (N7426, N7407, N2989);
nand NAND4 (N7427, N7417, N6707, N4152, N4534);
not NOT1 (N7428, N7415);
nand NAND2 (N7429, N7421, N3705);
nor NOR2 (N7430, N7410, N3830);
nand NAND3 (N7431, N7427, N1537, N1435);
xor XOR2 (N7432, N7426, N415);
nand NAND3 (N7433, N7395, N6723, N4955);
or OR4 (N7434, N7433, N4892, N5130, N308);
and AND3 (N7435, N7424, N1919, N5167);
buf BUF1 (N7436, N7435);
xor XOR2 (N7437, N7430, N1922);
xor XOR2 (N7438, N7431, N7247);
nor NOR3 (N7439, N7436, N348, N5454);
xor XOR2 (N7440, N7434, N7343);
not NOT1 (N7441, N7439);
or OR4 (N7442, N7388, N3492, N2991, N3414);
nor NOR3 (N7443, N7428, N6394, N6760);
nor NOR4 (N7444, N7437, N3793, N394, N797);
not NOT1 (N7445, N7429);
buf BUF1 (N7446, N7444);
buf BUF1 (N7447, N7446);
nor NOR2 (N7448, N7445, N5073);
and AND3 (N7449, N7443, N200, N1391);
nand NAND2 (N7450, N7441, N875);
or OR4 (N7451, N7440, N4260, N2234, N1683);
xor XOR2 (N7452, N7438, N5049);
nor NOR4 (N7453, N7448, N6713, N2971, N1029);
nor NOR3 (N7454, N7451, N5515, N7373);
not NOT1 (N7455, N7432);
or OR2 (N7456, N7450, N6143);
and AND3 (N7457, N7425, N2599, N1528);
and AND3 (N7458, N7453, N4106, N6345);
nor NOR3 (N7459, N7454, N4021, N4106);
or OR3 (N7460, N7455, N6700, N2506);
and AND4 (N7461, N7456, N1401, N4177, N3518);
xor XOR2 (N7462, N7460, N719);
not NOT1 (N7463, N7458);
nor NOR4 (N7464, N7457, N4304, N7432, N2122);
or OR4 (N7465, N7452, N2300, N169, N1206);
xor XOR2 (N7466, N7459, N5483);
or OR4 (N7467, N7449, N1962, N311, N1006);
not NOT1 (N7468, N7447);
xor XOR2 (N7469, N7468, N3028);
nor NOR3 (N7470, N7419, N6919, N7046);
nor NOR3 (N7471, N7463, N3888, N5622);
or OR2 (N7472, N7470, N6879);
and AND2 (N7473, N7466, N3300);
nor NOR3 (N7474, N7465, N5745, N1742);
and AND3 (N7475, N7474, N849, N5952);
xor XOR2 (N7476, N7467, N1161);
xor XOR2 (N7477, N7442, N470);
nand NAND4 (N7478, N7461, N7022, N1861, N7435);
nand NAND4 (N7479, N7473, N2075, N7114, N7270);
nand NAND2 (N7480, N7476, N7278);
and AND4 (N7481, N7462, N2246, N3875, N7252);
nand NAND3 (N7482, N7471, N183, N3035);
nor NOR4 (N7483, N7469, N6420, N3806, N4833);
buf BUF1 (N7484, N7481);
nor NOR3 (N7485, N7482, N3608, N1860);
and AND3 (N7486, N7478, N1377, N6595);
not NOT1 (N7487, N7472);
and AND4 (N7488, N7477, N6523, N4280, N7132);
nand NAND3 (N7489, N7480, N6445, N84);
or OR2 (N7490, N7486, N6039);
and AND3 (N7491, N7479, N2370, N2624);
nor NOR4 (N7492, N7464, N4126, N2968, N6137);
and AND3 (N7493, N7475, N5396, N4231);
xor XOR2 (N7494, N7488, N328);
buf BUF1 (N7495, N7487);
nand NAND3 (N7496, N7489, N4368, N7191);
nor NOR2 (N7497, N7492, N59);
not NOT1 (N7498, N7483);
not NOT1 (N7499, N7496);
xor XOR2 (N7500, N7484, N5226);
xor XOR2 (N7501, N7490, N6355);
nor NOR2 (N7502, N7485, N5885);
and AND4 (N7503, N7498, N797, N1348, N2196);
not NOT1 (N7504, N7497);
or OR3 (N7505, N7500, N1459, N908);
buf BUF1 (N7506, N7502);
buf BUF1 (N7507, N7499);
nor NOR4 (N7508, N7501, N6676, N3517, N5770);
xor XOR2 (N7509, N7505, N6395);
nand NAND3 (N7510, N7495, N1460, N4829);
nor NOR4 (N7511, N7494, N1692, N412, N406);
nand NAND3 (N7512, N7509, N1655, N102);
or OR3 (N7513, N7511, N754, N875);
or OR3 (N7514, N7513, N1308, N3680);
and AND2 (N7515, N7514, N1658);
nand NAND4 (N7516, N7503, N477, N2927, N3431);
and AND4 (N7517, N7491, N1282, N4346, N3126);
buf BUF1 (N7518, N7516);
xor XOR2 (N7519, N7512, N2625);
nor NOR4 (N7520, N7508, N4208, N4822, N6382);
xor XOR2 (N7521, N7507, N5173);
buf BUF1 (N7522, N7515);
buf BUF1 (N7523, N7522);
nor NOR3 (N7524, N7506, N5962, N1236);
or OR2 (N7525, N7518, N7490);
nor NOR2 (N7526, N7517, N7409);
or OR4 (N7527, N7504, N2316, N3068, N6083);
and AND3 (N7528, N7493, N5860, N5782);
nor NOR3 (N7529, N7528, N3681, N4054);
and AND2 (N7530, N7510, N1382);
not NOT1 (N7531, N7521);
xor XOR2 (N7532, N7520, N1882);
nor NOR4 (N7533, N7526, N1172, N5641, N1690);
not NOT1 (N7534, N7519);
not NOT1 (N7535, N7530);
xor XOR2 (N7536, N7533, N2756);
xor XOR2 (N7537, N7523, N7256);
or OR2 (N7538, N7536, N6290);
not NOT1 (N7539, N7537);
not NOT1 (N7540, N7539);
buf BUF1 (N7541, N7540);
buf BUF1 (N7542, N7527);
nand NAND4 (N7543, N7524, N5003, N1486, N5211);
not NOT1 (N7544, N7529);
nand NAND3 (N7545, N7535, N3331, N805);
nor NOR2 (N7546, N7542, N3090);
xor XOR2 (N7547, N7538, N412);
nand NAND2 (N7548, N7541, N2021);
buf BUF1 (N7549, N7534);
not NOT1 (N7550, N7545);
and AND4 (N7551, N7543, N2156, N1208, N502);
buf BUF1 (N7552, N7551);
or OR3 (N7553, N7544, N6912, N2544);
and AND4 (N7554, N7531, N1677, N2354, N4802);
or OR2 (N7555, N7552, N6552);
nor NOR4 (N7556, N7553, N2261, N4000, N737);
not NOT1 (N7557, N7548);
xor XOR2 (N7558, N7550, N2490);
buf BUF1 (N7559, N7546);
xor XOR2 (N7560, N7557, N1481);
or OR2 (N7561, N7532, N538);
nor NOR3 (N7562, N7561, N1239, N4353);
or OR2 (N7563, N7525, N979);
xor XOR2 (N7564, N7547, N4293);
nand NAND3 (N7565, N7559, N7032, N3186);
xor XOR2 (N7566, N7554, N1759);
or OR4 (N7567, N7556, N5553, N4600, N4128);
xor XOR2 (N7568, N7558, N3678);
or OR2 (N7569, N7549, N2499);
xor XOR2 (N7570, N7568, N6112);
buf BUF1 (N7571, N7562);
and AND3 (N7572, N7570, N6692, N7293);
xor XOR2 (N7573, N7563, N5562);
and AND2 (N7574, N7567, N837);
nor NOR3 (N7575, N7569, N947, N1161);
nand NAND4 (N7576, N7574, N697, N5147, N2651);
not NOT1 (N7577, N7566);
or OR3 (N7578, N7573, N840, N5769);
and AND4 (N7579, N7572, N1058, N503, N6065);
xor XOR2 (N7580, N7564, N2521);
not NOT1 (N7581, N7565);
nor NOR3 (N7582, N7581, N1660, N4001);
buf BUF1 (N7583, N7580);
or OR4 (N7584, N7578, N2683, N3374, N3292);
buf BUF1 (N7585, N7577);
nand NAND3 (N7586, N7585, N6054, N7546);
buf BUF1 (N7587, N7560);
xor XOR2 (N7588, N7575, N878);
xor XOR2 (N7589, N7588, N7387);
buf BUF1 (N7590, N7583);
or OR2 (N7591, N7586, N2283);
buf BUF1 (N7592, N7589);
xor XOR2 (N7593, N7576, N4597);
xor XOR2 (N7594, N7582, N2285);
buf BUF1 (N7595, N7590);
nor NOR4 (N7596, N7587, N267, N1274, N5150);
or OR3 (N7597, N7594, N6275, N2467);
xor XOR2 (N7598, N7596, N2862);
and AND4 (N7599, N7593, N861, N3362, N6562);
xor XOR2 (N7600, N7584, N5168);
nand NAND3 (N7601, N7595, N1317, N618);
buf BUF1 (N7602, N7599);
nor NOR2 (N7603, N7598, N5048);
buf BUF1 (N7604, N7579);
xor XOR2 (N7605, N7602, N3152);
or OR3 (N7606, N7600, N7047, N3352);
or OR2 (N7607, N7597, N5045);
nor NOR2 (N7608, N7601, N6187);
nor NOR2 (N7609, N7604, N2180);
xor XOR2 (N7610, N7571, N1785);
or OR2 (N7611, N7606, N1734);
nor NOR2 (N7612, N7605, N4392);
nor NOR4 (N7613, N7610, N522, N2813, N6724);
xor XOR2 (N7614, N7607, N6910);
or OR4 (N7615, N7611, N550, N3944, N4197);
xor XOR2 (N7616, N7603, N3352);
nor NOR3 (N7617, N7614, N1095, N4005);
or OR3 (N7618, N7555, N530, N3108);
nor NOR4 (N7619, N7617, N5528, N7108, N3181);
buf BUF1 (N7620, N7615);
and AND3 (N7621, N7616, N4459, N6478);
not NOT1 (N7622, N7613);
nor NOR2 (N7623, N7612, N5080);
nor NOR2 (N7624, N7622, N2795);
buf BUF1 (N7625, N7592);
not NOT1 (N7626, N7620);
nor NOR4 (N7627, N7624, N31, N6127, N6738);
xor XOR2 (N7628, N7627, N1104);
nand NAND4 (N7629, N7623, N6953, N2495, N3005);
or OR4 (N7630, N7618, N429, N7208, N1134);
or OR4 (N7631, N7591, N653, N2122, N4911);
nand NAND4 (N7632, N7630, N708, N6849, N3584);
and AND3 (N7633, N7626, N5852, N7454);
or OR2 (N7634, N7632, N7276);
or OR3 (N7635, N7631, N3346, N5555);
buf BUF1 (N7636, N7609);
not NOT1 (N7637, N7621);
and AND3 (N7638, N7634, N3780, N4827);
not NOT1 (N7639, N7608);
or OR4 (N7640, N7638, N1992, N1904, N5583);
not NOT1 (N7641, N7625);
buf BUF1 (N7642, N7633);
nor NOR2 (N7643, N7628, N5516);
nor NOR4 (N7644, N7619, N5870, N5473, N185);
or OR2 (N7645, N7636, N1223);
or OR2 (N7646, N7639, N1349);
and AND4 (N7647, N7637, N1547, N6980, N2137);
or OR3 (N7648, N7644, N7537, N5611);
nor NOR3 (N7649, N7641, N4464, N644);
buf BUF1 (N7650, N7645);
nor NOR3 (N7651, N7646, N3257, N4123);
nand NAND4 (N7652, N7649, N6104, N447, N7522);
nor NOR3 (N7653, N7643, N5979, N2765);
or OR2 (N7654, N7635, N4531);
not NOT1 (N7655, N7629);
nor NOR4 (N7656, N7647, N4902, N2786, N6285);
or OR4 (N7657, N7656, N6271, N4716, N3254);
not NOT1 (N7658, N7640);
not NOT1 (N7659, N7654);
nand NAND3 (N7660, N7650, N4222, N4322);
xor XOR2 (N7661, N7652, N5812);
not NOT1 (N7662, N7660);
buf BUF1 (N7663, N7662);
xor XOR2 (N7664, N7642, N4035);
or OR4 (N7665, N7658, N6879, N2373, N6248);
or OR4 (N7666, N7664, N3100, N7434, N3636);
and AND2 (N7667, N7663, N6299);
not NOT1 (N7668, N7655);
buf BUF1 (N7669, N7648);
and AND4 (N7670, N7653, N2440, N115, N6054);
buf BUF1 (N7671, N7666);
or OR4 (N7672, N7659, N5131, N2419, N4894);
nor NOR2 (N7673, N7665, N662);
buf BUF1 (N7674, N7651);
not NOT1 (N7675, N7673);
not NOT1 (N7676, N7669);
or OR3 (N7677, N7667, N4579, N545);
not NOT1 (N7678, N7661);
nand NAND4 (N7679, N7676, N610, N6384, N754);
nand NAND3 (N7680, N7657, N6606, N339);
nand NAND4 (N7681, N7680, N7057, N5345, N4231);
buf BUF1 (N7682, N7670);
or OR2 (N7683, N7674, N6533);
nand NAND4 (N7684, N7668, N6416, N4956, N4025);
buf BUF1 (N7685, N7678);
nand NAND4 (N7686, N7679, N7589, N7593, N7352);
not NOT1 (N7687, N7683);
nor NOR4 (N7688, N7677, N4427, N3896, N5812);
not NOT1 (N7689, N7671);
xor XOR2 (N7690, N7686, N5253);
xor XOR2 (N7691, N7687, N2193);
nand NAND2 (N7692, N7691, N3404);
or OR3 (N7693, N7689, N1408, N5980);
xor XOR2 (N7694, N7692, N2673);
nor NOR2 (N7695, N7690, N2916);
nand NAND4 (N7696, N7672, N7019, N7472, N118);
nand NAND2 (N7697, N7684, N7148);
or OR4 (N7698, N7688, N6654, N3921, N6075);
xor XOR2 (N7699, N7698, N7302);
nor NOR4 (N7700, N7697, N3323, N5876, N3971);
xor XOR2 (N7701, N7685, N1272);
xor XOR2 (N7702, N7675, N2846);
xor XOR2 (N7703, N7682, N3659);
and AND4 (N7704, N7703, N6171, N2860, N4875);
not NOT1 (N7705, N7695);
nand NAND2 (N7706, N7702, N3247);
buf BUF1 (N7707, N7681);
buf BUF1 (N7708, N7696);
xor XOR2 (N7709, N7694, N623);
buf BUF1 (N7710, N7704);
nor NOR4 (N7711, N7699, N6318, N5209, N7446);
or OR4 (N7712, N7709, N1081, N6114, N159);
or OR2 (N7713, N7711, N1500);
buf BUF1 (N7714, N7708);
or OR3 (N7715, N7707, N2065, N3503);
xor XOR2 (N7716, N7705, N2232);
nor NOR4 (N7717, N7712, N5289, N3245, N7453);
and AND2 (N7718, N7715, N4524);
nor NOR2 (N7719, N7716, N4880);
buf BUF1 (N7720, N7700);
buf BUF1 (N7721, N7720);
nand NAND2 (N7722, N7706, N3618);
or OR3 (N7723, N7693, N4622, N5588);
xor XOR2 (N7724, N7714, N1522);
xor XOR2 (N7725, N7713, N654);
xor XOR2 (N7726, N7722, N936);
buf BUF1 (N7727, N7726);
nand NAND2 (N7728, N7725, N7472);
xor XOR2 (N7729, N7718, N7298);
not NOT1 (N7730, N7723);
or OR4 (N7731, N7724, N3368, N2689, N4757);
nand NAND2 (N7732, N7717, N3332);
not NOT1 (N7733, N7731);
or OR3 (N7734, N7710, N5074, N585);
buf BUF1 (N7735, N7730);
nor NOR4 (N7736, N7701, N3178, N4164, N3584);
not NOT1 (N7737, N7719);
nor NOR3 (N7738, N7734, N7207, N7328);
xor XOR2 (N7739, N7721, N1140);
xor XOR2 (N7740, N7736, N6430);
nor NOR4 (N7741, N7732, N2504, N4592, N4227);
or OR4 (N7742, N7739, N3809, N6847, N6294);
buf BUF1 (N7743, N7737);
and AND3 (N7744, N7741, N224, N442);
not NOT1 (N7745, N7742);
nor NOR4 (N7746, N7745, N1598, N6276, N1625);
nand NAND3 (N7747, N7729, N2115, N5783);
not NOT1 (N7748, N7747);
not NOT1 (N7749, N7733);
buf BUF1 (N7750, N7735);
nand NAND4 (N7751, N7727, N5194, N67, N66);
buf BUF1 (N7752, N7751);
and AND3 (N7753, N7744, N6584, N1173);
buf BUF1 (N7754, N7752);
buf BUF1 (N7755, N7740);
nor NOR2 (N7756, N7754, N3221);
xor XOR2 (N7757, N7756, N7056);
buf BUF1 (N7758, N7750);
and AND4 (N7759, N7743, N7401, N1652, N4002);
nor NOR2 (N7760, N7755, N159);
and AND2 (N7761, N7738, N453);
nand NAND4 (N7762, N7759, N784, N3159, N833);
buf BUF1 (N7763, N7762);
nor NOR3 (N7764, N7753, N753, N7383);
not NOT1 (N7765, N7749);
nor NOR4 (N7766, N7760, N6529, N2999, N4531);
nor NOR3 (N7767, N7757, N74, N2566);
nor NOR2 (N7768, N7765, N4285);
or OR2 (N7769, N7761, N770);
and AND2 (N7770, N7769, N690);
or OR4 (N7771, N7728, N6176, N4116, N223);
nor NOR3 (N7772, N7770, N7018, N4220);
xor XOR2 (N7773, N7772, N2846);
xor XOR2 (N7774, N7766, N5346);
and AND2 (N7775, N7758, N3538);
xor XOR2 (N7776, N7767, N3593);
not NOT1 (N7777, N7774);
and AND4 (N7778, N7773, N5608, N4886, N5103);
nand NAND2 (N7779, N7768, N5517);
or OR3 (N7780, N7778, N19, N5918);
not NOT1 (N7781, N7771);
buf BUF1 (N7782, N7776);
and AND3 (N7783, N7781, N1587, N7120);
and AND3 (N7784, N7779, N5646, N7197);
xor XOR2 (N7785, N7746, N5067);
nor NOR3 (N7786, N7780, N6741, N3685);
nand NAND3 (N7787, N7748, N6366, N7067);
buf BUF1 (N7788, N7775);
nor NOR4 (N7789, N7782, N4122, N3558, N4160);
nand NAND3 (N7790, N7785, N7782, N4993);
xor XOR2 (N7791, N7783, N1632);
nor NOR4 (N7792, N7789, N71, N5040, N2418);
xor XOR2 (N7793, N7792, N4429);
nor NOR3 (N7794, N7763, N6197, N7547);
or OR3 (N7795, N7790, N4512, N1064);
not NOT1 (N7796, N7764);
buf BUF1 (N7797, N7796);
nand NAND3 (N7798, N7793, N3664, N2788);
not NOT1 (N7799, N7788);
not NOT1 (N7800, N7791);
not NOT1 (N7801, N7794);
nor NOR3 (N7802, N7798, N1642, N7485);
nor NOR3 (N7803, N7777, N5098, N5624);
xor XOR2 (N7804, N7802, N281);
nand NAND4 (N7805, N7799, N5855, N4699, N2729);
or OR3 (N7806, N7801, N3312, N3285);
or OR2 (N7807, N7806, N476);
not NOT1 (N7808, N7797);
and AND3 (N7809, N7804, N1989, N7616);
xor XOR2 (N7810, N7809, N2537);
not NOT1 (N7811, N7784);
and AND2 (N7812, N7787, N492);
nand NAND2 (N7813, N7812, N4615);
xor XOR2 (N7814, N7800, N2853);
or OR3 (N7815, N7811, N1964, N3395);
and AND2 (N7816, N7815, N3488);
not NOT1 (N7817, N7803);
not NOT1 (N7818, N7795);
nor NOR2 (N7819, N7808, N1730);
nand NAND4 (N7820, N7810, N7678, N2881, N6252);
nand NAND3 (N7821, N7814, N4770, N3974);
or OR4 (N7822, N7816, N7608, N1794, N3397);
xor XOR2 (N7823, N7818, N6354);
or OR3 (N7824, N7807, N1548, N1920);
not NOT1 (N7825, N7822);
xor XOR2 (N7826, N7821, N6571);
buf BUF1 (N7827, N7786);
not NOT1 (N7828, N7820);
and AND3 (N7829, N7817, N4547, N2653);
and AND2 (N7830, N7827, N5285);
not NOT1 (N7831, N7805);
or OR4 (N7832, N7825, N605, N272, N7353);
and AND4 (N7833, N7823, N7672, N3221, N1421);
not NOT1 (N7834, N7819);
xor XOR2 (N7835, N7813, N2135);
or OR2 (N7836, N7830, N1326);
and AND4 (N7837, N7824, N6281, N3448, N2436);
or OR2 (N7838, N7828, N1196);
and AND2 (N7839, N7837, N7611);
xor XOR2 (N7840, N7835, N2032);
and AND3 (N7841, N7838, N7301, N6849);
and AND3 (N7842, N7831, N4767, N5174);
not NOT1 (N7843, N7832);
not NOT1 (N7844, N7833);
and AND4 (N7845, N7844, N6653, N7690, N7096);
not NOT1 (N7846, N7843);
and AND4 (N7847, N7845, N5514, N4206, N6232);
or OR3 (N7848, N7846, N6823, N6735);
xor XOR2 (N7849, N7839, N456);
or OR3 (N7850, N7840, N5932, N2396);
xor XOR2 (N7851, N7834, N6963);
and AND2 (N7852, N7848, N6514);
or OR2 (N7853, N7851, N6853);
and AND3 (N7854, N7847, N7718, N6383);
nand NAND2 (N7855, N7829, N5477);
and AND3 (N7856, N7826, N4979, N6478);
nand NAND3 (N7857, N7836, N3235, N332);
buf BUF1 (N7858, N7849);
not NOT1 (N7859, N7856);
nand NAND3 (N7860, N7841, N1244, N260);
or OR4 (N7861, N7859, N1677, N415, N2126);
not NOT1 (N7862, N7853);
buf BUF1 (N7863, N7861);
not NOT1 (N7864, N7852);
nand NAND3 (N7865, N7863, N7621, N7404);
or OR2 (N7866, N7858, N2714);
nand NAND4 (N7867, N7854, N3134, N1580, N4614);
buf BUF1 (N7868, N7864);
not NOT1 (N7869, N7860);
xor XOR2 (N7870, N7866, N5345);
xor XOR2 (N7871, N7870, N7760);
not NOT1 (N7872, N7842);
not NOT1 (N7873, N7872);
xor XOR2 (N7874, N7850, N4057);
nor NOR4 (N7875, N7874, N18, N7783, N4045);
not NOT1 (N7876, N7857);
xor XOR2 (N7877, N7871, N7613);
xor XOR2 (N7878, N7867, N5455);
xor XOR2 (N7879, N7878, N5185);
nand NAND3 (N7880, N7873, N2636, N3116);
buf BUF1 (N7881, N7879);
not NOT1 (N7882, N7865);
xor XOR2 (N7883, N7869, N4508);
and AND3 (N7884, N7876, N4584, N3557);
or OR3 (N7885, N7881, N3988, N6136);
nand NAND3 (N7886, N7883, N7578, N528);
nor NOR4 (N7887, N7885, N2114, N5485, N6678);
and AND3 (N7888, N7887, N5784, N307);
and AND3 (N7889, N7884, N4445, N2872);
not NOT1 (N7890, N7882);
and AND2 (N7891, N7889, N4962);
xor XOR2 (N7892, N7877, N4582);
and AND3 (N7893, N7892, N1502, N7437);
xor XOR2 (N7894, N7862, N2864);
not NOT1 (N7895, N7868);
nand NAND4 (N7896, N7895, N7821, N4759, N767);
not NOT1 (N7897, N7894);
and AND2 (N7898, N7855, N5045);
nand NAND2 (N7899, N7896, N4722);
and AND3 (N7900, N7898, N5196, N118);
and AND2 (N7901, N7900, N7374);
nand NAND4 (N7902, N7901, N1800, N4165, N736);
nand NAND4 (N7903, N7899, N7824, N1530, N3154);
not NOT1 (N7904, N7891);
and AND3 (N7905, N7888, N5323, N7774);
buf BUF1 (N7906, N7880);
or OR3 (N7907, N7903, N3828, N3020);
xor XOR2 (N7908, N7907, N3202);
and AND4 (N7909, N7886, N4046, N7461, N5851);
or OR2 (N7910, N7905, N3611);
nor NOR3 (N7911, N7904, N7482, N5472);
or OR4 (N7912, N7893, N2989, N151, N862);
and AND2 (N7913, N7910, N3047);
nor NOR2 (N7914, N7908, N17);
not NOT1 (N7915, N7909);
and AND4 (N7916, N7911, N4917, N933, N2973);
nor NOR2 (N7917, N7906, N1447);
or OR2 (N7918, N7916, N999);
nor NOR3 (N7919, N7913, N690, N7291);
and AND3 (N7920, N7918, N1256, N7762);
not NOT1 (N7921, N7914);
or OR4 (N7922, N7902, N7102, N4705, N1780);
or OR4 (N7923, N7920, N4946, N1168, N5798);
and AND4 (N7924, N7875, N2283, N4918, N5363);
xor XOR2 (N7925, N7912, N1692);
nand NAND3 (N7926, N7923, N5923, N7533);
not NOT1 (N7927, N7917);
or OR2 (N7928, N7919, N4359);
not NOT1 (N7929, N7915);
and AND3 (N7930, N7897, N5230, N5718);
nand NAND2 (N7931, N7928, N313);
not NOT1 (N7932, N7890);
or OR2 (N7933, N7931, N4264);
buf BUF1 (N7934, N7927);
and AND3 (N7935, N7922, N1172, N3136);
buf BUF1 (N7936, N7929);
xor XOR2 (N7937, N7930, N7011);
xor XOR2 (N7938, N7921, N2448);
not NOT1 (N7939, N7932);
buf BUF1 (N7940, N7925);
nand NAND4 (N7941, N7926, N1300, N3420, N352);
nand NAND4 (N7942, N7940, N5868, N6275, N1643);
xor XOR2 (N7943, N7941, N5483);
and AND4 (N7944, N7943, N15, N3421, N2332);
xor XOR2 (N7945, N7924, N7344);
nor NOR4 (N7946, N7939, N3718, N5790, N4326);
and AND4 (N7947, N7942, N2817, N461, N2923);
buf BUF1 (N7948, N7934);
or OR2 (N7949, N7944, N3900);
xor XOR2 (N7950, N7945, N6111);
buf BUF1 (N7951, N7937);
xor XOR2 (N7952, N7950, N1352);
nand NAND2 (N7953, N7947, N2719);
nor NOR4 (N7954, N7933, N4621, N6777, N1406);
xor XOR2 (N7955, N7953, N3432);
or OR3 (N7956, N7936, N5543, N653);
and AND2 (N7957, N7952, N3109);
xor XOR2 (N7958, N7949, N582);
or OR4 (N7959, N7951, N1241, N4975, N5475);
or OR2 (N7960, N7946, N6492);
buf BUF1 (N7961, N7959);
not NOT1 (N7962, N7948);
nor NOR4 (N7963, N7958, N2038, N1467, N7062);
xor XOR2 (N7964, N7954, N3596);
and AND3 (N7965, N7956, N1054, N923);
and AND4 (N7966, N7935, N2085, N6378, N4555);
or OR4 (N7967, N7962, N6183, N1133, N2858);
or OR3 (N7968, N7955, N7543, N5572);
nor NOR3 (N7969, N7964, N3539, N3550);
nor NOR2 (N7970, N7938, N6814);
nand NAND3 (N7971, N7968, N5959, N7129);
or OR2 (N7972, N7970, N7432);
nor NOR3 (N7973, N7966, N2239, N4613);
or OR2 (N7974, N7960, N6996);
not NOT1 (N7975, N7963);
and AND2 (N7976, N7965, N5067);
or OR2 (N7977, N7975, N4104);
nor NOR3 (N7978, N7977, N4233, N2083);
and AND3 (N7979, N7961, N4857, N6376);
buf BUF1 (N7980, N7967);
nand NAND3 (N7981, N7978, N2705, N4221);
nand NAND3 (N7982, N7972, N6676, N2572);
buf BUF1 (N7983, N7969);
xor XOR2 (N7984, N7976, N559);
not NOT1 (N7985, N7982);
buf BUF1 (N7986, N7983);
xor XOR2 (N7987, N7985, N4625);
and AND3 (N7988, N7979, N7906, N4949);
nor NOR4 (N7989, N7971, N2530, N1844, N7721);
nand NAND3 (N7990, N7984, N5757, N5818);
nor NOR3 (N7991, N7989, N5090, N3105);
xor XOR2 (N7992, N7990, N1964);
or OR2 (N7993, N7986, N468);
not NOT1 (N7994, N7988);
or OR4 (N7995, N7991, N6080, N6400, N7401);
not NOT1 (N7996, N7973);
and AND3 (N7997, N7996, N6185, N6132);
and AND3 (N7998, N7995, N4248, N4215);
buf BUF1 (N7999, N7981);
buf BUF1 (N8000, N7987);
buf BUF1 (N8001, N7957);
buf BUF1 (N8002, N7974);
buf BUF1 (N8003, N7997);
or OR2 (N8004, N7992, N7005);
or OR4 (N8005, N7999, N4442, N2185, N4386);
and AND2 (N8006, N7998, N3048);
buf BUF1 (N8007, N8002);
and AND4 (N8008, N8007, N442, N3926, N6647);
nor NOR2 (N8009, N8004, N6265);
or OR3 (N8010, N7980, N2161, N7591);
not NOT1 (N8011, N8009);
nand NAND3 (N8012, N7994, N1663, N763);
xor XOR2 (N8013, N8005, N5466);
not NOT1 (N8014, N8000);
or OR3 (N8015, N8014, N4012, N3012);
not NOT1 (N8016, N8010);
nor NOR4 (N8017, N8012, N693, N1051, N4138);
or OR2 (N8018, N7993, N4896);
not NOT1 (N8019, N8003);
not NOT1 (N8020, N8017);
buf BUF1 (N8021, N8018);
nor NOR4 (N8022, N8008, N1820, N678, N8014);
nand NAND2 (N8023, N8016, N7354);
xor XOR2 (N8024, N8021, N4684);
not NOT1 (N8025, N8024);
buf BUF1 (N8026, N8020);
nand NAND2 (N8027, N8013, N2261);
buf BUF1 (N8028, N8026);
and AND2 (N8029, N8006, N4709);
buf BUF1 (N8030, N8025);
not NOT1 (N8031, N8029);
or OR3 (N8032, N8028, N183, N604);
xor XOR2 (N8033, N8023, N6664);
buf BUF1 (N8034, N8030);
nor NOR2 (N8035, N8034, N1207);
or OR2 (N8036, N8022, N1874);
nand NAND3 (N8037, N8033, N7541, N6425);
and AND4 (N8038, N8011, N2380, N5478, N247);
xor XOR2 (N8039, N8035, N1737);
nand NAND4 (N8040, N8001, N6908, N1783, N4884);
or OR4 (N8041, N8039, N5576, N320, N3753);
nor NOR2 (N8042, N8027, N5253);
or OR3 (N8043, N8032, N460, N6763);
buf BUF1 (N8044, N8031);
not NOT1 (N8045, N8044);
or OR2 (N8046, N8037, N7109);
or OR2 (N8047, N8046, N4407);
nor NOR4 (N8048, N8041, N6115, N6391, N1564);
nand NAND2 (N8049, N8040, N6149);
buf BUF1 (N8050, N8042);
nand NAND4 (N8051, N8036, N1851, N1784, N6044);
not NOT1 (N8052, N8048);
not NOT1 (N8053, N8050);
or OR2 (N8054, N8038, N6048);
buf BUF1 (N8055, N8043);
and AND3 (N8056, N8051, N6503, N3492);
xor XOR2 (N8057, N8053, N4632);
and AND4 (N8058, N8049, N3265, N7368, N2717);
nor NOR4 (N8059, N8056, N436, N7041, N3356);
or OR3 (N8060, N8052, N7646, N167);
xor XOR2 (N8061, N8057, N3163);
nor NOR2 (N8062, N8055, N2842);
nor NOR4 (N8063, N8054, N4234, N2408, N3328);
nand NAND2 (N8064, N8047, N1343);
and AND4 (N8065, N8058, N2198, N6642, N5016);
nor NOR2 (N8066, N8064, N4438);
nor NOR3 (N8067, N8065, N3469, N1141);
and AND4 (N8068, N8061, N2239, N7829, N2125);
not NOT1 (N8069, N8015);
not NOT1 (N8070, N8066);
nand NAND4 (N8071, N8069, N3710, N424, N929);
xor XOR2 (N8072, N8063, N6267);
nand NAND2 (N8073, N8070, N84);
or OR3 (N8074, N8068, N6177, N7784);
xor XOR2 (N8075, N8062, N6776);
buf BUF1 (N8076, N8072);
and AND4 (N8077, N8067, N2388, N2833, N8009);
buf BUF1 (N8078, N8075);
or OR3 (N8079, N8073, N331, N3967);
not NOT1 (N8080, N8060);
or OR2 (N8081, N8059, N1552);
not NOT1 (N8082, N8076);
not NOT1 (N8083, N8045);
not NOT1 (N8084, N8077);
not NOT1 (N8085, N8084);
and AND3 (N8086, N8083, N5090, N5869);
and AND2 (N8087, N8086, N5767);
not NOT1 (N8088, N8071);
nand NAND4 (N8089, N8074, N7120, N5277, N2008);
or OR3 (N8090, N8078, N7499, N6392);
or OR4 (N8091, N8085, N3699, N1767, N6377);
and AND3 (N8092, N8091, N4125, N1037);
or OR2 (N8093, N8081, N6199);
and AND4 (N8094, N8093, N5667, N625, N3629);
buf BUF1 (N8095, N8088);
xor XOR2 (N8096, N8082, N6799);
buf BUF1 (N8097, N8090);
nor NOR2 (N8098, N8092, N3681);
and AND4 (N8099, N8089, N2690, N2746, N7335);
nand NAND4 (N8100, N8098, N3981, N7488, N1886);
xor XOR2 (N8101, N8096, N497);
nand NAND4 (N8102, N8087, N7243, N1867, N6633);
xor XOR2 (N8103, N8080, N4642);
nand NAND4 (N8104, N8101, N7843, N1633, N6704);
xor XOR2 (N8105, N8097, N3935);
or OR3 (N8106, N8102, N4039, N5542);
buf BUF1 (N8107, N8103);
nor NOR4 (N8108, N8104, N4288, N521, N857);
nor NOR3 (N8109, N8079, N4808, N5395);
nand NAND2 (N8110, N8094, N6173);
not NOT1 (N8111, N8100);
nor NOR3 (N8112, N8099, N6567, N94);
and AND2 (N8113, N8111, N4460);
or OR4 (N8114, N8105, N4385, N5751, N5996);
buf BUF1 (N8115, N8106);
xor XOR2 (N8116, N8095, N3433);
not NOT1 (N8117, N8114);
not NOT1 (N8118, N8107);
not NOT1 (N8119, N8108);
xor XOR2 (N8120, N8109, N5597);
and AND4 (N8121, N8113, N5904, N6421, N2040);
nor NOR4 (N8122, N8115, N7929, N2537, N7644);
xor XOR2 (N8123, N8122, N1345);
buf BUF1 (N8124, N8118);
xor XOR2 (N8125, N8121, N5884);
or OR4 (N8126, N8117, N5119, N64, N928);
nand NAND2 (N8127, N8126, N1456);
nand NAND2 (N8128, N8112, N4498);
nor NOR2 (N8129, N8120, N3650);
buf BUF1 (N8130, N8019);
nand NAND3 (N8131, N8128, N6021, N3838);
nor NOR3 (N8132, N8110, N1635, N2072);
nand NAND4 (N8133, N8127, N7796, N4687, N3950);
xor XOR2 (N8134, N8129, N2634);
buf BUF1 (N8135, N8123);
and AND4 (N8136, N8119, N777, N5294, N4419);
not NOT1 (N8137, N8132);
buf BUF1 (N8138, N8134);
and AND4 (N8139, N8116, N3352, N3611, N94);
and AND2 (N8140, N8135, N1467);
nor NOR4 (N8141, N8139, N6847, N5521, N5089);
nor NOR2 (N8142, N8131, N2478);
not NOT1 (N8143, N8133);
xor XOR2 (N8144, N8124, N2476);
nand NAND3 (N8145, N8142, N5619, N2059);
or OR2 (N8146, N8144, N2788);
or OR4 (N8147, N8140, N5979, N8099, N2172);
or OR4 (N8148, N8145, N7926, N5135, N7508);
or OR3 (N8149, N8137, N382, N3534);
and AND4 (N8150, N8147, N6136, N6483, N5078);
or OR2 (N8151, N8136, N3492);
or OR2 (N8152, N8150, N6806);
nand NAND3 (N8153, N8151, N3063, N2159);
xor XOR2 (N8154, N8149, N7292);
nand NAND3 (N8155, N8141, N1578, N1278);
buf BUF1 (N8156, N8154);
or OR3 (N8157, N8138, N2833, N866);
buf BUF1 (N8158, N8155);
nand NAND2 (N8159, N8152, N6347);
not NOT1 (N8160, N8143);
buf BUF1 (N8161, N8158);
buf BUF1 (N8162, N8130);
or OR2 (N8163, N8161, N419);
nand NAND3 (N8164, N8160, N384, N6139);
and AND4 (N8165, N8163, N2704, N7113, N3951);
and AND4 (N8166, N8165, N1646, N748, N5453);
and AND2 (N8167, N8157, N4012);
nand NAND2 (N8168, N8159, N5284);
buf BUF1 (N8169, N8146);
and AND4 (N8170, N8148, N950, N4578, N3393);
nor NOR2 (N8171, N8125, N5745);
nor NOR3 (N8172, N8166, N5401, N3002);
and AND3 (N8173, N8156, N7629, N4208);
nor NOR3 (N8174, N8169, N5685, N3295);
and AND2 (N8175, N8167, N4306);
xor XOR2 (N8176, N8162, N7925);
nor NOR3 (N8177, N8172, N571, N2075);
not NOT1 (N8178, N8153);
nand NAND2 (N8179, N8173, N2693);
not NOT1 (N8180, N8174);
xor XOR2 (N8181, N8179, N7045);
xor XOR2 (N8182, N8176, N5065);
buf BUF1 (N8183, N8168);
nand NAND4 (N8184, N8171, N4936, N6004, N5713);
and AND4 (N8185, N8164, N6685, N687, N6706);
not NOT1 (N8186, N8175);
or OR2 (N8187, N8186, N4761);
not NOT1 (N8188, N8184);
nor NOR2 (N8189, N8180, N250);
nor NOR4 (N8190, N8185, N367, N2836, N1300);
xor XOR2 (N8191, N8178, N1184);
or OR4 (N8192, N8183, N5179, N3800, N6569);
xor XOR2 (N8193, N8191, N5698);
buf BUF1 (N8194, N8181);
not NOT1 (N8195, N8194);
or OR4 (N8196, N8190, N1317, N7201, N1034);
and AND3 (N8197, N8195, N5912, N6422);
nand NAND4 (N8198, N8196, N1045, N2032, N4591);
nand NAND3 (N8199, N8188, N171, N190);
and AND3 (N8200, N8198, N5307, N2985);
nand NAND4 (N8201, N8177, N2140, N6970, N5777);
and AND4 (N8202, N8192, N1909, N2859, N3516);
xor XOR2 (N8203, N8189, N341);
buf BUF1 (N8204, N8182);
buf BUF1 (N8205, N8199);
xor XOR2 (N8206, N8203, N3434);
nand NAND2 (N8207, N8205, N1724);
not NOT1 (N8208, N8197);
and AND3 (N8209, N8170, N7222, N156);
xor XOR2 (N8210, N8187, N4525);
xor XOR2 (N8211, N8208, N6517);
nand NAND4 (N8212, N8209, N2944, N555, N2419);
xor XOR2 (N8213, N8204, N1429);
not NOT1 (N8214, N8193);
and AND4 (N8215, N8213, N2733, N656, N1484);
nand NAND4 (N8216, N8202, N3816, N594, N1874);
nor NOR2 (N8217, N8210, N3018);
not NOT1 (N8218, N8200);
or OR2 (N8219, N8206, N6168);
or OR3 (N8220, N8219, N5277, N663);
not NOT1 (N8221, N8217);
nand NAND4 (N8222, N8201, N6238, N6916, N503);
not NOT1 (N8223, N8215);
or OR2 (N8224, N8220, N741);
xor XOR2 (N8225, N8224, N4609);
and AND3 (N8226, N8212, N5158, N1450);
or OR4 (N8227, N8216, N1652, N1433, N3264);
xor XOR2 (N8228, N8222, N398);
or OR2 (N8229, N8214, N8198);
not NOT1 (N8230, N8211);
nor NOR4 (N8231, N8218, N7419, N1512, N3184);
nor NOR3 (N8232, N8228, N1007, N3495);
and AND4 (N8233, N8225, N5660, N3254, N4461);
nor NOR3 (N8234, N8230, N3037, N7196);
nor NOR2 (N8235, N8232, N8063);
xor XOR2 (N8236, N8223, N8107);
not NOT1 (N8237, N8207);
nor NOR3 (N8238, N8227, N6965, N1842);
nor NOR2 (N8239, N8233, N6414);
and AND2 (N8240, N8234, N124);
buf BUF1 (N8241, N8221);
buf BUF1 (N8242, N8236);
buf BUF1 (N8243, N8231);
or OR2 (N8244, N8240, N154);
or OR3 (N8245, N8244, N6787, N3885);
or OR2 (N8246, N8241, N1600);
or OR4 (N8247, N8246, N4215, N1963, N5020);
nor NOR4 (N8248, N8243, N2145, N6302, N5858);
nand NAND3 (N8249, N8238, N6678, N8012);
not NOT1 (N8250, N8249);
not NOT1 (N8251, N8237);
xor XOR2 (N8252, N8235, N6644);
buf BUF1 (N8253, N8251);
or OR4 (N8254, N8248, N2650, N7095, N5707);
not NOT1 (N8255, N8239);
nand NAND4 (N8256, N8245, N7584, N8196, N155);
and AND3 (N8257, N8255, N7691, N867);
or OR2 (N8258, N8247, N4872);
xor XOR2 (N8259, N8254, N7581);
xor XOR2 (N8260, N8229, N2190);
nand NAND2 (N8261, N8226, N4865);
buf BUF1 (N8262, N8260);
buf BUF1 (N8263, N8256);
xor XOR2 (N8264, N8258, N6801);
xor XOR2 (N8265, N8242, N579);
not NOT1 (N8266, N8252);
xor XOR2 (N8267, N8253, N1555);
nor NOR4 (N8268, N8257, N2474, N2862, N6407);
nor NOR4 (N8269, N8267, N1652, N6424, N3039);
not NOT1 (N8270, N8266);
xor XOR2 (N8271, N8259, N7333);
nor NOR3 (N8272, N8264, N1046, N2860);
or OR3 (N8273, N8269, N6127, N5407);
not NOT1 (N8274, N8271);
or OR4 (N8275, N8261, N7391, N158, N4657);
or OR4 (N8276, N8250, N6131, N1132, N2672);
and AND2 (N8277, N8265, N108);
xor XOR2 (N8278, N8277, N4255);
not NOT1 (N8279, N8274);
nor NOR2 (N8280, N8262, N7320);
nand NAND2 (N8281, N8275, N7701);
and AND2 (N8282, N8268, N2656);
not NOT1 (N8283, N8278);
buf BUF1 (N8284, N8283);
buf BUF1 (N8285, N8281);
buf BUF1 (N8286, N8273);
or OR2 (N8287, N8272, N1792);
and AND2 (N8288, N8276, N5114);
nand NAND4 (N8289, N8282, N2115, N6252, N1830);
xor XOR2 (N8290, N8287, N1408);
buf BUF1 (N8291, N8286);
nor NOR4 (N8292, N8289, N7667, N6424, N8072);
xor XOR2 (N8293, N8280, N1293);
not NOT1 (N8294, N8270);
not NOT1 (N8295, N8279);
or OR4 (N8296, N8293, N7628, N5511, N5536);
or OR4 (N8297, N8291, N4996, N4572, N1004);
and AND3 (N8298, N8285, N7950, N190);
nor NOR2 (N8299, N8298, N2077);
not NOT1 (N8300, N8297);
not NOT1 (N8301, N8263);
xor XOR2 (N8302, N8301, N7461);
nor NOR2 (N8303, N8295, N74);
xor XOR2 (N8304, N8303, N6055);
or OR3 (N8305, N8296, N3484, N7477);
and AND3 (N8306, N8292, N1612, N6809);
and AND4 (N8307, N8304, N5538, N2542, N8048);
xor XOR2 (N8308, N8300, N6775);
not NOT1 (N8309, N8308);
or OR2 (N8310, N8288, N4973);
or OR2 (N8311, N8310, N2115);
nor NOR3 (N8312, N8309, N4701, N4314);
not NOT1 (N8313, N8311);
not NOT1 (N8314, N8306);
buf BUF1 (N8315, N8305);
and AND2 (N8316, N8290, N6141);
not NOT1 (N8317, N8284);
and AND2 (N8318, N8315, N4438);
nand NAND2 (N8319, N8302, N6865);
xor XOR2 (N8320, N8299, N7932);
nor NOR3 (N8321, N8314, N2914, N2177);
nand NAND2 (N8322, N8313, N7752);
or OR3 (N8323, N8307, N5056, N1923);
and AND3 (N8324, N8323, N291, N4715);
not NOT1 (N8325, N8321);
or OR3 (N8326, N8316, N5325, N8214);
not NOT1 (N8327, N8318);
buf BUF1 (N8328, N8319);
and AND4 (N8329, N8322, N66, N588, N2467);
nor NOR2 (N8330, N8317, N2512);
and AND4 (N8331, N8326, N5194, N5995, N4910);
xor XOR2 (N8332, N8327, N4370);
not NOT1 (N8333, N8320);
nor NOR3 (N8334, N8331, N1123, N6468);
not NOT1 (N8335, N8325);
nand NAND4 (N8336, N8329, N2745, N1898, N5637);
xor XOR2 (N8337, N8332, N6664);
and AND2 (N8338, N8324, N3968);
nand NAND3 (N8339, N8334, N7979, N1205);
not NOT1 (N8340, N8335);
or OR2 (N8341, N8328, N6386);
and AND4 (N8342, N8312, N7355, N5007, N7377);
nand NAND3 (N8343, N8333, N4209, N4863);
and AND2 (N8344, N8336, N7211);
or OR4 (N8345, N8330, N6765, N5298, N502);
not NOT1 (N8346, N8342);
nor NOR3 (N8347, N8294, N1774, N1355);
buf BUF1 (N8348, N8343);
or OR4 (N8349, N8340, N3635, N1190, N2838);
and AND4 (N8350, N8345, N4686, N4435, N3436);
and AND3 (N8351, N8349, N75, N7685);
buf BUF1 (N8352, N8351);
nor NOR4 (N8353, N8348, N181, N7138, N2142);
xor XOR2 (N8354, N8344, N4050);
and AND3 (N8355, N8346, N2841, N3123);
nor NOR2 (N8356, N8350, N7186);
or OR2 (N8357, N8353, N6929);
buf BUF1 (N8358, N8347);
or OR2 (N8359, N8339, N1383);
nand NAND4 (N8360, N8337, N5265, N2659, N5);
nand NAND3 (N8361, N8358, N1863, N3175);
nor NOR3 (N8362, N8361, N1087, N3320);
or OR4 (N8363, N8341, N5298, N2430, N7905);
not NOT1 (N8364, N8363);
and AND4 (N8365, N8362, N4274, N2118, N1697);
nand NAND2 (N8366, N8355, N8364);
xor XOR2 (N8367, N7402, N1562);
xor XOR2 (N8368, N8366, N7681);
or OR2 (N8369, N8338, N5589);
and AND3 (N8370, N8359, N4072, N387);
not NOT1 (N8371, N8354);
and AND4 (N8372, N8368, N5843, N2858, N7698);
xor XOR2 (N8373, N8372, N3698);
not NOT1 (N8374, N8370);
nand NAND3 (N8375, N8367, N1206, N8103);
or OR3 (N8376, N8369, N1303, N667);
or OR2 (N8377, N8352, N7925);
nand NAND4 (N8378, N8376, N6399, N8222, N2100);
not NOT1 (N8379, N8357);
buf BUF1 (N8380, N8377);
and AND3 (N8381, N8356, N927, N7562);
nor NOR4 (N8382, N8380, N7372, N1581, N6820);
buf BUF1 (N8383, N8379);
not NOT1 (N8384, N8360);
xor XOR2 (N8385, N8381, N5371);
or OR4 (N8386, N8374, N8083, N4831, N4095);
or OR3 (N8387, N8383, N4108, N1266);
nand NAND2 (N8388, N8375, N6270);
or OR4 (N8389, N8386, N5281, N5275, N824);
not NOT1 (N8390, N8378);
buf BUF1 (N8391, N8382);
buf BUF1 (N8392, N8390);
xor XOR2 (N8393, N8384, N4833);
or OR3 (N8394, N8371, N3325, N6138);
nand NAND4 (N8395, N8392, N7074, N1009, N4774);
and AND3 (N8396, N8385, N7224, N2105);
and AND2 (N8397, N8387, N5726);
nand NAND2 (N8398, N8395, N7935);
nor NOR4 (N8399, N8391, N7641, N6974, N7423);
and AND4 (N8400, N8396, N2705, N225, N6900);
xor XOR2 (N8401, N8398, N2290);
or OR3 (N8402, N8394, N8394, N3101);
nor NOR4 (N8403, N8393, N8174, N3806, N5779);
nand NAND3 (N8404, N8401, N5513, N152);
buf BUF1 (N8405, N8388);
xor XOR2 (N8406, N8399, N4430);
buf BUF1 (N8407, N8402);
and AND4 (N8408, N8407, N4173, N7758, N7126);
or OR2 (N8409, N8365, N2813);
buf BUF1 (N8410, N8406);
nand NAND3 (N8411, N8405, N7641, N4997);
or OR4 (N8412, N8373, N2299, N6480, N663);
xor XOR2 (N8413, N8410, N2887);
and AND2 (N8414, N8400, N6041);
not NOT1 (N8415, N8404);
xor XOR2 (N8416, N8389, N1708);
or OR3 (N8417, N8413, N2212, N2963);
buf BUF1 (N8418, N8415);
not NOT1 (N8419, N8411);
nand NAND4 (N8420, N8417, N3398, N2381, N5443);
or OR4 (N8421, N8420, N2041, N5167, N6575);
not NOT1 (N8422, N8408);
xor XOR2 (N8423, N8403, N1044);
or OR3 (N8424, N8418, N3946, N4346);
xor XOR2 (N8425, N8397, N5997);
nor NOR2 (N8426, N8425, N5920);
nand NAND4 (N8427, N8409, N583, N4380, N6849);
or OR2 (N8428, N8421, N1966);
and AND2 (N8429, N8416, N5948);
nand NAND2 (N8430, N8422, N7893);
xor XOR2 (N8431, N8423, N6245);
and AND2 (N8432, N8424, N5428);
nand NAND4 (N8433, N8419, N5641, N4903, N4419);
nor NOR3 (N8434, N8433, N2384, N3866);
buf BUF1 (N8435, N8414);
nand NAND2 (N8436, N8434, N3424);
buf BUF1 (N8437, N8412);
xor XOR2 (N8438, N8431, N4226);
or OR3 (N8439, N8429, N2888, N5655);
buf BUF1 (N8440, N8427);
xor XOR2 (N8441, N8430, N6032);
or OR2 (N8442, N8440, N8043);
nor NOR2 (N8443, N8426, N1303);
nor NOR3 (N8444, N8435, N4860, N7686);
and AND2 (N8445, N8428, N7504);
not NOT1 (N8446, N8436);
not NOT1 (N8447, N8438);
nand NAND2 (N8448, N8432, N8043);
nand NAND2 (N8449, N8437, N1933);
or OR3 (N8450, N8445, N178, N7866);
nor NOR2 (N8451, N8443, N4210);
or OR4 (N8452, N8444, N2032, N3517, N1555);
or OR4 (N8453, N8447, N3929, N7810, N1508);
xor XOR2 (N8454, N8442, N7534);
nor NOR3 (N8455, N8450, N7358, N5397);
buf BUF1 (N8456, N8449);
xor XOR2 (N8457, N8448, N2196);
buf BUF1 (N8458, N8455);
xor XOR2 (N8459, N8458, N1555);
and AND4 (N8460, N8456, N2777, N5725, N7040);
not NOT1 (N8461, N8457);
not NOT1 (N8462, N8459);
and AND4 (N8463, N8451, N5816, N6767, N77);
not NOT1 (N8464, N8460);
buf BUF1 (N8465, N8454);
nand NAND3 (N8466, N8464, N3240, N1063);
nand NAND2 (N8467, N8465, N4604);
and AND3 (N8468, N8441, N8265, N7585);
or OR3 (N8469, N8466, N8320, N7456);
nand NAND2 (N8470, N8446, N7973);
xor XOR2 (N8471, N8470, N8234);
nand NAND4 (N8472, N8439, N2694, N4884, N6958);
not NOT1 (N8473, N8461);
or OR2 (N8474, N8467, N7288);
nand NAND4 (N8475, N8468, N4395, N1306, N993);
or OR3 (N8476, N8462, N5321, N7284);
xor XOR2 (N8477, N8472, N194);
and AND2 (N8478, N8453, N3190);
or OR3 (N8479, N8473, N8336, N4997);
xor XOR2 (N8480, N8452, N7278);
buf BUF1 (N8481, N8479);
or OR2 (N8482, N8476, N3167);
nand NAND2 (N8483, N8463, N3877);
xor XOR2 (N8484, N8471, N6505);
buf BUF1 (N8485, N8478);
and AND2 (N8486, N8469, N1478);
not NOT1 (N8487, N8474);
nor NOR4 (N8488, N8483, N4992, N4838, N7114);
or OR3 (N8489, N8477, N8064, N4884);
buf BUF1 (N8490, N8481);
nor NOR4 (N8491, N8480, N2861, N5235, N2825);
buf BUF1 (N8492, N8486);
and AND4 (N8493, N8490, N4587, N6170, N2668);
nand NAND4 (N8494, N8492, N6722, N5256, N7921);
and AND3 (N8495, N8475, N636, N4036);
buf BUF1 (N8496, N8491);
and AND4 (N8497, N8493, N441, N5524, N3090);
nand NAND4 (N8498, N8485, N2341, N3710, N591);
nor NOR4 (N8499, N8495, N1297, N5771, N1809);
nand NAND4 (N8500, N8484, N5007, N6548, N7766);
or OR3 (N8501, N8500, N2271, N8385);
and AND4 (N8502, N8499, N1736, N5829, N3132);
or OR2 (N8503, N8496, N6825);
nand NAND3 (N8504, N8489, N5667, N2937);
buf BUF1 (N8505, N8502);
buf BUF1 (N8506, N8488);
buf BUF1 (N8507, N8501);
buf BUF1 (N8508, N8506);
nand NAND4 (N8509, N8482, N2030, N1680, N732);
xor XOR2 (N8510, N8498, N2950);
xor XOR2 (N8511, N8504, N4087);
nor NOR2 (N8512, N8487, N4270);
or OR3 (N8513, N8510, N2718, N6853);
not NOT1 (N8514, N8503);
not NOT1 (N8515, N8507);
not NOT1 (N8516, N8494);
xor XOR2 (N8517, N8514, N1233);
nand NAND3 (N8518, N8497, N4964, N7235);
or OR4 (N8519, N8518, N1860, N2470, N7550);
and AND4 (N8520, N8509, N4630, N607, N4240);
not NOT1 (N8521, N8508);
xor XOR2 (N8522, N8521, N7427);
buf BUF1 (N8523, N8520);
or OR4 (N8524, N8515, N3556, N8055, N5949);
nand NAND2 (N8525, N8523, N4796);
xor XOR2 (N8526, N8522, N5279);
buf BUF1 (N8527, N8524);
and AND2 (N8528, N8519, N2386);
buf BUF1 (N8529, N8517);
nand NAND3 (N8530, N8526, N1668, N7925);
nor NOR2 (N8531, N8513, N2442);
not NOT1 (N8532, N8530);
not NOT1 (N8533, N8525);
xor XOR2 (N8534, N8531, N4212);
and AND2 (N8535, N8532, N7244);
nor NOR2 (N8536, N8511, N2072);
not NOT1 (N8537, N8505);
nor NOR4 (N8538, N8512, N8415, N7532, N1339);
nand NAND4 (N8539, N8527, N389, N122, N7134);
not NOT1 (N8540, N8529);
not NOT1 (N8541, N8534);
nand NAND2 (N8542, N8538, N7917);
nor NOR3 (N8543, N8537, N2307, N265);
xor XOR2 (N8544, N8539, N7733);
xor XOR2 (N8545, N8541, N4089);
nor NOR3 (N8546, N8542, N2918, N4227);
not NOT1 (N8547, N8545);
nor NOR3 (N8548, N8535, N2096, N7194);
not NOT1 (N8549, N8547);
nand NAND4 (N8550, N8540, N4399, N148, N6583);
nand NAND4 (N8551, N8544, N3479, N4730, N4645);
nor NOR2 (N8552, N8533, N1148);
or OR2 (N8553, N8516, N1249);
nand NAND4 (N8554, N8528, N125, N428, N7695);
and AND3 (N8555, N8548, N8052, N6832);
xor XOR2 (N8556, N8536, N2825);
not NOT1 (N8557, N8553);
not NOT1 (N8558, N8549);
buf BUF1 (N8559, N8550);
not NOT1 (N8560, N8559);
nand NAND4 (N8561, N8543, N6984, N1867, N5901);
nor NOR2 (N8562, N8552, N2434);
xor XOR2 (N8563, N8561, N1030);
xor XOR2 (N8564, N8556, N5628);
nor NOR3 (N8565, N8563, N5429, N5274);
nor NOR2 (N8566, N8546, N2027);
nor NOR2 (N8567, N8564, N548);
not NOT1 (N8568, N8565);
xor XOR2 (N8569, N8557, N8517);
and AND3 (N8570, N8566, N3491, N7008);
nand NAND2 (N8571, N8569, N1595);
buf BUF1 (N8572, N8551);
and AND4 (N8573, N8570, N6185, N8249, N3042);
nor NOR4 (N8574, N8568, N4647, N2925, N393);
and AND3 (N8575, N8562, N7118, N4505);
nor NOR3 (N8576, N8560, N7471, N2686);
xor XOR2 (N8577, N8576, N5983);
buf BUF1 (N8578, N8573);
buf BUF1 (N8579, N8555);
not NOT1 (N8580, N8571);
buf BUF1 (N8581, N8579);
and AND4 (N8582, N8567, N2881, N6173, N581);
nand NAND2 (N8583, N8580, N7672);
or OR4 (N8584, N8574, N8398, N7011, N7485);
nor NOR3 (N8585, N8558, N8385, N8301);
nor NOR4 (N8586, N8575, N7703, N428, N3810);
and AND4 (N8587, N8582, N3739, N6219, N5971);
nand NAND3 (N8588, N8581, N7549, N891);
or OR2 (N8589, N8572, N2496);
nor NOR3 (N8590, N8585, N2260, N5527);
nor NOR2 (N8591, N8578, N7189);
nand NAND2 (N8592, N8577, N6975);
xor XOR2 (N8593, N8586, N8275);
or OR4 (N8594, N8590, N5706, N8232, N2737);
nor NOR3 (N8595, N8588, N2406, N142);
or OR4 (N8596, N8589, N3971, N96, N6110);
buf BUF1 (N8597, N8594);
xor XOR2 (N8598, N8596, N7444);
nand NAND4 (N8599, N8593, N5581, N6349, N5903);
not NOT1 (N8600, N8591);
buf BUF1 (N8601, N8554);
or OR4 (N8602, N8599, N5754, N5894, N6862);
or OR3 (N8603, N8602, N1303, N2627);
xor XOR2 (N8604, N8584, N7661);
buf BUF1 (N8605, N8604);
nor NOR4 (N8606, N8583, N1405, N3788, N4321);
or OR2 (N8607, N8605, N5572);
buf BUF1 (N8608, N8597);
or OR2 (N8609, N8587, N815);
and AND2 (N8610, N8608, N5887);
and AND4 (N8611, N8595, N2369, N7368, N4976);
xor XOR2 (N8612, N8611, N2116);
and AND3 (N8613, N8598, N6108, N617);
nor NOR3 (N8614, N8601, N7698, N5098);
xor XOR2 (N8615, N8606, N8227);
nand NAND2 (N8616, N8612, N4926);
buf BUF1 (N8617, N8607);
nand NAND3 (N8618, N8614, N3248, N2060);
nand NAND3 (N8619, N8618, N640, N4457);
buf BUF1 (N8620, N8609);
or OR4 (N8621, N8600, N4353, N960, N2394);
nor NOR2 (N8622, N8615, N4152);
nand NAND4 (N8623, N8613, N1551, N3887, N5680);
buf BUF1 (N8624, N8619);
buf BUF1 (N8625, N8617);
and AND2 (N8626, N8620, N6822);
and AND2 (N8627, N8616, N6145);
buf BUF1 (N8628, N8610);
buf BUF1 (N8629, N8603);
nand NAND2 (N8630, N8629, N1690);
not NOT1 (N8631, N8623);
and AND3 (N8632, N8625, N1423, N2944);
and AND3 (N8633, N8626, N3081, N1532);
and AND4 (N8634, N8621, N4065, N3761, N8616);
xor XOR2 (N8635, N8624, N1785);
nand NAND3 (N8636, N8630, N535, N8468);
xor XOR2 (N8637, N8627, N746);
xor XOR2 (N8638, N8632, N2670);
or OR4 (N8639, N8631, N1320, N4249, N2946);
and AND4 (N8640, N8636, N2541, N4796, N6762);
not NOT1 (N8641, N8592);
or OR4 (N8642, N8633, N6480, N7227, N4642);
nand NAND3 (N8643, N8622, N7362, N4426);
and AND2 (N8644, N8635, N5725);
nor NOR4 (N8645, N8642, N6793, N3858, N4965);
xor XOR2 (N8646, N8640, N2843);
or OR4 (N8647, N8638, N2180, N4443, N839);
xor XOR2 (N8648, N8643, N2302);
xor XOR2 (N8649, N8646, N4251);
or OR4 (N8650, N8634, N8212, N3686, N8366);
not NOT1 (N8651, N8628);
and AND2 (N8652, N8649, N4121);
xor XOR2 (N8653, N8637, N2595);
nor NOR4 (N8654, N8648, N3733, N6552, N1252);
and AND3 (N8655, N8654, N4816, N7833);
nand NAND2 (N8656, N8650, N547);
nand NAND4 (N8657, N8645, N4308, N4103, N2618);
not NOT1 (N8658, N8647);
and AND2 (N8659, N8644, N780);
nand NAND3 (N8660, N8653, N1770, N3700);
and AND2 (N8661, N8655, N7838);
and AND2 (N8662, N8656, N1625);
or OR4 (N8663, N8659, N5991, N7430, N3092);
and AND2 (N8664, N8652, N5967);
buf BUF1 (N8665, N8641);
xor XOR2 (N8666, N8661, N2010);
buf BUF1 (N8667, N8662);
nand NAND2 (N8668, N8657, N911);
nor NOR3 (N8669, N8660, N5017, N61);
xor XOR2 (N8670, N8668, N5691);
buf BUF1 (N8671, N8651);
or OR2 (N8672, N8663, N4377);
buf BUF1 (N8673, N8666);
or OR3 (N8674, N8673, N4401, N4416);
nand NAND2 (N8675, N8664, N2727);
and AND3 (N8676, N8670, N8400, N8257);
nor NOR2 (N8677, N8639, N6894);
and AND4 (N8678, N8665, N100, N7599, N6140);
nor NOR2 (N8679, N8678, N6038);
or OR2 (N8680, N8679, N256);
and AND3 (N8681, N8672, N2208, N8332);
not NOT1 (N8682, N8681);
not NOT1 (N8683, N8676);
or OR2 (N8684, N8658, N8414);
or OR3 (N8685, N8675, N509, N1705);
or OR4 (N8686, N8669, N2947, N8647, N4784);
or OR4 (N8687, N8684, N4270, N3710, N677);
and AND3 (N8688, N8680, N180, N3945);
nor NOR2 (N8689, N8687, N1488);
or OR2 (N8690, N8667, N5825);
and AND3 (N8691, N8685, N4653, N5083);
nor NOR2 (N8692, N8689, N7915);
buf BUF1 (N8693, N8691);
nand NAND3 (N8694, N8682, N5267, N5998);
xor XOR2 (N8695, N8683, N4511);
not NOT1 (N8696, N8671);
not NOT1 (N8697, N8693);
buf BUF1 (N8698, N8690);
xor XOR2 (N8699, N8696, N6298);
nor NOR4 (N8700, N8686, N5571, N7824, N8267);
not NOT1 (N8701, N8700);
not NOT1 (N8702, N8701);
and AND2 (N8703, N8674, N5864);
not NOT1 (N8704, N8695);
nand NAND3 (N8705, N8677, N1376, N5734);
nor NOR4 (N8706, N8688, N1570, N3917, N2152);
nand NAND3 (N8707, N8699, N2193, N1344);
or OR3 (N8708, N8702, N5568, N5146);
or OR2 (N8709, N8704, N5898);
xor XOR2 (N8710, N8697, N2149);
xor XOR2 (N8711, N8694, N3929);
xor XOR2 (N8712, N8705, N7435);
and AND4 (N8713, N8709, N6746, N264, N6481);
and AND3 (N8714, N8711, N4586, N1536);
nor NOR3 (N8715, N8707, N8353, N3254);
and AND3 (N8716, N8708, N5062, N4158);
nand NAND3 (N8717, N8710, N5795, N7351);
nor NOR4 (N8718, N8698, N6813, N6541, N1925);
not NOT1 (N8719, N8713);
nor NOR2 (N8720, N8706, N1535);
nor NOR2 (N8721, N8712, N5139);
nand NAND2 (N8722, N8715, N8230);
not NOT1 (N8723, N8703);
not NOT1 (N8724, N8721);
not NOT1 (N8725, N8720);
and AND4 (N8726, N8722, N1392, N4665, N4221);
nor NOR3 (N8727, N8718, N23, N6334);
nand NAND2 (N8728, N8717, N8109);
and AND2 (N8729, N8719, N4753);
nand NAND3 (N8730, N8723, N5123, N4029);
buf BUF1 (N8731, N8714);
buf BUF1 (N8732, N8728);
nand NAND3 (N8733, N8724, N4673, N7747);
not NOT1 (N8734, N8726);
xor XOR2 (N8735, N8733, N6822);
nand NAND4 (N8736, N8729, N4153, N5693, N675);
or OR2 (N8737, N8727, N3977);
or OR4 (N8738, N8732, N2887, N4253, N8311);
and AND3 (N8739, N8736, N4295, N1807);
not NOT1 (N8740, N8739);
or OR4 (N8741, N8730, N3098, N4858, N8032);
and AND2 (N8742, N8738, N2948);
xor XOR2 (N8743, N8716, N432);
xor XOR2 (N8744, N8743, N2167);
nor NOR4 (N8745, N8692, N5403, N7549, N4943);
nor NOR3 (N8746, N8734, N7754, N4454);
or OR2 (N8747, N8746, N5289);
or OR3 (N8748, N8725, N2467, N476);
nor NOR4 (N8749, N8744, N7872, N2503, N2263);
and AND4 (N8750, N8731, N600, N6455, N2015);
nor NOR4 (N8751, N8745, N1487, N6129, N2799);
and AND2 (N8752, N8741, N336);
not NOT1 (N8753, N8737);
nor NOR4 (N8754, N8749, N267, N8550, N4879);
and AND3 (N8755, N8752, N5019, N4183);
buf BUF1 (N8756, N8753);
nand NAND2 (N8757, N8750, N5993);
not NOT1 (N8758, N8757);
or OR4 (N8759, N8751, N93, N3945, N4827);
nand NAND4 (N8760, N8747, N4276, N1974, N198);
nor NOR4 (N8761, N8735, N6811, N3987, N6730);
nor NOR4 (N8762, N8761, N6872, N2012, N7151);
or OR2 (N8763, N8756, N8402);
nand NAND2 (N8764, N8759, N1193);
or OR4 (N8765, N8762, N3270, N2267, N1289);
nand NAND2 (N8766, N8763, N5766);
xor XOR2 (N8767, N8765, N5918);
and AND2 (N8768, N8754, N3831);
xor XOR2 (N8769, N8758, N6370);
nand NAND3 (N8770, N8748, N7070, N3744);
nor NOR2 (N8771, N8768, N641);
and AND4 (N8772, N8770, N3992, N6664, N7661);
nand NAND2 (N8773, N8740, N2423);
nor NOR3 (N8774, N8764, N3329, N6405);
nor NOR4 (N8775, N8742, N2754, N978, N1395);
xor XOR2 (N8776, N8774, N885);
nand NAND3 (N8777, N8769, N2766, N23);
buf BUF1 (N8778, N8766);
or OR4 (N8779, N8776, N1927, N7172, N1598);
nand NAND2 (N8780, N8773, N8051);
nand NAND4 (N8781, N8780, N7591, N160, N3320);
or OR4 (N8782, N8771, N479, N2806, N6940);
nand NAND3 (N8783, N8755, N917, N7889);
nor NOR4 (N8784, N8782, N416, N5210, N2693);
nand NAND4 (N8785, N8779, N1379, N4428, N6426);
and AND4 (N8786, N8772, N4289, N7228, N2114);
not NOT1 (N8787, N8767);
or OR3 (N8788, N8785, N4292, N3503);
not NOT1 (N8789, N8787);
nand NAND2 (N8790, N8786, N8511);
nor NOR4 (N8791, N8783, N3842, N6442, N7919);
nor NOR3 (N8792, N8790, N321, N5915);
not NOT1 (N8793, N8788);
and AND4 (N8794, N8781, N2615, N69, N7636);
not NOT1 (N8795, N8791);
buf BUF1 (N8796, N8760);
nor NOR4 (N8797, N8796, N8543, N7722, N3272);
not NOT1 (N8798, N8793);
and AND2 (N8799, N8784, N602);
nand NAND3 (N8800, N8795, N1431, N4957);
not NOT1 (N8801, N8800);
and AND2 (N8802, N8778, N7701);
and AND4 (N8803, N8775, N874, N2949, N7184);
xor XOR2 (N8804, N8792, N747);
not NOT1 (N8805, N8801);
xor XOR2 (N8806, N8804, N1286);
or OR4 (N8807, N8789, N1196, N174, N7006);
or OR2 (N8808, N8805, N7791);
nand NAND2 (N8809, N8798, N3110);
nor NOR2 (N8810, N8777, N8510);
nand NAND4 (N8811, N8806, N4080, N3402, N4139);
or OR2 (N8812, N8810, N1877);
not NOT1 (N8813, N8794);
xor XOR2 (N8814, N8802, N8351);
nor NOR4 (N8815, N8812, N4455, N3613, N7999);
not NOT1 (N8816, N8813);
buf BUF1 (N8817, N8809);
nand NAND3 (N8818, N8817, N3153, N2510);
or OR2 (N8819, N8811, N5439);
buf BUF1 (N8820, N8819);
and AND4 (N8821, N8799, N1084, N3924, N7558);
and AND4 (N8822, N8816, N1988, N4324, N3590);
xor XOR2 (N8823, N8815, N5765);
nand NAND4 (N8824, N8818, N1234, N3477, N2364);
nor NOR4 (N8825, N8807, N8052, N3727, N7649);
buf BUF1 (N8826, N8808);
buf BUF1 (N8827, N8825);
or OR4 (N8828, N8822, N2329, N4037, N7773);
buf BUF1 (N8829, N8824);
and AND2 (N8830, N8803, N7964);
nor NOR3 (N8831, N8828, N5676, N5555);
and AND2 (N8832, N8831, N765);
xor XOR2 (N8833, N8797, N1610);
nand NAND2 (N8834, N8829, N3370);
and AND4 (N8835, N8814, N6948, N4167, N6037);
nand NAND4 (N8836, N8821, N7434, N2603, N622);
not NOT1 (N8837, N8832);
not NOT1 (N8838, N8820);
xor XOR2 (N8839, N8826, N372);
or OR3 (N8840, N8838, N8437, N1049);
nand NAND4 (N8841, N8823, N2766, N5662, N8014);
nor NOR2 (N8842, N8833, N2038);
xor XOR2 (N8843, N8841, N4677);
nand NAND4 (N8844, N8837, N3711, N7619, N3607);
or OR4 (N8845, N8843, N3361, N6943, N2536);
and AND4 (N8846, N8842, N7888, N3473, N996);
buf BUF1 (N8847, N8830);
nand NAND3 (N8848, N8834, N2462, N8233);
xor XOR2 (N8849, N8840, N571);
nand NAND3 (N8850, N8846, N1343, N6551);
xor XOR2 (N8851, N8839, N2333);
xor XOR2 (N8852, N8849, N4064);
or OR4 (N8853, N8848, N7752, N8805, N6262);
and AND2 (N8854, N8847, N6432);
buf BUF1 (N8855, N8850);
nand NAND3 (N8856, N8835, N8105, N3371);
buf BUF1 (N8857, N8844);
not NOT1 (N8858, N8854);
not NOT1 (N8859, N8851);
and AND3 (N8860, N8852, N2419, N4872);
or OR2 (N8861, N8855, N8070);
xor XOR2 (N8862, N8860, N2043);
nor NOR4 (N8863, N8845, N3702, N1349, N4886);
and AND4 (N8864, N8853, N7713, N1820, N8717);
not NOT1 (N8865, N8836);
nor NOR4 (N8866, N8858, N6689, N6932, N5303);
nand NAND2 (N8867, N8864, N1609);
buf BUF1 (N8868, N8827);
nor NOR2 (N8869, N8865, N4935);
buf BUF1 (N8870, N8862);
nor NOR2 (N8871, N8866, N29);
not NOT1 (N8872, N8857);
or OR2 (N8873, N8869, N4003);
xor XOR2 (N8874, N8867, N3491);
not NOT1 (N8875, N8871);
not NOT1 (N8876, N8875);
nand NAND2 (N8877, N8876, N1351);
nand NAND4 (N8878, N8874, N183, N7845, N3618);
not NOT1 (N8879, N8861);
or OR2 (N8880, N8870, N4359);
and AND2 (N8881, N8873, N2174);
buf BUF1 (N8882, N8863);
buf BUF1 (N8883, N8881);
xor XOR2 (N8884, N8859, N1763);
and AND3 (N8885, N8879, N48, N8328);
or OR2 (N8886, N8882, N4723);
buf BUF1 (N8887, N8883);
not NOT1 (N8888, N8880);
nor NOR3 (N8889, N8868, N6769, N3057);
buf BUF1 (N8890, N8878);
not NOT1 (N8891, N8877);
buf BUF1 (N8892, N8884);
not NOT1 (N8893, N8891);
nand NAND3 (N8894, N8892, N5025, N5801);
not NOT1 (N8895, N8893);
xor XOR2 (N8896, N8888, N3097);
nor NOR2 (N8897, N8885, N6633);
not NOT1 (N8898, N8856);
nand NAND3 (N8899, N8897, N7596, N5897);
nand NAND4 (N8900, N8895, N398, N3487, N349);
not NOT1 (N8901, N8887);
not NOT1 (N8902, N8889);
and AND2 (N8903, N8898, N4174);
and AND3 (N8904, N8872, N6221, N2685);
xor XOR2 (N8905, N8903, N185);
nor NOR3 (N8906, N8886, N6782, N7778);
not NOT1 (N8907, N8902);
nor NOR4 (N8908, N8901, N715, N2537, N2434);
nand NAND4 (N8909, N8906, N3806, N7139, N3117);
or OR4 (N8910, N8904, N7942, N714, N5461);
or OR4 (N8911, N8890, N1784, N7132, N4393);
and AND4 (N8912, N8908, N5802, N7487, N7062);
xor XOR2 (N8913, N8910, N5076);
buf BUF1 (N8914, N8912);
or OR4 (N8915, N8911, N1629, N3174, N4139);
nand NAND4 (N8916, N8894, N4103, N5771, N2525);
or OR2 (N8917, N8913, N223);
nand NAND2 (N8918, N8900, N4221);
buf BUF1 (N8919, N8914);
not NOT1 (N8920, N8915);
buf BUF1 (N8921, N8896);
or OR3 (N8922, N8916, N984, N441);
xor XOR2 (N8923, N8899, N1721);
xor XOR2 (N8924, N8909, N1682);
and AND2 (N8925, N8924, N4117);
xor XOR2 (N8926, N8925, N4363);
nand NAND2 (N8927, N8919, N512);
not NOT1 (N8928, N8921);
and AND2 (N8929, N8905, N3517);
buf BUF1 (N8930, N8917);
nor NOR2 (N8931, N8926, N2998);
xor XOR2 (N8932, N8930, N2909);
xor XOR2 (N8933, N8927, N1068);
xor XOR2 (N8934, N8923, N356);
and AND3 (N8935, N8928, N1955, N8508);
nand NAND3 (N8936, N8931, N4834, N54);
nand NAND3 (N8937, N8935, N2251, N1277);
xor XOR2 (N8938, N8920, N340);
or OR3 (N8939, N8933, N329, N5636);
nor NOR2 (N8940, N8936, N7240);
and AND4 (N8941, N8934, N1889, N8312, N8448);
and AND3 (N8942, N8929, N3272, N1496);
xor XOR2 (N8943, N8940, N4983);
nor NOR4 (N8944, N8937, N7578, N5136, N2984);
and AND2 (N8945, N8939, N5115);
nor NOR2 (N8946, N8932, N1662);
nor NOR4 (N8947, N8946, N8761, N4465, N2815);
nand NAND2 (N8948, N8941, N7004);
and AND3 (N8949, N8918, N1954, N775);
or OR4 (N8950, N8944, N1729, N3353, N6066);
xor XOR2 (N8951, N8948, N5885);
nor NOR4 (N8952, N8938, N3345, N5721, N1576);
buf BUF1 (N8953, N8922);
and AND4 (N8954, N8951, N7192, N5010, N6314);
buf BUF1 (N8955, N8949);
nor NOR2 (N8956, N8943, N7192);
and AND2 (N8957, N8952, N8648);
and AND3 (N8958, N8957, N8496, N5506);
and AND3 (N8959, N8942, N4679, N4692);
or OR3 (N8960, N8947, N6863, N3473);
xor XOR2 (N8961, N8958, N4109);
not NOT1 (N8962, N8950);
xor XOR2 (N8963, N8945, N7995);
and AND4 (N8964, N8959, N3109, N4717, N6473);
and AND2 (N8965, N8964, N3155);
nor NOR2 (N8966, N8953, N8536);
not NOT1 (N8967, N8956);
or OR4 (N8968, N8960, N3691, N951, N6684);
xor XOR2 (N8969, N8962, N4181);
xor XOR2 (N8970, N8907, N6707);
or OR2 (N8971, N8970, N2441);
not NOT1 (N8972, N8965);
nor NOR2 (N8973, N8963, N3361);
and AND4 (N8974, N8954, N5821, N4535, N4147);
nand NAND4 (N8975, N8961, N3039, N7892, N372);
or OR2 (N8976, N8969, N3698);
or OR2 (N8977, N8967, N4695);
and AND4 (N8978, N8971, N4544, N4387, N8458);
or OR2 (N8979, N8955, N4069);
and AND3 (N8980, N8974, N936, N5535);
and AND4 (N8981, N8976, N5517, N434, N7101);
not NOT1 (N8982, N8979);
and AND2 (N8983, N8966, N8606);
not NOT1 (N8984, N8983);
and AND2 (N8985, N8968, N5338);
xor XOR2 (N8986, N8978, N7316);
nor NOR2 (N8987, N8981, N7441);
buf BUF1 (N8988, N8977);
xor XOR2 (N8989, N8986, N771);
xor XOR2 (N8990, N8980, N5496);
nand NAND3 (N8991, N8984, N4944, N5564);
or OR4 (N8992, N8982, N4337, N861, N3734);
buf BUF1 (N8993, N8975);
xor XOR2 (N8994, N8990, N8244);
and AND3 (N8995, N8989, N5821, N285);
and AND4 (N8996, N8973, N2106, N3162, N8769);
nand NAND4 (N8997, N8995, N194, N6521, N6339);
buf BUF1 (N8998, N8993);
buf BUF1 (N8999, N8991);
nand NAND2 (N9000, N8994, N816);
nand NAND3 (N9001, N8999, N8513, N6195);
and AND2 (N9002, N8998, N6558);
buf BUF1 (N9003, N9001);
nand NAND3 (N9004, N8996, N7357, N6468);
or OR4 (N9005, N8997, N2558, N2938, N6745);
not NOT1 (N9006, N8985);
buf BUF1 (N9007, N8988);
nand NAND3 (N9008, N9007, N1691, N2760);
and AND4 (N9009, N8972, N7914, N8555, N7963);
and AND2 (N9010, N9004, N1344);
xor XOR2 (N9011, N9006, N1355);
xor XOR2 (N9012, N9009, N3208);
xor XOR2 (N9013, N9010, N8480);
nand NAND4 (N9014, N9003, N6120, N4832, N380);
buf BUF1 (N9015, N9008);
or OR2 (N9016, N9011, N8863);
not NOT1 (N9017, N8987);
xor XOR2 (N9018, N9014, N7248);
buf BUF1 (N9019, N9002);
nor NOR3 (N9020, N9015, N5820, N4661);
and AND3 (N9021, N9013, N685, N5894);
nand NAND3 (N9022, N9012, N2901, N4256);
nand NAND2 (N9023, N9020, N8176);
nor NOR3 (N9024, N9023, N2936, N2868);
buf BUF1 (N9025, N9021);
or OR2 (N9026, N8992, N3714);
buf BUF1 (N9027, N9018);
xor XOR2 (N9028, N9025, N4891);
xor XOR2 (N9029, N9019, N1423);
xor XOR2 (N9030, N9000, N6100);
nand NAND3 (N9031, N9030, N5887, N7773);
nor NOR2 (N9032, N9031, N7640);
nor NOR2 (N9033, N9032, N176);
or OR3 (N9034, N9005, N8677, N7654);
nor NOR4 (N9035, N9022, N8066, N3387, N688);
nor NOR4 (N9036, N9029, N1436, N201, N3348);
nor NOR3 (N9037, N9024, N3700, N5317);
xor XOR2 (N9038, N9033, N4658);
and AND3 (N9039, N9034, N6822, N4119);
xor XOR2 (N9040, N9038, N6551);
buf BUF1 (N9041, N9036);
and AND2 (N9042, N9037, N2821);
xor XOR2 (N9043, N9028, N2715);
nand NAND4 (N9044, N9017, N166, N4995, N7754);
nand NAND4 (N9045, N9035, N3058, N686, N5774);
and AND3 (N9046, N9042, N3830, N5300);
xor XOR2 (N9047, N9027, N4353);
nor NOR2 (N9048, N9016, N7729);
or OR2 (N9049, N9044, N2465);
and AND2 (N9050, N9039, N957);
nand NAND2 (N9051, N9049, N4476);
nand NAND4 (N9052, N9050, N3814, N607, N3840);
xor XOR2 (N9053, N9043, N8647);
not NOT1 (N9054, N9040);
not NOT1 (N9055, N9047);
xor XOR2 (N9056, N9053, N6112);
not NOT1 (N9057, N9048);
nand NAND4 (N9058, N9054, N5443, N4530, N1542);
not NOT1 (N9059, N9041);
or OR3 (N9060, N9045, N7410, N4778);
and AND2 (N9061, N9060, N1291);
xor XOR2 (N9062, N9061, N2326);
xor XOR2 (N9063, N9056, N8981);
nor NOR3 (N9064, N9057, N1570, N3993);
or OR4 (N9065, N9051, N5375, N506, N3907);
nand NAND2 (N9066, N9055, N849);
not NOT1 (N9067, N9062);
and AND2 (N9068, N9052, N7925);
or OR2 (N9069, N9067, N5775);
buf BUF1 (N9070, N9059);
nand NAND3 (N9071, N9058, N2901, N3899);
buf BUF1 (N9072, N9069);
or OR2 (N9073, N9046, N6480);
or OR3 (N9074, N9066, N1232, N2937);
and AND4 (N9075, N9064, N846, N4779, N5305);
or OR2 (N9076, N9071, N8116);
and AND2 (N9077, N9073, N6388);
not NOT1 (N9078, N9072);
buf BUF1 (N9079, N9026);
xor XOR2 (N9080, N9078, N8876);
xor XOR2 (N9081, N9063, N5234);
or OR4 (N9082, N9075, N2188, N2333, N4644);
not NOT1 (N9083, N9068);
or OR4 (N9084, N9076, N60, N3914, N8113);
not NOT1 (N9085, N9083);
not NOT1 (N9086, N9085);
nand NAND3 (N9087, N9074, N9063, N4589);
nor NOR4 (N9088, N9077, N708, N3180, N3323);
and AND2 (N9089, N9080, N1601);
not NOT1 (N9090, N9086);
nand NAND3 (N9091, N9090, N4427, N4782);
xor XOR2 (N9092, N9084, N7186);
nor NOR2 (N9093, N9082, N4997);
xor XOR2 (N9094, N9092, N5836);
and AND2 (N9095, N9087, N8424);
not NOT1 (N9096, N9091);
xor XOR2 (N9097, N9096, N2142);
not NOT1 (N9098, N9089);
not NOT1 (N9099, N9095);
or OR4 (N9100, N9094, N4041, N1295, N2600);
not NOT1 (N9101, N9079);
nor NOR3 (N9102, N9088, N5560, N1608);
buf BUF1 (N9103, N9093);
or OR2 (N9104, N9100, N8419);
nand NAND3 (N9105, N9099, N3631, N1703);
and AND3 (N9106, N9098, N49, N7539);
xor XOR2 (N9107, N9081, N2248);
buf BUF1 (N9108, N9103);
buf BUF1 (N9109, N9107);
nand NAND4 (N9110, N9106, N4039, N8270, N2302);
and AND3 (N9111, N9110, N6492, N5707);
nand NAND4 (N9112, N9104, N2917, N6442, N1678);
buf BUF1 (N9113, N9108);
xor XOR2 (N9114, N9070, N2110);
or OR3 (N9115, N9065, N6920, N6380);
and AND3 (N9116, N9114, N4000, N4864);
or OR2 (N9117, N9097, N2939);
not NOT1 (N9118, N9115);
and AND3 (N9119, N9101, N5399, N752);
or OR2 (N9120, N9111, N4708);
or OR4 (N9121, N9109, N721, N5301, N5403);
nor NOR3 (N9122, N9102, N4428, N6301);
nor NOR3 (N9123, N9120, N351, N44);
nand NAND4 (N9124, N9122, N680, N4661, N5386);
buf BUF1 (N9125, N9117);
xor XOR2 (N9126, N9105, N1261);
nand NAND2 (N9127, N9123, N3182);
nor NOR4 (N9128, N9121, N4278, N6645, N7472);
nand NAND2 (N9129, N9113, N4871);
or OR3 (N9130, N9116, N89, N7153);
and AND4 (N9131, N9118, N1389, N7992, N2533);
buf BUF1 (N9132, N9126);
nand NAND4 (N9133, N9119, N1858, N6182, N6750);
xor XOR2 (N9134, N9131, N154);
nand NAND4 (N9135, N9129, N8145, N8872, N6227);
nor NOR4 (N9136, N9125, N7366, N5053, N6003);
or OR2 (N9137, N9135, N2255);
buf BUF1 (N9138, N9130);
buf BUF1 (N9139, N9137);
and AND3 (N9140, N9139, N3638, N2245);
not NOT1 (N9141, N9132);
nand NAND4 (N9142, N9136, N4455, N6934, N7568);
or OR2 (N9143, N9141, N8976);
buf BUF1 (N9144, N9124);
not NOT1 (N9145, N9127);
xor XOR2 (N9146, N9140, N3992);
buf BUF1 (N9147, N9145);
not NOT1 (N9148, N9147);
nor NOR2 (N9149, N9148, N3605);
not NOT1 (N9150, N9143);
nor NOR2 (N9151, N9133, N2141);
xor XOR2 (N9152, N9144, N8837);
not NOT1 (N9153, N9128);
nor NOR2 (N9154, N9150, N7534);
and AND4 (N9155, N9153, N2647, N3767, N3666);
not NOT1 (N9156, N9151);
not NOT1 (N9157, N9146);
xor XOR2 (N9158, N9155, N7424);
not NOT1 (N9159, N9154);
nor NOR2 (N9160, N9134, N3116);
nand NAND4 (N9161, N9152, N9126, N6055, N4090);
or OR4 (N9162, N9112, N6788, N2104, N7698);
or OR2 (N9163, N9161, N4551);
buf BUF1 (N9164, N9138);
buf BUF1 (N9165, N9164);
or OR2 (N9166, N9160, N6035);
buf BUF1 (N9167, N9149);
xor XOR2 (N9168, N9166, N948);
buf BUF1 (N9169, N9159);
nor NOR3 (N9170, N9168, N3886, N4228);
nor NOR2 (N9171, N9157, N3150);
buf BUF1 (N9172, N9158);
nor NOR4 (N9173, N9165, N4235, N1876, N4956);
or OR3 (N9174, N9162, N6447, N864);
or OR4 (N9175, N9173, N169, N5408, N2337);
or OR4 (N9176, N9169, N2873, N7516, N3836);
not NOT1 (N9177, N9156);
nor NOR2 (N9178, N9170, N4922);
or OR3 (N9179, N9172, N5319, N8869);
not NOT1 (N9180, N9142);
buf BUF1 (N9181, N9171);
not NOT1 (N9182, N9176);
or OR3 (N9183, N9182, N5412, N2107);
nand NAND2 (N9184, N9181, N822);
nand NAND3 (N9185, N9177, N64, N2616);
nor NOR2 (N9186, N9163, N2996);
nand NAND2 (N9187, N9178, N6887);
nor NOR4 (N9188, N9186, N8788, N5653, N88);
nand NAND4 (N9189, N9179, N8596, N2186, N8647);
xor XOR2 (N9190, N9188, N4863);
nor NOR4 (N9191, N9189, N7005, N8850, N6889);
or OR4 (N9192, N9180, N6028, N1034, N8994);
nor NOR4 (N9193, N9185, N7346, N6562, N2133);
xor XOR2 (N9194, N9192, N7487);
buf BUF1 (N9195, N9184);
not NOT1 (N9196, N9195);
xor XOR2 (N9197, N9194, N624);
not NOT1 (N9198, N9196);
or OR3 (N9199, N9190, N645, N6502);
or OR3 (N9200, N9193, N3048, N7530);
nand NAND4 (N9201, N9200, N1012, N3505, N36);
buf BUF1 (N9202, N9197);
or OR3 (N9203, N9167, N5213, N3548);
or OR2 (N9204, N9203, N463);
xor XOR2 (N9205, N9204, N3580);
nand NAND3 (N9206, N9198, N2100, N3381);
nand NAND4 (N9207, N9187, N9087, N5780, N8185);
nor NOR2 (N9208, N9205, N5508);
nand NAND2 (N9209, N9206, N6732);
buf BUF1 (N9210, N9183);
or OR4 (N9211, N9174, N8852, N5585, N3362);
nor NOR4 (N9212, N9207, N1400, N2020, N16);
nor NOR3 (N9213, N9210, N4363, N6704);
not NOT1 (N9214, N9202);
nand NAND2 (N9215, N9199, N682);
not NOT1 (N9216, N9209);
not NOT1 (N9217, N9211);
and AND4 (N9218, N9191, N4016, N6974, N7105);
or OR2 (N9219, N9212, N5240);
nor NOR4 (N9220, N9216, N2841, N4004, N2040);
or OR2 (N9221, N9214, N6478);
or OR3 (N9222, N9201, N910, N7944);
and AND3 (N9223, N9222, N6520, N5710);
nand NAND3 (N9224, N9219, N2441, N1620);
or OR2 (N9225, N9221, N5212);
nand NAND3 (N9226, N9215, N3692, N5203);
and AND4 (N9227, N9213, N1722, N6086, N6354);
nand NAND4 (N9228, N9175, N4991, N4995, N9004);
and AND4 (N9229, N9228, N7014, N6134, N320);
and AND3 (N9230, N9220, N2426, N235);
or OR3 (N9231, N9223, N9075, N1635);
not NOT1 (N9232, N9230);
not NOT1 (N9233, N9217);
nor NOR4 (N9234, N9232, N1071, N2291, N6207);
nand NAND2 (N9235, N9229, N7337);
not NOT1 (N9236, N9218);
buf BUF1 (N9237, N9236);
or OR3 (N9238, N9208, N3983, N5369);
nor NOR3 (N9239, N9235, N1467, N6882);
or OR3 (N9240, N9238, N642, N7598);
xor XOR2 (N9241, N9240, N7799);
not NOT1 (N9242, N9225);
and AND3 (N9243, N9226, N2466, N8574);
and AND4 (N9244, N9233, N2260, N1767, N6492);
buf BUF1 (N9245, N9237);
not NOT1 (N9246, N9244);
and AND4 (N9247, N9241, N1478, N9216, N6571);
nand NAND4 (N9248, N9231, N6947, N8572, N8288);
buf BUF1 (N9249, N9242);
not NOT1 (N9250, N9239);
or OR3 (N9251, N9234, N8464, N2460);
buf BUF1 (N9252, N9243);
xor XOR2 (N9253, N9249, N2762);
xor XOR2 (N9254, N9252, N6168);
and AND4 (N9255, N9227, N5336, N6862, N5396);
xor XOR2 (N9256, N9224, N7467);
or OR4 (N9257, N9251, N44, N5745, N3007);
buf BUF1 (N9258, N9250);
xor XOR2 (N9259, N9255, N4870);
nor NOR4 (N9260, N9254, N8976, N5503, N3140);
not NOT1 (N9261, N9245);
xor XOR2 (N9262, N9258, N2771);
and AND2 (N9263, N9248, N3102);
or OR2 (N9264, N9253, N8123);
and AND3 (N9265, N9264, N3801, N2447);
xor XOR2 (N9266, N9247, N7869);
xor XOR2 (N9267, N9266, N8109);
or OR4 (N9268, N9260, N7141, N6155, N2594);
xor XOR2 (N9269, N9265, N3860);
xor XOR2 (N9270, N9267, N3294);
and AND2 (N9271, N9256, N149);
nor NOR2 (N9272, N9270, N7858);
or OR3 (N9273, N9262, N5296, N3717);
buf BUF1 (N9274, N9263);
not NOT1 (N9275, N9261);
xor XOR2 (N9276, N9246, N2290);
nand NAND3 (N9277, N9275, N8424, N8654);
nor NOR3 (N9278, N9272, N8210, N617);
or OR3 (N9279, N9278, N392, N3144);
buf BUF1 (N9280, N9257);
buf BUF1 (N9281, N9280);
xor XOR2 (N9282, N9277, N7396);
buf BUF1 (N9283, N9271);
buf BUF1 (N9284, N9268);
xor XOR2 (N9285, N9284, N7940);
and AND3 (N9286, N9283, N1868, N458);
buf BUF1 (N9287, N9276);
nand NAND2 (N9288, N9269, N6656);
nand NAND4 (N9289, N9273, N504, N800, N8413);
buf BUF1 (N9290, N9282);
nor NOR4 (N9291, N9281, N5733, N5978, N9127);
xor XOR2 (N9292, N9259, N2718);
buf BUF1 (N9293, N9291);
not NOT1 (N9294, N9293);
nand NAND2 (N9295, N9279, N2355);
nor NOR3 (N9296, N9290, N3272, N5005);
and AND3 (N9297, N9295, N5075, N6162);
or OR2 (N9298, N9297, N5898);
not NOT1 (N9299, N9294);
xor XOR2 (N9300, N9298, N117);
or OR3 (N9301, N9287, N4979, N8743);
not NOT1 (N9302, N9299);
buf BUF1 (N9303, N9296);
and AND2 (N9304, N9300, N1399);
or OR2 (N9305, N9304, N2491);
nor NOR2 (N9306, N9292, N6888);
nand NAND3 (N9307, N9301, N5649, N3580);
not NOT1 (N9308, N9305);
or OR4 (N9309, N9307, N5468, N3172, N3088);
and AND3 (N9310, N9302, N2437, N3600);
nand NAND3 (N9311, N9308, N62, N1488);
xor XOR2 (N9312, N9286, N6252);
nor NOR2 (N9313, N9289, N6590);
or OR2 (N9314, N9313, N9080);
or OR3 (N9315, N9274, N3904, N3675);
nor NOR3 (N9316, N9315, N5549, N7128);
buf BUF1 (N9317, N9309);
buf BUF1 (N9318, N9303);
xor XOR2 (N9319, N9317, N6814);
buf BUF1 (N9320, N9306);
not NOT1 (N9321, N9310);
buf BUF1 (N9322, N9320);
or OR3 (N9323, N9318, N4872, N3732);
or OR3 (N9324, N9312, N3665, N8443);
and AND4 (N9325, N9285, N8408, N3561, N8939);
not NOT1 (N9326, N9325);
and AND3 (N9327, N9321, N4505, N1776);
nor NOR4 (N9328, N9311, N4687, N392, N1661);
xor XOR2 (N9329, N9326, N1130);
nand NAND4 (N9330, N9316, N4992, N3313, N4820);
nand NAND4 (N9331, N9314, N9028, N1194, N8171);
xor XOR2 (N9332, N9329, N9288);
buf BUF1 (N9333, N4035);
and AND2 (N9334, N9322, N1775);
buf BUF1 (N9335, N9332);
xor XOR2 (N9336, N9328, N952);
buf BUF1 (N9337, N9331);
nand NAND3 (N9338, N9336, N7825, N8419);
not NOT1 (N9339, N9324);
or OR3 (N9340, N9334, N1087, N4860);
xor XOR2 (N9341, N9323, N6871);
nand NAND3 (N9342, N9341, N6792, N2165);
nor NOR2 (N9343, N9342, N1146);
nand NAND2 (N9344, N9327, N6360);
nand NAND4 (N9345, N9343, N371, N5083, N617);
buf BUF1 (N9346, N9344);
and AND2 (N9347, N9345, N6663);
buf BUF1 (N9348, N9347);
xor XOR2 (N9349, N9330, N2881);
nor NOR4 (N9350, N9338, N7684, N8809, N7720);
nand NAND3 (N9351, N9348, N5322, N1208);
xor XOR2 (N9352, N9350, N2152);
nand NAND3 (N9353, N9335, N8920, N8882);
not NOT1 (N9354, N9340);
or OR3 (N9355, N9319, N2380, N9341);
buf BUF1 (N9356, N9337);
buf BUF1 (N9357, N9354);
not NOT1 (N9358, N9346);
xor XOR2 (N9359, N9339, N1672);
buf BUF1 (N9360, N9357);
nor NOR2 (N9361, N9360, N5734);
nor NOR2 (N9362, N9351, N3598);
buf BUF1 (N9363, N9356);
and AND4 (N9364, N9362, N3559, N5637, N4810);
or OR3 (N9365, N9349, N5905, N8068);
buf BUF1 (N9366, N9363);
or OR2 (N9367, N9361, N851);
buf BUF1 (N9368, N9358);
or OR2 (N9369, N9364, N4321);
buf BUF1 (N9370, N9366);
not NOT1 (N9371, N9367);
buf BUF1 (N9372, N9365);
not NOT1 (N9373, N9372);
nand NAND3 (N9374, N9369, N3174, N7728);
or OR4 (N9375, N9352, N8903, N7894, N4305);
nand NAND4 (N9376, N9374, N199, N3907, N6858);
buf BUF1 (N9377, N9333);
not NOT1 (N9378, N9355);
buf BUF1 (N9379, N9377);
and AND3 (N9380, N9376, N7598, N8154);
nand NAND3 (N9381, N9379, N299, N5732);
xor XOR2 (N9382, N9353, N6281);
not NOT1 (N9383, N9381);
or OR3 (N9384, N9368, N6997, N2670);
nor NOR4 (N9385, N9382, N2480, N8236, N4487);
buf BUF1 (N9386, N9370);
or OR4 (N9387, N9385, N795, N5291, N5283);
nand NAND2 (N9388, N9373, N4632);
or OR3 (N9389, N9383, N3438, N3181);
nand NAND4 (N9390, N9386, N4007, N8988, N3059);
or OR3 (N9391, N9387, N4495, N9200);
nor NOR2 (N9392, N9388, N767);
xor XOR2 (N9393, N9380, N6731);
buf BUF1 (N9394, N9391);
not NOT1 (N9395, N9375);
not NOT1 (N9396, N9393);
and AND2 (N9397, N9390, N8187);
nand NAND3 (N9398, N9394, N7666, N9005);
nand NAND3 (N9399, N9389, N4736, N3725);
not NOT1 (N9400, N9359);
not NOT1 (N9401, N9399);
not NOT1 (N9402, N9371);
or OR4 (N9403, N9392, N5719, N5164, N3505);
not NOT1 (N9404, N9395);
not NOT1 (N9405, N9384);
or OR4 (N9406, N9400, N584, N2400, N5796);
buf BUF1 (N9407, N9402);
buf BUF1 (N9408, N9398);
nor NOR2 (N9409, N9406, N4427);
xor XOR2 (N9410, N9403, N6801);
xor XOR2 (N9411, N9409, N1848);
xor XOR2 (N9412, N9404, N9335);
xor XOR2 (N9413, N9411, N628);
buf BUF1 (N9414, N9408);
nand NAND2 (N9415, N9412, N7497);
and AND4 (N9416, N9415, N7289, N2988, N5315);
buf BUF1 (N9417, N9413);
nand NAND4 (N9418, N9396, N7879, N7640, N7467);
or OR4 (N9419, N9401, N1694, N9228, N8239);
nor NOR3 (N9420, N9414, N4155, N2051);
buf BUF1 (N9421, N9410);
xor XOR2 (N9422, N9418, N4182);
nor NOR3 (N9423, N9422, N4596, N7723);
not NOT1 (N9424, N9420);
buf BUF1 (N9425, N9424);
or OR3 (N9426, N9416, N6894, N3814);
xor XOR2 (N9427, N9419, N7234);
and AND4 (N9428, N9407, N8825, N7687, N2508);
nor NOR4 (N9429, N9417, N6876, N7586, N50);
or OR4 (N9430, N9378, N4255, N3784, N8159);
not NOT1 (N9431, N9428);
and AND3 (N9432, N9405, N6672, N5775);
buf BUF1 (N9433, N9425);
nor NOR4 (N9434, N9431, N5089, N2596, N1464);
nor NOR3 (N9435, N9429, N3744, N5585);
nor NOR4 (N9436, N9397, N4313, N2929, N8577);
not NOT1 (N9437, N9427);
and AND4 (N9438, N9433, N5611, N8132, N6361);
xor XOR2 (N9439, N9438, N8989);
nand NAND2 (N9440, N9437, N9434);
or OR2 (N9441, N5613, N7554);
nor NOR3 (N9442, N9440, N4465, N1149);
nand NAND4 (N9443, N9442, N6030, N1958, N5751);
not NOT1 (N9444, N9432);
xor XOR2 (N9445, N9436, N9041);
buf BUF1 (N9446, N9426);
or OR3 (N9447, N9444, N7692, N90);
buf BUF1 (N9448, N9439);
nand NAND3 (N9449, N9448, N9398, N6569);
and AND2 (N9450, N9430, N7856);
and AND3 (N9451, N9450, N8733, N5202);
and AND2 (N9452, N9435, N6881);
and AND4 (N9453, N9451, N2057, N4707, N4155);
or OR4 (N9454, N9447, N3287, N5384, N4358);
buf BUF1 (N9455, N9443);
and AND4 (N9456, N9453, N4246, N8290, N1444);
xor XOR2 (N9457, N9421, N3349);
not NOT1 (N9458, N9452);
buf BUF1 (N9459, N9457);
xor XOR2 (N9460, N9423, N3410);
xor XOR2 (N9461, N9455, N7646);
nor NOR3 (N9462, N9454, N4522, N6152);
or OR3 (N9463, N9441, N205, N5044);
xor XOR2 (N9464, N9446, N1084);
not NOT1 (N9465, N9463);
not NOT1 (N9466, N9461);
buf BUF1 (N9467, N9445);
not NOT1 (N9468, N9449);
buf BUF1 (N9469, N9467);
buf BUF1 (N9470, N9459);
not NOT1 (N9471, N9458);
buf BUF1 (N9472, N9468);
xor XOR2 (N9473, N9469, N1762);
nand NAND3 (N9474, N9473, N906, N6901);
buf BUF1 (N9475, N9474);
nor NOR4 (N9476, N9465, N1078, N8331, N6445);
nand NAND3 (N9477, N9460, N6892, N2168);
or OR4 (N9478, N9470, N7111, N6618, N2193);
xor XOR2 (N9479, N9472, N9329);
nand NAND3 (N9480, N9478, N9236, N2004);
nand NAND4 (N9481, N9456, N8056, N403, N5080);
and AND4 (N9482, N9479, N4166, N4451, N6240);
nor NOR3 (N9483, N9475, N3403, N4923);
not NOT1 (N9484, N9477);
nand NAND2 (N9485, N9482, N743);
nand NAND3 (N9486, N9476, N3937, N2911);
or OR3 (N9487, N9485, N2379, N7246);
buf BUF1 (N9488, N9480);
or OR2 (N9489, N9488, N3493);
or OR4 (N9490, N9464, N3782, N3332, N7803);
xor XOR2 (N9491, N9486, N5632);
xor XOR2 (N9492, N9481, N2454);
and AND3 (N9493, N9483, N718, N4761);
nand NAND2 (N9494, N9493, N958);
nor NOR3 (N9495, N9492, N543, N1824);
nand NAND3 (N9496, N9494, N1700, N9076);
and AND4 (N9497, N9466, N8586, N748, N6813);
or OR3 (N9498, N9487, N5199, N1805);
or OR4 (N9499, N9471, N2638, N3078, N1305);
nand NAND2 (N9500, N9490, N4738);
not NOT1 (N9501, N9500);
not NOT1 (N9502, N9462);
nand NAND2 (N9503, N9497, N5209);
nor NOR3 (N9504, N9498, N6170, N6211);
and AND2 (N9505, N9503, N5099);
nor NOR2 (N9506, N9499, N2370);
or OR2 (N9507, N9502, N6304);
or OR2 (N9508, N9507, N3442);
buf BUF1 (N9509, N9505);
buf BUF1 (N9510, N9504);
or OR4 (N9511, N9501, N5768, N8171, N4393);
nand NAND2 (N9512, N9496, N9151);
nand NAND4 (N9513, N9511, N1171, N5753, N5255);
nor NOR4 (N9514, N9506, N6964, N3922, N3039);
buf BUF1 (N9515, N9510);
and AND4 (N9516, N9489, N4743, N7399, N3772);
or OR2 (N9517, N9508, N906);
or OR3 (N9518, N9495, N6826, N5553);
nor NOR2 (N9519, N9484, N8292);
not NOT1 (N9520, N9516);
or OR2 (N9521, N9519, N9453);
and AND4 (N9522, N9520, N1941, N8672, N4082);
and AND2 (N9523, N9522, N5976);
not NOT1 (N9524, N9491);
xor XOR2 (N9525, N9509, N3193);
nor NOR4 (N9526, N9515, N1680, N2450, N3569);
buf BUF1 (N9527, N9521);
and AND3 (N9528, N9527, N7916, N328);
nor NOR4 (N9529, N9528, N7359, N8905, N1400);
or OR2 (N9530, N9529, N6258);
buf BUF1 (N9531, N9512);
xor XOR2 (N9532, N9514, N5361);
nor NOR3 (N9533, N9532, N9258, N5804);
nor NOR4 (N9534, N9517, N978, N7404, N3998);
nand NAND4 (N9535, N9518, N1489, N5458, N5800);
nand NAND2 (N9536, N9531, N4385);
nor NOR3 (N9537, N9523, N7666, N6608);
and AND3 (N9538, N9526, N6429, N8777);
or OR3 (N9539, N9535, N8043, N4331);
buf BUF1 (N9540, N9539);
buf BUF1 (N9541, N9530);
xor XOR2 (N9542, N9524, N6942);
nand NAND3 (N9543, N9538, N6923, N5055);
nand NAND4 (N9544, N9537, N4495, N2985, N5071);
nand NAND2 (N9545, N9536, N837);
and AND2 (N9546, N9542, N7575);
nor NOR2 (N9547, N9525, N603);
or OR4 (N9548, N9546, N1931, N1628, N1874);
or OR2 (N9549, N9533, N3246);
buf BUF1 (N9550, N9541);
not NOT1 (N9551, N9544);
and AND2 (N9552, N9543, N5761);
buf BUF1 (N9553, N9547);
nand NAND4 (N9554, N9513, N1246, N4482, N8002);
or OR2 (N9555, N9550, N3034);
or OR4 (N9556, N9552, N8052, N61, N1156);
not NOT1 (N9557, N9545);
not NOT1 (N9558, N9540);
not NOT1 (N9559, N9534);
buf BUF1 (N9560, N9555);
nor NOR2 (N9561, N9559, N6235);
not NOT1 (N9562, N9551);
not NOT1 (N9563, N9549);
xor XOR2 (N9564, N9553, N6837);
and AND3 (N9565, N9557, N1564, N8879);
buf BUF1 (N9566, N9556);
buf BUF1 (N9567, N9560);
and AND3 (N9568, N9565, N485, N2015);
nor NOR4 (N9569, N9566, N4092, N4047, N4147);
xor XOR2 (N9570, N9562, N9102);
and AND3 (N9571, N9558, N4675, N1467);
or OR3 (N9572, N9564, N5155, N1536);
or OR4 (N9573, N9561, N9166, N2813, N3035);
and AND3 (N9574, N9568, N9207, N6024);
xor XOR2 (N9575, N9574, N9438);
nor NOR4 (N9576, N9571, N9252, N5299, N2608);
not NOT1 (N9577, N9575);
not NOT1 (N9578, N9576);
xor XOR2 (N9579, N9567, N3888);
xor XOR2 (N9580, N9563, N7871);
or OR3 (N9581, N9572, N8067, N1581);
nand NAND2 (N9582, N9569, N5938);
buf BUF1 (N9583, N9573);
buf BUF1 (N9584, N9582);
buf BUF1 (N9585, N9581);
nor NOR2 (N9586, N9577, N6101);
nand NAND2 (N9587, N9585, N7837);
and AND3 (N9588, N9586, N1112, N9328);
or OR4 (N9589, N9583, N5422, N8499, N3408);
and AND3 (N9590, N9588, N4808, N269);
nand NAND2 (N9591, N9579, N8815);
xor XOR2 (N9592, N9580, N5);
nor NOR4 (N9593, N9590, N304, N8435, N9337);
nor NOR3 (N9594, N9578, N9516, N4975);
and AND4 (N9595, N9593, N1085, N5298, N1401);
nor NOR2 (N9596, N9594, N453);
buf BUF1 (N9597, N9592);
not NOT1 (N9598, N9570);
nor NOR3 (N9599, N9591, N24, N9032);
buf BUF1 (N9600, N9595);
buf BUF1 (N9601, N9587);
nor NOR3 (N9602, N9598, N969, N633);
nor NOR4 (N9603, N9584, N6093, N3890, N2703);
or OR3 (N9604, N9548, N7425, N2213);
and AND4 (N9605, N9589, N6867, N8500, N6119);
and AND3 (N9606, N9602, N3596, N5121);
buf BUF1 (N9607, N9601);
xor XOR2 (N9608, N9606, N3214);
and AND2 (N9609, N9604, N4034);
nand NAND2 (N9610, N9603, N6025);
or OR2 (N9611, N9600, N6134);
xor XOR2 (N9612, N9597, N4545);
buf BUF1 (N9613, N9612);
or OR4 (N9614, N9554, N5441, N4285, N4602);
or OR4 (N9615, N9614, N7819, N5939, N3737);
and AND2 (N9616, N9605, N3);
xor XOR2 (N9617, N9607, N550);
nor NOR3 (N9618, N9608, N8400, N6249);
nor NOR4 (N9619, N9616, N4247, N4426, N5371);
xor XOR2 (N9620, N9611, N6881);
xor XOR2 (N9621, N9617, N796);
xor XOR2 (N9622, N9596, N6844);
or OR2 (N9623, N9610, N3056);
buf BUF1 (N9624, N9615);
xor XOR2 (N9625, N9619, N9455);
xor XOR2 (N9626, N9621, N3770);
or OR4 (N9627, N9623, N3407, N7522, N7346);
and AND3 (N9628, N9620, N9006, N6929);
or OR4 (N9629, N9627, N635, N6341, N7146);
buf BUF1 (N9630, N9622);
buf BUF1 (N9631, N9609);
nand NAND3 (N9632, N9625, N3102, N2772);
not NOT1 (N9633, N9629);
and AND4 (N9634, N9630, N2403, N2469, N297);
nand NAND4 (N9635, N9632, N1011, N111, N2356);
xor XOR2 (N9636, N9599, N4616);
nor NOR4 (N9637, N9631, N5337, N5886, N1583);
nor NOR3 (N9638, N9637, N2002, N3626);
xor XOR2 (N9639, N9628, N1912);
nand NAND2 (N9640, N9633, N8591);
xor XOR2 (N9641, N9624, N3737);
nand NAND2 (N9642, N9636, N4265);
buf BUF1 (N9643, N9638);
xor XOR2 (N9644, N9640, N1717);
not NOT1 (N9645, N9639);
nand NAND4 (N9646, N9618, N1309, N1834, N4838);
nor NOR2 (N9647, N9642, N410);
and AND3 (N9648, N9613, N528, N9515);
and AND3 (N9649, N9646, N3527, N5044);
buf BUF1 (N9650, N9643);
xor XOR2 (N9651, N9650, N7931);
buf BUF1 (N9652, N9645);
not NOT1 (N9653, N9626);
nor NOR3 (N9654, N9648, N7645, N7681);
not NOT1 (N9655, N9654);
not NOT1 (N9656, N9651);
buf BUF1 (N9657, N9655);
or OR2 (N9658, N9641, N25);
not NOT1 (N9659, N9658);
nand NAND3 (N9660, N9647, N8030, N6226);
xor XOR2 (N9661, N9657, N8884);
nand NAND4 (N9662, N9652, N9486, N3174, N2127);
or OR3 (N9663, N9660, N5608, N4455);
or OR2 (N9664, N9644, N9038);
nand NAND3 (N9665, N9659, N7250, N7343);
and AND3 (N9666, N9649, N5813, N3158);
and AND4 (N9667, N9666, N1085, N2708, N710);
buf BUF1 (N9668, N9634);
xor XOR2 (N9669, N9664, N573);
nand NAND3 (N9670, N9656, N5204, N7643);
or OR4 (N9671, N9665, N8638, N450, N674);
and AND2 (N9672, N9670, N5764);
nand NAND2 (N9673, N9671, N4541);
and AND2 (N9674, N9673, N607);
buf BUF1 (N9675, N9635);
buf BUF1 (N9676, N9667);
not NOT1 (N9677, N9675);
and AND3 (N9678, N9676, N3292, N1762);
xor XOR2 (N9679, N9669, N3566);
or OR3 (N9680, N9679, N1157, N5821);
not NOT1 (N9681, N9677);
nor NOR4 (N9682, N9680, N6597, N6117, N9234);
buf BUF1 (N9683, N9668);
nor NOR2 (N9684, N9681, N214);
xor XOR2 (N9685, N9682, N616);
or OR3 (N9686, N9662, N6026, N2751);
nand NAND4 (N9687, N9663, N3385, N3666, N4271);
or OR4 (N9688, N9653, N9166, N6260, N9666);
buf BUF1 (N9689, N9674);
buf BUF1 (N9690, N9684);
and AND2 (N9691, N9687, N2804);
and AND4 (N9692, N9672, N9240, N7682, N2004);
nor NOR3 (N9693, N9686, N8408, N8833);
or OR2 (N9694, N9691, N407);
buf BUF1 (N9695, N9694);
nor NOR4 (N9696, N9690, N5432, N1569, N3042);
nor NOR3 (N9697, N9689, N3846, N112);
nand NAND4 (N9698, N9661, N1508, N5267, N3752);
and AND3 (N9699, N9685, N6668, N9453);
buf BUF1 (N9700, N9699);
or OR2 (N9701, N9698, N9043);
xor XOR2 (N9702, N9700, N3427);
xor XOR2 (N9703, N9683, N7137);
or OR2 (N9704, N9692, N8487);
nor NOR3 (N9705, N9696, N6548, N4055);
and AND3 (N9706, N9693, N3582, N578);
and AND2 (N9707, N9702, N4901);
or OR2 (N9708, N9704, N246);
and AND3 (N9709, N9708, N5345, N238);
nand NAND3 (N9710, N9705, N1392, N7375);
and AND2 (N9711, N9710, N4938);
xor XOR2 (N9712, N9688, N8114);
nand NAND2 (N9713, N9711, N6538);
buf BUF1 (N9714, N9713);
not NOT1 (N9715, N9706);
buf BUF1 (N9716, N9715);
not NOT1 (N9717, N9709);
buf BUF1 (N9718, N9695);
not NOT1 (N9719, N9717);
buf BUF1 (N9720, N9697);
or OR2 (N9721, N9720, N3885);
xor XOR2 (N9722, N9718, N8257);
not NOT1 (N9723, N9678);
or OR3 (N9724, N9716, N3850, N3585);
and AND3 (N9725, N9719, N6007, N4875);
and AND3 (N9726, N9723, N3062, N8502);
buf BUF1 (N9727, N9722);
not NOT1 (N9728, N9707);
nor NOR3 (N9729, N9703, N1780, N8180);
or OR2 (N9730, N9724, N6726);
nor NOR4 (N9731, N9726, N8860, N7599, N318);
nor NOR2 (N9732, N9701, N5233);
buf BUF1 (N9733, N9714);
and AND4 (N9734, N9732, N8087, N714, N3360);
buf BUF1 (N9735, N9721);
nor NOR2 (N9736, N9727, N6548);
not NOT1 (N9737, N9734);
and AND3 (N9738, N9736, N5847, N1970);
nor NOR4 (N9739, N9729, N1849, N1786, N2025);
xor XOR2 (N9740, N9733, N8028);
nand NAND2 (N9741, N9737, N7373);
xor XOR2 (N9742, N9735, N6296);
nor NOR4 (N9743, N9712, N7027, N725, N6508);
xor XOR2 (N9744, N9738, N3674);
or OR2 (N9745, N9725, N3155);
nor NOR3 (N9746, N9744, N8586, N3189);
nand NAND2 (N9747, N9743, N7552);
xor XOR2 (N9748, N9747, N94);
nor NOR3 (N9749, N9740, N8227, N2470);
and AND3 (N9750, N9730, N2381, N2408);
buf BUF1 (N9751, N9745);
xor XOR2 (N9752, N9751, N8678);
or OR4 (N9753, N9748, N3696, N689, N4484);
and AND3 (N9754, N9741, N9580, N257);
nand NAND3 (N9755, N9753, N6477, N6443);
buf BUF1 (N9756, N9752);
or OR2 (N9757, N9731, N9604);
nand NAND2 (N9758, N9742, N3067);
nand NAND3 (N9759, N9749, N7031, N3866);
buf BUF1 (N9760, N9759);
buf BUF1 (N9761, N9750);
buf BUF1 (N9762, N9757);
nor NOR2 (N9763, N9758, N1828);
xor XOR2 (N9764, N9761, N2710);
not NOT1 (N9765, N9754);
nand NAND3 (N9766, N9755, N5642, N9624);
xor XOR2 (N9767, N9762, N2339);
or OR2 (N9768, N9746, N2277);
or OR3 (N9769, N9765, N1179, N58);
nand NAND2 (N9770, N9728, N9574);
or OR2 (N9771, N9769, N563);
nand NAND4 (N9772, N9764, N5494, N1577, N2838);
not NOT1 (N9773, N9763);
nor NOR3 (N9774, N9756, N1541, N3333);
nor NOR4 (N9775, N9772, N8404, N1566, N8690);
not NOT1 (N9776, N9775);
nor NOR4 (N9777, N9771, N6835, N4585, N7013);
or OR3 (N9778, N9774, N9439, N8183);
not NOT1 (N9779, N9773);
not NOT1 (N9780, N9776);
and AND4 (N9781, N9766, N7254, N5067, N9612);
and AND3 (N9782, N9760, N8362, N5407);
nand NAND2 (N9783, N9768, N7878);
or OR4 (N9784, N9781, N2714, N5015, N3336);
and AND3 (N9785, N9779, N9387, N8389);
not NOT1 (N9786, N9778);
buf BUF1 (N9787, N9739);
nand NAND2 (N9788, N9782, N6925);
and AND2 (N9789, N9770, N1655);
and AND3 (N9790, N9788, N2809, N689);
xor XOR2 (N9791, N9786, N8773);
and AND3 (N9792, N9780, N7128, N4900);
buf BUF1 (N9793, N9791);
buf BUF1 (N9794, N9785);
not NOT1 (N9795, N9794);
buf BUF1 (N9796, N9784);
or OR3 (N9797, N9795, N1477, N6150);
xor XOR2 (N9798, N9797, N4894);
nor NOR4 (N9799, N9798, N6216, N790, N9524);
and AND4 (N9800, N9767, N6643, N7209, N9246);
not NOT1 (N9801, N9787);
nor NOR2 (N9802, N9793, N8812);
nor NOR2 (N9803, N9792, N51);
or OR2 (N9804, N9796, N7707);
buf BUF1 (N9805, N9777);
or OR4 (N9806, N9805, N7301, N9318, N891);
or OR2 (N9807, N9790, N7687);
xor XOR2 (N9808, N9802, N5749);
xor XOR2 (N9809, N9789, N3055);
and AND3 (N9810, N9807, N8993, N6084);
not NOT1 (N9811, N9806);
nand NAND3 (N9812, N9809, N4313, N6674);
nand NAND4 (N9813, N9812, N4003, N3985, N2649);
buf BUF1 (N9814, N9803);
nand NAND2 (N9815, N9811, N3278);
xor XOR2 (N9816, N9813, N3190);
nor NOR4 (N9817, N9783, N8269, N7494, N7089);
buf BUF1 (N9818, N9816);
xor XOR2 (N9819, N9804, N3229);
or OR3 (N9820, N9799, N7012, N7250);
nor NOR3 (N9821, N9820, N1795, N9219);
or OR2 (N9822, N9815, N4659);
not NOT1 (N9823, N9801);
nand NAND2 (N9824, N9822, N1061);
xor XOR2 (N9825, N9821, N2035);
buf BUF1 (N9826, N9824);
or OR4 (N9827, N9800, N8547, N1125, N5575);
not NOT1 (N9828, N9819);
buf BUF1 (N9829, N9825);
and AND2 (N9830, N9808, N2488);
nor NOR4 (N9831, N9818, N7417, N5717, N4565);
or OR3 (N9832, N9830, N8039, N7766);
and AND3 (N9833, N9832, N1478, N6939);
buf BUF1 (N9834, N9829);
and AND4 (N9835, N9827, N215, N3704, N3250);
not NOT1 (N9836, N9826);
not NOT1 (N9837, N9834);
xor XOR2 (N9838, N9837, N8420);
nand NAND2 (N9839, N9831, N7459);
buf BUF1 (N9840, N9823);
and AND3 (N9841, N9814, N743, N831);
nand NAND4 (N9842, N9839, N844, N4326, N5464);
and AND2 (N9843, N9833, N4184);
or OR3 (N9844, N9840, N4377, N5983);
or OR2 (N9845, N9842, N5678);
and AND3 (N9846, N9817, N1959, N3242);
not NOT1 (N9847, N9810);
or OR4 (N9848, N9846, N41, N2811, N1655);
not NOT1 (N9849, N9844);
and AND3 (N9850, N9845, N4020, N9617);
nor NOR2 (N9851, N9841, N1035);
not NOT1 (N9852, N9843);
nor NOR3 (N9853, N9838, N8519, N6172);
xor XOR2 (N9854, N9835, N6390);
buf BUF1 (N9855, N9854);
nor NOR4 (N9856, N9850, N2733, N5094, N2129);
or OR4 (N9857, N9851, N7318, N429, N8409);
not NOT1 (N9858, N9849);
buf BUF1 (N9859, N9855);
nand NAND4 (N9860, N9848, N5151, N8104, N6851);
nand NAND3 (N9861, N9852, N8856, N6722);
not NOT1 (N9862, N9857);
and AND3 (N9863, N9828, N927, N2179);
and AND2 (N9864, N9836, N4875);
or OR4 (N9865, N9856, N538, N9677, N639);
and AND3 (N9866, N9861, N4720, N8732);
xor XOR2 (N9867, N9865, N3660);
nand NAND3 (N9868, N9863, N4342, N1633);
nor NOR4 (N9869, N9858, N8317, N4936, N5944);
xor XOR2 (N9870, N9860, N5699);
nor NOR3 (N9871, N9868, N4959, N3571);
nor NOR3 (N9872, N9862, N2698, N5936);
nand NAND4 (N9873, N9847, N2510, N6016, N8254);
nor NOR2 (N9874, N9871, N1789);
buf BUF1 (N9875, N9872);
or OR3 (N9876, N9869, N8185, N2626);
and AND3 (N9877, N9874, N2454, N9329);
xor XOR2 (N9878, N9877, N3820);
or OR2 (N9879, N9859, N6374);
not NOT1 (N9880, N9879);
xor XOR2 (N9881, N9873, N6821);
buf BUF1 (N9882, N9881);
nand NAND3 (N9883, N9878, N2624, N217);
nand NAND2 (N9884, N9875, N1511);
or OR3 (N9885, N9866, N1995, N176);
not NOT1 (N9886, N9884);
and AND2 (N9887, N9880, N7488);
nand NAND2 (N9888, N9867, N652);
not NOT1 (N9889, N9853);
buf BUF1 (N9890, N9882);
nand NAND3 (N9891, N9886, N9133, N3390);
or OR3 (N9892, N9876, N5955, N3368);
nor NOR2 (N9893, N9870, N6823);
xor XOR2 (N9894, N9890, N4043);
not NOT1 (N9895, N9888);
buf BUF1 (N9896, N9893);
xor XOR2 (N9897, N9896, N4201);
xor XOR2 (N9898, N9892, N4452);
nor NOR3 (N9899, N9885, N2373, N6348);
nand NAND3 (N9900, N9891, N75, N1677);
not NOT1 (N9901, N9894);
nor NOR4 (N9902, N9895, N2162, N8748, N6233);
xor XOR2 (N9903, N9900, N470);
xor XOR2 (N9904, N9889, N3094);
not NOT1 (N9905, N9903);
nor NOR2 (N9906, N9898, N2995);
buf BUF1 (N9907, N9901);
or OR2 (N9908, N9883, N5936);
or OR3 (N9909, N9887, N5386, N4945);
and AND3 (N9910, N9897, N5078, N953);
or OR3 (N9911, N9909, N9619, N8608);
buf BUF1 (N9912, N9911);
nor NOR2 (N9913, N9910, N1374);
buf BUF1 (N9914, N9864);
and AND4 (N9915, N9907, N264, N1305, N6597);
or OR4 (N9916, N9913, N1129, N7106, N3954);
or OR2 (N9917, N9899, N6010);
or OR4 (N9918, N9904, N9534, N7635, N2360);
and AND3 (N9919, N9917, N123, N7905);
and AND3 (N9920, N9919, N6366, N1796);
nand NAND3 (N9921, N9916, N1746, N3627);
nand NAND3 (N9922, N9905, N9803, N7337);
xor XOR2 (N9923, N9912, N5840);
not NOT1 (N9924, N9914);
or OR3 (N9925, N9906, N8889, N9767);
nor NOR4 (N9926, N9915, N4695, N8478, N472);
nand NAND2 (N9927, N9918, N3534);
nand NAND2 (N9928, N9926, N5584);
and AND3 (N9929, N9921, N6382, N6761);
or OR3 (N9930, N9902, N6428, N4874);
nor NOR4 (N9931, N9920, N2445, N9746, N4556);
nand NAND4 (N9932, N9931, N3579, N3863, N1817);
not NOT1 (N9933, N9928);
or OR2 (N9934, N9929, N7471);
buf BUF1 (N9935, N9924);
nor NOR2 (N9936, N9922, N563);
or OR3 (N9937, N9930, N9454, N7562);
buf BUF1 (N9938, N9933);
or OR4 (N9939, N9927, N3448, N729, N9323);
xor XOR2 (N9940, N9934, N4572);
not NOT1 (N9941, N9908);
buf BUF1 (N9942, N9940);
nor NOR3 (N9943, N9923, N5173, N3799);
or OR4 (N9944, N9935, N4672, N698, N84);
buf BUF1 (N9945, N9932);
buf BUF1 (N9946, N9937);
nand NAND3 (N9947, N9945, N5609, N2957);
nor NOR4 (N9948, N9936, N7032, N6918, N5986);
not NOT1 (N9949, N9944);
not NOT1 (N9950, N9942);
nand NAND2 (N9951, N9948, N3778);
not NOT1 (N9952, N9925);
or OR4 (N9953, N9947, N8000, N3678, N5505);
nor NOR4 (N9954, N9946, N2062, N1273, N3835);
or OR2 (N9955, N9938, N9041);
nor NOR3 (N9956, N9950, N9182, N7530);
nor NOR2 (N9957, N9951, N6479);
xor XOR2 (N9958, N9956, N1829);
and AND4 (N9959, N9954, N2382, N1061, N4641);
nand NAND3 (N9960, N9955, N4288, N5486);
and AND3 (N9961, N9949, N4215, N4381);
not NOT1 (N9962, N9958);
buf BUF1 (N9963, N9961);
not NOT1 (N9964, N9953);
and AND4 (N9965, N9959, N2745, N7064, N962);
nor NOR2 (N9966, N9957, N8969);
xor XOR2 (N9967, N9939, N8241);
not NOT1 (N9968, N9941);
xor XOR2 (N9969, N9960, N758);
xor XOR2 (N9970, N9964, N5983);
nor NOR4 (N9971, N9952, N6133, N398, N7396);
and AND4 (N9972, N9969, N8602, N7301, N1438);
nor NOR3 (N9973, N9968, N6019, N8688);
nor NOR4 (N9974, N9943, N3274, N5911, N6951);
buf BUF1 (N9975, N9966);
not NOT1 (N9976, N9971);
xor XOR2 (N9977, N9975, N7907);
and AND3 (N9978, N9963, N4819, N1715);
and AND3 (N9979, N9978, N3205, N141);
or OR3 (N9980, N9965, N5390, N9742);
buf BUF1 (N9981, N9962);
or OR3 (N9982, N9973, N7353, N475);
and AND4 (N9983, N9974, N5248, N4895, N6524);
nor NOR3 (N9984, N9979, N9494, N3326);
and AND2 (N9985, N9983, N644);
buf BUF1 (N9986, N9977);
nand NAND2 (N9987, N9984, N9053);
nor NOR4 (N9988, N9986, N1003, N8861, N3966);
and AND3 (N9989, N9987, N5665, N4845);
not NOT1 (N9990, N9982);
and AND2 (N9991, N9972, N1457);
and AND4 (N9992, N9985, N316, N773, N7921);
nor NOR4 (N9993, N9989, N4984, N5908, N3208);
not NOT1 (N9994, N9980);
nand NAND4 (N9995, N9993, N5592, N6272, N5036);
nand NAND4 (N9996, N9992, N2887, N3364, N9550);
nor NOR2 (N9997, N9976, N8032);
nand NAND4 (N9998, N9967, N7188, N805, N9221);
not NOT1 (N9999, N9996);
and AND4 (N10000, N9997, N6314, N2937, N2199);
nand NAND3 (N10001, N9970, N7793, N9952);
nor NOR4 (N10002, N10001, N6748, N7659, N4605);
and AND4 (N10003, N9998, N452, N6957, N7912);
or OR4 (N10004, N9990, N1191, N431, N6785);
not NOT1 (N10005, N9991);
nor NOR4 (N10006, N10005, N5810, N6587, N813);
not NOT1 (N10007, N10000);
nand NAND3 (N10008, N10003, N8702, N3455);
not NOT1 (N10009, N9999);
xor XOR2 (N10010, N10008, N1998);
xor XOR2 (N10011, N9981, N5205);
not NOT1 (N10012, N10002);
nor NOR3 (N10013, N9988, N5532, N3032);
and AND2 (N10014, N10006, N5830);
buf BUF1 (N10015, N10014);
nor NOR3 (N10016, N10012, N1011, N8864);
and AND2 (N10017, N10016, N9054);
nor NOR3 (N10018, N10007, N7807, N16);
nand NAND3 (N10019, N10017, N5633, N1246);
xor XOR2 (N10020, N10009, N6449);
and AND2 (N10021, N10004, N1694);
nor NOR2 (N10022, N10013, N2176);
or OR3 (N10023, N10018, N2394, N2793);
nand NAND3 (N10024, N10022, N8169, N4260);
nand NAND4 (N10025, N10015, N5300, N2643, N5626);
and AND3 (N10026, N10011, N9018, N7769);
buf BUF1 (N10027, N9995);
or OR4 (N10028, N10020, N7024, N4141, N2819);
or OR3 (N10029, N10023, N241, N1096);
xor XOR2 (N10030, N10026, N5638);
buf BUF1 (N10031, N10010);
not NOT1 (N10032, N10028);
buf BUF1 (N10033, N10029);
and AND3 (N10034, N10032, N3254, N4432);
buf BUF1 (N10035, N10019);
nand NAND4 (N10036, N10033, N529, N1431, N632);
or OR4 (N10037, N10025, N7161, N814, N139);
not NOT1 (N10038, N10030);
nor NOR2 (N10039, N10036, N9766);
xor XOR2 (N10040, N10034, N1177);
not NOT1 (N10041, N10024);
and AND4 (N10042, N10031, N5366, N7756, N1384);
not NOT1 (N10043, N10038);
xor XOR2 (N10044, N10042, N1664);
xor XOR2 (N10045, N10044, N302);
nand NAND2 (N10046, N10043, N8354);
and AND3 (N10047, N10045, N309, N3932);
nor NOR4 (N10048, N10039, N7348, N7025, N4028);
not NOT1 (N10049, N10048);
not NOT1 (N10050, N9994);
nor NOR4 (N10051, N10027, N221, N2711, N4562);
nor NOR2 (N10052, N10021, N3719);
nand NAND2 (N10053, N10037, N5167);
not NOT1 (N10054, N10051);
nor NOR2 (N10055, N10052, N129);
or OR3 (N10056, N10041, N4372, N1388);
and AND4 (N10057, N10040, N9520, N9077, N6632);
nand NAND2 (N10058, N10057, N580);
nor NOR2 (N10059, N10053, N3777);
xor XOR2 (N10060, N10054, N6002);
nand NAND4 (N10061, N10046, N369, N6294, N1347);
not NOT1 (N10062, N10035);
not NOT1 (N10063, N10050);
xor XOR2 (N10064, N10063, N2319);
not NOT1 (N10065, N10064);
nand NAND2 (N10066, N10060, N1443);
nand NAND3 (N10067, N10056, N2750, N3376);
not NOT1 (N10068, N10058);
or OR2 (N10069, N10068, N626);
and AND4 (N10070, N10067, N5843, N5988, N7830);
nor NOR4 (N10071, N10066, N2977, N2481, N236);
nand NAND3 (N10072, N10049, N150, N6945);
buf BUF1 (N10073, N10070);
not NOT1 (N10074, N10061);
buf BUF1 (N10075, N10047);
or OR4 (N10076, N10062, N2562, N7999, N3048);
nand NAND4 (N10077, N10055, N10061, N9082, N3073);
nor NOR3 (N10078, N10069, N5668, N6548);
xor XOR2 (N10079, N10078, N1720);
or OR2 (N10080, N10071, N825);
buf BUF1 (N10081, N10075);
not NOT1 (N10082, N10081);
nand NAND4 (N10083, N10082, N3701, N2177, N5575);
not NOT1 (N10084, N10059);
or OR4 (N10085, N10083, N4457, N7550, N5750);
nor NOR2 (N10086, N10076, N6225);
nor NOR2 (N10087, N10072, N4884);
nand NAND4 (N10088, N10079, N9403, N4318, N3501);
and AND3 (N10089, N10084, N4544, N2886);
and AND2 (N10090, N10088, N210);
xor XOR2 (N10091, N10074, N5165);
xor XOR2 (N10092, N10085, N7779);
nor NOR3 (N10093, N10080, N1477, N7223);
xor XOR2 (N10094, N10087, N9484);
and AND2 (N10095, N10093, N4135);
and AND4 (N10096, N10086, N915, N9075, N5586);
buf BUF1 (N10097, N10089);
or OR4 (N10098, N10096, N3337, N3652, N6506);
nor NOR3 (N10099, N10094, N4718, N7732);
or OR3 (N10100, N10098, N7422, N7549);
buf BUF1 (N10101, N10091);
not NOT1 (N10102, N10073);
and AND4 (N10103, N10090, N398, N6481, N2488);
nand NAND2 (N10104, N10077, N5771);
xor XOR2 (N10105, N10092, N8306);
or OR4 (N10106, N10100, N5818, N6641, N1327);
buf BUF1 (N10107, N10101);
nor NOR2 (N10108, N10065, N8382);
nand NAND3 (N10109, N10108, N2483, N6585);
xor XOR2 (N10110, N10104, N5040);
nand NAND2 (N10111, N10102, N1923);
buf BUF1 (N10112, N10109);
not NOT1 (N10113, N10099);
nor NOR4 (N10114, N10103, N8110, N4803, N5250);
or OR3 (N10115, N10097, N3963, N3979);
not NOT1 (N10116, N10112);
nand NAND3 (N10117, N10115, N7299, N1837);
and AND3 (N10118, N10105, N6673, N4759);
buf BUF1 (N10119, N10118);
and AND3 (N10120, N10111, N8719, N2556);
and AND4 (N10121, N10095, N5373, N1283, N1243);
buf BUF1 (N10122, N10107);
and AND3 (N10123, N10116, N8913, N9005);
not NOT1 (N10124, N10117);
and AND3 (N10125, N10113, N7503, N4922);
nor NOR4 (N10126, N10120, N5400, N3147, N7159);
nor NOR2 (N10127, N10123, N8825);
xor XOR2 (N10128, N10114, N8880);
or OR2 (N10129, N10106, N5324);
xor XOR2 (N10130, N10128, N1873);
nand NAND4 (N10131, N10126, N3466, N2353, N5169);
xor XOR2 (N10132, N10127, N4465);
or OR3 (N10133, N10110, N8957, N4855);
buf BUF1 (N10134, N10119);
nor NOR4 (N10135, N10133, N8172, N2682, N3234);
buf BUF1 (N10136, N10124);
nand NAND4 (N10137, N10136, N3444, N8853, N4479);
buf BUF1 (N10138, N10121);
xor XOR2 (N10139, N10122, N397);
not NOT1 (N10140, N10132);
and AND3 (N10141, N10135, N4692, N168);
buf BUF1 (N10142, N10141);
buf BUF1 (N10143, N10138);
nor NOR3 (N10144, N10143, N7414, N9481);
or OR4 (N10145, N10140, N346, N44, N4973);
or OR4 (N10146, N10142, N3693, N2497, N5476);
buf BUF1 (N10147, N10146);
and AND4 (N10148, N10147, N9115, N7404, N8486);
xor XOR2 (N10149, N10130, N6524);
and AND4 (N10150, N10129, N5790, N8670, N7062);
not NOT1 (N10151, N10137);
not NOT1 (N10152, N10131);
xor XOR2 (N10153, N10139, N3301);
and AND4 (N10154, N10151, N7818, N7773, N1378);
buf BUF1 (N10155, N10153);
or OR3 (N10156, N10154, N694, N6598);
nor NOR2 (N10157, N10148, N4185);
or OR3 (N10158, N10155, N8733, N1538);
and AND4 (N10159, N10158, N5847, N1770, N1935);
nor NOR4 (N10160, N10134, N141, N7626, N1028);
nor NOR4 (N10161, N10125, N3868, N1806, N1254);
and AND4 (N10162, N10145, N5877, N964, N3951);
and AND4 (N10163, N10152, N8498, N8764, N352);
not NOT1 (N10164, N10150);
buf BUF1 (N10165, N10162);
nand NAND3 (N10166, N10165, N8394, N2620);
and AND3 (N10167, N10149, N991, N8894);
nor NOR2 (N10168, N10144, N8601);
buf BUF1 (N10169, N10163);
not NOT1 (N10170, N10160);
nor NOR2 (N10171, N10168, N7223);
not NOT1 (N10172, N10161);
and AND4 (N10173, N10157, N8279, N2171, N7488);
nor NOR4 (N10174, N10156, N9401, N5292, N10104);
xor XOR2 (N10175, N10171, N2200);
nand NAND3 (N10176, N10166, N1475, N1732);
buf BUF1 (N10177, N10167);
nand NAND2 (N10178, N10169, N2158);
or OR3 (N10179, N10172, N5078, N2969);
or OR2 (N10180, N10176, N10068);
and AND4 (N10181, N10179, N2314, N8845, N129);
or OR2 (N10182, N10175, N10097);
nor NOR2 (N10183, N10173, N7219);
buf BUF1 (N10184, N10180);
nand NAND3 (N10185, N10184, N1893, N2316);
nor NOR3 (N10186, N10177, N3172, N5295);
buf BUF1 (N10187, N10178);
and AND4 (N10188, N10159, N3039, N4775, N8490);
nor NOR2 (N10189, N10174, N7943);
not NOT1 (N10190, N10188);
not NOT1 (N10191, N10190);
and AND2 (N10192, N10183, N2029);
not NOT1 (N10193, N10191);
and AND4 (N10194, N10164, N3236, N9630, N9198);
not NOT1 (N10195, N10192);
nor NOR3 (N10196, N10170, N7657, N2050);
or OR3 (N10197, N10182, N7108, N601);
and AND4 (N10198, N10186, N813, N2982, N523);
and AND3 (N10199, N10194, N3204, N6948);
nand NAND3 (N10200, N10197, N385, N1230);
or OR4 (N10201, N10193, N4295, N7271, N2476);
nand NAND2 (N10202, N10185, N1517);
and AND4 (N10203, N10201, N4609, N1615, N9938);
nor NOR2 (N10204, N10187, N7296);
xor XOR2 (N10205, N10181, N7569);
not NOT1 (N10206, N10203);
nor NOR3 (N10207, N10200, N1363, N1422);
xor XOR2 (N10208, N10204, N2560);
and AND3 (N10209, N10195, N9979, N7297);
buf BUF1 (N10210, N10199);
not NOT1 (N10211, N10205);
nand NAND2 (N10212, N10208, N7699);
xor XOR2 (N10213, N10207, N4952);
xor XOR2 (N10214, N10212, N186);
not NOT1 (N10215, N10196);
and AND2 (N10216, N10206, N8397);
or OR2 (N10217, N10209, N3499);
or OR3 (N10218, N10198, N1980, N6618);
xor XOR2 (N10219, N10214, N9768);
and AND4 (N10220, N10189, N2807, N2006, N839);
and AND3 (N10221, N10211, N3172, N8305);
not NOT1 (N10222, N10202);
not NOT1 (N10223, N10213);
xor XOR2 (N10224, N10216, N6876);
and AND3 (N10225, N10217, N8767, N183);
xor XOR2 (N10226, N10219, N1231);
nand NAND2 (N10227, N10224, N8299);
nor NOR2 (N10228, N10225, N641);
not NOT1 (N10229, N10215);
not NOT1 (N10230, N10223);
or OR3 (N10231, N10228, N3929, N6639);
and AND2 (N10232, N10230, N8773);
buf BUF1 (N10233, N10218);
and AND2 (N10234, N10231, N7966);
and AND3 (N10235, N10227, N3328, N4351);
not NOT1 (N10236, N10234);
and AND3 (N10237, N10210, N9268, N9986);
nor NOR2 (N10238, N10237, N6504);
buf BUF1 (N10239, N10238);
nand NAND3 (N10240, N10221, N7327, N9343);
and AND2 (N10241, N10220, N9311);
and AND3 (N10242, N10239, N7741, N6482);
nand NAND3 (N10243, N10242, N7994, N9040);
buf BUF1 (N10244, N10243);
nand NAND2 (N10245, N10233, N5978);
nand NAND3 (N10246, N10241, N8438, N4276);
nor NOR4 (N10247, N10245, N7398, N6925, N9136);
xor XOR2 (N10248, N10226, N5633);
buf BUF1 (N10249, N10232);
not NOT1 (N10250, N10236);
not NOT1 (N10251, N10246);
and AND4 (N10252, N10251, N6963, N6695, N3949);
not NOT1 (N10253, N10250);
buf BUF1 (N10254, N10247);
nand NAND2 (N10255, N10252, N1182);
or OR4 (N10256, N10244, N7649, N2570, N66);
not NOT1 (N10257, N10253);
not NOT1 (N10258, N10240);
and AND2 (N10259, N10255, N5268);
buf BUF1 (N10260, N10249);
nor NOR3 (N10261, N10248, N4926, N6789);
nor NOR3 (N10262, N10256, N10218, N6418);
nor NOR4 (N10263, N10258, N9234, N874, N3599);
not NOT1 (N10264, N10259);
and AND2 (N10265, N10264, N4153);
not NOT1 (N10266, N10222);
nand NAND3 (N10267, N10229, N5249, N7668);
nor NOR3 (N10268, N10265, N3688, N196);
xor XOR2 (N10269, N10266, N4374);
xor XOR2 (N10270, N10261, N8907);
or OR2 (N10271, N10254, N7811);
and AND3 (N10272, N10260, N8675, N9293);
or OR2 (N10273, N10262, N629);
or OR4 (N10274, N10271, N7834, N7472, N4591);
nand NAND3 (N10275, N10235, N5370, N1178);
xor XOR2 (N10276, N10268, N1707);
buf BUF1 (N10277, N10270);
buf BUF1 (N10278, N10277);
buf BUF1 (N10279, N10273);
buf BUF1 (N10280, N10263);
nand NAND3 (N10281, N10274, N2491, N14);
xor XOR2 (N10282, N10278, N156);
not NOT1 (N10283, N10282);
nand NAND3 (N10284, N10280, N8412, N833);
and AND4 (N10285, N10279, N2449, N6700, N9703);
or OR4 (N10286, N10272, N6047, N6613, N2395);
not NOT1 (N10287, N10269);
nand NAND3 (N10288, N10276, N3644, N979);
not NOT1 (N10289, N10283);
or OR4 (N10290, N10287, N9362, N1206, N3803);
buf BUF1 (N10291, N10286);
buf BUF1 (N10292, N10267);
not NOT1 (N10293, N10257);
xor XOR2 (N10294, N10290, N5015);
not NOT1 (N10295, N10294);
nor NOR4 (N10296, N10292, N1585, N4530, N1386);
and AND2 (N10297, N10295, N3215);
buf BUF1 (N10298, N10288);
not NOT1 (N10299, N10285);
and AND4 (N10300, N10297, N5161, N5658, N39);
and AND3 (N10301, N10300, N3320, N8371);
nor NOR4 (N10302, N10291, N8627, N60, N9727);
nor NOR3 (N10303, N10275, N4350, N9835);
or OR2 (N10304, N10302, N6773);
or OR3 (N10305, N10299, N9335, N6965);
nand NAND4 (N10306, N10281, N345, N3551, N7988);
buf BUF1 (N10307, N10304);
and AND2 (N10308, N10301, N7783);
buf BUF1 (N10309, N10305);
or OR2 (N10310, N10306, N9443);
buf BUF1 (N10311, N10309);
buf BUF1 (N10312, N10289);
or OR4 (N10313, N10308, N3487, N399, N5461);
nand NAND3 (N10314, N10296, N383, N6821);
nor NOR2 (N10315, N10310, N9805);
buf BUF1 (N10316, N10284);
xor XOR2 (N10317, N10303, N9115);
nor NOR4 (N10318, N10312, N3035, N9687, N5897);
xor XOR2 (N10319, N10313, N8316);
and AND2 (N10320, N10319, N7903);
buf BUF1 (N10321, N10314);
or OR3 (N10322, N10315, N10081, N7818);
buf BUF1 (N10323, N10311);
nand NAND2 (N10324, N10323, N2347);
buf BUF1 (N10325, N10320);
nand NAND2 (N10326, N10307, N3349);
and AND2 (N10327, N10325, N1572);
and AND4 (N10328, N10321, N5518, N837, N8207);
not NOT1 (N10329, N10293);
not NOT1 (N10330, N10318);
buf BUF1 (N10331, N10328);
nor NOR3 (N10332, N10316, N3111, N6791);
xor XOR2 (N10333, N10331, N593);
buf BUF1 (N10334, N10332);
and AND2 (N10335, N10329, N5681);
buf BUF1 (N10336, N10335);
buf BUF1 (N10337, N10317);
nand NAND2 (N10338, N10327, N5865);
nor NOR3 (N10339, N10337, N9566, N8381);
not NOT1 (N10340, N10333);
nand NAND3 (N10341, N10298, N9920, N1560);
buf BUF1 (N10342, N10341);
nand NAND4 (N10343, N10324, N3460, N8154, N6213);
nand NAND2 (N10344, N10330, N7222);
and AND2 (N10345, N10326, N2399);
and AND4 (N10346, N10336, N9994, N3654, N2266);
buf BUF1 (N10347, N10338);
or OR3 (N10348, N10342, N3399, N9860);
and AND3 (N10349, N10343, N3303, N1840);
or OR4 (N10350, N10344, N2712, N5008, N5002);
not NOT1 (N10351, N10348);
xor XOR2 (N10352, N10351, N1773);
not NOT1 (N10353, N10339);
and AND2 (N10354, N10349, N7911);
xor XOR2 (N10355, N10346, N4680);
buf BUF1 (N10356, N10350);
nand NAND4 (N10357, N10355, N5687, N8715, N1374);
or OR3 (N10358, N10334, N8726, N6782);
xor XOR2 (N10359, N10345, N3345);
buf BUF1 (N10360, N10357);
or OR3 (N10361, N10353, N3136, N8022);
not NOT1 (N10362, N10340);
or OR4 (N10363, N10362, N1917, N186, N6907);
nor NOR2 (N10364, N10359, N6164);
not NOT1 (N10365, N10322);
nand NAND4 (N10366, N10358, N5627, N8529, N7668);
buf BUF1 (N10367, N10361);
buf BUF1 (N10368, N10364);
nand NAND3 (N10369, N10366, N7177, N6012);
and AND3 (N10370, N10367, N7659, N312);
buf BUF1 (N10371, N10356);
xor XOR2 (N10372, N10370, N6550);
buf BUF1 (N10373, N10347);
not NOT1 (N10374, N10354);
not NOT1 (N10375, N10365);
or OR3 (N10376, N10363, N9670, N353);
or OR2 (N10377, N10373, N6964);
xor XOR2 (N10378, N10372, N3971);
nand NAND4 (N10379, N10374, N7625, N795, N3950);
not NOT1 (N10380, N10379);
nor NOR3 (N10381, N10378, N6919, N793);
or OR3 (N10382, N10380, N7671, N8046);
or OR3 (N10383, N10352, N1012, N4178);
not NOT1 (N10384, N10376);
or OR4 (N10385, N10371, N2470, N507, N9906);
nor NOR4 (N10386, N10383, N3821, N3758, N6823);
and AND3 (N10387, N10360, N6961, N7323);
nand NAND3 (N10388, N10375, N2980, N9854);
buf BUF1 (N10389, N10388);
not NOT1 (N10390, N10382);
nor NOR2 (N10391, N10368, N5090);
and AND2 (N10392, N10391, N6416);
buf BUF1 (N10393, N10389);
buf BUF1 (N10394, N10384);
nor NOR2 (N10395, N10369, N5811);
xor XOR2 (N10396, N10392, N2267);
or OR4 (N10397, N10393, N165, N2344, N4010);
not NOT1 (N10398, N10390);
and AND4 (N10399, N10381, N9099, N153, N2172);
or OR4 (N10400, N10397, N6842, N4819, N7422);
and AND4 (N10401, N10385, N2337, N1281, N780);
and AND4 (N10402, N10399, N4794, N7498, N5550);
xor XOR2 (N10403, N10394, N3520);
nand NAND3 (N10404, N10402, N147, N1172);
or OR3 (N10405, N10395, N10064, N2973);
or OR3 (N10406, N10377, N8203, N8699);
buf BUF1 (N10407, N10396);
nor NOR3 (N10408, N10400, N7795, N4214);
and AND2 (N10409, N10407, N2373);
not NOT1 (N10410, N10406);
nor NOR4 (N10411, N10405, N1725, N2684, N7385);
not NOT1 (N10412, N10411);
nor NOR4 (N10413, N10410, N7255, N9211, N8517);
nand NAND4 (N10414, N10412, N435, N5935, N9752);
xor XOR2 (N10415, N10401, N2297);
and AND2 (N10416, N10414, N8122);
and AND4 (N10417, N10404, N1401, N7708, N6327);
nand NAND4 (N10418, N10415, N4178, N2360, N4055);
xor XOR2 (N10419, N10418, N7449);
nor NOR2 (N10420, N10387, N2016);
not NOT1 (N10421, N10386);
not NOT1 (N10422, N10398);
and AND2 (N10423, N10420, N7822);
xor XOR2 (N10424, N10421, N7063);
xor XOR2 (N10425, N10419, N4632);
or OR3 (N10426, N10416, N2493, N5049);
and AND4 (N10427, N10424, N926, N1224, N6094);
buf BUF1 (N10428, N10417);
buf BUF1 (N10429, N10422);
or OR2 (N10430, N10413, N4295);
not NOT1 (N10431, N10425);
buf BUF1 (N10432, N10423);
nor NOR2 (N10433, N10431, N3305);
xor XOR2 (N10434, N10409, N3298);
buf BUF1 (N10435, N10434);
or OR4 (N10436, N10427, N8230, N2975, N9170);
nor NOR3 (N10437, N10433, N1422, N3490);
not NOT1 (N10438, N10426);
or OR2 (N10439, N10435, N239);
buf BUF1 (N10440, N10432);
not NOT1 (N10441, N10408);
and AND2 (N10442, N10403, N10408);
buf BUF1 (N10443, N10430);
and AND4 (N10444, N10442, N8154, N4776, N476);
or OR3 (N10445, N10429, N4155, N3252);
and AND3 (N10446, N10436, N7856, N1694);
and AND4 (N10447, N10441, N655, N2475, N5416);
nor NOR4 (N10448, N10446, N172, N1475, N4841);
nand NAND3 (N10449, N10437, N10255, N3338);
nor NOR4 (N10450, N10448, N4984, N9734, N159);
or OR2 (N10451, N10449, N1712);
not NOT1 (N10452, N10440);
not NOT1 (N10453, N10447);
not NOT1 (N10454, N10450);
not NOT1 (N10455, N10428);
xor XOR2 (N10456, N10451, N9616);
not NOT1 (N10457, N10445);
and AND4 (N10458, N10439, N10226, N10372, N9304);
nand NAND4 (N10459, N10457, N9989, N3155, N3156);
nand NAND4 (N10460, N10455, N3045, N4873, N753);
not NOT1 (N10461, N10460);
not NOT1 (N10462, N10458);
not NOT1 (N10463, N10459);
or OR2 (N10464, N10461, N1270);
nor NOR3 (N10465, N10456, N7584, N5895);
not NOT1 (N10466, N10465);
xor XOR2 (N10467, N10444, N6859);
nand NAND4 (N10468, N10438, N2039, N7771, N314);
buf BUF1 (N10469, N10468);
or OR2 (N10470, N10464, N1295);
nand NAND3 (N10471, N10462, N4567, N8411);
or OR3 (N10472, N10453, N4790, N10367);
and AND2 (N10473, N10472, N6124);
nor NOR2 (N10474, N10469, N7047);
xor XOR2 (N10475, N10443, N1385);
nand NAND3 (N10476, N10474, N6103, N4580);
nand NAND3 (N10477, N10471, N2851, N7382);
xor XOR2 (N10478, N10476, N7307);
buf BUF1 (N10479, N10452);
nor NOR4 (N10480, N10454, N274, N8426, N4683);
xor XOR2 (N10481, N10479, N9043);
nor NOR4 (N10482, N10470, N7359, N1130, N3542);
xor XOR2 (N10483, N10477, N6574);
or OR3 (N10484, N10480, N2593, N8262);
not NOT1 (N10485, N10484);
and AND2 (N10486, N10473, N1480);
and AND2 (N10487, N10466, N6171);
nand NAND4 (N10488, N10483, N9251, N2821, N2499);
or OR2 (N10489, N10481, N3900);
buf BUF1 (N10490, N10489);
not NOT1 (N10491, N10487);
nor NOR4 (N10492, N10463, N8722, N8777, N8809);
or OR4 (N10493, N10478, N7626, N9298, N1861);
xor XOR2 (N10494, N10486, N4458);
xor XOR2 (N10495, N10482, N4691);
or OR2 (N10496, N10467, N2696);
buf BUF1 (N10497, N10493);
buf BUF1 (N10498, N10496);
xor XOR2 (N10499, N10490, N7075);
xor XOR2 (N10500, N10498, N4439);
not NOT1 (N10501, N10500);
xor XOR2 (N10502, N10494, N1041);
not NOT1 (N10503, N10501);
xor XOR2 (N10504, N10492, N2908);
or OR4 (N10505, N10502, N1714, N5887, N5234);
xor XOR2 (N10506, N10488, N2985);
nor NOR3 (N10507, N10504, N7249, N4625);
not NOT1 (N10508, N10506);
not NOT1 (N10509, N10499);
not NOT1 (N10510, N10507);
nor NOR3 (N10511, N10485, N7520, N10343);
buf BUF1 (N10512, N10508);
not NOT1 (N10513, N10497);
and AND2 (N10514, N10503, N8858);
nand NAND2 (N10515, N10491, N5029);
and AND3 (N10516, N10510, N1934, N3158);
or OR4 (N10517, N10509, N6588, N10463, N2448);
xor XOR2 (N10518, N10513, N2506);
not NOT1 (N10519, N10515);
or OR3 (N10520, N10516, N3287, N1795);
nand NAND3 (N10521, N10517, N5401, N7618);
or OR2 (N10522, N10505, N6630);
not NOT1 (N10523, N10512);
xor XOR2 (N10524, N10495, N3792);
xor XOR2 (N10525, N10523, N7787);
nor NOR2 (N10526, N10475, N100);
nor NOR4 (N10527, N10521, N547, N4246, N5073);
nor NOR4 (N10528, N10522, N2001, N7662, N8948);
nor NOR2 (N10529, N10528, N1454);
xor XOR2 (N10530, N10519, N4986);
and AND3 (N10531, N10518, N3716, N8208);
nor NOR2 (N10532, N10527, N9031);
not NOT1 (N10533, N10511);
buf BUF1 (N10534, N10514);
buf BUF1 (N10535, N10531);
xor XOR2 (N10536, N10532, N4225);
buf BUF1 (N10537, N10520);
nand NAND2 (N10538, N10530, N679);
nor NOR3 (N10539, N10524, N6892, N5674);
or OR4 (N10540, N10537, N1716, N6200, N7410);
buf BUF1 (N10541, N10538);
not NOT1 (N10542, N10525);
nor NOR3 (N10543, N10526, N10481, N10029);
buf BUF1 (N10544, N10540);
nand NAND4 (N10545, N10544, N7942, N974, N9714);
nor NOR3 (N10546, N10545, N2598, N9396);
or OR3 (N10547, N10535, N3779, N2247);
buf BUF1 (N10548, N10543);
nor NOR2 (N10549, N10529, N9753);
nor NOR2 (N10550, N10541, N7475);
nand NAND4 (N10551, N10550, N5384, N3953, N10027);
and AND4 (N10552, N10534, N1130, N6992, N3760);
nor NOR2 (N10553, N10542, N6850);
xor XOR2 (N10554, N10547, N9074);
nand NAND2 (N10555, N10549, N7362);
not NOT1 (N10556, N10554);
buf BUF1 (N10557, N10552);
and AND2 (N10558, N10548, N4908);
nand NAND3 (N10559, N10533, N6883, N4562);
or OR3 (N10560, N10559, N9612, N3253);
or OR3 (N10561, N10556, N8, N1930);
not NOT1 (N10562, N10539);
xor XOR2 (N10563, N10551, N6592);
not NOT1 (N10564, N10536);
not NOT1 (N10565, N10555);
nand NAND3 (N10566, N10564, N421, N3252);
xor XOR2 (N10567, N10563, N5750);
and AND4 (N10568, N10562, N1803, N9236, N146);
or OR3 (N10569, N10546, N7471, N1634);
nand NAND3 (N10570, N10560, N7703, N6859);
xor XOR2 (N10571, N10567, N8638);
nand NAND4 (N10572, N10568, N8319, N4755, N806);
nor NOR2 (N10573, N10572, N4996);
xor XOR2 (N10574, N10569, N672);
and AND2 (N10575, N10561, N5793);
xor XOR2 (N10576, N10566, N3783);
buf BUF1 (N10577, N10571);
nor NOR4 (N10578, N10574, N8103, N3304, N6522);
nor NOR3 (N10579, N10573, N9703, N2053);
or OR4 (N10580, N10553, N6354, N7731, N1065);
xor XOR2 (N10581, N10575, N6220);
nand NAND4 (N10582, N10578, N2246, N3867, N2487);
not NOT1 (N10583, N10570);
not NOT1 (N10584, N10558);
or OR4 (N10585, N10577, N10537, N1436, N10151);
nor NOR3 (N10586, N10565, N1762, N3266);
and AND2 (N10587, N10586, N2966);
nor NOR3 (N10588, N10582, N4953, N5609);
buf BUF1 (N10589, N10581);
and AND2 (N10590, N10585, N6187);
buf BUF1 (N10591, N10583);
xor XOR2 (N10592, N10588, N4979);
or OR2 (N10593, N10590, N4613);
nor NOR4 (N10594, N10576, N996, N9630, N5424);
nor NOR4 (N10595, N10594, N4839, N10370, N5918);
not NOT1 (N10596, N10595);
nand NAND2 (N10597, N10584, N2648);
or OR3 (N10598, N10597, N1012, N7245);
nand NAND2 (N10599, N10591, N3757);
xor XOR2 (N10600, N10599, N7159);
nor NOR4 (N10601, N10596, N10230, N3888, N2405);
xor XOR2 (N10602, N10592, N8632);
and AND2 (N10603, N10601, N2780);
not NOT1 (N10604, N10603);
or OR3 (N10605, N10557, N8373, N9639);
nand NAND2 (N10606, N10605, N878);
and AND2 (N10607, N10579, N9161);
nand NAND4 (N10608, N10593, N5524, N3052, N556);
or OR4 (N10609, N10604, N3740, N4679, N8749);
xor XOR2 (N10610, N10580, N10203);
or OR4 (N10611, N10606, N7149, N3771, N7159);
not NOT1 (N10612, N10602);
xor XOR2 (N10613, N10607, N8206);
nor NOR4 (N10614, N10609, N6521, N6256, N5604);
not NOT1 (N10615, N10589);
buf BUF1 (N10616, N10587);
nor NOR2 (N10617, N10598, N3143);
nand NAND2 (N10618, N10617, N2139);
and AND4 (N10619, N10613, N6550, N2676, N6794);
nor NOR4 (N10620, N10610, N2157, N6169, N2516);
buf BUF1 (N10621, N10608);
xor XOR2 (N10622, N10619, N1062);
not NOT1 (N10623, N10621);
xor XOR2 (N10624, N10612, N5879);
buf BUF1 (N10625, N10624);
and AND4 (N10626, N10622, N3553, N2760, N5898);
nand NAND4 (N10627, N10611, N4670, N2165, N3296);
and AND4 (N10628, N10625, N4549, N7017, N4280);
buf BUF1 (N10629, N10626);
nand NAND3 (N10630, N10618, N6277, N9803);
or OR2 (N10631, N10614, N3570);
nand NAND3 (N10632, N10629, N4942, N4864);
or OR2 (N10633, N10632, N8777);
xor XOR2 (N10634, N10627, N2093);
or OR4 (N10635, N10620, N8281, N922, N6334);
nor NOR3 (N10636, N10616, N10273, N7945);
buf BUF1 (N10637, N10630);
and AND3 (N10638, N10637, N4855, N9120);
buf BUF1 (N10639, N10638);
xor XOR2 (N10640, N10600, N4031);
buf BUF1 (N10641, N10623);
buf BUF1 (N10642, N10628);
not NOT1 (N10643, N10615);
nor NOR3 (N10644, N10640, N6191, N8331);
nor NOR3 (N10645, N10633, N25, N2298);
not NOT1 (N10646, N10641);
nand NAND3 (N10647, N10631, N1419, N7987);
not NOT1 (N10648, N10643);
nor NOR2 (N10649, N10636, N2969);
or OR4 (N10650, N10635, N6841, N6548, N1413);
not NOT1 (N10651, N10648);
and AND4 (N10652, N10639, N10502, N8910, N2577);
buf BUF1 (N10653, N10645);
or OR2 (N10654, N10651, N8339);
not NOT1 (N10655, N10654);
xor XOR2 (N10656, N10634, N7775);
and AND3 (N10657, N10647, N4574, N7857);
buf BUF1 (N10658, N10652);
buf BUF1 (N10659, N10642);
nand NAND2 (N10660, N10644, N4849);
and AND4 (N10661, N10649, N1682, N9651, N6453);
nor NOR2 (N10662, N10657, N2381);
and AND4 (N10663, N10656, N4394, N3558, N8991);
and AND3 (N10664, N10650, N965, N6106);
nor NOR4 (N10665, N10662, N785, N3834, N9151);
not NOT1 (N10666, N10659);
and AND2 (N10667, N10663, N10235);
or OR2 (N10668, N10658, N7165);
xor XOR2 (N10669, N10668, N8474);
nand NAND3 (N10670, N10664, N8077, N5412);
nand NAND2 (N10671, N10665, N3923);
xor XOR2 (N10672, N10655, N4325);
and AND3 (N10673, N10671, N10280, N1937);
nor NOR4 (N10674, N10661, N4057, N8634, N10268);
xor XOR2 (N10675, N10646, N8432);
or OR3 (N10676, N10660, N7436, N1897);
xor XOR2 (N10677, N10667, N1518);
nor NOR3 (N10678, N10669, N6009, N440);
or OR2 (N10679, N10653, N2224);
xor XOR2 (N10680, N10674, N4416);
or OR2 (N10681, N10670, N7842);
and AND4 (N10682, N10677, N2852, N6534, N525);
nor NOR2 (N10683, N10679, N2562);
xor XOR2 (N10684, N10672, N4769);
buf BUF1 (N10685, N10676);
buf BUF1 (N10686, N10675);
and AND2 (N10687, N10666, N9862);
xor XOR2 (N10688, N10687, N8868);
nand NAND4 (N10689, N10673, N5987, N5780, N2129);
and AND2 (N10690, N10683, N10552);
or OR3 (N10691, N10681, N1568, N9425);
or OR2 (N10692, N10688, N1940);
xor XOR2 (N10693, N10689, N9649);
nand NAND3 (N10694, N10680, N951, N2535);
buf BUF1 (N10695, N10684);
not NOT1 (N10696, N10693);
not NOT1 (N10697, N10685);
nand NAND4 (N10698, N10690, N7400, N7035, N6883);
not NOT1 (N10699, N10695);
not NOT1 (N10700, N10686);
or OR3 (N10701, N10700, N1202, N2421);
not NOT1 (N10702, N10692);
and AND2 (N10703, N10699, N8636);
xor XOR2 (N10704, N10682, N3287);
xor XOR2 (N10705, N10696, N2106);
nand NAND3 (N10706, N10704, N1829, N9066);
nor NOR3 (N10707, N10702, N9559, N4327);
buf BUF1 (N10708, N10703);
and AND3 (N10709, N10707, N2870, N10662);
xor XOR2 (N10710, N10708, N704);
xor XOR2 (N10711, N10710, N1557);
buf BUF1 (N10712, N10705);
or OR2 (N10713, N10709, N51);
xor XOR2 (N10714, N10712, N3105);
or OR4 (N10715, N10713, N5681, N10640, N3195);
and AND2 (N10716, N10701, N7636);
buf BUF1 (N10717, N10706);
nand NAND3 (N10718, N10691, N8117, N4534);
not NOT1 (N10719, N10715);
nor NOR3 (N10720, N10716, N6528, N2214);
nor NOR4 (N10721, N10720, N8240, N5229, N3339);
nand NAND3 (N10722, N10678, N7159, N475);
xor XOR2 (N10723, N10694, N3900);
xor XOR2 (N10724, N10717, N148);
and AND4 (N10725, N10718, N1776, N8993, N2274);
xor XOR2 (N10726, N10723, N3508);
nor NOR4 (N10727, N10711, N8176, N6007, N7236);
buf BUF1 (N10728, N10726);
nor NOR4 (N10729, N10698, N10192, N8600, N3564);
and AND4 (N10730, N10719, N9351, N2616, N4621);
xor XOR2 (N10731, N10724, N2049);
not NOT1 (N10732, N10731);
or OR2 (N10733, N10728, N9085);
nor NOR2 (N10734, N10697, N7839);
and AND2 (N10735, N10732, N10310);
buf BUF1 (N10736, N10730);
nor NOR3 (N10737, N10722, N2866, N2918);
and AND2 (N10738, N10721, N311);
buf BUF1 (N10739, N10725);
not NOT1 (N10740, N10733);
or OR3 (N10741, N10740, N157, N4199);
nand NAND3 (N10742, N10736, N5723, N9756);
not NOT1 (N10743, N10742);
not NOT1 (N10744, N10737);
nand NAND4 (N10745, N10743, N8718, N4987, N6907);
buf BUF1 (N10746, N10729);
nor NOR3 (N10747, N10746, N6665, N951);
xor XOR2 (N10748, N10739, N1859);
or OR4 (N10749, N10744, N10320, N9602, N3467);
and AND3 (N10750, N10748, N4727, N8596);
nand NAND4 (N10751, N10735, N1565, N5407, N7787);
or OR2 (N10752, N10738, N9742);
nand NAND4 (N10753, N10750, N1490, N8324, N9059);
and AND2 (N10754, N10734, N2027);
or OR4 (N10755, N10754, N8409, N8561, N8106);
not NOT1 (N10756, N10753);
and AND4 (N10757, N10727, N650, N7157, N2545);
or OR4 (N10758, N10751, N10539, N7944, N322);
or OR4 (N10759, N10747, N8303, N5990, N8298);
not NOT1 (N10760, N10745);
buf BUF1 (N10761, N10759);
or OR3 (N10762, N10755, N7107, N8461);
and AND2 (N10763, N10756, N1019);
nor NOR3 (N10764, N10752, N6735, N7619);
nand NAND2 (N10765, N10757, N685);
xor XOR2 (N10766, N10764, N4719);
nor NOR3 (N10767, N10760, N219, N110);
buf BUF1 (N10768, N10765);
nor NOR2 (N10769, N10741, N9535);
nand NAND3 (N10770, N10769, N8535, N7626);
xor XOR2 (N10771, N10749, N851);
and AND4 (N10772, N10766, N3072, N4802, N10441);
xor XOR2 (N10773, N10714, N2576);
nand NAND2 (N10774, N10768, N5047);
or OR3 (N10775, N10772, N9495, N1047);
not NOT1 (N10776, N10773);
or OR4 (N10777, N10775, N9608, N3114, N5032);
or OR2 (N10778, N10770, N4423);
not NOT1 (N10779, N10771);
or OR2 (N10780, N10774, N7570);
nand NAND3 (N10781, N10763, N4839, N4183);
nand NAND2 (N10782, N10761, N1396);
and AND4 (N10783, N10780, N8930, N5187, N9034);
not NOT1 (N10784, N10781);
buf BUF1 (N10785, N10782);
nor NOR3 (N10786, N10777, N4997, N968);
and AND3 (N10787, N10776, N2, N34);
or OR4 (N10788, N10758, N6238, N10742, N3549);
xor XOR2 (N10789, N10787, N6936);
not NOT1 (N10790, N10788);
and AND3 (N10791, N10783, N5623, N163);
xor XOR2 (N10792, N10791, N7061);
and AND4 (N10793, N10784, N10124, N7069, N8345);
buf BUF1 (N10794, N10793);
not NOT1 (N10795, N10785);
and AND2 (N10796, N10762, N8176);
and AND3 (N10797, N10789, N7861, N5769);
not NOT1 (N10798, N10795);
or OR2 (N10799, N10786, N7511);
nand NAND3 (N10800, N10779, N6624, N8453);
nand NAND4 (N10801, N10796, N4273, N3044, N3174);
buf BUF1 (N10802, N10798);
buf BUF1 (N10803, N10797);
not NOT1 (N10804, N10799);
buf BUF1 (N10805, N10803);
and AND2 (N10806, N10802, N7808);
not NOT1 (N10807, N10805);
xor XOR2 (N10808, N10767, N8002);
nand NAND3 (N10809, N10792, N7324, N3563);
or OR2 (N10810, N10800, N6924);
nand NAND3 (N10811, N10806, N1989, N7076);
not NOT1 (N10812, N10809);
buf BUF1 (N10813, N10778);
and AND3 (N10814, N10808, N8257, N2622);
nand NAND3 (N10815, N10811, N10021, N7755);
not NOT1 (N10816, N10813);
or OR4 (N10817, N10810, N6089, N6309, N5280);
not NOT1 (N10818, N10815);
and AND4 (N10819, N10814, N8282, N4206, N5353);
nor NOR3 (N10820, N10790, N9784, N10112);
nand NAND2 (N10821, N10816, N6943);
nand NAND2 (N10822, N10820, N10545);
and AND4 (N10823, N10817, N10110, N1300, N278);
not NOT1 (N10824, N10804);
and AND2 (N10825, N10807, N7048);
nor NOR4 (N10826, N10825, N6876, N3730, N6445);
nand NAND2 (N10827, N10818, N266);
xor XOR2 (N10828, N10819, N9791);
nand NAND3 (N10829, N10828, N4134, N1205);
nor NOR4 (N10830, N10821, N6922, N222, N5702);
or OR3 (N10831, N10827, N9931, N10247);
nand NAND2 (N10832, N10826, N8509);
not NOT1 (N10833, N10812);
and AND3 (N10834, N10831, N7056, N3893);
not NOT1 (N10835, N10830);
not NOT1 (N10836, N10824);
not NOT1 (N10837, N10832);
nor NOR4 (N10838, N10836, N9487, N6730, N1369);
not NOT1 (N10839, N10838);
buf BUF1 (N10840, N10835);
xor XOR2 (N10841, N10794, N3753);
and AND4 (N10842, N10833, N6251, N115, N2760);
or OR2 (N10843, N10822, N185);
nand NAND4 (N10844, N10834, N2774, N4860, N3389);
or OR2 (N10845, N10841, N1065);
nor NOR2 (N10846, N10840, N1361);
buf BUF1 (N10847, N10845);
and AND4 (N10848, N10846, N7043, N3135, N5703);
nor NOR4 (N10849, N10829, N9971, N10803, N2734);
or OR4 (N10850, N10848, N1525, N6027, N7363);
xor XOR2 (N10851, N10842, N3732);
buf BUF1 (N10852, N10847);
buf BUF1 (N10853, N10843);
nor NOR3 (N10854, N10849, N3193, N2870);
xor XOR2 (N10855, N10850, N2681);
or OR4 (N10856, N10855, N6862, N1828, N906);
not NOT1 (N10857, N10823);
nand NAND2 (N10858, N10853, N5488);
nor NOR2 (N10859, N10852, N626);
not NOT1 (N10860, N10837);
nor NOR2 (N10861, N10844, N3201);
and AND2 (N10862, N10858, N2071);
nor NOR4 (N10863, N10801, N6838, N7730, N9242);
and AND4 (N10864, N10860, N5183, N3532, N1535);
xor XOR2 (N10865, N10839, N9634);
or OR3 (N10866, N10864, N1122, N5098);
nor NOR4 (N10867, N10856, N10612, N6862, N7813);
buf BUF1 (N10868, N10865);
and AND4 (N10869, N10851, N8809, N6718, N2239);
and AND3 (N10870, N10862, N7438, N3815);
not NOT1 (N10871, N10867);
xor XOR2 (N10872, N10868, N8586);
and AND4 (N10873, N10854, N8874, N3398, N1886);
not NOT1 (N10874, N10859);
xor XOR2 (N10875, N10857, N10081);
or OR3 (N10876, N10873, N4214, N9416);
not NOT1 (N10877, N10872);
buf BUF1 (N10878, N10871);
xor XOR2 (N10879, N10878, N1259);
not NOT1 (N10880, N10874);
and AND3 (N10881, N10866, N940, N195);
nand NAND4 (N10882, N10881, N10410, N155, N2971);
not NOT1 (N10883, N10875);
not NOT1 (N10884, N10870);
nor NOR3 (N10885, N10879, N7860, N8657);
nor NOR3 (N10886, N10876, N8826, N3231);
nor NOR3 (N10887, N10863, N2876, N4868);
and AND4 (N10888, N10861, N2121, N3123, N6656);
and AND4 (N10889, N10882, N2192, N9648, N10538);
or OR4 (N10890, N10884, N5354, N6460, N4957);
nand NAND2 (N10891, N10880, N7908);
not NOT1 (N10892, N10889);
and AND4 (N10893, N10888, N723, N4714, N6114);
nor NOR2 (N10894, N10892, N5678);
not NOT1 (N10895, N10869);
or OR3 (N10896, N10887, N6502, N4514);
xor XOR2 (N10897, N10893, N7018);
nor NOR4 (N10898, N10890, N961, N4359, N1032);
nor NOR3 (N10899, N10886, N9037, N4202);
or OR4 (N10900, N10897, N4986, N463, N7450);
buf BUF1 (N10901, N10896);
xor XOR2 (N10902, N10891, N4988);
and AND3 (N10903, N10885, N2053, N5158);
buf BUF1 (N10904, N10902);
nor NOR4 (N10905, N10900, N3908, N4229, N4046);
xor XOR2 (N10906, N10895, N9218);
and AND3 (N10907, N10904, N1485, N7225);
and AND3 (N10908, N10883, N1480, N9362);
nor NOR3 (N10909, N10908, N208, N4290);
nand NAND3 (N10910, N10898, N5266, N6816);
not NOT1 (N10911, N10899);
nor NOR2 (N10912, N10901, N4802);
and AND4 (N10913, N10909, N4283, N3719, N2148);
xor XOR2 (N10914, N10903, N1864);
not NOT1 (N10915, N10911);
or OR4 (N10916, N10906, N6614, N4329, N7429);
or OR3 (N10917, N10913, N8140, N9112);
nand NAND2 (N10918, N10894, N1647);
buf BUF1 (N10919, N10912);
buf BUF1 (N10920, N10915);
or OR2 (N10921, N10910, N6679);
xor XOR2 (N10922, N10916, N6526);
xor XOR2 (N10923, N10877, N10867);
buf BUF1 (N10924, N10907);
and AND4 (N10925, N10917, N8847, N1256, N9955);
nor NOR2 (N10926, N10914, N7004);
buf BUF1 (N10927, N10921);
xor XOR2 (N10928, N10926, N10443);
nor NOR2 (N10929, N10925, N4160);
not NOT1 (N10930, N10927);
or OR4 (N10931, N10918, N10590, N8217, N7343);
xor XOR2 (N10932, N10924, N10410);
xor XOR2 (N10933, N10922, N120);
xor XOR2 (N10934, N10928, N3644);
buf BUF1 (N10935, N10929);
nand NAND4 (N10936, N10933, N9280, N5151, N9175);
and AND4 (N10937, N10920, N4291, N273, N726);
buf BUF1 (N10938, N10937);
buf BUF1 (N10939, N10935);
and AND3 (N10940, N10919, N10197, N5277);
and AND4 (N10941, N10931, N10291, N10543, N10277);
and AND3 (N10942, N10930, N2691, N9345);
xor XOR2 (N10943, N10923, N9052);
nor NOR3 (N10944, N10934, N4038, N9977);
or OR2 (N10945, N10941, N672);
nand NAND2 (N10946, N10936, N10586);
nand NAND2 (N10947, N10938, N2820);
and AND4 (N10948, N10943, N9207, N8313, N10354);
nand NAND2 (N10949, N10905, N6297);
nand NAND2 (N10950, N10932, N9732);
xor XOR2 (N10951, N10947, N2321);
nor NOR3 (N10952, N10939, N1030, N5755);
xor XOR2 (N10953, N10944, N9370);
and AND2 (N10954, N10949, N5764);
xor XOR2 (N10955, N10951, N8053);
or OR2 (N10956, N10953, N8330);
not NOT1 (N10957, N10952);
buf BUF1 (N10958, N10954);
nand NAND4 (N10959, N10940, N6092, N7887, N4053);
not NOT1 (N10960, N10955);
or OR2 (N10961, N10960, N10750);
nor NOR3 (N10962, N10959, N6017, N5012);
nor NOR3 (N10963, N10961, N6013, N2498);
nor NOR2 (N10964, N10958, N409);
nand NAND3 (N10965, N10964, N1020, N5327);
xor XOR2 (N10966, N10945, N5590);
and AND2 (N10967, N10950, N7885);
xor XOR2 (N10968, N10962, N1697);
nor NOR4 (N10969, N10942, N4104, N9755, N8150);
xor XOR2 (N10970, N10957, N773);
xor XOR2 (N10971, N10969, N2621);
nor NOR2 (N10972, N10948, N8410);
not NOT1 (N10973, N10965);
xor XOR2 (N10974, N10970, N1467);
not NOT1 (N10975, N10974);
nand NAND4 (N10976, N10972, N9080, N4309, N10027);
and AND3 (N10977, N10946, N8346, N1002);
xor XOR2 (N10978, N10975, N8874);
buf BUF1 (N10979, N10971);
not NOT1 (N10980, N10973);
xor XOR2 (N10981, N10963, N8144);
xor XOR2 (N10982, N10978, N174);
and AND2 (N10983, N10966, N9382);
or OR3 (N10984, N10983, N8020, N5801);
not NOT1 (N10985, N10982);
and AND3 (N10986, N10980, N497, N4528);
nor NOR4 (N10987, N10986, N8996, N9230, N8449);
xor XOR2 (N10988, N10985, N8420);
and AND3 (N10989, N10987, N8395, N680);
buf BUF1 (N10990, N10977);
nand NAND4 (N10991, N10979, N10677, N4372, N7469);
buf BUF1 (N10992, N10981);
xor XOR2 (N10993, N10967, N4284);
nor NOR3 (N10994, N10988, N5297, N7273);
and AND3 (N10995, N10991, N10433, N8203);
and AND2 (N10996, N10995, N69);
and AND3 (N10997, N10968, N210, N1620);
nand NAND4 (N10998, N10997, N1178, N8172, N2969);
or OR4 (N10999, N10956, N1149, N7720, N8988);
xor XOR2 (N11000, N10990, N10567);
not NOT1 (N11001, N10976);
xor XOR2 (N11002, N10998, N3966);
xor XOR2 (N11003, N10993, N6153);
nor NOR3 (N11004, N10984, N1859, N10505);
buf BUF1 (N11005, N10996);
nand NAND3 (N11006, N11001, N4142, N2240);
buf BUF1 (N11007, N11006);
and AND2 (N11008, N10999, N6220);
and AND2 (N11009, N11003, N7498);
nor NOR3 (N11010, N10992, N8577, N8169);
xor XOR2 (N11011, N11005, N5860);
not NOT1 (N11012, N11000);
and AND3 (N11013, N11010, N4103, N743);
or OR4 (N11014, N11004, N4802, N2774, N3312);
not NOT1 (N11015, N11002);
not NOT1 (N11016, N11009);
or OR2 (N11017, N10994, N2167);
buf BUF1 (N11018, N11008);
or OR2 (N11019, N11011, N716);
or OR4 (N11020, N11017, N10717, N1039, N4512);
and AND2 (N11021, N11012, N1511);
nand NAND3 (N11022, N11014, N6870, N5109);
or OR2 (N11023, N11020, N6603);
buf BUF1 (N11024, N11018);
not NOT1 (N11025, N11007);
xor XOR2 (N11026, N11022, N9112);
not NOT1 (N11027, N11013);
not NOT1 (N11028, N11024);
or OR4 (N11029, N11016, N3855, N5939, N2290);
nor NOR4 (N11030, N11023, N6726, N7119, N836);
nor NOR4 (N11031, N11028, N9013, N10127, N1779);
nand NAND3 (N11032, N10989, N10683, N5581);
not NOT1 (N11033, N11031);
nor NOR4 (N11034, N11030, N7145, N7320, N3384);
or OR3 (N11035, N11025, N7546, N9348);
xor XOR2 (N11036, N11033, N7234);
or OR2 (N11037, N11036, N9275);
nor NOR3 (N11038, N11015, N3509, N5771);
or OR4 (N11039, N11032, N8937, N3072, N3252);
and AND3 (N11040, N11034, N10913, N2411);
or OR3 (N11041, N11037, N9064, N8322);
not NOT1 (N11042, N11029);
and AND2 (N11043, N11035, N7343);
xor XOR2 (N11044, N11027, N9268);
or OR2 (N11045, N11044, N5101);
xor XOR2 (N11046, N11021, N9809);
nand NAND4 (N11047, N11040, N6240, N4511, N2422);
xor XOR2 (N11048, N11046, N9944);
xor XOR2 (N11049, N11019, N6178);
xor XOR2 (N11050, N11039, N3736);
buf BUF1 (N11051, N11050);
or OR3 (N11052, N11047, N4118, N2695);
nor NOR2 (N11053, N11049, N6122);
buf BUF1 (N11054, N11052);
buf BUF1 (N11055, N11042);
buf BUF1 (N11056, N11045);
not NOT1 (N11057, N11053);
nand NAND2 (N11058, N11048, N4152);
xor XOR2 (N11059, N11026, N10848);
xor XOR2 (N11060, N11058, N7294);
nor NOR3 (N11061, N11055, N4424, N6947);
nor NOR3 (N11062, N11043, N6466, N47);
xor XOR2 (N11063, N11041, N7676);
and AND4 (N11064, N11060, N5147, N4485, N3557);
nor NOR3 (N11065, N11056, N9545, N8693);
and AND2 (N11066, N11062, N7703);
nor NOR2 (N11067, N11064, N10819);
or OR3 (N11068, N11061, N8354, N7389);
xor XOR2 (N11069, N11066, N9482);
not NOT1 (N11070, N11057);
not NOT1 (N11071, N11069);
nor NOR2 (N11072, N11071, N5412);
xor XOR2 (N11073, N11063, N8156);
xor XOR2 (N11074, N11065, N10789);
nor NOR4 (N11075, N11038, N7727, N8222, N3230);
nor NOR4 (N11076, N11051, N6148, N6358, N6326);
and AND2 (N11077, N11070, N1581);
nor NOR3 (N11078, N11073, N7156, N9618);
not NOT1 (N11079, N11074);
nor NOR3 (N11080, N11068, N9060, N10829);
and AND2 (N11081, N11054, N5709);
or OR4 (N11082, N11077, N1485, N8930, N2227);
buf BUF1 (N11083, N11081);
or OR4 (N11084, N11080, N4553, N4146, N9533);
or OR4 (N11085, N11083, N8626, N9169, N4952);
not NOT1 (N11086, N11085);
and AND3 (N11087, N11059, N10936, N10692);
xor XOR2 (N11088, N11072, N314);
nand NAND3 (N11089, N11084, N920, N9678);
or OR3 (N11090, N11079, N8854, N9215);
and AND4 (N11091, N11067, N3968, N4461, N5584);
and AND2 (N11092, N11091, N4181);
and AND4 (N11093, N11082, N10960, N4978, N8194);
buf BUF1 (N11094, N11088);
buf BUF1 (N11095, N11090);
nand NAND4 (N11096, N11086, N5547, N3103, N2325);
buf BUF1 (N11097, N11096);
xor XOR2 (N11098, N11095, N4490);
or OR4 (N11099, N11094, N6446, N3521, N8048);
and AND3 (N11100, N11097, N6590, N9313);
nor NOR4 (N11101, N11076, N6829, N2933, N10689);
not NOT1 (N11102, N11092);
not NOT1 (N11103, N11100);
or OR3 (N11104, N11099, N3377, N9403);
and AND3 (N11105, N11102, N8377, N2923);
and AND3 (N11106, N11087, N3898, N172);
not NOT1 (N11107, N11103);
not NOT1 (N11108, N11105);
nor NOR4 (N11109, N11104, N649, N8781, N5897);
buf BUF1 (N11110, N11089);
nand NAND4 (N11111, N11106, N9353, N8090, N2604);
xor XOR2 (N11112, N11111, N3562);
buf BUF1 (N11113, N11078);
xor XOR2 (N11114, N11110, N4957);
nor NOR4 (N11115, N11108, N8915, N5990, N5933);
buf BUF1 (N11116, N11112);
nand NAND3 (N11117, N11116, N6224, N6124);
buf BUF1 (N11118, N11075);
and AND2 (N11119, N11098, N3949);
or OR2 (N11120, N11107, N8243);
and AND4 (N11121, N11118, N1548, N341, N6454);
not NOT1 (N11122, N11121);
xor XOR2 (N11123, N11109, N763);
xor XOR2 (N11124, N11122, N608);
nand NAND3 (N11125, N11093, N7826, N2696);
buf BUF1 (N11126, N11124);
xor XOR2 (N11127, N11113, N8324);
not NOT1 (N11128, N11127);
not NOT1 (N11129, N11126);
buf BUF1 (N11130, N11123);
not NOT1 (N11131, N11119);
nand NAND3 (N11132, N11115, N755, N3959);
xor XOR2 (N11133, N11101, N2197);
not NOT1 (N11134, N11132);
buf BUF1 (N11135, N11125);
xor XOR2 (N11136, N11114, N1978);
and AND4 (N11137, N11134, N8497, N8380, N4587);
nor NOR2 (N11138, N11129, N8740);
nor NOR4 (N11139, N11135, N3512, N5546, N1870);
nand NAND2 (N11140, N11137, N10824);
buf BUF1 (N11141, N11136);
xor XOR2 (N11142, N11120, N10285);
nand NAND2 (N11143, N11140, N494);
or OR4 (N11144, N11139, N9868, N7161, N1294);
and AND4 (N11145, N11142, N51, N4434, N5754);
or OR2 (N11146, N11143, N8000);
not NOT1 (N11147, N11117);
nand NAND2 (N11148, N11141, N10183);
buf BUF1 (N11149, N11128);
or OR2 (N11150, N11130, N3506);
or OR3 (N11151, N11148, N7069, N6475);
xor XOR2 (N11152, N11151, N1994);
not NOT1 (N11153, N11138);
not NOT1 (N11154, N11145);
nand NAND4 (N11155, N11144, N2653, N8068, N460);
xor XOR2 (N11156, N11152, N3368);
and AND3 (N11157, N11146, N9882, N3673);
and AND2 (N11158, N11156, N44);
and AND2 (N11159, N11155, N2110);
nor NOR3 (N11160, N11153, N4910, N4432);
xor XOR2 (N11161, N11147, N9009);
nor NOR2 (N11162, N11154, N1191);
nand NAND3 (N11163, N11161, N9814, N6767);
or OR4 (N11164, N11157, N449, N11002, N7847);
nor NOR3 (N11165, N11158, N214, N9912);
or OR2 (N11166, N11150, N6009);
xor XOR2 (N11167, N11149, N3180);
nand NAND3 (N11168, N11165, N6983, N10105);
xor XOR2 (N11169, N11164, N4057);
nor NOR2 (N11170, N11169, N376);
or OR2 (N11171, N11170, N2083);
nor NOR3 (N11172, N11166, N10375, N3121);
not NOT1 (N11173, N11172);
nor NOR2 (N11174, N11162, N4803);
and AND2 (N11175, N11160, N6968);
nor NOR4 (N11176, N11131, N7150, N8573, N6860);
xor XOR2 (N11177, N11168, N6345);
nand NAND2 (N11178, N11173, N4617);
buf BUF1 (N11179, N11178);
or OR2 (N11180, N11175, N8900);
nand NAND4 (N11181, N11133, N3213, N2726, N2535);
not NOT1 (N11182, N11163);
or OR3 (N11183, N11179, N1084, N209);
not NOT1 (N11184, N11177);
or OR3 (N11185, N11180, N4662, N9768);
buf BUF1 (N11186, N11185);
nand NAND2 (N11187, N11159, N11030);
nand NAND3 (N11188, N11183, N3104, N8171);
nand NAND2 (N11189, N11176, N1776);
nand NAND2 (N11190, N11171, N7544);
nor NOR2 (N11191, N11186, N9831);
nand NAND2 (N11192, N11188, N7587);
not NOT1 (N11193, N11174);
nand NAND4 (N11194, N11190, N4980, N3659, N2776);
nand NAND3 (N11195, N11184, N408, N4124);
and AND4 (N11196, N11187, N2830, N6212, N1251);
xor XOR2 (N11197, N11192, N10706);
buf BUF1 (N11198, N11181);
nor NOR3 (N11199, N11195, N4773, N2189);
not NOT1 (N11200, N11182);
xor XOR2 (N11201, N11194, N9028);
xor XOR2 (N11202, N11199, N1492);
or OR4 (N11203, N11198, N1764, N4568, N5783);
buf BUF1 (N11204, N11202);
or OR2 (N11205, N11193, N9128);
xor XOR2 (N11206, N11191, N10811);
nor NOR2 (N11207, N11205, N7735);
nand NAND4 (N11208, N11206, N9806, N3408, N8264);
buf BUF1 (N11209, N11207);
and AND4 (N11210, N11197, N2781, N8437, N9181);
xor XOR2 (N11211, N11209, N9625);
or OR4 (N11212, N11200, N6491, N5188, N9459);
xor XOR2 (N11213, N11210, N1651);
nand NAND4 (N11214, N11201, N1437, N6280, N4694);
xor XOR2 (N11215, N11167, N1670);
xor XOR2 (N11216, N11212, N956);
xor XOR2 (N11217, N11216, N1655);
nand NAND4 (N11218, N11203, N931, N6411, N9448);
or OR4 (N11219, N11214, N4998, N3613, N789);
buf BUF1 (N11220, N11215);
and AND4 (N11221, N11219, N615, N1421, N2889);
not NOT1 (N11222, N11213);
not NOT1 (N11223, N11220);
nor NOR2 (N11224, N11222, N8962);
or OR4 (N11225, N11211, N7696, N10780, N2359);
not NOT1 (N11226, N11221);
nor NOR3 (N11227, N11196, N2824, N8296);
xor XOR2 (N11228, N11217, N5699);
nand NAND4 (N11229, N11208, N3618, N2899, N6676);
buf BUF1 (N11230, N11226);
nand NAND4 (N11231, N11227, N5436, N5517, N2299);
and AND3 (N11232, N11231, N7714, N3043);
or OR2 (N11233, N11223, N3551);
xor XOR2 (N11234, N11230, N6173);
nand NAND2 (N11235, N11218, N5104);
nor NOR2 (N11236, N11233, N10070);
not NOT1 (N11237, N11234);
xor XOR2 (N11238, N11237, N6125);
nand NAND3 (N11239, N11235, N7876, N584);
nand NAND4 (N11240, N11224, N3806, N7718, N3805);
not NOT1 (N11241, N11229);
and AND2 (N11242, N11228, N7633);
buf BUF1 (N11243, N11189);
nand NAND2 (N11244, N11236, N4505);
xor XOR2 (N11245, N11243, N6883);
xor XOR2 (N11246, N11238, N1028);
buf BUF1 (N11247, N11246);
or OR2 (N11248, N11242, N7401);
nor NOR4 (N11249, N11248, N731, N1288, N5340);
xor XOR2 (N11250, N11225, N703);
or OR2 (N11251, N11239, N11238);
nor NOR2 (N11252, N11251, N4136);
nand NAND2 (N11253, N11204, N7115);
not NOT1 (N11254, N11249);
or OR3 (N11255, N11247, N2308, N3363);
xor XOR2 (N11256, N11240, N11034);
not NOT1 (N11257, N11254);
not NOT1 (N11258, N11257);
not NOT1 (N11259, N11252);
buf BUF1 (N11260, N11250);
buf BUF1 (N11261, N11244);
nor NOR4 (N11262, N11261, N7399, N4679, N10148);
and AND3 (N11263, N11260, N3492, N9467);
buf BUF1 (N11264, N11232);
not NOT1 (N11265, N11259);
nand NAND4 (N11266, N11264, N3149, N3536, N4808);
nor NOR3 (N11267, N11258, N4324, N3486);
or OR2 (N11268, N11266, N2177);
not NOT1 (N11269, N11245);
not NOT1 (N11270, N11256);
or OR4 (N11271, N11255, N393, N711, N4049);
not NOT1 (N11272, N11241);
buf BUF1 (N11273, N11271);
buf BUF1 (N11274, N11273);
buf BUF1 (N11275, N11262);
not NOT1 (N11276, N11265);
or OR4 (N11277, N11263, N1231, N9544, N10503);
not NOT1 (N11278, N11276);
xor XOR2 (N11279, N11270, N7831);
or OR3 (N11280, N11269, N5420, N10201);
nor NOR4 (N11281, N11278, N805, N10309, N6739);
buf BUF1 (N11282, N11279);
xor XOR2 (N11283, N11277, N9143);
xor XOR2 (N11284, N11253, N10820);
nand NAND3 (N11285, N11282, N9262, N2357);
or OR2 (N11286, N11274, N2335);
not NOT1 (N11287, N11280);
not NOT1 (N11288, N11283);
xor XOR2 (N11289, N11281, N7292);
buf BUF1 (N11290, N11286);
buf BUF1 (N11291, N11287);
not NOT1 (N11292, N11288);
nand NAND4 (N11293, N11290, N5350, N1626, N2297);
or OR2 (N11294, N11267, N6918);
xor XOR2 (N11295, N11291, N6079);
buf BUF1 (N11296, N11275);
and AND4 (N11297, N11284, N9394, N1589, N10303);
nor NOR4 (N11298, N11293, N4283, N10474, N8017);
xor XOR2 (N11299, N11297, N10100);
nor NOR4 (N11300, N11292, N10077, N5642, N7539);
nand NAND4 (N11301, N11295, N11013, N9416, N9415);
nand NAND4 (N11302, N11285, N100, N906, N9695);
or OR4 (N11303, N11302, N1438, N9896, N7484);
nor NOR3 (N11304, N11298, N3578, N11216);
buf BUF1 (N11305, N11299);
buf BUF1 (N11306, N11301);
nand NAND3 (N11307, N11306, N9640, N6942);
and AND3 (N11308, N11307, N8658, N2893);
and AND4 (N11309, N11308, N3012, N1844, N6146);
nor NOR2 (N11310, N11272, N4276);
not NOT1 (N11311, N11289);
xor XOR2 (N11312, N11309, N2295);
buf BUF1 (N11313, N11300);
nor NOR2 (N11314, N11305, N3433);
xor XOR2 (N11315, N11304, N3220);
nor NOR3 (N11316, N11303, N1847, N7787);
xor XOR2 (N11317, N11312, N7569);
xor XOR2 (N11318, N11268, N858);
xor XOR2 (N11319, N11315, N3525);
xor XOR2 (N11320, N11296, N1665);
xor XOR2 (N11321, N11314, N6851);
xor XOR2 (N11322, N11311, N9337);
not NOT1 (N11323, N11294);
or OR2 (N11324, N11319, N4895);
not NOT1 (N11325, N11324);
or OR3 (N11326, N11325, N9201, N5770);
nor NOR4 (N11327, N11310, N490, N2725, N8201);
xor XOR2 (N11328, N11321, N6740);
buf BUF1 (N11329, N11313);
buf BUF1 (N11330, N11327);
or OR2 (N11331, N11326, N1625);
nand NAND2 (N11332, N11320, N1367);
nor NOR2 (N11333, N11328, N7363);
buf BUF1 (N11334, N11323);
buf BUF1 (N11335, N11331);
buf BUF1 (N11336, N11322);
nand NAND2 (N11337, N11332, N5493);
or OR3 (N11338, N11318, N1365, N10551);
and AND2 (N11339, N11330, N8808);
nor NOR3 (N11340, N11336, N142, N9827);
not NOT1 (N11341, N11316);
nand NAND2 (N11342, N11339, N8427);
not NOT1 (N11343, N11317);
nor NOR2 (N11344, N11333, N1236);
or OR2 (N11345, N11329, N3658);
not NOT1 (N11346, N11342);
and AND2 (N11347, N11344, N6485);
nor NOR2 (N11348, N11346, N9749);
not NOT1 (N11349, N11348);
nand NAND3 (N11350, N11341, N5603, N227);
or OR3 (N11351, N11335, N7553, N9205);
xor XOR2 (N11352, N11349, N1164);
and AND2 (N11353, N11350, N10847);
nor NOR4 (N11354, N11352, N6515, N5084, N10403);
nor NOR3 (N11355, N11351, N9665, N1237);
buf BUF1 (N11356, N11338);
or OR3 (N11357, N11355, N3999, N5326);
or OR2 (N11358, N11343, N11313);
not NOT1 (N11359, N11354);
or OR4 (N11360, N11334, N9857, N207, N5528);
nor NOR3 (N11361, N11359, N9881, N5328);
nor NOR2 (N11362, N11337, N2717);
and AND3 (N11363, N11353, N1087, N8208);
not NOT1 (N11364, N11340);
and AND2 (N11365, N11356, N9103);
nor NOR3 (N11366, N11364, N10328, N7032);
nor NOR3 (N11367, N11362, N8750, N9696);
nor NOR2 (N11368, N11365, N10211);
nand NAND4 (N11369, N11366, N9229, N7896, N240);
xor XOR2 (N11370, N11347, N3184);
nand NAND3 (N11371, N11363, N1015, N4001);
xor XOR2 (N11372, N11345, N5693);
xor XOR2 (N11373, N11360, N9305);
nor NOR4 (N11374, N11370, N7469, N2700, N914);
and AND2 (N11375, N11361, N2820);
xor XOR2 (N11376, N11367, N6282);
buf BUF1 (N11377, N11374);
nand NAND3 (N11378, N11373, N2692, N6845);
not NOT1 (N11379, N11378);
xor XOR2 (N11380, N11376, N1703);
nand NAND4 (N11381, N11375, N3320, N9679, N1534);
xor XOR2 (N11382, N11377, N10342);
nand NAND2 (N11383, N11358, N2513);
and AND4 (N11384, N11380, N4193, N2662, N2673);
xor XOR2 (N11385, N11371, N8463);
or OR3 (N11386, N11385, N7618, N1685);
buf BUF1 (N11387, N11379);
not NOT1 (N11388, N11387);
buf BUF1 (N11389, N11384);
buf BUF1 (N11390, N11368);
and AND2 (N11391, N11388, N3195);
and AND2 (N11392, N11382, N11188);
or OR4 (N11393, N11390, N9135, N7537, N1178);
not NOT1 (N11394, N11357);
nand NAND2 (N11395, N11372, N9718);
nand NAND2 (N11396, N11395, N1221);
nor NOR3 (N11397, N11383, N9858, N2534);
xor XOR2 (N11398, N11396, N9889);
nand NAND2 (N11399, N11389, N9081);
buf BUF1 (N11400, N11398);
nor NOR2 (N11401, N11391, N9947);
buf BUF1 (N11402, N11394);
nor NOR4 (N11403, N11402, N3325, N9065, N10295);
or OR3 (N11404, N11393, N6707, N4579);
and AND4 (N11405, N11386, N6598, N3559, N7953);
or OR3 (N11406, N11392, N2259, N544);
xor XOR2 (N11407, N11381, N8431);
buf BUF1 (N11408, N11401);
xor XOR2 (N11409, N11369, N9859);
not NOT1 (N11410, N11397);
nand NAND3 (N11411, N11405, N437, N5560);
nor NOR2 (N11412, N11400, N1825);
nand NAND4 (N11413, N11404, N7012, N6783, N7953);
buf BUF1 (N11414, N11412);
not NOT1 (N11415, N11410);
xor XOR2 (N11416, N11411, N7366);
xor XOR2 (N11417, N11415, N6511);
nor NOR2 (N11418, N11417, N2172);
or OR3 (N11419, N11416, N5796, N4729);
nor NOR2 (N11420, N11408, N3806);
not NOT1 (N11421, N11419);
or OR4 (N11422, N11421, N6480, N1755, N6033);
buf BUF1 (N11423, N11407);
buf BUF1 (N11424, N11418);
and AND2 (N11425, N11403, N7962);
nand NAND4 (N11426, N11413, N6540, N4766, N2542);
and AND4 (N11427, N11424, N10390, N4651, N1733);
xor XOR2 (N11428, N11427, N10757);
buf BUF1 (N11429, N11428);
nor NOR3 (N11430, N11409, N3586, N8702);
buf BUF1 (N11431, N11422);
and AND4 (N11432, N11429, N7857, N5100, N565);
nand NAND3 (N11433, N11420, N5074, N6591);
and AND3 (N11434, N11433, N395, N8673);
not NOT1 (N11435, N11431);
not NOT1 (N11436, N11425);
buf BUF1 (N11437, N11436);
or OR3 (N11438, N11414, N6123, N2579);
buf BUF1 (N11439, N11437);
not NOT1 (N11440, N11423);
nor NOR4 (N11441, N11399, N7305, N976, N3465);
xor XOR2 (N11442, N11434, N6958);
and AND4 (N11443, N11432, N10294, N7225, N10411);
not NOT1 (N11444, N11443);
or OR2 (N11445, N11440, N7500);
buf BUF1 (N11446, N11426);
nor NOR3 (N11447, N11438, N1906, N1255);
not NOT1 (N11448, N11447);
buf BUF1 (N11449, N11445);
nor NOR4 (N11450, N11448, N10906, N7331, N11006);
not NOT1 (N11451, N11430);
not NOT1 (N11452, N11439);
and AND2 (N11453, N11435, N9954);
nand NAND2 (N11454, N11452, N386);
and AND4 (N11455, N11442, N8102, N1076, N10907);
not NOT1 (N11456, N11441);
xor XOR2 (N11457, N11444, N7292);
or OR3 (N11458, N11454, N9690, N1959);
nor NOR2 (N11459, N11453, N2241);
or OR2 (N11460, N11451, N306);
or OR3 (N11461, N11406, N2579, N9904);
nand NAND2 (N11462, N11456, N3732);
and AND2 (N11463, N11461, N10583);
buf BUF1 (N11464, N11455);
nor NOR4 (N11465, N11463, N10617, N4092, N1596);
and AND2 (N11466, N11462, N4228);
and AND2 (N11467, N11458, N2005);
xor XOR2 (N11468, N11449, N2414);
nor NOR4 (N11469, N11457, N2618, N331, N3977);
nand NAND4 (N11470, N11467, N8726, N5302, N8102);
buf BUF1 (N11471, N11450);
or OR2 (N11472, N11464, N7119);
nand NAND4 (N11473, N11470, N1796, N908, N7332);
nand NAND2 (N11474, N11446, N10482);
nor NOR4 (N11475, N11460, N134, N8100, N6680);
or OR3 (N11476, N11469, N9361, N7456);
buf BUF1 (N11477, N11468);
not NOT1 (N11478, N11473);
or OR3 (N11479, N11476, N4001, N672);
buf BUF1 (N11480, N11472);
nand NAND4 (N11481, N11478, N7740, N383, N4951);
xor XOR2 (N11482, N11481, N6008);
and AND4 (N11483, N11479, N9957, N11185, N4739);
not NOT1 (N11484, N11471);
buf BUF1 (N11485, N11483);
and AND4 (N11486, N11480, N1505, N4108, N6825);
or OR4 (N11487, N11485, N8820, N5596, N9880);
nor NOR2 (N11488, N11486, N1368);
xor XOR2 (N11489, N11466, N5441);
and AND3 (N11490, N11477, N2279, N9707);
nor NOR4 (N11491, N11474, N10746, N10607, N2555);
not NOT1 (N11492, N11488);
nor NOR2 (N11493, N11490, N7000);
nor NOR4 (N11494, N11492, N7579, N7706, N6556);
nand NAND3 (N11495, N11491, N3850, N2195);
not NOT1 (N11496, N11475);
nand NAND4 (N11497, N11496, N655, N10793, N1527);
and AND2 (N11498, N11459, N7532);
nand NAND3 (N11499, N11498, N435, N8491);
xor XOR2 (N11500, N11493, N6127);
or OR4 (N11501, N11494, N3179, N7878, N3857);
nand NAND2 (N11502, N11465, N112);
nor NOR2 (N11503, N11487, N6735);
xor XOR2 (N11504, N11489, N5084);
not NOT1 (N11505, N11482);
xor XOR2 (N11506, N11497, N8495);
nor NOR3 (N11507, N11500, N6051, N2575);
nor NOR3 (N11508, N11507, N6334, N8691);
nand NAND2 (N11509, N11501, N10814);
or OR3 (N11510, N11502, N595, N809);
or OR2 (N11511, N11508, N1549);
nor NOR3 (N11512, N11484, N2407, N1545);
buf BUF1 (N11513, N11503);
or OR4 (N11514, N11513, N7705, N8564, N10760);
buf BUF1 (N11515, N11504);
nor NOR3 (N11516, N11514, N10830, N3852);
buf BUF1 (N11517, N11505);
nand NAND2 (N11518, N11512, N4164);
not NOT1 (N11519, N11509);
nand NAND4 (N11520, N11517, N7172, N4166, N2869);
or OR4 (N11521, N11499, N2973, N6050, N1223);
nor NOR2 (N11522, N11520, N5994);
and AND4 (N11523, N11521, N4099, N10784, N889);
nand NAND4 (N11524, N11515, N8250, N4978, N8776);
xor XOR2 (N11525, N11519, N5409);
xor XOR2 (N11526, N11516, N4091);
nor NOR2 (N11527, N11524, N6571);
and AND2 (N11528, N11522, N1729);
or OR2 (N11529, N11526, N2013);
buf BUF1 (N11530, N11529);
not NOT1 (N11531, N11527);
nand NAND3 (N11532, N11511, N2843, N3849);
not NOT1 (N11533, N11530);
nand NAND2 (N11534, N11518, N1939);
nor NOR2 (N11535, N11531, N5403);
buf BUF1 (N11536, N11510);
and AND2 (N11537, N11532, N3206);
nor NOR4 (N11538, N11495, N469, N10358, N11042);
nand NAND2 (N11539, N11535, N10725);
buf BUF1 (N11540, N11528);
or OR3 (N11541, N11523, N10754, N4042);
and AND4 (N11542, N11534, N9616, N7641, N10222);
buf BUF1 (N11543, N11539);
buf BUF1 (N11544, N11543);
xor XOR2 (N11545, N11541, N5332);
and AND2 (N11546, N11540, N9438);
nand NAND4 (N11547, N11537, N4298, N7232, N8305);
buf BUF1 (N11548, N11536);
nand NAND2 (N11549, N11545, N8921);
xor XOR2 (N11550, N11549, N10432);
nor NOR4 (N11551, N11548, N11088, N3710, N1537);
nand NAND4 (N11552, N11506, N1031, N682, N5197);
or OR3 (N11553, N11547, N4153, N1980);
or OR3 (N11554, N11546, N11304, N3680);
not NOT1 (N11555, N11554);
xor XOR2 (N11556, N11553, N5490);
or OR4 (N11557, N11533, N2897, N8644, N8483);
or OR3 (N11558, N11538, N10453, N9120);
not NOT1 (N11559, N11550);
xor XOR2 (N11560, N11544, N2402);
or OR2 (N11561, N11551, N3877);
nand NAND2 (N11562, N11558, N6364);
nand NAND4 (N11563, N11542, N2700, N3939, N7789);
nor NOR4 (N11564, N11556, N729, N7940, N1138);
not NOT1 (N11565, N11557);
or OR2 (N11566, N11525, N5721);
nand NAND2 (N11567, N11564, N6195);
and AND2 (N11568, N11555, N6283);
nor NOR2 (N11569, N11559, N5100);
xor XOR2 (N11570, N11568, N6836);
and AND4 (N11571, N11552, N8369, N1071, N1892);
or OR3 (N11572, N11569, N4219, N5306);
xor XOR2 (N11573, N11571, N10045);
buf BUF1 (N11574, N11562);
xor XOR2 (N11575, N11570, N8604);
not NOT1 (N11576, N11574);
buf BUF1 (N11577, N11576);
nand NAND3 (N11578, N11567, N2443, N7854);
not NOT1 (N11579, N11573);
nor NOR2 (N11580, N11563, N773);
nor NOR3 (N11581, N11579, N4623, N3734);
or OR2 (N11582, N11566, N9789);
buf BUF1 (N11583, N11565);
or OR2 (N11584, N11578, N6016);
buf BUF1 (N11585, N11560);
buf BUF1 (N11586, N11580);
and AND4 (N11587, N11585, N3031, N9198, N3615);
or OR4 (N11588, N11581, N1998, N7125, N2981);
buf BUF1 (N11589, N11588);
nor NOR2 (N11590, N11561, N7541);
and AND4 (N11591, N11582, N20, N5091, N2968);
not NOT1 (N11592, N11586);
nor NOR4 (N11593, N11577, N3247, N5634, N10395);
or OR3 (N11594, N11589, N8445, N2981);
nand NAND3 (N11595, N11590, N10164, N3966);
nor NOR3 (N11596, N11583, N5901, N10407);
nor NOR3 (N11597, N11593, N9868, N6920);
nand NAND4 (N11598, N11572, N3566, N1115, N6946);
xor XOR2 (N11599, N11591, N4077);
nor NOR2 (N11600, N11594, N8770);
buf BUF1 (N11601, N11592);
and AND4 (N11602, N11598, N10803, N29, N2973);
buf BUF1 (N11603, N11596);
xor XOR2 (N11604, N11602, N3232);
nand NAND3 (N11605, N11595, N1237, N8205);
buf BUF1 (N11606, N11587);
or OR4 (N11607, N11603, N3501, N9619, N7964);
nor NOR3 (N11608, N11606, N242, N9016);
nand NAND3 (N11609, N11584, N2100, N11234);
xor XOR2 (N11610, N11600, N8269);
and AND3 (N11611, N11604, N5201, N11479);
and AND3 (N11612, N11605, N8767, N499);
nor NOR3 (N11613, N11607, N4188, N3702);
xor XOR2 (N11614, N11613, N7760);
xor XOR2 (N11615, N11612, N3871);
not NOT1 (N11616, N11611);
buf BUF1 (N11617, N11599);
nor NOR2 (N11618, N11608, N7728);
nand NAND4 (N11619, N11618, N3866, N9588, N2676);
xor XOR2 (N11620, N11614, N6766);
nor NOR2 (N11621, N11617, N3536);
buf BUF1 (N11622, N11619);
not NOT1 (N11623, N11615);
xor XOR2 (N11624, N11622, N1570);
nor NOR3 (N11625, N11616, N10717, N9628);
and AND2 (N11626, N11625, N3283);
not NOT1 (N11627, N11610);
nor NOR4 (N11628, N11575, N57, N7692, N7068);
nor NOR4 (N11629, N11620, N7751, N7858, N1792);
xor XOR2 (N11630, N11629, N4249);
buf BUF1 (N11631, N11628);
and AND2 (N11632, N11621, N10971);
nand NAND3 (N11633, N11623, N6116, N8888);
and AND4 (N11634, N11627, N8294, N3754, N7649);
nor NOR2 (N11635, N11624, N9271);
nor NOR3 (N11636, N11630, N7883, N1552);
buf BUF1 (N11637, N11609);
nand NAND4 (N11638, N11597, N7980, N5291, N4513);
nor NOR3 (N11639, N11632, N10575, N5975);
xor XOR2 (N11640, N11636, N934);
or OR4 (N11641, N11640, N7760, N6712, N9612);
nor NOR2 (N11642, N11635, N3995);
or OR4 (N11643, N11641, N814, N1204, N10353);
nor NOR3 (N11644, N11601, N5635, N7117);
or OR3 (N11645, N11631, N9379, N6581);
nor NOR4 (N11646, N11633, N9269, N3661, N2065);
nand NAND3 (N11647, N11645, N11164, N6065);
not NOT1 (N11648, N11626);
xor XOR2 (N11649, N11637, N1483);
not NOT1 (N11650, N11639);
nor NOR2 (N11651, N11648, N5948);
nand NAND2 (N11652, N11647, N9937);
nor NOR4 (N11653, N11634, N1612, N4781, N5911);
nor NOR2 (N11654, N11644, N3490);
and AND2 (N11655, N11649, N9834);
buf BUF1 (N11656, N11646);
and AND4 (N11657, N11650, N3446, N9094, N1907);
not NOT1 (N11658, N11653);
and AND4 (N11659, N11658, N7753, N9949, N826);
or OR4 (N11660, N11638, N9272, N2200, N598);
not NOT1 (N11661, N11652);
not NOT1 (N11662, N11661);
nor NOR2 (N11663, N11654, N10792);
nand NAND4 (N11664, N11663, N2899, N7421, N3116);
not NOT1 (N11665, N11642);
xor XOR2 (N11666, N11651, N6879);
and AND4 (N11667, N11655, N328, N408, N4649);
nand NAND4 (N11668, N11643, N6993, N6320, N4280);
buf BUF1 (N11669, N11659);
or OR3 (N11670, N11660, N7946, N9090);
nor NOR4 (N11671, N11665, N5816, N9834, N7448);
nand NAND3 (N11672, N11666, N3533, N10095);
not NOT1 (N11673, N11664);
nor NOR3 (N11674, N11668, N969, N4186);
not NOT1 (N11675, N11674);
and AND4 (N11676, N11670, N6210, N10112, N2761);
not NOT1 (N11677, N11656);
or OR4 (N11678, N11677, N11672, N8343, N2568);
nand NAND2 (N11679, N2446, N3823);
nor NOR4 (N11680, N11678, N7101, N10498, N6358);
or OR4 (N11681, N11676, N10440, N3349, N8817);
not NOT1 (N11682, N11673);
buf BUF1 (N11683, N11681);
nand NAND3 (N11684, N11657, N3880, N11232);
or OR4 (N11685, N11679, N6600, N7859, N7228);
and AND2 (N11686, N11680, N10723);
buf BUF1 (N11687, N11682);
and AND4 (N11688, N11675, N8234, N3079, N3106);
buf BUF1 (N11689, N11685);
nor NOR3 (N11690, N11671, N6018, N10344);
nand NAND2 (N11691, N11669, N452);
xor XOR2 (N11692, N11688, N2915);
buf BUF1 (N11693, N11690);
not NOT1 (N11694, N11687);
or OR2 (N11695, N11683, N4395);
nand NAND3 (N11696, N11684, N2066, N1906);
nand NAND4 (N11697, N11689, N2475, N626, N9733);
buf BUF1 (N11698, N11696);
not NOT1 (N11699, N11691);
buf BUF1 (N11700, N11692);
or OR3 (N11701, N11686, N2491, N7383);
xor XOR2 (N11702, N11667, N5288);
nor NOR3 (N11703, N11695, N7444, N6765);
buf BUF1 (N11704, N11703);
buf BUF1 (N11705, N11701);
or OR2 (N11706, N11697, N9569);
nor NOR3 (N11707, N11706, N7083, N570);
nand NAND3 (N11708, N11662, N5328, N1818);
not NOT1 (N11709, N11707);
not NOT1 (N11710, N11709);
nor NOR4 (N11711, N11698, N11193, N10470, N11168);
not NOT1 (N11712, N11693);
xor XOR2 (N11713, N11702, N2674);
or OR3 (N11714, N11708, N6651, N6891);
not NOT1 (N11715, N11694);
buf BUF1 (N11716, N11710);
and AND2 (N11717, N11711, N9079);
or OR3 (N11718, N11714, N2020, N11108);
nand NAND2 (N11719, N11717, N3839);
and AND4 (N11720, N11719, N8670, N2543, N11699);
and AND4 (N11721, N1941, N6833, N8749, N5028);
or OR2 (N11722, N11713, N1333);
or OR4 (N11723, N11712, N9805, N9436, N9421);
not NOT1 (N11724, N11718);
not NOT1 (N11725, N11705);
nand NAND3 (N11726, N11722, N4309, N9122);
not NOT1 (N11727, N11723);
and AND3 (N11728, N11704, N11349, N11017);
xor XOR2 (N11729, N11727, N8113);
xor XOR2 (N11730, N11715, N2973);
or OR2 (N11731, N11726, N8588);
nand NAND4 (N11732, N11720, N2131, N3519, N1883);
not NOT1 (N11733, N11700);
and AND4 (N11734, N11721, N459, N5728, N4361);
and AND4 (N11735, N11734, N268, N6755, N11182);
not NOT1 (N11736, N11731);
and AND4 (N11737, N11730, N11000, N4673, N9824);
buf BUF1 (N11738, N11737);
nand NAND3 (N11739, N11732, N6378, N9280);
not NOT1 (N11740, N11725);
and AND3 (N11741, N11740, N8793, N8575);
not NOT1 (N11742, N11733);
nor NOR2 (N11743, N11728, N818);
buf BUF1 (N11744, N11738);
and AND2 (N11745, N11735, N5165);
and AND2 (N11746, N11724, N7777);
xor XOR2 (N11747, N11739, N3524);
nand NAND4 (N11748, N11741, N11192, N47, N377);
nand NAND4 (N11749, N11745, N10805, N6357, N7883);
xor XOR2 (N11750, N11746, N7922);
not NOT1 (N11751, N11743);
nand NAND4 (N11752, N11716, N3022, N10347, N8479);
not NOT1 (N11753, N11736);
nor NOR3 (N11754, N11753, N2254, N670);
buf BUF1 (N11755, N11747);
and AND3 (N11756, N11752, N1501, N10387);
xor XOR2 (N11757, N11755, N5781);
buf BUF1 (N11758, N11744);
nand NAND2 (N11759, N11751, N10470);
buf BUF1 (N11760, N11729);
or OR2 (N11761, N11758, N1587);
not NOT1 (N11762, N11757);
nor NOR4 (N11763, N11748, N8682, N10563, N1102);
and AND4 (N11764, N11763, N9518, N5433, N11625);
nor NOR2 (N11765, N11762, N3125);
and AND2 (N11766, N11756, N1560);
not NOT1 (N11767, N11754);
not NOT1 (N11768, N11750);
or OR4 (N11769, N11766, N6566, N6181, N1915);
nand NAND3 (N11770, N11761, N6209, N11165);
and AND4 (N11771, N11742, N4265, N3553, N8371);
nor NOR3 (N11772, N11764, N5639, N6644);
not NOT1 (N11773, N11768);
xor XOR2 (N11774, N11765, N5919);
or OR2 (N11775, N11772, N9942);
and AND3 (N11776, N11769, N3492, N10943);
nor NOR4 (N11777, N11774, N1945, N872, N9132);
or OR3 (N11778, N11749, N4279, N11471);
or OR4 (N11779, N11773, N11301, N7969, N10093);
and AND3 (N11780, N11779, N193, N7888);
buf BUF1 (N11781, N11760);
nor NOR2 (N11782, N11770, N3555);
or OR2 (N11783, N11759, N7440);
and AND2 (N11784, N11767, N9683);
or OR4 (N11785, N11776, N11484, N2781, N3208);
nor NOR4 (N11786, N11771, N7334, N6611, N11230);
not NOT1 (N11787, N11780);
nand NAND2 (N11788, N11778, N2838);
and AND4 (N11789, N11785, N9239, N6106, N2745);
nand NAND3 (N11790, N11781, N8703, N10281);
xor XOR2 (N11791, N11786, N149);
buf BUF1 (N11792, N11782);
buf BUF1 (N11793, N11775);
xor XOR2 (N11794, N11790, N2998);
or OR4 (N11795, N11777, N4251, N11355, N2690);
buf BUF1 (N11796, N11792);
or OR3 (N11797, N11783, N7248, N4415);
and AND2 (N11798, N11784, N6563);
and AND4 (N11799, N11787, N1436, N368, N4607);
nand NAND2 (N11800, N11799, N6977);
xor XOR2 (N11801, N11794, N7136);
and AND3 (N11802, N11791, N11137, N10066);
buf BUF1 (N11803, N11798);
buf BUF1 (N11804, N11796);
and AND2 (N11805, N11801, N10751);
or OR3 (N11806, N11795, N3357, N8342);
or OR2 (N11807, N11793, N3390);
xor XOR2 (N11808, N11788, N434);
not NOT1 (N11809, N11808);
xor XOR2 (N11810, N11806, N668);
or OR3 (N11811, N11804, N3248, N4170);
nand NAND4 (N11812, N11805, N2033, N3872, N9889);
and AND2 (N11813, N11811, N1879);
xor XOR2 (N11814, N11797, N1388);
xor XOR2 (N11815, N11800, N1636);
buf BUF1 (N11816, N11812);
nor NOR2 (N11817, N11816, N9362);
xor XOR2 (N11818, N11807, N6589);
nand NAND3 (N11819, N11810, N5931, N9831);
nor NOR3 (N11820, N11789, N9413, N6277);
buf BUF1 (N11821, N11809);
nand NAND3 (N11822, N11803, N2552, N10181);
nand NAND3 (N11823, N11814, N5928, N887);
or OR2 (N11824, N11823, N5857);
not NOT1 (N11825, N11813);
nor NOR4 (N11826, N11821, N11702, N6576, N492);
buf BUF1 (N11827, N11817);
buf BUF1 (N11828, N11818);
buf BUF1 (N11829, N11824);
or OR4 (N11830, N11828, N8387, N1313, N1049);
nor NOR3 (N11831, N11819, N6839, N6544);
buf BUF1 (N11832, N11822);
buf BUF1 (N11833, N11829);
xor XOR2 (N11834, N11827, N4662);
or OR2 (N11835, N11831, N3500);
buf BUF1 (N11836, N11820);
not NOT1 (N11837, N11830);
or OR2 (N11838, N11825, N1811);
xor XOR2 (N11839, N11833, N5115);
not NOT1 (N11840, N11802);
xor XOR2 (N11841, N11840, N5633);
or OR3 (N11842, N11815, N553, N8514);
not NOT1 (N11843, N11839);
and AND2 (N11844, N11842, N5024);
nand NAND2 (N11845, N11826, N8239);
not NOT1 (N11846, N11837);
nor NOR2 (N11847, N11844, N9699);
buf BUF1 (N11848, N11841);
xor XOR2 (N11849, N11832, N9577);
nor NOR3 (N11850, N11843, N1004, N10692);
or OR2 (N11851, N11835, N5658);
buf BUF1 (N11852, N11834);
not NOT1 (N11853, N11849);
nor NOR3 (N11854, N11848, N11388, N2375);
or OR2 (N11855, N11847, N9362);
nand NAND2 (N11856, N11851, N5009);
or OR2 (N11857, N11838, N391);
or OR4 (N11858, N11853, N6159, N7325, N4851);
buf BUF1 (N11859, N11858);
nor NOR4 (N11860, N11854, N10496, N5288, N4291);
buf BUF1 (N11861, N11846);
or OR4 (N11862, N11856, N3518, N521, N4114);
xor XOR2 (N11863, N11862, N10522);
nand NAND4 (N11864, N11861, N10870, N11557, N7021);
nand NAND3 (N11865, N11855, N1871, N8977);
nand NAND4 (N11866, N11852, N8931, N10566, N3929);
or OR2 (N11867, N11850, N3995);
and AND2 (N11868, N11867, N523);
and AND4 (N11869, N11836, N5992, N897, N9442);
buf BUF1 (N11870, N11869);
xor XOR2 (N11871, N11868, N46);
not NOT1 (N11872, N11863);
or OR4 (N11873, N11864, N11053, N1866, N1781);
and AND2 (N11874, N11866, N10975);
nand NAND3 (N11875, N11865, N5746, N773);
xor XOR2 (N11876, N11860, N10827);
not NOT1 (N11877, N11859);
xor XOR2 (N11878, N11874, N8558);
nand NAND2 (N11879, N11875, N10318);
nor NOR4 (N11880, N11870, N1142, N5308, N7498);
not NOT1 (N11881, N11871);
or OR4 (N11882, N11880, N10121, N1631, N4989);
nor NOR3 (N11883, N11878, N9355, N5437);
not NOT1 (N11884, N11883);
nand NAND3 (N11885, N11857, N2963, N1473);
not NOT1 (N11886, N11876);
or OR2 (N11887, N11845, N5341);
xor XOR2 (N11888, N11877, N10749);
not NOT1 (N11889, N11881);
xor XOR2 (N11890, N11879, N11572);
and AND2 (N11891, N11873, N11272);
or OR2 (N11892, N11891, N4504);
xor XOR2 (N11893, N11872, N9865);
buf BUF1 (N11894, N11885);
and AND3 (N11895, N11889, N5202, N7582);
buf BUF1 (N11896, N11894);
or OR3 (N11897, N11888, N2031, N7012);
or OR3 (N11898, N11887, N11657, N3291);
nor NOR2 (N11899, N11896, N2566);
not NOT1 (N11900, N11884);
buf BUF1 (N11901, N11893);
not NOT1 (N11902, N11898);
and AND4 (N11903, N11895, N10459, N9959, N10884);
and AND2 (N11904, N11902, N2192);
nand NAND4 (N11905, N11882, N2940, N6843, N4034);
xor XOR2 (N11906, N11901, N5524);
nor NOR2 (N11907, N11905, N1116);
nor NOR4 (N11908, N11907, N1795, N8277, N9073);
nand NAND3 (N11909, N11904, N10106, N6536);
nor NOR4 (N11910, N11892, N10571, N331, N11441);
nand NAND3 (N11911, N11897, N11361, N3370);
nor NOR2 (N11912, N11890, N11197);
and AND3 (N11913, N11908, N6908, N791);
and AND2 (N11914, N11911, N63);
and AND3 (N11915, N11899, N6570, N7451);
not NOT1 (N11916, N11913);
not NOT1 (N11917, N11916);
not NOT1 (N11918, N11900);
or OR4 (N11919, N11914, N3101, N10806, N7602);
nand NAND3 (N11920, N11917, N7650, N8363);
not NOT1 (N11921, N11903);
buf BUF1 (N11922, N11920);
and AND2 (N11923, N11915, N9728);
nand NAND3 (N11924, N11922, N5571, N5654);
not NOT1 (N11925, N11923);
nand NAND3 (N11926, N11906, N8140, N5612);
xor XOR2 (N11927, N11910, N6704);
not NOT1 (N11928, N11918);
buf BUF1 (N11929, N11924);
xor XOR2 (N11930, N11919, N3730);
nor NOR4 (N11931, N11929, N10107, N504, N8811);
xor XOR2 (N11932, N11921, N11582);
or OR2 (N11933, N11912, N630);
nand NAND3 (N11934, N11933, N2854, N5287);
xor XOR2 (N11935, N11926, N7231);
or OR3 (N11936, N11935, N55, N4499);
nor NOR4 (N11937, N11930, N9015, N4104, N5575);
nor NOR4 (N11938, N11934, N8229, N2495, N10570);
and AND2 (N11939, N11909, N6229);
buf BUF1 (N11940, N11936);
or OR3 (N11941, N11886, N8697, N9486);
nand NAND4 (N11942, N11939, N8753, N264, N7431);
nor NOR4 (N11943, N11937, N3833, N9282, N11271);
xor XOR2 (N11944, N11940, N5309);
and AND4 (N11945, N11932, N4790, N7286, N4417);
buf BUF1 (N11946, N11927);
or OR4 (N11947, N11941, N2651, N1711, N10584);
and AND2 (N11948, N11943, N8264);
xor XOR2 (N11949, N11944, N11022);
buf BUF1 (N11950, N11925);
nor NOR4 (N11951, N11947, N7230, N1500, N6695);
nand NAND3 (N11952, N11938, N1883, N7125);
nor NOR2 (N11953, N11931, N6940);
not NOT1 (N11954, N11942);
nand NAND3 (N11955, N11954, N2347, N1356);
nand NAND3 (N11956, N11953, N5613, N324);
or OR2 (N11957, N11950, N10263);
nand NAND4 (N11958, N11949, N674, N4570, N968);
or OR3 (N11959, N11952, N6039, N1141);
nor NOR3 (N11960, N11951, N1719, N7011);
nor NOR3 (N11961, N11955, N6552, N1051);
xor XOR2 (N11962, N11948, N11862);
nand NAND4 (N11963, N11945, N97, N7227, N9087);
and AND2 (N11964, N11960, N10716);
nor NOR4 (N11965, N11958, N8652, N3422, N11841);
nand NAND3 (N11966, N11964, N1952, N10492);
nand NAND3 (N11967, N11962, N3575, N2160);
buf BUF1 (N11968, N11966);
nand NAND4 (N11969, N11965, N6238, N3591, N9686);
and AND3 (N11970, N11946, N251, N5571);
nand NAND3 (N11971, N11959, N9526, N4861);
or OR4 (N11972, N11961, N9611, N4729, N6351);
xor XOR2 (N11973, N11967, N484);
nand NAND3 (N11974, N11970, N1434, N1179);
nor NOR3 (N11975, N11971, N4610, N2854);
not NOT1 (N11976, N11973);
or OR3 (N11977, N11956, N10832, N3693);
nand NAND3 (N11978, N11968, N2984, N1648);
nand NAND3 (N11979, N11978, N7541, N5962);
not NOT1 (N11980, N11963);
xor XOR2 (N11981, N11969, N6267);
nand NAND4 (N11982, N11975, N843, N10953, N4520);
or OR4 (N11983, N11928, N6827, N1911, N905);
nor NOR3 (N11984, N11974, N11590, N11704);
nor NOR2 (N11985, N11982, N8508);
buf BUF1 (N11986, N11979);
nor NOR2 (N11987, N11985, N3077);
not NOT1 (N11988, N11984);
and AND4 (N11989, N11957, N8813, N11732, N10738);
buf BUF1 (N11990, N11977);
not NOT1 (N11991, N11988);
xor XOR2 (N11992, N11981, N6618);
not NOT1 (N11993, N11983);
xor XOR2 (N11994, N11972, N3509);
not NOT1 (N11995, N11993);
xor XOR2 (N11996, N11994, N8110);
nand NAND4 (N11997, N11987, N2134, N10973, N6443);
not NOT1 (N11998, N11995);
nor NOR4 (N11999, N11990, N8902, N8917, N6888);
xor XOR2 (N12000, N11989, N5891);
nand NAND2 (N12001, N11992, N2294);
xor XOR2 (N12002, N11996, N3078);
nand NAND3 (N12003, N12000, N182, N11600);
nand NAND2 (N12004, N11980, N10838);
and AND4 (N12005, N12004, N8349, N7428, N6700);
or OR3 (N12006, N11976, N10970, N4361);
nor NOR3 (N12007, N11998, N3578, N6008);
buf BUF1 (N12008, N11991);
xor XOR2 (N12009, N12001, N9549);
not NOT1 (N12010, N12009);
not NOT1 (N12011, N12003);
buf BUF1 (N12012, N12006);
or OR3 (N12013, N12008, N1422, N1224);
not NOT1 (N12014, N12012);
nor NOR4 (N12015, N12011, N6651, N491, N677);
nand NAND4 (N12016, N11997, N5507, N7973, N10441);
nand NAND3 (N12017, N12013, N2032, N10077);
and AND3 (N12018, N12010, N11492, N4487);
nor NOR3 (N12019, N12007, N9221, N8207);
not NOT1 (N12020, N12017);
buf BUF1 (N12021, N12014);
nand NAND2 (N12022, N12002, N5215);
and AND3 (N12023, N12022, N12006, N9489);
not NOT1 (N12024, N12019);
buf BUF1 (N12025, N12024);
nand NAND4 (N12026, N12023, N6853, N1939, N1081);
buf BUF1 (N12027, N12018);
buf BUF1 (N12028, N12026);
and AND4 (N12029, N11986, N1637, N10693, N6681);
nand NAND3 (N12030, N12016, N5670, N10088);
xor XOR2 (N12031, N12029, N10176);
or OR3 (N12032, N11999, N6436, N1222);
xor XOR2 (N12033, N12032, N1588);
buf BUF1 (N12034, N12025);
nand NAND4 (N12035, N12015, N9249, N1294, N1220);
and AND2 (N12036, N12033, N6247);
buf BUF1 (N12037, N12028);
not NOT1 (N12038, N12031);
and AND3 (N12039, N12035, N3549, N436);
not NOT1 (N12040, N12005);
buf BUF1 (N12041, N12034);
nor NOR3 (N12042, N12040, N10266, N11960);
nor NOR4 (N12043, N12021, N1813, N5306, N3109);
and AND3 (N12044, N12036, N2396, N3373);
or OR2 (N12045, N12039, N4173);
and AND3 (N12046, N12041, N6162, N6165);
not NOT1 (N12047, N12044);
xor XOR2 (N12048, N12027, N6173);
or OR4 (N12049, N12037, N11949, N3553, N461);
and AND4 (N12050, N12047, N3799, N9056, N1330);
or OR4 (N12051, N12038, N10729, N4750, N12038);
nand NAND4 (N12052, N12020, N9313, N9143, N9936);
buf BUF1 (N12053, N12042);
or OR2 (N12054, N12045, N2885);
or OR2 (N12055, N12053, N6567);
not NOT1 (N12056, N12052);
and AND2 (N12057, N12030, N2592);
and AND3 (N12058, N12046, N278, N10705);
not NOT1 (N12059, N12043);
xor XOR2 (N12060, N12056, N3025);
and AND3 (N12061, N12054, N4380, N2367);
and AND4 (N12062, N12059, N9856, N9055, N7890);
or OR2 (N12063, N12058, N5729);
not NOT1 (N12064, N12062);
xor XOR2 (N12065, N12050, N12004);
not NOT1 (N12066, N12051);
and AND3 (N12067, N12048, N5389, N6663);
xor XOR2 (N12068, N12055, N1569);
and AND2 (N12069, N12061, N11691);
buf BUF1 (N12070, N12060);
buf BUF1 (N12071, N12066);
nand NAND3 (N12072, N12064, N11280, N6382);
or OR3 (N12073, N12071, N9091, N10848);
xor XOR2 (N12074, N12068, N11957);
not NOT1 (N12075, N12072);
not NOT1 (N12076, N12074);
or OR3 (N12077, N12057, N7865, N9954);
nor NOR3 (N12078, N12067, N4878, N4005);
not NOT1 (N12079, N12073);
not NOT1 (N12080, N12079);
xor XOR2 (N12081, N12049, N6672);
nor NOR3 (N12082, N12075, N6132, N9068);
xor XOR2 (N12083, N12070, N7079);
nand NAND3 (N12084, N12069, N11547, N11718);
or OR2 (N12085, N12078, N8506);
nor NOR2 (N12086, N12065, N138);
not NOT1 (N12087, N12086);
not NOT1 (N12088, N12063);
nor NOR2 (N12089, N12076, N8971);
nand NAND4 (N12090, N12089, N5482, N11517, N11125);
not NOT1 (N12091, N12084);
and AND4 (N12092, N12087, N654, N7680, N5736);
xor XOR2 (N12093, N12092, N10490);
nand NAND3 (N12094, N12083, N8503, N1446);
nand NAND2 (N12095, N12093, N7393);
nor NOR4 (N12096, N12081, N10752, N10316, N900);
not NOT1 (N12097, N12088);
and AND3 (N12098, N12090, N3470, N1014);
xor XOR2 (N12099, N12097, N10002);
buf BUF1 (N12100, N12080);
not NOT1 (N12101, N12085);
xor XOR2 (N12102, N12082, N2573);
nand NAND4 (N12103, N12095, N9109, N4800, N9601);
nand NAND4 (N12104, N12096, N3687, N7941, N11257);
not NOT1 (N12105, N12102);
and AND2 (N12106, N12101, N5150);
nor NOR4 (N12107, N12091, N6825, N9389, N9952);
nand NAND3 (N12108, N12104, N3527, N8005);
nor NOR2 (N12109, N12107, N1613);
or OR2 (N12110, N12098, N3772);
xor XOR2 (N12111, N12094, N9065);
xor XOR2 (N12112, N12109, N6345);
not NOT1 (N12113, N12110);
or OR3 (N12114, N12108, N10984, N10940);
and AND2 (N12115, N12100, N6854);
or OR3 (N12116, N12105, N375, N2955);
nor NOR4 (N12117, N12113, N2548, N6555, N8809);
or OR4 (N12118, N12117, N7695, N6954, N6240);
buf BUF1 (N12119, N12106);
not NOT1 (N12120, N12118);
buf BUF1 (N12121, N12111);
not NOT1 (N12122, N12103);
xor XOR2 (N12123, N12077, N5208);
xor XOR2 (N12124, N12123, N11799);
buf BUF1 (N12125, N12124);
nand NAND3 (N12126, N12122, N1895, N5424);
nor NOR3 (N12127, N12099, N7440, N2509);
and AND4 (N12128, N12120, N2593, N5709, N2494);
xor XOR2 (N12129, N12119, N7599);
xor XOR2 (N12130, N12128, N1599);
nand NAND4 (N12131, N12126, N5192, N10397, N11200);
xor XOR2 (N12132, N12116, N9796);
buf BUF1 (N12133, N12115);
and AND2 (N12134, N12130, N12115);
and AND4 (N12135, N12129, N837, N11904, N3626);
and AND2 (N12136, N12112, N9112);
not NOT1 (N12137, N12136);
and AND4 (N12138, N12135, N6338, N8136, N7519);
buf BUF1 (N12139, N12138);
not NOT1 (N12140, N12134);
or OR4 (N12141, N12132, N11909, N2661, N4463);
or OR2 (N12142, N12127, N6451);
xor XOR2 (N12143, N12133, N2483);
not NOT1 (N12144, N12125);
xor XOR2 (N12145, N12131, N2528);
not NOT1 (N12146, N12143);
or OR3 (N12147, N12145, N7991, N6355);
or OR4 (N12148, N12140, N4597, N10432, N7723);
xor XOR2 (N12149, N12146, N5334);
or OR4 (N12150, N12141, N4560, N10789, N9942);
and AND4 (N12151, N12148, N2894, N9269, N1813);
or OR4 (N12152, N12114, N716, N1944, N3510);
and AND2 (N12153, N12149, N7614);
or OR2 (N12154, N12150, N439);
or OR3 (N12155, N12121, N3608, N1908);
and AND4 (N12156, N12154, N11075, N5049, N3422);
and AND3 (N12157, N12155, N11625, N406);
not NOT1 (N12158, N12156);
xor XOR2 (N12159, N12139, N10266);
or OR4 (N12160, N12147, N2542, N6444, N11849);
xor XOR2 (N12161, N12160, N10811);
and AND3 (N12162, N12142, N8507, N4478);
xor XOR2 (N12163, N12158, N3342);
buf BUF1 (N12164, N12152);
not NOT1 (N12165, N12162);
nor NOR3 (N12166, N12159, N2449, N9322);
buf BUF1 (N12167, N12164);
not NOT1 (N12168, N12166);
and AND2 (N12169, N12151, N11483);
xor XOR2 (N12170, N12167, N3801);
nand NAND2 (N12171, N12153, N11354);
nor NOR4 (N12172, N12171, N5251, N3623, N7588);
nor NOR2 (N12173, N12157, N3288);
xor XOR2 (N12174, N12170, N2633);
xor XOR2 (N12175, N12168, N2249);
and AND3 (N12176, N12144, N2915, N9025);
xor XOR2 (N12177, N12161, N8644);
and AND4 (N12178, N12177, N2818, N1452, N10808);
buf BUF1 (N12179, N12172);
or OR2 (N12180, N12176, N3075);
not NOT1 (N12181, N12179);
xor XOR2 (N12182, N12169, N2561);
buf BUF1 (N12183, N12181);
xor XOR2 (N12184, N12178, N10532);
and AND2 (N12185, N12183, N11316);
not NOT1 (N12186, N12173);
or OR4 (N12187, N12186, N3789, N6881, N5831);
nor NOR2 (N12188, N12182, N3542);
or OR4 (N12189, N12187, N5712, N4841, N346);
or OR2 (N12190, N12175, N3328);
buf BUF1 (N12191, N12165);
buf BUF1 (N12192, N12180);
and AND2 (N12193, N12137, N1156);
buf BUF1 (N12194, N12184);
nor NOR4 (N12195, N12163, N4951, N1464, N634);
or OR3 (N12196, N12185, N5653, N668);
xor XOR2 (N12197, N12188, N4004);
xor XOR2 (N12198, N12190, N435);
xor XOR2 (N12199, N12194, N11113);
nor NOR4 (N12200, N12199, N11020, N10856, N3955);
not NOT1 (N12201, N12198);
nand NAND2 (N12202, N12192, N7652);
not NOT1 (N12203, N12193);
xor XOR2 (N12204, N12200, N10757);
nor NOR3 (N12205, N12189, N11003, N10321);
or OR4 (N12206, N12174, N995, N2993, N11029);
xor XOR2 (N12207, N12201, N10165);
nand NAND4 (N12208, N12197, N6898, N4151, N4481);
and AND2 (N12209, N12205, N9017);
or OR2 (N12210, N12206, N5990);
or OR2 (N12211, N12191, N9816);
and AND4 (N12212, N12209, N1470, N2820, N5805);
or OR2 (N12213, N12203, N10053);
and AND2 (N12214, N12195, N8186);
nor NOR2 (N12215, N12196, N12137);
xor XOR2 (N12216, N12207, N9423);
and AND2 (N12217, N12216, N10575);
buf BUF1 (N12218, N12211);
nand NAND4 (N12219, N12202, N6498, N244, N7614);
or OR4 (N12220, N12217, N1036, N10854, N7102);
nor NOR2 (N12221, N12212, N8679);
not NOT1 (N12222, N12214);
not NOT1 (N12223, N12213);
not NOT1 (N12224, N12218);
xor XOR2 (N12225, N12221, N2127);
or OR3 (N12226, N12224, N9133, N8047);
buf BUF1 (N12227, N12223);
and AND3 (N12228, N12226, N7894, N400);
or OR2 (N12229, N12208, N5770);
and AND3 (N12230, N12204, N1248, N7158);
and AND3 (N12231, N12220, N8346, N7308);
nor NOR2 (N12232, N12227, N1499);
xor XOR2 (N12233, N12230, N4729);
nand NAND3 (N12234, N12210, N3731, N11696);
buf BUF1 (N12235, N12233);
xor XOR2 (N12236, N12225, N10657);
or OR2 (N12237, N12236, N11137);
or OR2 (N12238, N12215, N4882);
and AND3 (N12239, N12219, N6238, N11337);
nor NOR4 (N12240, N12222, N3469, N8144, N704);
not NOT1 (N12241, N12232);
xor XOR2 (N12242, N12238, N11199);
or OR2 (N12243, N12234, N4377);
not NOT1 (N12244, N12231);
or OR4 (N12245, N12229, N6470, N9305, N3590);
nor NOR3 (N12246, N12235, N7602, N3677);
not NOT1 (N12247, N12237);
buf BUF1 (N12248, N12246);
nor NOR3 (N12249, N12242, N4404, N5801);
and AND4 (N12250, N12247, N8516, N5561, N9472);
and AND3 (N12251, N12243, N9041, N498);
not NOT1 (N12252, N12249);
nor NOR4 (N12253, N12241, N7585, N7986, N3642);
xor XOR2 (N12254, N12252, N5648);
nor NOR2 (N12255, N12239, N1709);
nor NOR3 (N12256, N12250, N2715, N5642);
not NOT1 (N12257, N12228);
and AND3 (N12258, N12253, N10331, N9318);
xor XOR2 (N12259, N12254, N7331);
nor NOR4 (N12260, N12245, N4431, N5981, N9792);
and AND4 (N12261, N12244, N6736, N12206, N12163);
or OR3 (N12262, N12261, N3607, N235);
nand NAND3 (N12263, N12260, N8196, N8857);
nor NOR3 (N12264, N12263, N10818, N6966);
xor XOR2 (N12265, N12255, N4215);
buf BUF1 (N12266, N12258);
buf BUF1 (N12267, N12248);
or OR3 (N12268, N12266, N4745, N6222);
xor XOR2 (N12269, N12268, N120);
and AND2 (N12270, N12269, N9643);
and AND3 (N12271, N12240, N2208, N8392);
or OR4 (N12272, N12264, N10895, N4272, N8187);
buf BUF1 (N12273, N12271);
xor XOR2 (N12274, N12265, N5159);
or OR4 (N12275, N12267, N12130, N3034, N5706);
not NOT1 (N12276, N12259);
not NOT1 (N12277, N12276);
nor NOR3 (N12278, N12262, N8316, N8530);
buf BUF1 (N12279, N12270);
xor XOR2 (N12280, N12273, N9030);
nand NAND4 (N12281, N12275, N11884, N11530, N1854);
nor NOR3 (N12282, N12278, N2459, N4228);
nor NOR4 (N12283, N12282, N7872, N7457, N11452);
or OR4 (N12284, N12251, N990, N2457, N2809);
not NOT1 (N12285, N12280);
xor XOR2 (N12286, N12277, N5975);
xor XOR2 (N12287, N12272, N3349);
nor NOR3 (N12288, N12274, N4143, N8003);
nor NOR4 (N12289, N12288, N4225, N6034, N8293);
or OR3 (N12290, N12285, N10805, N1913);
nor NOR2 (N12291, N12287, N8610);
buf BUF1 (N12292, N12283);
buf BUF1 (N12293, N12286);
xor XOR2 (N12294, N12284, N10510);
not NOT1 (N12295, N12290);
not NOT1 (N12296, N12279);
nor NOR3 (N12297, N12257, N8867, N5477);
xor XOR2 (N12298, N12289, N5250);
or OR3 (N12299, N12256, N4236, N7267);
not NOT1 (N12300, N12295);
or OR4 (N12301, N12293, N3242, N8219, N5186);
xor XOR2 (N12302, N12300, N6517);
nor NOR4 (N12303, N12301, N1707, N2911, N2268);
nor NOR2 (N12304, N12303, N11916);
nor NOR3 (N12305, N12294, N11752, N451);
and AND3 (N12306, N12291, N10175, N10610);
and AND4 (N12307, N12297, N8907, N4727, N6427);
not NOT1 (N12308, N12281);
not NOT1 (N12309, N12296);
nand NAND4 (N12310, N12308, N11426, N7632, N4795);
not NOT1 (N12311, N12298);
nor NOR4 (N12312, N12306, N7867, N3188, N8217);
xor XOR2 (N12313, N12304, N9398);
nor NOR4 (N12314, N12299, N1149, N1033, N10453);
buf BUF1 (N12315, N12309);
not NOT1 (N12316, N12302);
or OR2 (N12317, N12310, N3647);
and AND3 (N12318, N12311, N10893, N1347);
not NOT1 (N12319, N12312);
or OR2 (N12320, N12305, N8758);
buf BUF1 (N12321, N12313);
nor NOR3 (N12322, N12321, N3376, N8417);
buf BUF1 (N12323, N12320);
and AND4 (N12324, N12314, N8546, N11042, N739);
buf BUF1 (N12325, N12318);
xor XOR2 (N12326, N12317, N957);
or OR3 (N12327, N12315, N5674, N2087);
or OR3 (N12328, N12322, N9445, N605);
xor XOR2 (N12329, N12327, N6318);
buf BUF1 (N12330, N12324);
nand NAND4 (N12331, N12316, N430, N2734, N7469);
and AND3 (N12332, N12319, N7377, N3860);
xor XOR2 (N12333, N12328, N5327);
not NOT1 (N12334, N12332);
and AND4 (N12335, N12331, N8528, N945, N11660);
nor NOR3 (N12336, N12292, N10165, N4263);
buf BUF1 (N12337, N12325);
buf BUF1 (N12338, N12323);
not NOT1 (N12339, N12338);
and AND2 (N12340, N12330, N7721);
nor NOR3 (N12341, N12333, N8654, N2663);
and AND4 (N12342, N12329, N9341, N2596, N5930);
buf BUF1 (N12343, N12341);
not NOT1 (N12344, N12334);
or OR3 (N12345, N12337, N1486, N11015);
nor NOR3 (N12346, N12326, N5565, N8986);
and AND3 (N12347, N12344, N7096, N8207);
and AND3 (N12348, N12342, N5179, N10314);
buf BUF1 (N12349, N12336);
nor NOR4 (N12350, N12339, N8387, N1034, N8272);
not NOT1 (N12351, N12347);
not NOT1 (N12352, N12345);
buf BUF1 (N12353, N12351);
nand NAND4 (N12354, N12348, N11196, N8901, N7638);
not NOT1 (N12355, N12346);
and AND3 (N12356, N12335, N1583, N5350);
not NOT1 (N12357, N12343);
and AND2 (N12358, N12340, N8559);
xor XOR2 (N12359, N12358, N10775);
buf BUF1 (N12360, N12359);
nand NAND2 (N12361, N12356, N3021);
nor NOR2 (N12362, N12353, N10399);
xor XOR2 (N12363, N12349, N10529);
nand NAND4 (N12364, N12360, N8598, N2638, N6085);
or OR2 (N12365, N12354, N1738);
buf BUF1 (N12366, N12307);
not NOT1 (N12367, N12361);
nor NOR4 (N12368, N12352, N4666, N7947, N1971);
or OR4 (N12369, N12364, N1479, N7550, N3799);
or OR2 (N12370, N12362, N9259);
and AND2 (N12371, N12369, N2713);
buf BUF1 (N12372, N12371);
not NOT1 (N12373, N12365);
nor NOR4 (N12374, N12366, N399, N6076, N1979);
buf BUF1 (N12375, N12370);
or OR4 (N12376, N12350, N7858, N589, N7447);
nand NAND3 (N12377, N12355, N7308, N7911);
nand NAND3 (N12378, N12374, N10486, N5903);
or OR3 (N12379, N12357, N2984, N4751);
or OR2 (N12380, N12377, N8287);
nand NAND2 (N12381, N12373, N9771);
not NOT1 (N12382, N12372);
nand NAND4 (N12383, N12376, N6030, N8699, N5011);
nor NOR3 (N12384, N12382, N1827, N8098);
nand NAND3 (N12385, N12367, N1968, N10185);
and AND3 (N12386, N12363, N1645, N3312);
or OR3 (N12387, N12380, N6698, N12021);
buf BUF1 (N12388, N12375);
and AND4 (N12389, N12383, N5090, N5043, N4055);
buf BUF1 (N12390, N12381);
and AND4 (N12391, N12384, N9335, N2521, N627);
nand NAND3 (N12392, N12386, N12296, N9189);
nor NOR2 (N12393, N12387, N1918);
xor XOR2 (N12394, N12393, N8246);
nor NOR4 (N12395, N12391, N7521, N3995, N5212);
and AND3 (N12396, N12368, N1511, N7617);
or OR4 (N12397, N12394, N2551, N5324, N2055);
or OR4 (N12398, N12385, N292, N1624, N1225);
not NOT1 (N12399, N12398);
nor NOR4 (N12400, N12399, N2842, N9806, N11244);
buf BUF1 (N12401, N12379);
and AND3 (N12402, N12388, N7992, N1919);
nor NOR3 (N12403, N12402, N5648, N2312);
nand NAND3 (N12404, N12400, N11303, N5557);
xor XOR2 (N12405, N12378, N6687);
and AND3 (N12406, N12396, N12072, N39);
not NOT1 (N12407, N12397);
and AND2 (N12408, N12406, N9592);
buf BUF1 (N12409, N12405);
buf BUF1 (N12410, N12392);
nor NOR4 (N12411, N12389, N1767, N11475, N2366);
or OR3 (N12412, N12409, N1688, N3138);
and AND2 (N12413, N12390, N10020);
nor NOR2 (N12414, N12412, N2202);
nand NAND4 (N12415, N12408, N6069, N8208, N2559);
buf BUF1 (N12416, N12407);
buf BUF1 (N12417, N12416);
buf BUF1 (N12418, N12415);
nand NAND4 (N12419, N12411, N7532, N6432, N1538);
nor NOR3 (N12420, N12401, N12038, N8400);
nor NOR2 (N12421, N12418, N6887);
or OR4 (N12422, N12413, N11941, N11620, N1259);
or OR3 (N12423, N12403, N12282, N9599);
or OR4 (N12424, N12395, N7498, N10846, N263);
not NOT1 (N12425, N12424);
or OR2 (N12426, N12417, N376);
nor NOR4 (N12427, N12422, N308, N1807, N8677);
and AND4 (N12428, N12426, N7710, N1619, N5415);
and AND2 (N12429, N12428, N7191);
not NOT1 (N12430, N12429);
nand NAND4 (N12431, N12425, N4774, N10809, N3827);
xor XOR2 (N12432, N12419, N3034);
nand NAND3 (N12433, N12427, N7059, N12069);
not NOT1 (N12434, N12410);
and AND2 (N12435, N12430, N11214);
buf BUF1 (N12436, N12414);
nor NOR4 (N12437, N12432, N360, N9967, N11206);
or OR2 (N12438, N12434, N401);
not NOT1 (N12439, N12436);
and AND2 (N12440, N12421, N2465);
xor XOR2 (N12441, N12423, N4190);
nor NOR2 (N12442, N12433, N6413);
and AND2 (N12443, N12437, N2842);
or OR3 (N12444, N12431, N2427, N7138);
and AND2 (N12445, N12435, N10826);
or OR3 (N12446, N12439, N5650, N5380);
not NOT1 (N12447, N12441);
buf BUF1 (N12448, N12447);
buf BUF1 (N12449, N12420);
buf BUF1 (N12450, N12440);
nor NOR3 (N12451, N12450, N11210, N10853);
nand NAND2 (N12452, N12448, N529);
and AND3 (N12453, N12404, N9771, N4420);
or OR3 (N12454, N12449, N1318, N10970);
buf BUF1 (N12455, N12438);
xor XOR2 (N12456, N12451, N4154);
buf BUF1 (N12457, N12442);
and AND3 (N12458, N12456, N4809, N1494);
nand NAND3 (N12459, N12452, N8551, N9116);
nor NOR3 (N12460, N12454, N9730, N2925);
and AND2 (N12461, N12443, N9204);
nor NOR4 (N12462, N12455, N10398, N9628, N7099);
xor XOR2 (N12463, N12446, N2689);
buf BUF1 (N12464, N12445);
and AND3 (N12465, N12464, N7165, N962);
nand NAND2 (N12466, N12462, N5972);
xor XOR2 (N12467, N12458, N54);
buf BUF1 (N12468, N12444);
not NOT1 (N12469, N12463);
buf BUF1 (N12470, N12453);
not NOT1 (N12471, N12466);
xor XOR2 (N12472, N12459, N5427);
nand NAND4 (N12473, N12470, N6951, N6066, N2916);
xor XOR2 (N12474, N12461, N478);
not NOT1 (N12475, N12471);
and AND2 (N12476, N12468, N12314);
xor XOR2 (N12477, N12473, N11399);
not NOT1 (N12478, N12474);
nor NOR3 (N12479, N12478, N7507, N8190);
and AND2 (N12480, N12457, N2627);
or OR3 (N12481, N12472, N5808, N12096);
buf BUF1 (N12482, N12475);
and AND2 (N12483, N12479, N1206);
xor XOR2 (N12484, N12465, N11599);
buf BUF1 (N12485, N12480);
buf BUF1 (N12486, N12485);
not NOT1 (N12487, N12483);
xor XOR2 (N12488, N12460, N2485);
nor NOR3 (N12489, N12488, N10516, N1088);
xor XOR2 (N12490, N12482, N11989);
and AND2 (N12491, N12477, N5435);
nor NOR4 (N12492, N12469, N6598, N10555, N6776);
not NOT1 (N12493, N12476);
nand NAND2 (N12494, N12490, N11583);
xor XOR2 (N12495, N12492, N9197);
nand NAND3 (N12496, N12493, N350, N1500);
nand NAND3 (N12497, N12495, N6500, N10084);
or OR3 (N12498, N12496, N5808, N5834);
xor XOR2 (N12499, N12484, N10393);
nor NOR4 (N12500, N12499, N2036, N1688, N6373);
or OR3 (N12501, N12481, N5788, N3961);
buf BUF1 (N12502, N12486);
nor NOR4 (N12503, N12489, N26, N6773, N8868);
or OR3 (N12504, N12487, N6648, N2939);
xor XOR2 (N12505, N12502, N6918);
nor NOR4 (N12506, N12503, N5917, N609, N646);
and AND3 (N12507, N12467, N149, N7110);
nand NAND4 (N12508, N12498, N4015, N10930, N8612);
xor XOR2 (N12509, N12508, N11745);
buf BUF1 (N12510, N12500);
xor XOR2 (N12511, N12510, N9239);
buf BUF1 (N12512, N12504);
nor NOR2 (N12513, N12506, N4514);
not NOT1 (N12514, N12509);
not NOT1 (N12515, N12511);
buf BUF1 (N12516, N12513);
and AND4 (N12517, N12516, N1806, N2793, N12307);
buf BUF1 (N12518, N12501);
xor XOR2 (N12519, N12507, N8091);
or OR4 (N12520, N12512, N12403, N11425, N8970);
or OR2 (N12521, N12517, N8463);
buf BUF1 (N12522, N12521);
nor NOR2 (N12523, N12497, N4781);
buf BUF1 (N12524, N12522);
nor NOR4 (N12525, N12524, N5905, N12223, N5411);
or OR4 (N12526, N12523, N12202, N10818, N5818);
or OR4 (N12527, N12505, N10505, N8178, N5270);
buf BUF1 (N12528, N12525);
buf BUF1 (N12529, N12519);
and AND2 (N12530, N12518, N2718);
buf BUF1 (N12531, N12530);
or OR2 (N12532, N12491, N5571);
buf BUF1 (N12533, N12531);
buf BUF1 (N12534, N12532);
nand NAND2 (N12535, N12533, N8360);
buf BUF1 (N12536, N12534);
xor XOR2 (N12537, N12515, N2369);
nand NAND4 (N12538, N12494, N8962, N4017, N1527);
buf BUF1 (N12539, N12529);
and AND2 (N12540, N12538, N996);
nand NAND4 (N12541, N12527, N8781, N2459, N4422);
not NOT1 (N12542, N12514);
or OR3 (N12543, N12537, N7163, N7463);
or OR3 (N12544, N12541, N10710, N4608);
buf BUF1 (N12545, N12528);
not NOT1 (N12546, N12544);
nor NOR4 (N12547, N12546, N2644, N2264, N6564);
nand NAND3 (N12548, N12535, N4842, N6353);
or OR3 (N12549, N12539, N6479, N407);
not NOT1 (N12550, N12542);
nand NAND3 (N12551, N12548, N9391, N6099);
xor XOR2 (N12552, N12536, N8014);
and AND4 (N12553, N12549, N10153, N11285, N5430);
nor NOR3 (N12554, N12540, N7690, N9689);
and AND4 (N12555, N12520, N2957, N4390, N12273);
xor XOR2 (N12556, N12543, N12126);
or OR4 (N12557, N12547, N8294, N12077, N4535);
nand NAND2 (N12558, N12526, N9666);
nand NAND3 (N12559, N12545, N3147, N325);
or OR2 (N12560, N12556, N11232);
xor XOR2 (N12561, N12554, N5856);
buf BUF1 (N12562, N12561);
not NOT1 (N12563, N12562);
and AND4 (N12564, N12550, N10007, N905, N7921);
or OR2 (N12565, N12560, N3138);
nand NAND2 (N12566, N12557, N2237);
xor XOR2 (N12567, N12565, N10917);
nand NAND2 (N12568, N12566, N2868);
nand NAND4 (N12569, N12555, N9866, N4226, N10459);
nand NAND4 (N12570, N12552, N4833, N11131, N3563);
nand NAND4 (N12571, N12551, N6625, N11991, N8480);
buf BUF1 (N12572, N12563);
and AND2 (N12573, N12569, N4356);
or OR2 (N12574, N12573, N8573);
and AND4 (N12575, N12564, N5215, N8045, N5824);
or OR3 (N12576, N12571, N4256, N4381);
and AND2 (N12577, N12570, N8608);
not NOT1 (N12578, N12567);
nor NOR3 (N12579, N12568, N528, N3953);
nor NOR3 (N12580, N12553, N9526, N2);
or OR3 (N12581, N12580, N4078, N4294);
and AND2 (N12582, N12578, N3821);
buf BUF1 (N12583, N12581);
not NOT1 (N12584, N12579);
not NOT1 (N12585, N12583);
and AND4 (N12586, N12572, N1750, N2630, N6120);
nand NAND3 (N12587, N12559, N4379, N12156);
not NOT1 (N12588, N12577);
xor XOR2 (N12589, N12575, N5134);
or OR4 (N12590, N12574, N4013, N8206, N4130);
not NOT1 (N12591, N12576);
not NOT1 (N12592, N12587);
nor NOR2 (N12593, N12584, N567);
or OR2 (N12594, N12591, N10352);
not NOT1 (N12595, N12558);
buf BUF1 (N12596, N12595);
or OR4 (N12597, N12588, N5786, N9874, N11294);
buf BUF1 (N12598, N12597);
nand NAND3 (N12599, N12590, N8484, N10706);
buf BUF1 (N12600, N12596);
xor XOR2 (N12601, N12594, N1035);
xor XOR2 (N12602, N12601, N3216);
xor XOR2 (N12603, N12599, N11757);
not NOT1 (N12604, N12586);
or OR4 (N12605, N12582, N1441, N2727, N8135);
or OR2 (N12606, N12602, N4916);
nor NOR4 (N12607, N12605, N11593, N11219, N4449);
xor XOR2 (N12608, N12598, N11602);
nor NOR2 (N12609, N12603, N12078);
xor XOR2 (N12610, N12600, N1321);
buf BUF1 (N12611, N12609);
not NOT1 (N12612, N12610);
buf BUF1 (N12613, N12612);
buf BUF1 (N12614, N12604);
nand NAND2 (N12615, N12606, N641);
nand NAND2 (N12616, N12589, N6755);
or OR2 (N12617, N12614, N6770);
buf BUF1 (N12618, N12615);
nor NOR4 (N12619, N12592, N5979, N5412, N3182);
nand NAND3 (N12620, N12585, N1063, N226);
nand NAND4 (N12621, N12617, N5536, N10697, N9147);
or OR3 (N12622, N12620, N10292, N12416);
or OR2 (N12623, N12611, N8616);
xor XOR2 (N12624, N12593, N1838);
and AND3 (N12625, N12619, N2033, N6022);
buf BUF1 (N12626, N12613);
nor NOR4 (N12627, N12621, N2651, N1760, N6246);
buf BUF1 (N12628, N12626);
not NOT1 (N12629, N12625);
nand NAND3 (N12630, N12618, N8830, N4789);
nor NOR3 (N12631, N12608, N608, N29);
nor NOR2 (N12632, N12630, N1263);
buf BUF1 (N12633, N12627);
nand NAND3 (N12634, N12623, N4019, N3076);
nand NAND2 (N12635, N12631, N3799);
and AND3 (N12636, N12632, N11397, N10826);
or OR3 (N12637, N12616, N10305, N2630);
and AND4 (N12638, N12634, N2078, N11245, N5141);
buf BUF1 (N12639, N12624);
nor NOR3 (N12640, N12629, N2234, N12417);
not NOT1 (N12641, N12622);
or OR3 (N12642, N12637, N8344, N4023);
nor NOR2 (N12643, N12628, N6644);
not NOT1 (N12644, N12643);
or OR2 (N12645, N12639, N6200);
nand NAND3 (N12646, N12638, N3220, N8782);
buf BUF1 (N12647, N12635);
nor NOR4 (N12648, N12641, N7102, N2642, N12568);
nor NOR2 (N12649, N12640, N4035);
or OR2 (N12650, N12647, N5510);
or OR4 (N12651, N12636, N7408, N2936, N2351);
or OR4 (N12652, N12645, N11084, N10104, N3693);
or OR3 (N12653, N12633, N2522, N12309);
nand NAND3 (N12654, N12653, N5478, N8998);
buf BUF1 (N12655, N12607);
nand NAND3 (N12656, N12654, N7137, N3454);
not NOT1 (N12657, N12655);
and AND3 (N12658, N12657, N11137, N12523);
not NOT1 (N12659, N12650);
nor NOR2 (N12660, N12651, N10233);
xor XOR2 (N12661, N12642, N6649);
xor XOR2 (N12662, N12644, N6122);
nand NAND4 (N12663, N12646, N5053, N8102, N3448);
not NOT1 (N12664, N12656);
not NOT1 (N12665, N12649);
and AND4 (N12666, N12659, N6540, N7559, N3083);
or OR2 (N12667, N12648, N3757);
xor XOR2 (N12668, N12658, N2354);
or OR3 (N12669, N12660, N226, N7241);
not NOT1 (N12670, N12668);
not NOT1 (N12671, N12666);
nor NOR3 (N12672, N12652, N6149, N6965);
not NOT1 (N12673, N12669);
buf BUF1 (N12674, N12664);
buf BUF1 (N12675, N12663);
nor NOR3 (N12676, N12665, N5301, N146);
and AND2 (N12677, N12671, N5874);
not NOT1 (N12678, N12675);
not NOT1 (N12679, N12670);
buf BUF1 (N12680, N12674);
nand NAND3 (N12681, N12679, N2942, N1838);
xor XOR2 (N12682, N12678, N378);
or OR4 (N12683, N12682, N6913, N7595, N1481);
nor NOR2 (N12684, N12662, N10228);
not NOT1 (N12685, N12681);
xor XOR2 (N12686, N12673, N4676);
nor NOR4 (N12687, N12677, N5662, N7849, N8284);
buf BUF1 (N12688, N12685);
not NOT1 (N12689, N12684);
not NOT1 (N12690, N12689);
not NOT1 (N12691, N12687);
nor NOR3 (N12692, N12661, N5284, N112);
and AND2 (N12693, N12683, N3730);
or OR4 (N12694, N12691, N5912, N1508, N5490);
or OR2 (N12695, N12672, N4210);
or OR3 (N12696, N12680, N9436, N5408);
nor NOR4 (N12697, N12696, N2219, N8097, N9880);
or OR4 (N12698, N12690, N9847, N12103, N10678);
and AND2 (N12699, N12698, N3793);
nand NAND4 (N12700, N12699, N7811, N8964, N3074);
or OR2 (N12701, N12694, N10680);
not NOT1 (N12702, N12700);
and AND3 (N12703, N12693, N8067, N7637);
buf BUF1 (N12704, N12701);
not NOT1 (N12705, N12667);
nor NOR4 (N12706, N12704, N4602, N12359, N2034);
not NOT1 (N12707, N12702);
buf BUF1 (N12708, N12707);
nor NOR3 (N12709, N12692, N615, N5775);
nor NOR4 (N12710, N12695, N10719, N4414, N3902);
nor NOR2 (N12711, N12703, N607);
nor NOR4 (N12712, N12706, N11535, N3729, N1380);
or OR4 (N12713, N12712, N2280, N5369, N3743);
nand NAND2 (N12714, N12697, N4809);
not NOT1 (N12715, N12708);
and AND2 (N12716, N12714, N12085);
xor XOR2 (N12717, N12710, N11143);
nand NAND2 (N12718, N12686, N3020);
and AND3 (N12719, N12705, N8859, N1696);
not NOT1 (N12720, N12716);
nand NAND2 (N12721, N12709, N6436);
xor XOR2 (N12722, N12721, N1568);
nor NOR2 (N12723, N12688, N1308);
xor XOR2 (N12724, N12713, N1398);
nand NAND4 (N12725, N12717, N11837, N2219, N12599);
xor XOR2 (N12726, N12720, N6689);
nand NAND3 (N12727, N12725, N9437, N5636);
not NOT1 (N12728, N12723);
buf BUF1 (N12729, N12718);
nor NOR4 (N12730, N12722, N3039, N6101, N10177);
nand NAND4 (N12731, N12728, N4147, N4210, N12240);
xor XOR2 (N12732, N12730, N4083);
or OR3 (N12733, N12731, N5478, N12028);
nor NOR3 (N12734, N12729, N3019, N12661);
xor XOR2 (N12735, N12719, N208);
or OR2 (N12736, N12724, N5182);
xor XOR2 (N12737, N12733, N383);
nand NAND2 (N12738, N12736, N7034);
nor NOR2 (N12739, N12735, N3390);
not NOT1 (N12740, N12726);
nand NAND2 (N12741, N12676, N6893);
and AND4 (N12742, N12727, N3176, N7320, N10955);
nand NAND3 (N12743, N12711, N444, N159);
xor XOR2 (N12744, N12739, N5372);
xor XOR2 (N12745, N12737, N10631);
nor NOR3 (N12746, N12745, N12185, N10838);
and AND3 (N12747, N12740, N5264, N2229);
and AND4 (N12748, N12738, N2245, N10049, N971);
xor XOR2 (N12749, N12742, N10902);
or OR2 (N12750, N12732, N8940);
not NOT1 (N12751, N12746);
or OR2 (N12752, N12734, N1956);
buf BUF1 (N12753, N12744);
or OR4 (N12754, N12751, N8490, N4136, N3071);
nand NAND2 (N12755, N12747, N8854);
or OR4 (N12756, N12749, N8898, N6924, N12179);
and AND2 (N12757, N12715, N10059);
and AND2 (N12758, N12756, N5689);
or OR4 (N12759, N12748, N1639, N4535, N6602);
not NOT1 (N12760, N12741);
not NOT1 (N12761, N12754);
not NOT1 (N12762, N12758);
or OR3 (N12763, N12755, N7026, N11332);
and AND2 (N12764, N12762, N11825);
or OR3 (N12765, N12753, N3547, N5227);
nand NAND3 (N12766, N12763, N2554, N7852);
or OR3 (N12767, N12757, N7337, N1797);
or OR4 (N12768, N12760, N7960, N10760, N3242);
xor XOR2 (N12769, N12768, N4739);
or OR4 (N12770, N12752, N4789, N1039, N7105);
xor XOR2 (N12771, N12767, N3491);
nor NOR4 (N12772, N12743, N11240, N27, N4637);
nor NOR3 (N12773, N12765, N3574, N11414);
buf BUF1 (N12774, N12761);
nor NOR3 (N12775, N12772, N2317, N2310);
nand NAND4 (N12776, N12773, N5903, N7421, N74);
xor XOR2 (N12777, N12775, N10311);
and AND3 (N12778, N12771, N11735, N1480);
not NOT1 (N12779, N12778);
nor NOR4 (N12780, N12770, N6030, N245, N9454);
nand NAND4 (N12781, N12774, N5223, N10155, N6256);
not NOT1 (N12782, N12764);
nor NOR3 (N12783, N12782, N3213, N8616);
xor XOR2 (N12784, N12759, N8512);
or OR4 (N12785, N12750, N7458, N3881, N7657);
xor XOR2 (N12786, N12784, N2519);
or OR3 (N12787, N12766, N1913, N8825);
not NOT1 (N12788, N12781);
not NOT1 (N12789, N12777);
buf BUF1 (N12790, N12785);
nand NAND3 (N12791, N12783, N5463, N4241);
buf BUF1 (N12792, N12769);
not NOT1 (N12793, N12779);
and AND3 (N12794, N12792, N2501, N1158);
or OR3 (N12795, N12776, N10874, N11315);
xor XOR2 (N12796, N12791, N6199);
not NOT1 (N12797, N12780);
and AND3 (N12798, N12793, N436, N6246);
not NOT1 (N12799, N12795);
and AND3 (N12800, N12786, N8666, N12024);
and AND3 (N12801, N12790, N8083, N4230);
and AND3 (N12802, N12794, N1606, N8083);
buf BUF1 (N12803, N12788);
xor XOR2 (N12804, N12800, N4058);
nor NOR4 (N12805, N12798, N2479, N6967, N3534);
and AND4 (N12806, N12801, N3758, N1297, N7371);
and AND3 (N12807, N12804, N4899, N7569);
and AND3 (N12808, N12797, N1254, N3614);
xor XOR2 (N12809, N12799, N6939);
xor XOR2 (N12810, N12789, N5196);
or OR3 (N12811, N12806, N9636, N4708);
xor XOR2 (N12812, N12808, N2498);
nor NOR2 (N12813, N12810, N5048);
not NOT1 (N12814, N12805);
buf BUF1 (N12815, N12802);
and AND2 (N12816, N12807, N1736);
nand NAND2 (N12817, N12811, N11015);
not NOT1 (N12818, N12812);
and AND2 (N12819, N12817, N11511);
nand NAND2 (N12820, N12813, N567);
or OR2 (N12821, N12816, N9213);
and AND3 (N12822, N12796, N8711, N10540);
and AND3 (N12823, N12815, N2187, N11781);
nand NAND2 (N12824, N12820, N9295);
nand NAND3 (N12825, N12822, N10434, N6930);
or OR3 (N12826, N12809, N220, N1982);
and AND4 (N12827, N12803, N5080, N10009, N3096);
xor XOR2 (N12828, N12827, N5403);
xor XOR2 (N12829, N12823, N7376);
buf BUF1 (N12830, N12824);
and AND2 (N12831, N12826, N11738);
and AND3 (N12832, N12818, N5598, N11859);
or OR2 (N12833, N12829, N9418);
or OR3 (N12834, N12832, N12372, N6411);
nand NAND2 (N12835, N12831, N3386);
nand NAND3 (N12836, N12828, N2422, N1048);
xor XOR2 (N12837, N12825, N5160);
not NOT1 (N12838, N12814);
and AND2 (N12839, N12787, N10746);
not NOT1 (N12840, N12838);
and AND2 (N12841, N12819, N8554);
xor XOR2 (N12842, N12834, N8916);
not NOT1 (N12843, N12842);
nand NAND2 (N12844, N12841, N5987);
xor XOR2 (N12845, N12835, N2915);
nor NOR4 (N12846, N12833, N9123, N12595, N7163);
xor XOR2 (N12847, N12843, N12377);
and AND3 (N12848, N12830, N9861, N7697);
buf BUF1 (N12849, N12840);
or OR4 (N12850, N12821, N9422, N1703, N11588);
nor NOR3 (N12851, N12849, N2938, N4597);
nand NAND4 (N12852, N12846, N7390, N226, N4625);
or OR4 (N12853, N12848, N3151, N4269, N6867);
buf BUF1 (N12854, N12839);
and AND2 (N12855, N12845, N12157);
nand NAND3 (N12856, N12852, N5120, N5774);
or OR2 (N12857, N12856, N3821);
buf BUF1 (N12858, N12836);
nor NOR4 (N12859, N12851, N7053, N10510, N3595);
xor XOR2 (N12860, N12855, N3757);
nand NAND3 (N12861, N12859, N2351, N244);
nor NOR4 (N12862, N12844, N9773, N8868, N7696);
not NOT1 (N12863, N12857);
or OR3 (N12864, N12863, N4404, N1759);
nor NOR4 (N12865, N12847, N1374, N2360, N9769);
nand NAND4 (N12866, N12853, N6794, N3802, N1120);
buf BUF1 (N12867, N12850);
buf BUF1 (N12868, N12865);
xor XOR2 (N12869, N12854, N9773);
not NOT1 (N12870, N12869);
xor XOR2 (N12871, N12861, N3062);
buf BUF1 (N12872, N12866);
nand NAND3 (N12873, N12858, N6867, N4654);
xor XOR2 (N12874, N12864, N3077);
nor NOR3 (N12875, N12874, N11868, N11804);
nor NOR3 (N12876, N12868, N9328, N4642);
or OR3 (N12877, N12862, N10737, N12241);
nor NOR4 (N12878, N12871, N566, N491, N12699);
buf BUF1 (N12879, N12837);
nand NAND2 (N12880, N12878, N5248);
nand NAND2 (N12881, N12873, N9397);
and AND2 (N12882, N12872, N5279);
nor NOR4 (N12883, N12860, N6095, N214, N3206);
buf BUF1 (N12884, N12876);
nor NOR2 (N12885, N12870, N6609);
xor XOR2 (N12886, N12885, N5313);
nor NOR4 (N12887, N12879, N8625, N6306, N3076);
and AND2 (N12888, N12886, N3486);
buf BUF1 (N12889, N12880);
and AND4 (N12890, N12875, N11083, N4643, N7236);
and AND2 (N12891, N12884, N11875);
and AND3 (N12892, N12891, N11831, N11562);
not NOT1 (N12893, N12892);
nor NOR4 (N12894, N12881, N3032, N2003, N4185);
nor NOR2 (N12895, N12893, N1135);
nand NAND3 (N12896, N12889, N9701, N3989);
and AND2 (N12897, N12877, N8817);
nand NAND3 (N12898, N12882, N6967, N5302);
and AND2 (N12899, N12897, N9889);
nand NAND4 (N12900, N12895, N2902, N12631, N3213);
or OR4 (N12901, N12899, N9987, N10701, N10271);
and AND2 (N12902, N12901, N10922);
buf BUF1 (N12903, N12902);
nor NOR3 (N12904, N12887, N4077, N7375);
nand NAND2 (N12905, N12888, N805);
or OR3 (N12906, N12883, N12553, N454);
or OR4 (N12907, N12904, N9343, N5450, N10529);
buf BUF1 (N12908, N12903);
or OR3 (N12909, N12896, N4126, N10224);
xor XOR2 (N12910, N12908, N2375);
nor NOR2 (N12911, N12907, N9885);
xor XOR2 (N12912, N12894, N11560);
nor NOR2 (N12913, N12909, N12209);
not NOT1 (N12914, N12900);
xor XOR2 (N12915, N12898, N8384);
nor NOR4 (N12916, N12915, N12794, N5207, N8782);
not NOT1 (N12917, N12906);
and AND3 (N12918, N12914, N5557, N6864);
nor NOR2 (N12919, N12905, N6441);
not NOT1 (N12920, N12910);
or OR4 (N12921, N12890, N17, N7707, N4813);
buf BUF1 (N12922, N12917);
nor NOR3 (N12923, N12922, N8915, N2154);
and AND2 (N12924, N12916, N6974);
buf BUF1 (N12925, N12918);
and AND2 (N12926, N12920, N8399);
nor NOR4 (N12927, N12926, N11648, N9993, N10932);
and AND2 (N12928, N12919, N2779);
xor XOR2 (N12929, N12923, N4949);
buf BUF1 (N12930, N12911);
nor NOR3 (N12931, N12925, N3528, N3160);
nor NOR4 (N12932, N12929, N932, N2021, N548);
nand NAND3 (N12933, N12913, N3521, N5539);
nand NAND4 (N12934, N12932, N4058, N11808, N3884);
xor XOR2 (N12935, N12924, N7488);
nor NOR3 (N12936, N12867, N2729, N12338);
or OR2 (N12937, N12912, N10265);
or OR4 (N12938, N12921, N12659, N7677, N2584);
buf BUF1 (N12939, N12935);
not NOT1 (N12940, N12933);
nor NOR3 (N12941, N12939, N3446, N6511);
nand NAND3 (N12942, N12931, N7500, N10405);
buf BUF1 (N12943, N12934);
or OR4 (N12944, N12936, N3482, N11517, N3259);
or OR2 (N12945, N12944, N9642);
not NOT1 (N12946, N12938);
or OR4 (N12947, N12946, N8469, N4089, N10956);
not NOT1 (N12948, N12942);
nor NOR3 (N12949, N12941, N1870, N3017);
or OR3 (N12950, N12930, N8175, N5673);
buf BUF1 (N12951, N12927);
not NOT1 (N12952, N12937);
xor XOR2 (N12953, N12948, N4581);
buf BUF1 (N12954, N12928);
xor XOR2 (N12955, N12952, N5769);
nor NOR2 (N12956, N12945, N11478);
xor XOR2 (N12957, N12953, N7958);
and AND4 (N12958, N12955, N10219, N1131, N12163);
buf BUF1 (N12959, N12956);
or OR2 (N12960, N12949, N841);
and AND2 (N12961, N12954, N2315);
buf BUF1 (N12962, N12951);
nor NOR4 (N12963, N12960, N12290, N11374, N9314);
nor NOR3 (N12964, N12961, N10818, N3803);
not NOT1 (N12965, N12962);
nor NOR2 (N12966, N12958, N4211);
buf BUF1 (N12967, N12964);
and AND2 (N12968, N12957, N6401);
buf BUF1 (N12969, N12947);
or OR3 (N12970, N12969, N6969, N2981);
and AND2 (N12971, N12940, N10301);
nand NAND3 (N12972, N12959, N9484, N9582);
not NOT1 (N12973, N12950);
not NOT1 (N12974, N12972);
not NOT1 (N12975, N12970);
not NOT1 (N12976, N12971);
or OR3 (N12977, N12965, N1625, N10541);
nand NAND4 (N12978, N12967, N7342, N4020, N12040);
buf BUF1 (N12979, N12963);
nor NOR2 (N12980, N12976, N1878);
not NOT1 (N12981, N12979);
nor NOR2 (N12982, N12975, N12587);
nand NAND2 (N12983, N12981, N9481);
not NOT1 (N12984, N12977);
nand NAND4 (N12985, N12968, N3796, N5848, N5140);
buf BUF1 (N12986, N12983);
buf BUF1 (N12987, N12980);
and AND3 (N12988, N12987, N59, N8077);
and AND4 (N12989, N12943, N1550, N12784, N6790);
buf BUF1 (N12990, N12982);
and AND3 (N12991, N12988, N9053, N11443);
or OR4 (N12992, N12978, N7650, N6163, N1302);
xor XOR2 (N12993, N12992, N2449);
buf BUF1 (N12994, N12984);
or OR3 (N12995, N12985, N9118, N12088);
xor XOR2 (N12996, N12994, N7842);
nor NOR3 (N12997, N12973, N7573, N1831);
and AND2 (N12998, N12986, N3063);
not NOT1 (N12999, N12993);
or OR3 (N13000, N12974, N10553, N3453);
buf BUF1 (N13001, N12990);
and AND4 (N13002, N12997, N3398, N8423, N12916);
nor NOR2 (N13003, N12995, N1907);
xor XOR2 (N13004, N12991, N8678);
xor XOR2 (N13005, N13000, N12136);
nand NAND2 (N13006, N13004, N5645);
nand NAND3 (N13007, N13005, N4934, N2287);
and AND4 (N13008, N13001, N9875, N11661, N3009);
buf BUF1 (N13009, N12996);
and AND3 (N13010, N13006, N8825, N10090);
xor XOR2 (N13011, N13007, N2541);
and AND2 (N13012, N12966, N12443);
nor NOR2 (N13013, N12989, N12679);
buf BUF1 (N13014, N13012);
or OR4 (N13015, N12999, N12872, N1105, N1894);
or OR4 (N13016, N13009, N7457, N10090, N812);
nand NAND3 (N13017, N12998, N11073, N2606);
or OR3 (N13018, N13008, N5972, N11855);
or OR4 (N13019, N13015, N2307, N3933, N5996);
not NOT1 (N13020, N13014);
xor XOR2 (N13021, N13011, N10940);
nor NOR2 (N13022, N13010, N8075);
xor XOR2 (N13023, N13002, N12219);
and AND3 (N13024, N13023, N11064, N8556);
nor NOR3 (N13025, N13016, N6931, N5614);
not NOT1 (N13026, N13013);
and AND3 (N13027, N13017, N6612, N7410);
xor XOR2 (N13028, N13025, N12371);
nand NAND2 (N13029, N13020, N3348);
nor NOR3 (N13030, N13021, N2142, N8086);
buf BUF1 (N13031, N13030);
or OR3 (N13032, N13018, N1360, N4222);
nand NAND2 (N13033, N13003, N9312);
or OR4 (N13034, N13019, N12559, N3092, N11945);
buf BUF1 (N13035, N13022);
or OR2 (N13036, N13034, N6142);
nor NOR3 (N13037, N13027, N5324, N2618);
buf BUF1 (N13038, N13028);
or OR4 (N13039, N13037, N7825, N12632, N12428);
or OR3 (N13040, N13038, N1255, N12420);
and AND3 (N13041, N13036, N7121, N1783);
buf BUF1 (N13042, N13040);
not NOT1 (N13043, N13041);
or OR4 (N13044, N13024, N4434, N7189, N6159);
or OR4 (N13045, N13031, N10505, N8980, N11440);
xor XOR2 (N13046, N13044, N7855);
or OR2 (N13047, N13043, N695);
xor XOR2 (N13048, N13026, N3626);
and AND4 (N13049, N13035, N7450, N5547, N8278);
xor XOR2 (N13050, N13048, N7961);
buf BUF1 (N13051, N13029);
or OR2 (N13052, N13050, N7996);
or OR2 (N13053, N13046, N9967);
nor NOR4 (N13054, N13053, N5954, N6620, N5322);
and AND4 (N13055, N13054, N8076, N2383, N6072);
nand NAND2 (N13056, N13032, N4263);
or OR4 (N13057, N13039, N9331, N109, N5194);
and AND4 (N13058, N13049, N9197, N8905, N8287);
not NOT1 (N13059, N13056);
and AND4 (N13060, N13042, N549, N7973, N4879);
or OR2 (N13061, N13052, N1600);
buf BUF1 (N13062, N13045);
not NOT1 (N13063, N13058);
and AND2 (N13064, N13047, N1024);
or OR3 (N13065, N13061, N10863, N2280);
not NOT1 (N13066, N13062);
nand NAND4 (N13067, N13066, N2007, N8727, N3243);
or OR2 (N13068, N13067, N7943);
buf BUF1 (N13069, N13033);
or OR4 (N13070, N13064, N8048, N2002, N7066);
nor NOR4 (N13071, N13063, N4683, N9992, N10224);
not NOT1 (N13072, N13068);
buf BUF1 (N13073, N13055);
nand NAND2 (N13074, N13057, N12487);
nor NOR3 (N13075, N13060, N318, N9191);
buf BUF1 (N13076, N13070);
or OR2 (N13077, N13076, N9635);
or OR2 (N13078, N13069, N7972);
nand NAND2 (N13079, N13059, N12863);
buf BUF1 (N13080, N13073);
nand NAND2 (N13081, N13079, N4722);
nand NAND2 (N13082, N13081, N11361);
buf BUF1 (N13083, N13071);
nand NAND4 (N13084, N13078, N9746, N3207, N12355);
or OR2 (N13085, N13080, N77);
nor NOR2 (N13086, N13085, N3807);
and AND2 (N13087, N13072, N4069);
or OR3 (N13088, N13065, N8300, N12667);
buf BUF1 (N13089, N13082);
buf BUF1 (N13090, N13051);
xor XOR2 (N13091, N13083, N1455);
nand NAND2 (N13092, N13087, N10240);
buf BUF1 (N13093, N13074);
nor NOR4 (N13094, N13092, N7478, N11588, N5138);
nand NAND3 (N13095, N13086, N10373, N6711);
and AND2 (N13096, N13088, N581);
buf BUF1 (N13097, N13091);
buf BUF1 (N13098, N13075);
xor XOR2 (N13099, N13098, N9327);
nor NOR3 (N13100, N13093, N7782, N993);
not NOT1 (N13101, N13097);
nand NAND2 (N13102, N13094, N1109);
buf BUF1 (N13103, N13102);
xor XOR2 (N13104, N13096, N3612);
buf BUF1 (N13105, N13103);
buf BUF1 (N13106, N13077);
xor XOR2 (N13107, N13095, N5669);
nor NOR3 (N13108, N13106, N10850, N9590);
nor NOR3 (N13109, N13101, N3014, N6076);
xor XOR2 (N13110, N13104, N8790);
not NOT1 (N13111, N13099);
or OR4 (N13112, N13105, N5484, N12193, N3767);
or OR3 (N13113, N13110, N7333, N8714);
or OR3 (N13114, N13113, N4072, N8693);
nand NAND4 (N13115, N13109, N1328, N9779, N2196);
xor XOR2 (N13116, N13112, N5960);
and AND2 (N13117, N13100, N594);
nor NOR3 (N13118, N13111, N2591, N220);
nor NOR2 (N13119, N13108, N7652);
buf BUF1 (N13120, N13116);
nand NAND3 (N13121, N13084, N5426, N12551);
and AND3 (N13122, N13118, N2261, N4455);
and AND2 (N13123, N13115, N421);
not NOT1 (N13124, N13114);
nor NOR2 (N13125, N13117, N4972);
not NOT1 (N13126, N13124);
buf BUF1 (N13127, N13119);
xor XOR2 (N13128, N13122, N5183);
buf BUF1 (N13129, N13123);
nor NOR2 (N13130, N13121, N9332);
not NOT1 (N13131, N13129);
or OR3 (N13132, N13126, N4269, N109);
or OR3 (N13133, N13090, N7281, N304);
or OR2 (N13134, N13125, N333);
buf BUF1 (N13135, N13107);
not NOT1 (N13136, N13130);
xor XOR2 (N13137, N13132, N7558);
and AND4 (N13138, N13120, N5890, N10517, N753);
nor NOR3 (N13139, N13127, N11372, N2743);
or OR4 (N13140, N13139, N148, N10692, N7425);
xor XOR2 (N13141, N13140, N8741);
nand NAND3 (N13142, N13131, N10587, N4203);
nand NAND3 (N13143, N13133, N8628, N6403);
and AND4 (N13144, N13136, N7305, N6873, N6490);
and AND2 (N13145, N13135, N7948);
nand NAND3 (N13146, N13144, N10212, N10557);
nor NOR2 (N13147, N13146, N9845);
nor NOR2 (N13148, N13145, N6477);
buf BUF1 (N13149, N13141);
and AND3 (N13150, N13134, N6413, N9219);
buf BUF1 (N13151, N13138);
or OR2 (N13152, N13148, N10955);
nor NOR2 (N13153, N13149, N464);
or OR2 (N13154, N13151, N3284);
not NOT1 (N13155, N13147);
or OR2 (N13156, N13143, N6690);
nor NOR4 (N13157, N13128, N3377, N11132, N4380);
buf BUF1 (N13158, N13089);
nor NOR3 (N13159, N13137, N10971, N5600);
nor NOR2 (N13160, N13152, N9403);
buf BUF1 (N13161, N13157);
or OR3 (N13162, N13150, N11017, N397);
nand NAND4 (N13163, N13155, N3356, N12113, N3196);
nor NOR4 (N13164, N13161, N5996, N203, N949);
nand NAND2 (N13165, N13163, N8325);
and AND2 (N13166, N13154, N9891);
buf BUF1 (N13167, N13162);
nand NAND4 (N13168, N13165, N4180, N10225, N12820);
not NOT1 (N13169, N13156);
nor NOR2 (N13170, N13153, N10011);
not NOT1 (N13171, N13168);
buf BUF1 (N13172, N13167);
xor XOR2 (N13173, N13159, N4376);
or OR3 (N13174, N13164, N1768, N13152);
and AND3 (N13175, N13169, N2724, N5514);
not NOT1 (N13176, N13174);
xor XOR2 (N13177, N13166, N8086);
and AND2 (N13178, N13170, N1520);
nor NOR4 (N13179, N13171, N4360, N2947, N11471);
nor NOR3 (N13180, N13175, N12914, N1937);
xor XOR2 (N13181, N13158, N671);
and AND4 (N13182, N13181, N12653, N9471, N4190);
nor NOR4 (N13183, N13172, N8406, N10225, N7595);
xor XOR2 (N13184, N13180, N290);
xor XOR2 (N13185, N13178, N12746);
nor NOR3 (N13186, N13184, N1483, N3943);
xor XOR2 (N13187, N13177, N1615);
not NOT1 (N13188, N13142);
xor XOR2 (N13189, N13160, N8951);
xor XOR2 (N13190, N13189, N1431);
nand NAND4 (N13191, N13187, N9444, N10820, N463);
nand NAND3 (N13192, N13186, N9753, N6086);
or OR4 (N13193, N13173, N10406, N4158, N10717);
xor XOR2 (N13194, N13193, N7029);
xor XOR2 (N13195, N13179, N2542);
not NOT1 (N13196, N13182);
nand NAND3 (N13197, N13190, N10261, N3649);
nor NOR4 (N13198, N13185, N12623, N268, N12312);
or OR3 (N13199, N13188, N8391, N8962);
not NOT1 (N13200, N13192);
buf BUF1 (N13201, N13196);
and AND4 (N13202, N13200, N10206, N9308, N7325);
or OR4 (N13203, N13176, N4426, N7772, N3962);
xor XOR2 (N13204, N13202, N7966);
or OR2 (N13205, N13203, N8656);
or OR3 (N13206, N13201, N11211, N3463);
and AND2 (N13207, N13199, N11386);
not NOT1 (N13208, N13206);
not NOT1 (N13209, N13207);
nand NAND3 (N13210, N13205, N6032, N9778);
xor XOR2 (N13211, N13204, N2159);
nand NAND2 (N13212, N13211, N8548);
nor NOR3 (N13213, N13183, N3929, N10031);
and AND3 (N13214, N13212, N10335, N4280);
nor NOR4 (N13215, N13214, N6326, N8466, N11574);
xor XOR2 (N13216, N13210, N4270);
not NOT1 (N13217, N13194);
nand NAND4 (N13218, N13195, N5154, N5264, N4794);
nand NAND4 (N13219, N13217, N5837, N3321, N4292);
nor NOR2 (N13220, N13191, N11194);
nand NAND4 (N13221, N13197, N8369, N1526, N12999);
not NOT1 (N13222, N13221);
buf BUF1 (N13223, N13208);
not NOT1 (N13224, N13215);
and AND2 (N13225, N13209, N3108);
or OR4 (N13226, N13216, N1979, N7187, N9681);
and AND3 (N13227, N13198, N11816, N11041);
nand NAND4 (N13228, N13213, N7301, N11981, N1263);
nand NAND3 (N13229, N13226, N7061, N4650);
or OR4 (N13230, N13224, N4887, N10126, N8055);
and AND3 (N13231, N13223, N414, N7591);
buf BUF1 (N13232, N13225);
or OR4 (N13233, N13220, N4825, N8933, N3471);
nand NAND3 (N13234, N13231, N9110, N9987);
buf BUF1 (N13235, N13232);
nand NAND2 (N13236, N13227, N12222);
and AND4 (N13237, N13236, N9591, N12277, N743);
not NOT1 (N13238, N13233);
and AND3 (N13239, N13222, N10734, N2768);
buf BUF1 (N13240, N13238);
not NOT1 (N13241, N13235);
nand NAND4 (N13242, N13230, N5999, N11514, N6154);
and AND4 (N13243, N13242, N4390, N1676, N2939);
nand NAND3 (N13244, N13219, N11331, N9717);
nor NOR2 (N13245, N13218, N13016);
not NOT1 (N13246, N13234);
or OR3 (N13247, N13244, N9758, N11353);
buf BUF1 (N13248, N13247);
buf BUF1 (N13249, N13243);
and AND3 (N13250, N13228, N10435, N12878);
xor XOR2 (N13251, N13229, N3134);
and AND3 (N13252, N13249, N11540, N6750);
or OR4 (N13253, N13241, N10748, N1068, N3653);
and AND4 (N13254, N13240, N2366, N1526, N3183);
nand NAND3 (N13255, N13239, N5387, N7088);
and AND4 (N13256, N13250, N11125, N10119, N12052);
nor NOR3 (N13257, N13237, N13005, N3918);
buf BUF1 (N13258, N13257);
and AND3 (N13259, N13253, N1876, N6580);
and AND2 (N13260, N13256, N7760);
nand NAND3 (N13261, N13246, N12655, N4415);
buf BUF1 (N13262, N13255);
not NOT1 (N13263, N13260);
xor XOR2 (N13264, N13261, N2937);
nor NOR3 (N13265, N13264, N667, N4470);
buf BUF1 (N13266, N13262);
nor NOR2 (N13267, N13254, N6662);
nor NOR3 (N13268, N13258, N3959, N3516);
nand NAND4 (N13269, N13245, N6899, N7770, N1184);
nand NAND2 (N13270, N13251, N5697);
or OR3 (N13271, N13268, N1587, N4048);
not NOT1 (N13272, N13266);
nor NOR4 (N13273, N13271, N2810, N2988, N8911);
not NOT1 (N13274, N13272);
buf BUF1 (N13275, N13274);
or OR4 (N13276, N13267, N2541, N12260, N3485);
buf BUF1 (N13277, N13248);
buf BUF1 (N13278, N13252);
not NOT1 (N13279, N13273);
and AND2 (N13280, N13270, N12495);
nor NOR2 (N13281, N13279, N5749);
not NOT1 (N13282, N13263);
not NOT1 (N13283, N13278);
nor NOR2 (N13284, N13275, N12311);
or OR3 (N13285, N13276, N9281, N6333);
nand NAND2 (N13286, N13281, N1013);
not NOT1 (N13287, N13280);
nor NOR3 (N13288, N13287, N4017, N2836);
nand NAND4 (N13289, N13277, N4139, N11358, N6400);
buf BUF1 (N13290, N13259);
and AND4 (N13291, N13283, N1009, N1111, N10014);
and AND3 (N13292, N13285, N2260, N7629);
or OR3 (N13293, N13289, N11897, N7093);
and AND4 (N13294, N13293, N1199, N9595, N11935);
xor XOR2 (N13295, N13294, N2077);
not NOT1 (N13296, N13269);
or OR3 (N13297, N13296, N6662, N12474);
buf BUF1 (N13298, N13282);
nor NOR2 (N13299, N13290, N11628);
or OR2 (N13300, N13288, N2152);
nand NAND4 (N13301, N13292, N199, N9058, N9332);
nor NOR3 (N13302, N13297, N6687, N11259);
buf BUF1 (N13303, N13284);
nand NAND4 (N13304, N13265, N1841, N9421, N13194);
and AND2 (N13305, N13286, N10809);
buf BUF1 (N13306, N13302);
and AND3 (N13307, N13300, N13246, N10602);
and AND2 (N13308, N13305, N12542);
xor XOR2 (N13309, N13301, N5434);
nand NAND4 (N13310, N13309, N7987, N5034, N13002);
not NOT1 (N13311, N13304);
xor XOR2 (N13312, N13291, N5645);
or OR3 (N13313, N13307, N4239, N6429);
nand NAND2 (N13314, N13310, N7044);
nand NAND3 (N13315, N13313, N12107, N12032);
xor XOR2 (N13316, N13314, N11261);
not NOT1 (N13317, N13303);
not NOT1 (N13318, N13311);
buf BUF1 (N13319, N13312);
nand NAND3 (N13320, N13318, N290, N6907);
nor NOR3 (N13321, N13320, N10512, N12359);
or OR3 (N13322, N13316, N2995, N4625);
nand NAND3 (N13323, N13322, N11651, N3017);
nand NAND3 (N13324, N13308, N2774, N7217);
xor XOR2 (N13325, N13306, N9233);
buf BUF1 (N13326, N13315);
buf BUF1 (N13327, N13295);
or OR4 (N13328, N13321, N6931, N5087, N2217);
or OR2 (N13329, N13324, N8784);
not NOT1 (N13330, N13326);
xor XOR2 (N13331, N13325, N6587);
not NOT1 (N13332, N13319);
buf BUF1 (N13333, N13329);
or OR4 (N13334, N13331, N1360, N10906, N10896);
nand NAND2 (N13335, N13298, N497);
buf BUF1 (N13336, N13335);
and AND2 (N13337, N13336, N8626);
not NOT1 (N13338, N13337);
nor NOR4 (N13339, N13317, N6621, N96, N2192);
and AND4 (N13340, N13334, N7445, N2109, N1574);
buf BUF1 (N13341, N13299);
buf BUF1 (N13342, N13327);
nand NAND3 (N13343, N13341, N12204, N9595);
xor XOR2 (N13344, N13340, N484);
buf BUF1 (N13345, N13323);
xor XOR2 (N13346, N13345, N7283);
not NOT1 (N13347, N13343);
not NOT1 (N13348, N13339);
nor NOR3 (N13349, N13348, N2990, N588);
nand NAND4 (N13350, N13328, N7487, N641, N5862);
buf BUF1 (N13351, N13349);
nor NOR3 (N13352, N13347, N3233, N7174);
or OR3 (N13353, N13351, N5577, N4907);
nor NOR2 (N13354, N13344, N5264);
nand NAND4 (N13355, N13330, N10723, N2235, N7253);
not NOT1 (N13356, N13338);
xor XOR2 (N13357, N13354, N1250);
xor XOR2 (N13358, N13355, N213);
buf BUF1 (N13359, N13333);
not NOT1 (N13360, N13353);
or OR4 (N13361, N13357, N12672, N9215, N2981);
nand NAND4 (N13362, N13332, N6126, N11781, N11701);
xor XOR2 (N13363, N13361, N256);
xor XOR2 (N13364, N13356, N4374);
and AND3 (N13365, N13362, N12792, N6766);
and AND4 (N13366, N13346, N10578, N6955, N9266);
and AND4 (N13367, N13358, N174, N7301, N6895);
nand NAND2 (N13368, N13364, N12364);
nand NAND3 (N13369, N13342, N4349, N2154);
buf BUF1 (N13370, N13365);
nor NOR2 (N13371, N13366, N6305);
nand NAND2 (N13372, N13370, N3575);
and AND2 (N13373, N13372, N10483);
xor XOR2 (N13374, N13371, N1070);
not NOT1 (N13375, N13360);
and AND2 (N13376, N13368, N7655);
nand NAND4 (N13377, N13369, N5327, N7189, N13129);
or OR4 (N13378, N13374, N7791, N7856, N12415);
and AND4 (N13379, N13350, N1315, N6625, N3229);
not NOT1 (N13380, N13379);
not NOT1 (N13381, N13363);
nor NOR4 (N13382, N13359, N8661, N2339, N699);
buf BUF1 (N13383, N13378);
and AND3 (N13384, N13376, N4298, N11570);
nor NOR2 (N13385, N13384, N371);
nor NOR3 (N13386, N13373, N12934, N2255);
and AND2 (N13387, N13380, N6012);
nand NAND3 (N13388, N13377, N6659, N1571);
nor NOR4 (N13389, N13387, N11979, N7169, N1728);
nand NAND2 (N13390, N13389, N10754);
nor NOR4 (N13391, N13352, N10868, N2556, N723);
nand NAND2 (N13392, N13390, N9812);
nor NOR4 (N13393, N13388, N10587, N10063, N10539);
nand NAND4 (N13394, N13392, N8807, N12787, N11166);
nor NOR4 (N13395, N13385, N701, N8706, N4931);
not NOT1 (N13396, N13383);
nor NOR2 (N13397, N13381, N5548);
buf BUF1 (N13398, N13394);
nor NOR3 (N13399, N13396, N2746, N4335);
nor NOR3 (N13400, N13382, N7932, N1820);
nor NOR2 (N13401, N13399, N12857);
or OR3 (N13402, N13393, N10093, N4150);
or OR2 (N13403, N13386, N11090);
and AND2 (N13404, N13401, N7041);
and AND2 (N13405, N13398, N1045);
buf BUF1 (N13406, N13403);
buf BUF1 (N13407, N13404);
and AND3 (N13408, N13367, N1334, N11662);
not NOT1 (N13409, N13406);
xor XOR2 (N13410, N13400, N12767);
and AND4 (N13411, N13397, N10900, N5068, N836);
buf BUF1 (N13412, N13411);
nand NAND3 (N13413, N13410, N140, N9598);
buf BUF1 (N13414, N13407);
not NOT1 (N13415, N13412);
not NOT1 (N13416, N13395);
or OR2 (N13417, N13402, N6967);
xor XOR2 (N13418, N13408, N4663);
nand NAND3 (N13419, N13375, N10850, N957);
not NOT1 (N13420, N13413);
or OR3 (N13421, N13418, N13295, N4676);
or OR4 (N13422, N13421, N5100, N846, N8707);
and AND4 (N13423, N13414, N12045, N8303, N11980);
and AND2 (N13424, N13419, N11882);
buf BUF1 (N13425, N13409);
nand NAND3 (N13426, N13420, N7064, N5125);
and AND3 (N13427, N13415, N145, N6136);
xor XOR2 (N13428, N13417, N8516);
not NOT1 (N13429, N13391);
nand NAND4 (N13430, N13405, N10422, N7031, N2303);
nor NOR2 (N13431, N13424, N3627);
buf BUF1 (N13432, N13431);
and AND4 (N13433, N13423, N7915, N714, N8166);
nor NOR2 (N13434, N13430, N10216);
nor NOR2 (N13435, N13425, N12842);
nor NOR4 (N13436, N13435, N6232, N8135, N5282);
and AND3 (N13437, N13422, N7063, N9396);
and AND4 (N13438, N13434, N1501, N3981, N10359);
xor XOR2 (N13439, N13426, N4420);
or OR2 (N13440, N13429, N11528);
or OR3 (N13441, N13436, N2733, N11260);
buf BUF1 (N13442, N13440);
xor XOR2 (N13443, N13432, N10912);
and AND4 (N13444, N13441, N9664, N12860, N11318);
or OR4 (N13445, N13416, N431, N9948, N12602);
nor NOR3 (N13446, N13428, N11158, N2604);
nand NAND2 (N13447, N13445, N2489);
or OR2 (N13448, N13439, N1028);
buf BUF1 (N13449, N13448);
and AND3 (N13450, N13449, N2547, N243);
nand NAND3 (N13451, N13442, N4629, N2760);
not NOT1 (N13452, N13437);
nand NAND3 (N13453, N13427, N6711, N9976);
nor NOR2 (N13454, N13443, N8781);
or OR2 (N13455, N13433, N4259);
and AND3 (N13456, N13438, N11897, N3030);
and AND2 (N13457, N13455, N8889);
nand NAND3 (N13458, N13447, N8927, N12353);
nand NAND2 (N13459, N13446, N12926);
nor NOR4 (N13460, N13459, N8825, N2864, N4100);
nand NAND4 (N13461, N13453, N5314, N6733, N10820);
xor XOR2 (N13462, N13452, N2802);
and AND4 (N13463, N13444, N11129, N2493, N4221);
buf BUF1 (N13464, N13460);
nand NAND3 (N13465, N13457, N2376, N9718);
or OR3 (N13466, N13454, N10655, N6931);
nand NAND4 (N13467, N13462, N2239, N6034, N3663);
xor XOR2 (N13468, N13456, N9516);
not NOT1 (N13469, N13467);
not NOT1 (N13470, N13463);
or OR4 (N13471, N13458, N11037, N1078, N3729);
not NOT1 (N13472, N13466);
or OR3 (N13473, N13470, N4626, N3869);
xor XOR2 (N13474, N13465, N7384);
nor NOR2 (N13475, N13474, N3525);
nand NAND4 (N13476, N13451, N1845, N13344, N8246);
not NOT1 (N13477, N13450);
and AND3 (N13478, N13461, N6686, N4508);
nand NAND3 (N13479, N13478, N8282, N12866);
nand NAND2 (N13480, N13464, N12216);
nand NAND3 (N13481, N13475, N11720, N9710);
xor XOR2 (N13482, N13479, N1653);
nand NAND2 (N13483, N13482, N10579);
or OR3 (N13484, N13483, N10044, N6213);
nand NAND2 (N13485, N13484, N143);
and AND2 (N13486, N13468, N7373);
xor XOR2 (N13487, N13469, N6076);
nand NAND3 (N13488, N13481, N10145, N13247);
or OR4 (N13489, N13486, N6515, N9548, N1825);
not NOT1 (N13490, N13472);
buf BUF1 (N13491, N13488);
xor XOR2 (N13492, N13485, N2657);
or OR2 (N13493, N13480, N2588);
or OR3 (N13494, N13492, N5708, N5201);
xor XOR2 (N13495, N13491, N4048);
buf BUF1 (N13496, N13489);
nor NOR2 (N13497, N13495, N6082);
nand NAND3 (N13498, N13490, N9401, N11638);
nand NAND3 (N13499, N13493, N10553, N7366);
and AND2 (N13500, N13499, N6068);
nor NOR4 (N13501, N13477, N10942, N12964, N7305);
buf BUF1 (N13502, N13487);
xor XOR2 (N13503, N13471, N12122);
or OR3 (N13504, N13502, N13430, N2390);
or OR3 (N13505, N13501, N3717, N5946);
not NOT1 (N13506, N13494);
buf BUF1 (N13507, N13506);
nand NAND2 (N13508, N13497, N11363);
or OR3 (N13509, N13508, N10985, N11709);
nor NOR4 (N13510, N13505, N8233, N1083, N6825);
or OR3 (N13511, N13473, N9676, N6227);
and AND2 (N13512, N13500, N12786);
or OR4 (N13513, N13512, N9848, N5168, N3601);
not NOT1 (N13514, N13509);
or OR2 (N13515, N13498, N10573);
xor XOR2 (N13516, N13511, N1511);
not NOT1 (N13517, N13516);
xor XOR2 (N13518, N13517, N3471);
nor NOR2 (N13519, N13518, N10998);
xor XOR2 (N13520, N13515, N3877);
xor XOR2 (N13521, N13476, N4719);
buf BUF1 (N13522, N13507);
and AND2 (N13523, N13520, N11898);
nand NAND3 (N13524, N13504, N7155, N4687);
or OR2 (N13525, N13523, N981);
buf BUF1 (N13526, N13496);
and AND3 (N13527, N13514, N3739, N10003);
xor XOR2 (N13528, N13510, N9075);
xor XOR2 (N13529, N13519, N9540);
not NOT1 (N13530, N13529);
nor NOR3 (N13531, N13530, N693, N1101);
nor NOR2 (N13532, N13522, N1262);
nor NOR3 (N13533, N13528, N5208, N6081);
not NOT1 (N13534, N13527);
not NOT1 (N13535, N13513);
buf BUF1 (N13536, N13521);
xor XOR2 (N13537, N13503, N4457);
xor XOR2 (N13538, N13524, N411);
nor NOR4 (N13539, N13532, N7695, N6759, N9393);
xor XOR2 (N13540, N13537, N3813);
nor NOR3 (N13541, N13535, N4117, N5995);
nor NOR3 (N13542, N13531, N13393, N3954);
and AND3 (N13543, N13533, N2589, N8098);
nand NAND2 (N13544, N13539, N7020);
and AND2 (N13545, N13542, N4225);
nor NOR2 (N13546, N13541, N8902);
and AND4 (N13547, N13526, N6338, N3884, N4615);
xor XOR2 (N13548, N13538, N3796);
nand NAND3 (N13549, N13547, N7856, N6233);
nand NAND2 (N13550, N13548, N8031);
and AND4 (N13551, N13525, N2347, N7965, N4982);
not NOT1 (N13552, N13534);
xor XOR2 (N13553, N13536, N1933);
or OR4 (N13554, N13550, N700, N3789, N3474);
xor XOR2 (N13555, N13551, N1565);
nand NAND3 (N13556, N13545, N10237, N6780);
and AND2 (N13557, N13543, N8547);
xor XOR2 (N13558, N13556, N3236);
not NOT1 (N13559, N13549);
nand NAND4 (N13560, N13557, N7720, N11225, N9684);
and AND3 (N13561, N13560, N5952, N8913);
nand NAND2 (N13562, N13554, N9813);
and AND2 (N13563, N13559, N7509);
and AND4 (N13564, N13546, N3300, N13179, N116);
buf BUF1 (N13565, N13561);
nand NAND3 (N13566, N13540, N1450, N12250);
nor NOR4 (N13567, N13555, N8124, N4124, N10292);
not NOT1 (N13568, N13567);
xor XOR2 (N13569, N13544, N10894);
not NOT1 (N13570, N13552);
not NOT1 (N13571, N13558);
not NOT1 (N13572, N13565);
nand NAND4 (N13573, N13563, N13115, N6133, N187);
buf BUF1 (N13574, N13553);
not NOT1 (N13575, N13564);
and AND2 (N13576, N13568, N4110);
buf BUF1 (N13577, N13573);
not NOT1 (N13578, N13571);
buf BUF1 (N13579, N13570);
xor XOR2 (N13580, N13566, N1720);
and AND4 (N13581, N13580, N1248, N9630, N9164);
xor XOR2 (N13582, N13576, N4257);
nor NOR4 (N13583, N13577, N157, N11898, N10588);
and AND2 (N13584, N13582, N3803);
buf BUF1 (N13585, N13579);
xor XOR2 (N13586, N13585, N296);
and AND4 (N13587, N13572, N12510, N3835, N7342);
xor XOR2 (N13588, N13587, N1152);
and AND4 (N13589, N13578, N982, N4322, N2228);
nor NOR3 (N13590, N13575, N12259, N6612);
not NOT1 (N13591, N13574);
and AND3 (N13592, N13583, N9823, N10350);
xor XOR2 (N13593, N13589, N6599);
not NOT1 (N13594, N13586);
buf BUF1 (N13595, N13569);
nor NOR4 (N13596, N13581, N4294, N11424, N744);
nor NOR2 (N13597, N13596, N1751);
buf BUF1 (N13598, N13588);
and AND3 (N13599, N13598, N7290, N8580);
and AND3 (N13600, N13594, N8211, N1432);
nor NOR2 (N13601, N13584, N7104);
nand NAND4 (N13602, N13592, N8755, N10006, N13377);
or OR3 (N13603, N13601, N2233, N7021);
nor NOR4 (N13604, N13591, N6699, N7570, N1327);
or OR4 (N13605, N13604, N153, N1649, N11326);
nand NAND4 (N13606, N13590, N9045, N9720, N7164);
nand NAND4 (N13607, N13606, N4722, N5589, N12828);
buf BUF1 (N13608, N13605);
nor NOR4 (N13609, N13599, N5456, N6586, N6154);
xor XOR2 (N13610, N13600, N12054);
and AND2 (N13611, N13597, N5361);
xor XOR2 (N13612, N13595, N3170);
nor NOR3 (N13613, N13593, N10843, N11237);
nand NAND4 (N13614, N13613, N9900, N156, N6);
nor NOR2 (N13615, N13562, N742);
nand NAND4 (N13616, N13609, N5700, N13178, N7070);
xor XOR2 (N13617, N13614, N6120);
nor NOR3 (N13618, N13607, N2714, N4966);
not NOT1 (N13619, N13616);
buf BUF1 (N13620, N13608);
nand NAND4 (N13621, N13612, N788, N4517, N7481);
nor NOR2 (N13622, N13621, N603);
nor NOR3 (N13623, N13610, N128, N2483);
and AND4 (N13624, N13615, N8024, N12722, N110);
or OR2 (N13625, N13624, N2875);
not NOT1 (N13626, N13611);
not NOT1 (N13627, N13619);
nor NOR3 (N13628, N13625, N8785, N1061);
xor XOR2 (N13629, N13618, N8166);
not NOT1 (N13630, N13602);
or OR3 (N13631, N13628, N13205, N4713);
buf BUF1 (N13632, N13627);
nor NOR2 (N13633, N13623, N499);
xor XOR2 (N13634, N13617, N1355);
xor XOR2 (N13635, N13633, N9095);
not NOT1 (N13636, N13622);
xor XOR2 (N13637, N13603, N2552);
buf BUF1 (N13638, N13626);
or OR4 (N13639, N13620, N5974, N1963, N2436);
nand NAND3 (N13640, N13635, N7789, N220);
not NOT1 (N13641, N13640);
or OR4 (N13642, N13631, N11333, N830, N56);
and AND2 (N13643, N13639, N11026);
and AND4 (N13644, N13641, N3328, N11477, N5510);
and AND4 (N13645, N13642, N12643, N5802, N4060);
nor NOR2 (N13646, N13630, N5068);
nor NOR3 (N13647, N13634, N2995, N13086);
buf BUF1 (N13648, N13638);
and AND3 (N13649, N13637, N3400, N8289);
nor NOR4 (N13650, N13648, N9683, N11884, N6189);
not NOT1 (N13651, N13636);
and AND4 (N13652, N13629, N11141, N35, N8200);
and AND2 (N13653, N13643, N5769);
nor NOR4 (N13654, N13651, N9398, N6335, N8772);
buf BUF1 (N13655, N13652);
buf BUF1 (N13656, N13654);
nor NOR4 (N13657, N13655, N12515, N3522, N12654);
not NOT1 (N13658, N13653);
and AND3 (N13659, N13656, N5266, N316);
and AND4 (N13660, N13647, N6668, N13540, N5145);
or OR2 (N13661, N13632, N9072);
buf BUF1 (N13662, N13658);
nand NAND3 (N13663, N13650, N9574, N1611);
nand NAND3 (N13664, N13645, N5963, N1906);
buf BUF1 (N13665, N13664);
not NOT1 (N13666, N13660);
xor XOR2 (N13667, N13665, N2392);
and AND4 (N13668, N13646, N3240, N4569, N860);
not NOT1 (N13669, N13666);
buf BUF1 (N13670, N13669);
nor NOR2 (N13671, N13670, N9813);
nand NAND2 (N13672, N13667, N8843);
nand NAND4 (N13673, N13671, N2365, N10377, N7469);
or OR4 (N13674, N13649, N8429, N7874, N9738);
nand NAND3 (N13675, N13661, N8906, N6865);
and AND4 (N13676, N13673, N457, N9816, N4876);
xor XOR2 (N13677, N13657, N7850);
or OR2 (N13678, N13677, N990);
buf BUF1 (N13679, N13676);
not NOT1 (N13680, N13662);
nor NOR3 (N13681, N13678, N12487, N204);
xor XOR2 (N13682, N13680, N2758);
xor XOR2 (N13683, N13681, N7046);
buf BUF1 (N13684, N13672);
and AND2 (N13685, N13684, N12828);
not NOT1 (N13686, N13663);
or OR3 (N13687, N13668, N9785, N989);
nand NAND4 (N13688, N13682, N11439, N627, N13100);
nor NOR3 (N13689, N13687, N9431, N8427);
nor NOR2 (N13690, N13674, N10961);
or OR4 (N13691, N13683, N10889, N4953, N10857);
and AND4 (N13692, N13679, N6454, N3014, N2374);
and AND3 (N13693, N13689, N8315, N13448);
and AND3 (N13694, N13644, N1382, N9669);
not NOT1 (N13695, N13685);
nor NOR3 (N13696, N13695, N11658, N5912);
nor NOR2 (N13697, N13692, N10884);
not NOT1 (N13698, N13691);
xor XOR2 (N13699, N13675, N452);
nand NAND4 (N13700, N13699, N11857, N492, N1948);
and AND3 (N13701, N13688, N5213, N1670);
xor XOR2 (N13702, N13693, N2715);
or OR2 (N13703, N13686, N11674);
xor XOR2 (N13704, N13700, N9640);
nor NOR3 (N13705, N13703, N10594, N13472);
nor NOR3 (N13706, N13704, N7439, N9439);
buf BUF1 (N13707, N13697);
nand NAND3 (N13708, N13702, N1901, N2678);
nand NAND3 (N13709, N13701, N3106, N11204);
nand NAND2 (N13710, N13706, N10194);
xor XOR2 (N13711, N13707, N4645);
xor XOR2 (N13712, N13708, N10106);
buf BUF1 (N13713, N13698);
not NOT1 (N13714, N13709);
or OR3 (N13715, N13712, N215, N3283);
not NOT1 (N13716, N13705);
buf BUF1 (N13717, N13711);
and AND4 (N13718, N13713, N5077, N2802, N6284);
not NOT1 (N13719, N13690);
buf BUF1 (N13720, N13694);
or OR2 (N13721, N13714, N5799);
and AND2 (N13722, N13719, N6151);
nor NOR3 (N13723, N13715, N4553, N2178);
nor NOR2 (N13724, N13723, N8743);
and AND3 (N13725, N13710, N9351, N5864);
and AND4 (N13726, N13724, N3443, N5332, N3336);
nor NOR3 (N13727, N13726, N1466, N5189);
and AND4 (N13728, N13721, N3148, N6953, N4747);
and AND2 (N13729, N13717, N12410);
xor XOR2 (N13730, N13722, N13071);
not NOT1 (N13731, N13728);
not NOT1 (N13732, N13727);
nand NAND4 (N13733, N13725, N9087, N1401, N3761);
xor XOR2 (N13734, N13730, N2886);
or OR4 (N13735, N13734, N5728, N12950, N791);
not NOT1 (N13736, N13731);
or OR2 (N13737, N13733, N4556);
buf BUF1 (N13738, N13659);
nand NAND3 (N13739, N13735, N3022, N11289);
not NOT1 (N13740, N13739);
or OR3 (N13741, N13696, N5453, N12452);
not NOT1 (N13742, N13740);
buf BUF1 (N13743, N13737);
and AND4 (N13744, N13742, N986, N13326, N260);
and AND4 (N13745, N13743, N163, N5122, N9629);
not NOT1 (N13746, N13741);
and AND3 (N13747, N13729, N8599, N9782);
nand NAND4 (N13748, N13732, N7097, N13720, N10781);
nor NOR3 (N13749, N5851, N5965, N3565);
nor NOR4 (N13750, N13749, N11497, N7517, N8485);
nor NOR3 (N13751, N13716, N3060, N9757);
and AND3 (N13752, N13747, N9942, N990);
or OR3 (N13753, N13718, N11194, N4493);
nand NAND4 (N13754, N13736, N11233, N9929, N13640);
nor NOR2 (N13755, N13746, N12887);
and AND4 (N13756, N13738, N2770, N3202, N86);
not NOT1 (N13757, N13756);
nand NAND3 (N13758, N13745, N11887, N3792);
nor NOR3 (N13759, N13752, N7115, N3292);
buf BUF1 (N13760, N13755);
buf BUF1 (N13761, N13759);
nor NOR4 (N13762, N13754, N1108, N6613, N12127);
or OR2 (N13763, N13762, N8425);
nor NOR3 (N13764, N13763, N10001, N124);
nor NOR3 (N13765, N13753, N6856, N3821);
and AND3 (N13766, N13765, N990, N12812);
buf BUF1 (N13767, N13744);
nand NAND2 (N13768, N13766, N1504);
or OR3 (N13769, N13748, N8033, N11836);
buf BUF1 (N13770, N13769);
not NOT1 (N13771, N13757);
and AND3 (N13772, N13767, N10474, N4929);
xor XOR2 (N13773, N13768, N99);
nor NOR4 (N13774, N13761, N244, N4026, N13199);
nor NOR2 (N13775, N13772, N12707);
buf BUF1 (N13776, N13771);
nand NAND2 (N13777, N13764, N11650);
nand NAND4 (N13778, N13758, N12315, N6895, N3027);
buf BUF1 (N13779, N13774);
and AND2 (N13780, N13775, N840);
and AND3 (N13781, N13751, N9889, N12995);
not NOT1 (N13782, N13777);
and AND2 (N13783, N13750, N8036);
and AND3 (N13784, N13782, N4003, N5321);
or OR3 (N13785, N13776, N9066, N523);
not NOT1 (N13786, N13784);
not NOT1 (N13787, N13779);
xor XOR2 (N13788, N13770, N1309);
or OR2 (N13789, N13781, N11332);
nand NAND3 (N13790, N13780, N12283, N2601);
buf BUF1 (N13791, N13786);
and AND3 (N13792, N13789, N12738, N6193);
xor XOR2 (N13793, N13788, N10308);
nor NOR2 (N13794, N13791, N5825);
nand NAND4 (N13795, N13773, N13321, N6500, N4022);
and AND4 (N13796, N13794, N11522, N3054, N12666);
nand NAND2 (N13797, N13796, N8693);
buf BUF1 (N13798, N13778);
nand NAND3 (N13799, N13790, N3096, N6329);
nor NOR3 (N13800, N13795, N4260, N9252);
xor XOR2 (N13801, N13797, N5639);
nor NOR2 (N13802, N13787, N13014);
and AND2 (N13803, N13802, N9493);
and AND4 (N13804, N13783, N12769, N8523, N11013);
not NOT1 (N13805, N13793);
or OR3 (N13806, N13760, N806, N9668);
buf BUF1 (N13807, N13798);
and AND2 (N13808, N13806, N239);
not NOT1 (N13809, N13803);
buf BUF1 (N13810, N13808);
not NOT1 (N13811, N13785);
and AND2 (N13812, N13811, N12101);
not NOT1 (N13813, N13809);
and AND2 (N13814, N13792, N13114);
nor NOR4 (N13815, N13801, N5080, N7058, N13054);
xor XOR2 (N13816, N13812, N793);
xor XOR2 (N13817, N13814, N10477);
nor NOR3 (N13818, N13799, N11996, N9112);
not NOT1 (N13819, N13807);
or OR2 (N13820, N13815, N13073);
nand NAND4 (N13821, N13804, N12296, N5581, N12465);
and AND2 (N13822, N13817, N11904);
or OR4 (N13823, N13820, N13589, N13504, N2606);
nor NOR4 (N13824, N13819, N6746, N12161, N9386);
nor NOR4 (N13825, N13810, N3473, N2085, N7033);
nand NAND4 (N13826, N13818, N244, N7738, N5963);
and AND2 (N13827, N13825, N12979);
not NOT1 (N13828, N13827);
and AND3 (N13829, N13805, N12914, N322);
nand NAND4 (N13830, N13828, N1014, N9775, N6252);
buf BUF1 (N13831, N13816);
nand NAND3 (N13832, N13830, N6868, N5001);
xor XOR2 (N13833, N13813, N5635);
or OR3 (N13834, N13821, N12671, N5433);
and AND2 (N13835, N13831, N4689);
buf BUF1 (N13836, N13824);
nand NAND3 (N13837, N13826, N11767, N11432);
xor XOR2 (N13838, N13834, N3786);
not NOT1 (N13839, N13837);
not NOT1 (N13840, N13823);
nand NAND4 (N13841, N13839, N1210, N6167, N5626);
not NOT1 (N13842, N13838);
or OR4 (N13843, N13835, N3670, N11733, N12163);
or OR2 (N13844, N13833, N9294);
or OR2 (N13845, N13822, N12774);
nand NAND4 (N13846, N13845, N8219, N9688, N10349);
nor NOR3 (N13847, N13829, N4264, N8428);
not NOT1 (N13848, N13832);
xor XOR2 (N13849, N13843, N4883);
nor NOR3 (N13850, N13849, N2052, N2495);
nor NOR2 (N13851, N13842, N7957);
and AND2 (N13852, N13848, N5780);
or OR4 (N13853, N13800, N12767, N10850, N12818);
or OR3 (N13854, N13850, N11221, N12012);
nand NAND4 (N13855, N13841, N11874, N8798, N4229);
not NOT1 (N13856, N13847);
xor XOR2 (N13857, N13851, N13375);
not NOT1 (N13858, N13844);
and AND4 (N13859, N13846, N7195, N1090, N6497);
or OR3 (N13860, N13852, N12210, N8758);
nor NOR2 (N13861, N13857, N6054);
buf BUF1 (N13862, N13861);
nand NAND3 (N13863, N13855, N9141, N6669);
not NOT1 (N13864, N13856);
and AND2 (N13865, N13864, N1266);
nand NAND3 (N13866, N13854, N6373, N12391);
not NOT1 (N13867, N13865);
or OR3 (N13868, N13840, N385, N1921);
not NOT1 (N13869, N13859);
buf BUF1 (N13870, N13836);
xor XOR2 (N13871, N13867, N13459);
buf BUF1 (N13872, N13869);
buf BUF1 (N13873, N13853);
or OR3 (N13874, N13863, N13474, N4764);
not NOT1 (N13875, N13874);
and AND4 (N13876, N13862, N10946, N12423, N389);
xor XOR2 (N13877, N13875, N9369);
not NOT1 (N13878, N13871);
nor NOR4 (N13879, N13873, N524, N308, N317);
or OR3 (N13880, N13858, N9017, N13201);
xor XOR2 (N13881, N13870, N11361);
nand NAND3 (N13882, N13866, N5775, N13024);
nor NOR2 (N13883, N13876, N11580);
xor XOR2 (N13884, N13872, N9269);
and AND3 (N13885, N13880, N2978, N1763);
nor NOR4 (N13886, N13881, N3874, N8518, N4483);
and AND3 (N13887, N13884, N12861, N5169);
nand NAND3 (N13888, N13882, N1203, N7874);
nand NAND2 (N13889, N13878, N4226);
or OR4 (N13890, N13860, N225, N4469, N6145);
not NOT1 (N13891, N13883);
xor XOR2 (N13892, N13877, N3136);
buf BUF1 (N13893, N13889);
and AND2 (N13894, N13892, N4611);
nor NOR4 (N13895, N13891, N2997, N8007, N13347);
buf BUF1 (N13896, N13886);
or OR2 (N13897, N13894, N243);
or OR4 (N13898, N13888, N12203, N3863, N12679);
or OR2 (N13899, N13879, N5135);
not NOT1 (N13900, N13896);
xor XOR2 (N13901, N13885, N6068);
nand NAND3 (N13902, N13895, N4735, N6317);
nor NOR3 (N13903, N13898, N11916, N4821);
xor XOR2 (N13904, N13901, N322);
or OR2 (N13905, N13903, N12055);
not NOT1 (N13906, N13897);
nand NAND4 (N13907, N13900, N31, N8156, N11691);
or OR3 (N13908, N13906, N843, N702);
and AND4 (N13909, N13905, N13319, N12704, N1219);
xor XOR2 (N13910, N13868, N11008);
nor NOR3 (N13911, N13909, N13266, N13747);
or OR4 (N13912, N13893, N6384, N11013, N1907);
buf BUF1 (N13913, N13907);
nand NAND3 (N13914, N13902, N10179, N12250);
and AND2 (N13915, N13908, N5055);
xor XOR2 (N13916, N13913, N13622);
buf BUF1 (N13917, N13914);
buf BUF1 (N13918, N13899);
xor XOR2 (N13919, N13904, N13735);
and AND2 (N13920, N13910, N11127);
or OR3 (N13921, N13887, N896, N2793);
nor NOR3 (N13922, N13912, N756, N8961);
nand NAND2 (N13923, N13916, N9638);
or OR2 (N13924, N13890, N8544);
xor XOR2 (N13925, N13923, N5265);
or OR2 (N13926, N13924, N12217);
nor NOR4 (N13927, N13926, N8121, N7117, N10869);
not NOT1 (N13928, N13918);
buf BUF1 (N13929, N13921);
and AND3 (N13930, N13928, N6531, N2504);
or OR2 (N13931, N13927, N4635);
buf BUF1 (N13932, N13915);
nand NAND2 (N13933, N13925, N5444);
nand NAND2 (N13934, N13920, N10961);
not NOT1 (N13935, N13919);
buf BUF1 (N13936, N13929);
nand NAND2 (N13937, N13931, N3443);
nor NOR2 (N13938, N13917, N11311);
and AND2 (N13939, N13922, N6773);
not NOT1 (N13940, N13933);
xor XOR2 (N13941, N13935, N9898);
or OR4 (N13942, N13941, N5445, N590, N10558);
nand NAND2 (N13943, N13937, N1281);
and AND2 (N13944, N13939, N13058);
nand NAND2 (N13945, N13938, N8215);
buf BUF1 (N13946, N13940);
not NOT1 (N13947, N13945);
nor NOR2 (N13948, N13946, N3743);
or OR3 (N13949, N13932, N13794, N13338);
not NOT1 (N13950, N13936);
xor XOR2 (N13951, N13942, N4231);
nand NAND3 (N13952, N13934, N7600, N7090);
xor XOR2 (N13953, N13952, N1762);
nor NOR2 (N13954, N13953, N10908);
and AND3 (N13955, N13911, N6, N11343);
nor NOR2 (N13956, N13951, N9091);
or OR4 (N13957, N13950, N11792, N12083, N8402);
not NOT1 (N13958, N13956);
nor NOR2 (N13959, N13955, N509);
or OR2 (N13960, N13954, N6007);
and AND3 (N13961, N13959, N5482, N11413);
nor NOR4 (N13962, N13957, N6725, N2998, N7883);
or OR4 (N13963, N13961, N7568, N4085, N8032);
xor XOR2 (N13964, N13930, N11734);
nor NOR2 (N13965, N13963, N629);
not NOT1 (N13966, N13947);
buf BUF1 (N13967, N13962);
xor XOR2 (N13968, N13943, N11986);
not NOT1 (N13969, N13944);
or OR2 (N13970, N13968, N7488);
or OR3 (N13971, N13967, N5974, N1074);
xor XOR2 (N13972, N13971, N2411);
buf BUF1 (N13973, N13972);
and AND3 (N13974, N13970, N1472, N8477);
nor NOR2 (N13975, N13965, N13410);
nor NOR2 (N13976, N13966, N5830);
nor NOR3 (N13977, N13969, N4223, N1294);
and AND4 (N13978, N13964, N9257, N9195, N1249);
nand NAND2 (N13979, N13960, N1098);
nand NAND4 (N13980, N13949, N1060, N4250, N6114);
nand NAND2 (N13981, N13976, N11027);
or OR4 (N13982, N13980, N7368, N1311, N360);
or OR3 (N13983, N13948, N8142, N217);
nand NAND3 (N13984, N13983, N1014, N6229);
buf BUF1 (N13985, N13977);
buf BUF1 (N13986, N13974);
nor NOR2 (N13987, N13982, N10538);
and AND3 (N13988, N13986, N3470, N5598);
buf BUF1 (N13989, N13988);
xor XOR2 (N13990, N13978, N1174);
xor XOR2 (N13991, N13981, N9581);
nor NOR2 (N13992, N13990, N12973);
not NOT1 (N13993, N13958);
or OR2 (N13994, N13987, N853);
not NOT1 (N13995, N13979);
not NOT1 (N13996, N13994);
or OR2 (N13997, N13989, N2306);
buf BUF1 (N13998, N13996);
not NOT1 (N13999, N13984);
not NOT1 (N14000, N13999);
or OR4 (N14001, N14000, N9550, N3722, N5557);
xor XOR2 (N14002, N13995, N4323);
xor XOR2 (N14003, N13975, N10004);
nor NOR4 (N14004, N13973, N9767, N9466, N4751);
not NOT1 (N14005, N14001);
nand NAND4 (N14006, N13998, N177, N8634, N8056);
and AND2 (N14007, N14003, N3372);
not NOT1 (N14008, N13997);
and AND4 (N14009, N14008, N5163, N11168, N1814);
buf BUF1 (N14010, N14004);
or OR3 (N14011, N14009, N6168, N3961);
buf BUF1 (N14012, N14010);
xor XOR2 (N14013, N13993, N10397);
or OR2 (N14014, N13985, N9575);
or OR2 (N14015, N13991, N5621);
or OR2 (N14016, N14014, N4806);
buf BUF1 (N14017, N14002);
nor NOR2 (N14018, N14012, N11387);
and AND2 (N14019, N13992, N10274);
not NOT1 (N14020, N14015);
not NOT1 (N14021, N14007);
xor XOR2 (N14022, N14005, N4106);
buf BUF1 (N14023, N14019);
or OR3 (N14024, N14023, N1435, N3801);
nand NAND2 (N14025, N14016, N198);
nor NOR4 (N14026, N14024, N464, N1451, N8285);
or OR2 (N14027, N14025, N12323);
and AND3 (N14028, N14022, N2032, N11618);
buf BUF1 (N14029, N14011);
nor NOR3 (N14030, N14017, N529, N6563);
nor NOR3 (N14031, N14028, N4740, N1372);
nand NAND4 (N14032, N14018, N11756, N11852, N10193);
xor XOR2 (N14033, N14027, N8935);
xor XOR2 (N14034, N14013, N5893);
nand NAND3 (N14035, N14006, N11154, N7953);
nand NAND3 (N14036, N14033, N6748, N9421);
xor XOR2 (N14037, N14030, N10068);
nand NAND2 (N14038, N14020, N510);
not NOT1 (N14039, N14026);
buf BUF1 (N14040, N14034);
and AND2 (N14041, N14040, N12960);
nand NAND2 (N14042, N14037, N9681);
nor NOR3 (N14043, N14029, N10234, N7901);
nand NAND4 (N14044, N14032, N7713, N9581, N1979);
nand NAND3 (N14045, N14035, N1530, N4654);
xor XOR2 (N14046, N14036, N1814);
nor NOR2 (N14047, N14041, N6347);
xor XOR2 (N14048, N14021, N12863);
nand NAND2 (N14049, N14043, N3644);
nor NOR4 (N14050, N14047, N12842, N12269, N6442);
xor XOR2 (N14051, N14039, N220);
nand NAND4 (N14052, N14048, N12759, N1185, N6082);
or OR4 (N14053, N14045, N12343, N4598, N5306);
buf BUF1 (N14054, N14049);
xor XOR2 (N14055, N14054, N4385);
nand NAND3 (N14056, N14052, N2200, N12461);
and AND4 (N14057, N14056, N8605, N10630, N4519);
or OR2 (N14058, N14031, N12533);
buf BUF1 (N14059, N14051);
nor NOR3 (N14060, N14053, N11950, N3308);
not NOT1 (N14061, N14038);
nand NAND4 (N14062, N14058, N10061, N10477, N12947);
xor XOR2 (N14063, N14059, N2939);
xor XOR2 (N14064, N14055, N9576);
xor XOR2 (N14065, N14046, N13731);
or OR2 (N14066, N14061, N7218);
buf BUF1 (N14067, N14044);
nand NAND3 (N14068, N14066, N5368, N12599);
buf BUF1 (N14069, N14060);
not NOT1 (N14070, N14069);
not NOT1 (N14071, N14065);
or OR4 (N14072, N14062, N7066, N2828, N9465);
nor NOR4 (N14073, N14050, N11778, N10667, N7590);
xor XOR2 (N14074, N14067, N4350);
xor XOR2 (N14075, N14073, N6888);
not NOT1 (N14076, N14072);
nor NOR3 (N14077, N14074, N13475, N12663);
or OR2 (N14078, N14076, N9683);
or OR4 (N14079, N14075, N11821, N12001, N13339);
buf BUF1 (N14080, N14079);
nand NAND2 (N14081, N14063, N7128);
not NOT1 (N14082, N14064);
not NOT1 (N14083, N14071);
not NOT1 (N14084, N14078);
or OR2 (N14085, N14077, N6686);
not NOT1 (N14086, N14082);
xor XOR2 (N14087, N14084, N8950);
nand NAND4 (N14088, N14042, N12795, N3951, N13070);
xor XOR2 (N14089, N14086, N2291);
buf BUF1 (N14090, N14088);
not NOT1 (N14091, N14083);
nand NAND3 (N14092, N14057, N12992, N3075);
xor XOR2 (N14093, N14085, N12544);
or OR4 (N14094, N14070, N11042, N10531, N14092);
nor NOR2 (N14095, N10398, N443);
nand NAND3 (N14096, N14081, N4437, N338);
nor NOR2 (N14097, N14068, N234);
and AND3 (N14098, N14097, N7028, N9157);
buf BUF1 (N14099, N14098);
and AND3 (N14100, N14091, N10218, N9130);
xor XOR2 (N14101, N14099, N9593);
not NOT1 (N14102, N14096);
not NOT1 (N14103, N14094);
xor XOR2 (N14104, N14095, N7766);
nand NAND2 (N14105, N14101, N12720);
not NOT1 (N14106, N14089);
buf BUF1 (N14107, N14093);
nor NOR4 (N14108, N14080, N5248, N8649, N2021);
xor XOR2 (N14109, N14106, N11874);
xor XOR2 (N14110, N14100, N3937);
and AND3 (N14111, N14090, N13347, N2065);
and AND2 (N14112, N14109, N13136);
not NOT1 (N14113, N14111);
and AND2 (N14114, N14110, N2829);
nor NOR3 (N14115, N14107, N6774, N588);
nand NAND2 (N14116, N14105, N2105);
xor XOR2 (N14117, N14087, N9385);
nand NAND4 (N14118, N14113, N929, N13343, N12347);
and AND4 (N14119, N14115, N364, N2545, N12544);
xor XOR2 (N14120, N14116, N3145);
or OR3 (N14121, N14102, N6829, N2748);
xor XOR2 (N14122, N14121, N615);
buf BUF1 (N14123, N14112);
not NOT1 (N14124, N14114);
xor XOR2 (N14125, N14118, N3730);
or OR4 (N14126, N14123, N55, N12538, N10089);
buf BUF1 (N14127, N14122);
buf BUF1 (N14128, N14120);
not NOT1 (N14129, N14127);
nand NAND2 (N14130, N14126, N7737);
nor NOR3 (N14131, N14129, N228, N6385);
xor XOR2 (N14132, N14103, N9281);
and AND3 (N14133, N14117, N8899, N8371);
and AND3 (N14134, N14104, N9314, N550);
xor XOR2 (N14135, N14133, N3746);
buf BUF1 (N14136, N14131);
buf BUF1 (N14137, N14130);
nand NAND3 (N14138, N14124, N5432, N3046);
buf BUF1 (N14139, N14136);
buf BUF1 (N14140, N14125);
not NOT1 (N14141, N14135);
nor NOR3 (N14142, N14139, N9476, N2616);
nor NOR2 (N14143, N14138, N13221);
or OR2 (N14144, N14128, N3112);
or OR2 (N14145, N14108, N6256);
and AND2 (N14146, N14145, N6469);
buf BUF1 (N14147, N14141);
and AND4 (N14148, N14147, N12861, N12140, N2481);
buf BUF1 (N14149, N14146);
or OR3 (N14150, N14144, N10686, N4112);
or OR2 (N14151, N14148, N8800);
not NOT1 (N14152, N14149);
or OR4 (N14153, N14134, N1882, N4241, N12415);
and AND4 (N14154, N14152, N12310, N6307, N671);
xor XOR2 (N14155, N14150, N13456);
and AND3 (N14156, N14132, N6422, N11620);
xor XOR2 (N14157, N14153, N6347);
nor NOR3 (N14158, N14142, N5299, N1838);
nand NAND3 (N14159, N14158, N11762, N9574);
nor NOR4 (N14160, N14143, N2847, N4881, N909);
xor XOR2 (N14161, N14119, N7618);
not NOT1 (N14162, N14137);
or OR4 (N14163, N14140, N6827, N5555, N11087);
or OR3 (N14164, N14156, N7408, N5382);
buf BUF1 (N14165, N14155);
nand NAND4 (N14166, N14159, N1374, N505, N10974);
xor XOR2 (N14167, N14162, N4842);
not NOT1 (N14168, N14151);
and AND4 (N14169, N14160, N1482, N14165, N9676);
nand NAND3 (N14170, N11255, N12251, N4931);
nand NAND3 (N14171, N14166, N1343, N2402);
nor NOR2 (N14172, N14157, N8715);
nor NOR2 (N14173, N14169, N6145);
xor XOR2 (N14174, N14167, N7091);
and AND4 (N14175, N14164, N11556, N9808, N12226);
nor NOR3 (N14176, N14168, N9564, N1102);
nor NOR3 (N14177, N14154, N10440, N502);
nor NOR3 (N14178, N14161, N6118, N1719);
or OR3 (N14179, N14163, N2993, N8758);
nand NAND3 (N14180, N14170, N10048, N7567);
nand NAND2 (N14181, N14175, N12893);
xor XOR2 (N14182, N14172, N1537);
nor NOR3 (N14183, N14171, N11812, N6668);
or OR4 (N14184, N14181, N13808, N6438, N2484);
nor NOR4 (N14185, N14173, N11203, N3559, N9482);
and AND3 (N14186, N14179, N12280, N3812);
buf BUF1 (N14187, N14180);
buf BUF1 (N14188, N14176);
xor XOR2 (N14189, N14182, N771);
not NOT1 (N14190, N14187);
xor XOR2 (N14191, N14178, N3836);
buf BUF1 (N14192, N14185);
nand NAND2 (N14193, N14186, N2581);
or OR2 (N14194, N14183, N11221);
or OR3 (N14195, N14177, N3861, N226);
or OR3 (N14196, N14193, N4148, N804);
and AND3 (N14197, N14196, N12944, N884);
buf BUF1 (N14198, N14192);
or OR3 (N14199, N14194, N10600, N9401);
nor NOR4 (N14200, N14198, N4676, N187, N4343);
buf BUF1 (N14201, N14200);
nand NAND3 (N14202, N14174, N9584, N11040);
and AND4 (N14203, N14199, N473, N2026, N2187);
or OR4 (N14204, N14201, N4577, N2570, N10370);
not NOT1 (N14205, N14203);
and AND2 (N14206, N14202, N1649);
nand NAND2 (N14207, N14205, N9711);
buf BUF1 (N14208, N14189);
buf BUF1 (N14209, N14207);
or OR2 (N14210, N14209, N9677);
buf BUF1 (N14211, N14190);
buf BUF1 (N14212, N14197);
nor NOR2 (N14213, N14212, N1684);
not NOT1 (N14214, N14195);
xor XOR2 (N14215, N14214, N9731);
xor XOR2 (N14216, N14215, N7655);
buf BUF1 (N14217, N14206);
or OR4 (N14218, N14216, N7010, N1280, N9189);
xor XOR2 (N14219, N14208, N12050);
nor NOR3 (N14220, N14217, N2834, N12212);
or OR3 (N14221, N14219, N3878, N215);
or OR2 (N14222, N14211, N13759);
xor XOR2 (N14223, N14221, N10815);
nand NAND2 (N14224, N14213, N4298);
buf BUF1 (N14225, N14184);
and AND2 (N14226, N14188, N1169);
not NOT1 (N14227, N14218);
nor NOR3 (N14228, N14225, N4477, N9238);
buf BUF1 (N14229, N14223);
or OR2 (N14230, N14229, N11650);
not NOT1 (N14231, N14222);
xor XOR2 (N14232, N14210, N10867);
buf BUF1 (N14233, N14230);
nand NAND3 (N14234, N14224, N12018, N13467);
xor XOR2 (N14235, N14227, N13187);
not NOT1 (N14236, N14235);
and AND4 (N14237, N14236, N9418, N11375, N5572);
or OR4 (N14238, N14191, N3300, N9985, N12592);
and AND4 (N14239, N14226, N2083, N4974, N4010);
nand NAND4 (N14240, N14238, N2655, N10291, N1566);
and AND3 (N14241, N14240, N6425, N4412);
xor XOR2 (N14242, N14231, N14042);
xor XOR2 (N14243, N14228, N7552);
nand NAND2 (N14244, N14220, N11840);
or OR3 (N14245, N14233, N11059, N669);
nor NOR3 (N14246, N14245, N7678, N1727);
not NOT1 (N14247, N14239);
xor XOR2 (N14248, N14246, N2140);
not NOT1 (N14249, N14247);
buf BUF1 (N14250, N14237);
not NOT1 (N14251, N14242);
buf BUF1 (N14252, N14232);
buf BUF1 (N14253, N14250);
not NOT1 (N14254, N14251);
or OR3 (N14255, N14234, N2508, N9869);
and AND3 (N14256, N14204, N11410, N3418);
nor NOR2 (N14257, N14248, N7585);
nor NOR4 (N14258, N14244, N12682, N3424, N4322);
not NOT1 (N14259, N14253);
not NOT1 (N14260, N14252);
nand NAND3 (N14261, N14255, N9399, N5409);
buf BUF1 (N14262, N14259);
not NOT1 (N14263, N14254);
or OR2 (N14264, N14261, N8411);
buf BUF1 (N14265, N14258);
nor NOR4 (N14266, N14249, N9943, N10018, N6323);
not NOT1 (N14267, N14266);
and AND2 (N14268, N14267, N7989);
xor XOR2 (N14269, N14268, N6576);
xor XOR2 (N14270, N14262, N7366);
buf BUF1 (N14271, N14263);
buf BUF1 (N14272, N14269);
nand NAND4 (N14273, N14241, N1566, N8814, N1636);
and AND4 (N14274, N14264, N3070, N514, N1196);
buf BUF1 (N14275, N14257);
or OR2 (N14276, N14272, N10052);
xor XOR2 (N14277, N14270, N9334);
nand NAND3 (N14278, N14276, N13643, N8937);
nor NOR3 (N14279, N14278, N895, N6151);
nor NOR4 (N14280, N14265, N10395, N3498, N8009);
buf BUF1 (N14281, N14271);
or OR4 (N14282, N14274, N2822, N11128, N710);
not NOT1 (N14283, N14277);
nor NOR2 (N14284, N14283, N7633);
not NOT1 (N14285, N14273);
or OR4 (N14286, N14281, N2279, N7017, N7913);
buf BUF1 (N14287, N14260);
not NOT1 (N14288, N14243);
buf BUF1 (N14289, N14286);
buf BUF1 (N14290, N14279);
nand NAND3 (N14291, N14288, N1272, N8105);
nand NAND3 (N14292, N14282, N6908, N905);
not NOT1 (N14293, N14289);
and AND3 (N14294, N14293, N3144, N2821);
nand NAND2 (N14295, N14280, N8428);
buf BUF1 (N14296, N14295);
buf BUF1 (N14297, N14256);
not NOT1 (N14298, N14275);
not NOT1 (N14299, N14298);
or OR2 (N14300, N14296, N11381);
and AND3 (N14301, N14290, N4308, N13032);
nor NOR3 (N14302, N14297, N9814, N6223);
not NOT1 (N14303, N14300);
nor NOR3 (N14304, N14303, N9370, N4535);
and AND2 (N14305, N14292, N12391);
buf BUF1 (N14306, N14299);
nand NAND2 (N14307, N14304, N13364);
or OR2 (N14308, N14301, N10309);
nand NAND2 (N14309, N14305, N10081);
or OR2 (N14310, N14306, N9829);
xor XOR2 (N14311, N14307, N1963);
and AND3 (N14312, N14308, N8571, N6802);
or OR4 (N14313, N14285, N1528, N11532, N2737);
buf BUF1 (N14314, N14309);
xor XOR2 (N14315, N14311, N1123);
nor NOR2 (N14316, N14291, N1982);
nor NOR3 (N14317, N14302, N461, N696);
or OR3 (N14318, N14284, N8345, N2728);
not NOT1 (N14319, N14317);
and AND4 (N14320, N14318, N2828, N7158, N7948);
or OR2 (N14321, N14294, N4948);
nor NOR4 (N14322, N14319, N12110, N2285, N6442);
nand NAND2 (N14323, N14320, N2281);
not NOT1 (N14324, N14314);
nand NAND4 (N14325, N14312, N11856, N10649, N5551);
nand NAND3 (N14326, N14310, N5379, N11011);
and AND2 (N14327, N14316, N9557);
and AND4 (N14328, N14324, N4982, N7417, N3056);
nand NAND4 (N14329, N14322, N1092, N3251, N5373);
or OR3 (N14330, N14327, N7462, N9933);
not NOT1 (N14331, N14321);
or OR4 (N14332, N14329, N106, N13588, N12191);
nand NAND2 (N14333, N14315, N6195);
nor NOR4 (N14334, N14323, N7162, N2234, N7573);
nand NAND2 (N14335, N14287, N1654);
nor NOR3 (N14336, N14333, N9995, N6964);
and AND3 (N14337, N14328, N248, N4053);
xor XOR2 (N14338, N14335, N5430);
not NOT1 (N14339, N14313);
nor NOR4 (N14340, N14332, N5535, N7712, N1816);
nand NAND4 (N14341, N14330, N9349, N9132, N9084);
xor XOR2 (N14342, N14341, N5253);
xor XOR2 (N14343, N14326, N12907);
nand NAND2 (N14344, N14337, N7984);
nor NOR4 (N14345, N14331, N6930, N12426, N10300);
xor XOR2 (N14346, N14342, N7483);
nand NAND4 (N14347, N14345, N6304, N10350, N3094);
nand NAND2 (N14348, N14339, N11013);
nand NAND4 (N14349, N14340, N4314, N9873, N2056);
or OR2 (N14350, N14349, N12971);
and AND4 (N14351, N14347, N3461, N13291, N7388);
not NOT1 (N14352, N14334);
or OR2 (N14353, N14336, N12300);
nand NAND4 (N14354, N14343, N2515, N8347, N6838);
nor NOR4 (N14355, N14351, N13340, N12222, N5053);
not NOT1 (N14356, N14352);
nor NOR3 (N14357, N14355, N1133, N785);
nor NOR2 (N14358, N14338, N7448);
or OR4 (N14359, N14354, N13346, N6764, N8330);
or OR2 (N14360, N14359, N13231);
and AND2 (N14361, N14358, N5621);
not NOT1 (N14362, N14348);
buf BUF1 (N14363, N14357);
or OR2 (N14364, N14361, N8950);
or OR3 (N14365, N14364, N12333, N10998);
buf BUF1 (N14366, N14353);
nand NAND2 (N14367, N14344, N10014);
not NOT1 (N14368, N14363);
xor XOR2 (N14369, N14350, N6543);
buf BUF1 (N14370, N14346);
and AND3 (N14371, N14367, N7064, N12673);
or OR3 (N14372, N14360, N5252, N9050);
and AND4 (N14373, N14372, N5030, N11782, N3488);
or OR2 (N14374, N14371, N4416);
or OR4 (N14375, N14366, N11896, N12257, N10757);
and AND3 (N14376, N14369, N4679, N6297);
or OR3 (N14377, N14373, N29, N1198);
nand NAND3 (N14378, N14325, N2472, N9712);
xor XOR2 (N14379, N14368, N13982);
nand NAND2 (N14380, N14356, N13038);
or OR2 (N14381, N14374, N8992);
and AND2 (N14382, N14378, N59);
and AND4 (N14383, N14370, N12287, N3041, N3420);
nor NOR3 (N14384, N14376, N14003, N6596);
and AND4 (N14385, N14365, N12805, N4922, N8224);
xor XOR2 (N14386, N14383, N10412);
not NOT1 (N14387, N14380);
not NOT1 (N14388, N14385);
not NOT1 (N14389, N14381);
nor NOR2 (N14390, N14388, N645);
buf BUF1 (N14391, N14389);
xor XOR2 (N14392, N14384, N10847);
nor NOR4 (N14393, N14386, N2837, N6132, N2115);
or OR4 (N14394, N14379, N6388, N7983, N4918);
or OR2 (N14395, N14392, N8037);
not NOT1 (N14396, N14393);
nor NOR2 (N14397, N14396, N11900);
and AND4 (N14398, N14382, N12072, N5365, N11660);
and AND2 (N14399, N14391, N13055);
xor XOR2 (N14400, N14362, N965);
or OR4 (N14401, N14397, N2253, N3963, N2115);
not NOT1 (N14402, N14401);
nand NAND3 (N14403, N14398, N5216, N1391);
or OR3 (N14404, N14375, N3100, N1653);
buf BUF1 (N14405, N14395);
nor NOR2 (N14406, N14387, N43);
nand NAND4 (N14407, N14404, N3504, N1883, N519);
buf BUF1 (N14408, N14405);
buf BUF1 (N14409, N14402);
and AND2 (N14410, N14390, N13245);
nor NOR2 (N14411, N14399, N9100);
nand NAND3 (N14412, N14406, N48, N10139);
and AND2 (N14413, N14411, N11824);
nor NOR4 (N14414, N14377, N4198, N126, N22);
not NOT1 (N14415, N14413);
xor XOR2 (N14416, N14415, N3966);
and AND2 (N14417, N14407, N10981);
xor XOR2 (N14418, N14412, N11527);
nand NAND3 (N14419, N14418, N4508, N2289);
and AND4 (N14420, N14410, N11639, N3154, N2211);
nor NOR3 (N14421, N14419, N11246, N7833);
or OR3 (N14422, N14409, N8955, N1226);
or OR2 (N14423, N14422, N7448);
xor XOR2 (N14424, N14414, N2989);
and AND4 (N14425, N14416, N12515, N14350, N12378);
nor NOR4 (N14426, N14423, N11752, N5722, N654);
not NOT1 (N14427, N14425);
xor XOR2 (N14428, N14417, N2755);
nor NOR4 (N14429, N14394, N7309, N7252, N6917);
nor NOR3 (N14430, N14427, N5734, N14213);
or OR4 (N14431, N14430, N12, N8499, N3600);
or OR2 (N14432, N14420, N11201);
buf BUF1 (N14433, N14408);
or OR3 (N14434, N14426, N8933, N7850);
buf BUF1 (N14435, N14421);
or OR4 (N14436, N14428, N8063, N7813, N3036);
and AND2 (N14437, N14435, N5116);
xor XOR2 (N14438, N14432, N7234);
nor NOR3 (N14439, N14403, N3998, N7175);
not NOT1 (N14440, N14434);
or OR4 (N14441, N14438, N10475, N14198, N13931);
or OR4 (N14442, N14436, N6325, N1253, N9753);
and AND2 (N14443, N14441, N14109);
not NOT1 (N14444, N14424);
not NOT1 (N14445, N14400);
or OR2 (N14446, N14444, N5657);
or OR2 (N14447, N14442, N14313);
buf BUF1 (N14448, N14439);
xor XOR2 (N14449, N14446, N1658);
or OR2 (N14450, N14437, N10600);
or OR2 (N14451, N14445, N2262);
not NOT1 (N14452, N14449);
nor NOR2 (N14453, N14447, N3520);
and AND3 (N14454, N14433, N9325, N6896);
xor XOR2 (N14455, N14440, N4797);
nor NOR4 (N14456, N14429, N1954, N4150, N14261);
or OR2 (N14457, N14431, N778);
nand NAND4 (N14458, N14456, N3367, N3772, N10796);
and AND2 (N14459, N14451, N7327);
nand NAND2 (N14460, N14455, N14127);
not NOT1 (N14461, N14457);
nand NAND4 (N14462, N14454, N6463, N11229, N2653);
buf BUF1 (N14463, N14459);
not NOT1 (N14464, N14461);
or OR3 (N14465, N14452, N2151, N10503);
xor XOR2 (N14466, N14460, N13151);
buf BUF1 (N14467, N14466);
not NOT1 (N14468, N14464);
buf BUF1 (N14469, N14465);
not NOT1 (N14470, N14453);
and AND3 (N14471, N14467, N11753, N7259);
not NOT1 (N14472, N14448);
xor XOR2 (N14473, N14450, N804);
nor NOR4 (N14474, N14469, N6865, N9288, N1567);
not NOT1 (N14475, N14470);
buf BUF1 (N14476, N14463);
nand NAND4 (N14477, N14476, N1725, N12632, N3213);
nand NAND4 (N14478, N14458, N13211, N8360, N10373);
xor XOR2 (N14479, N14474, N11927);
or OR2 (N14480, N14477, N5297);
nor NOR4 (N14481, N14475, N5593, N13588, N12185);
or OR2 (N14482, N14472, N10350);
nand NAND3 (N14483, N14478, N7375, N11215);
nand NAND4 (N14484, N14443, N12861, N4303, N5811);
and AND4 (N14485, N14471, N5788, N6496, N3845);
not NOT1 (N14486, N14484);
nor NOR3 (N14487, N14483, N6412, N10581);
and AND2 (N14488, N14486, N773);
nor NOR4 (N14489, N14487, N7436, N8188, N7579);
nor NOR4 (N14490, N14480, N7295, N5860, N10099);
not NOT1 (N14491, N14468);
and AND4 (N14492, N14491, N5450, N8695, N5984);
nand NAND2 (N14493, N14492, N8604);
buf BUF1 (N14494, N14473);
nand NAND2 (N14495, N14462, N11309);
nand NAND3 (N14496, N14481, N9293, N14032);
not NOT1 (N14497, N14489);
nor NOR2 (N14498, N14495, N7709);
nand NAND2 (N14499, N14488, N11039);
not NOT1 (N14500, N14496);
xor XOR2 (N14501, N14479, N7527);
buf BUF1 (N14502, N14493);
xor XOR2 (N14503, N14482, N3830);
buf BUF1 (N14504, N14503);
not NOT1 (N14505, N14490);
not NOT1 (N14506, N14502);
or OR4 (N14507, N14501, N11090, N2798, N4981);
nor NOR3 (N14508, N14500, N7985, N1381);
nand NAND3 (N14509, N14508, N12342, N10878);
xor XOR2 (N14510, N14504, N4041);
xor XOR2 (N14511, N14498, N10629);
and AND4 (N14512, N14511, N2368, N5856, N9522);
nor NOR2 (N14513, N14505, N12567);
not NOT1 (N14514, N14512);
xor XOR2 (N14515, N14514, N317);
not NOT1 (N14516, N14506);
nand NAND3 (N14517, N14507, N2454, N8728);
nand NAND2 (N14518, N14485, N9316);
nand NAND3 (N14519, N14518, N5389, N3857);
nand NAND2 (N14520, N14519, N10806);
nand NAND4 (N14521, N14516, N8863, N9913, N9435);
or OR3 (N14522, N14497, N9039, N12913);
and AND3 (N14523, N14494, N5221, N1508);
not NOT1 (N14524, N14517);
nor NOR4 (N14525, N14524, N13413, N937, N2689);
nor NOR3 (N14526, N14520, N4591, N5354);
and AND2 (N14527, N14522, N3672);
not NOT1 (N14528, N14525);
buf BUF1 (N14529, N14523);
xor XOR2 (N14530, N14509, N1827);
xor XOR2 (N14531, N14513, N11121);
not NOT1 (N14532, N14530);
and AND4 (N14533, N14515, N11226, N4294, N12444);
or OR2 (N14534, N14533, N114);
and AND2 (N14535, N14532, N2847);
buf BUF1 (N14536, N14526);
buf BUF1 (N14537, N14528);
and AND4 (N14538, N14510, N6916, N10318, N7641);
and AND2 (N14539, N14527, N10412);
buf BUF1 (N14540, N14538);
xor XOR2 (N14541, N14537, N2612);
buf BUF1 (N14542, N14499);
nand NAND2 (N14543, N14539, N7259);
buf BUF1 (N14544, N14534);
and AND2 (N14545, N14536, N5748);
xor XOR2 (N14546, N14531, N6682);
buf BUF1 (N14547, N14521);
nand NAND3 (N14548, N14535, N2668, N2314);
buf BUF1 (N14549, N14545);
nor NOR4 (N14550, N14549, N4392, N8580, N13537);
xor XOR2 (N14551, N14550, N3440);
nand NAND2 (N14552, N14548, N404);
not NOT1 (N14553, N14544);
buf BUF1 (N14554, N14542);
and AND2 (N14555, N14547, N14274);
buf BUF1 (N14556, N14529);
xor XOR2 (N14557, N14554, N5921);
not NOT1 (N14558, N14543);
nor NOR4 (N14559, N14555, N14015, N1614, N767);
xor XOR2 (N14560, N14553, N8997);
nor NOR4 (N14561, N14559, N6255, N3943, N9850);
xor XOR2 (N14562, N14560, N1304);
and AND3 (N14563, N14551, N2713, N3999);
and AND4 (N14564, N14541, N14156, N4416, N11894);
and AND4 (N14565, N14556, N8199, N11629, N9025);
or OR3 (N14566, N14562, N7152, N3578);
not NOT1 (N14567, N14552);
not NOT1 (N14568, N14558);
nor NOR2 (N14569, N14540, N5638);
buf BUF1 (N14570, N14566);
and AND2 (N14571, N14569, N9407);
not NOT1 (N14572, N14561);
xor XOR2 (N14573, N14564, N6680);
and AND3 (N14574, N14567, N12908, N6724);
or OR4 (N14575, N14574, N6290, N8899, N7668);
xor XOR2 (N14576, N14568, N685);
nand NAND4 (N14577, N14575, N10949, N410, N13943);
nor NOR2 (N14578, N14571, N14008);
not NOT1 (N14579, N14557);
or OR4 (N14580, N14573, N1721, N10312, N5833);
nand NAND2 (N14581, N14579, N8844);
nor NOR3 (N14582, N14580, N93, N1366);
and AND3 (N14583, N14581, N11895, N995);
buf BUF1 (N14584, N14576);
nor NOR3 (N14585, N14583, N1495, N5136);
nand NAND4 (N14586, N14565, N5439, N10910, N13683);
nand NAND4 (N14587, N14570, N12656, N7010, N8986);
nand NAND2 (N14588, N14582, N1427);
xor XOR2 (N14589, N14584, N13710);
buf BUF1 (N14590, N14577);
or OR4 (N14591, N14586, N3511, N10238, N710);
or OR4 (N14592, N14585, N10215, N14447, N7988);
nand NAND2 (N14593, N14589, N3224);
and AND3 (N14594, N14587, N11411, N1815);
xor XOR2 (N14595, N14592, N3136);
and AND4 (N14596, N14578, N5706, N1138, N12615);
nand NAND4 (N14597, N14563, N2608, N14463, N1480);
nor NOR3 (N14598, N14546, N555, N1254);
or OR2 (N14599, N14594, N9830);
buf BUF1 (N14600, N14597);
xor XOR2 (N14601, N14595, N6667);
nand NAND3 (N14602, N14601, N7265, N10849);
or OR2 (N14603, N14591, N12621);
nand NAND4 (N14604, N14603, N8047, N10757, N13368);
buf BUF1 (N14605, N14593);
buf BUF1 (N14606, N14590);
nand NAND4 (N14607, N14588, N995, N11002, N12711);
or OR2 (N14608, N14596, N4749);
nor NOR3 (N14609, N14608, N9450, N7209);
and AND2 (N14610, N14599, N2680);
and AND2 (N14611, N14610, N745);
not NOT1 (N14612, N14605);
xor XOR2 (N14613, N14606, N3842);
buf BUF1 (N14614, N14613);
or OR4 (N14615, N14607, N2421, N14086, N7222);
nor NOR4 (N14616, N14611, N6393, N5790, N6629);
or OR3 (N14617, N14615, N1373, N11957);
nor NOR4 (N14618, N14609, N1528, N500, N10908);
xor XOR2 (N14619, N14598, N9183);
and AND2 (N14620, N14619, N12541);
buf BUF1 (N14621, N14600);
nand NAND4 (N14622, N14604, N662, N13772, N4620);
xor XOR2 (N14623, N14622, N12401);
not NOT1 (N14624, N14617);
or OR4 (N14625, N14572, N12917, N916, N7610);
or OR2 (N14626, N14623, N3322);
or OR3 (N14627, N14602, N9449, N9757);
not NOT1 (N14628, N14612);
and AND2 (N14629, N14627, N5747);
not NOT1 (N14630, N14625);
and AND4 (N14631, N14629, N1013, N7381, N1409);
nor NOR3 (N14632, N14621, N9534, N1479);
or OR3 (N14633, N14616, N12109, N11942);
and AND4 (N14634, N14618, N10938, N8516, N4363);
buf BUF1 (N14635, N14634);
xor XOR2 (N14636, N14620, N7954);
not NOT1 (N14637, N14633);
xor XOR2 (N14638, N14632, N13662);
xor XOR2 (N14639, N14635, N274);
and AND3 (N14640, N14614, N1797, N9622);
nor NOR3 (N14641, N14640, N5653, N9819);
and AND3 (N14642, N14637, N10599, N10709);
or OR3 (N14643, N14626, N13118, N3482);
nand NAND2 (N14644, N14624, N8405);
buf BUF1 (N14645, N14639);
nor NOR2 (N14646, N14642, N2288);
nand NAND4 (N14647, N14641, N9808, N14371, N8923);
nor NOR3 (N14648, N14636, N7520, N8238);
and AND3 (N14649, N14630, N9834, N4010);
nand NAND2 (N14650, N14638, N11808);
nand NAND2 (N14651, N14650, N146);
or OR3 (N14652, N14631, N3137, N6859);
nor NOR3 (N14653, N14645, N6375, N14005);
not NOT1 (N14654, N14652);
nand NAND4 (N14655, N14654, N7696, N9543, N2809);
or OR3 (N14656, N14628, N8344, N703);
and AND4 (N14657, N14653, N1138, N12450, N9953);
nor NOR4 (N14658, N14646, N8660, N5618, N3197);
not NOT1 (N14659, N14643);
and AND4 (N14660, N14648, N13068, N9435, N9854);
xor XOR2 (N14661, N14660, N8074);
nand NAND2 (N14662, N14644, N7239);
buf BUF1 (N14663, N14662);
and AND3 (N14664, N14659, N13106, N5935);
nand NAND3 (N14665, N14658, N2355, N8688);
nor NOR2 (N14666, N14647, N7720);
nand NAND2 (N14667, N14656, N8112);
nor NOR2 (N14668, N14664, N2271);
buf BUF1 (N14669, N14651);
xor XOR2 (N14670, N14665, N8441);
not NOT1 (N14671, N14657);
xor XOR2 (N14672, N14671, N7726);
xor XOR2 (N14673, N14666, N13442);
not NOT1 (N14674, N14672);
buf BUF1 (N14675, N14670);
nor NOR3 (N14676, N14669, N4311, N13283);
or OR3 (N14677, N14667, N1770, N9601);
buf BUF1 (N14678, N14674);
or OR3 (N14679, N14673, N12859, N3832);
and AND2 (N14680, N14676, N2410);
or OR4 (N14681, N14678, N10211, N1601, N7702);
nand NAND2 (N14682, N14668, N13416);
not NOT1 (N14683, N14663);
and AND2 (N14684, N14661, N8020);
nor NOR3 (N14685, N14680, N6972, N8926);
or OR2 (N14686, N14675, N3053);
and AND3 (N14687, N14683, N10666, N5935);
nand NAND4 (N14688, N14655, N8952, N6961, N6482);
not NOT1 (N14689, N14679);
nor NOR4 (N14690, N14682, N1950, N8778, N5746);
and AND2 (N14691, N14677, N5767);
or OR2 (N14692, N14684, N10439);
xor XOR2 (N14693, N14689, N11125);
and AND2 (N14694, N14691, N10191);
or OR3 (N14695, N14649, N14428, N1268);
buf BUF1 (N14696, N14693);
buf BUF1 (N14697, N14681);
nand NAND2 (N14698, N14690, N7143);
buf BUF1 (N14699, N14688);
nor NOR3 (N14700, N14694, N14687, N8703);
nand NAND2 (N14701, N14146, N6784);
nor NOR4 (N14702, N14701, N9288, N4746, N7929);
xor XOR2 (N14703, N14698, N1984);
not NOT1 (N14704, N14702);
or OR2 (N14705, N14704, N5243);
not NOT1 (N14706, N14696);
nand NAND2 (N14707, N14699, N2919);
or OR4 (N14708, N14692, N781, N12670, N3583);
not NOT1 (N14709, N14700);
or OR2 (N14710, N14709, N14619);
not NOT1 (N14711, N14705);
not NOT1 (N14712, N14707);
not NOT1 (N14713, N14708);
nand NAND3 (N14714, N14685, N193, N6403);
buf BUF1 (N14715, N14703);
or OR4 (N14716, N14715, N4806, N2443, N9942);
not NOT1 (N14717, N14697);
nand NAND3 (N14718, N14716, N6548, N14714);
and AND2 (N14719, N1103, N1169);
and AND4 (N14720, N14686, N4077, N5149, N6900);
nor NOR4 (N14721, N14719, N14068, N2553, N3169);
not NOT1 (N14722, N14706);
or OR3 (N14723, N14695, N11303, N5008);
buf BUF1 (N14724, N14712);
nand NAND3 (N14725, N14713, N4033, N804);
not NOT1 (N14726, N14711);
buf BUF1 (N14727, N14724);
nand NAND2 (N14728, N14726, N8456);
or OR2 (N14729, N14717, N7960);
nand NAND4 (N14730, N14728, N13794, N2892, N5192);
or OR2 (N14731, N14730, N3432);
not NOT1 (N14732, N14720);
buf BUF1 (N14733, N14722);
xor XOR2 (N14734, N14732, N5933);
or OR4 (N14735, N14725, N10419, N8145, N11628);
buf BUF1 (N14736, N14735);
and AND2 (N14737, N14723, N11987);
xor XOR2 (N14738, N14733, N13165);
nor NOR4 (N14739, N14727, N13656, N6206, N10204);
buf BUF1 (N14740, N14734);
nor NOR3 (N14741, N14740, N6936, N5920);
nand NAND4 (N14742, N14718, N2478, N2921, N13897);
xor XOR2 (N14743, N14721, N8326);
not NOT1 (N14744, N14729);
not NOT1 (N14745, N14731);
or OR3 (N14746, N14744, N12031, N10443);
buf BUF1 (N14747, N14743);
nor NOR3 (N14748, N14746, N9544, N8752);
and AND4 (N14749, N14710, N8142, N3756, N9899);
and AND3 (N14750, N14747, N3633, N8631);
or OR4 (N14751, N14750, N51, N4273, N9545);
or OR2 (N14752, N14742, N2112);
and AND2 (N14753, N14738, N6670);
or OR4 (N14754, N14739, N11216, N4159, N6138);
not NOT1 (N14755, N14737);
or OR2 (N14756, N14753, N8416);
or OR3 (N14757, N14736, N10111, N4521);
or OR2 (N14758, N14745, N10976);
nor NOR3 (N14759, N14755, N1987, N1772);
buf BUF1 (N14760, N14758);
buf BUF1 (N14761, N14751);
nand NAND2 (N14762, N14756, N4068);
buf BUF1 (N14763, N14762);
or OR3 (N14764, N14749, N8064, N1529);
and AND2 (N14765, N14752, N10037);
xor XOR2 (N14766, N14760, N4831);
buf BUF1 (N14767, N14764);
and AND4 (N14768, N14767, N13661, N10704, N4551);
xor XOR2 (N14769, N14748, N3225);
xor XOR2 (N14770, N14761, N5267);
and AND4 (N14771, N14770, N10514, N13909, N5135);
or OR2 (N14772, N14771, N13995);
nor NOR2 (N14773, N14766, N10199);
and AND3 (N14774, N14769, N5307, N12139);
nand NAND3 (N14775, N14759, N9150, N10017);
buf BUF1 (N14776, N14754);
and AND2 (N14777, N14757, N13576);
nand NAND3 (N14778, N14768, N589, N1695);
and AND2 (N14779, N14776, N12701);
and AND3 (N14780, N14741, N4904, N9584);
nor NOR3 (N14781, N14774, N9689, N13622);
not NOT1 (N14782, N14779);
buf BUF1 (N14783, N14763);
nor NOR4 (N14784, N14781, N5517, N2377, N3948);
and AND2 (N14785, N14775, N14144);
nand NAND4 (N14786, N14777, N12816, N906, N12837);
or OR3 (N14787, N14773, N4873, N5089);
or OR3 (N14788, N14765, N3597, N9082);
and AND4 (N14789, N14786, N10432, N3813, N9842);
or OR3 (N14790, N14783, N11677, N1761);
or OR2 (N14791, N14787, N9608);
buf BUF1 (N14792, N14788);
or OR2 (N14793, N14785, N7387);
or OR3 (N14794, N14784, N11818, N5936);
and AND4 (N14795, N14780, N3771, N5591, N417);
or OR2 (N14796, N14782, N13018);
not NOT1 (N14797, N14789);
and AND4 (N14798, N14793, N569, N917, N7611);
buf BUF1 (N14799, N14796);
buf BUF1 (N14800, N14794);
or OR2 (N14801, N14799, N1213);
and AND3 (N14802, N14792, N13138, N6563);
and AND2 (N14803, N14790, N5001);
not NOT1 (N14804, N14803);
nor NOR2 (N14805, N14801, N7789);
nand NAND2 (N14806, N14802, N10019);
and AND2 (N14807, N14805, N14134);
nand NAND2 (N14808, N14806, N7045);
not NOT1 (N14809, N14800);
and AND3 (N14810, N14804, N14509, N11477);
buf BUF1 (N14811, N14807);
and AND4 (N14812, N14798, N94, N298, N14397);
nand NAND2 (N14813, N14772, N5391);
and AND2 (N14814, N14795, N2396);
buf BUF1 (N14815, N14813);
or OR4 (N14816, N14809, N7471, N561, N7177);
and AND3 (N14817, N14810, N1054, N2573);
nor NOR4 (N14818, N14808, N6133, N5695, N9634);
or OR3 (N14819, N14818, N7875, N9616);
nand NAND3 (N14820, N14791, N625, N5476);
xor XOR2 (N14821, N14819, N2425);
xor XOR2 (N14822, N14817, N13823);
not NOT1 (N14823, N14811);
and AND2 (N14824, N14816, N11017);
nand NAND4 (N14825, N14820, N14027, N12803, N1576);
nor NOR2 (N14826, N14824, N2945);
and AND4 (N14827, N14823, N6487, N4776, N504);
or OR4 (N14828, N14822, N3494, N13452, N11088);
or OR2 (N14829, N14828, N8413);
nand NAND4 (N14830, N14778, N14146, N12395, N3923);
buf BUF1 (N14831, N14814);
or OR2 (N14832, N14829, N4236);
buf BUF1 (N14833, N14815);
buf BUF1 (N14834, N14830);
nor NOR2 (N14835, N14812, N14773);
nor NOR2 (N14836, N14827, N12276);
or OR2 (N14837, N14797, N6619);
nand NAND2 (N14838, N14835, N13172);
nor NOR3 (N14839, N14821, N1208, N8170);
nor NOR4 (N14840, N14837, N14481, N9359, N4651);
nor NOR2 (N14841, N14832, N14326);
or OR3 (N14842, N14841, N6506, N1463);
xor XOR2 (N14843, N14833, N1319);
and AND2 (N14844, N14825, N2180);
not NOT1 (N14845, N14826);
nand NAND2 (N14846, N14836, N6301);
nor NOR2 (N14847, N14845, N2676);
not NOT1 (N14848, N14839);
xor XOR2 (N14849, N14844, N3280);
and AND3 (N14850, N14848, N8758, N3987);
not NOT1 (N14851, N14834);
nor NOR2 (N14852, N14846, N1369);
buf BUF1 (N14853, N14831);
xor XOR2 (N14854, N14850, N1814);
and AND4 (N14855, N14843, N4329, N8586, N12988);
or OR4 (N14856, N14840, N10726, N12564, N13996);
or OR4 (N14857, N14842, N2114, N2801, N1161);
nor NOR3 (N14858, N14854, N2932, N10982);
nand NAND2 (N14859, N14838, N10440);
not NOT1 (N14860, N14851);
xor XOR2 (N14861, N14849, N2623);
buf BUF1 (N14862, N14859);
nand NAND2 (N14863, N14852, N2952);
xor XOR2 (N14864, N14857, N10534);
buf BUF1 (N14865, N14860);
or OR3 (N14866, N14861, N8590, N13144);
xor XOR2 (N14867, N14866, N13468);
nor NOR3 (N14868, N14856, N9866, N2470);
or OR2 (N14869, N14847, N7429);
nand NAND4 (N14870, N14865, N7898, N4932, N11105);
nor NOR4 (N14871, N14869, N4623, N13748, N14482);
and AND3 (N14872, N14855, N8124, N12108);
and AND3 (N14873, N14863, N13529, N11864);
xor XOR2 (N14874, N14858, N6004);
nand NAND3 (N14875, N14873, N10805, N7949);
nand NAND4 (N14876, N14872, N998, N1237, N4610);
nor NOR4 (N14877, N14875, N12371, N6509, N14674);
or OR3 (N14878, N14874, N2008, N8289);
nor NOR3 (N14879, N14878, N10088, N7770);
buf BUF1 (N14880, N14870);
buf BUF1 (N14881, N14880);
and AND4 (N14882, N14868, N5711, N10095, N4606);
not NOT1 (N14883, N14867);
buf BUF1 (N14884, N14879);
and AND4 (N14885, N14862, N2501, N7316, N1120);
xor XOR2 (N14886, N14883, N3537);
buf BUF1 (N14887, N14864);
nand NAND4 (N14888, N14876, N7512, N5048, N5736);
nand NAND3 (N14889, N14886, N6330, N8567);
nand NAND2 (N14890, N14884, N12093);
not NOT1 (N14891, N14882);
and AND4 (N14892, N14877, N9564, N10795, N4646);
xor XOR2 (N14893, N14891, N14613);
nor NOR3 (N14894, N14893, N8444, N11811);
nand NAND4 (N14895, N14887, N14264, N6468, N7459);
not NOT1 (N14896, N14885);
buf BUF1 (N14897, N14895);
buf BUF1 (N14898, N14892);
or OR4 (N14899, N14889, N12610, N6173, N2054);
nand NAND2 (N14900, N14894, N13080);
buf BUF1 (N14901, N14890);
and AND4 (N14902, N14898, N10276, N14361, N6354);
xor XOR2 (N14903, N14881, N7387);
nand NAND3 (N14904, N14903, N11280, N955);
and AND3 (N14905, N14853, N14109, N8240);
and AND4 (N14906, N14897, N13610, N10124, N5448);
nand NAND3 (N14907, N14905, N1983, N450);
nor NOR2 (N14908, N14896, N7005);
or OR2 (N14909, N14900, N8868);
not NOT1 (N14910, N14904);
nand NAND2 (N14911, N14910, N341);
not NOT1 (N14912, N14888);
nand NAND2 (N14913, N14902, N1111);
and AND4 (N14914, N14871, N10391, N13370, N9173);
nand NAND2 (N14915, N14909, N11643);
nor NOR3 (N14916, N14912, N5154, N6406);
and AND3 (N14917, N14911, N10505, N1559);
nor NOR4 (N14918, N14916, N11729, N8305, N10291);
not NOT1 (N14919, N14901);
nand NAND3 (N14920, N14919, N113, N5541);
nand NAND3 (N14921, N14899, N2588, N9382);
not NOT1 (N14922, N14920);
nand NAND2 (N14923, N14922, N8518);
or OR3 (N14924, N14914, N8783, N14010);
not NOT1 (N14925, N14924);
xor XOR2 (N14926, N14913, N11021);
and AND4 (N14927, N14918, N2961, N6928, N9598);
not NOT1 (N14928, N14907);
buf BUF1 (N14929, N14921);
nor NOR4 (N14930, N14923, N14138, N3414, N787);
nand NAND3 (N14931, N14926, N2485, N1772);
not NOT1 (N14932, N14917);
or OR2 (N14933, N14932, N557);
buf BUF1 (N14934, N14908);
xor XOR2 (N14935, N14930, N14436);
nor NOR4 (N14936, N14933, N13636, N4061, N11888);
nand NAND4 (N14937, N14928, N7377, N6517, N8244);
buf BUF1 (N14938, N14925);
nor NOR4 (N14939, N14927, N10116, N3669, N11278);
or OR4 (N14940, N14935, N4008, N9103, N12747);
or OR4 (N14941, N14940, N6944, N1087, N5634);
nor NOR4 (N14942, N14938, N10554, N226, N3151);
and AND3 (N14943, N14934, N12643, N7201);
or OR2 (N14944, N14906, N3664);
or OR4 (N14945, N14943, N14515, N11907, N10274);
nor NOR4 (N14946, N14941, N7514, N1416, N5105);
xor XOR2 (N14947, N14939, N9024);
nand NAND4 (N14948, N14915, N14197, N3906, N11231);
xor XOR2 (N14949, N14931, N4596);
and AND4 (N14950, N14936, N5566, N8460, N13413);
or OR4 (N14951, N14937, N14021, N11654, N6499);
xor XOR2 (N14952, N14950, N7339);
or OR3 (N14953, N14929, N6752, N13440);
and AND3 (N14954, N14949, N5147, N3500);
and AND3 (N14955, N14944, N10442, N112);
not NOT1 (N14956, N14945);
xor XOR2 (N14957, N14955, N5216);
nor NOR3 (N14958, N14954, N8335, N6552);
and AND3 (N14959, N14957, N7794, N1753);
xor XOR2 (N14960, N14958, N6263);
buf BUF1 (N14961, N14948);
nor NOR4 (N14962, N14961, N11406, N13554, N540);
and AND2 (N14963, N14953, N14292);
nand NAND4 (N14964, N14942, N6348, N13074, N4913);
nand NAND3 (N14965, N14947, N7429, N10429);
nand NAND2 (N14966, N14956, N5566);
and AND3 (N14967, N14965, N12944, N3585);
and AND4 (N14968, N14966, N11573, N5221, N12100);
and AND4 (N14969, N14952, N914, N1921, N8727);
buf BUF1 (N14970, N14969);
nor NOR3 (N14971, N14959, N11957, N3736);
nand NAND3 (N14972, N14968, N7055, N8843);
and AND4 (N14973, N14962, N6309, N6556, N1412);
nor NOR3 (N14974, N14967, N10959, N4803);
or OR3 (N14975, N14972, N4982, N6086);
buf BUF1 (N14976, N14964);
not NOT1 (N14977, N14974);
buf BUF1 (N14978, N14973);
not NOT1 (N14979, N14960);
xor XOR2 (N14980, N14946, N4338);
xor XOR2 (N14981, N14970, N11169);
not NOT1 (N14982, N14951);
buf BUF1 (N14983, N14978);
nor NOR2 (N14984, N14982, N156);
not NOT1 (N14985, N14981);
nor NOR4 (N14986, N14984, N6222, N8121, N5765);
nor NOR4 (N14987, N14985, N3240, N12231, N11486);
xor XOR2 (N14988, N14979, N4818);
not NOT1 (N14989, N14976);
and AND4 (N14990, N14988, N7308, N5292, N1399);
buf BUF1 (N14991, N14989);
or OR2 (N14992, N14983, N9941);
not NOT1 (N14993, N14977);
buf BUF1 (N14994, N14963);
nand NAND4 (N14995, N14993, N12093, N711, N14546);
not NOT1 (N14996, N14975);
xor XOR2 (N14997, N14991, N7905);
and AND3 (N14998, N14971, N11086, N10405);
nor NOR3 (N14999, N14987, N12871, N11346);
or OR2 (N15000, N14992, N2351);
or OR4 (N15001, N14995, N11380, N13922, N2391);
nor NOR2 (N15002, N14986, N529);
xor XOR2 (N15003, N14996, N11808);
nand NAND4 (N15004, N14997, N8929, N12632, N6143);
and AND4 (N15005, N14998, N2624, N6230, N3814);
or OR4 (N15006, N14990, N4235, N6444, N6318);
nand NAND4 (N15007, N14994, N3025, N12512, N8457);
or OR3 (N15008, N15004, N1448, N2066);
or OR2 (N15009, N15006, N10163);
nand NAND2 (N15010, N15002, N9999);
buf BUF1 (N15011, N15000);
not NOT1 (N15012, N15008);
xor XOR2 (N15013, N15011, N7548);
or OR3 (N15014, N15012, N2556, N10276);
nor NOR4 (N15015, N15010, N14562, N14260, N2421);
or OR3 (N15016, N14980, N7922, N4145);
not NOT1 (N15017, N15013);
not NOT1 (N15018, N15005);
or OR4 (N15019, N15017, N8443, N649, N11456);
xor XOR2 (N15020, N14999, N314);
nand NAND4 (N15021, N15019, N12930, N7006, N5847);
nand NAND4 (N15022, N15016, N8736, N3307, N6782);
not NOT1 (N15023, N15020);
nand NAND2 (N15024, N15014, N13700);
nor NOR4 (N15025, N15003, N4899, N2479, N12025);
xor XOR2 (N15026, N15024, N5798);
xor XOR2 (N15027, N15023, N9745);
not NOT1 (N15028, N15001);
xor XOR2 (N15029, N15027, N14883);
buf BUF1 (N15030, N15026);
buf BUF1 (N15031, N15025);
nand NAND2 (N15032, N15009, N10168);
nor NOR3 (N15033, N15022, N9245, N9360);
xor XOR2 (N15034, N15018, N8346);
not NOT1 (N15035, N15015);
buf BUF1 (N15036, N15033);
not NOT1 (N15037, N15029);
nand NAND2 (N15038, N15035, N1593);
nor NOR4 (N15039, N15028, N3829, N14084, N12717);
nand NAND4 (N15040, N15038, N9243, N4468, N648);
xor XOR2 (N15041, N15037, N11615);
nor NOR2 (N15042, N15034, N6987);
xor XOR2 (N15043, N15032, N2993);
or OR4 (N15044, N15007, N1113, N5391, N3452);
not NOT1 (N15045, N15031);
or OR3 (N15046, N15039, N14691, N13192);
or OR4 (N15047, N15021, N5739, N4248, N13777);
not NOT1 (N15048, N15040);
and AND2 (N15049, N15041, N9800);
and AND2 (N15050, N15044, N2838);
and AND3 (N15051, N15050, N11187, N13963);
and AND3 (N15052, N15045, N11357, N8247);
buf BUF1 (N15053, N15048);
nor NOR4 (N15054, N15052, N13839, N562, N6720);
or OR4 (N15055, N15054, N14457, N253, N10305);
not NOT1 (N15056, N15053);
nor NOR3 (N15057, N15046, N4723, N5691);
and AND2 (N15058, N15049, N5748);
or OR4 (N15059, N15057, N456, N4535, N8706);
xor XOR2 (N15060, N15055, N3045);
and AND4 (N15061, N15047, N1786, N2694, N1278);
not NOT1 (N15062, N15060);
xor XOR2 (N15063, N15042, N6697);
or OR2 (N15064, N15059, N10385);
nand NAND2 (N15065, N15064, N3788);
buf BUF1 (N15066, N15061);
nor NOR4 (N15067, N15063, N12458, N4491, N6314);
or OR4 (N15068, N15065, N8975, N8263, N4193);
nand NAND3 (N15069, N15062, N9931, N12838);
xor XOR2 (N15070, N15043, N10254);
nor NOR4 (N15071, N15069, N8918, N13299, N1504);
not NOT1 (N15072, N15071);
buf BUF1 (N15073, N15030);
not NOT1 (N15074, N15067);
xor XOR2 (N15075, N15051, N10592);
or OR3 (N15076, N15072, N177, N13499);
nor NOR4 (N15077, N15056, N1568, N2178, N13629);
and AND3 (N15078, N15073, N14880, N11114);
not NOT1 (N15079, N15076);
nor NOR4 (N15080, N15075, N7964, N8011, N1853);
nand NAND2 (N15081, N15036, N3024);
or OR3 (N15082, N15058, N7084, N3635);
or OR2 (N15083, N15082, N4772);
buf BUF1 (N15084, N15068);
nor NOR3 (N15085, N15080, N470, N12582);
nand NAND2 (N15086, N15070, N9813);
nor NOR3 (N15087, N15084, N10300, N2394);
or OR3 (N15088, N15077, N9909, N11913);
xor XOR2 (N15089, N15086, N1967);
nand NAND2 (N15090, N15081, N11370);
nor NOR3 (N15091, N15078, N8962, N6288);
nand NAND2 (N15092, N15083, N11990);
not NOT1 (N15093, N15090);
nand NAND4 (N15094, N15092, N13931, N12162, N3568);
or OR2 (N15095, N15088, N7553);
xor XOR2 (N15096, N15093, N11420);
and AND2 (N15097, N15066, N14963);
nor NOR3 (N15098, N15089, N5774, N3533);
xor XOR2 (N15099, N15079, N8174);
buf BUF1 (N15100, N15097);
and AND3 (N15101, N15094, N4181, N9426);
buf BUF1 (N15102, N15085);
nor NOR4 (N15103, N15091, N5395, N5294, N4831);
xor XOR2 (N15104, N15103, N8163);
not NOT1 (N15105, N15087);
nor NOR3 (N15106, N15074, N4639, N6796);
not NOT1 (N15107, N15099);
or OR3 (N15108, N15106, N7989, N13804);
or OR3 (N15109, N15100, N4526, N6088);
or OR4 (N15110, N15109, N14113, N3656, N1832);
not NOT1 (N15111, N15095);
xor XOR2 (N15112, N15104, N428);
nand NAND2 (N15113, N15111, N9968);
nand NAND4 (N15114, N15113, N5894, N4314, N11343);
or OR4 (N15115, N15101, N6237, N7408, N12736);
xor XOR2 (N15116, N15098, N411);
buf BUF1 (N15117, N15107);
not NOT1 (N15118, N15112);
nor NOR3 (N15119, N15102, N3252, N2494);
xor XOR2 (N15120, N15117, N3020);
nor NOR2 (N15121, N15115, N779);
nor NOR2 (N15122, N15119, N12719);
buf BUF1 (N15123, N15108);
not NOT1 (N15124, N15110);
xor XOR2 (N15125, N15121, N7730);
buf BUF1 (N15126, N15114);
and AND2 (N15127, N15105, N7609);
nand NAND3 (N15128, N15122, N4463, N13230);
not NOT1 (N15129, N15125);
xor XOR2 (N15130, N15118, N13068);
and AND3 (N15131, N15096, N2826, N12475);
nor NOR3 (N15132, N15120, N14769, N14648);
or OR2 (N15133, N15127, N655);
nor NOR3 (N15134, N15129, N3764, N4992);
buf BUF1 (N15135, N15124);
nor NOR3 (N15136, N15123, N3, N4015);
nand NAND4 (N15137, N15128, N9160, N10992, N11093);
and AND4 (N15138, N15130, N14714, N11132, N12958);
nand NAND4 (N15139, N15116, N12981, N7563, N3702);
nor NOR2 (N15140, N15134, N6422);
not NOT1 (N15141, N15133);
buf BUF1 (N15142, N15138);
or OR2 (N15143, N15132, N4346);
or OR2 (N15144, N15126, N6287);
nand NAND3 (N15145, N15142, N12497, N11009);
not NOT1 (N15146, N15137);
or OR2 (N15147, N15143, N9874);
nand NAND2 (N15148, N15145, N14002);
nand NAND4 (N15149, N15131, N1458, N907, N4898);
buf BUF1 (N15150, N15136);
nand NAND2 (N15151, N15148, N8031);
nor NOR2 (N15152, N15135, N10370);
and AND2 (N15153, N15139, N10958);
and AND4 (N15154, N15147, N12318, N8841, N10368);
and AND2 (N15155, N15141, N11998);
nand NAND3 (N15156, N15155, N4759, N3458);
buf BUF1 (N15157, N15154);
and AND4 (N15158, N15149, N6423, N3564, N2236);
xor XOR2 (N15159, N15158, N8932);
xor XOR2 (N15160, N15140, N3865);
nand NAND2 (N15161, N15151, N4648);
nand NAND2 (N15162, N15161, N12644);
or OR2 (N15163, N15162, N431);
and AND4 (N15164, N15160, N12178, N13777, N12580);
nor NOR4 (N15165, N15152, N6302, N8583, N11707);
not NOT1 (N15166, N15144);
xor XOR2 (N15167, N15165, N11291);
and AND3 (N15168, N15150, N13224, N4413);
or OR2 (N15169, N15168, N12022);
or OR2 (N15170, N15163, N10153);
nor NOR3 (N15171, N15169, N2452, N10246);
not NOT1 (N15172, N15156);
xor XOR2 (N15173, N15172, N15069);
and AND2 (N15174, N15153, N12116);
nand NAND3 (N15175, N15166, N14239, N5786);
and AND4 (N15176, N15157, N9909, N13409, N4872);
or OR3 (N15177, N15175, N11356, N14268);
not NOT1 (N15178, N15173);
nor NOR3 (N15179, N15176, N14275, N7319);
xor XOR2 (N15180, N15174, N9148);
xor XOR2 (N15181, N15146, N14822);
buf BUF1 (N15182, N15177);
and AND4 (N15183, N15164, N8259, N10148, N5904);
or OR3 (N15184, N15180, N8035, N11598);
and AND3 (N15185, N15184, N7732, N1632);
xor XOR2 (N15186, N15185, N7069);
or OR4 (N15187, N15186, N3714, N4230, N4488);
and AND3 (N15188, N15187, N14620, N239);
nor NOR3 (N15189, N15181, N11236, N2540);
nor NOR3 (N15190, N15183, N10451, N5635);
or OR4 (N15191, N15179, N8415, N7484, N3711);
and AND2 (N15192, N15191, N2584);
or OR4 (N15193, N15192, N3093, N6247, N11885);
xor XOR2 (N15194, N15189, N5945);
xor XOR2 (N15195, N15193, N8196);
nor NOR3 (N15196, N15178, N15064, N5873);
and AND3 (N15197, N15167, N10574, N14264);
xor XOR2 (N15198, N15190, N1969);
or OR4 (N15199, N15195, N3645, N3179, N6954);
not NOT1 (N15200, N15199);
nand NAND2 (N15201, N15196, N5901);
and AND4 (N15202, N15201, N5129, N2284, N40);
nand NAND3 (N15203, N15182, N7553, N5486);
buf BUF1 (N15204, N15197);
or OR4 (N15205, N15188, N9792, N8638, N11283);
xor XOR2 (N15206, N15159, N14098);
not NOT1 (N15207, N15171);
nor NOR3 (N15208, N15200, N14795, N2039);
and AND3 (N15209, N15207, N5680, N7627);
buf BUF1 (N15210, N15205);
nand NAND4 (N15211, N15209, N4656, N7489, N7035);
buf BUF1 (N15212, N15211);
and AND4 (N15213, N15206, N6326, N5896, N6696);
not NOT1 (N15214, N15213);
or OR2 (N15215, N15170, N7981);
or OR2 (N15216, N15214, N9516);
and AND2 (N15217, N15212, N12510);
xor XOR2 (N15218, N15194, N5479);
or OR2 (N15219, N15217, N3112);
and AND3 (N15220, N15219, N9749, N6349);
nand NAND4 (N15221, N15216, N8574, N12213, N5529);
and AND4 (N15222, N15210, N397, N10808, N787);
buf BUF1 (N15223, N15202);
and AND2 (N15224, N15203, N4657);
or OR4 (N15225, N15215, N8168, N6913, N2562);
buf BUF1 (N15226, N15198);
buf BUF1 (N15227, N15208);
or OR3 (N15228, N15227, N13426, N2179);
and AND3 (N15229, N15225, N14215, N13377);
and AND4 (N15230, N15229, N11645, N11664, N1237);
nor NOR4 (N15231, N15221, N7518, N14066, N13145);
nand NAND4 (N15232, N15218, N1580, N12992, N6632);
xor XOR2 (N15233, N15204, N3206);
nor NOR2 (N15234, N15220, N3365);
nand NAND2 (N15235, N15233, N12059);
and AND4 (N15236, N15226, N1807, N12835, N4887);
not NOT1 (N15237, N15222);
xor XOR2 (N15238, N15232, N12859);
xor XOR2 (N15239, N15234, N2051);
buf BUF1 (N15240, N15239);
or OR3 (N15241, N15231, N642, N2095);
not NOT1 (N15242, N15241);
nand NAND2 (N15243, N15228, N2671);
buf BUF1 (N15244, N15236);
not NOT1 (N15245, N15240);
buf BUF1 (N15246, N15237);
xor XOR2 (N15247, N15246, N6854);
nand NAND4 (N15248, N15247, N10654, N10506, N1595);
nor NOR4 (N15249, N15243, N14437, N4799, N13266);
not NOT1 (N15250, N15244);
nor NOR3 (N15251, N15250, N9581, N13415);
xor XOR2 (N15252, N15230, N768);
not NOT1 (N15253, N15251);
or OR2 (N15254, N15249, N144);
not NOT1 (N15255, N15253);
nand NAND3 (N15256, N15235, N9318, N7790);
or OR4 (N15257, N15248, N14063, N2892, N10119);
buf BUF1 (N15258, N15255);
xor XOR2 (N15259, N15254, N14215);
or OR4 (N15260, N15223, N696, N11524, N12405);
or OR2 (N15261, N15238, N4642);
and AND2 (N15262, N15242, N6461);
nor NOR4 (N15263, N15245, N1920, N3623, N11028);
nand NAND4 (N15264, N15257, N11394, N14765, N2114);
buf BUF1 (N15265, N15259);
and AND3 (N15266, N15265, N14987, N14696);
not NOT1 (N15267, N15256);
not NOT1 (N15268, N15261);
buf BUF1 (N15269, N15268);
not NOT1 (N15270, N15262);
and AND3 (N15271, N15270, N875, N4989);
and AND3 (N15272, N15269, N15154, N6927);
buf BUF1 (N15273, N15266);
buf BUF1 (N15274, N15271);
and AND3 (N15275, N15263, N1672, N11035);
and AND2 (N15276, N15274, N7892);
buf BUF1 (N15277, N15224);
buf BUF1 (N15278, N15252);
xor XOR2 (N15279, N15260, N11634);
xor XOR2 (N15280, N15264, N3174);
xor XOR2 (N15281, N15276, N2303);
buf BUF1 (N15282, N15279);
nand NAND2 (N15283, N15258, N1536);
and AND4 (N15284, N15272, N14210, N3812, N1208);
nand NAND3 (N15285, N15284, N1503, N853);
or OR3 (N15286, N15275, N10059, N9808);
nor NOR3 (N15287, N15267, N7194, N10834);
not NOT1 (N15288, N15286);
xor XOR2 (N15289, N15287, N6048);
nor NOR4 (N15290, N15273, N13734, N10636, N12875);
nand NAND3 (N15291, N15289, N13173, N6297);
buf BUF1 (N15292, N15291);
and AND3 (N15293, N15290, N10881, N12922);
nor NOR2 (N15294, N15288, N5578);
and AND3 (N15295, N15282, N5816, N1900);
nor NOR4 (N15296, N15294, N9772, N11484, N13594);
or OR4 (N15297, N15292, N7129, N14666, N13667);
nor NOR3 (N15298, N15295, N1791, N3483);
nor NOR2 (N15299, N15298, N1567);
or OR4 (N15300, N15285, N5738, N9150, N7666);
and AND2 (N15301, N15299, N12004);
not NOT1 (N15302, N15281);
or OR4 (N15303, N15283, N4140, N1171, N8893);
buf BUF1 (N15304, N15303);
buf BUF1 (N15305, N15304);
nand NAND2 (N15306, N15301, N8373);
not NOT1 (N15307, N15277);
nor NOR2 (N15308, N15302, N2368);
or OR4 (N15309, N15308, N13274, N5896, N12166);
not NOT1 (N15310, N15280);
buf BUF1 (N15311, N15278);
or OR4 (N15312, N15310, N2115, N10002, N3006);
or OR2 (N15313, N15309, N15163);
or OR3 (N15314, N15307, N1006, N8441);
nand NAND4 (N15315, N15314, N12049, N14507, N14606);
not NOT1 (N15316, N15311);
or OR2 (N15317, N15296, N6489);
nor NOR3 (N15318, N15297, N10737, N11452);
or OR2 (N15319, N15305, N7125);
or OR2 (N15320, N15306, N11703);
nor NOR3 (N15321, N15320, N14287, N11898);
nand NAND2 (N15322, N15317, N5417);
not NOT1 (N15323, N15312);
nor NOR2 (N15324, N15323, N10092);
and AND3 (N15325, N15316, N6379, N8479);
buf BUF1 (N15326, N15300);
or OR4 (N15327, N15319, N13742, N14444, N10687);
or OR2 (N15328, N15326, N14200);
buf BUF1 (N15329, N15293);
or OR4 (N15330, N15318, N7434, N10331, N10731);
and AND3 (N15331, N15325, N8717, N8855);
xor XOR2 (N15332, N15329, N13127);
nand NAND3 (N15333, N15332, N12712, N7182);
and AND3 (N15334, N15333, N1122, N12067);
and AND4 (N15335, N15328, N5557, N6732, N11562);
xor XOR2 (N15336, N15330, N8423);
nand NAND3 (N15337, N15327, N9875, N3928);
xor XOR2 (N15338, N15337, N5864);
nand NAND2 (N15339, N15336, N2767);
xor XOR2 (N15340, N15315, N13270);
xor XOR2 (N15341, N15334, N1211);
xor XOR2 (N15342, N15339, N4617);
not NOT1 (N15343, N15331);
nor NOR4 (N15344, N15335, N13647, N10035, N14300);
and AND3 (N15345, N15343, N12730, N1367);
not NOT1 (N15346, N15344);
not NOT1 (N15347, N15346);
xor XOR2 (N15348, N15324, N9782);
and AND3 (N15349, N15340, N7618, N9962);
xor XOR2 (N15350, N15349, N10999);
buf BUF1 (N15351, N15347);
nor NOR3 (N15352, N15338, N13562, N10159);
nand NAND3 (N15353, N15341, N2771, N11190);
nand NAND3 (N15354, N15350, N10990, N9174);
not NOT1 (N15355, N15321);
not NOT1 (N15356, N15313);
xor XOR2 (N15357, N15352, N9585);
not NOT1 (N15358, N15354);
nand NAND2 (N15359, N15345, N374);
xor XOR2 (N15360, N15322, N5133);
nor NOR4 (N15361, N15358, N1172, N10303, N3679);
not NOT1 (N15362, N15353);
not NOT1 (N15363, N15362);
and AND2 (N15364, N15359, N13044);
xor XOR2 (N15365, N15356, N12049);
xor XOR2 (N15366, N15360, N4522);
not NOT1 (N15367, N15351);
not NOT1 (N15368, N15361);
buf BUF1 (N15369, N15367);
xor XOR2 (N15370, N15369, N4448);
xor XOR2 (N15371, N15368, N8847);
nor NOR2 (N15372, N15364, N11583);
not NOT1 (N15373, N15370);
not NOT1 (N15374, N15373);
nor NOR3 (N15375, N15372, N4362, N1462);
nor NOR2 (N15376, N15348, N10226);
nor NOR2 (N15377, N15363, N9591);
nand NAND3 (N15378, N15366, N12446, N4602);
xor XOR2 (N15379, N15377, N3398);
nand NAND3 (N15380, N15371, N7667, N14968);
not NOT1 (N15381, N15380);
not NOT1 (N15382, N15365);
nor NOR4 (N15383, N15382, N11894, N2970, N1724);
xor XOR2 (N15384, N15355, N13759);
and AND4 (N15385, N15383, N10931, N4570, N89);
and AND4 (N15386, N15374, N13388, N13640, N5950);
xor XOR2 (N15387, N15381, N7809);
or OR4 (N15388, N15387, N3875, N1575, N5664);
nor NOR2 (N15389, N15378, N716);
buf BUF1 (N15390, N15386);
buf BUF1 (N15391, N15385);
xor XOR2 (N15392, N15342, N12044);
buf BUF1 (N15393, N15384);
nand NAND3 (N15394, N15390, N9791, N13571);
nand NAND3 (N15395, N15393, N4236, N11411);
xor XOR2 (N15396, N15395, N1109);
or OR3 (N15397, N15375, N11484, N2389);
buf BUF1 (N15398, N15396);
or OR3 (N15399, N15392, N1415, N10861);
nand NAND3 (N15400, N15388, N4676, N2479);
or OR2 (N15401, N15397, N12571);
xor XOR2 (N15402, N15376, N9659);
or OR2 (N15403, N15400, N9767);
buf BUF1 (N15404, N15403);
nor NOR2 (N15405, N15398, N923);
buf BUF1 (N15406, N15394);
nand NAND3 (N15407, N15405, N12486, N10026);
not NOT1 (N15408, N15389);
nor NOR3 (N15409, N15357, N12302, N10493);
and AND4 (N15410, N15406, N14462, N7801, N1304);
not NOT1 (N15411, N15410);
nor NOR2 (N15412, N15408, N1422);
nor NOR4 (N15413, N15404, N4261, N7878, N14835);
xor XOR2 (N15414, N15399, N13179);
buf BUF1 (N15415, N15391);
not NOT1 (N15416, N15402);
buf BUF1 (N15417, N15414);
not NOT1 (N15418, N15379);
buf BUF1 (N15419, N15412);
or OR3 (N15420, N15418, N6742, N5376);
xor XOR2 (N15421, N15401, N14259);
nand NAND3 (N15422, N15411, N298, N11534);
xor XOR2 (N15423, N15415, N3744);
and AND4 (N15424, N15407, N1141, N12368, N4499);
and AND4 (N15425, N15409, N11395, N1595, N1770);
nand NAND4 (N15426, N15424, N95, N2685, N14416);
nor NOR4 (N15427, N15420, N4827, N948, N14733);
and AND4 (N15428, N15417, N8422, N9711, N9802);
and AND4 (N15429, N15425, N5915, N11296, N10544);
buf BUF1 (N15430, N15419);
xor XOR2 (N15431, N15421, N11346);
xor XOR2 (N15432, N15428, N13246);
nor NOR3 (N15433, N15427, N9580, N7003);
nor NOR4 (N15434, N15431, N6966, N13093, N8339);
buf BUF1 (N15435, N15433);
nor NOR2 (N15436, N15423, N4783);
or OR4 (N15437, N15422, N4004, N13853, N11312);
not NOT1 (N15438, N15416);
nor NOR4 (N15439, N15426, N7787, N7096, N14445);
not NOT1 (N15440, N15437);
or OR2 (N15441, N15436, N10047);
xor XOR2 (N15442, N15429, N6043);
nand NAND3 (N15443, N15434, N4795, N8973);
xor XOR2 (N15444, N15430, N7432);
buf BUF1 (N15445, N15444);
buf BUF1 (N15446, N15438);
or OR2 (N15447, N15413, N3010);
nor NOR4 (N15448, N15440, N13316, N8239, N8276);
nand NAND4 (N15449, N15435, N3435, N13996, N10293);
or OR4 (N15450, N15448, N8408, N14681, N6200);
xor XOR2 (N15451, N15441, N1467);
nor NOR3 (N15452, N15447, N9170, N8454);
xor XOR2 (N15453, N15432, N2571);
nand NAND3 (N15454, N15443, N4656, N14208);
or OR2 (N15455, N15451, N2872);
or OR4 (N15456, N15453, N2512, N8935, N771);
or OR2 (N15457, N15442, N6531);
buf BUF1 (N15458, N15449);
nand NAND3 (N15459, N15456, N7303, N8375);
not NOT1 (N15460, N15455);
not NOT1 (N15461, N15459);
xor XOR2 (N15462, N15452, N1007);
buf BUF1 (N15463, N15457);
or OR3 (N15464, N15454, N8518, N512);
nand NAND2 (N15465, N15464, N13065);
not NOT1 (N15466, N15462);
or OR4 (N15467, N15458, N14492, N3392, N7594);
or OR4 (N15468, N15467, N15409, N7548, N6781);
buf BUF1 (N15469, N15461);
nor NOR4 (N15470, N15465, N12014, N8614, N10500);
nand NAND4 (N15471, N15466, N8968, N13677, N3127);
nor NOR2 (N15472, N15460, N13917);
and AND3 (N15473, N15471, N14407, N3950);
xor XOR2 (N15474, N15439, N15089);
and AND2 (N15475, N15445, N3843);
and AND4 (N15476, N15473, N2380, N6767, N11978);
buf BUF1 (N15477, N15446);
nand NAND3 (N15478, N15463, N13072, N9435);
nor NOR4 (N15479, N15468, N10221, N5860, N10902);
or OR4 (N15480, N15479, N799, N11687, N12217);
or OR4 (N15481, N15475, N7871, N3453, N8651);
xor XOR2 (N15482, N15474, N10333);
nand NAND2 (N15483, N15450, N6836);
nor NOR3 (N15484, N15482, N5963, N3569);
and AND3 (N15485, N15469, N13110, N13208);
and AND4 (N15486, N15476, N11857, N10406, N13160);
nor NOR2 (N15487, N15486, N1573);
not NOT1 (N15488, N15481);
buf BUF1 (N15489, N15485);
and AND3 (N15490, N15483, N376, N7143);
nand NAND4 (N15491, N15489, N3317, N3981, N12889);
xor XOR2 (N15492, N15480, N11773);
nand NAND2 (N15493, N15491, N9132);
nand NAND3 (N15494, N15477, N12958, N9337);
or OR2 (N15495, N15492, N12389);
not NOT1 (N15496, N15493);
xor XOR2 (N15497, N15487, N5313);
nor NOR4 (N15498, N15478, N3684, N8087, N6597);
or OR3 (N15499, N15496, N454, N2849);
xor XOR2 (N15500, N15495, N9706);
xor XOR2 (N15501, N15500, N5424);
not NOT1 (N15502, N15497);
not NOT1 (N15503, N15472);
not NOT1 (N15504, N15502);
and AND3 (N15505, N15499, N2747, N2609);
and AND2 (N15506, N15484, N6409);
xor XOR2 (N15507, N15503, N661);
nor NOR3 (N15508, N15494, N12457, N4100);
or OR3 (N15509, N15498, N6297, N13747);
and AND4 (N15510, N15505, N12610, N10141, N12929);
xor XOR2 (N15511, N15501, N12676);
buf BUF1 (N15512, N15508);
or OR4 (N15513, N15470, N8408, N7978, N10335);
buf BUF1 (N15514, N15509);
nand NAND3 (N15515, N15514, N13412, N13709);
xor XOR2 (N15516, N15515, N2768);
xor XOR2 (N15517, N15516, N10211);
xor XOR2 (N15518, N15490, N7943);
or OR3 (N15519, N15488, N8799, N13341);
nor NOR2 (N15520, N15511, N3715);
or OR4 (N15521, N15517, N1847, N4074, N12127);
and AND2 (N15522, N15518, N5463);
buf BUF1 (N15523, N15513);
or OR3 (N15524, N15504, N11730, N4073);
nor NOR4 (N15525, N15510, N12535, N13796, N13263);
buf BUF1 (N15526, N15519);
nor NOR3 (N15527, N15524, N3287, N7158);
nand NAND3 (N15528, N15521, N9685, N7494);
and AND3 (N15529, N15512, N13784, N3143);
and AND3 (N15530, N15525, N4092, N10373);
xor XOR2 (N15531, N15526, N14768);
xor XOR2 (N15532, N15530, N6465);
nand NAND2 (N15533, N15506, N10226);
or OR2 (N15534, N15533, N9007);
nor NOR4 (N15535, N15520, N13964, N111, N3689);
xor XOR2 (N15536, N15507, N12303);
nand NAND4 (N15537, N15535, N3752, N10843, N9937);
xor XOR2 (N15538, N15532, N5421);
nand NAND3 (N15539, N15523, N9529, N8824);
nand NAND3 (N15540, N15536, N5253, N2789);
or OR2 (N15541, N15539, N12099);
buf BUF1 (N15542, N15527);
or OR3 (N15543, N15541, N9232, N10356);
or OR4 (N15544, N15538, N13437, N7867, N2829);
buf BUF1 (N15545, N15531);
nor NOR4 (N15546, N15543, N15052, N12947, N8006);
xor XOR2 (N15547, N15540, N7739);
xor XOR2 (N15548, N15544, N3923);
nand NAND3 (N15549, N15545, N8664, N5562);
or OR2 (N15550, N15529, N12735);
xor XOR2 (N15551, N15542, N12094);
or OR2 (N15552, N15549, N14589);
nand NAND3 (N15553, N15522, N2439, N9275);
nor NOR4 (N15554, N15537, N339, N5595, N10715);
not NOT1 (N15555, N15553);
and AND2 (N15556, N15528, N13903);
and AND2 (N15557, N15552, N11227);
nor NOR3 (N15558, N15548, N8341, N10338);
nand NAND2 (N15559, N15555, N3647);
or OR4 (N15560, N15534, N13912, N13890, N5573);
nor NOR2 (N15561, N15547, N4920);
nor NOR2 (N15562, N15550, N9760);
xor XOR2 (N15563, N15559, N11193);
and AND3 (N15564, N15558, N15448, N5414);
nor NOR2 (N15565, N15564, N12707);
nor NOR3 (N15566, N15565, N5061, N10629);
nand NAND2 (N15567, N15561, N246);
xor XOR2 (N15568, N15562, N9014);
xor XOR2 (N15569, N15568, N284);
nor NOR3 (N15570, N15556, N5905, N739);
or OR2 (N15571, N15563, N13591);
not NOT1 (N15572, N15571);
nor NOR2 (N15573, N15546, N718);
xor XOR2 (N15574, N15557, N2716);
and AND3 (N15575, N15569, N2593, N15197);
nor NOR4 (N15576, N15567, N3407, N8694, N4803);
nand NAND3 (N15577, N15575, N729, N8046);
buf BUF1 (N15578, N15560);
nand NAND4 (N15579, N15577, N4514, N15460, N9261);
not NOT1 (N15580, N15576);
nand NAND4 (N15581, N15554, N2839, N264, N9564);
nand NAND2 (N15582, N15566, N11296);
buf BUF1 (N15583, N15570);
not NOT1 (N15584, N15583);
or OR3 (N15585, N15581, N9401, N5606);
xor XOR2 (N15586, N15584, N12353);
and AND2 (N15587, N15586, N3514);
buf BUF1 (N15588, N15572);
not NOT1 (N15589, N15582);
nand NAND2 (N15590, N15579, N5909);
nor NOR2 (N15591, N15578, N10143);
nor NOR3 (N15592, N15585, N359, N2464);
and AND4 (N15593, N15580, N15177, N7883, N13142);
nor NOR2 (N15594, N15588, N4247);
nor NOR2 (N15595, N15592, N808);
or OR2 (N15596, N15595, N11697);
and AND2 (N15597, N15574, N6945);
or OR2 (N15598, N15591, N3261);
buf BUF1 (N15599, N15593);
or OR2 (N15600, N15589, N8098);
buf BUF1 (N15601, N15598);
and AND3 (N15602, N15551, N755, N108);
not NOT1 (N15603, N15594);
buf BUF1 (N15604, N15599);
xor XOR2 (N15605, N15602, N279);
not NOT1 (N15606, N15601);
buf BUF1 (N15607, N15600);
not NOT1 (N15608, N15604);
not NOT1 (N15609, N15590);
buf BUF1 (N15610, N15596);
nand NAND4 (N15611, N15587, N12228, N2253, N8432);
buf BUF1 (N15612, N15610);
buf BUF1 (N15613, N15605);
xor XOR2 (N15614, N15613, N11620);
xor XOR2 (N15615, N15606, N9170);
and AND3 (N15616, N15611, N12762, N4786);
xor XOR2 (N15617, N15609, N627);
buf BUF1 (N15618, N15603);
or OR2 (N15619, N15614, N4382);
and AND4 (N15620, N15597, N4869, N12881, N11263);
not NOT1 (N15621, N15615);
buf BUF1 (N15622, N15607);
or OR2 (N15623, N15620, N12013);
xor XOR2 (N15624, N15608, N2903);
not NOT1 (N15625, N15573);
nand NAND4 (N15626, N15621, N4795, N9815, N15328);
and AND4 (N15627, N15616, N8690, N14630, N5086);
or OR2 (N15628, N15618, N6409);
and AND4 (N15629, N15627, N10194, N10538, N786);
buf BUF1 (N15630, N15623);
xor XOR2 (N15631, N15630, N3071);
or OR4 (N15632, N15612, N3911, N13650, N8083);
nor NOR2 (N15633, N15628, N9133);
nor NOR2 (N15634, N15625, N12895);
nand NAND4 (N15635, N15624, N7263, N2246, N14151);
not NOT1 (N15636, N15634);
nor NOR2 (N15637, N15619, N527);
buf BUF1 (N15638, N15629);
not NOT1 (N15639, N15633);
nand NAND3 (N15640, N15639, N12886, N9257);
or OR2 (N15641, N15632, N8160);
and AND2 (N15642, N15635, N1780);
nor NOR4 (N15643, N15617, N11732, N11803, N4016);
or OR3 (N15644, N15626, N11070, N8271);
or OR3 (N15645, N15622, N15534, N12743);
not NOT1 (N15646, N15631);
nor NOR4 (N15647, N15644, N8242, N10093, N14572);
or OR2 (N15648, N15637, N4193);
or OR2 (N15649, N15642, N6986);
or OR2 (N15650, N15643, N2883);
nor NOR3 (N15651, N15645, N11431, N12818);
nand NAND2 (N15652, N15647, N3436);
nor NOR3 (N15653, N15641, N9520, N13667);
nor NOR3 (N15654, N15648, N9647, N3947);
buf BUF1 (N15655, N15653);
nand NAND4 (N15656, N15649, N3239, N4806, N10029);
nand NAND3 (N15657, N15654, N15147, N2240);
buf BUF1 (N15658, N15656);
buf BUF1 (N15659, N15651);
nor NOR2 (N15660, N15657, N5707);
not NOT1 (N15661, N15652);
xor XOR2 (N15662, N15650, N13691);
or OR2 (N15663, N15661, N12301);
xor XOR2 (N15664, N15638, N9434);
or OR3 (N15665, N15640, N7760, N8112);
or OR3 (N15666, N15636, N3771, N2360);
nor NOR4 (N15667, N15660, N8356, N2369, N14611);
xor XOR2 (N15668, N15662, N4003);
xor XOR2 (N15669, N15655, N12849);
not NOT1 (N15670, N15664);
and AND4 (N15671, N15670, N5587, N9977, N9319);
buf BUF1 (N15672, N15646);
nor NOR3 (N15673, N15659, N8013, N7398);
and AND3 (N15674, N15665, N8212, N11373);
and AND3 (N15675, N15663, N15174, N13324);
xor XOR2 (N15676, N15674, N4308);
buf BUF1 (N15677, N15669);
not NOT1 (N15678, N15671);
not NOT1 (N15679, N15673);
not NOT1 (N15680, N15666);
or OR3 (N15681, N15677, N10445, N11878);
or OR4 (N15682, N15676, N8324, N4726, N11373);
not NOT1 (N15683, N15668);
not NOT1 (N15684, N15679);
nor NOR3 (N15685, N15680, N3879, N6966);
and AND3 (N15686, N15678, N4872, N2989);
xor XOR2 (N15687, N15675, N7799);
nor NOR4 (N15688, N15658, N12981, N5710, N8403);
nand NAND3 (N15689, N15667, N9425, N7401);
and AND3 (N15690, N15686, N6260, N9689);
nand NAND2 (N15691, N15682, N5261);
nor NOR4 (N15692, N15689, N10881, N10622, N452);
nand NAND3 (N15693, N15690, N13911, N6173);
nor NOR2 (N15694, N15692, N13571);
and AND4 (N15695, N15684, N3514, N13063, N978);
buf BUF1 (N15696, N15693);
not NOT1 (N15697, N15691);
and AND4 (N15698, N15672, N9311, N7581, N1089);
or OR3 (N15699, N15683, N13692, N8948);
or OR4 (N15700, N15699, N468, N1426, N11692);
or OR3 (N15701, N15695, N2298, N224);
xor XOR2 (N15702, N15694, N8976);
or OR4 (N15703, N15702, N8228, N11914, N4572);
xor XOR2 (N15704, N15685, N10239);
not NOT1 (N15705, N15696);
and AND2 (N15706, N15698, N9321);
nand NAND2 (N15707, N15701, N10035);
xor XOR2 (N15708, N15706, N3858);
nor NOR4 (N15709, N15708, N7965, N13231, N725);
not NOT1 (N15710, N15681);
nand NAND2 (N15711, N15703, N3422);
or OR4 (N15712, N15688, N3165, N11540, N7299);
xor XOR2 (N15713, N15705, N15610);
xor XOR2 (N15714, N15687, N2195);
nor NOR2 (N15715, N15707, N5451);
nor NOR4 (N15716, N15704, N14233, N5696, N13342);
nor NOR2 (N15717, N15709, N11819);
not NOT1 (N15718, N15712);
not NOT1 (N15719, N15700);
nor NOR4 (N15720, N15717, N3531, N172, N760);
xor XOR2 (N15721, N15718, N12007);
buf BUF1 (N15722, N15697);
nor NOR4 (N15723, N15721, N9914, N12331, N8703);
and AND3 (N15724, N15714, N10993, N2471);
xor XOR2 (N15725, N15713, N15318);
or OR3 (N15726, N15719, N3479, N4298);
nor NOR4 (N15727, N15715, N15696, N7073, N5902);
and AND2 (N15728, N15726, N11327);
xor XOR2 (N15729, N15724, N4459);
xor XOR2 (N15730, N15711, N1457);
not NOT1 (N15731, N15727);
buf BUF1 (N15732, N15728);
and AND3 (N15733, N15732, N8299, N2953);
or OR3 (N15734, N15730, N14699, N15397);
or OR2 (N15735, N15710, N570);
buf BUF1 (N15736, N15720);
or OR4 (N15737, N15734, N5233, N11555, N8525);
xor XOR2 (N15738, N15737, N1242);
not NOT1 (N15739, N15735);
and AND2 (N15740, N15733, N7006);
nand NAND2 (N15741, N15722, N4663);
and AND4 (N15742, N15731, N12925, N14809, N1280);
not NOT1 (N15743, N15741);
nand NAND3 (N15744, N15725, N6067, N4912);
or OR2 (N15745, N15743, N3869);
nand NAND2 (N15746, N15729, N3527);
not NOT1 (N15747, N15742);
and AND2 (N15748, N15744, N11593);
nand NAND2 (N15749, N15736, N10866);
not NOT1 (N15750, N15739);
and AND2 (N15751, N15740, N2249);
or OR3 (N15752, N15716, N12436, N10304);
buf BUF1 (N15753, N15750);
nor NOR4 (N15754, N15753, N11731, N271, N2318);
xor XOR2 (N15755, N15748, N5105);
and AND2 (N15756, N15746, N1431);
xor XOR2 (N15757, N15751, N2651);
xor XOR2 (N15758, N15747, N6772);
not NOT1 (N15759, N15723);
nand NAND3 (N15760, N15738, N1899, N7516);
xor XOR2 (N15761, N15752, N13188);
not NOT1 (N15762, N15749);
and AND4 (N15763, N15758, N3960, N2419, N2390);
or OR2 (N15764, N15759, N1178);
and AND2 (N15765, N15756, N4703);
not NOT1 (N15766, N15745);
xor XOR2 (N15767, N15765, N14761);
not NOT1 (N15768, N15766);
or OR4 (N15769, N15760, N9866, N11433, N12556);
not NOT1 (N15770, N15767);
nor NOR2 (N15771, N15763, N8856);
nand NAND4 (N15772, N15755, N1304, N2782, N578);
nor NOR2 (N15773, N15768, N5714);
nor NOR3 (N15774, N15772, N1370, N9192);
nand NAND3 (N15775, N15761, N10436, N11651);
nand NAND3 (N15776, N15770, N13020, N10200);
and AND3 (N15777, N15757, N3818, N9800);
nand NAND3 (N15778, N15754, N15435, N8396);
nor NOR3 (N15779, N15775, N12320, N8864);
or OR3 (N15780, N15778, N312, N3667);
not NOT1 (N15781, N15773);
nand NAND4 (N15782, N15776, N9484, N11932, N4798);
or OR2 (N15783, N15769, N6438);
not NOT1 (N15784, N15771);
and AND2 (N15785, N15781, N15367);
and AND4 (N15786, N15780, N5939, N5839, N15437);
or OR4 (N15787, N15762, N14170, N9299, N13790);
xor XOR2 (N15788, N15764, N14576);
or OR3 (N15789, N15787, N10073, N7543);
or OR2 (N15790, N15789, N8536);
or OR4 (N15791, N15779, N15283, N14881, N13117);
buf BUF1 (N15792, N15782);
not NOT1 (N15793, N15792);
not NOT1 (N15794, N15777);
nor NOR2 (N15795, N15788, N108);
not NOT1 (N15796, N15791);
not NOT1 (N15797, N15785);
or OR2 (N15798, N15786, N10446);
not NOT1 (N15799, N15774);
nand NAND3 (N15800, N15795, N14153, N9537);
not NOT1 (N15801, N15783);
buf BUF1 (N15802, N15801);
and AND2 (N15803, N15800, N10247);
nor NOR3 (N15804, N15802, N6844, N2784);
nor NOR2 (N15805, N15794, N12245);
xor XOR2 (N15806, N15797, N5913);
or OR2 (N15807, N15804, N11116);
nand NAND2 (N15808, N15784, N6238);
not NOT1 (N15809, N15790);
nand NAND4 (N15810, N15793, N12862, N2962, N768);
xor XOR2 (N15811, N15809, N10471);
and AND4 (N15812, N15805, N12966, N1870, N3918);
buf BUF1 (N15813, N15807);
not NOT1 (N15814, N15798);
buf BUF1 (N15815, N15811);
xor XOR2 (N15816, N15808, N11502);
buf BUF1 (N15817, N15806);
nor NOR3 (N15818, N15810, N15193, N14801);
xor XOR2 (N15819, N15812, N351);
not NOT1 (N15820, N15818);
and AND2 (N15821, N15820, N5755);
and AND2 (N15822, N15817, N1029);
nor NOR2 (N15823, N15814, N2038);
buf BUF1 (N15824, N15816);
buf BUF1 (N15825, N15815);
buf BUF1 (N15826, N15813);
or OR2 (N15827, N15799, N4782);
buf BUF1 (N15828, N15826);
not NOT1 (N15829, N15824);
buf BUF1 (N15830, N15825);
not NOT1 (N15831, N15830);
not NOT1 (N15832, N15822);
nand NAND4 (N15833, N15823, N4620, N11825, N1678);
nor NOR4 (N15834, N15829, N11898, N6585, N11143);
xor XOR2 (N15835, N15833, N9293);
or OR3 (N15836, N15831, N8267, N8157);
nand NAND3 (N15837, N15796, N5961, N5894);
or OR2 (N15838, N15836, N15711);
nor NOR4 (N15839, N15832, N13305, N11884, N14355);
buf BUF1 (N15840, N15838);
nand NAND2 (N15841, N15803, N7107);
nor NOR4 (N15842, N15821, N14917, N7638, N4962);
nor NOR3 (N15843, N15834, N10290, N9432);
nor NOR4 (N15844, N15843, N8721, N7936, N14156);
or OR4 (N15845, N15840, N4787, N12050, N868);
nand NAND3 (N15846, N15842, N977, N11790);
or OR2 (N15847, N15837, N11050);
or OR3 (N15848, N15844, N861, N8567);
or OR3 (N15849, N15841, N11083, N9403);
nand NAND2 (N15850, N15819, N509);
nand NAND3 (N15851, N15845, N6498, N11119);
not NOT1 (N15852, N15835);
xor XOR2 (N15853, N15851, N5895);
and AND2 (N15854, N15853, N4264);
and AND2 (N15855, N15847, N1509);
xor XOR2 (N15856, N15850, N3007);
nor NOR3 (N15857, N15827, N3013, N6882);
or OR2 (N15858, N15828, N13445);
and AND4 (N15859, N15855, N9863, N15222, N4374);
buf BUF1 (N15860, N15848);
buf BUF1 (N15861, N15858);
and AND3 (N15862, N15852, N11166, N7927);
xor XOR2 (N15863, N15860, N13301);
and AND2 (N15864, N15857, N6390);
and AND2 (N15865, N15861, N13634);
xor XOR2 (N15866, N15863, N6406);
nand NAND4 (N15867, N15856, N1715, N404, N12462);
nand NAND2 (N15868, N15859, N8487);
nand NAND2 (N15869, N15868, N3857);
or OR2 (N15870, N15864, N12434);
xor XOR2 (N15871, N15849, N8212);
nor NOR4 (N15872, N15867, N1329, N3746, N103);
and AND2 (N15873, N15846, N13541);
nor NOR2 (N15874, N15862, N13332);
xor XOR2 (N15875, N15839, N8846);
or OR2 (N15876, N15872, N6490);
or OR2 (N15877, N15873, N7666);
not NOT1 (N15878, N15866);
buf BUF1 (N15879, N15876);
not NOT1 (N15880, N15879);
or OR4 (N15881, N15870, N14235, N7157, N12302);
xor XOR2 (N15882, N15854, N6838);
and AND4 (N15883, N15869, N6306, N12455, N1941);
and AND4 (N15884, N15880, N14832, N13250, N1224);
and AND4 (N15885, N15865, N10762, N5347, N6230);
buf BUF1 (N15886, N15875);
or OR2 (N15887, N15877, N7529);
and AND2 (N15888, N15885, N9043);
buf BUF1 (N15889, N15882);
buf BUF1 (N15890, N15878);
or OR2 (N15891, N15883, N12002);
nor NOR3 (N15892, N15881, N12933, N2328);
nor NOR3 (N15893, N15892, N3466, N3837);
nor NOR3 (N15894, N15884, N2799, N6498);
xor XOR2 (N15895, N15871, N6619);
and AND2 (N15896, N15895, N7216);
not NOT1 (N15897, N15888);
nand NAND2 (N15898, N15887, N14404);
nand NAND4 (N15899, N15896, N15267, N12689, N9666);
or OR2 (N15900, N15874, N8371);
nor NOR3 (N15901, N15890, N9994, N15829);
or OR3 (N15902, N15891, N251, N182);
or OR2 (N15903, N15889, N1081);
or OR2 (N15904, N15886, N1948);
nor NOR2 (N15905, N15902, N8063);
xor XOR2 (N15906, N15899, N8991);
buf BUF1 (N15907, N15901);
not NOT1 (N15908, N15894);
buf BUF1 (N15909, N15893);
buf BUF1 (N15910, N15904);
not NOT1 (N15911, N15907);
not NOT1 (N15912, N15909);
xor XOR2 (N15913, N15900, N855);
xor XOR2 (N15914, N15905, N1227);
buf BUF1 (N15915, N15897);
buf BUF1 (N15916, N15915);
xor XOR2 (N15917, N15913, N13685);
and AND3 (N15918, N15906, N9718, N1046);
xor XOR2 (N15919, N15917, N9910);
or OR2 (N15920, N15918, N5884);
nand NAND2 (N15921, N15912, N3470);
nand NAND4 (N15922, N15919, N5075, N9044, N12802);
nor NOR2 (N15923, N15922, N8625);
or OR2 (N15924, N15910, N5261);
nand NAND4 (N15925, N15921, N5713, N761, N11244);
nor NOR4 (N15926, N15914, N13864, N12533, N1512);
xor XOR2 (N15927, N15916, N12840);
and AND4 (N15928, N15911, N2528, N4392, N9081);
not NOT1 (N15929, N15923);
buf BUF1 (N15930, N15925);
nor NOR4 (N15931, N15920, N3962, N268, N10463);
not NOT1 (N15932, N15928);
not NOT1 (N15933, N15924);
nor NOR4 (N15934, N15927, N8769, N14476, N13652);
or OR2 (N15935, N15929, N8009);
and AND4 (N15936, N15935, N1271, N13831, N1711);
nor NOR4 (N15937, N15930, N4743, N2899, N6114);
nand NAND2 (N15938, N15926, N8695);
not NOT1 (N15939, N15934);
and AND3 (N15940, N15939, N12621, N5508);
nand NAND3 (N15941, N15903, N11250, N11903);
buf BUF1 (N15942, N15898);
not NOT1 (N15943, N15933);
buf BUF1 (N15944, N15908);
nor NOR4 (N15945, N15938, N2045, N6169, N13969);
nor NOR4 (N15946, N15942, N1592, N15597, N8148);
not NOT1 (N15947, N15946);
nand NAND3 (N15948, N15944, N8602, N7638);
buf BUF1 (N15949, N15948);
xor XOR2 (N15950, N15932, N13947);
xor XOR2 (N15951, N15950, N4214);
buf BUF1 (N15952, N15941);
and AND4 (N15953, N15937, N11788, N10851, N4557);
or OR2 (N15954, N15949, N120);
nor NOR4 (N15955, N15952, N3603, N12267, N4080);
or OR3 (N15956, N15936, N11306, N3896);
nand NAND4 (N15957, N15951, N10413, N12206, N3165);
not NOT1 (N15958, N15945);
buf BUF1 (N15959, N15958);
not NOT1 (N15960, N15959);
and AND4 (N15961, N15953, N5017, N6060, N9487);
nand NAND4 (N15962, N15957, N7631, N14710, N976);
not NOT1 (N15963, N15962);
or OR2 (N15964, N15960, N14275);
and AND3 (N15965, N15954, N5747, N7748);
buf BUF1 (N15966, N15963);
or OR3 (N15967, N15943, N6223, N1365);
not NOT1 (N15968, N15966);
xor XOR2 (N15969, N15961, N1015);
nor NOR3 (N15970, N15967, N6851, N15171);
nor NOR3 (N15971, N15931, N12118, N14990);
buf BUF1 (N15972, N15947);
and AND2 (N15973, N15964, N11407);
or OR4 (N15974, N15968, N10221, N4789, N5199);
xor XOR2 (N15975, N15969, N8984);
buf BUF1 (N15976, N15940);
buf BUF1 (N15977, N15975);
buf BUF1 (N15978, N15977);
not NOT1 (N15979, N15976);
nand NAND4 (N15980, N15970, N13100, N2979, N6580);
and AND2 (N15981, N15973, N2581);
xor XOR2 (N15982, N15965, N6959);
and AND4 (N15983, N15980, N7894, N7966, N12745);
nand NAND4 (N15984, N15983, N172, N13180, N9080);
nor NOR2 (N15985, N15956, N7032);
or OR2 (N15986, N15984, N13444);
and AND4 (N15987, N15979, N3970, N3216, N12250);
xor XOR2 (N15988, N15981, N3838);
or OR2 (N15989, N15971, N8785);
xor XOR2 (N15990, N15955, N8689);
xor XOR2 (N15991, N15972, N9543);
or OR4 (N15992, N15978, N12415, N6636, N1782);
xor XOR2 (N15993, N15989, N4973);
xor XOR2 (N15994, N15993, N15361);
and AND3 (N15995, N15990, N4203, N3803);
or OR3 (N15996, N15988, N6893, N360);
and AND2 (N15997, N15991, N4753);
buf BUF1 (N15998, N15995);
nor NOR3 (N15999, N15982, N7840, N12460);
and AND2 (N16000, N15999, N14621);
or OR4 (N16001, N15998, N8994, N1230, N4544);
xor XOR2 (N16002, N15997, N1552);
or OR2 (N16003, N15992, N3444);
buf BUF1 (N16004, N15996);
not NOT1 (N16005, N15994);
or OR3 (N16006, N15985, N12589, N8838);
nor NOR4 (N16007, N16002, N5945, N13504, N3541);
nand NAND4 (N16008, N15986, N6091, N5749, N139);
buf BUF1 (N16009, N16006);
buf BUF1 (N16010, N16001);
or OR3 (N16011, N16005, N297, N4946);
nand NAND3 (N16012, N16007, N3045, N5541);
or OR2 (N16013, N16004, N2004);
and AND2 (N16014, N16010, N12253);
xor XOR2 (N16015, N16009, N654);
nand NAND2 (N16016, N16012, N4588);
nor NOR2 (N16017, N15987, N4000);
not NOT1 (N16018, N16011);
buf BUF1 (N16019, N16013);
nor NOR4 (N16020, N16008, N15906, N13799, N11761);
xor XOR2 (N16021, N16000, N4646);
nand NAND3 (N16022, N16003, N9009, N6019);
not NOT1 (N16023, N16014);
buf BUF1 (N16024, N16016);
not NOT1 (N16025, N16017);
nand NAND4 (N16026, N16024, N12699, N8269, N7345);
nand NAND2 (N16027, N16026, N9303);
buf BUF1 (N16028, N16019);
and AND2 (N16029, N16025, N14623);
xor XOR2 (N16030, N16021, N14099);
nor NOR3 (N16031, N16023, N13038, N7185);
xor XOR2 (N16032, N16020, N7121);
nor NOR4 (N16033, N16031, N14173, N14646, N736);
or OR4 (N16034, N16015, N2781, N1864, N15139);
nor NOR2 (N16035, N16033, N1396);
nand NAND2 (N16036, N16030, N356);
or OR2 (N16037, N16029, N12073);
nand NAND2 (N16038, N16036, N1957);
not NOT1 (N16039, N16038);
buf BUF1 (N16040, N16035);
buf BUF1 (N16041, N16037);
or OR2 (N16042, N16018, N5391);
not NOT1 (N16043, N16039);
nand NAND4 (N16044, N15974, N14396, N9112, N15703);
or OR2 (N16045, N16042, N3597);
nand NAND3 (N16046, N16032, N1381, N8365);
and AND3 (N16047, N16040, N9713, N14470);
not NOT1 (N16048, N16046);
nand NAND2 (N16049, N16048, N5625);
buf BUF1 (N16050, N16027);
not NOT1 (N16051, N16041);
xor XOR2 (N16052, N16028, N1874);
or OR4 (N16053, N16050, N11284, N6879, N8317);
and AND4 (N16054, N16044, N7174, N3558, N12239);
or OR2 (N16055, N16054, N4621);
nor NOR4 (N16056, N16051, N11412, N14237, N3648);
and AND4 (N16057, N16043, N10449, N9517, N804);
not NOT1 (N16058, N16052);
or OR2 (N16059, N16034, N1077);
xor XOR2 (N16060, N16022, N218);
buf BUF1 (N16061, N16058);
xor XOR2 (N16062, N16053, N14373);
nand NAND3 (N16063, N16049, N7079, N2849);
nor NOR2 (N16064, N16055, N2418);
nor NOR2 (N16065, N16045, N2295);
nand NAND2 (N16066, N16059, N3654);
or OR3 (N16067, N16061, N2380, N2003);
nor NOR3 (N16068, N16056, N5976, N8932);
or OR3 (N16069, N16060, N10371, N248);
not NOT1 (N16070, N16057);
nor NOR4 (N16071, N16070, N12659, N15353, N7257);
nand NAND2 (N16072, N16047, N7135);
and AND4 (N16073, N16067, N15179, N13859, N9503);
and AND4 (N16074, N16071, N3731, N14515, N850);
xor XOR2 (N16075, N16074, N15710);
nand NAND4 (N16076, N16065, N4301, N11993, N4543);
xor XOR2 (N16077, N16072, N8174);
nand NAND3 (N16078, N16075, N12634, N6654);
buf BUF1 (N16079, N16078);
or OR3 (N16080, N16077, N1982, N12600);
not NOT1 (N16081, N16073);
xor XOR2 (N16082, N16068, N9428);
nor NOR2 (N16083, N16066, N5046);
nor NOR2 (N16084, N16082, N10072);
and AND3 (N16085, N16081, N9907, N15864);
xor XOR2 (N16086, N16084, N4064);
nor NOR3 (N16087, N16076, N7901, N132);
xor XOR2 (N16088, N16087, N15975);
nor NOR2 (N16089, N16086, N15009);
or OR4 (N16090, N16069, N14080, N4805, N12808);
or OR3 (N16091, N16089, N14059, N1879);
or OR4 (N16092, N16063, N11709, N11869, N11080);
or OR3 (N16093, N16079, N15235, N11535);
or OR2 (N16094, N16088, N11619);
buf BUF1 (N16095, N16092);
not NOT1 (N16096, N16062);
xor XOR2 (N16097, N16095, N9311);
or OR4 (N16098, N16080, N1556, N13571, N14603);
nand NAND4 (N16099, N16098, N6274, N13728, N7270);
xor XOR2 (N16100, N16097, N4939);
or OR2 (N16101, N16100, N10249);
or OR2 (N16102, N16099, N8772);
buf BUF1 (N16103, N16093);
xor XOR2 (N16104, N16103, N9833);
nand NAND2 (N16105, N16083, N610);
and AND3 (N16106, N16101, N10197, N2306);
and AND4 (N16107, N16102, N5315, N6014, N14808);
nor NOR2 (N16108, N16105, N7642);
and AND4 (N16109, N16090, N9035, N1272, N2386);
nand NAND4 (N16110, N16104, N12641, N12933, N12268);
buf BUF1 (N16111, N16064);
not NOT1 (N16112, N16094);
nand NAND2 (N16113, N16109, N12927);
and AND2 (N16114, N16107, N5497);
or OR3 (N16115, N16085, N49, N11337);
nor NOR2 (N16116, N16096, N9265);
nor NOR2 (N16117, N16091, N11011);
nand NAND4 (N16118, N16108, N3873, N13284, N12958);
buf BUF1 (N16119, N16118);
buf BUF1 (N16120, N16110);
nand NAND2 (N16121, N16115, N1791);
and AND2 (N16122, N16112, N546);
nor NOR4 (N16123, N16122, N6472, N13294, N14564);
not NOT1 (N16124, N16111);
or OR2 (N16125, N16116, N6422);
xor XOR2 (N16126, N16117, N5824);
nand NAND4 (N16127, N16120, N1796, N11910, N11709);
buf BUF1 (N16128, N16121);
or OR3 (N16129, N16128, N8954, N4137);
or OR4 (N16130, N16106, N10317, N6991, N3580);
xor XOR2 (N16131, N16125, N5611);
not NOT1 (N16132, N16126);
nand NAND2 (N16133, N16130, N11349);
and AND4 (N16134, N16124, N8545, N13480, N218);
nor NOR2 (N16135, N16123, N8882);
nor NOR2 (N16136, N16129, N14377);
or OR4 (N16137, N16131, N1039, N11743, N9306);
nor NOR2 (N16138, N16114, N2977);
nand NAND2 (N16139, N16135, N15920);
and AND3 (N16140, N16113, N10334, N8552);
xor XOR2 (N16141, N16127, N1720);
buf BUF1 (N16142, N16119);
buf BUF1 (N16143, N16133);
nor NOR4 (N16144, N16141, N2941, N13756, N14974);
and AND2 (N16145, N16144, N4176);
or OR2 (N16146, N16137, N2332);
nand NAND3 (N16147, N16134, N5043, N4385);
xor XOR2 (N16148, N16146, N15106);
buf BUF1 (N16149, N16143);
and AND2 (N16150, N16132, N86);
nand NAND2 (N16151, N16148, N14505);
not NOT1 (N16152, N16140);
nor NOR4 (N16153, N16138, N3805, N12472, N3513);
nand NAND3 (N16154, N16142, N2697, N15181);
nand NAND4 (N16155, N16145, N9179, N8186, N2415);
nor NOR2 (N16156, N16152, N9571);
nand NAND3 (N16157, N16136, N14305, N12443);
and AND3 (N16158, N16153, N12593, N3982);
and AND4 (N16159, N16154, N8055, N529, N6472);
buf BUF1 (N16160, N16158);
nand NAND2 (N16161, N16159, N13968);
or OR3 (N16162, N16160, N6598, N9842);
and AND2 (N16163, N16147, N14598);
xor XOR2 (N16164, N16162, N15544);
nor NOR3 (N16165, N16150, N1693, N3992);
nand NAND4 (N16166, N16139, N174, N14991, N14417);
nor NOR4 (N16167, N16161, N114, N11522, N1924);
xor XOR2 (N16168, N16166, N9175);
and AND4 (N16169, N16168, N2980, N9996, N2796);
nor NOR4 (N16170, N16163, N15369, N4499, N8910);
and AND3 (N16171, N16169, N14225, N8573);
buf BUF1 (N16172, N16170);
xor XOR2 (N16173, N16165, N11772);
xor XOR2 (N16174, N16155, N5537);
and AND3 (N16175, N16174, N10957, N4276);
nand NAND2 (N16176, N16149, N1945);
nand NAND2 (N16177, N16172, N12175);
or OR3 (N16178, N16156, N15847, N1581);
or OR4 (N16179, N16157, N530, N9732, N7013);
buf BUF1 (N16180, N16173);
not NOT1 (N16181, N16171);
and AND3 (N16182, N16180, N2515, N1072);
buf BUF1 (N16183, N16164);
buf BUF1 (N16184, N16178);
buf BUF1 (N16185, N16151);
xor XOR2 (N16186, N16179, N3000);
and AND3 (N16187, N16167, N8380, N6768);
buf BUF1 (N16188, N16177);
nor NOR2 (N16189, N16187, N14131);
xor XOR2 (N16190, N16186, N12767);
or OR3 (N16191, N16182, N2218, N8934);
xor XOR2 (N16192, N16188, N1215);
or OR2 (N16193, N16192, N7568);
or OR4 (N16194, N16185, N7174, N8628, N8228);
xor XOR2 (N16195, N16181, N3780);
xor XOR2 (N16196, N16184, N15568);
and AND4 (N16197, N16183, N12919, N6193, N3883);
nand NAND3 (N16198, N16197, N12062, N6015);
nor NOR3 (N16199, N16191, N7928, N12257);
nor NOR3 (N16200, N16189, N202, N10459);
nor NOR2 (N16201, N16193, N16000);
or OR4 (N16202, N16195, N8331, N9114, N13798);
nor NOR2 (N16203, N16190, N12845);
and AND4 (N16204, N16200, N10604, N10289, N7448);
and AND2 (N16205, N16203, N7154);
xor XOR2 (N16206, N16194, N10257);
buf BUF1 (N16207, N16201);
xor XOR2 (N16208, N16199, N1500);
buf BUF1 (N16209, N16205);
and AND4 (N16210, N16175, N12398, N1570, N11773);
not NOT1 (N16211, N16210);
not NOT1 (N16212, N16207);
buf BUF1 (N16213, N16198);
buf BUF1 (N16214, N16196);
nand NAND3 (N16215, N16208, N6753, N14766);
nor NOR2 (N16216, N16209, N15302);
nor NOR3 (N16217, N16212, N11615, N14794);
nor NOR4 (N16218, N16211, N7877, N13783, N7970);
nor NOR2 (N16219, N16218, N2499);
and AND4 (N16220, N16204, N13988, N13721, N902);
buf BUF1 (N16221, N16217);
buf BUF1 (N16222, N16219);
buf BUF1 (N16223, N16215);
xor XOR2 (N16224, N16176, N1938);
buf BUF1 (N16225, N16223);
buf BUF1 (N16226, N16214);
or OR2 (N16227, N16202, N7860);
xor XOR2 (N16228, N16216, N4005);
not NOT1 (N16229, N16227);
not NOT1 (N16230, N16206);
or OR3 (N16231, N16226, N16045, N11233);
buf BUF1 (N16232, N16224);
and AND3 (N16233, N16221, N14903, N431);
xor XOR2 (N16234, N16229, N6923);
and AND3 (N16235, N16222, N1564, N13285);
nand NAND2 (N16236, N16231, N5227);
and AND4 (N16237, N16233, N10683, N12613, N6372);
not NOT1 (N16238, N16234);
nor NOR2 (N16239, N16225, N4675);
buf BUF1 (N16240, N16230);
nor NOR4 (N16241, N16237, N14133, N15937, N2832);
or OR2 (N16242, N16241, N6946);
buf BUF1 (N16243, N16213);
nor NOR2 (N16244, N16236, N7144);
nand NAND4 (N16245, N16243, N9007, N4202, N15834);
or OR4 (N16246, N16220, N2091, N3427, N4255);
not NOT1 (N16247, N16240);
and AND4 (N16248, N16245, N4807, N11982, N14736);
nand NAND4 (N16249, N16235, N11670, N11300, N11529);
not NOT1 (N16250, N16239);
nor NOR3 (N16251, N16242, N7126, N9690);
not NOT1 (N16252, N16244);
nand NAND2 (N16253, N16228, N1196);
not NOT1 (N16254, N16232);
or OR3 (N16255, N16251, N14713, N615);
nand NAND3 (N16256, N16248, N13347, N4921);
not NOT1 (N16257, N16250);
or OR3 (N16258, N16256, N12794, N8789);
buf BUF1 (N16259, N16249);
or OR4 (N16260, N16254, N9206, N5650, N4334);
nand NAND3 (N16261, N16255, N11759, N2186);
nor NOR4 (N16262, N16259, N8437, N5578, N13253);
not NOT1 (N16263, N16260);
and AND2 (N16264, N16246, N578);
or OR3 (N16265, N16247, N2752, N14585);
nor NOR3 (N16266, N16261, N5036, N14372);
nor NOR4 (N16267, N16238, N12898, N6632, N16211);
and AND2 (N16268, N16262, N14500);
nand NAND4 (N16269, N16258, N14109, N9144, N13050);
nor NOR2 (N16270, N16268, N3080);
not NOT1 (N16271, N16270);
nor NOR3 (N16272, N16271, N4032, N7465);
xor XOR2 (N16273, N16267, N4579);
and AND3 (N16274, N16272, N13237, N213);
not NOT1 (N16275, N16265);
or OR3 (N16276, N16266, N6436, N7592);
xor XOR2 (N16277, N16264, N9953);
buf BUF1 (N16278, N16263);
and AND4 (N16279, N16252, N3681, N135, N5252);
and AND2 (N16280, N16274, N9278);
buf BUF1 (N16281, N16257);
or OR2 (N16282, N16278, N9166);
buf BUF1 (N16283, N16275);
nor NOR4 (N16284, N16273, N7473, N1614, N7219);
and AND2 (N16285, N16284, N1955);
and AND3 (N16286, N16283, N3243, N2826);
xor XOR2 (N16287, N16280, N14221);
buf BUF1 (N16288, N16286);
not NOT1 (N16289, N16281);
nand NAND4 (N16290, N16282, N10871, N13988, N16120);
or OR2 (N16291, N16287, N8422);
xor XOR2 (N16292, N16269, N9097);
xor XOR2 (N16293, N16291, N2857);
not NOT1 (N16294, N16285);
xor XOR2 (N16295, N16293, N14725);
xor XOR2 (N16296, N16289, N85);
or OR3 (N16297, N16295, N13930, N13930);
nor NOR4 (N16298, N16277, N15585, N13099, N13646);
nand NAND4 (N16299, N16297, N4304, N14373, N10308);
and AND4 (N16300, N16288, N7260, N10304, N7812);
buf BUF1 (N16301, N16294);
and AND4 (N16302, N16299, N7902, N15662, N7540);
buf BUF1 (N16303, N16290);
nor NOR4 (N16304, N16296, N5816, N12531, N15086);
nand NAND4 (N16305, N16276, N11412, N1297, N2729);
not NOT1 (N16306, N16301);
not NOT1 (N16307, N16304);
not NOT1 (N16308, N16292);
xor XOR2 (N16309, N16302, N13352);
nand NAND2 (N16310, N16279, N7676);
or OR3 (N16311, N16310, N16093, N8270);
and AND4 (N16312, N16298, N9339, N515, N15346);
or OR4 (N16313, N16306, N541, N1752, N11801);
buf BUF1 (N16314, N16308);
or OR2 (N16315, N16307, N676);
not NOT1 (N16316, N16312);
nand NAND4 (N16317, N16303, N6337, N3543, N13561);
xor XOR2 (N16318, N16313, N10824);
and AND3 (N16319, N16305, N2311, N5071);
or OR4 (N16320, N16316, N9059, N15365, N9968);
buf BUF1 (N16321, N16300);
xor XOR2 (N16322, N16321, N730);
nand NAND2 (N16323, N16315, N3395);
or OR3 (N16324, N16323, N4869, N2586);
nor NOR3 (N16325, N16253, N14050, N15508);
xor XOR2 (N16326, N16322, N7634);
buf BUF1 (N16327, N16319);
nor NOR3 (N16328, N16327, N52, N2859);
xor XOR2 (N16329, N16320, N7319);
nand NAND4 (N16330, N16325, N5750, N9476, N11223);
and AND2 (N16331, N16317, N13785);
and AND3 (N16332, N16324, N14919, N10473);
buf BUF1 (N16333, N16318);
nor NOR3 (N16334, N16314, N14411, N13127);
nand NAND3 (N16335, N16329, N10621, N7471);
nand NAND4 (N16336, N16332, N1763, N10750, N7488);
not NOT1 (N16337, N16328);
and AND4 (N16338, N16333, N15107, N2908, N8859);
and AND4 (N16339, N16331, N10196, N1669, N7179);
nand NAND2 (N16340, N16335, N5916);
not NOT1 (N16341, N16337);
or OR4 (N16342, N16334, N4901, N9469, N6849);
not NOT1 (N16343, N16340);
and AND2 (N16344, N16336, N9621);
nand NAND4 (N16345, N16311, N1206, N1187, N9280);
or OR3 (N16346, N16345, N1285, N15835);
nor NOR4 (N16347, N16326, N4758, N12411, N324);
nand NAND2 (N16348, N16342, N1433);
xor XOR2 (N16349, N16347, N6364);
and AND3 (N16350, N16339, N10529, N13228);
and AND3 (N16351, N16330, N7679, N15188);
nor NOR3 (N16352, N16348, N10380, N11655);
nand NAND2 (N16353, N16343, N9801);
buf BUF1 (N16354, N16353);
nor NOR2 (N16355, N16346, N6183);
not NOT1 (N16356, N16341);
and AND4 (N16357, N16351, N1578, N7749, N5630);
xor XOR2 (N16358, N16352, N6714);
buf BUF1 (N16359, N16354);
or OR3 (N16360, N16357, N10009, N5850);
not NOT1 (N16361, N16359);
buf BUF1 (N16362, N16350);
nand NAND3 (N16363, N16362, N5695, N12909);
nor NOR2 (N16364, N16355, N12636);
not NOT1 (N16365, N16363);
nand NAND3 (N16366, N16364, N14261, N4741);
nor NOR3 (N16367, N16360, N5936, N4545);
not NOT1 (N16368, N16365);
nor NOR2 (N16369, N16367, N15040);
nand NAND4 (N16370, N16369, N5999, N3287, N11858);
or OR4 (N16371, N16338, N3862, N8266, N7410);
or OR4 (N16372, N16370, N6473, N1805, N8871);
or OR2 (N16373, N16349, N2451);
or OR2 (N16374, N16309, N773);
buf BUF1 (N16375, N16356);
and AND4 (N16376, N16371, N418, N15211, N15617);
xor XOR2 (N16377, N16366, N4861);
nor NOR4 (N16378, N16344, N12704, N3852, N13386);
or OR4 (N16379, N16378, N12942, N7652, N1528);
and AND3 (N16380, N16372, N4210, N11614);
buf BUF1 (N16381, N16373);
nand NAND3 (N16382, N16368, N12981, N2299);
nand NAND2 (N16383, N16376, N13790);
nor NOR3 (N16384, N16375, N8966, N8974);
xor XOR2 (N16385, N16380, N15906);
nor NOR2 (N16386, N16385, N385);
not NOT1 (N16387, N16386);
not NOT1 (N16388, N16361);
nand NAND2 (N16389, N16387, N5727);
and AND4 (N16390, N16381, N14316, N1187, N4959);
nand NAND3 (N16391, N16358, N16034, N14395);
nor NOR2 (N16392, N16374, N3672);
or OR3 (N16393, N16388, N3810, N12540);
not NOT1 (N16394, N16389);
or OR4 (N16395, N16383, N11885, N8835, N13611);
nand NAND2 (N16396, N16384, N11518);
nand NAND3 (N16397, N16392, N5920, N11075);
nor NOR3 (N16398, N16397, N8177, N6955);
xor XOR2 (N16399, N16395, N10874);
not NOT1 (N16400, N16393);
or OR3 (N16401, N16391, N3048, N9994);
buf BUF1 (N16402, N16398);
not NOT1 (N16403, N16382);
xor XOR2 (N16404, N16379, N11190);
not NOT1 (N16405, N16404);
nor NOR2 (N16406, N16377, N9652);
xor XOR2 (N16407, N16390, N2415);
not NOT1 (N16408, N16399);
buf BUF1 (N16409, N16402);
nand NAND3 (N16410, N16394, N4784, N13301);
nand NAND3 (N16411, N16401, N7436, N3973);
nand NAND4 (N16412, N16396, N15271, N13892, N8710);
or OR3 (N16413, N16409, N744, N7229);
buf BUF1 (N16414, N16400);
or OR3 (N16415, N16407, N5354, N12455);
or OR4 (N16416, N16411, N16103, N2976, N7414);
and AND4 (N16417, N16412, N4923, N6390, N9442);
nor NOR3 (N16418, N16403, N3355, N13570);
or OR2 (N16419, N16405, N16285);
xor XOR2 (N16420, N16413, N9780);
xor XOR2 (N16421, N16417, N10670);
nor NOR4 (N16422, N16421, N5724, N379, N11788);
nand NAND3 (N16423, N16408, N4716, N4686);
not NOT1 (N16424, N16420);
xor XOR2 (N16425, N16416, N2628);
nand NAND2 (N16426, N16419, N12214);
not NOT1 (N16427, N16426);
or OR3 (N16428, N16418, N15258, N2416);
and AND4 (N16429, N16422, N8551, N8210, N3042);
and AND4 (N16430, N16425, N4922, N8649, N12107);
buf BUF1 (N16431, N16429);
and AND4 (N16432, N16415, N6069, N4953, N13388);
nor NOR2 (N16433, N16432, N4004);
and AND2 (N16434, N16406, N3967);
or OR4 (N16435, N16410, N11776, N12661, N1179);
nand NAND2 (N16436, N16423, N3299);
or OR4 (N16437, N16436, N2086, N4044, N14761);
or OR4 (N16438, N16424, N6375, N9826, N11783);
xor XOR2 (N16439, N16431, N14034);
xor XOR2 (N16440, N16437, N4438);
xor XOR2 (N16441, N16439, N6138);
nor NOR2 (N16442, N16433, N11587);
xor XOR2 (N16443, N16430, N9375);
or OR3 (N16444, N16438, N166, N1710);
and AND4 (N16445, N16443, N15553, N10081, N14214);
nor NOR3 (N16446, N16445, N2812, N16112);
and AND2 (N16447, N16441, N13948);
nor NOR4 (N16448, N16434, N5605, N15706, N10835);
not NOT1 (N16449, N16427);
not NOT1 (N16450, N16414);
xor XOR2 (N16451, N16448, N9579);
and AND3 (N16452, N16444, N8368, N7052);
or OR4 (N16453, N16447, N4171, N1116, N8753);
and AND3 (N16454, N16428, N15005, N9060);
and AND4 (N16455, N16453, N8468, N4893, N16060);
and AND3 (N16456, N16454, N12284, N11734);
and AND2 (N16457, N16446, N13474);
or OR4 (N16458, N16456, N2063, N4802, N391);
and AND2 (N16459, N16450, N12227);
xor XOR2 (N16460, N16458, N10869);
not NOT1 (N16461, N16452);
not NOT1 (N16462, N16440);
nor NOR4 (N16463, N16459, N6947, N8282, N2195);
buf BUF1 (N16464, N16442);
and AND4 (N16465, N16460, N6594, N12620, N8719);
nor NOR4 (N16466, N16465, N12032, N4543, N6309);
and AND4 (N16467, N16455, N3499, N10065, N10423);
nor NOR2 (N16468, N16435, N5358);
nor NOR2 (N16469, N16451, N6676);
or OR3 (N16470, N16461, N10960, N6300);
not NOT1 (N16471, N16466);
nor NOR4 (N16472, N16470, N13121, N1944, N12290);
xor XOR2 (N16473, N16472, N7076);
not NOT1 (N16474, N16467);
nand NAND4 (N16475, N16449, N8335, N11460, N14589);
and AND2 (N16476, N16474, N16086);
or OR2 (N16477, N16469, N14023);
xor XOR2 (N16478, N16457, N12069);
not NOT1 (N16479, N16473);
xor XOR2 (N16480, N16476, N7898);
buf BUF1 (N16481, N16475);
buf BUF1 (N16482, N16478);
not NOT1 (N16483, N16480);
or OR4 (N16484, N16482, N15642, N9829, N3827);
nand NAND2 (N16485, N16462, N436);
xor XOR2 (N16486, N16463, N13661);
buf BUF1 (N16487, N16479);
or OR2 (N16488, N16468, N12488);
not NOT1 (N16489, N16464);
xor XOR2 (N16490, N16471, N15434);
nor NOR3 (N16491, N16488, N8992, N7598);
xor XOR2 (N16492, N16487, N7738);
nor NOR4 (N16493, N16489, N2373, N8666, N11019);
nor NOR3 (N16494, N16486, N1341, N1124);
xor XOR2 (N16495, N16477, N942);
nor NOR4 (N16496, N16485, N832, N4352, N11862);
and AND2 (N16497, N16495, N7679);
or OR3 (N16498, N16483, N4672, N12321);
nor NOR3 (N16499, N16494, N1489, N15209);
nand NAND3 (N16500, N16498, N6068, N11590);
not NOT1 (N16501, N16492);
and AND4 (N16502, N16493, N8347, N10318, N13286);
xor XOR2 (N16503, N16500, N10819);
xor XOR2 (N16504, N16503, N1125);
or OR3 (N16505, N16496, N2898, N5404);
buf BUF1 (N16506, N16505);
and AND4 (N16507, N16504, N2697, N13367, N2912);
buf BUF1 (N16508, N16507);
xor XOR2 (N16509, N16508, N15206);
and AND3 (N16510, N16506, N14541, N11760);
or OR3 (N16511, N16510, N11079, N13848);
nand NAND3 (N16512, N16499, N15875, N5577);
not NOT1 (N16513, N16481);
nor NOR4 (N16514, N16502, N14826, N11346, N12231);
and AND2 (N16515, N16497, N4207);
buf BUF1 (N16516, N16490);
and AND2 (N16517, N16512, N11446);
nor NOR3 (N16518, N16515, N5765, N11920);
or OR4 (N16519, N16518, N9589, N1381, N11860);
or OR2 (N16520, N16513, N14710);
nor NOR4 (N16521, N16517, N14194, N16281, N11784);
or OR3 (N16522, N16520, N13332, N5534);
nand NAND2 (N16523, N16511, N7971);
or OR3 (N16524, N16519, N407, N3818);
xor XOR2 (N16525, N16522, N13743);
nand NAND3 (N16526, N16491, N9819, N14124);
nand NAND3 (N16527, N16521, N9661, N6543);
buf BUF1 (N16528, N16516);
not NOT1 (N16529, N16526);
nor NOR3 (N16530, N16509, N5471, N1107);
and AND4 (N16531, N16528, N6612, N10021, N12554);
xor XOR2 (N16532, N16524, N4704);
and AND2 (N16533, N16532, N15044);
or OR3 (N16534, N16525, N4705, N10624);
xor XOR2 (N16535, N16523, N5870);
and AND4 (N16536, N16529, N13646, N2130, N3907);
not NOT1 (N16537, N16535);
xor XOR2 (N16538, N16531, N13698);
or OR2 (N16539, N16484, N14423);
not NOT1 (N16540, N16536);
nand NAND2 (N16541, N16527, N1008);
and AND2 (N16542, N16540, N6963);
not NOT1 (N16543, N16542);
or OR3 (N16544, N16543, N1810, N1984);
and AND3 (N16545, N16530, N5308, N13899);
not NOT1 (N16546, N16541);
not NOT1 (N16547, N16534);
buf BUF1 (N16548, N16545);
nand NAND3 (N16549, N16514, N11386, N13452);
xor XOR2 (N16550, N16544, N9128);
xor XOR2 (N16551, N16546, N8912);
nor NOR2 (N16552, N16533, N8222);
xor XOR2 (N16553, N16538, N13924);
or OR3 (N16554, N16547, N2815, N4922);
or OR3 (N16555, N16550, N1666, N11941);
or OR4 (N16556, N16554, N14500, N8823, N2100);
xor XOR2 (N16557, N16501, N8967);
nor NOR3 (N16558, N16557, N11935, N9401);
and AND2 (N16559, N16539, N4917);
nor NOR3 (N16560, N16537, N14579, N9736);
nand NAND4 (N16561, N16549, N6599, N15002, N14855);
xor XOR2 (N16562, N16560, N5447);
buf BUF1 (N16563, N16553);
not NOT1 (N16564, N16551);
nand NAND4 (N16565, N16562, N842, N2245, N1511);
xor XOR2 (N16566, N16556, N13975);
not NOT1 (N16567, N16552);
buf BUF1 (N16568, N16567);
nand NAND2 (N16569, N16564, N6841);
and AND3 (N16570, N16569, N2024, N653);
or OR4 (N16571, N16561, N8753, N5033, N11892);
not NOT1 (N16572, N16563);
and AND4 (N16573, N16566, N1936, N1876, N4602);
buf BUF1 (N16574, N16573);
xor XOR2 (N16575, N16548, N13706);
not NOT1 (N16576, N16571);
or OR4 (N16577, N16570, N2092, N12617, N10754);
buf BUF1 (N16578, N16555);
nor NOR3 (N16579, N16558, N138, N11187);
buf BUF1 (N16580, N16575);
buf BUF1 (N16581, N16576);
nor NOR4 (N16582, N16568, N12259, N3710, N14129);
buf BUF1 (N16583, N16565);
buf BUF1 (N16584, N16574);
nand NAND4 (N16585, N16580, N6807, N1918, N14501);
not NOT1 (N16586, N16584);
not NOT1 (N16587, N16572);
xor XOR2 (N16588, N16583, N7041);
buf BUF1 (N16589, N16578);
and AND3 (N16590, N16577, N9073, N2657);
and AND4 (N16591, N16587, N1520, N11399, N1908);
not NOT1 (N16592, N16559);
not NOT1 (N16593, N16592);
xor XOR2 (N16594, N16582, N14204);
xor XOR2 (N16595, N16586, N12799);
not NOT1 (N16596, N16588);
xor XOR2 (N16597, N16594, N7573);
nand NAND3 (N16598, N16595, N14406, N16002);
and AND3 (N16599, N16581, N14880, N3270);
nor NOR4 (N16600, N16591, N9591, N14725, N3442);
buf BUF1 (N16601, N16597);
buf BUF1 (N16602, N16596);
nand NAND4 (N16603, N16602, N12525, N4409, N9246);
not NOT1 (N16604, N16590);
nor NOR4 (N16605, N16599, N5093, N7980, N5060);
or OR2 (N16606, N16598, N1261);
nor NOR3 (N16607, N16606, N11810, N8956);
and AND4 (N16608, N16603, N14870, N9305, N11060);
and AND4 (N16609, N16585, N6226, N629, N14654);
not NOT1 (N16610, N16600);
or OR2 (N16611, N16610, N7026);
or OR2 (N16612, N16607, N12642);
or OR4 (N16613, N16608, N5098, N10960, N5781);
or OR2 (N16614, N16609, N13964);
nor NOR3 (N16615, N16613, N14315, N4535);
and AND4 (N16616, N16601, N7284, N5048, N4948);
nand NAND3 (N16617, N16605, N12099, N5059);
nor NOR3 (N16618, N16589, N13766, N8729);
xor XOR2 (N16619, N16617, N4828);
xor XOR2 (N16620, N16619, N1737);
xor XOR2 (N16621, N16611, N6776);
not NOT1 (N16622, N16612);
not NOT1 (N16623, N16593);
or OR4 (N16624, N16622, N5957, N4013, N1377);
nand NAND2 (N16625, N16618, N244);
or OR2 (N16626, N16623, N4684);
buf BUF1 (N16627, N16624);
xor XOR2 (N16628, N16615, N11342);
nor NOR3 (N16629, N16627, N8703, N13391);
buf BUF1 (N16630, N16629);
or OR4 (N16631, N16620, N13209, N9859, N16439);
not NOT1 (N16632, N16626);
nand NAND3 (N16633, N16628, N8430, N7232);
xor XOR2 (N16634, N16621, N2630);
xor XOR2 (N16635, N16604, N12656);
or OR2 (N16636, N16630, N1983);
not NOT1 (N16637, N16634);
nor NOR2 (N16638, N16614, N7556);
or OR4 (N16639, N16635, N11243, N14909, N6274);
nand NAND2 (N16640, N16631, N15653);
xor XOR2 (N16641, N16640, N1357);
xor XOR2 (N16642, N16636, N16213);
or OR3 (N16643, N16639, N6715, N14551);
and AND2 (N16644, N16641, N6755);
and AND3 (N16645, N16616, N9729, N15005);
nand NAND2 (N16646, N16643, N12525);
buf BUF1 (N16647, N16642);
xor XOR2 (N16648, N16646, N5337);
xor XOR2 (N16649, N16645, N10529);
nand NAND2 (N16650, N16625, N3210);
and AND3 (N16651, N16649, N338, N7396);
not NOT1 (N16652, N16647);
nor NOR3 (N16653, N16644, N1842, N7020);
nand NAND2 (N16654, N16650, N6432);
xor XOR2 (N16655, N16652, N3116);
nor NOR3 (N16656, N16633, N13276, N9497);
buf BUF1 (N16657, N16654);
nor NOR2 (N16658, N16653, N13853);
nand NAND4 (N16659, N16657, N14214, N6916, N12596);
nand NAND4 (N16660, N16655, N13348, N12945, N16068);
and AND3 (N16661, N16648, N5723, N9894);
or OR4 (N16662, N16651, N8063, N11747, N11992);
buf BUF1 (N16663, N16659);
or OR2 (N16664, N16663, N2106);
xor XOR2 (N16665, N16637, N9258);
nand NAND4 (N16666, N16660, N9099, N6601, N14654);
xor XOR2 (N16667, N16662, N4460);
not NOT1 (N16668, N16638);
nand NAND4 (N16669, N16579, N5812, N6954, N3107);
or OR2 (N16670, N16669, N2573);
nor NOR3 (N16671, N16661, N9991, N10035);
xor XOR2 (N16672, N16656, N130);
buf BUF1 (N16673, N16658);
not NOT1 (N16674, N16670);
xor XOR2 (N16675, N16632, N6501);
buf BUF1 (N16676, N16674);
or OR3 (N16677, N16676, N16168, N12046);
buf BUF1 (N16678, N16677);
or OR2 (N16679, N16668, N9260);
nor NOR3 (N16680, N16679, N16167, N13685);
buf BUF1 (N16681, N16673);
buf BUF1 (N16682, N16666);
or OR4 (N16683, N16678, N5732, N956, N3911);
buf BUF1 (N16684, N16675);
nor NOR3 (N16685, N16667, N7181, N16343);
buf BUF1 (N16686, N16682);
not NOT1 (N16687, N16683);
or OR3 (N16688, N16684, N1411, N8279);
nor NOR3 (N16689, N16671, N4226, N103);
nor NOR4 (N16690, N16689, N9844, N2291, N9621);
nor NOR2 (N16691, N16685, N7044);
nor NOR3 (N16692, N16686, N14521, N9374);
nor NOR4 (N16693, N16692, N4660, N3977, N6010);
and AND2 (N16694, N16672, N8958);
xor XOR2 (N16695, N16680, N15034);
nor NOR2 (N16696, N16694, N11192);
not NOT1 (N16697, N16695);
nor NOR2 (N16698, N16691, N15733);
and AND2 (N16699, N16696, N14520);
not NOT1 (N16700, N16697);
nor NOR3 (N16701, N16681, N1172, N6038);
buf BUF1 (N16702, N16664);
nor NOR4 (N16703, N16702, N2853, N12371, N2015);
and AND4 (N16704, N16701, N13955, N4082, N15346);
nor NOR3 (N16705, N16704, N12822, N4968);
or OR3 (N16706, N16700, N5056, N8520);
and AND4 (N16707, N16706, N1861, N1118, N11590);
xor XOR2 (N16708, N16698, N5787);
buf BUF1 (N16709, N16699);
xor XOR2 (N16710, N16709, N1275);
buf BUF1 (N16711, N16665);
and AND4 (N16712, N16688, N6711, N13079, N7631);
or OR2 (N16713, N16687, N2004);
or OR3 (N16714, N16711, N11383, N2824);
and AND2 (N16715, N16710, N8520);
and AND2 (N16716, N16708, N13862);
and AND3 (N16717, N16716, N7647, N16636);
or OR2 (N16718, N16690, N12725);
nand NAND4 (N16719, N16703, N8827, N12221, N14512);
and AND2 (N16720, N16693, N4626);
buf BUF1 (N16721, N16720);
nor NOR3 (N16722, N16721, N13453, N13838);
or OR4 (N16723, N16714, N5306, N9653, N2175);
and AND3 (N16724, N16722, N1171, N8824);
not NOT1 (N16725, N16719);
and AND3 (N16726, N16717, N12420, N13763);
nand NAND4 (N16727, N16718, N12516, N1344, N2739);
nor NOR3 (N16728, N16713, N354, N4125);
buf BUF1 (N16729, N16715);
xor XOR2 (N16730, N16727, N12371);
xor XOR2 (N16731, N16707, N4160);
not NOT1 (N16732, N16730);
xor XOR2 (N16733, N16724, N8424);
not NOT1 (N16734, N16733);
xor XOR2 (N16735, N16726, N8796);
buf BUF1 (N16736, N16735);
nand NAND2 (N16737, N16734, N10522);
and AND3 (N16738, N16712, N9398, N2477);
nor NOR4 (N16739, N16705, N15671, N6887, N8911);
or OR2 (N16740, N16729, N15803);
buf BUF1 (N16741, N16732);
buf BUF1 (N16742, N16736);
xor XOR2 (N16743, N16731, N7327);
not NOT1 (N16744, N16742);
and AND4 (N16745, N16739, N4772, N1324, N8757);
buf BUF1 (N16746, N16741);
not NOT1 (N16747, N16743);
and AND4 (N16748, N16737, N8217, N6883, N13406);
buf BUF1 (N16749, N16747);
or OR4 (N16750, N16749, N12548, N4411, N11912);
nor NOR4 (N16751, N16738, N12306, N8209, N8862);
and AND3 (N16752, N16728, N16021, N3799);
nand NAND3 (N16753, N16740, N7079, N15358);
nor NOR4 (N16754, N16744, N7462, N5722, N2213);
or OR2 (N16755, N16745, N14462);
nand NAND2 (N16756, N16725, N6751);
nand NAND2 (N16757, N16756, N13951);
nor NOR4 (N16758, N16757, N2007, N3327, N5874);
and AND3 (N16759, N16748, N212, N3383);
not NOT1 (N16760, N16759);
or OR3 (N16761, N16754, N9955, N15233);
or OR3 (N16762, N16746, N477, N6348);
and AND2 (N16763, N16753, N15323);
buf BUF1 (N16764, N16758);
nor NOR3 (N16765, N16723, N5922, N12261);
buf BUF1 (N16766, N16763);
not NOT1 (N16767, N16766);
nor NOR2 (N16768, N16755, N6958);
or OR3 (N16769, N16762, N8233, N1100);
xor XOR2 (N16770, N16750, N4683);
xor XOR2 (N16771, N16764, N7731);
nand NAND2 (N16772, N16771, N367);
nand NAND2 (N16773, N16767, N8316);
nor NOR4 (N16774, N16765, N11268, N13270, N12858);
buf BUF1 (N16775, N16760);
not NOT1 (N16776, N16752);
and AND2 (N16777, N16775, N11113);
xor XOR2 (N16778, N16769, N7804);
not NOT1 (N16779, N16777);
nor NOR4 (N16780, N16768, N9074, N440, N10100);
nor NOR2 (N16781, N16772, N5549);
or OR4 (N16782, N16773, N12917, N37, N14308);
xor XOR2 (N16783, N16781, N6749);
buf BUF1 (N16784, N16782);
xor XOR2 (N16785, N16779, N6748);
buf BUF1 (N16786, N16770);
not NOT1 (N16787, N16784);
xor XOR2 (N16788, N16780, N15158);
nand NAND4 (N16789, N16761, N2773, N13028, N3823);
or OR3 (N16790, N16776, N12845, N12065);
buf BUF1 (N16791, N16774);
and AND4 (N16792, N16788, N1006, N3285, N12053);
xor XOR2 (N16793, N16787, N14926);
or OR4 (N16794, N16789, N4733, N10792, N9547);
or OR3 (N16795, N16793, N10921, N8572);
and AND4 (N16796, N16791, N11703, N6741, N12538);
or OR2 (N16797, N16795, N14145);
and AND3 (N16798, N16794, N2298, N2793);
xor XOR2 (N16799, N16783, N14563);
buf BUF1 (N16800, N16797);
xor XOR2 (N16801, N16796, N10416);
not NOT1 (N16802, N16800);
and AND4 (N16803, N16802, N8000, N12667, N5628);
not NOT1 (N16804, N16751);
nand NAND4 (N16805, N16778, N5130, N9157, N9673);
nor NOR3 (N16806, N16799, N11545, N1203);
nor NOR4 (N16807, N16798, N11326, N9706, N16425);
nor NOR2 (N16808, N16807, N7753);
and AND3 (N16809, N16808, N3226, N10213);
buf BUF1 (N16810, N16786);
or OR4 (N16811, N16801, N6011, N13247, N3461);
and AND2 (N16812, N16811, N15555);
nor NOR4 (N16813, N16785, N13914, N11388, N9591);
nand NAND4 (N16814, N16810, N12644, N8335, N11418);
nand NAND4 (N16815, N16813, N10850, N9039, N15476);
nor NOR2 (N16816, N16790, N7857);
nor NOR2 (N16817, N16809, N2333);
not NOT1 (N16818, N16805);
xor XOR2 (N16819, N16818, N5983);
xor XOR2 (N16820, N16816, N3873);
not NOT1 (N16821, N16814);
nand NAND3 (N16822, N16815, N6626, N5677);
not NOT1 (N16823, N16803);
nor NOR4 (N16824, N16819, N16437, N8577, N16191);
and AND4 (N16825, N16792, N13150, N4444, N13935);
not NOT1 (N16826, N16823);
nand NAND3 (N16827, N16804, N7095, N9520);
and AND4 (N16828, N16817, N9738, N3129, N4920);
nand NAND4 (N16829, N16822, N3480, N3593, N600);
nor NOR3 (N16830, N16825, N16221, N11798);
buf BUF1 (N16831, N16826);
nand NAND4 (N16832, N16820, N12608, N3017, N3449);
xor XOR2 (N16833, N16828, N6374);
and AND4 (N16834, N16812, N15127, N7666, N2940);
buf BUF1 (N16835, N16833);
buf BUF1 (N16836, N16830);
nor NOR2 (N16837, N16835, N14484);
nand NAND2 (N16838, N16824, N10950);
xor XOR2 (N16839, N16834, N14758);
not NOT1 (N16840, N16831);
not NOT1 (N16841, N16840);
xor XOR2 (N16842, N16806, N3549);
or OR2 (N16843, N16838, N11569);
nand NAND4 (N16844, N16821, N4764, N4656, N16001);
buf BUF1 (N16845, N16843);
nor NOR2 (N16846, N16839, N13668);
buf BUF1 (N16847, N16827);
nand NAND4 (N16848, N16844, N13674, N9221, N2167);
nor NOR3 (N16849, N16842, N14232, N3306);
not NOT1 (N16850, N16829);
nand NAND3 (N16851, N16841, N13865, N2462);
buf BUF1 (N16852, N16848);
or OR3 (N16853, N16837, N8120, N9207);
not NOT1 (N16854, N16847);
not NOT1 (N16855, N16852);
and AND2 (N16856, N16853, N5008);
nor NOR2 (N16857, N16845, N10922);
nor NOR2 (N16858, N16846, N4794);
buf BUF1 (N16859, N16857);
not NOT1 (N16860, N16836);
and AND3 (N16861, N16855, N3342, N517);
buf BUF1 (N16862, N16859);
and AND4 (N16863, N16861, N10442, N1889, N4112);
not NOT1 (N16864, N16832);
xor XOR2 (N16865, N16854, N6507);
not NOT1 (N16866, N16858);
nand NAND2 (N16867, N16862, N3002);
and AND3 (N16868, N16864, N11923, N333);
nand NAND2 (N16869, N16865, N1476);
and AND2 (N16870, N16851, N1963);
not NOT1 (N16871, N16860);
nand NAND2 (N16872, N16870, N14719);
nand NAND4 (N16873, N16869, N12914, N3790, N6263);
and AND4 (N16874, N16850, N11082, N2058, N5329);
nand NAND3 (N16875, N16849, N10831, N12683);
not NOT1 (N16876, N16875);
and AND2 (N16877, N16871, N13237);
or OR4 (N16878, N16872, N9549, N4828, N12318);
and AND3 (N16879, N16878, N1316, N8821);
not NOT1 (N16880, N16874);
or OR3 (N16881, N16866, N13323, N16384);
buf BUF1 (N16882, N16873);
xor XOR2 (N16883, N16881, N10173);
and AND3 (N16884, N16883, N2834, N15998);
buf BUF1 (N16885, N16856);
not NOT1 (N16886, N16863);
nor NOR4 (N16887, N16879, N3017, N228, N14707);
nand NAND4 (N16888, N16867, N7429, N5755, N8624);
buf BUF1 (N16889, N16887);
or OR4 (N16890, N16876, N15380, N11347, N11760);
not NOT1 (N16891, N16889);
nand NAND4 (N16892, N16880, N9333, N9197, N10324);
and AND3 (N16893, N16888, N5089, N1032);
not NOT1 (N16894, N16884);
nand NAND2 (N16895, N16868, N13766);
or OR3 (N16896, N16894, N636, N14283);
and AND3 (N16897, N16895, N10705, N15623);
buf BUF1 (N16898, N16877);
not NOT1 (N16899, N16886);
or OR3 (N16900, N16892, N11190, N995);
not NOT1 (N16901, N16899);
nor NOR2 (N16902, N16882, N2376);
nand NAND4 (N16903, N16897, N14219, N2344, N7404);
not NOT1 (N16904, N16898);
not NOT1 (N16905, N16902);
and AND2 (N16906, N16890, N1511);
nor NOR2 (N16907, N16904, N12258);
buf BUF1 (N16908, N16900);
buf BUF1 (N16909, N16896);
or OR2 (N16910, N16907, N11753);
nand NAND2 (N16911, N16903, N12902);
buf BUF1 (N16912, N16906);
or OR2 (N16913, N16908, N15365);
nor NOR4 (N16914, N16913, N3934, N1026, N4208);
not NOT1 (N16915, N16905);
not NOT1 (N16916, N16891);
and AND2 (N16917, N16915, N11577);
not NOT1 (N16918, N16917);
nor NOR2 (N16919, N16910, N13221);
not NOT1 (N16920, N16914);
buf BUF1 (N16921, N16916);
or OR3 (N16922, N16911, N345, N7696);
and AND4 (N16923, N16919, N10855, N15199, N12818);
nor NOR4 (N16924, N16901, N16314, N13226, N391);
xor XOR2 (N16925, N16912, N10825);
buf BUF1 (N16926, N16893);
nor NOR4 (N16927, N16923, N2719, N7897, N13878);
and AND2 (N16928, N16925, N11357);
or OR3 (N16929, N16921, N15754, N12439);
and AND4 (N16930, N16926, N10487, N11211, N5228);
buf BUF1 (N16931, N16924);
xor XOR2 (N16932, N16929, N3191);
not NOT1 (N16933, N16930);
nor NOR4 (N16934, N16927, N16444, N15683, N7996);
nor NOR4 (N16935, N16931, N14219, N9826, N4719);
nor NOR2 (N16936, N16932, N15473);
and AND4 (N16937, N16885, N8459, N3313, N68);
and AND3 (N16938, N16909, N5840, N12821);
not NOT1 (N16939, N16935);
nor NOR3 (N16940, N16937, N11608, N2421);
nand NAND2 (N16941, N16934, N12292);
not NOT1 (N16942, N16939);
and AND2 (N16943, N16940, N11722);
not NOT1 (N16944, N16922);
or OR2 (N16945, N16941, N12545);
and AND4 (N16946, N16944, N3317, N14936, N3954);
and AND2 (N16947, N16920, N6803);
and AND2 (N16948, N16936, N16447);
and AND3 (N16949, N16918, N8465, N1594);
nand NAND3 (N16950, N16933, N14624, N16672);
and AND3 (N16951, N16928, N12933, N10018);
xor XOR2 (N16952, N16949, N12451);
buf BUF1 (N16953, N16952);
xor XOR2 (N16954, N16950, N5007);
not NOT1 (N16955, N16948);
xor XOR2 (N16956, N16955, N12705);
or OR4 (N16957, N16956, N10420, N8442, N1976);
xor XOR2 (N16958, N16942, N4675);
nor NOR2 (N16959, N16958, N4039);
xor XOR2 (N16960, N16951, N3135);
or OR2 (N16961, N16960, N12613);
buf BUF1 (N16962, N16943);
not NOT1 (N16963, N16962);
buf BUF1 (N16964, N16961);
or OR4 (N16965, N16964, N11483, N6106, N11379);
not NOT1 (N16966, N16938);
buf BUF1 (N16967, N16966);
and AND4 (N16968, N16953, N13212, N5733, N13974);
not NOT1 (N16969, N16965);
or OR2 (N16970, N16969, N10780);
nand NAND3 (N16971, N16957, N442, N5138);
or OR2 (N16972, N16945, N5391);
nor NOR3 (N16973, N16971, N15227, N11719);
or OR3 (N16974, N16947, N1722, N2341);
and AND2 (N16975, N16963, N7622);
buf BUF1 (N16976, N16974);
not NOT1 (N16977, N16959);
not NOT1 (N16978, N16976);
xor XOR2 (N16979, N16972, N1097);
xor XOR2 (N16980, N16968, N12085);
and AND3 (N16981, N16967, N15288, N8266);
buf BUF1 (N16982, N16975);
or OR4 (N16983, N16977, N7349, N5340, N9498);
not NOT1 (N16984, N16980);
nand NAND2 (N16985, N16973, N3431);
and AND4 (N16986, N16982, N11665, N12714, N14116);
xor XOR2 (N16987, N16970, N10238);
nor NOR3 (N16988, N16986, N2955, N9473);
or OR3 (N16989, N16985, N13063, N12452);
nand NAND3 (N16990, N16981, N13175, N4755);
nand NAND4 (N16991, N16954, N2468, N4440, N306);
nor NOR2 (N16992, N16983, N1503);
buf BUF1 (N16993, N16988);
not NOT1 (N16994, N16990);
or OR4 (N16995, N16946, N10806, N4010, N8412);
nand NAND3 (N16996, N16984, N7574, N7602);
xor XOR2 (N16997, N16989, N169);
and AND3 (N16998, N16991, N16927, N8022);
or OR3 (N16999, N16995, N1555, N3948);
or OR3 (N17000, N16992, N14736, N9628);
xor XOR2 (N17001, N16993, N15836);
buf BUF1 (N17002, N16996);
and AND4 (N17003, N17001, N15819, N12420, N11645);
xor XOR2 (N17004, N17000, N3535);
or OR3 (N17005, N16997, N13454, N2527);
buf BUF1 (N17006, N16978);
or OR3 (N17007, N16994, N14897, N10669);
and AND3 (N17008, N16999, N1063, N15989);
xor XOR2 (N17009, N17002, N6083);
not NOT1 (N17010, N16979);
or OR3 (N17011, N17003, N16405, N14107);
nand NAND3 (N17012, N17010, N4406, N4252);
nand NAND2 (N17013, N17008, N5479);
nor NOR3 (N17014, N17013, N2345, N11728);
nand NAND4 (N17015, N17014, N7481, N6908, N4011);
nand NAND4 (N17016, N16998, N1608, N15297, N6717);
nor NOR3 (N17017, N16987, N8819, N8304);
buf BUF1 (N17018, N17005);
or OR3 (N17019, N17011, N4523, N1607);
buf BUF1 (N17020, N17007);
nor NOR3 (N17021, N17019, N11324, N1767);
nor NOR4 (N17022, N17021, N11429, N15675, N14949);
nand NAND3 (N17023, N17012, N11667, N7565);
nor NOR3 (N17024, N17023, N4918, N3835);
nand NAND2 (N17025, N17006, N15967);
or OR2 (N17026, N17017, N11664);
nand NAND3 (N17027, N17024, N13204, N4700);
xor XOR2 (N17028, N17026, N7229);
nor NOR2 (N17029, N17022, N12386);
or OR3 (N17030, N17009, N9515, N5313);
nand NAND2 (N17031, N17015, N7736);
or OR2 (N17032, N17004, N498);
or OR3 (N17033, N17029, N4629, N8497);
or OR2 (N17034, N17028, N15697);
and AND2 (N17035, N17020, N793);
nor NOR2 (N17036, N17025, N5941);
xor XOR2 (N17037, N17033, N11010);
nor NOR3 (N17038, N17037, N14271, N2812);
buf BUF1 (N17039, N17027);
nand NAND4 (N17040, N17039, N12860, N5862, N3376);
nor NOR2 (N17041, N17031, N10209);
nand NAND4 (N17042, N17035, N7668, N10407, N6676);
nand NAND2 (N17043, N17036, N5946);
xor XOR2 (N17044, N17018, N8116);
nand NAND4 (N17045, N17044, N13134, N3882, N3525);
buf BUF1 (N17046, N17045);
xor XOR2 (N17047, N17041, N5322);
buf BUF1 (N17048, N17032);
nor NOR4 (N17049, N17030, N10917, N1550, N3021);
xor XOR2 (N17050, N17038, N12617);
buf BUF1 (N17051, N17048);
nand NAND2 (N17052, N17046, N9160);
nand NAND2 (N17053, N17042, N5136);
xor XOR2 (N17054, N17049, N7987);
xor XOR2 (N17055, N17053, N12308);
not NOT1 (N17056, N17054);
nand NAND4 (N17057, N17040, N16377, N12499, N16549);
not NOT1 (N17058, N17050);
or OR4 (N17059, N17016, N3867, N14335, N16324);
not NOT1 (N17060, N17055);
and AND4 (N17061, N17034, N5518, N15934, N14562);
buf BUF1 (N17062, N17043);
nor NOR3 (N17063, N17062, N477, N6073);
not NOT1 (N17064, N17059);
not NOT1 (N17065, N17060);
and AND4 (N17066, N17052, N9913, N4687, N5302);
and AND3 (N17067, N17051, N189, N15528);
nor NOR3 (N17068, N17064, N5395, N10244);
or OR3 (N17069, N17061, N5207, N11574);
not NOT1 (N17070, N17058);
or OR4 (N17071, N17057, N14953, N4977, N6081);
xor XOR2 (N17072, N17070, N16291);
nand NAND3 (N17073, N17068, N9388, N5941);
or OR3 (N17074, N17066, N4570, N15093);
or OR3 (N17075, N17063, N11430, N15885);
nor NOR2 (N17076, N17072, N6401);
and AND4 (N17077, N17074, N1990, N3799, N11368);
or OR3 (N17078, N17069, N14831, N11990);
and AND4 (N17079, N17075, N1546, N15803, N8862);
buf BUF1 (N17080, N17079);
xor XOR2 (N17081, N17078, N14588);
or OR4 (N17082, N17065, N5290, N12206, N5520);
nor NOR4 (N17083, N17080, N5546, N731, N15202);
buf BUF1 (N17084, N17073);
nor NOR3 (N17085, N17081, N11198, N5786);
or OR3 (N17086, N17084, N3380, N4014);
nand NAND4 (N17087, N17076, N4026, N12763, N8618);
or OR2 (N17088, N17067, N12847);
not NOT1 (N17089, N17088);
nand NAND2 (N17090, N17085, N4112);
or OR2 (N17091, N17090, N2718);
nand NAND2 (N17092, N17082, N15564);
nor NOR4 (N17093, N17092, N12395, N15612, N5411);
or OR2 (N17094, N17083, N7899);
xor XOR2 (N17095, N17077, N1641);
xor XOR2 (N17096, N17089, N12332);
nor NOR2 (N17097, N17047, N7304);
or OR4 (N17098, N17086, N13923, N12354, N4282);
nand NAND2 (N17099, N17095, N4192);
not NOT1 (N17100, N17099);
nand NAND4 (N17101, N17056, N11804, N9584, N12263);
nand NAND2 (N17102, N17101, N3241);
nand NAND3 (N17103, N17087, N3922, N918);
or OR2 (N17104, N17094, N3736);
nand NAND3 (N17105, N17103, N3894, N15631);
nor NOR2 (N17106, N17104, N11122);
or OR4 (N17107, N17091, N8141, N1091, N4517);
or OR4 (N17108, N17071, N11333, N1858, N9191);
and AND4 (N17109, N17107, N13188, N15976, N9439);
not NOT1 (N17110, N17100);
nor NOR3 (N17111, N17105, N8105, N11804);
and AND4 (N17112, N17098, N4987, N14604, N6527);
and AND2 (N17113, N17111, N9216);
xor XOR2 (N17114, N17096, N13609);
nor NOR3 (N17115, N17108, N2059, N4051);
buf BUF1 (N17116, N17110);
or OR2 (N17117, N17114, N17018);
buf BUF1 (N17118, N17102);
buf BUF1 (N17119, N17115);
nand NAND3 (N17120, N17112, N9417, N4425);
xor XOR2 (N17121, N17097, N13041);
nand NAND4 (N17122, N17106, N10434, N11318, N10897);
xor XOR2 (N17123, N17120, N10129);
nor NOR2 (N17124, N17121, N12103);
and AND4 (N17125, N17122, N7900, N8288, N2871);
xor XOR2 (N17126, N17109, N861);
nand NAND4 (N17127, N17113, N8943, N12065, N9220);
and AND3 (N17128, N17116, N14657, N14118);
or OR2 (N17129, N17126, N11947);
not NOT1 (N17130, N17127);
not NOT1 (N17131, N17130);
not NOT1 (N17132, N17118);
not NOT1 (N17133, N17124);
xor XOR2 (N17134, N17119, N13304);
not NOT1 (N17135, N17132);
xor XOR2 (N17136, N17129, N5291);
nor NOR2 (N17137, N17117, N509);
buf BUF1 (N17138, N17093);
and AND2 (N17139, N17128, N7043);
nor NOR2 (N17140, N17131, N16199);
or OR3 (N17141, N17135, N12758, N11405);
nor NOR4 (N17142, N17139, N10140, N9236, N7105);
not NOT1 (N17143, N17123);
nand NAND2 (N17144, N17143, N1589);
nor NOR2 (N17145, N17138, N4863);
xor XOR2 (N17146, N17125, N9101);
xor XOR2 (N17147, N17141, N70);
or OR2 (N17148, N17136, N8601);
nand NAND3 (N17149, N17148, N10262, N4396);
or OR2 (N17150, N17144, N15509);
nand NAND3 (N17151, N17145, N15921, N209);
buf BUF1 (N17152, N17133);
xor XOR2 (N17153, N17151, N13637);
nand NAND4 (N17154, N17142, N4707, N11961, N6271);
or OR2 (N17155, N17149, N8762);
or OR3 (N17156, N17147, N14910, N10596);
or OR4 (N17157, N17156, N16988, N3255, N2257);
and AND2 (N17158, N17157, N9578);
or OR3 (N17159, N17158, N8329, N232);
buf BUF1 (N17160, N17137);
not NOT1 (N17161, N17152);
not NOT1 (N17162, N17155);
buf BUF1 (N17163, N17153);
xor XOR2 (N17164, N17161, N13341);
or OR2 (N17165, N17160, N3198);
and AND4 (N17166, N17154, N4537, N12277, N4411);
nand NAND3 (N17167, N17140, N10288, N2609);
nor NOR3 (N17168, N17162, N11317, N17150);
nor NOR2 (N17169, N11674, N10581);
and AND3 (N17170, N17159, N1948, N4237);
not NOT1 (N17171, N17170);
nand NAND2 (N17172, N17166, N14443);
and AND2 (N17173, N17172, N8430);
not NOT1 (N17174, N17171);
nand NAND2 (N17175, N17169, N4826);
and AND2 (N17176, N17174, N14169);
or OR2 (N17177, N17164, N15945);
or OR3 (N17178, N17134, N5908, N8573);
and AND3 (N17179, N17165, N8080, N2969);
buf BUF1 (N17180, N17163);
not NOT1 (N17181, N17179);
not NOT1 (N17182, N17181);
nand NAND2 (N17183, N17173, N9131);
xor XOR2 (N17184, N17176, N1290);
nor NOR4 (N17185, N17183, N12840, N7289, N10276);
xor XOR2 (N17186, N17168, N8396);
and AND4 (N17187, N17167, N6094, N6173, N8335);
or OR3 (N17188, N17184, N15431, N16710);
or OR2 (N17189, N17175, N11878);
and AND3 (N17190, N17180, N14613, N2670);
nor NOR3 (N17191, N17177, N13620, N5910);
or OR2 (N17192, N17146, N11131);
nand NAND2 (N17193, N17178, N6270);
buf BUF1 (N17194, N17186);
nand NAND3 (N17195, N17191, N15764, N14478);
or OR2 (N17196, N17192, N12430);
buf BUF1 (N17197, N17195);
xor XOR2 (N17198, N17188, N6339);
nor NOR4 (N17199, N17197, N14958, N8504, N13673);
nand NAND3 (N17200, N17194, N129, N7826);
buf BUF1 (N17201, N17196);
xor XOR2 (N17202, N17187, N2844);
buf BUF1 (N17203, N17200);
nor NOR4 (N17204, N17201, N2288, N242, N5913);
and AND3 (N17205, N17203, N9661, N8533);
nor NOR2 (N17206, N17190, N11417);
nor NOR4 (N17207, N17204, N13096, N4089, N15031);
or OR3 (N17208, N17199, N704, N14008);
not NOT1 (N17209, N17207);
nand NAND2 (N17210, N17182, N5551);
or OR4 (N17211, N17206, N11867, N11805, N5825);
or OR3 (N17212, N17211, N8112, N6023);
or OR3 (N17213, N17205, N11891, N9919);
or OR4 (N17214, N17185, N11178, N9659, N6384);
xor XOR2 (N17215, N17212, N1009);
xor XOR2 (N17216, N17193, N15778);
nor NOR2 (N17217, N17202, N14738);
nand NAND3 (N17218, N17198, N4552, N10569);
nor NOR2 (N17219, N17209, N7479);
or OR3 (N17220, N17216, N4730, N7715);
or OR2 (N17221, N17218, N16304);
not NOT1 (N17222, N17213);
not NOT1 (N17223, N17214);
buf BUF1 (N17224, N17221);
buf BUF1 (N17225, N17208);
nor NOR4 (N17226, N17222, N3763, N6394, N3401);
buf BUF1 (N17227, N17215);
xor XOR2 (N17228, N17217, N10679);
nor NOR3 (N17229, N17219, N4164, N10845);
buf BUF1 (N17230, N17189);
buf BUF1 (N17231, N17230);
nand NAND4 (N17232, N17228, N5274, N578, N16277);
nor NOR2 (N17233, N17232, N8736);
or OR3 (N17234, N17229, N7357, N12895);
nand NAND2 (N17235, N17220, N5033);
buf BUF1 (N17236, N17227);
and AND3 (N17237, N17224, N5997, N14266);
not NOT1 (N17238, N17225);
nand NAND2 (N17239, N17238, N13703);
and AND3 (N17240, N17226, N15272, N9417);
buf BUF1 (N17241, N17237);
buf BUF1 (N17242, N17231);
xor XOR2 (N17243, N17236, N8275);
buf BUF1 (N17244, N17233);
nand NAND2 (N17245, N17241, N435);
nor NOR2 (N17246, N17245, N13268);
nand NAND3 (N17247, N17234, N7810, N13441);
not NOT1 (N17248, N17244);
and AND4 (N17249, N17247, N6848, N16006, N7321);
not NOT1 (N17250, N17249);
nor NOR2 (N17251, N17239, N14135);
not NOT1 (N17252, N17243);
xor XOR2 (N17253, N17240, N15436);
not NOT1 (N17254, N17223);
xor XOR2 (N17255, N17210, N597);
nand NAND3 (N17256, N17252, N7007, N3650);
and AND4 (N17257, N17251, N13767, N12401, N17087);
nor NOR2 (N17258, N17253, N5207);
xor XOR2 (N17259, N17250, N5352);
not NOT1 (N17260, N17259);
nor NOR3 (N17261, N17235, N11440, N13415);
nor NOR3 (N17262, N17242, N5547, N686);
or OR4 (N17263, N17257, N13737, N5378, N13541);
nand NAND2 (N17264, N17246, N5131);
not NOT1 (N17265, N17263);
nor NOR2 (N17266, N17261, N2295);
nand NAND3 (N17267, N17248, N6837, N10852);
nor NOR2 (N17268, N17256, N16681);
not NOT1 (N17269, N17267);
and AND3 (N17270, N17269, N14715, N15656);
xor XOR2 (N17271, N17258, N6407);
xor XOR2 (N17272, N17254, N6588);
xor XOR2 (N17273, N17260, N2290);
or OR4 (N17274, N17273, N4973, N16963, N1628);
nor NOR3 (N17275, N17270, N5213, N16977);
xor XOR2 (N17276, N17264, N6671);
nor NOR2 (N17277, N17266, N1721);
not NOT1 (N17278, N17255);
buf BUF1 (N17279, N17262);
or OR4 (N17280, N17277, N16796, N12731, N11856);
or OR3 (N17281, N17271, N1706, N13031);
or OR3 (N17282, N17278, N13979, N15823);
or OR2 (N17283, N17274, N1223);
and AND4 (N17284, N17282, N11816, N16880, N2505);
buf BUF1 (N17285, N17276);
and AND4 (N17286, N17279, N7210, N4044, N6650);
buf BUF1 (N17287, N17275);
and AND2 (N17288, N17287, N4878);
nor NOR4 (N17289, N17272, N3645, N4159, N14962);
not NOT1 (N17290, N17289);
and AND4 (N17291, N17280, N14269, N14565, N116);
or OR2 (N17292, N17290, N14509);
xor XOR2 (N17293, N17286, N4642);
xor XOR2 (N17294, N17283, N10344);
xor XOR2 (N17295, N17294, N14552);
nand NAND2 (N17296, N17285, N13493);
and AND4 (N17297, N17281, N15224, N12402, N2590);
not NOT1 (N17298, N17284);
xor XOR2 (N17299, N17268, N7736);
and AND2 (N17300, N17293, N10389);
buf BUF1 (N17301, N17296);
or OR3 (N17302, N17300, N5599, N2709);
not NOT1 (N17303, N17302);
nand NAND2 (N17304, N17265, N3502);
buf BUF1 (N17305, N17295);
buf BUF1 (N17306, N17301);
or OR3 (N17307, N17288, N13174, N11235);
nand NAND2 (N17308, N17303, N8040);
or OR4 (N17309, N17299, N16697, N9474, N12831);
and AND3 (N17310, N17298, N6304, N11081);
or OR3 (N17311, N17306, N11774, N15966);
xor XOR2 (N17312, N17307, N6219);
and AND3 (N17313, N17309, N12308, N11702);
buf BUF1 (N17314, N17312);
not NOT1 (N17315, N17313);
not NOT1 (N17316, N17314);
and AND2 (N17317, N17310, N7520);
nand NAND2 (N17318, N17315, N4215);
or OR3 (N17319, N17318, N3459, N3799);
nand NAND3 (N17320, N17317, N962, N15307);
or OR4 (N17321, N17311, N819, N9354, N8757);
or OR2 (N17322, N17320, N11154);
and AND2 (N17323, N17308, N16292);
not NOT1 (N17324, N17305);
or OR4 (N17325, N17324, N11569, N17119, N3519);
xor XOR2 (N17326, N17291, N599);
xor XOR2 (N17327, N17316, N9011);
buf BUF1 (N17328, N17321);
xor XOR2 (N17329, N17327, N3631);
buf BUF1 (N17330, N17292);
and AND4 (N17331, N17304, N11527, N6370, N5767);
or OR4 (N17332, N17325, N7406, N15728, N9884);
buf BUF1 (N17333, N17297);
or OR2 (N17334, N17326, N2334);
nand NAND4 (N17335, N17331, N2614, N263, N3762);
nor NOR3 (N17336, N17335, N13279, N11352);
nor NOR4 (N17337, N17334, N3718, N9678, N9165);
or OR2 (N17338, N17333, N15496);
nor NOR3 (N17339, N17336, N11814, N8787);
xor XOR2 (N17340, N17329, N10598);
nor NOR3 (N17341, N17322, N12857, N425);
and AND4 (N17342, N17338, N14196, N2829, N2373);
nor NOR2 (N17343, N17319, N5168);
buf BUF1 (N17344, N17323);
not NOT1 (N17345, N17342);
not NOT1 (N17346, N17328);
xor XOR2 (N17347, N17345, N7794);
buf BUF1 (N17348, N17347);
buf BUF1 (N17349, N17337);
or OR4 (N17350, N17349, N14445, N11398, N13594);
nand NAND2 (N17351, N17341, N2626);
nand NAND2 (N17352, N17339, N757);
nand NAND2 (N17353, N17346, N275);
nand NAND2 (N17354, N17344, N12270);
and AND2 (N17355, N17348, N4462);
or OR4 (N17356, N17354, N5021, N14541, N7183);
xor XOR2 (N17357, N17352, N4391);
and AND3 (N17358, N17332, N8359, N7879);
nand NAND3 (N17359, N17358, N12999, N11698);
buf BUF1 (N17360, N17357);
xor XOR2 (N17361, N17350, N16655);
not NOT1 (N17362, N17356);
nor NOR2 (N17363, N17343, N10772);
nand NAND2 (N17364, N17359, N1246);
nand NAND3 (N17365, N17360, N16602, N6438);
buf BUF1 (N17366, N17363);
or OR3 (N17367, N17365, N2521, N12295);
and AND3 (N17368, N17361, N7461, N16245);
nand NAND2 (N17369, N17367, N9807);
or OR4 (N17370, N17340, N14420, N8468, N2454);
and AND4 (N17371, N17364, N6733, N2234, N7476);
nand NAND3 (N17372, N17330, N15932, N9399);
xor XOR2 (N17373, N17368, N8);
xor XOR2 (N17374, N17362, N10063);
or OR4 (N17375, N17369, N819, N3465, N2782);
buf BUF1 (N17376, N17366);
not NOT1 (N17377, N17373);
nand NAND2 (N17378, N17372, N6617);
not NOT1 (N17379, N17374);
and AND4 (N17380, N17378, N6980, N11428, N2681);
nand NAND2 (N17381, N17379, N5188);
xor XOR2 (N17382, N17376, N2141);
nand NAND4 (N17383, N17381, N1416, N8445, N16979);
nor NOR3 (N17384, N17355, N4090, N8801);
nand NAND2 (N17385, N17382, N15667);
and AND4 (N17386, N17353, N7410, N5185, N9723);
nor NOR4 (N17387, N17375, N12874, N6792, N4686);
and AND3 (N17388, N17370, N5866, N141);
nor NOR4 (N17389, N17377, N13499, N12512, N4356);
xor XOR2 (N17390, N17389, N8658);
and AND2 (N17391, N17383, N5963);
and AND3 (N17392, N17380, N7062, N16965);
buf BUF1 (N17393, N17392);
and AND2 (N17394, N17391, N17087);
and AND2 (N17395, N17386, N12357);
and AND2 (N17396, N17385, N10663);
and AND2 (N17397, N17387, N16681);
or OR4 (N17398, N17390, N6311, N6726, N17340);
or OR2 (N17399, N17395, N4037);
nand NAND4 (N17400, N17396, N1559, N1477, N1014);
buf BUF1 (N17401, N17384);
buf BUF1 (N17402, N17393);
nand NAND3 (N17403, N17399, N17296, N7871);
or OR4 (N17404, N17398, N4950, N16917, N8126);
not NOT1 (N17405, N17403);
or OR2 (N17406, N17404, N4004);
nor NOR4 (N17407, N17402, N1168, N10879, N7408);
nor NOR3 (N17408, N17397, N16761, N4213);
buf BUF1 (N17409, N17388);
xor XOR2 (N17410, N17406, N8684);
nand NAND2 (N17411, N17410, N10884);
and AND4 (N17412, N17407, N4521, N12233, N13419);
nor NOR2 (N17413, N17405, N13385);
not NOT1 (N17414, N17351);
nand NAND2 (N17415, N17371, N8189);
or OR3 (N17416, N17412, N8337, N17181);
not NOT1 (N17417, N17411);
xor XOR2 (N17418, N17416, N17152);
buf BUF1 (N17419, N17413);
nand NAND2 (N17420, N17400, N7084);
and AND3 (N17421, N17414, N14740, N13579);
buf BUF1 (N17422, N17394);
not NOT1 (N17423, N17409);
nor NOR4 (N17424, N17421, N12894, N2585, N13284);
not NOT1 (N17425, N17424);
nor NOR4 (N17426, N17419, N9378, N7597, N11119);
not NOT1 (N17427, N17418);
buf BUF1 (N17428, N17427);
xor XOR2 (N17429, N17426, N13525);
buf BUF1 (N17430, N17408);
or OR3 (N17431, N17417, N3611, N5661);
nand NAND3 (N17432, N17425, N13692, N12594);
buf BUF1 (N17433, N17431);
nand NAND4 (N17434, N17423, N13143, N9658, N17050);
nand NAND4 (N17435, N17430, N2691, N12512, N13184);
nor NOR4 (N17436, N17435, N3555, N17398, N420);
nand NAND4 (N17437, N17436, N13201, N4872, N16314);
nor NOR3 (N17438, N17420, N8385, N16300);
xor XOR2 (N17439, N17438, N1860);
not NOT1 (N17440, N17429);
or OR2 (N17441, N17428, N694);
not NOT1 (N17442, N17433);
not NOT1 (N17443, N17434);
or OR4 (N17444, N17401, N17112, N6082, N888);
or OR2 (N17445, N17415, N12742);
and AND4 (N17446, N17439, N9831, N15227, N8427);
nor NOR3 (N17447, N17432, N6320, N8729);
nand NAND4 (N17448, N17447, N17105, N4778, N5127);
and AND3 (N17449, N17445, N1654, N2381);
or OR2 (N17450, N17444, N3416);
and AND4 (N17451, N17422, N7928, N7111, N3138);
or OR2 (N17452, N17449, N2488);
nor NOR2 (N17453, N17446, N1320);
buf BUF1 (N17454, N17442);
buf BUF1 (N17455, N17450);
xor XOR2 (N17456, N17455, N15069);
or OR2 (N17457, N17448, N4872);
or OR2 (N17458, N17454, N15064);
or OR3 (N17459, N17452, N7855, N256);
or OR3 (N17460, N17457, N4855, N7854);
and AND4 (N17461, N17437, N8210, N13220, N8321);
buf BUF1 (N17462, N17459);
or OR3 (N17463, N17458, N14555, N6267);
nand NAND3 (N17464, N17441, N14936, N7289);
xor XOR2 (N17465, N17443, N7142);
nand NAND3 (N17466, N17465, N15848, N3938);
xor XOR2 (N17467, N17453, N8900);
and AND2 (N17468, N17456, N571);
nor NOR2 (N17469, N17466, N138);
and AND4 (N17470, N17464, N4884, N3515, N5416);
xor XOR2 (N17471, N17469, N10752);
xor XOR2 (N17472, N17467, N8815);
and AND2 (N17473, N17468, N3584);
not NOT1 (N17474, N17472);
and AND4 (N17475, N17462, N8227, N10336, N14132);
not NOT1 (N17476, N17451);
buf BUF1 (N17477, N17475);
xor XOR2 (N17478, N17463, N4560);
buf BUF1 (N17479, N17476);
buf BUF1 (N17480, N17473);
not NOT1 (N17481, N17474);
buf BUF1 (N17482, N17478);
nor NOR4 (N17483, N17471, N10039, N13372, N2993);
nor NOR3 (N17484, N17461, N6952, N2269);
nor NOR3 (N17485, N17482, N6659, N10129);
and AND4 (N17486, N17485, N6654, N4756, N557);
buf BUF1 (N17487, N17484);
or OR4 (N17488, N17479, N16681, N9265, N956);
or OR2 (N17489, N17470, N6212);
buf BUF1 (N17490, N17477);
or OR3 (N17491, N17490, N14183, N913);
nor NOR2 (N17492, N17486, N468);
buf BUF1 (N17493, N17487);
nor NOR3 (N17494, N17480, N11307, N16632);
and AND4 (N17495, N17488, N13306, N9963, N14673);
nand NAND3 (N17496, N17493, N4606, N5311);
nor NOR3 (N17497, N17494, N5441, N15080);
buf BUF1 (N17498, N17495);
buf BUF1 (N17499, N17498);
xor XOR2 (N17500, N17483, N15458);
xor XOR2 (N17501, N17491, N13165);
xor XOR2 (N17502, N17492, N15986);
xor XOR2 (N17503, N17501, N5451);
or OR2 (N17504, N17481, N16106);
xor XOR2 (N17505, N17499, N9577);
not NOT1 (N17506, N17460);
not NOT1 (N17507, N17503);
xor XOR2 (N17508, N17507, N2066);
nor NOR2 (N17509, N17489, N11802);
nor NOR4 (N17510, N17440, N368, N12512, N13562);
and AND4 (N17511, N17505, N12916, N2576, N3591);
buf BUF1 (N17512, N17504);
and AND4 (N17513, N17496, N12807, N13045, N1703);
xor XOR2 (N17514, N17506, N8655);
not NOT1 (N17515, N17509);
nand NAND3 (N17516, N17511, N13015, N2190);
nand NAND3 (N17517, N17513, N4524, N9120);
buf BUF1 (N17518, N17515);
or OR2 (N17519, N17502, N7506);
not NOT1 (N17520, N17516);
xor XOR2 (N17521, N17497, N2252);
buf BUF1 (N17522, N17512);
and AND3 (N17523, N17522, N5114, N15050);
or OR4 (N17524, N17500, N15934, N12502, N290);
xor XOR2 (N17525, N17510, N12558);
nor NOR4 (N17526, N17521, N15637, N10906, N3214);
or OR2 (N17527, N17508, N15069);
xor XOR2 (N17528, N17514, N7785);
nand NAND4 (N17529, N17519, N12114, N11928, N1262);
xor XOR2 (N17530, N17518, N6585);
and AND4 (N17531, N17523, N2815, N4904, N2490);
xor XOR2 (N17532, N17520, N6719);
xor XOR2 (N17533, N17531, N7057);
nor NOR2 (N17534, N17532, N13821);
or OR3 (N17535, N17530, N10436, N9173);
xor XOR2 (N17536, N17529, N10857);
or OR2 (N17537, N17535, N1853);
and AND4 (N17538, N17517, N8117, N2119, N2250);
not NOT1 (N17539, N17536);
nand NAND2 (N17540, N17533, N5650);
not NOT1 (N17541, N17525);
or OR2 (N17542, N17527, N1834);
buf BUF1 (N17543, N17528);
xor XOR2 (N17544, N17543, N11095);
buf BUF1 (N17545, N17544);
or OR3 (N17546, N17540, N5121, N16446);
xor XOR2 (N17547, N17524, N16777);
or OR2 (N17548, N17534, N13817);
not NOT1 (N17549, N17539);
xor XOR2 (N17550, N17545, N11533);
xor XOR2 (N17551, N17547, N1235);
nand NAND4 (N17552, N17546, N11380, N14167, N9600);
xor XOR2 (N17553, N17552, N11615);
or OR2 (N17554, N17553, N9412);
or OR2 (N17555, N17550, N10898);
not NOT1 (N17556, N17542);
xor XOR2 (N17557, N17541, N91);
nand NAND2 (N17558, N17548, N15207);
not NOT1 (N17559, N17551);
nor NOR3 (N17560, N17555, N4428, N7338);
or OR4 (N17561, N17558, N11922, N17337, N15908);
or OR2 (N17562, N17559, N9714);
or OR2 (N17563, N17537, N11396);
nand NAND2 (N17564, N17562, N14097);
nor NOR2 (N17565, N17560, N5696);
not NOT1 (N17566, N17557);
or OR3 (N17567, N17566, N14824, N5071);
and AND4 (N17568, N17554, N15543, N1592, N10206);
buf BUF1 (N17569, N17561);
nand NAND4 (N17570, N17526, N14757, N10199, N1510);
nand NAND3 (N17571, N17569, N6715, N13869);
nand NAND2 (N17572, N17567, N14955);
nor NOR2 (N17573, N17549, N5801);
or OR3 (N17574, N17556, N16690, N7949);
or OR4 (N17575, N17565, N7869, N10075, N8515);
xor XOR2 (N17576, N17572, N7724);
or OR2 (N17577, N17575, N3681);
nand NAND3 (N17578, N17538, N10884, N2726);
and AND3 (N17579, N17577, N8863, N14574);
nor NOR4 (N17580, N17573, N8372, N13936, N13366);
nor NOR4 (N17581, N17579, N9655, N6464, N15279);
nand NAND3 (N17582, N17581, N10497, N14790);
buf BUF1 (N17583, N17568);
buf BUF1 (N17584, N17582);
not NOT1 (N17585, N17570);
nor NOR3 (N17586, N17574, N8484, N16616);
xor XOR2 (N17587, N17564, N11320);
and AND4 (N17588, N17578, N17376, N16597, N12502);
buf BUF1 (N17589, N17585);
or OR2 (N17590, N17587, N1799);
or OR2 (N17591, N17580, N8742);
xor XOR2 (N17592, N17591, N2380);
xor XOR2 (N17593, N17590, N17343);
nand NAND4 (N17594, N17586, N10279, N16517, N1132);
xor XOR2 (N17595, N17594, N8991);
or OR3 (N17596, N17563, N4822, N11224);
not NOT1 (N17597, N17592);
buf BUF1 (N17598, N17593);
not NOT1 (N17599, N17597);
buf BUF1 (N17600, N17596);
nand NAND4 (N17601, N17595, N10384, N7673, N5045);
or OR2 (N17602, N17583, N10485);
nand NAND3 (N17603, N17589, N17274, N7267);
or OR2 (N17604, N17602, N771);
xor XOR2 (N17605, N17599, N1824);
or OR2 (N17606, N17571, N15249);
xor XOR2 (N17607, N17576, N15960);
and AND4 (N17608, N17607, N4811, N13919, N17532);
nor NOR4 (N17609, N17604, N13096, N12428, N14301);
xor XOR2 (N17610, N17603, N14222);
not NOT1 (N17611, N17600);
nor NOR4 (N17612, N17598, N5751, N1949, N9657);
xor XOR2 (N17613, N17584, N59);
and AND2 (N17614, N17588, N9944);
nor NOR3 (N17615, N17605, N10218, N2422);
or OR2 (N17616, N17606, N10335);
buf BUF1 (N17617, N17613);
nand NAND2 (N17618, N17617, N1081);
and AND2 (N17619, N17615, N8462);
buf BUF1 (N17620, N17616);
xor XOR2 (N17621, N17601, N264);
xor XOR2 (N17622, N17609, N1878);
and AND3 (N17623, N17620, N370, N5786);
nand NAND3 (N17624, N17618, N8701, N9607);
nor NOR4 (N17625, N17622, N2213, N2010, N17220);
nor NOR3 (N17626, N17611, N9832, N7572);
and AND3 (N17627, N17608, N75, N16467);
nand NAND3 (N17628, N17610, N6489, N449);
buf BUF1 (N17629, N17614);
not NOT1 (N17630, N17623);
nor NOR3 (N17631, N17626, N6052, N1587);
buf BUF1 (N17632, N17631);
nor NOR4 (N17633, N17630, N632, N4663, N6772);
not NOT1 (N17634, N17633);
nor NOR3 (N17635, N17628, N2285, N16382);
xor XOR2 (N17636, N17627, N8262);
xor XOR2 (N17637, N17635, N5415);
and AND2 (N17638, N17621, N16609);
not NOT1 (N17639, N17638);
not NOT1 (N17640, N17637);
not NOT1 (N17641, N17629);
nand NAND3 (N17642, N17624, N13434, N78);
and AND3 (N17643, N17639, N6779, N350);
or OR3 (N17644, N17625, N9447, N1305);
xor XOR2 (N17645, N17636, N10832);
not NOT1 (N17646, N17640);
nor NOR3 (N17647, N17642, N5491, N6085);
and AND2 (N17648, N17612, N8586);
nand NAND2 (N17649, N17619, N2466);
not NOT1 (N17650, N17643);
nand NAND3 (N17651, N17644, N5338, N15759);
or OR2 (N17652, N17634, N7941);
xor XOR2 (N17653, N17646, N2394);
or OR2 (N17654, N17641, N13287);
nor NOR3 (N17655, N17649, N4444, N6115);
nor NOR2 (N17656, N17632, N14682);
or OR2 (N17657, N17655, N1414);
buf BUF1 (N17658, N17651);
nor NOR4 (N17659, N17653, N1597, N6562, N8326);
nor NOR2 (N17660, N17648, N14235);
buf BUF1 (N17661, N17652);
not NOT1 (N17662, N17656);
or OR3 (N17663, N17658, N12753, N7927);
or OR3 (N17664, N17663, N9048, N8302);
nor NOR2 (N17665, N17657, N10524);
buf BUF1 (N17666, N17659);
buf BUF1 (N17667, N17650);
or OR4 (N17668, N17654, N15716, N8791, N4599);
xor XOR2 (N17669, N17661, N11711);
nand NAND2 (N17670, N17669, N16471);
or OR2 (N17671, N17645, N6683);
or OR3 (N17672, N17668, N4780, N13822);
xor XOR2 (N17673, N17660, N13968);
buf BUF1 (N17674, N17662);
or OR4 (N17675, N17664, N16285, N16664, N3544);
xor XOR2 (N17676, N17675, N15788);
nor NOR4 (N17677, N17665, N431, N4429, N17182);
nand NAND2 (N17678, N17666, N4808);
and AND3 (N17679, N17672, N6033, N1334);
nor NOR2 (N17680, N17674, N16155);
xor XOR2 (N17681, N17671, N6756);
nor NOR3 (N17682, N17673, N3999, N8745);
and AND2 (N17683, N17680, N15965);
nor NOR2 (N17684, N17678, N16229);
buf BUF1 (N17685, N17684);
xor XOR2 (N17686, N17679, N9836);
nand NAND2 (N17687, N17667, N11174);
or OR4 (N17688, N17676, N11196, N11464, N12741);
buf BUF1 (N17689, N17686);
buf BUF1 (N17690, N17647);
xor XOR2 (N17691, N17687, N17481);
and AND2 (N17692, N17677, N11713);
and AND2 (N17693, N17691, N2502);
buf BUF1 (N17694, N17682);
xor XOR2 (N17695, N17694, N634);
xor XOR2 (N17696, N17690, N5316);
or OR4 (N17697, N17689, N10538, N6669, N16140);
buf BUF1 (N17698, N17696);
xor XOR2 (N17699, N17688, N1188);
or OR4 (N17700, N17697, N6884, N17208, N8734);
buf BUF1 (N17701, N17692);
or OR2 (N17702, N17701, N3058);
or OR2 (N17703, N17683, N14332);
not NOT1 (N17704, N17693);
xor XOR2 (N17705, N17699, N15768);
xor XOR2 (N17706, N17704, N15355);
and AND3 (N17707, N17700, N13533, N13493);
nor NOR3 (N17708, N17702, N3389, N6012);
xor XOR2 (N17709, N17670, N3740);
buf BUF1 (N17710, N17681);
buf BUF1 (N17711, N17705);
or OR3 (N17712, N17711, N3725, N2210);
not NOT1 (N17713, N17708);
nand NAND2 (N17714, N17710, N3047);
xor XOR2 (N17715, N17714, N11916);
nor NOR2 (N17716, N17713, N12761);
xor XOR2 (N17717, N17716, N6068);
nand NAND2 (N17718, N17712, N11720);
nand NAND2 (N17719, N17709, N15279);
or OR4 (N17720, N17707, N2252, N8978, N17420);
or OR4 (N17721, N17717, N8554, N3535, N13024);
and AND4 (N17722, N17685, N15925, N9523, N3816);
nand NAND3 (N17723, N17698, N14473, N16945);
not NOT1 (N17724, N17722);
buf BUF1 (N17725, N17695);
buf BUF1 (N17726, N17719);
nor NOR2 (N17727, N17718, N10463);
nor NOR4 (N17728, N17724, N14456, N1600, N15971);
or OR2 (N17729, N17715, N2490);
nor NOR4 (N17730, N17729, N16916, N66, N5334);
or OR4 (N17731, N17728, N11330, N2320, N5368);
or OR3 (N17732, N17721, N9169, N15210);
nand NAND3 (N17733, N17720, N4698, N6438);
xor XOR2 (N17734, N17733, N3157);
xor XOR2 (N17735, N17734, N12164);
and AND4 (N17736, N17723, N965, N16419, N9500);
buf BUF1 (N17737, N17703);
xor XOR2 (N17738, N17730, N7341);
xor XOR2 (N17739, N17737, N12028);
nand NAND4 (N17740, N17706, N16364, N5553, N8277);
nor NOR4 (N17741, N17726, N7784, N5664, N1832);
not NOT1 (N17742, N17741);
or OR2 (N17743, N17732, N11739);
not NOT1 (N17744, N17731);
nand NAND4 (N17745, N17742, N10538, N1621, N2968);
xor XOR2 (N17746, N17738, N8330);
and AND3 (N17747, N17745, N13512, N3172);
not NOT1 (N17748, N17736);
nand NAND4 (N17749, N17740, N10102, N8477, N11106);
nand NAND2 (N17750, N17743, N11387);
and AND3 (N17751, N17750, N16982, N2240);
and AND4 (N17752, N17744, N10852, N6803, N255);
or OR4 (N17753, N17748, N9985, N13199, N11902);
nand NAND3 (N17754, N17727, N6717, N286);
buf BUF1 (N17755, N17751);
and AND2 (N17756, N17735, N8136);
nand NAND4 (N17757, N17752, N15768, N8526, N4055);
not NOT1 (N17758, N17755);
not NOT1 (N17759, N17746);
nor NOR3 (N17760, N17749, N258, N4411);
and AND3 (N17761, N17753, N6929, N812);
or OR3 (N17762, N17725, N15922, N3300);
not NOT1 (N17763, N17757);
nor NOR4 (N17764, N17739, N5410, N16321, N1739);
or OR4 (N17765, N17761, N13251, N10409, N1655);
nand NAND3 (N17766, N17758, N7224, N2037);
xor XOR2 (N17767, N17754, N7196);
not NOT1 (N17768, N17767);
not NOT1 (N17769, N17759);
or OR2 (N17770, N17756, N3943);
or OR4 (N17771, N17765, N14963, N9699, N11441);
nor NOR4 (N17772, N17747, N736, N5062, N17361);
not NOT1 (N17773, N17771);
buf BUF1 (N17774, N17763);
and AND3 (N17775, N17766, N12677, N16230);
not NOT1 (N17776, N17762);
not NOT1 (N17777, N17772);
xor XOR2 (N17778, N17764, N5169);
or OR4 (N17779, N17778, N2628, N13022, N15101);
or OR4 (N17780, N17775, N17075, N15938, N9173);
or OR3 (N17781, N17773, N11055, N108);
nand NAND4 (N17782, N17780, N2320, N8546, N12388);
and AND2 (N17783, N17770, N16870);
and AND3 (N17784, N17768, N13276, N12602);
or OR4 (N17785, N17776, N11162, N13754, N382);
buf BUF1 (N17786, N17785);
buf BUF1 (N17787, N17777);
nor NOR3 (N17788, N17774, N15435, N2642);
buf BUF1 (N17789, N17788);
nand NAND2 (N17790, N17786, N16136);
xor XOR2 (N17791, N17790, N11419);
nand NAND4 (N17792, N17781, N2618, N8997, N3690);
nand NAND3 (N17793, N17792, N5976, N12920);
and AND4 (N17794, N17791, N3009, N4295, N7216);
nor NOR2 (N17795, N17794, N8840);
or OR3 (N17796, N17779, N7223, N2992);
xor XOR2 (N17797, N17783, N1581);
buf BUF1 (N17798, N17793);
nor NOR2 (N17799, N17789, N14553);
not NOT1 (N17800, N17782);
xor XOR2 (N17801, N17799, N3550);
xor XOR2 (N17802, N17801, N1400);
or OR2 (N17803, N17796, N14590);
xor XOR2 (N17804, N17797, N6237);
or OR4 (N17805, N17795, N7237, N17556, N14285);
nand NAND3 (N17806, N17800, N15322, N12909);
nor NOR3 (N17807, N17802, N6622, N4380);
and AND4 (N17808, N17787, N7350, N9763, N5895);
and AND2 (N17809, N17798, N877);
buf BUF1 (N17810, N17803);
and AND4 (N17811, N17806, N3216, N10060, N3147);
xor XOR2 (N17812, N17810, N1369);
nand NAND2 (N17813, N17812, N11389);
buf BUF1 (N17814, N17811);
or OR4 (N17815, N17760, N2113, N1851, N10812);
and AND2 (N17816, N17769, N4417);
xor XOR2 (N17817, N17814, N5791);
xor XOR2 (N17818, N17784, N6439);
nand NAND3 (N17819, N17807, N5238, N4884);
buf BUF1 (N17820, N17817);
not NOT1 (N17821, N17815);
xor XOR2 (N17822, N17821, N3393);
and AND4 (N17823, N17819, N16354, N7262, N11739);
nand NAND3 (N17824, N17808, N15493, N9456);
not NOT1 (N17825, N17809);
and AND3 (N17826, N17818, N2432, N8279);
buf BUF1 (N17827, N17822);
or OR2 (N17828, N17804, N12597);
or OR2 (N17829, N17816, N150);
buf BUF1 (N17830, N17828);
buf BUF1 (N17831, N17827);
or OR4 (N17832, N17830, N7034, N10403, N14640);
not NOT1 (N17833, N17831);
not NOT1 (N17834, N17820);
and AND4 (N17835, N17813, N3559, N16338, N9561);
and AND2 (N17836, N17834, N6882);
or OR4 (N17837, N17823, N7108, N15133, N16230);
not NOT1 (N17838, N17835);
and AND3 (N17839, N17824, N10667, N9301);
xor XOR2 (N17840, N17805, N14007);
buf BUF1 (N17841, N17839);
not NOT1 (N17842, N17826);
nor NOR2 (N17843, N17829, N13667);
nor NOR3 (N17844, N17837, N17719, N15968);
xor XOR2 (N17845, N17843, N9884);
not NOT1 (N17846, N17842);
nand NAND2 (N17847, N17845, N15405);
nand NAND3 (N17848, N17847, N10041, N2242);
not NOT1 (N17849, N17825);
not NOT1 (N17850, N17844);
or OR3 (N17851, N17849, N13846, N16348);
or OR3 (N17852, N17836, N3136, N4678);
nor NOR3 (N17853, N17851, N912, N14299);
nand NAND3 (N17854, N17841, N12639, N5055);
or OR2 (N17855, N17848, N14904);
buf BUF1 (N17856, N17832);
not NOT1 (N17857, N17838);
nor NOR4 (N17858, N17856, N13812, N14563, N7078);
nand NAND2 (N17859, N17853, N9646);
nor NOR4 (N17860, N17854, N5725, N6357, N3797);
and AND3 (N17861, N17833, N1020, N6817);
xor XOR2 (N17862, N17860, N13462);
xor XOR2 (N17863, N17846, N3423);
and AND2 (N17864, N17862, N245);
nand NAND2 (N17865, N17852, N17059);
nor NOR3 (N17866, N17855, N17148, N8630);
buf BUF1 (N17867, N17865);
nand NAND4 (N17868, N17863, N15487, N6078, N12956);
nand NAND3 (N17869, N17868, N121, N10068);
nand NAND2 (N17870, N17866, N14741);
not NOT1 (N17871, N17861);
buf BUF1 (N17872, N17869);
buf BUF1 (N17873, N17867);
not NOT1 (N17874, N17872);
not NOT1 (N17875, N17857);
nor NOR3 (N17876, N17864, N15403, N12991);
nor NOR2 (N17877, N17840, N2384);
buf BUF1 (N17878, N17871);
not NOT1 (N17879, N17878);
nand NAND4 (N17880, N17876, N437, N11584, N1798);
nand NAND4 (N17881, N17880, N10608, N7369, N6845);
nand NAND3 (N17882, N17858, N1303, N11421);
buf BUF1 (N17883, N17870);
or OR3 (N17884, N17881, N9108, N3837);
nand NAND3 (N17885, N17850, N9644, N14765);
not NOT1 (N17886, N17877);
or OR3 (N17887, N17885, N14684, N2091);
or OR2 (N17888, N17873, N896);
xor XOR2 (N17889, N17874, N5652);
or OR2 (N17890, N17882, N1187);
or OR3 (N17891, N17884, N2781, N3907);
and AND2 (N17892, N17890, N7347);
nor NOR3 (N17893, N17887, N4528, N1108);
nand NAND4 (N17894, N17888, N1359, N253, N120);
nor NOR2 (N17895, N17859, N13833);
nor NOR2 (N17896, N17895, N5115);
nor NOR3 (N17897, N17886, N5984, N13138);
xor XOR2 (N17898, N17891, N10547);
xor XOR2 (N17899, N17898, N13096);
xor XOR2 (N17900, N17883, N503);
and AND4 (N17901, N17893, N3496, N7501, N14979);
and AND4 (N17902, N17889, N15118, N4377, N10508);
buf BUF1 (N17903, N17896);
buf BUF1 (N17904, N17894);
nor NOR4 (N17905, N17901, N17710, N17492, N13843);
nor NOR4 (N17906, N17903, N9316, N17500, N10813);
not NOT1 (N17907, N17904);
nor NOR2 (N17908, N17879, N3262);
nand NAND4 (N17909, N17907, N15922, N17207, N6314);
or OR3 (N17910, N17909, N13724, N6185);
not NOT1 (N17911, N17897);
not NOT1 (N17912, N17875);
or OR4 (N17913, N17899, N13240, N7428, N17334);
not NOT1 (N17914, N17908);
nor NOR4 (N17915, N17914, N1759, N3069, N1318);
or OR2 (N17916, N17912, N2241);
buf BUF1 (N17917, N17910);
nand NAND3 (N17918, N17892, N1356, N2959);
nor NOR2 (N17919, N17902, N10418);
and AND2 (N17920, N17919, N42);
nor NOR2 (N17921, N17905, N4937);
nand NAND2 (N17922, N17921, N15173);
or OR2 (N17923, N17920, N9389);
nor NOR4 (N17924, N17915, N13226, N15113, N16182);
or OR3 (N17925, N17923, N11097, N6184);
xor XOR2 (N17926, N17922, N11085);
nand NAND4 (N17927, N17911, N5664, N10545, N1311);
xor XOR2 (N17928, N17924, N2156);
xor XOR2 (N17929, N17925, N2877);
nand NAND2 (N17930, N17928, N3222);
not NOT1 (N17931, N17929);
buf BUF1 (N17932, N17931);
buf BUF1 (N17933, N17932);
or OR2 (N17934, N17926, N15614);
not NOT1 (N17935, N17933);
nor NOR3 (N17936, N17906, N12443, N5001);
xor XOR2 (N17937, N17936, N9810);
nor NOR3 (N17938, N17900, N4406, N15777);
xor XOR2 (N17939, N17938, N3544);
not NOT1 (N17940, N17935);
and AND3 (N17941, N17939, N14041, N12353);
xor XOR2 (N17942, N17937, N9640);
buf BUF1 (N17943, N17942);
buf BUF1 (N17944, N17916);
and AND4 (N17945, N17913, N11404, N791, N6574);
not NOT1 (N17946, N17930);
nand NAND4 (N17947, N17918, N4186, N1846, N14956);
not NOT1 (N17948, N17917);
or OR2 (N17949, N17941, N7215);
buf BUF1 (N17950, N17949);
nand NAND4 (N17951, N17945, N10192, N12787, N16941);
and AND4 (N17952, N17943, N1752, N205, N9890);
nand NAND2 (N17953, N17934, N6501);
nor NOR3 (N17954, N17951, N4005, N1072);
nor NOR3 (N17955, N17944, N14146, N3230);
xor XOR2 (N17956, N17953, N4814);
nor NOR4 (N17957, N17955, N792, N13260, N15107);
nor NOR3 (N17958, N17950, N3238, N7530);
xor XOR2 (N17959, N17948, N14120);
and AND2 (N17960, N17956, N13518);
nand NAND2 (N17961, N17952, N13443);
nor NOR2 (N17962, N17946, N7611);
and AND2 (N17963, N17959, N2601);
and AND2 (N17964, N17927, N1558);
or OR2 (N17965, N17962, N5820);
or OR4 (N17966, N17958, N16181, N6990, N10096);
nand NAND3 (N17967, N17966, N8950, N13379);
xor XOR2 (N17968, N17965, N14183);
not NOT1 (N17969, N17967);
not NOT1 (N17970, N17964);
nor NOR3 (N17971, N17963, N3128, N9861);
buf BUF1 (N17972, N17969);
xor XOR2 (N17973, N17960, N4627);
buf BUF1 (N17974, N17957);
xor XOR2 (N17975, N17970, N5304);
nor NOR2 (N17976, N17947, N15166);
nor NOR2 (N17977, N17971, N6190);
not NOT1 (N17978, N17974);
nor NOR4 (N17979, N17977, N3243, N15983, N9318);
nor NOR3 (N17980, N17975, N13779, N2680);
nand NAND2 (N17981, N17940, N9104);
not NOT1 (N17982, N17980);
nor NOR4 (N17983, N17954, N16299, N14119, N6501);
and AND4 (N17984, N17979, N14261, N1960, N12432);
or OR4 (N17985, N17961, N17221, N17352, N1120);
or OR2 (N17986, N17982, N13525);
or OR3 (N17987, N17972, N10870, N16325);
nand NAND3 (N17988, N17978, N12013, N8809);
or OR4 (N17989, N17973, N17191, N10474, N9217);
not NOT1 (N17990, N17981);
nand NAND3 (N17991, N17989, N7197, N237);
not NOT1 (N17992, N17976);
not NOT1 (N17993, N17987);
buf BUF1 (N17994, N17992);
and AND2 (N17995, N17993, N11047);
and AND2 (N17996, N17968, N4657);
buf BUF1 (N17997, N17988);
and AND4 (N17998, N17996, N17947, N10155, N15696);
and AND3 (N17999, N17997, N2449, N3258);
not NOT1 (N18000, N17990);
and AND4 (N18001, N17986, N4712, N10159, N5962);
or OR2 (N18002, N17985, N12949);
nor NOR3 (N18003, N17994, N14841, N8831);
and AND3 (N18004, N18003, N13835, N16307);
buf BUF1 (N18005, N18004);
nor NOR4 (N18006, N17983, N1723, N14231, N5885);
nor NOR2 (N18007, N17995, N897);
buf BUF1 (N18008, N18000);
buf BUF1 (N18009, N18008);
nor NOR4 (N18010, N18005, N14101, N14601, N117);
and AND4 (N18011, N18001, N3207, N2533, N5923);
buf BUF1 (N18012, N18010);
or OR2 (N18013, N18007, N8558);
not NOT1 (N18014, N18013);
nor NOR2 (N18015, N18006, N14703);
xor XOR2 (N18016, N18009, N14215);
buf BUF1 (N18017, N17984);
nor NOR4 (N18018, N18011, N840, N11232, N11559);
nor NOR3 (N18019, N18002, N10021, N11953);
nand NAND3 (N18020, N17998, N365, N341);
xor XOR2 (N18021, N18014, N231);
nor NOR4 (N18022, N18019, N4697, N15430, N2311);
or OR2 (N18023, N18016, N13233);
not NOT1 (N18024, N18021);
nor NOR2 (N18025, N17999, N8331);
buf BUF1 (N18026, N18012);
nand NAND3 (N18027, N18018, N11640, N11889);
buf BUF1 (N18028, N18027);
and AND4 (N18029, N18023, N9562, N17631, N4722);
xor XOR2 (N18030, N17991, N1726);
xor XOR2 (N18031, N18024, N6977);
buf BUF1 (N18032, N18025);
not NOT1 (N18033, N18029);
nand NAND4 (N18034, N18032, N5867, N12752, N8812);
xor XOR2 (N18035, N18030, N15368);
nand NAND2 (N18036, N18026, N16977);
or OR4 (N18037, N18033, N17336, N12995, N10645);
and AND4 (N18038, N18028, N12725, N15409, N13290);
not NOT1 (N18039, N18031);
not NOT1 (N18040, N18035);
nand NAND4 (N18041, N18034, N6993, N1315, N5026);
not NOT1 (N18042, N18041);
or OR3 (N18043, N18017, N8017, N5463);
buf BUF1 (N18044, N18039);
xor XOR2 (N18045, N18022, N2689);
not NOT1 (N18046, N18042);
nor NOR3 (N18047, N18020, N17274, N7893);
xor XOR2 (N18048, N18038, N10392);
nor NOR2 (N18049, N18040, N13759);
not NOT1 (N18050, N18046);
buf BUF1 (N18051, N18043);
nor NOR3 (N18052, N18047, N16786, N17194);
and AND3 (N18053, N18037, N4151, N2651);
nor NOR2 (N18054, N18048, N16050);
xor XOR2 (N18055, N18049, N649);
and AND4 (N18056, N18045, N13206, N14160, N14490);
not NOT1 (N18057, N18054);
or OR4 (N18058, N18052, N2615, N7983, N5558);
nand NAND3 (N18059, N18058, N1434, N12544);
and AND3 (N18060, N18057, N3088, N12071);
buf BUF1 (N18061, N18044);
buf BUF1 (N18062, N18051);
xor XOR2 (N18063, N18036, N15096);
and AND2 (N18064, N18063, N11964);
not NOT1 (N18065, N18062);
xor XOR2 (N18066, N18056, N5484);
or OR2 (N18067, N18064, N5467);
not NOT1 (N18068, N18050);
buf BUF1 (N18069, N18065);
or OR4 (N18070, N18068, N12051, N12384, N13502);
or OR2 (N18071, N18060, N796);
nor NOR3 (N18072, N18067, N7808, N4797);
xor XOR2 (N18073, N18015, N12328);
nor NOR2 (N18074, N18072, N4197);
nand NAND2 (N18075, N18059, N9457);
and AND2 (N18076, N18070, N5164);
nand NAND2 (N18077, N18073, N15708);
xor XOR2 (N18078, N18069, N11549);
nor NOR4 (N18079, N18078, N7143, N5309, N8068);
nor NOR4 (N18080, N18055, N4757, N12667, N579);
not NOT1 (N18081, N18075);
nor NOR2 (N18082, N18077, N10894);
buf BUF1 (N18083, N18076);
nor NOR4 (N18084, N18083, N5515, N15069, N5261);
and AND2 (N18085, N18084, N11266);
nor NOR4 (N18086, N18071, N7010, N269, N10275);
and AND2 (N18087, N18066, N14596);
buf BUF1 (N18088, N18079);
xor XOR2 (N18089, N18085, N6423);
buf BUF1 (N18090, N18082);
nor NOR2 (N18091, N18088, N2230);
xor XOR2 (N18092, N18053, N4233);
nor NOR3 (N18093, N18086, N11339, N614);
nor NOR3 (N18094, N18090, N12758, N16227);
xor XOR2 (N18095, N18094, N14280);
and AND3 (N18096, N18095, N17220, N3787);
and AND2 (N18097, N18092, N10051);
nand NAND2 (N18098, N18093, N10169);
not NOT1 (N18099, N18080);
xor XOR2 (N18100, N18061, N4776);
buf BUF1 (N18101, N18087);
not NOT1 (N18102, N18074);
nor NOR3 (N18103, N18091, N6186, N10060);
nand NAND2 (N18104, N18097, N10280);
buf BUF1 (N18105, N18096);
or OR4 (N18106, N18089, N8906, N14138, N5963);
and AND4 (N18107, N18106, N14053, N1624, N8760);
or OR4 (N18108, N18107, N17526, N9998, N6987);
xor XOR2 (N18109, N18100, N7250);
buf BUF1 (N18110, N18098);
nor NOR2 (N18111, N18099, N908);
nor NOR2 (N18112, N18108, N8259);
not NOT1 (N18113, N18105);
xor XOR2 (N18114, N18110, N10696);
nand NAND2 (N18115, N18111, N5323);
xor XOR2 (N18116, N18102, N4810);
and AND4 (N18117, N18109, N14984, N566, N9018);
and AND2 (N18118, N18113, N12980);
nand NAND4 (N18119, N18104, N2619, N8720, N11838);
not NOT1 (N18120, N18115);
not NOT1 (N18121, N18120);
and AND3 (N18122, N18118, N14095, N8612);
buf BUF1 (N18123, N18117);
buf BUF1 (N18124, N18121);
and AND2 (N18125, N18123, N1762);
buf BUF1 (N18126, N18103);
not NOT1 (N18127, N18114);
nand NAND3 (N18128, N18116, N7421, N10161);
and AND2 (N18129, N18124, N7470);
or OR2 (N18130, N18126, N15227);
nand NAND3 (N18131, N18125, N3014, N1438);
and AND2 (N18132, N18129, N12987);
nand NAND3 (N18133, N18131, N7423, N7239);
not NOT1 (N18134, N18112);
and AND4 (N18135, N18122, N8074, N15325, N9715);
buf BUF1 (N18136, N18134);
and AND4 (N18137, N18132, N17351, N7864, N12650);
xor XOR2 (N18138, N18128, N10160);
nand NAND3 (N18139, N18119, N2002, N7241);
not NOT1 (N18140, N18127);
nand NAND4 (N18141, N18130, N12127, N7194, N9404);
nor NOR2 (N18142, N18135, N7372);
nand NAND2 (N18143, N18139, N10246);
and AND4 (N18144, N18137, N10461, N8041, N14877);
nor NOR4 (N18145, N18144, N475, N12192, N11388);
nor NOR3 (N18146, N18133, N15693, N5374);
xor XOR2 (N18147, N18142, N15442);
xor XOR2 (N18148, N18136, N15700);
buf BUF1 (N18149, N18145);
nand NAND3 (N18150, N18140, N9344, N7875);
buf BUF1 (N18151, N18146);
nor NOR4 (N18152, N18081, N2858, N12950, N9457);
nor NOR3 (N18153, N18147, N16391, N8359);
buf BUF1 (N18154, N18151);
nand NAND2 (N18155, N18143, N15218);
and AND2 (N18156, N18148, N1786);
and AND2 (N18157, N18149, N6761);
buf BUF1 (N18158, N18154);
or OR4 (N18159, N18153, N6395, N3140, N18007);
buf BUF1 (N18160, N18156);
xor XOR2 (N18161, N18141, N1898);
and AND2 (N18162, N18150, N11047);
and AND3 (N18163, N18158, N15798, N9150);
and AND3 (N18164, N18152, N10957, N744);
not NOT1 (N18165, N18159);
xor XOR2 (N18166, N18161, N15188);
and AND4 (N18167, N18163, N15881, N14630, N5811);
or OR4 (N18168, N18160, N10783, N12854, N8105);
xor XOR2 (N18169, N18155, N11375);
not NOT1 (N18170, N18169);
buf BUF1 (N18171, N18170);
and AND4 (N18172, N18162, N17739, N4272, N15621);
buf BUF1 (N18173, N18171);
not NOT1 (N18174, N18173);
not NOT1 (N18175, N18172);
xor XOR2 (N18176, N18138, N8944);
nand NAND4 (N18177, N18176, N15786, N9145, N1425);
nor NOR4 (N18178, N18157, N14435, N4946, N16768);
nand NAND2 (N18179, N18164, N16693);
nand NAND2 (N18180, N18178, N8499);
xor XOR2 (N18181, N18167, N11105);
nor NOR2 (N18182, N18174, N12708);
buf BUF1 (N18183, N18179);
or OR4 (N18184, N18182, N14739, N4547, N4221);
buf BUF1 (N18185, N18175);
nor NOR4 (N18186, N18181, N8344, N6496, N270);
nor NOR3 (N18187, N18166, N2573, N4643);
or OR2 (N18188, N18168, N9517);
buf BUF1 (N18189, N18185);
not NOT1 (N18190, N18186);
buf BUF1 (N18191, N18101);
buf BUF1 (N18192, N18177);
not NOT1 (N18193, N18187);
buf BUF1 (N18194, N18188);
xor XOR2 (N18195, N18183, N15994);
xor XOR2 (N18196, N18193, N13128);
and AND3 (N18197, N18189, N16780, N11226);
xor XOR2 (N18198, N18195, N2213);
and AND4 (N18199, N18197, N570, N6550, N4760);
and AND2 (N18200, N18192, N4114);
or OR2 (N18201, N18200, N17631);
nand NAND3 (N18202, N18194, N6205, N1915);
nor NOR2 (N18203, N18202, N4014);
xor XOR2 (N18204, N18184, N761);
and AND3 (N18205, N18204, N8065, N12869);
buf BUF1 (N18206, N18196);
not NOT1 (N18207, N18201);
buf BUF1 (N18208, N18198);
and AND2 (N18209, N18205, N12916);
or OR4 (N18210, N18208, N14273, N11733, N13796);
not NOT1 (N18211, N18180);
not NOT1 (N18212, N18207);
or OR3 (N18213, N18190, N8585, N1210);
nor NOR4 (N18214, N18191, N17361, N7357, N351);
buf BUF1 (N18215, N18165);
xor XOR2 (N18216, N18206, N9335);
not NOT1 (N18217, N18211);
nand NAND2 (N18218, N18203, N7401);
nor NOR4 (N18219, N18213, N5149, N789, N8902);
and AND2 (N18220, N18209, N10956);
buf BUF1 (N18221, N18214);
or OR3 (N18222, N18220, N5220, N11163);
xor XOR2 (N18223, N18210, N11795);
buf BUF1 (N18224, N18223);
and AND3 (N18225, N18199, N17633, N9327);
buf BUF1 (N18226, N18212);
xor XOR2 (N18227, N18216, N12065);
not NOT1 (N18228, N18227);
or OR4 (N18229, N18228, N10112, N12264, N15229);
xor XOR2 (N18230, N18224, N18015);
xor XOR2 (N18231, N18222, N17082);
not NOT1 (N18232, N18225);
nand NAND3 (N18233, N18217, N17599, N10087);
not NOT1 (N18234, N18229);
nor NOR4 (N18235, N18232, N4877, N534, N12204);
xor XOR2 (N18236, N18215, N10875);
nor NOR4 (N18237, N18226, N8273, N7904, N4157);
and AND4 (N18238, N18231, N11826, N969, N14459);
buf BUF1 (N18239, N18218);
xor XOR2 (N18240, N18237, N6690);
xor XOR2 (N18241, N18239, N6876);
and AND4 (N18242, N18241, N3781, N14445, N14692);
buf BUF1 (N18243, N18240);
and AND3 (N18244, N18219, N4979, N15690);
or OR3 (N18245, N18244, N7806, N17971);
nor NOR2 (N18246, N18238, N3035);
buf BUF1 (N18247, N18242);
xor XOR2 (N18248, N18230, N1990);
or OR2 (N18249, N18236, N1212);
nand NAND4 (N18250, N18246, N2127, N4015, N17485);
xor XOR2 (N18251, N18249, N8824);
not NOT1 (N18252, N18243);
nor NOR2 (N18253, N18233, N7471);
buf BUF1 (N18254, N18250);
not NOT1 (N18255, N18247);
nand NAND4 (N18256, N18235, N7824, N15288, N698);
nand NAND3 (N18257, N18253, N11362, N5392);
not NOT1 (N18258, N18245);
nand NAND2 (N18259, N18234, N14545);
nor NOR3 (N18260, N18255, N1216, N692);
or OR4 (N18261, N18254, N6587, N12604, N8055);
and AND4 (N18262, N18251, N5254, N12641, N1408);
xor XOR2 (N18263, N18262, N16034);
or OR4 (N18264, N18256, N8744, N7630, N2980);
nor NOR3 (N18265, N18260, N4941, N14461);
nor NOR3 (N18266, N18252, N1819, N1433);
and AND4 (N18267, N18264, N12095, N7074, N3619);
not NOT1 (N18268, N18267);
xor XOR2 (N18269, N18248, N3376);
buf BUF1 (N18270, N18265);
nor NOR4 (N18271, N18268, N7488, N8910, N1904);
or OR4 (N18272, N18259, N16528, N1462, N8658);
nor NOR4 (N18273, N18272, N10334, N5615, N9407);
buf BUF1 (N18274, N18261);
and AND3 (N18275, N18221, N5830, N8383);
buf BUF1 (N18276, N18274);
not NOT1 (N18277, N18275);
xor XOR2 (N18278, N18270, N16286);
and AND4 (N18279, N18273, N13889, N1335, N5481);
or OR3 (N18280, N18279, N9267, N725);
and AND2 (N18281, N18278, N8830);
or OR2 (N18282, N18277, N5231);
xor XOR2 (N18283, N18257, N7201);
and AND3 (N18284, N18276, N4294, N11049);
nor NOR4 (N18285, N18284, N11469, N8750, N10530);
not NOT1 (N18286, N18269);
nand NAND3 (N18287, N18280, N6397, N4654);
and AND2 (N18288, N18258, N17250);
and AND2 (N18289, N18282, N10842);
nand NAND4 (N18290, N18281, N14530, N16698, N5547);
and AND2 (N18291, N18288, N9430);
nand NAND4 (N18292, N18271, N7830, N1308, N13422);
xor XOR2 (N18293, N18287, N6613);
buf BUF1 (N18294, N18289);
xor XOR2 (N18295, N18294, N17526);
nor NOR4 (N18296, N18286, N7376, N10361, N2473);
not NOT1 (N18297, N18263);
xor XOR2 (N18298, N18285, N2423);
and AND4 (N18299, N18298, N10551, N6215, N14622);
buf BUF1 (N18300, N18295);
xor XOR2 (N18301, N18299, N17281);
nor NOR4 (N18302, N18290, N18160, N14527, N15832);
and AND3 (N18303, N18300, N5845, N13548);
or OR3 (N18304, N18296, N7322, N17264);
and AND3 (N18305, N18283, N3324, N14758);
not NOT1 (N18306, N18304);
nand NAND4 (N18307, N18291, N5298, N1629, N13164);
nand NAND2 (N18308, N18307, N13583);
nand NAND4 (N18309, N18308, N7892, N17385, N433);
not NOT1 (N18310, N18303);
buf BUF1 (N18311, N18266);
and AND3 (N18312, N18292, N4935, N16482);
xor XOR2 (N18313, N18306, N5454);
and AND4 (N18314, N18313, N5816, N14507, N1324);
xor XOR2 (N18315, N18293, N1004);
nand NAND2 (N18316, N18302, N12595);
not NOT1 (N18317, N18309);
or OR3 (N18318, N18317, N7903, N7282);
and AND3 (N18319, N18311, N2519, N14579);
nand NAND3 (N18320, N18314, N6831, N9416);
xor XOR2 (N18321, N18310, N16946);
and AND4 (N18322, N18312, N8433, N9207, N859);
nor NOR3 (N18323, N18315, N1123, N4170);
xor XOR2 (N18324, N18321, N1604);
not NOT1 (N18325, N18323);
nor NOR4 (N18326, N18320, N9272, N8106, N672);
or OR4 (N18327, N18324, N13899, N17590, N5286);
or OR3 (N18328, N18326, N14223, N3676);
xor XOR2 (N18329, N18325, N837);
not NOT1 (N18330, N18301);
xor XOR2 (N18331, N18319, N1894);
or OR2 (N18332, N18322, N10694);
nor NOR4 (N18333, N18305, N11778, N15194, N11049);
or OR3 (N18334, N18328, N10749, N5875);
xor XOR2 (N18335, N18318, N306);
and AND2 (N18336, N18330, N8791);
or OR2 (N18337, N18316, N3007);
xor XOR2 (N18338, N18327, N10826);
xor XOR2 (N18339, N18329, N14986);
and AND3 (N18340, N18332, N5644, N918);
nand NAND3 (N18341, N18338, N17123, N17776);
or OR4 (N18342, N18333, N916, N12512, N15303);
xor XOR2 (N18343, N18342, N4054);
not NOT1 (N18344, N18336);
nand NAND4 (N18345, N18334, N8440, N7910, N2414);
not NOT1 (N18346, N18345);
or OR2 (N18347, N18335, N12578);
buf BUF1 (N18348, N18344);
not NOT1 (N18349, N18341);
nor NOR2 (N18350, N18346, N808);
and AND2 (N18351, N18349, N7294);
nor NOR3 (N18352, N18337, N1671, N17722);
and AND2 (N18353, N18347, N14755);
not NOT1 (N18354, N18340);
nand NAND3 (N18355, N18297, N13108, N6869);
not NOT1 (N18356, N18351);
not NOT1 (N18357, N18355);
nand NAND4 (N18358, N18356, N10659, N381, N15366);
not NOT1 (N18359, N18352);
nor NOR2 (N18360, N18339, N7193);
xor XOR2 (N18361, N18343, N3145);
xor XOR2 (N18362, N18359, N16062);
nor NOR4 (N18363, N18353, N8861, N14899, N10513);
not NOT1 (N18364, N18354);
or OR2 (N18365, N18362, N10589);
not NOT1 (N18366, N18365);
nor NOR3 (N18367, N18357, N3144, N17172);
or OR2 (N18368, N18363, N13104);
or OR4 (N18369, N18364, N236, N755, N7561);
and AND4 (N18370, N18331, N17977, N11189, N17739);
nand NAND2 (N18371, N18367, N9205);
not NOT1 (N18372, N18369);
nand NAND4 (N18373, N18368, N9863, N16344, N14874);
or OR2 (N18374, N18372, N9327);
nand NAND3 (N18375, N18360, N8866, N10909);
nor NOR3 (N18376, N18373, N11820, N3544);
nand NAND3 (N18377, N18350, N14163, N8713);
or OR2 (N18378, N18371, N890);
nor NOR2 (N18379, N18377, N7262);
buf BUF1 (N18380, N18375);
xor XOR2 (N18381, N18380, N1958);
buf BUF1 (N18382, N18376);
xor XOR2 (N18383, N18370, N4247);
buf BUF1 (N18384, N18379);
buf BUF1 (N18385, N18383);
nand NAND2 (N18386, N18348, N11952);
buf BUF1 (N18387, N18385);
xor XOR2 (N18388, N18374, N9304);
or OR3 (N18389, N18388, N17723, N1354);
or OR2 (N18390, N18382, N10178);
buf BUF1 (N18391, N18361);
nor NOR4 (N18392, N18387, N3667, N15136, N8245);
not NOT1 (N18393, N18381);
buf BUF1 (N18394, N18378);
nor NOR3 (N18395, N18390, N11209, N2357);
xor XOR2 (N18396, N18389, N10868);
nand NAND3 (N18397, N18366, N379, N16824);
not NOT1 (N18398, N18396);
and AND4 (N18399, N18395, N15232, N15987, N3056);
not NOT1 (N18400, N18398);
and AND2 (N18401, N18391, N15715);
nand NAND4 (N18402, N18397, N9763, N6409, N16648);
not NOT1 (N18403, N18358);
nor NOR4 (N18404, N18399, N796, N894, N1905);
buf BUF1 (N18405, N18401);
nor NOR2 (N18406, N18402, N7048);
xor XOR2 (N18407, N18386, N11277);
buf BUF1 (N18408, N18393);
buf BUF1 (N18409, N18392);
and AND2 (N18410, N18394, N1354);
and AND2 (N18411, N18409, N9584);
nor NOR4 (N18412, N18411, N15246, N16814, N17826);
xor XOR2 (N18413, N18410, N1618);
buf BUF1 (N18414, N18403);
or OR3 (N18415, N18408, N158, N12915);
nand NAND2 (N18416, N18407, N3919);
not NOT1 (N18417, N18405);
xor XOR2 (N18418, N18416, N10958);
or OR2 (N18419, N18415, N14041);
nand NAND4 (N18420, N18384, N6902, N3895, N7388);
xor XOR2 (N18421, N18419, N7118);
xor XOR2 (N18422, N18414, N16488);
xor XOR2 (N18423, N18421, N16350);
xor XOR2 (N18424, N18400, N4590);
or OR4 (N18425, N18418, N702, N13933, N9913);
nor NOR3 (N18426, N18412, N3033, N15897);
nor NOR4 (N18427, N18426, N1268, N8426, N5260);
and AND4 (N18428, N18417, N18196, N8663, N12483);
nor NOR4 (N18429, N18428, N17073, N5880, N8210);
nor NOR2 (N18430, N18425, N5386);
and AND2 (N18431, N18406, N17437);
not NOT1 (N18432, N18413);
nand NAND2 (N18433, N18430, N13568);
and AND3 (N18434, N18433, N9130, N8276);
and AND2 (N18435, N18422, N11878);
xor XOR2 (N18436, N18424, N773);
nor NOR2 (N18437, N18435, N1560);
and AND4 (N18438, N18423, N16648, N6646, N9871);
not NOT1 (N18439, N18427);
not NOT1 (N18440, N18404);
and AND4 (N18441, N18420, N16626, N6741, N12268);
nand NAND2 (N18442, N18432, N7796);
not NOT1 (N18443, N18442);
buf BUF1 (N18444, N18441);
xor XOR2 (N18445, N18436, N12746);
not NOT1 (N18446, N18437);
buf BUF1 (N18447, N18443);
and AND2 (N18448, N18445, N11330);
not NOT1 (N18449, N18429);
xor XOR2 (N18450, N18439, N6063);
or OR4 (N18451, N18449, N12876, N540, N4459);
xor XOR2 (N18452, N18431, N12882);
buf BUF1 (N18453, N18434);
nand NAND4 (N18454, N18444, N9076, N8459, N18087);
and AND2 (N18455, N18440, N2082);
xor XOR2 (N18456, N18446, N3364);
and AND2 (N18457, N18447, N16084);
or OR3 (N18458, N18450, N17872, N2476);
nand NAND4 (N18459, N18451, N5804, N2451, N17034);
xor XOR2 (N18460, N18457, N17670);
xor XOR2 (N18461, N18456, N2413);
not NOT1 (N18462, N18461);
xor XOR2 (N18463, N18448, N16800);
buf BUF1 (N18464, N18462);
buf BUF1 (N18465, N18459);
buf BUF1 (N18466, N18454);
and AND3 (N18467, N18438, N3422, N15921);
buf BUF1 (N18468, N18464);
nor NOR4 (N18469, N18463, N1596, N10569, N8970);
and AND3 (N18470, N18467, N13482, N14454);
buf BUF1 (N18471, N18465);
and AND4 (N18472, N18458, N9936, N16528, N11562);
nand NAND3 (N18473, N18472, N12183, N5347);
xor XOR2 (N18474, N18453, N18230);
xor XOR2 (N18475, N18473, N7812);
buf BUF1 (N18476, N18455);
xor XOR2 (N18477, N18460, N5115);
xor XOR2 (N18478, N18452, N7420);
or OR2 (N18479, N18475, N1099);
and AND3 (N18480, N18476, N18370, N4816);
nand NAND4 (N18481, N18478, N13840, N7451, N2266);
nand NAND3 (N18482, N18481, N11456, N1668);
nand NAND3 (N18483, N18471, N5634, N17246);
xor XOR2 (N18484, N18469, N9375);
buf BUF1 (N18485, N18477);
nand NAND2 (N18486, N18474, N4775);
nor NOR2 (N18487, N18483, N13285);
and AND4 (N18488, N18485, N15165, N15358, N6642);
and AND3 (N18489, N18487, N14693, N1084);
nor NOR2 (N18490, N18489, N1259);
and AND3 (N18491, N18488, N1451, N1737);
nand NAND2 (N18492, N18466, N11927);
nand NAND4 (N18493, N18479, N14340, N1068, N10933);
buf BUF1 (N18494, N18480);
or OR3 (N18495, N18491, N12062, N18280);
nor NOR2 (N18496, N18493, N13431);
nor NOR3 (N18497, N18494, N4130, N8260);
xor XOR2 (N18498, N18495, N1824);
nor NOR2 (N18499, N18490, N8477);
xor XOR2 (N18500, N18492, N5210);
and AND2 (N18501, N18499, N12803);
buf BUF1 (N18502, N18468);
or OR2 (N18503, N18497, N18340);
not NOT1 (N18504, N18503);
and AND2 (N18505, N18502, N8093);
nand NAND3 (N18506, N18498, N14033, N4021);
and AND4 (N18507, N18482, N9739, N4189, N11616);
nand NAND3 (N18508, N18505, N16754, N11760);
xor XOR2 (N18509, N18508, N18136);
nor NOR4 (N18510, N18509, N4200, N14031, N7777);
xor XOR2 (N18511, N18504, N12915);
and AND4 (N18512, N18501, N6092, N17267, N1645);
nand NAND3 (N18513, N18507, N2391, N4696);
not NOT1 (N18514, N18512);
nand NAND3 (N18515, N18486, N3096, N13426);
buf BUF1 (N18516, N18510);
nor NOR2 (N18517, N18484, N13908);
nand NAND2 (N18518, N18496, N8851);
not NOT1 (N18519, N18516);
not NOT1 (N18520, N18519);
nor NOR3 (N18521, N18520, N7928, N13472);
or OR2 (N18522, N18500, N12522);
or OR4 (N18523, N18521, N8333, N6927, N16423);
not NOT1 (N18524, N18522);
xor XOR2 (N18525, N18517, N13942);
not NOT1 (N18526, N18506);
nand NAND3 (N18527, N18518, N17230, N5179);
not NOT1 (N18528, N18524);
and AND4 (N18529, N18470, N8879, N6052, N16940);
nand NAND2 (N18530, N18529, N3408);
xor XOR2 (N18531, N18511, N7876);
xor XOR2 (N18532, N18523, N18447);
and AND3 (N18533, N18531, N15558, N12792);
not NOT1 (N18534, N18525);
xor XOR2 (N18535, N18515, N371);
nand NAND2 (N18536, N18535, N9671);
or OR3 (N18537, N18528, N9549, N16406);
xor XOR2 (N18538, N18537, N14436);
or OR3 (N18539, N18536, N7334, N15535);
not NOT1 (N18540, N18539);
or OR4 (N18541, N18526, N9796, N1512, N17797);
and AND3 (N18542, N18534, N2796, N11046);
buf BUF1 (N18543, N18542);
nand NAND4 (N18544, N18540, N7602, N15425, N4811);
not NOT1 (N18545, N18514);
nor NOR4 (N18546, N18532, N14288, N11762, N12474);
nor NOR2 (N18547, N18543, N15012);
xor XOR2 (N18548, N18513, N17914);
xor XOR2 (N18549, N18538, N11429);
buf BUF1 (N18550, N18546);
buf BUF1 (N18551, N18545);
or OR2 (N18552, N18548, N14754);
nor NOR3 (N18553, N18527, N7600, N10414);
nand NAND3 (N18554, N18551, N3504, N8518);
buf BUF1 (N18555, N18541);
buf BUF1 (N18556, N18554);
nand NAND3 (N18557, N18553, N14339, N9983);
buf BUF1 (N18558, N18555);
nand NAND3 (N18559, N18556, N5499, N14561);
buf BUF1 (N18560, N18559);
buf BUF1 (N18561, N18558);
buf BUF1 (N18562, N18530);
buf BUF1 (N18563, N18562);
not NOT1 (N18564, N18544);
and AND2 (N18565, N18552, N3815);
and AND3 (N18566, N18563, N16831, N11776);
buf BUF1 (N18567, N18565);
and AND3 (N18568, N18550, N4227, N4003);
nand NAND3 (N18569, N18547, N1880, N8255);
nor NOR3 (N18570, N18564, N8715, N12031);
nor NOR2 (N18571, N18561, N15295);
nor NOR3 (N18572, N18567, N3088, N4735);
xor XOR2 (N18573, N18549, N4496);
not NOT1 (N18574, N18571);
not NOT1 (N18575, N18572);
xor XOR2 (N18576, N18557, N17892);
and AND2 (N18577, N18533, N3630);
buf BUF1 (N18578, N18569);
nor NOR3 (N18579, N18560, N17289, N12195);
and AND3 (N18580, N18573, N4230, N13191);
xor XOR2 (N18581, N18576, N12430);
or OR2 (N18582, N18570, N10043);
buf BUF1 (N18583, N18581);
xor XOR2 (N18584, N18583, N2325);
or OR4 (N18585, N18568, N13064, N15932, N4827);
nor NOR4 (N18586, N18574, N15307, N15890, N8507);
nor NOR3 (N18587, N18580, N15324, N4011);
nor NOR2 (N18588, N18582, N6408);
xor XOR2 (N18589, N18577, N1519);
not NOT1 (N18590, N18579);
not NOT1 (N18591, N18590);
nand NAND4 (N18592, N18589, N11220, N1746, N71);
and AND3 (N18593, N18578, N9699, N10361);
or OR4 (N18594, N18592, N8627, N488, N18336);
nor NOR2 (N18595, N18586, N11644);
or OR2 (N18596, N18575, N15975);
xor XOR2 (N18597, N18584, N8362);
nand NAND4 (N18598, N18596, N13551, N5469, N11871);
nand NAND3 (N18599, N18585, N10079, N17320);
xor XOR2 (N18600, N18591, N1315);
nand NAND2 (N18601, N18587, N677);
or OR2 (N18602, N18594, N10285);
or OR3 (N18603, N18595, N3089, N15254);
buf BUF1 (N18604, N18566);
nor NOR4 (N18605, N18588, N18555, N6477, N7930);
or OR4 (N18606, N18598, N7655, N10227, N16663);
nand NAND2 (N18607, N18606, N8737);
or OR4 (N18608, N18597, N3860, N7257, N4771);
nor NOR2 (N18609, N18593, N9089);
nor NOR2 (N18610, N18605, N6833);
nor NOR2 (N18611, N18607, N1417);
or OR2 (N18612, N18610, N17810);
buf BUF1 (N18613, N18599);
not NOT1 (N18614, N18611);
nor NOR4 (N18615, N18601, N9390, N18516, N8033);
or OR2 (N18616, N18609, N1606);
or OR3 (N18617, N18616, N1705, N14306);
nand NAND2 (N18618, N18617, N18004);
nand NAND3 (N18619, N18614, N360, N206);
xor XOR2 (N18620, N18608, N8600);
or OR3 (N18621, N18615, N7879, N3683);
not NOT1 (N18622, N18621);
nand NAND3 (N18623, N18613, N250, N13585);
and AND4 (N18624, N18619, N13890, N12786, N17977);
or OR3 (N18625, N18603, N6510, N1359);
or OR3 (N18626, N18600, N13708, N5472);
and AND2 (N18627, N18622, N12693);
and AND2 (N18628, N18620, N15360);
and AND3 (N18629, N18618, N15857, N159);
nand NAND4 (N18630, N18602, N13913, N16976, N6829);
or OR3 (N18631, N18630, N13286, N9469);
nor NOR3 (N18632, N18612, N3410, N17618);
not NOT1 (N18633, N18624);
nor NOR4 (N18634, N18632, N16215, N2920, N10600);
and AND3 (N18635, N18623, N676, N18204);
xor XOR2 (N18636, N18604, N1119);
buf BUF1 (N18637, N18635);
nor NOR3 (N18638, N18631, N12124, N10345);
buf BUF1 (N18639, N18638);
xor XOR2 (N18640, N18637, N13302);
or OR3 (N18641, N18636, N11941, N4678);
nand NAND3 (N18642, N18626, N2448, N11133);
and AND4 (N18643, N18625, N15636, N81, N6973);
not NOT1 (N18644, N18643);
xor XOR2 (N18645, N18627, N18293);
xor XOR2 (N18646, N18639, N12392);
and AND4 (N18647, N18641, N2591, N8419, N5670);
nand NAND4 (N18648, N18634, N9128, N6190, N8603);
and AND4 (N18649, N18640, N5936, N17120, N2260);
and AND3 (N18650, N18649, N948, N7391);
not NOT1 (N18651, N18628);
xor XOR2 (N18652, N18646, N17270);
buf BUF1 (N18653, N18650);
not NOT1 (N18654, N18648);
and AND2 (N18655, N18642, N4359);
nand NAND2 (N18656, N18654, N16929);
nor NOR3 (N18657, N18633, N11626, N12124);
and AND3 (N18658, N18629, N3205, N4833);
buf BUF1 (N18659, N18657);
buf BUF1 (N18660, N18645);
and AND2 (N18661, N18659, N12874);
and AND4 (N18662, N18660, N9195, N15530, N16866);
nand NAND4 (N18663, N18644, N7939, N641, N512);
and AND3 (N18664, N18653, N18021, N5823);
or OR3 (N18665, N18652, N13207, N4699);
nand NAND4 (N18666, N18655, N4369, N4132, N11530);
nand NAND4 (N18667, N18661, N6078, N15212, N13766);
nor NOR4 (N18668, N18665, N15889, N14814, N11989);
and AND4 (N18669, N18666, N9637, N11946, N6943);
and AND2 (N18670, N18669, N2362);
or OR2 (N18671, N18668, N15304);
buf BUF1 (N18672, N18670);
xor XOR2 (N18673, N18663, N5431);
nand NAND4 (N18674, N18673, N9879, N9680, N6906);
buf BUF1 (N18675, N18672);
nor NOR2 (N18676, N18664, N1049);
nand NAND3 (N18677, N18671, N18407, N17098);
xor XOR2 (N18678, N18647, N4365);
nor NOR3 (N18679, N18675, N17437, N12804);
nor NOR3 (N18680, N18667, N18079, N18630);
xor XOR2 (N18681, N18674, N8438);
nor NOR2 (N18682, N18662, N13426);
or OR4 (N18683, N18651, N15267, N3945, N15498);
and AND2 (N18684, N18682, N14544);
buf BUF1 (N18685, N18656);
nor NOR2 (N18686, N18683, N3412);
not NOT1 (N18687, N18681);
nor NOR4 (N18688, N18684, N2380, N3867, N1309);
nor NOR2 (N18689, N18676, N12510);
nand NAND2 (N18690, N18679, N15678);
not NOT1 (N18691, N18686);
xor XOR2 (N18692, N18677, N2402);
nand NAND4 (N18693, N18688, N11608, N670, N2994);
nor NOR3 (N18694, N18658, N14394, N11308);
nor NOR3 (N18695, N18680, N3913, N16240);
nor NOR2 (N18696, N18693, N6462);
nor NOR2 (N18697, N18695, N14190);
nand NAND4 (N18698, N18687, N13307, N9059, N5381);
buf BUF1 (N18699, N18690);
and AND3 (N18700, N18699, N15565, N11810);
and AND4 (N18701, N18697, N133, N9135, N8423);
and AND4 (N18702, N18698, N7124, N18037, N10807);
nand NAND2 (N18703, N18685, N7153);
xor XOR2 (N18704, N18700, N11415);
nor NOR2 (N18705, N18704, N545);
xor XOR2 (N18706, N18678, N15358);
not NOT1 (N18707, N18691);
not NOT1 (N18708, N18692);
buf BUF1 (N18709, N18689);
nand NAND2 (N18710, N18701, N5195);
not NOT1 (N18711, N18702);
buf BUF1 (N18712, N18710);
or OR4 (N18713, N18712, N5250, N10060, N17984);
not NOT1 (N18714, N18696);
xor XOR2 (N18715, N18711, N5000);
nor NOR4 (N18716, N18708, N13922, N8735, N2256);
xor XOR2 (N18717, N18714, N12878);
or OR2 (N18718, N18709, N13694);
and AND4 (N18719, N18716, N918, N10222, N8147);
buf BUF1 (N18720, N18715);
nor NOR3 (N18721, N18720, N11396, N2027);
not NOT1 (N18722, N18707);
nand NAND2 (N18723, N18722, N842);
and AND3 (N18724, N18721, N17997, N12589);
not NOT1 (N18725, N18723);
nand NAND2 (N18726, N18706, N686);
buf BUF1 (N18727, N18726);
xor XOR2 (N18728, N18713, N1220);
not NOT1 (N18729, N18719);
not NOT1 (N18730, N18694);
or OR4 (N18731, N18725, N1079, N16743, N17000);
buf BUF1 (N18732, N18728);
nand NAND3 (N18733, N18703, N16773, N6034);
not NOT1 (N18734, N18705);
or OR2 (N18735, N18724, N1190);
nand NAND2 (N18736, N18727, N9947);
not NOT1 (N18737, N18734);
not NOT1 (N18738, N18736);
nand NAND2 (N18739, N18730, N5987);
buf BUF1 (N18740, N18735);
not NOT1 (N18741, N18729);
nor NOR3 (N18742, N18741, N8951, N17127);
xor XOR2 (N18743, N18739, N6702);
buf BUF1 (N18744, N18740);
nand NAND3 (N18745, N18731, N17930, N582);
xor XOR2 (N18746, N18745, N373);
not NOT1 (N18747, N18732);
not NOT1 (N18748, N18742);
nor NOR3 (N18749, N18746, N9528, N9151);
and AND4 (N18750, N18738, N18033, N12761, N1252);
nor NOR4 (N18751, N18737, N9876, N3517, N6840);
and AND4 (N18752, N18750, N6435, N1254, N4762);
nor NOR4 (N18753, N18718, N149, N5929, N3067);
nand NAND4 (N18754, N18744, N3565, N15801, N6308);
buf BUF1 (N18755, N18751);
or OR3 (N18756, N18755, N17102, N11537);
not NOT1 (N18757, N18747);
nor NOR4 (N18758, N18756, N16878, N2002, N1742);
or OR3 (N18759, N18754, N11567, N2967);
and AND4 (N18760, N18717, N976, N1483, N4322);
nor NOR4 (N18761, N18759, N2403, N13127, N6986);
nand NAND3 (N18762, N18753, N3151, N8972);
buf BUF1 (N18763, N18743);
buf BUF1 (N18764, N18760);
or OR3 (N18765, N18763, N2038, N12246);
and AND2 (N18766, N18764, N6253);
nand NAND2 (N18767, N18762, N5036);
buf BUF1 (N18768, N18748);
or OR3 (N18769, N18766, N11394, N11971);
not NOT1 (N18770, N18768);
xor XOR2 (N18771, N18758, N9187);
buf BUF1 (N18772, N18765);
not NOT1 (N18773, N18749);
or OR3 (N18774, N18761, N4441, N1214);
or OR2 (N18775, N18767, N11720);
xor XOR2 (N18776, N18757, N3131);
nor NOR3 (N18777, N18775, N5876, N11712);
and AND2 (N18778, N18769, N5786);
xor XOR2 (N18779, N18777, N18277);
buf BUF1 (N18780, N18774);
and AND4 (N18781, N18752, N18339, N9505, N15197);
buf BUF1 (N18782, N18779);
nand NAND3 (N18783, N18778, N7146, N2753);
nor NOR4 (N18784, N18783, N18468, N581, N14805);
xor XOR2 (N18785, N18780, N7807);
not NOT1 (N18786, N18772);
nand NAND2 (N18787, N18782, N1004);
and AND2 (N18788, N18784, N3586);
buf BUF1 (N18789, N18786);
nand NAND3 (N18790, N18773, N14386, N4361);
xor XOR2 (N18791, N18771, N1420);
nand NAND3 (N18792, N18770, N8080, N7954);
nand NAND2 (N18793, N18789, N9334);
or OR3 (N18794, N18792, N5753, N4433);
xor XOR2 (N18795, N18790, N7070);
not NOT1 (N18796, N18793);
xor XOR2 (N18797, N18787, N6642);
xor XOR2 (N18798, N18794, N5480);
nor NOR4 (N18799, N18796, N6030, N18647, N11016);
and AND4 (N18800, N18788, N15739, N6644, N10673);
or OR4 (N18801, N18797, N15016, N15085, N5363);
xor XOR2 (N18802, N18801, N1730);
not NOT1 (N18803, N18791);
not NOT1 (N18804, N18798);
and AND4 (N18805, N18781, N8535, N6542, N4681);
xor XOR2 (N18806, N18802, N276);
or OR4 (N18807, N18795, N11678, N6465, N4588);
and AND2 (N18808, N18804, N13304);
nor NOR3 (N18809, N18785, N16450, N8177);
buf BUF1 (N18810, N18733);
nor NOR3 (N18811, N18808, N12767, N5596);
and AND2 (N18812, N18806, N11748);
buf BUF1 (N18813, N18810);
not NOT1 (N18814, N18809);
or OR3 (N18815, N18803, N10110, N3968);
not NOT1 (N18816, N18799);
or OR3 (N18817, N18814, N14195, N8488);
buf BUF1 (N18818, N18807);
nand NAND4 (N18819, N18800, N6880, N10737, N3343);
buf BUF1 (N18820, N18812);
not NOT1 (N18821, N18813);
and AND2 (N18822, N18818, N18780);
not NOT1 (N18823, N18811);
nand NAND4 (N18824, N18823, N8860, N12262, N12111);
not NOT1 (N18825, N18815);
xor XOR2 (N18826, N18817, N15453);
buf BUF1 (N18827, N18826);
nand NAND3 (N18828, N18822, N5142, N1907);
and AND3 (N18829, N18827, N12215, N13292);
buf BUF1 (N18830, N18819);
nand NAND2 (N18831, N18820, N6148);
and AND3 (N18832, N18828, N1646, N9503);
buf BUF1 (N18833, N18821);
not NOT1 (N18834, N18805);
xor XOR2 (N18835, N18829, N6719);
and AND4 (N18836, N18776, N17809, N6067, N6764);
or OR2 (N18837, N18835, N6109);
buf BUF1 (N18838, N18825);
or OR3 (N18839, N18830, N7481, N3880);
or OR3 (N18840, N18824, N8446, N3627);
not NOT1 (N18841, N18837);
not NOT1 (N18842, N18836);
xor XOR2 (N18843, N18832, N13197);
xor XOR2 (N18844, N18834, N3837);
and AND4 (N18845, N18842, N12576, N18280, N2989);
buf BUF1 (N18846, N18845);
nor NOR3 (N18847, N18840, N2139, N16622);
not NOT1 (N18848, N18841);
and AND4 (N18849, N18839, N8342, N6908, N18641);
or OR4 (N18850, N18847, N6908, N16009, N14098);
not NOT1 (N18851, N18848);
and AND4 (N18852, N18849, N15585, N8736, N12712);
nand NAND4 (N18853, N18851, N14075, N6455, N16408);
nand NAND2 (N18854, N18844, N18518);
nand NAND2 (N18855, N18831, N542);
or OR2 (N18856, N18843, N12081);
xor XOR2 (N18857, N18838, N18307);
and AND3 (N18858, N18856, N2706, N12376);
and AND3 (N18859, N18833, N6471, N12505);
or OR3 (N18860, N18852, N9106, N15198);
buf BUF1 (N18861, N18816);
or OR2 (N18862, N18850, N2963);
and AND3 (N18863, N18859, N13000, N10194);
buf BUF1 (N18864, N18853);
or OR4 (N18865, N18855, N16947, N16171, N10535);
nand NAND3 (N18866, N18857, N9987, N8932);
nor NOR2 (N18867, N18866, N3807);
nand NAND2 (N18868, N18867, N11041);
buf BUF1 (N18869, N18863);
not NOT1 (N18870, N18862);
xor XOR2 (N18871, N18858, N7168);
nand NAND3 (N18872, N18870, N5339, N14143);
or OR2 (N18873, N18865, N11633);
nor NOR4 (N18874, N18861, N5563, N3593, N17640);
buf BUF1 (N18875, N18864);
and AND4 (N18876, N18872, N15458, N4709, N7790);
and AND3 (N18877, N18876, N14854, N8470);
and AND4 (N18878, N18860, N5643, N5596, N13631);
nor NOR3 (N18879, N18871, N16868, N14811);
nand NAND2 (N18880, N18869, N18263);
buf BUF1 (N18881, N18854);
not NOT1 (N18882, N18878);
nor NOR4 (N18883, N18881, N10607, N8703, N14190);
not NOT1 (N18884, N18846);
nand NAND3 (N18885, N18880, N4037, N254);
and AND4 (N18886, N18873, N7641, N11648, N16944);
xor XOR2 (N18887, N18883, N16721);
or OR4 (N18888, N18877, N7463, N15908, N17202);
buf BUF1 (N18889, N18885);
xor XOR2 (N18890, N18888, N4278);
and AND2 (N18891, N18879, N1100);
or OR3 (N18892, N18875, N14013, N14605);
and AND4 (N18893, N18874, N11751, N16127, N16354);
and AND4 (N18894, N18891, N2899, N14297, N13472);
or OR3 (N18895, N18884, N3335, N10803);
nor NOR4 (N18896, N18892, N17344, N11926, N16552);
or OR4 (N18897, N18882, N18077, N10715, N11309);
buf BUF1 (N18898, N18887);
not NOT1 (N18899, N18898);
xor XOR2 (N18900, N18889, N13556);
or OR2 (N18901, N18899, N1803);
buf BUF1 (N18902, N18886);
or OR2 (N18903, N18897, N8829);
and AND3 (N18904, N18900, N2847, N10756);
nor NOR2 (N18905, N18895, N11674);
nand NAND3 (N18906, N18903, N17229, N8876);
not NOT1 (N18907, N18902);
not NOT1 (N18908, N18904);
nor NOR4 (N18909, N18896, N13211, N12071, N12503);
nor NOR3 (N18910, N18906, N15001, N6516);
or OR3 (N18911, N18890, N14963, N18469);
buf BUF1 (N18912, N18909);
or OR2 (N18913, N18910, N18703);
buf BUF1 (N18914, N18894);
and AND4 (N18915, N18912, N2355, N18537, N11518);
buf BUF1 (N18916, N18905);
or OR2 (N18917, N18893, N15399);
and AND2 (N18918, N18915, N1336);
nor NOR2 (N18919, N18868, N11982);
buf BUF1 (N18920, N18919);
xor XOR2 (N18921, N18911, N14450);
xor XOR2 (N18922, N18918, N12023);
nor NOR3 (N18923, N18913, N12114, N4759);
or OR2 (N18924, N18917, N12116);
nand NAND3 (N18925, N18923, N17919, N9235);
and AND3 (N18926, N18907, N13006, N9268);
and AND2 (N18927, N18924, N1002);
or OR4 (N18928, N18921, N13537, N14256, N881);
nand NAND4 (N18929, N18925, N1942, N13556, N9681);
and AND3 (N18930, N18901, N11966, N2829);
not NOT1 (N18931, N18916);
nor NOR4 (N18932, N18929, N13251, N15888, N9003);
nor NOR4 (N18933, N18928, N2225, N3734, N17942);
not NOT1 (N18934, N18920);
nand NAND3 (N18935, N18926, N12369, N14970);
nor NOR2 (N18936, N18922, N12292);
not NOT1 (N18937, N18930);
or OR3 (N18938, N18931, N1148, N4192);
buf BUF1 (N18939, N18937);
not NOT1 (N18940, N18935);
nor NOR3 (N18941, N18936, N2635, N3150);
or OR4 (N18942, N18939, N1897, N5866, N3636);
not NOT1 (N18943, N18914);
and AND3 (N18944, N18927, N4002, N5257);
or OR4 (N18945, N18908, N14687, N18882, N16628);
nand NAND3 (N18946, N18943, N16908, N3940);
buf BUF1 (N18947, N18938);
and AND4 (N18948, N18940, N9662, N4004, N2814);
buf BUF1 (N18949, N18947);
nand NAND4 (N18950, N18944, N4041, N6354, N3698);
or OR4 (N18951, N18945, N15966, N5202, N10848);
xor XOR2 (N18952, N18934, N17972);
buf BUF1 (N18953, N18933);
or OR3 (N18954, N18948, N5522, N8159);
xor XOR2 (N18955, N18952, N14922);
and AND3 (N18956, N18955, N17464, N13436);
not NOT1 (N18957, N18951);
nand NAND3 (N18958, N18949, N6322, N10984);
nand NAND4 (N18959, N18950, N1504, N6106, N9903);
or OR3 (N18960, N18959, N12356, N13505);
not NOT1 (N18961, N18957);
not NOT1 (N18962, N18961);
nor NOR3 (N18963, N18932, N8320, N4741);
nor NOR4 (N18964, N18953, N5999, N3857, N375);
not NOT1 (N18965, N18954);
or OR4 (N18966, N18958, N9023, N18040, N9458);
not NOT1 (N18967, N18966);
and AND4 (N18968, N18962, N17879, N16599, N10290);
or OR4 (N18969, N18965, N2678, N5069, N12408);
not NOT1 (N18970, N18964);
buf BUF1 (N18971, N18963);
not NOT1 (N18972, N18970);
or OR4 (N18973, N18972, N18562, N4176, N2197);
and AND3 (N18974, N18968, N14942, N3445);
and AND4 (N18975, N18974, N5004, N9406, N1780);
or OR2 (N18976, N18956, N12327);
buf BUF1 (N18977, N18975);
buf BUF1 (N18978, N18941);
buf BUF1 (N18979, N18946);
and AND3 (N18980, N18967, N2587, N16754);
nor NOR3 (N18981, N18978, N14246, N4337);
buf BUF1 (N18982, N18969);
nor NOR4 (N18983, N18979, N3970, N5085, N42);
nand NAND4 (N18984, N18982, N15848, N2439, N1561);
not NOT1 (N18985, N18983);
not NOT1 (N18986, N18960);
buf BUF1 (N18987, N18977);
or OR2 (N18988, N18976, N11453);
xor XOR2 (N18989, N18985, N12781);
xor XOR2 (N18990, N18980, N15599);
xor XOR2 (N18991, N18988, N2561);
buf BUF1 (N18992, N18986);
or OR3 (N18993, N18973, N11492, N18553);
or OR2 (N18994, N18984, N18835);
nand NAND4 (N18995, N18981, N11759, N2428, N5420);
not NOT1 (N18996, N18990);
nand NAND4 (N18997, N18991, N930, N14570, N9516);
or OR2 (N18998, N18996, N7680);
not NOT1 (N18999, N18992);
not NOT1 (N19000, N18971);
not NOT1 (N19001, N18998);
and AND2 (N19002, N18989, N2147);
buf BUF1 (N19003, N18987);
nor NOR2 (N19004, N18995, N11290);
nand NAND4 (N19005, N18994, N219, N12170, N18516);
not NOT1 (N19006, N18997);
not NOT1 (N19007, N18942);
nand NAND4 (N19008, N19005, N695, N11747, N2736);
xor XOR2 (N19009, N19006, N16103);
or OR4 (N19010, N18993, N10174, N7139, N3052);
and AND4 (N19011, N19001, N7372, N16309, N1581);
buf BUF1 (N19012, N19004);
not NOT1 (N19013, N19002);
and AND4 (N19014, N19013, N7122, N11595, N16772);
not NOT1 (N19015, N19003);
buf BUF1 (N19016, N19012);
or OR2 (N19017, N18999, N11973);
or OR4 (N19018, N19008, N13490, N18746, N120);
or OR2 (N19019, N19011, N7615);
not NOT1 (N19020, N19015);
xor XOR2 (N19021, N19018, N18553);
or OR3 (N19022, N19000, N10652, N11806);
nor NOR2 (N19023, N19021, N4583);
or OR2 (N19024, N19009, N2471);
buf BUF1 (N19025, N19016);
and AND4 (N19026, N19014, N8428, N12649, N15322);
and AND4 (N19027, N19022, N212, N539, N10968);
buf BUF1 (N19028, N19027);
nand NAND2 (N19029, N19023, N16786);
buf BUF1 (N19030, N19017);
buf BUF1 (N19031, N19026);
or OR4 (N19032, N19031, N16076, N12744, N18476);
buf BUF1 (N19033, N19020);
nor NOR3 (N19034, N19007, N5541, N4088);
and AND3 (N19035, N19030, N465, N2801);
nand NAND2 (N19036, N19033, N6791);
or OR3 (N19037, N19028, N12218, N8673);
xor XOR2 (N19038, N19010, N10017);
nand NAND3 (N19039, N19032, N12019, N10335);
nor NOR4 (N19040, N19025, N16543, N11751, N12580);
and AND3 (N19041, N19034, N2260, N3746);
nand NAND4 (N19042, N19029, N6824, N12091, N681);
nand NAND4 (N19043, N19041, N52, N10675, N18234);
xor XOR2 (N19044, N19040, N17003);
or OR2 (N19045, N19043, N13790);
not NOT1 (N19046, N19037);
nand NAND2 (N19047, N19044, N7519);
or OR4 (N19048, N19047, N12495, N3951, N15144);
xor XOR2 (N19049, N19019, N13799);
nor NOR3 (N19050, N19049, N11381, N8983);
not NOT1 (N19051, N19050);
nand NAND2 (N19052, N19035, N15459);
and AND3 (N19053, N19024, N18583, N7739);
xor XOR2 (N19054, N19052, N11505);
and AND3 (N19055, N19051, N122, N9021);
not NOT1 (N19056, N19042);
nand NAND2 (N19057, N19054, N7647);
not NOT1 (N19058, N19039);
nor NOR4 (N19059, N19053, N1057, N7729, N11993);
or OR2 (N19060, N19059, N16592);
buf BUF1 (N19061, N19038);
and AND4 (N19062, N19046, N5473, N9907, N3626);
nand NAND2 (N19063, N19060, N14773);
not NOT1 (N19064, N19048);
not NOT1 (N19065, N19062);
not NOT1 (N19066, N19056);
and AND2 (N19067, N19057, N16265);
or OR4 (N19068, N19065, N17101, N7100, N13906);
not NOT1 (N19069, N19067);
buf BUF1 (N19070, N19063);
xor XOR2 (N19071, N19068, N8834);
or OR2 (N19072, N19064, N1759);
xor XOR2 (N19073, N19069, N15785);
buf BUF1 (N19074, N19066);
nand NAND4 (N19075, N19055, N9898, N18997, N6480);
buf BUF1 (N19076, N19075);
buf BUF1 (N19077, N19071);
nand NAND4 (N19078, N19045, N6110, N61, N15244);
not NOT1 (N19079, N19078);
or OR3 (N19080, N19070, N16468, N11692);
xor XOR2 (N19081, N19077, N14093);
or OR3 (N19082, N19061, N1577, N13100);
or OR3 (N19083, N19036, N8700, N904);
nor NOR3 (N19084, N19073, N14066, N14054);
buf BUF1 (N19085, N19081);
not NOT1 (N19086, N19085);
buf BUF1 (N19087, N19074);
xor XOR2 (N19088, N19076, N11072);
or OR3 (N19089, N19080, N7696, N7921);
buf BUF1 (N19090, N19084);
or OR4 (N19091, N19090, N8518, N5072, N18960);
buf BUF1 (N19092, N19072);
or OR3 (N19093, N19089, N479, N1125);
not NOT1 (N19094, N19083);
or OR2 (N19095, N19092, N8361);
nor NOR4 (N19096, N19086, N3818, N444, N17088);
buf BUF1 (N19097, N19058);
not NOT1 (N19098, N19093);
xor XOR2 (N19099, N19091, N1336);
xor XOR2 (N19100, N19094, N9226);
and AND2 (N19101, N19098, N5046);
nor NOR3 (N19102, N19079, N7541, N16944);
or OR4 (N19103, N19102, N5650, N7315, N7261);
and AND2 (N19104, N19100, N14944);
not NOT1 (N19105, N19104);
and AND3 (N19106, N19097, N9641, N750);
buf BUF1 (N19107, N19082);
nand NAND2 (N19108, N19106, N18429);
nor NOR2 (N19109, N19105, N13157);
buf BUF1 (N19110, N19087);
or OR3 (N19111, N19088, N906, N787);
not NOT1 (N19112, N19095);
and AND2 (N19113, N19111, N9790);
not NOT1 (N19114, N19108);
and AND4 (N19115, N19101, N6305, N10866, N10821);
or OR3 (N19116, N19110, N9366, N9870);
or OR3 (N19117, N19109, N2487, N4731);
and AND3 (N19118, N19099, N6764, N12207);
nand NAND4 (N19119, N19114, N4464, N17905, N13388);
buf BUF1 (N19120, N19096);
nand NAND2 (N19121, N19115, N2084);
nand NAND4 (N19122, N19118, N13684, N3034, N3036);
buf BUF1 (N19123, N19112);
buf BUF1 (N19124, N19122);
and AND2 (N19125, N19116, N3174);
and AND2 (N19126, N19125, N2377);
xor XOR2 (N19127, N19126, N9627);
buf BUF1 (N19128, N19121);
not NOT1 (N19129, N19127);
nand NAND2 (N19130, N19103, N11645);
or OR2 (N19131, N19130, N15343);
and AND3 (N19132, N19123, N9679, N11310);
buf BUF1 (N19133, N19132);
or OR4 (N19134, N19107, N18192, N6750, N14068);
buf BUF1 (N19135, N19124);
nor NOR3 (N19136, N19129, N16832, N12742);
or OR4 (N19137, N19119, N14589, N1019, N12369);
and AND2 (N19138, N19136, N10419);
buf BUF1 (N19139, N19131);
xor XOR2 (N19140, N19113, N1638);
and AND4 (N19141, N19139, N3369, N2350, N8484);
nor NOR3 (N19142, N19135, N8603, N1167);
xor XOR2 (N19143, N19134, N3664);
xor XOR2 (N19144, N19141, N12006);
or OR2 (N19145, N19143, N6443);
not NOT1 (N19146, N19117);
not NOT1 (N19147, N19146);
and AND2 (N19148, N19140, N5231);
nand NAND3 (N19149, N19120, N26, N15959);
not NOT1 (N19150, N19138);
or OR2 (N19151, N19149, N495);
nor NOR4 (N19152, N19151, N18336, N531, N6278);
buf BUF1 (N19153, N19150);
buf BUF1 (N19154, N19133);
xor XOR2 (N19155, N19148, N14731);
xor XOR2 (N19156, N19152, N591);
buf BUF1 (N19157, N19137);
and AND3 (N19158, N19155, N9672, N3904);
nor NOR2 (N19159, N19157, N1103);
nor NOR3 (N19160, N19158, N456, N1225);
and AND3 (N19161, N19142, N7663, N5506);
nor NOR3 (N19162, N19154, N16514, N12120);
buf BUF1 (N19163, N19162);
or OR2 (N19164, N19128, N18500);
and AND4 (N19165, N19145, N10394, N15004, N9645);
buf BUF1 (N19166, N19147);
not NOT1 (N19167, N19165);
buf BUF1 (N19168, N19159);
nor NOR3 (N19169, N19163, N371, N1410);
buf BUF1 (N19170, N19168);
or OR4 (N19171, N19153, N8815, N1515, N9307);
not NOT1 (N19172, N19167);
not NOT1 (N19173, N19164);
nor NOR4 (N19174, N19161, N13534, N9851, N17444);
xor XOR2 (N19175, N19169, N15687);
and AND2 (N19176, N19166, N4183);
nand NAND2 (N19177, N19176, N14855);
or OR2 (N19178, N19172, N18775);
xor XOR2 (N19179, N19175, N5849);
xor XOR2 (N19180, N19156, N7601);
buf BUF1 (N19181, N19180);
buf BUF1 (N19182, N19144);
and AND4 (N19183, N19177, N11026, N12670, N2614);
xor XOR2 (N19184, N19179, N5572);
and AND2 (N19185, N19174, N16003);
nand NAND4 (N19186, N19182, N7322, N1067, N10851);
or OR4 (N19187, N19173, N10806, N18035, N18672);
or OR2 (N19188, N19160, N17744);
and AND3 (N19189, N19188, N3136, N3652);
nand NAND3 (N19190, N19187, N9278, N14081);
nand NAND3 (N19191, N19178, N13554, N6476);
and AND3 (N19192, N19189, N7111, N5965);
buf BUF1 (N19193, N19192);
nor NOR3 (N19194, N19181, N15303, N5070);
nand NAND2 (N19195, N19183, N11894);
nand NAND3 (N19196, N19171, N16472, N10122);
xor XOR2 (N19197, N19170, N12644);
not NOT1 (N19198, N19186);
not NOT1 (N19199, N19196);
xor XOR2 (N19200, N19199, N4336);
not NOT1 (N19201, N19190);
nor NOR3 (N19202, N19201, N12143, N4167);
nand NAND3 (N19203, N19202, N14307, N12034);
xor XOR2 (N19204, N19185, N18493);
or OR2 (N19205, N19204, N8338);
not NOT1 (N19206, N19203);
nand NAND3 (N19207, N19191, N9695, N2190);
buf BUF1 (N19208, N19197);
xor XOR2 (N19209, N19195, N4814);
nand NAND2 (N19210, N19207, N8915);
nand NAND3 (N19211, N19205, N156, N12983);
nor NOR3 (N19212, N19194, N11794, N16848);
buf BUF1 (N19213, N19208);
buf BUF1 (N19214, N19213);
nor NOR4 (N19215, N19184, N18103, N3119, N5558);
buf BUF1 (N19216, N19215);
not NOT1 (N19217, N19212);
buf BUF1 (N19218, N19210);
nor NOR4 (N19219, N19214, N16337, N5663, N953);
or OR2 (N19220, N19211, N998);
buf BUF1 (N19221, N19220);
or OR4 (N19222, N19198, N13297, N8563, N4171);
not NOT1 (N19223, N19217);
xor XOR2 (N19224, N19209, N16174);
not NOT1 (N19225, N19221);
buf BUF1 (N19226, N19206);
or OR3 (N19227, N19200, N8611, N19078);
and AND2 (N19228, N19218, N3265);
or OR2 (N19229, N19226, N2567);
xor XOR2 (N19230, N19229, N1698);
nand NAND4 (N19231, N19216, N13963, N15281, N33);
not NOT1 (N19232, N19193);
nor NOR2 (N19233, N19219, N9826);
not NOT1 (N19234, N19225);
and AND2 (N19235, N19223, N18304);
xor XOR2 (N19236, N19234, N2666);
nand NAND4 (N19237, N19233, N16654, N18473, N7065);
buf BUF1 (N19238, N19232);
xor XOR2 (N19239, N19231, N8283);
buf BUF1 (N19240, N19222);
xor XOR2 (N19241, N19239, N12008);
xor XOR2 (N19242, N19227, N5935);
not NOT1 (N19243, N19238);
and AND3 (N19244, N19241, N17612, N8911);
nand NAND3 (N19245, N19240, N13159, N15430);
not NOT1 (N19246, N19244);
or OR2 (N19247, N19246, N10);
and AND3 (N19248, N19242, N17255, N11325);
or OR2 (N19249, N19245, N11327);
nor NOR2 (N19250, N19235, N10594);
not NOT1 (N19251, N19236);
nand NAND2 (N19252, N19224, N6893);
or OR2 (N19253, N19251, N18930);
or OR2 (N19254, N19247, N14026);
or OR2 (N19255, N19237, N13253);
buf BUF1 (N19256, N19255);
or OR4 (N19257, N19249, N16355, N5894, N16296);
nand NAND3 (N19258, N19256, N10157, N5096);
nor NOR3 (N19259, N19258, N15949, N10335);
xor XOR2 (N19260, N19248, N13429);
or OR3 (N19261, N19257, N14930, N9832);
and AND2 (N19262, N19254, N8890);
nor NOR4 (N19263, N19230, N12844, N6157, N12674);
or OR3 (N19264, N19253, N2907, N15373);
xor XOR2 (N19265, N19243, N12550);
not NOT1 (N19266, N19263);
or OR2 (N19267, N19265, N18330);
and AND2 (N19268, N19252, N9149);
xor XOR2 (N19269, N19228, N19105);
nand NAND2 (N19270, N19268, N883);
not NOT1 (N19271, N19264);
not NOT1 (N19272, N19261);
nand NAND3 (N19273, N19272, N10870, N332);
and AND3 (N19274, N19259, N10227, N16295);
xor XOR2 (N19275, N19273, N6900);
not NOT1 (N19276, N19267);
or OR3 (N19277, N19270, N5212, N1749);
buf BUF1 (N19278, N19274);
or OR2 (N19279, N19271, N9007);
not NOT1 (N19280, N19260);
nand NAND4 (N19281, N19280, N15118, N15790, N4027);
buf BUF1 (N19282, N19278);
xor XOR2 (N19283, N19275, N4598);
nand NAND2 (N19284, N19281, N16338);
nand NAND4 (N19285, N19250, N17711, N3112, N2175);
not NOT1 (N19286, N19266);
nand NAND2 (N19287, N19284, N6595);
and AND2 (N19288, N19279, N7963);
xor XOR2 (N19289, N19287, N9373);
buf BUF1 (N19290, N19262);
and AND3 (N19291, N19289, N4447, N11486);
buf BUF1 (N19292, N19276);
not NOT1 (N19293, N19282);
nand NAND2 (N19294, N19291, N16441);
nand NAND2 (N19295, N19286, N6124);
or OR3 (N19296, N19283, N10673, N16011);
and AND4 (N19297, N19290, N4813, N2720, N9882);
not NOT1 (N19298, N19294);
nand NAND3 (N19299, N19296, N6681, N11436);
and AND2 (N19300, N19288, N16158);
or OR2 (N19301, N19269, N11866);
nand NAND4 (N19302, N19301, N5725, N7743, N14192);
xor XOR2 (N19303, N19277, N3647);
or OR3 (N19304, N19302, N12605, N9367);
not NOT1 (N19305, N19304);
or OR4 (N19306, N19292, N10950, N11921, N3081);
or OR2 (N19307, N19295, N13681);
or OR4 (N19308, N19300, N15327, N10810, N2728);
or OR2 (N19309, N19298, N2089);
not NOT1 (N19310, N19299);
xor XOR2 (N19311, N19310, N17200);
or OR2 (N19312, N19311, N4985);
and AND2 (N19313, N19308, N515);
buf BUF1 (N19314, N19306);
buf BUF1 (N19315, N19293);
or OR2 (N19316, N19285, N10715);
nand NAND4 (N19317, N19303, N3327, N1167, N7729);
not NOT1 (N19318, N19315);
or OR4 (N19319, N19317, N9923, N8895, N583);
xor XOR2 (N19320, N19307, N10017);
not NOT1 (N19321, N19297);
nand NAND2 (N19322, N19320, N1323);
buf BUF1 (N19323, N19314);
and AND3 (N19324, N19323, N10025, N8666);
nor NOR4 (N19325, N19321, N12055, N14287, N5563);
and AND3 (N19326, N19325, N8756, N10961);
nor NOR3 (N19327, N19324, N17680, N8410);
nor NOR2 (N19328, N19326, N15362);
buf BUF1 (N19329, N19327);
xor XOR2 (N19330, N19309, N6573);
nand NAND2 (N19331, N19316, N3865);
not NOT1 (N19332, N19330);
xor XOR2 (N19333, N19318, N18229);
not NOT1 (N19334, N19332);
not NOT1 (N19335, N19333);
buf BUF1 (N19336, N19335);
nor NOR4 (N19337, N19313, N6532, N2926, N13504);
nand NAND3 (N19338, N19319, N16954, N18036);
or OR2 (N19339, N19322, N5585);
xor XOR2 (N19340, N19334, N15174);
and AND2 (N19341, N19305, N17854);
not NOT1 (N19342, N19338);
nor NOR4 (N19343, N19339, N14853, N15490, N12830);
and AND3 (N19344, N19336, N1476, N2173);
not NOT1 (N19345, N19337);
or OR2 (N19346, N19342, N10150);
not NOT1 (N19347, N19312);
nor NOR3 (N19348, N19341, N13988, N1544);
not NOT1 (N19349, N19348);
nand NAND4 (N19350, N19331, N12291, N26, N10741);
or OR4 (N19351, N19346, N11689, N15725, N5016);
nand NAND3 (N19352, N19329, N6215, N16262);
nand NAND4 (N19353, N19347, N17976, N9282, N5846);
not NOT1 (N19354, N19352);
nand NAND3 (N19355, N19345, N12679, N2989);
nand NAND2 (N19356, N19355, N12778);
not NOT1 (N19357, N19349);
or OR4 (N19358, N19350, N16350, N12416, N17168);
buf BUF1 (N19359, N19351);
or OR4 (N19360, N19340, N12975, N10920, N18212);
buf BUF1 (N19361, N19343);
nor NOR2 (N19362, N19328, N19337);
xor XOR2 (N19363, N19354, N3924);
not NOT1 (N19364, N19363);
xor XOR2 (N19365, N19356, N9684);
xor XOR2 (N19366, N19361, N6953);
or OR2 (N19367, N19344, N13844);
nand NAND4 (N19368, N19359, N3520, N12734, N13375);
not NOT1 (N19369, N19364);
nand NAND4 (N19370, N19366, N12800, N13187, N10813);
and AND3 (N19371, N19362, N8704, N8956);
not NOT1 (N19372, N19357);
not NOT1 (N19373, N19367);
and AND3 (N19374, N19369, N16419, N330);
xor XOR2 (N19375, N19365, N13966);
and AND2 (N19376, N19373, N846);
nand NAND4 (N19377, N19372, N9438, N4553, N9578);
and AND2 (N19378, N19368, N6949);
and AND2 (N19379, N19374, N4441);
nor NOR2 (N19380, N19360, N7770);
nand NAND4 (N19381, N19358, N10725, N13773, N8332);
xor XOR2 (N19382, N19379, N3521);
buf BUF1 (N19383, N19370);
xor XOR2 (N19384, N19377, N15370);
nand NAND2 (N19385, N19375, N16083);
or OR3 (N19386, N19378, N10, N14924);
nor NOR2 (N19387, N19386, N1080);
nand NAND3 (N19388, N19384, N17181, N11992);
nand NAND4 (N19389, N19388, N17023, N611, N3668);
and AND4 (N19390, N19376, N2550, N4391, N3484);
and AND3 (N19391, N19389, N4914, N16674);
buf BUF1 (N19392, N19353);
nand NAND4 (N19393, N19391, N6803, N8114, N13430);
nor NOR2 (N19394, N19383, N3417);
or OR2 (N19395, N19392, N5608);
xor XOR2 (N19396, N19385, N13530);
and AND3 (N19397, N19394, N15366, N11308);
xor XOR2 (N19398, N19395, N8932);
buf BUF1 (N19399, N19381);
buf BUF1 (N19400, N19380);
or OR2 (N19401, N19371, N19154);
nor NOR3 (N19402, N19387, N11395, N15096);
nand NAND2 (N19403, N19400, N11174);
or OR2 (N19404, N19382, N18222);
nor NOR3 (N19405, N19401, N12462, N13127);
and AND4 (N19406, N19390, N11192, N14866, N4210);
nor NOR2 (N19407, N19405, N18460);
xor XOR2 (N19408, N19407, N4658);
nand NAND3 (N19409, N19403, N9395, N7153);
nor NOR4 (N19410, N19398, N18707, N16732, N8768);
not NOT1 (N19411, N19406);
xor XOR2 (N19412, N19411, N11197);
and AND4 (N19413, N19399, N7434, N8320, N18749);
nand NAND2 (N19414, N19408, N18071);
and AND2 (N19415, N19397, N767);
and AND4 (N19416, N19412, N18175, N11918, N1501);
nand NAND3 (N19417, N19415, N5609, N1828);
nand NAND3 (N19418, N19417, N17039, N3395);
or OR2 (N19419, N19410, N8590);
and AND2 (N19420, N19396, N15205);
nand NAND2 (N19421, N19419, N9622);
nand NAND3 (N19422, N19414, N10082, N14734);
or OR4 (N19423, N19404, N2668, N286, N3271);
and AND3 (N19424, N19423, N14244, N926);
buf BUF1 (N19425, N19393);
nor NOR3 (N19426, N19413, N14167, N16875);
xor XOR2 (N19427, N19409, N4880);
nand NAND4 (N19428, N19427, N10889, N17013, N18764);
or OR2 (N19429, N19418, N8361);
and AND3 (N19430, N19424, N2185, N4111);
buf BUF1 (N19431, N19425);
or OR3 (N19432, N19420, N6987, N2356);
xor XOR2 (N19433, N19422, N17630);
and AND2 (N19434, N19432, N1546);
buf BUF1 (N19435, N19433);
or OR4 (N19436, N19429, N14110, N16677, N1584);
buf BUF1 (N19437, N19428);
or OR3 (N19438, N19421, N937, N3953);
xor XOR2 (N19439, N19430, N6338);
nand NAND4 (N19440, N19438, N13711, N2003, N10471);
buf BUF1 (N19441, N19402);
xor XOR2 (N19442, N19439, N14291);
or OR3 (N19443, N19435, N4005, N11535);
nand NAND3 (N19444, N19437, N5066, N2422);
and AND4 (N19445, N19434, N10710, N1445, N10305);
nor NOR3 (N19446, N19416, N3620, N18063);
and AND4 (N19447, N19445, N1480, N1879, N17013);
buf BUF1 (N19448, N19436);
nand NAND2 (N19449, N19426, N12756);
buf BUF1 (N19450, N19443);
nand NAND3 (N19451, N19444, N15989, N11660);
or OR4 (N19452, N19431, N814, N10085, N14809);
nand NAND3 (N19453, N19446, N2796, N5188);
buf BUF1 (N19454, N19451);
nand NAND4 (N19455, N19440, N7445, N2756, N6160);
and AND4 (N19456, N19441, N13627, N17030, N13722);
nand NAND3 (N19457, N19442, N9536, N4699);
nor NOR2 (N19458, N19450, N19007);
buf BUF1 (N19459, N19455);
and AND4 (N19460, N19459, N13481, N8330, N3642);
nor NOR4 (N19461, N19448, N8546, N11231, N4353);
buf BUF1 (N19462, N19452);
nor NOR2 (N19463, N19462, N12758);
or OR2 (N19464, N19449, N4780);
not NOT1 (N19465, N19461);
buf BUF1 (N19466, N19460);
buf BUF1 (N19467, N19463);
not NOT1 (N19468, N19453);
and AND2 (N19469, N19447, N15147);
nor NOR4 (N19470, N19454, N10859, N5578, N4494);
nor NOR2 (N19471, N19465, N7683);
nand NAND3 (N19472, N19456, N2978, N16135);
or OR2 (N19473, N19464, N15555);
buf BUF1 (N19474, N19458);
nand NAND3 (N19475, N19467, N15334, N929);
or OR4 (N19476, N19471, N12331, N3800, N18871);
and AND2 (N19477, N19457, N17031);
not NOT1 (N19478, N19472);
buf BUF1 (N19479, N19473);
or OR4 (N19480, N19475, N5121, N9111, N2049);
not NOT1 (N19481, N19479);
xor XOR2 (N19482, N19478, N693);
nor NOR4 (N19483, N19476, N11318, N18332, N169);
or OR2 (N19484, N19480, N17543);
nor NOR3 (N19485, N19468, N173, N4916);
and AND4 (N19486, N19485, N4386, N6718, N384);
buf BUF1 (N19487, N19477);
and AND2 (N19488, N19474, N14287);
buf BUF1 (N19489, N19488);
xor XOR2 (N19490, N19489, N16740);
nor NOR3 (N19491, N19470, N11469, N6396);
buf BUF1 (N19492, N19487);
or OR4 (N19493, N19484, N1531, N12372, N11395);
buf BUF1 (N19494, N19492);
nor NOR2 (N19495, N19491, N6641);
not NOT1 (N19496, N19466);
and AND3 (N19497, N19481, N6493, N16502);
xor XOR2 (N19498, N19490, N4819);
and AND2 (N19499, N19486, N17861);
nand NAND3 (N19500, N19499, N1631, N14145);
not NOT1 (N19501, N19483);
and AND3 (N19502, N19498, N11564, N13051);
and AND2 (N19503, N19493, N6955);
nand NAND2 (N19504, N19494, N3325);
not NOT1 (N19505, N19482);
xor XOR2 (N19506, N19502, N18998);
nor NOR2 (N19507, N19503, N17349);
buf BUF1 (N19508, N19507);
nor NOR3 (N19509, N19469, N637, N1983);
or OR4 (N19510, N19496, N18976, N12620, N5137);
xor XOR2 (N19511, N19510, N19172);
nand NAND3 (N19512, N19508, N7260, N4503);
nand NAND4 (N19513, N19501, N10838, N13557, N9546);
nand NAND3 (N19514, N19504, N12925, N17457);
and AND2 (N19515, N19495, N337);
nand NAND3 (N19516, N19512, N1924, N14680);
nand NAND4 (N19517, N19500, N10428, N4633, N17775);
and AND3 (N19518, N19514, N2852, N13913);
xor XOR2 (N19519, N19509, N141);
xor XOR2 (N19520, N19518, N3304);
or OR3 (N19521, N19511, N15837, N11238);
xor XOR2 (N19522, N19520, N2630);
and AND3 (N19523, N19515, N16828, N12715);
and AND4 (N19524, N19517, N9923, N15083, N16632);
not NOT1 (N19525, N19505);
and AND2 (N19526, N19523, N18580);
xor XOR2 (N19527, N19516, N4953);
not NOT1 (N19528, N19513);
or OR3 (N19529, N19506, N7672, N5903);
not NOT1 (N19530, N19526);
nor NOR3 (N19531, N19529, N15959, N17430);
not NOT1 (N19532, N19530);
nor NOR3 (N19533, N19531, N1134, N10186);
and AND3 (N19534, N19528, N8051, N7152);
and AND4 (N19535, N19527, N17620, N15788, N13505);
nor NOR2 (N19536, N19532, N875);
or OR3 (N19537, N19521, N8460, N7963);
nand NAND3 (N19538, N19522, N10840, N16242);
nor NOR4 (N19539, N19537, N12163, N19502, N3330);
not NOT1 (N19540, N19525);
and AND4 (N19541, N19540, N9722, N15226, N13326);
or OR3 (N19542, N19538, N17395, N4374);
not NOT1 (N19543, N19519);
not NOT1 (N19544, N19536);
nor NOR3 (N19545, N19542, N1217, N19133);
or OR3 (N19546, N19524, N6255, N18609);
nor NOR4 (N19547, N19544, N8696, N4397, N4506);
nand NAND2 (N19548, N19545, N3807);
xor XOR2 (N19549, N19539, N14927);
buf BUF1 (N19550, N19549);
xor XOR2 (N19551, N19546, N2649);
nor NOR3 (N19552, N19497, N12527, N3840);
and AND3 (N19553, N19533, N1680, N12532);
nor NOR2 (N19554, N19551, N8915);
and AND2 (N19555, N19543, N683);
buf BUF1 (N19556, N19550);
not NOT1 (N19557, N19535);
nand NAND3 (N19558, N19552, N8687, N17800);
or OR2 (N19559, N19554, N11389);
buf BUF1 (N19560, N19547);
xor XOR2 (N19561, N19558, N9454);
nand NAND4 (N19562, N19556, N5157, N13411, N11973);
and AND3 (N19563, N19553, N17755, N14697);
buf BUF1 (N19564, N19559);
nor NOR3 (N19565, N19561, N16955, N16541);
and AND3 (N19566, N19557, N12219, N11276);
and AND4 (N19567, N19564, N16119, N10478, N8319);
nor NOR3 (N19568, N19555, N17382, N12872);
buf BUF1 (N19569, N19565);
nand NAND2 (N19570, N19534, N1846);
nand NAND2 (N19571, N19568, N2632);
and AND3 (N19572, N19562, N5284, N2937);
xor XOR2 (N19573, N19560, N3483);
buf BUF1 (N19574, N19572);
or OR4 (N19575, N19569, N3534, N14605, N19144);
not NOT1 (N19576, N19573);
buf BUF1 (N19577, N19548);
and AND4 (N19578, N19576, N2714, N12214, N4419);
nor NOR2 (N19579, N19577, N13403);
or OR3 (N19580, N19579, N3249, N998);
and AND3 (N19581, N19541, N16349, N16997);
xor XOR2 (N19582, N19575, N373);
or OR4 (N19583, N19574, N2059, N1262, N15583);
nor NOR4 (N19584, N19582, N15004, N13850, N18106);
xor XOR2 (N19585, N19578, N13038);
nand NAND2 (N19586, N19583, N12304);
or OR4 (N19587, N19570, N2057, N13438, N6224);
buf BUF1 (N19588, N19567);
and AND3 (N19589, N19586, N13664, N13217);
nand NAND4 (N19590, N19571, N12238, N676, N5802);
xor XOR2 (N19591, N19580, N5589);
not NOT1 (N19592, N19581);
and AND2 (N19593, N19589, N12348);
not NOT1 (N19594, N19588);
nand NAND2 (N19595, N19590, N16204);
not NOT1 (N19596, N19563);
nand NAND3 (N19597, N19593, N14446, N6295);
nand NAND2 (N19598, N19595, N18685);
buf BUF1 (N19599, N19587);
and AND4 (N19600, N19591, N9044, N6663, N13274);
nand NAND4 (N19601, N19585, N5837, N16234, N11439);
buf BUF1 (N19602, N19596);
nand NAND4 (N19603, N19599, N4905, N6234, N19586);
nand NAND3 (N19604, N19592, N4898, N17370);
buf BUF1 (N19605, N19601);
or OR3 (N19606, N19600, N1729, N10226);
nor NOR4 (N19607, N19602, N2351, N1519, N8490);
not NOT1 (N19608, N19598);
and AND4 (N19609, N19597, N6056, N13713, N13810);
xor XOR2 (N19610, N19584, N14369);
not NOT1 (N19611, N19608);
nor NOR2 (N19612, N19607, N1338);
or OR3 (N19613, N19604, N17803, N2822);
and AND4 (N19614, N19613, N4303, N2149, N14428);
xor XOR2 (N19615, N19614, N17153);
or OR3 (N19616, N19603, N12342, N14730);
and AND2 (N19617, N19606, N6921);
and AND2 (N19618, N19617, N4677);
nand NAND4 (N19619, N19615, N17008, N16406, N10023);
nand NAND3 (N19620, N19616, N6295, N1914);
or OR2 (N19621, N19612, N3618);
nand NAND2 (N19622, N19620, N13855);
or OR3 (N19623, N19610, N6991, N6511);
nor NOR2 (N19624, N19609, N9395);
buf BUF1 (N19625, N19611);
xor XOR2 (N19626, N19621, N15780);
nor NOR2 (N19627, N19624, N11914);
nor NOR4 (N19628, N19605, N10619, N18056, N11122);
buf BUF1 (N19629, N19618);
nor NOR2 (N19630, N19566, N13379);
nand NAND2 (N19631, N19628, N18684);
not NOT1 (N19632, N19626);
buf BUF1 (N19633, N19623);
or OR2 (N19634, N19632, N11375);
nand NAND3 (N19635, N19594, N744, N16355);
nor NOR2 (N19636, N19629, N8402);
buf BUF1 (N19637, N19636);
not NOT1 (N19638, N19631);
nand NAND3 (N19639, N19622, N18697, N15518);
buf BUF1 (N19640, N19627);
not NOT1 (N19641, N19633);
xor XOR2 (N19642, N19639, N4687);
or OR3 (N19643, N19638, N13914, N13932);
or OR3 (N19644, N19625, N11119, N11165);
nand NAND4 (N19645, N19640, N9280, N3611, N2404);
buf BUF1 (N19646, N19644);
nand NAND4 (N19647, N19642, N13279, N5969, N717);
xor XOR2 (N19648, N19646, N8632);
or OR2 (N19649, N19637, N7924);
nor NOR2 (N19650, N19648, N1697);
and AND2 (N19651, N19619, N6592);
or OR4 (N19652, N19643, N5911, N3926, N2855);
buf BUF1 (N19653, N19649);
not NOT1 (N19654, N19652);
and AND4 (N19655, N19650, N17373, N6441, N10002);
buf BUF1 (N19656, N19651);
nand NAND4 (N19657, N19635, N10148, N2025, N8095);
or OR4 (N19658, N19656, N19064, N12578, N12283);
nand NAND2 (N19659, N19655, N12851);
and AND4 (N19660, N19647, N9623, N16734, N10493);
and AND3 (N19661, N19653, N305, N17322);
xor XOR2 (N19662, N19661, N8863);
nor NOR2 (N19663, N19658, N18162);
or OR2 (N19664, N19645, N3045);
nand NAND4 (N19665, N19659, N9268, N1302, N5016);
buf BUF1 (N19666, N19665);
not NOT1 (N19667, N19663);
xor XOR2 (N19668, N19630, N17068);
nor NOR3 (N19669, N19654, N17939, N2007);
or OR2 (N19670, N19634, N16428);
nor NOR4 (N19671, N19670, N18904, N11528, N185);
xor XOR2 (N19672, N19657, N19499);
or OR2 (N19673, N19668, N9748);
not NOT1 (N19674, N19672);
or OR2 (N19675, N19641, N12745);
buf BUF1 (N19676, N19666);
nand NAND4 (N19677, N19674, N475, N18583, N5610);
not NOT1 (N19678, N19667);
xor XOR2 (N19679, N19676, N15374);
nor NOR3 (N19680, N19677, N8831, N1309);
nor NOR2 (N19681, N19680, N9813);
nor NOR2 (N19682, N19678, N19551);
or OR3 (N19683, N19669, N8055, N17150);
and AND4 (N19684, N19664, N1776, N5306, N2163);
and AND2 (N19685, N19660, N17796);
nor NOR2 (N19686, N19673, N13166);
nor NOR4 (N19687, N19671, N105, N866, N19106);
xor XOR2 (N19688, N19684, N8434);
not NOT1 (N19689, N19686);
buf BUF1 (N19690, N19681);
not NOT1 (N19691, N19688);
xor XOR2 (N19692, N19689, N2449);
or OR2 (N19693, N19662, N10321);
nor NOR3 (N19694, N19692, N818, N19032);
or OR2 (N19695, N19693, N14173);
and AND2 (N19696, N19687, N536);
or OR4 (N19697, N19683, N2044, N7897, N19464);
or OR3 (N19698, N19697, N8888, N6228);
nand NAND3 (N19699, N19694, N17298, N263);
or OR4 (N19700, N19695, N3987, N13525, N12191);
xor XOR2 (N19701, N19682, N8465);
or OR4 (N19702, N19675, N14995, N2562, N12495);
nand NAND3 (N19703, N19685, N4110, N9612);
buf BUF1 (N19704, N19679);
or OR2 (N19705, N19691, N3793);
or OR2 (N19706, N19705, N10441);
nor NOR4 (N19707, N19698, N6268, N6516, N4549);
buf BUF1 (N19708, N19699);
nand NAND3 (N19709, N19704, N6944, N19);
and AND3 (N19710, N19703, N3558, N4705);
or OR3 (N19711, N19701, N19481, N15965);
nor NOR3 (N19712, N19708, N8124, N274);
and AND3 (N19713, N19709, N16201, N7648);
and AND2 (N19714, N19690, N7391);
or OR3 (N19715, N19700, N18202, N2086);
buf BUF1 (N19716, N19707);
nand NAND3 (N19717, N19711, N6593, N16174);
and AND3 (N19718, N19712, N862, N9840);
and AND2 (N19719, N19706, N3620);
and AND2 (N19720, N19719, N18901);
nand NAND2 (N19721, N19714, N10802);
not NOT1 (N19722, N19717);
buf BUF1 (N19723, N19720);
and AND3 (N19724, N19696, N8085, N16532);
nor NOR3 (N19725, N19713, N9351, N2726);
and AND4 (N19726, N19715, N16648, N7527, N5800);
nor NOR3 (N19727, N19718, N5555, N1196);
or OR4 (N19728, N19725, N13225, N9055, N11351);
buf BUF1 (N19729, N19710);
or OR2 (N19730, N19721, N8813);
nor NOR3 (N19731, N19728, N18451, N6527);
buf BUF1 (N19732, N19724);
or OR3 (N19733, N19730, N16179, N5616);
nor NOR3 (N19734, N19732, N10587, N10109);
not NOT1 (N19735, N19702);
xor XOR2 (N19736, N19726, N18274);
nor NOR3 (N19737, N19731, N1800, N11743);
buf BUF1 (N19738, N19734);
xor XOR2 (N19739, N19733, N13505);
and AND3 (N19740, N19737, N10290, N5913);
and AND4 (N19741, N19736, N709, N15480, N2895);
buf BUF1 (N19742, N19727);
or OR2 (N19743, N19741, N8753);
nand NAND3 (N19744, N19743, N18501, N10125);
xor XOR2 (N19745, N19722, N13212);
nand NAND4 (N19746, N19738, N9974, N18119, N5616);
and AND2 (N19747, N19716, N11640);
or OR3 (N19748, N19744, N15377, N18714);
or OR4 (N19749, N19748, N8363, N14863, N14955);
xor XOR2 (N19750, N19742, N11357);
buf BUF1 (N19751, N19747);
xor XOR2 (N19752, N19729, N11912);
nor NOR3 (N19753, N19751, N4111, N4286);
buf BUF1 (N19754, N19750);
nand NAND2 (N19755, N19754, N8787);
nor NOR3 (N19756, N19755, N16482, N3944);
not NOT1 (N19757, N19749);
not NOT1 (N19758, N19723);
nor NOR4 (N19759, N19752, N16745, N8885, N5608);
nor NOR3 (N19760, N19740, N18335, N11866);
xor XOR2 (N19761, N19739, N13575);
nand NAND4 (N19762, N19758, N8957, N6055, N976);
and AND2 (N19763, N19759, N2733);
or OR2 (N19764, N19760, N3702);
nand NAND3 (N19765, N19763, N2254, N18800);
xor XOR2 (N19766, N19756, N6363);
or OR3 (N19767, N19746, N11544, N9229);
and AND4 (N19768, N19767, N14402, N4634, N17204);
buf BUF1 (N19769, N19753);
or OR4 (N19770, N19757, N11293, N7303, N15572);
not NOT1 (N19771, N19769);
nor NOR2 (N19772, N19768, N11577);
or OR3 (N19773, N19762, N18414, N4890);
xor XOR2 (N19774, N19770, N5836);
and AND2 (N19775, N19764, N9561);
xor XOR2 (N19776, N19772, N5498);
buf BUF1 (N19777, N19773);
nand NAND3 (N19778, N19774, N19524, N900);
buf BUF1 (N19779, N19765);
and AND3 (N19780, N19776, N11017, N5955);
and AND2 (N19781, N19735, N17910);
or OR4 (N19782, N19780, N13512, N5427, N7619);
nand NAND2 (N19783, N19782, N7709);
nand NAND2 (N19784, N19783, N13797);
nor NOR3 (N19785, N19775, N14946, N9447);
buf BUF1 (N19786, N19785);
not NOT1 (N19787, N19781);
not NOT1 (N19788, N19761);
or OR4 (N19789, N19777, N8636, N917, N4355);
buf BUF1 (N19790, N19771);
and AND3 (N19791, N19745, N14121, N12615);
nor NOR4 (N19792, N19766, N5184, N19253, N15639);
or OR4 (N19793, N19789, N9872, N137, N5303);
not NOT1 (N19794, N19788);
nor NOR4 (N19795, N19787, N11994, N16491, N15949);
and AND2 (N19796, N19795, N1648);
buf BUF1 (N19797, N19794);
and AND4 (N19798, N19791, N14655, N14552, N18367);
nand NAND3 (N19799, N19786, N1883, N1935);
and AND3 (N19800, N19793, N2649, N7129);
nand NAND4 (N19801, N19790, N15948, N1657, N12338);
xor XOR2 (N19802, N19778, N9751);
buf BUF1 (N19803, N19797);
nor NOR3 (N19804, N19779, N8641, N4104);
not NOT1 (N19805, N19800);
xor XOR2 (N19806, N19804, N1083);
nor NOR2 (N19807, N19796, N7608);
xor XOR2 (N19808, N19801, N12693);
nand NAND2 (N19809, N19807, N267);
nand NAND4 (N19810, N19806, N1295, N14191, N13643);
not NOT1 (N19811, N19798);
nor NOR4 (N19812, N19799, N3243, N18235, N8587);
buf BUF1 (N19813, N19805);
nor NOR2 (N19814, N19803, N13603);
buf BUF1 (N19815, N19812);
nand NAND4 (N19816, N19792, N5456, N14536, N17133);
buf BUF1 (N19817, N19811);
not NOT1 (N19818, N19784);
and AND2 (N19819, N19814, N16244);
or OR4 (N19820, N19819, N8057, N9014, N6795);
or OR2 (N19821, N19808, N18929);
not NOT1 (N19822, N19815);
not NOT1 (N19823, N19817);
nor NOR3 (N19824, N19802, N11666, N6566);
not NOT1 (N19825, N19821);
and AND4 (N19826, N19824, N17179, N10688, N12968);
nor NOR3 (N19827, N19826, N18089, N11456);
xor XOR2 (N19828, N19825, N9661);
xor XOR2 (N19829, N19813, N8031);
nor NOR4 (N19830, N19816, N2101, N945, N11443);
nand NAND3 (N19831, N19809, N2614, N11859);
nand NAND4 (N19832, N19828, N15881, N16770, N9798);
nor NOR4 (N19833, N19818, N10829, N18180, N8645);
xor XOR2 (N19834, N19827, N15196);
or OR2 (N19835, N19832, N10388);
not NOT1 (N19836, N19822);
xor XOR2 (N19837, N19833, N16178);
xor XOR2 (N19838, N19835, N6830);
and AND4 (N19839, N19810, N4297, N4685, N15051);
not NOT1 (N19840, N19829);
nor NOR2 (N19841, N19836, N8572);
not NOT1 (N19842, N19840);
nand NAND3 (N19843, N19830, N3798, N12119);
buf BUF1 (N19844, N19831);
not NOT1 (N19845, N19843);
nand NAND2 (N19846, N19837, N4729);
xor XOR2 (N19847, N19823, N8683);
not NOT1 (N19848, N19844);
not NOT1 (N19849, N19838);
or OR2 (N19850, N19839, N10879);
not NOT1 (N19851, N19834);
buf BUF1 (N19852, N19846);
or OR4 (N19853, N19851, N13055, N16197, N13508);
buf BUF1 (N19854, N19849);
xor XOR2 (N19855, N19847, N18342);
not NOT1 (N19856, N19852);
xor XOR2 (N19857, N19856, N6850);
not NOT1 (N19858, N19850);
not NOT1 (N19859, N19842);
nor NOR2 (N19860, N19854, N17555);
nand NAND4 (N19861, N19860, N3994, N17188, N14565);
and AND3 (N19862, N19841, N12146, N6004);
not NOT1 (N19863, N19820);
buf BUF1 (N19864, N19855);
or OR3 (N19865, N19857, N17891, N14178);
xor XOR2 (N19866, N19865, N3833);
not NOT1 (N19867, N19864);
and AND2 (N19868, N19867, N13314);
xor XOR2 (N19869, N19862, N12934);
xor XOR2 (N19870, N19848, N12854);
nand NAND4 (N19871, N19868, N3516, N5064, N7585);
nand NAND2 (N19872, N19870, N19541);
xor XOR2 (N19873, N19845, N5371);
nand NAND4 (N19874, N19871, N14048, N18313, N6839);
nor NOR4 (N19875, N19866, N12093, N1760, N15757);
xor XOR2 (N19876, N19859, N16037);
nand NAND2 (N19877, N19872, N4477);
xor XOR2 (N19878, N19877, N4459);
not NOT1 (N19879, N19861);
not NOT1 (N19880, N19858);
or OR2 (N19881, N19875, N1967);
and AND4 (N19882, N19879, N10788, N1125, N7010);
and AND4 (N19883, N19882, N10679, N19283, N9350);
not NOT1 (N19884, N19863);
buf BUF1 (N19885, N19878);
nand NAND4 (N19886, N19869, N15694, N8278, N15614);
not NOT1 (N19887, N19884);
or OR4 (N19888, N19887, N8676, N9478, N1074);
nand NAND2 (N19889, N19853, N12023);
and AND3 (N19890, N19880, N17226, N8857);
not NOT1 (N19891, N19873);
nor NOR2 (N19892, N19885, N14312);
buf BUF1 (N19893, N19892);
nor NOR4 (N19894, N19888, N2491, N3826, N1442);
nand NAND2 (N19895, N19890, N12553);
buf BUF1 (N19896, N19881);
nor NOR4 (N19897, N19896, N10407, N5290, N5295);
and AND4 (N19898, N19883, N7790, N5393, N14966);
buf BUF1 (N19899, N19876);
and AND3 (N19900, N19895, N1252, N15997);
buf BUF1 (N19901, N19891);
nand NAND3 (N19902, N19874, N10239, N9194);
buf BUF1 (N19903, N19893);
and AND2 (N19904, N19899, N228);
nand NAND3 (N19905, N19897, N5274, N14871);
or OR4 (N19906, N19894, N14940, N3236, N3775);
and AND3 (N19907, N19902, N8062, N8906);
xor XOR2 (N19908, N19906, N3342);
xor XOR2 (N19909, N19901, N1493);
or OR3 (N19910, N19898, N6373, N15167);
buf BUF1 (N19911, N19886);
not NOT1 (N19912, N19909);
xor XOR2 (N19913, N19904, N14840);
nor NOR4 (N19914, N19908, N16166, N14190, N7432);
nand NAND4 (N19915, N19900, N9180, N14588, N9920);
nor NOR2 (N19916, N19912, N8893);
nand NAND2 (N19917, N19905, N7605);
and AND4 (N19918, N19913, N11061, N12510, N7852);
nand NAND4 (N19919, N19915, N9602, N18774, N18742);
nand NAND3 (N19920, N19911, N11216, N18169);
buf BUF1 (N19921, N19889);
not NOT1 (N19922, N19917);
xor XOR2 (N19923, N19907, N9693);
buf BUF1 (N19924, N19916);
nand NAND4 (N19925, N19903, N12595, N154, N19523);
or OR2 (N19926, N19925, N11334);
and AND3 (N19927, N19919, N8166, N16334);
not NOT1 (N19928, N19922);
or OR3 (N19929, N19923, N19443, N15529);
not NOT1 (N19930, N19927);
nand NAND2 (N19931, N19921, N9616);
not NOT1 (N19932, N19918);
buf BUF1 (N19933, N19931);
nand NAND3 (N19934, N19926, N17707, N7084);
or OR4 (N19935, N19933, N4233, N17229, N10763);
and AND2 (N19936, N19920, N4750);
not NOT1 (N19937, N19924);
buf BUF1 (N19938, N19928);
not NOT1 (N19939, N19935);
nand NAND2 (N19940, N19939, N11373);
nand NAND4 (N19941, N19930, N799, N6301, N15991);
not NOT1 (N19942, N19938);
not NOT1 (N19943, N19941);
or OR3 (N19944, N19937, N16847, N3357);
and AND3 (N19945, N19910, N18223, N1311);
or OR2 (N19946, N19929, N7273);
buf BUF1 (N19947, N19945);
buf BUF1 (N19948, N19944);
nand NAND2 (N19949, N19946, N14046);
not NOT1 (N19950, N19942);
not NOT1 (N19951, N19932);
or OR4 (N19952, N19950, N18613, N5816, N12528);
nand NAND4 (N19953, N19934, N18351, N12635, N7964);
or OR2 (N19954, N19943, N6444);
xor XOR2 (N19955, N19936, N15614);
xor XOR2 (N19956, N19954, N9005);
or OR4 (N19957, N19952, N17350, N19820, N724);
or OR4 (N19958, N19956, N1512, N139, N2341);
xor XOR2 (N19959, N19947, N12822);
nand NAND3 (N19960, N19948, N19306, N8758);
not NOT1 (N19961, N19960);
and AND2 (N19962, N19940, N14106);
xor XOR2 (N19963, N19961, N2108);
buf BUF1 (N19964, N19959);
not NOT1 (N19965, N19957);
nand NAND2 (N19966, N19951, N3888);
buf BUF1 (N19967, N19962);
nand NAND2 (N19968, N19958, N14844);
xor XOR2 (N19969, N19964, N479);
nand NAND2 (N19970, N19968, N18699);
nor NOR3 (N19971, N19914, N16817, N12679);
buf BUF1 (N19972, N19949);
nand NAND3 (N19973, N19971, N5192, N6570);
or OR2 (N19974, N19972, N2352);
buf BUF1 (N19975, N19953);
nand NAND2 (N19976, N19975, N17394);
nand NAND4 (N19977, N19965, N603, N6932, N1851);
and AND3 (N19978, N19969, N1789, N14856);
or OR2 (N19979, N19967, N18231);
xor XOR2 (N19980, N19955, N13689);
xor XOR2 (N19981, N19966, N10573);
not NOT1 (N19982, N19980);
or OR2 (N19983, N19977, N19079);
or OR2 (N19984, N19978, N19144);
xor XOR2 (N19985, N19976, N10919);
nand NAND2 (N19986, N19985, N17346);
nand NAND4 (N19987, N19979, N19351, N15591, N12660);
nor NOR3 (N19988, N19970, N7612, N18389);
nand NAND3 (N19989, N19987, N8826, N3165);
not NOT1 (N19990, N19973);
not NOT1 (N19991, N19990);
buf BUF1 (N19992, N19982);
or OR3 (N19993, N19989, N8457, N5147);
buf BUF1 (N19994, N19993);
or OR2 (N19995, N19983, N586);
nand NAND3 (N19996, N19974, N16694, N18293);
not NOT1 (N19997, N19992);
not NOT1 (N19998, N19981);
nand NAND3 (N19999, N19996, N17793, N8403);
xor XOR2 (N20000, N19999, N10981);
nand NAND2 (N20001, N19995, N2943);
xor XOR2 (N20002, N19984, N2873);
nand NAND4 (N20003, N20002, N11078, N12019, N8498);
or OR4 (N20004, N19991, N19918, N17210, N15112);
not NOT1 (N20005, N20003);
and AND2 (N20006, N20005, N10565);
or OR4 (N20007, N19986, N12266, N8199, N17270);
and AND4 (N20008, N19997, N8862, N14006, N18869);
not NOT1 (N20009, N19998);
nor NOR3 (N20010, N19988, N7997, N8633);
not NOT1 (N20011, N20004);
nand NAND4 (N20012, N20000, N13861, N14380, N17237);
nand NAND2 (N20013, N20009, N15036);
and AND2 (N20014, N20010, N15421);
xor XOR2 (N20015, N20001, N13379);
xor XOR2 (N20016, N20015, N3686);
xor XOR2 (N20017, N20013, N9780);
or OR3 (N20018, N20016, N13142, N3429);
or OR3 (N20019, N20012, N8481, N11508);
xor XOR2 (N20020, N20017, N14459);
xor XOR2 (N20021, N19994, N14746);
and AND2 (N20022, N20011, N16091);
not NOT1 (N20023, N20014);
buf BUF1 (N20024, N20019);
not NOT1 (N20025, N20021);
not NOT1 (N20026, N20020);
xor XOR2 (N20027, N19963, N8473);
and AND2 (N20028, N20026, N5121);
not NOT1 (N20029, N20018);
buf BUF1 (N20030, N20024);
nor NOR4 (N20031, N20029, N5840, N8242, N6991);
nand NAND4 (N20032, N20022, N16337, N5587, N15596);
or OR3 (N20033, N20031, N16472, N14940);
xor XOR2 (N20034, N20030, N3399);
xor XOR2 (N20035, N20032, N10535);
not NOT1 (N20036, N20008);
buf BUF1 (N20037, N20036);
nand NAND4 (N20038, N20025, N3783, N1531, N4074);
xor XOR2 (N20039, N20035, N10686);
buf BUF1 (N20040, N20033);
nand NAND3 (N20041, N20037, N9618, N13701);
not NOT1 (N20042, N20038);
not NOT1 (N20043, N20040);
or OR3 (N20044, N20027, N12465, N6554);
nor NOR3 (N20045, N20043, N15446, N16230);
or OR3 (N20046, N20045, N3982, N5449);
nor NOR4 (N20047, N20006, N13768, N14089, N10027);
not NOT1 (N20048, N20046);
nand NAND3 (N20049, N20034, N5418, N2495);
nand NAND2 (N20050, N20042, N18422);
buf BUF1 (N20051, N20007);
nor NOR4 (N20052, N20028, N19836, N15352, N10009);
and AND4 (N20053, N20047, N16529, N8917, N11421);
or OR2 (N20054, N20023, N1257);
xor XOR2 (N20055, N20054, N6174);
nand NAND2 (N20056, N20051, N7997);
buf BUF1 (N20057, N20048);
xor XOR2 (N20058, N20055, N2183);
nor NOR2 (N20059, N20052, N15237);
nor NOR4 (N20060, N20059, N1274, N19773, N5209);
or OR2 (N20061, N20053, N19026);
xor XOR2 (N20062, N20058, N7513);
or OR4 (N20063, N20039, N12077, N16027, N15205);
nand NAND3 (N20064, N20060, N17759, N15211);
nor NOR2 (N20065, N20063, N17311);
buf BUF1 (N20066, N20056);
nor NOR2 (N20067, N20065, N12805);
not NOT1 (N20068, N20067);
not NOT1 (N20069, N20068);
nand NAND3 (N20070, N20057, N11630, N7234);
nor NOR4 (N20071, N20066, N15530, N5633, N2536);
buf BUF1 (N20072, N20061);
nor NOR3 (N20073, N20050, N19525, N12233);
nand NAND4 (N20074, N20049, N14048, N10984, N17975);
nand NAND3 (N20075, N20041, N2128, N19517);
buf BUF1 (N20076, N20071);
nand NAND4 (N20077, N20070, N8090, N9809, N6210);
or OR3 (N20078, N20076, N8080, N3169);
not NOT1 (N20079, N20075);
xor XOR2 (N20080, N20073, N5385);
nor NOR2 (N20081, N20044, N10884);
and AND4 (N20082, N20078, N5337, N12078, N2957);
or OR4 (N20083, N20077, N13226, N3943, N15075);
not NOT1 (N20084, N20083);
or OR4 (N20085, N20072, N1855, N12565, N3601);
and AND4 (N20086, N20064, N11362, N12014, N4472);
and AND2 (N20087, N20062, N7514);
and AND2 (N20088, N20079, N17846);
xor XOR2 (N20089, N20074, N10757);
and AND4 (N20090, N20084, N7203, N5383, N14281);
nand NAND3 (N20091, N20080, N7364, N11870);
and AND2 (N20092, N20069, N6205);
nand NAND3 (N20093, N20081, N13934, N3190);
or OR2 (N20094, N20086, N6268);
or OR4 (N20095, N20092, N4672, N14621, N522);
nand NAND4 (N20096, N20087, N650, N16612, N2704);
not NOT1 (N20097, N20093);
nor NOR3 (N20098, N20082, N8429, N18394);
xor XOR2 (N20099, N20090, N2802);
xor XOR2 (N20100, N20085, N1243);
or OR4 (N20101, N20091, N7771, N15634, N4191);
nor NOR3 (N20102, N20094, N8424, N2386);
nor NOR4 (N20103, N20100, N2523, N3531, N1854);
nor NOR4 (N20104, N20097, N18824, N3392, N12816);
not NOT1 (N20105, N20101);
xor XOR2 (N20106, N20105, N15135);
nor NOR2 (N20107, N20098, N14721);
buf BUF1 (N20108, N20088);
or OR4 (N20109, N20095, N647, N13747, N16616);
xor XOR2 (N20110, N20109, N2921);
nand NAND2 (N20111, N20089, N15450);
and AND3 (N20112, N20110, N2374, N11287);
and AND4 (N20113, N20104, N17620, N10280, N11083);
not NOT1 (N20114, N20112);
or OR3 (N20115, N20113, N14058, N16919);
buf BUF1 (N20116, N20114);
nor NOR4 (N20117, N20102, N11299, N9131, N4985);
and AND4 (N20118, N20108, N19322, N3587, N17396);
nor NOR4 (N20119, N20115, N5105, N7766, N19907);
xor XOR2 (N20120, N20119, N1411);
xor XOR2 (N20121, N20118, N5180);
or OR4 (N20122, N20120, N18624, N6786, N13340);
nand NAND4 (N20123, N20096, N9538, N6174, N14208);
nor NOR2 (N20124, N20107, N17198);
and AND4 (N20125, N20106, N6309, N17708, N2978);
and AND4 (N20126, N20122, N3197, N7369, N19718);
xor XOR2 (N20127, N20126, N7972);
nor NOR2 (N20128, N20121, N19092);
nor NOR2 (N20129, N20123, N19708);
or OR2 (N20130, N20099, N14191);
nor NOR2 (N20131, N20125, N1917);
nor NOR4 (N20132, N20103, N4247, N4019, N2971);
nand NAND3 (N20133, N20111, N13340, N11247);
and AND2 (N20134, N20124, N19999);
xor XOR2 (N20135, N20130, N15632);
not NOT1 (N20136, N20134);
not NOT1 (N20137, N20135);
and AND2 (N20138, N20132, N12327);
buf BUF1 (N20139, N20117);
nand NAND2 (N20140, N20139, N14128);
or OR4 (N20141, N20138, N11040, N19941, N5007);
buf BUF1 (N20142, N20133);
and AND4 (N20143, N20140, N3305, N7576, N8407);
nand NAND2 (N20144, N20136, N14271);
or OR3 (N20145, N20142, N16787, N13359);
xor XOR2 (N20146, N20128, N3374);
not NOT1 (N20147, N20116);
or OR2 (N20148, N20127, N3940);
buf BUF1 (N20149, N20143);
or OR2 (N20150, N20149, N5700);
not NOT1 (N20151, N20150);
buf BUF1 (N20152, N20129);
and AND4 (N20153, N20146, N2036, N8961, N6446);
nor NOR4 (N20154, N20153, N8541, N7543, N18076);
and AND3 (N20155, N20131, N3825, N186);
buf BUF1 (N20156, N20148);
nand NAND4 (N20157, N20144, N18798, N442, N14995);
nand NAND2 (N20158, N20145, N12461);
and AND2 (N20159, N20151, N5029);
xor XOR2 (N20160, N20152, N18410);
xor XOR2 (N20161, N20137, N17528);
and AND4 (N20162, N20156, N1949, N15132, N680);
nor NOR2 (N20163, N20154, N190);
xor XOR2 (N20164, N20147, N7692);
buf BUF1 (N20165, N20162);
xor XOR2 (N20166, N20155, N6367);
xor XOR2 (N20167, N20160, N560);
or OR4 (N20168, N20165, N8404, N13319, N13800);
not NOT1 (N20169, N20164);
xor XOR2 (N20170, N20163, N3154);
or OR2 (N20171, N20158, N14585);
not NOT1 (N20172, N20171);
not NOT1 (N20173, N20166);
and AND2 (N20174, N20141, N13519);
not NOT1 (N20175, N20169);
not NOT1 (N20176, N20174);
or OR3 (N20177, N20173, N18781, N1781);
or OR4 (N20178, N20167, N15743, N4357, N12455);
xor XOR2 (N20179, N20177, N153);
buf BUF1 (N20180, N20178);
not NOT1 (N20181, N20179);
and AND4 (N20182, N20175, N9673, N11934, N796);
nor NOR4 (N20183, N20161, N2466, N9627, N5615);
nor NOR2 (N20184, N20157, N14830);
nor NOR3 (N20185, N20183, N16191, N9860);
nor NOR2 (N20186, N20180, N1426);
and AND2 (N20187, N20181, N19645);
xor XOR2 (N20188, N20182, N15332);
xor XOR2 (N20189, N20185, N15203);
nand NAND3 (N20190, N20188, N11000, N3825);
not NOT1 (N20191, N20172);
not NOT1 (N20192, N20168);
or OR2 (N20193, N20186, N1728);
not NOT1 (N20194, N20184);
not NOT1 (N20195, N20194);
nor NOR2 (N20196, N20187, N16170);
buf BUF1 (N20197, N20159);
nand NAND3 (N20198, N20176, N19129, N153);
or OR2 (N20199, N20170, N19157);
and AND2 (N20200, N20196, N690);
buf BUF1 (N20201, N20197);
nor NOR4 (N20202, N20191, N6424, N10847, N17183);
and AND2 (N20203, N20200, N6794);
buf BUF1 (N20204, N20199);
not NOT1 (N20205, N20202);
nor NOR4 (N20206, N20192, N7747, N18690, N2530);
buf BUF1 (N20207, N20190);
and AND4 (N20208, N20189, N3001, N7091, N15788);
nor NOR3 (N20209, N20198, N19129, N3494);
and AND3 (N20210, N20203, N18384, N6941);
not NOT1 (N20211, N20210);
buf BUF1 (N20212, N20204);
buf BUF1 (N20213, N20205);
nand NAND2 (N20214, N20201, N1861);
buf BUF1 (N20215, N20211);
nor NOR3 (N20216, N20206, N2615, N978);
nor NOR2 (N20217, N20215, N13183);
buf BUF1 (N20218, N20214);
nor NOR2 (N20219, N20209, N14546);
buf BUF1 (N20220, N20195);
xor XOR2 (N20221, N20207, N15087);
xor XOR2 (N20222, N20213, N1118);
nand NAND4 (N20223, N20218, N983, N13421, N16215);
not NOT1 (N20224, N20221);
and AND2 (N20225, N20224, N6009);
nand NAND3 (N20226, N20217, N17921, N11148);
and AND4 (N20227, N20219, N17847, N12377, N12216);
not NOT1 (N20228, N20212);
not NOT1 (N20229, N20225);
or OR4 (N20230, N20216, N12834, N9473, N17788);
buf BUF1 (N20231, N20222);
not NOT1 (N20232, N20220);
not NOT1 (N20233, N20223);
xor XOR2 (N20234, N20227, N2508);
and AND3 (N20235, N20230, N1590, N17496);
or OR2 (N20236, N20193, N16310);
not NOT1 (N20237, N20231);
or OR3 (N20238, N20234, N12676, N1096);
nor NOR3 (N20239, N20228, N4866, N2984);
or OR4 (N20240, N20238, N5957, N3242, N15340);
nor NOR3 (N20241, N20235, N15690, N11928);
nand NAND3 (N20242, N20233, N294, N6620);
or OR2 (N20243, N20208, N10628);
or OR4 (N20244, N20237, N7010, N4657, N6276);
buf BUF1 (N20245, N20236);
buf BUF1 (N20246, N20239);
nand NAND3 (N20247, N20245, N2673, N883);
or OR4 (N20248, N20243, N1955, N15247, N17381);
buf BUF1 (N20249, N20246);
nor NOR2 (N20250, N20229, N11479);
buf BUF1 (N20251, N20241);
xor XOR2 (N20252, N20248, N7307);
not NOT1 (N20253, N20240);
xor XOR2 (N20254, N20249, N6510);
or OR2 (N20255, N20251, N4995);
nand NAND3 (N20256, N20226, N1100, N17799);
buf BUF1 (N20257, N20254);
or OR4 (N20258, N20257, N13446, N18009, N6276);
nand NAND3 (N20259, N20253, N11610, N3137);
xor XOR2 (N20260, N20258, N2201);
not NOT1 (N20261, N20244);
and AND4 (N20262, N20260, N14438, N7532, N11106);
xor XOR2 (N20263, N20242, N17948);
nor NOR2 (N20264, N20256, N1909);
buf BUF1 (N20265, N20232);
buf BUF1 (N20266, N20250);
not NOT1 (N20267, N20264);
buf BUF1 (N20268, N20263);
or OR3 (N20269, N20265, N5761, N9333);
nor NOR2 (N20270, N20252, N11346);
and AND4 (N20271, N20270, N18994, N18552, N16307);
buf BUF1 (N20272, N20271);
nand NAND2 (N20273, N20269, N10560);
nand NAND4 (N20274, N20262, N9832, N10352, N3155);
or OR3 (N20275, N20268, N11447, N591);
xor XOR2 (N20276, N20275, N874);
or OR4 (N20277, N20255, N10418, N415, N18595);
buf BUF1 (N20278, N20272);
and AND3 (N20279, N20261, N18491, N19416);
buf BUF1 (N20280, N20276);
xor XOR2 (N20281, N20273, N1031);
nor NOR3 (N20282, N20267, N17704, N3199);
nor NOR3 (N20283, N20274, N4486, N10431);
nor NOR2 (N20284, N20247, N12743);
nand NAND4 (N20285, N20277, N18745, N5280, N7900);
and AND3 (N20286, N20284, N4393, N7486);
nor NOR2 (N20287, N20281, N9903);
or OR3 (N20288, N20282, N5422, N13377);
not NOT1 (N20289, N20266);
or OR3 (N20290, N20279, N18507, N10397);
xor XOR2 (N20291, N20280, N17311);
and AND2 (N20292, N20259, N18695);
xor XOR2 (N20293, N20283, N13061);
nand NAND3 (N20294, N20289, N11477, N14040);
nand NAND4 (N20295, N20286, N125, N19479, N17476);
or OR2 (N20296, N20295, N2252);
not NOT1 (N20297, N20278);
and AND3 (N20298, N20290, N16738, N8284);
xor XOR2 (N20299, N20287, N9751);
and AND4 (N20300, N20297, N2088, N9839, N18794);
or OR4 (N20301, N20299, N6399, N17766, N6250);
xor XOR2 (N20302, N20300, N10616);
nor NOR3 (N20303, N20296, N9104, N3274);
nor NOR3 (N20304, N20292, N14576, N16710);
or OR2 (N20305, N20298, N249);
and AND3 (N20306, N20288, N2456, N9254);
not NOT1 (N20307, N20291);
xor XOR2 (N20308, N20293, N15092);
or OR4 (N20309, N20305, N11366, N14845, N10283);
nor NOR4 (N20310, N20301, N15896, N15229, N14580);
nand NAND4 (N20311, N20307, N3919, N17171, N15470);
nand NAND2 (N20312, N20303, N3614);
and AND2 (N20313, N20308, N6889);
xor XOR2 (N20314, N20313, N937);
nor NOR4 (N20315, N20310, N19156, N4211, N19163);
and AND4 (N20316, N20314, N2007, N13625, N14743);
and AND2 (N20317, N20312, N13012);
xor XOR2 (N20318, N20302, N17325);
not NOT1 (N20319, N20304);
xor XOR2 (N20320, N20319, N20078);
nand NAND2 (N20321, N20309, N1534);
or OR2 (N20322, N20317, N7520);
and AND4 (N20323, N20322, N7371, N1390, N14328);
and AND2 (N20324, N20306, N5380);
xor XOR2 (N20325, N20324, N10908);
nand NAND2 (N20326, N20321, N4312);
buf BUF1 (N20327, N20320);
buf BUF1 (N20328, N20326);
xor XOR2 (N20329, N20316, N3380);
xor XOR2 (N20330, N20329, N12077);
xor XOR2 (N20331, N20311, N10619);
xor XOR2 (N20332, N20323, N5802);
nor NOR2 (N20333, N20332, N12358);
nor NOR2 (N20334, N20315, N5384);
and AND3 (N20335, N20331, N10849, N11721);
buf BUF1 (N20336, N20327);
and AND2 (N20337, N20294, N12184);
or OR4 (N20338, N20336, N11698, N12322, N7919);
and AND4 (N20339, N20334, N11131, N4631, N18374);
and AND3 (N20340, N20328, N18224, N11437);
or OR2 (N20341, N20339, N12639);
xor XOR2 (N20342, N20318, N750);
and AND2 (N20343, N20341, N11573);
and AND3 (N20344, N20325, N18462, N12239);
buf BUF1 (N20345, N20338);
or OR2 (N20346, N20343, N15287);
buf BUF1 (N20347, N20333);
and AND4 (N20348, N20337, N8238, N16681, N15191);
or OR3 (N20349, N20346, N4078, N9752);
buf BUF1 (N20350, N20340);
or OR4 (N20351, N20342, N18173, N2961, N803);
xor XOR2 (N20352, N20344, N1873);
buf BUF1 (N20353, N20350);
not NOT1 (N20354, N20351);
buf BUF1 (N20355, N20335);
buf BUF1 (N20356, N20347);
nor NOR4 (N20357, N20353, N17282, N10678, N16725);
xor XOR2 (N20358, N20345, N4861);
nand NAND3 (N20359, N20348, N6722, N14584);
or OR2 (N20360, N20285, N981);
not NOT1 (N20361, N20356);
nor NOR4 (N20362, N20361, N18655, N20161, N13920);
buf BUF1 (N20363, N20360);
buf BUF1 (N20364, N20357);
or OR2 (N20365, N20359, N1212);
and AND4 (N20366, N20358, N442, N5724, N16908);
nand NAND2 (N20367, N20330, N13136);
xor XOR2 (N20368, N20367, N19069);
nand NAND2 (N20369, N20354, N13753);
xor XOR2 (N20370, N20365, N9465);
nor NOR4 (N20371, N20363, N6962, N17147, N2615);
or OR3 (N20372, N20364, N15932, N17372);
or OR4 (N20373, N20371, N12374, N877, N15217);
xor XOR2 (N20374, N20349, N2534);
and AND3 (N20375, N20373, N11322, N5840);
not NOT1 (N20376, N20355);
nor NOR3 (N20377, N20376, N17311, N15142);
nor NOR4 (N20378, N20377, N12100, N943, N15922);
not NOT1 (N20379, N20362);
nor NOR2 (N20380, N20379, N2899);
nor NOR4 (N20381, N20352, N5, N7093, N15667);
buf BUF1 (N20382, N20378);
and AND4 (N20383, N20374, N14092, N14442, N923);
nor NOR4 (N20384, N20375, N9918, N9017, N11695);
nor NOR2 (N20385, N20380, N16409);
nor NOR3 (N20386, N20385, N12242, N1375);
xor XOR2 (N20387, N20370, N3707);
xor XOR2 (N20388, N20386, N6200);
xor XOR2 (N20389, N20384, N19497);
buf BUF1 (N20390, N20369);
buf BUF1 (N20391, N20390);
and AND3 (N20392, N20387, N20267, N15033);
nor NOR2 (N20393, N20391, N20356);
and AND2 (N20394, N20393, N283);
nand NAND4 (N20395, N20389, N484, N20260, N8668);
and AND4 (N20396, N20368, N16657, N8246, N20252);
not NOT1 (N20397, N20396);
xor XOR2 (N20398, N20388, N11721);
nand NAND3 (N20399, N20392, N992, N20002);
nor NOR4 (N20400, N20372, N6174, N20397, N16882);
nor NOR4 (N20401, N6384, N7986, N7511, N13661);
xor XOR2 (N20402, N20400, N4395);
nor NOR4 (N20403, N20381, N7809, N9475, N2973);
xor XOR2 (N20404, N20383, N9296);
nand NAND3 (N20405, N20404, N18102, N16072);
buf BUF1 (N20406, N20402);
buf BUF1 (N20407, N20382);
nand NAND2 (N20408, N20401, N3670);
buf BUF1 (N20409, N20403);
not NOT1 (N20410, N20394);
or OR4 (N20411, N20407, N6706, N5245, N5248);
not NOT1 (N20412, N20411);
not NOT1 (N20413, N20410);
or OR3 (N20414, N20413, N11993, N8668);
nand NAND4 (N20415, N20412, N6924, N20382, N5472);
nor NOR2 (N20416, N20409, N11670);
buf BUF1 (N20417, N20366);
and AND4 (N20418, N20398, N17295, N6076, N4956);
not NOT1 (N20419, N20414);
nor NOR2 (N20420, N20406, N11771);
and AND4 (N20421, N20408, N14102, N15655, N2537);
and AND2 (N20422, N20416, N19924);
and AND4 (N20423, N20421, N18626, N9621, N16171);
nand NAND3 (N20424, N20423, N5647, N19350);
or OR3 (N20425, N20422, N562, N7494);
and AND2 (N20426, N20417, N16609);
buf BUF1 (N20427, N20399);
nand NAND3 (N20428, N20420, N14827, N10392);
or OR4 (N20429, N20415, N10511, N4053, N9134);
nor NOR4 (N20430, N20426, N58, N8999, N16513);
nor NOR3 (N20431, N20425, N4123, N11804);
not NOT1 (N20432, N20419);
and AND2 (N20433, N20405, N3123);
and AND4 (N20434, N20431, N12479, N18312, N15802);
nor NOR4 (N20435, N20432, N6695, N8165, N7176);
nand NAND4 (N20436, N20433, N16759, N13830, N3750);
and AND2 (N20437, N20430, N9311);
not NOT1 (N20438, N20434);
and AND2 (N20439, N20395, N20106);
or OR4 (N20440, N20436, N202, N16495, N6338);
nand NAND3 (N20441, N20428, N20269, N11193);
xor XOR2 (N20442, N20437, N7173);
nand NAND3 (N20443, N20429, N7435, N2876);
not NOT1 (N20444, N20424);
nand NAND3 (N20445, N20439, N6373, N20092);
buf BUF1 (N20446, N20444);
and AND3 (N20447, N20441, N1148, N16186);
nand NAND4 (N20448, N20418, N8678, N13960, N10705);
nor NOR4 (N20449, N20445, N2371, N1245, N4019);
and AND4 (N20450, N20427, N14736, N12381, N12596);
and AND2 (N20451, N20450, N11346);
nand NAND4 (N20452, N20451, N10263, N19604, N15913);
or OR3 (N20453, N20435, N16690, N17369);
or OR3 (N20454, N20443, N12383, N15885);
buf BUF1 (N20455, N20438);
xor XOR2 (N20456, N20440, N17458);
and AND4 (N20457, N20456, N1087, N16927, N13271);
not NOT1 (N20458, N20453);
buf BUF1 (N20459, N20447);
nand NAND2 (N20460, N20458, N258);
nor NOR4 (N20461, N20455, N10113, N3162, N18906);
nor NOR2 (N20462, N20442, N2422);
buf BUF1 (N20463, N20454);
nand NAND2 (N20464, N20446, N15648);
not NOT1 (N20465, N20464);
xor XOR2 (N20466, N20449, N5348);
not NOT1 (N20467, N20448);
xor XOR2 (N20468, N20461, N13498);
and AND2 (N20469, N20467, N11123);
xor XOR2 (N20470, N20469, N2771);
xor XOR2 (N20471, N20465, N10428);
or OR2 (N20472, N20470, N13437);
and AND2 (N20473, N20460, N15976);
buf BUF1 (N20474, N20452);
or OR3 (N20475, N20468, N10188, N6419);
xor XOR2 (N20476, N20475, N13552);
buf BUF1 (N20477, N20472);
not NOT1 (N20478, N20466);
and AND2 (N20479, N20463, N1227);
nand NAND2 (N20480, N20479, N13461);
xor XOR2 (N20481, N20478, N1328);
buf BUF1 (N20482, N20459);
and AND2 (N20483, N20476, N19083);
nor NOR2 (N20484, N20480, N12209);
or OR4 (N20485, N20471, N4876, N13772, N6588);
not NOT1 (N20486, N20473);
nand NAND4 (N20487, N20486, N14644, N7063, N11202);
buf BUF1 (N20488, N20483);
buf BUF1 (N20489, N20484);
buf BUF1 (N20490, N20477);
nand NAND4 (N20491, N20485, N17322, N20194, N7548);
or OR4 (N20492, N20488, N19843, N12102, N13475);
and AND3 (N20493, N20492, N1871, N7151);
nor NOR2 (N20494, N20489, N4086);
or OR2 (N20495, N20482, N18563);
nand NAND2 (N20496, N20491, N19200);
and AND2 (N20497, N20474, N20487);
and AND2 (N20498, N5075, N5442);
and AND2 (N20499, N20457, N7371);
nor NOR3 (N20500, N20495, N4076, N11075);
xor XOR2 (N20501, N20493, N3697);
xor XOR2 (N20502, N20499, N12218);
and AND4 (N20503, N20497, N14550, N3226, N13281);
buf BUF1 (N20504, N20494);
nand NAND3 (N20505, N20462, N15326, N15793);
or OR2 (N20506, N20490, N390);
or OR4 (N20507, N20498, N16609, N2360, N1267);
nand NAND3 (N20508, N20501, N4204, N8399);
not NOT1 (N20509, N20503);
nand NAND2 (N20510, N20496, N17609);
and AND2 (N20511, N20508, N1659);
xor XOR2 (N20512, N20506, N18843);
not NOT1 (N20513, N20507);
buf BUF1 (N20514, N20500);
not NOT1 (N20515, N20511);
and AND2 (N20516, N20512, N12833);
buf BUF1 (N20517, N20510);
nand NAND4 (N20518, N20481, N15051, N14573, N296);
not NOT1 (N20519, N20518);
buf BUF1 (N20520, N20519);
buf BUF1 (N20521, N20514);
not NOT1 (N20522, N20515);
or OR4 (N20523, N20509, N17030, N630, N18424);
not NOT1 (N20524, N20517);
nor NOR3 (N20525, N20520, N20498, N4014);
or OR2 (N20526, N20504, N11303);
buf BUF1 (N20527, N20526);
xor XOR2 (N20528, N20523, N5446);
xor XOR2 (N20529, N20524, N10662);
and AND3 (N20530, N20522, N1027, N13324);
nor NOR2 (N20531, N20505, N16318);
or OR2 (N20532, N20502, N3651);
buf BUF1 (N20533, N20532);
and AND2 (N20534, N20530, N7694);
nor NOR4 (N20535, N20531, N12352, N6360, N5661);
nand NAND4 (N20536, N20533, N9272, N1684, N19866);
or OR4 (N20537, N20527, N2714, N10697, N17653);
or OR3 (N20538, N20534, N16467, N12006);
and AND2 (N20539, N20513, N16759);
buf BUF1 (N20540, N20539);
nand NAND4 (N20541, N20538, N11916, N2333, N16524);
nor NOR3 (N20542, N20529, N12915, N2814);
and AND2 (N20543, N20516, N293);
not NOT1 (N20544, N20540);
xor XOR2 (N20545, N20544, N7178);
or OR3 (N20546, N20521, N7371, N6117);
and AND3 (N20547, N20543, N8589, N14088);
and AND3 (N20548, N20546, N12362, N457);
nor NOR4 (N20549, N20547, N14084, N11057, N5776);
or OR3 (N20550, N20525, N15085, N3591);
or OR2 (N20551, N20542, N17336);
nand NAND4 (N20552, N20549, N20234, N5886, N2622);
buf BUF1 (N20553, N20537);
not NOT1 (N20554, N20528);
buf BUF1 (N20555, N20552);
or OR2 (N20556, N20555, N13773);
or OR2 (N20557, N20553, N16256);
not NOT1 (N20558, N20535);
or OR2 (N20559, N20548, N12783);
nor NOR4 (N20560, N20558, N2108, N12835, N8025);
nand NAND2 (N20561, N20550, N9582);
not NOT1 (N20562, N20560);
or OR4 (N20563, N20562, N15384, N18721, N6395);
xor XOR2 (N20564, N20541, N8237);
or OR2 (N20565, N20557, N2997);
and AND2 (N20566, N20564, N14728);
buf BUF1 (N20567, N20545);
and AND3 (N20568, N20566, N14546, N16344);
nor NOR4 (N20569, N20563, N13830, N18721, N13351);
and AND3 (N20570, N20561, N6636, N17935);
nand NAND2 (N20571, N20554, N12243);
xor XOR2 (N20572, N20551, N14525);
and AND2 (N20573, N20567, N20131);
buf BUF1 (N20574, N20569);
buf BUF1 (N20575, N20571);
not NOT1 (N20576, N20568);
and AND4 (N20577, N20559, N9316, N2177, N8963);
not NOT1 (N20578, N20574);
nor NOR3 (N20579, N20556, N2235, N11577);
not NOT1 (N20580, N20576);
and AND2 (N20581, N20565, N15723);
nor NOR3 (N20582, N20573, N15332, N6446);
buf BUF1 (N20583, N20581);
and AND3 (N20584, N20580, N2012, N9949);
nand NAND4 (N20585, N20582, N4348, N3886, N12836);
not NOT1 (N20586, N20570);
and AND4 (N20587, N20572, N9342, N6392, N19327);
not NOT1 (N20588, N20584);
buf BUF1 (N20589, N20587);
nor NOR4 (N20590, N20577, N8738, N742, N12056);
and AND4 (N20591, N20585, N16621, N15898, N12829);
buf BUF1 (N20592, N20591);
buf BUF1 (N20593, N20588);
buf BUF1 (N20594, N20579);
nor NOR2 (N20595, N20594, N15001);
nand NAND2 (N20596, N20589, N4385);
not NOT1 (N20597, N20575);
not NOT1 (N20598, N20536);
not NOT1 (N20599, N20595);
not NOT1 (N20600, N20599);
nor NOR2 (N20601, N20600, N7500);
not NOT1 (N20602, N20592);
nand NAND2 (N20603, N20596, N3074);
nor NOR2 (N20604, N20603, N18221);
and AND4 (N20605, N20578, N14164, N11908, N6793);
or OR3 (N20606, N20602, N18190, N10110);
nand NAND3 (N20607, N20606, N6613, N19823);
and AND2 (N20608, N20590, N2492);
buf BUF1 (N20609, N20593);
xor XOR2 (N20610, N20607, N17285);
and AND3 (N20611, N20586, N1568, N9502);
nand NAND4 (N20612, N20597, N15703, N11859, N16713);
and AND2 (N20613, N20598, N19830);
not NOT1 (N20614, N20608);
nor NOR2 (N20615, N20613, N12001);
buf BUF1 (N20616, N20614);
xor XOR2 (N20617, N20610, N3338);
buf BUF1 (N20618, N20605);
not NOT1 (N20619, N20583);
xor XOR2 (N20620, N20612, N1728);
xor XOR2 (N20621, N20617, N19146);
or OR4 (N20622, N20621, N10650, N5845, N9455);
nor NOR3 (N20623, N20604, N3426, N10441);
not NOT1 (N20624, N20611);
nand NAND2 (N20625, N20623, N10198);
nand NAND2 (N20626, N20615, N13152);
xor XOR2 (N20627, N20609, N6459);
nor NOR3 (N20628, N20616, N13544, N7955);
or OR3 (N20629, N20620, N18170, N12418);
or OR4 (N20630, N20625, N16470, N1520, N6508);
and AND4 (N20631, N20629, N18420, N10454, N5551);
xor XOR2 (N20632, N20626, N13070);
buf BUF1 (N20633, N20601);
buf BUF1 (N20634, N20630);
or OR2 (N20635, N20628, N17035);
or OR4 (N20636, N20624, N14639, N12904, N19769);
nor NOR3 (N20637, N20619, N13888, N17655);
and AND3 (N20638, N20627, N6044, N1070);
and AND4 (N20639, N20637, N4927, N9018, N171);
nor NOR2 (N20640, N20639, N2944);
nand NAND2 (N20641, N20632, N4448);
nand NAND4 (N20642, N20638, N4920, N13595, N6328);
not NOT1 (N20643, N20642);
nand NAND4 (N20644, N20631, N13113, N5523, N2748);
nand NAND3 (N20645, N20622, N8107, N5050);
or OR2 (N20646, N20633, N14822);
not NOT1 (N20647, N20643);
or OR3 (N20648, N20636, N12156, N1425);
or OR4 (N20649, N20635, N1578, N7997, N1566);
buf BUF1 (N20650, N20618);
and AND2 (N20651, N20644, N1197);
buf BUF1 (N20652, N20634);
buf BUF1 (N20653, N20650);
buf BUF1 (N20654, N20646);
nor NOR3 (N20655, N20647, N12554, N18552);
nand NAND3 (N20656, N20641, N8413, N3498);
nand NAND3 (N20657, N20656, N12625, N1938);
and AND2 (N20658, N20640, N16545);
nand NAND4 (N20659, N20645, N10586, N11247, N10847);
nor NOR4 (N20660, N20657, N9092, N14419, N19287);
and AND4 (N20661, N20655, N4658, N19400, N5262);
or OR4 (N20662, N20654, N16803, N475, N3731);
and AND2 (N20663, N20660, N11990);
or OR4 (N20664, N20663, N18090, N18378, N5626);
xor XOR2 (N20665, N20658, N6326);
and AND4 (N20666, N20648, N8435, N16053, N10567);
buf BUF1 (N20667, N20662);
xor XOR2 (N20668, N20664, N13006);
and AND3 (N20669, N20659, N16589, N6767);
and AND2 (N20670, N20649, N16768);
buf BUF1 (N20671, N20653);
nand NAND2 (N20672, N20671, N11574);
or OR3 (N20673, N20669, N1650, N4196);
nor NOR4 (N20674, N20670, N18417, N10880, N69);
buf BUF1 (N20675, N20672);
buf BUF1 (N20676, N20675);
or OR3 (N20677, N20673, N14974, N18210);
buf BUF1 (N20678, N20652);
buf BUF1 (N20679, N20678);
not NOT1 (N20680, N20674);
nand NAND4 (N20681, N20665, N14259, N18745, N4603);
nand NAND2 (N20682, N20651, N8136);
nand NAND2 (N20683, N20661, N8475);
or OR4 (N20684, N20668, N3529, N7220, N15556);
or OR3 (N20685, N20667, N11869, N891);
not NOT1 (N20686, N20676);
or OR2 (N20687, N20680, N3072);
buf BUF1 (N20688, N20677);
buf BUF1 (N20689, N20688);
buf BUF1 (N20690, N20689);
nor NOR4 (N20691, N20690, N14582, N17095, N5718);
nand NAND3 (N20692, N20685, N7026, N18904);
nand NAND2 (N20693, N20692, N20117);
buf BUF1 (N20694, N20684);
xor XOR2 (N20695, N20679, N7877);
nand NAND4 (N20696, N20683, N9695, N13676, N2477);
xor XOR2 (N20697, N20691, N9668);
nor NOR2 (N20698, N20681, N12856);
nand NAND2 (N20699, N20682, N8423);
xor XOR2 (N20700, N20666, N1765);
and AND2 (N20701, N20687, N19512);
nor NOR2 (N20702, N20699, N19586);
and AND4 (N20703, N20686, N8321, N14154, N10652);
or OR4 (N20704, N20703, N17347, N7022, N20203);
nand NAND2 (N20705, N20697, N10358);
and AND4 (N20706, N20694, N15685, N15892, N7560);
buf BUF1 (N20707, N20693);
nor NOR4 (N20708, N20700, N4179, N12383, N17167);
xor XOR2 (N20709, N20696, N16949);
or OR3 (N20710, N20695, N9000, N3449);
not NOT1 (N20711, N20704);
buf BUF1 (N20712, N20708);
nor NOR2 (N20713, N20709, N12579);
nand NAND3 (N20714, N20705, N19902, N14596);
xor XOR2 (N20715, N20702, N2113);
not NOT1 (N20716, N20712);
not NOT1 (N20717, N20716);
nor NOR2 (N20718, N20701, N2587);
and AND4 (N20719, N20698, N13304, N12221, N5062);
or OR4 (N20720, N20713, N20613, N10541, N14674);
and AND2 (N20721, N20711, N9949);
or OR3 (N20722, N20707, N15956, N3875);
not NOT1 (N20723, N20717);
nor NOR2 (N20724, N20723, N18549);
or OR4 (N20725, N20719, N13636, N1731, N17149);
nor NOR2 (N20726, N20720, N2304);
nand NAND2 (N20727, N20715, N5405);
and AND3 (N20728, N20727, N17889, N1583);
nand NAND4 (N20729, N20706, N2735, N2626, N1511);
nand NAND4 (N20730, N20729, N11385, N5076, N1307);
and AND3 (N20731, N20730, N8512, N10515);
xor XOR2 (N20732, N20714, N11311);
xor XOR2 (N20733, N20722, N19439);
and AND3 (N20734, N20725, N8033, N4221);
buf BUF1 (N20735, N20734);
nand NAND4 (N20736, N20731, N8648, N9593, N18191);
nand NAND4 (N20737, N20718, N8170, N9547, N11707);
buf BUF1 (N20738, N20721);
buf BUF1 (N20739, N20724);
and AND3 (N20740, N20736, N7587, N15043);
nand NAND2 (N20741, N20726, N10184);
nor NOR3 (N20742, N20737, N136, N15994);
and AND4 (N20743, N20738, N14094, N9272, N9964);
not NOT1 (N20744, N20743);
not NOT1 (N20745, N20732);
nand NAND2 (N20746, N20735, N2868);
and AND2 (N20747, N20728, N9420);
buf BUF1 (N20748, N20744);
buf BUF1 (N20749, N20742);
xor XOR2 (N20750, N20748, N13640);
nor NOR2 (N20751, N20739, N16153);
buf BUF1 (N20752, N20751);
nor NOR2 (N20753, N20747, N11187);
nor NOR2 (N20754, N20733, N7216);
nand NAND2 (N20755, N20745, N9716);
not NOT1 (N20756, N20752);
nand NAND2 (N20757, N20756, N15076);
and AND4 (N20758, N20755, N20470, N7263, N7896);
buf BUF1 (N20759, N20710);
nand NAND4 (N20760, N20754, N12950, N1394, N7366);
xor XOR2 (N20761, N20759, N9553);
nor NOR3 (N20762, N20753, N2805, N5097);
nor NOR4 (N20763, N20757, N260, N8300, N7610);
xor XOR2 (N20764, N20750, N9463);
nor NOR3 (N20765, N20762, N10823, N15654);
buf BUF1 (N20766, N20760);
nor NOR2 (N20767, N20764, N2547);
buf BUF1 (N20768, N20758);
not NOT1 (N20769, N20761);
nand NAND4 (N20770, N20740, N15080, N17542, N4733);
and AND4 (N20771, N20746, N13376, N1182, N17606);
xor XOR2 (N20772, N20770, N2592);
nor NOR3 (N20773, N20766, N11558, N15238);
and AND3 (N20774, N20769, N13597, N4979);
nor NOR4 (N20775, N20768, N837, N4308, N15438);
xor XOR2 (N20776, N20775, N14930);
and AND3 (N20777, N20774, N10517, N10418);
or OR2 (N20778, N20771, N2027);
xor XOR2 (N20779, N20767, N18231);
buf BUF1 (N20780, N20765);
not NOT1 (N20781, N20741);
xor XOR2 (N20782, N20772, N17299);
nand NAND2 (N20783, N20777, N9565);
and AND4 (N20784, N20778, N13562, N1990, N11775);
or OR4 (N20785, N20781, N8622, N18522, N11384);
or OR4 (N20786, N20783, N7576, N15685, N13344);
or OR3 (N20787, N20763, N7792, N4809);
xor XOR2 (N20788, N20780, N6482);
nand NAND3 (N20789, N20786, N17975, N3929);
nor NOR3 (N20790, N20789, N8633, N4029);
buf BUF1 (N20791, N20779);
and AND4 (N20792, N20785, N14978, N6165, N4770);
or OR2 (N20793, N20791, N2815);
buf BUF1 (N20794, N20773);
or OR4 (N20795, N20776, N12212, N17527, N12796);
xor XOR2 (N20796, N20792, N17228);
nand NAND2 (N20797, N20796, N17633);
and AND4 (N20798, N20793, N6720, N9643, N6143);
and AND2 (N20799, N20784, N3525);
xor XOR2 (N20800, N20749, N6650);
nor NOR3 (N20801, N20800, N9774, N16762);
xor XOR2 (N20802, N20795, N3992);
or OR3 (N20803, N20798, N17283, N7511);
nand NAND4 (N20804, N20803, N9542, N490, N17339);
not NOT1 (N20805, N20797);
not NOT1 (N20806, N20802);
nor NOR2 (N20807, N20788, N2586);
and AND2 (N20808, N20806, N6600);
nor NOR3 (N20809, N20799, N3998, N6627);
and AND3 (N20810, N20808, N9537, N14096);
xor XOR2 (N20811, N20790, N14442);
buf BUF1 (N20812, N20804);
or OR2 (N20813, N20787, N5106);
xor XOR2 (N20814, N20810, N14858);
nand NAND4 (N20815, N20794, N1492, N6632, N39);
buf BUF1 (N20816, N20807);
not NOT1 (N20817, N20811);
xor XOR2 (N20818, N20814, N751);
xor XOR2 (N20819, N20816, N5525);
buf BUF1 (N20820, N20809);
buf BUF1 (N20821, N20805);
xor XOR2 (N20822, N20818, N11245);
nand NAND4 (N20823, N20817, N1004, N849, N13556);
buf BUF1 (N20824, N20782);
or OR2 (N20825, N20824, N6349);
xor XOR2 (N20826, N20825, N15885);
and AND4 (N20827, N20821, N13185, N9791, N11876);
xor XOR2 (N20828, N20815, N2694);
and AND2 (N20829, N20822, N8676);
and AND4 (N20830, N20826, N7172, N18404, N4934);
and AND4 (N20831, N20823, N8008, N14376, N5143);
buf BUF1 (N20832, N20819);
nand NAND4 (N20833, N20827, N9694, N4942, N19368);
or OR4 (N20834, N20820, N17239, N11899, N10733);
nor NOR4 (N20835, N20830, N12370, N7759, N12384);
not NOT1 (N20836, N20828);
nor NOR4 (N20837, N20834, N18295, N8053, N7481);
and AND3 (N20838, N20813, N14543, N5286);
xor XOR2 (N20839, N20832, N9443);
nor NOR4 (N20840, N20838, N619, N574, N11761);
buf BUF1 (N20841, N20837);
or OR3 (N20842, N20840, N19143, N12450);
and AND2 (N20843, N20839, N1434);
xor XOR2 (N20844, N20843, N7546);
nor NOR4 (N20845, N20836, N15465, N12026, N20293);
nand NAND3 (N20846, N20812, N7866, N507);
and AND2 (N20847, N20835, N18004);
nor NOR3 (N20848, N20846, N13427, N13681);
nor NOR2 (N20849, N20801, N2134);
nand NAND4 (N20850, N20844, N15275, N12862, N17381);
not NOT1 (N20851, N20850);
nand NAND4 (N20852, N20847, N14918, N3814, N17853);
nand NAND2 (N20853, N20841, N18235);
and AND2 (N20854, N20852, N437);
not NOT1 (N20855, N20829);
nand NAND3 (N20856, N20854, N11357, N18371);
buf BUF1 (N20857, N20833);
nor NOR3 (N20858, N20851, N4607, N15336);
not NOT1 (N20859, N20849);
nand NAND2 (N20860, N20859, N4101);
nand NAND4 (N20861, N20848, N14844, N11156, N6447);
xor XOR2 (N20862, N20853, N7039);
nand NAND2 (N20863, N20855, N11257);
nor NOR4 (N20864, N20842, N8892, N11018, N1035);
not NOT1 (N20865, N20857);
not NOT1 (N20866, N20858);
and AND2 (N20867, N20860, N720);
and AND4 (N20868, N20861, N9508, N1635, N8742);
nand NAND2 (N20869, N20856, N11902);
nor NOR2 (N20870, N20865, N16200);
nor NOR4 (N20871, N20866, N11118, N16021, N19852);
not NOT1 (N20872, N20862);
or OR3 (N20873, N20870, N1872, N11267);
xor XOR2 (N20874, N20863, N18287);
xor XOR2 (N20875, N20871, N10607);
nor NOR3 (N20876, N20872, N12545, N19052);
buf BUF1 (N20877, N20873);
or OR3 (N20878, N20875, N3791, N8521);
or OR3 (N20879, N20869, N2260, N18793);
and AND4 (N20880, N20831, N20665, N7602, N13631);
not NOT1 (N20881, N20868);
or OR4 (N20882, N20874, N15244, N10416, N11830);
buf BUF1 (N20883, N20845);
nand NAND3 (N20884, N20882, N5097, N10829);
or OR3 (N20885, N20880, N10490, N17644);
buf BUF1 (N20886, N20885);
buf BUF1 (N20887, N20876);
xor XOR2 (N20888, N20883, N5038);
xor XOR2 (N20889, N20879, N3327);
nor NOR3 (N20890, N20889, N17083, N12944);
nor NOR2 (N20891, N20881, N5034);
buf BUF1 (N20892, N20867);
not NOT1 (N20893, N20884);
and AND4 (N20894, N20891, N17330, N7961, N9742);
nor NOR2 (N20895, N20887, N15958);
nor NOR4 (N20896, N20892, N18647, N6212, N9564);
buf BUF1 (N20897, N20895);
buf BUF1 (N20898, N20877);
and AND3 (N20899, N20894, N18452, N19454);
and AND4 (N20900, N20893, N17658, N9814, N6271);
and AND3 (N20901, N20878, N3893, N4703);
not NOT1 (N20902, N20900);
nand NAND2 (N20903, N20899, N10574);
and AND2 (N20904, N20897, N2986);
xor XOR2 (N20905, N20864, N11481);
and AND4 (N20906, N20898, N7063, N12101, N10454);
nand NAND4 (N20907, N20904, N10711, N1047, N10514);
nand NAND4 (N20908, N20896, N672, N10333, N118);
not NOT1 (N20909, N20903);
or OR2 (N20910, N20908, N20559);
nor NOR4 (N20911, N20910, N20567, N6070, N7578);
not NOT1 (N20912, N20909);
not NOT1 (N20913, N20911);
xor XOR2 (N20914, N20905, N14023);
nand NAND3 (N20915, N20913, N18461, N17902);
xor XOR2 (N20916, N20914, N15991);
or OR3 (N20917, N20907, N3505, N19226);
and AND3 (N20918, N20901, N2615, N7453);
buf BUF1 (N20919, N20912);
xor XOR2 (N20920, N20916, N2026);
xor XOR2 (N20921, N20902, N3083);
nand NAND4 (N20922, N20919, N1902, N4115, N7147);
or OR4 (N20923, N20917, N2427, N10823, N8880);
nand NAND4 (N20924, N20923, N13174, N13528, N19977);
xor XOR2 (N20925, N20886, N5707);
not NOT1 (N20926, N20920);
nand NAND2 (N20927, N20888, N7477);
not NOT1 (N20928, N20890);
and AND3 (N20929, N20927, N17580, N1976);
not NOT1 (N20930, N20926);
nand NAND3 (N20931, N20930, N14007, N2642);
nor NOR2 (N20932, N20921, N7842);
or OR4 (N20933, N20929, N9455, N8720, N9137);
or OR4 (N20934, N20931, N17489, N7006, N6559);
xor XOR2 (N20935, N20918, N9030);
buf BUF1 (N20936, N20906);
xor XOR2 (N20937, N20915, N133);
nor NOR3 (N20938, N20924, N6779, N11653);
not NOT1 (N20939, N20925);
and AND4 (N20940, N20936, N11058, N19422, N20236);
xor XOR2 (N20941, N20937, N16400);
nand NAND4 (N20942, N20940, N830, N5581, N13210);
buf BUF1 (N20943, N20939);
not NOT1 (N20944, N20934);
or OR2 (N20945, N20944, N15191);
xor XOR2 (N20946, N20935, N13522);
nor NOR3 (N20947, N20928, N15377, N9907);
nor NOR2 (N20948, N20933, N4883);
xor XOR2 (N20949, N20943, N8738);
xor XOR2 (N20950, N20949, N17840);
nand NAND3 (N20951, N20942, N4864, N2021);
nor NOR3 (N20952, N20941, N15726, N9943);
buf BUF1 (N20953, N20948);
and AND4 (N20954, N20945, N20306, N16211, N6989);
nor NOR3 (N20955, N20932, N8353, N5461);
and AND4 (N20956, N20951, N11526, N14752, N768);
nand NAND4 (N20957, N20946, N15331, N17490, N15575);
nand NAND4 (N20958, N20938, N9088, N5557, N13495);
nand NAND2 (N20959, N20955, N15994);
nand NAND3 (N20960, N20959, N17596, N7808);
or OR4 (N20961, N20953, N17750, N18856, N4131);
nand NAND2 (N20962, N20947, N17907);
nor NOR2 (N20963, N20922, N4718);
or OR2 (N20964, N20958, N10711);
or OR2 (N20965, N20960, N5521);
and AND4 (N20966, N20956, N10718, N19721, N15144);
not NOT1 (N20967, N20964);
and AND2 (N20968, N20963, N17133);
and AND3 (N20969, N20950, N17403, N10449);
nor NOR3 (N20970, N20965, N14389, N19076);
nor NOR4 (N20971, N20968, N9728, N9181, N2529);
not NOT1 (N20972, N20966);
nor NOR2 (N20973, N20972, N5797);
xor XOR2 (N20974, N20952, N12623);
nand NAND2 (N20975, N20957, N13062);
or OR4 (N20976, N20970, N657, N11430, N3675);
and AND2 (N20977, N20976, N8778);
not NOT1 (N20978, N20969);
not NOT1 (N20979, N20967);
and AND4 (N20980, N20961, N10995, N4152, N322);
nor NOR4 (N20981, N20971, N7365, N13911, N11400);
or OR2 (N20982, N20975, N10487);
nor NOR3 (N20983, N20979, N4440, N15207);
xor XOR2 (N20984, N20981, N14129);
not NOT1 (N20985, N20954);
or OR4 (N20986, N20980, N12953, N18800, N1015);
and AND3 (N20987, N20974, N9984, N12572);
xor XOR2 (N20988, N20984, N1737);
buf BUF1 (N20989, N20985);
nor NOR3 (N20990, N20962, N8341, N2803);
nand NAND3 (N20991, N20973, N8431, N17378);
nor NOR3 (N20992, N20990, N20632, N14016);
nor NOR3 (N20993, N20992, N3253, N9045);
not NOT1 (N20994, N20989);
or OR4 (N20995, N20978, N2069, N11496, N20986);
buf BUF1 (N20996, N9661);
nand NAND4 (N20997, N20977, N3963, N14266, N9714);
nand NAND2 (N20998, N20987, N304);
nand NAND2 (N20999, N20995, N808);
and AND4 (N21000, N20993, N4181, N3661, N4690);
xor XOR2 (N21001, N20994, N16504);
or OR4 (N21002, N20983, N18538, N6465, N12208);
buf BUF1 (N21003, N20991);
buf BUF1 (N21004, N21003);
nor NOR3 (N21005, N20988, N5568, N11796);
or OR3 (N21006, N20998, N9068, N3136);
and AND2 (N21007, N21006, N1503);
xor XOR2 (N21008, N21001, N2872);
buf BUF1 (N21009, N21005);
nor NOR2 (N21010, N21000, N13630);
not NOT1 (N21011, N20982);
nor NOR3 (N21012, N20996, N460, N13465);
or OR4 (N21013, N20997, N20369, N1537, N17967);
nor NOR3 (N21014, N21011, N14072, N2421);
nor NOR2 (N21015, N21008, N1702);
nand NAND2 (N21016, N21002, N19711);
not NOT1 (N21017, N21010);
xor XOR2 (N21018, N21014, N2269);
nor NOR3 (N21019, N21018, N4897, N20620);
buf BUF1 (N21020, N20999);
not NOT1 (N21021, N21009);
or OR3 (N21022, N21020, N6857, N19992);
and AND2 (N21023, N21015, N2481);
not NOT1 (N21024, N21016);
or OR2 (N21025, N21021, N10729);
xor XOR2 (N21026, N21012, N19867);
buf BUF1 (N21027, N21024);
or OR2 (N21028, N21017, N9267);
xor XOR2 (N21029, N21028, N16208);
buf BUF1 (N21030, N21013);
not NOT1 (N21031, N21019);
nor NOR3 (N21032, N21026, N18709, N20575);
nand NAND3 (N21033, N21031, N12299, N19227);
or OR2 (N21034, N21025, N5898);
buf BUF1 (N21035, N21033);
buf BUF1 (N21036, N21034);
not NOT1 (N21037, N21022);
buf BUF1 (N21038, N21032);
buf BUF1 (N21039, N21007);
buf BUF1 (N21040, N21036);
nand NAND3 (N21041, N21039, N20988, N15669);
and AND3 (N21042, N21029, N8756, N17588);
and AND4 (N21043, N21035, N17323, N16734, N13333);
nor NOR4 (N21044, N21038, N7253, N18190, N20467);
nor NOR3 (N21045, N21023, N1648, N93);
xor XOR2 (N21046, N21040, N15689);
nor NOR4 (N21047, N21037, N18419, N918, N19106);
or OR2 (N21048, N21047, N11068);
or OR3 (N21049, N21046, N9370, N5550);
nor NOR4 (N21050, N21044, N4324, N16725, N11589);
nand NAND2 (N21051, N21050, N6103);
and AND4 (N21052, N21043, N15217, N5132, N12853);
not NOT1 (N21053, N21004);
xor XOR2 (N21054, N21048, N14151);
and AND4 (N21055, N21041, N18534, N8324, N18112);
nor NOR2 (N21056, N21053, N5197);
and AND4 (N21057, N21055, N18089, N15842, N13628);
nor NOR3 (N21058, N21057, N8569, N19297);
not NOT1 (N21059, N21054);
and AND2 (N21060, N21059, N14656);
and AND3 (N21061, N21049, N11091, N10075);
xor XOR2 (N21062, N21027, N14217);
not NOT1 (N21063, N21052);
xor XOR2 (N21064, N21056, N11749);
xor XOR2 (N21065, N21058, N2833);
not NOT1 (N21066, N21065);
and AND2 (N21067, N21051, N5323);
nor NOR2 (N21068, N21063, N600);
nor NOR2 (N21069, N21061, N7002);
nor NOR4 (N21070, N21062, N7846, N3122, N11371);
or OR2 (N21071, N21042, N8288);
nor NOR2 (N21072, N21067, N10264);
buf BUF1 (N21073, N21064);
not NOT1 (N21074, N21069);
nor NOR3 (N21075, N21045, N15858, N17952);
xor XOR2 (N21076, N21075, N16082);
nor NOR4 (N21077, N21074, N6260, N8884, N7108);
nor NOR4 (N21078, N21071, N575, N11298, N7770);
and AND2 (N21079, N21030, N6798);
and AND3 (N21080, N21066, N1461, N820);
nor NOR4 (N21081, N21070, N548, N6883, N6929);
buf BUF1 (N21082, N21079);
not NOT1 (N21083, N21077);
and AND4 (N21084, N21080, N930, N4919, N7892);
xor XOR2 (N21085, N21083, N6980);
nor NOR3 (N21086, N21082, N6146, N7752);
xor XOR2 (N21087, N21084, N14638);
or OR2 (N21088, N21087, N11056);
not NOT1 (N21089, N21081);
and AND4 (N21090, N21078, N10386, N13029, N14427);
and AND2 (N21091, N21089, N9551);
nand NAND3 (N21092, N21073, N13415, N14130);
or OR3 (N21093, N21086, N4940, N13850);
xor XOR2 (N21094, N21085, N2767);
or OR3 (N21095, N21092, N9216, N8867);
buf BUF1 (N21096, N21094);
not NOT1 (N21097, N21095);
and AND4 (N21098, N21088, N12897, N20522, N10545);
xor XOR2 (N21099, N21091, N18084);
buf BUF1 (N21100, N21096);
or OR2 (N21101, N21098, N19149);
buf BUF1 (N21102, N21090);
and AND3 (N21103, N21102, N7976, N16319);
not NOT1 (N21104, N21100);
not NOT1 (N21105, N21104);
xor XOR2 (N21106, N21101, N4238);
nand NAND4 (N21107, N21072, N8718, N12782, N14220);
buf BUF1 (N21108, N21076);
buf BUF1 (N21109, N21093);
xor XOR2 (N21110, N21106, N14322);
nand NAND2 (N21111, N21103, N1422);
not NOT1 (N21112, N21107);
nor NOR3 (N21113, N21111, N6408, N4248);
or OR3 (N21114, N21109, N7854, N20213);
not NOT1 (N21115, N21105);
or OR2 (N21116, N21108, N2494);
xor XOR2 (N21117, N21110, N9603);
not NOT1 (N21118, N21116);
or OR2 (N21119, N21099, N17777);
not NOT1 (N21120, N21060);
xor XOR2 (N21121, N21119, N5886);
and AND3 (N21122, N21113, N5373, N17731);
and AND4 (N21123, N21115, N16377, N20582, N17029);
xor XOR2 (N21124, N21118, N15609);
xor XOR2 (N21125, N21114, N7996);
nand NAND3 (N21126, N21121, N17400, N4817);
nor NOR4 (N21127, N21123, N18311, N9670, N1041);
nor NOR3 (N21128, N21126, N19777, N3660);
nor NOR4 (N21129, N21125, N13027, N2474, N9300);
xor XOR2 (N21130, N21129, N632);
nor NOR2 (N21131, N21128, N14652);
and AND2 (N21132, N21117, N19902);
nor NOR3 (N21133, N21120, N8357, N13688);
xor XOR2 (N21134, N21130, N8698);
xor XOR2 (N21135, N21122, N19294);
nand NAND4 (N21136, N21127, N12009, N17567, N19810);
or OR3 (N21137, N21097, N9453, N13608);
and AND3 (N21138, N21135, N16735, N8780);
buf BUF1 (N21139, N21136);
not NOT1 (N21140, N21132);
nand NAND2 (N21141, N21137, N20413);
xor XOR2 (N21142, N21124, N21110);
and AND3 (N21143, N21140, N1924, N345);
or OR4 (N21144, N21133, N6896, N7661, N19850);
nor NOR4 (N21145, N21142, N5598, N15957, N2875);
not NOT1 (N21146, N21068);
nand NAND4 (N21147, N21139, N4102, N7659, N10026);
and AND3 (N21148, N21147, N12954, N11078);
nand NAND4 (N21149, N21143, N2673, N5942, N4698);
buf BUF1 (N21150, N21145);
buf BUF1 (N21151, N21138);
not NOT1 (N21152, N21144);
or OR4 (N21153, N21141, N17846, N4219, N21083);
and AND4 (N21154, N21112, N15471, N13136, N9286);
buf BUF1 (N21155, N21149);
not NOT1 (N21156, N21131);
and AND3 (N21157, N21146, N7826, N8114);
not NOT1 (N21158, N21156);
not NOT1 (N21159, N21152);
not NOT1 (N21160, N21158);
buf BUF1 (N21161, N21155);
xor XOR2 (N21162, N21134, N14578);
nor NOR3 (N21163, N21153, N16257, N14863);
or OR4 (N21164, N21150, N5829, N20284, N20526);
and AND4 (N21165, N21157, N1281, N20420, N18171);
not NOT1 (N21166, N21154);
buf BUF1 (N21167, N21151);
nor NOR3 (N21168, N21162, N8335, N10137);
xor XOR2 (N21169, N21168, N11157);
nor NOR4 (N21170, N21165, N7568, N19051, N16405);
and AND3 (N21171, N21169, N16668, N13102);
xor XOR2 (N21172, N21163, N14550);
or OR3 (N21173, N21161, N1446, N19460);
nor NOR4 (N21174, N21173, N21098, N3890, N530);
buf BUF1 (N21175, N21164);
and AND3 (N21176, N21174, N2159, N16297);
not NOT1 (N21177, N21160);
buf BUF1 (N21178, N21167);
buf BUF1 (N21179, N21166);
and AND4 (N21180, N21171, N9989, N7860, N17094);
nand NAND2 (N21181, N21176, N2459);
nor NOR4 (N21182, N21178, N5681, N13772, N1602);
or OR3 (N21183, N21177, N2462, N7729);
nor NOR3 (N21184, N21183, N20760, N3103);
or OR2 (N21185, N21175, N18317);
not NOT1 (N21186, N21182);
not NOT1 (N21187, N21170);
xor XOR2 (N21188, N21181, N8342);
and AND4 (N21189, N21188, N14119, N10722, N11064);
or OR4 (N21190, N21172, N2855, N16997, N1294);
and AND3 (N21191, N21180, N19323, N13539);
and AND3 (N21192, N21148, N17845, N9216);
or OR4 (N21193, N21159, N2522, N7910, N4692);
xor XOR2 (N21194, N21186, N4087);
xor XOR2 (N21195, N21187, N12176);
xor XOR2 (N21196, N21185, N7667);
nand NAND2 (N21197, N21193, N1144);
nand NAND4 (N21198, N21184, N9931, N14430, N6992);
buf BUF1 (N21199, N21192);
nor NOR3 (N21200, N21195, N4295, N18697);
not NOT1 (N21201, N21199);
nand NAND3 (N21202, N21194, N8254, N10735);
not NOT1 (N21203, N21197);
or OR3 (N21204, N21202, N20599, N20218);
xor XOR2 (N21205, N21200, N16265);
xor XOR2 (N21206, N21191, N7715);
nand NAND4 (N21207, N21189, N18264, N8222, N16991);
or OR2 (N21208, N21201, N8707);
or OR2 (N21209, N21204, N14720);
not NOT1 (N21210, N21179);
nand NAND2 (N21211, N21190, N155);
and AND2 (N21212, N21210, N1361);
buf BUF1 (N21213, N21209);
buf BUF1 (N21214, N21211);
buf BUF1 (N21215, N21196);
xor XOR2 (N21216, N21205, N14609);
nor NOR4 (N21217, N21215, N3371, N7557, N19049);
nor NOR2 (N21218, N21206, N17193);
and AND2 (N21219, N21212, N9826);
buf BUF1 (N21220, N21198);
nand NAND3 (N21221, N21219, N20726, N4552);
and AND3 (N21222, N21217, N16447, N18331);
nor NOR2 (N21223, N21203, N4505);
nor NOR2 (N21224, N21213, N1903);
nor NOR2 (N21225, N21222, N503);
nor NOR2 (N21226, N21214, N1573);
buf BUF1 (N21227, N21216);
not NOT1 (N21228, N21220);
nor NOR4 (N21229, N21208, N15265, N9959, N631);
or OR4 (N21230, N21207, N21210, N13327, N3836);
or OR3 (N21231, N21230, N7247, N12863);
or OR2 (N21232, N21229, N12838);
nand NAND2 (N21233, N21218, N11563);
nand NAND3 (N21234, N21232, N950, N9061);
nand NAND4 (N21235, N21226, N9065, N11282, N3631);
nand NAND2 (N21236, N21231, N14210);
xor XOR2 (N21237, N21233, N931);
nor NOR4 (N21238, N21223, N5109, N10640, N10216);
nor NOR4 (N21239, N21236, N993, N2464, N20129);
buf BUF1 (N21240, N21239);
nand NAND2 (N21241, N21238, N2188);
and AND4 (N21242, N21221, N5316, N7293, N16140);
not NOT1 (N21243, N21227);
nor NOR3 (N21244, N21242, N11098, N2433);
buf BUF1 (N21245, N21234);
nor NOR3 (N21246, N21245, N18370, N18615);
nor NOR2 (N21247, N21246, N7921);
and AND4 (N21248, N21225, N9115, N21242, N11103);
not NOT1 (N21249, N21228);
buf BUF1 (N21250, N21240);
not NOT1 (N21251, N21235);
buf BUF1 (N21252, N21247);
nand NAND2 (N21253, N21251, N18579);
buf BUF1 (N21254, N21241);
or OR4 (N21255, N21252, N10747, N20523, N19321);
nand NAND3 (N21256, N21243, N17019, N20569);
nand NAND3 (N21257, N21249, N6065, N3397);
nor NOR2 (N21258, N21237, N1973);
and AND4 (N21259, N21256, N2816, N11505, N133);
buf BUF1 (N21260, N21244);
or OR3 (N21261, N21258, N7388, N9370);
nor NOR4 (N21262, N21248, N21147, N13379, N10886);
xor XOR2 (N21263, N21255, N13218);
and AND2 (N21264, N21263, N7074);
nand NAND4 (N21265, N21261, N2481, N6368, N14908);
or OR3 (N21266, N21260, N13014, N18683);
xor XOR2 (N21267, N21266, N13788);
or OR3 (N21268, N21259, N20888, N13103);
buf BUF1 (N21269, N21250);
not NOT1 (N21270, N21267);
nor NOR2 (N21271, N21254, N17287);
nand NAND2 (N21272, N21265, N1344);
nor NOR3 (N21273, N21268, N5140, N20931);
not NOT1 (N21274, N21269);
nand NAND2 (N21275, N21273, N20271);
xor XOR2 (N21276, N21262, N9198);
xor XOR2 (N21277, N21257, N142);
nor NOR4 (N21278, N21271, N131, N15374, N2400);
buf BUF1 (N21279, N21270);
or OR3 (N21280, N21275, N5806, N17178);
nor NOR4 (N21281, N21224, N12899, N14113, N20668);
buf BUF1 (N21282, N21280);
xor XOR2 (N21283, N21282, N14065);
or OR4 (N21284, N21279, N12420, N11776, N11285);
nand NAND2 (N21285, N21264, N14399);
not NOT1 (N21286, N21277);
buf BUF1 (N21287, N21281);
nor NOR4 (N21288, N21274, N15065, N13133, N4262);
buf BUF1 (N21289, N21253);
nand NAND2 (N21290, N21289, N17362);
not NOT1 (N21291, N21283);
xor XOR2 (N21292, N21287, N12859);
not NOT1 (N21293, N21291);
buf BUF1 (N21294, N21276);
xor XOR2 (N21295, N21286, N9121);
or OR4 (N21296, N21272, N3006, N12348, N2361);
or OR3 (N21297, N21294, N1751, N1667);
not NOT1 (N21298, N21296);
xor XOR2 (N21299, N21284, N5245);
or OR2 (N21300, N21292, N11635);
nor NOR4 (N21301, N21293, N21098, N18295, N5894);
xor XOR2 (N21302, N21285, N20011);
not NOT1 (N21303, N21295);
not NOT1 (N21304, N21278);
and AND4 (N21305, N21290, N4975, N20336, N15293);
nor NOR3 (N21306, N21299, N11160, N102);
not NOT1 (N21307, N21301);
xor XOR2 (N21308, N21298, N17118);
and AND2 (N21309, N21306, N1718);
and AND2 (N21310, N21297, N6999);
nand NAND2 (N21311, N21309, N1532);
or OR3 (N21312, N21302, N5814, N7200);
buf BUF1 (N21313, N21312);
nand NAND3 (N21314, N21307, N15015, N15675);
not NOT1 (N21315, N21313);
buf BUF1 (N21316, N21314);
or OR2 (N21317, N21308, N7786);
nand NAND3 (N21318, N21317, N16460, N7045);
or OR3 (N21319, N21300, N19969, N11150);
buf BUF1 (N21320, N21305);
not NOT1 (N21321, N21310);
xor XOR2 (N21322, N21303, N4697);
not NOT1 (N21323, N21318);
and AND3 (N21324, N21311, N14988, N8082);
nor NOR2 (N21325, N21304, N10720);
xor XOR2 (N21326, N21323, N10586);
nand NAND3 (N21327, N21321, N7003, N865);
or OR3 (N21328, N21316, N12082, N2820);
nor NOR3 (N21329, N21325, N449, N19544);
xor XOR2 (N21330, N21324, N14997);
nand NAND4 (N21331, N21319, N18677, N6737, N20052);
nand NAND4 (N21332, N21329, N7962, N1000, N12058);
xor XOR2 (N21333, N21332, N18453);
and AND3 (N21334, N21315, N21031, N14058);
buf BUF1 (N21335, N21322);
xor XOR2 (N21336, N21330, N14578);
buf BUF1 (N21337, N21326);
xor XOR2 (N21338, N21333, N1288);
buf BUF1 (N21339, N21338);
nor NOR2 (N21340, N21328, N13651);
and AND4 (N21341, N21327, N5474, N2781, N12017);
nand NAND3 (N21342, N21334, N10757, N4894);
nor NOR2 (N21343, N21336, N7152);
not NOT1 (N21344, N21320);
or OR3 (N21345, N21288, N11696, N9004);
or OR3 (N21346, N21341, N2610, N10115);
and AND2 (N21347, N21331, N11147);
nand NAND4 (N21348, N21337, N18829, N16061, N4139);
xor XOR2 (N21349, N21343, N17071);
not NOT1 (N21350, N21342);
xor XOR2 (N21351, N21346, N8635);
xor XOR2 (N21352, N21340, N7193);
or OR4 (N21353, N21347, N6886, N14527, N3466);
and AND2 (N21354, N21339, N17877);
or OR3 (N21355, N21354, N18, N13602);
nor NOR3 (N21356, N21349, N727, N13432);
xor XOR2 (N21357, N21353, N13802);
not NOT1 (N21358, N21352);
or OR4 (N21359, N21356, N13102, N13527, N2873);
buf BUF1 (N21360, N21348);
not NOT1 (N21361, N21344);
nor NOR2 (N21362, N21361, N106);
nand NAND3 (N21363, N21351, N17918, N14607);
and AND3 (N21364, N21360, N16722, N17804);
or OR2 (N21365, N21335, N833);
buf BUF1 (N21366, N21355);
or OR4 (N21367, N21363, N7185, N15935, N10680);
buf BUF1 (N21368, N21345);
nor NOR2 (N21369, N21368, N8810);
buf BUF1 (N21370, N21364);
not NOT1 (N21371, N21358);
or OR2 (N21372, N21369, N2111);
not NOT1 (N21373, N21357);
or OR4 (N21374, N21359, N14380, N3824, N2683);
or OR3 (N21375, N21365, N4797, N13400);
not NOT1 (N21376, N21370);
and AND4 (N21377, N21376, N8972, N9293, N20608);
not NOT1 (N21378, N21350);
and AND4 (N21379, N21378, N8382, N16920, N21155);
and AND3 (N21380, N21372, N10812, N14705);
xor XOR2 (N21381, N21371, N18591);
xor XOR2 (N21382, N21380, N3289);
and AND4 (N21383, N21366, N20436, N11986, N17795);
or OR3 (N21384, N21373, N9072, N19334);
nand NAND2 (N21385, N21384, N5415);
nand NAND3 (N21386, N21377, N8694, N16565);
nor NOR4 (N21387, N21374, N5938, N4001, N2138);
nor NOR4 (N21388, N21382, N1584, N15264, N5199);
nand NAND4 (N21389, N21388, N13443, N20801, N13993);
not NOT1 (N21390, N21379);
buf BUF1 (N21391, N21390);
xor XOR2 (N21392, N21367, N8821);
not NOT1 (N21393, N21387);
buf BUF1 (N21394, N21393);
or OR4 (N21395, N21391, N11584, N15764, N11323);
nor NOR3 (N21396, N21362, N5143, N15532);
or OR2 (N21397, N21395, N18339);
buf BUF1 (N21398, N21397);
or OR3 (N21399, N21392, N17667, N2952);
nor NOR2 (N21400, N21396, N4602);
buf BUF1 (N21401, N21386);
nor NOR4 (N21402, N21381, N14730, N16818, N12854);
and AND4 (N21403, N21383, N14830, N7329, N4835);
nand NAND4 (N21404, N21398, N12621, N14579, N14819);
not NOT1 (N21405, N21400);
buf BUF1 (N21406, N21375);
or OR2 (N21407, N21394, N9981);
not NOT1 (N21408, N21401);
buf BUF1 (N21409, N21389);
nand NAND2 (N21410, N21404, N16071);
xor XOR2 (N21411, N21409, N16989);
not NOT1 (N21412, N21385);
xor XOR2 (N21413, N21402, N17128);
xor XOR2 (N21414, N21413, N5518);
and AND3 (N21415, N21407, N3975, N3132);
not NOT1 (N21416, N21408);
buf BUF1 (N21417, N21416);
and AND2 (N21418, N21403, N10644);
not NOT1 (N21419, N21405);
nor NOR3 (N21420, N21417, N16119, N11085);
or OR4 (N21421, N21406, N9169, N1025, N10521);
not NOT1 (N21422, N21412);
buf BUF1 (N21423, N21419);
or OR2 (N21424, N21420, N12933);
buf BUF1 (N21425, N21424);
nor NOR3 (N21426, N21422, N11864, N6800);
or OR3 (N21427, N21411, N4217, N18800);
xor XOR2 (N21428, N21423, N13564);
nor NOR4 (N21429, N21414, N19970, N16896, N8395);
or OR2 (N21430, N21410, N7038);
xor XOR2 (N21431, N21429, N3242);
nor NOR3 (N21432, N21431, N1711, N9272);
buf BUF1 (N21433, N21428);
nand NAND3 (N21434, N21425, N12349, N9996);
or OR2 (N21435, N21418, N9742);
and AND3 (N21436, N21426, N11801, N18769);
and AND3 (N21437, N21430, N8183, N3167);
xor XOR2 (N21438, N21437, N2943);
or OR3 (N21439, N21436, N19799, N13840);
buf BUF1 (N21440, N21434);
buf BUF1 (N21441, N21439);
not NOT1 (N21442, N21441);
and AND2 (N21443, N21440, N19131);
and AND3 (N21444, N21421, N1633, N7051);
and AND4 (N21445, N21435, N1737, N14825, N9575);
or OR4 (N21446, N21442, N4324, N51, N7798);
not NOT1 (N21447, N21444);
xor XOR2 (N21448, N21438, N1187);
nor NOR2 (N21449, N21443, N2789);
or OR3 (N21450, N21445, N9158, N10002);
not NOT1 (N21451, N21415);
or OR4 (N21452, N21399, N14013, N7273, N8294);
nor NOR4 (N21453, N21452, N8666, N693, N9587);
and AND2 (N21454, N21433, N6307);
xor XOR2 (N21455, N21446, N16041);
nand NAND2 (N21456, N21450, N18405);
nand NAND4 (N21457, N21456, N9157, N9181, N15379);
not NOT1 (N21458, N21451);
nor NOR3 (N21459, N21449, N7715, N17124);
buf BUF1 (N21460, N21459);
not NOT1 (N21461, N21457);
and AND4 (N21462, N21447, N14155, N20580, N11492);
nand NAND2 (N21463, N21460, N20672);
or OR3 (N21464, N21461, N10725, N2781);
not NOT1 (N21465, N21455);
not NOT1 (N21466, N21454);
nand NAND3 (N21467, N21463, N16358, N12940);
nor NOR2 (N21468, N21427, N2822);
or OR3 (N21469, N21468, N6880, N18350);
and AND3 (N21470, N21458, N10042, N8591);
xor XOR2 (N21471, N21453, N796);
not NOT1 (N21472, N21467);
not NOT1 (N21473, N21470);
buf BUF1 (N21474, N21432);
or OR4 (N21475, N21472, N390, N6052, N18112);
nand NAND4 (N21476, N21465, N3137, N21046, N15372);
buf BUF1 (N21477, N21475);
and AND2 (N21478, N21471, N17367);
nand NAND4 (N21479, N21464, N11438, N900, N165);
nand NAND3 (N21480, N21448, N20026, N12875);
and AND4 (N21481, N21473, N21205, N12678, N6649);
not NOT1 (N21482, N21469);
buf BUF1 (N21483, N21480);
not NOT1 (N21484, N21478);
buf BUF1 (N21485, N21481);
nand NAND2 (N21486, N21485, N6235);
buf BUF1 (N21487, N21482);
not NOT1 (N21488, N21466);
nand NAND2 (N21489, N21479, N7582);
buf BUF1 (N21490, N21476);
and AND4 (N21491, N21462, N5630, N3223, N262);
nand NAND3 (N21492, N21491, N6343, N17631);
xor XOR2 (N21493, N21477, N8801);
nor NOR2 (N21494, N21488, N10399);
or OR4 (N21495, N21494, N12177, N17267, N2256);
xor XOR2 (N21496, N21493, N21191);
and AND4 (N21497, N21490, N6026, N12499, N20219);
nor NOR3 (N21498, N21492, N19895, N18916);
xor XOR2 (N21499, N21484, N18000);
and AND2 (N21500, N21496, N1338);
xor XOR2 (N21501, N21483, N20294);
not NOT1 (N21502, N21489);
not NOT1 (N21503, N21486);
or OR4 (N21504, N21500, N15070, N16268, N20906);
nor NOR4 (N21505, N21501, N17908, N11668, N16751);
buf BUF1 (N21506, N21505);
buf BUF1 (N21507, N21499);
not NOT1 (N21508, N21504);
not NOT1 (N21509, N21507);
nor NOR4 (N21510, N21498, N19750, N21406, N11772);
and AND2 (N21511, N21487, N5773);
xor XOR2 (N21512, N21511, N15290);
nand NAND4 (N21513, N21474, N20195, N18915, N12692);
nor NOR2 (N21514, N21503, N9328);
nor NOR2 (N21515, N21508, N6959);
or OR3 (N21516, N21514, N17321, N5377);
nor NOR3 (N21517, N21497, N3261, N17383);
or OR2 (N21518, N21495, N4213);
nor NOR2 (N21519, N21512, N10764);
nand NAND3 (N21520, N21510, N14677, N16315);
nor NOR3 (N21521, N21502, N16665, N2987);
and AND2 (N21522, N21518, N17617);
nand NAND2 (N21523, N21506, N19412);
buf BUF1 (N21524, N21520);
or OR3 (N21525, N21523, N18415, N12737);
not NOT1 (N21526, N21521);
and AND2 (N21527, N21517, N9932);
nand NAND3 (N21528, N21527, N13969, N5913);
nand NAND3 (N21529, N21528, N5747, N6340);
or OR3 (N21530, N21519, N5164, N6918);
not NOT1 (N21531, N21524);
nor NOR3 (N21532, N21525, N7300, N12029);
nor NOR2 (N21533, N21530, N12077);
or OR2 (N21534, N21529, N1894);
not NOT1 (N21535, N21509);
or OR2 (N21536, N21516, N10831);
not NOT1 (N21537, N21515);
xor XOR2 (N21538, N21534, N11468);
not NOT1 (N21539, N21533);
nor NOR4 (N21540, N21536, N1279, N2884, N12978);
or OR3 (N21541, N21535, N10873, N10098);
nand NAND2 (N21542, N21541, N7242);
or OR4 (N21543, N21522, N15393, N8073, N12227);
xor XOR2 (N21544, N21542, N306);
buf BUF1 (N21545, N21544);
buf BUF1 (N21546, N21532);
not NOT1 (N21547, N21539);
and AND4 (N21548, N21513, N18822, N1086, N12413);
or OR2 (N21549, N21538, N8796);
not NOT1 (N21550, N21531);
not NOT1 (N21551, N21549);
xor XOR2 (N21552, N21545, N3249);
and AND4 (N21553, N21550, N10010, N4999, N3932);
xor XOR2 (N21554, N21551, N4235);
buf BUF1 (N21555, N21537);
xor XOR2 (N21556, N21546, N12631);
and AND4 (N21557, N21552, N3374, N20025, N20154);
not NOT1 (N21558, N21553);
xor XOR2 (N21559, N21554, N3934);
nand NAND3 (N21560, N21559, N15969, N18441);
nor NOR4 (N21561, N21555, N3968, N7207, N15882);
not NOT1 (N21562, N21543);
nand NAND3 (N21563, N21557, N20031, N11691);
xor XOR2 (N21564, N21526, N14429);
buf BUF1 (N21565, N21547);
not NOT1 (N21566, N21540);
nand NAND3 (N21567, N21558, N17215, N10926);
and AND2 (N21568, N21566, N1957);
xor XOR2 (N21569, N21560, N5994);
not NOT1 (N21570, N21563);
buf BUF1 (N21571, N21562);
and AND4 (N21572, N21567, N16659, N10216, N16899);
nor NOR2 (N21573, N21556, N12059);
nor NOR3 (N21574, N21561, N3726, N9390);
or OR4 (N21575, N21570, N2028, N18439, N16025);
nand NAND3 (N21576, N21571, N21220, N353);
nor NOR2 (N21577, N21574, N19911);
or OR3 (N21578, N21575, N990, N15015);
buf BUF1 (N21579, N21573);
and AND3 (N21580, N21577, N12727, N18608);
not NOT1 (N21581, N21572);
nand NAND2 (N21582, N21564, N10215);
not NOT1 (N21583, N21568);
buf BUF1 (N21584, N21569);
xor XOR2 (N21585, N21580, N20118);
buf BUF1 (N21586, N21565);
and AND2 (N21587, N21579, N3417);
and AND2 (N21588, N21584, N16926);
nor NOR3 (N21589, N21548, N62, N4533);
not NOT1 (N21590, N21582);
xor XOR2 (N21591, N21578, N17815);
nor NOR2 (N21592, N21586, N16554);
nand NAND2 (N21593, N21588, N16448);
and AND3 (N21594, N21593, N1425, N17517);
nor NOR2 (N21595, N21594, N11751);
xor XOR2 (N21596, N21591, N1993);
xor XOR2 (N21597, N21585, N20480);
xor XOR2 (N21598, N21590, N4677);
and AND3 (N21599, N21581, N20389, N11948);
xor XOR2 (N21600, N21583, N5062);
buf BUF1 (N21601, N21596);
or OR4 (N21602, N21597, N14692, N16309, N5567);
xor XOR2 (N21603, N21599, N1464);
buf BUF1 (N21604, N21602);
and AND4 (N21605, N21587, N11048, N18284, N668);
xor XOR2 (N21606, N21603, N1405);
buf BUF1 (N21607, N21595);
xor XOR2 (N21608, N21576, N1025);
nor NOR4 (N21609, N21601, N5152, N17585, N15208);
buf BUF1 (N21610, N21592);
nand NAND4 (N21611, N21610, N5393, N15800, N3091);
buf BUF1 (N21612, N21605);
nor NOR2 (N21613, N21607, N9995);
xor XOR2 (N21614, N21604, N16593);
and AND4 (N21615, N21611, N20372, N750, N7289);
not NOT1 (N21616, N21609);
nor NOR2 (N21617, N21589, N21072);
nand NAND3 (N21618, N21617, N1813, N10002);
nor NOR4 (N21619, N21613, N10453, N10540, N20412);
nor NOR4 (N21620, N21616, N7226, N10681, N4713);
nor NOR3 (N21621, N21619, N7158, N5256);
not NOT1 (N21622, N21612);
nand NAND2 (N21623, N21615, N13345);
nand NAND2 (N21624, N21623, N811);
xor XOR2 (N21625, N21606, N18417);
nor NOR4 (N21626, N21618, N1563, N14817, N19812);
not NOT1 (N21627, N21624);
xor XOR2 (N21628, N21598, N6911);
buf BUF1 (N21629, N21608);
buf BUF1 (N21630, N21622);
nand NAND2 (N21631, N21614, N4222);
or OR4 (N21632, N21600, N14350, N12354, N18853);
buf BUF1 (N21633, N21631);
nor NOR2 (N21634, N21629, N1514);
xor XOR2 (N21635, N21620, N19570);
and AND4 (N21636, N21625, N6894, N14402, N11319);
or OR3 (N21637, N21636, N13127, N6523);
xor XOR2 (N21638, N21630, N3278);
buf BUF1 (N21639, N21635);
not NOT1 (N21640, N21628);
and AND3 (N21641, N21634, N4836, N1619);
nand NAND4 (N21642, N21626, N4769, N5616, N13224);
not NOT1 (N21643, N21627);
nor NOR4 (N21644, N21638, N2291, N13789, N13724);
not NOT1 (N21645, N21637);
nand NAND3 (N21646, N21621, N1617, N12361);
nor NOR4 (N21647, N21643, N8714, N9739, N18108);
buf BUF1 (N21648, N21632);
nand NAND2 (N21649, N21639, N14761);
or OR4 (N21650, N21642, N1759, N13542, N8932);
nand NAND3 (N21651, N21650, N14596, N21103);
nor NOR2 (N21652, N21645, N17118);
nor NOR4 (N21653, N21640, N929, N21094, N17477);
and AND2 (N21654, N21648, N11574);
nand NAND2 (N21655, N21644, N13644);
not NOT1 (N21656, N21649);
buf BUF1 (N21657, N21656);
nor NOR4 (N21658, N21651, N21039, N7773, N3154);
nand NAND2 (N21659, N21647, N21528);
or OR3 (N21660, N21657, N9910, N12194);
not NOT1 (N21661, N21653);
nor NOR2 (N21662, N21641, N1156);
or OR3 (N21663, N21652, N3991, N16401);
nor NOR3 (N21664, N21654, N558, N12980);
or OR2 (N21665, N21662, N1732);
nor NOR3 (N21666, N21646, N14916, N6291);
or OR3 (N21667, N21666, N6418, N11910);
and AND2 (N21668, N21655, N13728);
or OR3 (N21669, N21659, N5173, N15167);
not NOT1 (N21670, N21667);
xor XOR2 (N21671, N21658, N11144);
and AND3 (N21672, N21663, N18141, N12569);
nor NOR3 (N21673, N21668, N20924, N12471);
nand NAND4 (N21674, N21671, N9181, N2357, N18591);
nand NAND4 (N21675, N21670, N7182, N18168, N17704);
or OR2 (N21676, N21664, N8742);
nor NOR3 (N21677, N21673, N17922, N17515);
nand NAND3 (N21678, N21660, N10181, N13033);
not NOT1 (N21679, N21661);
buf BUF1 (N21680, N21665);
and AND4 (N21681, N21678, N6610, N19214, N3153);
or OR4 (N21682, N21669, N13144, N626, N18717);
buf BUF1 (N21683, N21633);
nand NAND2 (N21684, N21675, N12961);
and AND2 (N21685, N21683, N7439);
nor NOR2 (N21686, N21685, N19670);
buf BUF1 (N21687, N21680);
nand NAND3 (N21688, N21686, N4933, N4877);
xor XOR2 (N21689, N21674, N135);
buf BUF1 (N21690, N21679);
nand NAND3 (N21691, N21687, N18295, N12696);
and AND2 (N21692, N21689, N21600);
nand NAND3 (N21693, N21690, N7657, N21536);
buf BUF1 (N21694, N21681);
not NOT1 (N21695, N21684);
xor XOR2 (N21696, N21672, N17006);
nor NOR3 (N21697, N21688, N1817, N13103);
xor XOR2 (N21698, N21696, N17835);
nand NAND4 (N21699, N21695, N3098, N180, N15415);
not NOT1 (N21700, N21682);
and AND4 (N21701, N21697, N2202, N13922, N17249);
not NOT1 (N21702, N21701);
and AND3 (N21703, N21693, N18690, N17881);
nand NAND2 (N21704, N21676, N3846);
and AND3 (N21705, N21694, N9639, N16268);
nand NAND2 (N21706, N21700, N4635);
not NOT1 (N21707, N21702);
not NOT1 (N21708, N21705);
or OR4 (N21709, N21708, N2923, N14600, N19411);
and AND2 (N21710, N21704, N13241);
not NOT1 (N21711, N21709);
nand NAND3 (N21712, N21703, N6708, N11812);
and AND3 (N21713, N21710, N293, N17663);
nor NOR3 (N21714, N21692, N16230, N21150);
and AND4 (N21715, N21707, N1475, N15222, N10311);
buf BUF1 (N21716, N21712);
nand NAND3 (N21717, N21691, N21232, N16654);
nand NAND2 (N21718, N21713, N20862);
and AND4 (N21719, N21718, N21105, N20327, N1430);
or OR2 (N21720, N21716, N7563);
and AND4 (N21721, N21706, N14836, N3078, N6882);
nor NOR2 (N21722, N21715, N5167);
and AND2 (N21723, N21721, N14238);
xor XOR2 (N21724, N21699, N12858);
xor XOR2 (N21725, N21717, N11286);
and AND2 (N21726, N21711, N21230);
or OR2 (N21727, N21725, N20110);
and AND2 (N21728, N21726, N2736);
buf BUF1 (N21729, N21723);
or OR4 (N21730, N21719, N8042, N3849, N17121);
nand NAND4 (N21731, N21728, N15229, N807, N11376);
not NOT1 (N21732, N21727);
not NOT1 (N21733, N21732);
nor NOR3 (N21734, N21722, N15851, N4011);
not NOT1 (N21735, N21729);
not NOT1 (N21736, N21730);
nand NAND2 (N21737, N21735, N21048);
buf BUF1 (N21738, N21724);
nor NOR3 (N21739, N21720, N2813, N5324);
buf BUF1 (N21740, N21734);
nor NOR2 (N21741, N21677, N1948);
or OR3 (N21742, N21714, N4522, N4659);
not NOT1 (N21743, N21737);
nand NAND4 (N21744, N21741, N9077, N3819, N934);
nor NOR4 (N21745, N21740, N8210, N18850, N7910);
not NOT1 (N21746, N21745);
nand NAND4 (N21747, N21746, N1062, N19181, N18888);
not NOT1 (N21748, N21742);
and AND4 (N21749, N21733, N6821, N9955, N18294);
xor XOR2 (N21750, N21739, N1195);
and AND4 (N21751, N21750, N5758, N21249, N9080);
and AND4 (N21752, N21736, N13950, N1318, N19569);
not NOT1 (N21753, N21738);
nand NAND4 (N21754, N21748, N14755, N5035, N14345);
buf BUF1 (N21755, N21698);
buf BUF1 (N21756, N21731);
or OR3 (N21757, N21751, N18781, N7562);
and AND2 (N21758, N21754, N10956);
buf BUF1 (N21759, N21755);
buf BUF1 (N21760, N21744);
nand NAND2 (N21761, N21749, N10365);
or OR4 (N21762, N21756, N17888, N10415, N9127);
not NOT1 (N21763, N21752);
xor XOR2 (N21764, N21753, N12686);
and AND4 (N21765, N21762, N3571, N20721, N12969);
xor XOR2 (N21766, N21761, N9301);
nand NAND4 (N21767, N21743, N423, N8588, N2283);
buf BUF1 (N21768, N21759);
xor XOR2 (N21769, N21763, N16991);
buf BUF1 (N21770, N21769);
buf BUF1 (N21771, N21757);
nand NAND3 (N21772, N21768, N15832, N17676);
buf BUF1 (N21773, N21760);
or OR3 (N21774, N21747, N21190, N2959);
buf BUF1 (N21775, N21773);
not NOT1 (N21776, N21764);
nand NAND2 (N21777, N21765, N20021);
buf BUF1 (N21778, N21777);
buf BUF1 (N21779, N21774);
and AND2 (N21780, N21776, N5951);
or OR2 (N21781, N21775, N17358);
buf BUF1 (N21782, N21771);
xor XOR2 (N21783, N21778, N2408);
nor NOR3 (N21784, N21779, N8346, N710);
not NOT1 (N21785, N21766);
and AND3 (N21786, N21772, N35, N19718);
xor XOR2 (N21787, N21785, N4019);
not NOT1 (N21788, N21787);
buf BUF1 (N21789, N21780);
and AND3 (N21790, N21758, N10333, N7800);
buf BUF1 (N21791, N21784);
buf BUF1 (N21792, N21786);
buf BUF1 (N21793, N21782);
or OR3 (N21794, N21793, N1364, N3346);
nand NAND2 (N21795, N21770, N18814);
or OR2 (N21796, N21791, N772);
not NOT1 (N21797, N21788);
nor NOR3 (N21798, N21796, N669, N8291);
nand NAND2 (N21799, N21797, N19230);
not NOT1 (N21800, N21789);
nand NAND4 (N21801, N21783, N17610, N7357, N8466);
buf BUF1 (N21802, N21781);
nand NAND3 (N21803, N21801, N2756, N14862);
xor XOR2 (N21804, N21792, N18064);
nand NAND2 (N21805, N21798, N16723);
or OR2 (N21806, N21799, N8068);
nor NOR4 (N21807, N21803, N17740, N16400, N20011);
and AND4 (N21808, N21790, N18142, N10988, N2793);
xor XOR2 (N21809, N21807, N6288);
xor XOR2 (N21810, N21802, N21391);
xor XOR2 (N21811, N21767, N9953);
and AND3 (N21812, N21794, N4458, N11108);
buf BUF1 (N21813, N21811);
not NOT1 (N21814, N21795);
and AND3 (N21815, N21804, N19480, N15859);
or OR3 (N21816, N21812, N16932, N247);
not NOT1 (N21817, N21808);
and AND2 (N21818, N21800, N6588);
xor XOR2 (N21819, N21817, N5644);
or OR2 (N21820, N21805, N18670);
and AND2 (N21821, N21818, N18953);
xor XOR2 (N21822, N21821, N9428);
xor XOR2 (N21823, N21819, N2410);
buf BUF1 (N21824, N21806);
xor XOR2 (N21825, N21822, N13708);
nor NOR4 (N21826, N21814, N16114, N21652, N5740);
not NOT1 (N21827, N21813);
xor XOR2 (N21828, N21824, N17728);
nand NAND3 (N21829, N21815, N4365, N15676);
nand NAND3 (N21830, N21828, N19071, N19720);
or OR4 (N21831, N21829, N13984, N21230, N4065);
nor NOR4 (N21832, N21827, N16411, N17571, N2161);
xor XOR2 (N21833, N21831, N15160);
not NOT1 (N21834, N21809);
xor XOR2 (N21835, N21834, N13777);
and AND2 (N21836, N21835, N13089);
xor XOR2 (N21837, N21830, N19766);
not NOT1 (N21838, N21832);
nand NAND3 (N21839, N21837, N18919, N9968);
nand NAND3 (N21840, N21836, N18164, N946);
and AND4 (N21841, N21838, N12926, N17306, N10294);
nand NAND3 (N21842, N21839, N17188, N21468);
xor XOR2 (N21843, N21816, N8838);
not NOT1 (N21844, N21820);
and AND4 (N21845, N21823, N8784, N5165, N3680);
nor NOR3 (N21846, N21844, N5570, N17158);
xor XOR2 (N21847, N21846, N16136);
nand NAND2 (N21848, N21833, N10045);
or OR4 (N21849, N21847, N16609, N17943, N5684);
and AND3 (N21850, N21843, N12870, N18031);
buf BUF1 (N21851, N21840);
nand NAND3 (N21852, N21825, N9728, N15330);
not NOT1 (N21853, N21842);
nand NAND3 (N21854, N21851, N12075, N17624);
not NOT1 (N21855, N21841);
nand NAND2 (N21856, N21853, N3297);
buf BUF1 (N21857, N21849);
xor XOR2 (N21858, N21845, N19552);
not NOT1 (N21859, N21850);
not NOT1 (N21860, N21856);
and AND2 (N21861, N21857, N16144);
not NOT1 (N21862, N21855);
nand NAND3 (N21863, N21859, N20576, N19866);
nor NOR3 (N21864, N21852, N21220, N672);
and AND4 (N21865, N21861, N15999, N19335, N16513);
and AND4 (N21866, N21865, N16518, N1378, N10917);
buf BUF1 (N21867, N21848);
xor XOR2 (N21868, N21826, N2378);
nor NOR3 (N21869, N21862, N14001, N15003);
not NOT1 (N21870, N21866);
and AND3 (N21871, N21868, N16696, N7113);
buf BUF1 (N21872, N21871);
and AND2 (N21873, N21854, N1521);
not NOT1 (N21874, N21869);
not NOT1 (N21875, N21860);
and AND3 (N21876, N21863, N18500, N15975);
nor NOR4 (N21877, N21858, N2005, N13413, N19251);
nand NAND2 (N21878, N21877, N4782);
xor XOR2 (N21879, N21810, N18619);
nor NOR4 (N21880, N21872, N8866, N18571, N11427);
nor NOR2 (N21881, N21867, N17949);
nor NOR3 (N21882, N21875, N1678, N21880);
or OR4 (N21883, N12301, N14953, N312, N10430);
xor XOR2 (N21884, N21864, N4956);
or OR2 (N21885, N21870, N1386);
nand NAND2 (N21886, N21882, N3339);
buf BUF1 (N21887, N21874);
xor XOR2 (N21888, N21887, N5486);
xor XOR2 (N21889, N21879, N6236);
not NOT1 (N21890, N21881);
xor XOR2 (N21891, N21883, N12040);
buf BUF1 (N21892, N21891);
xor XOR2 (N21893, N21885, N15506);
not NOT1 (N21894, N21876);
buf BUF1 (N21895, N21878);
nor NOR3 (N21896, N21888, N14073, N19152);
buf BUF1 (N21897, N21889);
or OR2 (N21898, N21897, N16008);
not NOT1 (N21899, N21893);
or OR3 (N21900, N21892, N9170, N14734);
or OR3 (N21901, N21899, N699, N8140);
and AND3 (N21902, N21896, N11943, N12493);
not NOT1 (N21903, N21895);
nand NAND3 (N21904, N21884, N14968, N21616);
xor XOR2 (N21905, N21901, N13392);
buf BUF1 (N21906, N21905);
buf BUF1 (N21907, N21894);
buf BUF1 (N21908, N21890);
not NOT1 (N21909, N21907);
not NOT1 (N21910, N21873);
buf BUF1 (N21911, N21903);
xor XOR2 (N21912, N21908, N12009);
not NOT1 (N21913, N21906);
or OR2 (N21914, N21886, N20238);
nor NOR4 (N21915, N21912, N5846, N6743, N18813);
or OR2 (N21916, N21904, N1850);
or OR4 (N21917, N21900, N15236, N9318, N20693);
xor XOR2 (N21918, N21913, N706);
or OR4 (N21919, N21915, N8194, N17124, N10039);
and AND2 (N21920, N21916, N3965);
and AND4 (N21921, N21918, N1529, N18990, N4299);
xor XOR2 (N21922, N21921, N5890);
nor NOR4 (N21923, N21902, N3762, N16985, N14859);
nor NOR2 (N21924, N21909, N4455);
buf BUF1 (N21925, N21923);
and AND4 (N21926, N21925, N19057, N16341, N10394);
nand NAND3 (N21927, N21914, N12970, N20278);
not NOT1 (N21928, N21924);
or OR2 (N21929, N21928, N17806);
nor NOR4 (N21930, N21929, N19468, N11971, N11732);
xor XOR2 (N21931, N21911, N7751);
xor XOR2 (N21932, N21927, N6405);
buf BUF1 (N21933, N21917);
not NOT1 (N21934, N21932);
nand NAND4 (N21935, N21898, N12761, N18379, N8081);
or OR4 (N21936, N21933, N13845, N21632, N672);
xor XOR2 (N21937, N21930, N16746);
or OR4 (N21938, N21920, N17334, N2788, N4184);
or OR3 (N21939, N21931, N10668, N2446);
not NOT1 (N21940, N21910);
nand NAND3 (N21941, N21922, N16674, N8210);
nand NAND3 (N21942, N21939, N9353, N16740);
buf BUF1 (N21943, N21937);
and AND3 (N21944, N21942, N21448, N21672);
buf BUF1 (N21945, N21941);
and AND2 (N21946, N21936, N12292);
not NOT1 (N21947, N21926);
and AND3 (N21948, N21945, N16097, N13546);
not NOT1 (N21949, N21934);
or OR2 (N21950, N21944, N15337);
buf BUF1 (N21951, N21940);
buf BUF1 (N21952, N21949);
not NOT1 (N21953, N21935);
nor NOR2 (N21954, N21950, N840);
not NOT1 (N21955, N21947);
xor XOR2 (N21956, N21946, N11522);
not NOT1 (N21957, N21943);
xor XOR2 (N21958, N21948, N14562);
not NOT1 (N21959, N21952);
not NOT1 (N21960, N21955);
buf BUF1 (N21961, N21919);
nand NAND2 (N21962, N21961, N14774);
xor XOR2 (N21963, N21951, N15421);
nand NAND2 (N21964, N21957, N2703);
not NOT1 (N21965, N21959);
buf BUF1 (N21966, N21953);
not NOT1 (N21967, N21954);
buf BUF1 (N21968, N21966);
nand NAND3 (N21969, N21958, N787, N17124);
nor NOR2 (N21970, N21963, N5523);
nand NAND4 (N21971, N21960, N13874, N17218, N10307);
or OR3 (N21972, N21967, N17963, N13357);
not NOT1 (N21973, N21964);
xor XOR2 (N21974, N21973, N7628);
or OR2 (N21975, N21962, N8207);
or OR2 (N21976, N21968, N15111);
nand NAND2 (N21977, N21938, N10824);
xor XOR2 (N21978, N21976, N12898);
buf BUF1 (N21979, N21956);
buf BUF1 (N21980, N21975);
nor NOR3 (N21981, N21979, N10200, N19760);
nand NAND2 (N21982, N21981, N15158);
or OR3 (N21983, N21977, N18067, N15945);
xor XOR2 (N21984, N21974, N11833);
nor NOR4 (N21985, N21982, N15891, N20770, N9673);
xor XOR2 (N21986, N21980, N8377);
not NOT1 (N21987, N21970);
nand NAND2 (N21988, N21985, N9126);
not NOT1 (N21989, N21971);
xor XOR2 (N21990, N21969, N15200);
xor XOR2 (N21991, N21988, N1620);
nor NOR4 (N21992, N21989, N8433, N371, N10474);
xor XOR2 (N21993, N21983, N8311);
and AND2 (N21994, N21987, N20699);
not NOT1 (N21995, N21991);
or OR2 (N21996, N21995, N11658);
buf BUF1 (N21997, N21990);
not NOT1 (N21998, N21984);
not NOT1 (N21999, N21978);
not NOT1 (N22000, N21972);
nor NOR3 (N22001, N21998, N14712, N4045);
nor NOR3 (N22002, N21997, N3094, N11796);
nor NOR4 (N22003, N22000, N6284, N2463, N1708);
not NOT1 (N22004, N21996);
xor XOR2 (N22005, N21999, N17632);
nand NAND4 (N22006, N22004, N5148, N17561, N16200);
xor XOR2 (N22007, N21965, N14812);
nor NOR2 (N22008, N22007, N11321);
or OR4 (N22009, N22006, N1024, N13363, N2492);
buf BUF1 (N22010, N21986);
buf BUF1 (N22011, N21992);
nor NOR4 (N22012, N22002, N5944, N11318, N4519);
or OR2 (N22013, N22005, N21725);
buf BUF1 (N22014, N22008);
and AND4 (N22015, N22013, N21362, N17879, N17397);
and AND2 (N22016, N22011, N4766);
and AND3 (N22017, N22012, N3551, N13175);
not NOT1 (N22018, N22001);
not NOT1 (N22019, N22009);
nor NOR2 (N22020, N22003, N8154);
xor XOR2 (N22021, N22015, N547);
xor XOR2 (N22022, N21994, N565);
not NOT1 (N22023, N22017);
xor XOR2 (N22024, N22022, N11857);
nor NOR4 (N22025, N22021, N483, N12395, N13155);
or OR4 (N22026, N22023, N5264, N2983, N21716);
and AND2 (N22027, N22024, N13673);
not NOT1 (N22028, N22026);
buf BUF1 (N22029, N22020);
nand NAND3 (N22030, N22014, N3275, N19591);
xor XOR2 (N22031, N22019, N19079);
and AND2 (N22032, N22027, N6478);
not NOT1 (N22033, N22028);
and AND3 (N22034, N22031, N106, N19746);
or OR2 (N22035, N22029, N5122);
nand NAND2 (N22036, N22025, N10611);
nand NAND2 (N22037, N22018, N14956);
not NOT1 (N22038, N22035);
buf BUF1 (N22039, N21993);
xor XOR2 (N22040, N22037, N5210);
or OR4 (N22041, N22038, N8479, N9850, N5222);
nor NOR4 (N22042, N22030, N2574, N15636, N280);
or OR2 (N22043, N22040, N6671);
or OR2 (N22044, N22042, N9525);
xor XOR2 (N22045, N22034, N13300);
nor NOR3 (N22046, N22044, N5745, N11831);
not NOT1 (N22047, N22036);
nor NOR3 (N22048, N22043, N1952, N8354);
nand NAND4 (N22049, N22041, N8324, N1276, N1655);
not NOT1 (N22050, N22045);
or OR3 (N22051, N22032, N9294, N7181);
buf BUF1 (N22052, N22046);
not NOT1 (N22053, N22048);
or OR4 (N22054, N22039, N17935, N18191, N1588);
and AND3 (N22055, N22049, N6453, N11222);
not NOT1 (N22056, N22016);
nand NAND2 (N22057, N22056, N10810);
buf BUF1 (N22058, N22010);
nor NOR4 (N22059, N22057, N16988, N14591, N16848);
not NOT1 (N22060, N22051);
xor XOR2 (N22061, N22047, N1466);
xor XOR2 (N22062, N22033, N3751);
not NOT1 (N22063, N22062);
nor NOR2 (N22064, N22063, N3514);
and AND3 (N22065, N22059, N2333, N6683);
xor XOR2 (N22066, N22065, N5761);
and AND3 (N22067, N22058, N475, N13489);
xor XOR2 (N22068, N22060, N14743);
buf BUF1 (N22069, N22067);
buf BUF1 (N22070, N22066);
not NOT1 (N22071, N22053);
not NOT1 (N22072, N22069);
or OR2 (N22073, N22072, N11303);
buf BUF1 (N22074, N22073);
buf BUF1 (N22075, N22064);
or OR2 (N22076, N22052, N20418);
not NOT1 (N22077, N22071);
buf BUF1 (N22078, N22075);
xor XOR2 (N22079, N22055, N1733);
or OR4 (N22080, N22077, N13368, N3832, N13317);
nand NAND3 (N22081, N22050, N9154, N17173);
or OR4 (N22082, N22080, N21495, N17764, N15262);
nand NAND3 (N22083, N22054, N15148, N17722);
buf BUF1 (N22084, N22070);
xor XOR2 (N22085, N22081, N8568);
xor XOR2 (N22086, N22079, N2514);
nor NOR2 (N22087, N22074, N5567);
nand NAND4 (N22088, N22061, N20570, N6746, N20992);
or OR2 (N22089, N22082, N8010);
buf BUF1 (N22090, N22089);
nor NOR3 (N22091, N22078, N16826, N11734);
xor XOR2 (N22092, N22083, N6023);
nand NAND4 (N22093, N22084, N10972, N13479, N11730);
not NOT1 (N22094, N22093);
nand NAND3 (N22095, N22087, N17030, N13539);
buf BUF1 (N22096, N22088);
xor XOR2 (N22097, N22092, N20916);
and AND2 (N22098, N22068, N6509);
buf BUF1 (N22099, N22085);
buf BUF1 (N22100, N22094);
nor NOR4 (N22101, N22096, N4389, N13427, N14716);
or OR4 (N22102, N22076, N8918, N7284, N17848);
xor XOR2 (N22103, N22098, N1206);
and AND4 (N22104, N22100, N11450, N18044, N13141);
nor NOR3 (N22105, N22103, N4396, N7162);
and AND4 (N22106, N22095, N17710, N14130, N19628);
nand NAND4 (N22107, N22091, N8579, N7115, N8682);
or OR2 (N22108, N22101, N10066);
and AND2 (N22109, N22086, N9687);
not NOT1 (N22110, N22102);
nor NOR2 (N22111, N22104, N21421);
nand NAND4 (N22112, N22110, N3844, N5792, N15893);
xor XOR2 (N22113, N22105, N12104);
not NOT1 (N22114, N22108);
nor NOR4 (N22115, N22090, N11751, N11223, N14754);
not NOT1 (N22116, N22115);
or OR3 (N22117, N22111, N21766, N16996);
xor XOR2 (N22118, N22107, N9060);
and AND3 (N22119, N22109, N20208, N16256);
nand NAND4 (N22120, N22106, N10667, N9985, N11171);
nand NAND2 (N22121, N22097, N811);
nand NAND4 (N22122, N22119, N8276, N18822, N19967);
xor XOR2 (N22123, N22122, N11978);
and AND3 (N22124, N22117, N3916, N7593);
nand NAND4 (N22125, N22121, N1047, N3358, N16225);
and AND4 (N22126, N22120, N605, N7684, N19942);
not NOT1 (N22127, N22123);
buf BUF1 (N22128, N22126);
not NOT1 (N22129, N22113);
or OR3 (N22130, N22116, N15727, N3246);
nand NAND4 (N22131, N22114, N16803, N11884, N2246);
and AND4 (N22132, N22118, N21243, N19587, N13405);
or OR2 (N22133, N22125, N6963);
buf BUF1 (N22134, N22124);
nor NOR2 (N22135, N22130, N19347);
xor XOR2 (N22136, N22128, N20379);
or OR4 (N22137, N22133, N15897, N21676, N13579);
nor NOR2 (N22138, N22136, N984);
buf BUF1 (N22139, N22137);
and AND4 (N22140, N22127, N15485, N21388, N2036);
xor XOR2 (N22141, N22132, N22083);
and AND2 (N22142, N22139, N16270);
nand NAND2 (N22143, N22129, N20659);
nand NAND3 (N22144, N22141, N6838, N11542);
and AND2 (N22145, N22138, N13452);
or OR4 (N22146, N22135, N8549, N8505, N7018);
not NOT1 (N22147, N22131);
nor NOR4 (N22148, N22099, N10987, N19935, N19712);
buf BUF1 (N22149, N22143);
xor XOR2 (N22150, N22149, N950);
xor XOR2 (N22151, N22145, N547);
buf BUF1 (N22152, N22140);
buf BUF1 (N22153, N22147);
nor NOR3 (N22154, N22153, N16527, N7901);
xor XOR2 (N22155, N22151, N8918);
and AND4 (N22156, N22148, N16657, N10660, N8545);
and AND2 (N22157, N22155, N7769);
buf BUF1 (N22158, N22156);
or OR2 (N22159, N22112, N8641);
xor XOR2 (N22160, N22134, N15053);
and AND3 (N22161, N22150, N15643, N14769);
and AND4 (N22162, N22146, N20604, N4056, N21401);
xor XOR2 (N22163, N22157, N11676);
buf BUF1 (N22164, N22162);
or OR4 (N22165, N22158, N8751, N9296, N10459);
nand NAND3 (N22166, N22165, N10321, N11588);
xor XOR2 (N22167, N22160, N12097);
buf BUF1 (N22168, N22161);
nor NOR4 (N22169, N22167, N21450, N18015, N19798);
not NOT1 (N22170, N22166);
nand NAND4 (N22171, N22169, N3772, N1065, N9936);
not NOT1 (N22172, N22171);
nor NOR2 (N22173, N22164, N17343);
not NOT1 (N22174, N22170);
buf BUF1 (N22175, N22154);
and AND2 (N22176, N22144, N19263);
nor NOR3 (N22177, N22173, N18514, N6038);
not NOT1 (N22178, N22176);
buf BUF1 (N22179, N22159);
buf BUF1 (N22180, N22172);
xor XOR2 (N22181, N22174, N10344);
not NOT1 (N22182, N22179);
buf BUF1 (N22183, N22168);
buf BUF1 (N22184, N22175);
xor XOR2 (N22185, N22184, N1632);
or OR3 (N22186, N22182, N2027, N11933);
xor XOR2 (N22187, N22181, N5772);
buf BUF1 (N22188, N22152);
xor XOR2 (N22189, N22177, N13373);
nand NAND4 (N22190, N22178, N9461, N7201, N8987);
and AND2 (N22191, N22183, N16686);
and AND3 (N22192, N22190, N18927, N20948);
nor NOR3 (N22193, N22180, N21541, N7322);
xor XOR2 (N22194, N22163, N19778);
or OR2 (N22195, N22189, N20692);
or OR3 (N22196, N22194, N3466, N13016);
or OR4 (N22197, N22188, N9192, N6995, N4069);
not NOT1 (N22198, N22197);
not NOT1 (N22199, N22198);
nand NAND3 (N22200, N22142, N9279, N8332);
and AND3 (N22201, N22191, N10497, N22147);
nand NAND4 (N22202, N22201, N5682, N2732, N13013);
xor XOR2 (N22203, N22200, N3866);
buf BUF1 (N22204, N22187);
nor NOR4 (N22205, N22203, N13980, N21649, N18865);
xor XOR2 (N22206, N22192, N16907);
and AND3 (N22207, N22204, N10314, N7470);
xor XOR2 (N22208, N22196, N15557);
xor XOR2 (N22209, N22199, N795);
not NOT1 (N22210, N22208);
nor NOR4 (N22211, N22210, N15092, N7113, N11042);
not NOT1 (N22212, N22205);
and AND2 (N22213, N22185, N11180);
nand NAND4 (N22214, N22207, N7565, N3934, N18595);
xor XOR2 (N22215, N22213, N2086);
nor NOR4 (N22216, N22209, N11690, N16022, N16247);
xor XOR2 (N22217, N22214, N5958);
and AND3 (N22218, N22212, N10722, N16879);
buf BUF1 (N22219, N22206);
xor XOR2 (N22220, N22215, N966);
buf BUF1 (N22221, N22220);
nor NOR2 (N22222, N22218, N10870);
not NOT1 (N22223, N22217);
nand NAND3 (N22224, N22195, N8321, N15909);
and AND3 (N22225, N22216, N10401, N9453);
xor XOR2 (N22226, N22211, N1788);
and AND4 (N22227, N22223, N10153, N9115, N12226);
not NOT1 (N22228, N22227);
xor XOR2 (N22229, N22219, N12104);
nand NAND3 (N22230, N22186, N18151, N2324);
nor NOR2 (N22231, N22229, N17471);
nand NAND3 (N22232, N22193, N1936, N11439);
not NOT1 (N22233, N22226);
and AND3 (N22234, N22232, N2912, N19325);
and AND3 (N22235, N22225, N17070, N13279);
not NOT1 (N22236, N22202);
nand NAND2 (N22237, N22230, N1880);
not NOT1 (N22238, N22237);
and AND2 (N22239, N22236, N10678);
or OR3 (N22240, N22233, N9600, N18414);
nor NOR3 (N22241, N22234, N17713, N11509);
and AND4 (N22242, N22222, N1094, N20209, N10787);
nor NOR4 (N22243, N22238, N5473, N4601, N9243);
buf BUF1 (N22244, N22231);
or OR2 (N22245, N22241, N14892);
or OR2 (N22246, N22235, N8825);
and AND3 (N22247, N22245, N6803, N1704);
and AND3 (N22248, N22243, N8361, N17977);
nor NOR4 (N22249, N22246, N3362, N15529, N9156);
xor XOR2 (N22250, N22240, N3998);
xor XOR2 (N22251, N22250, N8449);
nand NAND3 (N22252, N22224, N13051, N16327);
xor XOR2 (N22253, N22239, N6545);
nor NOR3 (N22254, N22244, N18284, N3383);
nor NOR3 (N22255, N22249, N10902, N12877);
or OR3 (N22256, N22242, N11093, N4590);
nor NOR2 (N22257, N22255, N12938);
or OR3 (N22258, N22252, N3728, N18836);
and AND3 (N22259, N22256, N16048, N5022);
not NOT1 (N22260, N22228);
and AND4 (N22261, N22251, N18113, N21929, N14532);
and AND2 (N22262, N22254, N15513);
buf BUF1 (N22263, N22248);
not NOT1 (N22264, N22262);
nand NAND2 (N22265, N22264, N4081);
buf BUF1 (N22266, N22261);
and AND2 (N22267, N22259, N9314);
nand NAND4 (N22268, N22221, N19642, N18283, N14257);
and AND4 (N22269, N22258, N11019, N16957, N7673);
nor NOR4 (N22270, N22253, N13083, N12668, N15445);
and AND4 (N22271, N22270, N16390, N11218, N20422);
and AND3 (N22272, N22263, N19652, N9722);
nor NOR3 (N22273, N22271, N21334, N8265);
nand NAND4 (N22274, N22247, N21928, N1903, N7651);
nor NOR4 (N22275, N22267, N4743, N2488, N2719);
nand NAND2 (N22276, N22260, N7148);
nor NOR3 (N22277, N22269, N8040, N9652);
buf BUF1 (N22278, N22273);
nand NAND4 (N22279, N22274, N18480, N18593, N336);
or OR4 (N22280, N22257, N3788, N5819, N6960);
buf BUF1 (N22281, N22276);
not NOT1 (N22282, N22281);
and AND3 (N22283, N22268, N4569, N11854);
and AND2 (N22284, N22275, N8444);
and AND3 (N22285, N22283, N4724, N10405);
and AND4 (N22286, N22279, N19007, N17496, N9790);
not NOT1 (N22287, N22266);
xor XOR2 (N22288, N22280, N19979);
buf BUF1 (N22289, N22286);
and AND4 (N22290, N22285, N7653, N20411, N21025);
not NOT1 (N22291, N22288);
or OR2 (N22292, N22282, N4675);
buf BUF1 (N22293, N22265);
not NOT1 (N22294, N22289);
and AND3 (N22295, N22290, N13265, N12787);
buf BUF1 (N22296, N22272);
buf BUF1 (N22297, N22291);
nor NOR4 (N22298, N22293, N20613, N1979, N7491);
nor NOR4 (N22299, N22292, N3518, N5961, N21684);
xor XOR2 (N22300, N22294, N5226);
or OR4 (N22301, N22300, N9030, N17218, N18823);
xor XOR2 (N22302, N22278, N1144);
buf BUF1 (N22303, N22277);
xor XOR2 (N22304, N22303, N18161);
or OR4 (N22305, N22297, N21454, N3839, N17758);
not NOT1 (N22306, N22287);
xor XOR2 (N22307, N22298, N3746);
and AND3 (N22308, N22305, N92, N1901);
nand NAND4 (N22309, N22302, N12099, N6292, N991);
xor XOR2 (N22310, N22306, N20467);
xor XOR2 (N22311, N22307, N19234);
nor NOR4 (N22312, N22284, N5706, N2260, N21645);
nand NAND2 (N22313, N22301, N21939);
or OR3 (N22314, N22299, N7491, N3754);
not NOT1 (N22315, N22314);
buf BUF1 (N22316, N22295);
nor NOR3 (N22317, N22308, N3731, N3041);
not NOT1 (N22318, N22313);
xor XOR2 (N22319, N22309, N15632);
xor XOR2 (N22320, N22304, N20168);
or OR4 (N22321, N22320, N11463, N19447, N5210);
not NOT1 (N22322, N22310);
and AND4 (N22323, N22322, N177, N3861, N19425);
not NOT1 (N22324, N22315);
not NOT1 (N22325, N22321);
nor NOR4 (N22326, N22316, N12425, N16835, N20386);
or OR2 (N22327, N22326, N13769);
nand NAND3 (N22328, N22323, N18663, N11092);
not NOT1 (N22329, N22327);
xor XOR2 (N22330, N22329, N7138);
and AND4 (N22331, N22311, N16394, N11651, N13864);
or OR4 (N22332, N22296, N18132, N13833, N8025);
buf BUF1 (N22333, N22328);
nand NAND3 (N22334, N22325, N327, N19220);
or OR4 (N22335, N22317, N10220, N4441, N11913);
nand NAND4 (N22336, N22319, N17882, N14254, N11892);
buf BUF1 (N22337, N22335);
buf BUF1 (N22338, N22312);
and AND2 (N22339, N22333, N9705);
xor XOR2 (N22340, N22337, N20521);
and AND2 (N22341, N22318, N9997);
nand NAND4 (N22342, N22341, N6263, N8228, N5545);
nor NOR2 (N22343, N22339, N2007);
xor XOR2 (N22344, N22343, N7539);
xor XOR2 (N22345, N22342, N1203);
or OR4 (N22346, N22334, N12977, N8440, N5937);
nor NOR4 (N22347, N22324, N2931, N17474, N14819);
buf BUF1 (N22348, N22345);
buf BUF1 (N22349, N22330);
nand NAND3 (N22350, N22332, N5882, N1517);
nand NAND3 (N22351, N22349, N17427, N21939);
nor NOR2 (N22352, N22350, N9580);
not NOT1 (N22353, N22346);
buf BUF1 (N22354, N22340);
and AND3 (N22355, N22352, N14345, N22011);
xor XOR2 (N22356, N22347, N14059);
or OR2 (N22357, N22351, N14992);
or OR2 (N22358, N22336, N12967);
nor NOR2 (N22359, N22338, N14048);
nand NAND2 (N22360, N22357, N10653);
and AND3 (N22361, N22331, N16513, N8043);
or OR3 (N22362, N22348, N7620, N7847);
or OR4 (N22363, N22358, N12478, N16254, N16690);
or OR4 (N22364, N22360, N2766, N10470, N2802);
or OR4 (N22365, N22355, N6224, N19736, N4506);
buf BUF1 (N22366, N22344);
buf BUF1 (N22367, N22356);
or OR4 (N22368, N22362, N20279, N11402, N19546);
and AND4 (N22369, N22354, N21514, N4162, N17044);
buf BUF1 (N22370, N22364);
buf BUF1 (N22371, N22366);
or OR2 (N22372, N22359, N4211);
buf BUF1 (N22373, N22365);
xor XOR2 (N22374, N22363, N21978);
and AND4 (N22375, N22361, N19562, N6932, N22178);
not NOT1 (N22376, N22374);
nand NAND4 (N22377, N22370, N10454, N7741, N9300);
not NOT1 (N22378, N22371);
and AND2 (N22379, N22353, N8476);
or OR3 (N22380, N22368, N15017, N11244);
buf BUF1 (N22381, N22379);
and AND3 (N22382, N22376, N13449, N10355);
not NOT1 (N22383, N22372);
nand NAND2 (N22384, N22378, N5862);
xor XOR2 (N22385, N22373, N17627);
buf BUF1 (N22386, N22369);
nand NAND3 (N22387, N22377, N21776, N3203);
nand NAND3 (N22388, N22367, N1209, N13522);
or OR4 (N22389, N22375, N10150, N15992, N10387);
not NOT1 (N22390, N22388);
nand NAND4 (N22391, N22381, N3333, N20035, N2629);
nand NAND4 (N22392, N22390, N19657, N11471, N21450);
and AND2 (N22393, N22380, N15408);
xor XOR2 (N22394, N22384, N8665);
not NOT1 (N22395, N22386);
buf BUF1 (N22396, N22389);
nor NOR2 (N22397, N22392, N2303);
xor XOR2 (N22398, N22387, N21801);
nand NAND3 (N22399, N22398, N10913, N17613);
nor NOR2 (N22400, N22397, N246);
xor XOR2 (N22401, N22393, N15575);
xor XOR2 (N22402, N22400, N242);
nor NOR4 (N22403, N22402, N14809, N17605, N21402);
buf BUF1 (N22404, N22394);
or OR4 (N22405, N22403, N3172, N20940, N13528);
nor NOR2 (N22406, N22382, N21152);
and AND3 (N22407, N22391, N14239, N8798);
nand NAND3 (N22408, N22399, N454, N9438);
nor NOR4 (N22409, N22404, N9150, N11465, N14058);
and AND4 (N22410, N22401, N17796, N1302, N19189);
nor NOR3 (N22411, N22409, N18854, N12166);
nor NOR3 (N22412, N22408, N5002, N11768);
nor NOR4 (N22413, N22411, N14611, N18087, N3657);
and AND3 (N22414, N22405, N17987, N6586);
xor XOR2 (N22415, N22396, N5486);
and AND3 (N22416, N22415, N9103, N22393);
and AND3 (N22417, N22413, N13525, N16098);
nand NAND4 (N22418, N22412, N15728, N18642, N16898);
and AND2 (N22419, N22395, N9305);
nor NOR2 (N22420, N22416, N12396);
not NOT1 (N22421, N22407);
and AND3 (N22422, N22406, N9104, N3190);
nand NAND4 (N22423, N22417, N8016, N7990, N1577);
nor NOR2 (N22424, N22418, N11932);
or OR4 (N22425, N22410, N21194, N3062, N3993);
and AND3 (N22426, N22423, N17555, N11193);
nor NOR3 (N22427, N22385, N6846, N2751);
nand NAND3 (N22428, N22421, N6493, N340);
buf BUF1 (N22429, N22414);
and AND4 (N22430, N22420, N311, N6722, N2945);
nor NOR2 (N22431, N22425, N17677);
buf BUF1 (N22432, N22426);
not NOT1 (N22433, N22419);
nand NAND3 (N22434, N22429, N14341, N14898);
or OR3 (N22435, N22431, N12992, N4258);
and AND3 (N22436, N22430, N10401, N15402);
or OR4 (N22437, N22424, N18442, N18447, N19710);
and AND4 (N22438, N22422, N301, N14729, N7808);
nor NOR4 (N22439, N22434, N4017, N4886, N17297);
nand NAND4 (N22440, N22428, N13230, N15174, N13253);
nor NOR3 (N22441, N22439, N12714, N21002);
or OR2 (N22442, N22433, N13507);
xor XOR2 (N22443, N22427, N7169);
and AND3 (N22444, N22440, N999, N18692);
or OR2 (N22445, N22436, N18567);
and AND3 (N22446, N22443, N17382, N8349);
buf BUF1 (N22447, N22446);
and AND3 (N22448, N22435, N4057, N16164);
not NOT1 (N22449, N22442);
xor XOR2 (N22450, N22445, N15222);
buf BUF1 (N22451, N22444);
nand NAND2 (N22452, N22447, N13885);
nor NOR2 (N22453, N22438, N21837);
nand NAND3 (N22454, N22383, N3816, N4528);
xor XOR2 (N22455, N22432, N20595);
nand NAND4 (N22456, N22451, N15197, N12487, N4598);
nand NAND3 (N22457, N22452, N9393, N1956);
buf BUF1 (N22458, N22437);
and AND2 (N22459, N22457, N13075);
nor NOR2 (N22460, N22453, N18658);
nand NAND3 (N22461, N22455, N20062, N4050);
xor XOR2 (N22462, N22460, N18486);
nand NAND4 (N22463, N22462, N14077, N14924, N20879);
buf BUF1 (N22464, N22456);
xor XOR2 (N22465, N22459, N8002);
not NOT1 (N22466, N22458);
nor NOR2 (N22467, N22466, N536);
buf BUF1 (N22468, N22464);
or OR4 (N22469, N22441, N15041, N2524, N6403);
nand NAND4 (N22470, N22468, N8546, N9303, N14210);
nand NAND2 (N22471, N22463, N5708);
or OR2 (N22472, N22454, N18346);
xor XOR2 (N22473, N22465, N3131);
xor XOR2 (N22474, N22449, N8523);
xor XOR2 (N22475, N22472, N3916);
nor NOR2 (N22476, N22471, N2906);
nand NAND3 (N22477, N22473, N4204, N9864);
buf BUF1 (N22478, N22474);
buf BUF1 (N22479, N22478);
xor XOR2 (N22480, N22475, N19986);
or OR4 (N22481, N22450, N12559, N142, N17638);
not NOT1 (N22482, N22467);
buf BUF1 (N22483, N22479);
or OR4 (N22484, N22481, N10015, N5419, N11436);
nand NAND3 (N22485, N22469, N14198, N8674);
nand NAND3 (N22486, N22477, N5010, N477);
not NOT1 (N22487, N22483);
buf BUF1 (N22488, N22482);
nor NOR2 (N22489, N22485, N19037);
or OR3 (N22490, N22489, N18789, N10368);
not NOT1 (N22491, N22476);
buf BUF1 (N22492, N22488);
or OR3 (N22493, N22490, N16971, N19874);
or OR2 (N22494, N22486, N1721);
not NOT1 (N22495, N22491);
not NOT1 (N22496, N22492);
xor XOR2 (N22497, N22494, N4122);
or OR3 (N22498, N22493, N16956, N16407);
nand NAND2 (N22499, N22497, N1501);
nand NAND3 (N22500, N22499, N12996, N11510);
or OR2 (N22501, N22487, N904);
and AND2 (N22502, N22496, N18071);
and AND2 (N22503, N22502, N9953);
nand NAND4 (N22504, N22501, N9845, N21899, N15847);
and AND4 (N22505, N22495, N18148, N3089, N12783);
xor XOR2 (N22506, N22505, N9593);
or OR3 (N22507, N22498, N7749, N1937);
not NOT1 (N22508, N22503);
nor NOR4 (N22509, N22506, N4809, N7781, N5032);
not NOT1 (N22510, N22470);
or OR4 (N22511, N22484, N2655, N19860, N8789);
buf BUF1 (N22512, N22510);
and AND3 (N22513, N22507, N15018, N2211);
buf BUF1 (N22514, N22511);
nand NAND4 (N22515, N22509, N8392, N15560, N7682);
xor XOR2 (N22516, N22508, N8977);
xor XOR2 (N22517, N22516, N3851);
nor NOR3 (N22518, N22448, N940, N14233);
nand NAND4 (N22519, N22480, N569, N12082, N9510);
buf BUF1 (N22520, N22514);
and AND2 (N22521, N22461, N5595);
not NOT1 (N22522, N22520);
or OR3 (N22523, N22519, N18365, N16696);
buf BUF1 (N22524, N22517);
and AND4 (N22525, N22515, N8021, N4365, N21983);
or OR2 (N22526, N22522, N7792);
nand NAND3 (N22527, N22526, N3715, N1377);
xor XOR2 (N22528, N22523, N20435);
xor XOR2 (N22529, N22525, N13812);
not NOT1 (N22530, N22521);
or OR4 (N22531, N22527, N21159, N1915, N2480);
nand NAND3 (N22532, N22513, N1430, N6212);
or OR2 (N22533, N22530, N19234);
not NOT1 (N22534, N22500);
nor NOR3 (N22535, N22504, N6733, N10242);
nor NOR4 (N22536, N22512, N21675, N10728, N17015);
and AND4 (N22537, N22536, N10356, N3034, N22449);
xor XOR2 (N22538, N22537, N582);
not NOT1 (N22539, N22524);
buf BUF1 (N22540, N22532);
xor XOR2 (N22541, N22529, N4548);
nor NOR2 (N22542, N22538, N16305);
nor NOR3 (N22543, N22541, N15154, N20367);
nor NOR4 (N22544, N22528, N721, N19390, N15354);
nand NAND2 (N22545, N22542, N21342);
nor NOR4 (N22546, N22543, N1317, N14652, N18470);
and AND3 (N22547, N22531, N18691, N5651);
nor NOR4 (N22548, N22540, N17771, N9090, N11684);
xor XOR2 (N22549, N22545, N9975);
or OR4 (N22550, N22518, N8139, N8956, N14683);
xor XOR2 (N22551, N22535, N7125);
and AND2 (N22552, N22544, N14096);
or OR2 (N22553, N22547, N6208);
nand NAND4 (N22554, N22553, N14986, N11802, N5588);
or OR4 (N22555, N22552, N14221, N12146, N3265);
nand NAND4 (N22556, N22549, N8926, N13691, N17904);
not NOT1 (N22557, N22546);
buf BUF1 (N22558, N22548);
and AND4 (N22559, N22539, N15165, N7, N20300);
not NOT1 (N22560, N22533);
nand NAND2 (N22561, N22550, N3100);
or OR4 (N22562, N22560, N13966, N12224, N4872);
and AND3 (N22563, N22555, N12906, N20955);
nor NOR2 (N22564, N22556, N12703);
buf BUF1 (N22565, N22554);
not NOT1 (N22566, N22559);
not NOT1 (N22567, N22551);
buf BUF1 (N22568, N22557);
and AND2 (N22569, N22567, N18405);
or OR2 (N22570, N22558, N17961);
not NOT1 (N22571, N22562);
and AND2 (N22572, N22568, N19588);
or OR2 (N22573, N22570, N950);
or OR3 (N22574, N22573, N19733, N13655);
or OR4 (N22575, N22572, N3945, N8490, N12930);
or OR4 (N22576, N22575, N1295, N1228, N16910);
xor XOR2 (N22577, N22563, N7947);
and AND2 (N22578, N22534, N19363);
nand NAND2 (N22579, N22561, N6718);
and AND4 (N22580, N22566, N15241, N3920, N6546);
and AND3 (N22581, N22578, N17505, N2349);
and AND4 (N22582, N22580, N17664, N21225, N3397);
and AND2 (N22583, N22576, N11582);
xor XOR2 (N22584, N22581, N6390);
nor NOR3 (N22585, N22579, N6428, N875);
or OR2 (N22586, N22585, N11499);
buf BUF1 (N22587, N22582);
not NOT1 (N22588, N22565);
nor NOR2 (N22589, N22574, N2813);
and AND2 (N22590, N22564, N1654);
nor NOR3 (N22591, N22584, N15004, N15281);
not NOT1 (N22592, N22591);
buf BUF1 (N22593, N22588);
buf BUF1 (N22594, N22577);
xor XOR2 (N22595, N22587, N14628);
nand NAND2 (N22596, N22583, N6069);
nor NOR2 (N22597, N22592, N7775);
buf BUF1 (N22598, N22569);
buf BUF1 (N22599, N22589);
nor NOR3 (N22600, N22586, N12065, N15457);
nand NAND3 (N22601, N22595, N17688, N875);
not NOT1 (N22602, N22597);
nand NAND3 (N22603, N22596, N18056, N22148);
buf BUF1 (N22604, N22599);
not NOT1 (N22605, N22603);
not NOT1 (N22606, N22601);
nor NOR4 (N22607, N22604, N13270, N261, N18825);
or OR4 (N22608, N22598, N12932, N5413, N9985);
and AND3 (N22609, N22571, N283, N5418);
or OR3 (N22610, N22608, N7232, N3905);
nand NAND2 (N22611, N22610, N6017);
nand NAND4 (N22612, N22600, N3707, N7587, N9430);
and AND4 (N22613, N22612, N16445, N5505, N19135);
nand NAND2 (N22614, N22593, N8494);
nand NAND2 (N22615, N22609, N18471);
not NOT1 (N22616, N22590);
and AND4 (N22617, N22614, N3377, N19484, N11443);
or OR3 (N22618, N22594, N13292, N3710);
or OR4 (N22619, N22615, N17839, N3341, N2398);
or OR2 (N22620, N22606, N3677);
nor NOR2 (N22621, N22602, N14248);
nor NOR4 (N22622, N22616, N16970, N16920, N16860);
or OR4 (N22623, N22621, N20289, N17929, N7300);
not NOT1 (N22624, N22623);
xor XOR2 (N22625, N22622, N7701);
xor XOR2 (N22626, N22607, N142);
xor XOR2 (N22627, N22619, N811);
nor NOR2 (N22628, N22626, N16151);
not NOT1 (N22629, N22605);
buf BUF1 (N22630, N22628);
xor XOR2 (N22631, N22624, N16793);
and AND3 (N22632, N22618, N20972, N4035);
xor XOR2 (N22633, N22630, N16514);
nand NAND3 (N22634, N22613, N636, N17444);
nor NOR4 (N22635, N22625, N2548, N5214, N4565);
nor NOR3 (N22636, N22611, N13055, N17586);
nor NOR4 (N22637, N22627, N20258, N5126, N21874);
nand NAND3 (N22638, N22617, N14254, N10310);
not NOT1 (N22639, N22633);
buf BUF1 (N22640, N22620);
nand NAND4 (N22641, N22636, N19132, N4378, N12141);
not NOT1 (N22642, N22638);
xor XOR2 (N22643, N22640, N18897);
and AND3 (N22644, N22632, N10410, N7532);
nand NAND3 (N22645, N22637, N9886, N13498);
and AND2 (N22646, N22639, N9493);
and AND4 (N22647, N22646, N4621, N22381, N21462);
nand NAND3 (N22648, N22634, N17659, N9169);
and AND2 (N22649, N22641, N9117);
xor XOR2 (N22650, N22645, N13000);
nand NAND4 (N22651, N22650, N14377, N3829, N11197);
nand NAND2 (N22652, N22647, N12430);
not NOT1 (N22653, N22649);
not NOT1 (N22654, N22651);
or OR4 (N22655, N22642, N5181, N22067, N5233);
not NOT1 (N22656, N22643);
nor NOR2 (N22657, N22648, N12410);
buf BUF1 (N22658, N22631);
nor NOR2 (N22659, N22629, N7182);
nand NAND2 (N22660, N22652, N5061);
xor XOR2 (N22661, N22660, N11018);
or OR4 (N22662, N22657, N4373, N15036, N18803);
nand NAND2 (N22663, N22659, N952);
not NOT1 (N22664, N22635);
or OR2 (N22665, N22662, N21355);
or OR3 (N22666, N22664, N1263, N13522);
buf BUF1 (N22667, N22656);
xor XOR2 (N22668, N22661, N6194);
not NOT1 (N22669, N22654);
and AND2 (N22670, N22669, N15680);
xor XOR2 (N22671, N22665, N20641);
nand NAND3 (N22672, N22667, N10516, N11812);
not NOT1 (N22673, N22644);
not NOT1 (N22674, N22655);
and AND2 (N22675, N22672, N13119);
xor XOR2 (N22676, N22675, N7039);
and AND3 (N22677, N22676, N8910, N16290);
nor NOR4 (N22678, N22668, N9193, N6872, N3461);
nand NAND2 (N22679, N22673, N6307);
buf BUF1 (N22680, N22670);
and AND4 (N22681, N22674, N5708, N9867, N15786);
not NOT1 (N22682, N22658);
xor XOR2 (N22683, N22681, N8670);
nand NAND3 (N22684, N22666, N17975, N8536);
or OR2 (N22685, N22671, N6576);
nor NOR4 (N22686, N22685, N16266, N20954, N16985);
xor XOR2 (N22687, N22653, N17273);
not NOT1 (N22688, N22677);
not NOT1 (N22689, N22687);
or OR2 (N22690, N22678, N16133);
nor NOR4 (N22691, N22684, N13447, N9403, N8866);
buf BUF1 (N22692, N22690);
nand NAND2 (N22693, N22682, N623);
nand NAND3 (N22694, N22683, N9666, N661);
nor NOR4 (N22695, N22688, N19556, N11956, N16313);
or OR3 (N22696, N22691, N9362, N21357);
nor NOR2 (N22697, N22694, N17299);
and AND3 (N22698, N22693, N18567, N13316);
buf BUF1 (N22699, N22680);
nor NOR3 (N22700, N22663, N18919, N777);
xor XOR2 (N22701, N22679, N22278);
or OR2 (N22702, N22692, N9774);
buf BUF1 (N22703, N22702);
or OR2 (N22704, N22699, N11493);
xor XOR2 (N22705, N22704, N2360);
nor NOR4 (N22706, N22703, N12512, N1135, N17421);
buf BUF1 (N22707, N22698);
not NOT1 (N22708, N22689);
nor NOR2 (N22709, N22706, N872);
nor NOR4 (N22710, N22696, N6094, N1156, N4859);
and AND2 (N22711, N22707, N6282);
and AND2 (N22712, N22697, N10632);
and AND2 (N22713, N22709, N19791);
nor NOR4 (N22714, N22686, N13025, N18465, N15826);
and AND4 (N22715, N22713, N21929, N11570, N8086);
nor NOR3 (N22716, N22712, N20134, N3285);
not NOT1 (N22717, N22710);
nor NOR4 (N22718, N22705, N551, N18302, N4137);
xor XOR2 (N22719, N22716, N3478);
not NOT1 (N22720, N22718);
nor NOR3 (N22721, N22719, N12704, N22595);
nand NAND4 (N22722, N22720, N1973, N4167, N4008);
and AND3 (N22723, N22714, N8109, N1234);
and AND4 (N22724, N22722, N9169, N7296, N3008);
not NOT1 (N22725, N22717);
xor XOR2 (N22726, N22701, N9664);
nand NAND3 (N22727, N22721, N4502, N7874);
nor NOR3 (N22728, N22724, N2333, N11740);
nor NOR3 (N22729, N22715, N6543, N9299);
nor NOR2 (N22730, N22708, N19150);
buf BUF1 (N22731, N22725);
nand NAND3 (N22732, N22731, N3786, N18173);
buf BUF1 (N22733, N22695);
or OR4 (N22734, N22700, N21247, N22527, N1104);
not NOT1 (N22735, N22733);
nor NOR2 (N22736, N22727, N19177);
buf BUF1 (N22737, N22730);
not NOT1 (N22738, N22736);
buf BUF1 (N22739, N22728);
nand NAND3 (N22740, N22734, N4914, N3355);
not NOT1 (N22741, N22726);
not NOT1 (N22742, N22735);
or OR4 (N22743, N22732, N20940, N981, N8776);
and AND2 (N22744, N22741, N2274);
or OR3 (N22745, N22743, N5528, N16553);
nand NAND4 (N22746, N22738, N21856, N17405, N14667);
nand NAND4 (N22747, N22746, N9400, N9020, N6290);
or OR4 (N22748, N22737, N11130, N9138, N1883);
nand NAND2 (N22749, N22723, N20979);
buf BUF1 (N22750, N22749);
xor XOR2 (N22751, N22745, N8616);
nor NOR3 (N22752, N22739, N21867, N13533);
buf BUF1 (N22753, N22747);
and AND2 (N22754, N22748, N13619);
and AND3 (N22755, N22751, N19432, N7358);
nand NAND4 (N22756, N22742, N20323, N4547, N9463);
and AND2 (N22757, N22752, N3622);
nand NAND2 (N22758, N22740, N5850);
not NOT1 (N22759, N22729);
not NOT1 (N22760, N22755);
buf BUF1 (N22761, N22758);
nor NOR4 (N22762, N22757, N19301, N9970, N2435);
nand NAND2 (N22763, N22759, N18307);
and AND4 (N22764, N22711, N8059, N12086, N9944);
not NOT1 (N22765, N22760);
buf BUF1 (N22766, N22756);
nor NOR4 (N22767, N22754, N22042, N15436, N17286);
xor XOR2 (N22768, N22744, N8289);
nand NAND2 (N22769, N22762, N1394);
xor XOR2 (N22770, N22764, N2347);
or OR2 (N22771, N22753, N16807);
buf BUF1 (N22772, N22767);
xor XOR2 (N22773, N22770, N1128);
not NOT1 (N22774, N22763);
buf BUF1 (N22775, N22772);
nor NOR2 (N22776, N22750, N15154);
or OR2 (N22777, N22769, N3244);
buf BUF1 (N22778, N22768);
and AND2 (N22779, N22776, N21618);
nand NAND4 (N22780, N22775, N22535, N19838, N8392);
or OR3 (N22781, N22779, N5105, N7664);
xor XOR2 (N22782, N22780, N17382);
and AND2 (N22783, N22774, N6605);
not NOT1 (N22784, N22783);
nor NOR4 (N22785, N22761, N15983, N20387, N2538);
xor XOR2 (N22786, N22773, N6270);
nand NAND2 (N22787, N22786, N17272);
buf BUF1 (N22788, N22784);
xor XOR2 (N22789, N22787, N18924);
nand NAND4 (N22790, N22781, N1016, N6293, N14762);
and AND2 (N22791, N22790, N19716);
not NOT1 (N22792, N22778);
and AND3 (N22793, N22777, N15937, N4494);
nand NAND2 (N22794, N22782, N4575);
buf BUF1 (N22795, N22785);
nand NAND4 (N22796, N22766, N1856, N9535, N4691);
or OR3 (N22797, N22771, N18639, N10241);
nor NOR4 (N22798, N22792, N13962, N444, N9275);
xor XOR2 (N22799, N22794, N15671);
nand NAND3 (N22800, N22799, N10836, N861);
not NOT1 (N22801, N22796);
buf BUF1 (N22802, N22801);
not NOT1 (N22803, N22798);
xor XOR2 (N22804, N22765, N9678);
nand NAND4 (N22805, N22791, N11368, N1684, N21167);
or OR3 (N22806, N22800, N9248, N11651);
not NOT1 (N22807, N22789);
xor XOR2 (N22808, N22802, N2891);
or OR4 (N22809, N22795, N21425, N19902, N7613);
and AND2 (N22810, N22808, N478);
nor NOR3 (N22811, N22793, N22782, N17977);
xor XOR2 (N22812, N22811, N20963);
nor NOR3 (N22813, N22804, N2988, N18367);
not NOT1 (N22814, N22812);
nand NAND3 (N22815, N22803, N7649, N11094);
buf BUF1 (N22816, N22815);
and AND3 (N22817, N22814, N2186, N18879);
buf BUF1 (N22818, N22788);
or OR3 (N22819, N22816, N15726, N10520);
nor NOR4 (N22820, N22809, N8105, N14497, N5712);
and AND3 (N22821, N22819, N20578, N1508);
xor XOR2 (N22822, N22818, N15364);
buf BUF1 (N22823, N22822);
or OR4 (N22824, N22797, N22195, N3206, N2162);
xor XOR2 (N22825, N22805, N6428);
or OR4 (N22826, N22806, N9847, N15378, N15134);
buf BUF1 (N22827, N22823);
xor XOR2 (N22828, N22817, N19169);
xor XOR2 (N22829, N22826, N13416);
buf BUF1 (N22830, N22807);
xor XOR2 (N22831, N22820, N20139);
nand NAND4 (N22832, N22821, N11216, N13409, N22366);
and AND4 (N22833, N22825, N22348, N12874, N15686);
not NOT1 (N22834, N22833);
not NOT1 (N22835, N22832);
nor NOR3 (N22836, N22827, N10651, N16002);
buf BUF1 (N22837, N22824);
or OR4 (N22838, N22813, N21016, N1046, N10703);
nor NOR4 (N22839, N22837, N17520, N10510, N5922);
nor NOR4 (N22840, N22838, N2857, N18930, N10881);
buf BUF1 (N22841, N22829);
nor NOR4 (N22842, N22830, N21292, N3885, N10765);
nand NAND2 (N22843, N22839, N4680);
and AND2 (N22844, N22842, N14426);
xor XOR2 (N22845, N22828, N9541);
or OR4 (N22846, N22843, N18971, N5042, N7692);
and AND4 (N22847, N22845, N11981, N6048, N1048);
xor XOR2 (N22848, N22831, N20436);
buf BUF1 (N22849, N22836);
not NOT1 (N22850, N22848);
buf BUF1 (N22851, N22844);
and AND4 (N22852, N22847, N22576, N16855, N3873);
and AND2 (N22853, N22834, N6119);
nand NAND2 (N22854, N22852, N18740);
xor XOR2 (N22855, N22854, N12801);
xor XOR2 (N22856, N22846, N22276);
not NOT1 (N22857, N22856);
or OR2 (N22858, N22857, N6262);
buf BUF1 (N22859, N22841);
xor XOR2 (N22860, N22835, N22277);
or OR2 (N22861, N22810, N5990);
xor XOR2 (N22862, N22851, N2701);
or OR3 (N22863, N22853, N7078, N12354);
nand NAND2 (N22864, N22862, N14984);
buf BUF1 (N22865, N22864);
xor XOR2 (N22866, N22858, N6096);
or OR2 (N22867, N22863, N9591);
xor XOR2 (N22868, N22860, N15117);
not NOT1 (N22869, N22850);
not NOT1 (N22870, N22849);
not NOT1 (N22871, N22867);
nand NAND2 (N22872, N22871, N9680);
and AND3 (N22873, N22870, N17617, N10889);
or OR2 (N22874, N22873, N18736);
xor XOR2 (N22875, N22872, N4132);
not NOT1 (N22876, N22840);
nand NAND2 (N22877, N22869, N9486);
buf BUF1 (N22878, N22877);
and AND3 (N22879, N22855, N16781, N9724);
xor XOR2 (N22880, N22876, N10322);
nand NAND3 (N22881, N22879, N7592, N3893);
xor XOR2 (N22882, N22865, N14854);
not NOT1 (N22883, N22861);
nand NAND4 (N22884, N22880, N3839, N7774, N22792);
xor XOR2 (N22885, N22859, N9908);
not NOT1 (N22886, N22878);
nor NOR3 (N22887, N22868, N18331, N5342);
nand NAND2 (N22888, N22886, N2889);
nor NOR3 (N22889, N22866, N21837, N12915);
or OR2 (N22890, N22875, N18054);
nand NAND4 (N22891, N22882, N18166, N6670, N17585);
and AND4 (N22892, N22888, N12645, N8985, N3994);
buf BUF1 (N22893, N22889);
and AND4 (N22894, N22874, N3349, N10329, N19899);
xor XOR2 (N22895, N22893, N21481);
buf BUF1 (N22896, N22885);
xor XOR2 (N22897, N22890, N10661);
xor XOR2 (N22898, N22894, N13965);
nor NOR2 (N22899, N22896, N9069);
nor NOR2 (N22900, N22898, N3493);
nand NAND4 (N22901, N22900, N323, N15843, N10725);
and AND2 (N22902, N22891, N15404);
buf BUF1 (N22903, N22897);
not NOT1 (N22904, N22901);
xor XOR2 (N22905, N22904, N13713);
nor NOR4 (N22906, N22905, N18870, N17105, N11992);
not NOT1 (N22907, N22892);
xor XOR2 (N22908, N22903, N16215);
buf BUF1 (N22909, N22906);
buf BUF1 (N22910, N22908);
xor XOR2 (N22911, N22909, N9157);
nand NAND3 (N22912, N22911, N18024, N16908);
nand NAND4 (N22913, N22895, N21027, N21339, N22492);
xor XOR2 (N22914, N22887, N5544);
or OR4 (N22915, N22899, N19564, N20694, N18745);
or OR3 (N22916, N22907, N6692, N22817);
not NOT1 (N22917, N22884);
nor NOR2 (N22918, N22881, N14920);
buf BUF1 (N22919, N22916);
nand NAND2 (N22920, N22915, N2666);
buf BUF1 (N22921, N22883);
buf BUF1 (N22922, N22918);
buf BUF1 (N22923, N22922);
nand NAND2 (N22924, N22919, N432);
xor XOR2 (N22925, N22924, N8347);
xor XOR2 (N22926, N22921, N8417);
or OR3 (N22927, N22902, N496, N16256);
nand NAND2 (N22928, N22913, N19572);
xor XOR2 (N22929, N22910, N7639);
and AND3 (N22930, N22923, N9430, N18666);
buf BUF1 (N22931, N22914);
not NOT1 (N22932, N22925);
nor NOR4 (N22933, N22932, N12656, N7954, N9087);
nor NOR4 (N22934, N22917, N11366, N13588, N13532);
and AND3 (N22935, N22930, N6420, N701);
nand NAND3 (N22936, N22926, N1586, N3921);
buf BUF1 (N22937, N22933);
not NOT1 (N22938, N22935);
buf BUF1 (N22939, N22920);
or OR3 (N22940, N22939, N11271, N14780);
buf BUF1 (N22941, N22912);
buf BUF1 (N22942, N22936);
nand NAND2 (N22943, N22927, N15425);
buf BUF1 (N22944, N22941);
nor NOR4 (N22945, N22934, N13622, N9038, N21318);
nand NAND4 (N22946, N22945, N22441, N14786, N18482);
nor NOR4 (N22947, N22940, N12319, N21881, N9363);
xor XOR2 (N22948, N22943, N799);
not NOT1 (N22949, N22944);
not NOT1 (N22950, N22946);
buf BUF1 (N22951, N22948);
and AND4 (N22952, N22929, N12205, N1110, N13552);
xor XOR2 (N22953, N22928, N19022);
nand NAND2 (N22954, N22950, N19972);
not NOT1 (N22955, N22947);
nor NOR2 (N22956, N22938, N12069);
or OR3 (N22957, N22956, N6697, N14557);
buf BUF1 (N22958, N22931);
not NOT1 (N22959, N22951);
not NOT1 (N22960, N22949);
not NOT1 (N22961, N22955);
buf BUF1 (N22962, N22953);
nor NOR4 (N22963, N22937, N8594, N5482, N19392);
buf BUF1 (N22964, N22963);
nor NOR4 (N22965, N22952, N12695, N4620, N142);
and AND2 (N22966, N22954, N506);
buf BUF1 (N22967, N22960);
buf BUF1 (N22968, N22942);
xor XOR2 (N22969, N22957, N6563);
and AND2 (N22970, N22961, N9307);
nor NOR4 (N22971, N22962, N20565, N21814, N13135);
or OR3 (N22972, N22966, N8156, N5684);
nor NOR4 (N22973, N22970, N16573, N17920, N7136);
and AND2 (N22974, N22959, N14963);
and AND4 (N22975, N22958, N3080, N22209, N22187);
buf BUF1 (N22976, N22968);
not NOT1 (N22977, N22965);
not NOT1 (N22978, N22964);
or OR3 (N22979, N22976, N12030, N11536);
nor NOR4 (N22980, N22973, N4972, N17310, N3938);
and AND2 (N22981, N22974, N3746);
or OR3 (N22982, N22980, N3641, N18976);
and AND4 (N22983, N22967, N20410, N22245, N14045);
and AND3 (N22984, N22969, N2261, N18742);
xor XOR2 (N22985, N22983, N18096);
and AND3 (N22986, N22975, N20023, N17346);
not NOT1 (N22987, N22984);
not NOT1 (N22988, N22972);
not NOT1 (N22989, N22981);
buf BUF1 (N22990, N22977);
or OR2 (N22991, N22986, N11087);
xor XOR2 (N22992, N22989, N6980);
and AND4 (N22993, N22978, N15910, N2254, N21648);
nand NAND2 (N22994, N22991, N15818);
nand NAND2 (N22995, N22990, N8136);
xor XOR2 (N22996, N22979, N7360);
or OR4 (N22997, N22995, N4881, N12099, N19795);
nand NAND2 (N22998, N22993, N16444);
nand NAND4 (N22999, N22998, N5393, N17340, N11239);
xor XOR2 (N23000, N22997, N22954);
xor XOR2 (N23001, N22982, N262);
xor XOR2 (N23002, N22992, N8990);
buf BUF1 (N23003, N22994);
or OR3 (N23004, N23003, N598, N4722);
nand NAND3 (N23005, N22996, N19923, N17636);
and AND3 (N23006, N23001, N20014, N9905);
buf BUF1 (N23007, N23005);
or OR3 (N23008, N23002, N1512, N6235);
nor NOR4 (N23009, N22988, N7166, N15641, N4103);
or OR2 (N23010, N22971, N1604);
or OR2 (N23011, N23009, N20245);
nand NAND4 (N23012, N23008, N4655, N3782, N5399);
nor NOR2 (N23013, N23012, N1519);
nor NOR3 (N23014, N23010, N22353, N12069);
nor NOR3 (N23015, N22985, N18332, N19791);
not NOT1 (N23016, N23006);
nand NAND4 (N23017, N23000, N4193, N16829, N21269);
and AND4 (N23018, N23011, N10709, N8089, N13159);
nand NAND3 (N23019, N23007, N22988, N12427);
nand NAND4 (N23020, N23017, N20237, N22318, N9501);
xor XOR2 (N23021, N22987, N22252);
not NOT1 (N23022, N23014);
not NOT1 (N23023, N23020);
or OR4 (N23024, N23004, N6325, N4225, N14317);
and AND3 (N23025, N23018, N17226, N11644);
or OR2 (N23026, N23016, N15989);
xor XOR2 (N23027, N23019, N16965);
xor XOR2 (N23028, N23022, N19534);
xor XOR2 (N23029, N23026, N13775);
nor NOR4 (N23030, N22999, N11787, N18163, N22584);
nand NAND2 (N23031, N23027, N18072);
buf BUF1 (N23032, N23013);
and AND2 (N23033, N23030, N10446);
or OR2 (N23034, N23028, N3352);
buf BUF1 (N23035, N23032);
or OR3 (N23036, N23021, N6212, N18238);
nor NOR3 (N23037, N23023, N11416, N12036);
and AND3 (N23038, N23031, N18855, N13879);
and AND2 (N23039, N23038, N10388);
not NOT1 (N23040, N23025);
nor NOR2 (N23041, N23029, N15995);
nand NAND2 (N23042, N23036, N19578);
and AND4 (N23043, N23034, N3311, N19252, N7234);
xor XOR2 (N23044, N23037, N10386);
or OR3 (N23045, N23043, N5874, N20816);
not NOT1 (N23046, N23015);
buf BUF1 (N23047, N23041);
nand NAND4 (N23048, N23042, N21076, N10645, N11522);
not NOT1 (N23049, N23044);
or OR3 (N23050, N23024, N730, N13406);
nand NAND4 (N23051, N23040, N22549, N7441, N18049);
nand NAND3 (N23052, N23033, N3754, N22112);
and AND2 (N23053, N23045, N1189);
nor NOR3 (N23054, N23046, N19010, N15713);
buf BUF1 (N23055, N23039);
nand NAND3 (N23056, N23053, N18283, N14682);
not NOT1 (N23057, N23049);
and AND2 (N23058, N23056, N19357);
nor NOR3 (N23059, N23035, N14923, N20563);
buf BUF1 (N23060, N23048);
not NOT1 (N23061, N23051);
nor NOR3 (N23062, N23047, N20102, N22998);
or OR3 (N23063, N23062, N15159, N5662);
buf BUF1 (N23064, N23059);
nand NAND2 (N23065, N23063, N6161);
buf BUF1 (N23066, N23050);
and AND3 (N23067, N23061, N16778, N16253);
xor XOR2 (N23068, N23052, N19589);
buf BUF1 (N23069, N23057);
and AND3 (N23070, N23058, N21751, N4505);
buf BUF1 (N23071, N23055);
and AND2 (N23072, N23067, N11453);
buf BUF1 (N23073, N23068);
nand NAND2 (N23074, N23054, N727);
buf BUF1 (N23075, N23069);
nand NAND4 (N23076, N23075, N12653, N6437, N6255);
or OR2 (N23077, N23060, N591);
not NOT1 (N23078, N23074);
not NOT1 (N23079, N23071);
and AND2 (N23080, N23076, N4566);
xor XOR2 (N23081, N23077, N287);
not NOT1 (N23082, N23081);
nand NAND2 (N23083, N23066, N10260);
buf BUF1 (N23084, N23072);
nand NAND4 (N23085, N23083, N570, N7451, N618);
or OR2 (N23086, N23079, N6334);
nand NAND2 (N23087, N23064, N20878);
nand NAND3 (N23088, N23070, N10664, N17590);
and AND2 (N23089, N23082, N10562);
buf BUF1 (N23090, N23078);
buf BUF1 (N23091, N23065);
buf BUF1 (N23092, N23080);
xor XOR2 (N23093, N23073, N21992);
not NOT1 (N23094, N23093);
and AND4 (N23095, N23092, N20675, N16344, N7800);
nor NOR3 (N23096, N23086, N5822, N8565);
xor XOR2 (N23097, N23084, N21375);
not NOT1 (N23098, N23094);
and AND3 (N23099, N23097, N14463, N6646);
nor NOR2 (N23100, N23088, N14632);
and AND2 (N23101, N23085, N22665);
nor NOR4 (N23102, N23098, N16659, N18837, N7122);
buf BUF1 (N23103, N23096);
buf BUF1 (N23104, N23099);
nand NAND4 (N23105, N23090, N7365, N13814, N6652);
xor XOR2 (N23106, N23103, N15591);
xor XOR2 (N23107, N23104, N14846);
xor XOR2 (N23108, N23095, N4846);
nand NAND3 (N23109, N23101, N11585, N3029);
xor XOR2 (N23110, N23087, N19416);
nand NAND3 (N23111, N23089, N10337, N19307);
buf BUF1 (N23112, N23110);
and AND4 (N23113, N23109, N17465, N21071, N11588);
nand NAND3 (N23114, N23105, N5408, N19520);
xor XOR2 (N23115, N23107, N19141);
buf BUF1 (N23116, N23111);
not NOT1 (N23117, N23115);
buf BUF1 (N23118, N23102);
not NOT1 (N23119, N23118);
nand NAND4 (N23120, N23117, N4029, N10071, N8973);
buf BUF1 (N23121, N23114);
xor XOR2 (N23122, N23116, N4429);
not NOT1 (N23123, N23120);
nor NOR4 (N23124, N23113, N14511, N26, N10838);
buf BUF1 (N23125, N23106);
nor NOR3 (N23126, N23121, N4773, N16796);
nor NOR4 (N23127, N23123, N226, N15643, N15840);
not NOT1 (N23128, N23091);
or OR3 (N23129, N23122, N13235, N22802);
nand NAND2 (N23130, N23100, N6068);
not NOT1 (N23131, N23108);
and AND2 (N23132, N23129, N1794);
nand NAND2 (N23133, N23112, N19901);
nor NOR3 (N23134, N23124, N3621, N20853);
xor XOR2 (N23135, N23126, N12416);
nand NAND3 (N23136, N23128, N3338, N17965);
and AND4 (N23137, N23134, N15127, N21222, N5216);
or OR2 (N23138, N23131, N558);
xor XOR2 (N23139, N23137, N10138);
not NOT1 (N23140, N23127);
or OR3 (N23141, N23138, N7856, N13746);
xor XOR2 (N23142, N23119, N20896);
xor XOR2 (N23143, N23136, N4944);
not NOT1 (N23144, N23132);
nor NOR4 (N23145, N23143, N2862, N5320, N2185);
not NOT1 (N23146, N23135);
not NOT1 (N23147, N23140);
buf BUF1 (N23148, N23146);
nor NOR2 (N23149, N23148, N20764);
buf BUF1 (N23150, N23147);
and AND3 (N23151, N23150, N8352, N18755);
xor XOR2 (N23152, N23125, N563);
not NOT1 (N23153, N23149);
nand NAND2 (N23154, N23144, N22871);
or OR2 (N23155, N23130, N491);
not NOT1 (N23156, N23154);
nand NAND2 (N23157, N23139, N8877);
and AND4 (N23158, N23145, N14140, N8034, N9114);
buf BUF1 (N23159, N23142);
and AND4 (N23160, N23153, N4408, N3702, N16240);
nand NAND4 (N23161, N23152, N15195, N22256, N16567);
or OR2 (N23162, N23157, N1903);
or OR2 (N23163, N23141, N2256);
not NOT1 (N23164, N23156);
nand NAND2 (N23165, N23160, N11182);
or OR3 (N23166, N23151, N15856, N9061);
and AND2 (N23167, N23161, N18623);
nand NAND4 (N23168, N23158, N20007, N9283, N22735);
not NOT1 (N23169, N23163);
buf BUF1 (N23170, N23166);
and AND3 (N23171, N23155, N7586, N4313);
or OR4 (N23172, N23169, N3574, N16805, N17446);
not NOT1 (N23173, N23167);
not NOT1 (N23174, N23168);
xor XOR2 (N23175, N23133, N986);
buf BUF1 (N23176, N23165);
not NOT1 (N23177, N23173);
buf BUF1 (N23178, N23164);
buf BUF1 (N23179, N23162);
and AND4 (N23180, N23174, N8922, N13138, N13454);
xor XOR2 (N23181, N23172, N142);
nand NAND2 (N23182, N23159, N3014);
not NOT1 (N23183, N23176);
or OR3 (N23184, N23175, N20370, N2713);
nand NAND4 (N23185, N23171, N6145, N4564, N9223);
xor XOR2 (N23186, N23177, N16707);
xor XOR2 (N23187, N23185, N22777);
or OR3 (N23188, N23181, N313, N3442);
buf BUF1 (N23189, N23188);
not NOT1 (N23190, N23186);
not NOT1 (N23191, N23184);
or OR3 (N23192, N23190, N8171, N13597);
xor XOR2 (N23193, N23183, N22945);
and AND3 (N23194, N23191, N21545, N13206);
buf BUF1 (N23195, N23180);
or OR4 (N23196, N23192, N14568, N16262, N9593);
not NOT1 (N23197, N23194);
nand NAND4 (N23198, N23197, N20549, N19295, N12325);
xor XOR2 (N23199, N23198, N15833);
or OR3 (N23200, N23179, N10505, N6837);
or OR4 (N23201, N23193, N10949, N5772, N701);
nor NOR2 (N23202, N23201, N20800);
xor XOR2 (N23203, N23189, N18283);
nor NOR4 (N23204, N23196, N1645, N9043, N3615);
not NOT1 (N23205, N23199);
nor NOR2 (N23206, N23200, N3743);
nand NAND3 (N23207, N23203, N22188, N15844);
buf BUF1 (N23208, N23206);
xor XOR2 (N23209, N23208, N16751);
nand NAND2 (N23210, N23178, N21162);
not NOT1 (N23211, N23170);
xor XOR2 (N23212, N23187, N15673);
or OR2 (N23213, N23207, N6500);
buf BUF1 (N23214, N23209);
xor XOR2 (N23215, N23204, N7069);
nor NOR3 (N23216, N23202, N1134, N14104);
not NOT1 (N23217, N23211);
not NOT1 (N23218, N23216);
not NOT1 (N23219, N23215);
or OR2 (N23220, N23214, N1350);
buf BUF1 (N23221, N23205);
nand NAND4 (N23222, N23219, N13877, N20253, N9899);
and AND2 (N23223, N23217, N8587);
buf BUF1 (N23224, N23220);
and AND3 (N23225, N23182, N13776, N7312);
nor NOR3 (N23226, N23223, N277, N8660);
or OR4 (N23227, N23212, N5762, N10689, N19474);
buf BUF1 (N23228, N23226);
buf BUF1 (N23229, N23210);
xor XOR2 (N23230, N23225, N6763);
not NOT1 (N23231, N23221);
xor XOR2 (N23232, N23228, N5837);
not NOT1 (N23233, N23222);
nand NAND3 (N23234, N23227, N12584, N6502);
or OR2 (N23235, N23195, N2492);
buf BUF1 (N23236, N23213);
or OR2 (N23237, N23218, N2090);
and AND3 (N23238, N23232, N12241, N18730);
xor XOR2 (N23239, N23229, N21637);
nand NAND3 (N23240, N23233, N15931, N15275);
buf BUF1 (N23241, N23237);
buf BUF1 (N23242, N23236);
buf BUF1 (N23243, N23234);
not NOT1 (N23244, N23224);
and AND2 (N23245, N23241, N13644);
not NOT1 (N23246, N23242);
not NOT1 (N23247, N23245);
nand NAND4 (N23248, N23235, N952, N10844, N23214);
xor XOR2 (N23249, N23230, N4263);
not NOT1 (N23250, N23240);
buf BUF1 (N23251, N23243);
and AND3 (N23252, N23238, N20590, N16201);
nor NOR4 (N23253, N23244, N698, N10296, N8631);
xor XOR2 (N23254, N23249, N13805);
buf BUF1 (N23255, N23253);
nor NOR4 (N23256, N23231, N11069, N16250, N10162);
and AND4 (N23257, N23248, N18432, N3066, N12470);
nand NAND2 (N23258, N23239, N18432);
nor NOR4 (N23259, N23246, N16620, N18653, N19105);
not NOT1 (N23260, N23254);
nand NAND2 (N23261, N23247, N21271);
buf BUF1 (N23262, N23260);
nand NAND4 (N23263, N23259, N8328, N22928, N16203);
nor NOR4 (N23264, N23250, N12643, N13456, N13060);
and AND2 (N23265, N23255, N19228);
nand NAND4 (N23266, N23261, N21443, N2852, N14371);
nand NAND3 (N23267, N23262, N6939, N11983);
not NOT1 (N23268, N23266);
not NOT1 (N23269, N23256);
or OR2 (N23270, N23258, N21063);
buf BUF1 (N23271, N23265);
nor NOR2 (N23272, N23267, N11823);
not NOT1 (N23273, N23270);
buf BUF1 (N23274, N23269);
not NOT1 (N23275, N23268);
nand NAND4 (N23276, N23251, N9508, N3289, N2740);
and AND4 (N23277, N23273, N19444, N20558, N20868);
nand NAND3 (N23278, N23252, N20973, N17242);
nand NAND2 (N23279, N23272, N20077);
not NOT1 (N23280, N23257);
and AND2 (N23281, N23277, N20926);
nor NOR4 (N23282, N23280, N21701, N19192, N3425);
xor XOR2 (N23283, N23282, N3234);
xor XOR2 (N23284, N23263, N5840);
or OR2 (N23285, N23281, N13552);
nor NOR4 (N23286, N23276, N15238, N14056, N15563);
buf BUF1 (N23287, N23274);
not NOT1 (N23288, N23286);
buf BUF1 (N23289, N23285);
nand NAND2 (N23290, N23278, N20953);
xor XOR2 (N23291, N23283, N5255);
buf BUF1 (N23292, N23290);
nand NAND2 (N23293, N23279, N20255);
nand NAND2 (N23294, N23293, N6752);
and AND2 (N23295, N23287, N22998);
xor XOR2 (N23296, N23264, N8108);
or OR4 (N23297, N23289, N4502, N19609, N6736);
not NOT1 (N23298, N23271);
nor NOR3 (N23299, N23292, N3301, N19707);
not NOT1 (N23300, N23294);
xor XOR2 (N23301, N23291, N12400);
nand NAND4 (N23302, N23284, N19006, N6828, N8346);
not NOT1 (N23303, N23302);
buf BUF1 (N23304, N23296);
not NOT1 (N23305, N23298);
not NOT1 (N23306, N23297);
xor XOR2 (N23307, N23275, N15744);
buf BUF1 (N23308, N23299);
buf BUF1 (N23309, N23308);
nor NOR4 (N23310, N23304, N13548, N19044, N15471);
not NOT1 (N23311, N23307);
nand NAND4 (N23312, N23288, N9775, N3502, N22536);
not NOT1 (N23313, N23310);
not NOT1 (N23314, N23305);
not NOT1 (N23315, N23306);
nor NOR2 (N23316, N23301, N8098);
and AND2 (N23317, N23309, N6545);
and AND3 (N23318, N23303, N39, N2580);
xor XOR2 (N23319, N23315, N1577);
buf BUF1 (N23320, N23312);
nor NOR3 (N23321, N23313, N23167, N7790);
xor XOR2 (N23322, N23319, N15498);
and AND2 (N23323, N23320, N8647);
nor NOR2 (N23324, N23323, N12673);
not NOT1 (N23325, N23316);
nor NOR2 (N23326, N23300, N997);
xor XOR2 (N23327, N23314, N21261);
nand NAND3 (N23328, N23321, N10088, N22073);
and AND3 (N23329, N23295, N20545, N2170);
xor XOR2 (N23330, N23325, N15580);
buf BUF1 (N23331, N23326);
nand NAND4 (N23332, N23328, N4169, N22371, N8998);
buf BUF1 (N23333, N23324);
nand NAND4 (N23334, N23327, N17214, N9930, N12056);
buf BUF1 (N23335, N23334);
xor XOR2 (N23336, N23317, N13504);
not NOT1 (N23337, N23336);
nor NOR4 (N23338, N23332, N16259, N3312, N20531);
and AND3 (N23339, N23337, N5182, N18238);
or OR3 (N23340, N23331, N21373, N3912);
or OR3 (N23341, N23330, N20059, N18490);
and AND4 (N23342, N23311, N2969, N19279, N16753);
or OR2 (N23343, N23318, N21096);
nor NOR3 (N23344, N23335, N2686, N2315);
and AND3 (N23345, N23322, N12352, N322);
not NOT1 (N23346, N23345);
nor NOR4 (N23347, N23329, N22644, N2645, N1892);
and AND4 (N23348, N23346, N9664, N6025, N6285);
xor XOR2 (N23349, N23348, N246);
or OR2 (N23350, N23349, N19078);
and AND2 (N23351, N23350, N18641);
buf BUF1 (N23352, N23351);
and AND2 (N23353, N23342, N4308);
xor XOR2 (N23354, N23338, N2169);
not NOT1 (N23355, N23333);
not NOT1 (N23356, N23353);
buf BUF1 (N23357, N23355);
and AND2 (N23358, N23356, N8356);
xor XOR2 (N23359, N23341, N15591);
nor NOR4 (N23360, N23347, N1087, N5289, N6712);
buf BUF1 (N23361, N23360);
xor XOR2 (N23362, N23340, N21590);
buf BUF1 (N23363, N23343);
not NOT1 (N23364, N23339);
not NOT1 (N23365, N23344);
xor XOR2 (N23366, N23359, N21101);
nor NOR3 (N23367, N23363, N22350, N22721);
nand NAND2 (N23368, N23362, N9514);
nand NAND4 (N23369, N23368, N14052, N20468, N15358);
nor NOR4 (N23370, N23361, N17084, N7649, N8940);
xor XOR2 (N23371, N23366, N4678);
and AND4 (N23372, N23365, N8974, N10046, N3674);
nor NOR2 (N23373, N23371, N2255);
and AND3 (N23374, N23373, N20148, N4864);
xor XOR2 (N23375, N23370, N2180);
buf BUF1 (N23376, N23364);
nor NOR2 (N23377, N23375, N2754);
buf BUF1 (N23378, N23358);
or OR2 (N23379, N23354, N15194);
buf BUF1 (N23380, N23357);
and AND4 (N23381, N23352, N5509, N13177, N9178);
not NOT1 (N23382, N23381);
buf BUF1 (N23383, N23379);
buf BUF1 (N23384, N23378);
not NOT1 (N23385, N23374);
buf BUF1 (N23386, N23382);
nand NAND4 (N23387, N23380, N5163, N18924, N14739);
nor NOR4 (N23388, N23372, N21137, N11523, N2763);
nor NOR2 (N23389, N23386, N4873);
nand NAND4 (N23390, N23369, N19110, N4760, N18065);
xor XOR2 (N23391, N23388, N20333);
and AND3 (N23392, N23389, N18483, N11505);
or OR3 (N23393, N23367, N11326, N9827);
nor NOR4 (N23394, N23376, N5019, N21515, N9086);
not NOT1 (N23395, N23383);
not NOT1 (N23396, N23393);
nor NOR4 (N23397, N23396, N11307, N270, N14008);
nor NOR3 (N23398, N23391, N22426, N21886);
not NOT1 (N23399, N23390);
nand NAND3 (N23400, N23394, N11395, N23149);
nor NOR4 (N23401, N23387, N15798, N16736, N18521);
or OR2 (N23402, N23400, N13372);
or OR4 (N23403, N23399, N19454, N5068, N6808);
nor NOR4 (N23404, N23402, N3330, N4234, N19021);
nand NAND4 (N23405, N23401, N12015, N10484, N18916);
nor NOR4 (N23406, N23395, N7562, N4433, N1289);
and AND3 (N23407, N23377, N19273, N115);
not NOT1 (N23408, N23385);
not NOT1 (N23409, N23404);
nand NAND2 (N23410, N23398, N22041);
xor XOR2 (N23411, N23409, N11817);
nand NAND2 (N23412, N23405, N23342);
nor NOR3 (N23413, N23408, N3256, N10989);
nand NAND2 (N23414, N23397, N2904);
xor XOR2 (N23415, N23384, N20954);
xor XOR2 (N23416, N23413, N11126);
xor XOR2 (N23417, N23410, N851);
nand NAND3 (N23418, N23416, N5687, N1284);
and AND2 (N23419, N23406, N17301);
nor NOR2 (N23420, N23417, N16705);
nand NAND4 (N23421, N23411, N22549, N13462, N2902);
nand NAND4 (N23422, N23392, N5641, N31, N13917);
xor XOR2 (N23423, N23412, N16995);
nor NOR4 (N23424, N23414, N3549, N2597, N4239);
buf BUF1 (N23425, N23420);
or OR2 (N23426, N23424, N18652);
buf BUF1 (N23427, N23425);
and AND4 (N23428, N23423, N16209, N7648, N15646);
or OR2 (N23429, N23426, N6744);
nand NAND3 (N23430, N23419, N12315, N10138);
buf BUF1 (N23431, N23430);
or OR3 (N23432, N23415, N17209, N15932);
or OR4 (N23433, N23429, N15527, N19597, N9303);
or OR4 (N23434, N23407, N5323, N9337, N6371);
nand NAND4 (N23435, N23421, N3901, N18891, N10830);
and AND2 (N23436, N23422, N19291);
and AND4 (N23437, N23432, N11805, N8254, N5452);
nand NAND3 (N23438, N23418, N12839, N17366);
and AND4 (N23439, N23433, N4796, N6154, N17657);
xor XOR2 (N23440, N23427, N15015);
nand NAND2 (N23441, N23440, N16425);
buf BUF1 (N23442, N23438);
xor XOR2 (N23443, N23434, N13393);
buf BUF1 (N23444, N23443);
or OR3 (N23445, N23441, N13349, N18571);
nor NOR4 (N23446, N23435, N7733, N13556, N8061);
or OR3 (N23447, N23437, N18525, N11869);
and AND2 (N23448, N23442, N9191);
or OR4 (N23449, N23431, N14333, N12110, N5310);
or OR2 (N23450, N23448, N1988);
or OR2 (N23451, N23449, N4837);
buf BUF1 (N23452, N23450);
buf BUF1 (N23453, N23444);
nor NOR2 (N23454, N23445, N9348);
not NOT1 (N23455, N23403);
nor NOR4 (N23456, N23452, N4757, N1585, N16899);
nand NAND2 (N23457, N23428, N12890);
or OR3 (N23458, N23456, N2832, N568);
nor NOR4 (N23459, N23454, N9672, N55, N2602);
nand NAND4 (N23460, N23453, N9504, N5431, N1868);
buf BUF1 (N23461, N23447);
nand NAND2 (N23462, N23439, N18054);
xor XOR2 (N23463, N23459, N11014);
buf BUF1 (N23464, N23436);
nor NOR4 (N23465, N23461, N21970, N7945, N15365);
or OR3 (N23466, N23446, N8740, N23216);
nor NOR2 (N23467, N23463, N3092);
and AND3 (N23468, N23458, N11966, N1345);
xor XOR2 (N23469, N23457, N4702);
xor XOR2 (N23470, N23451, N2612);
or OR3 (N23471, N23466, N8629, N23100);
not NOT1 (N23472, N23462);
nand NAND2 (N23473, N23468, N12529);
nand NAND2 (N23474, N23471, N7855);
nor NOR4 (N23475, N23470, N22416, N6055, N11190);
or OR2 (N23476, N23465, N18171);
xor XOR2 (N23477, N23476, N10677);
xor XOR2 (N23478, N23473, N1372);
not NOT1 (N23479, N23464);
and AND4 (N23480, N23474, N19838, N6273, N12433);
nand NAND3 (N23481, N23480, N13238, N17867);
buf BUF1 (N23482, N23469);
and AND2 (N23483, N23460, N6012);
buf BUF1 (N23484, N23483);
buf BUF1 (N23485, N23478);
and AND4 (N23486, N23477, N14524, N5813, N17041);
nor NOR3 (N23487, N23481, N7337, N18252);
nor NOR2 (N23488, N23485, N14314);
xor XOR2 (N23489, N23484, N1237);
or OR4 (N23490, N23487, N17980, N23260, N13666);
or OR2 (N23491, N23486, N23297);
buf BUF1 (N23492, N23479);
buf BUF1 (N23493, N23467);
buf BUF1 (N23494, N23490);
or OR4 (N23495, N23492, N6537, N10056, N12377);
nand NAND3 (N23496, N23491, N19826, N3668);
nand NAND2 (N23497, N23495, N16929);
not NOT1 (N23498, N23475);
and AND3 (N23499, N23494, N14818, N21637);
and AND4 (N23500, N23455, N5156, N20143, N15705);
or OR4 (N23501, N23497, N19377, N20590, N3327);
or OR4 (N23502, N23499, N10191, N22931, N11533);
and AND4 (N23503, N23502, N3471, N4638, N13431);
buf BUF1 (N23504, N23496);
nor NOR3 (N23505, N23500, N10139, N11346);
nor NOR4 (N23506, N23472, N2807, N15675, N18325);
nor NOR4 (N23507, N23501, N8506, N949, N14287);
not NOT1 (N23508, N23498);
and AND2 (N23509, N23493, N16245);
or OR2 (N23510, N23508, N12649);
and AND3 (N23511, N23505, N13278, N6046);
and AND4 (N23512, N23509, N21958, N4620, N145);
nor NOR2 (N23513, N23507, N20023);
buf BUF1 (N23514, N23482);
not NOT1 (N23515, N23510);
nor NOR2 (N23516, N23512, N12680);
and AND3 (N23517, N23506, N7302, N10537);
xor XOR2 (N23518, N23503, N10412);
buf BUF1 (N23519, N23517);
nand NAND4 (N23520, N23513, N6485, N749, N15247);
xor XOR2 (N23521, N23488, N13618);
and AND4 (N23522, N23489, N16675, N12066, N20060);
buf BUF1 (N23523, N23518);
buf BUF1 (N23524, N23515);
and AND2 (N23525, N23520, N20112);
not NOT1 (N23526, N23524);
nor NOR3 (N23527, N23519, N3932, N13859);
buf BUF1 (N23528, N23516);
nor NOR2 (N23529, N23526, N2403);
xor XOR2 (N23530, N23527, N3953);
buf BUF1 (N23531, N23521);
nor NOR4 (N23532, N23511, N11175, N21372, N4124);
nor NOR4 (N23533, N23529, N5777, N10431, N2338);
and AND2 (N23534, N23522, N3984);
xor XOR2 (N23535, N23504, N2039);
or OR3 (N23536, N23523, N11357, N13580);
and AND3 (N23537, N23525, N21539, N12448);
nand NAND3 (N23538, N23537, N8948, N18655);
nor NOR4 (N23539, N23535, N10657, N20059, N11039);
or OR3 (N23540, N23531, N22322, N12683);
buf BUF1 (N23541, N23530);
nor NOR4 (N23542, N23539, N8226, N2853, N1116);
nand NAND3 (N23543, N23532, N2114, N19186);
buf BUF1 (N23544, N23536);
nand NAND4 (N23545, N23543, N7439, N9141, N20497);
buf BUF1 (N23546, N23534);
not NOT1 (N23547, N23538);
xor XOR2 (N23548, N23528, N19071);
and AND3 (N23549, N23545, N8847, N13583);
or OR4 (N23550, N23548, N21664, N19246, N1784);
xor XOR2 (N23551, N23544, N13501);
and AND2 (N23552, N23550, N19685);
and AND3 (N23553, N23514, N11823, N5089);
and AND2 (N23554, N23547, N1737);
not NOT1 (N23555, N23551);
nor NOR4 (N23556, N23542, N17764, N8679, N11814);
not NOT1 (N23557, N23546);
xor XOR2 (N23558, N23533, N1931);
buf BUF1 (N23559, N23549);
xor XOR2 (N23560, N23556, N92);
or OR3 (N23561, N23554, N9125, N5393);
not NOT1 (N23562, N23557);
and AND2 (N23563, N23559, N689);
nand NAND4 (N23564, N23562, N16919, N14822, N17950);
not NOT1 (N23565, N23563);
nand NAND2 (N23566, N23560, N23081);
nand NAND4 (N23567, N23564, N23227, N11109, N20244);
and AND2 (N23568, N23558, N223);
nor NOR3 (N23569, N23568, N17700, N15980);
and AND3 (N23570, N23561, N22332, N15288);
and AND3 (N23571, N23555, N5757, N16391);
nor NOR2 (N23572, N23571, N423);
not NOT1 (N23573, N23553);
nor NOR2 (N23574, N23566, N20045);
nand NAND2 (N23575, N23567, N8817);
or OR3 (N23576, N23552, N19457, N8010);
xor XOR2 (N23577, N23570, N1220);
not NOT1 (N23578, N23573);
xor XOR2 (N23579, N23577, N11100);
buf BUF1 (N23580, N23575);
nand NAND2 (N23581, N23574, N6811);
nor NOR4 (N23582, N23578, N3809, N12584, N16708);
buf BUF1 (N23583, N23540);
and AND4 (N23584, N23541, N19290, N142, N2170);
xor XOR2 (N23585, N23569, N2525);
and AND3 (N23586, N23580, N17451, N23290);
nand NAND4 (N23587, N23572, N7092, N8182, N10386);
nor NOR2 (N23588, N23587, N13335);
or OR4 (N23589, N23565, N3337, N2984, N565);
xor XOR2 (N23590, N23583, N5458);
nor NOR4 (N23591, N23581, N23260, N10697, N13819);
nor NOR3 (N23592, N23591, N1655, N23422);
or OR3 (N23593, N23590, N15142, N18308);
not NOT1 (N23594, N23586);
or OR3 (N23595, N23588, N12888, N11402);
and AND4 (N23596, N23594, N23494, N7999, N9464);
buf BUF1 (N23597, N23582);
nor NOR4 (N23598, N23596, N22542, N867, N2958);
buf BUF1 (N23599, N23585);
and AND4 (N23600, N23584, N16714, N18924, N9242);
buf BUF1 (N23601, N23589);
not NOT1 (N23602, N23598);
or OR2 (N23603, N23595, N22558);
xor XOR2 (N23604, N23597, N12880);
xor XOR2 (N23605, N23600, N16925);
or OR2 (N23606, N23603, N13278);
and AND2 (N23607, N23604, N21226);
nand NAND2 (N23608, N23593, N2264);
buf BUF1 (N23609, N23579);
or OR2 (N23610, N23602, N3309);
not NOT1 (N23611, N23592);
xor XOR2 (N23612, N23576, N3736);
or OR4 (N23613, N23610, N20234, N17871, N20932);
or OR3 (N23614, N23611, N14278, N14861);
not NOT1 (N23615, N23601);
nor NOR3 (N23616, N23606, N11887, N9493);
or OR2 (N23617, N23599, N10561);
and AND3 (N23618, N23609, N865, N8044);
xor XOR2 (N23619, N23614, N21446);
buf BUF1 (N23620, N23617);
xor XOR2 (N23621, N23607, N11246);
buf BUF1 (N23622, N23615);
nand NAND2 (N23623, N23605, N15866);
and AND4 (N23624, N23620, N3517, N11004, N16837);
not NOT1 (N23625, N23621);
not NOT1 (N23626, N23622);
not NOT1 (N23627, N23618);
or OR2 (N23628, N23608, N48);
xor XOR2 (N23629, N23626, N16312);
xor XOR2 (N23630, N23613, N9261);
buf BUF1 (N23631, N23627);
not NOT1 (N23632, N23623);
xor XOR2 (N23633, N23630, N9908);
not NOT1 (N23634, N23616);
or OR3 (N23635, N23634, N4457, N12587);
or OR4 (N23636, N23619, N2868, N23412, N3296);
xor XOR2 (N23637, N23629, N5290);
xor XOR2 (N23638, N23633, N22068);
and AND2 (N23639, N23628, N23417);
or OR2 (N23640, N23636, N3031);
not NOT1 (N23641, N23635);
nor NOR4 (N23642, N23632, N17476, N23287, N2095);
nor NOR3 (N23643, N23631, N2741, N5299);
buf BUF1 (N23644, N23625);
nand NAND2 (N23645, N23612, N9331);
nand NAND2 (N23646, N23640, N2594);
buf BUF1 (N23647, N23641);
nand NAND2 (N23648, N23645, N1150);
not NOT1 (N23649, N23644);
and AND2 (N23650, N23637, N21317);
xor XOR2 (N23651, N23648, N21056);
not NOT1 (N23652, N23643);
buf BUF1 (N23653, N23646);
nor NOR2 (N23654, N23649, N8860);
buf BUF1 (N23655, N23639);
and AND2 (N23656, N23652, N14235);
nor NOR4 (N23657, N23650, N3396, N16437, N5393);
not NOT1 (N23658, N23653);
nand NAND2 (N23659, N23657, N11779);
not NOT1 (N23660, N23654);
and AND3 (N23661, N23655, N16048, N1077);
or OR4 (N23662, N23656, N892, N6814, N23583);
and AND2 (N23663, N23638, N5058);
xor XOR2 (N23664, N23661, N13379);
not NOT1 (N23665, N23647);
nand NAND3 (N23666, N23659, N12555, N8605);
xor XOR2 (N23667, N23660, N17985);
xor XOR2 (N23668, N23666, N13515);
xor XOR2 (N23669, N23651, N18626);
not NOT1 (N23670, N23658);
nand NAND4 (N23671, N23665, N13555, N950, N11478);
and AND2 (N23672, N23670, N1066);
xor XOR2 (N23673, N23663, N19087);
nand NAND4 (N23674, N23673, N6286, N9827, N23013);
nor NOR2 (N23675, N23669, N16019);
nand NAND3 (N23676, N23642, N12007, N1563);
buf BUF1 (N23677, N23676);
nand NAND4 (N23678, N23671, N17361, N10395, N8600);
not NOT1 (N23679, N23668);
nor NOR2 (N23680, N23667, N6433);
xor XOR2 (N23681, N23678, N10049);
buf BUF1 (N23682, N23675);
not NOT1 (N23683, N23662);
not NOT1 (N23684, N23680);
nor NOR2 (N23685, N23681, N11459);
xor XOR2 (N23686, N23684, N6859);
nand NAND3 (N23687, N23664, N13402, N12087);
buf BUF1 (N23688, N23682);
nor NOR3 (N23689, N23683, N17000, N17454);
nor NOR3 (N23690, N23679, N19718, N7502);
and AND4 (N23691, N23688, N11596, N14696, N7536);
xor XOR2 (N23692, N23672, N502);
and AND2 (N23693, N23689, N9850);
nand NAND2 (N23694, N23624, N10253);
or OR4 (N23695, N23686, N17830, N17749, N4427);
not NOT1 (N23696, N23692);
buf BUF1 (N23697, N23677);
nor NOR2 (N23698, N23674, N7335);
nand NAND3 (N23699, N23698, N1992, N22696);
and AND2 (N23700, N23697, N8685);
xor XOR2 (N23701, N23690, N13347);
nand NAND4 (N23702, N23691, N15421, N23310, N10540);
buf BUF1 (N23703, N23696);
or OR2 (N23704, N23687, N13952);
or OR4 (N23705, N23700, N22583, N40, N21714);
not NOT1 (N23706, N23701);
nand NAND4 (N23707, N23685, N11241, N1421, N9960);
nor NOR4 (N23708, N23706, N17637, N12174, N6875);
xor XOR2 (N23709, N23703, N3199);
xor XOR2 (N23710, N23705, N987);
nor NOR3 (N23711, N23695, N22778, N15102);
or OR3 (N23712, N23709, N1388, N20561);
not NOT1 (N23713, N23704);
or OR3 (N23714, N23702, N14044, N3474);
and AND4 (N23715, N23694, N6518, N9017, N6889);
or OR4 (N23716, N23699, N18226, N11432, N18438);
or OR2 (N23717, N23713, N16219);
nor NOR3 (N23718, N23711, N1814, N4966);
and AND2 (N23719, N23708, N8939);
xor XOR2 (N23720, N23710, N20956);
not NOT1 (N23721, N23714);
nand NAND2 (N23722, N23719, N14535);
and AND4 (N23723, N23712, N23171, N3031, N4146);
not NOT1 (N23724, N23722);
and AND4 (N23725, N23715, N14847, N7056, N21144);
buf BUF1 (N23726, N23720);
and AND4 (N23727, N23721, N22925, N13481, N16690);
or OR3 (N23728, N23724, N14226, N21113);
buf BUF1 (N23729, N23716);
xor XOR2 (N23730, N23723, N5463);
nand NAND4 (N23731, N23718, N21590, N6152, N9975);
and AND3 (N23732, N23725, N22052, N4753);
not NOT1 (N23733, N23727);
nand NAND2 (N23734, N23717, N13510);
nor NOR4 (N23735, N23728, N18407, N15948, N14180);
and AND2 (N23736, N23729, N11778);
nor NOR2 (N23737, N23734, N9488);
not NOT1 (N23738, N23737);
nand NAND3 (N23739, N23733, N2769, N11211);
nor NOR2 (N23740, N23730, N19712);
nor NOR4 (N23741, N23736, N703, N1500, N16189);
and AND3 (N23742, N23739, N12373, N5245);
buf BUF1 (N23743, N23732);
and AND4 (N23744, N23693, N8290, N2321, N4914);
or OR4 (N23745, N23731, N7124, N6947, N15498);
not NOT1 (N23746, N23744);
xor XOR2 (N23747, N23735, N15256);
nand NAND4 (N23748, N23740, N1876, N10314, N17256);
not NOT1 (N23749, N23742);
buf BUF1 (N23750, N23738);
or OR3 (N23751, N23747, N13495, N4936);
xor XOR2 (N23752, N23743, N153);
and AND2 (N23753, N23751, N4931);
xor XOR2 (N23754, N23750, N6785);
not NOT1 (N23755, N23746);
or OR3 (N23756, N23748, N13893, N23657);
buf BUF1 (N23757, N23749);
xor XOR2 (N23758, N23757, N9380);
nand NAND3 (N23759, N23756, N19823, N11908);
not NOT1 (N23760, N23745);
buf BUF1 (N23761, N23752);
and AND3 (N23762, N23758, N5548, N8631);
and AND4 (N23763, N23760, N15054, N146, N9657);
or OR2 (N23764, N23759, N16518);
not NOT1 (N23765, N23726);
buf BUF1 (N23766, N23761);
or OR2 (N23767, N23754, N22569);
nor NOR4 (N23768, N23755, N22415, N14614, N21264);
nand NAND3 (N23769, N23741, N14243, N17723);
or OR2 (N23770, N23767, N3625);
xor XOR2 (N23771, N23768, N5210);
nand NAND3 (N23772, N23707, N17757, N18340);
nand NAND3 (N23773, N23769, N7799, N14122);
buf BUF1 (N23774, N23764);
and AND2 (N23775, N23762, N2514);
buf BUF1 (N23776, N23771);
not NOT1 (N23777, N23776);
xor XOR2 (N23778, N23753, N20129);
nand NAND4 (N23779, N23770, N1596, N19265, N18075);
and AND2 (N23780, N23766, N23778);
nand NAND4 (N23781, N1353, N14065, N17492, N16129);
xor XOR2 (N23782, N23765, N13095);
not NOT1 (N23783, N23782);
or OR4 (N23784, N23772, N771, N1257, N6105);
nor NOR3 (N23785, N23780, N11548, N14248);
or OR3 (N23786, N23783, N18027, N15340);
xor XOR2 (N23787, N23774, N13250);
buf BUF1 (N23788, N23763);
not NOT1 (N23789, N23786);
and AND4 (N23790, N23779, N8402, N17986, N18574);
and AND4 (N23791, N23785, N4543, N10662, N15253);
and AND4 (N23792, N23781, N13192, N8658, N16633);
not NOT1 (N23793, N23791);
nor NOR2 (N23794, N23787, N2373);
xor XOR2 (N23795, N23788, N7080);
nand NAND3 (N23796, N23794, N1651, N4578);
nand NAND4 (N23797, N23795, N3268, N5448, N22585);
and AND2 (N23798, N23797, N9375);
or OR3 (N23799, N23789, N11926, N12653);
nand NAND2 (N23800, N23792, N8791);
nor NOR2 (N23801, N23790, N3434);
nand NAND2 (N23802, N23784, N21676);
or OR4 (N23803, N23777, N23572, N10528, N8308);
xor XOR2 (N23804, N23802, N4419);
buf BUF1 (N23805, N23793);
nand NAND4 (N23806, N23773, N1181, N19608, N15584);
and AND2 (N23807, N23806, N7687);
and AND2 (N23808, N23800, N10346);
nor NOR2 (N23809, N23804, N1029);
not NOT1 (N23810, N23796);
or OR4 (N23811, N23809, N16921, N23082, N15830);
nand NAND3 (N23812, N23807, N10895, N12179);
xor XOR2 (N23813, N23799, N23424);
buf BUF1 (N23814, N23808);
nor NOR2 (N23815, N23803, N720);
buf BUF1 (N23816, N23805);
not NOT1 (N23817, N23812);
not NOT1 (N23818, N23817);
nor NOR2 (N23819, N23798, N23626);
and AND2 (N23820, N23813, N3838);
nor NOR4 (N23821, N23820, N21919, N10940, N21321);
and AND3 (N23822, N23819, N8757, N481);
not NOT1 (N23823, N23815);
nor NOR2 (N23824, N23823, N15665);
buf BUF1 (N23825, N23816);
nand NAND4 (N23826, N23825, N23022, N9411, N2524);
and AND2 (N23827, N23824, N14751);
and AND2 (N23828, N23822, N12533);
nand NAND2 (N23829, N23811, N2141);
and AND4 (N23830, N23818, N22769, N2595, N13184);
nand NAND2 (N23831, N23810, N4499);
xor XOR2 (N23832, N23828, N1906);
or OR3 (N23833, N23832, N6746, N10148);
nand NAND2 (N23834, N23814, N532);
or OR3 (N23835, N23831, N5850, N8366);
buf BUF1 (N23836, N23833);
or OR3 (N23837, N23835, N8764, N7534);
nand NAND3 (N23838, N23829, N12009, N5914);
not NOT1 (N23839, N23801);
or OR4 (N23840, N23830, N5322, N13766, N1784);
not NOT1 (N23841, N23821);
and AND2 (N23842, N23836, N16158);
or OR4 (N23843, N23775, N11853, N21057, N12143);
or OR4 (N23844, N23834, N11112, N527, N19131);
nor NOR2 (N23845, N23826, N2746);
not NOT1 (N23846, N23840);
and AND3 (N23847, N23845, N19642, N9572);
xor XOR2 (N23848, N23827, N22885);
or OR3 (N23849, N23843, N13706, N18762);
nor NOR3 (N23850, N23847, N13584, N16036);
buf BUF1 (N23851, N23844);
nand NAND4 (N23852, N23841, N17645, N20388, N20414);
not NOT1 (N23853, N23839);
nand NAND2 (N23854, N23838, N2739);
nand NAND3 (N23855, N23842, N1243, N3452);
or OR4 (N23856, N23852, N5347, N5316, N11772);
buf BUF1 (N23857, N23855);
nand NAND4 (N23858, N23850, N722, N1878, N22423);
xor XOR2 (N23859, N23851, N7353);
buf BUF1 (N23860, N23854);
nor NOR4 (N23861, N23857, N21339, N1181, N195);
and AND3 (N23862, N23846, N1167, N17940);
buf BUF1 (N23863, N23856);
xor XOR2 (N23864, N23853, N15450);
nor NOR4 (N23865, N23861, N15637, N4264, N1469);
not NOT1 (N23866, N23864);
or OR4 (N23867, N23837, N17919, N17018, N8794);
buf BUF1 (N23868, N23849);
nor NOR4 (N23869, N23860, N5354, N10832, N17567);
buf BUF1 (N23870, N23869);
nand NAND2 (N23871, N23867, N7435);
or OR2 (N23872, N23866, N23699);
or OR3 (N23873, N23859, N20969, N17060);
and AND4 (N23874, N23868, N10369, N203, N2893);
xor XOR2 (N23875, N23870, N12358);
and AND3 (N23876, N23873, N17862, N19409);
nor NOR3 (N23877, N23876, N3557, N4980);
buf BUF1 (N23878, N23848);
or OR4 (N23879, N23871, N2366, N18603, N6468);
buf BUF1 (N23880, N23862);
not NOT1 (N23881, N23875);
nor NOR3 (N23882, N23877, N15517, N18088);
or OR3 (N23883, N23872, N12875, N3098);
nor NOR4 (N23884, N23879, N33, N17892, N19087);
xor XOR2 (N23885, N23884, N20318);
nand NAND2 (N23886, N23878, N2078);
nor NOR2 (N23887, N23883, N7465);
nand NAND4 (N23888, N23865, N3895, N19455, N7612);
xor XOR2 (N23889, N23882, N5598);
xor XOR2 (N23890, N23885, N1014);
and AND4 (N23891, N23881, N19678, N19994, N20347);
not NOT1 (N23892, N23888);
and AND4 (N23893, N23892, N9373, N14511, N11823);
buf BUF1 (N23894, N23887);
xor XOR2 (N23895, N23893, N16663);
buf BUF1 (N23896, N23886);
not NOT1 (N23897, N23890);
and AND2 (N23898, N23894, N9838);
buf BUF1 (N23899, N23895);
nand NAND3 (N23900, N23874, N9252, N23843);
not NOT1 (N23901, N23880);
and AND3 (N23902, N23858, N14491, N7607);
and AND2 (N23903, N23897, N1889);
nor NOR4 (N23904, N23891, N3214, N10461, N13318);
not NOT1 (N23905, N23896);
nor NOR2 (N23906, N23902, N22569);
not NOT1 (N23907, N23905);
buf BUF1 (N23908, N23901);
nand NAND2 (N23909, N23908, N8498);
nand NAND2 (N23910, N23903, N19608);
buf BUF1 (N23911, N23906);
buf BUF1 (N23912, N23900);
nor NOR2 (N23913, N23904, N19251);
nand NAND2 (N23914, N23899, N22191);
and AND4 (N23915, N23889, N21242, N1133, N7889);
buf BUF1 (N23916, N23913);
or OR4 (N23917, N23915, N17485, N14132, N23898);
and AND4 (N23918, N15042, N2514, N15042, N10495);
and AND4 (N23919, N23907, N3552, N10689, N11371);
nand NAND2 (N23920, N23919, N17642);
or OR2 (N23921, N23909, N8117);
xor XOR2 (N23922, N23912, N22599);
nor NOR3 (N23923, N23921, N15289, N16185);
xor XOR2 (N23924, N23911, N243);
xor XOR2 (N23925, N23863, N472);
xor XOR2 (N23926, N23918, N20384);
nor NOR4 (N23927, N23917, N4077, N23258, N16278);
buf BUF1 (N23928, N23923);
nor NOR4 (N23929, N23925, N23248, N2192, N1647);
or OR2 (N23930, N23914, N9675);
buf BUF1 (N23931, N23922);
xor XOR2 (N23932, N23920, N4682);
or OR4 (N23933, N23924, N9163, N1120, N2695);
and AND4 (N23934, N23910, N6691, N12584, N20086);
not NOT1 (N23935, N23916);
nand NAND2 (N23936, N23931, N17);
not NOT1 (N23937, N23935);
nor NOR4 (N23938, N23928, N22456, N18772, N13080);
and AND4 (N23939, N23933, N8690, N9889, N6145);
buf BUF1 (N23940, N23939);
not NOT1 (N23941, N23929);
and AND3 (N23942, N23938, N13931, N18761);
nand NAND2 (N23943, N23940, N22535);
xor XOR2 (N23944, N23942, N18001);
xor XOR2 (N23945, N23941, N4424);
nor NOR3 (N23946, N23934, N4502, N18839);
nor NOR4 (N23947, N23930, N21445, N17288, N11886);
nand NAND3 (N23948, N23937, N3895, N7230);
not NOT1 (N23949, N23926);
buf BUF1 (N23950, N23927);
not NOT1 (N23951, N23943);
and AND3 (N23952, N23944, N15634, N10268);
nand NAND2 (N23953, N23936, N15725);
xor XOR2 (N23954, N23948, N15530);
buf BUF1 (N23955, N23952);
or OR2 (N23956, N23946, N6194);
and AND3 (N23957, N23947, N7780, N12964);
not NOT1 (N23958, N23932);
or OR4 (N23959, N23945, N15395, N6992, N18767);
and AND2 (N23960, N23953, N20951);
not NOT1 (N23961, N23956);
or OR4 (N23962, N23961, N21347, N21711, N14415);
nand NAND3 (N23963, N23957, N12283, N23071);
nor NOR4 (N23964, N23949, N532, N2715, N5137);
buf BUF1 (N23965, N23959);
buf BUF1 (N23966, N23963);
xor XOR2 (N23967, N23960, N3561);
buf BUF1 (N23968, N23950);
xor XOR2 (N23969, N23954, N8790);
and AND2 (N23970, N23955, N14166);
not NOT1 (N23971, N23969);
buf BUF1 (N23972, N23968);
not NOT1 (N23973, N23965);
nor NOR3 (N23974, N23964, N12158, N8559);
xor XOR2 (N23975, N23971, N23681);
and AND4 (N23976, N23958, N951, N2345, N2749);
and AND4 (N23977, N23973, N23675, N15005, N15458);
xor XOR2 (N23978, N23976, N16687);
buf BUF1 (N23979, N23970);
not NOT1 (N23980, N23962);
nand NAND4 (N23981, N23951, N23943, N6088, N18390);
nor NOR3 (N23982, N23980, N23806, N2902);
or OR3 (N23983, N23979, N373, N18192);
nand NAND4 (N23984, N23967, N15590, N7601, N16568);
xor XOR2 (N23985, N23966, N19299);
not NOT1 (N23986, N23982);
and AND4 (N23987, N23984, N21572, N6177, N5967);
or OR2 (N23988, N23983, N21509);
xor XOR2 (N23989, N23978, N2185);
or OR3 (N23990, N23975, N9062, N23664);
or OR2 (N23991, N23981, N17366);
nor NOR2 (N23992, N23988, N13137);
not NOT1 (N23993, N23991);
buf BUF1 (N23994, N23986);
not NOT1 (N23995, N23987);
buf BUF1 (N23996, N23990);
nor NOR2 (N23997, N23993, N23350);
and AND3 (N23998, N23992, N11762, N13866);
xor XOR2 (N23999, N23997, N22427);
or OR4 (N24000, N23994, N8714, N6616, N19905);
or OR2 (N24001, N23974, N2809);
xor XOR2 (N24002, N23977, N1445);
nand NAND2 (N24003, N23996, N13057);
buf BUF1 (N24004, N23999);
xor XOR2 (N24005, N23998, N22369);
and AND4 (N24006, N23995, N19128, N10408, N414);
not NOT1 (N24007, N24001);
nand NAND3 (N24008, N23989, N22404, N11855);
not NOT1 (N24009, N23972);
and AND3 (N24010, N24007, N7984, N13551);
nand NAND4 (N24011, N23985, N597, N6425, N10697);
xor XOR2 (N24012, N24009, N5585);
xor XOR2 (N24013, N24012, N5056);
or OR2 (N24014, N24000, N14540);
buf BUF1 (N24015, N24003);
xor XOR2 (N24016, N24006, N131);
or OR2 (N24017, N24014, N6328);
nor NOR4 (N24018, N24008, N22621, N11020, N9140);
and AND3 (N24019, N24015, N10639, N8470);
nand NAND3 (N24020, N24018, N16553, N4763);
or OR3 (N24021, N24020, N2712, N11573);
nor NOR3 (N24022, N24017, N9008, N19589);
not NOT1 (N24023, N24011);
not NOT1 (N24024, N24010);
buf BUF1 (N24025, N24023);
xor XOR2 (N24026, N24022, N16126);
nor NOR2 (N24027, N24021, N2861);
nand NAND4 (N24028, N24002, N23616, N2192, N5291);
nand NAND3 (N24029, N24026, N19123, N23856);
buf BUF1 (N24030, N24004);
and AND3 (N24031, N24028, N18181, N8972);
xor XOR2 (N24032, N24027, N21775);
nor NOR2 (N24033, N24031, N17704);
xor XOR2 (N24034, N24013, N18449);
and AND2 (N24035, N24030, N21943);
and AND4 (N24036, N24016, N20807, N17450, N6812);
buf BUF1 (N24037, N24029);
nor NOR4 (N24038, N24024, N3958, N9897, N15394);
buf BUF1 (N24039, N24033);
buf BUF1 (N24040, N24025);
nand NAND3 (N24041, N24034, N22638, N21863);
xor XOR2 (N24042, N24037, N10720);
nor NOR2 (N24043, N24040, N8120);
and AND4 (N24044, N24005, N2888, N6240, N3044);
buf BUF1 (N24045, N24036);
not NOT1 (N24046, N24035);
or OR4 (N24047, N24043, N18378, N16800, N2825);
and AND3 (N24048, N24039, N3840, N846);
or OR3 (N24049, N24047, N15900, N11864);
nor NOR2 (N24050, N24044, N20437);
nor NOR3 (N24051, N24049, N6311, N1025);
or OR3 (N24052, N24038, N20958, N22127);
nor NOR3 (N24053, N24041, N3602, N17711);
and AND3 (N24054, N24032, N15893, N13501);
buf BUF1 (N24055, N24053);
nand NAND3 (N24056, N24046, N23327, N19896);
or OR4 (N24057, N24019, N18756, N11319, N19079);
or OR4 (N24058, N24048, N18707, N3066, N3566);
or OR2 (N24059, N24056, N6438);
nor NOR2 (N24060, N24057, N22328);
nor NOR3 (N24061, N24059, N16929, N4264);
and AND2 (N24062, N24050, N12532);
nand NAND4 (N24063, N24055, N9618, N14096, N14875);
nand NAND4 (N24064, N24063, N20604, N1123, N13243);
xor XOR2 (N24065, N24064, N5186);
xor XOR2 (N24066, N24058, N11091);
nand NAND3 (N24067, N24066, N19424, N6549);
buf BUF1 (N24068, N24042);
nor NOR3 (N24069, N24062, N10796, N9498);
or OR2 (N24070, N24051, N21715);
xor XOR2 (N24071, N24068, N10674);
or OR2 (N24072, N24067, N16764);
buf BUF1 (N24073, N24054);
nand NAND2 (N24074, N24052, N4687);
not NOT1 (N24075, N24071);
nand NAND3 (N24076, N24061, N15413, N3839);
nor NOR3 (N24077, N24074, N5223, N22623);
not NOT1 (N24078, N24077);
xor XOR2 (N24079, N24069, N12699);
buf BUF1 (N24080, N24073);
buf BUF1 (N24081, N24060);
not NOT1 (N24082, N24075);
buf BUF1 (N24083, N24065);
nand NAND4 (N24084, N24045, N4725, N10895, N19703);
not NOT1 (N24085, N24083);
not NOT1 (N24086, N24084);
nor NOR3 (N24087, N24078, N20254, N2527);
buf BUF1 (N24088, N24079);
or OR3 (N24089, N24085, N12031, N14884);
xor XOR2 (N24090, N24080, N6034);
nor NOR2 (N24091, N24072, N3954);
buf BUF1 (N24092, N24091);
xor XOR2 (N24093, N24092, N18031);
not NOT1 (N24094, N24089);
and AND2 (N24095, N24094, N673);
nand NAND4 (N24096, N24093, N12789, N13298, N12330);
xor XOR2 (N24097, N24087, N14605);
not NOT1 (N24098, N24086);
buf BUF1 (N24099, N24095);
or OR3 (N24100, N24099, N8251, N2148);
and AND2 (N24101, N24096, N3966);
nor NOR3 (N24102, N24090, N951, N1829);
and AND3 (N24103, N24097, N6362, N23310);
nand NAND4 (N24104, N24076, N4282, N14680, N3460);
or OR2 (N24105, N24088, N19440);
nand NAND3 (N24106, N24101, N20846, N14957);
xor XOR2 (N24107, N24082, N13928);
nor NOR3 (N24108, N24102, N13207, N2129);
xor XOR2 (N24109, N24104, N20518);
nand NAND4 (N24110, N24081, N6716, N10048, N2012);
and AND2 (N24111, N24105, N6358);
and AND2 (N24112, N24109, N11770);
or OR2 (N24113, N24110, N2720);
and AND2 (N24114, N24070, N10699);
not NOT1 (N24115, N24103);
and AND4 (N24116, N24107, N8443, N18619, N22636);
xor XOR2 (N24117, N24115, N21815);
and AND4 (N24118, N24113, N14800, N23456, N1490);
or OR3 (N24119, N24117, N15159, N5015);
not NOT1 (N24120, N24114);
nor NOR2 (N24121, N24112, N11833);
not NOT1 (N24122, N24100);
xor XOR2 (N24123, N24120, N5536);
nor NOR2 (N24124, N24098, N14017);
xor XOR2 (N24125, N24108, N21830);
not NOT1 (N24126, N24125);
xor XOR2 (N24127, N24124, N6305);
or OR3 (N24128, N24106, N3858, N7601);
xor XOR2 (N24129, N24111, N21797);
nor NOR3 (N24130, N24126, N6308, N2784);
buf BUF1 (N24131, N24121);
not NOT1 (N24132, N24116);
buf BUF1 (N24133, N24122);
xor XOR2 (N24134, N24131, N11296);
not NOT1 (N24135, N24134);
nand NAND3 (N24136, N24132, N19864, N660);
nand NAND3 (N24137, N24130, N13087, N21474);
and AND4 (N24138, N24137, N3676, N2219, N11300);
xor XOR2 (N24139, N24118, N3635);
buf BUF1 (N24140, N24135);
not NOT1 (N24141, N24139);
not NOT1 (N24142, N24133);
and AND3 (N24143, N24138, N10884, N8165);
and AND2 (N24144, N24141, N7985);
buf BUF1 (N24145, N24140);
or OR4 (N24146, N24128, N20269, N8876, N14635);
xor XOR2 (N24147, N24123, N2218);
and AND2 (N24148, N24119, N1208);
and AND4 (N24149, N24146, N15327, N12504, N8873);
not NOT1 (N24150, N24127);
buf BUF1 (N24151, N24143);
not NOT1 (N24152, N24151);
nand NAND4 (N24153, N24149, N7245, N4248, N5662);
xor XOR2 (N24154, N24152, N23977);
nor NOR2 (N24155, N24147, N18770);
nor NOR3 (N24156, N24145, N11536, N14641);
nor NOR2 (N24157, N24155, N9083);
buf BUF1 (N24158, N24142);
and AND4 (N24159, N24153, N761, N23445, N20881);
nand NAND3 (N24160, N24144, N10230, N2511);
buf BUF1 (N24161, N24129);
nor NOR4 (N24162, N24159, N9494, N4581, N3720);
not NOT1 (N24163, N24148);
xor XOR2 (N24164, N24158, N10806);
buf BUF1 (N24165, N24157);
nor NOR2 (N24166, N24165, N5384);
not NOT1 (N24167, N24164);
buf BUF1 (N24168, N24150);
and AND3 (N24169, N24168, N12264, N17721);
not NOT1 (N24170, N24160);
or OR2 (N24171, N24161, N24115);
or OR3 (N24172, N24136, N17406, N18222);
and AND4 (N24173, N24163, N10277, N10716, N22739);
nor NOR3 (N24174, N24173, N8979, N3340);
or OR3 (N24175, N24170, N19603, N9590);
nand NAND2 (N24176, N24175, N22444);
not NOT1 (N24177, N24167);
and AND3 (N24178, N24171, N10008, N4754);
buf BUF1 (N24179, N24162);
and AND4 (N24180, N24176, N15892, N15606, N17954);
not NOT1 (N24181, N24178);
not NOT1 (N24182, N24166);
or OR4 (N24183, N24154, N12098, N24033, N5588);
nor NOR3 (N24184, N24179, N5760, N18178);
nor NOR3 (N24185, N24184, N2894, N15249);
and AND4 (N24186, N24169, N8158, N3339, N4818);
or OR4 (N24187, N24183, N11321, N23224, N13108);
or OR2 (N24188, N24186, N20335);
or OR2 (N24189, N24181, N14490);
xor XOR2 (N24190, N24177, N4242);
xor XOR2 (N24191, N24187, N5277);
and AND3 (N24192, N24189, N18698, N7851);
and AND3 (N24193, N24185, N14857, N23686);
nand NAND2 (N24194, N24192, N8814);
and AND3 (N24195, N24194, N12150, N18204);
or OR2 (N24196, N24193, N12526);
or OR2 (N24197, N24195, N4096);
xor XOR2 (N24198, N24190, N9958);
xor XOR2 (N24199, N24197, N7827);
and AND2 (N24200, N24191, N3166);
xor XOR2 (N24201, N24200, N7214);
or OR3 (N24202, N24198, N9714, N194);
nor NOR3 (N24203, N24199, N6559, N2464);
and AND2 (N24204, N24156, N16126);
not NOT1 (N24205, N24196);
or OR2 (N24206, N24172, N13282);
nand NAND4 (N24207, N24202, N9023, N16575, N7092);
and AND4 (N24208, N24204, N20260, N14257, N1494);
not NOT1 (N24209, N24180);
xor XOR2 (N24210, N24182, N6305);
xor XOR2 (N24211, N24208, N16725);
nor NOR3 (N24212, N24201, N18256, N10874);
buf BUF1 (N24213, N24188);
buf BUF1 (N24214, N24209);
xor XOR2 (N24215, N24211, N13991);
nand NAND2 (N24216, N24214, N4854);
buf BUF1 (N24217, N24207);
and AND2 (N24218, N24216, N23568);
not NOT1 (N24219, N24203);
buf BUF1 (N24220, N24205);
or OR4 (N24221, N24210, N18486, N18178, N24155);
nand NAND4 (N24222, N24215, N12418, N21581, N18893);
not NOT1 (N24223, N24174);
xor XOR2 (N24224, N24220, N8748);
nand NAND3 (N24225, N24217, N15092, N21770);
buf BUF1 (N24226, N24206);
not NOT1 (N24227, N24218);
buf BUF1 (N24228, N24225);
or OR4 (N24229, N24213, N17438, N8927, N1989);
nor NOR3 (N24230, N24212, N7816, N10531);
nor NOR2 (N24231, N24223, N20098);
nor NOR3 (N24232, N24221, N20070, N17247);
or OR2 (N24233, N24228, N23544);
and AND3 (N24234, N24224, N22559, N6069);
buf BUF1 (N24235, N24222);
and AND3 (N24236, N24233, N3027, N2182);
or OR4 (N24237, N24232, N6033, N9607, N8492);
nand NAND2 (N24238, N24226, N17848);
not NOT1 (N24239, N24237);
and AND4 (N24240, N24231, N17431, N16854, N19923);
not NOT1 (N24241, N24239);
buf BUF1 (N24242, N24227);
not NOT1 (N24243, N24219);
nand NAND2 (N24244, N24234, N16394);
and AND4 (N24245, N24243, N12189, N13146, N22041);
xor XOR2 (N24246, N24229, N12875);
buf BUF1 (N24247, N24230);
buf BUF1 (N24248, N24244);
nor NOR4 (N24249, N24238, N15634, N9846, N10064);
not NOT1 (N24250, N24242);
buf BUF1 (N24251, N24249);
nand NAND2 (N24252, N24235, N19461);
and AND3 (N24253, N24251, N15203, N7220);
not NOT1 (N24254, N24236);
and AND4 (N24255, N24247, N8513, N15195, N19503);
buf BUF1 (N24256, N24254);
nor NOR2 (N24257, N24253, N11954);
and AND4 (N24258, N24245, N19436, N17116, N14077);
xor XOR2 (N24259, N24252, N462);
and AND2 (N24260, N24258, N8300);
and AND4 (N24261, N24255, N2347, N17682, N14997);
buf BUF1 (N24262, N24257);
nand NAND3 (N24263, N24250, N22375, N8959);
nand NAND3 (N24264, N24241, N16182, N24078);
buf BUF1 (N24265, N24240);
and AND4 (N24266, N24256, N17879, N1786, N8786);
nand NAND4 (N24267, N24264, N6090, N15000, N14828);
not NOT1 (N24268, N24248);
buf BUF1 (N24269, N24246);
and AND3 (N24270, N24267, N8195, N8841);
or OR2 (N24271, N24259, N6391);
and AND4 (N24272, N24271, N3059, N9651, N14039);
xor XOR2 (N24273, N24266, N17091);
and AND4 (N24274, N24261, N23958, N19033, N1692);
nor NOR2 (N24275, N24273, N11798);
nand NAND4 (N24276, N24260, N8987, N13201, N18023);
nor NOR4 (N24277, N24275, N11730, N280, N8684);
xor XOR2 (N24278, N24268, N23831);
nand NAND3 (N24279, N24278, N22781, N285);
nand NAND2 (N24280, N24265, N10716);
or OR3 (N24281, N24263, N2133, N3499);
xor XOR2 (N24282, N24276, N16746);
xor XOR2 (N24283, N24272, N16913);
buf BUF1 (N24284, N24270);
buf BUF1 (N24285, N24269);
buf BUF1 (N24286, N24281);
and AND4 (N24287, N24285, N129, N23070, N16820);
or OR3 (N24288, N24283, N19472, N23538);
nor NOR3 (N24289, N24274, N966, N4215);
nand NAND4 (N24290, N24287, N997, N12726, N17286);
xor XOR2 (N24291, N24288, N275);
nand NAND2 (N24292, N24262, N18150);
not NOT1 (N24293, N24280);
not NOT1 (N24294, N24286);
nor NOR3 (N24295, N24289, N9453, N23843);
not NOT1 (N24296, N24282);
and AND2 (N24297, N24295, N13003);
buf BUF1 (N24298, N24296);
and AND4 (N24299, N24294, N11483, N14571, N15968);
nand NAND3 (N24300, N24292, N5787, N9347);
buf BUF1 (N24301, N24279);
nor NOR4 (N24302, N24291, N12673, N16813, N2335);
not NOT1 (N24303, N24300);
not NOT1 (N24304, N24303);
buf BUF1 (N24305, N24297);
and AND4 (N24306, N24284, N15250, N18740, N16613);
or OR4 (N24307, N24293, N552, N15808, N21428);
not NOT1 (N24308, N24307);
and AND4 (N24309, N24301, N17265, N14618, N6744);
xor XOR2 (N24310, N24277, N3779);
or OR4 (N24311, N24308, N19062, N1172, N3257);
not NOT1 (N24312, N24299);
xor XOR2 (N24313, N24304, N21620);
not NOT1 (N24314, N24313);
xor XOR2 (N24315, N24311, N9870);
buf BUF1 (N24316, N24315);
buf BUF1 (N24317, N24310);
nor NOR2 (N24318, N24298, N24211);
not NOT1 (N24319, N24314);
not NOT1 (N24320, N24316);
not NOT1 (N24321, N24312);
nand NAND4 (N24322, N24290, N23968, N2244, N19777);
not NOT1 (N24323, N24318);
buf BUF1 (N24324, N24306);
buf BUF1 (N24325, N24309);
xor XOR2 (N24326, N24321, N22581);
not NOT1 (N24327, N24322);
and AND3 (N24328, N24319, N6755, N11643);
xor XOR2 (N24329, N24323, N19515);
nor NOR3 (N24330, N24324, N15293, N9466);
buf BUF1 (N24331, N24328);
and AND3 (N24332, N24326, N739, N21111);
or OR2 (N24333, N24330, N5885);
not NOT1 (N24334, N24305);
nor NOR3 (N24335, N24334, N330, N11722);
nor NOR4 (N24336, N24335, N9505, N13771, N23766);
xor XOR2 (N24337, N24317, N19124);
xor XOR2 (N24338, N24336, N5274);
or OR2 (N24339, N24331, N468);
buf BUF1 (N24340, N24329);
and AND4 (N24341, N24337, N8541, N9427, N18545);
xor XOR2 (N24342, N24338, N9210);
buf BUF1 (N24343, N24332);
nand NAND2 (N24344, N24340, N3099);
not NOT1 (N24345, N24342);
and AND2 (N24346, N24341, N7991);
nor NOR4 (N24347, N24325, N12367, N14357, N24183);
or OR3 (N24348, N24346, N7296, N21213);
buf BUF1 (N24349, N24302);
nand NAND2 (N24350, N24339, N22360);
buf BUF1 (N24351, N24350);
buf BUF1 (N24352, N24344);
xor XOR2 (N24353, N24345, N23676);
nor NOR2 (N24354, N24352, N23152);
and AND4 (N24355, N24327, N16265, N23409, N3315);
xor XOR2 (N24356, N24355, N20570);
nand NAND4 (N24357, N24343, N8347, N12334, N18058);
buf BUF1 (N24358, N24356);
not NOT1 (N24359, N24320);
and AND2 (N24360, N24333, N20425);
and AND3 (N24361, N24359, N11471, N5380);
and AND2 (N24362, N24353, N22799);
xor XOR2 (N24363, N24348, N1478);
or OR2 (N24364, N24351, N21763);
or OR3 (N24365, N24354, N6196, N5745);
and AND4 (N24366, N24362, N2773, N6503, N5613);
not NOT1 (N24367, N24361);
buf BUF1 (N24368, N24358);
or OR3 (N24369, N24364, N4358, N1809);
xor XOR2 (N24370, N24360, N12263);
or OR4 (N24371, N24367, N6184, N583, N16667);
xor XOR2 (N24372, N24371, N17877);
xor XOR2 (N24373, N24366, N12067);
not NOT1 (N24374, N24368);
and AND4 (N24375, N24363, N16834, N16588, N7307);
xor XOR2 (N24376, N24365, N22973);
and AND2 (N24377, N24347, N17511);
or OR4 (N24378, N24373, N12143, N2111, N16669);
nand NAND3 (N24379, N24372, N6882, N14816);
nor NOR2 (N24380, N24376, N10744);
buf BUF1 (N24381, N24378);
and AND3 (N24382, N24381, N761, N8798);
and AND3 (N24383, N24349, N21775, N18839);
nor NOR2 (N24384, N24369, N12653);
xor XOR2 (N24385, N24375, N19929);
xor XOR2 (N24386, N24374, N8805);
or OR3 (N24387, N24386, N4395, N16516);
and AND3 (N24388, N24380, N238, N3878);
xor XOR2 (N24389, N24383, N19504);
or OR4 (N24390, N24389, N13926, N19882, N1023);
or OR4 (N24391, N24382, N9492, N7474, N5870);
nor NOR2 (N24392, N24388, N17554);
xor XOR2 (N24393, N24370, N13158);
xor XOR2 (N24394, N24390, N16735);
and AND2 (N24395, N24394, N7383);
buf BUF1 (N24396, N24392);
buf BUF1 (N24397, N24387);
nor NOR3 (N24398, N24396, N14788, N20575);
nand NAND4 (N24399, N24377, N21219, N21765, N4795);
xor XOR2 (N24400, N24357, N14360);
buf BUF1 (N24401, N24399);
nand NAND4 (N24402, N24401, N14860, N12984, N7619);
nor NOR2 (N24403, N24397, N15411);
and AND3 (N24404, N24398, N5744, N19087);
or OR2 (N24405, N24400, N22089);
and AND4 (N24406, N24403, N22959, N12789, N8335);
not NOT1 (N24407, N24393);
buf BUF1 (N24408, N24391);
nand NAND4 (N24409, N24402, N22954, N15930, N3480);
nand NAND4 (N24410, N24409, N13047, N14378, N10243);
buf BUF1 (N24411, N24385);
buf BUF1 (N24412, N24405);
buf BUF1 (N24413, N24406);
or OR2 (N24414, N24407, N16538);
buf BUF1 (N24415, N24379);
buf BUF1 (N24416, N24414);
buf BUF1 (N24417, N24416);
and AND3 (N24418, N24417, N22498, N21927);
not NOT1 (N24419, N24410);
or OR3 (N24420, N24419, N18101, N20892);
or OR2 (N24421, N24418, N23399);
not NOT1 (N24422, N24408);
buf BUF1 (N24423, N24415);
buf BUF1 (N24424, N24423);
or OR3 (N24425, N24413, N19882, N8585);
nor NOR3 (N24426, N24424, N10001, N5663);
and AND2 (N24427, N24421, N1740);
xor XOR2 (N24428, N24384, N20282);
and AND2 (N24429, N24412, N7260);
or OR3 (N24430, N24426, N18561, N18692);
not NOT1 (N24431, N24428);
xor XOR2 (N24432, N24427, N13752);
buf BUF1 (N24433, N24432);
and AND2 (N24434, N24422, N2177);
not NOT1 (N24435, N24433);
nor NOR2 (N24436, N24430, N809);
or OR4 (N24437, N24434, N23601, N19480, N3407);
or OR3 (N24438, N24411, N12864, N17166);
nand NAND4 (N24439, N24431, N4654, N13568, N17071);
nor NOR4 (N24440, N24425, N16609, N15282, N76);
nand NAND3 (N24441, N24436, N5421, N15111);
and AND3 (N24442, N24437, N5569, N24348);
nor NOR3 (N24443, N24438, N24102, N16215);
nand NAND4 (N24444, N24443, N10453, N12252, N24329);
not NOT1 (N24445, N24440);
nand NAND2 (N24446, N24442, N8762);
buf BUF1 (N24447, N24445);
not NOT1 (N24448, N24447);
nand NAND2 (N24449, N24439, N18574);
not NOT1 (N24450, N24429);
or OR3 (N24451, N24449, N3877, N22856);
nand NAND4 (N24452, N24446, N6830, N19419, N2382);
not NOT1 (N24453, N24441);
or OR3 (N24454, N24404, N5200, N19806);
nor NOR2 (N24455, N24451, N15457);
and AND4 (N24456, N24452, N20879, N10390, N3309);
or OR4 (N24457, N24420, N19854, N10692, N17463);
xor XOR2 (N24458, N24450, N14751);
nor NOR4 (N24459, N24454, N8636, N1783, N20584);
nor NOR4 (N24460, N24444, N19008, N20179, N5733);
nand NAND3 (N24461, N24453, N21573, N12389);
or OR2 (N24462, N24460, N19051);
nor NOR2 (N24463, N24456, N16685);
or OR4 (N24464, N24459, N11825, N22710, N18930);
xor XOR2 (N24465, N24462, N18921);
nand NAND2 (N24466, N24455, N22791);
buf BUF1 (N24467, N24435);
buf BUF1 (N24468, N24466);
or OR4 (N24469, N24467, N20123, N18005, N958);
and AND4 (N24470, N24463, N8444, N16926, N9734);
or OR4 (N24471, N24470, N15564, N16807, N19567);
buf BUF1 (N24472, N24461);
not NOT1 (N24473, N24448);
or OR4 (N24474, N24458, N877, N9201, N6891);
or OR3 (N24475, N24464, N541, N12241);
not NOT1 (N24476, N24457);
nor NOR3 (N24477, N24476, N22628, N23043);
not NOT1 (N24478, N24468);
nor NOR3 (N24479, N24469, N12274, N9102);
not NOT1 (N24480, N24474);
nand NAND3 (N24481, N24477, N13472, N10183);
nor NOR4 (N24482, N24472, N2576, N6541, N12106);
and AND4 (N24483, N24479, N8762, N9622, N22215);
or OR3 (N24484, N24471, N23662, N1079);
not NOT1 (N24485, N24483);
and AND2 (N24486, N24484, N9610);
xor XOR2 (N24487, N24482, N16370);
or OR4 (N24488, N24475, N3386, N9617, N20760);
and AND3 (N24489, N24395, N3054, N17596);
and AND4 (N24490, N24485, N1187, N4368, N17331);
nand NAND2 (N24491, N24488, N23865);
not NOT1 (N24492, N24486);
buf BUF1 (N24493, N24481);
and AND4 (N24494, N24490, N13079, N15856, N19684);
xor XOR2 (N24495, N24494, N10213);
nor NOR4 (N24496, N24465, N18407, N23692, N2454);
xor XOR2 (N24497, N24473, N22898);
not NOT1 (N24498, N24497);
nand NAND4 (N24499, N24495, N9531, N10296, N3787);
buf BUF1 (N24500, N24480);
not NOT1 (N24501, N24491);
buf BUF1 (N24502, N24496);
buf BUF1 (N24503, N24492);
xor XOR2 (N24504, N24501, N3497);
buf BUF1 (N24505, N24502);
or OR4 (N24506, N24505, N5152, N21750, N2447);
buf BUF1 (N24507, N24504);
buf BUF1 (N24508, N24500);
xor XOR2 (N24509, N24508, N13423);
nand NAND4 (N24510, N24509, N4234, N14809, N704);
xor XOR2 (N24511, N24478, N14704);
not NOT1 (N24512, N24489);
and AND4 (N24513, N24487, N23551, N3277, N21873);
not NOT1 (N24514, N24513);
nand NAND3 (N24515, N24503, N14888, N11287);
not NOT1 (N24516, N24499);
and AND2 (N24517, N24514, N2412);
buf BUF1 (N24518, N24516);
nor NOR4 (N24519, N24507, N20819, N9434, N10259);
xor XOR2 (N24520, N24512, N20280);
xor XOR2 (N24521, N24510, N19315);
not NOT1 (N24522, N24493);
xor XOR2 (N24523, N24518, N20120);
nor NOR4 (N24524, N24520, N5020, N1833, N1678);
nor NOR2 (N24525, N24521, N3620);
not NOT1 (N24526, N24511);
nand NAND4 (N24527, N24526, N7571, N23276, N21209);
xor XOR2 (N24528, N24517, N19883);
and AND4 (N24529, N24527, N20074, N20689, N3552);
not NOT1 (N24530, N24498);
and AND2 (N24531, N24523, N3531);
buf BUF1 (N24532, N24531);
nor NOR3 (N24533, N24532, N7856, N3014);
nor NOR3 (N24534, N24515, N21914, N19731);
xor XOR2 (N24535, N24528, N9285);
buf BUF1 (N24536, N24506);
xor XOR2 (N24537, N24536, N23661);
nand NAND3 (N24538, N24525, N6056, N18574);
buf BUF1 (N24539, N24538);
or OR2 (N24540, N24530, N7832);
xor XOR2 (N24541, N24534, N5025);
or OR2 (N24542, N24541, N15174);
nand NAND4 (N24543, N24524, N5218, N11785, N4793);
xor XOR2 (N24544, N24543, N8749);
xor XOR2 (N24545, N24537, N2283);
xor XOR2 (N24546, N24529, N18773);
nand NAND2 (N24547, N24542, N6392);
xor XOR2 (N24548, N24533, N11215);
and AND3 (N24549, N24522, N1522, N13135);
or OR4 (N24550, N24535, N14233, N1869, N2639);
buf BUF1 (N24551, N24546);
buf BUF1 (N24552, N24549);
nor NOR2 (N24553, N24544, N22022);
or OR2 (N24554, N24545, N13474);
xor XOR2 (N24555, N24539, N1295);
nand NAND4 (N24556, N24553, N7872, N21732, N16405);
buf BUF1 (N24557, N24551);
nand NAND4 (N24558, N24552, N1068, N10907, N14168);
nand NAND4 (N24559, N24519, N20538, N10651, N19867);
not NOT1 (N24560, N24554);
nand NAND4 (N24561, N24558, N19672, N22823, N18638);
and AND2 (N24562, N24548, N21462);
not NOT1 (N24563, N24559);
and AND2 (N24564, N24550, N21311);
xor XOR2 (N24565, N24547, N22064);
xor XOR2 (N24566, N24557, N14309);
buf BUF1 (N24567, N24565);
buf BUF1 (N24568, N24562);
not NOT1 (N24569, N24561);
xor XOR2 (N24570, N24563, N14521);
nand NAND4 (N24571, N24569, N16789, N15876, N13436);
xor XOR2 (N24572, N24568, N17174);
and AND3 (N24573, N24556, N8592, N9083);
buf BUF1 (N24574, N24566);
nor NOR4 (N24575, N24570, N11846, N15691, N464);
nor NOR2 (N24576, N24555, N15931);
xor XOR2 (N24577, N24573, N10147);
nor NOR3 (N24578, N24572, N7907, N16901);
or OR4 (N24579, N24576, N9193, N11340, N12923);
or OR4 (N24580, N24571, N22271, N11627, N15499);
not NOT1 (N24581, N24579);
nand NAND2 (N24582, N24580, N14783);
buf BUF1 (N24583, N24578);
xor XOR2 (N24584, N24564, N11733);
xor XOR2 (N24585, N24575, N16072);
buf BUF1 (N24586, N24585);
or OR3 (N24587, N24582, N10968, N10537);
and AND4 (N24588, N24560, N4895, N5330, N9876);
and AND2 (N24589, N24588, N12066);
buf BUF1 (N24590, N24586);
xor XOR2 (N24591, N24574, N9885);
buf BUF1 (N24592, N24591);
and AND3 (N24593, N24567, N11317, N10302);
not NOT1 (N24594, N24584);
nand NAND4 (N24595, N24587, N251, N378, N20230);
and AND4 (N24596, N24592, N15951, N6067, N17204);
xor XOR2 (N24597, N24590, N22076);
nand NAND3 (N24598, N24595, N22585, N309);
nand NAND3 (N24599, N24589, N23154, N12597);
nor NOR3 (N24600, N24593, N5176, N7024);
nor NOR2 (N24601, N24600, N5087);
nand NAND3 (N24602, N24577, N17878, N23072);
nor NOR3 (N24603, N24594, N21493, N9772);
nor NOR3 (N24604, N24602, N20986, N22115);
xor XOR2 (N24605, N24598, N9479);
nand NAND2 (N24606, N24597, N2913);
xor XOR2 (N24607, N24599, N6010);
or OR3 (N24608, N24607, N19271, N18856);
and AND2 (N24609, N24540, N19243);
not NOT1 (N24610, N24596);
xor XOR2 (N24611, N24581, N16118);
and AND2 (N24612, N24609, N7685);
and AND3 (N24613, N24605, N3255, N4271);
nand NAND3 (N24614, N24603, N20551, N23184);
nor NOR2 (N24615, N24614, N3237);
or OR2 (N24616, N24615, N11946);
not NOT1 (N24617, N24604);
buf BUF1 (N24618, N24606);
or OR3 (N24619, N24618, N19471, N7961);
nand NAND4 (N24620, N24611, N2689, N17612, N24012);
nor NOR4 (N24621, N24620, N10642, N3557, N19697);
buf BUF1 (N24622, N24619);
buf BUF1 (N24623, N24612);
and AND3 (N24624, N24622, N20404, N13212);
not NOT1 (N24625, N24617);
nor NOR3 (N24626, N24583, N22494, N10398);
nor NOR2 (N24627, N24616, N9358);
buf BUF1 (N24628, N24626);
nand NAND2 (N24629, N24601, N13881);
nor NOR3 (N24630, N24621, N4081, N18984);
xor XOR2 (N24631, N24624, N15739);
or OR2 (N24632, N24629, N8843);
nor NOR2 (N24633, N24630, N17852);
and AND2 (N24634, N24610, N9645);
nand NAND4 (N24635, N24627, N23847, N23212, N2110);
or OR2 (N24636, N24623, N10968);
not NOT1 (N24637, N24613);
nor NOR2 (N24638, N24608, N16505);
and AND2 (N24639, N24635, N11769);
xor XOR2 (N24640, N24628, N19694);
nand NAND2 (N24641, N24634, N22987);
or OR2 (N24642, N24637, N4941);
nand NAND2 (N24643, N24641, N19003);
or OR3 (N24644, N24639, N8956, N8993);
nand NAND3 (N24645, N24640, N2198, N20709);
or OR3 (N24646, N24625, N19170, N8634);
nand NAND3 (N24647, N24631, N12629, N13040);
xor XOR2 (N24648, N24636, N10455);
nor NOR2 (N24649, N24644, N18490);
and AND4 (N24650, N24638, N1684, N15476, N7206);
buf BUF1 (N24651, N24646);
xor XOR2 (N24652, N24645, N9312);
or OR3 (N24653, N24651, N5679, N22030);
buf BUF1 (N24654, N24652);
and AND3 (N24655, N24648, N14771, N3762);
and AND2 (N24656, N24632, N13966);
nor NOR4 (N24657, N24649, N5888, N13782, N8056);
not NOT1 (N24658, N24642);
xor XOR2 (N24659, N24654, N12630);
buf BUF1 (N24660, N24655);
nor NOR3 (N24661, N24650, N4371, N16654);
nor NOR2 (N24662, N24658, N9315);
or OR2 (N24663, N24633, N8932);
or OR2 (N24664, N24657, N12157);
buf BUF1 (N24665, N24664);
or OR3 (N24666, N24660, N14178, N4368);
xor XOR2 (N24667, N24661, N9093);
nor NOR3 (N24668, N24666, N6623, N22213);
buf BUF1 (N24669, N24643);
or OR4 (N24670, N24665, N23080, N24580, N8746);
nor NOR2 (N24671, N24662, N4114);
not NOT1 (N24672, N24656);
nand NAND4 (N24673, N24663, N10416, N7090, N15169);
or OR3 (N24674, N24672, N5905, N9818);
or OR4 (N24675, N24674, N15588, N10686, N789);
nor NOR2 (N24676, N24659, N21805);
or OR4 (N24677, N24653, N11758, N21391, N20473);
not NOT1 (N24678, N24667);
and AND4 (N24679, N24670, N14036, N15151, N3162);
not NOT1 (N24680, N24677);
xor XOR2 (N24681, N24678, N607);
not NOT1 (N24682, N24680);
not NOT1 (N24683, N24681);
nand NAND2 (N24684, N24671, N15646);
nand NAND2 (N24685, N24676, N21020);
buf BUF1 (N24686, N24669);
nor NOR3 (N24687, N24684, N19805, N18924);
and AND2 (N24688, N24673, N22138);
nand NAND4 (N24689, N24688, N24032, N3744, N24441);
buf BUF1 (N24690, N24675);
xor XOR2 (N24691, N24647, N460);
nand NAND3 (N24692, N24687, N5420, N21647);
not NOT1 (N24693, N24683);
buf BUF1 (N24694, N24668);
and AND4 (N24695, N24694, N5130, N1729, N3942);
nor NOR3 (N24696, N24689, N14185, N6030);
or OR2 (N24697, N24686, N8177);
and AND3 (N24698, N24693, N15111, N2330);
not NOT1 (N24699, N24696);
not NOT1 (N24700, N24679);
buf BUF1 (N24701, N24682);
buf BUF1 (N24702, N24692);
and AND3 (N24703, N24699, N22093, N9341);
xor XOR2 (N24704, N24697, N12889);
nor NOR4 (N24705, N24691, N19589, N6202, N22346);
or OR3 (N24706, N24703, N21908, N1869);
buf BUF1 (N24707, N24695);
or OR3 (N24708, N24700, N13196, N1114);
nand NAND3 (N24709, N24701, N12944, N15994);
and AND3 (N24710, N24702, N24549, N13573);
or OR3 (N24711, N24698, N4707, N11256);
buf BUF1 (N24712, N24710);
xor XOR2 (N24713, N24704, N24019);
xor XOR2 (N24714, N24708, N15686);
xor XOR2 (N24715, N24690, N4208);
nand NAND3 (N24716, N24685, N1324, N3646);
xor XOR2 (N24717, N24713, N17019);
not NOT1 (N24718, N24706);
buf BUF1 (N24719, N24717);
and AND4 (N24720, N24705, N361, N21657, N18008);
and AND3 (N24721, N24715, N15072, N5079);
xor XOR2 (N24722, N24719, N58);
nor NOR4 (N24723, N24712, N23359, N11262, N3682);
nor NOR2 (N24724, N24714, N7923);
or OR4 (N24725, N24722, N20759, N21688, N1727);
xor XOR2 (N24726, N24723, N13127);
nand NAND4 (N24727, N24718, N24306, N18332, N12006);
buf BUF1 (N24728, N24720);
xor XOR2 (N24729, N24707, N6492);
and AND3 (N24730, N24727, N15404, N24586);
or OR4 (N24731, N24725, N9246, N13453, N2583);
nand NAND4 (N24732, N24729, N17892, N14742, N2822);
nand NAND4 (N24733, N24728, N23014, N5828, N12267);
not NOT1 (N24734, N24709);
xor XOR2 (N24735, N24730, N10138);
xor XOR2 (N24736, N24724, N19978);
nand NAND2 (N24737, N24732, N7947);
buf BUF1 (N24738, N24726);
xor XOR2 (N24739, N24737, N1025);
xor XOR2 (N24740, N24711, N19423);
or OR3 (N24741, N24736, N4615, N6495);
nor NOR2 (N24742, N24721, N17187);
not NOT1 (N24743, N24716);
nand NAND4 (N24744, N24734, N885, N4912, N12425);
nor NOR3 (N24745, N24738, N4231, N405);
and AND3 (N24746, N24735, N3639, N15335);
nand NAND2 (N24747, N24745, N14013);
not NOT1 (N24748, N24741);
nor NOR4 (N24749, N24739, N16062, N20840, N6617);
nor NOR2 (N24750, N24746, N18813);
or OR4 (N24751, N24750, N12249, N24267, N9257);
buf BUF1 (N24752, N24744);
or OR2 (N24753, N24731, N22275);
and AND3 (N24754, N24742, N13870, N13175);
not NOT1 (N24755, N24753);
and AND4 (N24756, N24733, N16908, N13579, N301);
not NOT1 (N24757, N24755);
nor NOR4 (N24758, N24747, N12711, N23404, N8672);
nor NOR4 (N24759, N24752, N14782, N17817, N6605);
xor XOR2 (N24760, N24758, N15451);
buf BUF1 (N24761, N24756);
nand NAND2 (N24762, N24743, N17585);
nor NOR3 (N24763, N24759, N12513, N12767);
nand NAND2 (N24764, N24748, N22200);
or OR2 (N24765, N24763, N2292);
or OR2 (N24766, N24754, N3853);
and AND2 (N24767, N24757, N20040);
or OR2 (N24768, N24762, N7187);
and AND2 (N24769, N24760, N6271);
buf BUF1 (N24770, N24767);
buf BUF1 (N24771, N24765);
xor XOR2 (N24772, N24740, N5905);
nor NOR3 (N24773, N24770, N17664, N20623);
and AND3 (N24774, N24751, N4915, N7235);
buf BUF1 (N24775, N24749);
nor NOR4 (N24776, N24769, N20182, N10004, N24498);
nand NAND3 (N24777, N24766, N22400, N13038);
xor XOR2 (N24778, N24761, N7062);
nand NAND4 (N24779, N24777, N4590, N10728, N19532);
xor XOR2 (N24780, N24771, N23655);
xor XOR2 (N24781, N24772, N6700);
and AND2 (N24782, N24768, N6445);
xor XOR2 (N24783, N24778, N17028);
or OR3 (N24784, N24764, N6386, N16281);
and AND4 (N24785, N24781, N9939, N3296, N18700);
buf BUF1 (N24786, N24782);
xor XOR2 (N24787, N24785, N21617);
nand NAND4 (N24788, N24779, N17918, N596, N22645);
xor XOR2 (N24789, N24783, N11630);
xor XOR2 (N24790, N24784, N16238);
buf BUF1 (N24791, N24774);
xor XOR2 (N24792, N24773, N14151);
buf BUF1 (N24793, N24776);
and AND4 (N24794, N24792, N15681, N18643, N9273);
and AND2 (N24795, N24790, N302);
not NOT1 (N24796, N24795);
and AND2 (N24797, N24794, N14910);
xor XOR2 (N24798, N24797, N5429);
or OR4 (N24799, N24787, N10200, N11536, N7626);
or OR2 (N24800, N24791, N6720);
not NOT1 (N24801, N24780);
nor NOR4 (N24802, N24793, N23943, N11594, N15676);
nor NOR3 (N24803, N24798, N20792, N12628);
xor XOR2 (N24804, N24786, N17761);
not NOT1 (N24805, N24799);
and AND2 (N24806, N24802, N12188);
nand NAND3 (N24807, N24801, N10064, N20214);
not NOT1 (N24808, N24804);
nor NOR4 (N24809, N24789, N17759, N11259, N3624);
buf BUF1 (N24810, N24806);
and AND4 (N24811, N24775, N24452, N19695, N5569);
nor NOR3 (N24812, N24805, N9316, N22312);
nand NAND2 (N24813, N24811, N9444);
buf BUF1 (N24814, N24809);
nor NOR4 (N24815, N24807, N18165, N15501, N17691);
nand NAND4 (N24816, N24800, N22612, N15279, N14037);
nand NAND4 (N24817, N24810, N15199, N5328, N4783);
buf BUF1 (N24818, N24814);
xor XOR2 (N24819, N24803, N16733);
and AND2 (N24820, N24796, N18698);
or OR3 (N24821, N24815, N5689, N12524);
and AND4 (N24822, N24808, N4181, N13912, N24600);
buf BUF1 (N24823, N24822);
nand NAND3 (N24824, N24812, N15408, N15962);
or OR3 (N24825, N24820, N12297, N10177);
nor NOR3 (N24826, N24819, N4812, N12826);
nand NAND2 (N24827, N24821, N19433);
nand NAND2 (N24828, N24818, N11075);
or OR4 (N24829, N24788, N4346, N20433, N9782);
not NOT1 (N24830, N24816);
nand NAND3 (N24831, N24829, N17628, N2150);
xor XOR2 (N24832, N24826, N10896);
or OR3 (N24833, N24830, N4841, N19658);
nor NOR4 (N24834, N24833, N6671, N19340, N23535);
or OR4 (N24835, N24823, N10563, N12513, N13430);
buf BUF1 (N24836, N24824);
nor NOR2 (N24837, N24831, N18109);
xor XOR2 (N24838, N24817, N6378);
or OR4 (N24839, N24825, N9187, N10068, N13822);
not NOT1 (N24840, N24834);
or OR3 (N24841, N24839, N7079, N12138);
xor XOR2 (N24842, N24827, N15375);
nand NAND4 (N24843, N24835, N2608, N7755, N5844);
nor NOR3 (N24844, N24841, N10319, N2240);
nand NAND4 (N24845, N24844, N298, N15938, N9954);
nor NOR2 (N24846, N24845, N20250);
xor XOR2 (N24847, N24837, N15372);
or OR4 (N24848, N24813, N8009, N7533, N13224);
nand NAND2 (N24849, N24832, N19982);
and AND3 (N24850, N24840, N9607, N4746);
or OR3 (N24851, N24846, N733, N7743);
not NOT1 (N24852, N24849);
not NOT1 (N24853, N24842);
and AND2 (N24854, N24838, N15140);
buf BUF1 (N24855, N24853);
nor NOR4 (N24856, N24843, N7317, N5782, N17260);
nor NOR4 (N24857, N24836, N5049, N17888, N14555);
nor NOR3 (N24858, N24855, N23035, N21692);
not NOT1 (N24859, N24856);
and AND4 (N24860, N24828, N20606, N14159, N11228);
buf BUF1 (N24861, N24850);
buf BUF1 (N24862, N24851);
not NOT1 (N24863, N24857);
buf BUF1 (N24864, N24861);
xor XOR2 (N24865, N24852, N19682);
nand NAND4 (N24866, N24859, N13646, N23591, N18504);
buf BUF1 (N24867, N24854);
or OR3 (N24868, N24866, N3903, N22182);
xor XOR2 (N24869, N24848, N16221);
and AND4 (N24870, N24860, N5607, N5201, N15708);
nor NOR4 (N24871, N24847, N1995, N22891, N8680);
xor XOR2 (N24872, N24868, N5041);
buf BUF1 (N24873, N24858);
nand NAND3 (N24874, N24873, N20869, N9047);
nand NAND2 (N24875, N24862, N9195);
and AND3 (N24876, N24869, N2637, N19219);
nand NAND4 (N24877, N24871, N3749, N9213, N5010);
not NOT1 (N24878, N24874);
xor XOR2 (N24879, N24878, N12168);
not NOT1 (N24880, N24876);
or OR3 (N24881, N24863, N12819, N6250);
and AND3 (N24882, N24879, N19005, N1801);
xor XOR2 (N24883, N24880, N8798);
and AND2 (N24884, N24881, N9862);
or OR3 (N24885, N24872, N1049, N18164);
and AND4 (N24886, N24865, N2494, N81, N16796);
buf BUF1 (N24887, N24877);
or OR2 (N24888, N24864, N1312);
nand NAND4 (N24889, N24883, N18057, N20866, N20276);
nand NAND4 (N24890, N24885, N20965, N7453, N6147);
and AND2 (N24891, N24870, N11758);
nor NOR3 (N24892, N24888, N9160, N19733);
nor NOR3 (N24893, N24886, N7934, N13484);
nand NAND3 (N24894, N24887, N3654, N10407);
nor NOR2 (N24895, N24893, N19284);
not NOT1 (N24896, N24894);
buf BUF1 (N24897, N24882);
and AND2 (N24898, N24890, N20182);
buf BUF1 (N24899, N24895);
or OR3 (N24900, N24867, N16959, N16945);
or OR3 (N24901, N24897, N16878, N6740);
buf BUF1 (N24902, N24898);
buf BUF1 (N24903, N24884);
not NOT1 (N24904, N24875);
nand NAND3 (N24905, N24899, N16206, N6969);
nand NAND2 (N24906, N24889, N6165);
or OR2 (N24907, N24904, N3134);
and AND4 (N24908, N24900, N22232, N17794, N7482);
xor XOR2 (N24909, N24905, N10712);
nand NAND4 (N24910, N24909, N21556, N18134, N13439);
xor XOR2 (N24911, N24896, N14601);
xor XOR2 (N24912, N24906, N21755);
nor NOR4 (N24913, N24912, N5337, N13072, N15361);
nor NOR2 (N24914, N24892, N15150);
buf BUF1 (N24915, N24908);
not NOT1 (N24916, N24913);
and AND3 (N24917, N24891, N561, N26);
and AND4 (N24918, N24907, N17236, N10754, N17338);
nand NAND2 (N24919, N24915, N4244);
or OR3 (N24920, N24903, N3196, N18887);
nor NOR2 (N24921, N24910, N2564);
xor XOR2 (N24922, N24919, N20103);
or OR4 (N24923, N24902, N9680, N12815, N17409);
buf BUF1 (N24924, N24901);
buf BUF1 (N24925, N24921);
and AND4 (N24926, N24920, N19810, N10275, N2208);
not NOT1 (N24927, N24917);
nand NAND2 (N24928, N24914, N2718);
not NOT1 (N24929, N24924);
or OR3 (N24930, N24928, N7860, N22346);
xor XOR2 (N24931, N24927, N1376);
nand NAND2 (N24932, N24922, N19542);
or OR3 (N24933, N24911, N11313, N6401);
buf BUF1 (N24934, N24931);
or OR3 (N24935, N24929, N6180, N1203);
or OR4 (N24936, N24918, N21949, N719, N10366);
xor XOR2 (N24937, N24936, N10668);
nand NAND4 (N24938, N24933, N15745, N20956, N1299);
nor NOR3 (N24939, N24934, N9867, N17743);
buf BUF1 (N24940, N24938);
nand NAND4 (N24941, N24925, N14988, N682, N2795);
buf BUF1 (N24942, N24926);
nand NAND3 (N24943, N24937, N24848, N14139);
nor NOR4 (N24944, N24940, N22389, N15472, N24044);
and AND3 (N24945, N24930, N1291, N21900);
not NOT1 (N24946, N24943);
or OR2 (N24947, N24944, N6960);
xor XOR2 (N24948, N24935, N17522);
or OR2 (N24949, N24932, N7612);
not NOT1 (N24950, N24945);
not NOT1 (N24951, N24923);
not NOT1 (N24952, N24946);
xor XOR2 (N24953, N24948, N13715);
or OR4 (N24954, N24953, N14652, N5269, N22689);
or OR3 (N24955, N24939, N18503, N9069);
nor NOR2 (N24956, N24952, N5947);
nor NOR2 (N24957, N24947, N7588);
and AND4 (N24958, N24950, N19673, N523, N6417);
and AND4 (N24959, N24955, N1000, N14561, N22648);
not NOT1 (N24960, N24958);
not NOT1 (N24961, N24949);
or OR4 (N24962, N24959, N23672, N1575, N21841);
xor XOR2 (N24963, N24956, N2160);
or OR4 (N24964, N24942, N6434, N19314, N21658);
or OR2 (N24965, N24964, N6097);
not NOT1 (N24966, N24960);
or OR2 (N24967, N24961, N65);
or OR4 (N24968, N24967, N11190, N20854, N15962);
or OR3 (N24969, N24957, N1737, N14537);
xor XOR2 (N24970, N24966, N19777);
not NOT1 (N24971, N24954);
xor XOR2 (N24972, N24963, N8713);
not NOT1 (N24973, N24970);
not NOT1 (N24974, N24972);
and AND4 (N24975, N24973, N3886, N9507, N2672);
not NOT1 (N24976, N24974);
nand NAND3 (N24977, N24969, N6185, N19421);
not NOT1 (N24978, N24962);
not NOT1 (N24979, N24951);
or OR3 (N24980, N24941, N5639, N6870);
and AND3 (N24981, N24971, N15929, N6914);
or OR4 (N24982, N24975, N14572, N333, N14372);
nor NOR2 (N24983, N24979, N20373);
nand NAND4 (N24984, N24976, N16296, N5928, N10365);
nor NOR4 (N24985, N24978, N18067, N2060, N8132);
nor NOR3 (N24986, N24982, N23111, N24029);
buf BUF1 (N24987, N24916);
and AND4 (N24988, N24986, N17319, N18881, N12532);
buf BUF1 (N24989, N24980);
and AND3 (N24990, N24968, N5085, N10232);
nor NOR3 (N24991, N24988, N9869, N23356);
and AND2 (N24992, N24965, N491);
xor XOR2 (N24993, N24987, N5017);
and AND3 (N24994, N24993, N22547, N2228);
or OR3 (N24995, N24981, N2328, N15646);
nand NAND4 (N24996, N24995, N7472, N21716, N9315);
not NOT1 (N24997, N24990);
buf BUF1 (N24998, N24989);
xor XOR2 (N24999, N24991, N6251);
buf BUF1 (N25000, N24998);
or OR4 (N25001, N24984, N13298, N10094, N17259);
buf BUF1 (N25002, N24977);
buf BUF1 (N25003, N24997);
nand NAND4 (N25004, N25000, N18980, N9076, N17478);
nor NOR3 (N25005, N25002, N7300, N18127);
xor XOR2 (N25006, N24985, N8967);
or OR3 (N25007, N25003, N24544, N21185);
or OR2 (N25008, N24992, N11638);
and AND2 (N25009, N25001, N13903);
or OR3 (N25010, N24996, N5640, N5612);
xor XOR2 (N25011, N25006, N12819);
or OR3 (N25012, N25005, N13189, N6353);
and AND2 (N25013, N25011, N19368);
or OR2 (N25014, N25013, N22592);
xor XOR2 (N25015, N25014, N4864);
nor NOR4 (N25016, N25015, N22702, N13993, N3923);
and AND2 (N25017, N25007, N16442);
not NOT1 (N25018, N25016);
nor NOR2 (N25019, N24999, N20844);
nand NAND3 (N25020, N25009, N8388, N13456);
not NOT1 (N25021, N25017);
nand NAND2 (N25022, N25019, N8093);
xor XOR2 (N25023, N24994, N851);
and AND3 (N25024, N25023, N22768, N17315);
nand NAND3 (N25025, N25018, N14345, N2042);
nor NOR3 (N25026, N25025, N8216, N20067);
not NOT1 (N25027, N25021);
buf BUF1 (N25028, N25026);
buf BUF1 (N25029, N25024);
nor NOR2 (N25030, N25010, N24213);
nand NAND2 (N25031, N25008, N23933);
nor NOR2 (N25032, N25030, N4895);
not NOT1 (N25033, N25027);
not NOT1 (N25034, N25033);
nor NOR3 (N25035, N25004, N14841, N20649);
buf BUF1 (N25036, N25012);
and AND3 (N25037, N25020, N19701, N3339);
nor NOR4 (N25038, N25037, N6818, N12064, N11996);
or OR4 (N25039, N25035, N6226, N5002, N7042);
nand NAND4 (N25040, N25039, N21388, N21024, N15459);
buf BUF1 (N25041, N25032);
nor NOR4 (N25042, N25040, N19139, N6591, N24825);
nand NAND4 (N25043, N25042, N23838, N23118, N24393);
not NOT1 (N25044, N25041);
and AND4 (N25045, N25034, N699, N23737, N3309);
buf BUF1 (N25046, N25036);
nand NAND2 (N25047, N24983, N11020);
buf BUF1 (N25048, N25043);
or OR2 (N25049, N25044, N18618);
xor XOR2 (N25050, N25045, N18086);
xor XOR2 (N25051, N25047, N16797);
xor XOR2 (N25052, N25029, N1447);
and AND2 (N25053, N25046, N8027);
or OR2 (N25054, N25052, N6972);
and AND2 (N25055, N25054, N5831);
and AND3 (N25056, N25053, N8499, N7262);
nand NAND4 (N25057, N25050, N20373, N22572, N7804);
and AND2 (N25058, N25028, N3074);
not NOT1 (N25059, N25051);
xor XOR2 (N25060, N25048, N20759);
nor NOR2 (N25061, N25060, N4146);
buf BUF1 (N25062, N25057);
nand NAND3 (N25063, N25038, N9955, N14988);
or OR3 (N25064, N25059, N16621, N6678);
nand NAND3 (N25065, N25022, N991, N19782);
nand NAND4 (N25066, N25063, N2503, N8036, N738);
not NOT1 (N25067, N25049);
nand NAND4 (N25068, N25065, N17465, N13755, N16539);
nand NAND3 (N25069, N25066, N7339, N502);
or OR3 (N25070, N25067, N13090, N23387);
or OR2 (N25071, N25069, N1850);
or OR4 (N25072, N25055, N6289, N4502, N7339);
xor XOR2 (N25073, N25071, N5293);
nand NAND2 (N25074, N25073, N19427);
nand NAND3 (N25075, N25061, N24566, N13598);
or OR2 (N25076, N25068, N2827);
buf BUF1 (N25077, N25031);
and AND2 (N25078, N25056, N21981);
nand NAND2 (N25079, N25075, N14439);
or OR4 (N25080, N25062, N17711, N21685, N20447);
and AND4 (N25081, N25079, N2483, N24970, N12275);
not NOT1 (N25082, N25070);
nor NOR3 (N25083, N25082, N6148, N15526);
and AND2 (N25084, N25058, N20549);
or OR4 (N25085, N25077, N13763, N23113, N21878);
or OR4 (N25086, N25084, N6348, N20437, N23823);
nand NAND3 (N25087, N25074, N22225, N10826);
or OR4 (N25088, N25078, N12808, N24481, N6357);
xor XOR2 (N25089, N25080, N14045);
xor XOR2 (N25090, N25081, N13239);
xor XOR2 (N25091, N25083, N3633);
or OR4 (N25092, N25086, N9051, N3268, N11779);
nand NAND3 (N25093, N25087, N14658, N21469);
and AND2 (N25094, N25076, N21071);
or OR3 (N25095, N25072, N3521, N19064);
not NOT1 (N25096, N25093);
xor XOR2 (N25097, N25094, N16082);
nor NOR3 (N25098, N25090, N3653, N292);
or OR3 (N25099, N25064, N17141, N3391);
nor NOR3 (N25100, N25091, N8884, N9724);
buf BUF1 (N25101, N25097);
xor XOR2 (N25102, N25101, N16829);
nand NAND3 (N25103, N25100, N17539, N10403);
not NOT1 (N25104, N25089);
nand NAND4 (N25105, N25095, N13333, N23786, N8858);
nand NAND4 (N25106, N25098, N13211, N24798, N22549);
xor XOR2 (N25107, N25092, N9949);
nor NOR2 (N25108, N25088, N10495);
nor NOR3 (N25109, N25085, N3851, N8924);
nor NOR2 (N25110, N25108, N3374);
not NOT1 (N25111, N25103);
or OR4 (N25112, N25110, N11606, N18589, N14927);
xor XOR2 (N25113, N25104, N371);
nor NOR2 (N25114, N25105, N15030);
and AND2 (N25115, N25113, N21457);
nor NOR2 (N25116, N25109, N22167);
or OR3 (N25117, N25114, N5580, N19620);
or OR3 (N25118, N25116, N7584, N15019);
xor XOR2 (N25119, N25112, N16977);
nor NOR2 (N25120, N25102, N7092);
nand NAND4 (N25121, N25096, N10156, N19623, N4219);
nor NOR4 (N25122, N25111, N8456, N10809, N18404);
nor NOR3 (N25123, N25117, N20033, N8747);
xor XOR2 (N25124, N25123, N12441);
nor NOR4 (N25125, N25121, N20699, N388, N23824);
or OR4 (N25126, N25125, N14926, N3172, N16011);
nand NAND3 (N25127, N25118, N12954, N17152);
buf BUF1 (N25128, N25107);
xor XOR2 (N25129, N25124, N10900);
or OR3 (N25130, N25127, N7751, N11823);
buf BUF1 (N25131, N25129);
nor NOR3 (N25132, N25131, N1256, N24035);
nor NOR4 (N25133, N25128, N4340, N11812, N6170);
xor XOR2 (N25134, N25106, N5760);
nor NOR2 (N25135, N25119, N22981);
xor XOR2 (N25136, N25134, N5152);
or OR3 (N25137, N25126, N22120, N17380);
nand NAND4 (N25138, N25130, N16934, N8133, N10011);
nand NAND4 (N25139, N25132, N3717, N17340, N15902);
nor NOR3 (N25140, N25135, N3617, N5882);
or OR4 (N25141, N25115, N14875, N3979, N15596);
not NOT1 (N25142, N25136);
nor NOR4 (N25143, N25141, N7561, N20657, N23723);
xor XOR2 (N25144, N25143, N13733);
or OR2 (N25145, N25133, N25031);
nor NOR2 (N25146, N25122, N10790);
buf BUF1 (N25147, N25139);
not NOT1 (N25148, N25142);
and AND4 (N25149, N25138, N15163, N2421, N17392);
nor NOR4 (N25150, N25147, N10961, N2839, N9795);
not NOT1 (N25151, N25148);
nand NAND2 (N25152, N25120, N8047);
nor NOR4 (N25153, N25152, N433, N448, N20653);
not NOT1 (N25154, N25149);
or OR2 (N25155, N25151, N22376);
nor NOR3 (N25156, N25150, N19361, N2218);
nand NAND3 (N25157, N25146, N17783, N24299);
not NOT1 (N25158, N25154);
or OR2 (N25159, N25158, N25060);
not NOT1 (N25160, N25145);
not NOT1 (N25161, N25099);
xor XOR2 (N25162, N25156, N5913);
xor XOR2 (N25163, N25140, N126);
not NOT1 (N25164, N25161);
buf BUF1 (N25165, N25153);
nor NOR4 (N25166, N25157, N20600, N13244, N8485);
not NOT1 (N25167, N25144);
or OR4 (N25168, N25167, N17825, N21691, N1370);
nor NOR3 (N25169, N25168, N20164, N18026);
or OR4 (N25170, N25137, N20711, N23387, N20240);
not NOT1 (N25171, N25162);
nor NOR2 (N25172, N25171, N11713);
and AND4 (N25173, N25164, N19373, N14966, N17079);
or OR4 (N25174, N25159, N2541, N4575, N23830);
xor XOR2 (N25175, N25170, N12415);
not NOT1 (N25176, N25165);
not NOT1 (N25177, N25166);
nor NOR4 (N25178, N25176, N15208, N14906, N11848);
or OR4 (N25179, N25155, N1805, N3628, N6936);
or OR3 (N25180, N25173, N22419, N3048);
xor XOR2 (N25181, N25178, N11403);
and AND2 (N25182, N25169, N14938);
buf BUF1 (N25183, N25179);
and AND3 (N25184, N25160, N20649, N21818);
not NOT1 (N25185, N25175);
nor NOR4 (N25186, N25163, N2868, N19040, N8760);
nand NAND2 (N25187, N25177, N13139);
nor NOR3 (N25188, N25181, N6922, N16713);
nor NOR3 (N25189, N25184, N11060, N9015);
nand NAND4 (N25190, N25187, N9151, N549, N10516);
buf BUF1 (N25191, N25190);
nand NAND3 (N25192, N25186, N9065, N9980);
nand NAND4 (N25193, N25172, N13751, N9257, N4177);
nand NAND4 (N25194, N25174, N23744, N10596, N15887);
not NOT1 (N25195, N25185);
nor NOR2 (N25196, N25193, N23061);
or OR3 (N25197, N25180, N2424, N23919);
nand NAND2 (N25198, N25191, N11037);
xor XOR2 (N25199, N25197, N23731);
nor NOR4 (N25200, N25188, N8628, N5058, N24061);
or OR3 (N25201, N25198, N2705, N18784);
xor XOR2 (N25202, N25196, N23359);
nand NAND3 (N25203, N25200, N5258, N7884);
or OR4 (N25204, N25189, N20920, N25076, N8876);
not NOT1 (N25205, N25192);
xor XOR2 (N25206, N25205, N10027);
and AND2 (N25207, N25195, N19001);
xor XOR2 (N25208, N25194, N3144);
not NOT1 (N25209, N25203);
and AND4 (N25210, N25199, N5430, N20886, N9754);
not NOT1 (N25211, N25202);
buf BUF1 (N25212, N25206);
and AND3 (N25213, N25208, N19722, N14143);
nand NAND4 (N25214, N25209, N24365, N13550, N14473);
and AND3 (N25215, N25204, N23025, N13233);
nor NOR2 (N25216, N25211, N3375);
nor NOR4 (N25217, N25207, N13318, N2204, N13531);
nand NAND4 (N25218, N25215, N7407, N17027, N669);
buf BUF1 (N25219, N25183);
and AND2 (N25220, N25216, N1598);
or OR4 (N25221, N25218, N13130, N23279, N6048);
xor XOR2 (N25222, N25221, N789);
not NOT1 (N25223, N25182);
not NOT1 (N25224, N25213);
and AND2 (N25225, N25214, N24571);
not NOT1 (N25226, N25212);
xor XOR2 (N25227, N25210, N13674);
nand NAND3 (N25228, N25225, N23312, N24884);
not NOT1 (N25229, N25201);
buf BUF1 (N25230, N25227);
nor NOR2 (N25231, N25217, N4124);
xor XOR2 (N25232, N25223, N18077);
nor NOR3 (N25233, N25226, N9833, N4786);
or OR3 (N25234, N25222, N24593, N2970);
nor NOR2 (N25235, N25233, N7554);
not NOT1 (N25236, N25231);
buf BUF1 (N25237, N25230);
and AND4 (N25238, N25228, N16036, N21658, N11554);
nor NOR4 (N25239, N25238, N954, N19925, N14388);
or OR2 (N25240, N25224, N10186);
buf BUF1 (N25241, N25235);
not NOT1 (N25242, N25232);
nor NOR3 (N25243, N25219, N4990, N19961);
nor NOR3 (N25244, N25243, N16643, N21702);
xor XOR2 (N25245, N25241, N23656);
buf BUF1 (N25246, N25236);
not NOT1 (N25247, N25234);
nor NOR4 (N25248, N25242, N2088, N590, N14853);
not NOT1 (N25249, N25220);
or OR2 (N25250, N25248, N2196);
not NOT1 (N25251, N25244);
nand NAND2 (N25252, N25247, N22999);
buf BUF1 (N25253, N25246);
not NOT1 (N25254, N25245);
nor NOR3 (N25255, N25250, N2770, N9708);
buf BUF1 (N25256, N25253);
or OR4 (N25257, N25239, N1966, N6281, N19689);
xor XOR2 (N25258, N25240, N4363);
nand NAND2 (N25259, N25258, N10840);
not NOT1 (N25260, N25257);
nand NAND3 (N25261, N25251, N18337, N2227);
not NOT1 (N25262, N25259);
xor XOR2 (N25263, N25254, N10105);
buf BUF1 (N25264, N25237);
buf BUF1 (N25265, N25262);
not NOT1 (N25266, N25260);
xor XOR2 (N25267, N25264, N8578);
not NOT1 (N25268, N25249);
buf BUF1 (N25269, N25261);
nand NAND2 (N25270, N25267, N14392);
nand NAND4 (N25271, N25252, N18572, N14530, N11139);
xor XOR2 (N25272, N25263, N4271);
and AND4 (N25273, N25271, N13945, N8408, N15133);
buf BUF1 (N25274, N25256);
nor NOR3 (N25275, N25274, N23218, N17622);
and AND3 (N25276, N25272, N9763, N14760);
nand NAND3 (N25277, N25270, N2765, N10599);
and AND3 (N25278, N25277, N8841, N11663);
not NOT1 (N25279, N25268);
nand NAND4 (N25280, N25278, N22593, N1399, N21407);
and AND2 (N25281, N25279, N8653);
buf BUF1 (N25282, N25273);
xor XOR2 (N25283, N25265, N17969);
and AND2 (N25284, N25229, N5732);
nand NAND2 (N25285, N25284, N2442);
nand NAND2 (N25286, N25266, N23458);
buf BUF1 (N25287, N25281);
and AND3 (N25288, N25275, N10264, N17139);
nor NOR3 (N25289, N25276, N12404, N17763);
and AND3 (N25290, N25269, N18568, N21972);
buf BUF1 (N25291, N25287);
xor XOR2 (N25292, N25283, N1801);
or OR2 (N25293, N25292, N13212);
or OR4 (N25294, N25288, N23361, N14396, N2063);
xor XOR2 (N25295, N25290, N8372);
and AND2 (N25296, N25255, N6522);
buf BUF1 (N25297, N25291);
nor NOR3 (N25298, N25295, N1803, N4563);
xor XOR2 (N25299, N25298, N22520);
not NOT1 (N25300, N25285);
or OR2 (N25301, N25280, N8348);
buf BUF1 (N25302, N25286);
and AND2 (N25303, N25282, N3696);
buf BUF1 (N25304, N25302);
buf BUF1 (N25305, N25301);
nand NAND4 (N25306, N25296, N10528, N24968, N16441);
nand NAND2 (N25307, N25289, N459);
nor NOR4 (N25308, N25307, N16944, N16629, N6465);
nor NOR4 (N25309, N25293, N15354, N15390, N22953);
not NOT1 (N25310, N25294);
or OR3 (N25311, N25309, N1490, N16051);
buf BUF1 (N25312, N25304);
and AND4 (N25313, N25303, N1020, N8087, N13282);
nor NOR3 (N25314, N25305, N11097, N22639);
nor NOR3 (N25315, N25299, N11980, N13621);
buf BUF1 (N25316, N25308);
or OR4 (N25317, N25312, N21544, N893, N23905);
nor NOR2 (N25318, N25306, N2644);
buf BUF1 (N25319, N25310);
nand NAND2 (N25320, N25300, N16641);
and AND4 (N25321, N25319, N21053, N7878, N22623);
nor NOR4 (N25322, N25313, N845, N17415, N14860);
and AND2 (N25323, N25316, N12002);
or OR3 (N25324, N25297, N14533, N9699);
not NOT1 (N25325, N25314);
buf BUF1 (N25326, N25317);
and AND4 (N25327, N25322, N6592, N18385, N10293);
xor XOR2 (N25328, N25321, N10253);
not NOT1 (N25329, N25325);
or OR2 (N25330, N25324, N14847);
nor NOR3 (N25331, N25311, N5015, N14552);
nor NOR4 (N25332, N25318, N1120, N16495, N22458);
nand NAND2 (N25333, N25328, N10718);
nor NOR3 (N25334, N25333, N15286, N13666);
nor NOR4 (N25335, N25320, N12733, N13001, N8928);
not NOT1 (N25336, N25330);
and AND2 (N25337, N25323, N9999);
xor XOR2 (N25338, N25329, N20346);
xor XOR2 (N25339, N25334, N12542);
nor NOR4 (N25340, N25336, N14723, N17581, N22015);
not NOT1 (N25341, N25339);
not NOT1 (N25342, N25337);
and AND3 (N25343, N25326, N19466, N3135);
and AND3 (N25344, N25327, N11939, N4200);
nand NAND3 (N25345, N25335, N11607, N16704);
or OR4 (N25346, N25315, N4880, N9080, N9122);
and AND3 (N25347, N25331, N8496, N11601);
nand NAND4 (N25348, N25341, N7704, N6830, N18110);
and AND3 (N25349, N25344, N13897, N1179);
nand NAND3 (N25350, N25349, N7143, N19160);
or OR4 (N25351, N25348, N11506, N11500, N18222);
not NOT1 (N25352, N25343);
and AND2 (N25353, N25332, N20596);
not NOT1 (N25354, N25345);
and AND4 (N25355, N25346, N23109, N2437, N23343);
nor NOR3 (N25356, N25353, N12389, N10666);
buf BUF1 (N25357, N25340);
nand NAND4 (N25358, N25347, N6804, N6737, N2653);
nor NOR2 (N25359, N25342, N20774);
and AND4 (N25360, N25354, N14449, N3282, N2812);
not NOT1 (N25361, N25338);
or OR2 (N25362, N25361, N23802);
nand NAND3 (N25363, N25359, N11062, N1030);
buf BUF1 (N25364, N25350);
not NOT1 (N25365, N25351);
not NOT1 (N25366, N25364);
nor NOR4 (N25367, N25362, N11553, N12746, N17376);
buf BUF1 (N25368, N25360);
or OR2 (N25369, N25365, N782);
buf BUF1 (N25370, N25356);
and AND4 (N25371, N25368, N10788, N11194, N15223);
nand NAND4 (N25372, N25370, N15350, N18685, N14882);
nand NAND3 (N25373, N25363, N13045, N2803);
xor XOR2 (N25374, N25372, N10386);
or OR3 (N25375, N25374, N240, N12367);
buf BUF1 (N25376, N25371);
nand NAND3 (N25377, N25369, N15813, N22799);
nor NOR4 (N25378, N25355, N5882, N10454, N18192);
not NOT1 (N25379, N25357);
or OR3 (N25380, N25379, N835, N14358);
nand NAND4 (N25381, N25358, N7607, N23685, N24673);
nor NOR2 (N25382, N25380, N3850);
and AND3 (N25383, N25378, N20922, N14472);
or OR3 (N25384, N25373, N7325, N14184);
nor NOR4 (N25385, N25367, N20231, N6539, N1774);
nor NOR4 (N25386, N25382, N22985, N22003, N16911);
nor NOR4 (N25387, N25386, N22963, N15961, N21134);
not NOT1 (N25388, N25366);
nand NAND2 (N25389, N25376, N12719);
or OR2 (N25390, N25383, N24895);
and AND2 (N25391, N25377, N3150);
buf BUF1 (N25392, N25388);
and AND3 (N25393, N25390, N11057, N19643);
not NOT1 (N25394, N25393);
or OR4 (N25395, N25375, N24034, N4585, N14569);
not NOT1 (N25396, N25384);
and AND4 (N25397, N25396, N710, N2163, N13121);
xor XOR2 (N25398, N25397, N17891);
nand NAND3 (N25399, N25389, N24651, N15549);
or OR3 (N25400, N25395, N19885, N23314);
buf BUF1 (N25401, N25391);
nand NAND3 (N25402, N25387, N20388, N1588);
nand NAND2 (N25403, N25401, N18376);
and AND2 (N25404, N25352, N24937);
not NOT1 (N25405, N25402);
not NOT1 (N25406, N25381);
nor NOR2 (N25407, N25403, N11802);
nor NOR3 (N25408, N25404, N22798, N4242);
xor XOR2 (N25409, N25392, N486);
nand NAND2 (N25410, N25400, N12154);
buf BUF1 (N25411, N25408);
nor NOR3 (N25412, N25406, N14394, N13507);
nand NAND3 (N25413, N25410, N24062, N1370);
nor NOR3 (N25414, N25399, N10263, N20168);
nand NAND3 (N25415, N25414, N7533, N15400);
buf BUF1 (N25416, N25398);
and AND4 (N25417, N25405, N4903, N18693, N10120);
or OR3 (N25418, N25394, N16753, N20899);
nand NAND4 (N25419, N25407, N17058, N9435, N17261);
nand NAND2 (N25420, N25419, N2924);
not NOT1 (N25421, N25409);
nand NAND2 (N25422, N25412, N12883);
nand NAND4 (N25423, N25421, N3473, N24318, N6547);
xor XOR2 (N25424, N25418, N17067);
and AND2 (N25425, N25420, N681);
buf BUF1 (N25426, N25417);
buf BUF1 (N25427, N25422);
or OR2 (N25428, N25411, N16064);
or OR4 (N25429, N25424, N7843, N22203, N21423);
nand NAND4 (N25430, N25415, N3744, N24157, N18881);
not NOT1 (N25431, N25428);
not NOT1 (N25432, N25431);
and AND2 (N25433, N25427, N1577);
and AND4 (N25434, N25413, N5894, N17643, N20012);
or OR4 (N25435, N25429, N10040, N10702, N7274);
xor XOR2 (N25436, N25385, N15199);
nor NOR4 (N25437, N25423, N17681, N5452, N24232);
or OR3 (N25438, N25433, N5044, N1801);
and AND2 (N25439, N25416, N19405);
nor NOR2 (N25440, N25425, N11203);
nand NAND2 (N25441, N25426, N15578);
or OR2 (N25442, N25432, N6226);
not NOT1 (N25443, N25434);
and AND3 (N25444, N25442, N1381, N6261);
nor NOR3 (N25445, N25435, N4039, N7567);
nor NOR3 (N25446, N25436, N4137, N23210);
buf BUF1 (N25447, N25438);
and AND2 (N25448, N25437, N23709);
not NOT1 (N25449, N25440);
or OR2 (N25450, N25430, N1289);
buf BUF1 (N25451, N25450);
or OR2 (N25452, N25445, N14245);
xor XOR2 (N25453, N25447, N4429);
nand NAND4 (N25454, N25452, N15745, N4721, N20885);
nand NAND2 (N25455, N25439, N22460);
not NOT1 (N25456, N25446);
or OR3 (N25457, N25455, N19844, N4959);
xor XOR2 (N25458, N25441, N12322);
xor XOR2 (N25459, N25451, N15677);
xor XOR2 (N25460, N25443, N20476);
buf BUF1 (N25461, N25454);
buf BUF1 (N25462, N25457);
and AND3 (N25463, N25453, N10748, N22241);
buf BUF1 (N25464, N25461);
nand NAND2 (N25465, N25460, N1598);
or OR4 (N25466, N25463, N3227, N9300, N19980);
nor NOR2 (N25467, N25458, N4430);
and AND2 (N25468, N25449, N19691);
not NOT1 (N25469, N25467);
nand NAND3 (N25470, N25456, N947, N11109);
not NOT1 (N25471, N25448);
nand NAND2 (N25472, N25466, N6987);
and AND3 (N25473, N25459, N15456, N31);
xor XOR2 (N25474, N25444, N24844);
and AND3 (N25475, N25465, N22647, N11900);
xor XOR2 (N25476, N25474, N15383);
buf BUF1 (N25477, N25468);
nand NAND3 (N25478, N25472, N14118, N10262);
buf BUF1 (N25479, N25471);
nor NOR2 (N25480, N25462, N23696);
buf BUF1 (N25481, N25475);
not NOT1 (N25482, N25478);
and AND2 (N25483, N25480, N10145);
buf BUF1 (N25484, N25476);
or OR3 (N25485, N25482, N9560, N20684);
not NOT1 (N25486, N25483);
and AND2 (N25487, N25464, N18025);
nor NOR3 (N25488, N25473, N6605, N11564);
buf BUF1 (N25489, N25487);
xor XOR2 (N25490, N25489, N22709);
nand NAND2 (N25491, N25485, N15241);
or OR3 (N25492, N25484, N7006, N19478);
xor XOR2 (N25493, N25481, N3556);
not NOT1 (N25494, N25479);
buf BUF1 (N25495, N25490);
buf BUF1 (N25496, N25495);
and AND2 (N25497, N25486, N20265);
not NOT1 (N25498, N25469);
nand NAND3 (N25499, N25497, N16169, N15726);
buf BUF1 (N25500, N25470);
and AND3 (N25501, N25499, N18419, N403);
not NOT1 (N25502, N25477);
nand NAND4 (N25503, N25494, N2055, N24219, N11404);
or OR2 (N25504, N25498, N22526);
nand NAND4 (N25505, N25504, N23315, N21804, N21323);
xor XOR2 (N25506, N25503, N10138);
nand NAND3 (N25507, N25491, N21108, N21994);
nand NAND2 (N25508, N25502, N25240);
nor NOR4 (N25509, N25508, N9852, N1532, N6853);
and AND4 (N25510, N25507, N3193, N14442, N21729);
nor NOR3 (N25511, N25505, N7339, N19570);
or OR2 (N25512, N25496, N24991);
and AND3 (N25513, N25500, N7231, N17587);
nand NAND3 (N25514, N25512, N24375, N23578);
xor XOR2 (N25515, N25509, N23689);
not NOT1 (N25516, N25514);
nand NAND4 (N25517, N25511, N8839, N7230, N5110);
or OR3 (N25518, N25506, N10960, N82);
nand NAND2 (N25519, N25493, N8413);
nor NOR2 (N25520, N25517, N16905);
nand NAND4 (N25521, N25518, N22382, N9708, N6550);
or OR2 (N25522, N25513, N21459);
buf BUF1 (N25523, N25519);
xor XOR2 (N25524, N25521, N8000);
and AND4 (N25525, N25488, N9349, N9941, N6996);
or OR4 (N25526, N25501, N24172, N11267, N3353);
nor NOR2 (N25527, N25516, N22605);
or OR3 (N25528, N25520, N18553, N17443);
buf BUF1 (N25529, N25526);
not NOT1 (N25530, N25515);
nand NAND2 (N25531, N25530, N1852);
nand NAND2 (N25532, N25510, N1759);
not NOT1 (N25533, N25531);
nand NAND2 (N25534, N25524, N12303);
nor NOR3 (N25535, N25528, N16090, N7488);
or OR2 (N25536, N25534, N13105);
nand NAND2 (N25537, N25532, N14096);
buf BUF1 (N25538, N25527);
nor NOR2 (N25539, N25492, N12427);
buf BUF1 (N25540, N25536);
nand NAND3 (N25541, N25540, N8638, N13900);
and AND3 (N25542, N25541, N18409, N15774);
nand NAND4 (N25543, N25538, N2768, N20139, N17238);
or OR2 (N25544, N25523, N12959);
and AND4 (N25545, N25544, N9489, N17981, N11747);
nor NOR4 (N25546, N25537, N9823, N4613, N4253);
xor XOR2 (N25547, N25539, N19443);
or OR3 (N25548, N25529, N9967, N23986);
nor NOR2 (N25549, N25535, N15399);
nor NOR3 (N25550, N25543, N25414, N1295);
not NOT1 (N25551, N25522);
not NOT1 (N25552, N25551);
nor NOR2 (N25553, N25552, N12368);
not NOT1 (N25554, N25525);
xor XOR2 (N25555, N25549, N2333);
and AND2 (N25556, N25555, N1796);
nand NAND2 (N25557, N25556, N5471);
xor XOR2 (N25558, N25547, N8113);
not NOT1 (N25559, N25553);
or OR3 (N25560, N25548, N18582, N12693);
nor NOR2 (N25561, N25545, N15756);
nor NOR3 (N25562, N25559, N19664, N20491);
and AND4 (N25563, N25550, N977, N11138, N7615);
and AND4 (N25564, N25560, N10, N4, N18368);
xor XOR2 (N25565, N25546, N6173);
and AND3 (N25566, N25558, N21414, N4445);
not NOT1 (N25567, N25533);
xor XOR2 (N25568, N25565, N12799);
not NOT1 (N25569, N25561);
and AND4 (N25570, N25567, N4364, N1329, N10003);
nor NOR4 (N25571, N25570, N22118, N15231, N18990);
and AND4 (N25572, N25571, N7012, N24711, N5251);
buf BUF1 (N25573, N25568);
not NOT1 (N25574, N25554);
nand NAND3 (N25575, N25542, N24565, N2178);
not NOT1 (N25576, N25563);
nand NAND3 (N25577, N25562, N17277, N8238);
not NOT1 (N25578, N25576);
buf BUF1 (N25579, N25578);
and AND3 (N25580, N25577, N22200, N23349);
nor NOR4 (N25581, N25572, N18742, N25482, N22253);
buf BUF1 (N25582, N25574);
nor NOR4 (N25583, N25581, N10621, N18457, N2105);
and AND3 (N25584, N25564, N24147, N19603);
and AND3 (N25585, N25579, N7172, N21676);
nor NOR2 (N25586, N25557, N19782);
not NOT1 (N25587, N25575);
buf BUF1 (N25588, N25583);
and AND3 (N25589, N25566, N16130, N19599);
nor NOR2 (N25590, N25586, N23085);
buf BUF1 (N25591, N25585);
and AND4 (N25592, N25584, N14166, N21334, N11621);
xor XOR2 (N25593, N25590, N6520);
nand NAND4 (N25594, N25589, N6811, N13061, N14308);
nor NOR4 (N25595, N25580, N16814, N4527, N1377);
nand NAND2 (N25596, N25595, N13672);
nand NAND3 (N25597, N25596, N22435, N18924);
buf BUF1 (N25598, N25573);
not NOT1 (N25599, N25593);
not NOT1 (N25600, N25587);
buf BUF1 (N25601, N25588);
and AND4 (N25602, N25594, N22505, N5034, N1857);
or OR2 (N25603, N25597, N3856);
nor NOR2 (N25604, N25569, N17107);
nor NOR4 (N25605, N25604, N14529, N13460, N20825);
xor XOR2 (N25606, N25602, N23929);
not NOT1 (N25607, N25605);
nor NOR3 (N25608, N25599, N13588, N11861);
xor XOR2 (N25609, N25600, N6584);
nor NOR4 (N25610, N25606, N23402, N16996, N17217);
not NOT1 (N25611, N25592);
nand NAND2 (N25612, N25608, N9265);
buf BUF1 (N25613, N25611);
xor XOR2 (N25614, N25609, N6713);
nand NAND2 (N25615, N25582, N15274);
and AND2 (N25616, N25614, N18913);
and AND2 (N25617, N25615, N1771);
nor NOR2 (N25618, N25603, N14605);
endmodule