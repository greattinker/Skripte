// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14;

output N2513,N2509,N2508,N2512,N2505,N2507,N2504,N2481,N2503,N2514;

nor NOR3 (N15, N12, N5, N3);
nor NOR4 (N16, N1, N2, N5, N5);
nand NAND4 (N17, N14, N11, N10, N7);
nor NOR4 (N18, N10, N1, N4, N4);
or OR2 (N19, N14, N7);
nand NAND2 (N20, N10, N7);
buf BUF1 (N21, N2);
nor NOR3 (N22, N17, N15, N15);
nor NOR3 (N23, N12, N7, N15);
xor XOR2 (N24, N12, N1);
nand NAND4 (N25, N7, N21, N2, N22);
and AND4 (N26, N25, N10, N23, N1);
not NOT1 (N27, N21);
nand NAND3 (N28, N15, N21, N26);
buf BUF1 (N29, N7);
not NOT1 (N30, N26);
not NOT1 (N31, N7);
not NOT1 (N32, N20);
xor XOR2 (N33, N32, N5);
not NOT1 (N34, N16);
nor NOR2 (N35, N34, N11);
buf BUF1 (N36, N35);
nor NOR4 (N37, N19, N6, N34, N1);
xor XOR2 (N38, N37, N27);
nor NOR4 (N39, N4, N28, N29, N27);
or OR4 (N40, N19, N24, N22, N21);
and AND2 (N41, N37, N40);
nand NAND4 (N42, N14, N27, N25, N8);
and AND2 (N43, N6, N7);
buf BUF1 (N44, N42);
buf BUF1 (N45, N43);
nand NAND4 (N46, N41, N17, N32, N21);
nor NOR3 (N47, N30, N35, N4);
or OR2 (N48, N38, N36);
or OR3 (N49, N17, N1, N9);
nand NAND4 (N50, N33, N38, N6, N17);
buf BUF1 (N51, N49);
not NOT1 (N52, N47);
buf BUF1 (N53, N45);
xor XOR2 (N54, N48, N47);
nand NAND4 (N55, N18, N20, N2, N29);
not NOT1 (N56, N50);
nand NAND4 (N57, N52, N30, N22, N7);
nor NOR4 (N58, N56, N57, N12, N51);
or OR3 (N59, N54, N25, N16);
not NOT1 (N60, N18);
not NOT1 (N61, N11);
or OR4 (N62, N58, N18, N7, N61);
buf BUF1 (N63, N12);
and AND2 (N64, N60, N50);
buf BUF1 (N65, N62);
not NOT1 (N66, N59);
and AND2 (N67, N44, N2);
buf BUF1 (N68, N39);
xor XOR2 (N69, N68, N45);
not NOT1 (N70, N66);
nor NOR2 (N71, N46, N1);
or OR2 (N72, N64, N47);
nor NOR3 (N73, N31, N63, N2);
xor XOR2 (N74, N5, N69);
not NOT1 (N75, N52);
nand NAND4 (N76, N73, N45, N53, N2);
buf BUF1 (N77, N9);
nand NAND4 (N78, N65, N62, N48, N34);
or OR2 (N79, N77, N28);
buf BUF1 (N80, N76);
or OR2 (N81, N79, N4);
nor NOR3 (N82, N75, N35, N49);
xor XOR2 (N83, N72, N24);
nor NOR3 (N84, N74, N10, N56);
nor NOR3 (N85, N80, N72, N77);
or OR2 (N86, N82, N30);
buf BUF1 (N87, N86);
and AND4 (N88, N81, N67, N54, N14);
buf BUF1 (N89, N76);
and AND3 (N90, N85, N72, N22);
nor NOR4 (N91, N89, N38, N58, N49);
or OR2 (N92, N70, N70);
xor XOR2 (N93, N88, N72);
nand NAND4 (N94, N71, N88, N56, N51);
nor NOR3 (N95, N83, N2, N84);
and AND3 (N96, N73, N27, N17);
buf BUF1 (N97, N95);
nand NAND3 (N98, N97, N18, N95);
nand NAND2 (N99, N93, N40);
or OR4 (N100, N87, N66, N47, N95);
nor NOR4 (N101, N100, N10, N30, N90);
xor XOR2 (N102, N56, N72);
xor XOR2 (N103, N94, N51);
or OR4 (N104, N101, N16, N46, N103);
xor XOR2 (N105, N39, N53);
nand NAND4 (N106, N91, N9, N14, N51);
and AND4 (N107, N102, N39, N104, N86);
xor XOR2 (N108, N9, N50);
or OR4 (N109, N96, N4, N101, N24);
xor XOR2 (N110, N92, N44);
nand NAND4 (N111, N105, N24, N19, N16);
nor NOR2 (N112, N98, N52);
nand NAND3 (N113, N110, N14, N26);
not NOT1 (N114, N107);
buf BUF1 (N115, N55);
xor XOR2 (N116, N108, N104);
buf BUF1 (N117, N109);
xor XOR2 (N118, N114, N2);
nand NAND2 (N119, N115, N13);
xor XOR2 (N120, N119, N105);
nand NAND2 (N121, N120, N7);
and AND3 (N122, N121, N67, N5);
nor NOR3 (N123, N112, N96, N102);
xor XOR2 (N124, N113, N88);
not NOT1 (N125, N111);
not NOT1 (N126, N125);
nor NOR2 (N127, N124, N55);
and AND2 (N128, N127, N83);
not NOT1 (N129, N118);
nor NOR4 (N130, N126, N85, N113, N42);
not NOT1 (N131, N122);
or OR3 (N132, N78, N104, N101);
or OR4 (N133, N131, N33, N52, N9);
nand NAND3 (N134, N117, N30, N22);
not NOT1 (N135, N132);
not NOT1 (N136, N133);
xor XOR2 (N137, N134, N55);
nand NAND4 (N138, N137, N136, N115, N9);
buf BUF1 (N139, N49);
or OR2 (N140, N106, N122);
nor NOR4 (N141, N140, N127, N26, N85);
or OR3 (N142, N139, N128, N31);
buf BUF1 (N143, N135);
nor NOR3 (N144, N9, N21, N21);
and AND4 (N145, N130, N49, N89, N76);
xor XOR2 (N146, N142, N66);
buf BUF1 (N147, N145);
buf BUF1 (N148, N147);
not NOT1 (N149, N123);
xor XOR2 (N150, N138, N100);
xor XOR2 (N151, N144, N150);
nand NAND4 (N152, N89, N90, N17, N113);
not NOT1 (N153, N152);
and AND4 (N154, N146, N132, N17, N105);
xor XOR2 (N155, N151, N75);
xor XOR2 (N156, N148, N106);
xor XOR2 (N157, N155, N29);
nor NOR3 (N158, N116, N130, N28);
and AND3 (N159, N143, N123, N33);
xor XOR2 (N160, N153, N25);
nand NAND3 (N161, N154, N142, N63);
xor XOR2 (N162, N156, N54);
nor NOR2 (N163, N162, N141);
xor XOR2 (N164, N152, N90);
buf BUF1 (N165, N159);
xor XOR2 (N166, N164, N115);
and AND3 (N167, N99, N102, N160);
and AND3 (N168, N5, N154, N89);
buf BUF1 (N169, N129);
or OR3 (N170, N167, N11, N6);
nand NAND3 (N171, N166, N27, N6);
not NOT1 (N172, N149);
nand NAND2 (N173, N169, N72);
or OR4 (N174, N171, N66, N90, N67);
or OR3 (N175, N168, N119, N72);
xor XOR2 (N176, N172, N162);
xor XOR2 (N177, N173, N64);
or OR2 (N178, N161, N1);
and AND2 (N179, N170, N106);
and AND2 (N180, N157, N76);
nor NOR4 (N181, N177, N73, N146, N55);
buf BUF1 (N182, N179);
nand NAND2 (N183, N163, N126);
or OR4 (N184, N174, N181, N68, N4);
or OR3 (N185, N65, N25, N74);
nand NAND2 (N186, N184, N22);
nor NOR4 (N187, N185, N185, N42, N42);
or OR3 (N188, N178, N164, N134);
nor NOR3 (N189, N187, N182, N10);
and AND2 (N190, N117, N88);
buf BUF1 (N191, N190);
nor NOR3 (N192, N183, N22, N94);
nor NOR2 (N193, N186, N33);
nand NAND3 (N194, N193, N156, N129);
or OR3 (N195, N176, N110, N104);
xor XOR2 (N196, N191, N41);
nand NAND3 (N197, N192, N119, N72);
and AND4 (N198, N196, N122, N21, N25);
nor NOR4 (N199, N175, N156, N175, N163);
and AND2 (N200, N194, N86);
nor NOR4 (N201, N165, N108, N195, N46);
not NOT1 (N202, N144);
buf BUF1 (N203, N199);
buf BUF1 (N204, N197);
xor XOR2 (N205, N158, N108);
and AND2 (N206, N200, N173);
buf BUF1 (N207, N202);
nand NAND3 (N208, N207, N149, N123);
nand NAND4 (N209, N205, N145, N131, N139);
and AND4 (N210, N204, N31, N25, N195);
or OR2 (N211, N206, N171);
or OR2 (N212, N208, N128);
or OR4 (N213, N209, N20, N200, N22);
nand NAND3 (N214, N213, N124, N3);
nor NOR2 (N215, N180, N74);
and AND2 (N216, N201, N183);
nand NAND2 (N217, N189, N107);
and AND2 (N218, N212, N200);
or OR2 (N219, N211, N23);
not NOT1 (N220, N198);
nand NAND4 (N221, N203, N106, N159, N160);
nand NAND4 (N222, N221, N120, N64, N153);
or OR4 (N223, N219, N12, N4, N60);
nor NOR2 (N224, N222, N20);
or OR3 (N225, N220, N92, N70);
or OR3 (N226, N188, N214, N111);
xor XOR2 (N227, N202, N4);
not NOT1 (N228, N218);
nor NOR2 (N229, N210, N107);
and AND3 (N230, N227, N62, N147);
nor NOR3 (N231, N225, N167, N32);
not NOT1 (N232, N231);
buf BUF1 (N233, N232);
or OR2 (N234, N229, N53);
and AND4 (N235, N226, N146, N35, N16);
not NOT1 (N236, N235);
not NOT1 (N237, N223);
xor XOR2 (N238, N224, N177);
buf BUF1 (N239, N217);
not NOT1 (N240, N228);
nand NAND3 (N241, N240, N81, N109);
xor XOR2 (N242, N216, N182);
and AND4 (N243, N215, N22, N211, N60);
nor NOR3 (N244, N243, N185, N43);
nand NAND4 (N245, N236, N81, N223, N227);
and AND4 (N246, N233, N118, N77, N96);
or OR4 (N247, N230, N79, N39, N141);
or OR4 (N248, N238, N14, N220, N20);
or OR3 (N249, N244, N136, N5);
buf BUF1 (N250, N241);
nor NOR4 (N251, N242, N175, N36, N220);
nor NOR3 (N252, N237, N103, N119);
not NOT1 (N253, N251);
nand NAND3 (N254, N248, N71, N189);
and AND2 (N255, N239, N232);
not NOT1 (N256, N246);
nor NOR2 (N257, N234, N92);
not NOT1 (N258, N256);
xor XOR2 (N259, N258, N134);
nor NOR2 (N260, N259, N208);
nor NOR3 (N261, N260, N68, N9);
nor NOR3 (N262, N250, N144, N218);
nor NOR2 (N263, N253, N148);
not NOT1 (N264, N255);
nand NAND4 (N265, N254, N111, N218, N72);
buf BUF1 (N266, N245);
buf BUF1 (N267, N262);
or OR2 (N268, N265, N73);
nor NOR4 (N269, N249, N194, N127, N39);
xor XOR2 (N270, N269, N88);
nand NAND2 (N271, N247, N168);
nor NOR4 (N272, N263, N186, N25, N251);
nor NOR2 (N273, N267, N105);
buf BUF1 (N274, N270);
nor NOR4 (N275, N266, N56, N202, N223);
nor NOR4 (N276, N252, N96, N259, N165);
xor XOR2 (N277, N275, N34);
and AND3 (N278, N276, N190, N194);
not NOT1 (N279, N273);
buf BUF1 (N280, N264);
or OR4 (N281, N272, N241, N221, N21);
nand NAND4 (N282, N277, N243, N279, N82);
buf BUF1 (N283, N195);
nor NOR3 (N284, N274, N159, N24);
nor NOR2 (N285, N280, N280);
and AND3 (N286, N281, N256, N36);
nand NAND4 (N287, N257, N11, N240, N275);
nor NOR4 (N288, N286, N1, N85, N272);
buf BUF1 (N289, N271);
and AND4 (N290, N261, N249, N83, N265);
xor XOR2 (N291, N284, N90);
and AND3 (N292, N268, N64, N76);
xor XOR2 (N293, N282, N121);
xor XOR2 (N294, N285, N67);
not NOT1 (N295, N287);
or OR3 (N296, N292, N156, N93);
or OR3 (N297, N290, N166, N43);
nor NOR3 (N298, N289, N212, N33);
and AND4 (N299, N293, N252, N137, N83);
xor XOR2 (N300, N288, N20);
and AND2 (N301, N291, N29);
and AND4 (N302, N300, N142, N151, N271);
and AND3 (N303, N299, N101, N141);
or OR2 (N304, N296, N255);
buf BUF1 (N305, N283);
nand NAND4 (N306, N302, N111, N71, N257);
nand NAND4 (N307, N301, N185, N110, N141);
and AND4 (N308, N297, N221, N191, N113);
nand NAND3 (N309, N278, N183, N112);
not NOT1 (N310, N306);
not NOT1 (N311, N304);
nor NOR3 (N312, N298, N186, N42);
nand NAND2 (N313, N308, N277);
xor XOR2 (N314, N309, N246);
nor NOR2 (N315, N310, N40);
not NOT1 (N316, N313);
nor NOR2 (N317, N315, N176);
nor NOR2 (N318, N294, N102);
or OR3 (N319, N316, N218, N245);
buf BUF1 (N320, N305);
and AND2 (N321, N317, N269);
buf BUF1 (N322, N311);
xor XOR2 (N323, N307, N263);
not NOT1 (N324, N312);
or OR4 (N325, N319, N306, N283, N295);
not NOT1 (N326, N324);
not NOT1 (N327, N97);
or OR3 (N328, N326, N264, N130);
nor NOR3 (N329, N328, N303, N100);
or OR3 (N330, N257, N148, N54);
and AND4 (N331, N322, N308, N26, N264);
and AND3 (N332, N329, N187, N275);
and AND2 (N333, N318, N230);
and AND4 (N334, N325, N138, N292, N55);
and AND3 (N335, N331, N244, N116);
xor XOR2 (N336, N333, N40);
or OR3 (N337, N323, N32, N318);
not NOT1 (N338, N335);
or OR3 (N339, N332, N229, N115);
nand NAND4 (N340, N330, N70, N287, N253);
buf BUF1 (N341, N340);
or OR3 (N342, N314, N288, N20);
xor XOR2 (N343, N342, N178);
xor XOR2 (N344, N338, N122);
not NOT1 (N345, N327);
xor XOR2 (N346, N336, N227);
not NOT1 (N347, N344);
xor XOR2 (N348, N345, N19);
nand NAND3 (N349, N347, N136, N73);
or OR3 (N350, N337, N1, N34);
nor NOR2 (N351, N346, N34);
or OR2 (N352, N343, N269);
or OR3 (N353, N351, N134, N247);
buf BUF1 (N354, N350);
not NOT1 (N355, N352);
buf BUF1 (N356, N349);
and AND4 (N357, N353, N135, N252, N162);
buf BUF1 (N358, N354);
and AND2 (N359, N339, N135);
buf BUF1 (N360, N355);
buf BUF1 (N361, N360);
or OR3 (N362, N341, N216, N218);
and AND3 (N363, N361, N249, N240);
and AND2 (N364, N334, N203);
and AND2 (N365, N320, N182);
buf BUF1 (N366, N364);
xor XOR2 (N367, N359, N104);
nand NAND3 (N368, N321, N337, N121);
nand NAND3 (N369, N356, N122, N184);
not NOT1 (N370, N368);
buf BUF1 (N371, N369);
nor NOR4 (N372, N362, N343, N34, N45);
nor NOR3 (N373, N348, N25, N68);
buf BUF1 (N374, N372);
nor NOR2 (N375, N366, N348);
nand NAND3 (N376, N373, N258, N97);
xor XOR2 (N377, N365, N160);
xor XOR2 (N378, N358, N240);
buf BUF1 (N379, N370);
nor NOR3 (N380, N374, N358, N224);
not NOT1 (N381, N377);
buf BUF1 (N382, N363);
not NOT1 (N383, N379);
or OR2 (N384, N378, N209);
nor NOR2 (N385, N357, N237);
nand NAND3 (N386, N371, N103, N337);
and AND3 (N387, N381, N33, N315);
xor XOR2 (N388, N380, N383);
or OR2 (N389, N116, N365);
not NOT1 (N390, N376);
xor XOR2 (N391, N382, N85);
nor NOR2 (N392, N388, N87);
xor XOR2 (N393, N375, N376);
not NOT1 (N394, N367);
and AND4 (N395, N385, N105, N219, N93);
buf BUF1 (N396, N391);
nand NAND3 (N397, N387, N40, N213);
not NOT1 (N398, N389);
or OR3 (N399, N392, N385, N51);
buf BUF1 (N400, N398);
not NOT1 (N401, N397);
nor NOR3 (N402, N384, N68, N82);
and AND3 (N403, N400, N366, N266);
nand NAND2 (N404, N402, N32);
and AND3 (N405, N393, N79, N359);
xor XOR2 (N406, N401, N160);
not NOT1 (N407, N404);
nor NOR3 (N408, N403, N336, N66);
nor NOR2 (N409, N395, N56);
buf BUF1 (N410, N406);
buf BUF1 (N411, N407);
and AND2 (N412, N394, N36);
and AND4 (N413, N405, N35, N253, N68);
not NOT1 (N414, N411);
not NOT1 (N415, N399);
nand NAND3 (N416, N412, N24, N70);
nand NAND2 (N417, N414, N281);
xor XOR2 (N418, N409, N145);
xor XOR2 (N419, N396, N212);
nor NOR2 (N420, N386, N253);
nand NAND3 (N421, N408, N302, N89);
nand NAND3 (N422, N417, N212, N8);
nand NAND4 (N423, N415, N189, N352, N350);
nor NOR3 (N424, N416, N297, N30);
not NOT1 (N425, N422);
xor XOR2 (N426, N413, N237);
nor NOR2 (N427, N390, N394);
xor XOR2 (N428, N420, N34);
nor NOR4 (N429, N427, N7, N62, N307);
or OR3 (N430, N419, N142, N46);
xor XOR2 (N431, N421, N111);
xor XOR2 (N432, N430, N318);
xor XOR2 (N433, N429, N62);
xor XOR2 (N434, N432, N320);
buf BUF1 (N435, N431);
not NOT1 (N436, N423);
nand NAND4 (N437, N425, N412, N284, N352);
xor XOR2 (N438, N418, N224);
buf BUF1 (N439, N433);
or OR4 (N440, N435, N411, N418, N108);
nor NOR2 (N441, N410, N379);
nor NOR2 (N442, N440, N278);
buf BUF1 (N443, N442);
buf BUF1 (N444, N438);
nand NAND2 (N445, N444, N125);
not NOT1 (N446, N445);
and AND3 (N447, N437, N29, N238);
buf BUF1 (N448, N424);
not NOT1 (N449, N448);
xor XOR2 (N450, N426, N340);
and AND3 (N451, N428, N49, N111);
nor NOR3 (N452, N446, N79, N304);
not NOT1 (N453, N451);
nand NAND4 (N454, N452, N140, N223, N177);
xor XOR2 (N455, N447, N413);
and AND2 (N456, N439, N403);
buf BUF1 (N457, N436);
nor NOR4 (N458, N450, N425, N410, N75);
nand NAND2 (N459, N449, N144);
or OR4 (N460, N441, N311, N22, N205);
nand NAND2 (N461, N454, N293);
and AND3 (N462, N460, N29, N317);
nand NAND2 (N463, N434, N359);
buf BUF1 (N464, N462);
xor XOR2 (N465, N443, N280);
and AND4 (N466, N455, N441, N158, N443);
nor NOR4 (N467, N465, N50, N329, N367);
nor NOR2 (N468, N459, N244);
xor XOR2 (N469, N466, N448);
and AND3 (N470, N467, N48, N79);
or OR2 (N471, N463, N249);
not NOT1 (N472, N453);
xor XOR2 (N473, N456, N428);
nor NOR4 (N474, N458, N181, N311, N165);
not NOT1 (N475, N457);
not NOT1 (N476, N471);
and AND2 (N477, N461, N286);
and AND3 (N478, N475, N387, N181);
and AND3 (N479, N472, N424, N20);
or OR2 (N480, N478, N256);
nand NAND2 (N481, N470, N394);
not NOT1 (N482, N474);
and AND4 (N483, N481, N14, N250, N101);
nor NOR4 (N484, N477, N383, N37, N8);
nor NOR3 (N485, N482, N393, N405);
xor XOR2 (N486, N473, N114);
not NOT1 (N487, N476);
buf BUF1 (N488, N486);
xor XOR2 (N489, N488, N196);
not NOT1 (N490, N483);
buf BUF1 (N491, N469);
xor XOR2 (N492, N490, N291);
buf BUF1 (N493, N485);
nor NOR4 (N494, N491, N254, N178, N403);
xor XOR2 (N495, N492, N466);
and AND2 (N496, N480, N375);
buf BUF1 (N497, N493);
xor XOR2 (N498, N489, N213);
or OR2 (N499, N487, N82);
not NOT1 (N500, N484);
and AND4 (N501, N496, N342, N437, N67);
nand NAND3 (N502, N495, N185, N301);
nor NOR2 (N503, N501, N366);
buf BUF1 (N504, N497);
buf BUF1 (N505, N498);
not NOT1 (N506, N464);
nand NAND2 (N507, N500, N199);
not NOT1 (N508, N504);
nor NOR4 (N509, N506, N232, N57, N45);
not NOT1 (N510, N505);
nand NAND3 (N511, N479, N453, N225);
or OR3 (N512, N508, N276, N99);
or OR2 (N513, N510, N304);
or OR4 (N514, N513, N28, N439, N339);
nand NAND3 (N515, N494, N67, N332);
xor XOR2 (N516, N509, N312);
or OR4 (N517, N514, N169, N345, N194);
not NOT1 (N518, N503);
and AND3 (N519, N468, N115, N513);
xor XOR2 (N520, N518, N191);
and AND2 (N521, N520, N510);
nor NOR2 (N522, N507, N161);
xor XOR2 (N523, N499, N83);
not NOT1 (N524, N519);
or OR2 (N525, N511, N109);
not NOT1 (N526, N523);
not NOT1 (N527, N526);
or OR2 (N528, N521, N358);
nand NAND4 (N529, N515, N174, N299, N9);
xor XOR2 (N530, N529, N498);
nand NAND3 (N531, N527, N165, N511);
not NOT1 (N532, N531);
buf BUF1 (N533, N522);
nand NAND4 (N534, N502, N276, N401, N279);
and AND2 (N535, N517, N433);
not NOT1 (N536, N524);
xor XOR2 (N537, N530, N312);
nor NOR2 (N538, N512, N430);
nor NOR2 (N539, N538, N30);
and AND4 (N540, N535, N273, N16, N240);
or OR4 (N541, N539, N523, N201, N385);
nand NAND3 (N542, N541, N458, N49);
buf BUF1 (N543, N534);
xor XOR2 (N544, N536, N42);
or OR4 (N545, N528, N409, N505, N135);
xor XOR2 (N546, N516, N267);
not NOT1 (N547, N525);
or OR3 (N548, N543, N256, N247);
not NOT1 (N549, N544);
nand NAND4 (N550, N540, N180, N77, N196);
not NOT1 (N551, N547);
or OR4 (N552, N545, N24, N524, N374);
nor NOR3 (N553, N533, N114, N256);
not NOT1 (N554, N550);
or OR3 (N555, N553, N508, N406);
buf BUF1 (N556, N532);
xor XOR2 (N557, N555, N22);
xor XOR2 (N558, N552, N223);
nor NOR3 (N559, N537, N434, N297);
and AND3 (N560, N551, N358, N387);
nand NAND4 (N561, N558, N522, N308, N388);
nand NAND2 (N562, N559, N160);
or OR4 (N563, N548, N427, N346, N442);
and AND2 (N564, N557, N135);
nand NAND3 (N565, N563, N420, N304);
not NOT1 (N566, N542);
and AND4 (N567, N561, N420, N355, N527);
or OR4 (N568, N556, N234, N264, N187);
xor XOR2 (N569, N565, N279);
or OR3 (N570, N546, N107, N224);
not NOT1 (N571, N570);
nand NAND4 (N572, N560, N323, N136, N274);
or OR3 (N573, N549, N422, N324);
xor XOR2 (N574, N569, N382);
xor XOR2 (N575, N573, N381);
xor XOR2 (N576, N572, N123);
not NOT1 (N577, N575);
nor NOR2 (N578, N566, N391);
and AND3 (N579, N554, N254, N192);
nor NOR4 (N580, N568, N3, N428, N21);
and AND4 (N581, N579, N561, N57, N247);
xor XOR2 (N582, N578, N304);
buf BUF1 (N583, N581);
nor NOR3 (N584, N562, N370, N125);
or OR4 (N585, N564, N257, N12, N415);
and AND2 (N586, N582, N27);
or OR4 (N587, N577, N499, N42, N138);
not NOT1 (N588, N583);
or OR2 (N589, N567, N186);
or OR4 (N590, N574, N346, N347, N130);
buf BUF1 (N591, N586);
nor NOR3 (N592, N588, N59, N1);
xor XOR2 (N593, N589, N196);
or OR2 (N594, N585, N321);
nor NOR2 (N595, N571, N303);
and AND2 (N596, N580, N561);
and AND2 (N597, N595, N306);
xor XOR2 (N598, N590, N61);
and AND2 (N599, N597, N566);
and AND4 (N600, N584, N523, N485, N444);
nor NOR4 (N601, N600, N385, N598, N100);
not NOT1 (N602, N175);
xor XOR2 (N603, N599, N307);
and AND3 (N604, N602, N485, N468);
nor NOR4 (N605, N594, N87, N502, N242);
xor XOR2 (N606, N593, N44);
or OR3 (N607, N604, N22, N194);
xor XOR2 (N608, N607, N248);
and AND2 (N609, N608, N307);
buf BUF1 (N610, N603);
xor XOR2 (N611, N610, N422);
not NOT1 (N612, N611);
and AND4 (N613, N591, N333, N577, N552);
xor XOR2 (N614, N606, N165);
buf BUF1 (N615, N601);
nor NOR2 (N616, N612, N274);
or OR4 (N617, N609, N218, N378, N396);
not NOT1 (N618, N613);
or OR2 (N619, N605, N188);
nor NOR4 (N620, N616, N481, N609, N475);
and AND4 (N621, N614, N476, N320, N398);
and AND3 (N622, N617, N114, N185);
not NOT1 (N623, N615);
nand NAND4 (N624, N620, N52, N521, N450);
xor XOR2 (N625, N587, N64);
and AND4 (N626, N596, N177, N278, N454);
xor XOR2 (N627, N621, N215);
nor NOR4 (N628, N624, N134, N230, N462);
xor XOR2 (N629, N618, N615);
nand NAND4 (N630, N622, N312, N407, N329);
or OR2 (N631, N628, N542);
or OR2 (N632, N627, N103);
xor XOR2 (N633, N625, N448);
buf BUF1 (N634, N630);
not NOT1 (N635, N619);
and AND4 (N636, N633, N346, N487, N232);
not NOT1 (N637, N629);
nand NAND2 (N638, N576, N553);
and AND2 (N639, N623, N260);
and AND2 (N640, N635, N236);
or OR4 (N641, N638, N255, N154, N449);
not NOT1 (N642, N637);
buf BUF1 (N643, N640);
not NOT1 (N644, N626);
xor XOR2 (N645, N592, N175);
nand NAND2 (N646, N631, N542);
and AND2 (N647, N643, N7);
xor XOR2 (N648, N646, N526);
buf BUF1 (N649, N644);
nand NAND4 (N650, N641, N495, N33, N442);
nand NAND3 (N651, N650, N296, N500);
xor XOR2 (N652, N632, N179);
nor NOR4 (N653, N652, N114, N394, N13);
buf BUF1 (N654, N642);
nand NAND4 (N655, N653, N267, N164, N111);
or OR3 (N656, N654, N594, N461);
nor NOR3 (N657, N647, N61, N349);
and AND4 (N658, N649, N105, N91, N296);
buf BUF1 (N659, N657);
or OR3 (N660, N634, N224, N111);
xor XOR2 (N661, N636, N561);
nand NAND2 (N662, N661, N528);
nand NAND2 (N663, N662, N409);
xor XOR2 (N664, N660, N164);
not NOT1 (N665, N651);
or OR3 (N666, N659, N284, N520);
and AND4 (N667, N664, N76, N367, N380);
nor NOR4 (N668, N656, N123, N180, N381);
xor XOR2 (N669, N645, N41);
xor XOR2 (N670, N666, N649);
or OR2 (N671, N670, N593);
xor XOR2 (N672, N665, N159);
and AND4 (N673, N639, N619, N521, N305);
and AND2 (N674, N673, N512);
xor XOR2 (N675, N671, N266);
not NOT1 (N676, N663);
nor NOR2 (N677, N667, N132);
and AND4 (N678, N676, N670, N549, N306);
and AND4 (N679, N668, N458, N227, N568);
nor NOR4 (N680, N658, N222, N556, N647);
not NOT1 (N681, N648);
not NOT1 (N682, N669);
buf BUF1 (N683, N681);
or OR3 (N684, N683, N639, N338);
nor NOR4 (N685, N675, N254, N241, N265);
and AND4 (N686, N680, N216, N542, N250);
and AND4 (N687, N674, N189, N626, N241);
nor NOR2 (N688, N677, N547);
buf BUF1 (N689, N682);
nor NOR4 (N690, N679, N37, N196, N621);
and AND3 (N691, N685, N439, N609);
buf BUF1 (N692, N686);
and AND3 (N693, N678, N440, N569);
not NOT1 (N694, N672);
and AND2 (N695, N684, N444);
or OR3 (N696, N693, N571, N613);
xor XOR2 (N697, N687, N49);
nor NOR4 (N698, N694, N510, N269, N690);
nor NOR2 (N699, N43, N30);
nand NAND4 (N700, N655, N540, N444, N182);
nor NOR4 (N701, N689, N102, N59, N420);
and AND4 (N702, N699, N482, N73, N411);
and AND4 (N703, N702, N452, N40, N269);
and AND3 (N704, N703, N235, N253);
not NOT1 (N705, N701);
or OR2 (N706, N705, N454);
not NOT1 (N707, N696);
buf BUF1 (N708, N706);
not NOT1 (N709, N707);
nor NOR2 (N710, N691, N413);
and AND3 (N711, N708, N77, N409);
nand NAND4 (N712, N709, N683, N672, N540);
xor XOR2 (N713, N695, N72);
xor XOR2 (N714, N711, N294);
and AND2 (N715, N698, N110);
xor XOR2 (N716, N697, N500);
not NOT1 (N717, N700);
nand NAND3 (N718, N717, N303, N338);
xor XOR2 (N719, N712, N13);
buf BUF1 (N720, N688);
and AND2 (N721, N704, N624);
nand NAND4 (N722, N713, N653, N680, N404);
nand NAND4 (N723, N692, N500, N266, N329);
xor XOR2 (N724, N719, N519);
and AND4 (N725, N721, N352, N65, N384);
buf BUF1 (N726, N722);
and AND2 (N727, N710, N697);
nor NOR4 (N728, N725, N256, N679, N270);
nor NOR2 (N729, N727, N439);
and AND2 (N730, N728, N40);
and AND3 (N731, N718, N681, N439);
buf BUF1 (N732, N730);
or OR4 (N733, N731, N248, N227, N671);
buf BUF1 (N734, N723);
nand NAND4 (N735, N715, N478, N121, N615);
or OR4 (N736, N734, N338, N297, N260);
xor XOR2 (N737, N729, N40);
not NOT1 (N738, N726);
nand NAND4 (N739, N733, N361, N287, N611);
nor NOR3 (N740, N735, N239, N475);
and AND2 (N741, N724, N686);
nor NOR3 (N742, N732, N169, N701);
xor XOR2 (N743, N716, N322);
not NOT1 (N744, N742);
xor XOR2 (N745, N740, N500);
nand NAND2 (N746, N736, N533);
and AND4 (N747, N720, N745, N403, N329);
nor NOR2 (N748, N167, N3);
nor NOR2 (N749, N714, N356);
buf BUF1 (N750, N741);
or OR4 (N751, N746, N241, N652, N572);
nor NOR3 (N752, N739, N228, N716);
nor NOR2 (N753, N748, N460);
or OR4 (N754, N752, N590, N531, N237);
and AND4 (N755, N738, N381, N485, N601);
or OR4 (N756, N747, N656, N349, N152);
xor XOR2 (N757, N743, N476);
xor XOR2 (N758, N744, N491);
nor NOR3 (N759, N751, N747, N236);
nor NOR3 (N760, N758, N221, N7);
and AND4 (N761, N753, N604, N329, N555);
or OR3 (N762, N749, N236, N303);
or OR3 (N763, N757, N356, N601);
and AND2 (N764, N754, N101);
not NOT1 (N765, N763);
or OR3 (N766, N737, N550, N225);
buf BUF1 (N767, N762);
xor XOR2 (N768, N760, N455);
nor NOR4 (N769, N756, N337, N214, N375);
nor NOR2 (N770, N766, N733);
nor NOR2 (N771, N755, N567);
nor NOR3 (N772, N771, N102, N284);
buf BUF1 (N773, N769);
or OR4 (N774, N768, N63, N678, N345);
buf BUF1 (N775, N767);
xor XOR2 (N776, N770, N262);
nor NOR2 (N777, N765, N750);
nor NOR2 (N778, N485, N540);
or OR4 (N779, N764, N49, N696, N707);
xor XOR2 (N780, N775, N435);
or OR2 (N781, N774, N485);
not NOT1 (N782, N772);
or OR4 (N783, N759, N60, N432, N441);
nand NAND4 (N784, N778, N448, N755, N168);
nand NAND2 (N785, N779, N350);
buf BUF1 (N786, N777);
xor XOR2 (N787, N785, N389);
or OR4 (N788, N773, N104, N359, N685);
and AND3 (N789, N761, N443, N242);
buf BUF1 (N790, N782);
and AND4 (N791, N789, N226, N309, N426);
nor NOR2 (N792, N788, N239);
buf BUF1 (N793, N780);
nor NOR3 (N794, N781, N128, N635);
buf BUF1 (N795, N791);
buf BUF1 (N796, N792);
not NOT1 (N797, N787);
not NOT1 (N798, N784);
buf BUF1 (N799, N798);
xor XOR2 (N800, N786, N166);
nor NOR4 (N801, N799, N723, N31, N570);
buf BUF1 (N802, N800);
nor NOR2 (N803, N797, N304);
nor NOR2 (N804, N801, N727);
buf BUF1 (N805, N793);
nor NOR2 (N806, N776, N154);
nor NOR4 (N807, N783, N382, N432, N560);
or OR3 (N808, N806, N584, N542);
xor XOR2 (N809, N807, N62);
not NOT1 (N810, N796);
nor NOR4 (N811, N803, N110, N339, N172);
nor NOR4 (N812, N810, N796, N782, N663);
and AND4 (N813, N812, N222, N546, N126);
or OR4 (N814, N809, N730, N566, N493);
and AND3 (N815, N808, N186, N382);
buf BUF1 (N816, N815);
not NOT1 (N817, N811);
nor NOR2 (N818, N795, N511);
buf BUF1 (N819, N813);
or OR3 (N820, N819, N789, N228);
not NOT1 (N821, N820);
buf BUF1 (N822, N804);
nand NAND3 (N823, N818, N71, N99);
xor XOR2 (N824, N817, N403);
nand NAND2 (N825, N821, N341);
nand NAND2 (N826, N816, N214);
and AND3 (N827, N824, N385, N61);
or OR3 (N828, N794, N95, N28);
nand NAND4 (N829, N814, N177, N787, N562);
xor XOR2 (N830, N805, N359);
not NOT1 (N831, N829);
not NOT1 (N832, N825);
or OR4 (N833, N802, N438, N370, N218);
not NOT1 (N834, N826);
nor NOR3 (N835, N831, N831, N762);
nor NOR3 (N836, N790, N223, N457);
nand NAND3 (N837, N833, N520, N710);
xor XOR2 (N838, N828, N697);
or OR3 (N839, N822, N210, N190);
or OR3 (N840, N834, N284, N180);
nor NOR4 (N841, N832, N829, N726, N312);
buf BUF1 (N842, N827);
buf BUF1 (N843, N823);
and AND3 (N844, N840, N375, N137);
nor NOR4 (N845, N836, N599, N202, N8);
buf BUF1 (N846, N841);
nor NOR2 (N847, N846, N677);
or OR3 (N848, N847, N97, N359);
and AND4 (N849, N842, N613, N371, N639);
not NOT1 (N850, N844);
buf BUF1 (N851, N849);
or OR2 (N852, N845, N268);
nand NAND2 (N853, N839, N792);
nand NAND4 (N854, N835, N589, N696, N573);
buf BUF1 (N855, N852);
nand NAND3 (N856, N837, N517, N731);
not NOT1 (N857, N843);
and AND4 (N858, N855, N682, N182, N733);
buf BUF1 (N859, N830);
buf BUF1 (N860, N851);
nand NAND4 (N861, N848, N477, N606, N785);
or OR4 (N862, N853, N783, N489, N237);
xor XOR2 (N863, N862, N556);
buf BUF1 (N864, N838);
and AND4 (N865, N854, N848, N809, N453);
and AND2 (N866, N863, N209);
nor NOR3 (N867, N866, N418, N755);
and AND2 (N868, N865, N180);
xor XOR2 (N869, N868, N669);
nor NOR2 (N870, N861, N838);
nor NOR3 (N871, N850, N152, N343);
not NOT1 (N872, N867);
or OR2 (N873, N870, N210);
not NOT1 (N874, N860);
nor NOR3 (N875, N873, N29, N585);
nand NAND4 (N876, N874, N527, N547, N73);
nor NOR4 (N877, N859, N178, N163, N462);
not NOT1 (N878, N872);
and AND3 (N879, N858, N768, N272);
and AND2 (N880, N875, N113);
not NOT1 (N881, N880);
buf BUF1 (N882, N856);
not NOT1 (N883, N871);
or OR2 (N884, N857, N668);
and AND2 (N885, N881, N556);
and AND3 (N886, N877, N648, N148);
nand NAND4 (N887, N876, N511, N296, N406);
and AND2 (N888, N882, N29);
nor NOR4 (N889, N885, N736, N290, N601);
not NOT1 (N890, N869);
nor NOR4 (N891, N884, N190, N617, N497);
nand NAND4 (N892, N891, N593, N34, N241);
xor XOR2 (N893, N883, N96);
nand NAND3 (N894, N887, N623, N655);
or OR3 (N895, N893, N456, N626);
and AND2 (N896, N864, N426);
xor XOR2 (N897, N894, N377);
and AND2 (N898, N890, N649);
not NOT1 (N899, N892);
or OR3 (N900, N888, N3, N482);
nor NOR4 (N901, N900, N593, N658, N474);
nor NOR2 (N902, N896, N356);
xor XOR2 (N903, N886, N48);
or OR4 (N904, N902, N389, N668, N625);
nor NOR4 (N905, N879, N23, N609, N482);
and AND3 (N906, N901, N148, N654);
nor NOR3 (N907, N878, N328, N11);
nand NAND3 (N908, N904, N200, N351);
nand NAND3 (N909, N908, N869, N547);
or OR4 (N910, N895, N577, N67, N251);
or OR3 (N911, N889, N781, N865);
nand NAND4 (N912, N898, N230, N603, N708);
not NOT1 (N913, N899);
nor NOR4 (N914, N907, N545, N448, N648);
buf BUF1 (N915, N903);
or OR3 (N916, N905, N98, N406);
xor XOR2 (N917, N909, N791);
or OR3 (N918, N916, N816, N196);
or OR4 (N919, N912, N583, N536, N594);
nand NAND4 (N920, N915, N886, N261, N75);
or OR3 (N921, N917, N831, N220);
not NOT1 (N922, N911);
buf BUF1 (N923, N921);
not NOT1 (N924, N910);
and AND3 (N925, N913, N757, N595);
buf BUF1 (N926, N924);
buf BUF1 (N927, N926);
and AND4 (N928, N920, N269, N20, N684);
nand NAND4 (N929, N897, N42, N147, N412);
nand NAND4 (N930, N923, N108, N719, N617);
buf BUF1 (N931, N914);
nand NAND2 (N932, N906, N676);
and AND3 (N933, N927, N462, N235);
nand NAND4 (N934, N922, N10, N247, N292);
and AND2 (N935, N933, N77);
nand NAND4 (N936, N935, N381, N924, N470);
nor NOR2 (N937, N936, N106);
buf BUF1 (N938, N937);
or OR3 (N939, N931, N552, N176);
nor NOR2 (N940, N934, N1);
xor XOR2 (N941, N930, N712);
buf BUF1 (N942, N939);
not NOT1 (N943, N928);
nand NAND2 (N944, N943, N691);
xor XOR2 (N945, N925, N135);
buf BUF1 (N946, N938);
nor NOR2 (N947, N932, N798);
nand NAND4 (N948, N919, N905, N920, N239);
buf BUF1 (N949, N946);
buf BUF1 (N950, N948);
xor XOR2 (N951, N947, N635);
nand NAND4 (N952, N929, N289, N357, N311);
and AND2 (N953, N918, N405);
nand NAND3 (N954, N942, N279, N366);
or OR4 (N955, N941, N176, N235, N468);
xor XOR2 (N956, N950, N564);
or OR2 (N957, N944, N781);
nor NOR3 (N958, N956, N899, N521);
buf BUF1 (N959, N957);
or OR3 (N960, N958, N474, N103);
buf BUF1 (N961, N940);
buf BUF1 (N962, N955);
nor NOR2 (N963, N951, N609);
and AND2 (N964, N962, N42);
or OR2 (N965, N960, N783);
not NOT1 (N966, N963);
and AND3 (N967, N949, N566, N813);
and AND3 (N968, N961, N151, N805);
nor NOR3 (N969, N954, N796, N732);
buf BUF1 (N970, N953);
and AND3 (N971, N968, N563, N170);
or OR3 (N972, N971, N956, N208);
not NOT1 (N973, N966);
and AND2 (N974, N965, N160);
buf BUF1 (N975, N969);
not NOT1 (N976, N975);
not NOT1 (N977, N973);
and AND2 (N978, N964, N509);
and AND3 (N979, N945, N112, N310);
not NOT1 (N980, N979);
xor XOR2 (N981, N952, N480);
nor NOR4 (N982, N977, N936, N200, N731);
nand NAND3 (N983, N980, N302, N118);
and AND4 (N984, N983, N506, N889, N971);
buf BUF1 (N985, N984);
xor XOR2 (N986, N972, N426);
nor NOR4 (N987, N974, N562, N60, N758);
xor XOR2 (N988, N982, N124);
not NOT1 (N989, N985);
not NOT1 (N990, N976);
or OR2 (N991, N990, N797);
or OR2 (N992, N978, N636);
or OR3 (N993, N970, N383, N79);
xor XOR2 (N994, N992, N141);
nor NOR3 (N995, N987, N154, N51);
or OR4 (N996, N995, N682, N827, N111);
not NOT1 (N997, N967);
and AND4 (N998, N991, N899, N957, N165);
nand NAND3 (N999, N986, N506, N502);
and AND3 (N1000, N959, N215, N202);
or OR2 (N1001, N989, N688);
not NOT1 (N1002, N996);
not NOT1 (N1003, N988);
xor XOR2 (N1004, N1000, N170);
or OR2 (N1005, N997, N316);
and AND3 (N1006, N981, N249, N527);
buf BUF1 (N1007, N993);
or OR2 (N1008, N1005, N858);
nor NOR4 (N1009, N998, N412, N596, N308);
not NOT1 (N1010, N1006);
or OR2 (N1011, N994, N257);
nand NAND3 (N1012, N1010, N324, N968);
xor XOR2 (N1013, N1004, N734);
nor NOR2 (N1014, N1009, N610);
buf BUF1 (N1015, N1011);
xor XOR2 (N1016, N1014, N14);
nand NAND2 (N1017, N1016, N579);
nor NOR2 (N1018, N1001, N304);
or OR3 (N1019, N1017, N485, N456);
nand NAND3 (N1020, N1019, N788, N591);
buf BUF1 (N1021, N1018);
xor XOR2 (N1022, N1008, N819);
or OR4 (N1023, N1003, N459, N212, N541);
and AND2 (N1024, N1002, N3);
nand NAND3 (N1025, N1023, N681, N430);
nor NOR4 (N1026, N1012, N421, N27, N826);
and AND2 (N1027, N1007, N1018);
buf BUF1 (N1028, N1015);
or OR4 (N1029, N1020, N790, N341, N352);
nor NOR4 (N1030, N1027, N804, N71, N884);
not NOT1 (N1031, N1025);
xor XOR2 (N1032, N1022, N855);
and AND2 (N1033, N1030, N507);
nand NAND3 (N1034, N1013, N523, N208);
nor NOR2 (N1035, N1028, N381);
and AND3 (N1036, N1031, N103, N383);
not NOT1 (N1037, N1034);
xor XOR2 (N1038, N1026, N406);
xor XOR2 (N1039, N1029, N627);
buf BUF1 (N1040, N1035);
and AND3 (N1041, N1037, N680, N517);
not NOT1 (N1042, N1033);
nor NOR4 (N1043, N999, N880, N25, N958);
buf BUF1 (N1044, N1041);
xor XOR2 (N1045, N1032, N471);
not NOT1 (N1046, N1024);
and AND3 (N1047, N1038, N228, N848);
nand NAND3 (N1048, N1046, N767, N524);
buf BUF1 (N1049, N1036);
nor NOR3 (N1050, N1043, N371, N95);
or OR3 (N1051, N1039, N551, N695);
or OR3 (N1052, N1045, N252, N981);
and AND3 (N1053, N1042, N756, N197);
and AND4 (N1054, N1021, N678, N320, N137);
nor NOR3 (N1055, N1051, N275, N830);
nand NAND2 (N1056, N1044, N58);
nor NOR3 (N1057, N1056, N848, N137);
or OR3 (N1058, N1055, N126, N914);
and AND3 (N1059, N1050, N1044, N977);
buf BUF1 (N1060, N1048);
nor NOR3 (N1061, N1054, N545, N673);
not NOT1 (N1062, N1061);
buf BUF1 (N1063, N1040);
nor NOR4 (N1064, N1063, N219, N210, N752);
not NOT1 (N1065, N1058);
xor XOR2 (N1066, N1049, N174);
xor XOR2 (N1067, N1057, N828);
xor XOR2 (N1068, N1053, N126);
buf BUF1 (N1069, N1068);
or OR3 (N1070, N1059, N1024, N907);
or OR2 (N1071, N1060, N805);
nor NOR3 (N1072, N1067, N552, N438);
nor NOR4 (N1073, N1072, N492, N561, N369);
buf BUF1 (N1074, N1064);
not NOT1 (N1075, N1047);
nand NAND3 (N1076, N1074, N31, N157);
nor NOR3 (N1077, N1076, N675, N758);
nand NAND4 (N1078, N1066, N76, N519, N148);
xor XOR2 (N1079, N1071, N856);
not NOT1 (N1080, N1073);
nor NOR3 (N1081, N1079, N130, N134);
nand NAND3 (N1082, N1078, N536, N328);
and AND3 (N1083, N1052, N270, N732);
not NOT1 (N1084, N1080);
buf BUF1 (N1085, N1084);
nand NAND4 (N1086, N1081, N675, N512, N1049);
not NOT1 (N1087, N1082);
nand NAND2 (N1088, N1070, N959);
buf BUF1 (N1089, N1088);
nand NAND2 (N1090, N1087, N664);
nor NOR2 (N1091, N1062, N692);
xor XOR2 (N1092, N1065, N803);
not NOT1 (N1093, N1075);
not NOT1 (N1094, N1093);
and AND4 (N1095, N1086, N556, N459, N180);
buf BUF1 (N1096, N1089);
or OR2 (N1097, N1083, N124);
xor XOR2 (N1098, N1085, N789);
nor NOR3 (N1099, N1091, N1035, N442);
and AND4 (N1100, N1097, N79, N541, N134);
and AND3 (N1101, N1092, N358, N460);
buf BUF1 (N1102, N1101);
xor XOR2 (N1103, N1069, N839);
xor XOR2 (N1104, N1095, N254);
and AND4 (N1105, N1102, N309, N393, N810);
nor NOR3 (N1106, N1105, N1046, N581);
buf BUF1 (N1107, N1099);
xor XOR2 (N1108, N1090, N949);
nor NOR2 (N1109, N1107, N732);
not NOT1 (N1110, N1106);
not NOT1 (N1111, N1094);
or OR3 (N1112, N1110, N115, N1021);
nand NAND3 (N1113, N1096, N583, N981);
or OR2 (N1114, N1104, N470);
nor NOR2 (N1115, N1108, N207);
and AND4 (N1116, N1115, N735, N435, N198);
nand NAND4 (N1117, N1113, N485, N329, N1053);
or OR2 (N1118, N1109, N719);
xor XOR2 (N1119, N1100, N997);
not NOT1 (N1120, N1112);
or OR3 (N1121, N1077, N47, N77);
nor NOR2 (N1122, N1119, N696);
not NOT1 (N1123, N1118);
buf BUF1 (N1124, N1123);
and AND3 (N1125, N1117, N497, N143);
xor XOR2 (N1126, N1111, N1116);
not NOT1 (N1127, N333);
buf BUF1 (N1128, N1098);
or OR3 (N1129, N1124, N40, N824);
or OR4 (N1130, N1122, N603, N1055, N446);
not NOT1 (N1131, N1130);
not NOT1 (N1132, N1126);
nor NOR4 (N1133, N1125, N114, N962, N618);
or OR2 (N1134, N1131, N796);
and AND3 (N1135, N1120, N3, N932);
and AND3 (N1136, N1132, N833, N1013);
or OR3 (N1137, N1129, N580, N203);
xor XOR2 (N1138, N1135, N1131);
and AND4 (N1139, N1103, N115, N309, N207);
buf BUF1 (N1140, N1139);
and AND4 (N1141, N1127, N642, N987, N241);
buf BUF1 (N1142, N1114);
nor NOR2 (N1143, N1137, N956);
xor XOR2 (N1144, N1143, N142);
and AND2 (N1145, N1140, N1115);
buf BUF1 (N1146, N1136);
not NOT1 (N1147, N1121);
buf BUF1 (N1148, N1138);
or OR3 (N1149, N1145, N242, N554);
xor XOR2 (N1150, N1141, N746);
not NOT1 (N1151, N1150);
nor NOR3 (N1152, N1142, N354, N186);
nor NOR3 (N1153, N1147, N71, N281);
nor NOR2 (N1154, N1134, N481);
xor XOR2 (N1155, N1151, N856);
or OR4 (N1156, N1149, N448, N1124, N197);
xor XOR2 (N1157, N1152, N1069);
not NOT1 (N1158, N1148);
nor NOR4 (N1159, N1153, N5, N381, N466);
not NOT1 (N1160, N1146);
not NOT1 (N1161, N1158);
or OR4 (N1162, N1144, N839, N95, N1090);
not NOT1 (N1163, N1156);
and AND4 (N1164, N1133, N1100, N534, N549);
not NOT1 (N1165, N1161);
buf BUF1 (N1166, N1128);
and AND3 (N1167, N1162, N825, N14);
not NOT1 (N1168, N1154);
nand NAND4 (N1169, N1159, N765, N253, N576);
and AND2 (N1170, N1168, N620);
not NOT1 (N1171, N1170);
buf BUF1 (N1172, N1155);
xor XOR2 (N1173, N1171, N510);
not NOT1 (N1174, N1160);
nor NOR4 (N1175, N1166, N333, N283, N775);
nand NAND4 (N1176, N1172, N1018, N192, N999);
or OR3 (N1177, N1174, N180, N45);
not NOT1 (N1178, N1163);
or OR2 (N1179, N1173, N82);
not NOT1 (N1180, N1178);
xor XOR2 (N1181, N1167, N315);
and AND2 (N1182, N1165, N1041);
not NOT1 (N1183, N1169);
nor NOR2 (N1184, N1164, N1124);
or OR3 (N1185, N1183, N1038, N396);
or OR3 (N1186, N1157, N879, N825);
or OR2 (N1187, N1182, N356);
or OR3 (N1188, N1177, N95, N104);
xor XOR2 (N1189, N1176, N233);
or OR4 (N1190, N1188, N176, N798, N739);
nor NOR3 (N1191, N1185, N233, N1054);
nor NOR2 (N1192, N1187, N813);
nand NAND4 (N1193, N1192, N314, N165, N210);
buf BUF1 (N1194, N1189);
xor XOR2 (N1195, N1179, N1025);
xor XOR2 (N1196, N1193, N1162);
xor XOR2 (N1197, N1175, N311);
xor XOR2 (N1198, N1184, N601);
or OR2 (N1199, N1186, N197);
nor NOR3 (N1200, N1198, N396, N448);
or OR4 (N1201, N1196, N972, N354, N959);
not NOT1 (N1202, N1195);
xor XOR2 (N1203, N1180, N264);
or OR2 (N1204, N1191, N513);
buf BUF1 (N1205, N1201);
and AND4 (N1206, N1199, N6, N1135, N135);
nor NOR3 (N1207, N1190, N485, N361);
or OR4 (N1208, N1202, N231, N892, N335);
not NOT1 (N1209, N1205);
nor NOR2 (N1210, N1206, N1091);
nor NOR3 (N1211, N1208, N502, N632);
and AND3 (N1212, N1194, N920, N726);
and AND3 (N1213, N1210, N417, N388);
not NOT1 (N1214, N1212);
or OR4 (N1215, N1200, N319, N870, N633);
nand NAND2 (N1216, N1204, N873);
buf BUF1 (N1217, N1214);
buf BUF1 (N1218, N1181);
xor XOR2 (N1219, N1209, N1148);
buf BUF1 (N1220, N1203);
and AND3 (N1221, N1215, N949, N14);
or OR4 (N1222, N1207, N432, N1083, N401);
nor NOR2 (N1223, N1211, N1158);
or OR3 (N1224, N1197, N1126, N202);
or OR2 (N1225, N1213, N321);
xor XOR2 (N1226, N1218, N580);
buf BUF1 (N1227, N1224);
nor NOR2 (N1228, N1222, N588);
or OR4 (N1229, N1225, N520, N378, N232);
xor XOR2 (N1230, N1223, N103);
xor XOR2 (N1231, N1220, N943);
or OR2 (N1232, N1228, N880);
or OR2 (N1233, N1221, N703);
nand NAND3 (N1234, N1216, N485, N490);
nand NAND2 (N1235, N1217, N646);
buf BUF1 (N1236, N1234);
xor XOR2 (N1237, N1233, N364);
nor NOR2 (N1238, N1219, N520);
nand NAND4 (N1239, N1232, N1047, N29, N663);
xor XOR2 (N1240, N1226, N841);
and AND4 (N1241, N1237, N731, N792, N1128);
and AND2 (N1242, N1229, N288);
nor NOR2 (N1243, N1236, N974);
not NOT1 (N1244, N1235);
nand NAND2 (N1245, N1239, N922);
nor NOR4 (N1246, N1243, N1133, N360, N422);
buf BUF1 (N1247, N1227);
not NOT1 (N1248, N1230);
nor NOR3 (N1249, N1244, N378, N378);
nor NOR2 (N1250, N1247, N833);
xor XOR2 (N1251, N1240, N776);
nor NOR2 (N1252, N1242, N802);
or OR2 (N1253, N1231, N156);
not NOT1 (N1254, N1238);
and AND4 (N1255, N1241, N130, N1214, N336);
and AND4 (N1256, N1251, N516, N224, N1216);
nand NAND4 (N1257, N1245, N1255, N963, N371);
nor NOR2 (N1258, N783, N600);
nand NAND3 (N1259, N1256, N151, N303);
xor XOR2 (N1260, N1253, N667);
nand NAND4 (N1261, N1259, N1143, N1146, N425);
or OR4 (N1262, N1250, N635, N1023, N934);
buf BUF1 (N1263, N1260);
and AND3 (N1264, N1257, N474, N353);
nor NOR3 (N1265, N1249, N182, N1079);
xor XOR2 (N1266, N1261, N1067);
and AND3 (N1267, N1246, N1135, N35);
and AND2 (N1268, N1265, N1145);
not NOT1 (N1269, N1254);
nand NAND4 (N1270, N1263, N408, N419, N438);
buf BUF1 (N1271, N1258);
buf BUF1 (N1272, N1248);
not NOT1 (N1273, N1268);
not NOT1 (N1274, N1267);
and AND2 (N1275, N1271, N464);
nand NAND3 (N1276, N1272, N927, N780);
buf BUF1 (N1277, N1252);
and AND3 (N1278, N1276, N733, N158);
xor XOR2 (N1279, N1269, N68);
xor XOR2 (N1280, N1262, N1020);
not NOT1 (N1281, N1264);
buf BUF1 (N1282, N1274);
buf BUF1 (N1283, N1275);
xor XOR2 (N1284, N1273, N614);
buf BUF1 (N1285, N1283);
xor XOR2 (N1286, N1278, N489);
nand NAND4 (N1287, N1270, N616, N153, N44);
buf BUF1 (N1288, N1287);
and AND4 (N1289, N1286, N162, N1013, N1116);
buf BUF1 (N1290, N1288);
nand NAND4 (N1291, N1285, N919, N911, N637);
not NOT1 (N1292, N1279);
or OR2 (N1293, N1282, N160);
nor NOR4 (N1294, N1284, N754, N763, N235);
not NOT1 (N1295, N1289);
buf BUF1 (N1296, N1291);
and AND4 (N1297, N1296, N469, N143, N678);
xor XOR2 (N1298, N1292, N1009);
nor NOR4 (N1299, N1295, N1070, N1239, N1145);
buf BUF1 (N1300, N1298);
xor XOR2 (N1301, N1280, N322);
and AND2 (N1302, N1299, N83);
not NOT1 (N1303, N1281);
nor NOR3 (N1304, N1293, N726, N380);
and AND2 (N1305, N1297, N17);
not NOT1 (N1306, N1294);
nor NOR4 (N1307, N1302, N321, N1100, N781);
and AND4 (N1308, N1300, N565, N160, N349);
buf BUF1 (N1309, N1290);
nand NAND2 (N1310, N1307, N11);
nor NOR2 (N1311, N1277, N931);
or OR2 (N1312, N1309, N134);
xor XOR2 (N1313, N1305, N237);
buf BUF1 (N1314, N1266);
or OR2 (N1315, N1314, N342);
nand NAND2 (N1316, N1306, N73);
nand NAND2 (N1317, N1313, N724);
or OR4 (N1318, N1301, N717, N1173, N396);
or OR4 (N1319, N1304, N607, N1143, N1280);
not NOT1 (N1320, N1318);
nor NOR3 (N1321, N1303, N1178, N807);
or OR4 (N1322, N1320, N1193, N595, N336);
buf BUF1 (N1323, N1321);
buf BUF1 (N1324, N1312);
nor NOR2 (N1325, N1324, N798);
buf BUF1 (N1326, N1308);
not NOT1 (N1327, N1323);
and AND4 (N1328, N1325, N20, N949, N1198);
and AND4 (N1329, N1317, N1052, N16, N635);
nand NAND3 (N1330, N1326, N478, N696);
or OR4 (N1331, N1329, N669, N494, N842);
nor NOR4 (N1332, N1310, N606, N1204, N727);
buf BUF1 (N1333, N1316);
nand NAND3 (N1334, N1322, N539, N169);
nor NOR4 (N1335, N1332, N429, N596, N831);
nor NOR3 (N1336, N1311, N294, N238);
xor XOR2 (N1337, N1334, N692);
nor NOR3 (N1338, N1319, N755, N407);
xor XOR2 (N1339, N1336, N1187);
xor XOR2 (N1340, N1330, N689);
buf BUF1 (N1341, N1333);
nor NOR3 (N1342, N1315, N568, N87);
or OR3 (N1343, N1335, N1311, N381);
or OR4 (N1344, N1327, N258, N345, N178);
buf BUF1 (N1345, N1344);
nor NOR4 (N1346, N1341, N1148, N225, N497);
nor NOR2 (N1347, N1331, N541);
xor XOR2 (N1348, N1328, N709);
or OR4 (N1349, N1346, N408, N1244, N579);
or OR4 (N1350, N1343, N439, N743, N958);
not NOT1 (N1351, N1345);
nor NOR4 (N1352, N1348, N177, N392, N477);
not NOT1 (N1353, N1351);
nand NAND2 (N1354, N1339, N681);
or OR3 (N1355, N1349, N521, N819);
and AND2 (N1356, N1353, N208);
nand NAND2 (N1357, N1350, N393);
and AND2 (N1358, N1337, N22);
nor NOR2 (N1359, N1352, N78);
not NOT1 (N1360, N1355);
and AND3 (N1361, N1359, N1312, N1074);
and AND3 (N1362, N1361, N1198, N1185);
nor NOR3 (N1363, N1340, N483, N187);
and AND2 (N1364, N1358, N576);
nor NOR2 (N1365, N1342, N404);
or OR4 (N1366, N1360, N1001, N1052, N1236);
nor NOR3 (N1367, N1347, N297, N1127);
or OR2 (N1368, N1366, N1104);
nand NAND2 (N1369, N1338, N1183);
buf BUF1 (N1370, N1364);
buf BUF1 (N1371, N1367);
and AND2 (N1372, N1354, N1168);
nand NAND2 (N1373, N1356, N687);
buf BUF1 (N1374, N1371);
buf BUF1 (N1375, N1372);
nor NOR3 (N1376, N1368, N745, N410);
nor NOR4 (N1377, N1376, N544, N1017, N94);
not NOT1 (N1378, N1363);
and AND3 (N1379, N1375, N522, N596);
buf BUF1 (N1380, N1369);
nor NOR4 (N1381, N1379, N70, N877, N799);
nor NOR4 (N1382, N1381, N1093, N995, N1365);
buf BUF1 (N1383, N142);
buf BUF1 (N1384, N1380);
or OR2 (N1385, N1382, N510);
nor NOR3 (N1386, N1385, N30, N1299);
buf BUF1 (N1387, N1384);
not NOT1 (N1388, N1362);
buf BUF1 (N1389, N1383);
or OR2 (N1390, N1374, N737);
buf BUF1 (N1391, N1388);
nand NAND2 (N1392, N1386, N1112);
buf BUF1 (N1393, N1389);
not NOT1 (N1394, N1378);
and AND4 (N1395, N1390, N628, N810, N1045);
not NOT1 (N1396, N1373);
buf BUF1 (N1397, N1391);
nor NOR3 (N1398, N1395, N1029, N860);
buf BUF1 (N1399, N1396);
nor NOR4 (N1400, N1377, N1247, N1290, N930);
nand NAND4 (N1401, N1398, N640, N79, N143);
xor XOR2 (N1402, N1392, N582);
nor NOR4 (N1403, N1397, N730, N1292, N1303);
buf BUF1 (N1404, N1399);
buf BUF1 (N1405, N1357);
or OR3 (N1406, N1393, N1241, N586);
and AND2 (N1407, N1370, N618);
nor NOR4 (N1408, N1400, N1323, N723, N278);
nor NOR3 (N1409, N1406, N518, N1028);
or OR2 (N1410, N1401, N1228);
buf BUF1 (N1411, N1410);
nand NAND4 (N1412, N1387, N891, N1337, N522);
nand NAND2 (N1413, N1409, N1275);
xor XOR2 (N1414, N1411, N555);
buf BUF1 (N1415, N1404);
and AND2 (N1416, N1413, N1094);
and AND2 (N1417, N1416, N318);
xor XOR2 (N1418, N1394, N926);
nor NOR3 (N1419, N1402, N109, N842);
nor NOR3 (N1420, N1403, N756, N398);
buf BUF1 (N1421, N1414);
or OR3 (N1422, N1407, N738, N474);
xor XOR2 (N1423, N1417, N907);
nand NAND3 (N1424, N1412, N457, N83);
and AND3 (N1425, N1408, N382, N597);
nand NAND4 (N1426, N1418, N1309, N1123, N979);
nand NAND3 (N1427, N1425, N74, N893);
nand NAND4 (N1428, N1420, N960, N997, N437);
nor NOR3 (N1429, N1421, N670, N1312);
buf BUF1 (N1430, N1423);
nand NAND4 (N1431, N1424, N1385, N58, N133);
and AND4 (N1432, N1415, N1048, N1362, N1215);
nor NOR2 (N1433, N1427, N1254);
xor XOR2 (N1434, N1429, N586);
xor XOR2 (N1435, N1433, N366);
xor XOR2 (N1436, N1426, N1326);
buf BUF1 (N1437, N1435);
or OR4 (N1438, N1419, N192, N98, N869);
nor NOR4 (N1439, N1428, N468, N460, N850);
and AND2 (N1440, N1439, N148);
and AND2 (N1441, N1431, N774);
and AND3 (N1442, N1405, N872, N210);
nor NOR4 (N1443, N1422, N936, N398, N466);
or OR3 (N1444, N1434, N919, N594);
buf BUF1 (N1445, N1442);
nor NOR2 (N1446, N1444, N296);
nor NOR2 (N1447, N1440, N640);
xor XOR2 (N1448, N1441, N1302);
xor XOR2 (N1449, N1446, N325);
buf BUF1 (N1450, N1430);
nor NOR2 (N1451, N1443, N945);
not NOT1 (N1452, N1450);
and AND3 (N1453, N1432, N929, N848);
nand NAND2 (N1454, N1445, N279);
or OR2 (N1455, N1454, N1165);
nor NOR3 (N1456, N1447, N281, N936);
or OR2 (N1457, N1449, N83);
nor NOR3 (N1458, N1456, N11, N866);
and AND3 (N1459, N1436, N1312, N493);
not NOT1 (N1460, N1459);
xor XOR2 (N1461, N1455, N689);
nor NOR3 (N1462, N1448, N390, N1141);
or OR4 (N1463, N1452, N840, N513, N869);
buf BUF1 (N1464, N1457);
nor NOR2 (N1465, N1458, N266);
or OR3 (N1466, N1438, N1443, N8);
and AND3 (N1467, N1462, N1414, N433);
or OR4 (N1468, N1463, N533, N1334, N818);
and AND4 (N1469, N1468, N1346, N828, N1325);
or OR4 (N1470, N1467, N255, N889, N1319);
buf BUF1 (N1471, N1464);
or OR2 (N1472, N1461, N715);
nor NOR2 (N1473, N1453, N309);
buf BUF1 (N1474, N1466);
nor NOR3 (N1475, N1474, N1296, N183);
not NOT1 (N1476, N1471);
xor XOR2 (N1477, N1465, N1095);
or OR4 (N1478, N1469, N412, N183, N683);
or OR2 (N1479, N1437, N705);
not NOT1 (N1480, N1478);
and AND2 (N1481, N1470, N1085);
buf BUF1 (N1482, N1480);
or OR2 (N1483, N1477, N739);
buf BUF1 (N1484, N1482);
or OR3 (N1485, N1476, N453, N1316);
buf BUF1 (N1486, N1460);
buf BUF1 (N1487, N1481);
or OR3 (N1488, N1485, N556, N1010);
not NOT1 (N1489, N1472);
or OR4 (N1490, N1479, N1207, N1089, N532);
xor XOR2 (N1491, N1489, N716);
xor XOR2 (N1492, N1475, N775);
nor NOR3 (N1493, N1490, N620, N648);
xor XOR2 (N1494, N1491, N103);
nor NOR2 (N1495, N1486, N1453);
or OR3 (N1496, N1495, N372, N965);
xor XOR2 (N1497, N1487, N368);
nor NOR3 (N1498, N1497, N1392, N940);
and AND3 (N1499, N1484, N1286, N1345);
nor NOR3 (N1500, N1494, N1059, N683);
not NOT1 (N1501, N1496);
or OR4 (N1502, N1492, N1377, N1308, N533);
and AND4 (N1503, N1498, N598, N759, N631);
not NOT1 (N1504, N1501);
nand NAND2 (N1505, N1488, N231);
and AND2 (N1506, N1500, N1391);
and AND3 (N1507, N1483, N1345, N1023);
buf BUF1 (N1508, N1506);
nand NAND2 (N1509, N1505, N1351);
nor NOR2 (N1510, N1451, N605);
and AND3 (N1511, N1508, N793, N368);
and AND4 (N1512, N1499, N305, N996, N1384);
not NOT1 (N1513, N1511);
xor XOR2 (N1514, N1510, N581);
xor XOR2 (N1515, N1503, N713);
nand NAND3 (N1516, N1493, N866, N743);
and AND4 (N1517, N1512, N1118, N194, N875);
xor XOR2 (N1518, N1514, N861);
xor XOR2 (N1519, N1516, N684);
and AND4 (N1520, N1502, N1003, N199, N566);
and AND4 (N1521, N1504, N645, N1082, N281);
xor XOR2 (N1522, N1507, N909);
not NOT1 (N1523, N1513);
or OR3 (N1524, N1515, N715, N1477);
nand NAND3 (N1525, N1473, N1436, N648);
not NOT1 (N1526, N1517);
buf BUF1 (N1527, N1518);
buf BUF1 (N1528, N1509);
buf BUF1 (N1529, N1521);
buf BUF1 (N1530, N1522);
nor NOR2 (N1531, N1529, N866);
not NOT1 (N1532, N1524);
buf BUF1 (N1533, N1520);
not NOT1 (N1534, N1528);
xor XOR2 (N1535, N1523, N302);
nand NAND3 (N1536, N1519, N809, N479);
nor NOR2 (N1537, N1533, N348);
or OR2 (N1538, N1537, N721);
and AND3 (N1539, N1532, N1190, N1222);
buf BUF1 (N1540, N1536);
buf BUF1 (N1541, N1525);
and AND4 (N1542, N1535, N940, N1513, N350);
buf BUF1 (N1543, N1541);
buf BUF1 (N1544, N1527);
and AND2 (N1545, N1542, N1386);
xor XOR2 (N1546, N1530, N793);
xor XOR2 (N1547, N1534, N1340);
not NOT1 (N1548, N1540);
or OR3 (N1549, N1526, N1052, N1338);
or OR3 (N1550, N1543, N126, N1128);
xor XOR2 (N1551, N1531, N75);
or OR2 (N1552, N1546, N138);
not NOT1 (N1553, N1549);
and AND3 (N1554, N1545, N1524, N811);
xor XOR2 (N1555, N1550, N1386);
nor NOR2 (N1556, N1554, N671);
not NOT1 (N1557, N1551);
buf BUF1 (N1558, N1553);
buf BUF1 (N1559, N1539);
xor XOR2 (N1560, N1556, N1117);
xor XOR2 (N1561, N1548, N554);
nand NAND2 (N1562, N1538, N1316);
or OR4 (N1563, N1557, N368, N898, N1206);
nand NAND3 (N1564, N1552, N965, N328);
nand NAND2 (N1565, N1563, N1386);
buf BUF1 (N1566, N1555);
and AND3 (N1567, N1564, N106, N797);
nor NOR4 (N1568, N1566, N1477, N405, N521);
nor NOR2 (N1569, N1568, N116);
buf BUF1 (N1570, N1569);
and AND3 (N1571, N1562, N892, N926);
xor XOR2 (N1572, N1571, N462);
or OR2 (N1573, N1544, N853);
nor NOR2 (N1574, N1560, N1398);
buf BUF1 (N1575, N1558);
or OR4 (N1576, N1567, N1222, N460, N1074);
and AND4 (N1577, N1570, N166, N108, N41);
and AND4 (N1578, N1575, N1550, N1518, N736);
or OR3 (N1579, N1565, N1260, N715);
buf BUF1 (N1580, N1576);
or OR2 (N1581, N1572, N724);
and AND4 (N1582, N1578, N1097, N878, N1580);
nand NAND2 (N1583, N673, N1189);
and AND2 (N1584, N1574, N804);
and AND2 (N1585, N1579, N615);
or OR3 (N1586, N1577, N1353, N147);
nor NOR4 (N1587, N1581, N253, N1454, N336);
nand NAND2 (N1588, N1585, N1197);
and AND3 (N1589, N1559, N445, N1548);
buf BUF1 (N1590, N1561);
nand NAND2 (N1591, N1573, N847);
nor NOR4 (N1592, N1591, N1023, N1202, N584);
or OR2 (N1593, N1589, N568);
not NOT1 (N1594, N1582);
not NOT1 (N1595, N1592);
nand NAND3 (N1596, N1583, N1453, N319);
xor XOR2 (N1597, N1586, N1103);
nand NAND2 (N1598, N1596, N1333);
or OR4 (N1599, N1597, N717, N676, N835);
nor NOR2 (N1600, N1588, N757);
buf BUF1 (N1601, N1600);
nor NOR4 (N1602, N1595, N810, N1492, N532);
xor XOR2 (N1603, N1601, N417);
nand NAND2 (N1604, N1590, N794);
nand NAND4 (N1605, N1602, N922, N701, N1516);
xor XOR2 (N1606, N1599, N1333);
nand NAND2 (N1607, N1584, N605);
not NOT1 (N1608, N1607);
buf BUF1 (N1609, N1604);
and AND2 (N1610, N1587, N416);
xor XOR2 (N1611, N1603, N1025);
nand NAND4 (N1612, N1598, N1300, N1368, N619);
or OR4 (N1613, N1612, N637, N210, N1027);
and AND4 (N1614, N1593, N1083, N1442, N120);
xor XOR2 (N1615, N1609, N575);
and AND3 (N1616, N1613, N170, N1525);
and AND3 (N1617, N1610, N1582, N287);
nor NOR2 (N1618, N1611, N800);
not NOT1 (N1619, N1618);
or OR2 (N1620, N1605, N623);
buf BUF1 (N1621, N1547);
not NOT1 (N1622, N1621);
and AND3 (N1623, N1619, N414, N1252);
not NOT1 (N1624, N1622);
buf BUF1 (N1625, N1616);
or OR2 (N1626, N1606, N748);
nor NOR4 (N1627, N1617, N696, N1518, N622);
and AND2 (N1628, N1627, N153);
not NOT1 (N1629, N1614);
nand NAND3 (N1630, N1623, N379, N566);
xor XOR2 (N1631, N1594, N1543);
and AND3 (N1632, N1615, N1196, N246);
not NOT1 (N1633, N1608);
nand NAND3 (N1634, N1620, N632, N832);
buf BUF1 (N1635, N1633);
and AND4 (N1636, N1628, N1138, N197, N944);
not NOT1 (N1637, N1635);
and AND2 (N1638, N1626, N448);
nor NOR2 (N1639, N1637, N59);
nand NAND3 (N1640, N1630, N300, N544);
and AND3 (N1641, N1636, N1405, N1559);
nand NAND4 (N1642, N1638, N118, N99, N1317);
buf BUF1 (N1643, N1642);
and AND3 (N1644, N1631, N456, N1477);
not NOT1 (N1645, N1639);
xor XOR2 (N1646, N1625, N1072);
xor XOR2 (N1647, N1643, N771);
and AND2 (N1648, N1629, N1083);
nor NOR2 (N1649, N1641, N1181);
not NOT1 (N1650, N1644);
and AND3 (N1651, N1624, N974, N1190);
nand NAND2 (N1652, N1634, N1416);
not NOT1 (N1653, N1651);
buf BUF1 (N1654, N1649);
nand NAND3 (N1655, N1640, N1366, N212);
buf BUF1 (N1656, N1655);
not NOT1 (N1657, N1656);
xor XOR2 (N1658, N1632, N856);
not NOT1 (N1659, N1646);
nor NOR2 (N1660, N1653, N299);
not NOT1 (N1661, N1647);
not NOT1 (N1662, N1645);
buf BUF1 (N1663, N1652);
not NOT1 (N1664, N1660);
nor NOR2 (N1665, N1658, N435);
nand NAND3 (N1666, N1650, N957, N412);
buf BUF1 (N1667, N1666);
xor XOR2 (N1668, N1667, N157);
nand NAND4 (N1669, N1662, N748, N767, N29);
nor NOR3 (N1670, N1659, N949, N900);
nor NOR4 (N1671, N1669, N506, N387, N1372);
and AND3 (N1672, N1657, N583, N599);
and AND3 (N1673, N1663, N57, N889);
or OR2 (N1674, N1665, N338);
or OR4 (N1675, N1671, N1070, N250, N792);
xor XOR2 (N1676, N1674, N125);
buf BUF1 (N1677, N1670);
xor XOR2 (N1678, N1675, N260);
xor XOR2 (N1679, N1676, N1061);
and AND2 (N1680, N1654, N1525);
buf BUF1 (N1681, N1672);
nor NOR4 (N1682, N1681, N893, N1573, N627);
xor XOR2 (N1683, N1664, N148);
buf BUF1 (N1684, N1661);
or OR2 (N1685, N1684, N701);
nand NAND3 (N1686, N1685, N1378, N1234);
not NOT1 (N1687, N1686);
nor NOR4 (N1688, N1673, N81, N519, N1553);
or OR3 (N1689, N1668, N1562, N472);
nor NOR4 (N1690, N1687, N29, N1490, N1340);
and AND2 (N1691, N1690, N676);
nor NOR4 (N1692, N1682, N1020, N919, N796);
and AND2 (N1693, N1648, N715);
or OR4 (N1694, N1688, N550, N621, N618);
not NOT1 (N1695, N1693);
nand NAND4 (N1696, N1695, N262, N1332, N805);
nand NAND4 (N1697, N1680, N820, N1040, N618);
nor NOR4 (N1698, N1678, N1528, N1016, N156);
and AND4 (N1699, N1698, N81, N1533, N871);
and AND4 (N1700, N1692, N581, N1429, N1371);
xor XOR2 (N1701, N1700, N111);
buf BUF1 (N1702, N1697);
xor XOR2 (N1703, N1694, N275);
or OR4 (N1704, N1699, N526, N542, N905);
not NOT1 (N1705, N1701);
or OR2 (N1706, N1679, N1632);
or OR4 (N1707, N1683, N612, N317, N203);
and AND4 (N1708, N1691, N1250, N1576, N578);
not NOT1 (N1709, N1702);
not NOT1 (N1710, N1703);
or OR3 (N1711, N1704, N489, N621);
nor NOR3 (N1712, N1711, N380, N1559);
and AND2 (N1713, N1707, N903);
nand NAND4 (N1714, N1710, N158, N774, N1048);
or OR3 (N1715, N1709, N290, N329);
not NOT1 (N1716, N1708);
nand NAND4 (N1717, N1713, N718, N1215, N973);
nor NOR3 (N1718, N1716, N1665, N169);
nor NOR3 (N1719, N1706, N1182, N591);
and AND4 (N1720, N1717, N1305, N258, N639);
nor NOR2 (N1721, N1705, N803);
buf BUF1 (N1722, N1696);
nand NAND4 (N1723, N1719, N1276, N813, N1656);
buf BUF1 (N1724, N1718);
nand NAND4 (N1725, N1714, N783, N1094, N490);
xor XOR2 (N1726, N1720, N1708);
nor NOR4 (N1727, N1723, N1304, N1169, N351);
not NOT1 (N1728, N1677);
nor NOR3 (N1729, N1728, N920, N611);
nor NOR2 (N1730, N1729, N987);
not NOT1 (N1731, N1725);
not NOT1 (N1732, N1726);
buf BUF1 (N1733, N1712);
or OR3 (N1734, N1715, N1084, N1698);
or OR2 (N1735, N1731, N826);
nor NOR4 (N1736, N1689, N596, N1426, N1521);
or OR2 (N1737, N1733, N1432);
nor NOR3 (N1738, N1734, N1381, N78);
nand NAND3 (N1739, N1721, N104, N1058);
and AND3 (N1740, N1736, N1343, N1384);
and AND2 (N1741, N1739, N300);
xor XOR2 (N1742, N1740, N849);
buf BUF1 (N1743, N1727);
nor NOR3 (N1744, N1724, N905, N33);
buf BUF1 (N1745, N1738);
nand NAND4 (N1746, N1722, N715, N1439, N1215);
or OR2 (N1747, N1742, N1169);
nor NOR3 (N1748, N1744, N430, N1060);
nand NAND2 (N1749, N1737, N1315);
buf BUF1 (N1750, N1743);
not NOT1 (N1751, N1741);
xor XOR2 (N1752, N1730, N1066);
or OR2 (N1753, N1748, N1731);
xor XOR2 (N1754, N1732, N1674);
xor XOR2 (N1755, N1745, N506);
not NOT1 (N1756, N1735);
buf BUF1 (N1757, N1756);
not NOT1 (N1758, N1751);
nand NAND4 (N1759, N1750, N1370, N115, N376);
nand NAND3 (N1760, N1755, N627, N594);
or OR2 (N1761, N1757, N1091);
nand NAND4 (N1762, N1759, N339, N1424, N1394);
nand NAND4 (N1763, N1754, N976, N805, N1585);
nand NAND3 (N1764, N1752, N1671, N1467);
xor XOR2 (N1765, N1749, N1453);
nor NOR3 (N1766, N1746, N708, N1366);
buf BUF1 (N1767, N1762);
not NOT1 (N1768, N1753);
and AND3 (N1769, N1768, N1400, N1020);
or OR4 (N1770, N1763, N1545, N737, N1528);
nor NOR4 (N1771, N1767, N1638, N1764, N199);
and AND3 (N1772, N384, N1710, N385);
or OR4 (N1773, N1765, N553, N872, N1722);
not NOT1 (N1774, N1758);
and AND3 (N1775, N1747, N1430, N1202);
nand NAND3 (N1776, N1771, N36, N82);
nand NAND4 (N1777, N1773, N258, N578, N460);
nand NAND3 (N1778, N1776, N1268, N1456);
or OR2 (N1779, N1775, N1450);
and AND2 (N1780, N1769, N805);
not NOT1 (N1781, N1779);
buf BUF1 (N1782, N1780);
nor NOR3 (N1783, N1766, N1123, N922);
xor XOR2 (N1784, N1781, N1350);
and AND2 (N1785, N1761, N697);
xor XOR2 (N1786, N1783, N1764);
not NOT1 (N1787, N1770);
not NOT1 (N1788, N1760);
buf BUF1 (N1789, N1782);
not NOT1 (N1790, N1772);
buf BUF1 (N1791, N1777);
xor XOR2 (N1792, N1791, N1678);
and AND4 (N1793, N1790, N1719, N729, N1185);
not NOT1 (N1794, N1792);
buf BUF1 (N1795, N1789);
buf BUF1 (N1796, N1794);
or OR3 (N1797, N1785, N781, N1712);
or OR2 (N1798, N1796, N1212);
not NOT1 (N1799, N1784);
nor NOR2 (N1800, N1798, N1121);
and AND3 (N1801, N1799, N1610, N942);
or OR3 (N1802, N1800, N1499, N704);
nor NOR4 (N1803, N1793, N202, N1335, N1484);
buf BUF1 (N1804, N1801);
xor XOR2 (N1805, N1774, N1578);
nor NOR2 (N1806, N1797, N808);
not NOT1 (N1807, N1804);
or OR4 (N1808, N1806, N1753, N711, N220);
nor NOR2 (N1809, N1778, N993);
not NOT1 (N1810, N1805);
xor XOR2 (N1811, N1803, N1136);
not NOT1 (N1812, N1788);
nor NOR4 (N1813, N1812, N377, N242, N1539);
not NOT1 (N1814, N1810);
not NOT1 (N1815, N1787);
not NOT1 (N1816, N1814);
and AND3 (N1817, N1795, N1334, N1132);
buf BUF1 (N1818, N1815);
not NOT1 (N1819, N1816);
xor XOR2 (N1820, N1807, N1035);
nor NOR2 (N1821, N1786, N1669);
and AND4 (N1822, N1820, N753, N1133, N1127);
or OR4 (N1823, N1813, N379, N1340, N952);
not NOT1 (N1824, N1809);
xor XOR2 (N1825, N1823, N709);
or OR4 (N1826, N1825, N703, N1648, N229);
nand NAND4 (N1827, N1824, N1758, N33, N1058);
nand NAND2 (N1828, N1811, N1311);
nand NAND2 (N1829, N1817, N567);
not NOT1 (N1830, N1808);
buf BUF1 (N1831, N1828);
nand NAND2 (N1832, N1822, N28);
and AND2 (N1833, N1829, N1331);
nor NOR2 (N1834, N1818, N695);
and AND2 (N1835, N1827, N626);
nand NAND4 (N1836, N1821, N350, N762, N264);
xor XOR2 (N1837, N1830, N1789);
nand NAND4 (N1838, N1826, N1208, N1370, N547);
or OR2 (N1839, N1837, N340);
xor XOR2 (N1840, N1838, N1699);
or OR3 (N1841, N1802, N163, N1805);
or OR3 (N1842, N1836, N146, N448);
xor XOR2 (N1843, N1835, N1199);
not NOT1 (N1844, N1841);
buf BUF1 (N1845, N1833);
xor XOR2 (N1846, N1840, N522);
xor XOR2 (N1847, N1846, N279);
buf BUF1 (N1848, N1844);
buf BUF1 (N1849, N1831);
and AND4 (N1850, N1843, N510, N1456, N245);
or OR2 (N1851, N1848, N211);
xor XOR2 (N1852, N1832, N1555);
nand NAND2 (N1853, N1847, N199);
not NOT1 (N1854, N1853);
or OR3 (N1855, N1845, N642, N598);
or OR4 (N1856, N1850, N216, N1518, N528);
xor XOR2 (N1857, N1851, N1375);
or OR4 (N1858, N1842, N1218, N323, N1680);
nand NAND4 (N1859, N1855, N702, N879, N28);
or OR4 (N1860, N1849, N1746, N1283, N1558);
not NOT1 (N1861, N1819);
not NOT1 (N1862, N1861);
or OR4 (N1863, N1854, N1308, N251, N84);
buf BUF1 (N1864, N1863);
buf BUF1 (N1865, N1839);
xor XOR2 (N1866, N1864, N1253);
xor XOR2 (N1867, N1834, N716);
nand NAND4 (N1868, N1858, N1554, N1106, N153);
or OR2 (N1869, N1859, N1252);
buf BUF1 (N1870, N1862);
buf BUF1 (N1871, N1856);
buf BUF1 (N1872, N1865);
and AND4 (N1873, N1871, N1417, N1586, N286);
or OR2 (N1874, N1866, N1042);
buf BUF1 (N1875, N1873);
nand NAND4 (N1876, N1857, N1011, N1658, N1595);
or OR2 (N1877, N1875, N983);
not NOT1 (N1878, N1876);
not NOT1 (N1879, N1852);
nand NAND4 (N1880, N1867, N355, N316, N1577);
or OR4 (N1881, N1879, N1277, N1083, N203);
xor XOR2 (N1882, N1868, N844);
nand NAND3 (N1883, N1880, N1107, N1005);
buf BUF1 (N1884, N1870);
xor XOR2 (N1885, N1883, N841);
xor XOR2 (N1886, N1877, N162);
nand NAND3 (N1887, N1884, N756, N1826);
not NOT1 (N1888, N1886);
or OR2 (N1889, N1887, N1174);
nand NAND3 (N1890, N1882, N759, N837);
and AND3 (N1891, N1881, N102, N84);
nor NOR4 (N1892, N1860, N840, N385, N1064);
buf BUF1 (N1893, N1874);
or OR3 (N1894, N1878, N214, N151);
nand NAND2 (N1895, N1892, N682);
nor NOR4 (N1896, N1885, N1038, N1637, N829);
or OR4 (N1897, N1896, N995, N535, N44);
and AND2 (N1898, N1891, N1413);
buf BUF1 (N1899, N1895);
and AND2 (N1900, N1897, N1393);
xor XOR2 (N1901, N1869, N248);
and AND3 (N1902, N1893, N1556, N202);
buf BUF1 (N1903, N1888);
buf BUF1 (N1904, N1894);
xor XOR2 (N1905, N1872, N997);
not NOT1 (N1906, N1900);
nand NAND3 (N1907, N1904, N575, N216);
and AND4 (N1908, N1903, N1867, N1750, N1583);
nor NOR4 (N1909, N1908, N1240, N1160, N1758);
nor NOR3 (N1910, N1906, N279, N1290);
nand NAND4 (N1911, N1910, N898, N1292, N1269);
buf BUF1 (N1912, N1898);
xor XOR2 (N1913, N1899, N958);
nand NAND2 (N1914, N1890, N571);
or OR2 (N1915, N1909, N498);
or OR3 (N1916, N1915, N278, N830);
or OR2 (N1917, N1912, N1812);
nand NAND3 (N1918, N1911, N954, N772);
not NOT1 (N1919, N1905);
xor XOR2 (N1920, N1901, N1487);
xor XOR2 (N1921, N1907, N36);
nor NOR2 (N1922, N1918, N463);
xor XOR2 (N1923, N1916, N811);
or OR2 (N1924, N1921, N963);
nor NOR2 (N1925, N1917, N1369);
or OR3 (N1926, N1914, N473, N705);
xor XOR2 (N1927, N1925, N1659);
not NOT1 (N1928, N1919);
xor XOR2 (N1929, N1920, N228);
nand NAND4 (N1930, N1927, N1722, N552, N1629);
nor NOR2 (N1931, N1923, N908);
xor XOR2 (N1932, N1929, N64);
nand NAND4 (N1933, N1924, N1001, N1181, N1485);
buf BUF1 (N1934, N1889);
not NOT1 (N1935, N1922);
not NOT1 (N1936, N1913);
not NOT1 (N1937, N1936);
nor NOR3 (N1938, N1935, N503, N840);
buf BUF1 (N1939, N1938);
xor XOR2 (N1940, N1930, N1666);
xor XOR2 (N1941, N1926, N368);
buf BUF1 (N1942, N1932);
buf BUF1 (N1943, N1928);
nand NAND2 (N1944, N1940, N33);
or OR3 (N1945, N1931, N262, N108);
or OR4 (N1946, N1939, N682, N309, N1614);
and AND4 (N1947, N1946, N353, N5, N461);
nand NAND2 (N1948, N1937, N687);
or OR3 (N1949, N1948, N488, N133);
nor NOR4 (N1950, N1902, N1493, N411, N1825);
and AND2 (N1951, N1944, N117);
buf BUF1 (N1952, N1942);
xor XOR2 (N1953, N1941, N1321);
nand NAND2 (N1954, N1951, N1444);
or OR2 (N1955, N1953, N1954);
or OR3 (N1956, N448, N524, N1580);
xor XOR2 (N1957, N1956, N1485);
buf BUF1 (N1958, N1955);
nand NAND4 (N1959, N1949, N1127, N762, N1879);
buf BUF1 (N1960, N1933);
buf BUF1 (N1961, N1947);
and AND3 (N1962, N1960, N890, N1009);
nor NOR2 (N1963, N1952, N736);
or OR2 (N1964, N1943, N681);
not NOT1 (N1965, N1963);
not NOT1 (N1966, N1957);
xor XOR2 (N1967, N1950, N817);
nand NAND2 (N1968, N1934, N212);
and AND2 (N1969, N1968, N1633);
nand NAND3 (N1970, N1962, N1486, N438);
xor XOR2 (N1971, N1958, N109);
nor NOR2 (N1972, N1967, N579);
buf BUF1 (N1973, N1945);
nand NAND3 (N1974, N1965, N796, N703);
nor NOR3 (N1975, N1959, N265, N245);
nand NAND3 (N1976, N1969, N571, N282);
not NOT1 (N1977, N1970);
xor XOR2 (N1978, N1974, N647);
or OR2 (N1979, N1978, N1474);
not NOT1 (N1980, N1977);
xor XOR2 (N1981, N1980, N1575);
and AND3 (N1982, N1976, N403, N714);
buf BUF1 (N1983, N1971);
xor XOR2 (N1984, N1973, N1190);
nand NAND3 (N1985, N1982, N1763, N1819);
or OR4 (N1986, N1961, N1072, N780, N1488);
not NOT1 (N1987, N1983);
and AND2 (N1988, N1985, N874);
not NOT1 (N1989, N1987);
xor XOR2 (N1990, N1988, N173);
and AND3 (N1991, N1981, N1820, N1018);
not NOT1 (N1992, N1966);
and AND3 (N1993, N1972, N998, N1559);
nor NOR4 (N1994, N1964, N39, N109, N621);
not NOT1 (N1995, N1984);
nor NOR3 (N1996, N1989, N176, N860);
nand NAND4 (N1997, N1990, N1343, N305, N1042);
nand NAND2 (N1998, N1986, N1273);
buf BUF1 (N1999, N1979);
xor XOR2 (N2000, N1998, N777);
not NOT1 (N2001, N1991);
buf BUF1 (N2002, N1996);
or OR3 (N2003, N2001, N1813, N976);
buf BUF1 (N2004, N1997);
not NOT1 (N2005, N2004);
xor XOR2 (N2006, N1975, N876);
and AND3 (N2007, N2005, N168, N1942);
nor NOR4 (N2008, N1993, N894, N853, N46);
nor NOR2 (N2009, N2003, N1583);
buf BUF1 (N2010, N2002);
buf BUF1 (N2011, N2006);
buf BUF1 (N2012, N1999);
buf BUF1 (N2013, N1994);
or OR3 (N2014, N2007, N96, N702);
not NOT1 (N2015, N2014);
or OR3 (N2016, N2013, N511, N1529);
xor XOR2 (N2017, N2008, N1398);
nand NAND4 (N2018, N2011, N713, N316, N1817);
nand NAND4 (N2019, N1992, N663, N1664, N817);
buf BUF1 (N2020, N2012);
xor XOR2 (N2021, N2017, N1757);
xor XOR2 (N2022, N2020, N1656);
and AND4 (N2023, N2022, N533, N547, N1924);
buf BUF1 (N2024, N2021);
buf BUF1 (N2025, N2019);
nor NOR2 (N2026, N2010, N829);
nand NAND2 (N2027, N2025, N932);
nor NOR4 (N2028, N2026, N1192, N1463, N475);
buf BUF1 (N2029, N2015);
xor XOR2 (N2030, N2009, N1290);
and AND3 (N2031, N2029, N1806, N982);
not NOT1 (N2032, N2016);
nor NOR3 (N2033, N2031, N646, N960);
or OR4 (N2034, N2028, N1570, N1061, N905);
or OR3 (N2035, N1995, N1782, N253);
and AND2 (N2036, N2027, N1942);
nand NAND3 (N2037, N2033, N1023, N1492);
nand NAND2 (N2038, N2035, N317);
and AND3 (N2039, N2030, N889, N1722);
buf BUF1 (N2040, N2036);
or OR4 (N2041, N2000, N336, N1844, N1848);
nor NOR2 (N2042, N2034, N206);
nor NOR2 (N2043, N2042, N716);
nand NAND2 (N2044, N2023, N1830);
and AND4 (N2045, N2040, N1954, N1533, N58);
and AND4 (N2046, N2041, N1666, N1401, N1128);
nand NAND4 (N2047, N2037, N1566, N1752, N1734);
xor XOR2 (N2048, N2045, N23);
xor XOR2 (N2049, N2044, N1884);
not NOT1 (N2050, N2024);
buf BUF1 (N2051, N2047);
not NOT1 (N2052, N2038);
buf BUF1 (N2053, N2051);
nor NOR4 (N2054, N2052, N78, N1961, N892);
not NOT1 (N2055, N2043);
buf BUF1 (N2056, N2048);
xor XOR2 (N2057, N2055, N978);
nor NOR2 (N2058, N2032, N2034);
or OR4 (N2059, N2056, N611, N663, N189);
or OR3 (N2060, N2046, N112, N1718);
nand NAND4 (N2061, N2053, N1665, N761, N615);
or OR4 (N2062, N2054, N102, N922, N1004);
nor NOR3 (N2063, N2061, N1581, N123);
nor NOR4 (N2064, N2059, N2057, N847, N1804);
and AND4 (N2065, N1668, N1542, N1335, N1086);
not NOT1 (N2066, N2050);
nand NAND2 (N2067, N2063, N622);
xor XOR2 (N2068, N2058, N1999);
buf BUF1 (N2069, N2065);
buf BUF1 (N2070, N2060);
or OR2 (N2071, N2069, N899);
nand NAND2 (N2072, N2039, N184);
or OR2 (N2073, N2018, N1438);
xor XOR2 (N2074, N2068, N947);
buf BUF1 (N2075, N2073);
nand NAND4 (N2076, N2070, N1936, N737, N1100);
xor XOR2 (N2077, N2062, N1930);
nor NOR2 (N2078, N2076, N316);
or OR3 (N2079, N2078, N1163, N1462);
xor XOR2 (N2080, N2072, N1549);
not NOT1 (N2081, N2075);
or OR2 (N2082, N2064, N954);
xor XOR2 (N2083, N2077, N913);
buf BUF1 (N2084, N2083);
not NOT1 (N2085, N2049);
buf BUF1 (N2086, N2079);
and AND4 (N2087, N2067, N1832, N1067, N1845);
nor NOR3 (N2088, N2085, N1955, N278);
xor XOR2 (N2089, N2081, N1854);
xor XOR2 (N2090, N2087, N6);
nor NOR2 (N2091, N2088, N209);
nand NAND4 (N2092, N2089, N1475, N463, N1732);
buf BUF1 (N2093, N2092);
nor NOR4 (N2094, N2091, N1856, N1589, N1948);
or OR3 (N2095, N2080, N1289, N1859);
and AND4 (N2096, N2082, N713, N954, N145);
xor XOR2 (N2097, N2071, N1180);
nand NAND3 (N2098, N2095, N507, N1554);
xor XOR2 (N2099, N2090, N1594);
nor NOR3 (N2100, N2074, N1581, N1986);
xor XOR2 (N2101, N2098, N234);
nand NAND2 (N2102, N2086, N348);
xor XOR2 (N2103, N2094, N1154);
buf BUF1 (N2104, N2096);
not NOT1 (N2105, N2084);
not NOT1 (N2106, N2105);
buf BUF1 (N2107, N2066);
and AND3 (N2108, N2102, N584, N2021);
buf BUF1 (N2109, N2107);
xor XOR2 (N2110, N2100, N507);
and AND2 (N2111, N2101, N25);
not NOT1 (N2112, N2106);
not NOT1 (N2113, N2093);
nand NAND2 (N2114, N2099, N1409);
or OR2 (N2115, N2104, N458);
buf BUF1 (N2116, N2109);
xor XOR2 (N2117, N2112, N1550);
not NOT1 (N2118, N2110);
and AND4 (N2119, N2116, N1205, N1457, N1871);
nand NAND2 (N2120, N2111, N119);
nand NAND3 (N2121, N2115, N792, N382);
and AND2 (N2122, N2120, N1153);
and AND3 (N2123, N2097, N1446, N808);
xor XOR2 (N2124, N2114, N1402);
and AND4 (N2125, N2118, N172, N479, N438);
not NOT1 (N2126, N2119);
nor NOR4 (N2127, N2121, N1494, N1749, N608);
xor XOR2 (N2128, N2117, N120);
or OR4 (N2129, N2125, N577, N329, N626);
and AND4 (N2130, N2124, N1830, N1091, N433);
and AND3 (N2131, N2127, N1719, N1053);
nor NOR4 (N2132, N2123, N804, N1983, N891);
nand NAND3 (N2133, N2130, N103, N185);
and AND3 (N2134, N2113, N1371, N1125);
and AND3 (N2135, N2122, N729, N1516);
and AND3 (N2136, N2108, N252, N1772);
or OR2 (N2137, N2126, N914);
nor NOR4 (N2138, N2132, N1323, N707, N1296);
xor XOR2 (N2139, N2134, N1376);
or OR2 (N2140, N2135, N803);
not NOT1 (N2141, N2138);
nor NOR3 (N2142, N2103, N414, N1993);
xor XOR2 (N2143, N2129, N1416);
nor NOR4 (N2144, N2128, N1455, N1149, N1202);
buf BUF1 (N2145, N2139);
nor NOR3 (N2146, N2137, N1869, N1811);
buf BUF1 (N2147, N2131);
xor XOR2 (N2148, N2142, N1631);
buf BUF1 (N2149, N2148);
xor XOR2 (N2150, N2145, N1292);
and AND2 (N2151, N2144, N965);
xor XOR2 (N2152, N2151, N1435);
xor XOR2 (N2153, N2152, N976);
not NOT1 (N2154, N2133);
xor XOR2 (N2155, N2154, N166);
and AND2 (N2156, N2149, N728);
and AND3 (N2157, N2136, N814, N253);
not NOT1 (N2158, N2147);
or OR2 (N2159, N2157, N1471);
xor XOR2 (N2160, N2146, N1889);
or OR3 (N2161, N2159, N1406, N1833);
not NOT1 (N2162, N2155);
nand NAND4 (N2163, N2140, N1657, N1431, N501);
and AND3 (N2164, N2161, N2055, N1204);
not NOT1 (N2165, N2164);
and AND3 (N2166, N2156, N2068, N1436);
buf BUF1 (N2167, N2141);
nand NAND2 (N2168, N2162, N1905);
and AND4 (N2169, N2150, N76, N1487, N2144);
nand NAND3 (N2170, N2158, N1583, N1137);
nor NOR3 (N2171, N2166, N180, N1299);
xor XOR2 (N2172, N2165, N1555);
nor NOR2 (N2173, N2153, N1124);
xor XOR2 (N2174, N2169, N1632);
nor NOR4 (N2175, N2170, N2093, N2094, N2164);
nor NOR3 (N2176, N2168, N1570, N1472);
buf BUF1 (N2177, N2167);
or OR2 (N2178, N2175, N952);
and AND3 (N2179, N2176, N1072, N1843);
nand NAND2 (N2180, N2163, N1944);
not NOT1 (N2181, N2174);
or OR4 (N2182, N2172, N2019, N486, N530);
xor XOR2 (N2183, N2179, N1598);
or OR2 (N2184, N2173, N1224);
xor XOR2 (N2185, N2182, N1152);
not NOT1 (N2186, N2177);
xor XOR2 (N2187, N2186, N307);
buf BUF1 (N2188, N2180);
nor NOR2 (N2189, N2188, N2118);
buf BUF1 (N2190, N2171);
and AND3 (N2191, N2189, N452, N689);
not NOT1 (N2192, N2183);
and AND2 (N2193, N2184, N858);
or OR2 (N2194, N2193, N1043);
buf BUF1 (N2195, N2194);
nand NAND2 (N2196, N2181, N1738);
nor NOR2 (N2197, N2178, N1659);
and AND4 (N2198, N2185, N330, N1385, N1450);
or OR2 (N2199, N2197, N2180);
xor XOR2 (N2200, N2190, N1931);
not NOT1 (N2201, N2195);
nand NAND2 (N2202, N2200, N1122);
or OR2 (N2203, N2187, N499);
or OR4 (N2204, N2203, N209, N1821, N1739);
not NOT1 (N2205, N2198);
nor NOR3 (N2206, N2201, N1023, N1680);
nand NAND4 (N2207, N2202, N1594, N1385, N840);
nand NAND3 (N2208, N2206, N297, N1631);
or OR3 (N2209, N2191, N1955, N1412);
nand NAND4 (N2210, N2207, N1823, N2008, N2020);
nor NOR3 (N2211, N2208, N1917, N463);
nand NAND4 (N2212, N2160, N658, N980, N1287);
buf BUF1 (N2213, N2204);
nand NAND2 (N2214, N2205, N1834);
nor NOR4 (N2215, N2196, N1453, N1389, N1434);
xor XOR2 (N2216, N2214, N1201);
xor XOR2 (N2217, N2213, N810);
or OR4 (N2218, N2209, N965, N1375, N470);
nor NOR4 (N2219, N2212, N1487, N1800, N334);
not NOT1 (N2220, N2217);
or OR2 (N2221, N2219, N1944);
nor NOR2 (N2222, N2143, N2204);
nand NAND3 (N2223, N2222, N385, N2095);
nand NAND2 (N2224, N2218, N1937);
nand NAND3 (N2225, N2192, N2080, N1796);
nand NAND4 (N2226, N2210, N2103, N619, N1657);
xor XOR2 (N2227, N2211, N331);
or OR2 (N2228, N2227, N327);
or OR2 (N2229, N2223, N1812);
nor NOR2 (N2230, N2220, N259);
xor XOR2 (N2231, N2226, N1383);
nor NOR2 (N2232, N2199, N547);
and AND3 (N2233, N2229, N1575, N1785);
nand NAND3 (N2234, N2225, N1515, N1835);
nand NAND4 (N2235, N2228, N1341, N782, N2190);
nand NAND4 (N2236, N2221, N755, N593, N333);
nor NOR4 (N2237, N2215, N1861, N744, N588);
xor XOR2 (N2238, N2233, N1872);
nand NAND2 (N2239, N2237, N548);
buf BUF1 (N2240, N2238);
and AND3 (N2241, N2236, N1359, N549);
nand NAND3 (N2242, N2234, N2115, N2129);
or OR3 (N2243, N2231, N1426, N1201);
not NOT1 (N2244, N2242);
nor NOR3 (N2245, N2244, N1465, N1880);
or OR3 (N2246, N2224, N1173, N1121);
or OR2 (N2247, N2235, N2136);
buf BUF1 (N2248, N2230);
xor XOR2 (N2249, N2239, N1977);
and AND3 (N2250, N2232, N863, N1096);
nor NOR2 (N2251, N2250, N1864);
xor XOR2 (N2252, N2243, N2079);
buf BUF1 (N2253, N2241);
xor XOR2 (N2254, N2252, N542);
nand NAND3 (N2255, N2245, N547, N306);
or OR2 (N2256, N2255, N5);
or OR4 (N2257, N2216, N1261, N1999, N1644);
not NOT1 (N2258, N2240);
nor NOR3 (N2259, N2248, N1231, N2106);
and AND4 (N2260, N2249, N539, N1909, N731);
nand NAND3 (N2261, N2251, N871, N1304);
or OR2 (N2262, N2260, N1402);
xor XOR2 (N2263, N2258, N790);
nor NOR4 (N2264, N2246, N388, N196, N691);
nor NOR4 (N2265, N2259, N751, N1251, N1797);
or OR2 (N2266, N2256, N1457);
nand NAND3 (N2267, N2257, N1679, N1442);
nand NAND2 (N2268, N2264, N1125);
nor NOR4 (N2269, N2253, N1714, N429, N1599);
nand NAND4 (N2270, N2247, N74, N363, N1473);
not NOT1 (N2271, N2266);
or OR4 (N2272, N2269, N1591, N2168, N4);
nand NAND4 (N2273, N2263, N861, N834, N132);
xor XOR2 (N2274, N2270, N19);
not NOT1 (N2275, N2267);
xor XOR2 (N2276, N2262, N921);
or OR2 (N2277, N2276, N415);
nor NOR4 (N2278, N2274, N1607, N1253, N1);
not NOT1 (N2279, N2261);
nand NAND3 (N2280, N2268, N848, N2222);
or OR4 (N2281, N2278, N1687, N1857, N59);
or OR2 (N2282, N2277, N1267);
and AND3 (N2283, N2281, N2018, N1043);
buf BUF1 (N2284, N2283);
buf BUF1 (N2285, N2280);
buf BUF1 (N2286, N2272);
not NOT1 (N2287, N2275);
xor XOR2 (N2288, N2286, N1797);
buf BUF1 (N2289, N2265);
nor NOR3 (N2290, N2285, N1178, N245);
nor NOR4 (N2291, N2287, N628, N797, N1038);
nor NOR4 (N2292, N2290, N1745, N640, N2135);
xor XOR2 (N2293, N2273, N1829);
nand NAND2 (N2294, N2271, N1953);
nor NOR2 (N2295, N2254, N1502);
and AND4 (N2296, N2289, N259, N2073, N1206);
xor XOR2 (N2297, N2284, N1236);
nor NOR2 (N2298, N2296, N1802);
buf BUF1 (N2299, N2298);
xor XOR2 (N2300, N2293, N339);
xor XOR2 (N2301, N2299, N2044);
nand NAND4 (N2302, N2294, N829, N837, N889);
or OR2 (N2303, N2292, N736);
nor NOR4 (N2304, N2303, N1814, N1525, N1418);
nor NOR2 (N2305, N2300, N2096);
and AND2 (N2306, N2302, N1169);
and AND2 (N2307, N2288, N44);
or OR3 (N2308, N2291, N1594, N959);
nor NOR3 (N2309, N2282, N342, N1398);
not NOT1 (N2310, N2305);
nand NAND3 (N2311, N2310, N1357, N53);
nand NAND3 (N2312, N2301, N502, N687);
nand NAND3 (N2313, N2279, N1863, N2013);
nor NOR4 (N2314, N2309, N254, N2291, N14);
xor XOR2 (N2315, N2295, N1126);
buf BUF1 (N2316, N2311);
xor XOR2 (N2317, N2307, N923);
not NOT1 (N2318, N2312);
not NOT1 (N2319, N2314);
and AND3 (N2320, N2306, N405, N1012);
nand NAND3 (N2321, N2318, N2061, N277);
nand NAND3 (N2322, N2316, N150, N816);
and AND4 (N2323, N2308, N490, N1850, N1311);
and AND2 (N2324, N2304, N1142);
nand NAND3 (N2325, N2313, N1133, N2219);
and AND2 (N2326, N2321, N297);
nand NAND2 (N2327, N2320, N1246);
xor XOR2 (N2328, N2325, N2146);
or OR4 (N2329, N2297, N1571, N1101, N108);
xor XOR2 (N2330, N2317, N1115);
not NOT1 (N2331, N2328);
or OR2 (N2332, N2323, N1276);
xor XOR2 (N2333, N2332, N351);
xor XOR2 (N2334, N2319, N1197);
and AND4 (N2335, N2322, N332, N188, N1652);
not NOT1 (N2336, N2334);
xor XOR2 (N2337, N2315, N1349);
or OR2 (N2338, N2333, N691);
not NOT1 (N2339, N2326);
xor XOR2 (N2340, N2331, N1551);
and AND4 (N2341, N2330, N522, N486, N501);
nor NOR3 (N2342, N2327, N1480, N569);
or OR2 (N2343, N2339, N1815);
and AND3 (N2344, N2324, N1372, N1545);
nor NOR2 (N2345, N2341, N2181);
and AND4 (N2346, N2340, N2088, N1335, N1927);
and AND2 (N2347, N2337, N963);
xor XOR2 (N2348, N2338, N257);
buf BUF1 (N2349, N2342);
xor XOR2 (N2350, N2346, N481);
buf BUF1 (N2351, N2349);
or OR2 (N2352, N2351, N841);
buf BUF1 (N2353, N2329);
nor NOR3 (N2354, N2348, N820, N2092);
nand NAND3 (N2355, N2335, N585, N564);
or OR2 (N2356, N2352, N1462);
nor NOR2 (N2357, N2353, N1270);
nand NAND2 (N2358, N2350, N727);
not NOT1 (N2359, N2358);
buf BUF1 (N2360, N2344);
buf BUF1 (N2361, N2354);
nand NAND3 (N2362, N2345, N1913, N1236);
buf BUF1 (N2363, N2343);
nand NAND4 (N2364, N2336, N1410, N616, N567);
nand NAND3 (N2365, N2357, N1633, N1707);
or OR4 (N2366, N2364, N1095, N782, N384);
nor NOR4 (N2367, N2360, N823, N1549, N1023);
not NOT1 (N2368, N2355);
nor NOR3 (N2369, N2359, N337, N1250);
xor XOR2 (N2370, N2363, N85);
xor XOR2 (N2371, N2347, N207);
buf BUF1 (N2372, N2361);
nor NOR4 (N2373, N2372, N768, N1218, N583);
xor XOR2 (N2374, N2366, N946);
buf BUF1 (N2375, N2362);
not NOT1 (N2376, N2371);
nand NAND2 (N2377, N2374, N2146);
xor XOR2 (N2378, N2365, N1568);
and AND2 (N2379, N2368, N151);
and AND3 (N2380, N2375, N1002, N2331);
nand NAND3 (N2381, N2376, N1432, N1828);
and AND3 (N2382, N2373, N14, N1495);
and AND2 (N2383, N2367, N2170);
and AND3 (N2384, N2383, N291, N999);
not NOT1 (N2385, N2382);
nand NAND2 (N2386, N2380, N2267);
nor NOR3 (N2387, N2369, N1062, N889);
and AND3 (N2388, N2387, N726, N1755);
or OR4 (N2389, N2388, N110, N1860, N2097);
nor NOR2 (N2390, N2384, N1592);
or OR4 (N2391, N2381, N1282, N1757, N568);
or OR3 (N2392, N2385, N1576, N1929);
nand NAND3 (N2393, N2389, N2085, N447);
or OR4 (N2394, N2379, N715, N1521, N689);
buf BUF1 (N2395, N2377);
or OR4 (N2396, N2356, N681, N213, N1627);
not NOT1 (N2397, N2392);
nand NAND2 (N2398, N2396, N531);
nor NOR4 (N2399, N2391, N848, N696, N658);
or OR4 (N2400, N2386, N608, N808, N1224);
not NOT1 (N2401, N2395);
xor XOR2 (N2402, N2398, N2315);
and AND2 (N2403, N2370, N1);
and AND4 (N2404, N2399, N2393, N538, N1017);
nor NOR2 (N2405, N666, N831);
xor XOR2 (N2406, N2403, N1920);
buf BUF1 (N2407, N2406);
nor NOR3 (N2408, N2390, N824, N1036);
nor NOR2 (N2409, N2401, N391);
not NOT1 (N2410, N2378);
not NOT1 (N2411, N2394);
buf BUF1 (N2412, N2410);
or OR4 (N2413, N2400, N1939, N123, N1123);
or OR2 (N2414, N2411, N380);
nand NAND2 (N2415, N2413, N13);
nand NAND2 (N2416, N2404, N490);
buf BUF1 (N2417, N2412);
nand NAND2 (N2418, N2416, N1414);
xor XOR2 (N2419, N2415, N728);
buf BUF1 (N2420, N2405);
xor XOR2 (N2421, N2402, N1052);
and AND3 (N2422, N2409, N802, N65);
nand NAND4 (N2423, N2419, N440, N81, N1891);
nor NOR4 (N2424, N2423, N878, N136, N1867);
and AND2 (N2425, N2407, N1827);
xor XOR2 (N2426, N2422, N1321);
nor NOR3 (N2427, N2397, N1088, N1899);
nand NAND4 (N2428, N2427, N1305, N1393, N931);
buf BUF1 (N2429, N2428);
nand NAND3 (N2430, N2426, N2096, N1440);
nor NOR3 (N2431, N2414, N1798, N1090);
xor XOR2 (N2432, N2417, N898);
buf BUF1 (N2433, N2408);
or OR4 (N2434, N2421, N596, N1129, N431);
xor XOR2 (N2435, N2424, N383);
xor XOR2 (N2436, N2429, N1502);
xor XOR2 (N2437, N2430, N616);
nor NOR2 (N2438, N2433, N1898);
not NOT1 (N2439, N2435);
buf BUF1 (N2440, N2432);
not NOT1 (N2441, N2438);
and AND2 (N2442, N2418, N543);
or OR3 (N2443, N2440, N186, N1446);
or OR2 (N2444, N2434, N383);
nand NAND2 (N2445, N2431, N2292);
xor XOR2 (N2446, N2444, N1395);
not NOT1 (N2447, N2439);
buf BUF1 (N2448, N2437);
buf BUF1 (N2449, N2446);
xor XOR2 (N2450, N2436, N2098);
xor XOR2 (N2451, N2442, N2102);
and AND3 (N2452, N2420, N1502, N2010);
xor XOR2 (N2453, N2447, N1460);
nand NAND4 (N2454, N2449, N1806, N1963, N778);
not NOT1 (N2455, N2453);
or OR2 (N2456, N2441, N2326);
buf BUF1 (N2457, N2450);
buf BUF1 (N2458, N2454);
nand NAND3 (N2459, N2445, N561, N783);
nand NAND2 (N2460, N2452, N532);
nor NOR3 (N2461, N2425, N2162, N1562);
and AND3 (N2462, N2443, N1460, N1237);
buf BUF1 (N2463, N2459);
not NOT1 (N2464, N2460);
nor NOR2 (N2465, N2458, N305);
buf BUF1 (N2466, N2464);
xor XOR2 (N2467, N2466, N448);
xor XOR2 (N2468, N2463, N54);
and AND2 (N2469, N2455, N1775);
and AND3 (N2470, N2448, N1999, N1024);
buf BUF1 (N2471, N2467);
nor NOR3 (N2472, N2451, N737, N1353);
nor NOR4 (N2473, N2468, N1451, N2336, N466);
xor XOR2 (N2474, N2461, N2156);
buf BUF1 (N2475, N2473);
not NOT1 (N2476, N2475);
nand NAND2 (N2477, N2456, N1320);
not NOT1 (N2478, N2472);
xor XOR2 (N2479, N2465, N654);
not NOT1 (N2480, N2471);
buf BUF1 (N2481, N2479);
xor XOR2 (N2482, N2477, N343);
not NOT1 (N2483, N2482);
or OR3 (N2484, N2470, N1903, N2411);
and AND3 (N2485, N2457, N563, N602);
and AND3 (N2486, N2483, N569, N2235);
and AND4 (N2487, N2486, N1677, N1591, N2365);
and AND4 (N2488, N2469, N1471, N923, N688);
buf BUF1 (N2489, N2474);
buf BUF1 (N2490, N2478);
not NOT1 (N2491, N2462);
nand NAND4 (N2492, N2491, N1442, N1060, N1242);
nor NOR3 (N2493, N2480, N1434, N497);
or OR2 (N2494, N2488, N1534);
and AND2 (N2495, N2485, N635);
and AND2 (N2496, N2476, N790);
buf BUF1 (N2497, N2489);
not NOT1 (N2498, N2487);
not NOT1 (N2499, N2490);
not NOT1 (N2500, N2493);
nand NAND3 (N2501, N2498, N1828, N1679);
nand NAND3 (N2502, N2492, N382, N2386);
and AND2 (N2503, N2502, N1473);
and AND4 (N2504, N2497, N2425, N1058, N165);
or OR3 (N2505, N2501, N2135, N1323);
xor XOR2 (N2506, N2484, N2109);
or OR2 (N2507, N2499, N1441);
and AND3 (N2508, N2494, N2371, N1338);
and AND2 (N2509, N2500, N1288);
xor XOR2 (N2510, N2495, N1974);
nor NOR2 (N2511, N2510, N2177);
nor NOR2 (N2512, N2506, N1550);
nand NAND2 (N2513, N2496, N1020);
buf BUF1 (N2514, N2511);
endmodule