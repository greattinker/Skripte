// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13;

output N103,N112,N92,N95,N111,N99,N110,N108,N106,N113;

xor XOR2 (N14, N13, N5);
nand NAND4 (N15, N6, N5, N8, N6);
buf BUF1 (N16, N6);
nand NAND3 (N17, N9, N11, N8);
or OR2 (N18, N14, N16);
buf BUF1 (N19, N7);
xor XOR2 (N20, N3, N4);
or OR3 (N21, N11, N10, N3);
or OR3 (N22, N16, N15, N7);
xor XOR2 (N23, N1, N4);
and AND2 (N24, N22, N19);
or OR2 (N25, N10, N6);
buf BUF1 (N26, N1);
nor NOR2 (N27, N7, N13);
nand NAND3 (N28, N4, N22, N24);
buf BUF1 (N29, N23);
and AND3 (N30, N6, N13, N1);
or OR4 (N31, N17, N29, N20, N10);
nand NAND2 (N32, N29, N18);
and AND4 (N33, N15, N13, N16, N24);
buf BUF1 (N34, N10);
buf BUF1 (N35, N34);
nor NOR3 (N36, N30, N34, N4);
buf BUF1 (N37, N33);
and AND3 (N38, N36, N29, N13);
buf BUF1 (N39, N37);
and AND3 (N40, N35, N23, N31);
buf BUF1 (N41, N23);
or OR3 (N42, N40, N35, N27);
nand NAND4 (N43, N26, N37, N32, N24);
nand NAND3 (N44, N17, N25, N35);
nor NOR4 (N45, N39, N26, N29, N3);
nand NAND4 (N46, N44, N17, N37, N34);
and AND3 (N47, N26, N7, N29);
not NOT1 (N48, N21);
nand NAND2 (N49, N16, N8);
nor NOR3 (N50, N38, N12, N48);
buf BUF1 (N51, N12);
buf BUF1 (N52, N28);
or OR4 (N53, N41, N13, N32, N40);
xor XOR2 (N54, N49, N32);
xor XOR2 (N55, N53, N28);
nor NOR4 (N56, N52, N12, N20, N55);
buf BUF1 (N57, N33);
and AND3 (N58, N51, N26, N20);
and AND4 (N59, N43, N54, N47, N55);
and AND4 (N60, N55, N46, N40, N4);
and AND3 (N61, N13, N14, N40);
and AND2 (N62, N41, N8);
xor XOR2 (N63, N56, N7);
nand NAND4 (N64, N61, N58, N13, N27);
nor NOR2 (N65, N40, N48);
not NOT1 (N66, N63);
xor XOR2 (N67, N66, N44);
nand NAND4 (N68, N67, N16, N21, N47);
xor XOR2 (N69, N68, N59);
nand NAND3 (N70, N39, N29, N60);
or OR3 (N71, N2, N67, N63);
nand NAND2 (N72, N45, N52);
buf BUF1 (N73, N70);
or OR2 (N74, N42, N50);
not NOT1 (N75, N12);
or OR2 (N76, N65, N10);
nand NAND4 (N77, N74, N25, N49, N58);
buf BUF1 (N78, N76);
nor NOR3 (N79, N62, N61, N22);
nand NAND2 (N80, N57, N19);
and AND3 (N81, N79, N2, N32);
nor NOR4 (N82, N73, N35, N24, N26);
nor NOR4 (N83, N80, N10, N13, N22);
xor XOR2 (N84, N81, N57);
nor NOR4 (N85, N72, N15, N36, N50);
nand NAND2 (N86, N77, N66);
nand NAND4 (N87, N83, N31, N72, N69);
nor NOR3 (N88, N86, N83, N71);
or OR2 (N89, N88, N15);
buf BUF1 (N90, N73);
not NOT1 (N91, N71);
nor NOR2 (N92, N90, N62);
buf BUF1 (N93, N91);
and AND3 (N94, N64, N72, N54);
not NOT1 (N95, N75);
and AND3 (N96, N78, N11, N67);
xor XOR2 (N97, N94, N22);
xor XOR2 (N98, N96, N90);
nor NOR2 (N99, N89, N19);
nand NAND2 (N100, N85, N97);
or OR4 (N101, N38, N82, N34, N40);
nand NAND2 (N102, N15, N98);
and AND3 (N103, N100, N44, N72);
buf BUF1 (N104, N33);
and AND2 (N105, N87, N34);
nor NOR2 (N106, N105, N21);
nor NOR4 (N107, N101, N14, N98, N27);
buf BUF1 (N108, N84);
nor NOR2 (N109, N107, N60);
or OR2 (N110, N93, N64);
and AND4 (N111, N109, N50, N15, N85);
nor NOR3 (N112, N102, N50, N24);
not NOT1 (N113, N104);
endmodule