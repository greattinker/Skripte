// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11;

output N910,N908,N901,N880,N909,N907,N891,N906,N900,N911;

or OR3 (N12, N11, N3, N7);
not NOT1 (N13, N9);
or OR3 (N14, N1, N13, N3);
or OR2 (N15, N14, N8);
nor NOR4 (N16, N14, N2, N3, N14);
not NOT1 (N17, N5);
xor XOR2 (N18, N2, N6);
nor NOR2 (N19, N1, N9);
or OR2 (N20, N7, N16);
not NOT1 (N21, N4);
xor XOR2 (N22, N13, N19);
or OR3 (N23, N2, N11, N9);
and AND4 (N24, N21, N17, N9, N5);
buf BUF1 (N25, N9);
not NOT1 (N26, N9);
xor XOR2 (N27, N19, N26);
nand NAND2 (N28, N23, N27);
and AND3 (N29, N6, N26, N21);
and AND3 (N30, N16, N3, N13);
nor NOR4 (N31, N20, N7, N9, N15);
nor NOR2 (N32, N19, N13);
nand NAND2 (N33, N24, N14);
nand NAND2 (N34, N32, N17);
buf BUF1 (N35, N28);
buf BUF1 (N36, N25);
buf BUF1 (N37, N22);
nor NOR4 (N38, N18, N23, N18, N14);
or OR3 (N39, N29, N12, N2);
or OR3 (N40, N26, N39, N15);
buf BUF1 (N41, N31);
nor NOR2 (N42, N2, N19);
and AND3 (N43, N30, N32, N31);
and AND4 (N44, N42, N19, N2, N10);
and AND3 (N45, N33, N21, N26);
xor XOR2 (N46, N44, N44);
and AND2 (N47, N37, N25);
nor NOR3 (N48, N35, N41, N29);
or OR2 (N49, N24, N31);
buf BUF1 (N50, N47);
buf BUF1 (N51, N38);
and AND2 (N52, N34, N18);
and AND3 (N53, N36, N42, N24);
or OR3 (N54, N52, N17, N28);
and AND2 (N55, N48, N36);
or OR2 (N56, N43, N7);
or OR2 (N57, N56, N9);
xor XOR2 (N58, N53, N7);
nor NOR4 (N59, N57, N30, N31, N13);
or OR2 (N60, N45, N30);
and AND2 (N61, N50, N51);
nand NAND4 (N62, N36, N17, N13, N31);
nor NOR3 (N63, N54, N25, N62);
buf BUF1 (N64, N57);
buf BUF1 (N65, N59);
nand NAND4 (N66, N64, N24, N27, N28);
nand NAND4 (N67, N60, N40, N56, N35);
buf BUF1 (N68, N64);
xor XOR2 (N69, N63, N39);
and AND4 (N70, N66, N40, N19, N5);
nor NOR4 (N71, N46, N18, N27, N47);
nor NOR4 (N72, N69, N61, N44, N63);
nor NOR3 (N73, N30, N49, N36);
not NOT1 (N74, N26);
buf BUF1 (N75, N70);
xor XOR2 (N76, N71, N17);
not NOT1 (N77, N58);
not NOT1 (N78, N73);
nand NAND3 (N79, N55, N57, N77);
not NOT1 (N80, N2);
nor NOR4 (N81, N80, N6, N61, N27);
not NOT1 (N82, N74);
not NOT1 (N83, N68);
xor XOR2 (N84, N67, N14);
or OR3 (N85, N65, N22, N8);
nor NOR2 (N86, N81, N43);
buf BUF1 (N87, N72);
buf BUF1 (N88, N87);
not NOT1 (N89, N84);
or OR4 (N90, N83, N12, N49, N19);
and AND2 (N91, N88, N74);
nand NAND4 (N92, N91, N91, N86, N27);
xor XOR2 (N93, N89, N55);
xor XOR2 (N94, N49, N89);
or OR4 (N95, N85, N31, N39, N11);
buf BUF1 (N96, N82);
nand NAND2 (N97, N75, N60);
nand NAND4 (N98, N92, N41, N20, N5);
or OR2 (N99, N76, N37);
buf BUF1 (N100, N93);
not NOT1 (N101, N99);
not NOT1 (N102, N97);
xor XOR2 (N103, N95, N74);
and AND3 (N104, N100, N21, N22);
xor XOR2 (N105, N102, N72);
nor NOR3 (N106, N94, N58, N94);
and AND2 (N107, N96, N103);
or OR2 (N108, N100, N7);
or OR3 (N109, N79, N20, N42);
or OR4 (N110, N104, N87, N26, N73);
and AND2 (N111, N106, N94);
xor XOR2 (N112, N107, N30);
and AND3 (N113, N78, N39, N107);
nor NOR2 (N114, N112, N95);
or OR2 (N115, N90, N104);
nor NOR2 (N116, N114, N1);
buf BUF1 (N117, N110);
xor XOR2 (N118, N98, N79);
nand NAND4 (N119, N109, N75, N60, N51);
xor XOR2 (N120, N101, N83);
or OR2 (N121, N118, N100);
xor XOR2 (N122, N113, N2);
xor XOR2 (N123, N111, N95);
buf BUF1 (N124, N115);
buf BUF1 (N125, N105);
buf BUF1 (N126, N119);
and AND3 (N127, N108, N64, N68);
or OR3 (N128, N124, N74, N98);
not NOT1 (N129, N121);
buf BUF1 (N130, N129);
buf BUF1 (N131, N120);
xor XOR2 (N132, N126, N36);
or OR4 (N133, N123, N58, N94, N2);
buf BUF1 (N134, N131);
not NOT1 (N135, N116);
xor XOR2 (N136, N127, N44);
and AND3 (N137, N130, N72, N42);
xor XOR2 (N138, N135, N57);
nor NOR4 (N139, N133, N13, N42, N83);
nor NOR3 (N140, N132, N108, N15);
or OR3 (N141, N128, N23, N138);
or OR2 (N142, N84, N51);
xor XOR2 (N143, N140, N115);
xor XOR2 (N144, N139, N57);
not NOT1 (N145, N122);
xor XOR2 (N146, N145, N56);
nand NAND2 (N147, N141, N120);
nor NOR4 (N148, N142, N114, N108, N92);
buf BUF1 (N149, N148);
xor XOR2 (N150, N137, N125);
not NOT1 (N151, N124);
not NOT1 (N152, N149);
or OR3 (N153, N147, N130, N80);
xor XOR2 (N154, N136, N142);
and AND3 (N155, N153, N49, N24);
not NOT1 (N156, N155);
nor NOR3 (N157, N144, N144, N27);
not NOT1 (N158, N152);
nor NOR2 (N159, N146, N32);
and AND2 (N160, N156, N69);
nand NAND2 (N161, N160, N112);
or OR2 (N162, N158, N151);
xor XOR2 (N163, N50, N139);
nor NOR3 (N164, N159, N58, N9);
and AND2 (N165, N157, N117);
nor NOR3 (N166, N142, N151, N8);
nor NOR4 (N167, N166, N82, N56, N75);
nor NOR3 (N168, N134, N43, N88);
not NOT1 (N169, N165);
nand NAND2 (N170, N143, N12);
buf BUF1 (N171, N168);
not NOT1 (N172, N150);
nand NAND2 (N173, N170, N69);
buf BUF1 (N174, N161);
xor XOR2 (N175, N162, N156);
or OR3 (N176, N173, N116, N160);
not NOT1 (N177, N176);
nand NAND4 (N178, N171, N11, N42, N63);
xor XOR2 (N179, N178, N6);
and AND2 (N180, N177, N121);
or OR4 (N181, N169, N115, N9, N22);
not NOT1 (N182, N175);
and AND2 (N183, N180, N124);
not NOT1 (N184, N164);
and AND2 (N185, N172, N89);
and AND2 (N186, N183, N92);
or OR3 (N187, N154, N147, N122);
and AND2 (N188, N167, N174);
nor NOR4 (N189, N69, N74, N105, N82);
not NOT1 (N190, N182);
buf BUF1 (N191, N188);
nor NOR2 (N192, N190, N38);
not NOT1 (N193, N185);
buf BUF1 (N194, N189);
buf BUF1 (N195, N191);
xor XOR2 (N196, N194, N180);
or OR2 (N197, N179, N129);
not NOT1 (N198, N195);
or OR4 (N199, N184, N15, N116, N36);
buf BUF1 (N200, N198);
xor XOR2 (N201, N187, N176);
buf BUF1 (N202, N200);
or OR4 (N203, N196, N65, N23, N61);
or OR2 (N204, N192, N30);
nand NAND4 (N205, N204, N181, N116, N85);
nand NAND4 (N206, N90, N57, N16, N148);
buf BUF1 (N207, N206);
and AND4 (N208, N193, N75, N118, N105);
nor NOR4 (N209, N208, N13, N135, N37);
or OR4 (N210, N203, N107, N51, N52);
or OR2 (N211, N205, N62);
xor XOR2 (N212, N163, N103);
or OR4 (N213, N211, N103, N86, N2);
nand NAND4 (N214, N186, N184, N185, N7);
not NOT1 (N215, N199);
nor NOR3 (N216, N207, N213, N83);
not NOT1 (N217, N75);
and AND3 (N218, N209, N38, N49);
not NOT1 (N219, N217);
xor XOR2 (N220, N219, N9);
and AND3 (N221, N202, N23, N180);
or OR4 (N222, N212, N149, N137, N189);
xor XOR2 (N223, N220, N31);
and AND3 (N224, N221, N132, N105);
nor NOR2 (N225, N216, N141);
and AND4 (N226, N224, N6, N129, N196);
buf BUF1 (N227, N210);
nor NOR4 (N228, N197, N49, N18, N99);
xor XOR2 (N229, N214, N205);
and AND2 (N230, N226, N127);
buf BUF1 (N231, N218);
or OR3 (N232, N230, N93, N22);
not NOT1 (N233, N223);
nor NOR2 (N234, N215, N186);
or OR4 (N235, N228, N6, N81, N134);
not NOT1 (N236, N231);
or OR2 (N237, N227, N51);
not NOT1 (N238, N222);
buf BUF1 (N239, N234);
nor NOR3 (N240, N237, N141, N71);
and AND3 (N241, N238, N84, N51);
and AND3 (N242, N229, N203, N55);
buf BUF1 (N243, N240);
nand NAND2 (N244, N242, N111);
not NOT1 (N245, N239);
nand NAND2 (N246, N244, N135);
or OR2 (N247, N233, N126);
or OR4 (N248, N241, N160, N72, N172);
or OR2 (N249, N246, N92);
buf BUF1 (N250, N248);
not NOT1 (N251, N245);
xor XOR2 (N252, N235, N156);
nand NAND2 (N253, N201, N63);
or OR4 (N254, N247, N55, N227, N252);
not NOT1 (N255, N193);
not NOT1 (N256, N232);
buf BUF1 (N257, N236);
or OR4 (N258, N254, N91, N86, N3);
or OR3 (N259, N243, N67, N196);
or OR2 (N260, N258, N147);
nor NOR2 (N261, N225, N53);
not NOT1 (N262, N250);
or OR4 (N263, N256, N26, N61, N229);
nand NAND3 (N264, N260, N119, N177);
not NOT1 (N265, N253);
or OR3 (N266, N264, N131, N187);
or OR2 (N267, N251, N6);
and AND3 (N268, N257, N12, N149);
nor NOR3 (N269, N259, N55, N64);
xor XOR2 (N270, N269, N120);
nand NAND3 (N271, N270, N268, N145);
or OR2 (N272, N85, N80);
or OR3 (N273, N262, N220, N47);
not NOT1 (N274, N267);
nand NAND4 (N275, N263, N179, N130, N12);
or OR2 (N276, N272, N151);
nand NAND2 (N277, N274, N46);
nor NOR3 (N278, N275, N65, N273);
or OR3 (N279, N158, N72, N110);
and AND4 (N280, N255, N149, N13, N38);
xor XOR2 (N281, N278, N254);
nor NOR4 (N282, N265, N78, N33, N160);
nor NOR4 (N283, N249, N105, N39, N112);
or OR2 (N284, N282, N128);
xor XOR2 (N285, N279, N33);
nand NAND2 (N286, N284, N72);
or OR2 (N287, N281, N272);
and AND3 (N288, N266, N173, N8);
and AND2 (N289, N286, N273);
xor XOR2 (N290, N288, N152);
not NOT1 (N291, N283);
buf BUF1 (N292, N280);
or OR4 (N293, N289, N193, N233, N42);
and AND4 (N294, N292, N125, N248, N3);
buf BUF1 (N295, N293);
nand NAND3 (N296, N294, N164, N47);
or OR3 (N297, N261, N107, N15);
or OR3 (N298, N271, N213, N144);
and AND4 (N299, N295, N163, N35, N18);
and AND2 (N300, N287, N231);
xor XOR2 (N301, N276, N179);
nand NAND3 (N302, N296, N16, N155);
and AND4 (N303, N297, N82, N243, N111);
and AND3 (N304, N298, N241, N5);
not NOT1 (N305, N277);
not NOT1 (N306, N285);
nor NOR2 (N307, N302, N44);
xor XOR2 (N308, N300, N77);
or OR2 (N309, N308, N124);
buf BUF1 (N310, N290);
nor NOR3 (N311, N303, N46, N260);
or OR2 (N312, N304, N311);
xor XOR2 (N313, N90, N238);
buf BUF1 (N314, N305);
buf BUF1 (N315, N299);
nand NAND4 (N316, N313, N276, N88, N237);
buf BUF1 (N317, N306);
or OR2 (N318, N314, N218);
and AND3 (N319, N318, N47, N6);
and AND3 (N320, N316, N17, N22);
nand NAND4 (N321, N301, N204, N117, N234);
nand NAND4 (N322, N309, N284, N70, N90);
and AND3 (N323, N310, N94, N211);
and AND4 (N324, N320, N301, N143, N295);
and AND2 (N325, N317, N7);
buf BUF1 (N326, N319);
xor XOR2 (N327, N321, N153);
xor XOR2 (N328, N326, N153);
nand NAND4 (N329, N291, N274, N157, N35);
nor NOR3 (N330, N307, N255, N316);
and AND2 (N331, N328, N18);
xor XOR2 (N332, N331, N307);
not NOT1 (N333, N322);
nand NAND4 (N334, N323, N45, N282, N176);
and AND4 (N335, N332, N156, N122, N65);
and AND4 (N336, N333, N34, N90, N291);
nand NAND4 (N337, N329, N258, N158, N88);
not NOT1 (N338, N312);
buf BUF1 (N339, N327);
nand NAND2 (N340, N330, N165);
xor XOR2 (N341, N334, N250);
xor XOR2 (N342, N339, N5);
and AND2 (N343, N341, N271);
buf BUF1 (N344, N343);
buf BUF1 (N345, N336);
nand NAND2 (N346, N335, N281);
buf BUF1 (N347, N345);
buf BUF1 (N348, N342);
not NOT1 (N349, N325);
nor NOR3 (N350, N337, N175, N224);
or OR2 (N351, N349, N224);
and AND4 (N352, N348, N137, N272, N203);
buf BUF1 (N353, N340);
buf BUF1 (N354, N352);
or OR4 (N355, N344, N37, N6, N86);
or OR3 (N356, N354, N176, N20);
nor NOR4 (N357, N353, N32, N279, N95);
xor XOR2 (N358, N315, N249);
not NOT1 (N359, N351);
buf BUF1 (N360, N359);
buf BUF1 (N361, N347);
and AND3 (N362, N338, N113, N308);
buf BUF1 (N363, N324);
nand NAND3 (N364, N356, N363, N245);
nand NAND3 (N365, N346, N118, N162);
not NOT1 (N366, N260);
buf BUF1 (N367, N360);
xor XOR2 (N368, N365, N186);
and AND4 (N369, N367, N241, N358, N239);
xor XOR2 (N370, N14, N242);
and AND3 (N371, N369, N164, N293);
nor NOR3 (N372, N364, N65, N151);
buf BUF1 (N373, N372);
not NOT1 (N374, N355);
buf BUF1 (N375, N371);
nor NOR3 (N376, N362, N15, N348);
or OR2 (N377, N357, N195);
nand NAND4 (N378, N370, N242, N325, N184);
nor NOR4 (N379, N366, N24, N321, N272);
not NOT1 (N380, N376);
nand NAND3 (N381, N374, N354, N39);
and AND3 (N382, N361, N104, N69);
nor NOR4 (N383, N381, N203, N137, N132);
and AND3 (N384, N383, N333, N226);
and AND4 (N385, N377, N211, N54, N73);
buf BUF1 (N386, N385);
nor NOR2 (N387, N380, N384);
and AND4 (N388, N109, N321, N361, N81);
and AND3 (N389, N378, N220, N255);
or OR3 (N390, N387, N72, N255);
not NOT1 (N391, N388);
nand NAND4 (N392, N390, N344, N11, N352);
nor NOR3 (N393, N389, N26, N377);
or OR3 (N394, N350, N80, N73);
nand NAND4 (N395, N373, N99, N148, N338);
buf BUF1 (N396, N391);
xor XOR2 (N397, N375, N258);
nor NOR4 (N398, N382, N220, N310, N244);
not NOT1 (N399, N392);
not NOT1 (N400, N386);
not NOT1 (N401, N394);
and AND3 (N402, N396, N203, N360);
not NOT1 (N403, N393);
nor NOR4 (N404, N397, N88, N155, N371);
or OR4 (N405, N379, N144, N149, N293);
or OR4 (N406, N402, N5, N353, N125);
or OR2 (N407, N399, N45);
and AND2 (N408, N395, N74);
buf BUF1 (N409, N407);
not NOT1 (N410, N368);
not NOT1 (N411, N403);
nor NOR4 (N412, N411, N163, N249, N376);
or OR4 (N413, N410, N374, N105, N271);
not NOT1 (N414, N404);
buf BUF1 (N415, N406);
and AND2 (N416, N415, N201);
nor NOR3 (N417, N413, N70, N349);
nand NAND3 (N418, N414, N371, N278);
xor XOR2 (N419, N401, N164);
xor XOR2 (N420, N400, N207);
buf BUF1 (N421, N420);
nand NAND2 (N422, N405, N205);
or OR2 (N423, N422, N109);
xor XOR2 (N424, N412, N231);
nand NAND4 (N425, N398, N284, N229, N394);
nor NOR3 (N426, N424, N231, N29);
nand NAND3 (N427, N421, N194, N9);
nor NOR4 (N428, N416, N112, N187, N1);
or OR4 (N429, N425, N374, N31, N403);
xor XOR2 (N430, N426, N278);
or OR4 (N431, N418, N177, N320, N270);
and AND2 (N432, N428, N291);
nand NAND3 (N433, N423, N286, N294);
or OR2 (N434, N427, N290);
not NOT1 (N435, N433);
or OR2 (N436, N408, N39);
buf BUF1 (N437, N434);
or OR3 (N438, N432, N169, N35);
nor NOR3 (N439, N436, N33, N37);
nor NOR4 (N440, N431, N296, N94, N115);
not NOT1 (N441, N430);
xor XOR2 (N442, N440, N306);
xor XOR2 (N443, N442, N237);
nor NOR2 (N444, N429, N187);
nor NOR3 (N445, N439, N262, N313);
nor NOR4 (N446, N438, N288, N25, N150);
xor XOR2 (N447, N409, N244);
buf BUF1 (N448, N419);
nor NOR4 (N449, N437, N423, N382, N186);
or OR2 (N450, N447, N109);
not NOT1 (N451, N450);
xor XOR2 (N452, N449, N123);
buf BUF1 (N453, N417);
not NOT1 (N454, N452);
nor NOR2 (N455, N445, N25);
xor XOR2 (N456, N446, N99);
nand NAND4 (N457, N454, N376, N421, N30);
not NOT1 (N458, N457);
and AND3 (N459, N443, N72, N174);
xor XOR2 (N460, N453, N221);
xor XOR2 (N461, N458, N260);
nor NOR4 (N462, N448, N229, N460, N1);
buf BUF1 (N463, N294);
or OR2 (N464, N462, N352);
buf BUF1 (N465, N435);
not NOT1 (N466, N455);
not NOT1 (N467, N464);
not NOT1 (N468, N463);
nor NOR4 (N469, N444, N3, N53, N128);
buf BUF1 (N470, N461);
xor XOR2 (N471, N451, N426);
nor NOR2 (N472, N441, N374);
nor NOR2 (N473, N468, N84);
xor XOR2 (N474, N467, N50);
and AND2 (N475, N470, N417);
buf BUF1 (N476, N474);
nand NAND2 (N477, N466, N163);
nor NOR2 (N478, N475, N238);
and AND4 (N479, N478, N181, N222, N168);
buf BUF1 (N480, N476);
buf BUF1 (N481, N477);
xor XOR2 (N482, N471, N55);
xor XOR2 (N483, N480, N309);
buf BUF1 (N484, N469);
not NOT1 (N485, N482);
buf BUF1 (N486, N459);
xor XOR2 (N487, N481, N456);
nand NAND4 (N488, N454, N257, N336, N437);
and AND3 (N489, N465, N460, N276);
or OR2 (N490, N473, N135);
nor NOR3 (N491, N485, N300, N374);
nor NOR4 (N492, N491, N132, N103, N338);
nor NOR3 (N493, N490, N403, N334);
nor NOR2 (N494, N483, N77);
and AND3 (N495, N494, N451, N305);
and AND3 (N496, N495, N121, N191);
nor NOR2 (N497, N496, N276);
buf BUF1 (N498, N492);
buf BUF1 (N499, N493);
xor XOR2 (N500, N499, N288);
not NOT1 (N501, N472);
or OR4 (N502, N486, N208, N345, N175);
nor NOR3 (N503, N501, N401, N472);
and AND2 (N504, N498, N232);
buf BUF1 (N505, N500);
nand NAND4 (N506, N479, N337, N136, N447);
nand NAND4 (N507, N506, N46, N205, N452);
buf BUF1 (N508, N489);
xor XOR2 (N509, N487, N325);
nor NOR4 (N510, N503, N471, N233, N309);
buf BUF1 (N511, N488);
xor XOR2 (N512, N504, N274);
buf BUF1 (N513, N505);
xor XOR2 (N514, N502, N408);
xor XOR2 (N515, N497, N482);
and AND3 (N516, N513, N2, N105);
buf BUF1 (N517, N515);
or OR4 (N518, N507, N495, N57, N426);
buf BUF1 (N519, N514);
nor NOR4 (N520, N518, N39, N461, N244);
nor NOR3 (N521, N508, N333, N42);
or OR3 (N522, N517, N447, N390);
or OR4 (N523, N484, N289, N117, N78);
nor NOR3 (N524, N512, N511, N184);
nor NOR4 (N525, N289, N380, N358, N512);
and AND2 (N526, N520, N521);
xor XOR2 (N527, N325, N337);
nand NAND2 (N528, N523, N319);
nor NOR3 (N529, N522, N65, N106);
nor NOR3 (N530, N509, N403, N444);
nor NOR2 (N531, N530, N348);
or OR2 (N532, N519, N403);
not NOT1 (N533, N529);
nand NAND4 (N534, N528, N400, N112, N12);
nand NAND3 (N535, N516, N254, N432);
nor NOR2 (N536, N531, N375);
nand NAND4 (N537, N533, N379, N439, N225);
or OR2 (N538, N524, N127);
nor NOR3 (N539, N525, N434, N393);
and AND3 (N540, N537, N171, N139);
nand NAND3 (N541, N526, N248, N431);
or OR2 (N542, N534, N140);
or OR3 (N543, N510, N138, N186);
nor NOR2 (N544, N535, N288);
and AND2 (N545, N536, N516);
or OR4 (N546, N539, N234, N422, N104);
buf BUF1 (N547, N544);
buf BUF1 (N548, N527);
buf BUF1 (N549, N532);
buf BUF1 (N550, N538);
and AND2 (N551, N546, N520);
buf BUF1 (N552, N549);
buf BUF1 (N553, N551);
nand NAND2 (N554, N545, N89);
xor XOR2 (N555, N548, N463);
xor XOR2 (N556, N543, N332);
nand NAND4 (N557, N552, N80, N233, N240);
or OR2 (N558, N541, N323);
buf BUF1 (N559, N554);
buf BUF1 (N560, N550);
buf BUF1 (N561, N556);
nor NOR4 (N562, N559, N442, N307, N266);
nand NAND3 (N563, N561, N251, N469);
buf BUF1 (N564, N558);
not NOT1 (N565, N562);
nand NAND2 (N566, N540, N437);
and AND3 (N567, N565, N334, N488);
xor XOR2 (N568, N553, N286);
buf BUF1 (N569, N566);
nand NAND2 (N570, N569, N500);
and AND2 (N571, N547, N330);
and AND2 (N572, N570, N541);
nor NOR3 (N573, N571, N413, N511);
xor XOR2 (N574, N568, N515);
not NOT1 (N575, N542);
or OR2 (N576, N563, N495);
not NOT1 (N577, N576);
nand NAND3 (N578, N557, N93, N481);
and AND2 (N579, N574, N507);
and AND2 (N580, N572, N281);
or OR3 (N581, N560, N393, N168);
not NOT1 (N582, N577);
or OR4 (N583, N564, N289, N213, N450);
buf BUF1 (N584, N578);
and AND4 (N585, N573, N203, N288, N23);
not NOT1 (N586, N583);
nor NOR3 (N587, N581, N384, N91);
or OR2 (N588, N575, N396);
not NOT1 (N589, N587);
not NOT1 (N590, N580);
and AND2 (N591, N555, N63);
not NOT1 (N592, N591);
buf BUF1 (N593, N592);
nand NAND4 (N594, N567, N264, N190, N528);
nor NOR3 (N595, N586, N19, N297);
nor NOR3 (N596, N593, N91, N446);
buf BUF1 (N597, N584);
and AND3 (N598, N585, N374, N407);
nor NOR3 (N599, N595, N406, N231);
nor NOR3 (N600, N598, N331, N77);
buf BUF1 (N601, N582);
nor NOR3 (N602, N597, N294, N404);
buf BUF1 (N603, N600);
buf BUF1 (N604, N589);
buf BUF1 (N605, N599);
xor XOR2 (N606, N590, N464);
and AND4 (N607, N604, N543, N407, N406);
xor XOR2 (N608, N596, N164);
or OR3 (N609, N588, N170, N470);
or OR4 (N610, N605, N388, N344, N355);
not NOT1 (N611, N608);
nor NOR3 (N612, N601, N393, N435);
xor XOR2 (N613, N602, N569);
nand NAND4 (N614, N609, N222, N446, N141);
or OR4 (N615, N606, N352, N504, N533);
nand NAND3 (N616, N579, N294, N250);
nand NAND2 (N617, N610, N610);
xor XOR2 (N618, N614, N595);
or OR4 (N619, N613, N269, N36, N159);
not NOT1 (N620, N607);
nand NAND2 (N621, N612, N164);
nand NAND3 (N622, N619, N410, N40);
and AND3 (N623, N603, N241, N149);
nand NAND4 (N624, N617, N165, N244, N445);
nor NOR4 (N625, N618, N364, N200, N544);
and AND3 (N626, N611, N473, N409);
xor XOR2 (N627, N621, N599);
and AND3 (N628, N616, N585, N296);
xor XOR2 (N629, N625, N327);
not NOT1 (N630, N627);
or OR2 (N631, N628, N150);
or OR4 (N632, N615, N205, N625, N23);
and AND4 (N633, N622, N174, N75, N364);
buf BUF1 (N634, N626);
nand NAND2 (N635, N634, N507);
xor XOR2 (N636, N594, N469);
nor NOR3 (N637, N620, N129, N344);
not NOT1 (N638, N630);
buf BUF1 (N639, N633);
not NOT1 (N640, N636);
xor XOR2 (N641, N632, N635);
nor NOR2 (N642, N39, N352);
nand NAND3 (N643, N638, N455, N258);
nand NAND2 (N644, N623, N378);
and AND4 (N645, N637, N73, N100, N381);
nand NAND2 (N646, N639, N517);
buf BUF1 (N647, N644);
or OR4 (N648, N640, N163, N382, N28);
buf BUF1 (N649, N648);
or OR3 (N650, N631, N159, N151);
not NOT1 (N651, N649);
not NOT1 (N652, N642);
xor XOR2 (N653, N646, N52);
nor NOR3 (N654, N645, N99, N244);
or OR4 (N655, N654, N582, N444, N422);
not NOT1 (N656, N629);
not NOT1 (N657, N653);
nor NOR4 (N658, N641, N235, N125, N383);
xor XOR2 (N659, N647, N270);
nor NOR2 (N660, N651, N596);
not NOT1 (N661, N658);
or OR2 (N662, N624, N399);
not NOT1 (N663, N662);
nor NOR4 (N664, N663, N650, N261, N381);
buf BUF1 (N665, N648);
xor XOR2 (N666, N661, N29);
or OR4 (N667, N652, N391, N363, N125);
and AND2 (N668, N643, N609);
nor NOR3 (N669, N655, N360, N509);
buf BUF1 (N670, N668);
or OR3 (N671, N666, N501, N424);
not NOT1 (N672, N659);
not NOT1 (N673, N660);
xor XOR2 (N674, N657, N184);
not NOT1 (N675, N672);
nor NOR4 (N676, N670, N587, N474, N204);
xor XOR2 (N677, N671, N333);
and AND2 (N678, N656, N628);
buf BUF1 (N679, N678);
or OR3 (N680, N667, N275, N164);
and AND4 (N681, N676, N146, N481, N117);
nor NOR3 (N682, N669, N130, N244);
not NOT1 (N683, N664);
not NOT1 (N684, N673);
and AND2 (N685, N665, N109);
and AND4 (N686, N681, N679, N208, N163);
nor NOR3 (N687, N288, N195, N421);
nand NAND3 (N688, N675, N583, N273);
nand NAND4 (N689, N674, N56, N165, N60);
xor XOR2 (N690, N686, N617);
or OR3 (N691, N682, N469, N100);
nor NOR2 (N692, N690, N62);
not NOT1 (N693, N685);
buf BUF1 (N694, N692);
buf BUF1 (N695, N687);
and AND3 (N696, N693, N502, N274);
nor NOR2 (N697, N696, N620);
and AND4 (N698, N684, N351, N619, N392);
nor NOR2 (N699, N695, N68);
and AND4 (N700, N691, N288, N496, N672);
or OR3 (N701, N683, N650, N6);
or OR4 (N702, N701, N652, N452, N671);
and AND4 (N703, N677, N649, N426, N338);
or OR2 (N704, N689, N398);
nor NOR2 (N705, N700, N32);
nand NAND4 (N706, N702, N174, N4, N164);
or OR2 (N707, N694, N147);
and AND3 (N708, N680, N93, N84);
or OR4 (N709, N705, N226, N408, N561);
nand NAND4 (N710, N704, N176, N567, N678);
nand NAND4 (N711, N709, N645, N637, N653);
xor XOR2 (N712, N697, N3);
buf BUF1 (N713, N688);
xor XOR2 (N714, N698, N690);
nand NAND2 (N715, N713, N637);
nand NAND2 (N716, N706, N227);
xor XOR2 (N717, N708, N507);
and AND2 (N718, N717, N136);
or OR3 (N719, N711, N655, N568);
nand NAND3 (N720, N703, N441, N564);
xor XOR2 (N721, N720, N84);
or OR2 (N722, N714, N362);
xor XOR2 (N723, N699, N236);
nand NAND4 (N724, N707, N396, N590, N209);
not NOT1 (N725, N715);
or OR4 (N726, N718, N235, N717, N95);
and AND2 (N727, N726, N287);
and AND4 (N728, N712, N595, N485, N407);
nor NOR3 (N729, N721, N533, N708);
buf BUF1 (N730, N729);
nor NOR4 (N731, N722, N288, N275, N402);
xor XOR2 (N732, N728, N476);
and AND2 (N733, N716, N341);
not NOT1 (N734, N733);
or OR2 (N735, N710, N187);
nand NAND3 (N736, N734, N132, N663);
not NOT1 (N737, N732);
buf BUF1 (N738, N724);
nand NAND4 (N739, N735, N504, N626, N415);
xor XOR2 (N740, N723, N473);
not NOT1 (N741, N719);
and AND4 (N742, N738, N484, N692, N203);
not NOT1 (N743, N739);
buf BUF1 (N744, N731);
buf BUF1 (N745, N727);
or OR2 (N746, N743, N134);
xor XOR2 (N747, N745, N114);
xor XOR2 (N748, N730, N669);
nor NOR2 (N749, N736, N270);
xor XOR2 (N750, N742, N642);
not NOT1 (N751, N740);
not NOT1 (N752, N725);
buf BUF1 (N753, N741);
nor NOR3 (N754, N751, N62, N244);
and AND4 (N755, N748, N159, N626, N412);
nand NAND4 (N756, N737, N604, N55, N623);
nor NOR4 (N757, N756, N720, N367, N756);
nor NOR2 (N758, N747, N705);
or OR4 (N759, N750, N83, N449, N641);
nand NAND2 (N760, N749, N233);
nand NAND4 (N761, N752, N743, N76, N188);
nand NAND2 (N762, N755, N43);
or OR3 (N763, N761, N631, N436);
and AND2 (N764, N762, N335);
xor XOR2 (N765, N763, N271);
buf BUF1 (N766, N757);
xor XOR2 (N767, N760, N568);
not NOT1 (N768, N759);
buf BUF1 (N769, N754);
or OR4 (N770, N753, N329, N678, N279);
xor XOR2 (N771, N765, N385);
nor NOR3 (N772, N766, N150, N481);
xor XOR2 (N773, N768, N50);
not NOT1 (N774, N746);
nor NOR2 (N775, N769, N567);
nand NAND2 (N776, N767, N138);
and AND3 (N777, N770, N670, N764);
nand NAND3 (N778, N309, N371, N141);
buf BUF1 (N779, N744);
xor XOR2 (N780, N776, N15);
not NOT1 (N781, N775);
or OR3 (N782, N771, N493, N691);
buf BUF1 (N783, N780);
nand NAND3 (N784, N783, N217, N747);
not NOT1 (N785, N773);
and AND4 (N786, N774, N341, N356, N479);
nor NOR2 (N787, N786, N609);
nand NAND4 (N788, N782, N447, N729, N606);
nand NAND4 (N789, N777, N782, N153, N9);
nand NAND2 (N790, N758, N679);
nand NAND3 (N791, N779, N627, N350);
buf BUF1 (N792, N772);
nand NAND2 (N793, N784, N687);
nor NOR2 (N794, N785, N182);
xor XOR2 (N795, N792, N376);
nand NAND2 (N796, N791, N369);
buf BUF1 (N797, N787);
nor NOR3 (N798, N793, N393, N771);
xor XOR2 (N799, N790, N225);
and AND4 (N800, N794, N359, N507, N52);
buf BUF1 (N801, N788);
not NOT1 (N802, N796);
and AND4 (N803, N778, N469, N799, N519);
not NOT1 (N804, N554);
not NOT1 (N805, N797);
buf BUF1 (N806, N801);
and AND3 (N807, N789, N211, N463);
not NOT1 (N808, N802);
not NOT1 (N809, N795);
or OR4 (N810, N805, N414, N56, N681);
xor XOR2 (N811, N804, N631);
or OR4 (N812, N781, N599, N724, N226);
or OR3 (N813, N800, N456, N303);
nor NOR4 (N814, N806, N264, N489, N343);
nor NOR2 (N815, N807, N196);
and AND2 (N816, N798, N500);
nand NAND3 (N817, N814, N16, N672);
xor XOR2 (N818, N812, N654);
nor NOR4 (N819, N815, N502, N446, N699);
xor XOR2 (N820, N818, N387);
buf BUF1 (N821, N820);
and AND2 (N822, N810, N217);
nand NAND2 (N823, N813, N330);
nand NAND4 (N824, N821, N295, N172, N813);
or OR4 (N825, N817, N766, N645, N513);
xor XOR2 (N826, N822, N436);
and AND3 (N827, N803, N343, N494);
or OR3 (N828, N823, N234, N121);
buf BUF1 (N829, N827);
xor XOR2 (N830, N811, N640);
not NOT1 (N831, N825);
or OR2 (N832, N809, N192);
xor XOR2 (N833, N816, N126);
buf BUF1 (N834, N819);
buf BUF1 (N835, N832);
and AND2 (N836, N828, N244);
nand NAND2 (N837, N826, N518);
nand NAND2 (N838, N836, N599);
not NOT1 (N839, N833);
and AND3 (N840, N835, N557, N625);
buf BUF1 (N841, N831);
not NOT1 (N842, N808);
nand NAND3 (N843, N837, N720, N555);
not NOT1 (N844, N843);
or OR2 (N845, N834, N298);
nand NAND3 (N846, N830, N326, N667);
and AND4 (N847, N840, N202, N456, N372);
not NOT1 (N848, N824);
nor NOR4 (N849, N848, N414, N7, N806);
xor XOR2 (N850, N849, N417);
and AND4 (N851, N850, N689, N846, N830);
nor NOR3 (N852, N150, N788, N395);
not NOT1 (N853, N852);
xor XOR2 (N854, N845, N411);
xor XOR2 (N855, N839, N850);
nand NAND4 (N856, N854, N60, N331, N337);
or OR4 (N857, N856, N491, N186, N849);
xor XOR2 (N858, N857, N374);
xor XOR2 (N859, N844, N91);
not NOT1 (N860, N838);
or OR4 (N861, N829, N300, N416, N340);
buf BUF1 (N862, N855);
nand NAND3 (N863, N858, N213, N605);
not NOT1 (N864, N859);
nor NOR3 (N865, N864, N406, N169);
and AND4 (N866, N860, N551, N802, N807);
nand NAND3 (N867, N841, N568, N255);
xor XOR2 (N868, N842, N748);
or OR2 (N869, N851, N532);
nor NOR4 (N870, N863, N620, N301, N788);
buf BUF1 (N871, N847);
xor XOR2 (N872, N868, N734);
nand NAND4 (N873, N853, N699, N110, N51);
nor NOR2 (N874, N871, N515);
or OR2 (N875, N870, N625);
and AND4 (N876, N875, N288, N825, N158);
not NOT1 (N877, N873);
nor NOR3 (N878, N877, N193, N504);
xor XOR2 (N879, N867, N878);
buf BUF1 (N880, N62);
and AND4 (N881, N872, N770, N593, N726);
nor NOR3 (N882, N869, N311, N822);
not NOT1 (N883, N882);
not NOT1 (N884, N862);
nor NOR4 (N885, N883, N154, N747, N780);
nor NOR2 (N886, N885, N667);
or OR2 (N887, N865, N862);
or OR3 (N888, N886, N462, N497);
not NOT1 (N889, N879);
not NOT1 (N890, N889);
nand NAND4 (N891, N884, N50, N480, N818);
nor NOR4 (N892, N861, N51, N163, N866);
nand NAND2 (N893, N335, N121);
nand NAND4 (N894, N893, N849, N220, N403);
buf BUF1 (N895, N888);
not NOT1 (N896, N890);
not NOT1 (N897, N876);
buf BUF1 (N898, N896);
not NOT1 (N899, N894);
nand NAND3 (N900, N892, N765, N123);
not NOT1 (N901, N899);
buf BUF1 (N902, N898);
nand NAND2 (N903, N881, N622);
and AND3 (N904, N897, N596, N834);
xor XOR2 (N905, N903, N609);
or OR3 (N906, N887, N576, N75);
buf BUF1 (N907, N905);
buf BUF1 (N908, N904);
nor NOR2 (N909, N902, N741);
xor XOR2 (N910, N874, N410);
nand NAND2 (N911, N895, N455);
endmodule