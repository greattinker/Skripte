// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24;

output N799,N811,N821,N823,N822,N795,N819,N809,N806,N824;

not NOT1 (N25, N17);
nor NOR3 (N26, N3, N17, N12);
or OR4 (N27, N1, N22, N6, N7);
and AND2 (N28, N7, N27);
or OR4 (N29, N1, N13, N12, N3);
nand NAND4 (N30, N20, N3, N10, N26);
xor XOR2 (N31, N18, N3);
nor NOR2 (N32, N1, N10);
buf BUF1 (N33, N24);
and AND4 (N34, N28, N29, N14, N12);
buf BUF1 (N35, N10);
nand NAND2 (N36, N32, N22);
and AND4 (N37, N28, N27, N24, N8);
or OR2 (N38, N28, N18);
and AND2 (N39, N18, N6);
and AND4 (N40, N25, N31, N16, N32);
nand NAND4 (N41, N9, N17, N24, N20);
buf BUF1 (N42, N33);
nand NAND4 (N43, N41, N32, N37, N4);
nor NOR2 (N44, N30, N12);
or OR4 (N45, N44, N5, N13, N1);
xor XOR2 (N46, N20, N26);
not NOT1 (N47, N39);
or OR3 (N48, N34, N3, N6);
nor NOR4 (N49, N48, N28, N6, N24);
xor XOR2 (N50, N35, N19);
and AND2 (N51, N45, N19);
nand NAND4 (N52, N51, N25, N32, N46);
xor XOR2 (N53, N12, N40);
nor NOR3 (N54, N20, N4, N5);
or OR4 (N55, N38, N6, N5, N4);
or OR4 (N56, N43, N21, N44, N19);
not NOT1 (N57, N56);
and AND2 (N58, N52, N53);
buf BUF1 (N59, N56);
or OR3 (N60, N58, N47, N39);
not NOT1 (N61, N36);
buf BUF1 (N62, N45);
xor XOR2 (N63, N61, N35);
nor NOR3 (N64, N54, N31, N22);
nor NOR2 (N65, N62, N48);
nor NOR2 (N66, N55, N54);
nand NAND2 (N67, N65, N9);
or OR4 (N68, N67, N47, N9, N29);
nand NAND3 (N69, N59, N27, N50);
buf BUF1 (N70, N14);
nand NAND3 (N71, N42, N48, N70);
xor XOR2 (N72, N50, N58);
nand NAND2 (N73, N57, N19);
and AND3 (N74, N68, N9, N63);
nor NOR3 (N75, N24, N48, N16);
buf BUF1 (N76, N64);
xor XOR2 (N77, N74, N4);
and AND2 (N78, N49, N74);
nand NAND3 (N79, N72, N14, N42);
nand NAND4 (N80, N77, N68, N68, N51);
not NOT1 (N81, N60);
not NOT1 (N82, N80);
xor XOR2 (N83, N71, N80);
xor XOR2 (N84, N76, N79);
not NOT1 (N85, N49);
and AND2 (N86, N69, N24);
nand NAND3 (N87, N78, N37, N16);
or OR2 (N88, N66, N32);
nand NAND2 (N89, N82, N17);
nor NOR4 (N90, N88, N65, N78, N87);
and AND2 (N91, N76, N66);
not NOT1 (N92, N73);
and AND3 (N93, N86, N31, N16);
and AND3 (N94, N90, N92, N29);
buf BUF1 (N95, N19);
and AND2 (N96, N75, N58);
xor XOR2 (N97, N83, N64);
nand NAND4 (N98, N81, N19, N45, N10);
nor NOR2 (N99, N84, N93);
xor XOR2 (N100, N57, N97);
xor XOR2 (N101, N100, N55);
or OR4 (N102, N63, N17, N46, N9);
buf BUF1 (N103, N101);
and AND4 (N104, N103, N18, N10, N22);
and AND2 (N105, N99, N21);
or OR2 (N106, N96, N50);
or OR2 (N107, N105, N61);
xor XOR2 (N108, N89, N94);
not NOT1 (N109, N99);
and AND2 (N110, N109, N3);
nor NOR3 (N111, N91, N87, N73);
or OR4 (N112, N106, N37, N85, N70);
not NOT1 (N113, N42);
xor XOR2 (N114, N98, N35);
not NOT1 (N115, N113);
and AND4 (N116, N111, N34, N92, N32);
or OR4 (N117, N104, N22, N98, N82);
xor XOR2 (N118, N117, N112);
nor NOR3 (N119, N92, N24, N12);
not NOT1 (N120, N118);
buf BUF1 (N121, N95);
or OR4 (N122, N115, N70, N47, N38);
xor XOR2 (N123, N120, N34);
or OR3 (N124, N102, N55, N54);
nor NOR3 (N125, N114, N90, N42);
or OR2 (N126, N108, N104);
nand NAND2 (N127, N126, N54);
nor NOR4 (N128, N123, N35, N46, N27);
xor XOR2 (N129, N125, N10);
not NOT1 (N130, N116);
xor XOR2 (N131, N107, N78);
not NOT1 (N132, N124);
or OR3 (N133, N122, N64, N132);
and AND2 (N134, N45, N20);
nor NOR2 (N135, N119, N109);
buf BUF1 (N136, N110);
nor NOR2 (N137, N127, N54);
buf BUF1 (N138, N136);
xor XOR2 (N139, N128, N16);
nor NOR2 (N140, N137, N93);
and AND2 (N141, N134, N38);
nor NOR3 (N142, N129, N77, N121);
xor XOR2 (N143, N32, N118);
nand NAND3 (N144, N133, N40, N49);
not NOT1 (N145, N142);
nor NOR2 (N146, N130, N5);
not NOT1 (N147, N131);
nor NOR2 (N148, N143, N38);
xor XOR2 (N149, N145, N69);
nand NAND4 (N150, N144, N28, N16, N81);
or OR4 (N151, N141, N125, N84, N134);
and AND4 (N152, N138, N10, N53, N54);
nand NAND3 (N153, N139, N38, N3);
not NOT1 (N154, N147);
nand NAND3 (N155, N154, N69, N19);
nor NOR2 (N156, N146, N38);
not NOT1 (N157, N151);
buf BUF1 (N158, N149);
and AND3 (N159, N135, N125, N93);
nand NAND4 (N160, N155, N61, N31, N126);
and AND4 (N161, N153, N19, N37, N106);
and AND3 (N162, N159, N25, N76);
nand NAND4 (N163, N140, N126, N55, N154);
nand NAND2 (N164, N160, N110);
buf BUF1 (N165, N152);
xor XOR2 (N166, N165, N35);
xor XOR2 (N167, N148, N132);
nand NAND2 (N168, N150, N31);
nand NAND3 (N169, N167, N84, N155);
buf BUF1 (N170, N158);
and AND2 (N171, N161, N58);
nand NAND4 (N172, N168, N96, N92, N1);
and AND3 (N173, N157, N132, N51);
not NOT1 (N174, N164);
buf BUF1 (N175, N174);
and AND3 (N176, N166, N161, N123);
buf BUF1 (N177, N162);
buf BUF1 (N178, N170);
nand NAND3 (N179, N163, N49, N125);
and AND2 (N180, N176, N97);
nand NAND4 (N181, N171, N161, N23, N150);
or OR4 (N182, N179, N93, N137, N11);
nor NOR4 (N183, N173, N82, N84, N41);
nor NOR2 (N184, N180, N43);
not NOT1 (N185, N172);
and AND4 (N186, N182, N28, N126, N99);
or OR2 (N187, N175, N28);
and AND2 (N188, N178, N121);
xor XOR2 (N189, N177, N66);
or OR3 (N190, N183, N131, N142);
buf BUF1 (N191, N169);
nor NOR3 (N192, N190, N156, N125);
buf BUF1 (N193, N97);
and AND2 (N194, N181, N33);
nor NOR3 (N195, N186, N28, N85);
nor NOR4 (N196, N184, N176, N194, N176);
not NOT1 (N197, N112);
xor XOR2 (N198, N185, N33);
and AND3 (N199, N195, N79, N49);
nand NAND3 (N200, N187, N195, N47);
xor XOR2 (N201, N189, N138);
buf BUF1 (N202, N193);
buf BUF1 (N203, N200);
nor NOR3 (N204, N198, N113, N90);
xor XOR2 (N205, N196, N20);
nor NOR4 (N206, N203, N161, N135, N77);
buf BUF1 (N207, N202);
xor XOR2 (N208, N204, N84);
or OR2 (N209, N188, N203);
nor NOR3 (N210, N191, N132, N208);
nor NOR3 (N211, N20, N88, N201);
nor NOR4 (N212, N102, N31, N171, N31);
or OR3 (N213, N212, N4, N48);
or OR4 (N214, N197, N189, N83, N147);
xor XOR2 (N215, N199, N43);
and AND4 (N216, N211, N118, N64, N47);
nand NAND4 (N217, N206, N70, N183, N139);
buf BUF1 (N218, N216);
nand NAND2 (N219, N217, N200);
xor XOR2 (N220, N192, N163);
nand NAND2 (N221, N205, N177);
nor NOR3 (N222, N209, N100, N132);
nor NOR4 (N223, N218, N59, N159, N2);
nand NAND3 (N224, N221, N24, N68);
and AND2 (N225, N222, N188);
and AND2 (N226, N214, N105);
xor XOR2 (N227, N226, N151);
nand NAND4 (N228, N224, N184, N144, N201);
xor XOR2 (N229, N225, N11);
xor XOR2 (N230, N220, N152);
xor XOR2 (N231, N219, N135);
not NOT1 (N232, N210);
buf BUF1 (N233, N229);
not NOT1 (N234, N227);
nand NAND3 (N235, N231, N13, N12);
buf BUF1 (N236, N235);
nand NAND4 (N237, N233, N100, N8, N187);
not NOT1 (N238, N228);
not NOT1 (N239, N215);
and AND2 (N240, N223, N228);
and AND2 (N241, N236, N212);
nor NOR3 (N242, N237, N73, N111);
and AND4 (N243, N234, N4, N65, N133);
nor NOR2 (N244, N230, N27);
nor NOR2 (N245, N241, N17);
or OR3 (N246, N240, N94, N186);
nand NAND4 (N247, N245, N113, N224, N2);
not NOT1 (N248, N247);
or OR3 (N249, N213, N5, N92);
or OR2 (N250, N248, N48);
or OR3 (N251, N249, N16, N152);
buf BUF1 (N252, N246);
buf BUF1 (N253, N238);
xor XOR2 (N254, N207, N119);
nor NOR2 (N255, N239, N147);
xor XOR2 (N256, N243, N99);
nor NOR4 (N257, N256, N227, N82, N72);
nor NOR2 (N258, N253, N156);
not NOT1 (N259, N257);
xor XOR2 (N260, N259, N65);
nand NAND2 (N261, N255, N10);
or OR3 (N262, N251, N181, N239);
buf BUF1 (N263, N232);
nand NAND3 (N264, N254, N125, N108);
buf BUF1 (N265, N260);
xor XOR2 (N266, N262, N61);
and AND3 (N267, N258, N105, N203);
nand NAND2 (N268, N261, N232);
xor XOR2 (N269, N268, N67);
nor NOR2 (N270, N252, N145);
nor NOR3 (N271, N267, N26, N44);
nand NAND3 (N272, N271, N267, N270);
xor XOR2 (N273, N159, N96);
nor NOR3 (N274, N265, N72, N153);
xor XOR2 (N275, N264, N177);
nand NAND4 (N276, N242, N24, N251, N63);
nor NOR3 (N277, N250, N41, N112);
xor XOR2 (N278, N276, N135);
and AND2 (N279, N272, N30);
or OR3 (N280, N273, N174, N261);
nor NOR4 (N281, N277, N14, N209, N136);
nor NOR4 (N282, N281, N105, N250, N55);
and AND4 (N283, N263, N207, N112, N154);
nand NAND2 (N284, N269, N77);
xor XOR2 (N285, N244, N71);
buf BUF1 (N286, N284);
or OR2 (N287, N278, N246);
nor NOR4 (N288, N266, N92, N97, N247);
nor NOR4 (N289, N285, N206, N38, N92);
or OR4 (N290, N282, N227, N11, N188);
xor XOR2 (N291, N288, N127);
nor NOR2 (N292, N280, N125);
or OR2 (N293, N275, N270);
nand NAND4 (N294, N289, N100, N13, N144);
or OR4 (N295, N294, N218, N65, N87);
buf BUF1 (N296, N286);
buf BUF1 (N297, N296);
or OR3 (N298, N290, N153, N182);
nor NOR2 (N299, N283, N121);
nor NOR2 (N300, N291, N95);
nand NAND2 (N301, N295, N201);
xor XOR2 (N302, N301, N155);
or OR4 (N303, N287, N11, N94, N168);
xor XOR2 (N304, N298, N173);
nor NOR2 (N305, N279, N195);
and AND4 (N306, N302, N268, N114, N241);
not NOT1 (N307, N297);
nand NAND4 (N308, N293, N58, N99, N133);
nand NAND3 (N309, N305, N294, N9);
and AND3 (N310, N292, N115, N120);
nand NAND2 (N311, N303, N84);
and AND4 (N312, N308, N18, N73, N122);
buf BUF1 (N313, N306);
buf BUF1 (N314, N313);
not NOT1 (N315, N299);
and AND2 (N316, N310, N263);
or OR3 (N317, N307, N107, N67);
buf BUF1 (N318, N312);
not NOT1 (N319, N316);
or OR4 (N320, N311, N134, N262, N115);
and AND2 (N321, N319, N315);
or OR3 (N322, N160, N221, N263);
nand NAND4 (N323, N321, N314, N206, N227);
buf BUF1 (N324, N143);
nor NOR2 (N325, N324, N72);
or OR3 (N326, N304, N212, N287);
nor NOR2 (N327, N318, N137);
and AND4 (N328, N322, N150, N110, N89);
nand NAND3 (N329, N274, N203, N182);
buf BUF1 (N330, N325);
xor XOR2 (N331, N328, N103);
and AND4 (N332, N309, N65, N280, N277);
and AND2 (N333, N300, N74);
not NOT1 (N334, N332);
xor XOR2 (N335, N326, N112);
and AND4 (N336, N334, N105, N18, N278);
nand NAND3 (N337, N336, N34, N19);
or OR4 (N338, N333, N314, N285, N44);
nand NAND4 (N339, N331, N58, N291, N88);
buf BUF1 (N340, N335);
nand NAND4 (N341, N320, N245, N310, N310);
not NOT1 (N342, N340);
nand NAND4 (N343, N337, N184, N266, N165);
nor NOR4 (N344, N341, N161, N99, N343);
nand NAND4 (N345, N324, N211, N40, N256);
nand NAND4 (N346, N339, N105, N135, N26);
buf BUF1 (N347, N323);
nand NAND4 (N348, N344, N66, N183, N216);
or OR4 (N349, N317, N215, N179, N152);
and AND4 (N350, N330, N206, N248, N302);
xor XOR2 (N351, N350, N246);
xor XOR2 (N352, N351, N244);
nor NOR4 (N353, N345, N215, N78, N227);
buf BUF1 (N354, N342);
xor XOR2 (N355, N338, N245);
xor XOR2 (N356, N352, N159);
or OR3 (N357, N347, N58, N19);
or OR2 (N358, N356, N313);
and AND4 (N359, N327, N120, N126, N119);
nand NAND3 (N360, N359, N116, N275);
and AND2 (N361, N329, N320);
xor XOR2 (N362, N346, N44);
buf BUF1 (N363, N361);
and AND3 (N364, N360, N77, N88);
nor NOR3 (N365, N358, N193, N322);
and AND3 (N366, N362, N138, N129);
not NOT1 (N367, N355);
xor XOR2 (N368, N357, N152);
or OR4 (N369, N367, N44, N80, N313);
nand NAND2 (N370, N368, N345);
xor XOR2 (N371, N349, N229);
or OR2 (N372, N371, N279);
nor NOR2 (N373, N365, N11);
not NOT1 (N374, N372);
buf BUF1 (N375, N364);
xor XOR2 (N376, N353, N254);
xor XOR2 (N377, N366, N346);
and AND2 (N378, N370, N258);
nor NOR4 (N379, N373, N13, N143, N266);
xor XOR2 (N380, N378, N222);
xor XOR2 (N381, N354, N1);
not NOT1 (N382, N375);
or OR3 (N383, N380, N173, N343);
or OR3 (N384, N381, N379, N103);
or OR2 (N385, N46, N280);
and AND2 (N386, N383, N173);
or OR2 (N387, N376, N38);
nor NOR2 (N388, N348, N102);
xor XOR2 (N389, N388, N198);
not NOT1 (N390, N385);
nand NAND3 (N391, N377, N137, N66);
nor NOR4 (N392, N369, N282, N36, N295);
xor XOR2 (N393, N386, N303);
or OR2 (N394, N389, N310);
not NOT1 (N395, N392);
nand NAND3 (N396, N395, N315, N120);
nand NAND2 (N397, N391, N242);
nor NOR2 (N398, N393, N30);
and AND2 (N399, N374, N224);
nor NOR4 (N400, N387, N193, N204, N5);
nor NOR4 (N401, N396, N7, N183, N70);
nor NOR3 (N402, N398, N366, N40);
xor XOR2 (N403, N397, N139);
nand NAND3 (N404, N401, N60, N99);
xor XOR2 (N405, N384, N106);
and AND4 (N406, N399, N154, N246, N18);
or OR2 (N407, N403, N173);
not NOT1 (N408, N363);
and AND4 (N409, N400, N37, N125, N23);
xor XOR2 (N410, N409, N333);
not NOT1 (N411, N390);
nor NOR4 (N412, N405, N396, N306, N87);
not NOT1 (N413, N404);
nor NOR2 (N414, N412, N234);
nand NAND3 (N415, N411, N246, N117);
nand NAND2 (N416, N410, N23);
not NOT1 (N417, N382);
and AND3 (N418, N413, N38, N53);
buf BUF1 (N419, N418);
and AND2 (N420, N415, N355);
buf BUF1 (N421, N402);
nor NOR4 (N422, N419, N43, N23, N406);
xor XOR2 (N423, N194, N386);
not NOT1 (N424, N416);
nand NAND3 (N425, N423, N268, N74);
buf BUF1 (N426, N414);
nand NAND3 (N427, N394, N414, N366);
nor NOR2 (N428, N424, N336);
nand NAND2 (N429, N420, N412);
or OR3 (N430, N428, N409, N220);
or OR2 (N431, N425, N219);
not NOT1 (N432, N417);
or OR4 (N433, N430, N292, N24, N57);
nor NOR2 (N434, N427, N432);
xor XOR2 (N435, N113, N409);
and AND4 (N436, N433, N336, N271, N290);
nand NAND4 (N437, N421, N197, N51, N71);
xor XOR2 (N438, N426, N429);
and AND4 (N439, N189, N161, N32, N198);
or OR4 (N440, N436, N225, N2, N59);
nor NOR2 (N441, N440, N285);
xor XOR2 (N442, N422, N5);
buf BUF1 (N443, N434);
xor XOR2 (N444, N435, N17);
buf BUF1 (N445, N431);
not NOT1 (N446, N443);
xor XOR2 (N447, N442, N204);
nand NAND2 (N448, N439, N82);
nand NAND3 (N449, N448, N72, N336);
and AND4 (N450, N408, N401, N156, N192);
not NOT1 (N451, N446);
nor NOR3 (N452, N441, N121, N250);
not NOT1 (N453, N449);
and AND2 (N454, N437, N171);
buf BUF1 (N455, N444);
and AND4 (N456, N453, N302, N384, N288);
and AND3 (N457, N455, N249, N356);
and AND4 (N458, N454, N370, N127, N343);
nand NAND3 (N459, N438, N347, N110);
or OR2 (N460, N450, N165);
or OR3 (N461, N458, N436, N63);
or OR2 (N462, N460, N264);
or OR4 (N463, N452, N240, N16, N242);
nor NOR3 (N464, N447, N172, N268);
xor XOR2 (N465, N461, N5);
nor NOR4 (N466, N462, N113, N365, N303);
nand NAND2 (N467, N466, N22);
buf BUF1 (N468, N407);
and AND4 (N469, N457, N314, N237, N417);
nand NAND4 (N470, N469, N435, N67, N222);
not NOT1 (N471, N463);
or OR3 (N472, N471, N326, N265);
or OR4 (N473, N467, N95, N363, N304);
xor XOR2 (N474, N464, N11);
nor NOR2 (N475, N459, N362);
nor NOR3 (N476, N465, N132, N72);
buf BUF1 (N477, N468);
buf BUF1 (N478, N476);
or OR2 (N479, N477, N65);
nand NAND3 (N480, N474, N137, N284);
or OR3 (N481, N479, N171, N138);
or OR2 (N482, N481, N222);
buf BUF1 (N483, N451);
xor XOR2 (N484, N472, N117);
or OR3 (N485, N445, N235, N344);
and AND4 (N486, N484, N305, N219, N411);
xor XOR2 (N487, N470, N403);
buf BUF1 (N488, N478);
not NOT1 (N489, N483);
not NOT1 (N490, N482);
xor XOR2 (N491, N456, N13);
not NOT1 (N492, N491);
and AND2 (N493, N485, N293);
and AND4 (N494, N492, N362, N197, N127);
and AND4 (N495, N494, N402, N490, N81);
xor XOR2 (N496, N22, N83);
nor NOR2 (N497, N480, N2);
nor NOR2 (N498, N497, N366);
not NOT1 (N499, N493);
buf BUF1 (N500, N499);
buf BUF1 (N501, N500);
not NOT1 (N502, N501);
and AND2 (N503, N489, N384);
xor XOR2 (N504, N496, N430);
and AND4 (N505, N486, N169, N108, N356);
xor XOR2 (N506, N487, N178);
nor NOR2 (N507, N506, N262);
nand NAND4 (N508, N498, N385, N46, N348);
not NOT1 (N509, N473);
and AND2 (N510, N509, N123);
or OR4 (N511, N510, N228, N203, N417);
xor XOR2 (N512, N475, N341);
nand NAND2 (N513, N503, N426);
nor NOR4 (N514, N505, N406, N183, N451);
nand NAND2 (N515, N507, N219);
buf BUF1 (N516, N512);
not NOT1 (N517, N513);
and AND2 (N518, N514, N135);
buf BUF1 (N519, N517);
buf BUF1 (N520, N502);
nand NAND3 (N521, N508, N88, N155);
or OR2 (N522, N516, N147);
buf BUF1 (N523, N488);
nor NOR4 (N524, N504, N198, N10, N444);
nand NAND3 (N525, N521, N146, N463);
or OR2 (N526, N495, N28);
or OR3 (N527, N511, N159, N110);
and AND3 (N528, N519, N307, N317);
nand NAND3 (N529, N525, N472, N201);
and AND2 (N530, N515, N252);
not NOT1 (N531, N530);
or OR3 (N532, N523, N118, N332);
nand NAND3 (N533, N529, N443, N326);
not NOT1 (N534, N532);
nor NOR3 (N535, N534, N457, N351);
buf BUF1 (N536, N524);
nand NAND3 (N537, N536, N414, N169);
nand NAND4 (N538, N527, N4, N392, N526);
buf BUF1 (N539, N90);
or OR3 (N540, N535, N225, N44);
xor XOR2 (N541, N533, N329);
and AND3 (N542, N518, N10, N311);
or OR2 (N543, N528, N321);
nor NOR2 (N544, N543, N348);
nand NAND3 (N545, N540, N375, N148);
nor NOR4 (N546, N544, N406, N544, N41);
buf BUF1 (N547, N539);
and AND3 (N548, N541, N426, N130);
not NOT1 (N549, N537);
nand NAND3 (N550, N545, N423, N230);
xor XOR2 (N551, N522, N217);
not NOT1 (N552, N551);
xor XOR2 (N553, N531, N74);
nand NAND4 (N554, N547, N45, N235, N95);
not NOT1 (N555, N550);
nand NAND4 (N556, N554, N288, N323, N511);
xor XOR2 (N557, N553, N253);
buf BUF1 (N558, N538);
or OR2 (N559, N552, N147);
and AND3 (N560, N555, N130, N293);
nand NAND3 (N561, N549, N343, N232);
not NOT1 (N562, N548);
not NOT1 (N563, N559);
nand NAND4 (N564, N558, N203, N70, N450);
buf BUF1 (N565, N564);
nand NAND4 (N566, N556, N77, N378, N384);
buf BUF1 (N567, N566);
nand NAND3 (N568, N542, N196, N324);
nand NAND2 (N569, N560, N43);
or OR4 (N570, N568, N418, N139, N191);
xor XOR2 (N571, N565, N396);
or OR3 (N572, N569, N208, N26);
nand NAND4 (N573, N572, N221, N344, N413);
or OR3 (N574, N561, N118, N157);
not NOT1 (N575, N546);
not NOT1 (N576, N557);
not NOT1 (N577, N576);
nand NAND4 (N578, N520, N422, N339, N188);
and AND2 (N579, N577, N454);
nor NOR3 (N580, N562, N530, N403);
or OR4 (N581, N571, N50, N99, N65);
and AND4 (N582, N579, N155, N57, N513);
xor XOR2 (N583, N573, N274);
and AND4 (N584, N563, N173, N484, N360);
and AND3 (N585, N583, N405, N233);
xor XOR2 (N586, N575, N466);
and AND2 (N587, N574, N559);
nand NAND2 (N588, N567, N405);
buf BUF1 (N589, N587);
nor NOR3 (N590, N582, N325, N291);
not NOT1 (N591, N580);
buf BUF1 (N592, N586);
buf BUF1 (N593, N591);
buf BUF1 (N594, N589);
not NOT1 (N595, N590);
or OR3 (N596, N588, N591, N542);
nor NOR2 (N597, N592, N563);
buf BUF1 (N598, N593);
and AND2 (N599, N585, N290);
and AND3 (N600, N584, N285, N327);
nand NAND4 (N601, N596, N174, N133, N518);
and AND2 (N602, N581, N347);
or OR2 (N603, N600, N186);
nand NAND4 (N604, N601, N434, N43, N170);
or OR3 (N605, N599, N295, N376);
buf BUF1 (N606, N570);
xor XOR2 (N607, N597, N129);
nand NAND3 (N608, N606, N329, N588);
nor NOR4 (N609, N607, N496, N135, N383);
or OR3 (N610, N605, N62, N66);
or OR4 (N611, N604, N98, N584, N581);
nor NOR2 (N612, N608, N608);
xor XOR2 (N613, N612, N440);
buf BUF1 (N614, N611);
buf BUF1 (N615, N609);
xor XOR2 (N616, N602, N491);
xor XOR2 (N617, N578, N190);
nand NAND4 (N618, N610, N244, N407, N400);
and AND4 (N619, N603, N14, N298, N24);
or OR4 (N620, N619, N210, N545, N244);
nand NAND3 (N621, N598, N591, N566);
buf BUF1 (N622, N613);
xor XOR2 (N623, N617, N357);
buf BUF1 (N624, N623);
xor XOR2 (N625, N616, N478);
and AND3 (N626, N622, N314, N561);
nand NAND2 (N627, N595, N22);
and AND4 (N628, N624, N203, N329, N22);
buf BUF1 (N629, N627);
and AND2 (N630, N594, N476);
and AND4 (N631, N618, N437, N234, N444);
not NOT1 (N632, N620);
nand NAND2 (N633, N614, N518);
and AND2 (N634, N621, N527);
nand NAND2 (N635, N615, N163);
or OR4 (N636, N631, N428, N249, N175);
xor XOR2 (N637, N626, N303);
nor NOR2 (N638, N625, N49);
nand NAND4 (N639, N638, N423, N119, N152);
or OR2 (N640, N629, N131);
xor XOR2 (N641, N639, N230);
nand NAND2 (N642, N632, N512);
or OR3 (N643, N634, N189, N512);
and AND3 (N644, N628, N641, N250);
nor NOR3 (N645, N54, N424, N70);
and AND3 (N646, N635, N216, N36);
or OR2 (N647, N630, N194);
not NOT1 (N648, N644);
nor NOR3 (N649, N640, N191, N238);
xor XOR2 (N650, N649, N506);
nor NOR3 (N651, N643, N570, N209);
and AND2 (N652, N646, N321);
xor XOR2 (N653, N652, N168);
nor NOR4 (N654, N642, N433, N320, N553);
nor NOR3 (N655, N636, N381, N70);
nor NOR3 (N656, N651, N565, N84);
and AND4 (N657, N655, N271, N371, N434);
nor NOR2 (N658, N654, N327);
or OR3 (N659, N637, N88, N21);
not NOT1 (N660, N658);
buf BUF1 (N661, N656);
and AND3 (N662, N648, N230, N279);
buf BUF1 (N663, N661);
nor NOR2 (N664, N653, N360);
and AND2 (N665, N657, N615);
buf BUF1 (N666, N663);
nand NAND4 (N667, N660, N375, N358, N125);
nor NOR3 (N668, N666, N48, N617);
or OR3 (N669, N647, N130, N554);
xor XOR2 (N670, N633, N342);
or OR4 (N671, N645, N629, N643, N63);
buf BUF1 (N672, N659);
buf BUF1 (N673, N672);
or OR2 (N674, N662, N32);
not NOT1 (N675, N674);
and AND2 (N676, N664, N108);
and AND2 (N677, N668, N521);
and AND3 (N678, N675, N546, N675);
not NOT1 (N679, N673);
not NOT1 (N680, N670);
buf BUF1 (N681, N669);
buf BUF1 (N682, N667);
or OR4 (N683, N680, N588, N550, N403);
and AND3 (N684, N682, N141, N176);
or OR2 (N685, N683, N407);
nand NAND4 (N686, N676, N455, N331, N217);
and AND2 (N687, N650, N516);
nand NAND2 (N688, N677, N671);
or OR4 (N689, N634, N660, N337, N238);
or OR2 (N690, N679, N547);
or OR4 (N691, N687, N55, N242, N433);
xor XOR2 (N692, N690, N658);
nor NOR3 (N693, N686, N468, N647);
or OR3 (N694, N678, N292, N593);
nand NAND4 (N695, N684, N694, N315, N167);
nand NAND2 (N696, N693, N635);
buf BUF1 (N697, N669);
not NOT1 (N698, N689);
xor XOR2 (N699, N696, N600);
and AND3 (N700, N692, N384, N649);
nand NAND2 (N701, N698, N79);
or OR3 (N702, N701, N413, N689);
nor NOR4 (N703, N665, N488, N598, N330);
nand NAND3 (N704, N699, N178, N376);
nand NAND2 (N705, N703, N201);
xor XOR2 (N706, N691, N665);
not NOT1 (N707, N681);
or OR3 (N708, N700, N376, N510);
and AND4 (N709, N695, N487, N430, N151);
nor NOR3 (N710, N705, N491, N483);
nor NOR4 (N711, N685, N286, N244, N157);
or OR3 (N712, N707, N78, N273);
or OR4 (N713, N697, N664, N710, N577);
buf BUF1 (N714, N350);
and AND2 (N715, N714, N263);
buf BUF1 (N716, N704);
or OR2 (N717, N712, N530);
and AND3 (N718, N688, N715, N112);
buf BUF1 (N719, N18);
not NOT1 (N720, N718);
nand NAND2 (N721, N713, N634);
or OR2 (N722, N720, N146);
xor XOR2 (N723, N719, N465);
nor NOR3 (N724, N717, N401, N582);
not NOT1 (N725, N706);
nand NAND4 (N726, N711, N208, N291, N697);
or OR2 (N727, N702, N228);
or OR4 (N728, N709, N423, N173, N336);
buf BUF1 (N729, N725);
buf BUF1 (N730, N708);
not NOT1 (N731, N726);
not NOT1 (N732, N728);
or OR4 (N733, N727, N269, N366, N211);
and AND3 (N734, N730, N145, N424);
nor NOR3 (N735, N733, N367, N582);
nor NOR3 (N736, N722, N619, N671);
not NOT1 (N737, N716);
xor XOR2 (N738, N731, N123);
xor XOR2 (N739, N734, N488);
nand NAND2 (N740, N721, N559);
and AND2 (N741, N736, N131);
nor NOR4 (N742, N732, N48, N571, N133);
not NOT1 (N743, N723);
not NOT1 (N744, N740);
not NOT1 (N745, N737);
xor XOR2 (N746, N742, N38);
buf BUF1 (N747, N724);
not NOT1 (N748, N745);
not NOT1 (N749, N748);
and AND3 (N750, N735, N139, N484);
not NOT1 (N751, N738);
nand NAND3 (N752, N751, N585, N270);
not NOT1 (N753, N749);
not NOT1 (N754, N744);
nand NAND2 (N755, N746, N85);
and AND3 (N756, N754, N360, N577);
nor NOR2 (N757, N729, N726);
nand NAND2 (N758, N756, N724);
nor NOR2 (N759, N755, N565);
nand NAND4 (N760, N758, N619, N395, N342);
buf BUF1 (N761, N743);
and AND3 (N762, N757, N145, N430);
and AND3 (N763, N739, N305, N593);
or OR4 (N764, N759, N505, N641, N190);
and AND3 (N765, N763, N325, N139);
not NOT1 (N766, N764);
xor XOR2 (N767, N750, N145);
or OR2 (N768, N752, N426);
nand NAND3 (N769, N766, N302, N645);
or OR3 (N770, N769, N522, N574);
buf BUF1 (N771, N770);
or OR4 (N772, N767, N630, N86, N284);
not NOT1 (N773, N741);
buf BUF1 (N774, N747);
and AND2 (N775, N768, N99);
not NOT1 (N776, N771);
or OR2 (N777, N765, N505);
and AND4 (N778, N774, N682, N746, N466);
not NOT1 (N779, N775);
nor NOR2 (N780, N777, N154);
and AND2 (N781, N753, N595);
nand NAND4 (N782, N779, N145, N578, N319);
xor XOR2 (N783, N782, N494);
not NOT1 (N784, N773);
and AND4 (N785, N762, N455, N6, N708);
nand NAND3 (N786, N784, N274, N298);
xor XOR2 (N787, N781, N172);
xor XOR2 (N788, N778, N591);
buf BUF1 (N789, N761);
or OR3 (N790, N783, N506, N334);
buf BUF1 (N791, N780);
nand NAND3 (N792, N785, N169, N736);
buf BUF1 (N793, N786);
nand NAND2 (N794, N792, N106);
nor NOR3 (N795, N789, N261, N750);
buf BUF1 (N796, N794);
buf BUF1 (N797, N796);
xor XOR2 (N798, N776, N617);
buf BUF1 (N799, N787);
not NOT1 (N800, N788);
nor NOR2 (N801, N798, N576);
nand NAND2 (N802, N772, N779);
nor NOR3 (N803, N791, N404, N471);
not NOT1 (N804, N803);
xor XOR2 (N805, N797, N130);
buf BUF1 (N806, N801);
nor NOR3 (N807, N802, N57, N344);
nor NOR4 (N808, N805, N366, N715, N555);
nand NAND3 (N809, N790, N342, N421);
buf BUF1 (N810, N804);
nor NOR3 (N811, N807, N574, N240);
not NOT1 (N812, N760);
and AND2 (N813, N808, N263);
nand NAND4 (N814, N810, N654, N250, N274);
nor NOR4 (N815, N800, N460, N786, N672);
or OR3 (N816, N812, N485, N313);
and AND3 (N817, N793, N428, N429);
not NOT1 (N818, N814);
xor XOR2 (N819, N816, N368);
buf BUF1 (N820, N813);
or OR4 (N821, N818, N626, N147, N392);
buf BUF1 (N822, N817);
and AND2 (N823, N820, N17);
not NOT1 (N824, N815);
endmodule