// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15;

output N712,N682,N708,N706,N707,N713,N709,N703,N697,N715;

not NOT1 (N16, N8);
or OR3 (N17, N15, N1, N8);
xor XOR2 (N18, N11, N6);
nor NOR4 (N19, N14, N4, N1, N10);
nor NOR3 (N20, N1, N14, N15);
xor XOR2 (N21, N5, N16);
nand NAND3 (N22, N7, N5, N17);
nor NOR3 (N23, N22, N20, N9);
xor XOR2 (N24, N19, N15);
or OR3 (N25, N16, N15, N18);
not NOT1 (N26, N14);
nand NAND4 (N27, N1, N5, N22, N4);
or OR4 (N28, N11, N1, N7, N2);
and AND3 (N29, N7, N28, N18);
xor XOR2 (N30, N19, N20);
nor NOR4 (N31, N27, N20, N29, N3);
nor NOR3 (N32, N29, N15, N16);
and AND4 (N33, N23, N4, N10, N11);
or OR4 (N34, N9, N18, N24, N6);
nor NOR4 (N35, N4, N23, N9, N32);
or OR4 (N36, N12, N4, N22, N13);
not NOT1 (N37, N36);
nand NAND2 (N38, N34, N28);
or OR3 (N39, N30, N25, N7);
or OR2 (N40, N13, N36);
nand NAND4 (N41, N25, N11, N12, N2);
nand NAND2 (N42, N31, N36);
or OR2 (N43, N35, N15);
not NOT1 (N44, N38);
and AND2 (N45, N37, N12);
or OR2 (N46, N42, N23);
buf BUF1 (N47, N41);
not NOT1 (N48, N39);
buf BUF1 (N49, N44);
buf BUF1 (N50, N21);
buf BUF1 (N51, N46);
and AND2 (N52, N50, N1);
nand NAND4 (N53, N43, N27, N50, N44);
nor NOR2 (N54, N48, N42);
nor NOR3 (N55, N54, N7, N17);
not NOT1 (N56, N40);
not NOT1 (N57, N47);
and AND4 (N58, N57, N18, N42, N44);
nand NAND4 (N59, N49, N48, N34, N46);
xor XOR2 (N60, N52, N32);
or OR3 (N61, N60, N49, N56);
and AND3 (N62, N29, N14, N48);
or OR4 (N63, N58, N22, N57, N31);
not NOT1 (N64, N59);
xor XOR2 (N65, N26, N44);
not NOT1 (N66, N64);
buf BUF1 (N67, N51);
nand NAND2 (N68, N67, N6);
buf BUF1 (N69, N55);
nor NOR3 (N70, N69, N37, N45);
not NOT1 (N71, N30);
nand NAND4 (N72, N65, N30, N34, N15);
not NOT1 (N73, N62);
or OR2 (N74, N71, N38);
and AND4 (N75, N61, N4, N8, N11);
not NOT1 (N76, N75);
nand NAND3 (N77, N70, N48, N65);
buf BUF1 (N78, N63);
buf BUF1 (N79, N77);
or OR3 (N80, N33, N61, N12);
not NOT1 (N81, N73);
and AND2 (N82, N76, N7);
nor NOR4 (N83, N78, N53, N51, N49);
not NOT1 (N84, N59);
xor XOR2 (N85, N81, N45);
xor XOR2 (N86, N74, N18);
nand NAND4 (N87, N82, N78, N66, N36);
buf BUF1 (N88, N58);
or OR2 (N89, N86, N14);
buf BUF1 (N90, N88);
xor XOR2 (N91, N79, N1);
or OR3 (N92, N89, N42, N3);
buf BUF1 (N93, N84);
buf BUF1 (N94, N93);
or OR3 (N95, N87, N7, N76);
nor NOR3 (N96, N68, N82, N43);
and AND3 (N97, N91, N52, N42);
xor XOR2 (N98, N96, N93);
xor XOR2 (N99, N72, N87);
nor NOR2 (N100, N98, N5);
xor XOR2 (N101, N95, N100);
not NOT1 (N102, N83);
not NOT1 (N103, N61);
nor NOR4 (N104, N85, N42, N51, N50);
buf BUF1 (N105, N97);
nor NOR2 (N106, N90, N2);
or OR2 (N107, N105, N106);
xor XOR2 (N108, N62, N48);
or OR2 (N109, N108, N103);
xor XOR2 (N110, N35, N45);
or OR3 (N111, N109, N15, N74);
nand NAND3 (N112, N80, N75, N20);
not NOT1 (N113, N102);
buf BUF1 (N114, N101);
and AND3 (N115, N99, N76, N106);
or OR4 (N116, N115, N9, N47, N43);
or OR2 (N117, N111, N26);
and AND4 (N118, N107, N113, N55, N32);
or OR3 (N119, N102, N32, N93);
xor XOR2 (N120, N117, N4);
or OR2 (N121, N119, N72);
buf BUF1 (N122, N114);
not NOT1 (N123, N92);
nor NOR2 (N124, N104, N91);
nand NAND2 (N125, N122, N66);
buf BUF1 (N126, N120);
nor NOR2 (N127, N121, N66);
and AND4 (N128, N125, N58, N22, N82);
not NOT1 (N129, N126);
or OR4 (N130, N128, N105, N42, N19);
nand NAND4 (N131, N130, N57, N78, N78);
nor NOR2 (N132, N129, N59);
nor NOR2 (N133, N123, N118);
buf BUF1 (N134, N30);
buf BUF1 (N135, N134);
or OR3 (N136, N133, N126, N109);
not NOT1 (N137, N110);
nand NAND4 (N138, N136, N5, N103, N5);
or OR2 (N139, N132, N100);
nand NAND4 (N140, N135, N15, N20, N29);
buf BUF1 (N141, N124);
nand NAND2 (N142, N138, N43);
nand NAND4 (N143, N140, N31, N43, N40);
and AND4 (N144, N127, N83, N56, N106);
buf BUF1 (N145, N142);
xor XOR2 (N146, N143, N123);
not NOT1 (N147, N116);
xor XOR2 (N148, N145, N46);
or OR3 (N149, N94, N75, N85);
nor NOR2 (N150, N147, N101);
buf BUF1 (N151, N141);
and AND2 (N152, N151, N43);
and AND4 (N153, N146, N63, N114, N43);
and AND3 (N154, N137, N21, N30);
nor NOR4 (N155, N152, N58, N33, N9);
buf BUF1 (N156, N154);
buf BUF1 (N157, N148);
buf BUF1 (N158, N139);
nand NAND3 (N159, N158, N13, N12);
nor NOR2 (N160, N131, N149);
nand NAND4 (N161, N127, N105, N126, N52);
not NOT1 (N162, N161);
nor NOR3 (N163, N153, N8, N135);
nor NOR4 (N164, N157, N117, N102, N20);
buf BUF1 (N165, N156);
and AND4 (N166, N150, N152, N114, N90);
xor XOR2 (N167, N165, N80);
nor NOR4 (N168, N112, N140, N145, N76);
nor NOR3 (N169, N167, N66, N71);
and AND4 (N170, N164, N128, N110, N22);
nand NAND4 (N171, N170, N43, N41, N77);
nand NAND2 (N172, N159, N23);
or OR4 (N173, N169, N17, N55, N71);
buf BUF1 (N174, N144);
and AND4 (N175, N171, N80, N33, N148);
or OR2 (N176, N175, N88);
nand NAND2 (N177, N168, N92);
not NOT1 (N178, N155);
not NOT1 (N179, N177);
buf BUF1 (N180, N172);
not NOT1 (N181, N160);
xor XOR2 (N182, N166, N91);
nor NOR4 (N183, N176, N111, N26, N83);
or OR3 (N184, N173, N75, N159);
not NOT1 (N185, N182);
buf BUF1 (N186, N185);
and AND2 (N187, N178, N65);
xor XOR2 (N188, N180, N176);
and AND3 (N189, N184, N150, N155);
nor NOR2 (N190, N189, N103);
and AND4 (N191, N162, N162, N9, N98);
nor NOR2 (N192, N187, N44);
nand NAND4 (N193, N191, N59, N80, N80);
nor NOR2 (N194, N186, N10);
not NOT1 (N195, N194);
xor XOR2 (N196, N192, N86);
not NOT1 (N197, N190);
nand NAND2 (N198, N179, N68);
or OR3 (N199, N174, N24, N72);
nor NOR4 (N200, N197, N104, N174, N160);
not NOT1 (N201, N195);
nor NOR3 (N202, N199, N189, N50);
and AND4 (N203, N198, N85, N3, N74);
nand NAND2 (N204, N196, N194);
buf BUF1 (N205, N201);
not NOT1 (N206, N163);
nor NOR4 (N207, N203, N153, N56, N88);
nand NAND3 (N208, N202, N76, N174);
not NOT1 (N209, N206);
nand NAND3 (N210, N204, N77, N26);
not NOT1 (N211, N208);
or OR2 (N212, N210, N65);
nor NOR3 (N213, N181, N139, N128);
and AND2 (N214, N212, N68);
nor NOR3 (N215, N213, N107, N171);
not NOT1 (N216, N200);
not NOT1 (N217, N211);
and AND4 (N218, N209, N103, N196, N81);
not NOT1 (N219, N188);
nor NOR3 (N220, N215, N107, N24);
not NOT1 (N221, N217);
buf BUF1 (N222, N193);
buf BUF1 (N223, N214);
or OR2 (N224, N220, N174);
and AND2 (N225, N207, N59);
buf BUF1 (N226, N218);
nor NOR3 (N227, N205, N101, N63);
and AND3 (N228, N222, N113, N115);
buf BUF1 (N229, N183);
xor XOR2 (N230, N226, N182);
nand NAND2 (N231, N224, N15);
and AND3 (N232, N221, N50, N56);
or OR3 (N233, N228, N58, N21);
xor XOR2 (N234, N216, N196);
nand NAND2 (N235, N223, N131);
not NOT1 (N236, N231);
or OR3 (N237, N227, N151, N184);
nor NOR4 (N238, N236, N179, N123, N168);
and AND3 (N239, N238, N154, N140);
not NOT1 (N240, N237);
not NOT1 (N241, N235);
nor NOR3 (N242, N230, N134, N165);
not NOT1 (N243, N219);
xor XOR2 (N244, N243, N172);
and AND3 (N245, N239, N48, N21);
or OR4 (N246, N232, N130, N200, N188);
nand NAND4 (N247, N233, N61, N178, N17);
buf BUF1 (N248, N246);
not NOT1 (N249, N234);
nand NAND4 (N250, N244, N66, N181, N74);
nor NOR4 (N251, N240, N58, N187, N87);
nand NAND4 (N252, N225, N205, N183, N42);
xor XOR2 (N253, N229, N213);
buf BUF1 (N254, N248);
nand NAND2 (N255, N249, N193);
nand NAND3 (N256, N254, N125, N17);
buf BUF1 (N257, N245);
xor XOR2 (N258, N255, N42);
nand NAND3 (N259, N247, N161, N240);
nand NAND2 (N260, N253, N96);
buf BUF1 (N261, N260);
not NOT1 (N262, N258);
nand NAND2 (N263, N242, N161);
and AND2 (N264, N259, N152);
nor NOR4 (N265, N251, N56, N112, N5);
nor NOR4 (N266, N264, N4, N60, N255);
xor XOR2 (N267, N250, N192);
and AND3 (N268, N262, N226, N64);
not NOT1 (N269, N263);
not NOT1 (N270, N256);
nand NAND2 (N271, N252, N193);
nor NOR3 (N272, N266, N93, N20);
nor NOR4 (N273, N265, N101, N104, N189);
not NOT1 (N274, N268);
nor NOR3 (N275, N272, N201, N167);
or OR4 (N276, N267, N241, N46, N81);
or OR3 (N277, N163, N73, N212);
nand NAND4 (N278, N271, N148, N194, N263);
or OR3 (N279, N270, N21, N1);
nor NOR4 (N280, N261, N199, N202, N270);
or OR4 (N281, N257, N266, N241, N100);
buf BUF1 (N282, N275);
xor XOR2 (N283, N282, N173);
nor NOR2 (N284, N281, N274);
nor NOR3 (N285, N185, N56, N200);
xor XOR2 (N286, N283, N178);
or OR2 (N287, N284, N197);
or OR3 (N288, N280, N65, N276);
buf BUF1 (N289, N133);
not NOT1 (N290, N279);
or OR2 (N291, N289, N251);
and AND4 (N292, N269, N224, N118, N147);
buf BUF1 (N293, N286);
nor NOR2 (N294, N287, N292);
and AND2 (N295, N170, N156);
and AND3 (N296, N278, N4, N26);
and AND3 (N297, N293, N82, N176);
nor NOR4 (N298, N291, N97, N239, N28);
nor NOR2 (N299, N294, N97);
not NOT1 (N300, N273);
xor XOR2 (N301, N299, N272);
buf BUF1 (N302, N297);
nand NAND2 (N303, N285, N173);
and AND3 (N304, N298, N12, N59);
not NOT1 (N305, N302);
or OR3 (N306, N296, N117, N4);
or OR3 (N307, N290, N139, N94);
not NOT1 (N308, N307);
not NOT1 (N309, N308);
or OR2 (N310, N306, N229);
nor NOR4 (N311, N301, N29, N219, N52);
not NOT1 (N312, N277);
or OR4 (N313, N300, N281, N191, N87);
nor NOR2 (N314, N295, N7);
buf BUF1 (N315, N303);
xor XOR2 (N316, N305, N25);
nor NOR4 (N317, N311, N124, N73, N270);
and AND3 (N318, N315, N212, N129);
xor XOR2 (N319, N317, N213);
or OR2 (N320, N309, N201);
nand NAND4 (N321, N313, N249, N115, N243);
not NOT1 (N322, N314);
buf BUF1 (N323, N318);
or OR3 (N324, N323, N112, N251);
and AND3 (N325, N316, N307, N235);
or OR3 (N326, N319, N81, N199);
nand NAND2 (N327, N320, N118);
not NOT1 (N328, N304);
or OR4 (N329, N310, N188, N202, N179);
not NOT1 (N330, N321);
nor NOR4 (N331, N312, N80, N71, N295);
nand NAND2 (N332, N330, N137);
and AND3 (N333, N329, N80, N153);
not NOT1 (N334, N328);
not NOT1 (N335, N326);
nand NAND3 (N336, N334, N175, N90);
and AND3 (N337, N335, N187, N163);
nor NOR2 (N338, N333, N142);
xor XOR2 (N339, N337, N8);
nor NOR2 (N340, N331, N171);
and AND2 (N341, N325, N91);
xor XOR2 (N342, N288, N156);
nand NAND4 (N343, N339, N201, N147, N125);
buf BUF1 (N344, N332);
buf BUF1 (N345, N338);
not NOT1 (N346, N322);
not NOT1 (N347, N345);
not NOT1 (N348, N344);
xor XOR2 (N349, N346, N188);
not NOT1 (N350, N324);
nand NAND4 (N351, N341, N83, N78, N127);
buf BUF1 (N352, N336);
or OR3 (N353, N348, N137, N58);
xor XOR2 (N354, N352, N249);
nand NAND4 (N355, N340, N175, N325, N192);
nand NAND3 (N356, N351, N2, N189);
xor XOR2 (N357, N356, N48);
nor NOR4 (N358, N327, N259, N283, N285);
nor NOR3 (N359, N349, N190, N340);
nor NOR4 (N360, N350, N136, N112, N36);
and AND4 (N361, N358, N160, N151, N49);
or OR2 (N362, N343, N37);
or OR3 (N363, N362, N305, N205);
nand NAND3 (N364, N360, N211, N251);
buf BUF1 (N365, N364);
nor NOR3 (N366, N363, N18, N77);
and AND4 (N367, N342, N258, N271, N77);
and AND3 (N368, N367, N104, N191);
and AND3 (N369, N361, N45, N160);
not NOT1 (N370, N369);
nor NOR4 (N371, N368, N49, N201, N94);
and AND2 (N372, N357, N275);
nor NOR4 (N373, N366, N64, N251, N15);
buf BUF1 (N374, N370);
xor XOR2 (N375, N373, N162);
or OR2 (N376, N374, N85);
and AND3 (N377, N376, N129, N65);
nand NAND3 (N378, N359, N125, N214);
or OR4 (N379, N354, N332, N209, N244);
buf BUF1 (N380, N372);
xor XOR2 (N381, N377, N243);
and AND4 (N382, N371, N163, N177, N371);
not NOT1 (N383, N353);
xor XOR2 (N384, N381, N359);
buf BUF1 (N385, N347);
nor NOR3 (N386, N375, N337, N41);
nor NOR3 (N387, N379, N157, N298);
xor XOR2 (N388, N382, N186);
nor NOR2 (N389, N385, N104);
and AND3 (N390, N355, N22, N217);
nand NAND2 (N391, N388, N22);
and AND3 (N392, N389, N216, N96);
buf BUF1 (N393, N391);
nor NOR4 (N394, N365, N330, N143, N136);
buf BUF1 (N395, N390);
not NOT1 (N396, N383);
or OR2 (N397, N396, N77);
or OR2 (N398, N384, N106);
not NOT1 (N399, N392);
nand NAND2 (N400, N393, N317);
not NOT1 (N401, N386);
and AND3 (N402, N399, N104, N349);
nor NOR3 (N403, N387, N365, N182);
xor XOR2 (N404, N400, N300);
nor NOR3 (N405, N378, N130, N311);
or OR3 (N406, N394, N345, N265);
xor XOR2 (N407, N395, N41);
or OR3 (N408, N402, N324, N269);
nand NAND2 (N409, N397, N7);
buf BUF1 (N410, N407);
not NOT1 (N411, N410);
or OR2 (N412, N406, N69);
and AND2 (N413, N405, N263);
nand NAND3 (N414, N413, N80, N319);
and AND4 (N415, N412, N63, N364, N66);
nor NOR3 (N416, N403, N120, N187);
not NOT1 (N417, N380);
nand NAND4 (N418, N411, N106, N55, N371);
or OR2 (N419, N408, N256);
and AND3 (N420, N415, N52, N35);
nand NAND4 (N421, N414, N56, N420, N360);
and AND3 (N422, N61, N128, N108);
not NOT1 (N423, N404);
nand NAND3 (N424, N416, N341, N65);
and AND4 (N425, N398, N105, N140, N3);
or OR4 (N426, N409, N309, N385, N220);
or OR3 (N427, N421, N349, N200);
buf BUF1 (N428, N423);
nand NAND2 (N429, N419, N204);
nand NAND3 (N430, N422, N383, N20);
nand NAND3 (N431, N425, N131, N396);
and AND4 (N432, N427, N223, N333, N23);
or OR3 (N433, N429, N270, N90);
xor XOR2 (N434, N433, N76);
and AND2 (N435, N426, N277);
or OR2 (N436, N431, N205);
or OR4 (N437, N434, N250, N302, N125);
nand NAND2 (N438, N401, N15);
and AND4 (N439, N418, N282, N235, N47);
nor NOR2 (N440, N436, N229);
not NOT1 (N441, N424);
xor XOR2 (N442, N428, N122);
or OR2 (N443, N417, N90);
buf BUF1 (N444, N443);
not NOT1 (N445, N432);
nand NAND2 (N446, N442, N153);
xor XOR2 (N447, N437, N257);
nand NAND4 (N448, N435, N290, N127, N163);
not NOT1 (N449, N441);
and AND4 (N450, N440, N438, N423, N400);
not NOT1 (N451, N380);
nor NOR4 (N452, N447, N330, N146, N340);
buf BUF1 (N453, N446);
or OR4 (N454, N451, N253, N81, N219);
xor XOR2 (N455, N448, N362);
or OR4 (N456, N453, N25, N157, N386);
and AND3 (N457, N449, N210, N444);
nand NAND2 (N458, N173, N13);
xor XOR2 (N459, N458, N268);
xor XOR2 (N460, N450, N205);
not NOT1 (N461, N455);
xor XOR2 (N462, N459, N356);
nand NAND4 (N463, N430, N115, N319, N411);
not NOT1 (N464, N462);
not NOT1 (N465, N452);
nor NOR4 (N466, N463, N297, N267, N44);
xor XOR2 (N467, N445, N237);
nand NAND3 (N468, N457, N346, N63);
buf BUF1 (N469, N465);
xor XOR2 (N470, N460, N248);
and AND4 (N471, N439, N398, N232, N43);
buf BUF1 (N472, N471);
buf BUF1 (N473, N464);
nand NAND2 (N474, N472, N318);
nor NOR3 (N475, N470, N388, N138);
or OR4 (N476, N461, N320, N48, N372);
or OR4 (N477, N468, N382, N329, N246);
xor XOR2 (N478, N454, N82);
or OR3 (N479, N466, N217, N277);
or OR2 (N480, N475, N272);
and AND2 (N481, N476, N470);
nor NOR2 (N482, N474, N20);
buf BUF1 (N483, N482);
not NOT1 (N484, N478);
nand NAND3 (N485, N481, N240, N357);
nand NAND2 (N486, N467, N430);
buf BUF1 (N487, N486);
nand NAND4 (N488, N479, N185, N367, N360);
or OR4 (N489, N484, N147, N210, N52);
and AND2 (N490, N480, N338);
nor NOR3 (N491, N488, N52, N71);
not NOT1 (N492, N490);
xor XOR2 (N493, N491, N474);
xor XOR2 (N494, N485, N147);
or OR4 (N495, N456, N133, N44, N145);
nand NAND3 (N496, N469, N282, N119);
buf BUF1 (N497, N494);
not NOT1 (N498, N493);
nand NAND4 (N499, N477, N23, N458, N327);
buf BUF1 (N500, N495);
nor NOR3 (N501, N487, N392, N201);
xor XOR2 (N502, N492, N147);
or OR2 (N503, N496, N96);
nand NAND3 (N504, N501, N61, N6);
nor NOR4 (N505, N500, N67, N313, N78);
buf BUF1 (N506, N504);
not NOT1 (N507, N473);
and AND4 (N508, N502, N25, N479, N229);
buf BUF1 (N509, N489);
nand NAND3 (N510, N507, N480, N359);
nor NOR3 (N511, N503, N14, N479);
nand NAND4 (N512, N509, N271, N384, N126);
buf BUF1 (N513, N511);
and AND2 (N514, N512, N195);
xor XOR2 (N515, N510, N261);
nor NOR4 (N516, N498, N212, N221, N87);
not NOT1 (N517, N515);
or OR4 (N518, N506, N365, N458, N126);
or OR3 (N519, N514, N271, N434);
xor XOR2 (N520, N519, N272);
or OR2 (N521, N508, N94);
or OR2 (N522, N521, N426);
buf BUF1 (N523, N483);
and AND2 (N524, N523, N339);
nand NAND3 (N525, N516, N311, N264);
not NOT1 (N526, N520);
or OR4 (N527, N525, N428, N48, N235);
xor XOR2 (N528, N524, N351);
buf BUF1 (N529, N518);
not NOT1 (N530, N497);
and AND3 (N531, N529, N422, N384);
not NOT1 (N532, N530);
nor NOR2 (N533, N527, N191);
or OR3 (N534, N528, N249, N286);
not NOT1 (N535, N531);
not NOT1 (N536, N517);
and AND3 (N537, N522, N207, N75);
buf BUF1 (N538, N537);
and AND4 (N539, N534, N413, N128, N217);
nand NAND3 (N540, N536, N379, N279);
nand NAND2 (N541, N535, N367);
and AND4 (N542, N540, N345, N495, N477);
and AND2 (N543, N513, N282);
not NOT1 (N544, N543);
xor XOR2 (N545, N505, N104);
not NOT1 (N546, N499);
not NOT1 (N547, N544);
nor NOR4 (N548, N545, N540, N85, N361);
buf BUF1 (N549, N526);
not NOT1 (N550, N548);
and AND3 (N551, N541, N147, N257);
nor NOR3 (N552, N532, N506, N201);
xor XOR2 (N553, N533, N518);
xor XOR2 (N554, N547, N413);
buf BUF1 (N555, N551);
nand NAND3 (N556, N554, N154, N2);
not NOT1 (N557, N556);
buf BUF1 (N558, N546);
or OR2 (N559, N538, N394);
or OR3 (N560, N558, N527, N465);
xor XOR2 (N561, N550, N366);
not NOT1 (N562, N555);
not NOT1 (N563, N557);
xor XOR2 (N564, N559, N146);
not NOT1 (N565, N563);
not NOT1 (N566, N560);
buf BUF1 (N567, N552);
not NOT1 (N568, N549);
xor XOR2 (N569, N561, N168);
not NOT1 (N570, N539);
nor NOR2 (N571, N562, N481);
or OR2 (N572, N567, N176);
or OR4 (N573, N571, N214, N431, N421);
and AND3 (N574, N572, N41, N82);
not NOT1 (N575, N565);
xor XOR2 (N576, N542, N316);
and AND2 (N577, N553, N66);
and AND4 (N578, N574, N544, N82, N145);
buf BUF1 (N579, N570);
nor NOR3 (N580, N575, N199, N81);
or OR2 (N581, N576, N129);
and AND3 (N582, N573, N417, N580);
nor NOR2 (N583, N361, N282);
not NOT1 (N584, N569);
or OR3 (N585, N583, N423, N339);
nor NOR2 (N586, N579, N371);
nand NAND3 (N587, N578, N563, N582);
buf BUF1 (N588, N402);
and AND3 (N589, N585, N461, N57);
and AND2 (N590, N564, N204);
and AND3 (N591, N586, N60, N141);
not NOT1 (N592, N568);
nand NAND3 (N593, N584, N333, N429);
or OR3 (N594, N591, N194, N71);
nand NAND4 (N595, N588, N543, N426, N464);
nor NOR4 (N596, N566, N241, N182, N586);
nor NOR3 (N597, N587, N141, N323);
xor XOR2 (N598, N592, N373);
and AND2 (N599, N589, N478);
not NOT1 (N600, N595);
and AND2 (N601, N597, N259);
nand NAND2 (N602, N594, N109);
and AND2 (N603, N596, N573);
and AND4 (N604, N600, N127, N42, N15);
nor NOR4 (N605, N598, N600, N147, N314);
xor XOR2 (N606, N601, N414);
xor XOR2 (N607, N606, N464);
nand NAND4 (N608, N607, N219, N412, N489);
not NOT1 (N609, N590);
nor NOR2 (N610, N605, N61);
or OR2 (N611, N602, N450);
nor NOR4 (N612, N608, N225, N300, N588);
and AND2 (N613, N604, N56);
not NOT1 (N614, N613);
xor XOR2 (N615, N599, N595);
nand NAND2 (N616, N609, N181);
buf BUF1 (N617, N593);
not NOT1 (N618, N611);
nor NOR3 (N619, N603, N79, N285);
buf BUF1 (N620, N614);
nor NOR4 (N621, N610, N194, N408, N1);
nand NAND2 (N622, N617, N544);
nand NAND4 (N623, N618, N594, N510, N100);
not NOT1 (N624, N621);
buf BUF1 (N625, N624);
nor NOR2 (N626, N620, N394);
xor XOR2 (N627, N612, N48);
xor XOR2 (N628, N581, N54);
not NOT1 (N629, N625);
or OR3 (N630, N629, N151, N419);
nand NAND4 (N631, N628, N487, N4, N126);
buf BUF1 (N632, N622);
and AND3 (N633, N627, N248, N350);
buf BUF1 (N634, N577);
nor NOR3 (N635, N630, N590, N456);
and AND3 (N636, N623, N280, N171);
nor NOR2 (N637, N619, N56);
or OR3 (N638, N634, N444, N636);
buf BUF1 (N639, N319);
xor XOR2 (N640, N638, N105);
or OR3 (N641, N631, N376, N259);
xor XOR2 (N642, N640, N584);
and AND3 (N643, N639, N385, N530);
not NOT1 (N644, N643);
nor NOR2 (N645, N641, N39);
and AND3 (N646, N642, N5, N547);
not NOT1 (N647, N615);
nor NOR2 (N648, N633, N441);
buf BUF1 (N649, N632);
not NOT1 (N650, N616);
buf BUF1 (N651, N644);
nand NAND4 (N652, N650, N309, N497, N388);
nor NOR3 (N653, N635, N79, N484);
nand NAND3 (N654, N651, N100, N376);
and AND3 (N655, N653, N457, N219);
and AND4 (N656, N652, N406, N156, N81);
xor XOR2 (N657, N656, N196);
not NOT1 (N658, N646);
nor NOR4 (N659, N637, N554, N295, N565);
not NOT1 (N660, N654);
not NOT1 (N661, N659);
nand NAND4 (N662, N658, N525, N557, N9);
or OR4 (N663, N648, N36, N498, N287);
not NOT1 (N664, N657);
and AND3 (N665, N663, N571, N398);
or OR3 (N666, N655, N646, N637);
nor NOR3 (N667, N664, N60, N256);
buf BUF1 (N668, N660);
buf BUF1 (N669, N645);
not NOT1 (N670, N665);
or OR2 (N671, N661, N403);
nor NOR2 (N672, N662, N263);
xor XOR2 (N673, N666, N551);
and AND4 (N674, N649, N266, N253, N353);
and AND2 (N675, N647, N224);
buf BUF1 (N676, N674);
nor NOR3 (N677, N626, N434, N527);
and AND4 (N678, N672, N172, N465, N55);
xor XOR2 (N679, N675, N506);
nand NAND4 (N680, N677, N225, N11, N450);
and AND4 (N681, N673, N430, N270, N642);
buf BUF1 (N682, N671);
nand NAND3 (N683, N668, N668, N307);
xor XOR2 (N684, N678, N181);
buf BUF1 (N685, N680);
buf BUF1 (N686, N684);
and AND3 (N687, N667, N386, N483);
nor NOR2 (N688, N681, N456);
nor NOR2 (N689, N676, N174);
and AND4 (N690, N687, N211, N35, N70);
nand NAND4 (N691, N669, N319, N263, N150);
xor XOR2 (N692, N683, N125);
and AND4 (N693, N692, N436, N160, N208);
nor NOR4 (N694, N691, N494, N137, N482);
and AND2 (N695, N694, N125);
not NOT1 (N696, N689);
nor NOR3 (N697, N695, N309, N165);
nand NAND4 (N698, N686, N201, N276, N299);
nor NOR3 (N699, N693, N458, N650);
buf BUF1 (N700, N679);
not NOT1 (N701, N698);
or OR3 (N702, N688, N103, N46);
nor NOR2 (N703, N701, N89);
and AND2 (N704, N702, N103);
nor NOR2 (N705, N699, N469);
not NOT1 (N706, N696);
buf BUF1 (N707, N685);
or OR2 (N708, N704, N177);
not NOT1 (N709, N700);
buf BUF1 (N710, N705);
not NOT1 (N711, N670);
and AND2 (N712, N690, N194);
nand NAND2 (N713, N710, N639);
xor XOR2 (N714, N711, N24);
not NOT1 (N715, N714);
endmodule