// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19;

output N116,N103,N95,N118,N107,N108,N106,N99,N104,N119;

buf BUF1 (N20, N19);
not NOT1 (N21, N7);
not NOT1 (N22, N9);
or OR2 (N23, N8, N7);
and AND4 (N24, N12, N5, N15, N7);
nand NAND4 (N25, N14, N16, N15, N22);
or OR2 (N26, N12, N14);
nand NAND4 (N27, N18, N13, N1, N15);
or OR4 (N28, N15, N15, N12, N1);
buf BUF1 (N29, N20);
xor XOR2 (N30, N26, N22);
and AND2 (N31, N6, N4);
nand NAND4 (N32, N22, N13, N10, N12);
not NOT1 (N33, N25);
buf BUF1 (N34, N23);
or OR2 (N35, N30, N32);
nand NAND4 (N36, N20, N9, N32, N35);
xor XOR2 (N37, N2, N19);
and AND4 (N38, N34, N21, N4, N10);
nor NOR2 (N39, N16, N31);
nand NAND3 (N40, N28, N13, N15);
buf BUF1 (N41, N9);
and AND3 (N42, N39, N3, N4);
nor NOR2 (N43, N29, N40);
nor NOR3 (N44, N31, N19, N29);
and AND2 (N45, N24, N4);
and AND3 (N46, N43, N35, N6);
nor NOR3 (N47, N41, N38, N2);
buf BUF1 (N48, N16);
buf BUF1 (N49, N46);
nand NAND2 (N50, N42, N40);
and AND4 (N51, N48, N28, N21, N37);
xor XOR2 (N52, N18, N10);
or OR2 (N53, N51, N34);
not NOT1 (N54, N44);
nor NOR4 (N55, N50, N40, N11, N6);
nor NOR3 (N56, N52, N6, N6);
and AND2 (N57, N56, N43);
xor XOR2 (N58, N49, N57);
and AND2 (N59, N5, N7);
and AND3 (N60, N54, N54, N26);
not NOT1 (N61, N59);
not NOT1 (N62, N45);
nand NAND3 (N63, N36, N16, N54);
and AND4 (N64, N55, N61, N48, N35);
buf BUF1 (N65, N4);
not NOT1 (N66, N64);
and AND2 (N67, N27, N44);
nor NOR4 (N68, N66, N26, N22, N67);
or OR4 (N69, N34, N36, N12, N62);
buf BUF1 (N70, N47);
xor XOR2 (N71, N58, N44);
xor XOR2 (N72, N32, N38);
buf BUF1 (N73, N70);
buf BUF1 (N74, N72);
or OR3 (N75, N69, N22, N46);
xor XOR2 (N76, N71, N26);
not NOT1 (N77, N76);
xor XOR2 (N78, N73, N35);
and AND2 (N79, N68, N31);
nor NOR4 (N80, N79, N30, N39, N41);
xor XOR2 (N81, N53, N70);
buf BUF1 (N82, N75);
nand NAND2 (N83, N33, N15);
or OR4 (N84, N63, N35, N74, N1);
nand NAND3 (N85, N50, N36, N17);
or OR3 (N86, N81, N75, N68);
nor NOR3 (N87, N85, N35, N46);
xor XOR2 (N88, N77, N51);
buf BUF1 (N89, N65);
xor XOR2 (N90, N83, N64);
and AND3 (N91, N78, N25, N43);
nand NAND2 (N92, N80, N63);
or OR2 (N93, N84, N72);
and AND2 (N94, N89, N48);
or OR4 (N95, N93, N89, N48, N88);
or OR2 (N96, N4, N28);
xor XOR2 (N97, N92, N37);
and AND2 (N98, N96, N65);
and AND2 (N99, N90, N87);
xor XOR2 (N100, N89, N18);
nor NOR3 (N101, N98, N94, N5);
xor XOR2 (N102, N90, N26);
xor XOR2 (N103, N86, N59);
nand NAND4 (N104, N91, N10, N19, N6);
nor NOR4 (N105, N101, N60, N56, N41);
xor XOR2 (N106, N48, N44);
nor NOR2 (N107, N100, N42);
xor XOR2 (N108, N102, N96);
nor NOR2 (N109, N105, N32);
not NOT1 (N110, N109);
not NOT1 (N111, N97);
buf BUF1 (N112, N110);
or OR4 (N113, N82, N67, N87, N14);
buf BUF1 (N114, N112);
or OR4 (N115, N114, N63, N94, N52);
nand NAND3 (N116, N115, N7, N66);
and AND2 (N117, N113, N105);
buf BUF1 (N118, N111);
buf BUF1 (N119, N117);
endmodule