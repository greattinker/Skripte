// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17;

output N16009,N16011,N16015,N15982,N16014,N16016,N16003,N16006,N16007,N16017;

not NOT1 (N18, N10);
nand NAND2 (N19, N16, N15);
and AND4 (N20, N2, N18, N5, N6);
not NOT1 (N21, N9);
or OR4 (N22, N15, N5, N18, N8);
xor XOR2 (N23, N20, N16);
and AND3 (N24, N12, N6, N5);
or OR2 (N25, N10, N8);
nor NOR4 (N26, N4, N7, N7, N23);
nand NAND2 (N27, N16, N20);
and AND3 (N28, N3, N25, N18);
not NOT1 (N29, N18);
xor XOR2 (N30, N25, N26);
xor XOR2 (N31, N8, N17);
xor XOR2 (N32, N10, N8);
xor XOR2 (N33, N27, N15);
or OR3 (N34, N21, N16, N26);
not NOT1 (N35, N31);
nor NOR2 (N36, N35, N17);
and AND2 (N37, N29, N6);
nor NOR4 (N38, N36, N7, N28, N14);
nor NOR3 (N39, N26, N6, N25);
nor NOR3 (N40, N22, N19, N21);
buf BUF1 (N41, N15);
nand NAND2 (N42, N41, N14);
xor XOR2 (N43, N33, N42);
buf BUF1 (N44, N35);
xor XOR2 (N45, N32, N41);
nor NOR3 (N46, N38, N24, N28);
or OR2 (N47, N14, N17);
xor XOR2 (N48, N39, N45);
or OR4 (N49, N32, N39, N21, N36);
xor XOR2 (N50, N30, N1);
nor NOR3 (N51, N34, N16, N37);
or OR3 (N52, N33, N5, N38);
nor NOR4 (N53, N40, N25, N13, N11);
and AND4 (N54, N50, N38, N29, N21);
and AND3 (N55, N43, N42, N2);
buf BUF1 (N56, N55);
and AND2 (N57, N52, N56);
xor XOR2 (N58, N6, N32);
not NOT1 (N59, N57);
xor XOR2 (N60, N46, N32);
not NOT1 (N61, N48);
nor NOR3 (N62, N44, N19, N59);
nor NOR4 (N63, N26, N62, N41, N1);
and AND2 (N64, N53, N2);
xor XOR2 (N65, N18, N26);
buf BUF1 (N66, N47);
buf BUF1 (N67, N63);
or OR4 (N68, N67, N39, N23, N55);
nor NOR2 (N69, N49, N1);
nor NOR4 (N70, N64, N54, N21, N67);
buf BUF1 (N71, N57);
not NOT1 (N72, N61);
or OR4 (N73, N58, N51, N36, N36);
not NOT1 (N74, N41);
not NOT1 (N75, N69);
not NOT1 (N76, N66);
not NOT1 (N77, N74);
and AND2 (N78, N70, N31);
nor NOR2 (N79, N60, N54);
not NOT1 (N80, N65);
xor XOR2 (N81, N75, N58);
nor NOR2 (N82, N81, N34);
and AND2 (N83, N73, N17);
xor XOR2 (N84, N83, N22);
or OR3 (N85, N80, N83, N60);
not NOT1 (N86, N82);
nand NAND2 (N87, N76, N34);
or OR4 (N88, N72, N25, N65, N82);
or OR3 (N89, N86, N28, N16);
not NOT1 (N90, N87);
buf BUF1 (N91, N79);
not NOT1 (N92, N71);
and AND4 (N93, N92, N48, N75, N87);
nor NOR4 (N94, N85, N23, N4, N65);
not NOT1 (N95, N93);
xor XOR2 (N96, N77, N65);
xor XOR2 (N97, N88, N6);
or OR3 (N98, N84, N63, N83);
nor NOR4 (N99, N96, N41, N49, N3);
and AND2 (N100, N89, N87);
buf BUF1 (N101, N68);
not NOT1 (N102, N100);
nand NAND3 (N103, N99, N53, N37);
nand NAND3 (N104, N97, N43, N40);
or OR4 (N105, N104, N104, N49, N33);
buf BUF1 (N106, N91);
nor NOR3 (N107, N106, N8, N72);
nor NOR4 (N108, N78, N99, N82, N74);
and AND4 (N109, N108, N74, N86, N108);
buf BUF1 (N110, N109);
and AND2 (N111, N95, N103);
nand NAND3 (N112, N58, N33, N36);
nor NOR4 (N113, N101, N13, N15, N81);
not NOT1 (N114, N102);
or OR4 (N115, N114, N80, N37, N24);
nand NAND4 (N116, N110, N59, N55, N73);
nor NOR4 (N117, N115, N105, N101, N18);
nand NAND2 (N118, N110, N4);
and AND3 (N119, N107, N38, N1);
buf BUF1 (N120, N113);
buf BUF1 (N121, N94);
and AND2 (N122, N112, N16);
or OR3 (N123, N120, N59, N108);
and AND2 (N124, N98, N71);
not NOT1 (N125, N123);
or OR2 (N126, N117, N57);
xor XOR2 (N127, N124, N51);
and AND4 (N128, N90, N21, N120, N81);
not NOT1 (N129, N116);
not NOT1 (N130, N127);
not NOT1 (N131, N126);
not NOT1 (N132, N129);
and AND2 (N133, N125, N70);
nand NAND4 (N134, N131, N55, N47, N77);
xor XOR2 (N135, N119, N12);
or OR4 (N136, N118, N113, N74, N49);
not NOT1 (N137, N122);
or OR2 (N138, N111, N94);
buf BUF1 (N139, N128);
buf BUF1 (N140, N135);
not NOT1 (N141, N140);
and AND2 (N142, N132, N42);
and AND4 (N143, N133, N83, N103, N44);
or OR2 (N144, N143, N107);
nor NOR3 (N145, N136, N4, N122);
not NOT1 (N146, N141);
and AND3 (N147, N130, N9, N62);
xor XOR2 (N148, N138, N5);
or OR4 (N149, N147, N102, N74, N51);
and AND4 (N150, N149, N93, N117, N120);
not NOT1 (N151, N139);
and AND4 (N152, N137, N88, N13, N86);
xor XOR2 (N153, N142, N45);
nand NAND3 (N154, N144, N142, N68);
and AND2 (N155, N134, N85);
nor NOR3 (N156, N148, N117, N151);
xor XOR2 (N157, N61, N16);
buf BUF1 (N158, N152);
buf BUF1 (N159, N155);
xor XOR2 (N160, N121, N85);
buf BUF1 (N161, N158);
or OR3 (N162, N156, N140, N142);
buf BUF1 (N163, N157);
not NOT1 (N164, N161);
nor NOR4 (N165, N150, N126, N131, N163);
not NOT1 (N166, N65);
buf BUF1 (N167, N166);
not NOT1 (N168, N167);
buf BUF1 (N169, N154);
not NOT1 (N170, N169);
xor XOR2 (N171, N170, N23);
nand NAND2 (N172, N162, N21);
buf BUF1 (N173, N171);
nand NAND2 (N174, N172, N91);
and AND4 (N175, N164, N131, N122, N25);
and AND3 (N176, N145, N96, N20);
buf BUF1 (N177, N168);
nand NAND2 (N178, N165, N154);
not NOT1 (N179, N173);
or OR2 (N180, N176, N6);
not NOT1 (N181, N146);
buf BUF1 (N182, N153);
not NOT1 (N183, N180);
xor XOR2 (N184, N159, N112);
nor NOR2 (N185, N181, N86);
buf BUF1 (N186, N184);
nand NAND3 (N187, N175, N158, N44);
xor XOR2 (N188, N183, N146);
not NOT1 (N189, N177);
and AND4 (N190, N179, N140, N177, N131);
nand NAND3 (N191, N190, N142, N38);
nand NAND4 (N192, N189, N14, N43, N63);
buf BUF1 (N193, N188);
xor XOR2 (N194, N191, N79);
nor NOR4 (N195, N186, N31, N63, N188);
nor NOR2 (N196, N193, N166);
not NOT1 (N197, N185);
not NOT1 (N198, N174);
and AND3 (N199, N195, N29, N192);
and AND4 (N200, N37, N174, N90, N172);
not NOT1 (N201, N200);
nor NOR4 (N202, N198, N129, N165, N187);
xor XOR2 (N203, N131, N82);
and AND3 (N204, N160, N73, N42);
xor XOR2 (N205, N204, N198);
nand NAND3 (N206, N202, N82, N185);
nand NAND2 (N207, N199, N93);
or OR4 (N208, N194, N179, N14, N197);
not NOT1 (N209, N52);
buf BUF1 (N210, N207);
nor NOR2 (N211, N178, N175);
buf BUF1 (N212, N208);
and AND4 (N213, N182, N201, N32, N145);
and AND2 (N214, N96, N73);
buf BUF1 (N215, N206);
xor XOR2 (N216, N210, N206);
not NOT1 (N217, N203);
buf BUF1 (N218, N212);
and AND4 (N219, N213, N2, N199, N193);
and AND2 (N220, N218, N86);
nand NAND2 (N221, N219, N127);
nand NAND4 (N222, N209, N127, N52, N55);
nor NOR3 (N223, N217, N216, N178);
xor XOR2 (N224, N108, N67);
nand NAND3 (N225, N220, N45, N114);
xor XOR2 (N226, N196, N172);
not NOT1 (N227, N211);
nand NAND3 (N228, N225, N225, N72);
xor XOR2 (N229, N215, N137);
xor XOR2 (N230, N222, N92);
nand NAND3 (N231, N227, N152, N195);
xor XOR2 (N232, N223, N62);
or OR4 (N233, N214, N164, N207, N164);
nor NOR2 (N234, N231, N213);
not NOT1 (N235, N229);
or OR2 (N236, N235, N74);
xor XOR2 (N237, N230, N82);
and AND2 (N238, N236, N44);
buf BUF1 (N239, N224);
not NOT1 (N240, N234);
xor XOR2 (N241, N221, N180);
xor XOR2 (N242, N239, N228);
nor NOR3 (N243, N98, N65, N45);
nand NAND3 (N244, N226, N209, N93);
and AND4 (N245, N237, N220, N51, N244);
nor NOR3 (N246, N113, N214, N132);
and AND2 (N247, N205, N141);
nor NOR4 (N248, N247, N155, N197, N159);
buf BUF1 (N249, N238);
not NOT1 (N250, N245);
xor XOR2 (N251, N250, N139);
buf BUF1 (N252, N251);
nor NOR3 (N253, N240, N55, N163);
xor XOR2 (N254, N242, N16);
xor XOR2 (N255, N248, N35);
buf BUF1 (N256, N249);
nor NOR2 (N257, N241, N9);
nand NAND2 (N258, N256, N143);
nand NAND3 (N259, N255, N209, N104);
buf BUF1 (N260, N253);
not NOT1 (N261, N260);
or OR2 (N262, N232, N222);
nor NOR4 (N263, N246, N6, N258, N27);
not NOT1 (N264, N114);
and AND2 (N265, N263, N201);
nor NOR4 (N266, N243, N104, N263, N224);
nand NAND2 (N267, N264, N250);
xor XOR2 (N268, N265, N164);
and AND4 (N269, N266, N267, N224, N180);
buf BUF1 (N270, N202);
and AND4 (N271, N261, N254, N144, N140);
and AND4 (N272, N4, N244, N106, N11);
and AND3 (N273, N233, N112, N145);
xor XOR2 (N274, N252, N107);
not NOT1 (N275, N273);
nor NOR4 (N276, N257, N67, N273, N36);
and AND4 (N277, N274, N189, N168, N208);
xor XOR2 (N278, N259, N18);
and AND4 (N279, N269, N46, N156, N3);
nand NAND2 (N280, N275, N103);
nor NOR3 (N281, N277, N106, N248);
buf BUF1 (N282, N272);
and AND4 (N283, N268, N253, N177, N165);
xor XOR2 (N284, N279, N141);
xor XOR2 (N285, N280, N18);
or OR3 (N286, N262, N125, N59);
not NOT1 (N287, N271);
nor NOR4 (N288, N281, N163, N223, N142);
and AND2 (N289, N287, N174);
nand NAND3 (N290, N286, N148, N91);
buf BUF1 (N291, N290);
buf BUF1 (N292, N289);
or OR4 (N293, N292, N157, N124, N235);
nand NAND4 (N294, N293, N220, N95, N101);
buf BUF1 (N295, N288);
buf BUF1 (N296, N283);
or OR3 (N297, N282, N243, N92);
xor XOR2 (N298, N294, N116);
not NOT1 (N299, N296);
nor NOR2 (N300, N270, N93);
nand NAND2 (N301, N285, N243);
nor NOR3 (N302, N278, N210, N300);
buf BUF1 (N303, N62);
and AND4 (N304, N291, N12, N79, N193);
not NOT1 (N305, N298);
buf BUF1 (N306, N284);
buf BUF1 (N307, N306);
nor NOR4 (N308, N295, N136, N237, N238);
and AND2 (N309, N302, N227);
and AND2 (N310, N299, N277);
and AND2 (N311, N305, N305);
not NOT1 (N312, N304);
buf BUF1 (N313, N301);
buf BUF1 (N314, N297);
or OR3 (N315, N314, N227, N3);
or OR2 (N316, N315, N260);
buf BUF1 (N317, N313);
and AND2 (N318, N303, N259);
nor NOR2 (N319, N276, N126);
nor NOR4 (N320, N319, N298, N175, N281);
nand NAND4 (N321, N312, N31, N121, N213);
xor XOR2 (N322, N308, N212);
xor XOR2 (N323, N322, N246);
or OR4 (N324, N316, N272, N225, N111);
or OR4 (N325, N317, N268, N279, N320);
buf BUF1 (N326, N279);
or OR3 (N327, N326, N29, N159);
xor XOR2 (N328, N324, N87);
xor XOR2 (N329, N321, N107);
nor NOR3 (N330, N307, N84, N254);
xor XOR2 (N331, N328, N72);
xor XOR2 (N332, N325, N314);
nand NAND2 (N333, N327, N315);
buf BUF1 (N334, N311);
xor XOR2 (N335, N309, N137);
buf BUF1 (N336, N335);
nor NOR2 (N337, N333, N315);
buf BUF1 (N338, N336);
nor NOR2 (N339, N334, N127);
buf BUF1 (N340, N337);
or OR3 (N341, N332, N84, N183);
buf BUF1 (N342, N331);
and AND4 (N343, N330, N177, N288, N163);
and AND3 (N344, N323, N226, N99);
not NOT1 (N345, N338);
and AND3 (N346, N341, N102, N323);
not NOT1 (N347, N342);
nor NOR2 (N348, N339, N328);
and AND4 (N349, N340, N232, N158, N234);
not NOT1 (N350, N310);
nor NOR4 (N351, N344, N95, N167, N120);
not NOT1 (N352, N329);
xor XOR2 (N353, N352, N31);
and AND4 (N354, N347, N73, N54, N247);
buf BUF1 (N355, N348);
or OR3 (N356, N345, N158, N187);
xor XOR2 (N357, N350, N224);
nand NAND3 (N358, N354, N47, N207);
buf BUF1 (N359, N355);
xor XOR2 (N360, N359, N157);
xor XOR2 (N361, N318, N88);
and AND4 (N362, N356, N79, N68, N330);
nand NAND4 (N363, N353, N153, N90, N5);
or OR4 (N364, N351, N197, N144, N335);
not NOT1 (N365, N343);
xor XOR2 (N366, N346, N195);
nand NAND4 (N367, N364, N336, N227, N83);
xor XOR2 (N368, N360, N306);
or OR3 (N369, N357, N226, N67);
or OR3 (N370, N349, N9, N131);
not NOT1 (N371, N368);
xor XOR2 (N372, N361, N239);
nand NAND4 (N373, N365, N3, N311, N310);
buf BUF1 (N374, N362);
or OR4 (N375, N374, N93, N187, N20);
or OR3 (N376, N375, N124, N346);
xor XOR2 (N377, N367, N56);
nand NAND4 (N378, N358, N41, N121, N142);
buf BUF1 (N379, N370);
nor NOR4 (N380, N377, N213, N350, N222);
not NOT1 (N381, N378);
buf BUF1 (N382, N372);
or OR2 (N383, N382, N114);
buf BUF1 (N384, N376);
xor XOR2 (N385, N373, N364);
xor XOR2 (N386, N381, N135);
nor NOR3 (N387, N371, N288, N373);
nor NOR3 (N388, N369, N56, N204);
buf BUF1 (N389, N379);
not NOT1 (N390, N366);
xor XOR2 (N391, N385, N342);
and AND2 (N392, N388, N46);
xor XOR2 (N393, N391, N103);
or OR2 (N394, N390, N266);
nand NAND3 (N395, N384, N68, N253);
buf BUF1 (N396, N393);
not NOT1 (N397, N389);
and AND2 (N398, N394, N260);
and AND4 (N399, N383, N252, N263, N35);
nor NOR2 (N400, N386, N205);
xor XOR2 (N401, N363, N79);
and AND3 (N402, N380, N240, N33);
and AND3 (N403, N402, N394, N147);
or OR3 (N404, N396, N340, N263);
not NOT1 (N405, N398);
nand NAND2 (N406, N400, N47);
and AND3 (N407, N401, N310, N346);
xor XOR2 (N408, N403, N400);
buf BUF1 (N409, N407);
or OR3 (N410, N387, N310, N146);
xor XOR2 (N411, N405, N62);
or OR2 (N412, N399, N258);
nand NAND4 (N413, N411, N172, N379, N190);
or OR2 (N414, N412, N386);
nor NOR3 (N415, N404, N169, N169);
not NOT1 (N416, N392);
nor NOR3 (N417, N413, N3, N227);
or OR2 (N418, N410, N397);
buf BUF1 (N419, N269);
xor XOR2 (N420, N414, N67);
buf BUF1 (N421, N408);
nor NOR3 (N422, N415, N400, N263);
xor XOR2 (N423, N417, N91);
and AND4 (N424, N423, N41, N246, N359);
and AND2 (N425, N420, N393);
buf BUF1 (N426, N409);
nor NOR4 (N427, N421, N351, N365, N271);
nand NAND2 (N428, N416, N350);
or OR2 (N429, N419, N213);
not NOT1 (N430, N395);
and AND4 (N431, N425, N181, N299, N128);
and AND3 (N432, N427, N199, N122);
buf BUF1 (N433, N426);
buf BUF1 (N434, N418);
or OR4 (N435, N431, N206, N111, N219);
nand NAND3 (N436, N434, N230, N19);
nand NAND4 (N437, N435, N381, N306, N44);
and AND4 (N438, N424, N318, N70, N116);
or OR2 (N439, N433, N316);
nand NAND2 (N440, N406, N406);
nor NOR2 (N441, N437, N239);
not NOT1 (N442, N432);
buf BUF1 (N443, N440);
and AND2 (N444, N438, N2);
not NOT1 (N445, N429);
nand NAND3 (N446, N422, N100, N88);
nand NAND4 (N447, N446, N39, N69, N6);
or OR2 (N448, N444, N163);
not NOT1 (N449, N430);
xor XOR2 (N450, N439, N382);
and AND4 (N451, N441, N355, N413, N129);
nor NOR4 (N452, N447, N349, N199, N430);
and AND4 (N453, N445, N12, N90, N154);
nor NOR4 (N454, N442, N253, N106, N305);
xor XOR2 (N455, N448, N51);
xor XOR2 (N456, N454, N71);
nand NAND2 (N457, N428, N440);
not NOT1 (N458, N452);
buf BUF1 (N459, N456);
buf BUF1 (N460, N453);
buf BUF1 (N461, N460);
nor NOR3 (N462, N461, N339, N188);
not NOT1 (N463, N449);
nand NAND2 (N464, N459, N171);
or OR4 (N465, N443, N296, N67, N2);
nor NOR2 (N466, N458, N189);
and AND2 (N467, N457, N235);
or OR3 (N468, N463, N265, N390);
nor NOR2 (N469, N436, N275);
xor XOR2 (N470, N464, N196);
and AND2 (N471, N466, N346);
not NOT1 (N472, N471);
xor XOR2 (N473, N472, N69);
and AND4 (N474, N450, N267, N88, N377);
or OR2 (N475, N473, N263);
and AND3 (N476, N474, N244, N389);
xor XOR2 (N477, N467, N437);
buf BUF1 (N478, N455);
and AND4 (N479, N469, N314, N370, N331);
or OR2 (N480, N465, N422);
buf BUF1 (N481, N451);
or OR4 (N482, N478, N72, N87, N366);
nor NOR2 (N483, N482, N237);
xor XOR2 (N484, N480, N17);
buf BUF1 (N485, N484);
xor XOR2 (N486, N483, N344);
nor NOR3 (N487, N476, N283, N133);
xor XOR2 (N488, N468, N411);
xor XOR2 (N489, N486, N397);
xor XOR2 (N490, N481, N85);
nor NOR3 (N491, N490, N453, N420);
buf BUF1 (N492, N475);
nor NOR3 (N493, N477, N434, N301);
nor NOR4 (N494, N493, N391, N419, N202);
and AND2 (N495, N462, N2);
buf BUF1 (N496, N470);
not NOT1 (N497, N488);
xor XOR2 (N498, N485, N144);
or OR3 (N499, N494, N208, N470);
nand NAND3 (N500, N496, N278, N119);
buf BUF1 (N501, N479);
or OR4 (N502, N500, N49, N242, N108);
not NOT1 (N503, N487);
xor XOR2 (N504, N503, N307);
nand NAND2 (N505, N498, N499);
not NOT1 (N506, N136);
buf BUF1 (N507, N506);
xor XOR2 (N508, N502, N434);
buf BUF1 (N509, N501);
not NOT1 (N510, N495);
nand NAND3 (N511, N489, N261, N379);
or OR3 (N512, N510, N452, N201);
buf BUF1 (N513, N507);
not NOT1 (N514, N497);
xor XOR2 (N515, N512, N145);
buf BUF1 (N516, N492);
and AND4 (N517, N509, N125, N100, N51);
not NOT1 (N518, N513);
buf BUF1 (N519, N505);
buf BUF1 (N520, N517);
not NOT1 (N521, N519);
nand NAND2 (N522, N520, N115);
buf BUF1 (N523, N508);
xor XOR2 (N524, N523, N422);
or OR3 (N525, N522, N143, N288);
and AND3 (N526, N515, N26, N370);
buf BUF1 (N527, N516);
nand NAND4 (N528, N518, N142, N217, N255);
xor XOR2 (N529, N528, N373);
buf BUF1 (N530, N526);
buf BUF1 (N531, N504);
buf BUF1 (N532, N524);
not NOT1 (N533, N521);
xor XOR2 (N534, N511, N192);
xor XOR2 (N535, N514, N302);
or OR2 (N536, N530, N237);
buf BUF1 (N537, N536);
nand NAND2 (N538, N525, N523);
and AND4 (N539, N532, N317, N483, N233);
xor XOR2 (N540, N534, N164);
buf BUF1 (N541, N540);
buf BUF1 (N542, N538);
or OR3 (N543, N533, N508, N400);
xor XOR2 (N544, N543, N154);
not NOT1 (N545, N529);
xor XOR2 (N546, N541, N452);
not NOT1 (N547, N535);
nor NOR2 (N548, N546, N179);
nand NAND3 (N549, N542, N167, N464);
nor NOR2 (N550, N549, N153);
and AND3 (N551, N548, N377, N224);
nand NAND2 (N552, N547, N224);
not NOT1 (N553, N551);
or OR3 (N554, N531, N205, N60);
buf BUF1 (N555, N550);
nor NOR3 (N556, N491, N539, N348);
nand NAND3 (N557, N419, N492, N310);
not NOT1 (N558, N554);
buf BUF1 (N559, N544);
not NOT1 (N560, N555);
xor XOR2 (N561, N559, N187);
nor NOR2 (N562, N557, N138);
or OR2 (N563, N545, N455);
xor XOR2 (N564, N556, N155);
or OR2 (N565, N537, N289);
nor NOR2 (N566, N564, N155);
or OR3 (N567, N560, N177, N336);
nand NAND4 (N568, N565, N89, N192, N87);
xor XOR2 (N569, N527, N409);
nand NAND2 (N570, N563, N487);
or OR3 (N571, N568, N50, N94);
nor NOR4 (N572, N571, N419, N239, N152);
buf BUF1 (N573, N552);
not NOT1 (N574, N562);
xor XOR2 (N575, N573, N353);
nand NAND2 (N576, N553, N478);
or OR3 (N577, N570, N398, N477);
xor XOR2 (N578, N561, N61);
xor XOR2 (N579, N569, N202);
and AND2 (N580, N579, N79);
not NOT1 (N581, N574);
or OR2 (N582, N575, N476);
nor NOR3 (N583, N558, N480, N194);
xor XOR2 (N584, N582, N423);
not NOT1 (N585, N580);
buf BUF1 (N586, N576);
xor XOR2 (N587, N584, N475);
and AND2 (N588, N585, N464);
nand NAND3 (N589, N572, N84, N141);
nor NOR3 (N590, N588, N29, N490);
and AND4 (N591, N586, N100, N140, N453);
buf BUF1 (N592, N581);
and AND2 (N593, N578, N120);
not NOT1 (N594, N587);
nand NAND2 (N595, N594, N542);
buf BUF1 (N596, N595);
not NOT1 (N597, N596);
buf BUF1 (N598, N591);
buf BUF1 (N599, N567);
not NOT1 (N600, N583);
and AND4 (N601, N589, N244, N354, N262);
buf BUF1 (N602, N599);
not NOT1 (N603, N600);
or OR2 (N604, N592, N204);
and AND4 (N605, N597, N158, N188, N451);
and AND2 (N606, N593, N272);
nand NAND3 (N607, N601, N117, N13);
nand NAND3 (N608, N604, N482, N99);
nand NAND4 (N609, N566, N252, N183, N378);
or OR3 (N610, N598, N201, N579);
nand NAND2 (N611, N605, N219);
xor XOR2 (N612, N607, N380);
or OR2 (N613, N590, N294);
or OR3 (N614, N610, N70, N372);
buf BUF1 (N615, N612);
or OR2 (N616, N608, N412);
buf BUF1 (N617, N577);
nor NOR2 (N618, N603, N521);
or OR2 (N619, N606, N485);
and AND4 (N620, N615, N208, N467, N69);
nand NAND2 (N621, N614, N293);
and AND4 (N622, N620, N95, N32, N418);
nor NOR3 (N623, N613, N95, N293);
and AND4 (N624, N617, N187, N298, N49);
not NOT1 (N625, N619);
nor NOR4 (N626, N623, N591, N621, N64);
and AND2 (N627, N429, N299);
not NOT1 (N628, N624);
nand NAND4 (N629, N626, N253, N264, N46);
xor XOR2 (N630, N629, N431);
and AND4 (N631, N616, N396, N544, N206);
not NOT1 (N632, N609);
or OR4 (N633, N630, N22, N560, N558);
or OR3 (N634, N622, N94, N591);
or OR2 (N635, N632, N219);
not NOT1 (N636, N634);
and AND2 (N637, N618, N515);
buf BUF1 (N638, N631);
or OR2 (N639, N638, N200);
not NOT1 (N640, N627);
buf BUF1 (N641, N636);
nor NOR3 (N642, N639, N333, N327);
nor NOR3 (N643, N602, N92, N467);
xor XOR2 (N644, N633, N542);
and AND3 (N645, N637, N93, N459);
not NOT1 (N646, N645);
not NOT1 (N647, N646);
and AND3 (N648, N628, N50, N475);
or OR3 (N649, N647, N53, N414);
or OR3 (N650, N644, N63, N525);
nor NOR2 (N651, N611, N8);
buf BUF1 (N652, N651);
not NOT1 (N653, N642);
and AND3 (N654, N635, N580, N550);
nand NAND3 (N655, N643, N324, N289);
or OR2 (N656, N654, N522);
not NOT1 (N657, N649);
xor XOR2 (N658, N641, N124);
buf BUF1 (N659, N658);
buf BUF1 (N660, N640);
nor NOR4 (N661, N652, N184, N212, N49);
or OR3 (N662, N648, N418, N566);
not NOT1 (N663, N661);
buf BUF1 (N664, N653);
xor XOR2 (N665, N656, N27);
and AND4 (N666, N625, N105, N461, N29);
or OR2 (N667, N664, N217);
or OR3 (N668, N650, N595, N38);
buf BUF1 (N669, N667);
nand NAND3 (N670, N660, N162, N424);
xor XOR2 (N671, N655, N442);
xor XOR2 (N672, N657, N285);
or OR3 (N673, N665, N470, N513);
xor XOR2 (N674, N669, N254);
or OR2 (N675, N663, N212);
or OR3 (N676, N662, N361, N98);
not NOT1 (N677, N670);
and AND2 (N678, N676, N492);
nor NOR3 (N679, N659, N253, N439);
and AND2 (N680, N668, N135);
or OR2 (N681, N680, N9);
and AND2 (N682, N677, N482);
nand NAND2 (N683, N681, N345);
not NOT1 (N684, N671);
xor XOR2 (N685, N678, N60);
not NOT1 (N686, N679);
nor NOR4 (N687, N686, N159, N71, N246);
buf BUF1 (N688, N666);
or OR4 (N689, N684, N619, N602, N659);
buf BUF1 (N690, N675);
and AND3 (N691, N674, N33, N633);
or OR4 (N692, N683, N562, N130, N272);
nor NOR3 (N693, N673, N372, N624);
or OR4 (N694, N682, N455, N643, N676);
nand NAND3 (N695, N693, N42, N77);
or OR4 (N696, N690, N395, N152, N110);
or OR2 (N697, N689, N530);
nor NOR3 (N698, N688, N271, N406);
and AND2 (N699, N695, N455);
xor XOR2 (N700, N696, N193);
buf BUF1 (N701, N692);
and AND3 (N702, N687, N585, N133);
and AND2 (N703, N698, N276);
not NOT1 (N704, N697);
buf BUF1 (N705, N685);
or OR2 (N706, N701, N261);
not NOT1 (N707, N705);
buf BUF1 (N708, N703);
or OR4 (N709, N706, N277, N195, N195);
not NOT1 (N710, N707);
nand NAND3 (N711, N709, N244, N588);
xor XOR2 (N712, N700, N660);
nor NOR3 (N713, N704, N37, N687);
nand NAND4 (N714, N699, N525, N572, N504);
xor XOR2 (N715, N691, N693);
nor NOR4 (N716, N713, N615, N585, N403);
or OR3 (N717, N716, N334, N235);
nand NAND2 (N718, N672, N442);
nor NOR2 (N719, N711, N247);
not NOT1 (N720, N719);
nor NOR2 (N721, N702, N121);
or OR4 (N722, N717, N471, N704, N169);
or OR4 (N723, N715, N457, N31, N382);
and AND4 (N724, N714, N274, N13, N167);
nand NAND2 (N725, N722, N108);
nor NOR4 (N726, N721, N437, N508, N137);
xor XOR2 (N727, N725, N591);
buf BUF1 (N728, N712);
not NOT1 (N729, N726);
not NOT1 (N730, N718);
nor NOR4 (N731, N729, N482, N419, N511);
buf BUF1 (N732, N727);
nand NAND2 (N733, N708, N323);
not NOT1 (N734, N733);
and AND3 (N735, N720, N246, N111);
nor NOR4 (N736, N728, N545, N733, N59);
not NOT1 (N737, N723);
not NOT1 (N738, N724);
not NOT1 (N739, N730);
and AND2 (N740, N734, N369);
nor NOR2 (N741, N738, N407);
buf BUF1 (N742, N731);
or OR4 (N743, N742, N731, N397, N417);
xor XOR2 (N744, N737, N219);
nand NAND2 (N745, N739, N722);
and AND2 (N746, N736, N234);
nor NOR4 (N747, N746, N740, N553, N584);
xor XOR2 (N748, N138, N657);
nor NOR2 (N749, N735, N168);
and AND3 (N750, N745, N579, N718);
nand NAND4 (N751, N732, N645, N138, N620);
and AND4 (N752, N747, N732, N479, N466);
nor NOR2 (N753, N741, N121);
xor XOR2 (N754, N744, N361);
nor NOR2 (N755, N743, N366);
not NOT1 (N756, N751);
xor XOR2 (N757, N756, N249);
buf BUF1 (N758, N750);
nor NOR3 (N759, N749, N73, N90);
nand NAND4 (N760, N757, N424, N652, N591);
buf BUF1 (N761, N753);
and AND3 (N762, N760, N661, N90);
xor XOR2 (N763, N754, N438);
or OR4 (N764, N752, N136, N724, N50);
xor XOR2 (N765, N710, N75);
xor XOR2 (N766, N748, N486);
buf BUF1 (N767, N759);
and AND4 (N768, N767, N316, N608, N349);
nor NOR4 (N769, N762, N708, N732, N164);
xor XOR2 (N770, N766, N758);
and AND3 (N771, N234, N39, N225);
or OR2 (N772, N765, N52);
xor XOR2 (N773, N770, N186);
not NOT1 (N774, N763);
or OR2 (N775, N774, N142);
nand NAND3 (N776, N768, N106, N322);
and AND3 (N777, N761, N683, N213);
and AND2 (N778, N755, N659);
nor NOR2 (N779, N694, N290);
nand NAND4 (N780, N773, N762, N44, N221);
xor XOR2 (N781, N772, N51);
and AND4 (N782, N775, N337, N24, N541);
or OR4 (N783, N779, N429, N336, N244);
nand NAND2 (N784, N782, N292);
nor NOR2 (N785, N771, N438);
nand NAND3 (N786, N769, N19, N727);
and AND2 (N787, N776, N538);
buf BUF1 (N788, N784);
nand NAND2 (N789, N780, N295);
or OR2 (N790, N786, N106);
and AND4 (N791, N783, N669, N382, N205);
or OR4 (N792, N791, N120, N118, N198);
or OR3 (N793, N781, N593, N209);
not NOT1 (N794, N793);
buf BUF1 (N795, N787);
and AND2 (N796, N764, N59);
and AND2 (N797, N777, N109);
nand NAND4 (N798, N796, N604, N747, N132);
buf BUF1 (N799, N792);
buf BUF1 (N800, N794);
xor XOR2 (N801, N785, N767);
buf BUF1 (N802, N801);
nor NOR2 (N803, N799, N65);
or OR3 (N804, N778, N443, N10);
nor NOR3 (N805, N804, N229, N582);
nor NOR3 (N806, N789, N330, N702);
buf BUF1 (N807, N795);
nor NOR3 (N808, N790, N254, N154);
buf BUF1 (N809, N800);
xor XOR2 (N810, N808, N85);
nand NAND2 (N811, N805, N115);
or OR3 (N812, N811, N27, N112);
buf BUF1 (N813, N812);
and AND3 (N814, N809, N791, N591);
nor NOR3 (N815, N788, N522, N442);
nand NAND2 (N816, N803, N367);
or OR2 (N817, N802, N161);
nand NAND2 (N818, N816, N536);
or OR3 (N819, N815, N643, N625);
buf BUF1 (N820, N817);
nand NAND4 (N821, N814, N179, N178, N87);
xor XOR2 (N822, N820, N613);
xor XOR2 (N823, N798, N166);
nor NOR3 (N824, N821, N629, N159);
nand NAND4 (N825, N813, N792, N10, N156);
nand NAND2 (N826, N797, N694);
or OR4 (N827, N810, N748, N369, N370);
xor XOR2 (N828, N824, N594);
not NOT1 (N829, N819);
xor XOR2 (N830, N822, N455);
nor NOR2 (N831, N829, N131);
nand NAND3 (N832, N831, N646, N32);
not NOT1 (N833, N830);
buf BUF1 (N834, N823);
xor XOR2 (N835, N826, N343);
not NOT1 (N836, N832);
xor XOR2 (N837, N827, N61);
or OR2 (N838, N807, N598);
buf BUF1 (N839, N834);
buf BUF1 (N840, N835);
buf BUF1 (N841, N838);
buf BUF1 (N842, N837);
xor XOR2 (N843, N825, N352);
nand NAND4 (N844, N840, N469, N55, N527);
not NOT1 (N845, N828);
nor NOR3 (N846, N836, N187, N74);
and AND4 (N847, N833, N718, N235, N73);
and AND4 (N848, N843, N449, N19, N98);
nand NAND3 (N849, N818, N778, N481);
nor NOR4 (N850, N849, N703, N755, N639);
nor NOR4 (N851, N842, N533, N375, N84);
and AND4 (N852, N850, N813, N504, N53);
nand NAND2 (N853, N841, N318);
not NOT1 (N854, N839);
nor NOR4 (N855, N848, N203, N9, N147);
nor NOR3 (N856, N845, N646, N245);
xor XOR2 (N857, N853, N560);
nand NAND2 (N858, N806, N825);
buf BUF1 (N859, N847);
nand NAND4 (N860, N859, N821, N775, N148);
or OR2 (N861, N852, N68);
not NOT1 (N862, N860);
or OR4 (N863, N854, N311, N523, N66);
buf BUF1 (N864, N846);
nand NAND4 (N865, N856, N379, N840, N20);
nor NOR4 (N866, N864, N521, N127, N663);
and AND2 (N867, N858, N738);
and AND2 (N868, N844, N233);
xor XOR2 (N869, N866, N151);
or OR2 (N870, N863, N226);
buf BUF1 (N871, N870);
or OR3 (N872, N855, N136, N751);
and AND3 (N873, N868, N864, N199);
or OR4 (N874, N867, N54, N590, N383);
xor XOR2 (N875, N869, N739);
xor XOR2 (N876, N872, N281);
nand NAND4 (N877, N876, N502, N472, N420);
and AND3 (N878, N877, N21, N406);
xor XOR2 (N879, N871, N613);
not NOT1 (N880, N857);
xor XOR2 (N881, N873, N726);
buf BUF1 (N882, N874);
nor NOR3 (N883, N875, N330, N141);
or OR4 (N884, N878, N725, N648, N505);
or OR4 (N885, N880, N309, N283, N242);
and AND4 (N886, N882, N326, N175, N381);
nor NOR3 (N887, N851, N42, N369);
not NOT1 (N888, N886);
not NOT1 (N889, N881);
nor NOR3 (N890, N885, N693, N38);
or OR3 (N891, N879, N796, N194);
xor XOR2 (N892, N862, N108);
xor XOR2 (N893, N889, N448);
buf BUF1 (N894, N891);
buf BUF1 (N895, N861);
or OR2 (N896, N865, N712);
not NOT1 (N897, N883);
or OR2 (N898, N888, N145);
buf BUF1 (N899, N895);
and AND2 (N900, N894, N191);
or OR3 (N901, N892, N252, N224);
nor NOR3 (N902, N890, N635, N506);
and AND3 (N903, N899, N341, N792);
nand NAND2 (N904, N901, N159);
buf BUF1 (N905, N900);
nand NAND4 (N906, N905, N444, N79, N296);
buf BUF1 (N907, N887);
nand NAND4 (N908, N906, N768, N222, N651);
nand NAND4 (N909, N896, N95, N275, N291);
and AND2 (N910, N902, N591);
buf BUF1 (N911, N893);
buf BUF1 (N912, N884);
and AND2 (N913, N911, N694);
not NOT1 (N914, N912);
nor NOR4 (N915, N913, N67, N254, N642);
and AND3 (N916, N909, N288, N41);
buf BUF1 (N917, N898);
nor NOR3 (N918, N897, N457, N420);
nand NAND4 (N919, N908, N824, N298, N534);
not NOT1 (N920, N903);
buf BUF1 (N921, N919);
xor XOR2 (N922, N910, N821);
xor XOR2 (N923, N922, N124);
not NOT1 (N924, N918);
and AND3 (N925, N923, N489, N269);
buf BUF1 (N926, N907);
and AND3 (N927, N920, N855, N491);
not NOT1 (N928, N917);
or OR3 (N929, N926, N23, N656);
nor NOR4 (N930, N904, N206, N465, N576);
not NOT1 (N931, N914);
buf BUF1 (N932, N916);
and AND3 (N933, N932, N96, N423);
and AND2 (N934, N930, N231);
xor XOR2 (N935, N929, N81);
buf BUF1 (N936, N934);
nand NAND4 (N937, N928, N361, N651, N817);
buf BUF1 (N938, N933);
or OR2 (N939, N925, N272);
or OR2 (N940, N927, N428);
xor XOR2 (N941, N915, N761);
nand NAND4 (N942, N931, N899, N211, N237);
buf BUF1 (N943, N941);
nand NAND4 (N944, N937, N689, N748, N202);
nand NAND3 (N945, N924, N118, N417);
or OR3 (N946, N942, N887, N17);
and AND3 (N947, N935, N892, N195);
or OR2 (N948, N944, N919);
nor NOR4 (N949, N940, N662, N450, N474);
xor XOR2 (N950, N921, N91);
xor XOR2 (N951, N950, N131);
nand NAND3 (N952, N945, N161, N169);
nand NAND4 (N953, N946, N333, N374, N320);
xor XOR2 (N954, N949, N675);
buf BUF1 (N955, N954);
or OR4 (N956, N938, N432, N181, N740);
not NOT1 (N957, N948);
buf BUF1 (N958, N936);
or OR2 (N959, N939, N338);
nand NAND4 (N960, N959, N225, N193, N282);
nor NOR4 (N961, N960, N31, N204, N230);
and AND3 (N962, N952, N470, N603);
or OR4 (N963, N951, N424, N553, N794);
and AND4 (N964, N943, N430, N533, N190);
not NOT1 (N965, N953);
buf BUF1 (N966, N955);
and AND3 (N967, N963, N196, N846);
xor XOR2 (N968, N958, N209);
not NOT1 (N969, N967);
xor XOR2 (N970, N964, N268);
nand NAND2 (N971, N970, N800);
and AND2 (N972, N968, N626);
nand NAND2 (N973, N947, N850);
nor NOR3 (N974, N972, N60, N828);
or OR2 (N975, N962, N680);
nor NOR4 (N976, N966, N352, N496, N61);
buf BUF1 (N977, N965);
and AND4 (N978, N977, N16, N303, N746);
xor XOR2 (N979, N973, N32);
or OR3 (N980, N969, N452, N544);
not NOT1 (N981, N976);
buf BUF1 (N982, N979);
or OR3 (N983, N961, N272, N163);
or OR2 (N984, N978, N391);
or OR4 (N985, N971, N923, N841, N802);
nor NOR3 (N986, N956, N900, N263);
nor NOR3 (N987, N980, N318, N851);
nor NOR3 (N988, N957, N615, N414);
buf BUF1 (N989, N975);
and AND2 (N990, N989, N97);
nor NOR4 (N991, N981, N490, N505, N779);
or OR4 (N992, N990, N692, N522, N498);
xor XOR2 (N993, N987, N191);
not NOT1 (N994, N991);
buf BUF1 (N995, N992);
nand NAND4 (N996, N993, N541, N645, N651);
and AND2 (N997, N982, N914);
nor NOR2 (N998, N983, N252);
or OR2 (N999, N995, N431);
and AND4 (N1000, N984, N563, N306, N593);
and AND3 (N1001, N997, N453, N204);
or OR4 (N1002, N996, N494, N445, N891);
nand NAND2 (N1003, N986, N173);
nand NAND3 (N1004, N1002, N373, N460);
xor XOR2 (N1005, N985, N4);
and AND2 (N1006, N998, N666);
or OR3 (N1007, N1005, N425, N390);
nand NAND3 (N1008, N1003, N10, N193);
not NOT1 (N1009, N994);
buf BUF1 (N1010, N1006);
not NOT1 (N1011, N974);
or OR2 (N1012, N1000, N311);
xor XOR2 (N1013, N1009, N957);
buf BUF1 (N1014, N999);
and AND4 (N1015, N988, N436, N80, N763);
nor NOR3 (N1016, N1010, N138, N1003);
buf BUF1 (N1017, N1007);
buf BUF1 (N1018, N1001);
nor NOR3 (N1019, N1011, N79, N737);
not NOT1 (N1020, N1008);
buf BUF1 (N1021, N1019);
nand NAND4 (N1022, N1017, N264, N546, N166);
not NOT1 (N1023, N1014);
nand NAND3 (N1024, N1016, N219, N304);
nand NAND4 (N1025, N1012, N530, N26, N728);
nand NAND3 (N1026, N1023, N117, N612);
not NOT1 (N1027, N1022);
xor XOR2 (N1028, N1021, N1009);
not NOT1 (N1029, N1013);
nor NOR2 (N1030, N1004, N577);
buf BUF1 (N1031, N1029);
or OR3 (N1032, N1020, N952, N742);
nand NAND4 (N1033, N1025, N540, N322, N798);
buf BUF1 (N1034, N1026);
xor XOR2 (N1035, N1034, N470);
not NOT1 (N1036, N1015);
and AND4 (N1037, N1018, N685, N153, N179);
not NOT1 (N1038, N1035);
or OR3 (N1039, N1028, N552, N836);
xor XOR2 (N1040, N1031, N992);
not NOT1 (N1041, N1033);
xor XOR2 (N1042, N1030, N190);
or OR4 (N1043, N1037, N513, N1019, N804);
xor XOR2 (N1044, N1040, N72);
and AND3 (N1045, N1027, N851, N186);
nand NAND4 (N1046, N1042, N308, N182, N813);
nand NAND2 (N1047, N1043, N696);
and AND4 (N1048, N1047, N162, N160, N19);
nor NOR2 (N1049, N1032, N115);
buf BUF1 (N1050, N1044);
or OR3 (N1051, N1039, N759, N2);
buf BUF1 (N1052, N1046);
xor XOR2 (N1053, N1038, N607);
buf BUF1 (N1054, N1050);
and AND2 (N1055, N1052, N228);
xor XOR2 (N1056, N1051, N64);
and AND3 (N1057, N1024, N836, N172);
xor XOR2 (N1058, N1054, N196);
not NOT1 (N1059, N1055);
buf BUF1 (N1060, N1036);
not NOT1 (N1061, N1053);
or OR4 (N1062, N1041, N354, N908, N732);
buf BUF1 (N1063, N1049);
nand NAND4 (N1064, N1062, N206, N710, N554);
and AND3 (N1065, N1057, N850, N68);
or OR4 (N1066, N1058, N67, N984, N678);
or OR2 (N1067, N1060, N171);
nor NOR3 (N1068, N1061, N143, N606);
not NOT1 (N1069, N1064);
nor NOR2 (N1070, N1059, N736);
xor XOR2 (N1071, N1045, N459);
xor XOR2 (N1072, N1063, N620);
or OR3 (N1073, N1068, N410, N416);
buf BUF1 (N1074, N1070);
nand NAND4 (N1075, N1067, N592, N355, N581);
xor XOR2 (N1076, N1071, N613);
xor XOR2 (N1077, N1075, N630);
xor XOR2 (N1078, N1074, N35);
nand NAND3 (N1079, N1056, N534, N1039);
or OR3 (N1080, N1048, N1017, N358);
not NOT1 (N1081, N1069);
not NOT1 (N1082, N1080);
not NOT1 (N1083, N1072);
nor NOR2 (N1084, N1065, N572);
nor NOR4 (N1085, N1078, N1037, N802, N704);
and AND3 (N1086, N1066, N675, N273);
not NOT1 (N1087, N1076);
buf BUF1 (N1088, N1077);
or OR2 (N1089, N1088, N282);
nand NAND4 (N1090, N1079, N697, N642, N309);
buf BUF1 (N1091, N1085);
nor NOR3 (N1092, N1091, N365, N570);
nor NOR4 (N1093, N1084, N310, N84, N665);
and AND4 (N1094, N1092, N975, N213, N78);
buf BUF1 (N1095, N1093);
buf BUF1 (N1096, N1083);
nand NAND3 (N1097, N1095, N514, N923);
buf BUF1 (N1098, N1094);
or OR3 (N1099, N1098, N572, N289);
nand NAND3 (N1100, N1087, N907, N974);
nor NOR4 (N1101, N1089, N593, N158, N538);
not NOT1 (N1102, N1096);
not NOT1 (N1103, N1102);
buf BUF1 (N1104, N1082);
and AND3 (N1105, N1103, N893, N1011);
not NOT1 (N1106, N1101);
not NOT1 (N1107, N1100);
xor XOR2 (N1108, N1090, N671);
not NOT1 (N1109, N1086);
xor XOR2 (N1110, N1097, N498);
or OR2 (N1111, N1105, N117);
xor XOR2 (N1112, N1106, N1107);
buf BUF1 (N1113, N72);
nand NAND3 (N1114, N1113, N560, N852);
and AND4 (N1115, N1104, N1100, N671, N902);
not NOT1 (N1116, N1110);
not NOT1 (N1117, N1081);
nand NAND3 (N1118, N1111, N124, N770);
buf BUF1 (N1119, N1108);
buf BUF1 (N1120, N1119);
xor XOR2 (N1121, N1073, N914);
nor NOR4 (N1122, N1115, N334, N821, N108);
xor XOR2 (N1123, N1116, N914);
nand NAND4 (N1124, N1118, N592, N1047, N1100);
and AND2 (N1125, N1124, N253);
xor XOR2 (N1126, N1125, N942);
nand NAND3 (N1127, N1121, N732, N599);
buf BUF1 (N1128, N1120);
xor XOR2 (N1129, N1114, N470);
nor NOR4 (N1130, N1123, N283, N254, N748);
buf BUF1 (N1131, N1129);
buf BUF1 (N1132, N1130);
nor NOR2 (N1133, N1112, N454);
or OR3 (N1134, N1128, N1087, N356);
not NOT1 (N1135, N1126);
and AND3 (N1136, N1127, N883, N479);
xor XOR2 (N1137, N1117, N360);
xor XOR2 (N1138, N1135, N111);
not NOT1 (N1139, N1133);
nand NAND3 (N1140, N1136, N798, N734);
xor XOR2 (N1141, N1131, N156);
and AND3 (N1142, N1140, N136, N224);
or OR4 (N1143, N1132, N1125, N334, N379);
nand NAND3 (N1144, N1099, N297, N65);
or OR4 (N1145, N1109, N949, N252, N613);
xor XOR2 (N1146, N1145, N612);
nor NOR3 (N1147, N1139, N135, N210);
and AND4 (N1148, N1142, N1120, N524, N286);
xor XOR2 (N1149, N1146, N544);
and AND3 (N1150, N1137, N1146, N1016);
not NOT1 (N1151, N1143);
nand NAND2 (N1152, N1149, N520);
nor NOR2 (N1153, N1122, N554);
or OR3 (N1154, N1148, N236, N373);
buf BUF1 (N1155, N1141);
nor NOR2 (N1156, N1155, N171);
buf BUF1 (N1157, N1147);
xor XOR2 (N1158, N1151, N593);
nand NAND2 (N1159, N1158, N388);
nor NOR4 (N1160, N1154, N727, N179, N346);
xor XOR2 (N1161, N1156, N251);
and AND4 (N1162, N1134, N806, N721, N402);
buf BUF1 (N1163, N1153);
not NOT1 (N1164, N1138);
nand NAND2 (N1165, N1164, N792);
buf BUF1 (N1166, N1152);
nor NOR4 (N1167, N1166, N106, N839, N712);
xor XOR2 (N1168, N1160, N724);
xor XOR2 (N1169, N1157, N59);
xor XOR2 (N1170, N1167, N270);
nor NOR3 (N1171, N1161, N388, N604);
not NOT1 (N1172, N1162);
nand NAND2 (N1173, N1172, N1050);
or OR2 (N1174, N1169, N172);
xor XOR2 (N1175, N1159, N59);
buf BUF1 (N1176, N1150);
nor NOR3 (N1177, N1168, N257, N1153);
not NOT1 (N1178, N1173);
or OR4 (N1179, N1163, N394, N152, N432);
nand NAND3 (N1180, N1175, N487, N376);
buf BUF1 (N1181, N1174);
and AND3 (N1182, N1180, N527, N248);
not NOT1 (N1183, N1144);
nor NOR2 (N1184, N1181, N155);
not NOT1 (N1185, N1171);
nor NOR4 (N1186, N1179, N241, N726, N720);
buf BUF1 (N1187, N1178);
or OR2 (N1188, N1183, N1131);
and AND3 (N1189, N1165, N806, N31);
buf BUF1 (N1190, N1188);
nor NOR2 (N1191, N1189, N762);
nor NOR3 (N1192, N1176, N1023, N535);
buf BUF1 (N1193, N1190);
buf BUF1 (N1194, N1185);
buf BUF1 (N1195, N1184);
and AND4 (N1196, N1187, N969, N740, N464);
not NOT1 (N1197, N1195);
and AND3 (N1198, N1192, N709, N1066);
nor NOR3 (N1199, N1182, N454, N146);
xor XOR2 (N1200, N1170, N804);
not NOT1 (N1201, N1198);
nor NOR4 (N1202, N1194, N498, N1002, N783);
buf BUF1 (N1203, N1193);
nand NAND4 (N1204, N1191, N932, N681, N649);
nor NOR3 (N1205, N1177, N50, N504);
xor XOR2 (N1206, N1197, N401);
nand NAND4 (N1207, N1205, N1041, N773, N620);
buf BUF1 (N1208, N1206);
nand NAND2 (N1209, N1199, N472);
xor XOR2 (N1210, N1201, N576);
and AND2 (N1211, N1186, N1164);
xor XOR2 (N1212, N1207, N644);
or OR2 (N1213, N1210, N758);
xor XOR2 (N1214, N1203, N723);
or OR3 (N1215, N1212, N177, N171);
buf BUF1 (N1216, N1213);
buf BUF1 (N1217, N1200);
nand NAND2 (N1218, N1204, N459);
nand NAND4 (N1219, N1215, N248, N239, N1105);
xor XOR2 (N1220, N1202, N15);
nand NAND2 (N1221, N1219, N894);
xor XOR2 (N1222, N1208, N611);
buf BUF1 (N1223, N1221);
not NOT1 (N1224, N1217);
or OR4 (N1225, N1211, N60, N1101, N1214);
and AND2 (N1226, N65, N1194);
buf BUF1 (N1227, N1218);
nor NOR3 (N1228, N1223, N116, N361);
nor NOR3 (N1229, N1216, N910, N1149);
or OR2 (N1230, N1196, N16);
and AND2 (N1231, N1226, N1213);
nor NOR2 (N1232, N1227, N246);
and AND2 (N1233, N1232, N9);
and AND3 (N1234, N1230, N494, N44);
nand NAND2 (N1235, N1229, N317);
and AND2 (N1236, N1235, N175);
nand NAND3 (N1237, N1222, N156, N1031);
or OR2 (N1238, N1236, N715);
buf BUF1 (N1239, N1234);
buf BUF1 (N1240, N1238);
xor XOR2 (N1241, N1240, N452);
not NOT1 (N1242, N1209);
and AND2 (N1243, N1233, N87);
buf BUF1 (N1244, N1239);
nand NAND2 (N1245, N1220, N90);
nor NOR3 (N1246, N1243, N20, N60);
not NOT1 (N1247, N1242);
and AND4 (N1248, N1245, N858, N179, N225);
xor XOR2 (N1249, N1231, N1068);
or OR4 (N1250, N1228, N451, N571, N786);
not NOT1 (N1251, N1247);
or OR4 (N1252, N1241, N415, N830, N447);
and AND2 (N1253, N1252, N535);
nor NOR2 (N1254, N1237, N404);
buf BUF1 (N1255, N1248);
nor NOR2 (N1256, N1225, N705);
xor XOR2 (N1257, N1224, N713);
xor XOR2 (N1258, N1257, N989);
buf BUF1 (N1259, N1253);
and AND4 (N1260, N1258, N489, N234, N135);
or OR4 (N1261, N1250, N146, N717, N1042);
or OR2 (N1262, N1251, N247);
nand NAND4 (N1263, N1254, N643, N452, N142);
nor NOR4 (N1264, N1261, N818, N571, N1196);
nor NOR4 (N1265, N1262, N354, N787, N682);
or OR2 (N1266, N1244, N445);
nand NAND2 (N1267, N1246, N534);
buf BUF1 (N1268, N1260);
nand NAND3 (N1269, N1249, N193, N94);
and AND3 (N1270, N1263, N997, N1072);
or OR3 (N1271, N1259, N794, N638);
buf BUF1 (N1272, N1264);
nand NAND3 (N1273, N1256, N433, N358);
xor XOR2 (N1274, N1271, N772);
nand NAND3 (N1275, N1274, N953, N359);
and AND4 (N1276, N1255, N1040, N1255, N947);
nand NAND3 (N1277, N1267, N354, N282);
and AND3 (N1278, N1277, N1126, N924);
nand NAND3 (N1279, N1265, N484, N15);
buf BUF1 (N1280, N1278);
nand NAND3 (N1281, N1272, N1018, N177);
or OR4 (N1282, N1280, N191, N144, N590);
xor XOR2 (N1283, N1275, N700);
buf BUF1 (N1284, N1282);
buf BUF1 (N1285, N1273);
nand NAND3 (N1286, N1268, N263, N628);
nand NAND2 (N1287, N1284, N1016);
buf BUF1 (N1288, N1283);
not NOT1 (N1289, N1281);
not NOT1 (N1290, N1286);
xor XOR2 (N1291, N1285, N177);
nand NAND4 (N1292, N1266, N6, N151, N1056);
xor XOR2 (N1293, N1290, N135);
not NOT1 (N1294, N1269);
xor XOR2 (N1295, N1270, N1014);
nand NAND2 (N1296, N1279, N125);
nor NOR3 (N1297, N1294, N44, N1018);
and AND3 (N1298, N1288, N1265, N1025);
xor XOR2 (N1299, N1295, N1042);
or OR3 (N1300, N1292, N243, N932);
and AND2 (N1301, N1276, N165);
buf BUF1 (N1302, N1291);
xor XOR2 (N1303, N1301, N375);
nand NAND2 (N1304, N1296, N740);
xor XOR2 (N1305, N1289, N436);
buf BUF1 (N1306, N1303);
or OR2 (N1307, N1293, N472);
not NOT1 (N1308, N1287);
not NOT1 (N1309, N1304);
not NOT1 (N1310, N1299);
nand NAND4 (N1311, N1305, N1135, N304, N843);
nand NAND2 (N1312, N1302, N1043);
and AND3 (N1313, N1308, N391, N23);
not NOT1 (N1314, N1298);
nand NAND3 (N1315, N1306, N1106, N246);
buf BUF1 (N1316, N1312);
buf BUF1 (N1317, N1300);
not NOT1 (N1318, N1297);
or OR4 (N1319, N1317, N777, N78, N1067);
or OR2 (N1320, N1311, N447);
and AND4 (N1321, N1310, N1318, N130, N1284);
buf BUF1 (N1322, N419);
nand NAND4 (N1323, N1307, N203, N1050, N276);
and AND2 (N1324, N1321, N25);
or OR3 (N1325, N1320, N376, N1048);
buf BUF1 (N1326, N1313);
or OR3 (N1327, N1314, N583, N110);
nand NAND4 (N1328, N1322, N40, N255, N689);
nor NOR3 (N1329, N1327, N873, N1243);
or OR3 (N1330, N1325, N544, N29);
buf BUF1 (N1331, N1315);
or OR3 (N1332, N1309, N429, N648);
nand NAND3 (N1333, N1319, N862, N1039);
and AND3 (N1334, N1323, N515, N787);
or OR4 (N1335, N1334, N1173, N1263, N531);
or OR3 (N1336, N1329, N711, N301);
xor XOR2 (N1337, N1331, N472);
not NOT1 (N1338, N1332);
not NOT1 (N1339, N1335);
not NOT1 (N1340, N1316);
xor XOR2 (N1341, N1330, N971);
and AND3 (N1342, N1339, N927, N390);
nor NOR3 (N1343, N1340, N491, N956);
nor NOR3 (N1344, N1337, N1218, N688);
xor XOR2 (N1345, N1328, N320);
buf BUF1 (N1346, N1324);
nand NAND2 (N1347, N1336, N1109);
xor XOR2 (N1348, N1346, N569);
not NOT1 (N1349, N1326);
or OR3 (N1350, N1349, N315, N89);
xor XOR2 (N1351, N1347, N585);
and AND4 (N1352, N1351, N1155, N143, N389);
nand NAND2 (N1353, N1342, N471);
xor XOR2 (N1354, N1345, N1273);
nor NOR2 (N1355, N1348, N489);
and AND2 (N1356, N1352, N1137);
nor NOR2 (N1357, N1355, N757);
nand NAND2 (N1358, N1341, N427);
nand NAND3 (N1359, N1344, N1242, N236);
and AND4 (N1360, N1338, N553, N645, N963);
nor NOR4 (N1361, N1360, N527, N471, N2);
and AND4 (N1362, N1354, N234, N386, N358);
nand NAND2 (N1363, N1356, N697);
nor NOR3 (N1364, N1359, N14, N1289);
or OR2 (N1365, N1353, N617);
nand NAND3 (N1366, N1363, N1055, N289);
xor XOR2 (N1367, N1365, N35);
not NOT1 (N1368, N1362);
buf BUF1 (N1369, N1343);
nor NOR2 (N1370, N1357, N985);
and AND3 (N1371, N1369, N150, N582);
or OR4 (N1372, N1368, N91, N431, N1180);
nand NAND2 (N1373, N1371, N21);
not NOT1 (N1374, N1361);
and AND3 (N1375, N1372, N279, N331);
not NOT1 (N1376, N1358);
or OR3 (N1377, N1367, N661, N162);
xor XOR2 (N1378, N1375, N252);
buf BUF1 (N1379, N1370);
buf BUF1 (N1380, N1333);
or OR4 (N1381, N1379, N599, N1280, N548);
and AND4 (N1382, N1376, N1168, N506, N877);
xor XOR2 (N1383, N1374, N256);
nand NAND3 (N1384, N1382, N898, N1337);
or OR4 (N1385, N1383, N550, N410, N568);
buf BUF1 (N1386, N1384);
buf BUF1 (N1387, N1373);
and AND2 (N1388, N1385, N659);
buf BUF1 (N1389, N1364);
nor NOR2 (N1390, N1386, N1089);
and AND2 (N1391, N1378, N18);
nand NAND3 (N1392, N1350, N609, N660);
or OR3 (N1393, N1387, N555, N918);
nand NAND2 (N1394, N1381, N894);
or OR4 (N1395, N1377, N1392, N868, N778);
not NOT1 (N1396, N4);
nand NAND4 (N1397, N1389, N349, N623, N979);
xor XOR2 (N1398, N1394, N647);
nand NAND4 (N1399, N1388, N526, N361, N1145);
nand NAND2 (N1400, N1393, N172);
nand NAND2 (N1401, N1397, N941);
nor NOR3 (N1402, N1400, N579, N290);
nor NOR4 (N1403, N1401, N833, N199, N114);
nand NAND2 (N1404, N1398, N848);
xor XOR2 (N1405, N1403, N216);
buf BUF1 (N1406, N1405);
xor XOR2 (N1407, N1396, N1339);
nand NAND4 (N1408, N1399, N1338, N1255, N1318);
or OR2 (N1409, N1402, N560);
or OR2 (N1410, N1404, N366);
not NOT1 (N1411, N1391);
not NOT1 (N1412, N1408);
or OR3 (N1413, N1380, N850, N1200);
nand NAND2 (N1414, N1395, N134);
nor NOR3 (N1415, N1414, N1162, N29);
and AND4 (N1416, N1411, N937, N782, N1374);
xor XOR2 (N1417, N1410, N393);
buf BUF1 (N1418, N1409);
nand NAND2 (N1419, N1418, N654);
and AND2 (N1420, N1366, N344);
nor NOR2 (N1421, N1412, N476);
xor XOR2 (N1422, N1421, N330);
not NOT1 (N1423, N1390);
nand NAND2 (N1424, N1406, N1062);
nor NOR2 (N1425, N1415, N1243);
xor XOR2 (N1426, N1423, N223);
and AND3 (N1427, N1420, N318, N712);
nor NOR2 (N1428, N1419, N231);
or OR2 (N1429, N1416, N897);
nand NAND3 (N1430, N1425, N1333, N1412);
not NOT1 (N1431, N1429);
or OR4 (N1432, N1431, N1150, N678, N1054);
or OR2 (N1433, N1426, N555);
not NOT1 (N1434, N1407);
not NOT1 (N1435, N1434);
not NOT1 (N1436, N1428);
and AND4 (N1437, N1436, N271, N921, N716);
not NOT1 (N1438, N1413);
or OR2 (N1439, N1435, N547);
nand NAND2 (N1440, N1432, N858);
or OR4 (N1441, N1424, N3, N1268, N154);
buf BUF1 (N1442, N1417);
nand NAND4 (N1443, N1442, N329, N1400, N229);
nor NOR2 (N1444, N1427, N885);
xor XOR2 (N1445, N1433, N1156);
nand NAND2 (N1446, N1422, N1216);
xor XOR2 (N1447, N1446, N153);
xor XOR2 (N1448, N1440, N1212);
xor XOR2 (N1449, N1430, N344);
or OR4 (N1450, N1449, N107, N538, N843);
nand NAND3 (N1451, N1448, N610, N1438);
nand NAND4 (N1452, N634, N1350, N636, N505);
nor NOR3 (N1453, N1439, N207, N1246);
xor XOR2 (N1454, N1453, N532);
nand NAND2 (N1455, N1447, N84);
nor NOR2 (N1456, N1443, N333);
and AND4 (N1457, N1444, N336, N600, N296);
xor XOR2 (N1458, N1456, N610);
or OR2 (N1459, N1441, N633);
not NOT1 (N1460, N1459);
nand NAND2 (N1461, N1451, N191);
nand NAND2 (N1462, N1461, N116);
buf BUF1 (N1463, N1452);
and AND2 (N1464, N1457, N1086);
buf BUF1 (N1465, N1454);
and AND4 (N1466, N1455, N248, N1143, N87);
not NOT1 (N1467, N1437);
and AND2 (N1468, N1467, N673);
and AND4 (N1469, N1463, N230, N664, N19);
nor NOR4 (N1470, N1445, N621, N892, N299);
nand NAND2 (N1471, N1460, N416);
nor NOR2 (N1472, N1470, N494);
not NOT1 (N1473, N1468);
not NOT1 (N1474, N1458);
buf BUF1 (N1475, N1473);
nor NOR3 (N1476, N1466, N210, N396);
and AND4 (N1477, N1476, N859, N390, N1141);
xor XOR2 (N1478, N1472, N1372);
or OR4 (N1479, N1471, N198, N340, N280);
or OR2 (N1480, N1477, N1051);
buf BUF1 (N1481, N1479);
nand NAND4 (N1482, N1469, N294, N170, N925);
xor XOR2 (N1483, N1481, N879);
not NOT1 (N1484, N1480);
or OR3 (N1485, N1475, N1276, N288);
nor NOR3 (N1486, N1462, N1459, N12);
xor XOR2 (N1487, N1485, N1181);
or OR4 (N1488, N1464, N899, N1206, N977);
nand NAND3 (N1489, N1474, N1112, N1198);
not NOT1 (N1490, N1483);
buf BUF1 (N1491, N1482);
and AND3 (N1492, N1489, N459, N862);
nand NAND3 (N1493, N1450, N682, N315);
nor NOR4 (N1494, N1484, N2, N529, N1401);
not NOT1 (N1495, N1487);
or OR4 (N1496, N1491, N867, N831, N990);
nor NOR4 (N1497, N1486, N1490, N1212, N1448);
nor NOR2 (N1498, N173, N764);
or OR4 (N1499, N1498, N1133, N1395, N129);
xor XOR2 (N1500, N1493, N76);
nor NOR4 (N1501, N1465, N1130, N1364, N739);
and AND3 (N1502, N1497, N836, N1369);
buf BUF1 (N1503, N1488);
nor NOR4 (N1504, N1492, N1219, N898, N1441);
nand NAND2 (N1505, N1501, N684);
or OR2 (N1506, N1504, N253);
nand NAND3 (N1507, N1499, N633, N800);
not NOT1 (N1508, N1478);
nand NAND2 (N1509, N1502, N649);
xor XOR2 (N1510, N1506, N664);
xor XOR2 (N1511, N1507, N701);
nor NOR3 (N1512, N1500, N493, N1057);
xor XOR2 (N1513, N1511, N229);
nor NOR4 (N1514, N1513, N1451, N1463, N150);
xor XOR2 (N1515, N1512, N226);
xor XOR2 (N1516, N1494, N1367);
or OR3 (N1517, N1514, N1387, N373);
nor NOR3 (N1518, N1503, N988, N1383);
nor NOR3 (N1519, N1518, N408, N907);
xor XOR2 (N1520, N1517, N1375);
xor XOR2 (N1521, N1509, N997);
buf BUF1 (N1522, N1496);
or OR2 (N1523, N1495, N1478);
or OR4 (N1524, N1523, N577, N1223, N1114);
not NOT1 (N1525, N1522);
nand NAND4 (N1526, N1510, N1007, N734, N1172);
xor XOR2 (N1527, N1524, N1459);
and AND3 (N1528, N1525, N2, N1033);
and AND2 (N1529, N1505, N196);
or OR4 (N1530, N1520, N589, N1095, N1297);
and AND2 (N1531, N1526, N1036);
or OR4 (N1532, N1515, N1031, N478, N748);
nand NAND4 (N1533, N1532, N963, N1002, N741);
and AND2 (N1534, N1530, N180);
or OR2 (N1535, N1533, N306);
and AND3 (N1536, N1508, N954, N510);
buf BUF1 (N1537, N1535);
and AND4 (N1538, N1536, N863, N1330, N1221);
and AND4 (N1539, N1519, N1453, N120, N1038);
buf BUF1 (N1540, N1529);
or OR2 (N1541, N1534, N830);
xor XOR2 (N1542, N1531, N1393);
buf BUF1 (N1543, N1540);
nand NAND4 (N1544, N1521, N240, N34, N11);
nor NOR3 (N1545, N1528, N83, N122);
and AND4 (N1546, N1545, N1185, N834, N1009);
and AND4 (N1547, N1538, N1099, N1294, N195);
xor XOR2 (N1548, N1539, N782);
nor NOR3 (N1549, N1527, N375, N1527);
buf BUF1 (N1550, N1547);
xor XOR2 (N1551, N1548, N1193);
nor NOR3 (N1552, N1546, N340, N306);
or OR4 (N1553, N1552, N265, N973, N1477);
and AND2 (N1554, N1553, N383);
not NOT1 (N1555, N1541);
or OR2 (N1556, N1537, N192);
or OR3 (N1557, N1542, N527, N571);
nor NOR2 (N1558, N1557, N320);
xor XOR2 (N1559, N1550, N91);
nor NOR4 (N1560, N1555, N1504, N1103, N894);
buf BUF1 (N1561, N1558);
xor XOR2 (N1562, N1551, N1520);
buf BUF1 (N1563, N1544);
and AND3 (N1564, N1560, N1490, N571);
or OR3 (N1565, N1561, N1121, N467);
buf BUF1 (N1566, N1554);
xor XOR2 (N1567, N1549, N716);
not NOT1 (N1568, N1564);
and AND4 (N1569, N1566, N416, N489, N1534);
and AND4 (N1570, N1569, N189, N56, N914);
or OR4 (N1571, N1563, N1188, N1014, N1362);
and AND4 (N1572, N1565, N699, N43, N539);
and AND3 (N1573, N1543, N454, N707);
buf BUF1 (N1574, N1573);
or OR3 (N1575, N1559, N442, N751);
or OR3 (N1576, N1516, N1339, N1460);
or OR2 (N1577, N1576, N1523);
and AND3 (N1578, N1568, N372, N1018);
nand NAND3 (N1579, N1556, N703, N1138);
and AND2 (N1580, N1577, N840);
buf BUF1 (N1581, N1579);
nand NAND4 (N1582, N1562, N1423, N552, N491);
nor NOR4 (N1583, N1574, N1378, N1347, N688);
nor NOR3 (N1584, N1580, N1038, N118);
nor NOR3 (N1585, N1571, N1555, N1048);
or OR2 (N1586, N1570, N1372);
nand NAND3 (N1587, N1582, N1480, N1146);
or OR3 (N1588, N1586, N1215, N1381);
not NOT1 (N1589, N1575);
not NOT1 (N1590, N1584);
buf BUF1 (N1591, N1589);
not NOT1 (N1592, N1587);
xor XOR2 (N1593, N1591, N267);
nand NAND2 (N1594, N1578, N72);
not NOT1 (N1595, N1585);
nor NOR4 (N1596, N1588, N529, N997, N1547);
buf BUF1 (N1597, N1572);
nand NAND2 (N1598, N1583, N596);
xor XOR2 (N1599, N1593, N348);
nand NAND2 (N1600, N1598, N585);
buf BUF1 (N1601, N1581);
nand NAND2 (N1602, N1595, N583);
nand NAND4 (N1603, N1602, N1438, N509, N1015);
and AND2 (N1604, N1590, N1050);
not NOT1 (N1605, N1603);
nor NOR3 (N1606, N1594, N338, N1450);
not NOT1 (N1607, N1567);
buf BUF1 (N1608, N1600);
or OR2 (N1609, N1597, N52);
and AND4 (N1610, N1609, N1456, N952, N944);
buf BUF1 (N1611, N1601);
and AND3 (N1612, N1608, N1519, N1392);
not NOT1 (N1613, N1611);
nor NOR2 (N1614, N1599, N711);
buf BUF1 (N1615, N1596);
not NOT1 (N1616, N1612);
or OR2 (N1617, N1616, N1066);
buf BUF1 (N1618, N1606);
nand NAND2 (N1619, N1613, N1237);
nand NAND4 (N1620, N1618, N897, N906, N90);
nand NAND4 (N1621, N1620, N189, N550, N444);
buf BUF1 (N1622, N1621);
xor XOR2 (N1623, N1622, N1185);
not NOT1 (N1624, N1604);
nand NAND3 (N1625, N1619, N633, N976);
nand NAND3 (N1626, N1615, N867, N257);
or OR3 (N1627, N1625, N216, N1562);
nor NOR4 (N1628, N1627, N1445, N952, N1518);
and AND2 (N1629, N1614, N995);
nand NAND2 (N1630, N1607, N130);
or OR2 (N1631, N1630, N726);
nand NAND3 (N1632, N1610, N360, N414);
nand NAND3 (N1633, N1623, N235, N476);
or OR4 (N1634, N1632, N982, N1532, N894);
xor XOR2 (N1635, N1629, N1491);
and AND2 (N1636, N1631, N990);
buf BUF1 (N1637, N1605);
xor XOR2 (N1638, N1592, N1073);
nor NOR4 (N1639, N1633, N1384, N636, N1442);
buf BUF1 (N1640, N1626);
and AND2 (N1641, N1628, N1180);
buf BUF1 (N1642, N1634);
nor NOR3 (N1643, N1637, N1440, N224);
or OR2 (N1644, N1636, N65);
and AND4 (N1645, N1635, N884, N61, N308);
xor XOR2 (N1646, N1638, N970);
buf BUF1 (N1647, N1624);
xor XOR2 (N1648, N1642, N1645);
nand NAND3 (N1649, N1621, N1502, N1638);
nor NOR2 (N1650, N1640, N772);
and AND4 (N1651, N1643, N1493, N600, N56);
buf BUF1 (N1652, N1644);
and AND2 (N1653, N1649, N1498);
nor NOR4 (N1654, N1650, N1015, N755, N337);
nand NAND4 (N1655, N1653, N355, N1222, N1102);
nand NAND2 (N1656, N1641, N1333);
nor NOR3 (N1657, N1652, N1494, N1061);
nor NOR4 (N1658, N1656, N1338, N152, N78);
and AND2 (N1659, N1617, N171);
not NOT1 (N1660, N1651);
xor XOR2 (N1661, N1654, N517);
nand NAND3 (N1662, N1646, N1556, N537);
and AND4 (N1663, N1657, N336, N578, N240);
nand NAND3 (N1664, N1658, N1377, N1047);
not NOT1 (N1665, N1659);
or OR4 (N1666, N1648, N1387, N1200, N585);
nor NOR2 (N1667, N1660, N860);
not NOT1 (N1668, N1662);
and AND3 (N1669, N1667, N674, N1612);
xor XOR2 (N1670, N1639, N516);
nand NAND4 (N1671, N1669, N1513, N307, N454);
nor NOR4 (N1672, N1647, N1143, N813, N218);
nand NAND2 (N1673, N1661, N292);
buf BUF1 (N1674, N1672);
xor XOR2 (N1675, N1670, N87);
or OR3 (N1676, N1673, N584, N78);
nor NOR3 (N1677, N1664, N430, N87);
nand NAND2 (N1678, N1675, N276);
nor NOR3 (N1679, N1674, N729, N347);
buf BUF1 (N1680, N1676);
or OR4 (N1681, N1666, N632, N252, N846);
not NOT1 (N1682, N1677);
or OR2 (N1683, N1678, N453);
nand NAND2 (N1684, N1663, N1165);
or OR2 (N1685, N1671, N1330);
xor XOR2 (N1686, N1682, N824);
not NOT1 (N1687, N1668);
and AND4 (N1688, N1686, N1073, N773, N1536);
buf BUF1 (N1689, N1681);
or OR4 (N1690, N1655, N498, N995, N1508);
xor XOR2 (N1691, N1685, N425);
or OR2 (N1692, N1680, N1135);
buf BUF1 (N1693, N1683);
and AND2 (N1694, N1691, N365);
not NOT1 (N1695, N1693);
or OR3 (N1696, N1692, N1079, N342);
nor NOR2 (N1697, N1696, N1214);
xor XOR2 (N1698, N1687, N1239);
not NOT1 (N1699, N1695);
or OR2 (N1700, N1684, N712);
nand NAND2 (N1701, N1698, N882);
or OR3 (N1702, N1679, N228, N332);
or OR2 (N1703, N1699, N1436);
nand NAND3 (N1704, N1702, N1507, N446);
and AND2 (N1705, N1688, N351);
nand NAND3 (N1706, N1700, N1036, N575);
nor NOR3 (N1707, N1703, N299, N1665);
nand NAND3 (N1708, N1625, N1471, N913);
nand NAND2 (N1709, N1690, N479);
xor XOR2 (N1710, N1697, N435);
nor NOR2 (N1711, N1689, N686);
or OR2 (N1712, N1710, N1049);
xor XOR2 (N1713, N1707, N526);
or OR4 (N1714, N1706, N1644, N467, N1397);
and AND2 (N1715, N1694, N1499);
nand NAND2 (N1716, N1701, N749);
not NOT1 (N1717, N1713);
not NOT1 (N1718, N1711);
or OR2 (N1719, N1714, N1372);
nand NAND4 (N1720, N1717, N1045, N168, N1059);
nand NAND2 (N1721, N1708, N144);
xor XOR2 (N1722, N1709, N623);
buf BUF1 (N1723, N1712);
nand NAND3 (N1724, N1715, N438, N352);
nor NOR4 (N1725, N1705, N111, N874, N872);
and AND2 (N1726, N1725, N1227);
xor XOR2 (N1727, N1720, N899);
not NOT1 (N1728, N1724);
xor XOR2 (N1729, N1722, N1705);
nand NAND4 (N1730, N1721, N484, N339, N210);
xor XOR2 (N1731, N1729, N451);
xor XOR2 (N1732, N1731, N1480);
nand NAND4 (N1733, N1730, N606, N1038, N1128);
or OR2 (N1734, N1719, N1728);
xor XOR2 (N1735, N1216, N1382);
xor XOR2 (N1736, N1727, N1321);
not NOT1 (N1737, N1723);
or OR2 (N1738, N1736, N1282);
not NOT1 (N1739, N1726);
nor NOR4 (N1740, N1739, N1665, N475, N532);
nor NOR2 (N1741, N1732, N1335);
xor XOR2 (N1742, N1716, N736);
buf BUF1 (N1743, N1733);
not NOT1 (N1744, N1704);
or OR4 (N1745, N1744, N1164, N747, N686);
buf BUF1 (N1746, N1740);
xor XOR2 (N1747, N1738, N804);
or OR4 (N1748, N1745, N489, N1421, N1409);
and AND3 (N1749, N1742, N1116, N688);
and AND3 (N1750, N1743, N1705, N1129);
xor XOR2 (N1751, N1735, N163);
nor NOR3 (N1752, N1749, N1400, N1745);
or OR3 (N1753, N1751, N1227, N1138);
and AND4 (N1754, N1741, N275, N1443, N422);
xor XOR2 (N1755, N1747, N1091);
and AND2 (N1756, N1737, N367);
nand NAND3 (N1757, N1752, N1594, N1502);
nand NAND2 (N1758, N1734, N1741);
or OR3 (N1759, N1754, N611, N146);
xor XOR2 (N1760, N1746, N487);
or OR3 (N1761, N1759, N945, N903);
nor NOR3 (N1762, N1756, N510, N1322);
nor NOR2 (N1763, N1753, N811);
or OR3 (N1764, N1758, N1753, N1307);
buf BUF1 (N1765, N1718);
nor NOR4 (N1766, N1762, N960, N945, N1347);
not NOT1 (N1767, N1757);
buf BUF1 (N1768, N1765);
and AND2 (N1769, N1748, N967);
or OR2 (N1770, N1750, N983);
or OR2 (N1771, N1768, N992);
nand NAND4 (N1772, N1755, N1652, N1532, N1451);
xor XOR2 (N1773, N1764, N921);
xor XOR2 (N1774, N1770, N1013);
and AND2 (N1775, N1767, N944);
not NOT1 (N1776, N1766);
xor XOR2 (N1777, N1763, N1436);
nor NOR3 (N1778, N1775, N941, N191);
and AND3 (N1779, N1773, N1001, N781);
xor XOR2 (N1780, N1771, N556);
not NOT1 (N1781, N1769);
nor NOR2 (N1782, N1778, N1319);
nor NOR3 (N1783, N1777, N1339, N376);
nor NOR2 (N1784, N1760, N1494);
not NOT1 (N1785, N1782);
or OR3 (N1786, N1781, N926, N1089);
nand NAND4 (N1787, N1774, N28, N822, N1189);
xor XOR2 (N1788, N1780, N1658);
nor NOR3 (N1789, N1788, N893, N667);
nor NOR3 (N1790, N1784, N1654, N1688);
nand NAND4 (N1791, N1776, N1477, N248, N404);
or OR2 (N1792, N1761, N622);
buf BUF1 (N1793, N1789);
xor XOR2 (N1794, N1787, N624);
not NOT1 (N1795, N1785);
not NOT1 (N1796, N1791);
nor NOR2 (N1797, N1790, N1015);
nand NAND4 (N1798, N1795, N66, N639, N520);
nand NAND4 (N1799, N1779, N951, N476, N257);
and AND4 (N1800, N1794, N355, N43, N886);
buf BUF1 (N1801, N1796);
and AND4 (N1802, N1798, N1296, N220, N1146);
and AND4 (N1803, N1792, N162, N676, N915);
and AND4 (N1804, N1799, N556, N320, N311);
and AND3 (N1805, N1783, N534, N459);
nand NAND3 (N1806, N1797, N235, N1082);
nand NAND4 (N1807, N1803, N1272, N1650, N240);
and AND3 (N1808, N1804, N1082, N749);
not NOT1 (N1809, N1800);
not NOT1 (N1810, N1786);
buf BUF1 (N1811, N1807);
nand NAND3 (N1812, N1802, N1754, N423);
nor NOR3 (N1813, N1806, N775, N560);
xor XOR2 (N1814, N1793, N282);
or OR3 (N1815, N1808, N877, N595);
not NOT1 (N1816, N1815);
not NOT1 (N1817, N1772);
and AND2 (N1818, N1816, N1167);
xor XOR2 (N1819, N1813, N723);
buf BUF1 (N1820, N1819);
and AND3 (N1821, N1810, N1258, N141);
buf BUF1 (N1822, N1821);
or OR2 (N1823, N1817, N81);
not NOT1 (N1824, N1809);
buf BUF1 (N1825, N1805);
and AND4 (N1826, N1820, N1413, N1721, N646);
and AND2 (N1827, N1818, N1641);
nor NOR2 (N1828, N1814, N1123);
and AND3 (N1829, N1825, N436, N314);
buf BUF1 (N1830, N1812);
buf BUF1 (N1831, N1829);
not NOT1 (N1832, N1801);
nor NOR4 (N1833, N1826, N1077, N200, N521);
and AND2 (N1834, N1828, N657);
and AND2 (N1835, N1832, N48);
buf BUF1 (N1836, N1827);
xor XOR2 (N1837, N1811, N677);
xor XOR2 (N1838, N1834, N383);
or OR2 (N1839, N1824, N798);
or OR2 (N1840, N1837, N1190);
nor NOR3 (N1841, N1833, N1717, N909);
not NOT1 (N1842, N1836);
not NOT1 (N1843, N1831);
buf BUF1 (N1844, N1843);
buf BUF1 (N1845, N1842);
or OR3 (N1846, N1822, N1089, N264);
xor XOR2 (N1847, N1845, N641);
nand NAND4 (N1848, N1844, N874, N115, N1064);
nand NAND2 (N1849, N1838, N418);
not NOT1 (N1850, N1847);
and AND4 (N1851, N1848, N1022, N292, N1569);
nor NOR2 (N1852, N1850, N1547);
or OR2 (N1853, N1849, N1315);
buf BUF1 (N1854, N1830);
nor NOR3 (N1855, N1851, N246, N667);
nand NAND3 (N1856, N1835, N86, N1086);
nand NAND4 (N1857, N1823, N774, N1856, N400);
nand NAND4 (N1858, N1752, N1038, N1267, N1274);
buf BUF1 (N1859, N1852);
or OR4 (N1860, N1855, N1495, N1113, N1654);
not NOT1 (N1861, N1840);
nand NAND2 (N1862, N1858, N956);
nor NOR2 (N1863, N1859, N1418);
buf BUF1 (N1864, N1857);
not NOT1 (N1865, N1853);
or OR4 (N1866, N1839, N1232, N661, N185);
nor NOR4 (N1867, N1860, N1307, N1017, N461);
and AND3 (N1868, N1866, N507, N504);
xor XOR2 (N1869, N1867, N1647);
not NOT1 (N1870, N1865);
buf BUF1 (N1871, N1862);
xor XOR2 (N1872, N1854, N970);
not NOT1 (N1873, N1870);
nand NAND3 (N1874, N1846, N1009, N194);
nor NOR4 (N1875, N1873, N1309, N1682, N1148);
not NOT1 (N1876, N1864);
not NOT1 (N1877, N1874);
not NOT1 (N1878, N1869);
buf BUF1 (N1879, N1841);
and AND4 (N1880, N1863, N1486, N1429, N1121);
not NOT1 (N1881, N1872);
xor XOR2 (N1882, N1868, N1842);
buf BUF1 (N1883, N1875);
and AND4 (N1884, N1861, N484, N762, N1090);
nor NOR2 (N1885, N1878, N1089);
xor XOR2 (N1886, N1879, N71);
xor XOR2 (N1887, N1885, N1229);
or OR2 (N1888, N1881, N1492);
nand NAND2 (N1889, N1886, N1344);
not NOT1 (N1890, N1876);
nand NAND3 (N1891, N1880, N731, N546);
or OR3 (N1892, N1883, N1123, N1502);
or OR2 (N1893, N1891, N308);
buf BUF1 (N1894, N1890);
buf BUF1 (N1895, N1889);
or OR3 (N1896, N1882, N1871, N75);
buf BUF1 (N1897, N638);
nand NAND3 (N1898, N1892, N1642, N809);
xor XOR2 (N1899, N1893, N787);
nand NAND2 (N1900, N1898, N1757);
or OR4 (N1901, N1900, N315, N545, N1487);
nand NAND3 (N1902, N1894, N955, N536);
nand NAND3 (N1903, N1897, N1584, N393);
nand NAND4 (N1904, N1902, N1450, N1506, N268);
not NOT1 (N1905, N1896);
xor XOR2 (N1906, N1888, N1433);
not NOT1 (N1907, N1905);
nor NOR4 (N1908, N1895, N1129, N415, N1700);
nand NAND3 (N1909, N1901, N71, N870);
or OR3 (N1910, N1908, N729, N1675);
xor XOR2 (N1911, N1910, N1821);
or OR2 (N1912, N1903, N1133);
and AND4 (N1913, N1887, N1138, N21, N790);
nand NAND2 (N1914, N1911, N1626);
nor NOR3 (N1915, N1909, N1304, N1411);
and AND2 (N1916, N1906, N133);
buf BUF1 (N1917, N1912);
not NOT1 (N1918, N1884);
or OR4 (N1919, N1904, N270, N1552, N1152);
not NOT1 (N1920, N1907);
or OR2 (N1921, N1899, N97);
xor XOR2 (N1922, N1920, N500);
or OR2 (N1923, N1877, N714);
buf BUF1 (N1924, N1918);
nor NOR4 (N1925, N1917, N261, N267, N1708);
not NOT1 (N1926, N1921);
and AND4 (N1927, N1915, N783, N1385, N1576);
xor XOR2 (N1928, N1913, N1577);
buf BUF1 (N1929, N1925);
nor NOR2 (N1930, N1916, N779);
nand NAND4 (N1931, N1914, N850, N168, N1702);
nand NAND2 (N1932, N1931, N81);
and AND4 (N1933, N1930, N486, N1606, N1880);
nor NOR2 (N1934, N1922, N460);
nor NOR2 (N1935, N1927, N1032);
or OR2 (N1936, N1934, N690);
xor XOR2 (N1937, N1924, N391);
buf BUF1 (N1938, N1923);
and AND2 (N1939, N1933, N874);
nor NOR2 (N1940, N1937, N1287);
not NOT1 (N1941, N1935);
nor NOR2 (N1942, N1928, N1708);
or OR4 (N1943, N1926, N257, N1816, N1538);
and AND3 (N1944, N1941, N1089, N1434);
or OR2 (N1945, N1932, N95);
xor XOR2 (N1946, N1938, N1338);
buf BUF1 (N1947, N1940);
or OR4 (N1948, N1936, N922, N443, N647);
or OR4 (N1949, N1919, N483, N1756, N655);
buf BUF1 (N1950, N1942);
nor NOR4 (N1951, N1946, N1788, N1494, N196);
nand NAND2 (N1952, N1939, N731);
xor XOR2 (N1953, N1951, N472);
not NOT1 (N1954, N1952);
nor NOR3 (N1955, N1945, N1944, N894);
nand NAND4 (N1956, N1928, N1814, N301, N423);
xor XOR2 (N1957, N1943, N984);
buf BUF1 (N1958, N1949);
nand NAND3 (N1959, N1953, N1619, N1859);
xor XOR2 (N1960, N1957, N549);
not NOT1 (N1961, N1950);
buf BUF1 (N1962, N1960);
not NOT1 (N1963, N1956);
or OR2 (N1964, N1958, N756);
buf BUF1 (N1965, N1963);
and AND2 (N1966, N1961, N1568);
xor XOR2 (N1967, N1955, N191);
and AND3 (N1968, N1959, N794, N1639);
buf BUF1 (N1969, N1948);
or OR3 (N1970, N1967, N1889, N636);
or OR2 (N1971, N1947, N1074);
xor XOR2 (N1972, N1971, N1748);
xor XOR2 (N1973, N1966, N739);
nor NOR3 (N1974, N1970, N1346, N519);
or OR2 (N1975, N1929, N676);
not NOT1 (N1976, N1954);
not NOT1 (N1977, N1972);
nand NAND3 (N1978, N1973, N1666, N527);
or OR2 (N1979, N1977, N1468);
and AND2 (N1980, N1976, N1268);
xor XOR2 (N1981, N1965, N1373);
nor NOR3 (N1982, N1980, N851, N468);
nand NAND4 (N1983, N1975, N1583, N1391, N813);
not NOT1 (N1984, N1962);
or OR2 (N1985, N1969, N1535);
buf BUF1 (N1986, N1964);
buf BUF1 (N1987, N1979);
buf BUF1 (N1988, N1978);
xor XOR2 (N1989, N1988, N153);
not NOT1 (N1990, N1982);
buf BUF1 (N1991, N1984);
nor NOR4 (N1992, N1968, N1332, N1117, N599);
not NOT1 (N1993, N1991);
xor XOR2 (N1994, N1993, N1437);
and AND2 (N1995, N1992, N1669);
xor XOR2 (N1996, N1974, N1340);
or OR3 (N1997, N1983, N806, N986);
nand NAND3 (N1998, N1985, N809, N223);
and AND4 (N1999, N1996, N1102, N1253, N1754);
not NOT1 (N2000, N1998);
or OR4 (N2001, N2000, N675, N1967, N592);
not NOT1 (N2002, N1990);
or OR4 (N2003, N1981, N951, N943, N1129);
nor NOR4 (N2004, N1997, N543, N519, N1595);
nor NOR3 (N2005, N1987, N1611, N155);
buf BUF1 (N2006, N2002);
nor NOR3 (N2007, N1989, N253, N1949);
nor NOR3 (N2008, N2006, N1110, N460);
nor NOR2 (N2009, N2007, N1254);
not NOT1 (N2010, N1999);
nand NAND3 (N2011, N2009, N1816, N605);
not NOT1 (N2012, N2011);
buf BUF1 (N2013, N2004);
buf BUF1 (N2014, N2003);
nand NAND4 (N2015, N2014, N135, N1475, N491);
nand NAND3 (N2016, N2001, N712, N1168);
or OR4 (N2017, N1986, N791, N609, N250);
or OR3 (N2018, N2016, N1021, N293);
or OR3 (N2019, N2015, N1324, N1410);
nor NOR3 (N2020, N2013, N774, N1554);
xor XOR2 (N2021, N2012, N630);
xor XOR2 (N2022, N2018, N151);
or OR3 (N2023, N2017, N879, N1111);
xor XOR2 (N2024, N2008, N1201);
not NOT1 (N2025, N1995);
or OR3 (N2026, N2010, N736, N1155);
xor XOR2 (N2027, N2025, N304);
xor XOR2 (N2028, N2005, N1131);
and AND3 (N2029, N2019, N1301, N1752);
or OR4 (N2030, N1994, N484, N1228, N1653);
not NOT1 (N2031, N2024);
and AND3 (N2032, N2031, N1818, N56);
xor XOR2 (N2033, N2021, N456);
nor NOR2 (N2034, N2028, N1407);
not NOT1 (N2035, N2026);
not NOT1 (N2036, N2020);
buf BUF1 (N2037, N2029);
or OR4 (N2038, N2030, N1792, N783, N159);
xor XOR2 (N2039, N2037, N29);
nor NOR2 (N2040, N2035, N225);
buf BUF1 (N2041, N2039);
not NOT1 (N2042, N2034);
nand NAND4 (N2043, N2022, N1686, N342, N1168);
buf BUF1 (N2044, N2027);
buf BUF1 (N2045, N2023);
not NOT1 (N2046, N2033);
nand NAND3 (N2047, N2041, N1941, N1435);
nor NOR3 (N2048, N2036, N1812, N1479);
nand NAND3 (N2049, N2043, N857, N1924);
nor NOR2 (N2050, N2047, N119);
not NOT1 (N2051, N2050);
or OR3 (N2052, N2042, N295, N1977);
or OR2 (N2053, N2045, N679);
xor XOR2 (N2054, N2052, N1002);
xor XOR2 (N2055, N2046, N992);
buf BUF1 (N2056, N2053);
and AND3 (N2057, N2032, N771, N1675);
and AND2 (N2058, N2054, N1765);
buf BUF1 (N2059, N2057);
nand NAND3 (N2060, N2038, N1664, N124);
nand NAND3 (N2061, N2059, N1815, N614);
or OR3 (N2062, N2056, N655, N947);
or OR4 (N2063, N2061, N147, N1295, N2042);
nand NAND3 (N2064, N2049, N974, N1270);
nor NOR3 (N2065, N2051, N1851, N850);
nor NOR4 (N2066, N2055, N1518, N187, N953);
buf BUF1 (N2067, N2063);
nor NOR4 (N2068, N2062, N274, N719, N541);
nand NAND3 (N2069, N2064, N756, N1098);
nor NOR4 (N2070, N2040, N518, N596, N1070);
nor NOR4 (N2071, N2060, N266, N443, N1218);
buf BUF1 (N2072, N2048);
buf BUF1 (N2073, N2065);
nand NAND2 (N2074, N2069, N1592);
buf BUF1 (N2075, N2072);
xor XOR2 (N2076, N2058, N1712);
or OR2 (N2077, N2068, N1663);
nor NOR4 (N2078, N2070, N246, N1683, N52);
and AND4 (N2079, N2044, N1291, N686, N540);
xor XOR2 (N2080, N2071, N158);
xor XOR2 (N2081, N2076, N171);
not NOT1 (N2082, N2079);
not NOT1 (N2083, N2081);
nand NAND2 (N2084, N2074, N2017);
buf BUF1 (N2085, N2083);
nor NOR2 (N2086, N2073, N1883);
not NOT1 (N2087, N2077);
xor XOR2 (N2088, N2067, N1542);
nor NOR2 (N2089, N2075, N95);
xor XOR2 (N2090, N2082, N648);
and AND3 (N2091, N2080, N1104, N1347);
xor XOR2 (N2092, N2087, N1383);
or OR4 (N2093, N2092, N1634, N1417, N1687);
buf BUF1 (N2094, N2066);
not NOT1 (N2095, N2093);
not NOT1 (N2096, N2090);
and AND4 (N2097, N2091, N1323, N766, N1228);
and AND3 (N2098, N2084, N703, N1770);
and AND3 (N2099, N2096, N1744, N1855);
nand NAND2 (N2100, N2078, N1104);
nor NOR4 (N2101, N2086, N1524, N454, N572);
nand NAND4 (N2102, N2088, N1301, N175, N937);
and AND4 (N2103, N2099, N850, N1372, N1512);
not NOT1 (N2104, N2102);
and AND4 (N2105, N2098, N1938, N1598, N220);
and AND4 (N2106, N2095, N960, N1435, N41);
and AND4 (N2107, N2089, N1104, N865, N2101);
and AND4 (N2108, N920, N1125, N1179, N612);
not NOT1 (N2109, N2100);
xor XOR2 (N2110, N2107, N972);
buf BUF1 (N2111, N2097);
nor NOR4 (N2112, N2085, N2105, N343, N1987);
not NOT1 (N2113, N459);
and AND2 (N2114, N2111, N582);
xor XOR2 (N2115, N2104, N13);
and AND2 (N2116, N2108, N455);
nand NAND4 (N2117, N2115, N723, N666, N808);
buf BUF1 (N2118, N2094);
and AND3 (N2119, N2110, N1657, N1018);
buf BUF1 (N2120, N2116);
and AND3 (N2121, N2120, N1000, N1847);
nor NOR2 (N2122, N2103, N509);
or OR4 (N2123, N2117, N299, N1811, N654);
nand NAND3 (N2124, N2114, N1956, N1588);
buf BUF1 (N2125, N2119);
xor XOR2 (N2126, N2113, N812);
xor XOR2 (N2127, N2126, N933);
or OR4 (N2128, N2127, N1528, N1890, N268);
nor NOR2 (N2129, N2123, N265);
and AND3 (N2130, N2124, N1097, N512);
and AND4 (N2131, N2130, N1949, N622, N1756);
or OR2 (N2132, N2112, N2046);
and AND2 (N2133, N2106, N2087);
xor XOR2 (N2134, N2131, N626);
nor NOR2 (N2135, N2133, N663);
not NOT1 (N2136, N2122);
not NOT1 (N2137, N2128);
nand NAND3 (N2138, N2132, N378, N948);
not NOT1 (N2139, N2134);
nand NAND3 (N2140, N2121, N2031, N1531);
buf BUF1 (N2141, N2139);
not NOT1 (N2142, N2109);
or OR4 (N2143, N2136, N249, N1108, N829);
and AND2 (N2144, N2118, N225);
buf BUF1 (N2145, N2142);
or OR2 (N2146, N2138, N1950);
nor NOR4 (N2147, N2146, N1114, N705, N1980);
xor XOR2 (N2148, N2143, N823);
not NOT1 (N2149, N2129);
or OR4 (N2150, N2140, N2048, N1093, N889);
and AND3 (N2151, N2148, N1027, N602);
not NOT1 (N2152, N2145);
buf BUF1 (N2153, N2135);
and AND2 (N2154, N2153, N320);
nand NAND3 (N2155, N2125, N1520, N868);
nand NAND3 (N2156, N2151, N1108, N724);
nand NAND4 (N2157, N2149, N2062, N775, N1117);
nand NAND2 (N2158, N2155, N382);
xor XOR2 (N2159, N2152, N1295);
xor XOR2 (N2160, N2144, N961);
and AND4 (N2161, N2156, N1948, N740, N542);
not NOT1 (N2162, N2137);
nand NAND4 (N2163, N2162, N1364, N691, N281);
or OR3 (N2164, N2154, N2050, N1759);
nand NAND3 (N2165, N2158, N1934, N1392);
buf BUF1 (N2166, N2159);
and AND2 (N2167, N2166, N1137);
not NOT1 (N2168, N2163);
buf BUF1 (N2169, N2141);
not NOT1 (N2170, N2147);
buf BUF1 (N2171, N2170);
nor NOR4 (N2172, N2168, N170, N1667, N8);
and AND3 (N2173, N2169, N936, N332);
nand NAND3 (N2174, N2173, N357, N269);
and AND2 (N2175, N2171, N1827);
buf BUF1 (N2176, N2165);
or OR2 (N2177, N2172, N1829);
nand NAND3 (N2178, N2167, N647, N435);
and AND4 (N2179, N2178, N937, N1692, N796);
nor NOR2 (N2180, N2176, N1594);
or OR3 (N2181, N2175, N1166, N1194);
and AND3 (N2182, N2160, N1223, N493);
not NOT1 (N2183, N2182);
or OR2 (N2184, N2174, N588);
not NOT1 (N2185, N2164);
buf BUF1 (N2186, N2161);
xor XOR2 (N2187, N2186, N1203);
xor XOR2 (N2188, N2185, N20);
nor NOR2 (N2189, N2184, N987);
not NOT1 (N2190, N2189);
buf BUF1 (N2191, N2177);
not NOT1 (N2192, N2191);
buf BUF1 (N2193, N2180);
xor XOR2 (N2194, N2157, N2162);
buf BUF1 (N2195, N2193);
nand NAND4 (N2196, N2150, N1874, N893, N744);
not NOT1 (N2197, N2195);
buf BUF1 (N2198, N2188);
nor NOR2 (N2199, N2197, N2120);
nand NAND2 (N2200, N2192, N1997);
nand NAND4 (N2201, N2200, N1723, N1513, N1611);
buf BUF1 (N2202, N2187);
buf BUF1 (N2203, N2202);
nor NOR3 (N2204, N2181, N2121, N2192);
nand NAND2 (N2205, N2203, N92);
not NOT1 (N2206, N2198);
nor NOR3 (N2207, N2194, N2054, N2111);
not NOT1 (N2208, N2190);
xor XOR2 (N2209, N2179, N929);
buf BUF1 (N2210, N2201);
not NOT1 (N2211, N2204);
nor NOR4 (N2212, N2207, N957, N1467, N1064);
xor XOR2 (N2213, N2183, N1775);
not NOT1 (N2214, N2212);
or OR4 (N2215, N2213, N943, N2106, N777);
xor XOR2 (N2216, N2205, N472);
nor NOR4 (N2217, N2196, N853, N1795, N1176);
xor XOR2 (N2218, N2211, N1475);
not NOT1 (N2219, N2215);
nand NAND2 (N2220, N2216, N163);
buf BUF1 (N2221, N2209);
xor XOR2 (N2222, N2210, N872);
nor NOR2 (N2223, N2208, N1580);
and AND3 (N2224, N2223, N1318, N2067);
nor NOR4 (N2225, N2222, N2175, N700, N1068);
buf BUF1 (N2226, N2206);
nor NOR4 (N2227, N2224, N471, N994, N1604);
nand NAND2 (N2228, N2199, N2165);
nand NAND3 (N2229, N2225, N1191, N1127);
buf BUF1 (N2230, N2226);
or OR2 (N2231, N2221, N2032);
and AND2 (N2232, N2227, N983);
not NOT1 (N2233, N2214);
not NOT1 (N2234, N2229);
nor NOR2 (N2235, N2219, N2067);
nor NOR3 (N2236, N2232, N231, N498);
buf BUF1 (N2237, N2236);
nand NAND3 (N2238, N2220, N791, N1179);
xor XOR2 (N2239, N2234, N1767);
and AND3 (N2240, N2217, N192, N183);
and AND2 (N2241, N2233, N1785);
not NOT1 (N2242, N2231);
or OR2 (N2243, N2242, N1163);
or OR2 (N2244, N2218, N431);
nand NAND3 (N2245, N2230, N1108, N1917);
or OR4 (N2246, N2238, N1878, N1805, N1364);
or OR4 (N2247, N2241, N643, N272, N1901);
nand NAND2 (N2248, N2244, N989);
xor XOR2 (N2249, N2237, N466);
not NOT1 (N2250, N2240);
or OR4 (N2251, N2243, N439, N1035, N53);
or OR4 (N2252, N2235, N149, N936, N1012);
nand NAND4 (N2253, N2247, N1405, N363, N1658);
or OR2 (N2254, N2239, N1976);
or OR4 (N2255, N2252, N439, N738, N713);
xor XOR2 (N2256, N2249, N1723);
xor XOR2 (N2257, N2248, N78);
or OR3 (N2258, N2257, N1235, N1804);
nor NOR3 (N2259, N2251, N1475, N836);
or OR2 (N2260, N2253, N2078);
nand NAND2 (N2261, N2245, N1342);
nand NAND4 (N2262, N2246, N440, N141, N1359);
nor NOR2 (N2263, N2256, N481);
not NOT1 (N2264, N2250);
and AND3 (N2265, N2228, N317, N1807);
not NOT1 (N2266, N2258);
nor NOR2 (N2267, N2254, N462);
buf BUF1 (N2268, N2255);
buf BUF1 (N2269, N2262);
nand NAND4 (N2270, N2264, N185, N844, N1535);
nor NOR2 (N2271, N2267, N1247);
buf BUF1 (N2272, N2268);
buf BUF1 (N2273, N2263);
not NOT1 (N2274, N2265);
buf BUF1 (N2275, N2266);
or OR4 (N2276, N2273, N1644, N1671, N479);
or OR4 (N2277, N2269, N818, N1160, N1761);
buf BUF1 (N2278, N2271);
xor XOR2 (N2279, N2277, N1555);
buf BUF1 (N2280, N2261);
nand NAND4 (N2281, N2279, N2154, N180, N2214);
not NOT1 (N2282, N2278);
xor XOR2 (N2283, N2260, N1489);
or OR4 (N2284, N2272, N1940, N1879, N1666);
nand NAND2 (N2285, N2284, N1076);
and AND2 (N2286, N2280, N1589);
xor XOR2 (N2287, N2283, N311);
nor NOR2 (N2288, N2270, N1863);
nand NAND4 (N2289, N2259, N1794, N2065, N2102);
or OR2 (N2290, N2288, N701);
xor XOR2 (N2291, N2289, N2019);
xor XOR2 (N2292, N2275, N2004);
and AND4 (N2293, N2282, N435, N731, N2126);
not NOT1 (N2294, N2292);
buf BUF1 (N2295, N2274);
xor XOR2 (N2296, N2285, N415);
buf BUF1 (N2297, N2290);
buf BUF1 (N2298, N2276);
buf BUF1 (N2299, N2295);
nand NAND3 (N2300, N2293, N1479, N1422);
buf BUF1 (N2301, N2287);
and AND3 (N2302, N2297, N1350, N1038);
and AND2 (N2303, N2286, N2125);
and AND4 (N2304, N2291, N1646, N1795, N1910);
and AND4 (N2305, N2304, N214, N1006, N972);
buf BUF1 (N2306, N2294);
buf BUF1 (N2307, N2301);
not NOT1 (N2308, N2303);
nand NAND4 (N2309, N2281, N1029, N1912, N991);
nor NOR3 (N2310, N2296, N1662, N1474);
and AND4 (N2311, N2299, N240, N210, N824);
not NOT1 (N2312, N2305);
or OR4 (N2313, N2306, N614, N1060, N2008);
nor NOR2 (N2314, N2312, N2041);
nor NOR2 (N2315, N2307, N2198);
buf BUF1 (N2316, N2314);
and AND3 (N2317, N2300, N1607, N1409);
or OR4 (N2318, N2310, N1593, N325, N1024);
buf BUF1 (N2319, N2318);
nand NAND4 (N2320, N2316, N1443, N1773, N1985);
not NOT1 (N2321, N2311);
xor XOR2 (N2322, N2320, N645);
and AND3 (N2323, N2315, N717, N1369);
nor NOR4 (N2324, N2322, N1022, N948, N2035);
and AND2 (N2325, N2308, N1414);
xor XOR2 (N2326, N2325, N281);
and AND3 (N2327, N2323, N524, N1687);
nor NOR4 (N2328, N2309, N70, N1512, N1783);
buf BUF1 (N2329, N2317);
or OR4 (N2330, N2321, N1214, N1972, N1975);
not NOT1 (N2331, N2298);
nand NAND4 (N2332, N2324, N1105, N691, N59);
and AND2 (N2333, N2331, N66);
not NOT1 (N2334, N2327);
not NOT1 (N2335, N2332);
not NOT1 (N2336, N2328);
and AND2 (N2337, N2333, N9);
nor NOR3 (N2338, N2329, N968, N1799);
buf BUF1 (N2339, N2338);
not NOT1 (N2340, N2339);
buf BUF1 (N2341, N2313);
xor XOR2 (N2342, N2337, N35);
buf BUF1 (N2343, N2340);
buf BUF1 (N2344, N2336);
xor XOR2 (N2345, N2302, N1258);
nor NOR2 (N2346, N2330, N2087);
and AND4 (N2347, N2342, N1185, N2123, N972);
nor NOR4 (N2348, N2344, N173, N2066, N1203);
nand NAND3 (N2349, N2343, N2177, N419);
or OR2 (N2350, N2335, N492);
nor NOR2 (N2351, N2334, N966);
not NOT1 (N2352, N2348);
nor NOR4 (N2353, N2345, N759, N1000, N467);
or OR4 (N2354, N2349, N1523, N372, N1529);
not NOT1 (N2355, N2353);
or OR2 (N2356, N2347, N283);
nor NOR2 (N2357, N2356, N1368);
nand NAND4 (N2358, N2350, N166, N2286, N2138);
nor NOR4 (N2359, N2346, N2261, N1661, N2222);
buf BUF1 (N2360, N2326);
nor NOR3 (N2361, N2354, N489, N1631);
or OR4 (N2362, N2361, N589, N576, N851);
not NOT1 (N2363, N2351);
buf BUF1 (N2364, N2358);
or OR4 (N2365, N2319, N952, N540, N72);
not NOT1 (N2366, N2352);
nand NAND2 (N2367, N2355, N867);
not NOT1 (N2368, N2362);
nand NAND3 (N2369, N2366, N1498, N644);
nand NAND2 (N2370, N2360, N373);
and AND2 (N2371, N2370, N590);
buf BUF1 (N2372, N2368);
nand NAND4 (N2373, N2364, N1804, N499, N1433);
and AND2 (N2374, N2341, N407);
and AND3 (N2375, N2367, N1957, N1008);
nor NOR2 (N2376, N2373, N1605);
not NOT1 (N2377, N2365);
buf BUF1 (N2378, N2377);
nand NAND2 (N2379, N2371, N2273);
xor XOR2 (N2380, N2375, N1918);
buf BUF1 (N2381, N2369);
xor XOR2 (N2382, N2357, N153);
or OR3 (N2383, N2363, N1761, N97);
not NOT1 (N2384, N2380);
nand NAND3 (N2385, N2382, N803, N828);
nor NOR4 (N2386, N2372, N999, N376, N2100);
and AND4 (N2387, N2385, N286, N52, N607);
xor XOR2 (N2388, N2359, N688);
and AND4 (N2389, N2374, N1210, N2099, N2322);
nand NAND3 (N2390, N2379, N231, N313);
nand NAND3 (N2391, N2376, N1696, N324);
buf BUF1 (N2392, N2389);
xor XOR2 (N2393, N2387, N2227);
not NOT1 (N2394, N2381);
nand NAND4 (N2395, N2390, N906, N271, N1111);
nand NAND3 (N2396, N2395, N1605, N1877);
not NOT1 (N2397, N2391);
not NOT1 (N2398, N2394);
nor NOR2 (N2399, N2396, N211);
buf BUF1 (N2400, N2399);
and AND4 (N2401, N2397, N1454, N1728, N1446);
or OR2 (N2402, N2401, N371);
xor XOR2 (N2403, N2384, N330);
nor NOR2 (N2404, N2392, N1192);
nand NAND4 (N2405, N2393, N1075, N1793, N1078);
buf BUF1 (N2406, N2378);
xor XOR2 (N2407, N2398, N1161);
nor NOR3 (N2408, N2406, N102, N2337);
nand NAND2 (N2409, N2404, N776);
xor XOR2 (N2410, N2405, N115);
nand NAND2 (N2411, N2386, N1061);
or OR4 (N2412, N2388, N2257, N2372, N1969);
nor NOR4 (N2413, N2400, N1251, N367, N1068);
xor XOR2 (N2414, N2402, N906);
and AND3 (N2415, N2403, N1645, N1984);
and AND2 (N2416, N2415, N199);
nand NAND4 (N2417, N2413, N1491, N1156, N813);
or OR2 (N2418, N2412, N1093);
and AND4 (N2419, N2408, N492, N1535, N1563);
or OR4 (N2420, N2414, N752, N307, N2030);
and AND3 (N2421, N2417, N31, N1969);
buf BUF1 (N2422, N2421);
nor NOR3 (N2423, N2383, N2303, N1419);
buf BUF1 (N2424, N2411);
buf BUF1 (N2425, N2424);
nor NOR3 (N2426, N2419, N2336, N1446);
nor NOR3 (N2427, N2410, N2287, N245);
nand NAND4 (N2428, N2416, N863, N507, N1252);
or OR4 (N2429, N2425, N966, N2251, N957);
xor XOR2 (N2430, N2420, N473);
not NOT1 (N2431, N2422);
nand NAND3 (N2432, N2429, N77, N174);
or OR4 (N2433, N2427, N2002, N981, N656);
buf BUF1 (N2434, N2428);
buf BUF1 (N2435, N2409);
buf BUF1 (N2436, N2433);
xor XOR2 (N2437, N2426, N203);
not NOT1 (N2438, N2432);
nand NAND4 (N2439, N2434, N2173, N2363, N1338);
xor XOR2 (N2440, N2439, N1109);
and AND2 (N2441, N2430, N738);
buf BUF1 (N2442, N2431);
nor NOR2 (N2443, N2438, N2255);
buf BUF1 (N2444, N2418);
nor NOR4 (N2445, N2436, N784, N118, N2415);
buf BUF1 (N2446, N2442);
xor XOR2 (N2447, N2435, N762);
and AND2 (N2448, N2437, N926);
xor XOR2 (N2449, N2444, N429);
not NOT1 (N2450, N2446);
xor XOR2 (N2451, N2449, N2411);
nor NOR2 (N2452, N2440, N1965);
nor NOR3 (N2453, N2407, N1202, N204);
buf BUF1 (N2454, N2447);
nand NAND3 (N2455, N2451, N1933, N1193);
not NOT1 (N2456, N2441);
nor NOR2 (N2457, N2453, N1517);
and AND4 (N2458, N2443, N1388, N739, N1419);
xor XOR2 (N2459, N2423, N743);
xor XOR2 (N2460, N2445, N1434);
xor XOR2 (N2461, N2454, N1645);
nand NAND2 (N2462, N2450, N1794);
nand NAND3 (N2463, N2457, N1592, N570);
or OR4 (N2464, N2455, N1269, N268, N138);
or OR4 (N2465, N2459, N1680, N1910, N856);
or OR4 (N2466, N2456, N2220, N2068, N1300);
nor NOR4 (N2467, N2463, N2056, N2263, N1159);
nand NAND2 (N2468, N2462, N180);
nor NOR4 (N2469, N2458, N1203, N1223, N6);
nand NAND3 (N2470, N2466, N501, N458);
not NOT1 (N2471, N2467);
buf BUF1 (N2472, N2468);
xor XOR2 (N2473, N2464, N1026);
not NOT1 (N2474, N2465);
not NOT1 (N2475, N2461);
nand NAND3 (N2476, N2452, N1637, N1212);
xor XOR2 (N2477, N2470, N831);
and AND3 (N2478, N2473, N1753, N2456);
nand NAND4 (N2479, N2474, N37, N763, N2051);
buf BUF1 (N2480, N2469);
not NOT1 (N2481, N2478);
nand NAND4 (N2482, N2460, N1301, N1815, N414);
not NOT1 (N2483, N2481);
nor NOR2 (N2484, N2471, N1550);
xor XOR2 (N2485, N2479, N55);
xor XOR2 (N2486, N2477, N927);
buf BUF1 (N2487, N2485);
nor NOR3 (N2488, N2484, N1688, N1302);
and AND4 (N2489, N2483, N1107, N2236, N1513);
or OR4 (N2490, N2475, N1353, N1858, N20);
xor XOR2 (N2491, N2482, N885);
not NOT1 (N2492, N2488);
xor XOR2 (N2493, N2480, N817);
or OR4 (N2494, N2448, N1621, N2216, N2329);
nor NOR2 (N2495, N2472, N361);
nand NAND2 (N2496, N2486, N1253);
or OR3 (N2497, N2489, N1889, N616);
xor XOR2 (N2498, N2487, N287);
or OR3 (N2499, N2495, N1113, N226);
and AND3 (N2500, N2491, N2148, N1254);
nor NOR3 (N2501, N2500, N2326, N1045);
nor NOR3 (N2502, N2493, N1181, N190);
not NOT1 (N2503, N2497);
xor XOR2 (N2504, N2498, N153);
or OR4 (N2505, N2476, N2138, N2224, N104);
xor XOR2 (N2506, N2490, N803);
nor NOR4 (N2507, N2506, N2280, N536, N257);
nor NOR3 (N2508, N2496, N1845, N557);
nand NAND3 (N2509, N2503, N2040, N779);
and AND4 (N2510, N2507, N1443, N1565, N1984);
and AND2 (N2511, N2510, N1613);
buf BUF1 (N2512, N2494);
and AND3 (N2513, N2505, N1714, N1013);
and AND2 (N2514, N2504, N2385);
xor XOR2 (N2515, N2499, N656);
nand NAND3 (N2516, N2492, N1002, N1750);
not NOT1 (N2517, N2513);
and AND3 (N2518, N2501, N896, N342);
buf BUF1 (N2519, N2518);
and AND2 (N2520, N2515, N1274);
not NOT1 (N2521, N2514);
buf BUF1 (N2522, N2521);
nor NOR2 (N2523, N2517, N2031);
and AND3 (N2524, N2523, N1467, N1847);
and AND3 (N2525, N2512, N1953, N962);
and AND2 (N2526, N2519, N2226);
and AND2 (N2527, N2520, N298);
nor NOR3 (N2528, N2511, N539, N820);
buf BUF1 (N2529, N2522);
nand NAND2 (N2530, N2508, N747);
and AND4 (N2531, N2525, N1288, N2078, N1218);
not NOT1 (N2532, N2502);
nor NOR4 (N2533, N2527, N1517, N326, N1041);
xor XOR2 (N2534, N2526, N2067);
or OR4 (N2535, N2509, N1766, N135, N2118);
buf BUF1 (N2536, N2516);
not NOT1 (N2537, N2532);
buf BUF1 (N2538, N2531);
buf BUF1 (N2539, N2535);
buf BUF1 (N2540, N2529);
nand NAND4 (N2541, N2538, N1623, N2424, N451);
and AND4 (N2542, N2534, N2378, N415, N1443);
or OR2 (N2543, N2524, N1512);
not NOT1 (N2544, N2537);
not NOT1 (N2545, N2533);
or OR2 (N2546, N2542, N1007);
or OR2 (N2547, N2536, N1446);
buf BUF1 (N2548, N2546);
nor NOR3 (N2549, N2539, N913, N257);
nand NAND4 (N2550, N2544, N1632, N2066, N457);
nor NOR4 (N2551, N2550, N2244, N293, N1744);
xor XOR2 (N2552, N2541, N1570);
not NOT1 (N2553, N2545);
or OR2 (N2554, N2548, N759);
and AND2 (N2555, N2543, N2271);
nor NOR2 (N2556, N2549, N1149);
or OR3 (N2557, N2553, N2147, N1325);
buf BUF1 (N2558, N2528);
nand NAND3 (N2559, N2551, N401, N2377);
and AND3 (N2560, N2559, N959, N1426);
xor XOR2 (N2561, N2552, N2084);
or OR4 (N2562, N2556, N1786, N583, N272);
nor NOR2 (N2563, N2554, N1418);
buf BUF1 (N2564, N2563);
buf BUF1 (N2565, N2564);
nor NOR3 (N2566, N2560, N1874, N2311);
xor XOR2 (N2567, N2530, N996);
xor XOR2 (N2568, N2547, N73);
not NOT1 (N2569, N2558);
nor NOR4 (N2570, N2561, N1162, N1884, N298);
and AND3 (N2571, N2566, N1595, N78);
nor NOR2 (N2572, N2567, N1970);
and AND3 (N2573, N2557, N1715, N7);
and AND2 (N2574, N2573, N2459);
nand NAND3 (N2575, N2565, N333, N171);
or OR2 (N2576, N2555, N2194);
nor NOR4 (N2577, N2571, N2495, N2274, N287);
buf BUF1 (N2578, N2575);
nor NOR4 (N2579, N2576, N2016, N2333, N370);
nand NAND3 (N2580, N2578, N2308, N109);
or OR2 (N2581, N2568, N628);
buf BUF1 (N2582, N2572);
and AND3 (N2583, N2577, N776, N1467);
xor XOR2 (N2584, N2583, N1740);
not NOT1 (N2585, N2580);
nand NAND2 (N2586, N2574, N1433);
or OR3 (N2587, N2579, N509, N2332);
or OR4 (N2588, N2540, N1416, N1793, N1523);
and AND3 (N2589, N2570, N1300, N882);
nand NAND4 (N2590, N2589, N1803, N66, N514);
nand NAND4 (N2591, N2582, N2541, N2073, N2461);
xor XOR2 (N2592, N2588, N15);
or OR2 (N2593, N2584, N2121);
nor NOR3 (N2594, N2562, N864, N2332);
not NOT1 (N2595, N2590);
buf BUF1 (N2596, N2569);
nand NAND4 (N2597, N2595, N2431, N504, N188);
buf BUF1 (N2598, N2596);
or OR4 (N2599, N2597, N1175, N271, N194);
buf BUF1 (N2600, N2598);
and AND4 (N2601, N2587, N2055, N2184, N221);
xor XOR2 (N2602, N2599, N770);
nand NAND3 (N2603, N2601, N2300, N2239);
not NOT1 (N2604, N2602);
and AND2 (N2605, N2600, N2190);
or OR2 (N2606, N2585, N124);
buf BUF1 (N2607, N2591);
buf BUF1 (N2608, N2586);
buf BUF1 (N2609, N2603);
or OR2 (N2610, N2605, N310);
xor XOR2 (N2611, N2610, N1362);
or OR4 (N2612, N2592, N157, N1396, N1246);
nor NOR3 (N2613, N2606, N1022, N357);
xor XOR2 (N2614, N2611, N1259);
buf BUF1 (N2615, N2608);
not NOT1 (N2616, N2593);
nand NAND2 (N2617, N2615, N1584);
or OR4 (N2618, N2617, N1230, N2101, N278);
not NOT1 (N2619, N2609);
not NOT1 (N2620, N2619);
or OR4 (N2621, N2612, N2222, N112, N96);
or OR2 (N2622, N2621, N103);
nand NAND2 (N2623, N2581, N629);
nand NAND4 (N2624, N2618, N1017, N419, N373);
buf BUF1 (N2625, N2614);
and AND3 (N2626, N2624, N2085, N1759);
nor NOR4 (N2627, N2616, N1373, N2006, N1800);
not NOT1 (N2628, N2620);
or OR4 (N2629, N2604, N2286, N2515, N2378);
nor NOR2 (N2630, N2628, N2522);
not NOT1 (N2631, N2623);
nand NAND2 (N2632, N2594, N2358);
nor NOR3 (N2633, N2629, N1592, N1058);
not NOT1 (N2634, N2632);
or OR3 (N2635, N2633, N375, N2310);
nand NAND2 (N2636, N2613, N958);
not NOT1 (N2637, N2607);
nand NAND3 (N2638, N2627, N2583, N349);
or OR4 (N2639, N2637, N1935, N2173, N535);
xor XOR2 (N2640, N2636, N1147);
not NOT1 (N2641, N2638);
nor NOR2 (N2642, N2622, N797);
not NOT1 (N2643, N2625);
xor XOR2 (N2644, N2640, N289);
buf BUF1 (N2645, N2643);
xor XOR2 (N2646, N2634, N1039);
buf BUF1 (N2647, N2626);
nand NAND3 (N2648, N2641, N2073, N1697);
not NOT1 (N2649, N2646);
not NOT1 (N2650, N2630);
nand NAND4 (N2651, N2635, N1470, N1498, N1043);
xor XOR2 (N2652, N2639, N2096);
nor NOR3 (N2653, N2645, N1303, N2439);
nor NOR3 (N2654, N2651, N1097, N2311);
buf BUF1 (N2655, N2650);
and AND3 (N2656, N2642, N2389, N2063);
or OR3 (N2657, N2649, N887, N2112);
nand NAND4 (N2658, N2656, N652, N1837, N1761);
buf BUF1 (N2659, N2657);
not NOT1 (N2660, N2648);
xor XOR2 (N2661, N2659, N69);
not NOT1 (N2662, N2647);
xor XOR2 (N2663, N2661, N1370);
nor NOR4 (N2664, N2660, N2642, N698, N1544);
nand NAND4 (N2665, N2664, N2047, N1955, N562);
buf BUF1 (N2666, N2655);
nor NOR2 (N2667, N2631, N182);
buf BUF1 (N2668, N2665);
xor XOR2 (N2669, N2663, N556);
or OR2 (N2670, N2662, N72);
nor NOR3 (N2671, N2667, N2140, N2513);
nand NAND2 (N2672, N2658, N480);
nand NAND2 (N2673, N2669, N1125);
xor XOR2 (N2674, N2644, N2664);
and AND3 (N2675, N2654, N698, N1192);
not NOT1 (N2676, N2674);
xor XOR2 (N2677, N2671, N2121);
xor XOR2 (N2678, N2676, N2145);
not NOT1 (N2679, N2653);
nor NOR3 (N2680, N2679, N361, N983);
not NOT1 (N2681, N2666);
nand NAND2 (N2682, N2678, N61);
and AND2 (N2683, N2670, N2437);
nor NOR3 (N2684, N2668, N741, N1941);
xor XOR2 (N2685, N2682, N1690);
not NOT1 (N2686, N2685);
nor NOR2 (N2687, N2686, N822);
nor NOR2 (N2688, N2680, N1230);
and AND4 (N2689, N2672, N1477, N1531, N595);
xor XOR2 (N2690, N2681, N1119);
and AND3 (N2691, N2673, N801, N2078);
buf BUF1 (N2692, N2690);
xor XOR2 (N2693, N2692, N2036);
and AND3 (N2694, N2677, N1067, N475);
not NOT1 (N2695, N2683);
nor NOR3 (N2696, N2684, N1933, N716);
xor XOR2 (N2697, N2693, N308);
buf BUF1 (N2698, N2688);
and AND2 (N2699, N2695, N250);
xor XOR2 (N2700, N2697, N686);
nor NOR2 (N2701, N2699, N1745);
and AND4 (N2702, N2696, N203, N560, N604);
xor XOR2 (N2703, N2652, N2253);
nand NAND2 (N2704, N2675, N2629);
or OR2 (N2705, N2689, N1757);
or OR2 (N2706, N2704, N1676);
not NOT1 (N2707, N2706);
and AND3 (N2708, N2700, N915, N1648);
nand NAND3 (N2709, N2691, N1436, N2600);
or OR2 (N2710, N2702, N979);
xor XOR2 (N2711, N2709, N1166);
buf BUF1 (N2712, N2701);
xor XOR2 (N2713, N2707, N2230);
and AND3 (N2714, N2711, N2121, N202);
or OR3 (N2715, N2708, N2286, N1465);
or OR4 (N2716, N2687, N191, N1580, N751);
nand NAND2 (N2717, N2712, N1586);
and AND4 (N2718, N2717, N1963, N2146, N1375);
not NOT1 (N2719, N2715);
nand NAND4 (N2720, N2713, N393, N1318, N473);
buf BUF1 (N2721, N2710);
buf BUF1 (N2722, N2720);
nand NAND3 (N2723, N2694, N1805, N1366);
and AND4 (N2724, N2721, N1774, N137, N215);
nand NAND3 (N2725, N2722, N348, N2638);
nand NAND3 (N2726, N2698, N1694, N2232);
and AND2 (N2727, N2719, N606);
buf BUF1 (N2728, N2718);
and AND4 (N2729, N2724, N2647, N1077, N2313);
or OR2 (N2730, N2703, N824);
and AND2 (N2731, N2729, N637);
nand NAND2 (N2732, N2731, N571);
or OR2 (N2733, N2728, N1474);
nor NOR3 (N2734, N2723, N1503, N1555);
buf BUF1 (N2735, N2734);
not NOT1 (N2736, N2725);
not NOT1 (N2737, N2730);
or OR2 (N2738, N2726, N2456);
nand NAND3 (N2739, N2716, N13, N2264);
nor NOR3 (N2740, N2727, N1394, N996);
nor NOR3 (N2741, N2737, N935, N1399);
and AND4 (N2742, N2714, N1599, N1735, N1537);
and AND4 (N2743, N2705, N2379, N1101, N1446);
buf BUF1 (N2744, N2735);
nand NAND4 (N2745, N2744, N1729, N1248, N1785);
and AND4 (N2746, N2745, N1558, N654, N311);
or OR3 (N2747, N2739, N411, N1369);
nand NAND2 (N2748, N2743, N1728);
or OR4 (N2749, N2748, N2297, N2060, N2435);
and AND3 (N2750, N2742, N2213, N227);
nor NOR4 (N2751, N2736, N1871, N1630, N1701);
not NOT1 (N2752, N2732);
or OR3 (N2753, N2747, N1488, N776);
xor XOR2 (N2754, N2733, N1506);
and AND2 (N2755, N2746, N401);
nor NOR3 (N2756, N2741, N809, N2392);
nand NAND4 (N2757, N2738, N474, N702, N1457);
and AND4 (N2758, N2757, N704, N2386, N79);
xor XOR2 (N2759, N2750, N429);
and AND3 (N2760, N2756, N619, N1599);
nand NAND2 (N2761, N2740, N371);
xor XOR2 (N2762, N2753, N537);
and AND2 (N2763, N2749, N1535);
nand NAND3 (N2764, N2760, N1527, N394);
or OR3 (N2765, N2758, N1863, N1480);
nand NAND4 (N2766, N2765, N317, N1147, N1862);
and AND4 (N2767, N2755, N719, N194, N562);
nand NAND2 (N2768, N2754, N581);
xor XOR2 (N2769, N2764, N1154);
xor XOR2 (N2770, N2761, N1148);
not NOT1 (N2771, N2766);
not NOT1 (N2772, N2751);
nor NOR4 (N2773, N2771, N1966, N2441, N1900);
nand NAND2 (N2774, N2773, N1884);
buf BUF1 (N2775, N2759);
or OR3 (N2776, N2763, N2514, N458);
xor XOR2 (N2777, N2752, N697);
and AND2 (N2778, N2768, N525);
buf BUF1 (N2779, N2769);
and AND3 (N2780, N2776, N2435, N2237);
xor XOR2 (N2781, N2762, N1543);
nor NOR4 (N2782, N2767, N569, N1621, N514);
or OR2 (N2783, N2775, N2347);
xor XOR2 (N2784, N2770, N1264);
nand NAND4 (N2785, N2774, N1904, N1432, N1492);
not NOT1 (N2786, N2778);
buf BUF1 (N2787, N2772);
nor NOR4 (N2788, N2782, N1978, N1043, N116);
buf BUF1 (N2789, N2788);
nor NOR2 (N2790, N2785, N273);
xor XOR2 (N2791, N2777, N2053);
nor NOR2 (N2792, N2779, N2040);
xor XOR2 (N2793, N2786, N84);
not NOT1 (N2794, N2781);
and AND4 (N2795, N2787, N1259, N2754, N871);
not NOT1 (N2796, N2793);
or OR3 (N2797, N2783, N2339, N1217);
buf BUF1 (N2798, N2794);
or OR2 (N2799, N2796, N1370);
nor NOR4 (N2800, N2797, N1837, N1926, N1875);
not NOT1 (N2801, N2800);
nand NAND3 (N2802, N2791, N392, N222);
not NOT1 (N2803, N2798);
not NOT1 (N2804, N2799);
nor NOR2 (N2805, N2803, N2017);
xor XOR2 (N2806, N2789, N243);
nand NAND3 (N2807, N2784, N2802, N2086);
nor NOR4 (N2808, N1219, N765, N233, N2517);
xor XOR2 (N2809, N2804, N1375);
and AND4 (N2810, N2790, N21, N89, N2670);
or OR4 (N2811, N2807, N1636, N2405, N1678);
and AND4 (N2812, N2806, N1501, N362, N57);
or OR2 (N2813, N2801, N815);
xor XOR2 (N2814, N2812, N248);
nor NOR4 (N2815, N2780, N533, N2432, N2614);
and AND2 (N2816, N2792, N481);
nand NAND2 (N2817, N2815, N30);
not NOT1 (N2818, N2817);
buf BUF1 (N2819, N2808);
nor NOR2 (N2820, N2814, N282);
buf BUF1 (N2821, N2795);
not NOT1 (N2822, N2821);
or OR4 (N2823, N2810, N2786, N358, N2090);
not NOT1 (N2824, N2822);
and AND3 (N2825, N2811, N1057, N1825);
nand NAND2 (N2826, N2819, N2364);
not NOT1 (N2827, N2824);
nor NOR3 (N2828, N2805, N64, N2694);
and AND2 (N2829, N2813, N2248);
nor NOR4 (N2830, N2823, N1161, N2178, N17);
nand NAND2 (N2831, N2820, N1712);
nand NAND3 (N2832, N2818, N2313, N43);
and AND3 (N2833, N2809, N2627, N117);
nor NOR2 (N2834, N2830, N974);
not NOT1 (N2835, N2834);
buf BUF1 (N2836, N2827);
and AND2 (N2837, N2836, N376);
buf BUF1 (N2838, N2828);
nand NAND4 (N2839, N2838, N1957, N402, N1709);
and AND2 (N2840, N2837, N1104);
and AND3 (N2841, N2832, N1954, N1839);
nor NOR4 (N2842, N2840, N971, N1678, N2480);
nor NOR4 (N2843, N2829, N2545, N1709, N417);
and AND3 (N2844, N2833, N2804, N1634);
and AND3 (N2845, N2842, N366, N452);
not NOT1 (N2846, N2844);
buf BUF1 (N2847, N2831);
nor NOR3 (N2848, N2839, N753, N190);
xor XOR2 (N2849, N2835, N458);
xor XOR2 (N2850, N2841, N2354);
nor NOR3 (N2851, N2843, N2182, N754);
not NOT1 (N2852, N2848);
xor XOR2 (N2853, N2845, N1757);
buf BUF1 (N2854, N2826);
xor XOR2 (N2855, N2850, N665);
and AND3 (N2856, N2816, N444, N764);
nand NAND3 (N2857, N2851, N2439, N458);
nand NAND3 (N2858, N2847, N387, N534);
not NOT1 (N2859, N2852);
xor XOR2 (N2860, N2856, N1607);
xor XOR2 (N2861, N2859, N500);
and AND2 (N2862, N2858, N2550);
nor NOR3 (N2863, N2846, N1694, N2070);
nor NOR2 (N2864, N2825, N2225);
nor NOR2 (N2865, N2860, N2277);
buf BUF1 (N2866, N2865);
nand NAND2 (N2867, N2857, N720);
not NOT1 (N2868, N2849);
or OR4 (N2869, N2867, N1786, N346, N1809);
not NOT1 (N2870, N2853);
nand NAND2 (N2871, N2869, N1015);
nand NAND4 (N2872, N2861, N2564, N345, N717);
not NOT1 (N2873, N2871);
not NOT1 (N2874, N2863);
buf BUF1 (N2875, N2872);
and AND4 (N2876, N2866, N2606, N219, N1202);
not NOT1 (N2877, N2870);
or OR4 (N2878, N2868, N2104, N676, N1432);
or OR4 (N2879, N2873, N2708, N1838, N2472);
buf BUF1 (N2880, N2864);
xor XOR2 (N2881, N2877, N2826);
nor NOR4 (N2882, N2878, N1617, N908, N2875);
and AND2 (N2883, N1753, N2015);
xor XOR2 (N2884, N2881, N2652);
nor NOR3 (N2885, N2883, N879, N1773);
or OR4 (N2886, N2855, N2369, N1802, N1597);
nand NAND3 (N2887, N2854, N442, N1574);
and AND4 (N2888, N2862, N2320, N421, N2713);
and AND4 (N2889, N2876, N1937, N2542, N2666);
or OR4 (N2890, N2886, N1925, N2392, N236);
nand NAND4 (N2891, N2882, N1658, N898, N97);
xor XOR2 (N2892, N2879, N721);
xor XOR2 (N2893, N2874, N1218);
nand NAND2 (N2894, N2891, N142);
nor NOR4 (N2895, N2885, N157, N240, N114);
nand NAND4 (N2896, N2893, N1821, N2339, N461);
nand NAND3 (N2897, N2889, N2155, N2859);
xor XOR2 (N2898, N2880, N2718);
or OR3 (N2899, N2896, N2694, N2030);
or OR3 (N2900, N2895, N1984, N2406);
or OR3 (N2901, N2892, N2861, N891);
nor NOR3 (N2902, N2901, N837, N572);
nor NOR2 (N2903, N2898, N2673);
and AND2 (N2904, N2887, N2415);
buf BUF1 (N2905, N2899);
not NOT1 (N2906, N2894);
buf BUF1 (N2907, N2884);
nand NAND2 (N2908, N2907, N1898);
buf BUF1 (N2909, N2897);
nand NAND2 (N2910, N2902, N2573);
and AND3 (N2911, N2910, N857, N509);
and AND3 (N2912, N2888, N2740, N450);
or OR2 (N2913, N2903, N2022);
buf BUF1 (N2914, N2900);
nor NOR4 (N2915, N2904, N2414, N179, N2305);
nor NOR4 (N2916, N2890, N111, N1907, N1418);
nand NAND3 (N2917, N2915, N2845, N1203);
not NOT1 (N2918, N2909);
not NOT1 (N2919, N2908);
not NOT1 (N2920, N2916);
or OR3 (N2921, N2919, N1928, N2534);
xor XOR2 (N2922, N2906, N40);
and AND3 (N2923, N2914, N1436, N2145);
buf BUF1 (N2924, N2923);
buf BUF1 (N2925, N2911);
nor NOR3 (N2926, N2921, N838, N573);
and AND4 (N2927, N2912, N637, N564, N2253);
buf BUF1 (N2928, N2917);
or OR3 (N2929, N2913, N2109, N2497);
xor XOR2 (N2930, N2927, N1518);
not NOT1 (N2931, N2918);
xor XOR2 (N2932, N2931, N2642);
nand NAND3 (N2933, N2929, N721, N2387);
nor NOR3 (N2934, N2928, N1341, N68);
buf BUF1 (N2935, N2933);
buf BUF1 (N2936, N2924);
xor XOR2 (N2937, N2925, N882);
and AND3 (N2938, N2905, N560, N1061);
xor XOR2 (N2939, N2922, N1269);
xor XOR2 (N2940, N2926, N585);
and AND4 (N2941, N2934, N230, N464, N2004);
nand NAND3 (N2942, N2920, N2386, N189);
and AND3 (N2943, N2932, N474, N1056);
or OR2 (N2944, N2941, N1949);
not NOT1 (N2945, N2942);
nand NAND2 (N2946, N2937, N1091);
not NOT1 (N2947, N2946);
not NOT1 (N2948, N2930);
and AND4 (N2949, N2947, N1611, N2462, N1082);
nor NOR4 (N2950, N2939, N69, N927, N1136);
xor XOR2 (N2951, N2944, N2066);
or OR4 (N2952, N2940, N2780, N265, N487);
nand NAND2 (N2953, N2943, N381);
xor XOR2 (N2954, N2936, N145);
nand NAND3 (N2955, N2949, N133, N617);
or OR3 (N2956, N2950, N367, N1858);
not NOT1 (N2957, N2954);
or OR2 (N2958, N2938, N615);
not NOT1 (N2959, N2956);
or OR4 (N2960, N2953, N222, N734, N2089);
and AND3 (N2961, N2959, N651, N1193);
or OR3 (N2962, N2945, N1750, N1205);
and AND4 (N2963, N2952, N1136, N1361, N1710);
nand NAND3 (N2964, N2961, N1328, N813);
nor NOR3 (N2965, N2963, N1516, N1834);
nand NAND4 (N2966, N2957, N1010, N489, N2660);
nand NAND4 (N2967, N2955, N750, N48, N1567);
nor NOR3 (N2968, N2962, N699, N2007);
or OR2 (N2969, N2967, N771);
or OR2 (N2970, N2968, N2325);
xor XOR2 (N2971, N2966, N696);
not NOT1 (N2972, N2971);
nand NAND4 (N2973, N2972, N158, N1265, N2336);
or OR2 (N2974, N2969, N1504);
not NOT1 (N2975, N2951);
not NOT1 (N2976, N2964);
or OR4 (N2977, N2974, N1363, N2627, N2521);
buf BUF1 (N2978, N2958);
not NOT1 (N2979, N2976);
xor XOR2 (N2980, N2978, N535);
not NOT1 (N2981, N2965);
nor NOR4 (N2982, N2979, N673, N934, N1134);
buf BUF1 (N2983, N2977);
or OR2 (N2984, N2970, N2480);
buf BUF1 (N2985, N2982);
nand NAND3 (N2986, N2981, N329, N1744);
xor XOR2 (N2987, N2960, N1370);
buf BUF1 (N2988, N2986);
nand NAND4 (N2989, N2980, N2431, N2861, N567);
nor NOR4 (N2990, N2948, N2771, N1558, N1691);
and AND2 (N2991, N2975, N32);
nor NOR4 (N2992, N2987, N2542, N1614, N2929);
nor NOR4 (N2993, N2983, N845, N1915, N1886);
or OR4 (N2994, N2993, N2406, N2965, N2556);
nor NOR4 (N2995, N2994, N1646, N1875, N962);
and AND4 (N2996, N2995, N378, N1175, N771);
buf BUF1 (N2997, N2991);
not NOT1 (N2998, N2973);
and AND3 (N2999, N2990, N334, N419);
buf BUF1 (N3000, N2998);
and AND3 (N3001, N2984, N346, N328);
and AND4 (N3002, N2999, N1290, N2577, N37);
not NOT1 (N3003, N2935);
nor NOR3 (N3004, N2989, N2055, N2209);
nand NAND4 (N3005, N3004, N2766, N2329, N2998);
xor XOR2 (N3006, N2992, N1227);
nor NOR3 (N3007, N3000, N1722, N1119);
buf BUF1 (N3008, N3002);
nand NAND2 (N3009, N2997, N760);
nand NAND4 (N3010, N2985, N362, N2324, N1992);
or OR2 (N3011, N3001, N2254);
and AND4 (N3012, N2988, N2941, N2809, N807);
xor XOR2 (N3013, N3005, N2737);
or OR4 (N3014, N3011, N2662, N2215, N1716);
and AND3 (N3015, N3006, N1205, N379);
xor XOR2 (N3016, N3010, N757);
or OR4 (N3017, N3016, N2227, N2001, N1552);
not NOT1 (N3018, N3009);
not NOT1 (N3019, N3013);
xor XOR2 (N3020, N2996, N999);
and AND2 (N3021, N3020, N1214);
nand NAND2 (N3022, N3018, N147);
and AND4 (N3023, N3019, N2272, N4, N2548);
buf BUF1 (N3024, N3015);
not NOT1 (N3025, N3023);
nand NAND2 (N3026, N3012, N1333);
buf BUF1 (N3027, N3008);
or OR3 (N3028, N3022, N1314, N2091);
and AND4 (N3029, N3027, N2155, N1986, N2154);
nor NOR3 (N3030, N3007, N1971, N420);
or OR2 (N3031, N3030, N1071);
nand NAND4 (N3032, N3026, N87, N1966, N54);
nor NOR3 (N3033, N3021, N2849, N1972);
xor XOR2 (N3034, N3033, N2339);
and AND2 (N3035, N3031, N651);
buf BUF1 (N3036, N3034);
nand NAND2 (N3037, N3025, N2772);
nor NOR3 (N3038, N3029, N622, N1005);
xor XOR2 (N3039, N3028, N1961);
nand NAND3 (N3040, N3037, N541, N3026);
buf BUF1 (N3041, N3038);
not NOT1 (N3042, N3040);
not NOT1 (N3043, N3032);
nor NOR3 (N3044, N3036, N2204, N208);
xor XOR2 (N3045, N3044, N510);
or OR2 (N3046, N3039, N2724);
nor NOR4 (N3047, N3042, N604, N1673, N396);
nor NOR2 (N3048, N3045, N2176);
nor NOR4 (N3049, N3014, N2477, N570, N1632);
xor XOR2 (N3050, N3049, N292);
buf BUF1 (N3051, N3035);
not NOT1 (N3052, N3050);
or OR4 (N3053, N3043, N944, N1695, N2225);
nor NOR2 (N3054, N3048, N335);
xor XOR2 (N3055, N3047, N1427);
and AND4 (N3056, N3017, N2161, N2694, N2216);
xor XOR2 (N3057, N3024, N922);
not NOT1 (N3058, N3055);
buf BUF1 (N3059, N3054);
xor XOR2 (N3060, N3051, N1639);
or OR4 (N3061, N3060, N1905, N1812, N1093);
nor NOR2 (N3062, N3046, N1139);
nor NOR3 (N3063, N3059, N2183, N995);
nand NAND4 (N3064, N3062, N2789, N2842, N666);
nand NAND4 (N3065, N3064, N773, N706, N2324);
and AND4 (N3066, N3063, N306, N1762, N699);
nor NOR4 (N3067, N3065, N392, N2061, N1922);
and AND2 (N3068, N3003, N848);
and AND2 (N3069, N3056, N1214);
and AND3 (N3070, N3052, N11, N2543);
xor XOR2 (N3071, N3069, N678);
not NOT1 (N3072, N3070);
and AND4 (N3073, N3057, N2015, N3010, N1059);
and AND3 (N3074, N3071, N1109, N2861);
not NOT1 (N3075, N3074);
or OR4 (N3076, N3058, N310, N2215, N2846);
nand NAND3 (N3077, N3068, N2266, N1004);
nor NOR4 (N3078, N3076, N1051, N837, N1087);
nor NOR3 (N3079, N3066, N1001, N1977);
buf BUF1 (N3080, N3077);
nor NOR4 (N3081, N3067, N1705, N88, N1160);
xor XOR2 (N3082, N3080, N241);
buf BUF1 (N3083, N3072);
buf BUF1 (N3084, N3082);
or OR3 (N3085, N3053, N1086, N2753);
nor NOR4 (N3086, N3085, N244, N2315, N597);
not NOT1 (N3087, N3061);
not NOT1 (N3088, N3084);
xor XOR2 (N3089, N3083, N336);
nor NOR4 (N3090, N3041, N2222, N1502, N2166);
buf BUF1 (N3091, N3086);
xor XOR2 (N3092, N3078, N2832);
nand NAND3 (N3093, N3091, N894, N2414);
buf BUF1 (N3094, N3087);
not NOT1 (N3095, N3088);
not NOT1 (N3096, N3095);
nand NAND3 (N3097, N3094, N3089, N2976);
buf BUF1 (N3098, N2264);
xor XOR2 (N3099, N3092, N901);
not NOT1 (N3100, N3075);
nand NAND2 (N3101, N3081, N2043);
xor XOR2 (N3102, N3100, N132);
nor NOR2 (N3103, N3073, N414);
xor XOR2 (N3104, N3097, N2682);
or OR4 (N3105, N3090, N92, N2306, N3008);
or OR3 (N3106, N3101, N59, N1193);
xor XOR2 (N3107, N3106, N1801);
and AND4 (N3108, N3107, N1628, N1046, N1764);
not NOT1 (N3109, N3079);
nor NOR4 (N3110, N3105, N1473, N992, N677);
buf BUF1 (N3111, N3093);
xor XOR2 (N3112, N3108, N3014);
and AND3 (N3113, N3098, N788, N2677);
not NOT1 (N3114, N3096);
nor NOR4 (N3115, N3104, N2867, N1141, N269);
and AND4 (N3116, N3111, N2210, N443, N27);
not NOT1 (N3117, N3115);
and AND4 (N3118, N3117, N2933, N211, N2927);
not NOT1 (N3119, N3109);
xor XOR2 (N3120, N3114, N974);
nand NAND2 (N3121, N3099, N1938);
and AND4 (N3122, N3102, N1438, N1866, N133);
nand NAND4 (N3123, N3118, N1849, N2886, N1154);
nand NAND4 (N3124, N3121, N215, N2898, N1532);
buf BUF1 (N3125, N3124);
and AND3 (N3126, N3125, N1398, N1246);
nor NOR4 (N3127, N3103, N462, N471, N616);
xor XOR2 (N3128, N3110, N757);
not NOT1 (N3129, N3123);
xor XOR2 (N3130, N3126, N181);
not NOT1 (N3131, N3129);
nor NOR2 (N3132, N3131, N186);
not NOT1 (N3133, N3112);
and AND4 (N3134, N3119, N1130, N801, N2995);
not NOT1 (N3135, N3128);
xor XOR2 (N3136, N3127, N784);
buf BUF1 (N3137, N3113);
buf BUF1 (N3138, N3135);
and AND3 (N3139, N3134, N1870, N1933);
and AND3 (N3140, N3133, N2478, N1749);
nand NAND4 (N3141, N3122, N737, N1223, N1948);
and AND4 (N3142, N3138, N1127, N2104, N2237);
nand NAND2 (N3143, N3140, N2646);
xor XOR2 (N3144, N3137, N2203);
and AND3 (N3145, N3141, N1540, N2226);
buf BUF1 (N3146, N3144);
buf BUF1 (N3147, N3145);
nand NAND2 (N3148, N3143, N171);
buf BUF1 (N3149, N3147);
nor NOR3 (N3150, N3116, N1543, N1006);
not NOT1 (N3151, N3139);
not NOT1 (N3152, N3148);
nand NAND2 (N3153, N3132, N766);
nand NAND3 (N3154, N3142, N731, N2030);
or OR4 (N3155, N3136, N1187, N977, N1802);
not NOT1 (N3156, N3120);
or OR3 (N3157, N3153, N122, N2031);
xor XOR2 (N3158, N3149, N2994);
buf BUF1 (N3159, N3146);
not NOT1 (N3160, N3150);
xor XOR2 (N3161, N3155, N942);
not NOT1 (N3162, N3160);
not NOT1 (N3163, N3161);
nor NOR3 (N3164, N3162, N2822, N270);
buf BUF1 (N3165, N3151);
and AND4 (N3166, N3154, N999, N2941, N265);
nor NOR2 (N3167, N3158, N2652);
nand NAND3 (N3168, N3163, N3158, N1406);
xor XOR2 (N3169, N3164, N1871);
or OR2 (N3170, N3130, N1014);
buf BUF1 (N3171, N3165);
and AND4 (N3172, N3156, N1904, N1225, N2294);
nand NAND4 (N3173, N3159, N2492, N166, N2755);
and AND3 (N3174, N3168, N1273, N608);
not NOT1 (N3175, N3170);
nor NOR2 (N3176, N3169, N1392);
buf BUF1 (N3177, N3172);
or OR3 (N3178, N3174, N95, N2149);
and AND3 (N3179, N3173, N1067, N424);
not NOT1 (N3180, N3177);
and AND2 (N3181, N3171, N437);
nand NAND3 (N3182, N3181, N2636, N2894);
and AND2 (N3183, N3179, N2026);
nor NOR2 (N3184, N3152, N445);
nand NAND3 (N3185, N3175, N3104, N2755);
not NOT1 (N3186, N3167);
buf BUF1 (N3187, N3166);
not NOT1 (N3188, N3176);
buf BUF1 (N3189, N3183);
and AND3 (N3190, N3180, N1881, N2614);
nand NAND2 (N3191, N3178, N1521);
or OR3 (N3192, N3187, N951, N2581);
and AND3 (N3193, N3184, N2370, N1993);
nand NAND2 (N3194, N3189, N3013);
nand NAND4 (N3195, N3191, N1953, N1652, N1984);
nand NAND2 (N3196, N3185, N2400);
and AND3 (N3197, N3190, N2056, N1142);
nand NAND4 (N3198, N3157, N2097, N118, N2109);
nand NAND3 (N3199, N3192, N2814, N1202);
xor XOR2 (N3200, N3182, N1431);
nor NOR4 (N3201, N3196, N3107, N2181, N2407);
buf BUF1 (N3202, N3193);
buf BUF1 (N3203, N3200);
nand NAND3 (N3204, N3186, N414, N1431);
nor NOR3 (N3205, N3203, N2304, N854);
buf BUF1 (N3206, N3202);
nand NAND4 (N3207, N3198, N2489, N34, N274);
nor NOR3 (N3208, N3199, N76, N1034);
or OR2 (N3209, N3206, N353);
and AND4 (N3210, N3201, N1005, N479, N2265);
or OR2 (N3211, N3195, N2817);
nand NAND2 (N3212, N3211, N3159);
or OR4 (N3213, N3209, N2964, N2000, N423);
and AND2 (N3214, N3188, N910);
and AND3 (N3215, N3197, N811, N1279);
buf BUF1 (N3216, N3207);
nor NOR3 (N3217, N3194, N2672, N2059);
or OR3 (N3218, N3208, N529, N2469);
xor XOR2 (N3219, N3218, N438);
and AND4 (N3220, N3212, N1884, N2863, N3041);
xor XOR2 (N3221, N3205, N896);
xor XOR2 (N3222, N3210, N1166);
or OR2 (N3223, N3216, N1671);
or OR4 (N3224, N3217, N2027, N1978, N503);
not NOT1 (N3225, N3204);
not NOT1 (N3226, N3219);
or OR2 (N3227, N3220, N2512);
and AND4 (N3228, N3223, N2903, N778, N623);
buf BUF1 (N3229, N3213);
buf BUF1 (N3230, N3214);
or OR2 (N3231, N3226, N284);
and AND2 (N3232, N3230, N273);
and AND2 (N3233, N3215, N1337);
nand NAND4 (N3234, N3222, N1914, N1100, N2530);
and AND2 (N3235, N3225, N2221);
nor NOR3 (N3236, N3231, N771, N1836);
or OR3 (N3237, N3233, N361, N2298);
nand NAND4 (N3238, N3221, N1507, N271, N2219);
xor XOR2 (N3239, N3227, N960);
or OR3 (N3240, N3236, N2446, N2068);
not NOT1 (N3241, N3232);
nor NOR2 (N3242, N3241, N100);
nand NAND4 (N3243, N3234, N392, N775, N2278);
nor NOR2 (N3244, N3240, N1520);
xor XOR2 (N3245, N3235, N653);
nand NAND4 (N3246, N3239, N384, N2600, N2032);
xor XOR2 (N3247, N3243, N1315);
buf BUF1 (N3248, N3245);
xor XOR2 (N3249, N3247, N1832);
not NOT1 (N3250, N3244);
nand NAND2 (N3251, N3237, N1222);
xor XOR2 (N3252, N3250, N837);
not NOT1 (N3253, N3228);
not NOT1 (N3254, N3242);
xor XOR2 (N3255, N3224, N1722);
nor NOR2 (N3256, N3248, N382);
not NOT1 (N3257, N3256);
not NOT1 (N3258, N3253);
xor XOR2 (N3259, N3254, N653);
not NOT1 (N3260, N3255);
not NOT1 (N3261, N3252);
buf BUF1 (N3262, N3257);
xor XOR2 (N3263, N3238, N2575);
nor NOR4 (N3264, N3259, N2866, N2970, N2081);
not NOT1 (N3265, N3229);
nand NAND2 (N3266, N3249, N1651);
not NOT1 (N3267, N3264);
nand NAND3 (N3268, N3262, N1895, N2463);
not NOT1 (N3269, N3265);
nand NAND3 (N3270, N3251, N3264, N2932);
xor XOR2 (N3271, N3267, N2043);
nor NOR3 (N3272, N3263, N2877, N2216);
or OR3 (N3273, N3266, N3187, N1977);
buf BUF1 (N3274, N3270);
not NOT1 (N3275, N3261);
not NOT1 (N3276, N3246);
nand NAND2 (N3277, N3275, N2911);
or OR4 (N3278, N3272, N969, N894, N2112);
not NOT1 (N3279, N3268);
nand NAND3 (N3280, N3278, N1484, N1184);
and AND2 (N3281, N3279, N1063);
nand NAND3 (N3282, N3258, N2419, N528);
xor XOR2 (N3283, N3274, N2724);
not NOT1 (N3284, N3273);
and AND3 (N3285, N3280, N2486, N990);
nand NAND2 (N3286, N3276, N1095);
and AND3 (N3287, N3260, N452, N20);
not NOT1 (N3288, N3287);
and AND4 (N3289, N3288, N360, N3207, N1064);
not NOT1 (N3290, N3282);
nor NOR2 (N3291, N3290, N2346);
buf BUF1 (N3292, N3281);
not NOT1 (N3293, N3277);
or OR4 (N3294, N3293, N2453, N2726, N2920);
or OR3 (N3295, N3292, N2907, N334);
and AND3 (N3296, N3271, N799, N937);
nand NAND3 (N3297, N3269, N197, N2269);
or OR2 (N3298, N3286, N2664);
not NOT1 (N3299, N3289);
or OR2 (N3300, N3298, N1601);
or OR2 (N3301, N3283, N2500);
nor NOR2 (N3302, N3284, N1419);
xor XOR2 (N3303, N3299, N1984);
nor NOR4 (N3304, N3303, N2966, N2465, N2340);
nand NAND3 (N3305, N3295, N1353, N1876);
not NOT1 (N3306, N3297);
buf BUF1 (N3307, N3300);
and AND3 (N3308, N3302, N2802, N268);
and AND4 (N3309, N3294, N989, N662, N2325);
xor XOR2 (N3310, N3304, N422);
xor XOR2 (N3311, N3296, N1152);
or OR2 (N3312, N3301, N1559);
xor XOR2 (N3313, N3311, N2719);
xor XOR2 (N3314, N3313, N2405);
not NOT1 (N3315, N3312);
or OR3 (N3316, N3305, N3296, N704);
nand NAND4 (N3317, N3309, N3017, N2221, N1034);
or OR3 (N3318, N3291, N2924, N2738);
and AND4 (N3319, N3314, N806, N1858, N709);
nand NAND3 (N3320, N3285, N1191, N845);
not NOT1 (N3321, N3317);
nand NAND2 (N3322, N3316, N2691);
nor NOR3 (N3323, N3315, N1383, N45);
not NOT1 (N3324, N3306);
nand NAND3 (N3325, N3319, N187, N1486);
xor XOR2 (N3326, N3323, N2892);
or OR3 (N3327, N3320, N1604, N889);
not NOT1 (N3328, N3307);
not NOT1 (N3329, N3327);
xor XOR2 (N3330, N3321, N1163);
buf BUF1 (N3331, N3326);
nand NAND2 (N3332, N3325, N1706);
xor XOR2 (N3333, N3310, N1002);
nor NOR2 (N3334, N3331, N2394);
and AND4 (N3335, N3334, N2349, N2550, N356);
and AND2 (N3336, N3318, N2882);
and AND4 (N3337, N3330, N379, N738, N589);
not NOT1 (N3338, N3333);
not NOT1 (N3339, N3324);
nand NAND2 (N3340, N3338, N1684);
not NOT1 (N3341, N3322);
buf BUF1 (N3342, N3341);
nand NAND2 (N3343, N3332, N78);
nor NOR2 (N3344, N3335, N2719);
not NOT1 (N3345, N3308);
and AND4 (N3346, N3340, N2393, N2524, N2075);
buf BUF1 (N3347, N3337);
nor NOR2 (N3348, N3347, N2925);
and AND2 (N3349, N3344, N2871);
buf BUF1 (N3350, N3342);
xor XOR2 (N3351, N3346, N433);
buf BUF1 (N3352, N3349);
or OR3 (N3353, N3339, N2639, N2900);
nor NOR2 (N3354, N3343, N29);
not NOT1 (N3355, N3328);
nor NOR2 (N3356, N3348, N3059);
nor NOR3 (N3357, N3353, N1295, N35);
buf BUF1 (N3358, N3354);
not NOT1 (N3359, N3336);
or OR4 (N3360, N3358, N250, N3315, N1548);
nor NOR3 (N3361, N3345, N3253, N3197);
and AND4 (N3362, N3351, N454, N1621, N3355);
nor NOR2 (N3363, N2666, N1789);
or OR2 (N3364, N3356, N2017);
nor NOR3 (N3365, N3364, N2237, N1570);
or OR4 (N3366, N3361, N2655, N1424, N3100);
or OR4 (N3367, N3362, N2853, N3247, N1512);
nor NOR2 (N3368, N3350, N2728);
nor NOR3 (N3369, N3367, N402, N3075);
and AND4 (N3370, N3329, N2371, N2370, N2329);
nor NOR2 (N3371, N3369, N2572);
or OR3 (N3372, N3366, N2586, N219);
or OR3 (N3373, N3357, N2346, N826);
and AND4 (N3374, N3360, N3170, N1514, N904);
or OR3 (N3375, N3365, N479, N2961);
or OR2 (N3376, N3363, N1116);
xor XOR2 (N3377, N3372, N1263);
or OR3 (N3378, N3376, N1296, N1633);
and AND4 (N3379, N3359, N3056, N1373, N2435);
xor XOR2 (N3380, N3368, N100);
buf BUF1 (N3381, N3374);
xor XOR2 (N3382, N3381, N2606);
not NOT1 (N3383, N3378);
nand NAND2 (N3384, N3382, N621);
nand NAND2 (N3385, N3373, N912);
nor NOR4 (N3386, N3385, N991, N2140, N2724);
or OR2 (N3387, N3384, N876);
buf BUF1 (N3388, N3383);
buf BUF1 (N3389, N3370);
and AND2 (N3390, N3380, N3165);
not NOT1 (N3391, N3387);
nand NAND4 (N3392, N3375, N3284, N1117, N1496);
and AND2 (N3393, N3377, N570);
xor XOR2 (N3394, N3352, N416);
nor NOR3 (N3395, N3379, N1505, N1825);
or OR2 (N3396, N3390, N852);
not NOT1 (N3397, N3392);
nand NAND3 (N3398, N3395, N1222, N2491);
and AND3 (N3399, N3391, N1561, N1216);
not NOT1 (N3400, N3399);
nor NOR2 (N3401, N3394, N421);
or OR3 (N3402, N3400, N1949, N2743);
buf BUF1 (N3403, N3396);
buf BUF1 (N3404, N3402);
xor XOR2 (N3405, N3371, N1238);
or OR2 (N3406, N3398, N808);
nand NAND3 (N3407, N3386, N738, N1842);
xor XOR2 (N3408, N3405, N786);
nor NOR3 (N3409, N3407, N1061, N2122);
not NOT1 (N3410, N3401);
nand NAND3 (N3411, N3389, N1657, N617);
xor XOR2 (N3412, N3404, N3408);
xor XOR2 (N3413, N88, N2374);
buf BUF1 (N3414, N3413);
not NOT1 (N3415, N3410);
buf BUF1 (N3416, N3403);
not NOT1 (N3417, N3412);
nor NOR2 (N3418, N3411, N1276);
xor XOR2 (N3419, N3393, N1986);
or OR2 (N3420, N3414, N861);
nor NOR3 (N3421, N3397, N424, N644);
or OR4 (N3422, N3388, N970, N637, N3419);
nand NAND4 (N3423, N1752, N732, N2412, N84);
xor XOR2 (N3424, N3409, N3297);
or OR2 (N3425, N3415, N94);
nand NAND2 (N3426, N3423, N16);
nand NAND4 (N3427, N3406, N3079, N451, N1978);
xor XOR2 (N3428, N3421, N2237);
xor XOR2 (N3429, N3424, N713);
nand NAND4 (N3430, N3425, N3379, N1153, N1023);
nand NAND2 (N3431, N3426, N2713);
nor NOR3 (N3432, N3416, N2373, N173);
nor NOR3 (N3433, N3422, N59, N512);
not NOT1 (N3434, N3427);
not NOT1 (N3435, N3431);
nor NOR4 (N3436, N3418, N1881, N1845, N2154);
buf BUF1 (N3437, N3430);
xor XOR2 (N3438, N3417, N2729);
or OR4 (N3439, N3428, N523, N2378, N2015);
nand NAND3 (N3440, N3432, N2441, N1316);
nand NAND4 (N3441, N3434, N615, N3017, N1296);
not NOT1 (N3442, N3436);
and AND2 (N3443, N3441, N1315);
nand NAND4 (N3444, N3433, N1608, N757, N2309);
and AND2 (N3445, N3435, N2071);
nor NOR3 (N3446, N3443, N350, N538);
not NOT1 (N3447, N3439);
buf BUF1 (N3448, N3447);
xor XOR2 (N3449, N3445, N1579);
buf BUF1 (N3450, N3446);
and AND2 (N3451, N3450, N1377);
buf BUF1 (N3452, N3437);
buf BUF1 (N3453, N3442);
buf BUF1 (N3454, N3444);
buf BUF1 (N3455, N3448);
not NOT1 (N3456, N3452);
nor NOR4 (N3457, N3453, N2532, N1514, N982);
or OR4 (N3458, N3451, N767, N2100, N3087);
xor XOR2 (N3459, N3449, N1526);
or OR4 (N3460, N3420, N3311, N867, N1470);
buf BUF1 (N3461, N3429);
not NOT1 (N3462, N3460);
nor NOR4 (N3463, N3461, N1338, N2552, N2372);
and AND3 (N3464, N3457, N1442, N3388);
xor XOR2 (N3465, N3462, N320);
xor XOR2 (N3466, N3438, N2994);
not NOT1 (N3467, N3465);
or OR3 (N3468, N3440, N1838, N1380);
nor NOR3 (N3469, N3455, N2682, N518);
xor XOR2 (N3470, N3456, N1748);
nand NAND2 (N3471, N3470, N1171);
nand NAND3 (N3472, N3471, N2510, N1700);
buf BUF1 (N3473, N3459);
or OR2 (N3474, N3472, N1406);
nand NAND3 (N3475, N3474, N2831, N518);
nand NAND3 (N3476, N3463, N1533, N1896);
buf BUF1 (N3477, N3467);
nor NOR2 (N3478, N3466, N1106);
nor NOR3 (N3479, N3473, N1187, N538);
nand NAND2 (N3480, N3454, N992);
and AND3 (N3481, N3469, N55, N1769);
nand NAND3 (N3482, N3477, N1184, N1900);
buf BUF1 (N3483, N3476);
and AND4 (N3484, N3479, N953, N2828, N2009);
xor XOR2 (N3485, N3483, N1763);
buf BUF1 (N3486, N3458);
and AND4 (N3487, N3468, N157, N2384, N406);
xor XOR2 (N3488, N3475, N2231);
buf BUF1 (N3489, N3486);
nor NOR2 (N3490, N3484, N3135);
buf BUF1 (N3491, N3480);
buf BUF1 (N3492, N3464);
not NOT1 (N3493, N3487);
and AND3 (N3494, N3481, N1164, N1362);
or OR3 (N3495, N3482, N848, N823);
nand NAND2 (N3496, N3495, N2376);
nor NOR4 (N3497, N3488, N3331, N713, N638);
buf BUF1 (N3498, N3485);
xor XOR2 (N3499, N3497, N436);
or OR3 (N3500, N3494, N899, N1324);
nand NAND4 (N3501, N3492, N735, N2911, N1621);
xor XOR2 (N3502, N3489, N138);
xor XOR2 (N3503, N3499, N2665);
nand NAND3 (N3504, N3490, N2128, N646);
or OR3 (N3505, N3493, N1611, N1289);
xor XOR2 (N3506, N3500, N555);
or OR3 (N3507, N3478, N2010, N1647);
nand NAND2 (N3508, N3506, N2899);
nor NOR4 (N3509, N3501, N672, N1551, N3499);
or OR4 (N3510, N3498, N849, N2098, N168);
not NOT1 (N3511, N3504);
buf BUF1 (N3512, N3491);
not NOT1 (N3513, N3503);
buf BUF1 (N3514, N3502);
not NOT1 (N3515, N3496);
not NOT1 (N3516, N3515);
or OR3 (N3517, N3508, N541, N3257);
buf BUF1 (N3518, N3512);
nand NAND2 (N3519, N3509, N364);
and AND3 (N3520, N3507, N2513, N2491);
nor NOR2 (N3521, N3510, N628);
and AND3 (N3522, N3519, N496, N1067);
and AND2 (N3523, N3520, N873);
nand NAND4 (N3524, N3518, N538, N1164, N3354);
buf BUF1 (N3525, N3514);
xor XOR2 (N3526, N3522, N3112);
nor NOR3 (N3527, N3513, N825, N2862);
or OR2 (N3528, N3523, N2715);
xor XOR2 (N3529, N3521, N1835);
nand NAND4 (N3530, N3524, N3277, N790, N3286);
and AND2 (N3531, N3516, N555);
or OR4 (N3532, N3526, N2305, N1903, N2910);
not NOT1 (N3533, N3530);
and AND3 (N3534, N3527, N3125, N3065);
or OR2 (N3535, N3533, N2507);
xor XOR2 (N3536, N3511, N3117);
and AND2 (N3537, N3528, N1265);
or OR2 (N3538, N3537, N1360);
buf BUF1 (N3539, N3531);
or OR4 (N3540, N3517, N475, N751, N3139);
buf BUF1 (N3541, N3540);
xor XOR2 (N3542, N3539, N3437);
not NOT1 (N3543, N3525);
xor XOR2 (N3544, N3541, N3060);
nor NOR2 (N3545, N3536, N108);
not NOT1 (N3546, N3542);
buf BUF1 (N3547, N3544);
buf BUF1 (N3548, N3535);
and AND3 (N3549, N3545, N2931, N630);
xor XOR2 (N3550, N3546, N3297);
or OR4 (N3551, N3547, N937, N747, N589);
or OR4 (N3552, N3548, N1840, N3531, N3449);
or OR3 (N3553, N3532, N3410, N412);
nor NOR3 (N3554, N3543, N3325, N31);
or OR2 (N3555, N3553, N1988);
and AND3 (N3556, N3552, N2373, N3411);
xor XOR2 (N3557, N3529, N3184);
xor XOR2 (N3558, N3534, N1897);
and AND2 (N3559, N3554, N2326);
or OR4 (N3560, N3551, N2552, N1121, N1013);
not NOT1 (N3561, N3558);
not NOT1 (N3562, N3559);
nand NAND4 (N3563, N3538, N550, N1912, N2740);
xor XOR2 (N3564, N3556, N1849);
nand NAND2 (N3565, N3555, N3162);
or OR3 (N3566, N3564, N711, N3421);
and AND4 (N3567, N3557, N1355, N1380, N2437);
and AND3 (N3568, N3565, N3441, N320);
xor XOR2 (N3569, N3549, N3502);
or OR3 (N3570, N3561, N911, N3438);
or OR4 (N3571, N3563, N2920, N2601, N1306);
nor NOR2 (N3572, N3571, N2960);
not NOT1 (N3573, N3562);
not NOT1 (N3574, N3566);
nor NOR2 (N3575, N3550, N2475);
or OR4 (N3576, N3575, N2113, N570, N349);
nand NAND2 (N3577, N3573, N2383);
xor XOR2 (N3578, N3567, N1141);
xor XOR2 (N3579, N3568, N476);
and AND2 (N3580, N3572, N1994);
buf BUF1 (N3581, N3580);
buf BUF1 (N3582, N3569);
nand NAND3 (N3583, N3576, N2910, N2064);
or OR2 (N3584, N3582, N2757);
buf BUF1 (N3585, N3583);
nor NOR2 (N3586, N3585, N79);
and AND3 (N3587, N3578, N466, N862);
nor NOR4 (N3588, N3505, N1486, N2707, N2398);
buf BUF1 (N3589, N3586);
nand NAND3 (N3590, N3577, N2512, N1941);
xor XOR2 (N3591, N3587, N128);
nor NOR2 (N3592, N3579, N73);
not NOT1 (N3593, N3590);
nor NOR4 (N3594, N3584, N1246, N2261, N2358);
not NOT1 (N3595, N3594);
or OR2 (N3596, N3574, N2306);
nand NAND4 (N3597, N3595, N2148, N1202, N231);
buf BUF1 (N3598, N3593);
nor NOR4 (N3599, N3598, N1675, N2304, N2305);
nor NOR4 (N3600, N3588, N1848, N2387, N768);
xor XOR2 (N3601, N3589, N2852);
or OR3 (N3602, N3596, N1798, N3057);
nand NAND4 (N3603, N3601, N1060, N259, N488);
or OR4 (N3604, N3597, N3033, N113, N3598);
xor XOR2 (N3605, N3570, N1108);
or OR4 (N3606, N3591, N2463, N3331, N2105);
buf BUF1 (N3607, N3606);
nor NOR4 (N3608, N3605, N1758, N589, N940);
nand NAND4 (N3609, N3560, N2891, N1298, N485);
or OR4 (N3610, N3609, N1144, N94, N2835);
nor NOR4 (N3611, N3610, N1773, N1473, N3055);
buf BUF1 (N3612, N3599);
xor XOR2 (N3613, N3612, N2831);
nand NAND4 (N3614, N3611, N2501, N1617, N2518);
buf BUF1 (N3615, N3592);
and AND3 (N3616, N3602, N146, N1334);
xor XOR2 (N3617, N3607, N1333);
xor XOR2 (N3618, N3608, N2711);
nand NAND4 (N3619, N3617, N1802, N240, N1147);
nor NOR4 (N3620, N3616, N3528, N1464, N2093);
nor NOR2 (N3621, N3603, N2642);
nand NAND2 (N3622, N3613, N2265);
buf BUF1 (N3623, N3618);
xor XOR2 (N3624, N3621, N1936);
nand NAND3 (N3625, N3600, N3588, N2569);
nor NOR2 (N3626, N3622, N1984);
xor XOR2 (N3627, N3623, N3080);
xor XOR2 (N3628, N3626, N2475);
buf BUF1 (N3629, N3624);
and AND4 (N3630, N3615, N364, N2108, N3186);
nor NOR4 (N3631, N3614, N1944, N2809, N3625);
not NOT1 (N3632, N3097);
and AND4 (N3633, N3630, N1612, N1542, N2081);
xor XOR2 (N3634, N3628, N2220);
nand NAND4 (N3635, N3604, N1736, N388, N1413);
and AND3 (N3636, N3581, N1293, N2388);
or OR3 (N3637, N3629, N3583, N1262);
and AND3 (N3638, N3627, N2885, N3314);
nand NAND2 (N3639, N3638, N3049);
buf BUF1 (N3640, N3632);
nor NOR2 (N3641, N3619, N947);
and AND3 (N3642, N3636, N725, N3021);
xor XOR2 (N3643, N3640, N1151);
and AND4 (N3644, N3642, N3485, N1286, N1355);
or OR3 (N3645, N3633, N3574, N1398);
nand NAND2 (N3646, N3639, N1662);
not NOT1 (N3647, N3641);
nand NAND2 (N3648, N3646, N3620);
buf BUF1 (N3649, N1354);
buf BUF1 (N3650, N3635);
nor NOR4 (N3651, N3644, N2447, N54, N73);
and AND2 (N3652, N3649, N490);
nor NOR2 (N3653, N3634, N2409);
nand NAND2 (N3654, N3643, N1112);
and AND3 (N3655, N3648, N2751, N1020);
or OR2 (N3656, N3654, N1884);
xor XOR2 (N3657, N3656, N2368);
nand NAND4 (N3658, N3647, N1708, N2769, N579);
nand NAND4 (N3659, N3653, N1262, N2819, N2190);
nor NOR2 (N3660, N3651, N1182);
or OR4 (N3661, N3658, N924, N1789, N856);
xor XOR2 (N3662, N3631, N3250);
or OR3 (N3663, N3659, N670, N3352);
buf BUF1 (N3664, N3655);
xor XOR2 (N3665, N3661, N2437);
xor XOR2 (N3666, N3657, N3474);
and AND3 (N3667, N3652, N1775, N3049);
nor NOR2 (N3668, N3667, N3535);
nand NAND3 (N3669, N3665, N1773, N1866);
and AND2 (N3670, N3662, N771);
nand NAND4 (N3671, N3666, N3258, N3438, N977);
and AND4 (N3672, N3671, N1473, N2506, N1262);
and AND3 (N3673, N3668, N865, N1681);
not NOT1 (N3674, N3650);
or OR2 (N3675, N3674, N960);
nor NOR3 (N3676, N3670, N922, N1216);
xor XOR2 (N3677, N3669, N1574);
nand NAND4 (N3678, N3645, N2047, N1435, N1944);
buf BUF1 (N3679, N3663);
nand NAND2 (N3680, N3672, N2599);
nor NOR2 (N3681, N3678, N3530);
and AND3 (N3682, N3681, N3300, N2434);
buf BUF1 (N3683, N3664);
or OR2 (N3684, N3673, N715);
and AND2 (N3685, N3677, N502);
xor XOR2 (N3686, N3660, N418);
nand NAND2 (N3687, N3686, N478);
nor NOR3 (N3688, N3680, N794, N1741);
or OR3 (N3689, N3688, N3630, N129);
and AND3 (N3690, N3685, N3063, N1816);
xor XOR2 (N3691, N3690, N368);
nor NOR4 (N3692, N3689, N427, N1856, N3413);
and AND4 (N3693, N3683, N509, N3369, N3546);
or OR3 (N3694, N3675, N36, N3569);
nand NAND3 (N3695, N3637, N149, N1742);
nor NOR3 (N3696, N3687, N2195, N2261);
not NOT1 (N3697, N3691);
or OR2 (N3698, N3679, N192);
xor XOR2 (N3699, N3676, N2540);
buf BUF1 (N3700, N3695);
and AND3 (N3701, N3684, N1849, N1422);
buf BUF1 (N3702, N3693);
xor XOR2 (N3703, N3697, N860);
xor XOR2 (N3704, N3700, N42);
xor XOR2 (N3705, N3692, N342);
nor NOR3 (N3706, N3703, N228, N2346);
or OR2 (N3707, N3701, N2928);
and AND2 (N3708, N3699, N1481);
nor NOR2 (N3709, N3704, N2657);
nor NOR3 (N3710, N3705, N738, N363);
xor XOR2 (N3711, N3694, N3473);
and AND4 (N3712, N3706, N3077, N3580, N1458);
nor NOR2 (N3713, N3710, N3651);
nor NOR4 (N3714, N3713, N3297, N1458, N3378);
nor NOR3 (N3715, N3708, N1099, N2852);
not NOT1 (N3716, N3698);
nor NOR3 (N3717, N3709, N1115, N2623);
nor NOR2 (N3718, N3711, N3706);
xor XOR2 (N3719, N3712, N1904);
and AND4 (N3720, N3716, N463, N523, N1955);
or OR2 (N3721, N3715, N3196);
buf BUF1 (N3722, N3717);
and AND4 (N3723, N3721, N231, N3393, N3549);
nor NOR2 (N3724, N3714, N3619);
nor NOR4 (N3725, N3724, N629, N2328, N2701);
or OR2 (N3726, N3725, N1013);
nor NOR2 (N3727, N3719, N802);
nor NOR3 (N3728, N3722, N340, N3661);
and AND3 (N3729, N3702, N923, N87);
and AND2 (N3730, N3728, N396);
xor XOR2 (N3731, N3696, N3469);
nand NAND3 (N3732, N3727, N188, N2399);
not NOT1 (N3733, N3723);
buf BUF1 (N3734, N3732);
nor NOR2 (N3735, N3726, N3254);
xor XOR2 (N3736, N3682, N1643);
xor XOR2 (N3737, N3735, N3616);
xor XOR2 (N3738, N3720, N2763);
not NOT1 (N3739, N3730);
nor NOR2 (N3740, N3729, N3384);
nand NAND4 (N3741, N3734, N839, N2056, N3269);
and AND3 (N3742, N3740, N3419, N2713);
nand NAND2 (N3743, N3737, N2366);
nor NOR3 (N3744, N3736, N2670, N3096);
or OR4 (N3745, N3718, N523, N2860, N2445);
nand NAND2 (N3746, N3741, N2452);
nand NAND2 (N3747, N3733, N2267);
nor NOR2 (N3748, N3739, N3662);
buf BUF1 (N3749, N3747);
and AND3 (N3750, N3749, N2196, N1733);
or OR2 (N3751, N3744, N3342);
and AND3 (N3752, N3748, N3317, N273);
nor NOR2 (N3753, N3752, N3694);
or OR2 (N3754, N3707, N1348);
and AND3 (N3755, N3750, N236, N1329);
and AND2 (N3756, N3743, N1402);
xor XOR2 (N3757, N3731, N609);
or OR4 (N3758, N3753, N2354, N3688, N260);
or OR3 (N3759, N3746, N2015, N2512);
and AND3 (N3760, N3738, N515, N1583);
xor XOR2 (N3761, N3754, N2111);
and AND4 (N3762, N3757, N2344, N3549, N3726);
nor NOR3 (N3763, N3755, N2047, N1842);
nand NAND2 (N3764, N3742, N866);
nand NAND3 (N3765, N3751, N1031, N8);
nor NOR3 (N3766, N3764, N821, N192);
buf BUF1 (N3767, N3766);
and AND2 (N3768, N3745, N2714);
nand NAND3 (N3769, N3759, N2441, N190);
buf BUF1 (N3770, N3758);
or OR4 (N3771, N3760, N3357, N1206, N768);
not NOT1 (N3772, N3771);
xor XOR2 (N3773, N3765, N1977);
nand NAND4 (N3774, N3767, N2167, N665, N2624);
or OR3 (N3775, N3772, N409, N2408);
xor XOR2 (N3776, N3762, N3526);
not NOT1 (N3777, N3775);
not NOT1 (N3778, N3777);
nand NAND4 (N3779, N3770, N2669, N383, N556);
buf BUF1 (N3780, N3774);
nor NOR2 (N3781, N3773, N21);
or OR2 (N3782, N3778, N896);
xor XOR2 (N3783, N3769, N3227);
or OR3 (N3784, N3761, N2647, N3174);
not NOT1 (N3785, N3779);
buf BUF1 (N3786, N3780);
buf BUF1 (N3787, N3782);
buf BUF1 (N3788, N3768);
or OR3 (N3789, N3776, N1556, N3296);
nand NAND4 (N3790, N3788, N1517, N2230, N1035);
or OR3 (N3791, N3756, N1784, N216);
nor NOR2 (N3792, N3783, N2370);
and AND4 (N3793, N3790, N2737, N3410, N3407);
nand NAND2 (N3794, N3789, N1625);
nand NAND2 (N3795, N3786, N2353);
nor NOR3 (N3796, N3784, N1123, N1932);
or OR4 (N3797, N3785, N2367, N2204, N30);
not NOT1 (N3798, N3787);
xor XOR2 (N3799, N3793, N2118);
and AND3 (N3800, N3781, N539, N2899);
nand NAND3 (N3801, N3798, N2148, N1585);
xor XOR2 (N3802, N3795, N1358);
and AND2 (N3803, N3801, N3380);
xor XOR2 (N3804, N3802, N440);
buf BUF1 (N3805, N3792);
buf BUF1 (N3806, N3794);
not NOT1 (N3807, N3791);
not NOT1 (N3808, N3797);
nor NOR4 (N3809, N3805, N152, N3100, N1414);
nand NAND3 (N3810, N3807, N2672, N2191);
and AND4 (N3811, N3803, N3585, N2379, N3493);
buf BUF1 (N3812, N3808);
not NOT1 (N3813, N3810);
and AND2 (N3814, N3811, N2793);
or OR2 (N3815, N3809, N3636);
xor XOR2 (N3816, N3814, N532);
or OR2 (N3817, N3796, N431);
buf BUF1 (N3818, N3813);
or OR4 (N3819, N3815, N2849, N2881, N1902);
and AND3 (N3820, N3799, N397, N1585);
nor NOR4 (N3821, N3819, N2738, N2330, N3346);
xor XOR2 (N3822, N3820, N1421);
nor NOR3 (N3823, N3812, N1788, N172);
buf BUF1 (N3824, N3816);
nand NAND3 (N3825, N3824, N1330, N3331);
or OR4 (N3826, N3825, N3212, N1048, N739);
and AND4 (N3827, N3822, N2479, N2195, N1883);
and AND2 (N3828, N3826, N3215);
nor NOR3 (N3829, N3823, N1076, N53);
and AND4 (N3830, N3804, N354, N3020, N1166);
xor XOR2 (N3831, N3817, N1992);
not NOT1 (N3832, N3831);
or OR2 (N3833, N3830, N539);
not NOT1 (N3834, N3833);
buf BUF1 (N3835, N3832);
buf BUF1 (N3836, N3821);
nand NAND3 (N3837, N3834, N1045, N3657);
xor XOR2 (N3838, N3828, N1853);
and AND2 (N3839, N3827, N3531);
or OR2 (N3840, N3837, N3547);
or OR2 (N3841, N3818, N302);
xor XOR2 (N3842, N3835, N2247);
or OR4 (N3843, N3806, N2148, N2685, N2741);
buf BUF1 (N3844, N3800);
and AND4 (N3845, N3840, N2820, N3248, N317);
not NOT1 (N3846, N3841);
xor XOR2 (N3847, N3842, N3099);
nand NAND2 (N3848, N3763, N1976);
not NOT1 (N3849, N3848);
or OR4 (N3850, N3844, N326, N3033, N3666);
not NOT1 (N3851, N3849);
nor NOR4 (N3852, N3838, N495, N2016, N345);
or OR4 (N3853, N3847, N731, N121, N1310);
buf BUF1 (N3854, N3846);
or OR3 (N3855, N3845, N1361, N3393);
and AND2 (N3856, N3851, N350);
or OR4 (N3857, N3850, N1286, N2318, N880);
and AND2 (N3858, N3854, N1561);
nand NAND4 (N3859, N3836, N3447, N2438, N1772);
xor XOR2 (N3860, N3856, N3377);
xor XOR2 (N3861, N3843, N998);
nand NAND4 (N3862, N3860, N1625, N1997, N1520);
nand NAND4 (N3863, N3861, N376, N1493, N1386);
or OR2 (N3864, N3862, N1937);
buf BUF1 (N3865, N3857);
not NOT1 (N3866, N3863);
not NOT1 (N3867, N3865);
buf BUF1 (N3868, N3829);
or OR3 (N3869, N3864, N363, N1141);
or OR3 (N3870, N3855, N1165, N2201);
nor NOR3 (N3871, N3870, N958, N2128);
or OR3 (N3872, N3853, N2490, N2766);
xor XOR2 (N3873, N3858, N2166);
nor NOR4 (N3874, N3866, N1474, N3527, N3496);
xor XOR2 (N3875, N3867, N757);
and AND2 (N3876, N3852, N1684);
nor NOR3 (N3877, N3839, N5, N2053);
or OR3 (N3878, N3876, N3080, N3437);
nor NOR3 (N3879, N3871, N1562, N2549);
xor XOR2 (N3880, N3877, N2930);
xor XOR2 (N3881, N3880, N418);
not NOT1 (N3882, N3872);
nand NAND2 (N3883, N3878, N2612);
xor XOR2 (N3884, N3875, N3259);
or OR3 (N3885, N3883, N709, N2724);
nor NOR4 (N3886, N3882, N1828, N3850, N1952);
nor NOR4 (N3887, N3881, N363, N559, N1750);
and AND4 (N3888, N3879, N3027, N3858, N2540);
nand NAND4 (N3889, N3859, N3503, N2126, N3706);
nor NOR4 (N3890, N3889, N1937, N1351, N935);
and AND4 (N3891, N3885, N2425, N3067, N36);
buf BUF1 (N3892, N3884);
or OR2 (N3893, N3892, N2336);
xor XOR2 (N3894, N3887, N1617);
xor XOR2 (N3895, N3890, N2845);
and AND4 (N3896, N3893, N3660, N2143, N3021);
or OR3 (N3897, N3868, N72, N1012);
and AND3 (N3898, N3895, N3226, N3267);
nand NAND4 (N3899, N3896, N1795, N2968, N1053);
and AND4 (N3900, N3899, N1651, N315, N940);
buf BUF1 (N3901, N3888);
not NOT1 (N3902, N3897);
and AND2 (N3903, N3900, N1018);
nor NOR2 (N3904, N3886, N490);
xor XOR2 (N3905, N3894, N3191);
or OR4 (N3906, N3904, N2555, N2825, N436);
not NOT1 (N3907, N3902);
nand NAND2 (N3908, N3901, N3123);
nor NOR2 (N3909, N3907, N2133);
not NOT1 (N3910, N3874);
and AND3 (N3911, N3891, N3382, N496);
nor NOR4 (N3912, N3898, N1827, N2547, N513);
xor XOR2 (N3913, N3905, N3152);
and AND2 (N3914, N3903, N826);
nor NOR2 (N3915, N3914, N86);
xor XOR2 (N3916, N3915, N1013);
buf BUF1 (N3917, N3906);
or OR2 (N3918, N3869, N3734);
nor NOR2 (N3919, N3911, N280);
and AND4 (N3920, N3913, N3757, N3272, N2873);
nor NOR3 (N3921, N3919, N484, N282);
not NOT1 (N3922, N3873);
xor XOR2 (N3923, N3920, N3569);
not NOT1 (N3924, N3909);
or OR3 (N3925, N3910, N2925, N1538);
nand NAND4 (N3926, N3924, N2540, N3294, N25);
nor NOR4 (N3927, N3908, N635, N1490, N850);
and AND3 (N3928, N3926, N1153, N546);
not NOT1 (N3929, N3917);
and AND2 (N3930, N3912, N2377);
or OR4 (N3931, N3927, N2743, N3507, N1961);
nand NAND3 (N3932, N3929, N2800, N3765);
nand NAND2 (N3933, N3928, N3586);
not NOT1 (N3934, N3921);
nor NOR2 (N3935, N3930, N806);
nor NOR4 (N3936, N3918, N670, N1176, N2436);
and AND2 (N3937, N3933, N478);
buf BUF1 (N3938, N3922);
xor XOR2 (N3939, N3936, N3468);
buf BUF1 (N3940, N3916);
nand NAND4 (N3941, N3923, N2235, N931, N2128);
and AND2 (N3942, N3937, N213);
xor XOR2 (N3943, N3940, N136);
nand NAND4 (N3944, N3939, N3251, N3868, N1326);
nand NAND2 (N3945, N3934, N2925);
or OR4 (N3946, N3942, N2520, N622, N827);
not NOT1 (N3947, N3943);
and AND4 (N3948, N3938, N2413, N930, N1420);
or OR3 (N3949, N3941, N776, N3581);
nor NOR4 (N3950, N3945, N1995, N1460, N2326);
not NOT1 (N3951, N3947);
not NOT1 (N3952, N3948);
or OR3 (N3953, N3949, N350, N3388);
or OR3 (N3954, N3953, N3690, N3949);
nand NAND2 (N3955, N3950, N911);
or OR3 (N3956, N3931, N3846, N918);
buf BUF1 (N3957, N3955);
buf BUF1 (N3958, N3944);
nor NOR3 (N3959, N3925, N2371, N261);
and AND2 (N3960, N3932, N589);
buf BUF1 (N3961, N3952);
or OR4 (N3962, N3960, N3883, N3031, N267);
not NOT1 (N3963, N3958);
or OR2 (N3964, N3946, N3760);
or OR2 (N3965, N3959, N457);
nor NOR3 (N3966, N3962, N1102, N1498);
and AND4 (N3967, N3935, N2508, N942, N228);
nor NOR2 (N3968, N3954, N200);
nor NOR3 (N3969, N3963, N3027, N2850);
not NOT1 (N3970, N3966);
nor NOR3 (N3971, N3965, N2295, N551);
xor XOR2 (N3972, N3957, N3779);
and AND4 (N3973, N3971, N1675, N249, N1861);
and AND3 (N3974, N3951, N3567, N2941);
or OR4 (N3975, N3974, N1839, N1745, N68);
not NOT1 (N3976, N3973);
or OR3 (N3977, N3969, N2421, N287);
or OR3 (N3978, N3956, N2708, N238);
xor XOR2 (N3979, N3975, N2580);
buf BUF1 (N3980, N3977);
buf BUF1 (N3981, N3976);
and AND3 (N3982, N3961, N3582, N2311);
xor XOR2 (N3983, N3967, N2273);
and AND2 (N3984, N3978, N3150);
and AND3 (N3985, N3980, N2864, N325);
nor NOR2 (N3986, N3981, N3355);
nor NOR2 (N3987, N3964, N1582);
and AND4 (N3988, N3970, N194, N562, N2257);
nor NOR2 (N3989, N3983, N3436);
or OR3 (N3990, N3979, N2677, N1541);
and AND2 (N3991, N3990, N1814);
or OR4 (N3992, N3991, N1588, N1655, N755);
or OR3 (N3993, N3987, N2370, N2001);
not NOT1 (N3994, N3988);
xor XOR2 (N3995, N3992, N332);
buf BUF1 (N3996, N3993);
and AND2 (N3997, N3989, N633);
xor XOR2 (N3998, N3994, N567);
not NOT1 (N3999, N3998);
not NOT1 (N4000, N3984);
xor XOR2 (N4001, N3982, N394);
xor XOR2 (N4002, N3996, N1119);
or OR4 (N4003, N4000, N386, N510, N2599);
xor XOR2 (N4004, N3986, N3260);
or OR4 (N4005, N3985, N2855, N3159, N1568);
nand NAND2 (N4006, N4004, N3775);
nor NOR4 (N4007, N3968, N1865, N372, N1450);
and AND3 (N4008, N4007, N651, N3548);
nand NAND2 (N4009, N4006, N3571);
and AND4 (N4010, N3972, N2742, N151, N2264);
nor NOR4 (N4011, N4001, N884, N1757, N376);
buf BUF1 (N4012, N4002);
nor NOR2 (N4013, N3997, N516);
and AND2 (N4014, N4003, N726);
nand NAND2 (N4015, N4014, N1770);
or OR2 (N4016, N3995, N2006);
buf BUF1 (N4017, N4009);
xor XOR2 (N4018, N4013, N2136);
nand NAND4 (N4019, N4005, N1749, N3329, N33);
or OR4 (N4020, N4008, N966, N3657, N2531);
nor NOR4 (N4021, N3999, N2589, N2755, N512);
nor NOR4 (N4022, N4011, N1867, N1142, N1284);
nor NOR2 (N4023, N4010, N2827);
and AND2 (N4024, N4023, N2989);
or OR2 (N4025, N4020, N1551);
nand NAND4 (N4026, N4012, N704, N1669, N1982);
buf BUF1 (N4027, N4024);
or OR4 (N4028, N4017, N3937, N827, N2170);
xor XOR2 (N4029, N4018, N2636);
not NOT1 (N4030, N4016);
and AND4 (N4031, N4019, N3735, N2943, N1912);
not NOT1 (N4032, N4022);
buf BUF1 (N4033, N4027);
nand NAND3 (N4034, N4031, N723, N3440);
nand NAND3 (N4035, N4021, N1354, N1382);
nor NOR2 (N4036, N4033, N734);
nor NOR2 (N4037, N4025, N2068);
nand NAND2 (N4038, N4032, N727);
xor XOR2 (N4039, N4037, N89);
not NOT1 (N4040, N4029);
nor NOR2 (N4041, N4028, N3148);
buf BUF1 (N4042, N4026);
buf BUF1 (N4043, N4042);
nor NOR3 (N4044, N4043, N2232, N1095);
not NOT1 (N4045, N4038);
and AND4 (N4046, N4035, N1715, N625, N990);
xor XOR2 (N4047, N4039, N2119);
buf BUF1 (N4048, N4041);
nand NAND4 (N4049, N4040, N230, N986, N19);
and AND4 (N4050, N4049, N3463, N3275, N1458);
nor NOR3 (N4051, N4045, N3530, N3842);
nand NAND4 (N4052, N4044, N2670, N998, N1894);
xor XOR2 (N4053, N4051, N3294);
xor XOR2 (N4054, N4034, N1184);
buf BUF1 (N4055, N4046);
buf BUF1 (N4056, N4030);
nor NOR3 (N4057, N4055, N1962, N591);
and AND4 (N4058, N4050, N3704, N652, N2906);
nand NAND3 (N4059, N4036, N505, N563);
xor XOR2 (N4060, N4047, N952);
and AND2 (N4061, N4060, N265);
xor XOR2 (N4062, N4052, N14);
and AND2 (N4063, N4054, N3211);
nor NOR2 (N4064, N4061, N41);
nor NOR4 (N4065, N4058, N3621, N2023, N2325);
buf BUF1 (N4066, N4048);
nor NOR3 (N4067, N4059, N1313, N1679);
xor XOR2 (N4068, N4066, N2130);
or OR3 (N4069, N4062, N2150, N3159);
and AND4 (N4070, N4064, N153, N3460, N27);
or OR3 (N4071, N4056, N1653, N1027);
not NOT1 (N4072, N4063);
not NOT1 (N4073, N4069);
nor NOR2 (N4074, N4068, N2068);
or OR3 (N4075, N4074, N3135, N3248);
buf BUF1 (N4076, N4071);
nand NAND3 (N4077, N4065, N1629, N1841);
not NOT1 (N4078, N4015);
and AND2 (N4079, N4075, N1603);
and AND2 (N4080, N4076, N1008);
nor NOR3 (N4081, N4053, N1286, N97);
and AND2 (N4082, N4070, N3420);
buf BUF1 (N4083, N4078);
nor NOR4 (N4084, N4081, N1780, N1396, N3685);
nor NOR3 (N4085, N4079, N1789, N1946);
xor XOR2 (N4086, N4082, N1885);
nand NAND2 (N4087, N4083, N184);
buf BUF1 (N4088, N4080);
and AND4 (N4089, N4086, N864, N883, N76);
nand NAND4 (N4090, N4089, N2024, N3271, N504);
xor XOR2 (N4091, N4090, N2910);
buf BUF1 (N4092, N4088);
or OR3 (N4093, N4091, N2470, N177);
nand NAND3 (N4094, N4085, N2939, N730);
or OR2 (N4095, N4073, N1146);
nand NAND4 (N4096, N4095, N3307, N2032, N1602);
nand NAND2 (N4097, N4057, N3636);
and AND2 (N4098, N4097, N1028);
and AND2 (N4099, N4093, N2307);
xor XOR2 (N4100, N4094, N3300);
buf BUF1 (N4101, N4077);
nor NOR2 (N4102, N4092, N1285);
and AND3 (N4103, N4102, N2928, N2968);
buf BUF1 (N4104, N4087);
nand NAND4 (N4105, N4104, N3910, N1627, N2513);
nor NOR4 (N4106, N4103, N1652, N2222, N1572);
not NOT1 (N4107, N4106);
xor XOR2 (N4108, N4100, N1021);
xor XOR2 (N4109, N4096, N3383);
or OR4 (N4110, N4101, N2340, N866, N1183);
nor NOR2 (N4111, N4084, N3742);
xor XOR2 (N4112, N4110, N1652);
and AND4 (N4113, N4072, N3470, N3227, N3664);
nor NOR4 (N4114, N4098, N3047, N766, N3684);
nand NAND3 (N4115, N4107, N2296, N401);
nand NAND4 (N4116, N4067, N2540, N961, N1400);
not NOT1 (N4117, N4113);
or OR4 (N4118, N4116, N2056, N2221, N2862);
nand NAND2 (N4119, N4108, N2638);
xor XOR2 (N4120, N4105, N2678);
nor NOR3 (N4121, N4115, N2482, N2615);
nand NAND3 (N4122, N4117, N2214, N2164);
and AND3 (N4123, N4114, N1245, N3422);
buf BUF1 (N4124, N4123);
or OR4 (N4125, N4121, N2230, N1590, N2757);
nand NAND4 (N4126, N4119, N379, N1825, N2235);
buf BUF1 (N4127, N4126);
xor XOR2 (N4128, N4109, N1276);
nor NOR4 (N4129, N4125, N338, N3807, N3608);
xor XOR2 (N4130, N4118, N1104);
or OR3 (N4131, N4099, N1849, N654);
buf BUF1 (N4132, N4124);
and AND4 (N4133, N4120, N324, N1831, N398);
or OR4 (N4134, N4112, N767, N2416, N3147);
xor XOR2 (N4135, N4128, N2091);
xor XOR2 (N4136, N4134, N3994);
buf BUF1 (N4137, N4133);
or OR2 (N4138, N4111, N3105);
nor NOR3 (N4139, N4131, N3461, N693);
buf BUF1 (N4140, N4138);
nor NOR3 (N4141, N4136, N910, N881);
not NOT1 (N4142, N4141);
buf BUF1 (N4143, N4142);
not NOT1 (N4144, N4127);
nor NOR2 (N4145, N4122, N2971);
nor NOR2 (N4146, N4132, N1870);
nor NOR3 (N4147, N4145, N195, N219);
nand NAND2 (N4148, N4137, N1072);
nor NOR3 (N4149, N4148, N1759, N3316);
buf BUF1 (N4150, N4130);
and AND4 (N4151, N4143, N1398, N3552, N2180);
or OR3 (N4152, N4129, N513, N3885);
nand NAND4 (N4153, N4147, N3845, N648, N3711);
nor NOR2 (N4154, N4146, N3899);
not NOT1 (N4155, N4153);
nand NAND2 (N4156, N4140, N3219);
not NOT1 (N4157, N4150);
buf BUF1 (N4158, N4135);
buf BUF1 (N4159, N4156);
and AND2 (N4160, N4158, N3223);
and AND4 (N4161, N4154, N2231, N1408, N923);
nand NAND3 (N4162, N4157, N1179, N3566);
nor NOR3 (N4163, N4155, N2377, N771);
nand NAND3 (N4164, N4161, N3600, N1910);
nand NAND3 (N4165, N4163, N610, N2818);
not NOT1 (N4166, N4151);
buf BUF1 (N4167, N4164);
nor NOR3 (N4168, N4149, N674, N1981);
nor NOR2 (N4169, N4160, N1384);
xor XOR2 (N4170, N4167, N1701);
or OR2 (N4171, N4152, N1985);
not NOT1 (N4172, N4169);
or OR2 (N4173, N4159, N1831);
nor NOR2 (N4174, N4144, N1972);
not NOT1 (N4175, N4173);
or OR3 (N4176, N4170, N1988, N2799);
not NOT1 (N4177, N4176);
nor NOR4 (N4178, N4165, N1146, N733, N1140);
or OR2 (N4179, N4168, N1671);
nor NOR3 (N4180, N4175, N459, N1694);
buf BUF1 (N4181, N4166);
not NOT1 (N4182, N4177);
or OR2 (N4183, N4174, N135);
or OR4 (N4184, N4182, N3987, N3337, N4175);
xor XOR2 (N4185, N4181, N2828);
xor XOR2 (N4186, N4172, N632);
xor XOR2 (N4187, N4186, N1602);
or OR4 (N4188, N4171, N1311, N467, N3074);
not NOT1 (N4189, N4185);
or OR4 (N4190, N4188, N3057, N1964, N697);
nand NAND4 (N4191, N4189, N3229, N3222, N3690);
nor NOR2 (N4192, N4139, N2177);
nand NAND2 (N4193, N4187, N1477);
buf BUF1 (N4194, N4179);
and AND2 (N4195, N4193, N116);
nand NAND4 (N4196, N4162, N2925, N3584, N2765);
buf BUF1 (N4197, N4183);
and AND4 (N4198, N4178, N36, N3794, N403);
nand NAND2 (N4199, N4198, N3644);
nand NAND3 (N4200, N4195, N3399, N2301);
xor XOR2 (N4201, N4194, N4102);
xor XOR2 (N4202, N4200, N423);
xor XOR2 (N4203, N4192, N3796);
xor XOR2 (N4204, N4184, N398);
or OR2 (N4205, N4196, N2183);
nand NAND3 (N4206, N4205, N1833, N960);
not NOT1 (N4207, N4201);
and AND3 (N4208, N4204, N586, N741);
nor NOR3 (N4209, N4190, N325, N1207);
xor XOR2 (N4210, N4191, N162);
not NOT1 (N4211, N4209);
and AND3 (N4212, N4211, N2625, N1143);
nor NOR4 (N4213, N4212, N3662, N329, N1520);
not NOT1 (N4214, N4199);
nor NOR3 (N4215, N4214, N1857, N799);
nand NAND4 (N4216, N4215, N2056, N1641, N2114);
nand NAND4 (N4217, N4210, N3574, N1216, N490);
nor NOR4 (N4218, N4213, N2909, N3116, N707);
or OR2 (N4219, N4197, N2588);
nand NAND3 (N4220, N4218, N3751, N3387);
buf BUF1 (N4221, N4180);
xor XOR2 (N4222, N4203, N3590);
not NOT1 (N4223, N4222);
xor XOR2 (N4224, N4216, N1961);
nand NAND2 (N4225, N4217, N1086);
not NOT1 (N4226, N4207);
xor XOR2 (N4227, N4202, N4099);
and AND3 (N4228, N4225, N3308, N359);
nand NAND2 (N4229, N4220, N2787);
xor XOR2 (N4230, N4228, N1920);
nor NOR3 (N4231, N4223, N1180, N1990);
nor NOR4 (N4232, N4208, N3677, N2153, N2597);
nor NOR2 (N4233, N4227, N1060);
or OR3 (N4234, N4221, N2260, N2589);
nor NOR2 (N4235, N4224, N3648);
nor NOR4 (N4236, N4233, N1878, N3823, N451);
nand NAND3 (N4237, N4236, N2291, N3620);
buf BUF1 (N4238, N4226);
nand NAND4 (N4239, N4229, N2368, N2601, N2030);
buf BUF1 (N4240, N4230);
xor XOR2 (N4241, N4239, N3756);
nand NAND3 (N4242, N4240, N3511, N3063);
or OR3 (N4243, N4241, N2398, N2153);
xor XOR2 (N4244, N4242, N2797);
nor NOR3 (N4245, N4234, N3616, N2999);
buf BUF1 (N4246, N4238);
nor NOR2 (N4247, N4237, N4097);
nor NOR2 (N4248, N4245, N75);
nor NOR3 (N4249, N4232, N2952, N2834);
and AND3 (N4250, N4219, N1198, N548);
or OR4 (N4251, N4248, N870, N2707, N4016);
not NOT1 (N4252, N4250);
or OR4 (N4253, N4231, N2182, N3921, N1928);
or OR2 (N4254, N4244, N1963);
nor NOR2 (N4255, N4235, N2706);
xor XOR2 (N4256, N4247, N213);
xor XOR2 (N4257, N4256, N4135);
nand NAND3 (N4258, N4206, N1466, N2199);
buf BUF1 (N4259, N4257);
not NOT1 (N4260, N4253);
or OR3 (N4261, N4258, N855, N2334);
and AND4 (N4262, N4260, N2039, N2588, N4077);
buf BUF1 (N4263, N4262);
nand NAND3 (N4264, N4255, N4248, N1046);
xor XOR2 (N4265, N4251, N1687);
nor NOR3 (N4266, N4265, N3791, N3429);
buf BUF1 (N4267, N4263);
not NOT1 (N4268, N4259);
nor NOR3 (N4269, N4266, N1177, N1071);
buf BUF1 (N4270, N4269);
or OR2 (N4271, N4270, N3762);
not NOT1 (N4272, N4267);
nor NOR3 (N4273, N4271, N1847, N2491);
buf BUF1 (N4274, N4261);
nand NAND2 (N4275, N4273, N2214);
or OR2 (N4276, N4274, N2731);
xor XOR2 (N4277, N4254, N1609);
nor NOR4 (N4278, N4276, N1054, N2473, N2088);
xor XOR2 (N4279, N4268, N2119);
nand NAND4 (N4280, N4272, N2089, N4246, N887);
nand NAND2 (N4281, N4016, N1147);
buf BUF1 (N4282, N4279);
and AND4 (N4283, N4249, N410, N3994, N2485);
nor NOR2 (N4284, N4252, N3678);
and AND3 (N4285, N4281, N1394, N2743);
and AND2 (N4286, N4275, N353);
or OR3 (N4287, N4286, N1321, N2147);
or OR4 (N4288, N4283, N2128, N345, N411);
or OR2 (N4289, N4285, N2755);
xor XOR2 (N4290, N4243, N2102);
buf BUF1 (N4291, N4288);
and AND2 (N4292, N4287, N226);
buf BUF1 (N4293, N4290);
nand NAND2 (N4294, N4284, N3435);
not NOT1 (N4295, N4264);
nor NOR2 (N4296, N4289, N2124);
and AND3 (N4297, N4292, N3154, N1745);
xor XOR2 (N4298, N4280, N4056);
nor NOR2 (N4299, N4298, N1408);
not NOT1 (N4300, N4294);
not NOT1 (N4301, N4282);
xor XOR2 (N4302, N4301, N1630);
or OR3 (N4303, N4277, N113, N2493);
buf BUF1 (N4304, N4302);
buf BUF1 (N4305, N4304);
xor XOR2 (N4306, N4303, N3692);
or OR3 (N4307, N4306, N2672, N503);
nor NOR3 (N4308, N4291, N1934, N4240);
xor XOR2 (N4309, N4308, N1158);
buf BUF1 (N4310, N4305);
not NOT1 (N4311, N4295);
not NOT1 (N4312, N4310);
nand NAND2 (N4313, N4299, N1681);
xor XOR2 (N4314, N4293, N1747);
or OR3 (N4315, N4307, N2994, N1695);
and AND2 (N4316, N4296, N2778);
and AND3 (N4317, N4309, N1886, N185);
buf BUF1 (N4318, N4278);
or OR3 (N4319, N4318, N4097, N1896);
not NOT1 (N4320, N4315);
not NOT1 (N4321, N4320);
xor XOR2 (N4322, N4300, N616);
xor XOR2 (N4323, N4314, N3391);
nor NOR3 (N4324, N4317, N2614, N3562);
buf BUF1 (N4325, N4321);
not NOT1 (N4326, N4322);
nor NOR2 (N4327, N4323, N2487);
and AND3 (N4328, N4312, N473, N299);
and AND2 (N4329, N4325, N2797);
nor NOR3 (N4330, N4327, N4313, N2339);
not NOT1 (N4331, N4042);
nand NAND4 (N4332, N4328, N2087, N1145, N892);
buf BUF1 (N4333, N4332);
not NOT1 (N4334, N4316);
buf BUF1 (N4335, N4330);
buf BUF1 (N4336, N4319);
xor XOR2 (N4337, N4326, N2080);
buf BUF1 (N4338, N4333);
or OR2 (N4339, N4329, N881);
nor NOR3 (N4340, N4337, N1313, N960);
not NOT1 (N4341, N4331);
or OR2 (N4342, N4324, N3313);
buf BUF1 (N4343, N4334);
and AND2 (N4344, N4311, N3362);
or OR3 (N4345, N4340, N679, N1206);
not NOT1 (N4346, N4344);
and AND2 (N4347, N4336, N4255);
xor XOR2 (N4348, N4347, N2078);
nor NOR4 (N4349, N4341, N1918, N1574, N1342);
nor NOR4 (N4350, N4348, N196, N333, N1369);
xor XOR2 (N4351, N4335, N3823);
xor XOR2 (N4352, N4339, N3987);
or OR4 (N4353, N4351, N2050, N1031, N59);
or OR3 (N4354, N4349, N3304, N739);
nor NOR3 (N4355, N4297, N431, N3341);
xor XOR2 (N4356, N4346, N3177);
nand NAND2 (N4357, N4338, N1227);
xor XOR2 (N4358, N4352, N3190);
nand NAND2 (N4359, N4354, N1012);
buf BUF1 (N4360, N4358);
nor NOR4 (N4361, N4343, N3069, N4129, N741);
buf BUF1 (N4362, N4350);
buf BUF1 (N4363, N4360);
xor XOR2 (N4364, N4355, N2767);
not NOT1 (N4365, N4345);
or OR3 (N4366, N4353, N2861, N3370);
not NOT1 (N4367, N4366);
or OR3 (N4368, N4361, N2006, N2354);
nand NAND2 (N4369, N4367, N1903);
nor NOR2 (N4370, N4356, N2602);
nand NAND4 (N4371, N4342, N587, N559, N3150);
not NOT1 (N4372, N4363);
buf BUF1 (N4373, N4357);
not NOT1 (N4374, N4362);
xor XOR2 (N4375, N4368, N1712);
nand NAND2 (N4376, N4370, N2821);
not NOT1 (N4377, N4364);
xor XOR2 (N4378, N4369, N2451);
nor NOR3 (N4379, N4375, N3357, N3225);
nand NAND4 (N4380, N4365, N3985, N1421, N1312);
buf BUF1 (N4381, N4377);
nand NAND3 (N4382, N4371, N2131, N622);
nor NOR4 (N4383, N4374, N768, N3980, N963);
or OR2 (N4384, N4372, N537);
nor NOR2 (N4385, N4373, N2176);
nand NAND4 (N4386, N4379, N1872, N3097, N2515);
and AND2 (N4387, N4386, N1691);
and AND4 (N4388, N4383, N3845, N2570, N1497);
nor NOR4 (N4389, N4382, N2434, N716, N1159);
or OR4 (N4390, N4389, N365, N1590, N825);
not NOT1 (N4391, N4390);
or OR4 (N4392, N4381, N862, N2939, N2501);
nand NAND2 (N4393, N4391, N1623);
nand NAND2 (N4394, N4392, N1336);
nand NAND2 (N4395, N4394, N1396);
and AND2 (N4396, N4385, N697);
buf BUF1 (N4397, N4393);
buf BUF1 (N4398, N4378);
xor XOR2 (N4399, N4398, N2072);
not NOT1 (N4400, N4380);
nand NAND3 (N4401, N4387, N2929, N334);
nor NOR2 (N4402, N4396, N3441);
nand NAND4 (N4403, N4384, N1593, N2588, N1072);
xor XOR2 (N4404, N4388, N445);
and AND4 (N4405, N4376, N1150, N3239, N3218);
nand NAND3 (N4406, N4401, N3170, N2924);
nand NAND3 (N4407, N4359, N940, N4228);
nand NAND2 (N4408, N4402, N762);
nor NOR4 (N4409, N4404, N3862, N2529, N2912);
or OR2 (N4410, N4400, N1310);
and AND3 (N4411, N4409, N3747, N1622);
nand NAND3 (N4412, N4399, N2366, N881);
buf BUF1 (N4413, N4410);
nor NOR3 (N4414, N4405, N2245, N1341);
nor NOR3 (N4415, N4406, N4216, N367);
or OR3 (N4416, N4413, N1964, N3565);
buf BUF1 (N4417, N4397);
and AND2 (N4418, N4411, N46);
xor XOR2 (N4419, N4418, N2441);
xor XOR2 (N4420, N4395, N4025);
and AND4 (N4421, N4403, N1043, N2048, N2275);
or OR3 (N4422, N4420, N607, N432);
xor XOR2 (N4423, N4415, N1026);
nor NOR3 (N4424, N4407, N2472, N2268);
and AND3 (N4425, N4412, N874, N1970);
buf BUF1 (N4426, N4414);
and AND2 (N4427, N4417, N409);
or OR2 (N4428, N4408, N118);
not NOT1 (N4429, N4425);
nand NAND2 (N4430, N4416, N2278);
buf BUF1 (N4431, N4424);
nor NOR4 (N4432, N4419, N2204, N2053, N1437);
and AND4 (N4433, N4428, N564, N3714, N2832);
buf BUF1 (N4434, N4431);
nor NOR4 (N4435, N4427, N2815, N1734, N366);
buf BUF1 (N4436, N4423);
buf BUF1 (N4437, N4436);
and AND3 (N4438, N4421, N630, N2005);
not NOT1 (N4439, N4426);
not NOT1 (N4440, N4429);
nor NOR3 (N4441, N4434, N2311, N1419);
and AND4 (N4442, N4422, N3479, N351, N2439);
and AND4 (N4443, N4432, N4096, N3150, N895);
xor XOR2 (N4444, N4438, N222);
not NOT1 (N4445, N4439);
not NOT1 (N4446, N4435);
nor NOR2 (N4447, N4442, N3005);
xor XOR2 (N4448, N4445, N2611);
not NOT1 (N4449, N4437);
or OR2 (N4450, N4449, N2678);
xor XOR2 (N4451, N4447, N3558);
buf BUF1 (N4452, N4450);
or OR2 (N4453, N4430, N42);
nor NOR4 (N4454, N4433, N3298, N3891, N1525);
xor XOR2 (N4455, N4444, N199);
or OR2 (N4456, N4446, N2339);
or OR2 (N4457, N4455, N805);
not NOT1 (N4458, N4454);
or OR3 (N4459, N4452, N1984, N2504);
xor XOR2 (N4460, N4453, N2276);
nand NAND2 (N4461, N4443, N3972);
nand NAND3 (N4462, N4448, N2442, N513);
not NOT1 (N4463, N4459);
not NOT1 (N4464, N4462);
and AND4 (N4465, N4440, N3751, N646, N2575);
nor NOR4 (N4466, N4456, N1103, N2473, N1062);
or OR4 (N4467, N4465, N3553, N2170, N2347);
nor NOR2 (N4468, N4451, N929);
and AND3 (N4469, N4461, N387, N298);
not NOT1 (N4470, N4468);
nor NOR3 (N4471, N4458, N3603, N1087);
buf BUF1 (N4472, N4467);
not NOT1 (N4473, N4466);
nand NAND2 (N4474, N4441, N4395);
nor NOR3 (N4475, N4471, N3337, N1895);
or OR3 (N4476, N4457, N1505, N1838);
not NOT1 (N4477, N4472);
xor XOR2 (N4478, N4460, N427);
nand NAND4 (N4479, N4470, N2122, N1232, N2183);
nand NAND2 (N4480, N4478, N1279);
and AND2 (N4481, N4475, N2278);
or OR4 (N4482, N4481, N316, N3497, N1405);
not NOT1 (N4483, N4479);
or OR3 (N4484, N4469, N576, N2545);
xor XOR2 (N4485, N4476, N2189);
nor NOR3 (N4486, N4477, N3129, N2945);
not NOT1 (N4487, N4486);
nor NOR4 (N4488, N4464, N1809, N1569, N355);
or OR2 (N4489, N4463, N3692);
xor XOR2 (N4490, N4482, N1478);
xor XOR2 (N4491, N4487, N31);
or OR2 (N4492, N4491, N1515);
buf BUF1 (N4493, N4483);
nor NOR2 (N4494, N4488, N3171);
and AND4 (N4495, N4473, N1142, N3178, N705);
nor NOR4 (N4496, N4494, N4235, N2883, N1935);
xor XOR2 (N4497, N4496, N1312);
or OR3 (N4498, N4480, N1590, N2792);
or OR3 (N4499, N4498, N23, N485);
buf BUF1 (N4500, N4490);
and AND4 (N4501, N4489, N2040, N613, N515);
or OR4 (N4502, N4499, N1898, N1106, N21);
not NOT1 (N4503, N4495);
and AND2 (N4504, N4492, N3294);
not NOT1 (N4505, N4497);
not NOT1 (N4506, N4493);
or OR4 (N4507, N4503, N3412, N4465, N3555);
nand NAND4 (N4508, N4504, N4300, N32, N2090);
buf BUF1 (N4509, N4508);
nor NOR3 (N4510, N4484, N1438, N4289);
or OR2 (N4511, N4505, N1823);
nand NAND2 (N4512, N4501, N4244);
nor NOR3 (N4513, N4512, N3736, N1945);
and AND3 (N4514, N4474, N3777, N4456);
nand NAND4 (N4515, N4511, N2103, N159, N3991);
xor XOR2 (N4516, N4515, N80);
nor NOR3 (N4517, N4485, N4307, N2297);
buf BUF1 (N4518, N4514);
and AND3 (N4519, N4507, N1259, N2635);
nand NAND4 (N4520, N4516, N4072, N3321, N3572);
not NOT1 (N4521, N4513);
and AND3 (N4522, N4509, N1565, N3209);
nor NOR3 (N4523, N4510, N1026, N1403);
buf BUF1 (N4524, N4519);
nand NAND4 (N4525, N4500, N2075, N4001, N3211);
nand NAND4 (N4526, N4520, N3754, N1197, N810);
nand NAND2 (N4527, N4517, N295);
buf BUF1 (N4528, N4522);
or OR4 (N4529, N4528, N493, N2214, N632);
nand NAND2 (N4530, N4502, N3180);
buf BUF1 (N4531, N4530);
nand NAND3 (N4532, N4523, N3453, N3143);
nand NAND3 (N4533, N4532, N2059, N4013);
nor NOR3 (N4534, N4526, N270, N3071);
buf BUF1 (N4535, N4521);
xor XOR2 (N4536, N4533, N117);
buf BUF1 (N4537, N4536);
nor NOR4 (N4538, N4534, N3967, N1428, N1174);
xor XOR2 (N4539, N4506, N775);
and AND2 (N4540, N4535, N2414);
nor NOR2 (N4541, N4537, N708);
xor XOR2 (N4542, N4527, N3882);
not NOT1 (N4543, N4539);
not NOT1 (N4544, N4529);
buf BUF1 (N4545, N4524);
buf BUF1 (N4546, N4543);
nor NOR3 (N4547, N4541, N2863, N2325);
or OR3 (N4548, N4542, N4228, N3332);
nand NAND4 (N4549, N4540, N339, N1134, N3670);
and AND4 (N4550, N4548, N4431, N2788, N4403);
nand NAND3 (N4551, N4525, N3777, N2619);
nand NAND4 (N4552, N4538, N822, N2493, N2046);
and AND2 (N4553, N4551, N2937);
buf BUF1 (N4554, N4552);
buf BUF1 (N4555, N4553);
or OR4 (N4556, N4550, N4460, N930, N3774);
buf BUF1 (N4557, N4556);
nor NOR4 (N4558, N4531, N329, N1469, N1794);
buf BUF1 (N4559, N4549);
nand NAND4 (N4560, N4555, N2216, N304, N237);
not NOT1 (N4561, N4545);
not NOT1 (N4562, N4518);
nand NAND3 (N4563, N4562, N445, N3727);
not NOT1 (N4564, N4559);
and AND3 (N4565, N4564, N1500, N4103);
buf BUF1 (N4566, N4557);
buf BUF1 (N4567, N4546);
nand NAND3 (N4568, N4566, N4327, N1206);
xor XOR2 (N4569, N4567, N1641);
nand NAND4 (N4570, N4568, N4197, N1240, N3395);
and AND3 (N4571, N4544, N2116, N2055);
nand NAND2 (N4572, N4565, N3597);
or OR2 (N4573, N4572, N2467);
nand NAND2 (N4574, N4571, N2594);
buf BUF1 (N4575, N4563);
xor XOR2 (N4576, N4570, N3334);
nand NAND4 (N4577, N4547, N18, N2228, N2057);
nand NAND4 (N4578, N4577, N4141, N2431, N1076);
nor NOR4 (N4579, N4574, N1848, N512, N37);
nand NAND4 (N4580, N4560, N940, N3253, N2571);
buf BUF1 (N4581, N4579);
buf BUF1 (N4582, N4580);
and AND3 (N4583, N4576, N1170, N239);
not NOT1 (N4584, N4583);
and AND3 (N4585, N4561, N2102, N1723);
nand NAND3 (N4586, N4554, N1964, N4148);
and AND3 (N4587, N4581, N3889, N153);
nor NOR2 (N4588, N4586, N311);
and AND4 (N4589, N4578, N1788, N4327, N1536);
or OR3 (N4590, N4589, N4326, N3629);
nor NOR4 (N4591, N4573, N449, N2904, N1061);
nor NOR3 (N4592, N4588, N1148, N3783);
not NOT1 (N4593, N4584);
not NOT1 (N4594, N4591);
xor XOR2 (N4595, N4585, N4192);
nand NAND3 (N4596, N4558, N595, N2745);
not NOT1 (N4597, N4594);
xor XOR2 (N4598, N4569, N2111);
and AND2 (N4599, N4575, N1163);
xor XOR2 (N4600, N4587, N2560);
nor NOR4 (N4601, N4597, N702, N2152, N3302);
buf BUF1 (N4602, N4601);
and AND3 (N4603, N4599, N1322, N3807);
buf BUF1 (N4604, N4582);
nor NOR4 (N4605, N4604, N1252, N1701, N4254);
and AND3 (N4606, N4593, N1528, N1303);
not NOT1 (N4607, N4602);
nor NOR3 (N4608, N4600, N1710, N4542);
xor XOR2 (N4609, N4596, N1067);
xor XOR2 (N4610, N4606, N3241);
buf BUF1 (N4611, N4592);
and AND3 (N4612, N4598, N3610, N1587);
nand NAND3 (N4613, N4611, N2794, N262);
buf BUF1 (N4614, N4590);
nor NOR3 (N4615, N4595, N4444, N300);
and AND4 (N4616, N4603, N3336, N3118, N2483);
or OR4 (N4617, N4612, N3216, N3312, N1023);
xor XOR2 (N4618, N4605, N4185);
or OR2 (N4619, N4613, N2854);
xor XOR2 (N4620, N4614, N1812);
nor NOR3 (N4621, N4617, N1354, N877);
or OR2 (N4622, N4615, N2136);
nor NOR3 (N4623, N4609, N2581, N1236);
nand NAND3 (N4624, N4620, N73, N513);
not NOT1 (N4625, N4610);
buf BUF1 (N4626, N4624);
and AND4 (N4627, N4619, N512, N2210, N4190);
nor NOR2 (N4628, N4626, N3271);
xor XOR2 (N4629, N4628, N531);
xor XOR2 (N4630, N4627, N2222);
and AND2 (N4631, N4625, N3288);
xor XOR2 (N4632, N4618, N2884);
xor XOR2 (N4633, N4629, N888);
not NOT1 (N4634, N4607);
nor NOR3 (N4635, N4633, N134, N3944);
nand NAND2 (N4636, N4622, N963);
nand NAND3 (N4637, N4616, N6, N3951);
xor XOR2 (N4638, N4608, N4533);
buf BUF1 (N4639, N4634);
nor NOR3 (N4640, N4636, N3804, N638);
xor XOR2 (N4641, N4635, N3156);
nand NAND3 (N4642, N4639, N1507, N841);
and AND4 (N4643, N4638, N2856, N2185, N142);
nor NOR3 (N4644, N4623, N1098, N1156);
nor NOR3 (N4645, N4630, N1526, N4144);
or OR3 (N4646, N4645, N2806, N564);
and AND2 (N4647, N4641, N306);
not NOT1 (N4648, N4621);
xor XOR2 (N4649, N4637, N116);
nand NAND4 (N4650, N4649, N4493, N2419, N3906);
or OR4 (N4651, N4643, N2896, N2531, N3322);
and AND4 (N4652, N4650, N3771, N1544, N3479);
not NOT1 (N4653, N4632);
and AND3 (N4654, N4640, N299, N2099);
buf BUF1 (N4655, N4631);
xor XOR2 (N4656, N4646, N4504);
and AND4 (N4657, N4648, N4027, N614, N1699);
nand NAND3 (N4658, N4647, N3963, N1101);
buf BUF1 (N4659, N4653);
nor NOR4 (N4660, N4655, N4325, N2158, N2954);
and AND3 (N4661, N4652, N2078, N1627);
xor XOR2 (N4662, N4654, N1128);
nor NOR2 (N4663, N4658, N2408);
or OR4 (N4664, N4657, N702, N30, N137);
and AND3 (N4665, N4661, N1091, N2687);
and AND3 (N4666, N4651, N1502, N579);
and AND2 (N4667, N4664, N1871);
xor XOR2 (N4668, N4656, N396);
xor XOR2 (N4669, N4662, N1865);
nor NOR3 (N4670, N4663, N1108, N1969);
or OR2 (N4671, N4642, N1964);
xor XOR2 (N4672, N4671, N4260);
xor XOR2 (N4673, N4666, N3053);
buf BUF1 (N4674, N4669);
and AND3 (N4675, N4667, N1943, N627);
or OR2 (N4676, N4673, N2581);
not NOT1 (N4677, N4675);
xor XOR2 (N4678, N4644, N3989);
or OR4 (N4679, N4677, N3336, N4652, N3647);
or OR4 (N4680, N4659, N3097, N4081, N1190);
nor NOR4 (N4681, N4668, N2113, N1811, N4660);
nor NOR2 (N4682, N4253, N477);
and AND4 (N4683, N4670, N2185, N2775, N3001);
or OR3 (N4684, N4678, N4250, N1222);
not NOT1 (N4685, N4682);
nand NAND2 (N4686, N4672, N316);
or OR4 (N4687, N4679, N2090, N3286, N3996);
not NOT1 (N4688, N4687);
buf BUF1 (N4689, N4665);
not NOT1 (N4690, N4681);
not NOT1 (N4691, N4685);
buf BUF1 (N4692, N4684);
and AND3 (N4693, N4674, N1532, N1265);
not NOT1 (N4694, N4692);
nor NOR3 (N4695, N4694, N713, N801);
nor NOR4 (N4696, N4676, N1524, N545, N1312);
and AND2 (N4697, N4680, N2228);
buf BUF1 (N4698, N4693);
xor XOR2 (N4699, N4697, N267);
not NOT1 (N4700, N4683);
not NOT1 (N4701, N4688);
xor XOR2 (N4702, N4701, N2720);
and AND3 (N4703, N4699, N1976, N4009);
or OR3 (N4704, N4691, N620, N3183);
xor XOR2 (N4705, N4700, N977);
xor XOR2 (N4706, N4690, N2828);
not NOT1 (N4707, N4686);
or OR2 (N4708, N4696, N3694);
xor XOR2 (N4709, N4702, N2622);
or OR2 (N4710, N4703, N1893);
and AND4 (N4711, N4705, N104, N2755, N4253);
or OR4 (N4712, N4707, N1564, N2957, N2094);
not NOT1 (N4713, N4709);
and AND3 (N4714, N4710, N4477, N2375);
nand NAND4 (N4715, N4712, N3457, N334, N3578);
buf BUF1 (N4716, N4704);
xor XOR2 (N4717, N4698, N3079);
not NOT1 (N4718, N4708);
xor XOR2 (N4719, N4711, N1080);
xor XOR2 (N4720, N4718, N371);
not NOT1 (N4721, N4717);
nor NOR4 (N4722, N4716, N2089, N2832, N4387);
nand NAND2 (N4723, N4722, N2624);
xor XOR2 (N4724, N4713, N1314);
nor NOR3 (N4725, N4719, N874, N2048);
nand NAND3 (N4726, N4715, N2708, N993);
or OR3 (N4727, N4706, N2692, N4506);
and AND2 (N4728, N4727, N720);
not NOT1 (N4729, N4725);
buf BUF1 (N4730, N4724);
nand NAND4 (N4731, N4721, N2331, N4064, N317);
not NOT1 (N4732, N4714);
or OR3 (N4733, N4726, N4619, N2502);
xor XOR2 (N4734, N4731, N51);
nand NAND4 (N4735, N4695, N1034, N2544, N3829);
or OR3 (N4736, N4729, N3222, N4668);
buf BUF1 (N4737, N4736);
not NOT1 (N4738, N4723);
or OR3 (N4739, N4733, N3789, N1173);
and AND4 (N4740, N4737, N1638, N3017, N656);
nand NAND2 (N4741, N4740, N2482);
not NOT1 (N4742, N4689);
nor NOR3 (N4743, N4742, N3378, N4221);
or OR4 (N4744, N4730, N4307, N3621, N353);
or OR2 (N4745, N4743, N2011);
nand NAND4 (N4746, N4732, N2679, N950, N3941);
buf BUF1 (N4747, N4738);
nand NAND4 (N4748, N4735, N2593, N3420, N1286);
not NOT1 (N4749, N4744);
not NOT1 (N4750, N4720);
xor XOR2 (N4751, N4749, N4193);
and AND4 (N4752, N4747, N2517, N982, N62);
nor NOR3 (N4753, N4734, N2038, N4356);
and AND4 (N4754, N4750, N4152, N2288, N1242);
nand NAND4 (N4755, N4748, N4559, N2475, N1030);
not NOT1 (N4756, N4755);
not NOT1 (N4757, N4739);
and AND3 (N4758, N4752, N338, N3818);
xor XOR2 (N4759, N4754, N2582);
xor XOR2 (N4760, N4756, N2897);
nor NOR2 (N4761, N4760, N3256);
not NOT1 (N4762, N4759);
and AND2 (N4763, N4762, N1263);
nor NOR4 (N4764, N4763, N2302, N1859, N3339);
nor NOR4 (N4765, N4728, N91, N3835, N156);
not NOT1 (N4766, N4761);
or OR4 (N4767, N4745, N3960, N199, N1109);
nand NAND2 (N4768, N4746, N3530);
nand NAND3 (N4769, N4751, N3583, N129);
and AND2 (N4770, N4768, N3109);
not NOT1 (N4771, N4767);
not NOT1 (N4772, N4769);
or OR3 (N4773, N4757, N4721, N1519);
xor XOR2 (N4774, N4772, N4149);
nand NAND4 (N4775, N4765, N1061, N2326, N4115);
nor NOR3 (N4776, N4766, N2051, N3951);
or OR2 (N4777, N4764, N2046);
xor XOR2 (N4778, N4776, N2841);
xor XOR2 (N4779, N4771, N3095);
and AND3 (N4780, N4779, N4528, N1008);
and AND2 (N4781, N4758, N901);
not NOT1 (N4782, N4775);
nand NAND4 (N4783, N4773, N1780, N3382, N864);
not NOT1 (N4784, N4778);
and AND3 (N4785, N4753, N4230, N2069);
not NOT1 (N4786, N4781);
or OR2 (N4787, N4786, N4425);
and AND3 (N4788, N4782, N4223, N4143);
and AND3 (N4789, N4774, N214, N1218);
not NOT1 (N4790, N4780);
nor NOR3 (N4791, N4789, N527, N3137);
and AND2 (N4792, N4770, N3351);
and AND4 (N4793, N4784, N460, N4292, N1945);
not NOT1 (N4794, N4788);
or OR3 (N4795, N4787, N3399, N610);
buf BUF1 (N4796, N4785);
and AND3 (N4797, N4792, N3077, N1442);
and AND3 (N4798, N4796, N1276, N3496);
nor NOR3 (N4799, N4777, N954, N4749);
xor XOR2 (N4800, N4798, N4367);
or OR3 (N4801, N4793, N1086, N1491);
xor XOR2 (N4802, N4795, N2900);
or OR2 (N4803, N4790, N1996);
xor XOR2 (N4804, N4801, N2571);
and AND3 (N4805, N4797, N1764, N857);
nand NAND2 (N4806, N4783, N393);
xor XOR2 (N4807, N4741, N3309);
and AND3 (N4808, N4802, N56, N656);
nor NOR3 (N4809, N4800, N760, N356);
not NOT1 (N4810, N4805);
or OR3 (N4811, N4809, N6, N2621);
or OR4 (N4812, N4807, N3249, N123, N3694);
and AND2 (N4813, N4811, N1724);
xor XOR2 (N4814, N4813, N3567);
not NOT1 (N4815, N4808);
nand NAND2 (N4816, N4814, N948);
or OR4 (N4817, N4812, N961, N1413, N3670);
xor XOR2 (N4818, N4817, N1258);
nor NOR4 (N4819, N4818, N3910, N2091, N921);
xor XOR2 (N4820, N4799, N3225);
or OR2 (N4821, N4794, N2204);
nor NOR2 (N4822, N4820, N4253);
and AND2 (N4823, N4816, N2592);
buf BUF1 (N4824, N4806);
buf BUF1 (N4825, N4819);
and AND4 (N4826, N4824, N967, N270, N3596);
buf BUF1 (N4827, N4822);
or OR2 (N4828, N4827, N4775);
buf BUF1 (N4829, N4810);
xor XOR2 (N4830, N4803, N1678);
buf BUF1 (N4831, N4830);
not NOT1 (N4832, N4828);
nand NAND4 (N4833, N4831, N1661, N934, N3929);
not NOT1 (N4834, N4825);
xor XOR2 (N4835, N4829, N3959);
nor NOR4 (N4836, N4821, N3797, N1756, N1828);
buf BUF1 (N4837, N4833);
nor NOR2 (N4838, N4837, N3243);
not NOT1 (N4839, N4832);
nand NAND2 (N4840, N4815, N1823);
and AND4 (N4841, N4823, N929, N1699, N265);
nor NOR4 (N4842, N4835, N2930, N4416, N1453);
buf BUF1 (N4843, N4840);
not NOT1 (N4844, N4804);
buf BUF1 (N4845, N4791);
xor XOR2 (N4846, N4839, N128);
buf BUF1 (N4847, N4836);
buf BUF1 (N4848, N4834);
nor NOR4 (N4849, N4844, N1901, N376, N3136);
nor NOR2 (N4850, N4848, N1628);
buf BUF1 (N4851, N4846);
and AND4 (N4852, N4843, N1211, N428, N3979);
buf BUF1 (N4853, N4842);
not NOT1 (N4854, N4852);
nor NOR2 (N4855, N4826, N3069);
not NOT1 (N4856, N4853);
and AND4 (N4857, N4847, N2988, N2512, N2436);
buf BUF1 (N4858, N4856);
and AND4 (N4859, N4855, N4680, N3500, N4251);
or OR4 (N4860, N4845, N2097, N602, N3613);
buf BUF1 (N4861, N4851);
not NOT1 (N4862, N4854);
nand NAND4 (N4863, N4841, N3422, N752, N2312);
nand NAND2 (N4864, N4860, N2786);
nor NOR3 (N4865, N4862, N680, N4338);
nand NAND4 (N4866, N4859, N2248, N2092, N1757);
not NOT1 (N4867, N4857);
nor NOR2 (N4868, N4866, N172);
xor XOR2 (N4869, N4867, N600);
or OR2 (N4870, N4850, N1741);
and AND2 (N4871, N4868, N1043);
xor XOR2 (N4872, N4858, N2269);
or OR2 (N4873, N4871, N3994);
nor NOR4 (N4874, N4863, N3276, N1932, N3596);
not NOT1 (N4875, N4870);
buf BUF1 (N4876, N4849);
or OR2 (N4877, N4874, N3843);
not NOT1 (N4878, N4869);
or OR2 (N4879, N4864, N252);
or OR3 (N4880, N4875, N4508, N2176);
and AND4 (N4881, N4879, N5, N3091, N4431);
xor XOR2 (N4882, N4873, N2635);
nand NAND4 (N4883, N4878, N3593, N2208, N1690);
nor NOR3 (N4884, N4838, N2156, N2714);
xor XOR2 (N4885, N4876, N1127);
and AND4 (N4886, N4865, N2919, N2799, N3499);
or OR4 (N4887, N4881, N562, N3542, N1509);
or OR4 (N4888, N4877, N3318, N2947, N2565);
and AND2 (N4889, N4880, N776);
not NOT1 (N4890, N4889);
and AND4 (N4891, N4882, N3534, N1842, N3793);
or OR2 (N4892, N4885, N3371);
nand NAND4 (N4893, N4888, N3607, N3032, N2420);
nor NOR3 (N4894, N4892, N3371, N697);
buf BUF1 (N4895, N4887);
nor NOR2 (N4896, N4872, N4887);
not NOT1 (N4897, N4861);
buf BUF1 (N4898, N4890);
nor NOR3 (N4899, N4895, N3032, N705);
nand NAND2 (N4900, N4899, N1677);
nand NAND2 (N4901, N4891, N587);
buf BUF1 (N4902, N4900);
or OR3 (N4903, N4894, N4879, N4448);
or OR4 (N4904, N4901, N3166, N3644, N3806);
and AND3 (N4905, N4902, N3966, N2753);
buf BUF1 (N4906, N4898);
or OR3 (N4907, N4886, N2694, N3586);
nor NOR4 (N4908, N4883, N4019, N3298, N4068);
xor XOR2 (N4909, N4905, N3570);
and AND3 (N4910, N4907, N2366, N4730);
not NOT1 (N4911, N4908);
xor XOR2 (N4912, N4910, N2520);
or OR4 (N4913, N4903, N3648, N3034, N2468);
buf BUF1 (N4914, N4909);
xor XOR2 (N4915, N4911, N4891);
xor XOR2 (N4916, N4897, N3763);
nand NAND4 (N4917, N4912, N563, N2449, N4785);
xor XOR2 (N4918, N4904, N4397);
not NOT1 (N4919, N4913);
nand NAND2 (N4920, N4884, N199);
xor XOR2 (N4921, N4919, N599);
and AND4 (N4922, N4920, N4009, N1643, N3230);
nand NAND4 (N4923, N4918, N3314, N4433, N123);
or OR2 (N4924, N4916, N4438);
nor NOR4 (N4925, N4921, N1628, N463, N1115);
xor XOR2 (N4926, N4924, N4887);
and AND3 (N4927, N4923, N873, N4044);
xor XOR2 (N4928, N4927, N530);
and AND3 (N4929, N4915, N1686, N82);
and AND4 (N4930, N4926, N2548, N526, N3358);
and AND4 (N4931, N4893, N3403, N2670, N2516);
nand NAND3 (N4932, N4925, N4409, N2147);
nor NOR3 (N4933, N4917, N383, N1299);
or OR4 (N4934, N4928, N4926, N445, N3417);
buf BUF1 (N4935, N4922);
buf BUF1 (N4936, N4929);
buf BUF1 (N4937, N4930);
buf BUF1 (N4938, N4937);
xor XOR2 (N4939, N4935, N998);
not NOT1 (N4940, N4914);
or OR3 (N4941, N4906, N575, N2972);
nor NOR2 (N4942, N4941, N2555);
and AND2 (N4943, N4934, N1782);
nand NAND2 (N4944, N4943, N3107);
nor NOR2 (N4945, N4942, N4844);
nor NOR4 (N4946, N4936, N2083, N1453, N530);
and AND2 (N4947, N4933, N1003);
buf BUF1 (N4948, N4945);
not NOT1 (N4949, N4896);
not NOT1 (N4950, N4948);
nand NAND2 (N4951, N4944, N1327);
not NOT1 (N4952, N4949);
or OR2 (N4953, N4952, N2936);
not NOT1 (N4954, N4931);
and AND2 (N4955, N4946, N3578);
buf BUF1 (N4956, N4951);
xor XOR2 (N4957, N4939, N2270);
buf BUF1 (N4958, N4955);
buf BUF1 (N4959, N4950);
xor XOR2 (N4960, N4953, N2532);
or OR3 (N4961, N4959, N1370, N3358);
and AND3 (N4962, N4957, N1203, N4318);
xor XOR2 (N4963, N4961, N731);
xor XOR2 (N4964, N4958, N1938);
not NOT1 (N4965, N4962);
and AND3 (N4966, N4960, N3015, N4501);
buf BUF1 (N4967, N4938);
nand NAND4 (N4968, N4964, N1588, N186, N1953);
nand NAND3 (N4969, N4966, N3777, N64);
nand NAND2 (N4970, N4969, N4904);
nor NOR3 (N4971, N4954, N1038, N3046);
not NOT1 (N4972, N4940);
nand NAND2 (N4973, N4965, N1389);
xor XOR2 (N4974, N4972, N3260);
buf BUF1 (N4975, N4947);
and AND2 (N4976, N4973, N3439);
nor NOR4 (N4977, N4975, N2236, N602, N1025);
nand NAND4 (N4978, N4977, N486, N1227, N4297);
xor XOR2 (N4979, N4932, N79);
buf BUF1 (N4980, N4963);
or OR4 (N4981, N4979, N3886, N3411, N1014);
xor XOR2 (N4982, N4981, N1405);
or OR2 (N4983, N4976, N241);
xor XOR2 (N4984, N4982, N1258);
buf BUF1 (N4985, N4967);
or OR3 (N4986, N4974, N2791, N2745);
buf BUF1 (N4987, N4986);
or OR2 (N4988, N4968, N205);
nor NOR4 (N4989, N4987, N3918, N4895, N450);
and AND2 (N4990, N4988, N1222);
xor XOR2 (N4991, N4989, N2081);
nor NOR4 (N4992, N4980, N2875, N2137, N3055);
and AND2 (N4993, N4983, N3465);
nor NOR2 (N4994, N4984, N4006);
buf BUF1 (N4995, N4978);
nand NAND4 (N4996, N4992, N430, N4145, N3112);
nor NOR4 (N4997, N4956, N3410, N1493, N777);
nor NOR4 (N4998, N4971, N2637, N62, N3143);
buf BUF1 (N4999, N4995);
nor NOR4 (N5000, N4997, N3734, N365, N3599);
nand NAND3 (N5001, N5000, N1083, N708);
buf BUF1 (N5002, N4993);
not NOT1 (N5003, N4970);
not NOT1 (N5004, N4994);
and AND3 (N5005, N4990, N4706, N1280);
xor XOR2 (N5006, N5004, N3425);
nand NAND4 (N5007, N4998, N2905, N1415, N4283);
or OR4 (N5008, N5005, N3134, N3275, N922);
not NOT1 (N5009, N5003);
xor XOR2 (N5010, N5007, N3254);
xor XOR2 (N5011, N4991, N2746);
nand NAND2 (N5012, N5011, N4609);
not NOT1 (N5013, N5006);
xor XOR2 (N5014, N5002, N22);
nand NAND2 (N5015, N5009, N2407);
not NOT1 (N5016, N5013);
nor NOR4 (N5017, N5016, N4865, N1247, N768);
or OR2 (N5018, N5014, N2946);
nor NOR2 (N5019, N4996, N1800);
or OR2 (N5020, N5012, N2253);
not NOT1 (N5021, N5020);
and AND2 (N5022, N5015, N4599);
and AND2 (N5023, N5019, N2094);
or OR4 (N5024, N5021, N586, N1186, N3963);
buf BUF1 (N5025, N4985);
or OR4 (N5026, N5023, N3092, N3026, N319);
and AND2 (N5027, N5008, N3866);
nand NAND4 (N5028, N5022, N1280, N1879, N3530);
buf BUF1 (N5029, N5018);
and AND3 (N5030, N5024, N3407, N4895);
nor NOR2 (N5031, N5001, N4367);
buf BUF1 (N5032, N5010);
nand NAND2 (N5033, N5017, N4554);
not NOT1 (N5034, N5025);
nor NOR2 (N5035, N5033, N2695);
nand NAND3 (N5036, N5029, N186, N1827);
xor XOR2 (N5037, N5026, N2196);
and AND2 (N5038, N5037, N1796);
xor XOR2 (N5039, N5031, N672);
not NOT1 (N5040, N4999);
nor NOR2 (N5041, N5039, N1867);
xor XOR2 (N5042, N5041, N214);
and AND3 (N5043, N5032, N2152, N4019);
not NOT1 (N5044, N5040);
nor NOR3 (N5045, N5027, N3010, N880);
xor XOR2 (N5046, N5043, N1701);
or OR2 (N5047, N5030, N844);
or OR4 (N5048, N5028, N448, N5014, N4542);
nand NAND3 (N5049, N5036, N3168, N4707);
nor NOR3 (N5050, N5042, N1753, N4496);
buf BUF1 (N5051, N5046);
or OR3 (N5052, N5034, N3487, N4949);
and AND4 (N5053, N5052, N3450, N4671, N69);
and AND3 (N5054, N5047, N805, N4760);
xor XOR2 (N5055, N5038, N418);
nand NAND4 (N5056, N5048, N4474, N4840, N3483);
or OR2 (N5057, N5054, N1546);
nor NOR4 (N5058, N5044, N4021, N742, N3859);
and AND4 (N5059, N5035, N3886, N324, N1776);
nor NOR3 (N5060, N5053, N1009, N1151);
not NOT1 (N5061, N5050);
nor NOR2 (N5062, N5055, N52);
and AND2 (N5063, N5058, N201);
and AND3 (N5064, N5062, N1347, N4183);
and AND2 (N5065, N5064, N2711);
nor NOR2 (N5066, N5057, N3218);
not NOT1 (N5067, N5066);
nand NAND2 (N5068, N5045, N3232);
nand NAND2 (N5069, N5061, N2667);
or OR3 (N5070, N5063, N2977, N104);
and AND2 (N5071, N5060, N1724);
buf BUF1 (N5072, N5049);
nor NOR4 (N5073, N5068, N822, N3909, N2163);
buf BUF1 (N5074, N5051);
and AND4 (N5075, N5070, N5010, N4977, N4537);
or OR2 (N5076, N5067, N1516);
or OR4 (N5077, N5076, N3740, N244, N2394);
or OR2 (N5078, N5059, N4820);
buf BUF1 (N5079, N5075);
or OR2 (N5080, N5071, N525);
nor NOR3 (N5081, N5074, N4976, N309);
nor NOR4 (N5082, N5056, N2484, N4047, N2318);
buf BUF1 (N5083, N5080);
xor XOR2 (N5084, N5073, N969);
buf BUF1 (N5085, N5081);
or OR3 (N5086, N5078, N5005, N2706);
not NOT1 (N5087, N5084);
nand NAND3 (N5088, N5086, N3288, N4198);
nor NOR3 (N5089, N5088, N3007, N3670);
nor NOR2 (N5090, N5065, N136);
and AND3 (N5091, N5089, N17, N4487);
nand NAND4 (N5092, N5087, N4661, N4789, N955);
xor XOR2 (N5093, N5085, N409);
nor NOR2 (N5094, N5079, N736);
not NOT1 (N5095, N5093);
nor NOR3 (N5096, N5077, N4948, N3986);
nor NOR3 (N5097, N5069, N2933, N4877);
or OR2 (N5098, N5097, N4372);
not NOT1 (N5099, N5090);
nand NAND4 (N5100, N5099, N1693, N3667, N4885);
nand NAND2 (N5101, N5092, N106);
and AND2 (N5102, N5096, N2675);
xor XOR2 (N5103, N5095, N2386);
or OR4 (N5104, N5094, N2075, N1185, N4629);
or OR4 (N5105, N5072, N330, N527, N4637);
and AND4 (N5106, N5101, N4863, N3758, N3154);
and AND4 (N5107, N5091, N2155, N683, N2661);
and AND3 (N5108, N5107, N109, N1452);
and AND3 (N5109, N5100, N811, N1360);
xor XOR2 (N5110, N5104, N3449);
or OR3 (N5111, N5102, N2343, N5040);
not NOT1 (N5112, N5110);
nor NOR4 (N5113, N5103, N3716, N4349, N3455);
and AND3 (N5114, N5111, N3276, N724);
not NOT1 (N5115, N5114);
buf BUF1 (N5116, N5115);
nand NAND4 (N5117, N5116, N1283, N2716, N2517);
nand NAND2 (N5118, N5082, N279);
or OR3 (N5119, N5108, N4128, N3721);
buf BUF1 (N5120, N5118);
and AND4 (N5121, N5098, N396, N976, N2127);
buf BUF1 (N5122, N5112);
xor XOR2 (N5123, N5122, N1692);
nor NOR3 (N5124, N5119, N4785, N4833);
or OR3 (N5125, N5120, N382, N4926);
xor XOR2 (N5126, N5125, N5090);
not NOT1 (N5127, N5105);
or OR3 (N5128, N5083, N1803, N107);
xor XOR2 (N5129, N5117, N4394);
xor XOR2 (N5130, N5123, N3427);
not NOT1 (N5131, N5129);
not NOT1 (N5132, N5130);
and AND2 (N5133, N5121, N1849);
nand NAND4 (N5134, N5131, N1034, N4983, N1872);
or OR2 (N5135, N5113, N1737);
or OR3 (N5136, N5132, N2248, N69);
xor XOR2 (N5137, N5133, N2190);
nand NAND3 (N5138, N5134, N3631, N303);
and AND2 (N5139, N5136, N1323);
xor XOR2 (N5140, N5126, N2354);
and AND4 (N5141, N5138, N190, N417, N5021);
not NOT1 (N5142, N5139);
not NOT1 (N5143, N5142);
not NOT1 (N5144, N5140);
not NOT1 (N5145, N5109);
buf BUF1 (N5146, N5143);
and AND4 (N5147, N5128, N2258, N4436, N3908);
nand NAND4 (N5148, N5145, N4747, N3811, N551);
nor NOR3 (N5149, N5124, N643, N2855);
nor NOR3 (N5150, N5137, N4700, N1546);
nor NOR3 (N5151, N5135, N4256, N4787);
nand NAND4 (N5152, N5144, N1970, N3219, N975);
buf BUF1 (N5153, N5106);
not NOT1 (N5154, N5146);
not NOT1 (N5155, N5127);
buf BUF1 (N5156, N5141);
nand NAND4 (N5157, N5150, N1452, N1291, N1239);
or OR3 (N5158, N5149, N2697, N1532);
xor XOR2 (N5159, N5156, N3319);
nand NAND4 (N5160, N5157, N4921, N1684, N2451);
buf BUF1 (N5161, N5147);
nor NOR2 (N5162, N5155, N1577);
nor NOR3 (N5163, N5152, N4527, N3704);
nor NOR3 (N5164, N5162, N2821, N2732);
buf BUF1 (N5165, N5164);
or OR3 (N5166, N5148, N1524, N697);
not NOT1 (N5167, N5159);
and AND2 (N5168, N5163, N3702);
nand NAND3 (N5169, N5161, N5001, N253);
not NOT1 (N5170, N5166);
nor NOR3 (N5171, N5169, N1306, N2765);
buf BUF1 (N5172, N5153);
xor XOR2 (N5173, N5165, N3957);
and AND2 (N5174, N5170, N4165);
buf BUF1 (N5175, N5173);
not NOT1 (N5176, N5175);
and AND3 (N5177, N5151, N4511, N345);
xor XOR2 (N5178, N5160, N1088);
nand NAND4 (N5179, N5177, N3884, N491, N4219);
nor NOR4 (N5180, N5154, N1264, N3120, N1284);
xor XOR2 (N5181, N5167, N3951);
and AND3 (N5182, N5181, N2592, N1111);
nor NOR4 (N5183, N5172, N568, N462, N4972);
or OR2 (N5184, N5179, N100);
buf BUF1 (N5185, N5180);
buf BUF1 (N5186, N5185);
or OR3 (N5187, N5174, N878, N4759);
nor NOR3 (N5188, N5168, N2093, N3971);
not NOT1 (N5189, N5171);
and AND3 (N5190, N5187, N92, N1499);
xor XOR2 (N5191, N5188, N2873);
nor NOR2 (N5192, N5190, N2625);
or OR2 (N5193, N5182, N3442);
or OR4 (N5194, N5189, N1993, N502, N3828);
xor XOR2 (N5195, N5191, N4673);
nor NOR2 (N5196, N5192, N4023);
or OR2 (N5197, N5183, N683);
xor XOR2 (N5198, N5184, N1995);
not NOT1 (N5199, N5194);
not NOT1 (N5200, N5186);
buf BUF1 (N5201, N5176);
nor NOR3 (N5202, N5200, N851, N2575);
not NOT1 (N5203, N5202);
nor NOR2 (N5204, N5178, N4885);
or OR3 (N5205, N5193, N2592, N2821);
xor XOR2 (N5206, N5196, N609);
nor NOR3 (N5207, N5206, N261, N4070);
nand NAND3 (N5208, N5158, N14, N3199);
and AND4 (N5209, N5205, N2406, N1191, N2533);
not NOT1 (N5210, N5201);
or OR4 (N5211, N5198, N394, N1593, N4206);
nor NOR2 (N5212, N5204, N4041);
not NOT1 (N5213, N5212);
or OR3 (N5214, N5213, N1525, N1605);
xor XOR2 (N5215, N5197, N941);
nor NOR2 (N5216, N5203, N3471);
nand NAND4 (N5217, N5211, N225, N457, N4353);
nor NOR3 (N5218, N5208, N4435, N2002);
nor NOR3 (N5219, N5218, N3166, N1812);
and AND4 (N5220, N5215, N116, N2294, N3306);
and AND2 (N5221, N5219, N5005);
xor XOR2 (N5222, N5216, N1806);
nand NAND3 (N5223, N5214, N4849, N760);
buf BUF1 (N5224, N5199);
xor XOR2 (N5225, N5209, N306);
or OR2 (N5226, N5223, N2679);
not NOT1 (N5227, N5220);
not NOT1 (N5228, N5224);
not NOT1 (N5229, N5195);
xor XOR2 (N5230, N5227, N128);
xor XOR2 (N5231, N5221, N4147);
and AND4 (N5232, N5225, N3146, N5126, N1215);
nor NOR2 (N5233, N5232, N1103);
and AND4 (N5234, N5226, N1497, N555, N4925);
or OR2 (N5235, N5231, N1879);
xor XOR2 (N5236, N5207, N5176);
nand NAND3 (N5237, N5228, N752, N3823);
and AND2 (N5238, N5236, N2822);
nand NAND2 (N5239, N5234, N1514);
nand NAND3 (N5240, N5210, N119, N2254);
or OR2 (N5241, N5235, N4077);
or OR3 (N5242, N5241, N3774, N558);
or OR3 (N5243, N5230, N1108, N734);
not NOT1 (N5244, N5239);
or OR4 (N5245, N5238, N597, N2245, N602);
not NOT1 (N5246, N5244);
buf BUF1 (N5247, N5222);
nand NAND2 (N5248, N5246, N5173);
or OR3 (N5249, N5242, N4923, N951);
and AND3 (N5250, N5243, N1993, N1011);
nand NAND3 (N5251, N5247, N830, N198);
and AND3 (N5252, N5248, N4194, N3950);
xor XOR2 (N5253, N5229, N694);
nand NAND4 (N5254, N5252, N110, N3560, N3735);
and AND2 (N5255, N5250, N290);
and AND4 (N5256, N5253, N1434, N3125, N291);
buf BUF1 (N5257, N5217);
or OR4 (N5258, N5256, N3302, N4782, N2592);
not NOT1 (N5259, N5251);
and AND4 (N5260, N5233, N5097, N1242, N3471);
xor XOR2 (N5261, N5254, N4947);
not NOT1 (N5262, N5255);
or OR2 (N5263, N5257, N2664);
xor XOR2 (N5264, N5262, N4734);
not NOT1 (N5265, N5245);
not NOT1 (N5266, N5258);
xor XOR2 (N5267, N5240, N3378);
or OR3 (N5268, N5259, N2129, N5208);
nor NOR2 (N5269, N5267, N5080);
or OR2 (N5270, N5237, N18);
xor XOR2 (N5271, N5266, N1795);
not NOT1 (N5272, N5268);
buf BUF1 (N5273, N5264);
nor NOR3 (N5274, N5270, N2577, N3650);
nand NAND3 (N5275, N5273, N4039, N4219);
nand NAND2 (N5276, N5271, N1563);
not NOT1 (N5277, N5272);
xor XOR2 (N5278, N5269, N1013);
xor XOR2 (N5279, N5265, N2612);
not NOT1 (N5280, N5274);
xor XOR2 (N5281, N5278, N1440);
buf BUF1 (N5282, N5275);
nor NOR3 (N5283, N5281, N2937, N2213);
xor XOR2 (N5284, N5282, N2104);
or OR3 (N5285, N5260, N306, N5150);
not NOT1 (N5286, N5283);
and AND2 (N5287, N5261, N4871);
and AND2 (N5288, N5286, N1165);
nand NAND2 (N5289, N5249, N3918);
or OR2 (N5290, N5277, N1662);
or OR4 (N5291, N5289, N4193, N2044, N3171);
buf BUF1 (N5292, N5276);
and AND4 (N5293, N5263, N5022, N1183, N4);
xor XOR2 (N5294, N5284, N4047);
and AND4 (N5295, N5291, N4950, N5141, N2076);
nor NOR2 (N5296, N5292, N2050);
or OR3 (N5297, N5295, N4889, N1676);
xor XOR2 (N5298, N5290, N3893);
nor NOR4 (N5299, N5293, N3189, N4615, N2400);
and AND3 (N5300, N5299, N5139, N134);
xor XOR2 (N5301, N5287, N2929);
and AND2 (N5302, N5300, N1138);
buf BUF1 (N5303, N5279);
nor NOR4 (N5304, N5303, N5081, N3229, N365);
and AND3 (N5305, N5304, N429, N446);
or OR3 (N5306, N5301, N4501, N999);
buf BUF1 (N5307, N5297);
or OR3 (N5308, N5306, N763, N3942);
not NOT1 (N5309, N5298);
not NOT1 (N5310, N5305);
and AND2 (N5311, N5307, N3192);
xor XOR2 (N5312, N5296, N608);
nand NAND4 (N5313, N5310, N317, N5299, N3980);
or OR3 (N5314, N5288, N678, N657);
buf BUF1 (N5315, N5311);
and AND3 (N5316, N5294, N995, N4191);
buf BUF1 (N5317, N5285);
xor XOR2 (N5318, N5302, N3184);
xor XOR2 (N5319, N5316, N3043);
not NOT1 (N5320, N5319);
and AND4 (N5321, N5309, N188, N3659, N1617);
nor NOR3 (N5322, N5312, N3886, N794);
xor XOR2 (N5323, N5320, N205);
and AND3 (N5324, N5314, N3972, N5095);
or OR3 (N5325, N5324, N369, N423);
or OR4 (N5326, N5318, N1788, N1389, N5095);
and AND2 (N5327, N5280, N2807);
nand NAND2 (N5328, N5315, N3768);
nand NAND4 (N5329, N5327, N2781, N392, N4973);
or OR4 (N5330, N5308, N1564, N2524, N113);
nor NOR2 (N5331, N5328, N908);
nor NOR3 (N5332, N5325, N1383, N3781);
xor XOR2 (N5333, N5329, N4111);
not NOT1 (N5334, N5317);
xor XOR2 (N5335, N5330, N254);
xor XOR2 (N5336, N5323, N3750);
nor NOR3 (N5337, N5332, N1812, N2927);
buf BUF1 (N5338, N5321);
xor XOR2 (N5339, N5313, N3603);
nand NAND3 (N5340, N5335, N4382, N2899);
or OR3 (N5341, N5331, N848, N1858);
xor XOR2 (N5342, N5334, N1);
not NOT1 (N5343, N5341);
not NOT1 (N5344, N5336);
not NOT1 (N5345, N5338);
and AND2 (N5346, N5339, N2345);
and AND3 (N5347, N5337, N397, N106);
nor NOR2 (N5348, N5345, N5236);
or OR2 (N5349, N5322, N3873);
nand NAND3 (N5350, N5333, N2990, N1993);
nor NOR4 (N5351, N5348, N2932, N4729, N4745);
nand NAND3 (N5352, N5347, N4082, N2313);
xor XOR2 (N5353, N5350, N4891);
or OR4 (N5354, N5340, N4954, N1970, N1207);
not NOT1 (N5355, N5349);
nand NAND3 (N5356, N5343, N726, N2623);
buf BUF1 (N5357, N5356);
nand NAND3 (N5358, N5342, N1211, N668);
buf BUF1 (N5359, N5357);
nand NAND2 (N5360, N5326, N175);
not NOT1 (N5361, N5352);
or OR3 (N5362, N5355, N3188, N2390);
xor XOR2 (N5363, N5354, N1535);
and AND3 (N5364, N5359, N3064, N3690);
buf BUF1 (N5365, N5353);
buf BUF1 (N5366, N5358);
nor NOR3 (N5367, N5360, N2645, N200);
or OR3 (N5368, N5364, N3177, N3444);
buf BUF1 (N5369, N5361);
or OR3 (N5370, N5368, N1311, N982);
nand NAND2 (N5371, N5363, N3803);
or OR3 (N5372, N5369, N4658, N2655);
xor XOR2 (N5373, N5371, N2799);
or OR4 (N5374, N5372, N3040, N697, N846);
nand NAND4 (N5375, N5362, N2012, N3562, N4534);
xor XOR2 (N5376, N5370, N4029);
and AND2 (N5377, N5344, N1905);
and AND2 (N5378, N5351, N1606);
xor XOR2 (N5379, N5367, N3573);
and AND4 (N5380, N5375, N2190, N2581, N3940);
and AND2 (N5381, N5346, N4835);
xor XOR2 (N5382, N5366, N4229);
nor NOR4 (N5383, N5376, N4767, N5142, N3718);
and AND2 (N5384, N5383, N3381);
or OR3 (N5385, N5378, N2292, N4763);
xor XOR2 (N5386, N5374, N5233);
not NOT1 (N5387, N5384);
or OR4 (N5388, N5377, N5006, N1756, N3857);
nor NOR4 (N5389, N5388, N4324, N1816, N2851);
and AND3 (N5390, N5389, N2543, N4513);
xor XOR2 (N5391, N5365, N1099);
or OR2 (N5392, N5390, N920);
not NOT1 (N5393, N5373);
and AND2 (N5394, N5393, N68);
nor NOR3 (N5395, N5380, N2156, N1435);
nand NAND4 (N5396, N5392, N5032, N2649, N2995);
nor NOR4 (N5397, N5385, N3119, N200, N3046);
not NOT1 (N5398, N5395);
nor NOR3 (N5399, N5382, N1376, N403);
nand NAND3 (N5400, N5391, N4276, N3067);
nand NAND3 (N5401, N5396, N2306, N4402);
nand NAND3 (N5402, N5400, N2183, N3732);
buf BUF1 (N5403, N5379);
or OR2 (N5404, N5397, N4425);
xor XOR2 (N5405, N5402, N1575);
or OR3 (N5406, N5386, N4449, N1415);
and AND4 (N5407, N5399, N4924, N4633, N3364);
and AND3 (N5408, N5406, N2032, N4225);
or OR4 (N5409, N5403, N1438, N4243, N1123);
nor NOR4 (N5410, N5398, N3698, N2543, N1803);
xor XOR2 (N5411, N5405, N2153);
buf BUF1 (N5412, N5408);
or OR4 (N5413, N5410, N471, N1542, N1367);
or OR3 (N5414, N5412, N4719, N130);
xor XOR2 (N5415, N5404, N1194);
nand NAND4 (N5416, N5381, N5191, N2227, N3701);
nor NOR2 (N5417, N5394, N641);
xor XOR2 (N5418, N5407, N266);
xor XOR2 (N5419, N5413, N2380);
buf BUF1 (N5420, N5411);
xor XOR2 (N5421, N5401, N4127);
and AND3 (N5422, N5418, N1802, N3827);
nor NOR4 (N5423, N5416, N695, N1507, N3206);
not NOT1 (N5424, N5415);
nor NOR3 (N5425, N5419, N1043, N2457);
nor NOR3 (N5426, N5414, N3092, N366);
and AND3 (N5427, N5421, N1344, N4808);
buf BUF1 (N5428, N5409);
nor NOR3 (N5429, N5417, N888, N3105);
buf BUF1 (N5430, N5426);
xor XOR2 (N5431, N5423, N746);
nor NOR2 (N5432, N5429, N201);
buf BUF1 (N5433, N5428);
buf BUF1 (N5434, N5433);
xor XOR2 (N5435, N5427, N3953);
and AND3 (N5436, N5424, N3825, N4132);
and AND3 (N5437, N5430, N2651, N1303);
xor XOR2 (N5438, N5420, N5384);
nor NOR3 (N5439, N5438, N5075, N4171);
nand NAND4 (N5440, N5387, N2165, N954, N3356);
not NOT1 (N5441, N5437);
not NOT1 (N5442, N5436);
or OR3 (N5443, N5441, N1892, N1540);
not NOT1 (N5444, N5439);
xor XOR2 (N5445, N5422, N5415);
nand NAND2 (N5446, N5432, N1368);
and AND2 (N5447, N5425, N914);
not NOT1 (N5448, N5445);
buf BUF1 (N5449, N5444);
buf BUF1 (N5450, N5446);
and AND4 (N5451, N5448, N4093, N468, N1245);
nor NOR4 (N5452, N5449, N2469, N979, N2584);
nand NAND3 (N5453, N5443, N4571, N1628);
nand NAND4 (N5454, N5435, N1317, N5127, N5298);
and AND3 (N5455, N5440, N3398, N5179);
not NOT1 (N5456, N5447);
or OR2 (N5457, N5442, N2369);
nand NAND3 (N5458, N5454, N685, N770);
and AND2 (N5459, N5452, N827);
or OR2 (N5460, N5457, N288);
or OR4 (N5461, N5460, N4976, N124, N2706);
nand NAND4 (N5462, N5461, N5428, N149, N3172);
nor NOR2 (N5463, N5434, N4521);
nand NAND4 (N5464, N5451, N2389, N4167, N4208);
or OR2 (N5465, N5450, N3347);
not NOT1 (N5466, N5465);
nor NOR4 (N5467, N5466, N1065, N5165, N5286);
or OR3 (N5468, N5467, N4768, N458);
buf BUF1 (N5469, N5462);
and AND2 (N5470, N5458, N3015);
nand NAND3 (N5471, N5469, N3658, N394);
and AND3 (N5472, N5459, N857, N3349);
xor XOR2 (N5473, N5470, N4903);
or OR4 (N5474, N5464, N4973, N2045, N2886);
nand NAND4 (N5475, N5456, N4903, N4804, N134);
nand NAND4 (N5476, N5472, N4566, N2018, N777);
or OR2 (N5477, N5468, N708);
and AND3 (N5478, N5471, N4872, N3743);
nor NOR4 (N5479, N5473, N4416, N2906, N3683);
xor XOR2 (N5480, N5475, N4618);
and AND4 (N5481, N5431, N4833, N1820, N4249);
nor NOR2 (N5482, N5453, N1131);
nand NAND3 (N5483, N5463, N3885, N3894);
nor NOR3 (N5484, N5483, N1151, N647);
nand NAND3 (N5485, N5481, N1476, N2656);
nor NOR2 (N5486, N5476, N856);
xor XOR2 (N5487, N5480, N962);
nor NOR2 (N5488, N5478, N5329);
and AND2 (N5489, N5487, N3796);
and AND4 (N5490, N5485, N217, N4803, N1475);
or OR4 (N5491, N5488, N5043, N1464, N5356);
and AND4 (N5492, N5486, N2656, N2817, N36);
not NOT1 (N5493, N5482);
not NOT1 (N5494, N5455);
not NOT1 (N5495, N5493);
buf BUF1 (N5496, N5495);
not NOT1 (N5497, N5490);
or OR4 (N5498, N5484, N1553, N1207, N2539);
or OR2 (N5499, N5491, N943);
not NOT1 (N5500, N5489);
nor NOR3 (N5501, N5499, N4099, N1097);
or OR3 (N5502, N5474, N4849, N4569);
or OR4 (N5503, N5477, N4978, N313, N2438);
xor XOR2 (N5504, N5494, N3770);
or OR2 (N5505, N5500, N2348);
and AND4 (N5506, N5492, N2416, N1076, N2408);
nand NAND3 (N5507, N5479, N3971, N2364);
or OR2 (N5508, N5496, N1556);
not NOT1 (N5509, N5508);
buf BUF1 (N5510, N5503);
buf BUF1 (N5511, N5497);
and AND2 (N5512, N5507, N707);
nand NAND2 (N5513, N5505, N2157);
nor NOR2 (N5514, N5511, N3792);
nor NOR4 (N5515, N5502, N2303, N4383, N3099);
nor NOR4 (N5516, N5501, N835, N2556, N3329);
or OR3 (N5517, N5498, N2143, N1701);
buf BUF1 (N5518, N5512);
xor XOR2 (N5519, N5514, N2944);
and AND3 (N5520, N5504, N4599, N1545);
xor XOR2 (N5521, N5515, N2962);
nand NAND3 (N5522, N5521, N3365, N2635);
nor NOR2 (N5523, N5506, N4948);
nand NAND4 (N5524, N5510, N4945, N3089, N4774);
and AND4 (N5525, N5516, N497, N379, N946);
nor NOR4 (N5526, N5517, N2550, N3652, N826);
nor NOR3 (N5527, N5519, N2699, N1986);
xor XOR2 (N5528, N5509, N3831);
or OR2 (N5529, N5528, N3667);
and AND3 (N5530, N5513, N2965, N1086);
xor XOR2 (N5531, N5529, N3430);
or OR2 (N5532, N5531, N3964);
nor NOR2 (N5533, N5530, N2187);
or OR2 (N5534, N5524, N1833);
nand NAND4 (N5535, N5520, N934, N821, N2812);
not NOT1 (N5536, N5525);
nand NAND3 (N5537, N5533, N5435, N35);
buf BUF1 (N5538, N5536);
and AND4 (N5539, N5527, N3694, N1382, N178);
not NOT1 (N5540, N5534);
nand NAND4 (N5541, N5523, N5047, N4661, N2600);
xor XOR2 (N5542, N5532, N3426);
nand NAND4 (N5543, N5542, N148, N1559, N1036);
or OR2 (N5544, N5540, N1046);
nand NAND2 (N5545, N5522, N1677);
not NOT1 (N5546, N5543);
nor NOR4 (N5547, N5537, N4199, N352, N2961);
not NOT1 (N5548, N5541);
not NOT1 (N5549, N5548);
nor NOR3 (N5550, N5535, N2088, N3536);
and AND4 (N5551, N5539, N626, N737, N2557);
or OR4 (N5552, N5551, N4990, N1633, N5029);
xor XOR2 (N5553, N5538, N4083);
and AND4 (N5554, N5518, N2052, N3217, N3802);
buf BUF1 (N5555, N5553);
or OR2 (N5556, N5554, N5443);
buf BUF1 (N5557, N5549);
or OR3 (N5558, N5555, N3291, N4252);
and AND3 (N5559, N5558, N4689, N3454);
or OR3 (N5560, N5550, N4406, N2974);
not NOT1 (N5561, N5556);
nor NOR3 (N5562, N5557, N55, N1127);
buf BUF1 (N5563, N5561);
nand NAND3 (N5564, N5563, N3081, N2843);
nor NOR3 (N5565, N5559, N2143, N758);
xor XOR2 (N5566, N5526, N3055);
and AND3 (N5567, N5544, N2090, N2653);
nor NOR3 (N5568, N5567, N2897, N468);
nand NAND2 (N5569, N5547, N2636);
and AND3 (N5570, N5552, N3119, N2008);
nand NAND2 (N5571, N5565, N567);
and AND3 (N5572, N5562, N3966, N550);
not NOT1 (N5573, N5560);
not NOT1 (N5574, N5573);
nand NAND4 (N5575, N5572, N2118, N3812, N4820);
nand NAND2 (N5576, N5570, N1525);
or OR3 (N5577, N5574, N5556, N4732);
and AND2 (N5578, N5546, N5317);
nand NAND3 (N5579, N5571, N3294, N2476);
buf BUF1 (N5580, N5578);
and AND2 (N5581, N5579, N2502);
buf BUF1 (N5582, N5581);
not NOT1 (N5583, N5580);
nand NAND4 (N5584, N5569, N4403, N3637, N5389);
nand NAND4 (N5585, N5566, N3477, N4602, N2861);
nand NAND4 (N5586, N5585, N576, N2965, N1303);
xor XOR2 (N5587, N5577, N4249);
and AND4 (N5588, N5575, N3165, N4417, N1266);
and AND3 (N5589, N5587, N3858, N3128);
buf BUF1 (N5590, N5545);
not NOT1 (N5591, N5564);
nor NOR2 (N5592, N5591, N1391);
nand NAND2 (N5593, N5584, N3559);
nand NAND4 (N5594, N5568, N1312, N742, N3529);
nor NOR4 (N5595, N5589, N3741, N1115, N5040);
nor NOR2 (N5596, N5592, N5443);
or OR3 (N5597, N5586, N816, N1867);
and AND4 (N5598, N5595, N3035, N2934, N4267);
xor XOR2 (N5599, N5598, N1898);
and AND4 (N5600, N5593, N4567, N1632, N3628);
or OR3 (N5601, N5594, N5449, N3015);
not NOT1 (N5602, N5600);
nand NAND3 (N5603, N5602, N5271, N1656);
nand NAND2 (N5604, N5588, N3089);
xor XOR2 (N5605, N5597, N4788);
not NOT1 (N5606, N5583);
xor XOR2 (N5607, N5603, N1500);
xor XOR2 (N5608, N5596, N4457);
nand NAND4 (N5609, N5582, N4798, N3122, N1344);
and AND4 (N5610, N5608, N206, N1558, N2789);
nor NOR2 (N5611, N5576, N3224);
xor XOR2 (N5612, N5607, N162);
buf BUF1 (N5613, N5606);
nand NAND4 (N5614, N5612, N3830, N4084, N2829);
xor XOR2 (N5615, N5613, N4391);
not NOT1 (N5616, N5604);
or OR4 (N5617, N5610, N1084, N3588, N2100);
xor XOR2 (N5618, N5601, N1492);
and AND4 (N5619, N5615, N104, N5133, N4866);
nor NOR3 (N5620, N5605, N604, N592);
nor NOR2 (N5621, N5617, N1756);
and AND2 (N5622, N5614, N1564);
nand NAND2 (N5623, N5618, N659);
xor XOR2 (N5624, N5620, N5483);
nor NOR4 (N5625, N5624, N1617, N2198, N4304);
or OR2 (N5626, N5622, N2321);
not NOT1 (N5627, N5619);
and AND4 (N5628, N5626, N1876, N4642, N3658);
and AND3 (N5629, N5616, N3794, N881);
not NOT1 (N5630, N5609);
xor XOR2 (N5631, N5623, N4716);
buf BUF1 (N5632, N5621);
not NOT1 (N5633, N5630);
xor XOR2 (N5634, N5599, N2805);
nand NAND3 (N5635, N5590, N355, N3874);
not NOT1 (N5636, N5633);
not NOT1 (N5637, N5625);
buf BUF1 (N5638, N5611);
nand NAND2 (N5639, N5627, N2537);
xor XOR2 (N5640, N5637, N281);
xor XOR2 (N5641, N5635, N2706);
nand NAND3 (N5642, N5631, N5283, N5602);
nand NAND3 (N5643, N5628, N2033, N3363);
nand NAND4 (N5644, N5640, N3290, N5592, N2930);
nand NAND3 (N5645, N5639, N2929, N3262);
not NOT1 (N5646, N5636);
xor XOR2 (N5647, N5646, N4813);
xor XOR2 (N5648, N5642, N675);
xor XOR2 (N5649, N5648, N5617);
nand NAND4 (N5650, N5644, N4833, N1275, N3087);
nand NAND4 (N5651, N5645, N1980, N5245, N653);
or OR2 (N5652, N5638, N3808);
nor NOR2 (N5653, N5650, N4576);
buf BUF1 (N5654, N5641);
and AND2 (N5655, N5654, N416);
and AND2 (N5656, N5652, N2353);
or OR3 (N5657, N5651, N1852, N4400);
nor NOR2 (N5658, N5634, N4895);
or OR3 (N5659, N5653, N5175, N2213);
not NOT1 (N5660, N5658);
nor NOR3 (N5661, N5660, N1091, N1575);
and AND2 (N5662, N5647, N4343);
and AND3 (N5663, N5649, N4394, N4090);
and AND4 (N5664, N5663, N4007, N2757, N3928);
nor NOR3 (N5665, N5655, N1745, N4232);
buf BUF1 (N5666, N5643);
nor NOR2 (N5667, N5659, N4440);
and AND2 (N5668, N5665, N1355);
or OR4 (N5669, N5664, N5390, N84, N5326);
buf BUF1 (N5670, N5629);
nor NOR2 (N5671, N5669, N1379);
nor NOR2 (N5672, N5632, N3389);
xor XOR2 (N5673, N5666, N1907);
not NOT1 (N5674, N5668);
xor XOR2 (N5675, N5661, N5267);
or OR2 (N5676, N5657, N3999);
or OR4 (N5677, N5667, N1570, N464, N4541);
and AND2 (N5678, N5677, N1511);
nand NAND3 (N5679, N5675, N4825, N5015);
nor NOR3 (N5680, N5671, N5040, N2157);
xor XOR2 (N5681, N5670, N1538);
nor NOR4 (N5682, N5676, N4412, N4247, N5432);
nand NAND2 (N5683, N5656, N4045);
nand NAND4 (N5684, N5682, N3291, N1761, N5076);
and AND3 (N5685, N5662, N3523, N3048);
nor NOR2 (N5686, N5674, N4766);
not NOT1 (N5687, N5686);
nor NOR3 (N5688, N5673, N2210, N5266);
nor NOR2 (N5689, N5684, N1074);
nand NAND4 (N5690, N5687, N1957, N4800, N4640);
and AND3 (N5691, N5681, N715, N2798);
or OR2 (N5692, N5679, N3211);
not NOT1 (N5693, N5683);
buf BUF1 (N5694, N5672);
or OR2 (N5695, N5690, N2165);
and AND2 (N5696, N5678, N3859);
nand NAND2 (N5697, N5692, N3793);
nand NAND2 (N5698, N5689, N2019);
not NOT1 (N5699, N5685);
nand NAND3 (N5700, N5688, N590, N3514);
nor NOR3 (N5701, N5693, N2307, N3923);
not NOT1 (N5702, N5695);
and AND4 (N5703, N5697, N3361, N5533, N652);
not NOT1 (N5704, N5702);
xor XOR2 (N5705, N5703, N1148);
xor XOR2 (N5706, N5698, N782);
or OR3 (N5707, N5691, N5458, N5453);
not NOT1 (N5708, N5699);
nand NAND4 (N5709, N5704, N3326, N2118, N3869);
nor NOR4 (N5710, N5707, N4243, N2556, N2341);
xor XOR2 (N5711, N5700, N3928);
nor NOR2 (N5712, N5705, N2170);
and AND2 (N5713, N5706, N3811);
nand NAND2 (N5714, N5680, N5215);
xor XOR2 (N5715, N5708, N4385);
nor NOR3 (N5716, N5711, N3867, N1468);
xor XOR2 (N5717, N5712, N2632);
buf BUF1 (N5718, N5717);
xor XOR2 (N5719, N5709, N100);
not NOT1 (N5720, N5694);
not NOT1 (N5721, N5720);
or OR3 (N5722, N5715, N5134, N3454);
buf BUF1 (N5723, N5721);
or OR4 (N5724, N5696, N563, N3864, N1378);
nor NOR2 (N5725, N5713, N5500);
nand NAND2 (N5726, N5724, N2329);
xor XOR2 (N5727, N5710, N2129);
xor XOR2 (N5728, N5714, N4612);
nor NOR2 (N5729, N5723, N4241);
nand NAND3 (N5730, N5727, N2586, N4480);
and AND2 (N5731, N5725, N4048);
nor NOR2 (N5732, N5701, N518);
not NOT1 (N5733, N5729);
not NOT1 (N5734, N5722);
xor XOR2 (N5735, N5728, N3712);
buf BUF1 (N5736, N5718);
and AND4 (N5737, N5730, N5265, N4705, N851);
and AND2 (N5738, N5719, N4311);
nand NAND2 (N5739, N5735, N3601);
not NOT1 (N5740, N5733);
xor XOR2 (N5741, N5732, N506);
not NOT1 (N5742, N5738);
xor XOR2 (N5743, N5736, N558);
nand NAND2 (N5744, N5742, N1081);
or OR4 (N5745, N5716, N5700, N2130, N5440);
nor NOR2 (N5746, N5726, N3122);
nand NAND4 (N5747, N5743, N1705, N2783, N905);
nand NAND4 (N5748, N5737, N597, N3124, N2068);
buf BUF1 (N5749, N5747);
or OR3 (N5750, N5741, N3431, N2913);
xor XOR2 (N5751, N5746, N4162);
xor XOR2 (N5752, N5734, N3596);
nand NAND4 (N5753, N5751, N236, N3368, N4053);
and AND2 (N5754, N5748, N2606);
or OR3 (N5755, N5750, N4325, N1416);
xor XOR2 (N5756, N5744, N5092);
xor XOR2 (N5757, N5745, N1930);
and AND3 (N5758, N5739, N1425, N5395);
and AND3 (N5759, N5753, N3284, N1130);
or OR2 (N5760, N5749, N2049);
nand NAND2 (N5761, N5731, N4460);
xor XOR2 (N5762, N5755, N342);
buf BUF1 (N5763, N5760);
nor NOR3 (N5764, N5757, N1442, N4209);
nand NAND4 (N5765, N5754, N2254, N214, N399);
nor NOR4 (N5766, N5752, N2484, N3217, N4000);
not NOT1 (N5767, N5765);
or OR3 (N5768, N5756, N2463, N3044);
nor NOR4 (N5769, N5762, N5605, N2122, N5170);
not NOT1 (N5770, N5763);
nor NOR3 (N5771, N5767, N4828, N3794);
nor NOR4 (N5772, N5758, N2513, N3110, N4416);
not NOT1 (N5773, N5740);
xor XOR2 (N5774, N5770, N2691);
buf BUF1 (N5775, N5771);
nand NAND2 (N5776, N5774, N2961);
not NOT1 (N5777, N5769);
and AND2 (N5778, N5768, N3486);
xor XOR2 (N5779, N5759, N1268);
xor XOR2 (N5780, N5773, N4699);
nand NAND3 (N5781, N5776, N3376, N4081);
xor XOR2 (N5782, N5764, N1433);
nor NOR4 (N5783, N5761, N455, N2156, N2148);
and AND2 (N5784, N5777, N3937);
nand NAND4 (N5785, N5775, N697, N5199, N4838);
xor XOR2 (N5786, N5780, N3870);
xor XOR2 (N5787, N5766, N5529);
or OR3 (N5788, N5783, N4756, N3895);
or OR3 (N5789, N5782, N4510, N2341);
not NOT1 (N5790, N5785);
and AND2 (N5791, N5786, N464);
buf BUF1 (N5792, N5787);
nor NOR3 (N5793, N5778, N1214, N751);
nor NOR4 (N5794, N5788, N3958, N5431, N289);
not NOT1 (N5795, N5793);
nor NOR2 (N5796, N5791, N1903);
or OR4 (N5797, N5790, N3658, N2939, N2039);
buf BUF1 (N5798, N5781);
xor XOR2 (N5799, N5779, N2609);
or OR3 (N5800, N5792, N3827, N4394);
nand NAND2 (N5801, N5795, N2495);
xor XOR2 (N5802, N5796, N3441);
buf BUF1 (N5803, N5799);
and AND4 (N5804, N5802, N843, N4601, N4881);
xor XOR2 (N5805, N5772, N801);
nand NAND4 (N5806, N5804, N5243, N1709, N1148);
nor NOR3 (N5807, N5801, N1437, N4470);
nor NOR4 (N5808, N5803, N5584, N3416, N3975);
not NOT1 (N5809, N5805);
and AND4 (N5810, N5808, N4341, N5433, N5744);
buf BUF1 (N5811, N5797);
not NOT1 (N5812, N5789);
not NOT1 (N5813, N5800);
xor XOR2 (N5814, N5794, N1340);
buf BUF1 (N5815, N5784);
xor XOR2 (N5816, N5807, N5278);
xor XOR2 (N5817, N5806, N2762);
or OR2 (N5818, N5813, N5756);
and AND2 (N5819, N5809, N1258);
xor XOR2 (N5820, N5798, N3435);
xor XOR2 (N5821, N5814, N5261);
and AND3 (N5822, N5816, N2139, N3923);
and AND4 (N5823, N5821, N64, N3790, N3779);
nand NAND2 (N5824, N5819, N4764);
buf BUF1 (N5825, N5818);
nor NOR3 (N5826, N5817, N2415, N1174);
or OR3 (N5827, N5826, N1583, N4562);
nor NOR2 (N5828, N5823, N5394);
nand NAND2 (N5829, N5827, N787);
and AND3 (N5830, N5822, N1388, N3063);
buf BUF1 (N5831, N5830);
nand NAND2 (N5832, N5810, N897);
or OR3 (N5833, N5832, N95, N2437);
and AND3 (N5834, N5824, N1663, N4205);
buf BUF1 (N5835, N5829);
nand NAND2 (N5836, N5811, N4020);
nor NOR3 (N5837, N5835, N4434, N5085);
not NOT1 (N5838, N5836);
buf BUF1 (N5839, N5815);
xor XOR2 (N5840, N5837, N2269);
nor NOR4 (N5841, N5840, N2035, N3947, N602);
nor NOR3 (N5842, N5820, N2859, N427);
nand NAND3 (N5843, N5842, N4725, N1626);
nor NOR3 (N5844, N5839, N5662, N1773);
xor XOR2 (N5845, N5828, N1654);
and AND4 (N5846, N5843, N4233, N5375, N3691);
and AND2 (N5847, N5841, N2174);
nand NAND3 (N5848, N5844, N1560, N5805);
and AND2 (N5849, N5831, N3225);
xor XOR2 (N5850, N5848, N2286);
nor NOR4 (N5851, N5838, N4799, N5718, N4908);
or OR2 (N5852, N5833, N2860);
nor NOR2 (N5853, N5852, N1588);
buf BUF1 (N5854, N5845);
or OR3 (N5855, N5846, N3539, N1136);
or OR3 (N5856, N5812, N2200, N757);
nor NOR3 (N5857, N5855, N2480, N1183);
xor XOR2 (N5858, N5854, N3680);
not NOT1 (N5859, N5853);
and AND3 (N5860, N5825, N3748, N2518);
xor XOR2 (N5861, N5858, N3522);
xor XOR2 (N5862, N5834, N909);
and AND2 (N5863, N5851, N2325);
or OR4 (N5864, N5857, N1792, N5104, N5122);
and AND3 (N5865, N5860, N2304, N5730);
not NOT1 (N5866, N5863);
nor NOR2 (N5867, N5850, N3549);
xor XOR2 (N5868, N5865, N2778);
nand NAND3 (N5869, N5856, N2733, N2895);
buf BUF1 (N5870, N5869);
nor NOR2 (N5871, N5870, N2753);
and AND3 (N5872, N5867, N1481, N1489);
buf BUF1 (N5873, N5849);
nand NAND2 (N5874, N5868, N5772);
or OR4 (N5875, N5874, N2105, N3046, N585);
nand NAND4 (N5876, N5875, N3532, N4359, N286);
nor NOR3 (N5877, N5861, N2565, N2082);
and AND3 (N5878, N5866, N1296, N4284);
or OR3 (N5879, N5877, N5248, N245);
or OR3 (N5880, N5871, N2558, N3668);
not NOT1 (N5881, N5862);
buf BUF1 (N5882, N5876);
xor XOR2 (N5883, N5872, N3701);
and AND3 (N5884, N5882, N3758, N671);
not NOT1 (N5885, N5878);
and AND2 (N5886, N5879, N595);
buf BUF1 (N5887, N5880);
xor XOR2 (N5888, N5859, N5687);
nor NOR3 (N5889, N5886, N4301, N1482);
buf BUF1 (N5890, N5889);
nor NOR3 (N5891, N5884, N4587, N4759);
not NOT1 (N5892, N5883);
buf BUF1 (N5893, N5847);
or OR3 (N5894, N5891, N2060, N5229);
not NOT1 (N5895, N5873);
or OR4 (N5896, N5885, N5352, N4387, N5255);
nand NAND2 (N5897, N5896, N4535);
and AND4 (N5898, N5897, N265, N2122, N345);
buf BUF1 (N5899, N5892);
and AND2 (N5900, N5887, N32);
not NOT1 (N5901, N5890);
xor XOR2 (N5902, N5898, N125);
buf BUF1 (N5903, N5895);
nor NOR4 (N5904, N5881, N2182, N1315, N1991);
xor XOR2 (N5905, N5864, N5473);
nand NAND2 (N5906, N5900, N918);
buf BUF1 (N5907, N5888);
nor NOR4 (N5908, N5893, N5384, N3845, N2610);
and AND3 (N5909, N5907, N4802, N4309);
and AND4 (N5910, N5906, N5162, N315, N5253);
xor XOR2 (N5911, N5899, N1471);
and AND3 (N5912, N5902, N3987, N1457);
and AND2 (N5913, N5908, N1247);
nand NAND4 (N5914, N5894, N2879, N2523, N331);
xor XOR2 (N5915, N5911, N4440);
and AND3 (N5916, N5901, N5005, N4521);
not NOT1 (N5917, N5912);
and AND4 (N5918, N5917, N1323, N2152, N2442);
nand NAND3 (N5919, N5909, N2676, N2251);
xor XOR2 (N5920, N5904, N2216);
xor XOR2 (N5921, N5916, N2701);
nor NOR4 (N5922, N5903, N4259, N2385, N1831);
nor NOR4 (N5923, N5905, N821, N3953, N4361);
buf BUF1 (N5924, N5914);
xor XOR2 (N5925, N5924, N5053);
or OR4 (N5926, N5920, N2305, N1332, N228);
or OR2 (N5927, N5921, N4628);
buf BUF1 (N5928, N5918);
or OR3 (N5929, N5919, N427, N4);
nand NAND3 (N5930, N5927, N2085, N2145);
nand NAND3 (N5931, N5926, N3188, N5096);
and AND4 (N5932, N5931, N4215, N5277, N3705);
nor NOR4 (N5933, N5913, N47, N712, N818);
or OR2 (N5934, N5910, N4757);
or OR3 (N5935, N5929, N3891, N3293);
buf BUF1 (N5936, N5930);
xor XOR2 (N5937, N5923, N5846);
xor XOR2 (N5938, N5925, N5900);
xor XOR2 (N5939, N5915, N1675);
nand NAND2 (N5940, N5938, N3506);
or OR4 (N5941, N5940, N3113, N175, N4072);
not NOT1 (N5942, N5936);
buf BUF1 (N5943, N5934);
xor XOR2 (N5944, N5935, N4338);
xor XOR2 (N5945, N5922, N4401);
nand NAND2 (N5946, N5932, N5152);
nor NOR2 (N5947, N5937, N84);
nand NAND2 (N5948, N5945, N611);
nand NAND3 (N5949, N5933, N2792, N2197);
xor XOR2 (N5950, N5944, N285);
nor NOR3 (N5951, N5943, N4931, N3098);
not NOT1 (N5952, N5946);
not NOT1 (N5953, N5942);
nand NAND2 (N5954, N5950, N4191);
xor XOR2 (N5955, N5928, N502);
nor NOR4 (N5956, N5941, N2486, N5561, N5603);
nand NAND3 (N5957, N5949, N5568, N5387);
not NOT1 (N5958, N5956);
or OR4 (N5959, N5939, N2851, N5543, N3767);
xor XOR2 (N5960, N5953, N2629);
nand NAND2 (N5961, N5954, N3680);
and AND2 (N5962, N5960, N3186);
nor NOR4 (N5963, N5959, N3168, N5059, N2898);
nor NOR4 (N5964, N5962, N3703, N132, N1159);
nor NOR4 (N5965, N5948, N4190, N4032, N2374);
nand NAND2 (N5966, N5947, N5541);
xor XOR2 (N5967, N5952, N538);
or OR4 (N5968, N5951, N5214, N320, N1427);
buf BUF1 (N5969, N5964);
and AND3 (N5970, N5955, N3132, N815);
not NOT1 (N5971, N5963);
xor XOR2 (N5972, N5961, N3141);
or OR3 (N5973, N5971, N734, N3313);
buf BUF1 (N5974, N5966);
nor NOR3 (N5975, N5967, N1724, N2439);
buf BUF1 (N5976, N5968);
and AND2 (N5977, N5972, N632);
nand NAND4 (N5978, N5975, N5586, N2481, N3629);
and AND3 (N5979, N5965, N3605, N3281);
xor XOR2 (N5980, N5970, N718);
nand NAND4 (N5981, N5980, N2874, N5427, N4756);
not NOT1 (N5982, N5969);
nand NAND2 (N5983, N5981, N1405);
not NOT1 (N5984, N5982);
buf BUF1 (N5985, N5958);
nor NOR2 (N5986, N5957, N616);
xor XOR2 (N5987, N5983, N975);
xor XOR2 (N5988, N5976, N5435);
or OR4 (N5989, N5974, N2925, N5419, N4016);
nand NAND2 (N5990, N5989, N1781);
nand NAND3 (N5991, N5988, N1417, N5500);
nand NAND3 (N5992, N5991, N1528, N3549);
and AND4 (N5993, N5979, N5429, N1490, N1272);
nand NAND2 (N5994, N5990, N926);
and AND2 (N5995, N5978, N2978);
or OR2 (N5996, N5984, N4079);
xor XOR2 (N5997, N5987, N5296);
nor NOR4 (N5998, N5985, N3295, N4960, N396);
not NOT1 (N5999, N5986);
not NOT1 (N6000, N5996);
not NOT1 (N6001, N5997);
nor NOR3 (N6002, N5998, N1160, N3394);
not NOT1 (N6003, N5973);
nor NOR2 (N6004, N6003, N2744);
nand NAND4 (N6005, N5992, N5387, N5514, N4237);
nand NAND2 (N6006, N6000, N2178);
or OR3 (N6007, N6006, N3849, N3599);
xor XOR2 (N6008, N5993, N5953);
and AND4 (N6009, N6007, N5339, N3419, N3615);
or OR3 (N6010, N6002, N23, N670);
or OR3 (N6011, N6001, N3208, N1409);
nand NAND2 (N6012, N6005, N1575);
and AND2 (N6013, N6008, N3098);
nand NAND4 (N6014, N5977, N4852, N3907, N5383);
buf BUF1 (N6015, N6012);
not NOT1 (N6016, N6014);
nor NOR4 (N6017, N6010, N562, N3200, N2380);
nand NAND2 (N6018, N6015, N985);
xor XOR2 (N6019, N6018, N3297);
nor NOR4 (N6020, N5994, N1151, N3176, N5821);
nand NAND3 (N6021, N6013, N2960, N140);
not NOT1 (N6022, N6017);
or OR2 (N6023, N6011, N1579);
not NOT1 (N6024, N6019);
nand NAND4 (N6025, N6016, N1246, N5478, N3477);
xor XOR2 (N6026, N5999, N2050);
nand NAND4 (N6027, N6020, N585, N1591, N2108);
not NOT1 (N6028, N6022);
and AND2 (N6029, N5995, N5442);
buf BUF1 (N6030, N6029);
or OR2 (N6031, N6009, N2229);
nor NOR4 (N6032, N6024, N4483, N3103, N1658);
not NOT1 (N6033, N6032);
not NOT1 (N6034, N6026);
xor XOR2 (N6035, N6004, N3621);
buf BUF1 (N6036, N6023);
and AND4 (N6037, N6033, N2686, N3271, N1384);
buf BUF1 (N6038, N6027);
nand NAND2 (N6039, N6031, N4956);
or OR3 (N6040, N6037, N5790, N5391);
buf BUF1 (N6041, N6036);
nand NAND2 (N6042, N6041, N3997);
not NOT1 (N6043, N6039);
or OR4 (N6044, N6025, N5487, N4315, N4561);
nand NAND3 (N6045, N6043, N4333, N2733);
or OR3 (N6046, N6040, N3360, N1429);
nand NAND4 (N6047, N6038, N3546, N1266, N4365);
xor XOR2 (N6048, N6045, N3833);
not NOT1 (N6049, N6034);
or OR4 (N6050, N6048, N5268, N5888, N360);
buf BUF1 (N6051, N6047);
not NOT1 (N6052, N6046);
or OR3 (N6053, N6052, N2025, N1436);
nand NAND4 (N6054, N6035, N942, N5279, N1050);
xor XOR2 (N6055, N6054, N1755);
or OR3 (N6056, N6051, N506, N5968);
or OR4 (N6057, N6050, N2954, N1875, N2872);
and AND2 (N6058, N6042, N1147);
nand NAND3 (N6059, N6049, N4450, N1644);
xor XOR2 (N6060, N6057, N3089);
not NOT1 (N6061, N6021);
nand NAND2 (N6062, N6044, N1586);
xor XOR2 (N6063, N6055, N3802);
nand NAND4 (N6064, N6028, N4776, N4389, N2312);
nor NOR2 (N6065, N6060, N1538);
xor XOR2 (N6066, N6030, N5044);
buf BUF1 (N6067, N6063);
xor XOR2 (N6068, N6056, N1025);
xor XOR2 (N6069, N6065, N2488);
or OR4 (N6070, N6061, N4429, N1011, N4188);
buf BUF1 (N6071, N6068);
nand NAND3 (N6072, N6067, N3646, N5745);
nand NAND3 (N6073, N6072, N862, N3734);
or OR2 (N6074, N6058, N5088);
xor XOR2 (N6075, N6064, N5901);
or OR2 (N6076, N6074, N4190);
and AND4 (N6077, N6069, N5920, N2391, N513);
buf BUF1 (N6078, N6076);
buf BUF1 (N6079, N6075);
nor NOR4 (N6080, N6059, N3483, N631, N1996);
buf BUF1 (N6081, N6077);
xor XOR2 (N6082, N6081, N3837);
nor NOR2 (N6083, N6066, N1535);
nor NOR3 (N6084, N6080, N5230, N3401);
not NOT1 (N6085, N6073);
and AND4 (N6086, N6071, N3529, N6075, N4269);
or OR3 (N6087, N6062, N4896, N5915);
buf BUF1 (N6088, N6082);
nor NOR4 (N6089, N6079, N1879, N4182, N5508);
nor NOR2 (N6090, N6085, N5992);
and AND4 (N6091, N6087, N6053, N5547, N1286);
nor NOR3 (N6092, N4165, N6033, N63);
buf BUF1 (N6093, N6092);
not NOT1 (N6094, N6090);
or OR2 (N6095, N6070, N5183);
not NOT1 (N6096, N6083);
not NOT1 (N6097, N6088);
buf BUF1 (N6098, N6096);
buf BUF1 (N6099, N6089);
and AND3 (N6100, N6078, N483, N1203);
nand NAND4 (N6101, N6097, N4665, N4927, N37);
buf BUF1 (N6102, N6095);
xor XOR2 (N6103, N6101, N4670);
and AND4 (N6104, N6084, N678, N1940, N2473);
nor NOR3 (N6105, N6104, N4114, N3553);
and AND2 (N6106, N6094, N5807);
nor NOR2 (N6107, N6086, N5757);
nor NOR4 (N6108, N6107, N198, N4127, N4324);
nor NOR2 (N6109, N6103, N5316);
xor XOR2 (N6110, N6109, N3726);
and AND2 (N6111, N6099, N2876);
or OR4 (N6112, N6108, N5644, N5732, N3250);
and AND4 (N6113, N6110, N3006, N5329, N4992);
buf BUF1 (N6114, N6091);
not NOT1 (N6115, N6112);
and AND2 (N6116, N6105, N1726);
and AND3 (N6117, N6113, N4083, N388);
not NOT1 (N6118, N6093);
nor NOR3 (N6119, N6116, N2892, N3380);
nor NOR3 (N6120, N6102, N4037, N1473);
buf BUF1 (N6121, N6114);
xor XOR2 (N6122, N6115, N965);
xor XOR2 (N6123, N6121, N5113);
and AND2 (N6124, N6106, N2168);
and AND3 (N6125, N6124, N1150, N3204);
and AND3 (N6126, N6119, N5693, N6091);
nor NOR3 (N6127, N6125, N3307, N3365);
and AND4 (N6128, N6126, N5863, N4836, N1843);
xor XOR2 (N6129, N6118, N1851);
xor XOR2 (N6130, N6127, N4424);
nand NAND4 (N6131, N6129, N46, N5188, N5725);
nor NOR3 (N6132, N6111, N430, N3077);
xor XOR2 (N6133, N6130, N1655);
or OR3 (N6134, N6131, N2438, N1689);
not NOT1 (N6135, N6120);
buf BUF1 (N6136, N6133);
nor NOR4 (N6137, N6132, N1122, N1487, N4595);
nor NOR3 (N6138, N6098, N4144, N491);
nor NOR2 (N6139, N6137, N4708);
nand NAND2 (N6140, N6128, N1349);
nand NAND3 (N6141, N6123, N4795, N515);
nor NOR4 (N6142, N6135, N3018, N4550, N179);
nor NOR2 (N6143, N6138, N5969);
xor XOR2 (N6144, N6140, N1235);
or OR3 (N6145, N6139, N5691, N4819);
nand NAND3 (N6146, N6136, N126, N3656);
or OR4 (N6147, N6134, N4909, N2449, N2106);
nor NOR4 (N6148, N6142, N4425, N3687, N5457);
nor NOR2 (N6149, N6148, N4696);
and AND3 (N6150, N6100, N3629, N4508);
nand NAND3 (N6151, N6150, N1587, N552);
not NOT1 (N6152, N6145);
nor NOR4 (N6153, N6143, N4549, N6007, N3084);
or OR3 (N6154, N6149, N609, N2355);
not NOT1 (N6155, N6147);
not NOT1 (N6156, N6144);
nor NOR4 (N6157, N6153, N4158, N1795, N1516);
buf BUF1 (N6158, N6122);
xor XOR2 (N6159, N6158, N1694);
buf BUF1 (N6160, N6141);
nand NAND3 (N6161, N6152, N503, N2485);
xor XOR2 (N6162, N6154, N216);
or OR2 (N6163, N6156, N5386);
nand NAND4 (N6164, N6155, N6119, N4736, N3020);
and AND2 (N6165, N6146, N1083);
and AND2 (N6166, N6160, N1125);
nand NAND2 (N6167, N6151, N3434);
xor XOR2 (N6168, N6159, N2992);
buf BUF1 (N6169, N6117);
xor XOR2 (N6170, N6165, N4435);
or OR3 (N6171, N6167, N3185, N2820);
nor NOR3 (N6172, N6166, N1443, N139);
xor XOR2 (N6173, N6168, N5417);
buf BUF1 (N6174, N6171);
or OR4 (N6175, N6174, N3641, N4206, N3565);
xor XOR2 (N6176, N6173, N2446);
xor XOR2 (N6177, N6175, N4447);
buf BUF1 (N6178, N6172);
nand NAND3 (N6179, N6170, N4406, N5393);
xor XOR2 (N6180, N6169, N3476);
nor NOR3 (N6181, N6176, N1394, N924);
xor XOR2 (N6182, N6162, N5693);
and AND3 (N6183, N6157, N4020, N4476);
xor XOR2 (N6184, N6178, N4004);
and AND2 (N6185, N6177, N6057);
or OR4 (N6186, N6163, N4452, N5789, N4429);
nor NOR4 (N6187, N6182, N5317, N748, N3297);
or OR3 (N6188, N6181, N748, N5492);
not NOT1 (N6189, N6180);
nor NOR2 (N6190, N6186, N3101);
buf BUF1 (N6191, N6190);
not NOT1 (N6192, N6164);
or OR4 (N6193, N6161, N5849, N1637, N277);
buf BUF1 (N6194, N6187);
xor XOR2 (N6195, N6189, N1875);
buf BUF1 (N6196, N6194);
or OR4 (N6197, N6179, N5687, N4150, N5919);
xor XOR2 (N6198, N6183, N3565);
or OR2 (N6199, N6193, N1848);
not NOT1 (N6200, N6196);
nor NOR4 (N6201, N6184, N730, N3522, N4261);
nand NAND3 (N6202, N6188, N3660, N5623);
nand NAND4 (N6203, N6191, N5808, N5237, N183);
or OR2 (N6204, N6201, N777);
or OR4 (N6205, N6197, N4450, N3224, N313);
nor NOR3 (N6206, N6199, N2036, N1084);
and AND3 (N6207, N6203, N5468, N3184);
or OR3 (N6208, N6195, N983, N4408);
not NOT1 (N6209, N6206);
not NOT1 (N6210, N6204);
xor XOR2 (N6211, N6198, N6020);
nor NOR4 (N6212, N6192, N3679, N1454, N5606);
and AND4 (N6213, N6208, N4512, N2620, N5739);
buf BUF1 (N6214, N6200);
nand NAND2 (N6215, N6214, N1547);
or OR4 (N6216, N6215, N2670, N711, N1682);
xor XOR2 (N6217, N6209, N1742);
buf BUF1 (N6218, N6217);
buf BUF1 (N6219, N6185);
or OR3 (N6220, N6212, N950, N3830);
nor NOR2 (N6221, N6205, N1492);
not NOT1 (N6222, N6221);
not NOT1 (N6223, N6220);
and AND4 (N6224, N6211, N3469, N499, N2694);
nor NOR2 (N6225, N6224, N1931);
and AND2 (N6226, N6218, N1953);
or OR2 (N6227, N6213, N3174);
nand NAND2 (N6228, N6227, N1088);
nand NAND4 (N6229, N6202, N4293, N4923, N4468);
xor XOR2 (N6230, N6210, N2115);
nand NAND2 (N6231, N6229, N2894);
nor NOR4 (N6232, N6222, N395, N5056, N2420);
buf BUF1 (N6233, N6230);
not NOT1 (N6234, N6207);
or OR2 (N6235, N6225, N1217);
or OR2 (N6236, N6223, N5282);
or OR2 (N6237, N6216, N3409);
buf BUF1 (N6238, N6235);
nand NAND2 (N6239, N6238, N1396);
xor XOR2 (N6240, N6233, N3838);
not NOT1 (N6241, N6231);
not NOT1 (N6242, N6219);
or OR2 (N6243, N6236, N4017);
xor XOR2 (N6244, N6237, N4896);
and AND3 (N6245, N6228, N148, N1035);
nor NOR2 (N6246, N6241, N5865);
and AND4 (N6247, N6242, N2996, N4904, N4167);
nor NOR3 (N6248, N6246, N3055, N1812);
nand NAND3 (N6249, N6244, N3181, N742);
nand NAND2 (N6250, N6234, N660);
nor NOR4 (N6251, N6243, N164, N514, N1757);
nor NOR4 (N6252, N6226, N151, N765, N1902);
not NOT1 (N6253, N6249);
nand NAND3 (N6254, N6239, N432, N5879);
not NOT1 (N6255, N6254);
nand NAND3 (N6256, N6252, N935, N4567);
and AND4 (N6257, N6232, N2458, N5343, N3923);
xor XOR2 (N6258, N6240, N6144);
or OR2 (N6259, N6248, N4786);
xor XOR2 (N6260, N6245, N2595);
xor XOR2 (N6261, N6260, N531);
and AND3 (N6262, N6258, N3715, N507);
xor XOR2 (N6263, N6256, N2602);
nand NAND2 (N6264, N6250, N1666);
buf BUF1 (N6265, N6255);
xor XOR2 (N6266, N6257, N2313);
nand NAND2 (N6267, N6253, N4330);
buf BUF1 (N6268, N6265);
nand NAND4 (N6269, N6247, N5684, N4401, N4758);
xor XOR2 (N6270, N6269, N776);
xor XOR2 (N6271, N6259, N4616);
or OR2 (N6272, N6271, N1394);
nand NAND2 (N6273, N6270, N533);
nor NOR2 (N6274, N6273, N5859);
or OR2 (N6275, N6251, N344);
xor XOR2 (N6276, N6261, N4143);
not NOT1 (N6277, N6262);
nand NAND3 (N6278, N6276, N6048, N2061);
nand NAND2 (N6279, N6277, N2179);
nand NAND4 (N6280, N6278, N2744, N4117, N2996);
xor XOR2 (N6281, N6274, N6144);
and AND3 (N6282, N6272, N5291, N6115);
and AND4 (N6283, N6281, N338, N418, N1552);
xor XOR2 (N6284, N6279, N5213);
xor XOR2 (N6285, N6267, N4469);
or OR4 (N6286, N6266, N2003, N5986, N4458);
not NOT1 (N6287, N6280);
buf BUF1 (N6288, N6287);
not NOT1 (N6289, N6284);
or OR3 (N6290, N6263, N5654, N5290);
nand NAND2 (N6291, N6285, N80);
nor NOR2 (N6292, N6291, N308);
and AND3 (N6293, N6282, N4579, N2208);
or OR4 (N6294, N6289, N1153, N2825, N676);
not NOT1 (N6295, N6293);
nor NOR4 (N6296, N6288, N3704, N3284, N4008);
nor NOR3 (N6297, N6295, N4351, N2604);
and AND4 (N6298, N6296, N3221, N2497, N2877);
not NOT1 (N6299, N6275);
nand NAND4 (N6300, N6286, N2263, N332, N4430);
buf BUF1 (N6301, N6283);
nand NAND4 (N6302, N6300, N488, N2835, N423);
not NOT1 (N6303, N6301);
nand NAND4 (N6304, N6297, N924, N1409, N4834);
nand NAND3 (N6305, N6303, N103, N1552);
xor XOR2 (N6306, N6304, N4608);
or OR4 (N6307, N6268, N4890, N1161, N4082);
nand NAND3 (N6308, N6302, N2317, N5838);
nand NAND2 (N6309, N6264, N4069);
or OR4 (N6310, N6309, N1303, N146, N3613);
nor NOR2 (N6311, N6305, N3753);
xor XOR2 (N6312, N6299, N3047);
xor XOR2 (N6313, N6306, N2825);
and AND2 (N6314, N6312, N329);
buf BUF1 (N6315, N6310);
buf BUF1 (N6316, N6313);
buf BUF1 (N6317, N6311);
and AND2 (N6318, N6294, N3439);
nor NOR3 (N6319, N6308, N1043, N4260);
not NOT1 (N6320, N6298);
nand NAND4 (N6321, N6317, N2484, N6147, N2237);
xor XOR2 (N6322, N6315, N2988);
buf BUF1 (N6323, N6318);
or OR2 (N6324, N6320, N2094);
not NOT1 (N6325, N6290);
buf BUF1 (N6326, N6319);
xor XOR2 (N6327, N6323, N5764);
not NOT1 (N6328, N6324);
and AND2 (N6329, N6314, N707);
nor NOR3 (N6330, N6321, N5757, N2207);
not NOT1 (N6331, N6327);
buf BUF1 (N6332, N6307);
buf BUF1 (N6333, N6329);
and AND2 (N6334, N6328, N2874);
and AND4 (N6335, N6331, N2456, N4647, N4189);
or OR4 (N6336, N6333, N1567, N5089, N53);
nor NOR4 (N6337, N6336, N3771, N34, N2980);
not NOT1 (N6338, N6330);
nand NAND3 (N6339, N6322, N5025, N3460);
and AND2 (N6340, N6338, N3983);
not NOT1 (N6341, N6337);
not NOT1 (N6342, N6292);
not NOT1 (N6343, N6340);
xor XOR2 (N6344, N6341, N3013);
or OR4 (N6345, N6343, N6042, N625, N3183);
nor NOR2 (N6346, N6344, N3933);
not NOT1 (N6347, N6332);
xor XOR2 (N6348, N6339, N3459);
or OR2 (N6349, N6335, N2121);
nand NAND2 (N6350, N6342, N2027);
or OR3 (N6351, N6345, N808, N2908);
not NOT1 (N6352, N6325);
and AND3 (N6353, N6351, N5973, N206);
nor NOR4 (N6354, N6316, N3560, N4859, N825);
xor XOR2 (N6355, N6326, N1631);
buf BUF1 (N6356, N6348);
and AND3 (N6357, N6347, N1028, N344);
nand NAND3 (N6358, N6355, N1929, N6016);
xor XOR2 (N6359, N6334, N3551);
xor XOR2 (N6360, N6353, N6222);
or OR4 (N6361, N6350, N1712, N3362, N4626);
nor NOR3 (N6362, N6356, N5423, N5958);
nor NOR2 (N6363, N6362, N2669);
or OR3 (N6364, N6363, N3475, N6281);
buf BUF1 (N6365, N6354);
nand NAND3 (N6366, N6365, N5417, N985);
buf BUF1 (N6367, N6346);
buf BUF1 (N6368, N6352);
and AND2 (N6369, N6358, N3627);
and AND4 (N6370, N6349, N4973, N4193, N773);
and AND4 (N6371, N6359, N4037, N5032, N718);
not NOT1 (N6372, N6360);
or OR2 (N6373, N6372, N2089);
and AND2 (N6374, N6361, N2724);
xor XOR2 (N6375, N6371, N1816);
xor XOR2 (N6376, N6357, N5544);
nor NOR3 (N6377, N6367, N5585, N4863);
or OR3 (N6378, N6375, N36, N5608);
xor XOR2 (N6379, N6364, N3751);
xor XOR2 (N6380, N6368, N3080);
buf BUF1 (N6381, N6373);
and AND2 (N6382, N6376, N1897);
or OR3 (N6383, N6380, N5372, N3181);
nand NAND4 (N6384, N6378, N2460, N284, N5886);
or OR2 (N6385, N6381, N5472);
not NOT1 (N6386, N6369);
buf BUF1 (N6387, N6370);
buf BUF1 (N6388, N6385);
or OR3 (N6389, N6384, N4045, N2460);
xor XOR2 (N6390, N6387, N2423);
not NOT1 (N6391, N6379);
nand NAND4 (N6392, N6382, N76, N2544, N2660);
and AND3 (N6393, N6392, N5619, N5128);
nand NAND4 (N6394, N6374, N5382, N3079, N5399);
xor XOR2 (N6395, N6389, N4051);
nor NOR4 (N6396, N6377, N1383, N2572, N2668);
and AND4 (N6397, N6388, N6125, N6307, N5895);
nor NOR4 (N6398, N6366, N1275, N1811, N4405);
xor XOR2 (N6399, N6396, N4886);
xor XOR2 (N6400, N6399, N4746);
not NOT1 (N6401, N6390);
or OR3 (N6402, N6383, N6312, N1930);
nand NAND4 (N6403, N6402, N6083, N1778, N5019);
not NOT1 (N6404, N6397);
xor XOR2 (N6405, N6391, N2553);
or OR4 (N6406, N6395, N4994, N1526, N4019);
nor NOR4 (N6407, N6406, N4485, N1797, N1589);
nand NAND3 (N6408, N6407, N5729, N4218);
or OR4 (N6409, N6398, N2294, N5118, N3519);
buf BUF1 (N6410, N6404);
nand NAND2 (N6411, N6386, N6368);
xor XOR2 (N6412, N6401, N4577);
nand NAND4 (N6413, N6412, N4819, N4154, N4867);
nand NAND4 (N6414, N6408, N3128, N5222, N1205);
xor XOR2 (N6415, N6394, N5693);
or OR3 (N6416, N6400, N6120, N3301);
nand NAND3 (N6417, N6409, N4415, N2291);
buf BUF1 (N6418, N6403);
or OR4 (N6419, N6414, N4904, N437, N1501);
and AND3 (N6420, N6410, N3976, N1670);
not NOT1 (N6421, N6413);
or OR3 (N6422, N6393, N65, N2004);
and AND4 (N6423, N6419, N6195, N2875, N5495);
nor NOR4 (N6424, N6418, N349, N2799, N4394);
and AND3 (N6425, N6421, N2912, N1509);
or OR2 (N6426, N6411, N4176);
and AND4 (N6427, N6415, N371, N6176, N1014);
nand NAND2 (N6428, N6417, N931);
xor XOR2 (N6429, N6420, N4380);
nor NOR3 (N6430, N6427, N1835, N4794);
buf BUF1 (N6431, N6405);
and AND2 (N6432, N6429, N5254);
nor NOR4 (N6433, N6431, N5819, N317, N1818);
xor XOR2 (N6434, N6416, N3641);
and AND3 (N6435, N6423, N1457, N578);
buf BUF1 (N6436, N6428);
or OR3 (N6437, N6432, N4743, N6101);
nand NAND4 (N6438, N6435, N6279, N5189, N5452);
xor XOR2 (N6439, N6437, N1072);
not NOT1 (N6440, N6430);
nor NOR3 (N6441, N6434, N4032, N5214);
not NOT1 (N6442, N6422);
buf BUF1 (N6443, N6424);
buf BUF1 (N6444, N6441);
not NOT1 (N6445, N6426);
not NOT1 (N6446, N6440);
or OR2 (N6447, N6446, N2000);
nor NOR4 (N6448, N6439, N5602, N4061, N738);
buf BUF1 (N6449, N6445);
and AND4 (N6450, N6448, N124, N3157, N4783);
nor NOR2 (N6451, N6438, N2340);
or OR2 (N6452, N6443, N1774);
buf BUF1 (N6453, N6436);
nor NOR4 (N6454, N6449, N2109, N160, N2135);
and AND4 (N6455, N6433, N2884, N5253, N518);
nand NAND2 (N6456, N6451, N4384);
not NOT1 (N6457, N6453);
buf BUF1 (N6458, N6452);
nor NOR3 (N6459, N6444, N575, N6272);
not NOT1 (N6460, N6458);
buf BUF1 (N6461, N6447);
buf BUF1 (N6462, N6460);
not NOT1 (N6463, N6442);
nand NAND3 (N6464, N6459, N5834, N6254);
not NOT1 (N6465, N6450);
nand NAND2 (N6466, N6461, N6435);
xor XOR2 (N6467, N6456, N4737);
or OR3 (N6468, N6462, N4168, N6078);
nand NAND4 (N6469, N6464, N609, N1360, N3812);
or OR2 (N6470, N6457, N2227);
nand NAND4 (N6471, N6425, N4737, N917, N2015);
buf BUF1 (N6472, N6465);
buf BUF1 (N6473, N6471);
nor NOR4 (N6474, N6472, N4194, N4403, N6240);
not NOT1 (N6475, N6468);
or OR4 (N6476, N6474, N6054, N4189, N2290);
and AND2 (N6477, N6463, N2357);
not NOT1 (N6478, N6473);
and AND3 (N6479, N6469, N4814, N322);
or OR3 (N6480, N6475, N3247, N5267);
not NOT1 (N6481, N6454);
xor XOR2 (N6482, N6476, N5770);
buf BUF1 (N6483, N6480);
or OR4 (N6484, N6467, N6461, N3900, N1455);
and AND3 (N6485, N6483, N6416, N6464);
nand NAND2 (N6486, N6484, N3017);
buf BUF1 (N6487, N6482);
and AND3 (N6488, N6481, N6052, N2389);
xor XOR2 (N6489, N6485, N5202);
nor NOR3 (N6490, N6478, N4965, N1307);
xor XOR2 (N6491, N6455, N2210);
and AND4 (N6492, N6479, N4786, N1169, N3316);
nand NAND4 (N6493, N6492, N2090, N5617, N3972);
buf BUF1 (N6494, N6486);
xor XOR2 (N6495, N6487, N182);
nor NOR3 (N6496, N6489, N421, N2379);
or OR3 (N6497, N6491, N2246, N5258);
xor XOR2 (N6498, N6493, N6024);
not NOT1 (N6499, N6497);
nor NOR3 (N6500, N6477, N3376, N4230);
buf BUF1 (N6501, N6488);
xor XOR2 (N6502, N6495, N3275);
xor XOR2 (N6503, N6500, N4512);
buf BUF1 (N6504, N6503);
not NOT1 (N6505, N6502);
not NOT1 (N6506, N6490);
not NOT1 (N6507, N6501);
buf BUF1 (N6508, N6470);
buf BUF1 (N6509, N6504);
nor NOR3 (N6510, N6508, N5700, N1630);
buf BUF1 (N6511, N6510);
not NOT1 (N6512, N6494);
and AND2 (N6513, N6498, N4481);
xor XOR2 (N6514, N6505, N5783);
or OR3 (N6515, N6509, N1663, N4723);
and AND3 (N6516, N6512, N2963, N2035);
buf BUF1 (N6517, N6514);
not NOT1 (N6518, N6506);
not NOT1 (N6519, N6507);
and AND4 (N6520, N6516, N4596, N697, N6011);
or OR2 (N6521, N6466, N5133);
nand NAND4 (N6522, N6499, N1049, N88, N3832);
nand NAND2 (N6523, N6520, N4948);
nand NAND3 (N6524, N6521, N6512, N4262);
or OR3 (N6525, N6522, N3835, N6158);
nor NOR4 (N6526, N6517, N6126, N598, N2514);
xor XOR2 (N6527, N6496, N5463);
buf BUF1 (N6528, N6519);
nand NAND3 (N6529, N6524, N2602, N4675);
nand NAND4 (N6530, N6529, N3565, N3762, N394);
nand NAND3 (N6531, N6527, N5143, N3678);
and AND4 (N6532, N6518, N6421, N5016, N523);
not NOT1 (N6533, N6515);
nand NAND3 (N6534, N6525, N2015, N325);
buf BUF1 (N6535, N6531);
and AND4 (N6536, N6523, N3968, N6292, N1587);
nor NOR3 (N6537, N6532, N1192, N4820);
nor NOR3 (N6538, N6534, N4232, N164);
buf BUF1 (N6539, N6528);
nand NAND4 (N6540, N6526, N814, N5344, N6195);
xor XOR2 (N6541, N6539, N2328);
buf BUF1 (N6542, N6511);
or OR3 (N6543, N6536, N986, N2432);
xor XOR2 (N6544, N6543, N3585);
xor XOR2 (N6545, N6542, N3404);
or OR2 (N6546, N6530, N2414);
not NOT1 (N6547, N6544);
and AND3 (N6548, N6537, N5820, N3839);
xor XOR2 (N6549, N6513, N5371);
buf BUF1 (N6550, N6535);
and AND3 (N6551, N6547, N1931, N1525);
xor XOR2 (N6552, N6538, N2002);
nor NOR4 (N6553, N6540, N1810, N3213, N2513);
or OR3 (N6554, N6549, N2089, N1076);
nor NOR3 (N6555, N6551, N2605, N3609);
or OR2 (N6556, N6541, N4600);
and AND2 (N6557, N6546, N4231);
nand NAND3 (N6558, N6545, N1685, N2776);
buf BUF1 (N6559, N6533);
buf BUF1 (N6560, N6558);
buf BUF1 (N6561, N6554);
xor XOR2 (N6562, N6548, N3093);
nor NOR2 (N6563, N6560, N1275);
or OR2 (N6564, N6555, N5973);
nor NOR2 (N6565, N6563, N5723);
or OR2 (N6566, N6556, N6122);
not NOT1 (N6567, N6565);
xor XOR2 (N6568, N6562, N630);
nand NAND3 (N6569, N6559, N5813, N3018);
and AND2 (N6570, N6567, N5835);
or OR4 (N6571, N6550, N4641, N2657, N3357);
nor NOR2 (N6572, N6561, N1190);
nor NOR3 (N6573, N6572, N2475, N5362);
buf BUF1 (N6574, N6570);
nor NOR4 (N6575, N6574, N3032, N3842, N5116);
not NOT1 (N6576, N6566);
nor NOR4 (N6577, N6568, N6551, N5612, N5723);
or OR4 (N6578, N6557, N4377, N6219, N2308);
nor NOR3 (N6579, N6571, N3217, N74);
or OR4 (N6580, N6552, N397, N4470, N6485);
or OR3 (N6581, N6579, N3616, N6459);
nor NOR2 (N6582, N6564, N3357);
or OR3 (N6583, N6577, N2152, N4175);
xor XOR2 (N6584, N6578, N5402);
and AND2 (N6585, N6581, N3134);
and AND4 (N6586, N6575, N1529, N4672, N3279);
nor NOR3 (N6587, N6586, N4574, N1374);
and AND2 (N6588, N6576, N879);
xor XOR2 (N6589, N6580, N765);
nand NAND2 (N6590, N6585, N310);
or OR4 (N6591, N6584, N1959, N3129, N3070);
and AND3 (N6592, N6587, N3559, N4494);
buf BUF1 (N6593, N6583);
and AND4 (N6594, N6590, N5514, N3853, N2016);
or OR3 (N6595, N6573, N5732, N4046);
not NOT1 (N6596, N6595);
nor NOR3 (N6597, N6596, N6152, N3632);
xor XOR2 (N6598, N6569, N2295);
and AND3 (N6599, N6553, N3305, N3076);
buf BUF1 (N6600, N6592);
buf BUF1 (N6601, N6588);
and AND4 (N6602, N6594, N2364, N6295, N3000);
nand NAND3 (N6603, N6602, N2177, N3227);
buf BUF1 (N6604, N6593);
buf BUF1 (N6605, N6582);
not NOT1 (N6606, N6604);
and AND4 (N6607, N6606, N1505, N2267, N616);
buf BUF1 (N6608, N6598);
xor XOR2 (N6609, N6601, N1004);
buf BUF1 (N6610, N6607);
not NOT1 (N6611, N6600);
nand NAND4 (N6612, N6605, N505, N4626, N1260);
nor NOR3 (N6613, N6608, N2515, N5092);
nor NOR3 (N6614, N6597, N1558, N4779);
not NOT1 (N6615, N6611);
nor NOR2 (N6616, N6609, N430);
nand NAND2 (N6617, N6616, N1245);
not NOT1 (N6618, N6615);
nor NOR2 (N6619, N6610, N2823);
and AND3 (N6620, N6599, N1065, N110);
nor NOR2 (N6621, N6619, N3232);
xor XOR2 (N6622, N6617, N5496);
not NOT1 (N6623, N6612);
buf BUF1 (N6624, N6613);
and AND3 (N6625, N6622, N5644, N1126);
and AND2 (N6626, N6621, N4710);
buf BUF1 (N6627, N6618);
nor NOR3 (N6628, N6625, N5783, N3094);
or OR2 (N6629, N6626, N2103);
xor XOR2 (N6630, N6624, N21);
or OR4 (N6631, N6589, N6451, N648, N4854);
nor NOR2 (N6632, N6623, N1981);
nor NOR4 (N6633, N6631, N630, N2202, N5395);
buf BUF1 (N6634, N6629);
nor NOR3 (N6635, N6627, N3081, N5673);
or OR2 (N6636, N6632, N3724);
and AND2 (N6637, N6603, N3778);
buf BUF1 (N6638, N6636);
not NOT1 (N6639, N6614);
nand NAND3 (N6640, N6630, N4038, N1410);
xor XOR2 (N6641, N6591, N127);
and AND2 (N6642, N6641, N352);
nand NAND3 (N6643, N6635, N4027, N313);
xor XOR2 (N6644, N6628, N3780);
xor XOR2 (N6645, N6637, N4202);
nand NAND4 (N6646, N6633, N1713, N2304, N864);
and AND3 (N6647, N6645, N2023, N5172);
buf BUF1 (N6648, N6642);
nor NOR2 (N6649, N6638, N5137);
and AND3 (N6650, N6649, N1572, N6275);
buf BUF1 (N6651, N6648);
not NOT1 (N6652, N6647);
buf BUF1 (N6653, N6651);
nand NAND2 (N6654, N6634, N5063);
not NOT1 (N6655, N6639);
and AND2 (N6656, N6652, N3100);
xor XOR2 (N6657, N6650, N6015);
not NOT1 (N6658, N6643);
xor XOR2 (N6659, N6655, N1925);
nand NAND4 (N6660, N6620, N2538, N1807, N5679);
xor XOR2 (N6661, N6646, N552);
nand NAND3 (N6662, N6661, N3169, N5863);
not NOT1 (N6663, N6656);
nor NOR3 (N6664, N6663, N4671, N6258);
buf BUF1 (N6665, N6659);
and AND3 (N6666, N6658, N5402, N1504);
and AND2 (N6667, N6662, N2461);
buf BUF1 (N6668, N6666);
not NOT1 (N6669, N6657);
not NOT1 (N6670, N6654);
nand NAND3 (N6671, N6668, N1297, N4138);
not NOT1 (N6672, N6640);
xor XOR2 (N6673, N6670, N5536);
and AND3 (N6674, N6664, N6484, N4746);
or OR4 (N6675, N6671, N6621, N2753, N4628);
buf BUF1 (N6676, N6660);
xor XOR2 (N6677, N6672, N6363);
nor NOR2 (N6678, N6665, N3067);
not NOT1 (N6679, N6678);
and AND3 (N6680, N6676, N6619, N1630);
and AND4 (N6681, N6669, N1617, N4409, N2452);
nand NAND3 (N6682, N6673, N5613, N3934);
and AND4 (N6683, N6680, N4346, N4383, N231);
xor XOR2 (N6684, N6653, N4630);
not NOT1 (N6685, N6683);
nor NOR3 (N6686, N6667, N700, N3504);
or OR3 (N6687, N6679, N3653, N1460);
or OR2 (N6688, N6677, N1230);
nand NAND2 (N6689, N6682, N1663);
or OR2 (N6690, N6687, N5988);
or OR2 (N6691, N6684, N3990);
nand NAND3 (N6692, N6690, N1218, N456);
or OR3 (N6693, N6675, N1326, N3575);
or OR2 (N6694, N6692, N2441);
xor XOR2 (N6695, N6693, N2589);
or OR3 (N6696, N6681, N5922, N3591);
buf BUF1 (N6697, N6685);
buf BUF1 (N6698, N6697);
or OR4 (N6699, N6686, N1575, N5982, N4408);
nor NOR3 (N6700, N6695, N5112, N4849);
nand NAND2 (N6701, N6688, N2307);
buf BUF1 (N6702, N6689);
and AND4 (N6703, N6674, N64, N1467, N898);
nor NOR2 (N6704, N6703, N1648);
buf BUF1 (N6705, N6696);
nor NOR3 (N6706, N6704, N1835, N5835);
xor XOR2 (N6707, N6698, N4390);
nor NOR2 (N6708, N6701, N3362);
buf BUF1 (N6709, N6694);
and AND2 (N6710, N6644, N36);
nand NAND2 (N6711, N6706, N1639);
nor NOR4 (N6712, N6709, N2350, N3104, N170);
not NOT1 (N6713, N6702);
xor XOR2 (N6714, N6711, N4349);
or OR4 (N6715, N6710, N5062, N1777, N5497);
buf BUF1 (N6716, N6712);
not NOT1 (N6717, N6714);
not NOT1 (N6718, N6705);
buf BUF1 (N6719, N6713);
or OR3 (N6720, N6715, N2987, N4769);
not NOT1 (N6721, N6718);
buf BUF1 (N6722, N6699);
xor XOR2 (N6723, N6707, N1653);
and AND2 (N6724, N6708, N5746);
and AND4 (N6725, N6700, N3740, N5177, N4273);
and AND3 (N6726, N6716, N2445, N1521);
not NOT1 (N6727, N6717);
not NOT1 (N6728, N6724);
xor XOR2 (N6729, N6725, N6277);
or OR3 (N6730, N6691, N1194, N490);
nor NOR4 (N6731, N6726, N687, N978, N3961);
buf BUF1 (N6732, N6728);
xor XOR2 (N6733, N6727, N310);
buf BUF1 (N6734, N6730);
xor XOR2 (N6735, N6732, N1226);
nor NOR4 (N6736, N6735, N3706, N1207, N1082);
not NOT1 (N6737, N6736);
nand NAND3 (N6738, N6723, N4018, N3045);
buf BUF1 (N6739, N6733);
xor XOR2 (N6740, N6721, N1209);
nand NAND3 (N6741, N6719, N6599, N3472);
buf BUF1 (N6742, N6739);
xor XOR2 (N6743, N6738, N4215);
xor XOR2 (N6744, N6743, N5716);
nand NAND4 (N6745, N6722, N3856, N4303, N6619);
nor NOR2 (N6746, N6745, N6583);
xor XOR2 (N6747, N6741, N4314);
xor XOR2 (N6748, N6746, N3995);
xor XOR2 (N6749, N6747, N5567);
nor NOR2 (N6750, N6748, N1646);
and AND4 (N6751, N6734, N4063, N2129, N4040);
xor XOR2 (N6752, N6731, N1012);
or OR3 (N6753, N6744, N4101, N1227);
or OR3 (N6754, N6751, N6138, N6592);
nor NOR2 (N6755, N6749, N1636);
or OR3 (N6756, N6740, N812, N5410);
and AND3 (N6757, N6754, N6597, N570);
and AND4 (N6758, N6753, N564, N3163, N4957);
buf BUF1 (N6759, N6755);
or OR2 (N6760, N6720, N2408);
buf BUF1 (N6761, N6737);
nor NOR3 (N6762, N6756, N5745, N4352);
and AND4 (N6763, N6761, N6743, N6601, N3863);
not NOT1 (N6764, N6742);
not NOT1 (N6765, N6752);
nor NOR2 (N6766, N6750, N1018);
and AND2 (N6767, N6766, N3084);
or OR2 (N6768, N6767, N6571);
buf BUF1 (N6769, N6759);
or OR2 (N6770, N6764, N546);
buf BUF1 (N6771, N6758);
xor XOR2 (N6772, N6762, N1209);
nand NAND3 (N6773, N6768, N6238, N5121);
buf BUF1 (N6774, N6769);
xor XOR2 (N6775, N6774, N1787);
or OR3 (N6776, N6729, N3879, N5352);
and AND3 (N6777, N6757, N5674, N3167);
or OR2 (N6778, N6772, N6408);
nand NAND3 (N6779, N6760, N1100, N6695);
buf BUF1 (N6780, N6770);
xor XOR2 (N6781, N6771, N2470);
not NOT1 (N6782, N6781);
xor XOR2 (N6783, N6779, N5617);
nand NAND2 (N6784, N6775, N5194);
not NOT1 (N6785, N6776);
and AND2 (N6786, N6773, N6767);
nor NOR3 (N6787, N6778, N3820, N1189);
and AND3 (N6788, N6763, N2030, N480);
xor XOR2 (N6789, N6765, N2757);
and AND2 (N6790, N6789, N2227);
nor NOR4 (N6791, N6785, N6293, N1414, N3078);
nor NOR3 (N6792, N6791, N1536, N2640);
not NOT1 (N6793, N6782);
nand NAND2 (N6794, N6790, N2052);
or OR3 (N6795, N6777, N2248, N6121);
nand NAND3 (N6796, N6784, N1922, N5932);
or OR4 (N6797, N6787, N4869, N1503, N3553);
buf BUF1 (N6798, N6788);
xor XOR2 (N6799, N6795, N2018);
nor NOR3 (N6800, N6794, N6763, N5170);
xor XOR2 (N6801, N6796, N1293);
or OR3 (N6802, N6783, N3189, N3245);
buf BUF1 (N6803, N6802);
buf BUF1 (N6804, N6798);
buf BUF1 (N6805, N6800);
and AND2 (N6806, N6793, N18);
xor XOR2 (N6807, N6792, N4866);
not NOT1 (N6808, N6807);
xor XOR2 (N6809, N6805, N3564);
and AND2 (N6810, N6804, N554);
buf BUF1 (N6811, N6780);
not NOT1 (N6812, N6797);
and AND2 (N6813, N6786, N3766);
xor XOR2 (N6814, N6799, N1693);
buf BUF1 (N6815, N6814);
and AND2 (N6816, N6813, N329);
xor XOR2 (N6817, N6801, N815);
or OR2 (N6818, N6811, N4106);
nand NAND3 (N6819, N6809, N4684, N1670);
and AND3 (N6820, N6816, N1924, N1604);
xor XOR2 (N6821, N6817, N899);
nand NAND3 (N6822, N6821, N2933, N4172);
or OR2 (N6823, N6803, N5998);
and AND2 (N6824, N6822, N3203);
nand NAND3 (N6825, N6810, N5055, N5174);
nand NAND3 (N6826, N6818, N3175, N1752);
and AND3 (N6827, N6812, N85, N2170);
nor NOR4 (N6828, N6806, N2432, N690, N1091);
buf BUF1 (N6829, N6828);
nor NOR3 (N6830, N6808, N4713, N3214);
or OR3 (N6831, N6815, N2621, N168);
and AND3 (N6832, N6823, N5673, N4538);
not NOT1 (N6833, N6820);
or OR4 (N6834, N6819, N4446, N382, N1120);
xor XOR2 (N6835, N6827, N2704);
nor NOR2 (N6836, N6830, N4663);
buf BUF1 (N6837, N6825);
nand NAND4 (N6838, N6837, N2863, N6353, N5891);
buf BUF1 (N6839, N6834);
buf BUF1 (N6840, N6832);
or OR2 (N6841, N6824, N103);
nand NAND4 (N6842, N6831, N5911, N810, N1744);
nor NOR3 (N6843, N6836, N6615, N5030);
nand NAND3 (N6844, N6826, N3390, N3539);
and AND2 (N6845, N6838, N2294);
not NOT1 (N6846, N6833);
xor XOR2 (N6847, N6843, N3201);
and AND4 (N6848, N6844, N4493, N6575, N1022);
xor XOR2 (N6849, N6840, N5766);
nand NAND3 (N6850, N6842, N6143, N6015);
xor XOR2 (N6851, N6850, N6390);
or OR2 (N6852, N6846, N4732);
xor XOR2 (N6853, N6829, N6739);
nor NOR3 (N6854, N6835, N2080, N6750);
buf BUF1 (N6855, N6841);
and AND3 (N6856, N6851, N74, N5651);
nand NAND3 (N6857, N6848, N4004, N2845);
or OR3 (N6858, N6853, N1988, N5423);
xor XOR2 (N6859, N6849, N1060);
and AND2 (N6860, N6847, N276);
and AND3 (N6861, N6855, N821, N3524);
not NOT1 (N6862, N6860);
or OR3 (N6863, N6854, N5694, N121);
and AND4 (N6864, N6858, N2678, N4816, N841);
not NOT1 (N6865, N6859);
nor NOR2 (N6866, N6839, N1791);
nor NOR3 (N6867, N6857, N2932, N1851);
nor NOR3 (N6868, N6861, N908, N5959);
nand NAND2 (N6869, N6868, N3769);
buf BUF1 (N6870, N6863);
not NOT1 (N6871, N6845);
buf BUF1 (N6872, N6862);
nand NAND4 (N6873, N6867, N6393, N3195, N862);
not NOT1 (N6874, N6852);
nor NOR3 (N6875, N6873, N4687, N6500);
xor XOR2 (N6876, N6875, N5149);
xor XOR2 (N6877, N6876, N6359);
nand NAND3 (N6878, N6872, N5276, N6549);
nor NOR2 (N6879, N6866, N3522);
buf BUF1 (N6880, N6870);
nand NAND3 (N6881, N6880, N3613, N1613);
and AND2 (N6882, N6869, N4931);
or OR2 (N6883, N6856, N4423);
not NOT1 (N6884, N6883);
not NOT1 (N6885, N6881);
nor NOR3 (N6886, N6877, N1694, N4491);
xor XOR2 (N6887, N6882, N3303);
and AND3 (N6888, N6864, N2358, N6475);
buf BUF1 (N6889, N6888);
nand NAND4 (N6890, N6879, N6066, N1228, N489);
nor NOR3 (N6891, N6874, N6836, N3583);
xor XOR2 (N6892, N6884, N6239);
or OR2 (N6893, N6887, N2946);
not NOT1 (N6894, N6889);
not NOT1 (N6895, N6892);
nand NAND2 (N6896, N6890, N4057);
nor NOR3 (N6897, N6878, N1428, N2038);
nand NAND4 (N6898, N6896, N2319, N2626, N2285);
or OR2 (N6899, N6895, N5981);
xor XOR2 (N6900, N6893, N4103);
buf BUF1 (N6901, N6894);
buf BUF1 (N6902, N6899);
or OR2 (N6903, N6865, N2656);
or OR4 (N6904, N6902, N4143, N3593, N1649);
or OR4 (N6905, N6900, N1650, N5708, N4791);
and AND4 (N6906, N6905, N4126, N2062, N1513);
xor XOR2 (N6907, N6871, N4457);
nor NOR3 (N6908, N6891, N5805, N5849);
and AND4 (N6909, N6904, N594, N2028, N1990);
buf BUF1 (N6910, N6907);
not NOT1 (N6911, N6886);
nand NAND4 (N6912, N6909, N91, N5915, N5606);
buf BUF1 (N6913, N6898);
and AND2 (N6914, N6910, N4937);
not NOT1 (N6915, N6885);
nor NOR3 (N6916, N6906, N3333, N6207);
nand NAND2 (N6917, N6914, N5762);
nand NAND2 (N6918, N6901, N3914);
not NOT1 (N6919, N6916);
not NOT1 (N6920, N6912);
nand NAND4 (N6921, N6920, N1372, N3688, N4288);
buf BUF1 (N6922, N6921);
xor XOR2 (N6923, N6917, N4601);
nand NAND3 (N6924, N6911, N5045, N2442);
or OR2 (N6925, N6908, N5107);
nor NOR4 (N6926, N6913, N6171, N3004, N2705);
or OR2 (N6927, N6926, N3356);
and AND2 (N6928, N6919, N5413);
xor XOR2 (N6929, N6897, N388);
not NOT1 (N6930, N6924);
not NOT1 (N6931, N6903);
nand NAND4 (N6932, N6925, N400, N6684, N3715);
nor NOR3 (N6933, N6930, N3900, N167);
and AND4 (N6934, N6928, N3192, N5797, N6379);
nand NAND3 (N6935, N6923, N1972, N5858);
nand NAND3 (N6936, N6922, N5188, N6220);
and AND2 (N6937, N6929, N5607);
or OR4 (N6938, N6935, N6880, N1291, N3469);
nor NOR2 (N6939, N6915, N4381);
nand NAND2 (N6940, N6918, N4109);
buf BUF1 (N6941, N6927);
nand NAND2 (N6942, N6937, N6451);
xor XOR2 (N6943, N6939, N1961);
and AND4 (N6944, N6936, N5281, N4925, N6039);
nand NAND4 (N6945, N6942, N1326, N3722, N6258);
and AND3 (N6946, N6934, N5294, N1881);
and AND3 (N6947, N6931, N3059, N192);
or OR2 (N6948, N6933, N1448);
nand NAND3 (N6949, N6941, N5427, N53);
not NOT1 (N6950, N6943);
nand NAND4 (N6951, N6950, N1467, N6668, N3317);
and AND4 (N6952, N6944, N2538, N3877, N3225);
xor XOR2 (N6953, N6932, N2317);
or OR4 (N6954, N6951, N6232, N5595, N6887);
xor XOR2 (N6955, N6947, N6888);
nand NAND2 (N6956, N6954, N5186);
or OR2 (N6957, N6949, N4887);
not NOT1 (N6958, N6955);
not NOT1 (N6959, N6956);
xor XOR2 (N6960, N6946, N5143);
nor NOR2 (N6961, N6940, N6518);
nand NAND4 (N6962, N6958, N866, N756, N5591);
nand NAND3 (N6963, N6962, N3931, N5193);
xor XOR2 (N6964, N6957, N4747);
nand NAND2 (N6965, N6959, N834);
buf BUF1 (N6966, N6961);
and AND4 (N6967, N6945, N2209, N2882, N4140);
xor XOR2 (N6968, N6966, N1857);
and AND2 (N6969, N6964, N781);
or OR4 (N6970, N6965, N2809, N5874, N5619);
or OR2 (N6971, N6948, N3051);
nor NOR4 (N6972, N6967, N2736, N2439, N2030);
xor XOR2 (N6973, N6963, N4136);
xor XOR2 (N6974, N6938, N1695);
and AND2 (N6975, N6972, N1766);
nor NOR3 (N6976, N6975, N1480, N2747);
nand NAND2 (N6977, N6969, N6274);
buf BUF1 (N6978, N6970);
not NOT1 (N6979, N6952);
not NOT1 (N6980, N6971);
or OR4 (N6981, N6978, N4773, N3752, N1584);
buf BUF1 (N6982, N6976);
xor XOR2 (N6983, N6973, N2035);
nor NOR2 (N6984, N6974, N2749);
not NOT1 (N6985, N6968);
xor XOR2 (N6986, N6984, N2335);
nor NOR2 (N6987, N6960, N2680);
nand NAND2 (N6988, N6977, N1393);
and AND2 (N6989, N6981, N2259);
nand NAND3 (N6990, N6987, N3886, N3312);
nand NAND4 (N6991, N6986, N5416, N3926, N4792);
buf BUF1 (N6992, N6985);
and AND2 (N6993, N6988, N6052);
or OR4 (N6994, N6992, N3284, N2096, N696);
not NOT1 (N6995, N6982);
not NOT1 (N6996, N6983);
xor XOR2 (N6997, N6993, N580);
not NOT1 (N6998, N6996);
nand NAND4 (N6999, N6995, N2890, N1460, N3690);
xor XOR2 (N7000, N6989, N4814);
xor XOR2 (N7001, N6998, N6336);
or OR2 (N7002, N6991, N74);
and AND3 (N7003, N6953, N6943, N4970);
buf BUF1 (N7004, N7000);
xor XOR2 (N7005, N6997, N5461);
nor NOR3 (N7006, N7002, N4859, N5097);
buf BUF1 (N7007, N6999);
nand NAND2 (N7008, N7004, N400);
and AND2 (N7009, N7005, N459);
and AND3 (N7010, N6994, N4324, N5740);
nor NOR3 (N7011, N7010, N4420, N3074);
xor XOR2 (N7012, N7001, N4684);
not NOT1 (N7013, N7009);
nor NOR2 (N7014, N7003, N5668);
and AND3 (N7015, N7013, N4990, N3047);
or OR2 (N7016, N7008, N5337);
buf BUF1 (N7017, N7014);
not NOT1 (N7018, N7012);
nor NOR4 (N7019, N7015, N2201, N1462, N5652);
not NOT1 (N7020, N6980);
and AND2 (N7021, N7007, N1997);
xor XOR2 (N7022, N7006, N624);
xor XOR2 (N7023, N7020, N2421);
buf BUF1 (N7024, N7023);
and AND2 (N7025, N6979, N1064);
xor XOR2 (N7026, N7016, N5045);
xor XOR2 (N7027, N7011, N5263);
xor XOR2 (N7028, N7027, N3582);
nand NAND2 (N7029, N7026, N2789);
and AND4 (N7030, N7025, N1018, N6803, N4442);
or OR4 (N7031, N6990, N6112, N6321, N1398);
nand NAND3 (N7032, N7022, N1946, N3345);
nand NAND2 (N7033, N7031, N1904);
not NOT1 (N7034, N7028);
or OR3 (N7035, N7034, N6009, N4330);
xor XOR2 (N7036, N7032, N438);
xor XOR2 (N7037, N7024, N4800);
xor XOR2 (N7038, N7036, N838);
not NOT1 (N7039, N7030);
buf BUF1 (N7040, N7039);
not NOT1 (N7041, N7021);
nand NAND4 (N7042, N7035, N954, N1989, N94);
not NOT1 (N7043, N7018);
xor XOR2 (N7044, N7029, N193);
buf BUF1 (N7045, N7044);
buf BUF1 (N7046, N7017);
and AND3 (N7047, N7037, N1992, N164);
nor NOR3 (N7048, N7045, N4260, N1516);
or OR2 (N7049, N7041, N4471);
nand NAND2 (N7050, N7033, N3319);
xor XOR2 (N7051, N7043, N4612);
not NOT1 (N7052, N7049);
or OR3 (N7053, N7042, N4234, N4443);
not NOT1 (N7054, N7040);
nor NOR2 (N7055, N7050, N1914);
not NOT1 (N7056, N7038);
or OR4 (N7057, N7019, N2068, N5746, N1769);
or OR4 (N7058, N7051, N5841, N6780, N4441);
or OR2 (N7059, N7055, N6021);
nor NOR4 (N7060, N7056, N6416, N7046, N6175);
or OR2 (N7061, N5936, N413);
not NOT1 (N7062, N7058);
nor NOR2 (N7063, N7048, N439);
not NOT1 (N7064, N7062);
buf BUF1 (N7065, N7054);
not NOT1 (N7066, N7047);
xor XOR2 (N7067, N7066, N950);
xor XOR2 (N7068, N7052, N4702);
and AND3 (N7069, N7053, N2779, N2854);
buf BUF1 (N7070, N7064);
nand NAND3 (N7071, N7059, N483, N1531);
not NOT1 (N7072, N7065);
xor XOR2 (N7073, N7060, N4548);
nor NOR2 (N7074, N7069, N2317);
nand NAND4 (N7075, N7072, N1905, N3919, N713);
and AND4 (N7076, N7074, N5749, N497, N6048);
and AND2 (N7077, N7067, N539);
nand NAND2 (N7078, N7070, N877);
not NOT1 (N7079, N7068);
nand NAND2 (N7080, N7071, N1146);
xor XOR2 (N7081, N7075, N2690);
buf BUF1 (N7082, N7057);
or OR3 (N7083, N7077, N5612, N4776);
nand NAND2 (N7084, N7082, N1974);
or OR4 (N7085, N7078, N3478, N4872, N3602);
or OR2 (N7086, N7079, N3547);
buf BUF1 (N7087, N7085);
or OR3 (N7088, N7084, N3367, N4723);
buf BUF1 (N7089, N7073);
nor NOR3 (N7090, N7081, N4795, N3147);
buf BUF1 (N7091, N7086);
buf BUF1 (N7092, N7088);
or OR2 (N7093, N7090, N3354);
not NOT1 (N7094, N7093);
or OR2 (N7095, N7080, N415);
nand NAND2 (N7096, N7092, N1113);
or OR2 (N7097, N7091, N2852);
and AND2 (N7098, N7095, N4796);
or OR2 (N7099, N7076, N6453);
or OR4 (N7100, N7097, N26, N3866, N3822);
or OR4 (N7101, N7096, N5614, N6760, N2337);
nand NAND3 (N7102, N7094, N1293, N7009);
nor NOR2 (N7103, N7083, N4600);
nand NAND2 (N7104, N7087, N3072);
buf BUF1 (N7105, N7063);
not NOT1 (N7106, N7101);
buf BUF1 (N7107, N7106);
nor NOR4 (N7108, N7104, N4982, N6639, N2261);
and AND2 (N7109, N7107, N4991);
buf BUF1 (N7110, N7098);
xor XOR2 (N7111, N7061, N3751);
nand NAND2 (N7112, N7099, N4596);
and AND4 (N7113, N7112, N3547, N728, N6279);
not NOT1 (N7114, N7111);
or OR2 (N7115, N7103, N2592);
xor XOR2 (N7116, N7102, N2524);
nor NOR3 (N7117, N7114, N2538, N453);
nor NOR3 (N7118, N7116, N4886, N5055);
or OR2 (N7119, N7109, N606);
xor XOR2 (N7120, N7105, N4149);
nor NOR3 (N7121, N7113, N130, N1107);
and AND4 (N7122, N7089, N5550, N5772, N5928);
or OR4 (N7123, N7117, N6274, N3544, N2558);
nand NAND2 (N7124, N7115, N3446);
not NOT1 (N7125, N7122);
nor NOR2 (N7126, N7125, N5459);
xor XOR2 (N7127, N7123, N6567);
nand NAND4 (N7128, N7127, N3305, N396, N3942);
buf BUF1 (N7129, N7128);
not NOT1 (N7130, N7110);
or OR2 (N7131, N7108, N18);
buf BUF1 (N7132, N7124);
or OR2 (N7133, N7100, N1402);
buf BUF1 (N7134, N7130);
not NOT1 (N7135, N7133);
xor XOR2 (N7136, N7120, N3446);
buf BUF1 (N7137, N7118);
not NOT1 (N7138, N7119);
not NOT1 (N7139, N7136);
not NOT1 (N7140, N7137);
not NOT1 (N7141, N7140);
buf BUF1 (N7142, N7135);
nand NAND2 (N7143, N7134, N6014);
buf BUF1 (N7144, N7126);
nor NOR4 (N7145, N7141, N3971, N3105, N5168);
nor NOR4 (N7146, N7145, N6591, N2829, N2691);
or OR2 (N7147, N7132, N2386);
not NOT1 (N7148, N7131);
buf BUF1 (N7149, N7148);
buf BUF1 (N7150, N7146);
not NOT1 (N7151, N7147);
not NOT1 (N7152, N7139);
and AND4 (N7153, N7150, N1722, N4353, N6402);
nor NOR2 (N7154, N7143, N5900);
and AND4 (N7155, N7129, N507, N5095, N6190);
nand NAND4 (N7156, N7154, N6721, N2351, N2381);
nor NOR4 (N7157, N7153, N4307, N3038, N3535);
buf BUF1 (N7158, N7157);
xor XOR2 (N7159, N7121, N1609);
and AND2 (N7160, N7152, N5663);
not NOT1 (N7161, N7142);
or OR4 (N7162, N7160, N1553, N7087, N5068);
buf BUF1 (N7163, N7159);
xor XOR2 (N7164, N7138, N7094);
and AND2 (N7165, N7151, N6304);
nor NOR4 (N7166, N7165, N138, N2325, N2736);
xor XOR2 (N7167, N7158, N6486);
and AND2 (N7168, N7164, N953);
nor NOR3 (N7169, N7144, N5849, N204);
nand NAND3 (N7170, N7168, N5644, N6662);
not NOT1 (N7171, N7167);
nor NOR4 (N7172, N7162, N5968, N5958, N2384);
buf BUF1 (N7173, N7172);
not NOT1 (N7174, N7163);
or OR4 (N7175, N7174, N5066, N901, N7051);
nand NAND4 (N7176, N7155, N1735, N5108, N3215);
not NOT1 (N7177, N7169);
nor NOR3 (N7178, N7161, N4426, N4055);
or OR2 (N7179, N7166, N322);
xor XOR2 (N7180, N7178, N1525);
nor NOR2 (N7181, N7180, N2017);
xor XOR2 (N7182, N7177, N722);
nand NAND2 (N7183, N7179, N1985);
or OR2 (N7184, N7170, N1431);
buf BUF1 (N7185, N7181);
nor NOR3 (N7186, N7149, N2139, N3065);
or OR3 (N7187, N7182, N3614, N983);
and AND3 (N7188, N7175, N1152, N2227);
xor XOR2 (N7189, N7185, N3229);
xor XOR2 (N7190, N7171, N6653);
xor XOR2 (N7191, N7184, N5680);
not NOT1 (N7192, N7188);
not NOT1 (N7193, N7183);
nor NOR3 (N7194, N7173, N1721, N5294);
and AND2 (N7195, N7186, N4996);
not NOT1 (N7196, N7192);
buf BUF1 (N7197, N7196);
and AND4 (N7198, N7176, N3916, N1397, N1058);
buf BUF1 (N7199, N7191);
not NOT1 (N7200, N7199);
nor NOR4 (N7201, N7189, N2700, N4200, N1075);
nor NOR3 (N7202, N7156, N5330, N5879);
and AND3 (N7203, N7195, N1225, N1084);
buf BUF1 (N7204, N7187);
not NOT1 (N7205, N7204);
nand NAND2 (N7206, N7200, N3799);
buf BUF1 (N7207, N7198);
nor NOR2 (N7208, N7206, N4763);
nor NOR4 (N7209, N7193, N6968, N6824, N5452);
or OR2 (N7210, N7209, N2907);
nor NOR3 (N7211, N7190, N3532, N2445);
buf BUF1 (N7212, N7202);
not NOT1 (N7213, N7201);
xor XOR2 (N7214, N7213, N7144);
nor NOR4 (N7215, N7214, N5980, N6768, N6868);
buf BUF1 (N7216, N7194);
xor XOR2 (N7217, N7207, N59);
nor NOR4 (N7218, N7217, N4803, N3927, N3500);
xor XOR2 (N7219, N7205, N4781);
not NOT1 (N7220, N7197);
and AND3 (N7221, N7219, N3062, N2171);
and AND4 (N7222, N7208, N5105, N1255, N5860);
xor XOR2 (N7223, N7212, N5769);
and AND2 (N7224, N7222, N4862);
and AND2 (N7225, N7221, N3632);
or OR2 (N7226, N7210, N649);
buf BUF1 (N7227, N7226);
or OR4 (N7228, N7225, N7023, N378, N1543);
xor XOR2 (N7229, N7215, N1917);
not NOT1 (N7230, N7211);
nand NAND4 (N7231, N7224, N6803, N4986, N4720);
xor XOR2 (N7232, N7218, N421);
or OR3 (N7233, N7232, N2486, N2996);
or OR3 (N7234, N7231, N5503, N1733);
and AND3 (N7235, N7223, N5258, N6559);
and AND2 (N7236, N7233, N1986);
or OR2 (N7237, N7236, N6689);
not NOT1 (N7238, N7237);
or OR4 (N7239, N7227, N5576, N1956, N4081);
nand NAND2 (N7240, N7230, N741);
nand NAND4 (N7241, N7228, N1616, N5806, N3944);
nor NOR3 (N7242, N7238, N1248, N392);
not NOT1 (N7243, N7235);
xor XOR2 (N7244, N7220, N2183);
xor XOR2 (N7245, N7241, N6975);
and AND3 (N7246, N7242, N4083, N73);
not NOT1 (N7247, N7240);
xor XOR2 (N7248, N7244, N2485);
buf BUF1 (N7249, N7203);
xor XOR2 (N7250, N7243, N6865);
and AND2 (N7251, N7249, N4640);
not NOT1 (N7252, N7251);
xor XOR2 (N7253, N7229, N7169);
and AND3 (N7254, N7239, N1632, N5520);
nor NOR3 (N7255, N7248, N6, N218);
not NOT1 (N7256, N7253);
nand NAND4 (N7257, N7216, N7188, N3383, N3653);
or OR4 (N7258, N7254, N6343, N627, N4734);
and AND4 (N7259, N7255, N1610, N2302, N1621);
nand NAND2 (N7260, N7258, N1406);
nor NOR4 (N7261, N7250, N3171, N1949, N2331);
xor XOR2 (N7262, N7247, N6598);
or OR2 (N7263, N7256, N6192);
and AND3 (N7264, N7245, N6511, N281);
and AND2 (N7265, N7260, N45);
nor NOR2 (N7266, N7263, N2590);
and AND4 (N7267, N7259, N669, N2054, N3940);
nor NOR4 (N7268, N7261, N4245, N6902, N1042);
and AND4 (N7269, N7265, N4147, N5919, N3775);
and AND2 (N7270, N7264, N4811);
not NOT1 (N7271, N7266);
not NOT1 (N7272, N7234);
xor XOR2 (N7273, N7272, N1836);
xor XOR2 (N7274, N7271, N3717);
not NOT1 (N7275, N7268);
or OR4 (N7276, N7262, N2848, N195, N1031);
nand NAND4 (N7277, N7275, N3378, N4902, N3888);
not NOT1 (N7278, N7277);
xor XOR2 (N7279, N7276, N6803);
or OR2 (N7280, N7267, N3322);
not NOT1 (N7281, N7246);
and AND4 (N7282, N7280, N3163, N6787, N4890);
nand NAND3 (N7283, N7281, N610, N5914);
nand NAND2 (N7284, N7273, N5318);
buf BUF1 (N7285, N7279);
not NOT1 (N7286, N7270);
buf BUF1 (N7287, N7252);
xor XOR2 (N7288, N7257, N1936);
and AND4 (N7289, N7285, N2120, N2656, N5708);
xor XOR2 (N7290, N7282, N654);
nor NOR2 (N7291, N7284, N614);
xor XOR2 (N7292, N7291, N5953);
nor NOR4 (N7293, N7287, N2452, N5749, N5155);
nor NOR4 (N7294, N7289, N894, N281, N1132);
not NOT1 (N7295, N7283);
nor NOR4 (N7296, N7286, N5896, N6983, N789);
buf BUF1 (N7297, N7296);
nand NAND2 (N7298, N7278, N116);
or OR4 (N7299, N7297, N1316, N953, N4520);
nor NOR2 (N7300, N7299, N3787);
nand NAND3 (N7301, N7298, N3740, N4504);
xor XOR2 (N7302, N7295, N1194);
buf BUF1 (N7303, N7301);
xor XOR2 (N7304, N7303, N4414);
buf BUF1 (N7305, N7288);
or OR3 (N7306, N7293, N6983, N5135);
and AND4 (N7307, N7290, N2175, N3667, N4020);
nand NAND4 (N7308, N7307, N3551, N547, N6801);
nor NOR2 (N7309, N7305, N6723);
and AND4 (N7310, N7309, N821, N2638, N2442);
nand NAND2 (N7311, N7310, N6242);
nor NOR4 (N7312, N7302, N4997, N6804, N7265);
and AND4 (N7313, N7294, N1118, N5193, N701);
nor NOR4 (N7314, N7292, N209, N5802, N6153);
and AND4 (N7315, N7313, N3679, N5370, N1317);
and AND2 (N7316, N7274, N2448);
xor XOR2 (N7317, N7312, N5252);
and AND4 (N7318, N7308, N2355, N3078, N6878);
xor XOR2 (N7319, N7314, N6612);
nor NOR4 (N7320, N7269, N1555, N4997, N752);
nor NOR3 (N7321, N7316, N408, N6386);
xor XOR2 (N7322, N7321, N827);
not NOT1 (N7323, N7317);
not NOT1 (N7324, N7315);
and AND2 (N7325, N7311, N6308);
xor XOR2 (N7326, N7300, N4799);
xor XOR2 (N7327, N7325, N2541);
nor NOR4 (N7328, N7327, N2978, N4151, N1263);
and AND3 (N7329, N7304, N6311, N837);
and AND3 (N7330, N7319, N1082, N7088);
nor NOR2 (N7331, N7320, N1143);
xor XOR2 (N7332, N7318, N4086);
buf BUF1 (N7333, N7326);
xor XOR2 (N7334, N7331, N1818);
not NOT1 (N7335, N7322);
or OR2 (N7336, N7330, N2556);
not NOT1 (N7337, N7332);
xor XOR2 (N7338, N7334, N2702);
xor XOR2 (N7339, N7335, N912);
nand NAND3 (N7340, N7339, N140, N4743);
xor XOR2 (N7341, N7328, N4201);
nor NOR2 (N7342, N7324, N652);
buf BUF1 (N7343, N7337);
not NOT1 (N7344, N7342);
xor XOR2 (N7345, N7341, N339);
nand NAND3 (N7346, N7343, N52, N3397);
not NOT1 (N7347, N7340);
xor XOR2 (N7348, N7346, N2910);
nand NAND4 (N7349, N7336, N1370, N6851, N1704);
and AND4 (N7350, N7348, N2259, N2337, N4000);
buf BUF1 (N7351, N7323);
and AND4 (N7352, N7347, N5652, N4643, N2739);
nor NOR2 (N7353, N7338, N4171);
xor XOR2 (N7354, N7349, N5363);
nor NOR4 (N7355, N7345, N2138, N1399, N296);
buf BUF1 (N7356, N7351);
nand NAND2 (N7357, N7306, N4750);
buf BUF1 (N7358, N7329);
not NOT1 (N7359, N7353);
or OR4 (N7360, N7333, N3897, N4845, N402);
or OR3 (N7361, N7355, N3644, N326);
not NOT1 (N7362, N7344);
or OR4 (N7363, N7359, N1919, N3619, N1666);
not NOT1 (N7364, N7360);
and AND2 (N7365, N7363, N2722);
not NOT1 (N7366, N7365);
xor XOR2 (N7367, N7358, N5393);
or OR4 (N7368, N7364, N2185, N7352, N4206);
buf BUF1 (N7369, N3144);
and AND4 (N7370, N7362, N4894, N7331, N6844);
nor NOR3 (N7371, N7356, N5660, N5991);
or OR3 (N7372, N7350, N6411, N6572);
buf BUF1 (N7373, N7366);
nand NAND3 (N7374, N7361, N4889, N4919);
nand NAND3 (N7375, N7368, N543, N5342);
xor XOR2 (N7376, N7357, N530);
not NOT1 (N7377, N7371);
xor XOR2 (N7378, N7374, N995);
buf BUF1 (N7379, N7378);
not NOT1 (N7380, N7372);
nand NAND2 (N7381, N7370, N890);
not NOT1 (N7382, N7354);
or OR4 (N7383, N7373, N6044, N4286, N7330);
buf BUF1 (N7384, N7382);
and AND2 (N7385, N7377, N5356);
buf BUF1 (N7386, N7375);
not NOT1 (N7387, N7381);
nand NAND2 (N7388, N7379, N2774);
xor XOR2 (N7389, N7384, N5827);
xor XOR2 (N7390, N7376, N5531);
and AND4 (N7391, N7383, N2525, N2905, N5439);
nand NAND3 (N7392, N7380, N5491, N4588);
not NOT1 (N7393, N7387);
not NOT1 (N7394, N7390);
buf BUF1 (N7395, N7367);
not NOT1 (N7396, N7369);
or OR4 (N7397, N7391, N5282, N4553, N6989);
nor NOR4 (N7398, N7392, N3839, N107, N6083);
not NOT1 (N7399, N7386);
nor NOR4 (N7400, N7389, N5744, N1004, N2577);
not NOT1 (N7401, N7400);
and AND2 (N7402, N7393, N4021);
and AND3 (N7403, N7398, N1419, N5565);
or OR3 (N7404, N7399, N3083, N3770);
and AND4 (N7405, N7388, N2311, N5388, N6282);
buf BUF1 (N7406, N7405);
nand NAND4 (N7407, N7403, N1421, N2486, N2978);
or OR2 (N7408, N7394, N2826);
or OR2 (N7409, N7406, N5990);
buf BUF1 (N7410, N7395);
nor NOR3 (N7411, N7409, N5519, N4226);
nand NAND4 (N7412, N7385, N1556, N1802, N4404);
and AND4 (N7413, N7404, N458, N978, N6350);
and AND4 (N7414, N7408, N1195, N2411, N3053);
or OR2 (N7415, N7413, N1670);
buf BUF1 (N7416, N7412);
buf BUF1 (N7417, N7397);
and AND2 (N7418, N7417, N7218);
nand NAND3 (N7419, N7416, N2907, N1390);
nand NAND2 (N7420, N7407, N6295);
not NOT1 (N7421, N7418);
buf BUF1 (N7422, N7410);
nand NAND2 (N7423, N7414, N1070);
xor XOR2 (N7424, N7419, N7067);
xor XOR2 (N7425, N7415, N1076);
nor NOR2 (N7426, N7421, N4166);
not NOT1 (N7427, N7426);
nand NAND4 (N7428, N7420, N45, N6780, N3103);
nor NOR4 (N7429, N7396, N1229, N2148, N2921);
nand NAND4 (N7430, N7428, N6385, N1533, N3010);
and AND3 (N7431, N7429, N6479, N3633);
nand NAND4 (N7432, N7427, N2377, N1534, N53);
nor NOR4 (N7433, N7425, N6287, N3271, N3456);
or OR2 (N7434, N7401, N4353);
buf BUF1 (N7435, N7402);
not NOT1 (N7436, N7433);
nor NOR2 (N7437, N7422, N2079);
or OR3 (N7438, N7424, N1749, N1863);
buf BUF1 (N7439, N7411);
xor XOR2 (N7440, N7435, N6802);
nor NOR4 (N7441, N7438, N5270, N119, N6296);
and AND2 (N7442, N7430, N104);
xor XOR2 (N7443, N7434, N917);
or OR3 (N7444, N7439, N4528, N2045);
or OR4 (N7445, N7442, N6103, N1238, N5762);
nor NOR2 (N7446, N7437, N6698);
and AND2 (N7447, N7445, N4260);
or OR4 (N7448, N7444, N2009, N3882, N7179);
and AND4 (N7449, N7431, N2286, N3060, N4072);
or OR4 (N7450, N7436, N4940, N7294, N3201);
nor NOR2 (N7451, N7443, N5379);
xor XOR2 (N7452, N7447, N2088);
not NOT1 (N7453, N7452);
and AND4 (N7454, N7451, N4817, N3921, N7217);
not NOT1 (N7455, N7441);
or OR4 (N7456, N7446, N7155, N2130, N6153);
xor XOR2 (N7457, N7450, N5647);
and AND2 (N7458, N7455, N5872);
nand NAND3 (N7459, N7423, N4552, N2858);
and AND4 (N7460, N7432, N7370, N6777, N3887);
buf BUF1 (N7461, N7456);
xor XOR2 (N7462, N7453, N4431);
buf BUF1 (N7463, N7462);
and AND4 (N7464, N7449, N1955, N7250, N1447);
or OR4 (N7465, N7461, N1300, N4759, N3827);
nand NAND2 (N7466, N7454, N1776);
buf BUF1 (N7467, N7463);
not NOT1 (N7468, N7440);
not NOT1 (N7469, N7457);
not NOT1 (N7470, N7469);
nand NAND2 (N7471, N7448, N1210);
nand NAND4 (N7472, N7471, N2540, N510, N3287);
not NOT1 (N7473, N7460);
buf BUF1 (N7474, N7473);
buf BUF1 (N7475, N7466);
or OR3 (N7476, N7470, N6535, N3797);
not NOT1 (N7477, N7465);
buf BUF1 (N7478, N7464);
buf BUF1 (N7479, N7475);
buf BUF1 (N7480, N7474);
and AND4 (N7481, N7476, N3422, N810, N3789);
nand NAND2 (N7482, N7480, N3786);
or OR4 (N7483, N7478, N2059, N6389, N3596);
and AND2 (N7484, N7458, N2624);
or OR4 (N7485, N7468, N5104, N3313, N1534);
nor NOR3 (N7486, N7459, N807, N6906);
not NOT1 (N7487, N7485);
nor NOR4 (N7488, N7484, N3669, N7068, N4941);
buf BUF1 (N7489, N7487);
nor NOR4 (N7490, N7472, N6113, N5646, N4233);
or OR3 (N7491, N7467, N7266, N5774);
buf BUF1 (N7492, N7490);
nor NOR4 (N7493, N7477, N1370, N5728, N2289);
xor XOR2 (N7494, N7493, N792);
and AND4 (N7495, N7481, N4793, N5841, N6352);
nor NOR4 (N7496, N7486, N3758, N5811, N2691);
or OR4 (N7497, N7488, N178, N5824, N2460);
buf BUF1 (N7498, N7489);
not NOT1 (N7499, N7492);
and AND2 (N7500, N7491, N4282);
xor XOR2 (N7501, N7500, N3002);
or OR4 (N7502, N7497, N571, N573, N7021);
or OR2 (N7503, N7479, N3257);
nand NAND3 (N7504, N7501, N5547, N4178);
buf BUF1 (N7505, N7482);
nand NAND4 (N7506, N7498, N7320, N6643, N4306);
or OR4 (N7507, N7502, N4495, N2122, N1162);
xor XOR2 (N7508, N7505, N6490);
not NOT1 (N7509, N7503);
nor NOR3 (N7510, N7499, N5188, N1704);
not NOT1 (N7511, N7510);
and AND4 (N7512, N7494, N3125, N3973, N2534);
nor NOR4 (N7513, N7483, N3608, N6045, N4960);
xor XOR2 (N7514, N7506, N1493);
not NOT1 (N7515, N7507);
xor XOR2 (N7516, N7512, N6933);
or OR2 (N7517, N7496, N1605);
or OR2 (N7518, N7508, N3937);
or OR4 (N7519, N7515, N6450, N3140, N7116);
and AND2 (N7520, N7509, N878);
and AND3 (N7521, N7514, N5858, N432);
and AND2 (N7522, N7495, N1498);
xor XOR2 (N7523, N7513, N5551);
nor NOR4 (N7524, N7504, N7112, N5844, N2745);
not NOT1 (N7525, N7521);
nand NAND3 (N7526, N7524, N7049, N3531);
xor XOR2 (N7527, N7525, N4306);
buf BUF1 (N7528, N7518);
nor NOR3 (N7529, N7517, N6469, N4760);
buf BUF1 (N7530, N7519);
nand NAND4 (N7531, N7523, N7458, N4810, N5347);
and AND4 (N7532, N7528, N5058, N4317, N4001);
xor XOR2 (N7533, N7526, N6767);
nor NOR2 (N7534, N7530, N6027);
not NOT1 (N7535, N7531);
and AND3 (N7536, N7533, N4440, N5918);
nor NOR2 (N7537, N7534, N3079);
and AND2 (N7538, N7535, N4837);
and AND4 (N7539, N7529, N4959, N1626, N2507);
buf BUF1 (N7540, N7522);
or OR3 (N7541, N7511, N1158, N4158);
nor NOR3 (N7542, N7516, N4774, N1833);
buf BUF1 (N7543, N7539);
xor XOR2 (N7544, N7540, N5961);
xor XOR2 (N7545, N7538, N2813);
not NOT1 (N7546, N7536);
nor NOR3 (N7547, N7520, N5294, N2446);
nand NAND4 (N7548, N7547, N5341, N5155, N4872);
nand NAND2 (N7549, N7548, N7347);
and AND2 (N7550, N7537, N5171);
or OR3 (N7551, N7544, N1405, N1754);
nand NAND2 (N7552, N7543, N4062);
not NOT1 (N7553, N7549);
xor XOR2 (N7554, N7550, N5778);
buf BUF1 (N7555, N7551);
or OR3 (N7556, N7532, N4654, N4991);
and AND2 (N7557, N7542, N1102);
and AND2 (N7558, N7554, N3440);
buf BUF1 (N7559, N7545);
xor XOR2 (N7560, N7558, N4332);
buf BUF1 (N7561, N7546);
xor XOR2 (N7562, N7541, N4341);
nand NAND4 (N7563, N7561, N477, N2763, N2649);
nor NOR2 (N7564, N7552, N2684);
and AND2 (N7565, N7557, N4882);
and AND2 (N7566, N7553, N270);
not NOT1 (N7567, N7564);
xor XOR2 (N7568, N7562, N3487);
buf BUF1 (N7569, N7568);
nor NOR3 (N7570, N7527, N1324, N3069);
nand NAND3 (N7571, N7559, N3444, N6724);
or OR2 (N7572, N7565, N4633);
xor XOR2 (N7573, N7572, N607);
or OR2 (N7574, N7566, N5386);
xor XOR2 (N7575, N7573, N5806);
and AND3 (N7576, N7575, N1993, N5782);
buf BUF1 (N7577, N7560);
buf BUF1 (N7578, N7577);
not NOT1 (N7579, N7569);
xor XOR2 (N7580, N7563, N7354);
not NOT1 (N7581, N7567);
or OR4 (N7582, N7580, N3055, N7393, N3498);
nand NAND3 (N7583, N7574, N3313, N7551);
nor NOR2 (N7584, N7556, N2363);
and AND2 (N7585, N7581, N1457);
nand NAND4 (N7586, N7555, N5848, N446, N7323);
buf BUF1 (N7587, N7571);
buf BUF1 (N7588, N7584);
or OR4 (N7589, N7582, N4462, N247, N3257);
buf BUF1 (N7590, N7583);
xor XOR2 (N7591, N7588, N6077);
or OR2 (N7592, N7587, N7377);
and AND2 (N7593, N7590, N3815);
xor XOR2 (N7594, N7576, N2868);
not NOT1 (N7595, N7579);
nand NAND4 (N7596, N7595, N4578, N5504, N6544);
nor NOR4 (N7597, N7578, N5077, N964, N5865);
or OR4 (N7598, N7591, N5268, N4691, N5015);
nor NOR3 (N7599, N7570, N515, N3038);
or OR2 (N7600, N7585, N1683);
nor NOR2 (N7601, N7596, N7119);
and AND4 (N7602, N7601, N7215, N457, N197);
nand NAND2 (N7603, N7600, N4734);
xor XOR2 (N7604, N7593, N328);
nand NAND4 (N7605, N7594, N3461, N3909, N7569);
or OR4 (N7606, N7605, N3944, N499, N6086);
buf BUF1 (N7607, N7592);
or OR4 (N7608, N7598, N2224, N1541, N6904);
xor XOR2 (N7609, N7599, N1606);
nor NOR2 (N7610, N7589, N4115);
and AND2 (N7611, N7609, N3119);
nor NOR4 (N7612, N7608, N7490, N709, N1862);
xor XOR2 (N7613, N7611, N986);
xor XOR2 (N7614, N7612, N6948);
xor XOR2 (N7615, N7610, N2977);
xor XOR2 (N7616, N7614, N2092);
buf BUF1 (N7617, N7615);
and AND4 (N7618, N7604, N6342, N1271, N471);
nor NOR2 (N7619, N7606, N7064);
or OR2 (N7620, N7618, N5301);
or OR4 (N7621, N7616, N5029, N6698, N7438);
xor XOR2 (N7622, N7607, N6243);
nand NAND2 (N7623, N7586, N5013);
and AND4 (N7624, N7619, N1308, N1372, N491);
and AND4 (N7625, N7603, N5706, N4693, N3270);
not NOT1 (N7626, N7597);
buf BUF1 (N7627, N7623);
and AND2 (N7628, N7617, N6282);
nand NAND3 (N7629, N7620, N2720, N1752);
not NOT1 (N7630, N7622);
buf BUF1 (N7631, N7626);
nand NAND2 (N7632, N7628, N556);
nand NAND2 (N7633, N7631, N7418);
buf BUF1 (N7634, N7602);
nand NAND3 (N7635, N7632, N1639, N6295);
and AND2 (N7636, N7625, N3688);
buf BUF1 (N7637, N7621);
nor NOR3 (N7638, N7637, N3885, N2945);
buf BUF1 (N7639, N7629);
nor NOR4 (N7640, N7639, N4875, N1440, N1215);
not NOT1 (N7641, N7640);
nand NAND4 (N7642, N7635, N6610, N3959, N2359);
buf BUF1 (N7643, N7636);
not NOT1 (N7644, N7613);
buf BUF1 (N7645, N7641);
buf BUF1 (N7646, N7630);
and AND3 (N7647, N7638, N4499, N4080);
nand NAND2 (N7648, N7634, N1032);
buf BUF1 (N7649, N7642);
xor XOR2 (N7650, N7648, N232);
and AND3 (N7651, N7646, N6069, N7051);
nand NAND3 (N7652, N7627, N6441, N6874);
and AND4 (N7653, N7652, N5413, N4587, N1659);
xor XOR2 (N7654, N7653, N6712);
not NOT1 (N7655, N7650);
nand NAND3 (N7656, N7624, N1566, N5580);
not NOT1 (N7657, N7656);
or OR2 (N7658, N7654, N1709);
xor XOR2 (N7659, N7655, N5557);
nand NAND3 (N7660, N7649, N3852, N7481);
nand NAND2 (N7661, N7633, N4230);
and AND4 (N7662, N7647, N2371, N114, N6438);
buf BUF1 (N7663, N7659);
not NOT1 (N7664, N7645);
xor XOR2 (N7665, N7657, N5752);
nor NOR4 (N7666, N7665, N6933, N3821, N1980);
nand NAND2 (N7667, N7663, N1854);
nor NOR4 (N7668, N7664, N4220, N233, N6810);
or OR3 (N7669, N7658, N1954, N4303);
nand NAND4 (N7670, N7667, N5638, N2116, N4339);
nand NAND2 (N7671, N7643, N7349);
nor NOR2 (N7672, N7662, N7326);
nor NOR4 (N7673, N7669, N2898, N665, N3904);
or OR2 (N7674, N7671, N4905);
buf BUF1 (N7675, N7674);
or OR2 (N7676, N7675, N411);
nor NOR4 (N7677, N7644, N134, N597, N5413);
not NOT1 (N7678, N7670);
and AND4 (N7679, N7651, N6911, N4628, N2098);
nand NAND2 (N7680, N7678, N6085);
nand NAND4 (N7681, N7677, N1463, N1845, N6837);
nor NOR4 (N7682, N7672, N3484, N5632, N5888);
xor XOR2 (N7683, N7668, N6427);
buf BUF1 (N7684, N7680);
nand NAND3 (N7685, N7684, N882, N4070);
not NOT1 (N7686, N7681);
xor XOR2 (N7687, N7661, N278);
or OR4 (N7688, N7687, N7240, N1892, N6099);
buf BUF1 (N7689, N7666);
and AND3 (N7690, N7679, N4855, N4979);
xor XOR2 (N7691, N7690, N3472);
nor NOR4 (N7692, N7689, N705, N2779, N3177);
or OR4 (N7693, N7683, N2642, N6723, N6733);
not NOT1 (N7694, N7693);
xor XOR2 (N7695, N7673, N583);
or OR3 (N7696, N7691, N6133, N2484);
nor NOR2 (N7697, N7676, N1787);
or OR2 (N7698, N7682, N1732);
nand NAND4 (N7699, N7695, N4841, N7630, N6687);
xor XOR2 (N7700, N7686, N1949);
buf BUF1 (N7701, N7700);
not NOT1 (N7702, N7660);
not NOT1 (N7703, N7699);
not NOT1 (N7704, N7685);
or OR2 (N7705, N7697, N5927);
buf BUF1 (N7706, N7701);
buf BUF1 (N7707, N7703);
and AND3 (N7708, N7696, N3758, N6096);
or OR4 (N7709, N7705, N2543, N4767, N5830);
nand NAND2 (N7710, N7709, N1936);
and AND2 (N7711, N7707, N5347);
or OR2 (N7712, N7704, N1610);
not NOT1 (N7713, N7710);
buf BUF1 (N7714, N7688);
or OR2 (N7715, N7708, N4610);
nand NAND2 (N7716, N7698, N870);
nor NOR2 (N7717, N7712, N4685);
nand NAND3 (N7718, N7702, N7659, N2322);
or OR3 (N7719, N7718, N4287, N693);
xor XOR2 (N7720, N7694, N5734);
and AND2 (N7721, N7714, N3459);
nand NAND2 (N7722, N7717, N2674);
or OR4 (N7723, N7715, N2650, N1805, N6014);
and AND3 (N7724, N7711, N1214, N2487);
nand NAND3 (N7725, N7719, N3520, N3327);
or OR4 (N7726, N7722, N2039, N2163, N4553);
buf BUF1 (N7727, N7713);
not NOT1 (N7728, N7724);
nor NOR2 (N7729, N7725, N2608);
nor NOR4 (N7730, N7723, N2593, N1796, N558);
buf BUF1 (N7731, N7726);
xor XOR2 (N7732, N7731, N4649);
xor XOR2 (N7733, N7716, N5698);
not NOT1 (N7734, N7706);
not NOT1 (N7735, N7730);
xor XOR2 (N7736, N7728, N1912);
and AND2 (N7737, N7692, N4103);
xor XOR2 (N7738, N7737, N5734);
or OR4 (N7739, N7732, N3781, N6461, N4137);
xor XOR2 (N7740, N7720, N6562);
buf BUF1 (N7741, N7736);
nor NOR2 (N7742, N7734, N4770);
nand NAND2 (N7743, N7739, N3802);
or OR3 (N7744, N7742, N6407, N3211);
xor XOR2 (N7745, N7729, N1126);
or OR2 (N7746, N7744, N4564);
nor NOR4 (N7747, N7745, N7456, N5547, N3583);
not NOT1 (N7748, N7735);
xor XOR2 (N7749, N7738, N96);
and AND4 (N7750, N7743, N2309, N374, N7618);
nor NOR4 (N7751, N7749, N1968, N6388, N5182);
or OR4 (N7752, N7750, N2578, N7271, N5470);
not NOT1 (N7753, N7740);
nand NAND4 (N7754, N7747, N1441, N2202, N1851);
not NOT1 (N7755, N7733);
or OR3 (N7756, N7748, N3288, N921);
and AND4 (N7757, N7753, N6777, N3231, N3687);
or OR3 (N7758, N7721, N6081, N466);
or OR3 (N7759, N7757, N1323, N5163);
not NOT1 (N7760, N7758);
not NOT1 (N7761, N7752);
or OR3 (N7762, N7751, N5199, N1051);
buf BUF1 (N7763, N7727);
nor NOR4 (N7764, N7761, N6847, N6669, N5423);
and AND4 (N7765, N7754, N75, N6172, N3309);
not NOT1 (N7766, N7762);
nor NOR3 (N7767, N7763, N2178, N3689);
xor XOR2 (N7768, N7764, N3631);
and AND2 (N7769, N7759, N5876);
nor NOR3 (N7770, N7741, N5992, N3198);
or OR3 (N7771, N7766, N5499, N3154);
not NOT1 (N7772, N7760);
nand NAND4 (N7773, N7771, N2565, N6713, N6607);
and AND2 (N7774, N7773, N1349);
xor XOR2 (N7775, N7768, N6733);
and AND4 (N7776, N7775, N612, N6570, N221);
not NOT1 (N7777, N7765);
buf BUF1 (N7778, N7774);
or OR2 (N7779, N7772, N4878);
buf BUF1 (N7780, N7779);
xor XOR2 (N7781, N7776, N4816);
buf BUF1 (N7782, N7770);
nand NAND2 (N7783, N7767, N3094);
nor NOR3 (N7784, N7756, N2074, N2077);
nor NOR2 (N7785, N7769, N5772);
buf BUF1 (N7786, N7778);
xor XOR2 (N7787, N7782, N6718);
xor XOR2 (N7788, N7785, N7187);
nand NAND3 (N7789, N7788, N533, N6529);
not NOT1 (N7790, N7777);
or OR2 (N7791, N7781, N7443);
buf BUF1 (N7792, N7790);
not NOT1 (N7793, N7787);
buf BUF1 (N7794, N7783);
nand NAND3 (N7795, N7784, N6019, N1823);
buf BUF1 (N7796, N7780);
xor XOR2 (N7797, N7791, N1341);
nor NOR2 (N7798, N7793, N7204);
xor XOR2 (N7799, N7789, N4642);
nor NOR4 (N7800, N7795, N2653, N122, N3038);
xor XOR2 (N7801, N7800, N3790);
nand NAND3 (N7802, N7796, N3261, N4072);
nand NAND3 (N7803, N7801, N26, N4244);
xor XOR2 (N7804, N7797, N5810);
buf BUF1 (N7805, N7798);
nand NAND3 (N7806, N7805, N2906, N6738);
not NOT1 (N7807, N7804);
or OR3 (N7808, N7746, N1509, N3407);
and AND2 (N7809, N7806, N1644);
not NOT1 (N7810, N7799);
or OR4 (N7811, N7792, N7695, N6516, N5242);
xor XOR2 (N7812, N7803, N2760);
not NOT1 (N7813, N7755);
or OR4 (N7814, N7813, N4098, N3202, N6672);
and AND2 (N7815, N7808, N6500);
xor XOR2 (N7816, N7814, N6099);
nand NAND3 (N7817, N7809, N369, N5571);
not NOT1 (N7818, N7811);
and AND4 (N7819, N7794, N6376, N7592, N1123);
and AND2 (N7820, N7816, N2380);
nand NAND2 (N7821, N7820, N489);
buf BUF1 (N7822, N7812);
and AND4 (N7823, N7818, N6764, N60, N469);
and AND4 (N7824, N7807, N5897, N5845, N180);
nand NAND2 (N7825, N7815, N3379);
and AND3 (N7826, N7786, N2233, N7634);
nand NAND4 (N7827, N7825, N4021, N6223, N7106);
nor NOR4 (N7828, N7823, N5448, N5919, N1355);
nor NOR2 (N7829, N7822, N5067);
not NOT1 (N7830, N7827);
not NOT1 (N7831, N7824);
xor XOR2 (N7832, N7830, N7537);
not NOT1 (N7833, N7810);
nor NOR2 (N7834, N7829, N5990);
nor NOR3 (N7835, N7828, N1216, N2989);
nand NAND4 (N7836, N7819, N864, N3407, N3830);
not NOT1 (N7837, N7836);
nand NAND2 (N7838, N7834, N6338);
xor XOR2 (N7839, N7835, N1320);
xor XOR2 (N7840, N7832, N6148);
not NOT1 (N7841, N7840);
nand NAND2 (N7842, N7833, N5974);
nor NOR4 (N7843, N7817, N4295, N93, N507);
or OR4 (N7844, N7841, N1366, N3714, N5310);
nand NAND3 (N7845, N7831, N5285, N2803);
or OR2 (N7846, N7839, N6656);
or OR4 (N7847, N7843, N61, N872, N7349);
or OR3 (N7848, N7821, N6284, N7571);
nand NAND3 (N7849, N7845, N20, N4237);
or OR3 (N7850, N7837, N2678, N2668);
not NOT1 (N7851, N7846);
buf BUF1 (N7852, N7851);
xor XOR2 (N7853, N7844, N6808);
not NOT1 (N7854, N7852);
xor XOR2 (N7855, N7842, N3262);
and AND2 (N7856, N7854, N4175);
buf BUF1 (N7857, N7838);
and AND2 (N7858, N7848, N2717);
and AND3 (N7859, N7826, N4798, N6073);
or OR3 (N7860, N7856, N5419, N1157);
not NOT1 (N7861, N7853);
and AND3 (N7862, N7855, N4809, N1553);
nand NAND3 (N7863, N7847, N3250, N2063);
nor NOR4 (N7864, N7850, N6349, N7339, N1064);
and AND2 (N7865, N7859, N603);
or OR4 (N7866, N7862, N598, N494, N7213);
buf BUF1 (N7867, N7802);
nor NOR2 (N7868, N7849, N571);
nand NAND4 (N7869, N7860, N5428, N7711, N3974);
xor XOR2 (N7870, N7861, N1016);
buf BUF1 (N7871, N7857);
nor NOR3 (N7872, N7871, N1924, N4841);
xor XOR2 (N7873, N7870, N5039);
and AND3 (N7874, N7866, N311, N483);
nor NOR2 (N7875, N7863, N4086);
nand NAND2 (N7876, N7867, N7280);
and AND4 (N7877, N7876, N6097, N473, N7036);
and AND4 (N7878, N7875, N6991, N641, N4107);
nor NOR4 (N7879, N7874, N1619, N2843, N3037);
buf BUF1 (N7880, N7877);
nand NAND3 (N7881, N7880, N2645, N15);
nand NAND2 (N7882, N7858, N4874);
not NOT1 (N7883, N7881);
xor XOR2 (N7884, N7869, N557);
not NOT1 (N7885, N7878);
nor NOR3 (N7886, N7872, N3962, N5586);
xor XOR2 (N7887, N7884, N7129);
buf BUF1 (N7888, N7865);
or OR3 (N7889, N7887, N376, N3426);
xor XOR2 (N7890, N7879, N5556);
nand NAND3 (N7891, N7888, N3512, N5953);
buf BUF1 (N7892, N7868);
not NOT1 (N7893, N7885);
or OR2 (N7894, N7892, N3663);
nand NAND3 (N7895, N7891, N5748, N569);
nor NOR2 (N7896, N7873, N6015);
xor XOR2 (N7897, N7883, N4961);
and AND2 (N7898, N7896, N262);
or OR4 (N7899, N7894, N5198, N3297, N5490);
xor XOR2 (N7900, N7897, N1845);
and AND2 (N7901, N7899, N4240);
nand NAND3 (N7902, N7895, N2625, N7093);
or OR3 (N7903, N7898, N4041, N5300);
nor NOR3 (N7904, N7901, N803, N6364);
and AND3 (N7905, N7864, N6614, N5947);
buf BUF1 (N7906, N7900);
or OR2 (N7907, N7906, N5437);
nand NAND3 (N7908, N7889, N1648, N5617);
and AND2 (N7909, N7904, N5181);
nor NOR3 (N7910, N7882, N1909, N1139);
nor NOR3 (N7911, N7903, N7271, N7419);
nand NAND4 (N7912, N7910, N707, N4476, N1658);
nor NOR4 (N7913, N7886, N4682, N1577, N4693);
not NOT1 (N7914, N7902);
and AND2 (N7915, N7908, N2595);
or OR3 (N7916, N7905, N1389, N4080);
and AND3 (N7917, N7911, N6160, N7411);
buf BUF1 (N7918, N7917);
or OR4 (N7919, N7907, N4709, N7621, N4176);
nor NOR2 (N7920, N7915, N6336);
nor NOR3 (N7921, N7918, N6049, N1692);
xor XOR2 (N7922, N7890, N4673);
xor XOR2 (N7923, N7914, N4141);
nand NAND2 (N7924, N7913, N5859);
nand NAND3 (N7925, N7924, N1987, N5549);
not NOT1 (N7926, N7921);
buf BUF1 (N7927, N7925);
xor XOR2 (N7928, N7920, N19);
or OR3 (N7929, N7928, N2769, N2290);
not NOT1 (N7930, N7909);
nor NOR4 (N7931, N7893, N3199, N5050, N3072);
buf BUF1 (N7932, N7929);
xor XOR2 (N7933, N7926, N3796);
buf BUF1 (N7934, N7931);
xor XOR2 (N7935, N7919, N1374);
and AND2 (N7936, N7933, N4600);
not NOT1 (N7937, N7930);
nand NAND2 (N7938, N7916, N6143);
not NOT1 (N7939, N7912);
nand NAND3 (N7940, N7923, N3966, N1865);
xor XOR2 (N7941, N7938, N6511);
nor NOR4 (N7942, N7922, N7747, N5016, N6260);
not NOT1 (N7943, N7934);
xor XOR2 (N7944, N7936, N3569);
and AND4 (N7945, N7943, N5430, N4203, N3530);
not NOT1 (N7946, N7945);
xor XOR2 (N7947, N7946, N2145);
and AND4 (N7948, N7942, N4828, N1891, N4027);
and AND4 (N7949, N7932, N1440, N1324, N7332);
xor XOR2 (N7950, N7948, N3911);
buf BUF1 (N7951, N7937);
buf BUF1 (N7952, N7944);
and AND2 (N7953, N7952, N7781);
nor NOR3 (N7954, N7941, N8, N4994);
nor NOR3 (N7955, N7949, N166, N3576);
buf BUF1 (N7956, N7955);
buf BUF1 (N7957, N7950);
nand NAND2 (N7958, N7951, N2880);
xor XOR2 (N7959, N7954, N1423);
or OR2 (N7960, N7947, N4570);
not NOT1 (N7961, N7939);
and AND4 (N7962, N7957, N2009, N3252, N4810);
nand NAND4 (N7963, N7962, N2002, N6395, N4369);
nand NAND4 (N7964, N7956, N5230, N4475, N6495);
not NOT1 (N7965, N7964);
nor NOR4 (N7966, N7953, N7157, N2247, N1429);
nand NAND2 (N7967, N7959, N356);
buf BUF1 (N7968, N7958);
and AND4 (N7969, N7935, N3507, N7706, N5687);
and AND3 (N7970, N7961, N4874, N183);
not NOT1 (N7971, N7960);
buf BUF1 (N7972, N7927);
and AND4 (N7973, N7970, N3994, N3498, N1221);
nand NAND3 (N7974, N7968, N2391, N2991);
nand NAND4 (N7975, N7965, N1545, N4470, N2653);
buf BUF1 (N7976, N7974);
and AND3 (N7977, N7973, N4619, N4542);
xor XOR2 (N7978, N7969, N3003);
or OR3 (N7979, N7966, N2900, N7864);
nor NOR4 (N7980, N7976, N5828, N2488, N5250);
nand NAND2 (N7981, N7963, N2724);
and AND3 (N7982, N7977, N6273, N5577);
nand NAND3 (N7983, N7979, N3580, N4116);
xor XOR2 (N7984, N7967, N3239);
or OR3 (N7985, N7975, N5103, N3889);
xor XOR2 (N7986, N7971, N2153);
or OR2 (N7987, N7981, N4813);
xor XOR2 (N7988, N7985, N856);
xor XOR2 (N7989, N7987, N7417);
not NOT1 (N7990, N7972);
or OR2 (N7991, N7986, N3291);
xor XOR2 (N7992, N7940, N3613);
or OR4 (N7993, N7980, N4600, N2256, N3543);
and AND3 (N7994, N7991, N3903, N2776);
not NOT1 (N7995, N7989);
xor XOR2 (N7996, N7982, N2663);
buf BUF1 (N7997, N7988);
buf BUF1 (N7998, N7984);
or OR4 (N7999, N7978, N2080, N6253, N7159);
not NOT1 (N8000, N7983);
or OR4 (N8001, N7994, N285, N1974, N6144);
not NOT1 (N8002, N7993);
and AND2 (N8003, N7997, N3970);
nor NOR2 (N8004, N7992, N5969);
nor NOR3 (N8005, N8000, N4774, N3269);
buf BUF1 (N8006, N8004);
nand NAND4 (N8007, N8006, N6875, N2657, N1356);
nand NAND2 (N8008, N8005, N7134);
buf BUF1 (N8009, N8001);
xor XOR2 (N8010, N7999, N1058);
xor XOR2 (N8011, N8003, N6433);
nor NOR3 (N8012, N8011, N988, N4204);
xor XOR2 (N8013, N8007, N7757);
nor NOR2 (N8014, N7990, N1644);
not NOT1 (N8015, N8002);
or OR4 (N8016, N8015, N3275, N2289, N886);
or OR3 (N8017, N8016, N5378, N6564);
or OR4 (N8018, N8010, N6196, N4627, N5326);
or OR3 (N8019, N8008, N4678, N4880);
buf BUF1 (N8020, N8012);
not NOT1 (N8021, N8014);
nand NAND4 (N8022, N8009, N6502, N2499, N6577);
nor NOR4 (N8023, N8021, N5339, N4131, N1941);
nand NAND2 (N8024, N8019, N5132);
xor XOR2 (N8025, N8013, N759);
not NOT1 (N8026, N8023);
or OR4 (N8027, N8020, N4357, N1938, N1348);
xor XOR2 (N8028, N7998, N2880);
nor NOR3 (N8029, N8022, N2991, N472);
or OR3 (N8030, N8026, N3568, N4242);
not NOT1 (N8031, N8025);
nor NOR2 (N8032, N8030, N5856);
not NOT1 (N8033, N8029);
not NOT1 (N8034, N7995);
or OR2 (N8035, N8018, N2377);
buf BUF1 (N8036, N8024);
nor NOR2 (N8037, N8028, N5602);
not NOT1 (N8038, N8031);
not NOT1 (N8039, N8034);
nor NOR4 (N8040, N8017, N7054, N7512, N7871);
not NOT1 (N8041, N8039);
nor NOR3 (N8042, N8038, N4288, N1908);
xor XOR2 (N8043, N8035, N7914);
nor NOR3 (N8044, N8036, N6447, N3610);
not NOT1 (N8045, N8032);
and AND4 (N8046, N8041, N4277, N4171, N2486);
nor NOR3 (N8047, N8027, N1985, N6057);
or OR2 (N8048, N8042, N1223);
nand NAND4 (N8049, N8033, N3257, N4015, N5761);
or OR3 (N8050, N8037, N652, N525);
and AND3 (N8051, N8047, N495, N4514);
and AND3 (N8052, N8040, N7104, N2538);
xor XOR2 (N8053, N8043, N5780);
nand NAND4 (N8054, N8051, N3040, N7072, N60);
nand NAND2 (N8055, N8045, N1933);
nor NOR3 (N8056, N8048, N860, N383);
not NOT1 (N8057, N8044);
nand NAND4 (N8058, N8050, N3841, N8028, N2725);
not NOT1 (N8059, N8054);
or OR2 (N8060, N8055, N2802);
buf BUF1 (N8061, N8049);
buf BUF1 (N8062, N8061);
xor XOR2 (N8063, N8062, N7176);
buf BUF1 (N8064, N8052);
nand NAND2 (N8065, N7996, N7807);
nand NAND4 (N8066, N8053, N1546, N5669, N393);
xor XOR2 (N8067, N8058, N2793);
nor NOR2 (N8068, N8063, N4929);
or OR3 (N8069, N8064, N4838, N4003);
xor XOR2 (N8070, N8057, N2433);
xor XOR2 (N8071, N8046, N4116);
buf BUF1 (N8072, N8071);
buf BUF1 (N8073, N8060);
nor NOR3 (N8074, N8069, N4630, N2905);
not NOT1 (N8075, N8068);
and AND4 (N8076, N8075, N2232, N2895, N6043);
not NOT1 (N8077, N8056);
xor XOR2 (N8078, N8066, N1913);
buf BUF1 (N8079, N8065);
or OR4 (N8080, N8077, N7283, N7200, N6995);
nand NAND3 (N8081, N8079, N7768, N2026);
and AND3 (N8082, N8081, N6256, N1159);
nor NOR3 (N8083, N8072, N6505, N5488);
xor XOR2 (N8084, N8076, N2527);
not NOT1 (N8085, N8080);
xor XOR2 (N8086, N8059, N2796);
buf BUF1 (N8087, N8083);
or OR2 (N8088, N8067, N2138);
not NOT1 (N8089, N8070);
not NOT1 (N8090, N8085);
nor NOR4 (N8091, N8078, N539, N2150, N7334);
or OR3 (N8092, N8086, N6563, N3631);
buf BUF1 (N8093, N8092);
buf BUF1 (N8094, N8091);
or OR3 (N8095, N8093, N5723, N6185);
and AND2 (N8096, N8095, N5644);
and AND3 (N8097, N8089, N4399, N1204);
not NOT1 (N8098, N8096);
nor NOR2 (N8099, N8088, N7632);
not NOT1 (N8100, N8082);
buf BUF1 (N8101, N8094);
not NOT1 (N8102, N8098);
nand NAND4 (N8103, N8087, N4109, N5095, N138);
and AND3 (N8104, N8103, N2909, N6822);
buf BUF1 (N8105, N8073);
and AND2 (N8106, N8105, N2739);
not NOT1 (N8107, N8100);
not NOT1 (N8108, N8107);
or OR4 (N8109, N8106, N1296, N6142, N1317);
not NOT1 (N8110, N8101);
nor NOR3 (N8111, N8102, N3608, N8036);
or OR3 (N8112, N8099, N4008, N5112);
or OR2 (N8113, N8110, N425);
nand NAND3 (N8114, N8109, N3270, N3320);
xor XOR2 (N8115, N8111, N7138);
not NOT1 (N8116, N8108);
xor XOR2 (N8117, N8097, N7568);
nand NAND3 (N8118, N8074, N229, N1585);
and AND4 (N8119, N8113, N4917, N6137, N7916);
buf BUF1 (N8120, N8090);
nand NAND2 (N8121, N8114, N3863);
xor XOR2 (N8122, N8104, N7978);
not NOT1 (N8123, N8117);
nor NOR2 (N8124, N8116, N6784);
and AND4 (N8125, N8118, N5298, N3250, N1249);
nand NAND3 (N8126, N8120, N1822, N2824);
xor XOR2 (N8127, N8126, N5919);
nor NOR3 (N8128, N8127, N246, N3584);
nand NAND4 (N8129, N8119, N6463, N2358, N7472);
nand NAND4 (N8130, N8115, N5469, N199, N3);
buf BUF1 (N8131, N8084);
not NOT1 (N8132, N8128);
and AND2 (N8133, N8131, N6292);
nor NOR4 (N8134, N8121, N1752, N3200, N2812);
nand NAND4 (N8135, N8124, N5127, N7630, N61);
nor NOR3 (N8136, N8112, N7932, N120);
nor NOR2 (N8137, N8135, N6283);
nand NAND3 (N8138, N8130, N4824, N6571);
or OR2 (N8139, N8125, N7963);
nor NOR2 (N8140, N8138, N7979);
buf BUF1 (N8141, N8123);
xor XOR2 (N8142, N8132, N2285);
or OR2 (N8143, N8134, N7302);
nand NAND4 (N8144, N8137, N7462, N3399, N1857);
buf BUF1 (N8145, N8136);
nor NOR3 (N8146, N8133, N5877, N4626);
not NOT1 (N8147, N8145);
not NOT1 (N8148, N8141);
buf BUF1 (N8149, N8146);
not NOT1 (N8150, N8144);
nand NAND3 (N8151, N8122, N5226, N2295);
xor XOR2 (N8152, N8149, N3989);
buf BUF1 (N8153, N8151);
buf BUF1 (N8154, N8142);
nor NOR2 (N8155, N8143, N6763);
or OR3 (N8156, N8140, N6699, N1495);
nor NOR3 (N8157, N8152, N779, N5541);
or OR2 (N8158, N8155, N4604);
xor XOR2 (N8159, N8154, N5677);
buf BUF1 (N8160, N8150);
and AND2 (N8161, N8156, N125);
buf BUF1 (N8162, N8161);
not NOT1 (N8163, N8147);
not NOT1 (N8164, N8158);
and AND4 (N8165, N8153, N4958, N5668, N3887);
nor NOR2 (N8166, N8139, N3338);
nor NOR2 (N8167, N8166, N3358);
xor XOR2 (N8168, N8164, N5907);
nand NAND2 (N8169, N8163, N3853);
nor NOR2 (N8170, N8157, N449);
xor XOR2 (N8171, N8160, N560);
and AND2 (N8172, N8171, N6879);
buf BUF1 (N8173, N8168);
buf BUF1 (N8174, N8165);
or OR2 (N8175, N8167, N7369);
not NOT1 (N8176, N8169);
nor NOR3 (N8177, N8172, N4989, N679);
nand NAND2 (N8178, N8162, N3021);
xor XOR2 (N8179, N8178, N2116);
nor NOR3 (N8180, N8129, N4037, N4723);
and AND2 (N8181, N8175, N8133);
nand NAND4 (N8182, N8148, N4025, N6964, N628);
or OR4 (N8183, N8170, N4249, N4190, N2225);
buf BUF1 (N8184, N8177);
nor NOR2 (N8185, N8176, N4521);
xor XOR2 (N8186, N8173, N5446);
nor NOR4 (N8187, N8180, N5864, N6689, N4214);
nor NOR4 (N8188, N8183, N6499, N8185, N82);
nand NAND2 (N8189, N1941, N5742);
not NOT1 (N8190, N8187);
nand NAND2 (N8191, N8174, N764);
and AND3 (N8192, N8181, N5182, N39);
nor NOR2 (N8193, N8191, N8002);
nor NOR4 (N8194, N8179, N5774, N6137, N6822);
nand NAND2 (N8195, N8192, N5333);
and AND2 (N8196, N8194, N3187);
buf BUF1 (N8197, N8186);
xor XOR2 (N8198, N8195, N4931);
and AND3 (N8199, N8182, N1749, N4806);
and AND2 (N8200, N8193, N2816);
nor NOR2 (N8201, N8200, N5801);
or OR2 (N8202, N8159, N6071);
nor NOR4 (N8203, N8202, N5904, N410, N7440);
xor XOR2 (N8204, N8198, N5620);
xor XOR2 (N8205, N8190, N7149);
buf BUF1 (N8206, N8204);
nor NOR4 (N8207, N8184, N5211, N4140, N8160);
and AND3 (N8208, N8197, N5803, N7933);
buf BUF1 (N8209, N8196);
xor XOR2 (N8210, N8189, N1550);
nor NOR3 (N8211, N8201, N1728, N7329);
nor NOR2 (N8212, N8211, N3521);
buf BUF1 (N8213, N8209);
or OR4 (N8214, N8199, N52, N6694, N366);
and AND2 (N8215, N8203, N3066);
nand NAND3 (N8216, N8208, N1451, N7820);
nand NAND2 (N8217, N8188, N96);
nand NAND2 (N8218, N8210, N5165);
or OR4 (N8219, N8205, N5251, N70, N3676);
not NOT1 (N8220, N8206);
nor NOR2 (N8221, N8218, N627);
and AND2 (N8222, N8213, N6725);
nand NAND2 (N8223, N8207, N3029);
or OR2 (N8224, N8220, N2614);
xor XOR2 (N8225, N8219, N2661);
and AND2 (N8226, N8212, N1132);
and AND3 (N8227, N8215, N7534, N2224);
and AND2 (N8228, N8227, N1872);
buf BUF1 (N8229, N8217);
or OR3 (N8230, N8216, N1156, N5742);
and AND3 (N8231, N8226, N1431, N3387);
and AND4 (N8232, N8224, N1788, N8124, N5092);
or OR3 (N8233, N8231, N5229, N5466);
or OR4 (N8234, N8229, N6660, N2259, N2308);
buf BUF1 (N8235, N8221);
nor NOR2 (N8236, N8228, N163);
not NOT1 (N8237, N8225);
buf BUF1 (N8238, N8223);
and AND2 (N8239, N8237, N3467);
buf BUF1 (N8240, N8238);
or OR4 (N8241, N8239, N3116, N7872, N7170);
not NOT1 (N8242, N8240);
nor NOR4 (N8243, N8242, N5183, N836, N785);
buf BUF1 (N8244, N8230);
buf BUF1 (N8245, N8234);
not NOT1 (N8246, N8232);
nand NAND4 (N8247, N8246, N351, N325, N2813);
nor NOR3 (N8248, N8233, N426, N2669);
buf BUF1 (N8249, N8243);
and AND4 (N8250, N8236, N913, N2857, N935);
not NOT1 (N8251, N8248);
xor XOR2 (N8252, N8241, N6696);
buf BUF1 (N8253, N8251);
buf BUF1 (N8254, N8253);
and AND3 (N8255, N8214, N820, N6196);
nor NOR4 (N8256, N8254, N5148, N1320, N505);
and AND4 (N8257, N8222, N3428, N1879, N1967);
xor XOR2 (N8258, N8247, N987);
or OR4 (N8259, N8252, N2955, N7954, N7113);
nand NAND4 (N8260, N8249, N3797, N7435, N3112);
and AND3 (N8261, N8257, N5717, N4211);
not NOT1 (N8262, N8259);
buf BUF1 (N8263, N8245);
buf BUF1 (N8264, N8235);
xor XOR2 (N8265, N8255, N3132);
nor NOR4 (N8266, N8265, N2233, N1765, N7349);
and AND2 (N8267, N8263, N6878);
or OR2 (N8268, N8250, N1027);
xor XOR2 (N8269, N8268, N7724);
xor XOR2 (N8270, N8244, N7953);
or OR2 (N8271, N8270, N6711);
or OR2 (N8272, N8256, N1246);
not NOT1 (N8273, N8271);
nor NOR4 (N8274, N8262, N4661, N3558, N3442);
xor XOR2 (N8275, N8274, N3301);
nor NOR4 (N8276, N8258, N6982, N2809, N6476);
and AND3 (N8277, N8266, N323, N525);
and AND4 (N8278, N8267, N3650, N3520, N828);
nand NAND3 (N8279, N8273, N6252, N2553);
or OR4 (N8280, N8260, N431, N91, N8071);
nor NOR2 (N8281, N8276, N7282);
nor NOR3 (N8282, N8277, N4093, N3407);
not NOT1 (N8283, N8279);
and AND4 (N8284, N8261, N816, N3782, N3420);
or OR3 (N8285, N8264, N2565, N5713);
xor XOR2 (N8286, N8284, N8210);
nor NOR3 (N8287, N8280, N5973, N5016);
not NOT1 (N8288, N8283);
nor NOR3 (N8289, N8287, N3901, N5522);
nor NOR4 (N8290, N8289, N5698, N3436, N1973);
nor NOR4 (N8291, N8290, N7969, N7603, N2707);
nand NAND3 (N8292, N8282, N6488, N1331);
nor NOR2 (N8293, N8292, N7234);
nand NAND3 (N8294, N8281, N4423, N7412);
and AND3 (N8295, N8286, N191, N7690);
nand NAND4 (N8296, N8291, N7030, N4241, N2596);
and AND3 (N8297, N8269, N5629, N1258);
or OR3 (N8298, N8285, N4778, N2578);
not NOT1 (N8299, N8294);
nor NOR4 (N8300, N8297, N8018, N3428, N4200);
nor NOR4 (N8301, N8278, N2775, N6427, N1627);
and AND2 (N8302, N8295, N6054);
nand NAND2 (N8303, N8302, N5920);
xor XOR2 (N8304, N8272, N8041);
or OR4 (N8305, N8299, N4994, N923, N7393);
or OR2 (N8306, N8293, N1014);
not NOT1 (N8307, N8303);
not NOT1 (N8308, N8301);
nor NOR2 (N8309, N8298, N8202);
buf BUF1 (N8310, N8308);
buf BUF1 (N8311, N8307);
and AND2 (N8312, N8300, N3667);
and AND4 (N8313, N8311, N590, N1318, N2033);
xor XOR2 (N8314, N8275, N3872);
buf BUF1 (N8315, N8313);
or OR2 (N8316, N8288, N8270);
nor NOR2 (N8317, N8316, N1250);
or OR3 (N8318, N8315, N6484, N5485);
and AND4 (N8319, N8310, N4740, N1542, N393);
buf BUF1 (N8320, N8319);
nor NOR3 (N8321, N8312, N1993, N5328);
xor XOR2 (N8322, N8320, N7029);
xor XOR2 (N8323, N8296, N2113);
nor NOR2 (N8324, N8317, N906);
nand NAND4 (N8325, N8318, N4477, N1894, N723);
nand NAND3 (N8326, N8306, N3578, N4653);
nor NOR3 (N8327, N8325, N974, N5172);
buf BUF1 (N8328, N8323);
nand NAND2 (N8329, N8321, N6920);
nand NAND3 (N8330, N8322, N1433, N2766);
not NOT1 (N8331, N8326);
not NOT1 (N8332, N8329);
or OR4 (N8333, N8328, N5684, N4516, N7456);
xor XOR2 (N8334, N8330, N2281);
xor XOR2 (N8335, N8309, N816);
or OR2 (N8336, N8305, N3010);
or OR2 (N8337, N8336, N1360);
or OR3 (N8338, N8314, N2852, N5883);
nor NOR3 (N8339, N8335, N4071, N6543);
or OR4 (N8340, N8332, N464, N354, N7035);
buf BUF1 (N8341, N8339);
not NOT1 (N8342, N8340);
xor XOR2 (N8343, N8333, N4224);
xor XOR2 (N8344, N8341, N798);
buf BUF1 (N8345, N8334);
not NOT1 (N8346, N8344);
nand NAND3 (N8347, N8346, N1442, N7285);
not NOT1 (N8348, N8337);
nand NAND4 (N8349, N8345, N4591, N1740, N6363);
not NOT1 (N8350, N8347);
and AND3 (N8351, N8327, N5219, N3411);
and AND3 (N8352, N8351, N249, N1020);
not NOT1 (N8353, N8304);
xor XOR2 (N8354, N8324, N7827);
buf BUF1 (N8355, N8350);
and AND2 (N8356, N8331, N7108);
nand NAND2 (N8357, N8355, N4978);
nand NAND3 (N8358, N8342, N5410, N5230);
nor NOR2 (N8359, N8349, N1758);
buf BUF1 (N8360, N8356);
xor XOR2 (N8361, N8352, N2606);
not NOT1 (N8362, N8359);
not NOT1 (N8363, N8358);
and AND4 (N8364, N8360, N3203, N6417, N262);
xor XOR2 (N8365, N8354, N5455);
xor XOR2 (N8366, N8348, N1774);
not NOT1 (N8367, N8363);
and AND4 (N8368, N8353, N7559, N6305, N5418);
xor XOR2 (N8369, N8362, N4917);
not NOT1 (N8370, N8364);
nand NAND2 (N8371, N8370, N1080);
or OR3 (N8372, N8369, N3847, N1710);
not NOT1 (N8373, N8338);
xor XOR2 (N8374, N8357, N5893);
xor XOR2 (N8375, N8373, N3612);
and AND3 (N8376, N8365, N1934, N6188);
nor NOR2 (N8377, N8375, N7875);
xor XOR2 (N8378, N8366, N5815);
not NOT1 (N8379, N8372);
not NOT1 (N8380, N8378);
and AND4 (N8381, N8376, N1729, N2684, N7349);
nor NOR3 (N8382, N8377, N5768, N6993);
not NOT1 (N8383, N8367);
not NOT1 (N8384, N8381);
buf BUF1 (N8385, N8383);
nor NOR2 (N8386, N8379, N4412);
not NOT1 (N8387, N8374);
xor XOR2 (N8388, N8361, N4064);
buf BUF1 (N8389, N8385);
buf BUF1 (N8390, N8382);
not NOT1 (N8391, N8387);
xor XOR2 (N8392, N8371, N1305);
not NOT1 (N8393, N8390);
xor XOR2 (N8394, N8380, N3154);
or OR2 (N8395, N8388, N7538);
and AND2 (N8396, N8389, N5214);
nor NOR2 (N8397, N8393, N2048);
buf BUF1 (N8398, N8384);
nand NAND2 (N8399, N8395, N6937);
nand NAND2 (N8400, N8368, N1488);
nand NAND2 (N8401, N8392, N4258);
xor XOR2 (N8402, N8398, N3234);
nand NAND4 (N8403, N8394, N2163, N7800, N3945);
buf BUF1 (N8404, N8403);
or OR4 (N8405, N8391, N7903, N3421, N157);
xor XOR2 (N8406, N8343, N2829);
buf BUF1 (N8407, N8401);
or OR2 (N8408, N8404, N8205);
nand NAND3 (N8409, N8397, N4929, N5615);
or OR3 (N8410, N8406, N1756, N7423);
nor NOR2 (N8411, N8409, N3390);
buf BUF1 (N8412, N8396);
nor NOR3 (N8413, N8402, N7438, N4689);
xor XOR2 (N8414, N8413, N5013);
nand NAND2 (N8415, N8412, N8256);
xor XOR2 (N8416, N8405, N4400);
nand NAND4 (N8417, N8407, N2034, N6515, N3461);
not NOT1 (N8418, N8410);
and AND3 (N8419, N8386, N2843, N3146);
nand NAND3 (N8420, N8416, N3005, N5820);
nor NOR4 (N8421, N8420, N3017, N2101, N7564);
and AND3 (N8422, N8414, N119, N2030);
xor XOR2 (N8423, N8411, N3370);
not NOT1 (N8424, N8417);
nor NOR2 (N8425, N8419, N7711);
not NOT1 (N8426, N8399);
buf BUF1 (N8427, N8426);
not NOT1 (N8428, N8421);
nor NOR3 (N8429, N8400, N2895, N2605);
not NOT1 (N8430, N8423);
or OR2 (N8431, N8422, N7506);
buf BUF1 (N8432, N8424);
or OR2 (N8433, N8429, N4544);
not NOT1 (N8434, N8430);
buf BUF1 (N8435, N8428);
xor XOR2 (N8436, N8435, N4793);
xor XOR2 (N8437, N8431, N2239);
or OR3 (N8438, N8427, N84, N3083);
nand NAND4 (N8439, N8408, N2075, N6913, N8237);
xor XOR2 (N8440, N8434, N2271);
nor NOR3 (N8441, N8425, N3911, N7071);
buf BUF1 (N8442, N8438);
nor NOR4 (N8443, N8442, N5580, N1381, N4128);
nand NAND3 (N8444, N8433, N5537, N516);
xor XOR2 (N8445, N8439, N8189);
or OR4 (N8446, N8441, N6679, N1200, N7802);
nor NOR4 (N8447, N8440, N4593, N6633, N7546);
xor XOR2 (N8448, N8437, N1606);
nand NAND4 (N8449, N8415, N8128, N8043, N1162);
not NOT1 (N8450, N8444);
nand NAND3 (N8451, N8443, N5317, N7931);
or OR3 (N8452, N8418, N5291, N3977);
buf BUF1 (N8453, N8436);
and AND3 (N8454, N8432, N1720, N1191);
or OR4 (N8455, N8454, N3342, N8427, N4031);
buf BUF1 (N8456, N8445);
buf BUF1 (N8457, N8448);
nand NAND3 (N8458, N8449, N7715, N6446);
xor XOR2 (N8459, N8446, N6695);
xor XOR2 (N8460, N8452, N5623);
not NOT1 (N8461, N8459);
buf BUF1 (N8462, N8456);
and AND2 (N8463, N8455, N3912);
not NOT1 (N8464, N8462);
xor XOR2 (N8465, N8447, N2209);
not NOT1 (N8466, N8460);
nor NOR4 (N8467, N8451, N5547, N7699, N7498);
or OR3 (N8468, N8450, N1138, N2263);
not NOT1 (N8469, N8465);
nor NOR2 (N8470, N8469, N3861);
xor XOR2 (N8471, N8463, N4013);
buf BUF1 (N8472, N8467);
nand NAND4 (N8473, N8461, N787, N4631, N5354);
nor NOR4 (N8474, N8453, N781, N4544, N4739);
nand NAND3 (N8475, N8471, N1106, N3584);
xor XOR2 (N8476, N8466, N6125);
nand NAND4 (N8477, N8470, N1191, N5199, N3303);
not NOT1 (N8478, N8477);
nand NAND3 (N8479, N8474, N1632, N1514);
and AND2 (N8480, N8464, N3649);
and AND2 (N8481, N8458, N7985);
or OR2 (N8482, N8473, N5257);
not NOT1 (N8483, N8468);
not NOT1 (N8484, N8478);
nand NAND3 (N8485, N8457, N1084, N4443);
nor NOR4 (N8486, N8482, N1035, N5653, N1959);
nand NAND4 (N8487, N8485, N7443, N2521, N7329);
and AND3 (N8488, N8480, N8451, N4360);
not NOT1 (N8489, N8486);
nand NAND3 (N8490, N8483, N652, N463);
xor XOR2 (N8491, N8490, N6507);
buf BUF1 (N8492, N8472);
nor NOR4 (N8493, N8484, N5826, N8003, N5068);
buf BUF1 (N8494, N8479);
buf BUF1 (N8495, N8488);
buf BUF1 (N8496, N8481);
not NOT1 (N8497, N8489);
buf BUF1 (N8498, N8495);
nor NOR3 (N8499, N8496, N1371, N6059);
nor NOR2 (N8500, N8475, N5780);
and AND4 (N8501, N8492, N6900, N476, N2003);
or OR2 (N8502, N8501, N5164);
and AND3 (N8503, N8476, N1628, N3803);
nand NAND2 (N8504, N8503, N4753);
not NOT1 (N8505, N8502);
not NOT1 (N8506, N8497);
or OR2 (N8507, N8498, N7885);
and AND2 (N8508, N8491, N3820);
or OR4 (N8509, N8506, N745, N2356, N7937);
xor XOR2 (N8510, N8508, N2496);
or OR2 (N8511, N8509, N6608);
nor NOR4 (N8512, N8494, N1719, N503, N3696);
and AND3 (N8513, N8487, N4097, N1855);
not NOT1 (N8514, N8513);
nor NOR3 (N8515, N8505, N5325, N4164);
and AND2 (N8516, N8493, N4098);
nand NAND4 (N8517, N8507, N695, N3058, N7125);
or OR3 (N8518, N8499, N7542, N3430);
xor XOR2 (N8519, N8504, N818);
nand NAND2 (N8520, N8512, N6397);
buf BUF1 (N8521, N8514);
buf BUF1 (N8522, N8500);
or OR4 (N8523, N8510, N604, N7746, N7473);
nor NOR4 (N8524, N8515, N7191, N7031, N5826);
and AND3 (N8525, N8511, N2709, N6241);
not NOT1 (N8526, N8520);
buf BUF1 (N8527, N8526);
nor NOR3 (N8528, N8521, N8327, N3838);
buf BUF1 (N8529, N8525);
nor NOR2 (N8530, N8529, N6770);
nand NAND2 (N8531, N8524, N4550);
not NOT1 (N8532, N8528);
not NOT1 (N8533, N8532);
xor XOR2 (N8534, N8533, N247);
nor NOR2 (N8535, N8518, N841);
buf BUF1 (N8536, N8527);
nand NAND4 (N8537, N8519, N6174, N5016, N7101);
nand NAND4 (N8538, N8537, N635, N2486, N6323);
nand NAND3 (N8539, N8523, N7756, N3536);
or OR4 (N8540, N8516, N1999, N2183, N6499);
or OR3 (N8541, N8522, N6966, N141);
xor XOR2 (N8542, N8539, N5013);
nor NOR2 (N8543, N8531, N1801);
or OR2 (N8544, N8540, N6363);
not NOT1 (N8545, N8517);
nand NAND4 (N8546, N8541, N6782, N5704, N4441);
nor NOR3 (N8547, N8530, N4418, N7794);
nand NAND2 (N8548, N8538, N6503);
or OR4 (N8549, N8542, N7107, N5076, N3836);
nor NOR3 (N8550, N8549, N7982, N2339);
nor NOR3 (N8551, N8536, N3485, N4193);
and AND3 (N8552, N8547, N3702, N4525);
nor NOR4 (N8553, N8550, N2001, N5897, N212);
nor NOR4 (N8554, N8545, N1410, N6894, N4095);
buf BUF1 (N8555, N8544);
or OR3 (N8556, N8552, N5245, N6196);
nand NAND4 (N8557, N8556, N2284, N5397, N8213);
buf BUF1 (N8558, N8555);
and AND4 (N8559, N8546, N3426, N7656, N4435);
and AND4 (N8560, N8559, N7262, N2302, N6637);
and AND4 (N8561, N8534, N6405, N6823, N7296);
or OR3 (N8562, N8543, N6198, N7734);
nand NAND3 (N8563, N8554, N3518, N3932);
not NOT1 (N8564, N8548);
or OR2 (N8565, N8561, N6260);
nand NAND2 (N8566, N8553, N5126);
nor NOR3 (N8567, N8560, N7361, N7529);
nand NAND3 (N8568, N8558, N1925, N17);
xor XOR2 (N8569, N8568, N900);
nand NAND4 (N8570, N8563, N2192, N6555, N6915);
nor NOR2 (N8571, N8562, N6376);
and AND4 (N8572, N8571, N1551, N6264, N1579);
or OR3 (N8573, N8557, N7159, N5373);
nor NOR3 (N8574, N8573, N4657, N6248);
or OR4 (N8575, N8551, N7285, N579, N7021);
nor NOR4 (N8576, N8574, N7468, N7594, N4494);
or OR2 (N8577, N8566, N2951);
nand NAND2 (N8578, N8569, N1855);
buf BUF1 (N8579, N8572);
nand NAND3 (N8580, N8565, N1685, N983);
and AND3 (N8581, N8576, N7102, N457);
or OR2 (N8582, N8580, N7998);
and AND3 (N8583, N8564, N2966, N7053);
xor XOR2 (N8584, N8581, N1841);
not NOT1 (N8585, N8579);
nor NOR4 (N8586, N8578, N5262, N149, N7989);
or OR2 (N8587, N8577, N7785);
buf BUF1 (N8588, N8584);
xor XOR2 (N8589, N8587, N6283);
not NOT1 (N8590, N8585);
buf BUF1 (N8591, N8588);
and AND3 (N8592, N8575, N7519, N7901);
buf BUF1 (N8593, N8590);
and AND3 (N8594, N8592, N5976, N7135);
nand NAND4 (N8595, N8583, N7042, N2375, N7484);
xor XOR2 (N8596, N8591, N7617);
not NOT1 (N8597, N8567);
nor NOR3 (N8598, N8596, N1240, N1551);
buf BUF1 (N8599, N8582);
nor NOR2 (N8600, N8597, N668);
nor NOR3 (N8601, N8570, N5749, N2832);
buf BUF1 (N8602, N8589);
nor NOR3 (N8603, N8595, N482, N4966);
and AND4 (N8604, N8602, N4266, N3649, N2684);
nor NOR3 (N8605, N8586, N7995, N1016);
nor NOR2 (N8606, N8603, N3694);
or OR4 (N8607, N8604, N3998, N4755, N5154);
not NOT1 (N8608, N8605);
nand NAND3 (N8609, N8608, N4318, N1795);
not NOT1 (N8610, N8598);
and AND3 (N8611, N8610, N6980, N845);
nor NOR2 (N8612, N8594, N3877);
not NOT1 (N8613, N8600);
or OR2 (N8614, N8609, N2941);
not NOT1 (N8615, N8606);
not NOT1 (N8616, N8612);
buf BUF1 (N8617, N8599);
nand NAND2 (N8618, N8535, N5689);
xor XOR2 (N8619, N8607, N2847);
xor XOR2 (N8620, N8615, N4763);
xor XOR2 (N8621, N8616, N7821);
buf BUF1 (N8622, N8613);
and AND4 (N8623, N8617, N2234, N6309, N2487);
buf BUF1 (N8624, N8601);
xor XOR2 (N8625, N8593, N6614);
nor NOR2 (N8626, N8624, N2431);
nand NAND3 (N8627, N8621, N3229, N2247);
xor XOR2 (N8628, N8619, N4892);
and AND3 (N8629, N8614, N6170, N403);
or OR2 (N8630, N8623, N6821);
and AND4 (N8631, N8625, N1888, N7494, N6655);
buf BUF1 (N8632, N8618);
nand NAND2 (N8633, N8622, N5055);
nand NAND4 (N8634, N8627, N5002, N2438, N2903);
buf BUF1 (N8635, N8611);
and AND3 (N8636, N8620, N8404, N1767);
nor NOR4 (N8637, N8636, N2161, N187, N121);
nand NAND3 (N8638, N8637, N557, N3234);
not NOT1 (N8639, N8629);
xor XOR2 (N8640, N8632, N249);
and AND3 (N8641, N8633, N5631, N7935);
and AND3 (N8642, N8630, N5385, N7099);
nor NOR4 (N8643, N8641, N2362, N2531, N4016);
xor XOR2 (N8644, N8638, N4032);
nor NOR2 (N8645, N8639, N6834);
buf BUF1 (N8646, N8626);
buf BUF1 (N8647, N8635);
buf BUF1 (N8648, N8646);
nand NAND4 (N8649, N8647, N1868, N4656, N4285);
or OR2 (N8650, N8643, N4034);
xor XOR2 (N8651, N8640, N282);
nand NAND3 (N8652, N8628, N2646, N7270);
and AND3 (N8653, N8650, N3690, N8476);
nand NAND4 (N8654, N8645, N7830, N7907, N6443);
nand NAND4 (N8655, N8648, N6307, N6651, N2851);
xor XOR2 (N8656, N8653, N2760);
nor NOR3 (N8657, N8642, N5318, N6401);
nand NAND4 (N8658, N8631, N5719, N8433, N4478);
buf BUF1 (N8659, N8652);
xor XOR2 (N8660, N8634, N6791);
nand NAND2 (N8661, N8657, N4389);
and AND4 (N8662, N8654, N792, N5678, N6210);
not NOT1 (N8663, N8660);
buf BUF1 (N8664, N8658);
or OR2 (N8665, N8656, N4144);
xor XOR2 (N8666, N8663, N4948);
not NOT1 (N8667, N8664);
buf BUF1 (N8668, N8666);
nor NOR3 (N8669, N8667, N5637, N1687);
nor NOR4 (N8670, N8662, N2097, N8294, N6238);
buf BUF1 (N8671, N8644);
nand NAND2 (N8672, N8655, N7980);
or OR3 (N8673, N8659, N4564, N8549);
and AND3 (N8674, N8665, N2042, N7794);
buf BUF1 (N8675, N8668);
or OR2 (N8676, N8674, N4636);
xor XOR2 (N8677, N8670, N4452);
not NOT1 (N8678, N8649);
not NOT1 (N8679, N8661);
nand NAND4 (N8680, N8651, N3502, N4091, N4256);
or OR2 (N8681, N8671, N2895);
nand NAND4 (N8682, N8675, N6922, N1000, N4854);
not NOT1 (N8683, N8679);
and AND4 (N8684, N8677, N3324, N2079, N3846);
xor XOR2 (N8685, N8682, N301);
xor XOR2 (N8686, N8678, N5813);
buf BUF1 (N8687, N8669);
and AND3 (N8688, N8687, N8239, N2696);
buf BUF1 (N8689, N8685);
and AND2 (N8690, N8688, N4747);
and AND4 (N8691, N8684, N5955, N6618, N5168);
nand NAND2 (N8692, N8672, N6457);
or OR4 (N8693, N8689, N8557, N4758, N5252);
nand NAND2 (N8694, N8691, N1469);
and AND2 (N8695, N8692, N7158);
buf BUF1 (N8696, N8693);
xor XOR2 (N8697, N8681, N6753);
nand NAND3 (N8698, N8695, N6146, N6241);
not NOT1 (N8699, N8694);
xor XOR2 (N8700, N8686, N1828);
buf BUF1 (N8701, N8680);
xor XOR2 (N8702, N8696, N4176);
nor NOR3 (N8703, N8673, N591, N2876);
not NOT1 (N8704, N8698);
nor NOR2 (N8705, N8676, N2279);
xor XOR2 (N8706, N8704, N7271);
not NOT1 (N8707, N8699);
nor NOR4 (N8708, N8683, N5546, N6150, N3163);
or OR3 (N8709, N8697, N7745, N4881);
nand NAND4 (N8710, N8702, N2866, N3834, N3430);
not NOT1 (N8711, N8707);
xor XOR2 (N8712, N8710, N4613);
and AND4 (N8713, N8709, N1599, N5458, N611);
xor XOR2 (N8714, N8712, N7539);
nor NOR4 (N8715, N8708, N5471, N5002, N4967);
nor NOR3 (N8716, N8713, N5272, N6884);
xor XOR2 (N8717, N8706, N3578);
buf BUF1 (N8718, N8715);
buf BUF1 (N8719, N8717);
nor NOR2 (N8720, N8716, N4763);
xor XOR2 (N8721, N8711, N4955);
nor NOR3 (N8722, N8701, N1083, N3942);
buf BUF1 (N8723, N8718);
nor NOR4 (N8724, N8714, N1626, N1270, N4722);
nand NAND3 (N8725, N8705, N6053, N8021);
xor XOR2 (N8726, N8724, N8358);
not NOT1 (N8727, N8700);
nand NAND4 (N8728, N8726, N1151, N4485, N750);
nand NAND2 (N8729, N8722, N3272);
or OR2 (N8730, N8719, N1313);
not NOT1 (N8731, N8727);
nand NAND3 (N8732, N8725, N7841, N2666);
nand NAND3 (N8733, N8732, N8354, N7569);
nor NOR4 (N8734, N8728, N5027, N7513, N5956);
and AND3 (N8735, N8721, N7882, N2640);
nand NAND4 (N8736, N8730, N636, N5265, N216);
buf BUF1 (N8737, N8733);
or OR2 (N8738, N8736, N3447);
or OR3 (N8739, N8735, N2981, N801);
not NOT1 (N8740, N8734);
xor XOR2 (N8741, N8739, N3890);
buf BUF1 (N8742, N8737);
or OR2 (N8743, N8742, N2502);
xor XOR2 (N8744, N8738, N6159);
nand NAND2 (N8745, N8690, N3320);
nand NAND2 (N8746, N8729, N7647);
and AND3 (N8747, N8720, N1128, N8677);
and AND4 (N8748, N8747, N5621, N912, N5399);
and AND2 (N8749, N8731, N8724);
nor NOR3 (N8750, N8744, N8728, N2999);
nor NOR4 (N8751, N8750, N8625, N8351, N6711);
nand NAND2 (N8752, N8703, N3230);
buf BUF1 (N8753, N8749);
and AND3 (N8754, N8746, N7676, N2337);
xor XOR2 (N8755, N8748, N1341);
buf BUF1 (N8756, N8741);
and AND4 (N8757, N8754, N5917, N3692, N3001);
or OR2 (N8758, N8756, N136);
not NOT1 (N8759, N8740);
buf BUF1 (N8760, N8752);
xor XOR2 (N8761, N8755, N3365);
xor XOR2 (N8762, N8753, N122);
and AND4 (N8763, N8751, N2721, N6852, N4634);
and AND4 (N8764, N8761, N3342, N5134, N6876);
xor XOR2 (N8765, N8723, N8475);
not NOT1 (N8766, N8745);
and AND2 (N8767, N8757, N3337);
nor NOR4 (N8768, N8760, N6027, N8447, N7058);
and AND3 (N8769, N8743, N592, N2521);
nand NAND4 (N8770, N8758, N6756, N6760, N3609);
buf BUF1 (N8771, N8762);
nand NAND2 (N8772, N8765, N7090);
nand NAND4 (N8773, N8768, N6520, N684, N4648);
nand NAND3 (N8774, N8764, N526, N6486);
not NOT1 (N8775, N8766);
or OR2 (N8776, N8775, N6458);
xor XOR2 (N8777, N8771, N1969);
or OR3 (N8778, N8767, N140, N4532);
buf BUF1 (N8779, N8763);
nor NOR4 (N8780, N8759, N5673, N3691, N6967);
nor NOR2 (N8781, N8770, N2216);
or OR4 (N8782, N8779, N6140, N1046, N6532);
or OR4 (N8783, N8769, N139, N2964, N8729);
not NOT1 (N8784, N8781);
and AND3 (N8785, N8776, N941, N97);
not NOT1 (N8786, N8780);
nand NAND3 (N8787, N8785, N826, N5089);
nand NAND2 (N8788, N8778, N4777);
nand NAND4 (N8789, N8774, N4789, N6445, N5553);
nor NOR4 (N8790, N8782, N6844, N3600, N2915);
nor NOR4 (N8791, N8772, N4407, N7116, N4650);
nand NAND3 (N8792, N8786, N314, N3707);
xor XOR2 (N8793, N8789, N5967);
nor NOR3 (N8794, N8787, N2934, N6995);
buf BUF1 (N8795, N8793);
or OR2 (N8796, N8790, N7617);
nand NAND3 (N8797, N8773, N1285, N2796);
or OR3 (N8798, N8783, N5965, N3153);
or OR4 (N8799, N8792, N909, N5922, N5231);
buf BUF1 (N8800, N8798);
nor NOR4 (N8801, N8791, N5844, N2852, N5917);
and AND2 (N8802, N8796, N1614);
nor NOR3 (N8803, N8777, N7040, N6789);
xor XOR2 (N8804, N8794, N6032);
xor XOR2 (N8805, N8795, N6884);
buf BUF1 (N8806, N8800);
not NOT1 (N8807, N8802);
not NOT1 (N8808, N8797);
xor XOR2 (N8809, N8806, N4233);
xor XOR2 (N8810, N8788, N1416);
not NOT1 (N8811, N8809);
nor NOR4 (N8812, N8801, N4311, N2582, N7485);
and AND3 (N8813, N8804, N6889, N8655);
or OR3 (N8814, N8810, N5273, N5106);
and AND3 (N8815, N8803, N601, N5652);
or OR4 (N8816, N8812, N5515, N3514, N3810);
xor XOR2 (N8817, N8816, N8412);
buf BUF1 (N8818, N8807);
and AND3 (N8819, N8813, N1283, N5952);
nand NAND2 (N8820, N8819, N8333);
nand NAND4 (N8821, N8784, N7090, N1500, N2468);
not NOT1 (N8822, N8811);
xor XOR2 (N8823, N8805, N8184);
buf BUF1 (N8824, N8815);
buf BUF1 (N8825, N8821);
nand NAND2 (N8826, N8818, N5570);
nor NOR2 (N8827, N8825, N1179);
nor NOR4 (N8828, N8822, N2560, N3261, N11);
and AND3 (N8829, N8799, N2890, N7717);
and AND3 (N8830, N8828, N7269, N6600);
not NOT1 (N8831, N8814);
nor NOR4 (N8832, N8823, N1863, N1212, N5792);
nor NOR4 (N8833, N8824, N7109, N4078, N8460);
xor XOR2 (N8834, N8832, N6141);
or OR3 (N8835, N8829, N8635, N2964);
or OR3 (N8836, N8817, N6792, N6145);
and AND2 (N8837, N8820, N7325);
not NOT1 (N8838, N8808);
or OR3 (N8839, N8833, N6863, N3731);
and AND3 (N8840, N8830, N802, N1036);
or OR4 (N8841, N8837, N6937, N1642, N6557);
nand NAND2 (N8842, N8826, N7653);
buf BUF1 (N8843, N8841);
nor NOR2 (N8844, N8836, N1662);
and AND4 (N8845, N8827, N4815, N2501, N8224);
not NOT1 (N8846, N8840);
not NOT1 (N8847, N8845);
buf BUF1 (N8848, N8847);
nor NOR2 (N8849, N8835, N8154);
and AND2 (N8850, N8844, N1935);
and AND2 (N8851, N8848, N3904);
xor XOR2 (N8852, N8843, N5358);
or OR4 (N8853, N8846, N2258, N4107, N5793);
and AND4 (N8854, N8834, N3203, N2689, N356);
and AND4 (N8855, N8831, N8080, N2502, N4121);
nand NAND3 (N8856, N8853, N4868, N2641);
nand NAND2 (N8857, N8856, N300);
nand NAND3 (N8858, N8851, N1221, N8183);
xor XOR2 (N8859, N8852, N4238);
and AND3 (N8860, N8854, N4293, N7878);
not NOT1 (N8861, N8859);
not NOT1 (N8862, N8850);
buf BUF1 (N8863, N8839);
nor NOR3 (N8864, N8842, N3035, N3309);
not NOT1 (N8865, N8855);
and AND3 (N8866, N8860, N6947, N850);
nand NAND3 (N8867, N8864, N5503, N7154);
buf BUF1 (N8868, N8866);
and AND2 (N8869, N8867, N8181);
or OR3 (N8870, N8858, N8816, N8588);
and AND3 (N8871, N8861, N7488, N3834);
xor XOR2 (N8872, N8865, N59);
not NOT1 (N8873, N8863);
xor XOR2 (N8874, N8849, N4121);
xor XOR2 (N8875, N8838, N7551);
xor XOR2 (N8876, N8869, N2171);
and AND4 (N8877, N8870, N8783, N4950, N6279);
buf BUF1 (N8878, N8857);
not NOT1 (N8879, N8878);
buf BUF1 (N8880, N8879);
nand NAND2 (N8881, N8862, N4856);
nor NOR4 (N8882, N8873, N7094, N6564, N4923);
xor XOR2 (N8883, N8874, N2368);
buf BUF1 (N8884, N8871);
not NOT1 (N8885, N8868);
not NOT1 (N8886, N8885);
nand NAND4 (N8887, N8877, N6624, N4212, N6581);
xor XOR2 (N8888, N8880, N7327);
xor XOR2 (N8889, N8888, N6773);
nor NOR3 (N8890, N8886, N3446, N3346);
buf BUF1 (N8891, N8875);
and AND3 (N8892, N8884, N7880, N7376);
xor XOR2 (N8893, N8891, N4376);
and AND4 (N8894, N8882, N3633, N4428, N6883);
not NOT1 (N8895, N8889);
xor XOR2 (N8896, N8895, N1246);
buf BUF1 (N8897, N8890);
xor XOR2 (N8898, N8876, N7236);
not NOT1 (N8899, N8883);
or OR2 (N8900, N8898, N268);
or OR3 (N8901, N8897, N1602, N5172);
buf BUF1 (N8902, N8893);
and AND4 (N8903, N8901, N7057, N3905, N7412);
not NOT1 (N8904, N8887);
nand NAND2 (N8905, N8900, N7401);
or OR2 (N8906, N8903, N1063);
and AND2 (N8907, N8905, N4656);
nand NAND4 (N8908, N8881, N4178, N7567, N79);
not NOT1 (N8909, N8872);
nand NAND2 (N8910, N8896, N8885);
nand NAND4 (N8911, N8909, N4684, N7569, N3618);
or OR4 (N8912, N8892, N6972, N4814, N8448);
xor XOR2 (N8913, N8894, N712);
not NOT1 (N8914, N8899);
nor NOR4 (N8915, N8913, N4170, N5580, N7866);
not NOT1 (N8916, N8915);
buf BUF1 (N8917, N8911);
xor XOR2 (N8918, N8916, N2968);
xor XOR2 (N8919, N8918, N7418);
xor XOR2 (N8920, N8907, N7219);
nand NAND2 (N8921, N8917, N773);
not NOT1 (N8922, N8920);
nand NAND4 (N8923, N8904, N1003, N1072, N5120);
nand NAND2 (N8924, N8921, N1534);
or OR3 (N8925, N8912, N1063, N4914);
buf BUF1 (N8926, N8919);
nand NAND4 (N8927, N8908, N4646, N2157, N10);
not NOT1 (N8928, N8910);
or OR2 (N8929, N8923, N3127);
nor NOR3 (N8930, N8929, N4447, N3214);
nand NAND3 (N8931, N8925, N6175, N589);
and AND2 (N8932, N8927, N8666);
or OR3 (N8933, N8924, N8590, N4271);
not NOT1 (N8934, N8914);
not NOT1 (N8935, N8931);
nand NAND3 (N8936, N8902, N505, N2454);
nand NAND2 (N8937, N8932, N44);
or OR2 (N8938, N8934, N5172);
nor NOR2 (N8939, N8926, N3711);
not NOT1 (N8940, N8922);
buf BUF1 (N8941, N8937);
xor XOR2 (N8942, N8939, N565);
nand NAND3 (N8943, N8940, N2616, N6896);
buf BUF1 (N8944, N8930);
and AND3 (N8945, N8933, N1585, N194);
or OR3 (N8946, N8941, N2498, N380);
nor NOR2 (N8947, N8938, N6021);
nand NAND4 (N8948, N8946, N6941, N548, N3818);
buf BUF1 (N8949, N8942);
and AND3 (N8950, N8943, N4700, N3728);
buf BUF1 (N8951, N8950);
nor NOR4 (N8952, N8948, N4156, N1270, N4551);
xor XOR2 (N8953, N8947, N1187);
not NOT1 (N8954, N8952);
nor NOR3 (N8955, N8928, N3298, N5765);
buf BUF1 (N8956, N8954);
or OR4 (N8957, N8956, N7066, N3633, N5509);
nand NAND3 (N8958, N8951, N6824, N7709);
nand NAND2 (N8959, N8955, N7190);
nor NOR4 (N8960, N8936, N1253, N157, N4525);
or OR3 (N8961, N8945, N3902, N4535);
not NOT1 (N8962, N8960);
and AND3 (N8963, N8958, N3984, N7596);
buf BUF1 (N8964, N8906);
nor NOR3 (N8965, N8963, N5539, N629);
and AND2 (N8966, N8964, N5058);
and AND3 (N8967, N8959, N1366, N3823);
not NOT1 (N8968, N8965);
and AND4 (N8969, N8935, N2027, N7600, N6030);
nand NAND3 (N8970, N8957, N1644, N3645);
nor NOR3 (N8971, N8967, N2005, N3808);
nor NOR3 (N8972, N8966, N1695, N4038);
or OR2 (N8973, N8969, N7904);
not NOT1 (N8974, N8970);
nand NAND2 (N8975, N8968, N2468);
or OR4 (N8976, N8972, N270, N1386, N6666);
and AND4 (N8977, N8949, N1721, N2456, N1891);
nor NOR2 (N8978, N8944, N7759);
or OR4 (N8979, N8953, N3965, N1447, N4284);
and AND3 (N8980, N8971, N4034, N4159);
or OR3 (N8981, N8962, N600, N8039);
or OR2 (N8982, N8980, N5768);
not NOT1 (N8983, N8978);
and AND3 (N8984, N8961, N6267, N8586);
buf BUF1 (N8985, N8974);
xor XOR2 (N8986, N8973, N8479);
xor XOR2 (N8987, N8982, N8263);
not NOT1 (N8988, N8985);
nor NOR4 (N8989, N8984, N5116, N306, N8806);
buf BUF1 (N8990, N8976);
xor XOR2 (N8991, N8975, N5847);
and AND3 (N8992, N8983, N3760, N3319);
or OR3 (N8993, N8989, N3648, N647);
buf BUF1 (N8994, N8979);
or OR4 (N8995, N8987, N1933, N8415, N7606);
and AND3 (N8996, N8994, N1966, N8690);
or OR4 (N8997, N8996, N3480, N8972, N5369);
or OR2 (N8998, N8995, N666);
buf BUF1 (N8999, N8998);
buf BUF1 (N9000, N8991);
xor XOR2 (N9001, N8993, N5996);
nor NOR2 (N9002, N8992, N946);
xor XOR2 (N9003, N9001, N3825);
or OR3 (N9004, N8977, N8924, N7135);
nand NAND3 (N9005, N8997, N7425, N5528);
nand NAND4 (N9006, N9004, N5888, N8048, N4544);
or OR3 (N9007, N8981, N4756, N4345);
nand NAND3 (N9008, N8986, N3053, N8110);
nor NOR4 (N9009, N9006, N8755, N924, N4807);
or OR2 (N9010, N9008, N7448);
buf BUF1 (N9011, N8988);
and AND4 (N9012, N9002, N6381, N8482, N1860);
not NOT1 (N9013, N9010);
or OR3 (N9014, N9007, N7102, N5828);
and AND3 (N9015, N8999, N4529, N2444);
not NOT1 (N9016, N9005);
xor XOR2 (N9017, N9000, N1497);
nand NAND2 (N9018, N9009, N6092);
and AND2 (N9019, N9017, N3905);
nand NAND3 (N9020, N9018, N2539, N7532);
not NOT1 (N9021, N9011);
not NOT1 (N9022, N9012);
nand NAND4 (N9023, N8990, N5079, N8811, N5016);
buf BUF1 (N9024, N9021);
not NOT1 (N9025, N9014);
and AND4 (N9026, N9015, N2024, N4593, N6947);
nor NOR2 (N9027, N9026, N2944);
or OR2 (N9028, N9003, N503);
nor NOR3 (N9029, N9027, N8370, N4612);
xor XOR2 (N9030, N9023, N7523);
buf BUF1 (N9031, N9016);
not NOT1 (N9032, N9013);
xor XOR2 (N9033, N9029, N6236);
buf BUF1 (N9034, N9022);
xor XOR2 (N9035, N9031, N2396);
buf BUF1 (N9036, N9020);
xor XOR2 (N9037, N9024, N6589);
or OR4 (N9038, N9019, N1771, N7162, N8266);
buf BUF1 (N9039, N9032);
xor XOR2 (N9040, N9035, N2683);
nand NAND4 (N9041, N9038, N4899, N7468, N2441);
nand NAND2 (N9042, N9025, N6234);
buf BUF1 (N9043, N9034);
or OR4 (N9044, N9039, N1637, N477, N3109);
nand NAND3 (N9045, N9040, N4114, N8376);
xor XOR2 (N9046, N9037, N6374);
xor XOR2 (N9047, N9044, N731);
buf BUF1 (N9048, N9033);
xor XOR2 (N9049, N9046, N1158);
or OR2 (N9050, N9047, N8634);
and AND4 (N9051, N9042, N8266, N1498, N8547);
not NOT1 (N9052, N9036);
not NOT1 (N9053, N9045);
xor XOR2 (N9054, N9030, N7363);
xor XOR2 (N9055, N9043, N4853);
xor XOR2 (N9056, N9053, N404);
nand NAND3 (N9057, N9054, N294, N4354);
nand NAND4 (N9058, N9056, N8715, N7175, N157);
or OR2 (N9059, N9041, N8421);
nand NAND3 (N9060, N9028, N3716, N5713);
nor NOR2 (N9061, N9049, N2921);
and AND4 (N9062, N9059, N2421, N142, N363);
or OR4 (N9063, N9061, N1132, N5266, N1451);
nor NOR3 (N9064, N9057, N9017, N8978);
or OR3 (N9065, N9052, N7541, N5316);
nand NAND2 (N9066, N9060, N3622);
xor XOR2 (N9067, N9066, N3546);
and AND2 (N9068, N9050, N6197);
not NOT1 (N9069, N9048);
nand NAND2 (N9070, N9062, N3300);
nand NAND3 (N9071, N9068, N6577, N7124);
nor NOR4 (N9072, N9070, N3038, N5552, N2885);
xor XOR2 (N9073, N9067, N6001);
or OR2 (N9074, N9065, N1631);
not NOT1 (N9075, N9055);
and AND3 (N9076, N9074, N8406, N7064);
nor NOR2 (N9077, N9069, N6759);
and AND3 (N9078, N9064, N3526, N7827);
nand NAND2 (N9079, N9077, N5847);
nand NAND3 (N9080, N9075, N2519, N5845);
buf BUF1 (N9081, N9078);
and AND2 (N9082, N9051, N4510);
xor XOR2 (N9083, N9072, N3123);
nand NAND4 (N9084, N9079, N6745, N3105, N9074);
and AND2 (N9085, N9076, N966);
nand NAND2 (N9086, N9082, N3564);
buf BUF1 (N9087, N9086);
xor XOR2 (N9088, N9081, N6904);
not NOT1 (N9089, N9080);
or OR4 (N9090, N9058, N958, N4919, N3959);
xor XOR2 (N9091, N9090, N8824);
xor XOR2 (N9092, N9087, N4773);
xor XOR2 (N9093, N9091, N6743);
nor NOR4 (N9094, N9085, N1626, N3933, N8015);
and AND3 (N9095, N9083, N1851, N3623);
nand NAND4 (N9096, N9089, N4999, N4820, N5006);
not NOT1 (N9097, N9073);
not NOT1 (N9098, N9063);
or OR4 (N9099, N9094, N1900, N8432, N4083);
nand NAND2 (N9100, N9071, N2313);
xor XOR2 (N9101, N9098, N4831);
and AND2 (N9102, N9100, N8739);
not NOT1 (N9103, N9097);
and AND3 (N9104, N9101, N8936, N1355);
buf BUF1 (N9105, N9102);
and AND4 (N9106, N9105, N4362, N6240, N1183);
nor NOR3 (N9107, N9084, N6452, N3310);
xor XOR2 (N9108, N9096, N6300);
or OR4 (N9109, N9103, N8302, N3837, N6927);
or OR4 (N9110, N9108, N7306, N6604, N5154);
and AND3 (N9111, N9110, N1343, N1410);
nor NOR3 (N9112, N9092, N5799, N715);
or OR4 (N9113, N9106, N3452, N1177, N1906);
buf BUF1 (N9114, N9104);
and AND3 (N9115, N9095, N130, N2234);
not NOT1 (N9116, N9114);
nor NOR4 (N9117, N9113, N6704, N8672, N7370);
xor XOR2 (N9118, N9116, N4444);
buf BUF1 (N9119, N9112);
buf BUF1 (N9120, N9088);
nor NOR2 (N9121, N9119, N5666);
not NOT1 (N9122, N9120);
nand NAND3 (N9123, N9115, N3490, N3566);
and AND3 (N9124, N9121, N4772, N2223);
nor NOR2 (N9125, N9122, N6098);
buf BUF1 (N9126, N9109);
and AND2 (N9127, N9125, N877);
xor XOR2 (N9128, N9107, N4505);
not NOT1 (N9129, N9128);
or OR4 (N9130, N9127, N6969, N6839, N6560);
buf BUF1 (N9131, N9124);
or OR2 (N9132, N9117, N4783);
xor XOR2 (N9133, N9129, N3241);
nor NOR3 (N9134, N9133, N7094, N8439);
or OR2 (N9135, N9126, N5801);
nand NAND2 (N9136, N9132, N5909);
and AND2 (N9137, N9134, N2742);
buf BUF1 (N9138, N9123);
or OR3 (N9139, N9118, N3719, N3440);
nor NOR3 (N9140, N9111, N2739, N5456);
or OR2 (N9141, N9139, N7407);
and AND2 (N9142, N9130, N2940);
buf BUF1 (N9143, N9138);
nand NAND4 (N9144, N9131, N4901, N6321, N5696);
buf BUF1 (N9145, N9144);
nor NOR4 (N9146, N9140, N950, N5933, N7629);
buf BUF1 (N9147, N9143);
and AND3 (N9148, N9136, N3043, N2718);
buf BUF1 (N9149, N9146);
or OR3 (N9150, N9147, N1232, N1776);
nand NAND3 (N9151, N9141, N3124, N6473);
nand NAND3 (N9152, N9142, N596, N2275);
and AND3 (N9153, N9099, N7269, N2990);
xor XOR2 (N9154, N9152, N4552);
nand NAND3 (N9155, N9149, N455, N4052);
buf BUF1 (N9156, N9150);
not NOT1 (N9157, N9153);
not NOT1 (N9158, N9135);
xor XOR2 (N9159, N9157, N1086);
or OR2 (N9160, N9093, N1400);
buf BUF1 (N9161, N9159);
buf BUF1 (N9162, N9148);
nand NAND2 (N9163, N9154, N572);
or OR2 (N9164, N9163, N8834);
nand NAND4 (N9165, N9164, N5038, N5992, N3186);
xor XOR2 (N9166, N9151, N1774);
not NOT1 (N9167, N9160);
nor NOR2 (N9168, N9167, N854);
nand NAND2 (N9169, N9165, N3140);
and AND4 (N9170, N9158, N2709, N6964, N7239);
or OR2 (N9171, N9137, N1600);
buf BUF1 (N9172, N9171);
nand NAND4 (N9173, N9155, N2316, N1098, N6717);
or OR4 (N9174, N9162, N7157, N803, N596);
not NOT1 (N9175, N9166);
not NOT1 (N9176, N9172);
or OR3 (N9177, N9145, N8334, N7346);
or OR2 (N9178, N9176, N3415);
and AND2 (N9179, N9175, N2747);
xor XOR2 (N9180, N9178, N2482);
or OR3 (N9181, N9179, N1961, N3150);
buf BUF1 (N9182, N9161);
xor XOR2 (N9183, N9173, N1821);
buf BUF1 (N9184, N9181);
nand NAND4 (N9185, N9177, N4650, N5966, N6442);
buf BUF1 (N9186, N9156);
buf BUF1 (N9187, N9180);
xor XOR2 (N9188, N9182, N775);
buf BUF1 (N9189, N9184);
buf BUF1 (N9190, N9188);
and AND3 (N9191, N9169, N3302, N5413);
not NOT1 (N9192, N9186);
nor NOR2 (N9193, N9183, N8290);
buf BUF1 (N9194, N9191);
buf BUF1 (N9195, N9185);
nor NOR2 (N9196, N9194, N6752);
nor NOR3 (N9197, N9187, N2504, N8006);
nand NAND3 (N9198, N9192, N3287, N7754);
nor NOR2 (N9199, N9190, N6985);
or OR4 (N9200, N9196, N2037, N8058, N3156);
and AND4 (N9201, N9197, N7242, N6172, N4322);
xor XOR2 (N9202, N9170, N4868);
nor NOR2 (N9203, N9200, N8817);
nand NAND2 (N9204, N9174, N9101);
buf BUF1 (N9205, N9198);
nand NAND2 (N9206, N9204, N4452);
or OR2 (N9207, N9168, N1769);
not NOT1 (N9208, N9206);
buf BUF1 (N9209, N9202);
or OR4 (N9210, N9208, N1076, N5377, N4894);
xor XOR2 (N9211, N9193, N5568);
or OR3 (N9212, N9210, N8362, N8346);
or OR2 (N9213, N9211, N787);
or OR4 (N9214, N9195, N2937, N7350, N4604);
buf BUF1 (N9215, N9213);
nor NOR4 (N9216, N9205, N7239, N4610, N2558);
buf BUF1 (N9217, N9209);
nand NAND2 (N9218, N9216, N1665);
nor NOR3 (N9219, N9212, N4266, N6389);
xor XOR2 (N9220, N9214, N492);
or OR3 (N9221, N9219, N4585, N5777);
and AND4 (N9222, N9201, N8867, N339, N1474);
xor XOR2 (N9223, N9189, N4902);
and AND3 (N9224, N9220, N135, N6130);
not NOT1 (N9225, N9203);
buf BUF1 (N9226, N9207);
nor NOR3 (N9227, N9218, N1735, N4920);
buf BUF1 (N9228, N9217);
buf BUF1 (N9229, N9228);
xor XOR2 (N9230, N9227, N567);
nand NAND4 (N9231, N9221, N8639, N8100, N5632);
nand NAND2 (N9232, N9231, N8577);
nand NAND4 (N9233, N9226, N2180, N1027, N3841);
buf BUF1 (N9234, N9223);
and AND2 (N9235, N9222, N3120);
nand NAND4 (N9236, N9232, N7435, N5886, N7851);
buf BUF1 (N9237, N9230);
and AND2 (N9238, N9236, N1350);
nand NAND3 (N9239, N9224, N6363, N1263);
buf BUF1 (N9240, N9234);
buf BUF1 (N9241, N9240);
not NOT1 (N9242, N9241);
xor XOR2 (N9243, N9233, N3860);
and AND2 (N9244, N9243, N3648);
nand NAND4 (N9245, N9237, N7071, N8692, N2780);
and AND2 (N9246, N9199, N7565);
or OR2 (N9247, N9245, N3305);
and AND3 (N9248, N9244, N3277, N466);
or OR3 (N9249, N9235, N8362, N8353);
nand NAND2 (N9250, N9248, N8880);
nand NAND2 (N9251, N9238, N2240);
and AND3 (N9252, N9242, N7517, N7559);
xor XOR2 (N9253, N9225, N4739);
xor XOR2 (N9254, N9246, N2684);
buf BUF1 (N9255, N9247);
not NOT1 (N9256, N9215);
nand NAND4 (N9257, N9254, N316, N3337, N5364);
not NOT1 (N9258, N9255);
nand NAND4 (N9259, N9256, N5917, N7009, N334);
or OR2 (N9260, N9253, N3272);
or OR2 (N9261, N9258, N6398);
nor NOR3 (N9262, N9260, N4784, N1005);
xor XOR2 (N9263, N9249, N191);
nand NAND2 (N9264, N9250, N7154);
and AND3 (N9265, N9259, N6713, N3158);
xor XOR2 (N9266, N9252, N1357);
and AND2 (N9267, N9257, N6263);
buf BUF1 (N9268, N9266);
xor XOR2 (N9269, N9268, N8868);
xor XOR2 (N9270, N9267, N5410);
nand NAND3 (N9271, N9239, N9163, N3432);
nor NOR3 (N9272, N9251, N7501, N264);
and AND4 (N9273, N9264, N2657, N5649, N4150);
buf BUF1 (N9274, N9261);
not NOT1 (N9275, N9274);
buf BUF1 (N9276, N9262);
buf BUF1 (N9277, N9272);
buf BUF1 (N9278, N9277);
buf BUF1 (N9279, N9275);
nand NAND2 (N9280, N9270, N4326);
not NOT1 (N9281, N9265);
not NOT1 (N9282, N9271);
nand NAND3 (N9283, N9282, N7838, N6495);
or OR2 (N9284, N9263, N479);
not NOT1 (N9285, N9276);
xor XOR2 (N9286, N9280, N5343);
buf BUF1 (N9287, N9285);
and AND4 (N9288, N9286, N1786, N16, N6744);
nand NAND2 (N9289, N9273, N5049);
nor NOR4 (N9290, N9269, N4947, N8278, N8578);
and AND4 (N9291, N9278, N6448, N8293, N5352);
and AND3 (N9292, N9289, N6637, N4796);
not NOT1 (N9293, N9287);
xor XOR2 (N9294, N9284, N9194);
and AND2 (N9295, N9279, N703);
buf BUF1 (N9296, N9291);
nor NOR4 (N9297, N9283, N2425, N4304, N3712);
nor NOR2 (N9298, N9293, N6219);
xor XOR2 (N9299, N9281, N178);
xor XOR2 (N9300, N9288, N2893);
nor NOR2 (N9301, N9295, N8774);
or OR4 (N9302, N9292, N3073, N5549, N7295);
not NOT1 (N9303, N9299);
and AND3 (N9304, N9301, N1321, N4189);
not NOT1 (N9305, N9300);
not NOT1 (N9306, N9302);
nand NAND4 (N9307, N9297, N5775, N2642, N3491);
not NOT1 (N9308, N9306);
or OR2 (N9309, N9307, N5749);
xor XOR2 (N9310, N9294, N7645);
xor XOR2 (N9311, N9296, N8328);
and AND3 (N9312, N9304, N5838, N8660);
and AND3 (N9313, N9309, N4630, N4306);
and AND4 (N9314, N9311, N7945, N4051, N8760);
nor NOR2 (N9315, N9305, N6843);
nor NOR2 (N9316, N9303, N8252);
buf BUF1 (N9317, N9314);
xor XOR2 (N9318, N9316, N584);
and AND4 (N9319, N9308, N727, N8337, N858);
buf BUF1 (N9320, N9312);
nor NOR2 (N9321, N9315, N7656);
buf BUF1 (N9322, N9319);
not NOT1 (N9323, N9322);
and AND2 (N9324, N9318, N4094);
buf BUF1 (N9325, N9313);
not NOT1 (N9326, N9320);
buf BUF1 (N9327, N9317);
not NOT1 (N9328, N9310);
xor XOR2 (N9329, N9326, N4085);
and AND3 (N9330, N9229, N7236, N354);
buf BUF1 (N9331, N9290);
nor NOR4 (N9332, N9328, N5353, N8369, N8720);
not NOT1 (N9333, N9327);
xor XOR2 (N9334, N9321, N5479);
and AND4 (N9335, N9332, N3687, N8944, N82);
buf BUF1 (N9336, N9335);
or OR2 (N9337, N9329, N7457);
nand NAND2 (N9338, N9334, N6573);
or OR4 (N9339, N9298, N6435, N3106, N5575);
or OR4 (N9340, N9324, N8208, N3704, N4435);
nand NAND2 (N9341, N9337, N3586);
or OR3 (N9342, N9330, N7070, N1734);
and AND3 (N9343, N9339, N801, N8105);
nor NOR4 (N9344, N9338, N3845, N5414, N7072);
or OR4 (N9345, N9333, N3173, N818, N3410);
xor XOR2 (N9346, N9336, N4973);
xor XOR2 (N9347, N9342, N3681);
buf BUF1 (N9348, N9346);
and AND4 (N9349, N9340, N74, N8997, N3570);
xor XOR2 (N9350, N9345, N788);
and AND3 (N9351, N9350, N6556, N112);
or OR3 (N9352, N9351, N6597, N738);
not NOT1 (N9353, N9331);
or OR4 (N9354, N9349, N3898, N2874, N84);
xor XOR2 (N9355, N9354, N6753);
nor NOR4 (N9356, N9343, N8709, N3040, N2385);
or OR3 (N9357, N9323, N1581, N5365);
buf BUF1 (N9358, N9347);
not NOT1 (N9359, N9357);
nor NOR4 (N9360, N9325, N6539, N7530, N8455);
nand NAND4 (N9361, N9348, N6615, N2272, N53);
xor XOR2 (N9362, N9355, N796);
or OR3 (N9363, N9352, N8650, N5471);
nor NOR3 (N9364, N9341, N5575, N319);
not NOT1 (N9365, N9363);
and AND2 (N9366, N9361, N5657);
nor NOR4 (N9367, N9364, N3939, N6679, N8357);
not NOT1 (N9368, N9358);
xor XOR2 (N9369, N9367, N9039);
xor XOR2 (N9370, N9353, N2769);
not NOT1 (N9371, N9365);
not NOT1 (N9372, N9370);
xor XOR2 (N9373, N9344, N9293);
nor NOR4 (N9374, N9373, N7265, N6116, N1101);
and AND4 (N9375, N9360, N4268, N1305, N3453);
nor NOR2 (N9376, N9366, N2068);
and AND2 (N9377, N9376, N6147);
or OR3 (N9378, N9377, N7488, N8537);
not NOT1 (N9379, N9372);
xor XOR2 (N9380, N9359, N2345);
xor XOR2 (N9381, N9375, N3020);
or OR4 (N9382, N9374, N6927, N5315, N5442);
not NOT1 (N9383, N9362);
buf BUF1 (N9384, N9381);
not NOT1 (N9385, N9380);
xor XOR2 (N9386, N9385, N3392);
nor NOR2 (N9387, N9368, N8776);
and AND3 (N9388, N9369, N916, N2124);
and AND4 (N9389, N9388, N6915, N2700, N8701);
xor XOR2 (N9390, N9384, N3970);
buf BUF1 (N9391, N9371);
not NOT1 (N9392, N9382);
and AND4 (N9393, N9390, N4443, N773, N3247);
or OR4 (N9394, N9387, N7668, N1708, N7994);
buf BUF1 (N9395, N9383);
xor XOR2 (N9396, N9394, N3546);
not NOT1 (N9397, N9378);
buf BUF1 (N9398, N9379);
buf BUF1 (N9399, N9389);
not NOT1 (N9400, N9393);
nor NOR3 (N9401, N9356, N4057, N8329);
buf BUF1 (N9402, N9395);
buf BUF1 (N9403, N9399);
xor XOR2 (N9404, N9396, N3939);
not NOT1 (N9405, N9392);
nand NAND3 (N9406, N9403, N2318, N6153);
and AND4 (N9407, N9400, N9350, N7327, N7767);
and AND2 (N9408, N9406, N3488);
or OR2 (N9409, N9386, N8369);
and AND2 (N9410, N9402, N1);
and AND2 (N9411, N9398, N3672);
nand NAND4 (N9412, N9410, N9253, N5318, N6119);
or OR3 (N9413, N9408, N6758, N855);
buf BUF1 (N9414, N9413);
and AND2 (N9415, N9397, N978);
and AND3 (N9416, N9414, N5176, N4082);
not NOT1 (N9417, N9404);
xor XOR2 (N9418, N9417, N3565);
buf BUF1 (N9419, N9416);
or OR4 (N9420, N9405, N5571, N3486, N2803);
xor XOR2 (N9421, N9412, N2926);
nor NOR3 (N9422, N9420, N1576, N8090);
xor XOR2 (N9423, N9407, N7243);
nor NOR2 (N9424, N9415, N3567);
nand NAND4 (N9425, N9424, N8880, N4411, N8965);
nor NOR4 (N9426, N9422, N6016, N6796, N6641);
not NOT1 (N9427, N9426);
or OR3 (N9428, N9411, N9391, N3150);
and AND3 (N9429, N3763, N1633, N2568);
nand NAND3 (N9430, N9428, N856, N7366);
xor XOR2 (N9431, N9419, N2583);
nor NOR4 (N9432, N9401, N612, N211, N9275);
not NOT1 (N9433, N9421);
nor NOR3 (N9434, N9430, N5127, N4505);
buf BUF1 (N9435, N9434);
buf BUF1 (N9436, N9433);
nor NOR2 (N9437, N9431, N7223);
or OR3 (N9438, N9436, N2026, N2452);
nor NOR3 (N9439, N9409, N159, N6952);
or OR3 (N9440, N9438, N4588, N284);
and AND2 (N9441, N9423, N3522);
or OR2 (N9442, N9418, N920);
not NOT1 (N9443, N9427);
nor NOR4 (N9444, N9425, N4129, N3618, N5626);
and AND3 (N9445, N9435, N131, N2712);
not NOT1 (N9446, N9440);
buf BUF1 (N9447, N9442);
buf BUF1 (N9448, N9447);
not NOT1 (N9449, N9448);
not NOT1 (N9450, N9446);
buf BUF1 (N9451, N9443);
or OR4 (N9452, N9439, N4236, N7017, N4131);
nand NAND4 (N9453, N9452, N6401, N2343, N4784);
xor XOR2 (N9454, N9444, N4582);
buf BUF1 (N9455, N9429);
not NOT1 (N9456, N9445);
and AND4 (N9457, N9456, N2606, N50, N8771);
buf BUF1 (N9458, N9454);
nand NAND2 (N9459, N9457, N3923);
nor NOR3 (N9460, N9449, N4320, N8805);
not NOT1 (N9461, N9458);
xor XOR2 (N9462, N9441, N1078);
xor XOR2 (N9463, N9459, N7703);
and AND3 (N9464, N9455, N2248, N4116);
buf BUF1 (N9465, N9461);
nor NOR4 (N9466, N9450, N5434, N1589, N8124);
buf BUF1 (N9467, N9462);
not NOT1 (N9468, N9437);
not NOT1 (N9469, N9451);
nand NAND2 (N9470, N9432, N5087);
not NOT1 (N9471, N9470);
nor NOR3 (N9472, N9460, N691, N8963);
xor XOR2 (N9473, N9464, N7739);
buf BUF1 (N9474, N9463);
or OR3 (N9475, N9467, N8034, N1422);
nor NOR2 (N9476, N9474, N3024);
or OR2 (N9477, N9472, N2093);
not NOT1 (N9478, N9471);
xor XOR2 (N9479, N9465, N6143);
or OR4 (N9480, N9473, N7698, N7139, N588);
not NOT1 (N9481, N9477);
nor NOR4 (N9482, N9469, N3942, N9067, N1637);
nor NOR4 (N9483, N9481, N9343, N3654, N8896);
nor NOR2 (N9484, N9483, N5357);
nor NOR3 (N9485, N9476, N8796, N6066);
nor NOR2 (N9486, N9484, N2394);
not NOT1 (N9487, N9466);
or OR3 (N9488, N9487, N9134, N4260);
not NOT1 (N9489, N9488);
nor NOR2 (N9490, N9486, N6078);
and AND4 (N9491, N9482, N4914, N7690, N8515);
nor NOR3 (N9492, N9490, N3846, N3239);
nand NAND2 (N9493, N9489, N1069);
or OR2 (N9494, N9493, N5400);
not NOT1 (N9495, N9478);
not NOT1 (N9496, N9479);
and AND4 (N9497, N9494, N1966, N5702, N1714);
xor XOR2 (N9498, N9495, N5618);
not NOT1 (N9499, N9475);
nor NOR4 (N9500, N9498, N8691, N6373, N2800);
xor XOR2 (N9501, N9499, N1177);
nor NOR3 (N9502, N9497, N6708, N1285);
and AND2 (N9503, N9491, N2267);
nor NOR3 (N9504, N9496, N7510, N6967);
and AND3 (N9505, N9502, N8253, N5819);
nor NOR3 (N9506, N9492, N181, N2072);
not NOT1 (N9507, N9505);
not NOT1 (N9508, N9500);
nor NOR4 (N9509, N9503, N7389, N823, N2998);
xor XOR2 (N9510, N9501, N348);
not NOT1 (N9511, N9468);
and AND4 (N9512, N9511, N4157, N1213, N2791);
xor XOR2 (N9513, N9506, N3104);
not NOT1 (N9514, N9508);
not NOT1 (N9515, N9514);
or OR2 (N9516, N9504, N6637);
and AND2 (N9517, N9480, N1949);
xor XOR2 (N9518, N9510, N2419);
nor NOR3 (N9519, N9518, N4944, N4473);
and AND3 (N9520, N9517, N3235, N7910);
and AND2 (N9521, N9515, N5782);
nor NOR4 (N9522, N9513, N7883, N1140, N5625);
nand NAND2 (N9523, N9519, N1687);
nand NAND2 (N9524, N9520, N4386);
and AND2 (N9525, N9485, N5218);
not NOT1 (N9526, N9509);
buf BUF1 (N9527, N9453);
not NOT1 (N9528, N9526);
or OR4 (N9529, N9522, N4086, N7346, N1271);
xor XOR2 (N9530, N9524, N3351);
or OR2 (N9531, N9516, N6564);
and AND4 (N9532, N9512, N5513, N3234, N3129);
nand NAND2 (N9533, N9529, N7);
nand NAND3 (N9534, N9532, N301, N7456);
nand NAND4 (N9535, N9523, N4183, N6672, N5636);
nand NAND4 (N9536, N9533, N7811, N672, N7112);
nor NOR2 (N9537, N9534, N3659);
xor XOR2 (N9538, N9521, N2128);
nor NOR4 (N9539, N9531, N2963, N3703, N7252);
xor XOR2 (N9540, N9525, N8644);
not NOT1 (N9541, N9527);
xor XOR2 (N9542, N9538, N1563);
or OR3 (N9543, N9539, N6789, N321);
xor XOR2 (N9544, N9542, N7355);
nor NOR2 (N9545, N9536, N3880);
nand NAND4 (N9546, N9535, N5873, N8393, N6857);
nor NOR2 (N9547, N9530, N5863);
and AND3 (N9548, N9546, N1699, N7543);
and AND3 (N9549, N9545, N5582, N1207);
nor NOR3 (N9550, N9543, N5799, N3967);
nand NAND4 (N9551, N9537, N4470, N8383, N7515);
nor NOR2 (N9552, N9540, N6804);
xor XOR2 (N9553, N9528, N8227);
and AND4 (N9554, N9507, N8221, N729, N1979);
nor NOR4 (N9555, N9549, N7490, N9547, N3766);
xor XOR2 (N9556, N6644, N6499);
nand NAND4 (N9557, N9551, N3201, N2803, N4853);
not NOT1 (N9558, N9555);
xor XOR2 (N9559, N9553, N8218);
xor XOR2 (N9560, N9558, N5470);
and AND3 (N9561, N9548, N2271, N6951);
xor XOR2 (N9562, N9550, N4358);
and AND4 (N9563, N9554, N7886, N6414, N5974);
and AND2 (N9564, N9561, N9257);
not NOT1 (N9565, N9562);
xor XOR2 (N9566, N9544, N7484);
or OR3 (N9567, N9541, N7652, N5621);
and AND2 (N9568, N9564, N4520);
buf BUF1 (N9569, N9556);
and AND2 (N9570, N9552, N5080);
nor NOR3 (N9571, N9563, N3327, N800);
nor NOR2 (N9572, N9571, N5709);
nor NOR2 (N9573, N9567, N5321);
or OR4 (N9574, N9560, N7740, N5658, N2605);
and AND2 (N9575, N9569, N8727);
nand NAND3 (N9576, N9557, N5343, N9456);
or OR3 (N9577, N9565, N7792, N3890);
nor NOR3 (N9578, N9572, N203, N5705);
and AND4 (N9579, N9577, N5051, N5584, N2714);
nand NAND3 (N9580, N9579, N2539, N3223);
nand NAND3 (N9581, N9580, N6040, N6791);
nor NOR3 (N9582, N9566, N14, N7059);
nor NOR4 (N9583, N9582, N6153, N6922, N6164);
buf BUF1 (N9584, N9583);
nor NOR2 (N9585, N9575, N1827);
nand NAND4 (N9586, N9585, N3042, N904, N1203);
buf BUF1 (N9587, N9581);
nand NAND3 (N9588, N9586, N610, N4794);
not NOT1 (N9589, N9576);
nand NAND2 (N9590, N9578, N3017);
not NOT1 (N9591, N9590);
nand NAND3 (N9592, N9584, N4297, N2663);
not NOT1 (N9593, N9589);
and AND2 (N9594, N9570, N851);
buf BUF1 (N9595, N9587);
nand NAND4 (N9596, N9574, N8472, N6677, N537);
or OR3 (N9597, N9591, N1147, N5983);
not NOT1 (N9598, N9573);
nor NOR4 (N9599, N9597, N353, N3146, N5367);
nand NAND3 (N9600, N9593, N1422, N794);
xor XOR2 (N9601, N9568, N1789);
xor XOR2 (N9602, N9588, N6294);
not NOT1 (N9603, N9598);
or OR4 (N9604, N9601, N4086, N4008, N4004);
not NOT1 (N9605, N9602);
buf BUF1 (N9606, N9603);
nand NAND2 (N9607, N9600, N6469);
buf BUF1 (N9608, N9607);
nor NOR4 (N9609, N9604, N1360, N5760, N6908);
not NOT1 (N9610, N9594);
and AND2 (N9611, N9595, N1301);
nand NAND3 (N9612, N9605, N9496, N1357);
or OR2 (N9613, N9611, N6501);
or OR3 (N9614, N9613, N6431, N2072);
buf BUF1 (N9615, N9559);
nor NOR3 (N9616, N9614, N7274, N8227);
nand NAND3 (N9617, N9592, N4562, N855);
nand NAND3 (N9618, N9599, N8391, N99);
xor XOR2 (N9619, N9612, N3944);
and AND4 (N9620, N9610, N3738, N5787, N5798);
and AND2 (N9621, N9616, N8109);
xor XOR2 (N9622, N9618, N6218);
xor XOR2 (N9623, N9615, N4205);
buf BUF1 (N9624, N9608);
not NOT1 (N9625, N9609);
not NOT1 (N9626, N9619);
nor NOR3 (N9627, N9620, N6896, N3545);
nor NOR3 (N9628, N9596, N9212, N8461);
nor NOR2 (N9629, N9627, N520);
nand NAND4 (N9630, N9624, N3955, N6385, N648);
nand NAND3 (N9631, N9606, N2474, N2932);
nor NOR3 (N9632, N9626, N1668, N5150);
or OR3 (N9633, N9617, N2593, N3649);
not NOT1 (N9634, N9630);
nor NOR3 (N9635, N9625, N3868, N1139);
xor XOR2 (N9636, N9628, N5635);
or OR3 (N9637, N9622, N974, N3536);
and AND3 (N9638, N9631, N1918, N5475);
and AND2 (N9639, N9636, N4092);
buf BUF1 (N9640, N9638);
xor XOR2 (N9641, N9623, N7624);
buf BUF1 (N9642, N9621);
buf BUF1 (N9643, N9640);
buf BUF1 (N9644, N9633);
xor XOR2 (N9645, N9635, N7372);
nand NAND3 (N9646, N9639, N7371, N8289);
xor XOR2 (N9647, N9629, N5852);
or OR3 (N9648, N9644, N5178, N7775);
buf BUF1 (N9649, N9641);
not NOT1 (N9650, N9647);
or OR2 (N9651, N9648, N8635);
and AND3 (N9652, N9645, N2969, N1687);
not NOT1 (N9653, N9646);
not NOT1 (N9654, N9643);
not NOT1 (N9655, N9642);
not NOT1 (N9656, N9632);
xor XOR2 (N9657, N9637, N5646);
or OR4 (N9658, N9634, N5762, N4003, N4454);
and AND4 (N9659, N9649, N8386, N4760, N6760);
buf BUF1 (N9660, N9654);
and AND2 (N9661, N9655, N1010);
or OR4 (N9662, N9661, N4817, N726, N6821);
nand NAND4 (N9663, N9656, N7004, N8115, N2264);
buf BUF1 (N9664, N9658);
not NOT1 (N9665, N9653);
not NOT1 (N9666, N9664);
buf BUF1 (N9667, N9662);
buf BUF1 (N9668, N9665);
nor NOR4 (N9669, N9663, N8150, N3622, N7197);
not NOT1 (N9670, N9660);
nor NOR2 (N9671, N9650, N1850);
nor NOR4 (N9672, N9668, N8379, N4254, N4358);
nor NOR3 (N9673, N9659, N5272, N812);
or OR3 (N9674, N9666, N5439, N2721);
not NOT1 (N9675, N9657);
nand NAND4 (N9676, N9672, N5852, N6636, N6374);
or OR3 (N9677, N9671, N8209, N7198);
and AND4 (N9678, N9651, N1509, N2344, N5049);
not NOT1 (N9679, N9675);
not NOT1 (N9680, N9678);
nand NAND4 (N9681, N9673, N8398, N240, N4597);
buf BUF1 (N9682, N9674);
and AND4 (N9683, N9682, N6187, N2240, N6858);
xor XOR2 (N9684, N9680, N2304);
buf BUF1 (N9685, N9667);
buf BUF1 (N9686, N9681);
buf BUF1 (N9687, N9683);
nor NOR2 (N9688, N9676, N2454);
and AND4 (N9689, N9679, N743, N8651, N6443);
and AND3 (N9690, N9670, N2428, N8771);
buf BUF1 (N9691, N9689);
or OR3 (N9692, N9686, N8446, N4038);
nor NOR3 (N9693, N9669, N1386, N6955);
nand NAND2 (N9694, N9685, N6275);
nor NOR3 (N9695, N9687, N8077, N461);
buf BUF1 (N9696, N9652);
xor XOR2 (N9697, N9695, N614);
xor XOR2 (N9698, N9677, N524);
and AND4 (N9699, N9696, N2651, N1606, N7619);
and AND2 (N9700, N9684, N5425);
or OR2 (N9701, N9699, N1024);
or OR3 (N9702, N9694, N4238, N5130);
buf BUF1 (N9703, N9701);
nor NOR2 (N9704, N9702, N5517);
not NOT1 (N9705, N9693);
and AND2 (N9706, N9697, N9341);
nand NAND3 (N9707, N9705, N3353, N5388);
nor NOR4 (N9708, N9706, N1354, N4942, N8961);
nand NAND2 (N9709, N9692, N2005);
nor NOR4 (N9710, N9708, N641, N9333, N4540);
nor NOR4 (N9711, N9698, N8820, N7073, N95);
not NOT1 (N9712, N9707);
buf BUF1 (N9713, N9703);
buf BUF1 (N9714, N9700);
or OR3 (N9715, N9712, N5597, N2044);
xor XOR2 (N9716, N9704, N5906);
and AND4 (N9717, N9714, N848, N8497, N2571);
xor XOR2 (N9718, N9716, N2453);
xor XOR2 (N9719, N9690, N5775);
or OR2 (N9720, N9713, N690);
nor NOR2 (N9721, N9720, N453);
nor NOR4 (N9722, N9688, N7695, N1119, N2153);
or OR2 (N9723, N9709, N3549);
nor NOR3 (N9724, N9719, N85, N7834);
nor NOR3 (N9725, N9717, N8429, N9296);
buf BUF1 (N9726, N9725);
buf BUF1 (N9727, N9711);
not NOT1 (N9728, N9722);
and AND4 (N9729, N9726, N580, N1190, N8949);
nand NAND4 (N9730, N9710, N6068, N7944, N5143);
or OR4 (N9731, N9728, N3603, N6810, N424);
or OR4 (N9732, N9729, N6055, N2375, N6498);
nor NOR4 (N9733, N9718, N4474, N8587, N2670);
buf BUF1 (N9734, N9715);
buf BUF1 (N9735, N9731);
and AND3 (N9736, N9691, N1853, N6724);
and AND4 (N9737, N9735, N3510, N7279, N6668);
xor XOR2 (N9738, N9733, N3847);
or OR3 (N9739, N9736, N6547, N8852);
not NOT1 (N9740, N9737);
or OR3 (N9741, N9723, N838, N7229);
and AND2 (N9742, N9741, N1587);
and AND2 (N9743, N9740, N7458);
or OR2 (N9744, N9732, N4207);
not NOT1 (N9745, N9742);
not NOT1 (N9746, N9721);
and AND3 (N9747, N9744, N5228, N5241);
nand NAND4 (N9748, N9747, N4067, N8738, N8257);
nand NAND2 (N9749, N9724, N8600);
not NOT1 (N9750, N9745);
nor NOR4 (N9751, N9749, N9136, N4396, N8960);
buf BUF1 (N9752, N9751);
buf BUF1 (N9753, N9748);
nor NOR2 (N9754, N9730, N7567);
and AND4 (N9755, N9746, N6919, N5444, N277);
nand NAND4 (N9756, N9734, N1359, N7739, N126);
nand NAND3 (N9757, N9755, N1020, N2119);
xor XOR2 (N9758, N9750, N3738);
nand NAND4 (N9759, N9727, N3262, N3093, N9307);
nor NOR4 (N9760, N9743, N7362, N5118, N59);
buf BUF1 (N9761, N9753);
nor NOR3 (N9762, N9761, N2677, N3021);
xor XOR2 (N9763, N9754, N8405);
and AND3 (N9764, N9763, N9307, N5022);
not NOT1 (N9765, N9764);
nor NOR4 (N9766, N9757, N7095, N5763, N1168);
not NOT1 (N9767, N9765);
xor XOR2 (N9768, N9759, N7833);
not NOT1 (N9769, N9756);
not NOT1 (N9770, N9758);
and AND2 (N9771, N9770, N4975);
not NOT1 (N9772, N9768);
nand NAND3 (N9773, N9767, N7276, N4088);
nand NAND4 (N9774, N9773, N3439, N6409, N7790);
nor NOR2 (N9775, N9738, N8277);
or OR2 (N9776, N9739, N85);
buf BUF1 (N9777, N9766);
nand NAND3 (N9778, N9777, N8414, N2980);
or OR2 (N9779, N9776, N3070);
or OR4 (N9780, N9769, N4298, N7437, N7184);
nor NOR2 (N9781, N9780, N5142);
and AND3 (N9782, N9778, N7143, N262);
not NOT1 (N9783, N9772);
buf BUF1 (N9784, N9781);
not NOT1 (N9785, N9783);
buf BUF1 (N9786, N9762);
not NOT1 (N9787, N9786);
or OR2 (N9788, N9787, N8033);
not NOT1 (N9789, N9779);
nand NAND4 (N9790, N9760, N7853, N6652, N9559);
nand NAND2 (N9791, N9788, N9430);
nand NAND4 (N9792, N9785, N5771, N2896, N1651);
buf BUF1 (N9793, N9791);
nor NOR2 (N9794, N9752, N6362);
and AND4 (N9795, N9774, N9065, N8697, N8605);
xor XOR2 (N9796, N9790, N7629);
xor XOR2 (N9797, N9794, N1016);
or OR4 (N9798, N9775, N1241, N224, N2575);
and AND4 (N9799, N9784, N9034, N2940, N2574);
xor XOR2 (N9800, N9792, N6446);
xor XOR2 (N9801, N9800, N6333);
buf BUF1 (N9802, N9799);
buf BUF1 (N9803, N9797);
buf BUF1 (N9804, N9793);
nor NOR3 (N9805, N9795, N8887, N9602);
nor NOR4 (N9806, N9801, N5243, N3253, N3851);
and AND2 (N9807, N9796, N4557);
and AND3 (N9808, N9771, N7542, N7928);
nand NAND4 (N9809, N9806, N7647, N4822, N4192);
xor XOR2 (N9810, N9809, N5717);
nand NAND3 (N9811, N9807, N9105, N4213);
nor NOR4 (N9812, N9798, N6289, N4761, N8047);
nor NOR2 (N9813, N9812, N3159);
buf BUF1 (N9814, N9802);
not NOT1 (N9815, N9789);
buf BUF1 (N9816, N9808);
and AND2 (N9817, N9814, N4114);
or OR3 (N9818, N9805, N2946, N1682);
buf BUF1 (N9819, N9818);
nand NAND3 (N9820, N9815, N9050, N8885);
nor NOR2 (N9821, N9803, N7881);
and AND2 (N9822, N9813, N4418);
and AND2 (N9823, N9820, N2317);
not NOT1 (N9824, N9804);
nand NAND4 (N9825, N9822, N402, N2539, N5771);
nand NAND4 (N9826, N9821, N9709, N656, N2546);
and AND3 (N9827, N9819, N1189, N6020);
not NOT1 (N9828, N9817);
xor XOR2 (N9829, N9810, N3164);
nor NOR4 (N9830, N9816, N2419, N7487, N9116);
not NOT1 (N9831, N9824);
and AND3 (N9832, N9827, N1149, N7522);
nor NOR2 (N9833, N9826, N5881);
nor NOR4 (N9834, N9823, N3626, N9531, N7139);
nor NOR4 (N9835, N9829, N6620, N3838, N8373);
or OR4 (N9836, N9835, N8549, N6012, N7899);
buf BUF1 (N9837, N9836);
and AND2 (N9838, N9837, N2871);
not NOT1 (N9839, N9832);
nor NOR4 (N9840, N9782, N7522, N4872, N2050);
and AND3 (N9841, N9833, N2227, N1279);
nand NAND4 (N9842, N9840, N1177, N319, N6263);
and AND4 (N9843, N9830, N3250, N1368, N7956);
not NOT1 (N9844, N9831);
xor XOR2 (N9845, N9839, N3569);
or OR3 (N9846, N9834, N9036, N4975);
buf BUF1 (N9847, N9825);
xor XOR2 (N9848, N9838, N4293);
buf BUF1 (N9849, N9848);
nor NOR4 (N9850, N9828, N9236, N1731, N3862);
xor XOR2 (N9851, N9846, N7590);
xor XOR2 (N9852, N9844, N6161);
xor XOR2 (N9853, N9843, N4671);
nand NAND4 (N9854, N9841, N6603, N2617, N5637);
buf BUF1 (N9855, N9842);
or OR2 (N9856, N9845, N6467);
nand NAND3 (N9857, N9849, N6905, N2576);
buf BUF1 (N9858, N9853);
and AND4 (N9859, N9858, N4947, N7269, N3763);
nand NAND2 (N9860, N9856, N7394);
not NOT1 (N9861, N9859);
not NOT1 (N9862, N9811);
or OR2 (N9863, N9855, N7992);
nor NOR3 (N9864, N9863, N8214, N3818);
not NOT1 (N9865, N9860);
or OR3 (N9866, N9862, N1502, N7889);
and AND3 (N9867, N9865, N4643, N1981);
nor NOR2 (N9868, N9852, N3095);
xor XOR2 (N9869, N9866, N8102);
nor NOR4 (N9870, N9869, N6481, N3412, N645);
not NOT1 (N9871, N9847);
buf BUF1 (N9872, N9861);
and AND2 (N9873, N9854, N675);
not NOT1 (N9874, N9864);
nand NAND2 (N9875, N9868, N241);
or OR2 (N9876, N9850, N1667);
nor NOR4 (N9877, N9873, N1832, N5048, N9670);
or OR3 (N9878, N9871, N4890, N7356);
not NOT1 (N9879, N9876);
and AND2 (N9880, N9872, N9311);
xor XOR2 (N9881, N9851, N6940);
nor NOR3 (N9882, N9875, N1328, N2156);
buf BUF1 (N9883, N9874);
or OR2 (N9884, N9878, N3200);
xor XOR2 (N9885, N9884, N8092);
nand NAND3 (N9886, N9870, N3868, N7888);
nand NAND4 (N9887, N9857, N857, N5259, N5829);
and AND2 (N9888, N9877, N120);
nor NOR3 (N9889, N9888, N4334, N3103);
not NOT1 (N9890, N9882);
not NOT1 (N9891, N9889);
nand NAND2 (N9892, N9890, N6544);
nand NAND4 (N9893, N9880, N6922, N9838, N6873);
xor XOR2 (N9894, N9881, N9892);
xor XOR2 (N9895, N6836, N408);
and AND4 (N9896, N9895, N8528, N5284, N6721);
or OR4 (N9897, N9883, N2246, N7310, N681);
and AND4 (N9898, N9885, N370, N4709, N3425);
xor XOR2 (N9899, N9897, N6614);
or OR2 (N9900, N9879, N8804);
nor NOR3 (N9901, N9898, N8927, N22);
and AND3 (N9902, N9894, N3074, N8133);
not NOT1 (N9903, N9891);
nor NOR4 (N9904, N9886, N7263, N5763, N8406);
buf BUF1 (N9905, N9902);
and AND3 (N9906, N9893, N2398, N2811);
or OR4 (N9907, N9900, N227, N8087, N7686);
not NOT1 (N9908, N9887);
buf BUF1 (N9909, N9905);
or OR4 (N9910, N9896, N3381, N4285, N2583);
or OR3 (N9911, N9904, N3183, N7203);
not NOT1 (N9912, N9910);
not NOT1 (N9913, N9906);
and AND4 (N9914, N9908, N9566, N6666, N7683);
nand NAND3 (N9915, N9909, N8395, N6923);
nor NOR4 (N9916, N9912, N3221, N2053, N8388);
and AND2 (N9917, N9913, N4510);
not NOT1 (N9918, N9917);
nor NOR4 (N9919, N9918, N4690, N7563, N3991);
xor XOR2 (N9920, N9903, N4889);
or OR4 (N9921, N9915, N3555, N6062, N9047);
xor XOR2 (N9922, N9911, N6734);
not NOT1 (N9923, N9914);
nor NOR3 (N9924, N9901, N6898, N3156);
buf BUF1 (N9925, N9924);
not NOT1 (N9926, N9922);
not NOT1 (N9927, N9867);
nand NAND4 (N9928, N9899, N6653, N255, N8067);
xor XOR2 (N9929, N9927, N8207);
nor NOR2 (N9930, N9929, N6313);
or OR4 (N9931, N9907, N9826, N5918, N3894);
or OR4 (N9932, N9926, N4362, N758, N6696);
or OR3 (N9933, N9919, N8173, N6276);
not NOT1 (N9934, N9920);
not NOT1 (N9935, N9925);
buf BUF1 (N9936, N9923);
and AND3 (N9937, N9932, N564, N7214);
xor XOR2 (N9938, N9930, N1403);
xor XOR2 (N9939, N9938, N8794);
nor NOR4 (N9940, N9937, N5168, N8401, N1215);
buf BUF1 (N9941, N9935);
and AND4 (N9942, N9934, N3178, N2551, N9904);
and AND3 (N9943, N9942, N7236, N5145);
xor XOR2 (N9944, N9941, N8276);
not NOT1 (N9945, N9939);
nor NOR3 (N9946, N9943, N6757, N9642);
xor XOR2 (N9947, N9916, N3349);
xor XOR2 (N9948, N9947, N2256);
buf BUF1 (N9949, N9940);
or OR2 (N9950, N9949, N8217);
buf BUF1 (N9951, N9944);
nand NAND2 (N9952, N9921, N6563);
not NOT1 (N9953, N9948);
or OR4 (N9954, N9936, N4341, N3264, N8473);
nor NOR3 (N9955, N9952, N1324, N1537);
or OR4 (N9956, N9955, N4940, N2292, N856);
and AND3 (N9957, N9931, N1024, N1790);
xor XOR2 (N9958, N9933, N8577);
and AND2 (N9959, N9956, N3261);
nand NAND4 (N9960, N9953, N3802, N9390, N2498);
and AND3 (N9961, N9959, N5384, N3412);
xor XOR2 (N9962, N9928, N4308);
xor XOR2 (N9963, N9958, N781);
buf BUF1 (N9964, N9951);
xor XOR2 (N9965, N9954, N5871);
nand NAND4 (N9966, N9962, N8633, N6598, N6056);
not NOT1 (N9967, N9966);
or OR3 (N9968, N9965, N6197, N4355);
nand NAND4 (N9969, N9960, N4568, N3205, N583);
and AND2 (N9970, N9950, N9551);
xor XOR2 (N9971, N9968, N9040);
buf BUF1 (N9972, N9964);
nand NAND4 (N9973, N9972, N5152, N3427, N20);
or OR3 (N9974, N9961, N7455, N2);
nor NOR2 (N9975, N9970, N1327);
not NOT1 (N9976, N9946);
xor XOR2 (N9977, N9974, N2326);
buf BUF1 (N9978, N9973);
nand NAND2 (N9979, N9963, N504);
buf BUF1 (N9980, N9978);
nor NOR2 (N9981, N9976, N2612);
buf BUF1 (N9982, N9981);
nor NOR3 (N9983, N9945, N699, N2389);
nor NOR3 (N9984, N9957, N1253, N573);
or OR4 (N9985, N9984, N1940, N4069, N2920);
xor XOR2 (N9986, N9983, N3498);
nor NOR4 (N9987, N9986, N79, N9131, N8572);
nor NOR4 (N9988, N9977, N8655, N3508, N1963);
or OR3 (N9989, N9987, N8147, N4588);
nor NOR2 (N9990, N9971, N5963);
or OR4 (N9991, N9985, N2417, N4107, N8922);
buf BUF1 (N9992, N9990);
xor XOR2 (N9993, N9989, N2149);
nand NAND2 (N9994, N9980, N9409);
or OR4 (N9995, N9994, N4497, N8377, N8614);
and AND3 (N9996, N9975, N3801, N6183);
not NOT1 (N9997, N9995);
or OR2 (N9998, N9996, N5856);
and AND2 (N9999, N9992, N6513);
nor NOR3 (N10000, N9988, N8387, N8333);
or OR2 (N10001, N9998, N6868);
not NOT1 (N10002, N9982);
nor NOR2 (N10003, N9979, N2751);
and AND2 (N10004, N10001, N7439);
nor NOR3 (N10005, N9993, N94, N5900);
nor NOR2 (N10006, N10005, N6397);
not NOT1 (N10007, N9967);
not NOT1 (N10008, N10002);
buf BUF1 (N10009, N10006);
buf BUF1 (N10010, N9991);
or OR2 (N10011, N10009, N3339);
buf BUF1 (N10012, N10004);
not NOT1 (N10013, N10000);
buf BUF1 (N10014, N10012);
nand NAND3 (N10015, N10014, N9778, N1348);
xor XOR2 (N10016, N10015, N5790);
or OR3 (N10017, N10013, N2774, N1746);
buf BUF1 (N10018, N10017);
or OR4 (N10019, N10007, N6302, N3875, N5860);
not NOT1 (N10020, N10003);
buf BUF1 (N10021, N9997);
not NOT1 (N10022, N10016);
or OR2 (N10023, N9999, N898);
nor NOR3 (N10024, N9969, N8078, N3155);
or OR3 (N10025, N10023, N7905, N7493);
and AND3 (N10026, N10018, N8740, N9879);
buf BUF1 (N10027, N10008);
and AND3 (N10028, N10027, N5683, N5743);
buf BUF1 (N10029, N10011);
nand NAND2 (N10030, N10021, N664);
nand NAND2 (N10031, N10024, N8113);
or OR3 (N10032, N10029, N1431, N3281);
xor XOR2 (N10033, N10022, N5426);
or OR2 (N10034, N10010, N5628);
nand NAND4 (N10035, N10034, N8733, N1403, N6494);
not NOT1 (N10036, N10033);
not NOT1 (N10037, N10020);
buf BUF1 (N10038, N10019);
buf BUF1 (N10039, N10025);
nand NAND4 (N10040, N10036, N2961, N7993, N9140);
and AND3 (N10041, N10037, N8640, N3539);
xor XOR2 (N10042, N10032, N7577);
or OR3 (N10043, N10028, N3250, N9649);
nand NAND2 (N10044, N10026, N3516);
or OR2 (N10045, N10030, N8445);
or OR4 (N10046, N10041, N3725, N8258, N8178);
and AND2 (N10047, N10039, N5115);
and AND3 (N10048, N10038, N4853, N6389);
not NOT1 (N10049, N10035);
xor XOR2 (N10050, N10031, N4942);
or OR4 (N10051, N10049, N4490, N9255, N1329);
xor XOR2 (N10052, N10050, N9352);
or OR4 (N10053, N10044, N9710, N46, N2769);
and AND2 (N10054, N10048, N7027);
and AND2 (N10055, N10052, N793);
buf BUF1 (N10056, N10055);
and AND3 (N10057, N10040, N4696, N6699);
nor NOR2 (N10058, N10056, N8263);
or OR4 (N10059, N10042, N476, N3837, N6641);
not NOT1 (N10060, N10047);
or OR4 (N10061, N10057, N3033, N2767, N5067);
nand NAND2 (N10062, N10053, N415);
not NOT1 (N10063, N10060);
buf BUF1 (N10064, N10054);
xor XOR2 (N10065, N10045, N8395);
nand NAND4 (N10066, N10043, N6187, N5336, N5979);
not NOT1 (N10067, N10064);
nand NAND3 (N10068, N10065, N1846, N3778);
not NOT1 (N10069, N10066);
buf BUF1 (N10070, N10069);
xor XOR2 (N10071, N10046, N7301);
buf BUF1 (N10072, N10061);
not NOT1 (N10073, N10067);
or OR2 (N10074, N10059, N6939);
not NOT1 (N10075, N10072);
not NOT1 (N10076, N10070);
or OR3 (N10077, N10063, N6284, N4697);
not NOT1 (N10078, N10058);
xor XOR2 (N10079, N10073, N7276);
nand NAND3 (N10080, N10076, N6922, N6790);
nor NOR3 (N10081, N10051, N7161, N3831);
or OR3 (N10082, N10074, N7579, N5549);
or OR3 (N10083, N10080, N6629, N9231);
buf BUF1 (N10084, N10078);
nor NOR3 (N10085, N10081, N8851, N9508);
buf BUF1 (N10086, N10071);
nor NOR3 (N10087, N10084, N6271, N788);
and AND4 (N10088, N10077, N7970, N2649, N8538);
and AND3 (N10089, N10086, N4720, N6444);
nand NAND4 (N10090, N10085, N2016, N1110, N3562);
nand NAND3 (N10091, N10090, N3188, N5735);
nor NOR4 (N10092, N10089, N937, N9186, N6926);
or OR2 (N10093, N10087, N3848);
or OR2 (N10094, N10091, N6969);
not NOT1 (N10095, N10094);
nor NOR2 (N10096, N10093, N9813);
nor NOR2 (N10097, N10096, N2425);
and AND4 (N10098, N10083, N891, N836, N9996);
nand NAND4 (N10099, N10095, N9021, N8840, N8182);
xor XOR2 (N10100, N10088, N6753);
not NOT1 (N10101, N10100);
not NOT1 (N10102, N10079);
and AND4 (N10103, N10062, N3893, N7131, N2198);
or OR3 (N10104, N10103, N8484, N2905);
or OR4 (N10105, N10082, N3873, N2748, N8953);
and AND4 (N10106, N10098, N3475, N7984, N7560);
nor NOR2 (N10107, N10099, N1180);
not NOT1 (N10108, N10102);
nand NAND3 (N10109, N10092, N5476, N5839);
or OR4 (N10110, N10105, N7427, N9030, N9971);
nor NOR4 (N10111, N10109, N4328, N8754, N3964);
nor NOR4 (N10112, N10104, N3992, N3892, N5323);
buf BUF1 (N10113, N10110);
not NOT1 (N10114, N10112);
nand NAND3 (N10115, N10106, N7702, N790);
nand NAND2 (N10116, N10114, N8252);
nor NOR2 (N10117, N10113, N44);
nor NOR2 (N10118, N10111, N4827);
or OR2 (N10119, N10118, N8386);
nand NAND2 (N10120, N10108, N1624);
xor XOR2 (N10121, N10119, N2531);
nand NAND4 (N10122, N10101, N836, N8720, N9424);
or OR2 (N10123, N10116, N9832);
buf BUF1 (N10124, N10122);
nor NOR4 (N10125, N10068, N8737, N5951, N5882);
or OR3 (N10126, N10075, N2815, N5833);
and AND4 (N10127, N10107, N9881, N8845, N1297);
nand NAND3 (N10128, N10125, N7916, N2959);
buf BUF1 (N10129, N10120);
buf BUF1 (N10130, N10126);
buf BUF1 (N10131, N10130);
nand NAND4 (N10132, N10123, N9771, N2917, N5966);
nand NAND2 (N10133, N10127, N2135);
not NOT1 (N10134, N10132);
or OR2 (N10135, N10128, N2960);
xor XOR2 (N10136, N10131, N8065);
or OR2 (N10137, N10121, N6416);
nor NOR4 (N10138, N10117, N1069, N2491, N5702);
and AND3 (N10139, N10136, N5660, N4269);
xor XOR2 (N10140, N10137, N7214);
or OR3 (N10141, N10133, N5900, N7186);
not NOT1 (N10142, N10124);
or OR3 (N10143, N10129, N5148, N5531);
nor NOR3 (N10144, N10097, N606, N754);
nor NOR2 (N10145, N10138, N2518);
nand NAND3 (N10146, N10144, N3119, N4765);
and AND3 (N10147, N10139, N672, N3514);
buf BUF1 (N10148, N10143);
nand NAND3 (N10149, N10141, N1345, N9227);
nand NAND3 (N10150, N10135, N4592, N1268);
not NOT1 (N10151, N10115);
and AND2 (N10152, N10142, N8132);
nor NOR3 (N10153, N10134, N6803, N7830);
xor XOR2 (N10154, N10147, N1323);
buf BUF1 (N10155, N10150);
nand NAND4 (N10156, N10146, N2943, N8760, N7783);
nor NOR3 (N10157, N10149, N1738, N6084);
not NOT1 (N10158, N10153);
nand NAND4 (N10159, N10145, N6443, N9454, N5127);
xor XOR2 (N10160, N10157, N2557);
or OR3 (N10161, N10148, N9761, N2316);
or OR3 (N10162, N10155, N3995, N7225);
not NOT1 (N10163, N10156);
or OR4 (N10164, N10154, N1553, N4405, N8009);
not NOT1 (N10165, N10151);
and AND2 (N10166, N10161, N2907);
nor NOR4 (N10167, N10162, N1032, N494, N8626);
nand NAND3 (N10168, N10164, N8080, N7144);
nand NAND4 (N10169, N10160, N10085, N5397, N10014);
buf BUF1 (N10170, N10163);
xor XOR2 (N10171, N10169, N3795);
xor XOR2 (N10172, N10168, N6748);
nor NOR4 (N10173, N10158, N1498, N5218, N4218);
nand NAND2 (N10174, N10173, N8959);
and AND3 (N10175, N10170, N5064, N1938);
and AND3 (N10176, N10152, N1034, N1517);
nor NOR3 (N10177, N10175, N2088, N362);
xor XOR2 (N10178, N10174, N9824);
xor XOR2 (N10179, N10140, N5262);
buf BUF1 (N10180, N10176);
or OR3 (N10181, N10165, N5204, N3282);
not NOT1 (N10182, N10171);
and AND3 (N10183, N10166, N5835, N4);
nand NAND3 (N10184, N10183, N4961, N8826);
nand NAND3 (N10185, N10179, N6884, N3276);
buf BUF1 (N10186, N10180);
buf BUF1 (N10187, N10185);
or OR2 (N10188, N10187, N1108);
or OR4 (N10189, N10181, N7438, N8489, N9664);
and AND2 (N10190, N10184, N8095);
nor NOR3 (N10191, N10190, N9113, N1085);
nor NOR4 (N10192, N10172, N3174, N9332, N3049);
not NOT1 (N10193, N10177);
and AND2 (N10194, N10192, N31);
xor XOR2 (N10195, N10191, N5034);
xor XOR2 (N10196, N10189, N5307);
xor XOR2 (N10197, N10196, N9488);
nand NAND3 (N10198, N10182, N6731, N2857);
buf BUF1 (N10199, N10167);
nor NOR3 (N10200, N10159, N6106, N8541);
not NOT1 (N10201, N10199);
nand NAND4 (N10202, N10195, N3510, N1514, N4754);
nor NOR4 (N10203, N10193, N642, N4497, N1736);
not NOT1 (N10204, N10202);
nor NOR2 (N10205, N10198, N10201);
nand NAND3 (N10206, N4434, N3095, N9033);
buf BUF1 (N10207, N10186);
xor XOR2 (N10208, N10206, N933);
nand NAND2 (N10209, N10203, N9394);
or OR3 (N10210, N10207, N8478, N2553);
and AND4 (N10211, N10210, N10099, N6665, N5452);
or OR4 (N10212, N10204, N3539, N7221, N3963);
nand NAND4 (N10213, N10178, N1977, N5466, N4377);
and AND3 (N10214, N10194, N3329, N9481);
nor NOR2 (N10215, N10200, N6914);
not NOT1 (N10216, N10212);
nand NAND3 (N10217, N10211, N2809, N10145);
nand NAND4 (N10218, N10209, N4590, N9183, N7844);
xor XOR2 (N10219, N10197, N4890);
not NOT1 (N10220, N10218);
and AND2 (N10221, N10216, N6699);
nor NOR4 (N10222, N10215, N2942, N4435, N5655);
and AND2 (N10223, N10213, N4025);
nand NAND4 (N10224, N10208, N3562, N7806, N3275);
or OR2 (N10225, N10205, N6771);
nand NAND2 (N10226, N10225, N1904);
nor NOR3 (N10227, N10222, N4274, N2335);
not NOT1 (N10228, N10214);
and AND3 (N10229, N10217, N5649, N5913);
not NOT1 (N10230, N10221);
buf BUF1 (N10231, N10188);
and AND4 (N10232, N10220, N6661, N2329, N10140);
buf BUF1 (N10233, N10228);
and AND2 (N10234, N10227, N4304);
buf BUF1 (N10235, N10230);
buf BUF1 (N10236, N10235);
and AND2 (N10237, N10233, N7201);
xor XOR2 (N10238, N10236, N3102);
xor XOR2 (N10239, N10226, N6125);
and AND4 (N10240, N10219, N9581, N2092, N6246);
and AND3 (N10241, N10237, N9935, N1329);
nor NOR3 (N10242, N10238, N3989, N1030);
and AND4 (N10243, N10224, N4183, N1315, N8516);
buf BUF1 (N10244, N10234);
or OR2 (N10245, N10239, N959);
nand NAND3 (N10246, N10245, N3556, N1343);
nand NAND3 (N10247, N10223, N1626, N4741);
and AND4 (N10248, N10232, N8816, N7338, N8235);
xor XOR2 (N10249, N10229, N5596);
and AND2 (N10250, N10242, N9985);
and AND4 (N10251, N10241, N5759, N3815, N10090);
xor XOR2 (N10252, N10249, N335);
or OR2 (N10253, N10243, N210);
and AND3 (N10254, N10247, N8864, N6874);
buf BUF1 (N10255, N10248);
and AND2 (N10256, N10251, N8147);
nor NOR2 (N10257, N10256, N4201);
or OR2 (N10258, N10255, N331);
nand NAND2 (N10259, N10253, N757);
not NOT1 (N10260, N10252);
and AND3 (N10261, N10250, N5601, N8472);
nand NAND2 (N10262, N10246, N2217);
xor XOR2 (N10263, N10260, N4428);
nor NOR3 (N10264, N10254, N7023, N6643);
nand NAND2 (N10265, N10257, N5428);
or OR2 (N10266, N10264, N6043);
nand NAND2 (N10267, N10259, N3693);
or OR3 (N10268, N10258, N10221, N7836);
buf BUF1 (N10269, N10263);
not NOT1 (N10270, N10266);
xor XOR2 (N10271, N10267, N3356);
not NOT1 (N10272, N10244);
nand NAND2 (N10273, N10271, N9667);
nor NOR3 (N10274, N10273, N5723, N1541);
buf BUF1 (N10275, N10270);
and AND3 (N10276, N10272, N1270, N3508);
nor NOR3 (N10277, N10265, N1247, N8623);
not NOT1 (N10278, N10262);
xor XOR2 (N10279, N10240, N1148);
nand NAND3 (N10280, N10277, N5538, N1169);
not NOT1 (N10281, N10276);
nor NOR3 (N10282, N10261, N4848, N1502);
nand NAND3 (N10283, N10281, N6079, N4037);
not NOT1 (N10284, N10274);
and AND2 (N10285, N10279, N6973);
or OR2 (N10286, N10282, N1001);
not NOT1 (N10287, N10286);
not NOT1 (N10288, N10231);
or OR4 (N10289, N10280, N2791, N2093, N4165);
or OR4 (N10290, N10288, N6904, N4003, N1011);
or OR3 (N10291, N10289, N5816, N5812);
buf BUF1 (N10292, N10291);
not NOT1 (N10293, N10269);
nor NOR4 (N10294, N10293, N9435, N8808, N2674);
xor XOR2 (N10295, N10287, N641);
not NOT1 (N10296, N10285);
nand NAND4 (N10297, N10292, N10110, N154, N8663);
nor NOR3 (N10298, N10297, N10035, N5022);
xor XOR2 (N10299, N10298, N3406);
nand NAND2 (N10300, N10295, N6229);
xor XOR2 (N10301, N10294, N1125);
not NOT1 (N10302, N10290);
or OR3 (N10303, N10300, N3590, N5000);
or OR4 (N10304, N10283, N8327, N7803, N5023);
and AND2 (N10305, N10278, N2493);
or OR3 (N10306, N10303, N5731, N5637);
nor NOR4 (N10307, N10275, N4815, N1460, N9226);
xor XOR2 (N10308, N10296, N5364);
or OR4 (N10309, N10301, N4213, N7279, N5939);
nor NOR3 (N10310, N10308, N6895, N4977);
nand NAND4 (N10311, N10307, N4129, N6691, N6493);
xor XOR2 (N10312, N10309, N10000);
nor NOR4 (N10313, N10268, N6450, N451, N9393);
nor NOR4 (N10314, N10304, N7411, N7646, N5590);
and AND2 (N10315, N10312, N4579);
buf BUF1 (N10316, N10310);
not NOT1 (N10317, N10306);
and AND3 (N10318, N10317, N8006, N942);
and AND4 (N10319, N10314, N8547, N4893, N7218);
or OR3 (N10320, N10311, N1458, N8185);
xor XOR2 (N10321, N10320, N2584);
nand NAND4 (N10322, N10318, N273, N5553, N5040);
xor XOR2 (N10323, N10284, N8558);
nand NAND3 (N10324, N10305, N7850, N9387);
xor XOR2 (N10325, N10316, N233);
and AND2 (N10326, N10313, N9921);
nor NOR4 (N10327, N10319, N3579, N3529, N3828);
nor NOR4 (N10328, N10324, N6846, N6358, N1350);
nor NOR3 (N10329, N10327, N435, N1569);
not NOT1 (N10330, N10299);
or OR2 (N10331, N10325, N10022);
or OR2 (N10332, N10321, N300);
buf BUF1 (N10333, N10322);
nor NOR3 (N10334, N10333, N4828, N9590);
not NOT1 (N10335, N10326);
nand NAND2 (N10336, N10302, N9267);
or OR2 (N10337, N10336, N9912);
or OR2 (N10338, N10328, N9969);
not NOT1 (N10339, N10329);
or OR3 (N10340, N10323, N2774, N5429);
buf BUF1 (N10341, N10334);
not NOT1 (N10342, N10341);
not NOT1 (N10343, N10330);
nand NAND2 (N10344, N10331, N8386);
and AND4 (N10345, N10342, N3050, N10261, N1135);
nor NOR2 (N10346, N10335, N467);
xor XOR2 (N10347, N10345, N7691);
or OR3 (N10348, N10332, N2748, N10090);
nand NAND4 (N10349, N10340, N8938, N4108, N6234);
or OR4 (N10350, N10344, N4509, N6484, N7335);
or OR3 (N10351, N10347, N8094, N6152);
and AND4 (N10352, N10343, N7801, N4274, N5454);
nor NOR2 (N10353, N10338, N9680);
or OR4 (N10354, N10337, N9851, N8758, N153);
not NOT1 (N10355, N10315);
nand NAND2 (N10356, N10346, N6798);
xor XOR2 (N10357, N10355, N8771);
and AND4 (N10358, N10349, N6463, N7736, N8468);
buf BUF1 (N10359, N10356);
and AND2 (N10360, N10359, N532);
xor XOR2 (N10361, N10360, N993);
nor NOR2 (N10362, N10350, N4937);
or OR4 (N10363, N10358, N2444, N2887, N6629);
not NOT1 (N10364, N10362);
or OR2 (N10365, N10361, N2047);
nor NOR4 (N10366, N10351, N5661, N3350, N6279);
nand NAND2 (N10367, N10339, N8548);
and AND4 (N10368, N10348, N5443, N9476, N3186);
nand NAND4 (N10369, N10368, N1319, N1974, N6485);
buf BUF1 (N10370, N10369);
xor XOR2 (N10371, N10353, N4507);
nand NAND3 (N10372, N10364, N2278, N8258);
nor NOR3 (N10373, N10365, N7407, N1553);
xor XOR2 (N10374, N10357, N8502);
not NOT1 (N10375, N10373);
xor XOR2 (N10376, N10374, N778);
and AND2 (N10377, N10354, N5514);
nand NAND3 (N10378, N10377, N946, N8772);
and AND3 (N10379, N10363, N579, N7488);
and AND2 (N10380, N10378, N8013);
not NOT1 (N10381, N10366);
nand NAND2 (N10382, N10380, N4248);
xor XOR2 (N10383, N10367, N169);
nor NOR2 (N10384, N10371, N6127);
or OR4 (N10385, N10383, N7003, N1370, N858);
and AND4 (N10386, N10382, N3615, N1680, N9843);
not NOT1 (N10387, N10370);
nand NAND2 (N10388, N10352, N4440);
and AND3 (N10389, N10376, N1130, N8640);
and AND4 (N10390, N10388, N6943, N7563, N7899);
buf BUF1 (N10391, N10389);
nand NAND4 (N10392, N10391, N6442, N9574, N4492);
nand NAND2 (N10393, N10392, N8220);
or OR3 (N10394, N10372, N9860, N1981);
nor NOR4 (N10395, N10390, N4835, N7978, N6183);
or OR3 (N10396, N10386, N6986, N5364);
not NOT1 (N10397, N10387);
nor NOR3 (N10398, N10379, N9800, N6408);
buf BUF1 (N10399, N10394);
buf BUF1 (N10400, N10398);
not NOT1 (N10401, N10375);
xor XOR2 (N10402, N10397, N7439);
nand NAND4 (N10403, N10399, N3952, N2988, N667);
nand NAND4 (N10404, N10395, N7546, N4735, N1304);
xor XOR2 (N10405, N10384, N1555);
not NOT1 (N10406, N10404);
xor XOR2 (N10407, N10401, N779);
xor XOR2 (N10408, N10405, N8655);
buf BUF1 (N10409, N10408);
buf BUF1 (N10410, N10385);
xor XOR2 (N10411, N10402, N4058);
buf BUF1 (N10412, N10411);
nand NAND2 (N10413, N10407, N9049);
nor NOR4 (N10414, N10413, N6422, N4429, N4266);
xor XOR2 (N10415, N10406, N2918);
and AND2 (N10416, N10393, N3995);
or OR2 (N10417, N10414, N1307);
buf BUF1 (N10418, N10381);
and AND4 (N10419, N10418, N3464, N4349, N4634);
xor XOR2 (N10420, N10400, N8387);
nand NAND3 (N10421, N10419, N5844, N5687);
and AND2 (N10422, N10417, N4247);
xor XOR2 (N10423, N10422, N9117);
not NOT1 (N10424, N10410);
and AND4 (N10425, N10421, N3259, N3369, N5405);
nand NAND2 (N10426, N10420, N261);
xor XOR2 (N10427, N10425, N4996);
nand NAND4 (N10428, N10412, N8831, N652, N9648);
xor XOR2 (N10429, N10403, N1744);
xor XOR2 (N10430, N10409, N4399);
or OR4 (N10431, N10426, N3986, N3971, N4828);
nand NAND2 (N10432, N10396, N1573);
or OR2 (N10433, N10429, N1841);
not NOT1 (N10434, N10431);
buf BUF1 (N10435, N10430);
not NOT1 (N10436, N10433);
buf BUF1 (N10437, N10423);
not NOT1 (N10438, N10434);
nand NAND3 (N10439, N10416, N6089, N10047);
not NOT1 (N10440, N10438);
or OR3 (N10441, N10424, N5356, N1848);
nand NAND2 (N10442, N10436, N313);
nor NOR2 (N10443, N10432, N639);
and AND4 (N10444, N10437, N1348, N5305, N9520);
not NOT1 (N10445, N10442);
or OR3 (N10446, N10443, N5032, N5418);
nand NAND3 (N10447, N10439, N3710, N7153);
or OR4 (N10448, N10415, N2950, N3725, N8321);
buf BUF1 (N10449, N10448);
or OR3 (N10450, N10447, N6394, N3160);
not NOT1 (N10451, N10450);
xor XOR2 (N10452, N10451, N7386);
nor NOR2 (N10453, N10435, N1615);
buf BUF1 (N10454, N10445);
nor NOR4 (N10455, N10454, N2037, N6728, N2621);
nor NOR2 (N10456, N10444, N386);
nand NAND4 (N10457, N10441, N3894, N2110, N7339);
and AND3 (N10458, N10449, N4614, N2778);
or OR3 (N10459, N10446, N4320, N6620);
and AND2 (N10460, N10427, N9380);
buf BUF1 (N10461, N10459);
and AND4 (N10462, N10453, N379, N9321, N4762);
and AND2 (N10463, N10428, N3820);
or OR2 (N10464, N10460, N1339);
not NOT1 (N10465, N10461);
buf BUF1 (N10466, N10464);
xor XOR2 (N10467, N10452, N3280);
not NOT1 (N10468, N10455);
or OR4 (N10469, N10463, N8928, N3945, N8250);
nand NAND3 (N10470, N10467, N8296, N7153);
nor NOR2 (N10471, N10440, N3919);
or OR3 (N10472, N10468, N1118, N7847);
buf BUF1 (N10473, N10469);
xor XOR2 (N10474, N10471, N6998);
and AND2 (N10475, N10473, N10229);
buf BUF1 (N10476, N10475);
not NOT1 (N10477, N10466);
or OR2 (N10478, N10462, N10428);
xor XOR2 (N10479, N10476, N4547);
nand NAND2 (N10480, N10470, N6227);
and AND2 (N10481, N10478, N3951);
not NOT1 (N10482, N10477);
xor XOR2 (N10483, N10481, N921);
buf BUF1 (N10484, N10474);
not NOT1 (N10485, N10483);
buf BUF1 (N10486, N10458);
or OR2 (N10487, N10480, N2656);
nor NOR4 (N10488, N10479, N3174, N9491, N2464);
buf BUF1 (N10489, N10456);
and AND3 (N10490, N10487, N4250, N8686);
or OR3 (N10491, N10490, N4887, N6445);
or OR3 (N10492, N10491, N5670, N9281);
xor XOR2 (N10493, N10484, N4244);
and AND2 (N10494, N10472, N7132);
buf BUF1 (N10495, N10488);
nor NOR3 (N10496, N10493, N2337, N6690);
and AND3 (N10497, N10486, N8204, N8878);
xor XOR2 (N10498, N10485, N7886);
buf BUF1 (N10499, N10496);
nor NOR4 (N10500, N10499, N9796, N485, N4710);
xor XOR2 (N10501, N10497, N2540);
nor NOR4 (N10502, N10494, N3430, N3068, N9811);
or OR3 (N10503, N10482, N1021, N2470);
xor XOR2 (N10504, N10465, N8405);
and AND2 (N10505, N10500, N8316);
nand NAND3 (N10506, N10502, N10078, N4480);
not NOT1 (N10507, N10498);
nor NOR2 (N10508, N10501, N7556);
buf BUF1 (N10509, N10505);
nor NOR2 (N10510, N10504, N10147);
or OR4 (N10511, N10510, N3732, N6513, N10021);
nand NAND4 (N10512, N10457, N2311, N5955, N9886);
nor NOR4 (N10513, N10511, N2841, N9700, N5602);
or OR3 (N10514, N10489, N9785, N8185);
nor NOR3 (N10515, N10514, N6706, N7404);
and AND2 (N10516, N10513, N2423);
nand NAND4 (N10517, N10512, N4022, N37, N9974);
and AND3 (N10518, N10517, N7568, N6434);
nor NOR2 (N10519, N10492, N6238);
buf BUF1 (N10520, N10495);
buf BUF1 (N10521, N10516);
or OR2 (N10522, N10503, N9732);
or OR3 (N10523, N10507, N8816, N8916);
or OR2 (N10524, N10506, N869);
and AND2 (N10525, N10515, N9846);
nor NOR4 (N10526, N10523, N2245, N10357, N4661);
xor XOR2 (N10527, N10519, N6984);
xor XOR2 (N10528, N10518, N2104);
or OR2 (N10529, N10508, N1658);
not NOT1 (N10530, N10528);
nand NAND4 (N10531, N10525, N6797, N8471, N1179);
xor XOR2 (N10532, N10531, N8728);
buf BUF1 (N10533, N10509);
buf BUF1 (N10534, N10530);
or OR3 (N10535, N10532, N2680, N3249);
nand NAND2 (N10536, N10520, N5730);
nand NAND4 (N10537, N10534, N9559, N3800, N7758);
or OR3 (N10538, N10524, N3387, N9307);
nand NAND2 (N10539, N10535, N8945);
or OR4 (N10540, N10538, N8042, N7101, N905);
buf BUF1 (N10541, N10537);
buf BUF1 (N10542, N10539);
nor NOR4 (N10543, N10526, N6742, N8050, N7514);
not NOT1 (N10544, N10527);
buf BUF1 (N10545, N10540);
nand NAND4 (N10546, N10543, N9089, N2540, N4947);
xor XOR2 (N10547, N10521, N6524);
nor NOR2 (N10548, N10544, N4707);
or OR3 (N10549, N10546, N6909, N4123);
nand NAND2 (N10550, N10542, N8863);
nor NOR3 (N10551, N10522, N7375, N3776);
buf BUF1 (N10552, N10529);
nor NOR4 (N10553, N10545, N8505, N1276, N10461);
not NOT1 (N10554, N10551);
or OR3 (N10555, N10552, N3923, N8299);
nor NOR4 (N10556, N10550, N3516, N7, N9489);
buf BUF1 (N10557, N10556);
nand NAND2 (N10558, N10555, N5477);
buf BUF1 (N10559, N10547);
nand NAND4 (N10560, N10553, N3283, N113, N9603);
nor NOR4 (N10561, N10533, N10395, N9011, N3325);
not NOT1 (N10562, N10560);
nor NOR2 (N10563, N10554, N8793);
nor NOR4 (N10564, N10561, N2741, N7071, N6675);
or OR2 (N10565, N10562, N10237);
nand NAND3 (N10566, N10549, N9958, N3259);
xor XOR2 (N10567, N10541, N73);
nor NOR3 (N10568, N10557, N6590, N4652);
not NOT1 (N10569, N10548);
nor NOR3 (N10570, N10558, N7709, N2496);
and AND4 (N10571, N10559, N9738, N3592, N2495);
xor XOR2 (N10572, N10569, N5020);
xor XOR2 (N10573, N10572, N6928);
nor NOR3 (N10574, N10563, N10314, N3356);
and AND4 (N10575, N10570, N118, N9212, N3639);
and AND3 (N10576, N10536, N1328, N9365);
or OR3 (N10577, N10575, N6283, N678);
nor NOR3 (N10578, N10564, N7139, N1075);
not NOT1 (N10579, N10565);
nor NOR3 (N10580, N10573, N5701, N9540);
nor NOR4 (N10581, N10568, N3361, N9077, N2304);
nor NOR3 (N10582, N10574, N782, N4692);
not NOT1 (N10583, N10576);
and AND4 (N10584, N10583, N7608, N2209, N7977);
nor NOR4 (N10585, N10571, N5085, N3411, N7971);
not NOT1 (N10586, N10582);
nor NOR4 (N10587, N10578, N8422, N9308, N5093);
or OR3 (N10588, N10567, N6715, N1681);
nor NOR4 (N10589, N10587, N8706, N4179, N3946);
buf BUF1 (N10590, N10581);
nor NOR4 (N10591, N10577, N9177, N2831, N834);
and AND4 (N10592, N10584, N7770, N4776, N5296);
nor NOR4 (N10593, N10586, N5601, N4184, N3108);
nand NAND2 (N10594, N10566, N9049);
nor NOR2 (N10595, N10593, N207);
and AND2 (N10596, N10589, N8615);
nor NOR4 (N10597, N10579, N7519, N9393, N8530);
buf BUF1 (N10598, N10580);
not NOT1 (N10599, N10595);
or OR2 (N10600, N10590, N8833);
nor NOR4 (N10601, N10598, N7315, N3384, N1359);
nor NOR3 (N10602, N10592, N10474, N1881);
nor NOR2 (N10603, N10601, N2771);
nand NAND4 (N10604, N10588, N4545, N2548, N4548);
buf BUF1 (N10605, N10600);
buf BUF1 (N10606, N10605);
nor NOR3 (N10607, N10597, N4642, N7398);
nor NOR3 (N10608, N10607, N1159, N8374);
not NOT1 (N10609, N10596);
nand NAND3 (N10610, N10594, N4015, N9781);
and AND3 (N10611, N10609, N5352, N6038);
xor XOR2 (N10612, N10606, N731);
nand NAND2 (N10613, N10608, N4051);
buf BUF1 (N10614, N10612);
and AND4 (N10615, N10611, N6804, N9903, N3819);
not NOT1 (N10616, N10599);
buf BUF1 (N10617, N10615);
xor XOR2 (N10618, N10604, N641);
or OR4 (N10619, N10613, N9262, N4006, N3329);
or OR2 (N10620, N10591, N986);
or OR4 (N10621, N10619, N6542, N10155, N2500);
and AND3 (N10622, N10585, N8112, N8205);
not NOT1 (N10623, N10602);
or OR3 (N10624, N10614, N7342, N3993);
xor XOR2 (N10625, N10618, N1432);
buf BUF1 (N10626, N10603);
xor XOR2 (N10627, N10620, N2596);
xor XOR2 (N10628, N10616, N1237);
xor XOR2 (N10629, N10626, N3078);
or OR4 (N10630, N10628, N8143, N517, N6395);
not NOT1 (N10631, N10624);
and AND4 (N10632, N10610, N7823, N3696, N255);
and AND3 (N10633, N10631, N6325, N4026);
xor XOR2 (N10634, N10622, N5661);
nand NAND4 (N10635, N10623, N3279, N10516, N51);
not NOT1 (N10636, N10633);
not NOT1 (N10637, N10627);
not NOT1 (N10638, N10621);
not NOT1 (N10639, N10625);
nor NOR4 (N10640, N10632, N10560, N8258, N2);
buf BUF1 (N10641, N10637);
nor NOR2 (N10642, N10617, N5279);
xor XOR2 (N10643, N10630, N6692);
or OR4 (N10644, N10638, N8763, N6240, N2336);
or OR3 (N10645, N10641, N415, N8199);
and AND4 (N10646, N10640, N5400, N7218, N6268);
and AND4 (N10647, N10635, N8019, N8777, N8736);
and AND4 (N10648, N10636, N10132, N332, N2622);
nor NOR2 (N10649, N10639, N3268);
xor XOR2 (N10650, N10642, N1808);
nor NOR4 (N10651, N10648, N2287, N379, N7485);
buf BUF1 (N10652, N10644);
and AND4 (N10653, N10643, N1371, N8741, N10634);
nand NAND3 (N10654, N9593, N2324, N4484);
or OR2 (N10655, N10647, N6505);
not NOT1 (N10656, N10645);
not NOT1 (N10657, N10629);
not NOT1 (N10658, N10646);
or OR4 (N10659, N10658, N4837, N5867, N2796);
and AND4 (N10660, N10657, N2602, N6984, N7508);
nor NOR3 (N10661, N10653, N5543, N516);
not NOT1 (N10662, N10654);
xor XOR2 (N10663, N10661, N5131);
nor NOR3 (N10664, N10660, N7593, N9840);
and AND2 (N10665, N10659, N8986);
nor NOR2 (N10666, N10664, N1364);
buf BUF1 (N10667, N10651);
nor NOR4 (N10668, N10656, N438, N3509, N7042);
and AND4 (N10669, N10668, N8679, N6014, N8730);
nand NAND3 (N10670, N10666, N8044, N6360);
and AND4 (N10671, N10650, N7171, N10348, N10082);
not NOT1 (N10672, N10665);
and AND3 (N10673, N10649, N164, N94);
not NOT1 (N10674, N10671);
buf BUF1 (N10675, N10673);
not NOT1 (N10676, N10652);
nand NAND3 (N10677, N10674, N31, N10183);
xor XOR2 (N10678, N10669, N8907);
xor XOR2 (N10679, N10667, N10338);
or OR3 (N10680, N10679, N81, N3800);
and AND3 (N10681, N10678, N7712, N821);
or OR2 (N10682, N10681, N3308);
or OR4 (N10683, N10655, N4771, N5511, N2914);
xor XOR2 (N10684, N10676, N9933);
and AND3 (N10685, N10682, N7126, N9564);
not NOT1 (N10686, N10672);
and AND2 (N10687, N10685, N8778);
buf BUF1 (N10688, N10675);
or OR4 (N10689, N10670, N10029, N6041, N6110);
buf BUF1 (N10690, N10688);
nand NAND3 (N10691, N10687, N189, N1700);
nor NOR3 (N10692, N10680, N5653, N9568);
nor NOR2 (N10693, N10662, N5628);
nand NAND2 (N10694, N10693, N7315);
nand NAND4 (N10695, N10689, N884, N2716, N2981);
nand NAND3 (N10696, N10677, N8687, N7437);
buf BUF1 (N10697, N10695);
or OR3 (N10698, N10697, N1161, N7889);
buf BUF1 (N10699, N10698);
or OR3 (N10700, N10692, N1238, N4815);
buf BUF1 (N10701, N10699);
and AND4 (N10702, N10691, N4271, N129, N6947);
or OR4 (N10703, N10686, N4917, N8105, N10277);
and AND2 (N10704, N10702, N2512);
or OR4 (N10705, N10690, N5983, N1308, N5794);
nand NAND3 (N10706, N10696, N4290, N9404);
not NOT1 (N10707, N10700);
and AND2 (N10708, N10701, N4291);
or OR2 (N10709, N10703, N4317);
nand NAND2 (N10710, N10709, N454);
not NOT1 (N10711, N10710);
xor XOR2 (N10712, N10706, N2550);
buf BUF1 (N10713, N10705);
buf BUF1 (N10714, N10713);
xor XOR2 (N10715, N10694, N2353);
and AND3 (N10716, N10708, N7151, N9505);
nor NOR2 (N10717, N10711, N4868);
nand NAND3 (N10718, N10714, N3446, N8183);
xor XOR2 (N10719, N10707, N5111);
nor NOR4 (N10720, N10716, N1550, N4551, N354);
or OR3 (N10721, N10712, N10669, N9951);
not NOT1 (N10722, N10717);
nand NAND2 (N10723, N10715, N7966);
buf BUF1 (N10724, N10722);
nand NAND4 (N10725, N10720, N1935, N1440, N2785);
buf BUF1 (N10726, N10719);
buf BUF1 (N10727, N10725);
and AND2 (N10728, N10704, N3744);
not NOT1 (N10729, N10727);
or OR2 (N10730, N10728, N5108);
nor NOR4 (N10731, N10684, N6516, N322, N3916);
and AND2 (N10732, N10724, N4523);
not NOT1 (N10733, N10683);
nor NOR3 (N10734, N10723, N9770, N3876);
or OR4 (N10735, N10663, N10114, N645, N4384);
and AND4 (N10736, N10721, N386, N5469, N5768);
or OR4 (N10737, N10731, N5053, N8, N5109);
buf BUF1 (N10738, N10729);
nor NOR2 (N10739, N10738, N9988);
buf BUF1 (N10740, N10733);
nor NOR2 (N10741, N10726, N3297);
nand NAND2 (N10742, N10734, N8876);
nor NOR2 (N10743, N10735, N2708);
xor XOR2 (N10744, N10737, N6319);
and AND3 (N10745, N10742, N10367, N5837);
nor NOR3 (N10746, N10730, N8038, N8467);
not NOT1 (N10747, N10740);
nand NAND2 (N10748, N10745, N3651);
or OR2 (N10749, N10747, N8028);
not NOT1 (N10750, N10718);
or OR4 (N10751, N10749, N2937, N5373, N3417);
buf BUF1 (N10752, N10744);
nand NAND4 (N10753, N10741, N3426, N5490, N7167);
nand NAND3 (N10754, N10750, N2091, N5901);
or OR3 (N10755, N10754, N8597, N7143);
and AND3 (N10756, N10732, N151, N8329);
buf BUF1 (N10757, N10753);
xor XOR2 (N10758, N10739, N5906);
buf BUF1 (N10759, N10746);
nor NOR4 (N10760, N10757, N539, N7878, N51);
not NOT1 (N10761, N10756);
and AND4 (N10762, N10759, N7587, N3413, N9740);
and AND2 (N10763, N10748, N6161);
nor NOR3 (N10764, N10743, N2029, N3644);
xor XOR2 (N10765, N10762, N7979);
buf BUF1 (N10766, N10751);
not NOT1 (N10767, N10736);
xor XOR2 (N10768, N10766, N5757);
and AND2 (N10769, N10752, N3722);
nand NAND4 (N10770, N10765, N8483, N379, N5545);
not NOT1 (N10771, N10758);
and AND3 (N10772, N10763, N1881, N2152);
xor XOR2 (N10773, N10767, N6335);
not NOT1 (N10774, N10772);
xor XOR2 (N10775, N10760, N9103);
nor NOR3 (N10776, N10768, N10453, N9142);
nor NOR4 (N10777, N10761, N9061, N8722, N2720);
buf BUF1 (N10778, N10769);
nor NOR2 (N10779, N10777, N3267);
buf BUF1 (N10780, N10778);
buf BUF1 (N10781, N10779);
or OR2 (N10782, N10764, N854);
xor XOR2 (N10783, N10780, N7733);
not NOT1 (N10784, N10770);
buf BUF1 (N10785, N10783);
nand NAND3 (N10786, N10782, N710, N3028);
buf BUF1 (N10787, N10775);
not NOT1 (N10788, N10773);
not NOT1 (N10789, N10785);
and AND3 (N10790, N10774, N2116, N5549);
xor XOR2 (N10791, N10784, N8577);
or OR2 (N10792, N10790, N4193);
or OR4 (N10793, N10776, N3232, N2748, N8445);
buf BUF1 (N10794, N10793);
nand NAND3 (N10795, N10791, N4388, N9082);
not NOT1 (N10796, N10795);
not NOT1 (N10797, N10792);
buf BUF1 (N10798, N10755);
and AND3 (N10799, N10788, N7778, N723);
nand NAND4 (N10800, N10781, N2315, N849, N7025);
or OR3 (N10801, N10800, N8459, N5505);
xor XOR2 (N10802, N10796, N3252);
and AND2 (N10803, N10789, N8880);
nor NOR2 (N10804, N10801, N241);
or OR2 (N10805, N10804, N275);
not NOT1 (N10806, N10805);
or OR3 (N10807, N10803, N3599, N8535);
buf BUF1 (N10808, N10806);
nand NAND2 (N10809, N10798, N3766);
nor NOR4 (N10810, N10809, N10088, N6256, N2867);
not NOT1 (N10811, N10786);
not NOT1 (N10812, N10811);
or OR4 (N10813, N10810, N8098, N332, N1372);
buf BUF1 (N10814, N10807);
nand NAND4 (N10815, N10814, N8223, N7907, N3195);
nor NOR4 (N10816, N10808, N7402, N5554, N6706);
and AND4 (N10817, N10816, N6994, N6444, N3143);
buf BUF1 (N10818, N10794);
nand NAND3 (N10819, N10815, N10294, N5427);
and AND4 (N10820, N10817, N587, N5056, N10037);
xor XOR2 (N10821, N10812, N327);
not NOT1 (N10822, N10821);
buf BUF1 (N10823, N10799);
nor NOR4 (N10824, N10818, N62, N10427, N6415);
or OR4 (N10825, N10787, N9848, N9483, N964);
buf BUF1 (N10826, N10819);
nand NAND4 (N10827, N10825, N10537, N651, N3892);
or OR3 (N10828, N10802, N673, N8065);
and AND4 (N10829, N10826, N4564, N1539, N1934);
or OR2 (N10830, N10813, N1589);
xor XOR2 (N10831, N10822, N92);
or OR2 (N10832, N10827, N8142);
buf BUF1 (N10833, N10829);
not NOT1 (N10834, N10823);
not NOT1 (N10835, N10831);
or OR3 (N10836, N10835, N8120, N7459);
nor NOR3 (N10837, N10828, N10422, N3950);
xor XOR2 (N10838, N10832, N3533);
nand NAND4 (N10839, N10830, N5607, N7613, N10505);
nand NAND2 (N10840, N10797, N4384);
xor XOR2 (N10841, N10820, N6829);
buf BUF1 (N10842, N10834);
or OR3 (N10843, N10840, N4045, N2926);
nand NAND3 (N10844, N10824, N8952, N6204);
buf BUF1 (N10845, N10842);
xor XOR2 (N10846, N10771, N1222);
nor NOR4 (N10847, N10838, N9861, N2385, N8515);
nor NOR4 (N10848, N10839, N621, N4397, N10048);
nor NOR3 (N10849, N10836, N3605, N10744);
nor NOR3 (N10850, N10848, N8728, N9231);
xor XOR2 (N10851, N10843, N5052);
and AND3 (N10852, N10850, N2462, N376);
not NOT1 (N10853, N10841);
nand NAND4 (N10854, N10847, N6202, N7052, N4094);
or OR2 (N10855, N10845, N2607);
and AND3 (N10856, N10844, N7159, N6764);
buf BUF1 (N10857, N10856);
nor NOR3 (N10858, N10855, N3530, N5691);
buf BUF1 (N10859, N10849);
and AND3 (N10860, N10853, N4360, N9835);
nand NAND3 (N10861, N10860, N2474, N6083);
xor XOR2 (N10862, N10846, N3341);
or OR2 (N10863, N10862, N813);
or OR3 (N10864, N10858, N5611, N9332);
and AND2 (N10865, N10864, N9773);
not NOT1 (N10866, N10863);
nand NAND3 (N10867, N10865, N8281, N3108);
xor XOR2 (N10868, N10851, N6106);
buf BUF1 (N10869, N10852);
or OR3 (N10870, N10854, N8143, N4224);
or OR3 (N10871, N10861, N6807, N6920);
nor NOR3 (N10872, N10871, N5876, N1225);
or OR2 (N10873, N10866, N5519);
nand NAND3 (N10874, N10868, N10536, N3481);
nand NAND3 (N10875, N10867, N7526, N9895);
not NOT1 (N10876, N10837);
xor XOR2 (N10877, N10875, N259);
not NOT1 (N10878, N10857);
not NOT1 (N10879, N10859);
and AND3 (N10880, N10879, N10303, N7563);
nand NAND2 (N10881, N10874, N6113);
nand NAND2 (N10882, N10872, N3699);
buf BUF1 (N10883, N10873);
buf BUF1 (N10884, N10880);
nor NOR3 (N10885, N10833, N9991, N9701);
nor NOR4 (N10886, N10881, N3534, N812, N4341);
xor XOR2 (N10887, N10876, N10723);
buf BUF1 (N10888, N10869);
not NOT1 (N10889, N10882);
buf BUF1 (N10890, N10877);
nand NAND2 (N10891, N10888, N8286);
and AND3 (N10892, N10890, N468, N2681);
and AND4 (N10893, N10892, N8525, N4567, N1374);
nor NOR4 (N10894, N10884, N4926, N854, N880);
nand NAND4 (N10895, N10883, N1985, N8353, N1116);
buf BUF1 (N10896, N10893);
xor XOR2 (N10897, N10896, N8204);
and AND2 (N10898, N10886, N3270);
and AND4 (N10899, N10894, N10784, N3761, N421);
xor XOR2 (N10900, N10899, N1174);
xor XOR2 (N10901, N10897, N4809);
buf BUF1 (N10902, N10901);
nand NAND4 (N10903, N10891, N5582, N3812, N5547);
or OR4 (N10904, N10887, N4643, N5585, N9170);
xor XOR2 (N10905, N10903, N258);
and AND3 (N10906, N10870, N4384, N9316);
not NOT1 (N10907, N10885);
buf BUF1 (N10908, N10905);
not NOT1 (N10909, N10895);
not NOT1 (N10910, N10909);
or OR3 (N10911, N10878, N6145, N2428);
buf BUF1 (N10912, N10904);
buf BUF1 (N10913, N10910);
xor XOR2 (N10914, N10900, N6436);
nor NOR2 (N10915, N10912, N1357);
not NOT1 (N10916, N10898);
buf BUF1 (N10917, N10911);
xor XOR2 (N10918, N10907, N6387);
xor XOR2 (N10919, N10915, N6732);
or OR2 (N10920, N10914, N10547);
buf BUF1 (N10921, N10902);
buf BUF1 (N10922, N10918);
or OR4 (N10923, N10917, N5666, N6343, N9248);
nand NAND3 (N10924, N10920, N10316, N4543);
buf BUF1 (N10925, N10913);
nor NOR2 (N10926, N10906, N6376);
buf BUF1 (N10927, N10924);
not NOT1 (N10928, N10927);
xor XOR2 (N10929, N10908, N1065);
and AND3 (N10930, N10925, N8118, N7534);
not NOT1 (N10931, N10928);
not NOT1 (N10932, N10919);
or OR2 (N10933, N10929, N6089);
and AND4 (N10934, N10921, N3365, N10109, N251);
not NOT1 (N10935, N10930);
xor XOR2 (N10936, N10926, N1572);
xor XOR2 (N10937, N10935, N3389);
nand NAND2 (N10938, N10936, N8200);
and AND3 (N10939, N10922, N5730, N2140);
and AND4 (N10940, N10938, N1859, N2735, N3783);
and AND3 (N10941, N10931, N9038, N5171);
nor NOR3 (N10942, N10889, N4762, N5226);
not NOT1 (N10943, N10916);
nand NAND2 (N10944, N10942, N1260);
nand NAND4 (N10945, N10937, N4404, N4431, N180);
not NOT1 (N10946, N10932);
buf BUF1 (N10947, N10945);
buf BUF1 (N10948, N10934);
not NOT1 (N10949, N10941);
and AND4 (N10950, N10923, N3459, N4058, N5741);
or OR4 (N10951, N10939, N3338, N757, N7992);
nor NOR4 (N10952, N10944, N4884, N4457, N8965);
nand NAND2 (N10953, N10949, N6096);
and AND3 (N10954, N10940, N8934, N10253);
or OR4 (N10955, N10951, N3339, N6510, N5584);
nand NAND3 (N10956, N10953, N955, N5600);
nand NAND4 (N10957, N10946, N2869, N10861, N10904);
buf BUF1 (N10958, N10948);
not NOT1 (N10959, N10957);
not NOT1 (N10960, N10954);
nor NOR4 (N10961, N10950, N8566, N9417, N415);
and AND2 (N10962, N10959, N7414);
and AND2 (N10963, N10952, N7618);
nor NOR3 (N10964, N10943, N8240, N510);
nor NOR3 (N10965, N10955, N2371, N5953);
buf BUF1 (N10966, N10947);
not NOT1 (N10967, N10958);
and AND2 (N10968, N10962, N7696);
or OR3 (N10969, N10960, N7629, N8817);
buf BUF1 (N10970, N10966);
buf BUF1 (N10971, N10963);
nand NAND2 (N10972, N10969, N4833);
nor NOR4 (N10973, N10972, N10579, N926, N1156);
and AND4 (N10974, N10965, N10365, N5487, N3260);
not NOT1 (N10975, N10973);
xor XOR2 (N10976, N10974, N10640);
not NOT1 (N10977, N10964);
nor NOR4 (N10978, N10977, N5468, N1263, N3876);
nand NAND4 (N10979, N10967, N7757, N2150, N9678);
xor XOR2 (N10980, N10970, N6113);
nor NOR4 (N10981, N10980, N1934, N5298, N2856);
xor XOR2 (N10982, N10981, N8539);
buf BUF1 (N10983, N10971);
nand NAND4 (N10984, N10933, N746, N3975, N40);
or OR4 (N10985, N10983, N2162, N4524, N5710);
or OR3 (N10986, N10985, N3519, N2253);
buf BUF1 (N10987, N10986);
and AND2 (N10988, N10979, N10253);
xor XOR2 (N10989, N10987, N5516);
buf BUF1 (N10990, N10956);
not NOT1 (N10991, N10982);
not NOT1 (N10992, N10984);
nand NAND3 (N10993, N10961, N8471, N3630);
or OR2 (N10994, N10976, N460);
buf BUF1 (N10995, N10994);
and AND3 (N10996, N10968, N2331, N7458);
xor XOR2 (N10997, N10995, N3836);
and AND4 (N10998, N10996, N10434, N10339, N3209);
or OR3 (N10999, N10978, N10170, N6738);
xor XOR2 (N11000, N10993, N4528);
nor NOR4 (N11001, N11000, N5119, N1457, N1348);
or OR4 (N11002, N10998, N9177, N5143, N892);
and AND3 (N11003, N10989, N6687, N1063);
or OR3 (N11004, N10975, N7229, N2886);
not NOT1 (N11005, N10991);
nor NOR3 (N11006, N10990, N8791, N864);
and AND3 (N11007, N10997, N1397, N4240);
buf BUF1 (N11008, N11007);
and AND2 (N11009, N11005, N6017);
nor NOR4 (N11010, N10992, N853, N1283, N762);
and AND3 (N11011, N10988, N278, N9332);
buf BUF1 (N11012, N10999);
or OR2 (N11013, N11009, N5813);
buf BUF1 (N11014, N11013);
not NOT1 (N11015, N11010);
nor NOR4 (N11016, N11006, N2297, N4107, N10752);
nor NOR3 (N11017, N11011, N6695, N1231);
or OR2 (N11018, N11017, N2692);
buf BUF1 (N11019, N11001);
and AND4 (N11020, N11014, N8844, N8041, N4717);
xor XOR2 (N11021, N11019, N8248);
nor NOR2 (N11022, N11004, N6716);
or OR4 (N11023, N11012, N10326, N8558, N382);
and AND3 (N11024, N11023, N6112, N1510);
buf BUF1 (N11025, N11020);
xor XOR2 (N11026, N11008, N9818);
nand NAND3 (N11027, N11024, N1824, N1993);
not NOT1 (N11028, N11018);
or OR4 (N11029, N11022, N10382, N6850, N4898);
buf BUF1 (N11030, N11016);
and AND2 (N11031, N11003, N1298);
buf BUF1 (N11032, N11027);
buf BUF1 (N11033, N11029);
buf BUF1 (N11034, N11031);
nand NAND2 (N11035, N11025, N10212);
nor NOR2 (N11036, N11026, N8372);
nand NAND2 (N11037, N11028, N5907);
nor NOR4 (N11038, N11035, N2795, N2669, N6900);
nand NAND3 (N11039, N11033, N755, N2447);
xor XOR2 (N11040, N11032, N4534);
not NOT1 (N11041, N11036);
and AND2 (N11042, N11038, N4494);
buf BUF1 (N11043, N11015);
not NOT1 (N11044, N11041);
or OR2 (N11045, N11034, N5525);
or OR3 (N11046, N11042, N2957, N5190);
buf BUF1 (N11047, N11037);
and AND3 (N11048, N11002, N8302, N7713);
buf BUF1 (N11049, N11043);
nor NOR4 (N11050, N11039, N10146, N6223, N8841);
and AND3 (N11051, N11045, N1606, N6443);
not NOT1 (N11052, N11046);
buf BUF1 (N11053, N11044);
xor XOR2 (N11054, N11040, N8430);
nor NOR2 (N11055, N11053, N7762);
xor XOR2 (N11056, N11030, N4872);
xor XOR2 (N11057, N11055, N2103);
nor NOR2 (N11058, N11021, N2144);
and AND2 (N11059, N11054, N5835);
and AND3 (N11060, N11057, N1199, N6659);
buf BUF1 (N11061, N11047);
xor XOR2 (N11062, N11048, N2668);
and AND2 (N11063, N11051, N1392);
not NOT1 (N11064, N11060);
buf BUF1 (N11065, N11064);
and AND4 (N11066, N11061, N8337, N7674, N4253);
and AND3 (N11067, N11052, N2798, N2758);
xor XOR2 (N11068, N11065, N2640);
nand NAND3 (N11069, N11058, N8543, N3887);
or OR4 (N11070, N11062, N9455, N6400, N1374);
xor XOR2 (N11071, N11059, N7778);
xor XOR2 (N11072, N11067, N8936);
or OR2 (N11073, N11071, N10458);
buf BUF1 (N11074, N11068);
and AND3 (N11075, N11050, N2374, N2976);
not NOT1 (N11076, N11056);
or OR3 (N11077, N11063, N5071, N8548);
nand NAND3 (N11078, N11077, N4565, N5747);
buf BUF1 (N11079, N11075);
nand NAND3 (N11080, N11072, N4415, N637);
xor XOR2 (N11081, N11078, N10921);
xor XOR2 (N11082, N11081, N6154);
buf BUF1 (N11083, N11080);
not NOT1 (N11084, N11049);
not NOT1 (N11085, N11074);
and AND4 (N11086, N11070, N2401, N9361, N2205);
and AND4 (N11087, N11069, N6124, N9680, N9741);
nand NAND2 (N11088, N11087, N5034);
xor XOR2 (N11089, N11066, N7912);
xor XOR2 (N11090, N11083, N2414);
xor XOR2 (N11091, N11088, N5336);
or OR4 (N11092, N11073, N2173, N6114, N4329);
nand NAND4 (N11093, N11086, N10467, N1023, N3651);
buf BUF1 (N11094, N11091);
or OR2 (N11095, N11089, N8169);
nand NAND3 (N11096, N11082, N3885, N7681);
buf BUF1 (N11097, N11090);
buf BUF1 (N11098, N11076);
xor XOR2 (N11099, N11096, N10181);
not NOT1 (N11100, N11093);
xor XOR2 (N11101, N11084, N2161);
and AND2 (N11102, N11101, N290);
nand NAND2 (N11103, N11097, N6843);
buf BUF1 (N11104, N11098);
nand NAND3 (N11105, N11104, N9989, N9686);
buf BUF1 (N11106, N11095);
not NOT1 (N11107, N11103);
not NOT1 (N11108, N11085);
or OR4 (N11109, N11107, N2409, N2026, N4524);
or OR3 (N11110, N11100, N5085, N8986);
and AND3 (N11111, N11079, N6292, N9944);
or OR4 (N11112, N11106, N9752, N7763, N600);
nor NOR3 (N11113, N11102, N6638, N6662);
or OR4 (N11114, N11110, N9909, N2837, N2961);
not NOT1 (N11115, N11113);
or OR4 (N11116, N11099, N1176, N8882, N4643);
nand NAND3 (N11117, N11105, N8493, N7286);
and AND3 (N11118, N11111, N10016, N9358);
buf BUF1 (N11119, N11118);
buf BUF1 (N11120, N11108);
or OR4 (N11121, N11117, N7418, N3168, N10924);
buf BUF1 (N11122, N11109);
xor XOR2 (N11123, N11112, N7063);
nand NAND3 (N11124, N11123, N3673, N9011);
nor NOR2 (N11125, N11114, N9985);
xor XOR2 (N11126, N11115, N546);
not NOT1 (N11127, N11120);
or OR3 (N11128, N11124, N8450, N8369);
nand NAND2 (N11129, N11127, N3091);
nand NAND3 (N11130, N11121, N5574, N5908);
xor XOR2 (N11131, N11130, N458);
xor XOR2 (N11132, N11131, N3274);
and AND2 (N11133, N11092, N2669);
nand NAND2 (N11134, N11133, N6931);
buf BUF1 (N11135, N11126);
nor NOR3 (N11136, N11122, N2932, N1482);
and AND4 (N11137, N11135, N4116, N159, N8626);
buf BUF1 (N11138, N11094);
xor XOR2 (N11139, N11129, N1396);
xor XOR2 (N11140, N11132, N10510);
buf BUF1 (N11141, N11128);
and AND4 (N11142, N11125, N7632, N4244, N10925);
buf BUF1 (N11143, N11119);
nand NAND3 (N11144, N11137, N1368, N4799);
buf BUF1 (N11145, N11139);
or OR2 (N11146, N11140, N10805);
or OR3 (N11147, N11138, N5998, N7415);
nor NOR4 (N11148, N11145, N9755, N3125, N8011);
buf BUF1 (N11149, N11136);
nand NAND3 (N11150, N11142, N8716, N5044);
not NOT1 (N11151, N11134);
buf BUF1 (N11152, N11148);
xor XOR2 (N11153, N11146, N4407);
not NOT1 (N11154, N11143);
not NOT1 (N11155, N11150);
or OR4 (N11156, N11151, N148, N8227, N1674);
nor NOR4 (N11157, N11154, N8244, N9179, N6035);
nand NAND4 (N11158, N11156, N10513, N5017, N3717);
xor XOR2 (N11159, N11155, N5857);
buf BUF1 (N11160, N11159);
nor NOR4 (N11161, N11153, N7768, N5491, N3119);
or OR4 (N11162, N11160, N416, N8793, N2488);
buf BUF1 (N11163, N11141);
buf BUF1 (N11164, N11162);
and AND4 (N11165, N11164, N1732, N7990, N6407);
and AND3 (N11166, N11158, N6789, N7891);
xor XOR2 (N11167, N11152, N1363);
nand NAND3 (N11168, N11165, N10886, N4068);
nor NOR4 (N11169, N11149, N5129, N6913, N4913);
and AND4 (N11170, N11168, N2305, N2471, N2820);
nor NOR4 (N11171, N11163, N4441, N6903, N537);
nand NAND3 (N11172, N11161, N3585, N6981);
xor XOR2 (N11173, N11157, N6588);
not NOT1 (N11174, N11172);
nor NOR2 (N11175, N11144, N7321);
nor NOR3 (N11176, N11169, N1956, N8764);
buf BUF1 (N11177, N11116);
buf BUF1 (N11178, N11175);
nand NAND2 (N11179, N11171, N4829);
buf BUF1 (N11180, N11177);
nor NOR3 (N11181, N11176, N2010, N429);
or OR3 (N11182, N11178, N748, N9884);
or OR3 (N11183, N11166, N10760, N4710);
or OR4 (N11184, N11180, N3454, N2945, N832);
buf BUF1 (N11185, N11179);
xor XOR2 (N11186, N11173, N4639);
or OR4 (N11187, N11182, N9915, N424, N453);
or OR3 (N11188, N11185, N1625, N9170);
and AND3 (N11189, N11186, N7530, N5295);
nor NOR3 (N11190, N11184, N4016, N10764);
and AND3 (N11191, N11147, N6889, N1822);
nand NAND4 (N11192, N11191, N3998, N3898, N2817);
or OR3 (N11193, N11187, N3858, N8217);
buf BUF1 (N11194, N11188);
buf BUF1 (N11195, N11170);
or OR3 (N11196, N11195, N9319, N8501);
or OR3 (N11197, N11189, N8012, N10754);
and AND4 (N11198, N11196, N581, N8869, N8066);
and AND3 (N11199, N11190, N8233, N10787);
buf BUF1 (N11200, N11167);
and AND4 (N11201, N11174, N10139, N6624, N2722);
buf BUF1 (N11202, N11198);
and AND2 (N11203, N11197, N10655);
or OR2 (N11204, N11199, N4169);
nand NAND2 (N11205, N11204, N10819);
or OR2 (N11206, N11205, N8421);
xor XOR2 (N11207, N11201, N6990);
xor XOR2 (N11208, N11206, N484);
nor NOR4 (N11209, N11181, N3285, N8955, N976);
nand NAND4 (N11210, N11193, N7563, N4604, N3642);
or OR2 (N11211, N11203, N2303);
nand NAND4 (N11212, N11202, N7794, N2360, N1082);
buf BUF1 (N11213, N11194);
buf BUF1 (N11214, N11200);
buf BUF1 (N11215, N11208);
and AND3 (N11216, N11207, N7943, N343);
not NOT1 (N11217, N11192);
or OR4 (N11218, N11217, N4151, N9061, N2588);
xor XOR2 (N11219, N11214, N8246);
and AND4 (N11220, N11219, N10082, N9899, N10152);
buf BUF1 (N11221, N11210);
buf BUF1 (N11222, N11216);
not NOT1 (N11223, N11209);
not NOT1 (N11224, N11212);
xor XOR2 (N11225, N11215, N3932);
and AND2 (N11226, N11225, N8018);
and AND4 (N11227, N11213, N5409, N7340, N3590);
xor XOR2 (N11228, N11183, N652);
nor NOR2 (N11229, N11226, N2686);
or OR4 (N11230, N11228, N10519, N1892, N7249);
and AND2 (N11231, N11229, N8310);
or OR2 (N11232, N11220, N1947);
buf BUF1 (N11233, N11231);
or OR3 (N11234, N11232, N4121, N341);
buf BUF1 (N11235, N11221);
or OR2 (N11236, N11234, N2747);
not NOT1 (N11237, N11227);
nor NOR3 (N11238, N11218, N9255, N9721);
not NOT1 (N11239, N11224);
not NOT1 (N11240, N11237);
buf BUF1 (N11241, N11238);
and AND3 (N11242, N11211, N3984, N8052);
xor XOR2 (N11243, N11236, N2607);
and AND2 (N11244, N11230, N8551);
not NOT1 (N11245, N11244);
xor XOR2 (N11246, N11239, N9774);
or OR4 (N11247, N11233, N6134, N2468, N7885);
nand NAND2 (N11248, N11223, N9828);
nor NOR3 (N11249, N11246, N9695, N8555);
or OR4 (N11250, N11245, N7033, N3294, N7527);
buf BUF1 (N11251, N11235);
buf BUF1 (N11252, N11249);
buf BUF1 (N11253, N11250);
nor NOR4 (N11254, N11253, N4753, N5749, N4244);
xor XOR2 (N11255, N11252, N10306);
or OR2 (N11256, N11240, N1803);
or OR4 (N11257, N11251, N1399, N6768, N2536);
and AND2 (N11258, N11254, N7440);
or OR3 (N11259, N11241, N318, N3584);
xor XOR2 (N11260, N11243, N6404);
xor XOR2 (N11261, N11259, N10232);
nor NOR2 (N11262, N11242, N3773);
xor XOR2 (N11263, N11258, N7462);
or OR2 (N11264, N11257, N4978);
xor XOR2 (N11265, N11261, N5181);
xor XOR2 (N11266, N11247, N9814);
or OR3 (N11267, N11263, N6836, N1977);
and AND2 (N11268, N11260, N4921);
and AND2 (N11269, N11266, N8793);
or OR3 (N11270, N11265, N5173, N1406);
nor NOR2 (N11271, N11268, N622);
buf BUF1 (N11272, N11262);
buf BUF1 (N11273, N11271);
buf BUF1 (N11274, N11222);
nand NAND4 (N11275, N11270, N1541, N9106, N6764);
nand NAND2 (N11276, N11255, N432);
or OR3 (N11277, N11274, N1984, N5495);
or OR4 (N11278, N11276, N7544, N7304, N4953);
nand NAND2 (N11279, N11278, N5182);
xor XOR2 (N11280, N11248, N6181);
nor NOR4 (N11281, N11275, N2876, N2529, N3480);
and AND4 (N11282, N11264, N8208, N1898, N9107);
nor NOR3 (N11283, N11256, N289, N9530);
nand NAND2 (N11284, N11269, N6886);
xor XOR2 (N11285, N11281, N1003);
nor NOR2 (N11286, N11273, N8773);
buf BUF1 (N11287, N11283);
buf BUF1 (N11288, N11282);
not NOT1 (N11289, N11284);
and AND3 (N11290, N11286, N4299, N2875);
xor XOR2 (N11291, N11288, N7058);
nor NOR3 (N11292, N11289, N4515, N6745);
not NOT1 (N11293, N11272);
nand NAND2 (N11294, N11290, N5005);
or OR3 (N11295, N11293, N5709, N8556);
nand NAND2 (N11296, N11291, N1297);
nand NAND2 (N11297, N11287, N9815);
and AND3 (N11298, N11279, N5415, N7811);
xor XOR2 (N11299, N11298, N7752);
buf BUF1 (N11300, N11296);
buf BUF1 (N11301, N11300);
nand NAND2 (N11302, N11294, N9234);
nand NAND2 (N11303, N11299, N9038);
xor XOR2 (N11304, N11295, N5793);
nand NAND4 (N11305, N11280, N3293, N6636, N4541);
xor XOR2 (N11306, N11302, N6698);
and AND2 (N11307, N11292, N10499);
and AND3 (N11308, N11267, N3432, N9234);
not NOT1 (N11309, N11303);
and AND2 (N11310, N11304, N3435);
nor NOR2 (N11311, N11308, N5180);
buf BUF1 (N11312, N11306);
xor XOR2 (N11313, N11310, N9278);
nor NOR3 (N11314, N11307, N3931, N6330);
nor NOR3 (N11315, N11301, N7402, N5346);
and AND4 (N11316, N11309, N680, N96, N11017);
not NOT1 (N11317, N11316);
nand NAND4 (N11318, N11311, N9153, N5901, N6521);
not NOT1 (N11319, N11297);
not NOT1 (N11320, N11318);
or OR2 (N11321, N11317, N97);
nor NOR2 (N11322, N11277, N9528);
xor XOR2 (N11323, N11313, N7106);
nand NAND3 (N11324, N11320, N5489, N10032);
not NOT1 (N11325, N11285);
xor XOR2 (N11326, N11315, N2491);
buf BUF1 (N11327, N11322);
nor NOR2 (N11328, N11314, N7239);
or OR4 (N11329, N11327, N5186, N3746, N8757);
not NOT1 (N11330, N11326);
nor NOR2 (N11331, N11330, N2635);
and AND4 (N11332, N11321, N2302, N8258, N2129);
and AND3 (N11333, N11312, N8920, N10089);
not NOT1 (N11334, N11331);
buf BUF1 (N11335, N11319);
or OR4 (N11336, N11325, N4076, N6913, N3625);
xor XOR2 (N11337, N11328, N7680);
nor NOR4 (N11338, N11335, N6373, N9073, N6186);
and AND2 (N11339, N11334, N5871);
nor NOR4 (N11340, N11324, N8705, N1977, N7498);
or OR3 (N11341, N11336, N219, N1102);
buf BUF1 (N11342, N11338);
buf BUF1 (N11343, N11305);
xor XOR2 (N11344, N11341, N9405);
or OR3 (N11345, N11343, N2860, N6666);
or OR4 (N11346, N11332, N648, N4334, N5442);
nand NAND4 (N11347, N11346, N9821, N6072, N3395);
or OR3 (N11348, N11344, N5280, N9538);
nor NOR3 (N11349, N11345, N4094, N8617);
xor XOR2 (N11350, N11337, N3812);
nand NAND2 (N11351, N11347, N7372);
nand NAND2 (N11352, N11349, N3565);
buf BUF1 (N11353, N11350);
or OR2 (N11354, N11333, N3962);
or OR3 (N11355, N11329, N7814, N1278);
xor XOR2 (N11356, N11352, N1195);
nor NOR4 (N11357, N11356, N2246, N6734, N4572);
or OR4 (N11358, N11355, N5393, N1597, N7300);
nor NOR2 (N11359, N11358, N2942);
buf BUF1 (N11360, N11323);
not NOT1 (N11361, N11340);
and AND4 (N11362, N11339, N10627, N2487, N11153);
not NOT1 (N11363, N11357);
xor XOR2 (N11364, N11360, N7898);
xor XOR2 (N11365, N11348, N4860);
nor NOR2 (N11366, N11362, N11302);
nor NOR4 (N11367, N11354, N7189, N5343, N4673);
not NOT1 (N11368, N11361);
nor NOR2 (N11369, N11353, N1666);
buf BUF1 (N11370, N11365);
xor XOR2 (N11371, N11367, N10357);
or OR4 (N11372, N11363, N1103, N2193, N1428);
buf BUF1 (N11373, N11370);
nor NOR3 (N11374, N11372, N1794, N2703);
nor NOR4 (N11375, N11364, N10315, N7769, N6364);
nor NOR2 (N11376, N11369, N11258);
not NOT1 (N11377, N11342);
buf BUF1 (N11378, N11374);
nand NAND3 (N11379, N11366, N3015, N3174);
not NOT1 (N11380, N11377);
nor NOR2 (N11381, N11380, N8105);
or OR3 (N11382, N11371, N2782, N4939);
xor XOR2 (N11383, N11378, N5043);
nand NAND4 (N11384, N11359, N10776, N5680, N6326);
nor NOR2 (N11385, N11351, N4417);
nor NOR3 (N11386, N11376, N10504, N3449);
buf BUF1 (N11387, N11368);
and AND4 (N11388, N11386, N1409, N2662, N9737);
not NOT1 (N11389, N11379);
and AND4 (N11390, N11385, N1051, N2670, N3812);
or OR4 (N11391, N11381, N9165, N6246, N6113);
xor XOR2 (N11392, N11390, N8699);
nand NAND2 (N11393, N11391, N3003);
nand NAND2 (N11394, N11382, N541);
not NOT1 (N11395, N11393);
nand NAND3 (N11396, N11389, N8129, N5183);
nand NAND4 (N11397, N11387, N7668, N828, N9144);
not NOT1 (N11398, N11395);
or OR4 (N11399, N11375, N7770, N2000, N8333);
xor XOR2 (N11400, N11392, N266);
xor XOR2 (N11401, N11394, N4660);
and AND3 (N11402, N11397, N7974, N5811);
or OR3 (N11403, N11399, N11292, N9365);
not NOT1 (N11404, N11403);
or OR3 (N11405, N11400, N7276, N1356);
buf BUF1 (N11406, N11402);
and AND2 (N11407, N11401, N7500);
buf BUF1 (N11408, N11373);
not NOT1 (N11409, N11384);
or OR2 (N11410, N11404, N10248);
nand NAND2 (N11411, N11396, N1493);
and AND4 (N11412, N11409, N7825, N2947, N7356);
xor XOR2 (N11413, N11411, N9168);
nand NAND2 (N11414, N11413, N3175);
not NOT1 (N11415, N11407);
xor XOR2 (N11416, N11415, N7592);
xor XOR2 (N11417, N11406, N1226);
and AND3 (N11418, N11410, N4485, N3929);
nand NAND2 (N11419, N11388, N3132);
nor NOR3 (N11420, N11418, N7846, N9990);
xor XOR2 (N11421, N11416, N4065);
not NOT1 (N11422, N11414);
xor XOR2 (N11423, N11398, N2199);
nor NOR3 (N11424, N11419, N11144, N2175);
or OR3 (N11425, N11412, N3602, N5626);
and AND2 (N11426, N11408, N3013);
buf BUF1 (N11427, N11423);
xor XOR2 (N11428, N11383, N11205);
or OR2 (N11429, N11428, N5767);
nor NOR2 (N11430, N11420, N1393);
nor NOR2 (N11431, N11421, N10481);
xor XOR2 (N11432, N11427, N7295);
or OR2 (N11433, N11431, N773);
nand NAND3 (N11434, N11424, N5586, N8115);
xor XOR2 (N11435, N11433, N7988);
and AND4 (N11436, N11434, N7644, N306, N899);
not NOT1 (N11437, N11436);
buf BUF1 (N11438, N11422);
and AND4 (N11439, N11425, N3781, N10631, N8595);
xor XOR2 (N11440, N11439, N498);
and AND4 (N11441, N11429, N3308, N5952, N10327);
or OR3 (N11442, N11405, N3735, N3597);
nand NAND2 (N11443, N11432, N4252);
or OR4 (N11444, N11417, N4940, N5520, N9662);
buf BUF1 (N11445, N11430);
nor NOR3 (N11446, N11435, N1825, N7524);
nand NAND4 (N11447, N11438, N4382, N2840, N8425);
or OR2 (N11448, N11440, N8217);
or OR3 (N11449, N11444, N7564, N10123);
or OR4 (N11450, N11448, N3313, N1153, N4152);
or OR2 (N11451, N11441, N2728);
nand NAND4 (N11452, N11426, N3894, N1552, N4334);
xor XOR2 (N11453, N11451, N9997);
nand NAND3 (N11454, N11445, N5975, N5684);
or OR2 (N11455, N11446, N3285);
xor XOR2 (N11456, N11452, N1158);
xor XOR2 (N11457, N11453, N2327);
or OR4 (N11458, N11437, N5066, N6683, N6644);
and AND3 (N11459, N11457, N4931, N4869);
buf BUF1 (N11460, N11458);
xor XOR2 (N11461, N11450, N8877);
not NOT1 (N11462, N11447);
buf BUF1 (N11463, N11455);
not NOT1 (N11464, N11460);
buf BUF1 (N11465, N11462);
or OR4 (N11466, N11449, N2705, N6240, N7283);
xor XOR2 (N11467, N11461, N3434);
or OR4 (N11468, N11456, N10457, N9602, N1286);
nand NAND4 (N11469, N11464, N752, N10705, N726);
not NOT1 (N11470, N11459);
and AND3 (N11471, N11465, N7939, N8205);
not NOT1 (N11472, N11443);
or OR2 (N11473, N11442, N1959);
xor XOR2 (N11474, N11472, N1195);
and AND4 (N11475, N11466, N1677, N8598, N3106);
buf BUF1 (N11476, N11468);
not NOT1 (N11477, N11463);
xor XOR2 (N11478, N11475, N6054);
or OR2 (N11479, N11454, N1156);
not NOT1 (N11480, N11470);
buf BUF1 (N11481, N11474);
buf BUF1 (N11482, N11469);
nor NOR3 (N11483, N11481, N7466, N2673);
nor NOR3 (N11484, N11473, N9653, N1875);
nor NOR3 (N11485, N11480, N7469, N10691);
not NOT1 (N11486, N11484);
or OR2 (N11487, N11486, N10532);
buf BUF1 (N11488, N11479);
nand NAND3 (N11489, N11483, N7488, N7664);
or OR3 (N11490, N11485, N4894, N948);
xor XOR2 (N11491, N11489, N9499);
nor NOR3 (N11492, N11488, N4271, N798);
nand NAND2 (N11493, N11482, N4827);
and AND4 (N11494, N11491, N10371, N7160, N7394);
xor XOR2 (N11495, N11493, N1929);
nand NAND2 (N11496, N11471, N1);
nor NOR3 (N11497, N11492, N8268, N11015);
xor XOR2 (N11498, N11490, N10621);
buf BUF1 (N11499, N11496);
or OR4 (N11500, N11487, N2406, N7274, N7195);
xor XOR2 (N11501, N11500, N6922);
nand NAND4 (N11502, N11497, N2459, N98, N3566);
or OR2 (N11503, N11502, N6858);
and AND3 (N11504, N11501, N1906, N5443);
nor NOR4 (N11505, N11495, N2384, N10095, N4490);
not NOT1 (N11506, N11476);
nor NOR2 (N11507, N11506, N5297);
not NOT1 (N11508, N11504);
and AND4 (N11509, N11503, N8870, N10043, N4096);
and AND4 (N11510, N11505, N1273, N6334, N5509);
or OR3 (N11511, N11509, N8004, N227);
and AND3 (N11512, N11478, N7464, N342);
nor NOR3 (N11513, N11494, N7000, N7919);
xor XOR2 (N11514, N11498, N8121);
and AND3 (N11515, N11467, N7354, N1629);
xor XOR2 (N11516, N11513, N7797);
and AND2 (N11517, N11514, N3845);
nor NOR4 (N11518, N11511, N10747, N10962, N3434);
nor NOR3 (N11519, N11477, N11199, N3312);
nand NAND4 (N11520, N11510, N342, N7874, N3781);
and AND3 (N11521, N11517, N7680, N8196);
not NOT1 (N11522, N11499);
xor XOR2 (N11523, N11521, N10163);
or OR4 (N11524, N11508, N4074, N4436, N1680);
xor XOR2 (N11525, N11515, N4778);
not NOT1 (N11526, N11516);
not NOT1 (N11527, N11507);
buf BUF1 (N11528, N11524);
not NOT1 (N11529, N11518);
or OR2 (N11530, N11512, N9722);
nand NAND4 (N11531, N11527, N2218, N8885, N4754);
and AND4 (N11532, N11531, N182, N10749, N8984);
and AND3 (N11533, N11525, N4582, N8130);
nand NAND3 (N11534, N11530, N2095, N5061);
not NOT1 (N11535, N11533);
buf BUF1 (N11536, N11529);
buf BUF1 (N11537, N11523);
xor XOR2 (N11538, N11534, N10384);
not NOT1 (N11539, N11522);
and AND2 (N11540, N11535, N10175);
nor NOR2 (N11541, N11532, N356);
xor XOR2 (N11542, N11540, N5665);
and AND3 (N11543, N11520, N9452, N6165);
and AND2 (N11544, N11538, N9150);
and AND4 (N11545, N11541, N5187, N4946, N1195);
xor XOR2 (N11546, N11526, N2281);
nand NAND2 (N11547, N11545, N11092);
and AND3 (N11548, N11543, N3175, N7971);
buf BUF1 (N11549, N11539);
or OR4 (N11550, N11519, N4411, N8812, N4679);
and AND2 (N11551, N11528, N287);
nor NOR2 (N11552, N11544, N6466);
nor NOR4 (N11553, N11552, N8702, N8124, N6393);
nor NOR4 (N11554, N11537, N262, N5585, N7705);
not NOT1 (N11555, N11549);
not NOT1 (N11556, N11553);
nand NAND3 (N11557, N11547, N11151, N869);
xor XOR2 (N11558, N11546, N7624);
and AND2 (N11559, N11557, N11112);
and AND3 (N11560, N11558, N7381, N1089);
xor XOR2 (N11561, N11560, N4484);
or OR4 (N11562, N11556, N10470, N9846, N10008);
xor XOR2 (N11563, N11555, N5674);
buf BUF1 (N11564, N11561);
nor NOR3 (N11565, N11563, N264, N9423);
nor NOR2 (N11566, N11551, N7069);
not NOT1 (N11567, N11562);
nor NOR4 (N11568, N11554, N294, N11034, N4488);
and AND3 (N11569, N11548, N2543, N6586);
or OR2 (N11570, N11542, N5907);
and AND4 (N11571, N11570, N2573, N11298, N2095);
nor NOR4 (N11572, N11566, N8636, N6110, N11058);
not NOT1 (N11573, N11536);
nand NAND2 (N11574, N11568, N7511);
and AND4 (N11575, N11567, N9870, N737, N1588);
buf BUF1 (N11576, N11574);
nor NOR4 (N11577, N11550, N6451, N8766, N7677);
not NOT1 (N11578, N11559);
nand NAND2 (N11579, N11573, N7285);
nand NAND4 (N11580, N11577, N3693, N6606, N366);
xor XOR2 (N11581, N11564, N7525);
xor XOR2 (N11582, N11578, N4113);
xor XOR2 (N11583, N11580, N9681);
nand NAND4 (N11584, N11582, N8198, N3828, N4070);
buf BUF1 (N11585, N11575);
and AND2 (N11586, N11571, N11349);
not NOT1 (N11587, N11585);
buf BUF1 (N11588, N11565);
not NOT1 (N11589, N11586);
and AND4 (N11590, N11584, N3966, N3749, N10479);
and AND3 (N11591, N11569, N6863, N2027);
nor NOR3 (N11592, N11581, N4593, N9358);
buf BUF1 (N11593, N11587);
nand NAND2 (N11594, N11592, N7154);
or OR2 (N11595, N11572, N417);
and AND4 (N11596, N11593, N7838, N4399, N9449);
xor XOR2 (N11597, N11579, N11596);
and AND2 (N11598, N3386, N4796);
and AND4 (N11599, N11597, N4664, N3565, N7591);
xor XOR2 (N11600, N11598, N9439);
buf BUF1 (N11601, N11595);
xor XOR2 (N11602, N11601, N1613);
buf BUF1 (N11603, N11589);
and AND4 (N11604, N11594, N5287, N7067, N3944);
nand NAND4 (N11605, N11588, N7548, N8489, N9577);
or OR3 (N11606, N11602, N4779, N5173);
xor XOR2 (N11607, N11599, N3489);
nand NAND3 (N11608, N11606, N2974, N1995);
not NOT1 (N11609, N11605);
buf BUF1 (N11610, N11576);
buf BUF1 (N11611, N11600);
nor NOR2 (N11612, N11611, N2725);
buf BUF1 (N11613, N11610);
nor NOR2 (N11614, N11591, N1695);
xor XOR2 (N11615, N11607, N8370);
or OR4 (N11616, N11613, N8936, N10465, N5409);
or OR2 (N11617, N11612, N2098);
or OR2 (N11618, N11590, N9887);
xor XOR2 (N11619, N11583, N10557);
xor XOR2 (N11620, N11619, N3743);
buf BUF1 (N11621, N11620);
and AND3 (N11622, N11608, N3640, N4122);
nor NOR2 (N11623, N11618, N1511);
or OR4 (N11624, N11617, N4246, N4756, N2682);
not NOT1 (N11625, N11621);
nand NAND2 (N11626, N11609, N4908);
nand NAND2 (N11627, N11604, N809);
and AND4 (N11628, N11616, N941, N8260, N8144);
buf BUF1 (N11629, N11623);
not NOT1 (N11630, N11625);
not NOT1 (N11631, N11603);
and AND2 (N11632, N11629, N11005);
buf BUF1 (N11633, N11627);
and AND4 (N11634, N11630, N5881, N10081, N2780);
or OR3 (N11635, N11624, N8948, N1121);
nor NOR3 (N11636, N11634, N9901, N9123);
or OR4 (N11637, N11614, N11380, N7849, N1131);
and AND2 (N11638, N11615, N1345);
buf BUF1 (N11639, N11636);
or OR2 (N11640, N11637, N4981);
nand NAND3 (N11641, N11639, N6522, N5497);
nor NOR2 (N11642, N11632, N6426);
or OR2 (N11643, N11628, N2118);
buf BUF1 (N11644, N11638);
xor XOR2 (N11645, N11622, N10834);
nor NOR3 (N11646, N11644, N1776, N4644);
or OR4 (N11647, N11646, N853, N10317, N6712);
nor NOR2 (N11648, N11626, N797);
and AND2 (N11649, N11643, N9566);
or OR3 (N11650, N11645, N5961, N1514);
xor XOR2 (N11651, N11647, N3347);
not NOT1 (N11652, N11651);
nand NAND2 (N11653, N11650, N970);
or OR3 (N11654, N11653, N6050, N2835);
nand NAND3 (N11655, N11631, N4041, N6239);
xor XOR2 (N11656, N11633, N2410);
nor NOR4 (N11657, N11652, N4890, N4093, N8622);
nand NAND2 (N11658, N11649, N10803);
xor XOR2 (N11659, N11635, N9848);
nand NAND4 (N11660, N11656, N933, N6613, N538);
not NOT1 (N11661, N11641);
nand NAND2 (N11662, N11659, N7234);
and AND3 (N11663, N11642, N2828, N7081);
nand NAND2 (N11664, N11663, N219);
buf BUF1 (N11665, N11662);
or OR2 (N11666, N11660, N10949);
nor NOR2 (N11667, N11666, N4382);
buf BUF1 (N11668, N11664);
not NOT1 (N11669, N11661);
nand NAND4 (N11670, N11669, N55, N5151, N10385);
or OR2 (N11671, N11655, N8705);
not NOT1 (N11672, N11657);
and AND2 (N11673, N11658, N5682);
or OR3 (N11674, N11654, N1938, N10585);
xor XOR2 (N11675, N11674, N10987);
or OR3 (N11676, N11648, N4164, N1404);
xor XOR2 (N11677, N11670, N8504);
xor XOR2 (N11678, N11640, N6476);
nor NOR2 (N11679, N11668, N1743);
or OR3 (N11680, N11676, N9300, N3224);
xor XOR2 (N11681, N11665, N4697);
not NOT1 (N11682, N11681);
nor NOR2 (N11683, N11673, N9780);
nand NAND4 (N11684, N11667, N5627, N6905, N5294);
nor NOR3 (N11685, N11677, N4390, N9565);
not NOT1 (N11686, N11683);
xor XOR2 (N11687, N11672, N10949);
and AND2 (N11688, N11686, N11321);
not NOT1 (N11689, N11679);
xor XOR2 (N11690, N11689, N2831);
not NOT1 (N11691, N11678);
xor XOR2 (N11692, N11684, N11575);
nand NAND4 (N11693, N11675, N6042, N10333, N1838);
nor NOR4 (N11694, N11687, N1695, N647, N10635);
buf BUF1 (N11695, N11694);
nand NAND4 (N11696, N11690, N6810, N6218, N556);
nor NOR2 (N11697, N11691, N7445);
and AND2 (N11698, N11695, N429);
buf BUF1 (N11699, N11671);
nand NAND4 (N11700, N11698, N10834, N1329, N6582);
buf BUF1 (N11701, N11699);
not NOT1 (N11702, N11688);
or OR2 (N11703, N11693, N8527);
nand NAND4 (N11704, N11703, N104, N8621, N2744);
nor NOR2 (N11705, N11692, N7201);
not NOT1 (N11706, N11682);
xor XOR2 (N11707, N11704, N8151);
buf BUF1 (N11708, N11702);
nand NAND4 (N11709, N11696, N3162, N10404, N4041);
nor NOR3 (N11710, N11705, N10314, N10318);
nand NAND3 (N11711, N11685, N5080, N2205);
nand NAND3 (N11712, N11711, N9253, N937);
nand NAND4 (N11713, N11710, N7625, N11425, N6853);
not NOT1 (N11714, N11701);
xor XOR2 (N11715, N11707, N8358);
not NOT1 (N11716, N11708);
xor XOR2 (N11717, N11716, N7890);
not NOT1 (N11718, N11712);
nand NAND4 (N11719, N11706, N420, N4722, N1174);
nor NOR2 (N11720, N11713, N6593);
not NOT1 (N11721, N11697);
or OR4 (N11722, N11680, N2236, N7047, N9231);
xor XOR2 (N11723, N11714, N6583);
nand NAND2 (N11724, N11722, N2194);
xor XOR2 (N11725, N11719, N710);
and AND3 (N11726, N11721, N7625, N984);
and AND2 (N11727, N11709, N2936);
nand NAND4 (N11728, N11727, N8110, N9269, N1719);
or OR2 (N11729, N11720, N5062);
and AND3 (N11730, N11726, N9217, N623);
or OR2 (N11731, N11730, N4469);
and AND2 (N11732, N11700, N1135);
not NOT1 (N11733, N11724);
not NOT1 (N11734, N11717);
or OR3 (N11735, N11723, N10314, N11157);
nand NAND4 (N11736, N11718, N8251, N5011, N4928);
and AND3 (N11737, N11731, N1646, N9274);
xor XOR2 (N11738, N11737, N6022);
nor NOR3 (N11739, N11729, N2790, N3004);
buf BUF1 (N11740, N11738);
not NOT1 (N11741, N11728);
buf BUF1 (N11742, N11741);
not NOT1 (N11743, N11742);
buf BUF1 (N11744, N11715);
not NOT1 (N11745, N11735);
buf BUF1 (N11746, N11739);
or OR2 (N11747, N11736, N5546);
nor NOR4 (N11748, N11734, N1567, N7601, N6730);
nand NAND3 (N11749, N11733, N4915, N3673);
buf BUF1 (N11750, N11749);
buf BUF1 (N11751, N11725);
buf BUF1 (N11752, N11745);
nor NOR3 (N11753, N11744, N6739, N4221);
not NOT1 (N11754, N11740);
buf BUF1 (N11755, N11752);
and AND4 (N11756, N11753, N11635, N3935, N7829);
or OR2 (N11757, N11743, N2687);
not NOT1 (N11758, N11747);
or OR4 (N11759, N11746, N1874, N1672, N9885);
buf BUF1 (N11760, N11732);
nor NOR2 (N11761, N11754, N7935);
xor XOR2 (N11762, N11751, N1944);
and AND2 (N11763, N11757, N2843);
xor XOR2 (N11764, N11755, N5628);
nor NOR4 (N11765, N11750, N1176, N11651, N5018);
nand NAND2 (N11766, N11761, N6533);
nand NAND4 (N11767, N11763, N10483, N1111, N4057);
not NOT1 (N11768, N11756);
xor XOR2 (N11769, N11758, N3432);
nor NOR2 (N11770, N11748, N10801);
xor XOR2 (N11771, N11770, N9230);
nor NOR4 (N11772, N11765, N8152, N6498, N5480);
and AND4 (N11773, N11759, N7233, N5939, N7159);
xor XOR2 (N11774, N11769, N7379);
buf BUF1 (N11775, N11766);
nor NOR2 (N11776, N11767, N5729);
not NOT1 (N11777, N11762);
buf BUF1 (N11778, N11760);
nor NOR2 (N11779, N11764, N8924);
nand NAND2 (N11780, N11772, N4780);
and AND2 (N11781, N11768, N9945);
nand NAND2 (N11782, N11773, N3419);
buf BUF1 (N11783, N11775);
buf BUF1 (N11784, N11777);
and AND2 (N11785, N11774, N8241);
nor NOR2 (N11786, N11779, N7562);
not NOT1 (N11787, N11776);
and AND3 (N11788, N11771, N9229, N9410);
nor NOR3 (N11789, N11785, N5651, N3243);
and AND3 (N11790, N11783, N305, N2310);
buf BUF1 (N11791, N11781);
nor NOR3 (N11792, N11791, N1581, N3078);
and AND3 (N11793, N11787, N11783, N9208);
nor NOR4 (N11794, N11788, N3266, N2492, N5191);
not NOT1 (N11795, N11793);
buf BUF1 (N11796, N11786);
or OR4 (N11797, N11796, N392, N3782, N8062);
nand NAND4 (N11798, N11780, N7196, N8005, N1351);
xor XOR2 (N11799, N11792, N6243);
and AND4 (N11800, N11797, N3539, N9224, N9535);
nor NOR2 (N11801, N11778, N8062);
nand NAND3 (N11802, N11799, N3681, N2728);
or OR2 (N11803, N11800, N7481);
nand NAND2 (N11804, N11782, N10270);
nand NAND3 (N11805, N11784, N545, N9691);
nand NAND2 (N11806, N11802, N11801);
or OR3 (N11807, N3847, N1093, N3100);
nand NAND4 (N11808, N11807, N4429, N9215, N8315);
buf BUF1 (N11809, N11808);
nand NAND3 (N11810, N11790, N6067, N1597);
not NOT1 (N11811, N11804);
buf BUF1 (N11812, N11806);
not NOT1 (N11813, N11812);
xor XOR2 (N11814, N11789, N2547);
or OR3 (N11815, N11798, N11767, N3682);
nor NOR2 (N11816, N11803, N6160);
xor XOR2 (N11817, N11794, N4428);
xor XOR2 (N11818, N11809, N4444);
xor XOR2 (N11819, N11814, N4271);
xor XOR2 (N11820, N11805, N10527);
buf BUF1 (N11821, N11817);
and AND4 (N11822, N11813, N6154, N9346, N4721);
not NOT1 (N11823, N11821);
nand NAND4 (N11824, N11818, N10553, N10359, N10144);
or OR3 (N11825, N11824, N5995, N8586);
or OR4 (N11826, N11822, N180, N5805, N5774);
nand NAND2 (N11827, N11811, N9808);
and AND3 (N11828, N11795, N6421, N8671);
not NOT1 (N11829, N11827);
buf BUF1 (N11830, N11819);
and AND3 (N11831, N11825, N10646, N1013);
not NOT1 (N11832, N11831);
nand NAND3 (N11833, N11830, N4053, N3294);
and AND4 (N11834, N11810, N6955, N1101, N2449);
nor NOR3 (N11835, N11829, N3681, N8562);
xor XOR2 (N11836, N11834, N4762);
or OR2 (N11837, N11826, N8232);
xor XOR2 (N11838, N11837, N7521);
not NOT1 (N11839, N11832);
nor NOR4 (N11840, N11839, N6668, N2626, N6962);
nand NAND4 (N11841, N11828, N4781, N4259, N11432);
or OR2 (N11842, N11841, N9477);
xor XOR2 (N11843, N11815, N4011);
not NOT1 (N11844, N11840);
nand NAND4 (N11845, N11843, N9011, N10335, N9752);
xor XOR2 (N11846, N11838, N11042);
buf BUF1 (N11847, N11816);
or OR3 (N11848, N11844, N1556, N8940);
and AND2 (N11849, N11835, N3193);
or OR3 (N11850, N11833, N7545, N5347);
nor NOR4 (N11851, N11836, N5716, N4642, N2215);
nand NAND4 (N11852, N11851, N9256, N6708, N8473);
not NOT1 (N11853, N11820);
and AND2 (N11854, N11846, N11238);
xor XOR2 (N11855, N11848, N10271);
xor XOR2 (N11856, N11823, N3360);
and AND2 (N11857, N11854, N3240);
xor XOR2 (N11858, N11856, N11183);
or OR3 (N11859, N11849, N9453, N2564);
nand NAND4 (N11860, N11845, N9447, N511, N8895);
not NOT1 (N11861, N11858);
nand NAND2 (N11862, N11861, N10717);
or OR3 (N11863, N11852, N11779, N9869);
xor XOR2 (N11864, N11857, N3946);
or OR3 (N11865, N11863, N2859, N9362);
nor NOR3 (N11866, N11862, N3062, N9230);
xor XOR2 (N11867, N11855, N7163);
and AND3 (N11868, N11860, N3260, N9485);
or OR2 (N11869, N11847, N2987);
xor XOR2 (N11870, N11868, N7820);
buf BUF1 (N11871, N11859);
and AND3 (N11872, N11864, N10235, N692);
nor NOR2 (N11873, N11871, N6204);
nand NAND4 (N11874, N11853, N9752, N1087, N9323);
nor NOR4 (N11875, N11842, N996, N6241, N9128);
not NOT1 (N11876, N11865);
nor NOR4 (N11877, N11870, N6237, N3662, N7698);
not NOT1 (N11878, N11875);
xor XOR2 (N11879, N11867, N9676);
and AND2 (N11880, N11850, N421);
nor NOR3 (N11881, N11872, N3119, N3190);
not NOT1 (N11882, N11876);
nor NOR2 (N11883, N11878, N160);
or OR3 (N11884, N11883, N5945, N2011);
xor XOR2 (N11885, N11877, N10265);
not NOT1 (N11886, N11866);
xor XOR2 (N11887, N11884, N274);
or OR4 (N11888, N11882, N7998, N8898, N517);
not NOT1 (N11889, N11880);
nand NAND4 (N11890, N11887, N6984, N7832, N11612);
buf BUF1 (N11891, N11881);
buf BUF1 (N11892, N11874);
xor XOR2 (N11893, N11890, N6683);
or OR4 (N11894, N11886, N784, N11458, N8982);
nand NAND4 (N11895, N11888, N646, N7997, N10503);
or OR3 (N11896, N11869, N4913, N5612);
not NOT1 (N11897, N11892);
or OR3 (N11898, N11897, N10876, N169);
or OR2 (N11899, N11873, N6909);
xor XOR2 (N11900, N11896, N3268);
nand NAND2 (N11901, N11893, N3212);
or OR3 (N11902, N11901, N4234, N8057);
nor NOR3 (N11903, N11894, N4690, N9644);
or OR3 (N11904, N11891, N1557, N6057);
buf BUF1 (N11905, N11903);
and AND4 (N11906, N11889, N7804, N3196, N11548);
xor XOR2 (N11907, N11895, N270);
not NOT1 (N11908, N11907);
or OR3 (N11909, N11904, N3651, N9424);
not NOT1 (N11910, N11885);
and AND3 (N11911, N11900, N1346, N9073);
nand NAND3 (N11912, N11908, N9455, N3891);
or OR4 (N11913, N11879, N2753, N7566, N3844);
xor XOR2 (N11914, N11913, N5060);
xor XOR2 (N11915, N11898, N7915);
xor XOR2 (N11916, N11911, N252);
and AND4 (N11917, N11915, N1473, N7993, N3832);
and AND3 (N11918, N11906, N5367, N9154);
nor NOR2 (N11919, N11902, N8248);
and AND4 (N11920, N11909, N8216, N4557, N3508);
nand NAND2 (N11921, N11920, N4897);
and AND4 (N11922, N11910, N4511, N6719, N5130);
nand NAND3 (N11923, N11921, N3299, N8534);
or OR3 (N11924, N11919, N9232, N2541);
buf BUF1 (N11925, N11924);
or OR3 (N11926, N11914, N11875, N8312);
nand NAND2 (N11927, N11899, N2061);
buf BUF1 (N11928, N11922);
or OR2 (N11929, N11927, N10449);
xor XOR2 (N11930, N11928, N8015);
buf BUF1 (N11931, N11923);
nand NAND4 (N11932, N11917, N9361, N8640, N1938);
or OR3 (N11933, N11916, N3883, N11746);
nor NOR4 (N11934, N11925, N2514, N11022, N7006);
and AND3 (N11935, N11933, N11925, N6370);
nor NOR2 (N11936, N11932, N1140);
and AND3 (N11937, N11936, N2337, N11338);
xor XOR2 (N11938, N11931, N9583);
buf BUF1 (N11939, N11929);
buf BUF1 (N11940, N11918);
and AND4 (N11941, N11938, N2802, N8473, N8963);
buf BUF1 (N11942, N11935);
xor XOR2 (N11943, N11912, N3605);
not NOT1 (N11944, N11937);
and AND2 (N11945, N11944, N3268);
or OR2 (N11946, N11943, N3155);
not NOT1 (N11947, N11926);
xor XOR2 (N11948, N11905, N8890);
buf BUF1 (N11949, N11947);
buf BUF1 (N11950, N11942);
nand NAND2 (N11951, N11950, N6969);
or OR4 (N11952, N11934, N3852, N8135, N10816);
nand NAND2 (N11953, N11952, N2720);
nand NAND2 (N11954, N11951, N10764);
or OR4 (N11955, N11946, N4449, N5757, N3513);
xor XOR2 (N11956, N11930, N7673);
and AND2 (N11957, N11953, N1796);
nor NOR3 (N11958, N11954, N9677, N2797);
not NOT1 (N11959, N11957);
nor NOR4 (N11960, N11945, N8936, N2465, N10690);
xor XOR2 (N11961, N11939, N1985);
or OR2 (N11962, N11955, N4262);
not NOT1 (N11963, N11940);
xor XOR2 (N11964, N11960, N9331);
buf BUF1 (N11965, N11959);
buf BUF1 (N11966, N11941);
not NOT1 (N11967, N11962);
nand NAND4 (N11968, N11961, N11094, N1996, N3600);
or OR3 (N11969, N11966, N1705, N11913);
not NOT1 (N11970, N11948);
not NOT1 (N11971, N11968);
and AND3 (N11972, N11949, N9253, N2158);
not NOT1 (N11973, N11971);
buf BUF1 (N11974, N11969);
nor NOR3 (N11975, N11958, N11224, N8149);
and AND4 (N11976, N11975, N8323, N167, N7738);
not NOT1 (N11977, N11967);
or OR2 (N11978, N11964, N10010);
or OR4 (N11979, N11974, N70, N4154, N9434);
buf BUF1 (N11980, N11963);
or OR4 (N11981, N11956, N4134, N2153, N5875);
xor XOR2 (N11982, N11965, N11244);
nor NOR2 (N11983, N11981, N4053);
and AND4 (N11984, N11980, N11099, N5047, N1285);
xor XOR2 (N11985, N11982, N6125);
xor XOR2 (N11986, N11978, N3075);
not NOT1 (N11987, N11970);
buf BUF1 (N11988, N11984);
buf BUF1 (N11989, N11973);
or OR4 (N11990, N11972, N10730, N2909, N7859);
or OR2 (N11991, N11985, N5181);
and AND3 (N11992, N11986, N8649, N3002);
not NOT1 (N11993, N11983);
xor XOR2 (N11994, N11979, N2081);
and AND2 (N11995, N11991, N9281);
not NOT1 (N11996, N11987);
or OR3 (N11997, N11994, N2684, N1867);
xor XOR2 (N11998, N11989, N3961);
or OR4 (N11999, N11993, N597, N11722, N6350);
or OR4 (N12000, N11995, N5141, N4862, N1916);
nor NOR4 (N12001, N11988, N2399, N2585, N3240);
and AND3 (N12002, N12000, N454, N8208);
not NOT1 (N12003, N11996);
buf BUF1 (N12004, N11999);
not NOT1 (N12005, N12001);
nor NOR2 (N12006, N12003, N1242);
buf BUF1 (N12007, N12002);
and AND4 (N12008, N11977, N4303, N9229, N9122);
nor NOR4 (N12009, N12004, N270, N8361, N11721);
not NOT1 (N12010, N12005);
or OR4 (N12011, N12010, N4966, N788, N10282);
xor XOR2 (N12012, N12009, N4948);
buf BUF1 (N12013, N12006);
nand NAND2 (N12014, N12011, N1770);
buf BUF1 (N12015, N11997);
buf BUF1 (N12016, N12015);
xor XOR2 (N12017, N11992, N11612);
and AND4 (N12018, N12013, N3571, N11899, N2748);
not NOT1 (N12019, N12017);
nor NOR4 (N12020, N12018, N11542, N4520, N11517);
xor XOR2 (N12021, N11976, N4054);
not NOT1 (N12022, N11990);
nand NAND3 (N12023, N12021, N10073, N1020);
buf BUF1 (N12024, N11998);
or OR4 (N12025, N12024, N11755, N7069, N7824);
not NOT1 (N12026, N12012);
nor NOR2 (N12027, N12014, N3311);
nand NAND2 (N12028, N12007, N7937);
nor NOR4 (N12029, N12028, N11869, N7249, N3155);
not NOT1 (N12030, N12020);
or OR4 (N12031, N12025, N1384, N9108, N5410);
and AND3 (N12032, N12008, N10758, N7029);
and AND3 (N12033, N12023, N7122, N2034);
xor XOR2 (N12034, N12033, N11590);
nand NAND2 (N12035, N12034, N7327);
or OR2 (N12036, N12026, N2587);
or OR2 (N12037, N12022, N2623);
or OR2 (N12038, N12032, N6803);
and AND3 (N12039, N12029, N4868, N3879);
nand NAND3 (N12040, N12030, N9971, N10272);
nand NAND4 (N12041, N12038, N2514, N3732, N810);
xor XOR2 (N12042, N12027, N2231);
nor NOR3 (N12043, N12042, N500, N8629);
and AND4 (N12044, N12019, N2418, N8550, N6284);
and AND2 (N12045, N12036, N7453);
buf BUF1 (N12046, N12016);
and AND3 (N12047, N12041, N4903, N8844);
xor XOR2 (N12048, N12031, N11386);
nand NAND2 (N12049, N12039, N5733);
nor NOR4 (N12050, N12044, N11378, N11166, N11681);
nand NAND4 (N12051, N12046, N7721, N3991, N3563);
xor XOR2 (N12052, N12049, N10507);
nand NAND4 (N12053, N12045, N976, N5839, N1647);
not NOT1 (N12054, N12043);
or OR4 (N12055, N12047, N4700, N10426, N3065);
not NOT1 (N12056, N12051);
buf BUF1 (N12057, N12052);
not NOT1 (N12058, N12057);
not NOT1 (N12059, N12058);
buf BUF1 (N12060, N12037);
buf BUF1 (N12061, N12054);
buf BUF1 (N12062, N12056);
xor XOR2 (N12063, N12061, N4775);
nand NAND3 (N12064, N12062, N11728, N9594);
nand NAND2 (N12065, N12060, N7009);
and AND4 (N12066, N12035, N8414, N6982, N1087);
buf BUF1 (N12067, N12055);
xor XOR2 (N12068, N12064, N9183);
xor XOR2 (N12069, N12059, N11905);
buf BUF1 (N12070, N12065);
nand NAND2 (N12071, N12066, N5790);
xor XOR2 (N12072, N12050, N8391);
xor XOR2 (N12073, N12063, N2225);
or OR4 (N12074, N12072, N3375, N2647, N9364);
nand NAND4 (N12075, N12074, N6740, N5171, N6193);
nand NAND3 (N12076, N12048, N3176, N8913);
nand NAND4 (N12077, N12070, N10972, N3791, N1761);
xor XOR2 (N12078, N12040, N690);
not NOT1 (N12079, N12076);
nand NAND2 (N12080, N12069, N9012);
and AND3 (N12081, N12075, N6297, N7777);
buf BUF1 (N12082, N12080);
and AND2 (N12083, N12068, N8477);
xor XOR2 (N12084, N12077, N7068);
or OR3 (N12085, N12084, N1717, N4411);
xor XOR2 (N12086, N12053, N5603);
nor NOR3 (N12087, N12082, N1656, N979);
or OR2 (N12088, N12083, N4138);
not NOT1 (N12089, N12079);
or OR2 (N12090, N12088, N10995);
not NOT1 (N12091, N12078);
nand NAND4 (N12092, N12081, N3394, N7403, N10357);
nor NOR4 (N12093, N12087, N9397, N11149, N11225);
or OR4 (N12094, N12071, N4948, N4626, N7061);
and AND2 (N12095, N12092, N5312);
nor NOR4 (N12096, N12085, N11622, N1743, N7847);
and AND2 (N12097, N12095, N1774);
nand NAND4 (N12098, N12094, N520, N8460, N11217);
buf BUF1 (N12099, N12096);
buf BUF1 (N12100, N12098);
xor XOR2 (N12101, N12090, N8246);
not NOT1 (N12102, N12097);
or OR2 (N12103, N12099, N10794);
xor XOR2 (N12104, N12100, N7235);
or OR2 (N12105, N12067, N2909);
and AND2 (N12106, N12102, N7781);
not NOT1 (N12107, N12093);
buf BUF1 (N12108, N12104);
buf BUF1 (N12109, N12106);
nand NAND4 (N12110, N12073, N12028, N5309, N10237);
and AND2 (N12111, N12086, N4098);
not NOT1 (N12112, N12103);
not NOT1 (N12113, N12105);
and AND4 (N12114, N12107, N10292, N11697, N1708);
not NOT1 (N12115, N12108);
not NOT1 (N12116, N12111);
nand NAND4 (N12117, N12109, N5383, N9793, N9648);
xor XOR2 (N12118, N12091, N1393);
and AND3 (N12119, N12116, N3477, N3418);
buf BUF1 (N12120, N12089);
and AND4 (N12121, N12110, N10423, N9143, N3463);
and AND2 (N12122, N12121, N9223);
nor NOR2 (N12123, N12112, N4842);
nor NOR2 (N12124, N12123, N1781);
or OR3 (N12125, N12120, N3922, N1091);
nand NAND4 (N12126, N12115, N4595, N658, N9373);
and AND3 (N12127, N12101, N6719, N1537);
or OR4 (N12128, N12124, N1208, N3204, N841);
buf BUF1 (N12129, N12118);
nand NAND2 (N12130, N12126, N88);
nor NOR3 (N12131, N12114, N8916, N7110);
buf BUF1 (N12132, N12113);
and AND3 (N12133, N12130, N150, N7592);
nand NAND4 (N12134, N12128, N3243, N551, N6566);
buf BUF1 (N12135, N12119);
and AND3 (N12136, N12135, N1331, N7289);
not NOT1 (N12137, N12122);
not NOT1 (N12138, N12133);
or OR4 (N12139, N12134, N6406, N7790, N11523);
xor XOR2 (N12140, N12139, N5355);
nor NOR4 (N12141, N12131, N1304, N2540, N11893);
or OR2 (N12142, N12127, N7685);
or OR2 (N12143, N12125, N3001);
buf BUF1 (N12144, N12132);
nor NOR3 (N12145, N12144, N2901, N8320);
not NOT1 (N12146, N12145);
not NOT1 (N12147, N12140);
and AND3 (N12148, N12147, N1621, N11353);
buf BUF1 (N12149, N12136);
or OR3 (N12150, N12137, N8742, N10400);
buf BUF1 (N12151, N12138);
buf BUF1 (N12152, N12150);
xor XOR2 (N12153, N12141, N3661);
nand NAND4 (N12154, N12151, N4223, N6509, N343);
and AND4 (N12155, N12117, N6487, N5980, N7152);
xor XOR2 (N12156, N12129, N350);
nand NAND3 (N12157, N12155, N9174, N8495);
not NOT1 (N12158, N12153);
xor XOR2 (N12159, N12146, N4019);
or OR4 (N12160, N12152, N8809, N8606, N361);
buf BUF1 (N12161, N12157);
nand NAND4 (N12162, N12142, N6842, N7790, N5161);
not NOT1 (N12163, N12160);
or OR2 (N12164, N12163, N9121);
nand NAND4 (N12165, N12164, N2436, N7150, N11819);
buf BUF1 (N12166, N12148);
nor NOR4 (N12167, N12161, N11771, N10856, N4196);
and AND3 (N12168, N12149, N11620, N1621);
xor XOR2 (N12169, N12165, N10065);
not NOT1 (N12170, N12166);
not NOT1 (N12171, N12162);
nand NAND4 (N12172, N12170, N143, N7425, N11391);
buf BUF1 (N12173, N12159);
or OR3 (N12174, N12143, N1921, N4033);
buf BUF1 (N12175, N12174);
not NOT1 (N12176, N12158);
nor NOR2 (N12177, N12167, N6436);
nor NOR4 (N12178, N12156, N6006, N993, N790);
or OR2 (N12179, N12168, N3531);
nor NOR3 (N12180, N12154, N889, N1308);
not NOT1 (N12181, N12178);
xor XOR2 (N12182, N12177, N8657);
and AND2 (N12183, N12182, N6474);
and AND2 (N12184, N12171, N6845);
buf BUF1 (N12185, N12173);
buf BUF1 (N12186, N12179);
or OR3 (N12187, N12169, N10143, N5463);
not NOT1 (N12188, N12187);
buf BUF1 (N12189, N12185);
and AND2 (N12190, N12186, N9581);
and AND3 (N12191, N12172, N11171, N6543);
buf BUF1 (N12192, N12180);
xor XOR2 (N12193, N12183, N764);
nand NAND2 (N12194, N12191, N1426);
or OR2 (N12195, N12181, N5298);
nor NOR2 (N12196, N12192, N4180);
or OR4 (N12197, N12188, N6702, N8250, N5466);
nor NOR2 (N12198, N12176, N2843);
nor NOR2 (N12199, N12194, N11660);
nor NOR4 (N12200, N12175, N5502, N9099, N8537);
buf BUF1 (N12201, N12197);
buf BUF1 (N12202, N12198);
nand NAND3 (N12203, N12202, N8014, N6064);
not NOT1 (N12204, N12201);
xor XOR2 (N12205, N12184, N6025);
or OR3 (N12206, N12205, N914, N5566);
and AND3 (N12207, N12195, N7279, N7420);
nor NOR4 (N12208, N12199, N995, N11507, N9816);
buf BUF1 (N12209, N12190);
nor NOR2 (N12210, N12206, N2269);
xor XOR2 (N12211, N12210, N10239);
and AND2 (N12212, N12204, N7718);
not NOT1 (N12213, N12207);
not NOT1 (N12214, N12203);
nand NAND2 (N12215, N12214, N11375);
not NOT1 (N12216, N12215);
or OR4 (N12217, N12212, N8617, N5429, N7839);
or OR4 (N12218, N12211, N9009, N2054, N2511);
nor NOR3 (N12219, N12189, N9828, N8051);
not NOT1 (N12220, N12218);
buf BUF1 (N12221, N12209);
not NOT1 (N12222, N12200);
xor XOR2 (N12223, N12196, N10682);
buf BUF1 (N12224, N12216);
buf BUF1 (N12225, N12223);
buf BUF1 (N12226, N12222);
buf BUF1 (N12227, N12226);
nand NAND3 (N12228, N12213, N2381, N1824);
xor XOR2 (N12229, N12225, N3778);
nor NOR4 (N12230, N12227, N9892, N1986, N7371);
xor XOR2 (N12231, N12221, N9064);
or OR3 (N12232, N12231, N11303, N6914);
buf BUF1 (N12233, N12224);
or OR2 (N12234, N12208, N11104);
buf BUF1 (N12235, N12193);
nor NOR4 (N12236, N12228, N8354, N6185, N1234);
nor NOR4 (N12237, N12236, N5566, N4572, N3310);
and AND4 (N12238, N12235, N1252, N9779, N1415);
nand NAND3 (N12239, N12234, N4145, N12093);
buf BUF1 (N12240, N12230);
or OR3 (N12241, N12237, N11608, N3007);
and AND3 (N12242, N12239, N11932, N5323);
buf BUF1 (N12243, N12242);
nor NOR3 (N12244, N12217, N10655, N7425);
nor NOR2 (N12245, N12233, N10580);
nand NAND3 (N12246, N12232, N9815, N4293);
and AND3 (N12247, N12220, N330, N5426);
or OR4 (N12248, N12245, N10070, N1568, N2525);
xor XOR2 (N12249, N12238, N9378);
not NOT1 (N12250, N12243);
buf BUF1 (N12251, N12246);
buf BUF1 (N12252, N12229);
not NOT1 (N12253, N12248);
and AND3 (N12254, N12241, N3979, N5682);
and AND2 (N12255, N12244, N6545);
or OR4 (N12256, N12219, N5568, N1816, N7260);
xor XOR2 (N12257, N12250, N2175);
and AND4 (N12258, N12252, N7322, N2506, N3595);
and AND3 (N12259, N12254, N8212, N11100);
buf BUF1 (N12260, N12259);
buf BUF1 (N12261, N12257);
not NOT1 (N12262, N12253);
nand NAND3 (N12263, N12256, N12193, N574);
buf BUF1 (N12264, N12251);
nand NAND4 (N12265, N12249, N10086, N1827, N4197);
nor NOR3 (N12266, N12264, N578, N2768);
not NOT1 (N12267, N12255);
nor NOR4 (N12268, N12265, N4553, N1797, N561);
not NOT1 (N12269, N12268);
nand NAND2 (N12270, N12260, N7828);
not NOT1 (N12271, N12258);
nand NAND3 (N12272, N12270, N7878, N1494);
buf BUF1 (N12273, N12263);
or OR3 (N12274, N12269, N255, N969);
xor XOR2 (N12275, N12261, N9493);
or OR2 (N12276, N12267, N11257);
nand NAND2 (N12277, N12262, N12210);
not NOT1 (N12278, N12240);
and AND3 (N12279, N12278, N7484, N10098);
buf BUF1 (N12280, N12275);
nand NAND2 (N12281, N12279, N1972);
nand NAND4 (N12282, N12280, N10234, N4004, N10073);
nand NAND3 (N12283, N12247, N4376, N3593);
or OR3 (N12284, N12283, N3277, N4127);
nand NAND4 (N12285, N12266, N11440, N10601, N7539);
buf BUF1 (N12286, N12282);
and AND3 (N12287, N12277, N5152, N3604);
nor NOR2 (N12288, N12287, N1220);
nor NOR4 (N12289, N12274, N4767, N3737, N4035);
xor XOR2 (N12290, N12276, N10487);
and AND2 (N12291, N12271, N8487);
buf BUF1 (N12292, N12286);
and AND3 (N12293, N12289, N8522, N7038);
nand NAND4 (N12294, N12273, N9867, N10828, N9316);
nor NOR4 (N12295, N12291, N1777, N9629, N8148);
xor XOR2 (N12296, N12293, N6580);
nor NOR2 (N12297, N12285, N9598);
buf BUF1 (N12298, N12296);
buf BUF1 (N12299, N12295);
or OR2 (N12300, N12290, N1353);
nand NAND4 (N12301, N12300, N3990, N4898, N776);
xor XOR2 (N12302, N12294, N8634);
buf BUF1 (N12303, N12297);
buf BUF1 (N12304, N12298);
nand NAND4 (N12305, N12301, N400, N2455, N6517);
not NOT1 (N12306, N12288);
nor NOR2 (N12307, N12292, N5852);
or OR4 (N12308, N12281, N8786, N12100, N7101);
buf BUF1 (N12309, N12303);
not NOT1 (N12310, N12305);
buf BUF1 (N12311, N12284);
or OR4 (N12312, N12309, N10708, N6111, N11771);
or OR2 (N12313, N12311, N8231);
buf BUF1 (N12314, N12306);
or OR4 (N12315, N12302, N11742, N6024, N11322);
nand NAND2 (N12316, N12310, N9161);
nor NOR4 (N12317, N12316, N781, N5775, N9187);
not NOT1 (N12318, N12307);
nand NAND2 (N12319, N12272, N2716);
buf BUF1 (N12320, N12315);
not NOT1 (N12321, N12299);
nor NOR4 (N12322, N12314, N656, N6463, N6763);
nand NAND4 (N12323, N12320, N9529, N4250, N4334);
nand NAND2 (N12324, N12313, N8448);
and AND4 (N12325, N12308, N8141, N10079, N7136);
and AND2 (N12326, N12318, N8401);
nor NOR2 (N12327, N12326, N3582);
or OR4 (N12328, N12323, N8773, N3840, N8166);
not NOT1 (N12329, N12319);
buf BUF1 (N12330, N12304);
buf BUF1 (N12331, N12325);
and AND2 (N12332, N12321, N7164);
or OR3 (N12333, N12329, N11871, N5624);
and AND2 (N12334, N12322, N7431);
not NOT1 (N12335, N12328);
and AND3 (N12336, N12327, N7543, N8091);
nand NAND4 (N12337, N12331, N11099, N6641, N2366);
xor XOR2 (N12338, N12337, N8552);
or OR2 (N12339, N12332, N8067);
nand NAND3 (N12340, N12335, N5082, N11019);
and AND4 (N12341, N12312, N2022, N8452, N10787);
not NOT1 (N12342, N12333);
and AND3 (N12343, N12336, N10983, N4100);
buf BUF1 (N12344, N12341);
xor XOR2 (N12345, N12324, N4721);
xor XOR2 (N12346, N12340, N7397);
nand NAND2 (N12347, N12344, N6454);
nand NAND4 (N12348, N12334, N5610, N1013, N1680);
and AND3 (N12349, N12343, N703, N4265);
buf BUF1 (N12350, N12317);
or OR4 (N12351, N12330, N12333, N3506, N3563);
and AND2 (N12352, N12348, N4353);
and AND2 (N12353, N12339, N5793);
buf BUF1 (N12354, N12347);
xor XOR2 (N12355, N12353, N5513);
and AND3 (N12356, N12338, N6969, N2863);
or OR3 (N12357, N12352, N1061, N7422);
or OR3 (N12358, N12354, N5444, N3316);
nor NOR3 (N12359, N12350, N11357, N8373);
nor NOR3 (N12360, N12357, N6377, N8450);
nor NOR4 (N12361, N12349, N11927, N6045, N2696);
buf BUF1 (N12362, N12342);
buf BUF1 (N12363, N12359);
nand NAND3 (N12364, N12345, N11083, N1064);
xor XOR2 (N12365, N12351, N6277);
not NOT1 (N12366, N12356);
buf BUF1 (N12367, N12366);
not NOT1 (N12368, N12363);
nand NAND3 (N12369, N12360, N2315, N9032);
nand NAND3 (N12370, N12362, N11238, N2299);
buf BUF1 (N12371, N12364);
nor NOR2 (N12372, N12346, N3472);
not NOT1 (N12373, N12365);
buf BUF1 (N12374, N12369);
nand NAND3 (N12375, N12373, N3651, N7255);
nor NOR4 (N12376, N12375, N7773, N1737, N285);
not NOT1 (N12377, N12358);
buf BUF1 (N12378, N12370);
xor XOR2 (N12379, N12372, N2372);
nand NAND2 (N12380, N12367, N7033);
not NOT1 (N12381, N12376);
nand NAND4 (N12382, N12379, N5829, N1807, N12123);
and AND4 (N12383, N12374, N3607, N4622, N7366);
nand NAND4 (N12384, N12382, N2525, N8387, N9308);
buf BUF1 (N12385, N12378);
and AND2 (N12386, N12384, N8671);
and AND3 (N12387, N12385, N8543, N8122);
not NOT1 (N12388, N12380);
buf BUF1 (N12389, N12388);
xor XOR2 (N12390, N12386, N3398);
not NOT1 (N12391, N12387);
and AND2 (N12392, N12361, N5448);
or OR2 (N12393, N12377, N3545);
nor NOR2 (N12394, N12390, N3911);
nand NAND2 (N12395, N12355, N284);
or OR2 (N12396, N12383, N1168);
nand NAND2 (N12397, N12381, N4477);
xor XOR2 (N12398, N12392, N10986);
and AND4 (N12399, N12397, N6020, N2528, N4718);
or OR4 (N12400, N12394, N12279, N10898, N10199);
and AND4 (N12401, N12389, N11517, N8031, N2990);
xor XOR2 (N12402, N12398, N11428);
nor NOR3 (N12403, N12396, N10501, N8813);
or OR4 (N12404, N12395, N5823, N4721, N10889);
xor XOR2 (N12405, N12393, N9711);
or OR2 (N12406, N12368, N2576);
nand NAND2 (N12407, N12400, N8707);
buf BUF1 (N12408, N12404);
buf BUF1 (N12409, N12403);
nand NAND2 (N12410, N12401, N9976);
nor NOR2 (N12411, N12371, N10274);
xor XOR2 (N12412, N12407, N9343);
nor NOR3 (N12413, N12408, N4315, N9474);
not NOT1 (N12414, N12410);
xor XOR2 (N12415, N12411, N10360);
xor XOR2 (N12416, N12412, N5901);
nand NAND2 (N12417, N12406, N10086);
buf BUF1 (N12418, N12414);
nor NOR3 (N12419, N12417, N2845, N2808);
or OR4 (N12420, N12391, N9171, N1848, N12216);
or OR3 (N12421, N12399, N10098, N4673);
or OR4 (N12422, N12420, N10324, N5065, N3298);
and AND4 (N12423, N12421, N4434, N4726, N544);
and AND3 (N12424, N12416, N3008, N175);
nand NAND3 (N12425, N12409, N6365, N8740);
or OR2 (N12426, N12413, N4860);
not NOT1 (N12427, N12402);
nor NOR2 (N12428, N12427, N2803);
and AND4 (N12429, N12426, N8335, N4653, N2349);
not NOT1 (N12430, N12422);
or OR2 (N12431, N12418, N8180);
and AND3 (N12432, N12425, N6780, N284);
or OR3 (N12433, N12428, N8886, N277);
nor NOR3 (N12434, N12415, N8976, N7958);
xor XOR2 (N12435, N12424, N3598);
nor NOR2 (N12436, N12433, N11912);
or OR4 (N12437, N12434, N9008, N8910, N3083);
nor NOR2 (N12438, N12405, N11661);
nor NOR2 (N12439, N12437, N236);
nand NAND4 (N12440, N12436, N7054, N10568, N8342);
and AND3 (N12441, N12440, N8338, N9993);
and AND4 (N12442, N12430, N4590, N8207, N8156);
nor NOR4 (N12443, N12431, N7539, N5108, N9497);
and AND3 (N12444, N12438, N10588, N1019);
or OR3 (N12445, N12419, N2521, N7966);
buf BUF1 (N12446, N12435);
nand NAND4 (N12447, N12423, N10845, N3075, N4000);
not NOT1 (N12448, N12443);
and AND4 (N12449, N12447, N1161, N7093, N946);
not NOT1 (N12450, N12442);
and AND3 (N12451, N12449, N8139, N2958);
not NOT1 (N12452, N12441);
not NOT1 (N12453, N12432);
nand NAND2 (N12454, N12439, N1679);
nor NOR4 (N12455, N12448, N11143, N9118, N3251);
nand NAND4 (N12456, N12454, N9597, N4041, N11660);
or OR3 (N12457, N12446, N10218, N5367);
not NOT1 (N12458, N12457);
nor NOR3 (N12459, N12451, N11582, N1992);
buf BUF1 (N12460, N12456);
nand NAND2 (N12461, N12429, N11192);
xor XOR2 (N12462, N12461, N9208);
buf BUF1 (N12463, N12458);
and AND4 (N12464, N12462, N10038, N361, N976);
buf BUF1 (N12465, N12460);
buf BUF1 (N12466, N12445);
and AND2 (N12467, N12463, N10841);
nor NOR2 (N12468, N12465, N11855);
nor NOR4 (N12469, N12459, N8406, N6452, N4457);
nor NOR3 (N12470, N12444, N10842, N2095);
buf BUF1 (N12471, N12468);
not NOT1 (N12472, N12471);
not NOT1 (N12473, N12452);
not NOT1 (N12474, N12467);
buf BUF1 (N12475, N12474);
and AND3 (N12476, N12466, N10355, N2618);
xor XOR2 (N12477, N12469, N2007);
nand NAND3 (N12478, N12470, N8604, N2087);
or OR4 (N12479, N12475, N5456, N784, N3031);
buf BUF1 (N12480, N12476);
xor XOR2 (N12481, N12478, N12057);
not NOT1 (N12482, N12453);
and AND2 (N12483, N12455, N9056);
or OR3 (N12484, N12472, N8451, N3522);
xor XOR2 (N12485, N12450, N7235);
xor XOR2 (N12486, N12480, N10312);
nand NAND4 (N12487, N12484, N699, N6638, N7732);
xor XOR2 (N12488, N12483, N1212);
not NOT1 (N12489, N12488);
and AND2 (N12490, N12481, N4729);
and AND4 (N12491, N12477, N2300, N2161, N8834);
not NOT1 (N12492, N12485);
xor XOR2 (N12493, N12490, N4383);
or OR4 (N12494, N12489, N11215, N5796, N5863);
and AND3 (N12495, N12473, N7883, N4676);
not NOT1 (N12496, N12492);
or OR2 (N12497, N12482, N12484);
buf BUF1 (N12498, N12487);
nor NOR4 (N12499, N12498, N6141, N11267, N665);
xor XOR2 (N12500, N12494, N3505);
buf BUF1 (N12501, N12479);
buf BUF1 (N12502, N12499);
xor XOR2 (N12503, N12493, N6419);
or OR2 (N12504, N12497, N1072);
buf BUF1 (N12505, N12486);
xor XOR2 (N12506, N12496, N7142);
nor NOR4 (N12507, N12501, N10515, N1449, N5773);
nand NAND2 (N12508, N12505, N8668);
or OR3 (N12509, N12508, N7143, N11403);
and AND3 (N12510, N12506, N5077, N11937);
nor NOR4 (N12511, N12491, N1513, N10130, N5459);
xor XOR2 (N12512, N12500, N10836);
xor XOR2 (N12513, N12512, N1889);
nor NOR3 (N12514, N12511, N11835, N9950);
xor XOR2 (N12515, N12510, N10373);
nor NOR3 (N12516, N12502, N6112, N3238);
and AND3 (N12517, N12503, N11374, N7143);
or OR4 (N12518, N12504, N3446, N9389, N3925);
or OR4 (N12519, N12495, N6275, N3368, N8840);
nor NOR3 (N12520, N12515, N11450, N3499);
nor NOR3 (N12521, N12514, N10604, N10427);
nand NAND2 (N12522, N12507, N7261);
nand NAND4 (N12523, N12521, N8176, N9699, N5952);
not NOT1 (N12524, N12464);
buf BUF1 (N12525, N12517);
xor XOR2 (N12526, N12518, N8742);
or OR2 (N12527, N12520, N10867);
nor NOR4 (N12528, N12525, N10035, N5071, N826);
not NOT1 (N12529, N12528);
or OR4 (N12530, N12522, N11296, N3978, N6148);
not NOT1 (N12531, N12530);
buf BUF1 (N12532, N12529);
nand NAND2 (N12533, N12524, N3508);
buf BUF1 (N12534, N12531);
not NOT1 (N12535, N12509);
and AND3 (N12536, N12534, N526, N12106);
and AND2 (N12537, N12527, N4966);
not NOT1 (N12538, N12536);
not NOT1 (N12539, N12513);
xor XOR2 (N12540, N12523, N5517);
nor NOR2 (N12541, N12516, N7751);
not NOT1 (N12542, N12540);
xor XOR2 (N12543, N12538, N9187);
xor XOR2 (N12544, N12541, N4485);
not NOT1 (N12545, N12526);
buf BUF1 (N12546, N12519);
or OR2 (N12547, N12543, N451);
not NOT1 (N12548, N12546);
buf BUF1 (N12549, N12545);
buf BUF1 (N12550, N12547);
xor XOR2 (N12551, N12535, N2256);
or OR3 (N12552, N12537, N6422, N7314);
nor NOR4 (N12553, N12552, N6854, N4390, N10109);
buf BUF1 (N12554, N12550);
nand NAND3 (N12555, N12551, N1145, N2520);
xor XOR2 (N12556, N12548, N7727);
or OR2 (N12557, N12539, N8904);
xor XOR2 (N12558, N12556, N2580);
not NOT1 (N12559, N12549);
not NOT1 (N12560, N12532);
and AND3 (N12561, N12560, N9316, N6601);
xor XOR2 (N12562, N12558, N10084);
or OR2 (N12563, N12557, N3811);
nor NOR4 (N12564, N12544, N8859, N5819, N1573);
and AND4 (N12565, N12563, N3088, N11118, N5062);
and AND3 (N12566, N12542, N9643, N2437);
and AND4 (N12567, N12553, N11058, N8383, N7836);
not NOT1 (N12568, N12562);
nand NAND2 (N12569, N12564, N9125);
nand NAND4 (N12570, N12561, N5325, N6743, N11344);
and AND3 (N12571, N12570, N9561, N9499);
nor NOR3 (N12572, N12568, N11361, N9709);
buf BUF1 (N12573, N12567);
not NOT1 (N12574, N12571);
or OR3 (N12575, N12533, N6712, N10699);
and AND4 (N12576, N12565, N10053, N6605, N11312);
nand NAND4 (N12577, N12574, N10955, N4697, N7005);
xor XOR2 (N12578, N12577, N12128);
nor NOR3 (N12579, N12569, N5669, N3743);
nand NAND2 (N12580, N12576, N2237);
not NOT1 (N12581, N12578);
and AND3 (N12582, N12555, N6587, N2442);
xor XOR2 (N12583, N12554, N3611);
nor NOR2 (N12584, N12581, N5990);
not NOT1 (N12585, N12579);
buf BUF1 (N12586, N12584);
or OR3 (N12587, N12580, N10816, N11123);
not NOT1 (N12588, N12559);
buf BUF1 (N12589, N12572);
buf BUF1 (N12590, N12588);
or OR3 (N12591, N12585, N10979, N972);
xor XOR2 (N12592, N12591, N8766);
buf BUF1 (N12593, N12592);
buf BUF1 (N12594, N12590);
or OR4 (N12595, N12589, N3954, N6818, N1605);
xor XOR2 (N12596, N12595, N7579);
buf BUF1 (N12597, N12586);
nand NAND3 (N12598, N12594, N5519, N3750);
xor XOR2 (N12599, N12575, N10595);
and AND2 (N12600, N12582, N6672);
nand NAND3 (N12601, N12597, N7431, N3044);
nor NOR4 (N12602, N12601, N10168, N9774, N10124);
nor NOR3 (N12603, N12587, N9188, N5190);
not NOT1 (N12604, N12599);
and AND3 (N12605, N12566, N7803, N464);
and AND2 (N12606, N12583, N9557);
or OR4 (N12607, N12598, N7929, N7250, N12199);
buf BUF1 (N12608, N12600);
xor XOR2 (N12609, N12593, N625);
and AND2 (N12610, N12606, N5874);
and AND3 (N12611, N12608, N8495, N7076);
buf BUF1 (N12612, N12573);
or OR2 (N12613, N12596, N7427);
buf BUF1 (N12614, N12609);
or OR3 (N12615, N12607, N9512, N9871);
xor XOR2 (N12616, N12610, N6854);
xor XOR2 (N12617, N12613, N1625);
or OR2 (N12618, N12604, N1732);
buf BUF1 (N12619, N12617);
buf BUF1 (N12620, N12614);
nand NAND2 (N12621, N12602, N11380);
or OR2 (N12622, N12619, N4434);
nand NAND4 (N12623, N12618, N12285, N6302, N3521);
buf BUF1 (N12624, N12615);
nor NOR2 (N12625, N12624, N12407);
nand NAND2 (N12626, N12625, N10244);
nor NOR3 (N12627, N12612, N10774, N11027);
xor XOR2 (N12628, N12603, N6822);
or OR4 (N12629, N12621, N11720, N2010, N2044);
not NOT1 (N12630, N12627);
buf BUF1 (N12631, N12629);
xor XOR2 (N12632, N12620, N1956);
nor NOR2 (N12633, N12611, N9592);
nand NAND4 (N12634, N12622, N140, N3183, N10024);
nand NAND3 (N12635, N12631, N940, N10820);
not NOT1 (N12636, N12605);
or OR2 (N12637, N12623, N3354);
and AND4 (N12638, N12634, N744, N4038, N9248);
xor XOR2 (N12639, N12635, N5405);
not NOT1 (N12640, N12636);
buf BUF1 (N12641, N12632);
xor XOR2 (N12642, N12639, N5508);
xor XOR2 (N12643, N12640, N9243);
or OR3 (N12644, N12626, N906, N9531);
buf BUF1 (N12645, N12616);
nand NAND2 (N12646, N12645, N1637);
xor XOR2 (N12647, N12638, N8244);
not NOT1 (N12648, N12646);
or OR2 (N12649, N12633, N414);
not NOT1 (N12650, N12642);
nand NAND2 (N12651, N12648, N7388);
nand NAND4 (N12652, N12649, N12538, N8199, N4918);
xor XOR2 (N12653, N12652, N10556);
nand NAND4 (N12654, N12651, N5752, N6963, N11803);
or OR3 (N12655, N12630, N2149, N10821);
or OR3 (N12656, N12628, N6780, N5896);
nor NOR2 (N12657, N12656, N11837);
buf BUF1 (N12658, N12637);
buf BUF1 (N12659, N12654);
not NOT1 (N12660, N12650);
or OR2 (N12661, N12660, N7474);
buf BUF1 (N12662, N12658);
not NOT1 (N12663, N12644);
or OR2 (N12664, N12659, N602);
xor XOR2 (N12665, N12662, N829);
buf BUF1 (N12666, N12647);
not NOT1 (N12667, N12663);
nor NOR2 (N12668, N12664, N10182);
and AND4 (N12669, N12655, N8446, N6444, N9980);
buf BUF1 (N12670, N12657);
nand NAND2 (N12671, N12665, N8885);
not NOT1 (N12672, N12666);
nand NAND2 (N12673, N12668, N7717);
xor XOR2 (N12674, N12661, N11429);
and AND4 (N12675, N12672, N10022, N49, N10718);
xor XOR2 (N12676, N12675, N1794);
nor NOR4 (N12677, N12669, N5541, N1370, N6922);
and AND3 (N12678, N12643, N5200, N10624);
xor XOR2 (N12679, N12653, N2035);
and AND2 (N12680, N12641, N1839);
xor XOR2 (N12681, N12680, N7960);
nor NOR4 (N12682, N12676, N5926, N3828, N1852);
nor NOR3 (N12683, N12673, N12398, N10758);
xor XOR2 (N12684, N12674, N6710);
nand NAND4 (N12685, N12683, N6523, N9579, N3313);
not NOT1 (N12686, N12671);
buf BUF1 (N12687, N12681);
and AND4 (N12688, N12687, N2352, N10683, N9696);
not NOT1 (N12689, N12685);
nor NOR4 (N12690, N12677, N2502, N10640, N6732);
buf BUF1 (N12691, N12688);
nor NOR3 (N12692, N12684, N2304, N5788);
xor XOR2 (N12693, N12670, N5499);
and AND2 (N12694, N12689, N12391);
not NOT1 (N12695, N12682);
buf BUF1 (N12696, N12686);
nor NOR3 (N12697, N12678, N5094, N9329);
nand NAND2 (N12698, N12693, N5656);
buf BUF1 (N12699, N12679);
not NOT1 (N12700, N12690);
nor NOR4 (N12701, N12700, N10999, N11395, N1643);
nor NOR3 (N12702, N12667, N11102, N10848);
buf BUF1 (N12703, N12695);
not NOT1 (N12704, N12698);
nor NOR3 (N12705, N12701, N7951, N8514);
buf BUF1 (N12706, N12691);
xor XOR2 (N12707, N12705, N11459);
buf BUF1 (N12708, N12699);
nand NAND4 (N12709, N12694, N981, N8483, N7238);
and AND3 (N12710, N12708, N8800, N2668);
buf BUF1 (N12711, N12697);
or OR4 (N12712, N12711, N11745, N8539, N2600);
nor NOR2 (N12713, N12710, N3376);
xor XOR2 (N12714, N12702, N8287);
nor NOR3 (N12715, N12696, N3722, N12462);
and AND2 (N12716, N12713, N8957);
and AND4 (N12717, N12703, N739, N2424, N8143);
buf BUF1 (N12718, N12709);
nor NOR3 (N12719, N12712, N9948, N5209);
nor NOR4 (N12720, N12692, N4235, N12158, N3571);
not NOT1 (N12721, N12714);
not NOT1 (N12722, N12706);
xor XOR2 (N12723, N12721, N12027);
xor XOR2 (N12724, N12723, N6070);
not NOT1 (N12725, N12722);
xor XOR2 (N12726, N12718, N1333);
buf BUF1 (N12727, N12715);
nor NOR3 (N12728, N12707, N12442, N2040);
buf BUF1 (N12729, N12719);
and AND4 (N12730, N12728, N9851, N10386, N550);
not NOT1 (N12731, N12730);
nor NOR3 (N12732, N12724, N5062, N4617);
xor XOR2 (N12733, N12717, N8197);
and AND2 (N12734, N12720, N11134);
nand NAND3 (N12735, N12726, N235, N3674);
xor XOR2 (N12736, N12727, N2114);
and AND2 (N12737, N12729, N2959);
not NOT1 (N12738, N12731);
xor XOR2 (N12739, N12732, N5631);
buf BUF1 (N12740, N12739);
xor XOR2 (N12741, N12725, N8122);
nand NAND4 (N12742, N12733, N9244, N3991, N7571);
or OR2 (N12743, N12735, N3567);
not NOT1 (N12744, N12742);
or OR2 (N12745, N12743, N7033);
and AND2 (N12746, N12704, N8571);
nor NOR3 (N12747, N12736, N462, N6796);
nor NOR2 (N12748, N12741, N7351);
nand NAND2 (N12749, N12716, N6551);
nor NOR3 (N12750, N12748, N7883, N8869);
xor XOR2 (N12751, N12750, N4628);
xor XOR2 (N12752, N12749, N4907);
buf BUF1 (N12753, N12740);
buf BUF1 (N12754, N12734);
and AND2 (N12755, N12747, N1448);
not NOT1 (N12756, N12737);
and AND3 (N12757, N12753, N1530, N12564);
xor XOR2 (N12758, N12738, N2773);
nand NAND4 (N12759, N12751, N1654, N6009, N5013);
nor NOR4 (N12760, N12759, N2389, N436, N6132);
not NOT1 (N12761, N12746);
and AND3 (N12762, N12755, N8622, N4018);
or OR3 (N12763, N12756, N4845, N8362);
buf BUF1 (N12764, N12762);
xor XOR2 (N12765, N12744, N3562);
nor NOR2 (N12766, N12760, N1191);
nand NAND3 (N12767, N12764, N7788, N5255);
not NOT1 (N12768, N12761);
or OR4 (N12769, N12768, N8485, N54, N1594);
and AND2 (N12770, N12767, N2757);
not NOT1 (N12771, N12765);
or OR4 (N12772, N12758, N8412, N5263, N8355);
xor XOR2 (N12773, N12769, N4079);
nor NOR2 (N12774, N12754, N11973);
and AND2 (N12775, N12770, N1004);
nor NOR3 (N12776, N12771, N4665, N4765);
or OR3 (N12777, N12773, N2455, N9121);
and AND3 (N12778, N12752, N2792, N212);
buf BUF1 (N12779, N12763);
buf BUF1 (N12780, N12772);
not NOT1 (N12781, N12777);
nor NOR3 (N12782, N12781, N2134, N79);
xor XOR2 (N12783, N12780, N12567);
xor XOR2 (N12784, N12778, N11433);
buf BUF1 (N12785, N12766);
nor NOR2 (N12786, N12774, N8651);
not NOT1 (N12787, N12775);
not NOT1 (N12788, N12783);
buf BUF1 (N12789, N12785);
nand NAND4 (N12790, N12786, N9308, N2863, N1500);
xor XOR2 (N12791, N12787, N4456);
nor NOR4 (N12792, N12791, N4842, N12150, N2480);
and AND4 (N12793, N12757, N11828, N7829, N6999);
or OR3 (N12794, N12745, N3855, N6388);
nand NAND2 (N12795, N12789, N3970);
nand NAND4 (N12796, N12793, N7753, N5373, N1443);
and AND2 (N12797, N12795, N909);
buf BUF1 (N12798, N12776);
buf BUF1 (N12799, N12788);
buf BUF1 (N12800, N12779);
and AND2 (N12801, N12799, N3279);
not NOT1 (N12802, N12794);
and AND4 (N12803, N12801, N11572, N11257, N636);
or OR4 (N12804, N12797, N12749, N263, N12364);
nand NAND3 (N12805, N12792, N8637, N1916);
or OR3 (N12806, N12782, N6650, N5620);
not NOT1 (N12807, N12796);
nand NAND4 (N12808, N12800, N5244, N1052, N405);
nand NAND3 (N12809, N12798, N10381, N1673);
nand NAND2 (N12810, N12784, N8512);
or OR3 (N12811, N12806, N8729, N10752);
or OR3 (N12812, N12807, N4001, N10112);
not NOT1 (N12813, N12812);
buf BUF1 (N12814, N12809);
buf BUF1 (N12815, N12805);
buf BUF1 (N12816, N12813);
nor NOR4 (N12817, N12815, N682, N11145, N9153);
and AND2 (N12818, N12817, N8604);
nand NAND4 (N12819, N12802, N11186, N5105, N11547);
not NOT1 (N12820, N12816);
or OR4 (N12821, N12808, N235, N10983, N2748);
nor NOR4 (N12822, N12811, N5230, N463, N2466);
not NOT1 (N12823, N12804);
nand NAND4 (N12824, N12820, N9636, N6473, N11174);
xor XOR2 (N12825, N12810, N2566);
nand NAND2 (N12826, N12825, N5595);
or OR4 (N12827, N12814, N3833, N10064, N4413);
nand NAND2 (N12828, N12826, N5864);
and AND3 (N12829, N12828, N8979, N8576);
and AND2 (N12830, N12829, N8753);
xor XOR2 (N12831, N12821, N9667);
not NOT1 (N12832, N12819);
buf BUF1 (N12833, N12831);
buf BUF1 (N12834, N12827);
or OR2 (N12835, N12830, N2353);
nor NOR3 (N12836, N12790, N10700, N4199);
not NOT1 (N12837, N12822);
buf BUF1 (N12838, N12803);
buf BUF1 (N12839, N12837);
nor NOR3 (N12840, N12833, N7530, N8222);
nand NAND4 (N12841, N12823, N3247, N1794, N4086);
buf BUF1 (N12842, N12841);
not NOT1 (N12843, N12834);
nand NAND3 (N12844, N12839, N4904, N11115);
and AND4 (N12845, N12836, N10559, N8776, N11089);
or OR3 (N12846, N12832, N7365, N11971);
or OR3 (N12847, N12844, N7730, N1479);
xor XOR2 (N12848, N12845, N189);
or OR2 (N12849, N12835, N10309);
and AND3 (N12850, N12838, N5553, N7294);
buf BUF1 (N12851, N12843);
or OR2 (N12852, N12848, N6529);
nor NOR4 (N12853, N12818, N5789, N10273, N1611);
buf BUF1 (N12854, N12851);
not NOT1 (N12855, N12853);
or OR3 (N12856, N12854, N8207, N7006);
nor NOR4 (N12857, N12849, N12273, N5192, N2783);
not NOT1 (N12858, N12842);
not NOT1 (N12859, N12858);
not NOT1 (N12860, N12847);
xor XOR2 (N12861, N12857, N10032);
not NOT1 (N12862, N12846);
nor NOR4 (N12863, N12862, N6565, N1168, N12682);
or OR2 (N12864, N12856, N3431);
nor NOR3 (N12865, N12824, N10666, N2123);
nor NOR4 (N12866, N12852, N8405, N6285, N2210);
buf BUF1 (N12867, N12864);
or OR2 (N12868, N12867, N4361);
xor XOR2 (N12869, N12850, N5711);
nor NOR3 (N12870, N12865, N11624, N1637);
xor XOR2 (N12871, N12870, N1167);
nor NOR3 (N12872, N12871, N1259, N9746);
xor XOR2 (N12873, N12840, N5282);
buf BUF1 (N12874, N12872);
nor NOR4 (N12875, N12861, N8832, N9362, N4073);
and AND2 (N12876, N12860, N217);
or OR2 (N12877, N12868, N3160);
buf BUF1 (N12878, N12855);
nand NAND3 (N12879, N12874, N8921, N11177);
and AND3 (N12880, N12873, N1319, N3943);
not NOT1 (N12881, N12876);
xor XOR2 (N12882, N12859, N2794);
or OR4 (N12883, N12880, N2268, N58, N5368);
not NOT1 (N12884, N12882);
nor NOR2 (N12885, N12866, N7788);
nor NOR2 (N12886, N12875, N9065);
nor NOR2 (N12887, N12883, N4293);
not NOT1 (N12888, N12877);
nand NAND3 (N12889, N12863, N10403, N12220);
buf BUF1 (N12890, N12887);
or OR3 (N12891, N12885, N2573, N5117);
buf BUF1 (N12892, N12884);
not NOT1 (N12893, N12892);
and AND3 (N12894, N12878, N3379, N6871);
and AND3 (N12895, N12889, N3901, N1715);
buf BUF1 (N12896, N12879);
nand NAND4 (N12897, N12869, N6433, N8871, N9684);
nand NAND3 (N12898, N12891, N6359, N1108);
buf BUF1 (N12899, N12895);
or OR2 (N12900, N12896, N909);
or OR2 (N12901, N12897, N7534);
and AND2 (N12902, N12888, N6466);
and AND2 (N12903, N12902, N12505);
xor XOR2 (N12904, N12881, N257);
buf BUF1 (N12905, N12904);
nor NOR3 (N12906, N12901, N3566, N6324);
and AND3 (N12907, N12898, N6542, N10062);
and AND3 (N12908, N12907, N1189, N5778);
nor NOR4 (N12909, N12900, N6544, N12714, N10192);
xor XOR2 (N12910, N12886, N9623);
or OR2 (N12911, N12906, N9491);
not NOT1 (N12912, N12893);
nand NAND2 (N12913, N12899, N6896);
buf BUF1 (N12914, N12910);
not NOT1 (N12915, N12913);
not NOT1 (N12916, N12911);
buf BUF1 (N12917, N12909);
nor NOR3 (N12918, N12894, N3299, N3882);
buf BUF1 (N12919, N12914);
nor NOR4 (N12920, N12890, N11050, N3186, N6383);
not NOT1 (N12921, N12918);
and AND4 (N12922, N12912, N2669, N660, N149);
xor XOR2 (N12923, N12903, N705);
or OR3 (N12924, N12908, N11696, N7783);
and AND3 (N12925, N12905, N7958, N12886);
nand NAND3 (N12926, N12923, N299, N12448);
buf BUF1 (N12927, N12920);
not NOT1 (N12928, N12924);
buf BUF1 (N12929, N12915);
not NOT1 (N12930, N12925);
nor NOR4 (N12931, N12930, N3865, N7330, N6515);
nor NOR3 (N12932, N12916, N7906, N12666);
xor XOR2 (N12933, N12927, N6820);
xor XOR2 (N12934, N12928, N4190);
and AND3 (N12935, N12921, N7719, N1978);
xor XOR2 (N12936, N12932, N3264);
or OR3 (N12937, N12931, N11056, N10916);
not NOT1 (N12938, N12937);
nor NOR4 (N12939, N12926, N11018, N12000, N9321);
nand NAND3 (N12940, N12922, N7341, N6724);
buf BUF1 (N12941, N12934);
not NOT1 (N12942, N12939);
xor XOR2 (N12943, N12936, N12428);
or OR2 (N12944, N12943, N7519);
buf BUF1 (N12945, N12933);
nor NOR3 (N12946, N12919, N7689, N2175);
buf BUF1 (N12947, N12941);
buf BUF1 (N12948, N12938);
nor NOR2 (N12949, N12945, N4589);
and AND4 (N12950, N12935, N10983, N12796, N6096);
not NOT1 (N12951, N12949);
buf BUF1 (N12952, N12951);
and AND4 (N12953, N12947, N2215, N12865, N3559);
nand NAND3 (N12954, N12942, N7251, N8405);
xor XOR2 (N12955, N12946, N9571);
nor NOR2 (N12956, N12940, N5302);
not NOT1 (N12957, N12953);
nand NAND4 (N12958, N12944, N6004, N12731, N6214);
not NOT1 (N12959, N12956);
or OR2 (N12960, N12948, N9828);
buf BUF1 (N12961, N12952);
nor NOR2 (N12962, N12958, N3466);
buf BUF1 (N12963, N12917);
and AND4 (N12964, N12959, N10717, N4088, N3);
buf BUF1 (N12965, N12950);
not NOT1 (N12966, N12957);
xor XOR2 (N12967, N12955, N9289);
and AND3 (N12968, N12964, N9706, N11515);
xor XOR2 (N12969, N12963, N12072);
xor XOR2 (N12970, N12954, N4995);
or OR4 (N12971, N12961, N8351, N9970, N1764);
and AND2 (N12972, N12966, N4535);
buf BUF1 (N12973, N12971);
not NOT1 (N12974, N12962);
nor NOR4 (N12975, N12974, N556, N9299, N12336);
nand NAND4 (N12976, N12967, N8560, N12459, N858);
nor NOR4 (N12977, N12929, N3952, N12523, N6394);
and AND3 (N12978, N12970, N3590, N915);
or OR2 (N12979, N12975, N4267);
nor NOR3 (N12980, N12973, N5976, N7621);
not NOT1 (N12981, N12965);
buf BUF1 (N12982, N12977);
not NOT1 (N12983, N12969);
and AND4 (N12984, N12979, N4535, N5193, N5803);
nand NAND3 (N12985, N12968, N5298, N578);
not NOT1 (N12986, N12978);
buf BUF1 (N12987, N12981);
and AND2 (N12988, N12986, N11612);
nor NOR4 (N12989, N12980, N5977, N1721, N5124);
nor NOR4 (N12990, N12989, N8927, N2734, N4377);
nand NAND3 (N12991, N12990, N6818, N12276);
xor XOR2 (N12992, N12976, N575);
or OR2 (N12993, N12983, N9866);
and AND4 (N12994, N12960, N6002, N9830, N9551);
and AND4 (N12995, N12994, N5773, N10572, N4475);
not NOT1 (N12996, N12982);
nor NOR4 (N12997, N12996, N9965, N12966, N7702);
xor XOR2 (N12998, N12991, N8081);
and AND4 (N12999, N12997, N6615, N9610, N4722);
not NOT1 (N13000, N12984);
xor XOR2 (N13001, N12993, N11140);
and AND4 (N13002, N12987, N7914, N9781, N7698);
buf BUF1 (N13003, N12995);
and AND3 (N13004, N12985, N306, N891);
buf BUF1 (N13005, N12999);
buf BUF1 (N13006, N13001);
not NOT1 (N13007, N12972);
not NOT1 (N13008, N13005);
nor NOR4 (N13009, N12992, N6626, N9664, N784);
xor XOR2 (N13010, N12988, N3724);
nand NAND3 (N13011, N13010, N7281, N11420);
buf BUF1 (N13012, N13008);
not NOT1 (N13013, N13003);
or OR4 (N13014, N13013, N1733, N614, N12980);
buf BUF1 (N13015, N13012);
nand NAND3 (N13016, N13009, N8448, N3061);
buf BUF1 (N13017, N13000);
not NOT1 (N13018, N13002);
xor XOR2 (N13019, N13007, N607);
nand NAND4 (N13020, N13017, N7512, N8473, N4891);
or OR3 (N13021, N13011, N3158, N8575);
or OR2 (N13022, N13006, N7069);
xor XOR2 (N13023, N13015, N1028);
and AND4 (N13024, N13020, N9949, N4647, N2589);
nand NAND2 (N13025, N13004, N4748);
not NOT1 (N13026, N13025);
nor NOR4 (N13027, N13024, N1790, N7936, N9375);
and AND4 (N13028, N13021, N3863, N1499, N4463);
and AND4 (N13029, N13023, N11499, N1272, N8809);
or OR2 (N13030, N13027, N6725);
buf BUF1 (N13031, N13029);
nor NOR2 (N13032, N13031, N5837);
nor NOR3 (N13033, N12998, N11016, N5617);
buf BUF1 (N13034, N13022);
xor XOR2 (N13035, N13034, N4090);
not NOT1 (N13036, N13028);
nand NAND2 (N13037, N13014, N6431);
nand NAND2 (N13038, N13030, N11486);
and AND2 (N13039, N13016, N12570);
xor XOR2 (N13040, N13018, N8818);
nor NOR3 (N13041, N13037, N1175, N4400);
and AND4 (N13042, N13039, N9037, N11201, N3586);
xor XOR2 (N13043, N13019, N9235);
buf BUF1 (N13044, N13032);
xor XOR2 (N13045, N13026, N2474);
buf BUF1 (N13046, N13035);
not NOT1 (N13047, N13044);
xor XOR2 (N13048, N13033, N3532);
nand NAND4 (N13049, N13042, N4687, N1984, N6083);
nand NAND2 (N13050, N13046, N8461);
nor NOR4 (N13051, N13036, N10823, N12898, N10830);
nor NOR2 (N13052, N13041, N7244);
nor NOR4 (N13053, N13038, N1564, N2318, N2808);
buf BUF1 (N13054, N13048);
not NOT1 (N13055, N13049);
xor XOR2 (N13056, N13045, N8662);
nor NOR4 (N13057, N13047, N4030, N652, N4402);
xor XOR2 (N13058, N13053, N5033);
or OR4 (N13059, N13052, N6908, N7788, N8574);
and AND2 (N13060, N13040, N11099);
nand NAND3 (N13061, N13057, N8863, N3773);
and AND3 (N13062, N13060, N8947, N12571);
nand NAND3 (N13063, N13061, N1085, N6916);
and AND4 (N13064, N13063, N12795, N5336, N10346);
not NOT1 (N13065, N13064);
xor XOR2 (N13066, N13059, N6283);
xor XOR2 (N13067, N13065, N4207);
not NOT1 (N13068, N13051);
and AND3 (N13069, N13058, N6328, N3026);
nor NOR3 (N13070, N13043, N4380, N2596);
or OR4 (N13071, N13054, N3090, N12054, N2157);
or OR3 (N13072, N13069, N3570, N1110);
and AND3 (N13073, N13056, N12081, N8193);
buf BUF1 (N13074, N13071);
buf BUF1 (N13075, N13074);
nor NOR2 (N13076, N13050, N12132);
nand NAND2 (N13077, N13055, N8159);
nand NAND3 (N13078, N13066, N8712, N12163);
not NOT1 (N13079, N13072);
nor NOR3 (N13080, N13075, N4728, N11483);
buf BUF1 (N13081, N13079);
not NOT1 (N13082, N13068);
nor NOR3 (N13083, N13082, N6061, N7949);
xor XOR2 (N13084, N13083, N12215);
buf BUF1 (N13085, N13067);
xor XOR2 (N13086, N13070, N4171);
and AND3 (N13087, N13078, N127, N11342);
not NOT1 (N13088, N13076);
not NOT1 (N13089, N13084);
nand NAND2 (N13090, N13073, N4951);
buf BUF1 (N13091, N13077);
not NOT1 (N13092, N13080);
not NOT1 (N13093, N13086);
or OR3 (N13094, N13093, N11707, N284);
buf BUF1 (N13095, N13062);
nand NAND3 (N13096, N13085, N1646, N622);
buf BUF1 (N13097, N13081);
buf BUF1 (N13098, N13097);
or OR4 (N13099, N13089, N1118, N10305, N11600);
and AND3 (N13100, N13087, N4943, N10913);
or OR3 (N13101, N13094, N11777, N11670);
or OR2 (N13102, N13101, N4330);
and AND3 (N13103, N13099, N3104, N12728);
nor NOR3 (N13104, N13100, N82, N12787);
or OR4 (N13105, N13095, N2812, N11535, N7296);
not NOT1 (N13106, N13090);
buf BUF1 (N13107, N13088);
and AND3 (N13108, N13092, N8542, N9220);
buf BUF1 (N13109, N13102);
not NOT1 (N13110, N13104);
nand NAND4 (N13111, N13107, N10794, N3957, N9336);
xor XOR2 (N13112, N13096, N3642);
and AND4 (N13113, N13109, N11506, N1094, N1176);
not NOT1 (N13114, N13098);
nor NOR3 (N13115, N13111, N5320, N4781);
or OR3 (N13116, N13115, N2097, N12254);
not NOT1 (N13117, N13091);
buf BUF1 (N13118, N13103);
not NOT1 (N13119, N13106);
and AND3 (N13120, N13110, N7629, N5268);
nand NAND3 (N13121, N13112, N9022, N7672);
not NOT1 (N13122, N13113);
buf BUF1 (N13123, N13108);
xor XOR2 (N13124, N13117, N5557);
nor NOR2 (N13125, N13120, N11762);
buf BUF1 (N13126, N13105);
and AND3 (N13127, N13118, N4523, N192);
nor NOR2 (N13128, N13116, N8378);
or OR4 (N13129, N13122, N11472, N9525, N931);
not NOT1 (N13130, N13129);
buf BUF1 (N13131, N13126);
and AND2 (N13132, N13124, N9368);
and AND3 (N13133, N13114, N11223, N1192);
nand NAND2 (N13134, N13119, N6795);
not NOT1 (N13135, N13125);
xor XOR2 (N13136, N13131, N7665);
nand NAND2 (N13137, N13136, N1155);
and AND4 (N13138, N13128, N3356, N5178, N7132);
nand NAND2 (N13139, N13138, N4229);
not NOT1 (N13140, N13127);
xor XOR2 (N13141, N13135, N4808);
or OR4 (N13142, N13139, N11248, N4840, N7179);
xor XOR2 (N13143, N13132, N1837);
nand NAND2 (N13144, N13143, N2457);
not NOT1 (N13145, N13144);
and AND4 (N13146, N13134, N12573, N8790, N10097);
xor XOR2 (N13147, N13123, N3940);
nor NOR4 (N13148, N13146, N10335, N9893, N9385);
nor NOR2 (N13149, N13137, N11422);
not NOT1 (N13150, N13142);
and AND3 (N13151, N13130, N9059, N1856);
xor XOR2 (N13152, N13140, N5002);
nand NAND4 (N13153, N13149, N12990, N6578, N5464);
buf BUF1 (N13154, N13145);
buf BUF1 (N13155, N13154);
or OR4 (N13156, N13151, N7928, N3927, N8891);
and AND2 (N13157, N13156, N5663);
and AND3 (N13158, N13121, N6274, N5140);
and AND4 (N13159, N13148, N3599, N12277, N3915);
xor XOR2 (N13160, N13133, N2371);
nor NOR4 (N13161, N13155, N9021, N7951, N10470);
xor XOR2 (N13162, N13157, N11311);
not NOT1 (N13163, N13147);
nand NAND4 (N13164, N13141, N11046, N1781, N9912);
xor XOR2 (N13165, N13153, N3548);
or OR3 (N13166, N13164, N8745, N4742);
nor NOR4 (N13167, N13166, N9580, N974, N3591);
buf BUF1 (N13168, N13150);
buf BUF1 (N13169, N13152);
nor NOR4 (N13170, N13158, N6031, N11143, N2140);
not NOT1 (N13171, N13163);
nor NOR4 (N13172, N13168, N7162, N3916, N3775);
and AND4 (N13173, N13171, N10545, N7234, N3188);
or OR3 (N13174, N13162, N694, N1596);
and AND4 (N13175, N13170, N3507, N12510, N830);
buf BUF1 (N13176, N13160);
not NOT1 (N13177, N13159);
nor NOR2 (N13178, N13175, N5054);
and AND4 (N13179, N13169, N12634, N4119, N10510);
and AND3 (N13180, N13176, N508, N5514);
buf BUF1 (N13181, N13167);
buf BUF1 (N13182, N13174);
not NOT1 (N13183, N13182);
xor XOR2 (N13184, N13183, N5829);
or OR4 (N13185, N13184, N466, N1389, N6826);
or OR4 (N13186, N13172, N6266, N10975, N2917);
not NOT1 (N13187, N13179);
xor XOR2 (N13188, N13173, N5022);
or OR2 (N13189, N13188, N10490);
nand NAND3 (N13190, N13189, N5243, N2459);
buf BUF1 (N13191, N13177);
nand NAND3 (N13192, N13161, N1719, N5091);
xor XOR2 (N13193, N13180, N9255);
not NOT1 (N13194, N13193);
and AND4 (N13195, N13192, N9033, N145, N8936);
buf BUF1 (N13196, N13185);
and AND3 (N13197, N13191, N1487, N7816);
xor XOR2 (N13198, N13165, N3230);
xor XOR2 (N13199, N13186, N8071);
buf BUF1 (N13200, N13196);
nand NAND3 (N13201, N13199, N9057, N13);
buf BUF1 (N13202, N13194);
not NOT1 (N13203, N13200);
not NOT1 (N13204, N13197);
xor XOR2 (N13205, N13198, N11278);
xor XOR2 (N13206, N13205, N2105);
buf BUF1 (N13207, N13181);
or OR3 (N13208, N13178, N12782, N2460);
not NOT1 (N13209, N13187);
nand NAND3 (N13210, N13208, N10820, N10849);
buf BUF1 (N13211, N13210);
or OR2 (N13212, N13206, N5182);
and AND4 (N13213, N13212, N6063, N4385, N12140);
not NOT1 (N13214, N13190);
nand NAND4 (N13215, N13214, N4301, N12691, N944);
xor XOR2 (N13216, N13211, N12402);
nand NAND4 (N13217, N13213, N6258, N4639, N705);
not NOT1 (N13218, N13201);
nor NOR4 (N13219, N13218, N9592, N5508, N3970);
and AND3 (N13220, N13207, N3411, N2881);
nand NAND3 (N13221, N13204, N8288, N8623);
buf BUF1 (N13222, N13209);
or OR3 (N13223, N13203, N10539, N3850);
and AND2 (N13224, N13223, N5977);
or OR3 (N13225, N13219, N5615, N5429);
buf BUF1 (N13226, N13195);
and AND3 (N13227, N13215, N2262, N11694);
nand NAND2 (N13228, N13220, N8571);
nor NOR2 (N13229, N13225, N1908);
xor XOR2 (N13230, N13217, N1090);
or OR3 (N13231, N13228, N11708, N8337);
not NOT1 (N13232, N13224);
nor NOR3 (N13233, N13226, N6110, N11487);
or OR2 (N13234, N13233, N12464);
nand NAND4 (N13235, N13232, N13081, N1274, N3442);
nand NAND2 (N13236, N13231, N12822);
and AND3 (N13237, N13222, N2841, N10629);
nand NAND3 (N13238, N13236, N1395, N8332);
buf BUF1 (N13239, N13230);
buf BUF1 (N13240, N13229);
nor NOR2 (N13241, N13202, N7805);
nand NAND4 (N13242, N13237, N6285, N9595, N4877);
or OR4 (N13243, N13240, N12704, N7931, N106);
nor NOR3 (N13244, N13227, N6370, N4381);
nor NOR3 (N13245, N13242, N554, N5470);
buf BUF1 (N13246, N13239);
and AND2 (N13247, N13221, N12859);
or OR3 (N13248, N13244, N2614, N6590);
or OR4 (N13249, N13243, N12785, N1330, N1238);
nor NOR3 (N13250, N13216, N12517, N4714);
nor NOR3 (N13251, N13246, N2606, N13146);
buf BUF1 (N13252, N13251);
buf BUF1 (N13253, N13238);
nand NAND2 (N13254, N13248, N7213);
or OR3 (N13255, N13250, N119, N11649);
and AND3 (N13256, N13245, N9277, N3429);
or OR3 (N13257, N13254, N10110, N7801);
not NOT1 (N13258, N13249);
buf BUF1 (N13259, N13234);
xor XOR2 (N13260, N13255, N9269);
or OR2 (N13261, N13247, N12250);
and AND3 (N13262, N13235, N4033, N10423);
not NOT1 (N13263, N13262);
not NOT1 (N13264, N13263);
and AND4 (N13265, N13241, N8611, N9186, N514);
buf BUF1 (N13266, N13252);
nand NAND4 (N13267, N13259, N5123, N920, N5398);
nor NOR2 (N13268, N13266, N5621);
or OR2 (N13269, N13267, N855);
buf BUF1 (N13270, N13260);
and AND3 (N13271, N13261, N11361, N4892);
nand NAND4 (N13272, N13271, N1356, N11605, N6739);
xor XOR2 (N13273, N13257, N5837);
or OR4 (N13274, N13256, N219, N278, N1279);
nand NAND3 (N13275, N13269, N3516, N5778);
nor NOR4 (N13276, N13268, N1619, N1576, N4179);
nor NOR4 (N13277, N13253, N5800, N4612, N4596);
nand NAND2 (N13278, N13264, N6561);
not NOT1 (N13279, N13270);
nor NOR2 (N13280, N13274, N11937);
xor XOR2 (N13281, N13280, N3484);
nand NAND4 (N13282, N13275, N5005, N12831, N7095);
buf BUF1 (N13283, N13277);
and AND4 (N13284, N13265, N8792, N10162, N8492);
not NOT1 (N13285, N13273);
not NOT1 (N13286, N13279);
xor XOR2 (N13287, N13272, N388);
and AND4 (N13288, N13278, N11819, N6273, N11501);
xor XOR2 (N13289, N13281, N3235);
and AND3 (N13290, N13286, N12221, N9997);
not NOT1 (N13291, N13285);
or OR3 (N13292, N13283, N7124, N12995);
nand NAND4 (N13293, N13258, N12631, N4806, N8922);
or OR2 (N13294, N13284, N12664);
or OR4 (N13295, N13288, N6128, N11769, N5077);
and AND2 (N13296, N13293, N1714);
nor NOR4 (N13297, N13295, N10134, N9215, N9120);
or OR2 (N13298, N13296, N6048);
or OR4 (N13299, N13294, N4505, N7274, N6074);
and AND2 (N13300, N13297, N6934);
buf BUF1 (N13301, N13291);
buf BUF1 (N13302, N13300);
not NOT1 (N13303, N13290);
nand NAND4 (N13304, N13276, N10436, N11323, N4376);
or OR2 (N13305, N13289, N1449);
nor NOR2 (N13306, N13303, N3408);
buf BUF1 (N13307, N13304);
or OR4 (N13308, N13301, N10094, N30, N2117);
nor NOR3 (N13309, N13292, N1038, N7523);
nand NAND3 (N13310, N13307, N5527, N13102);
nand NAND3 (N13311, N13308, N2187, N1355);
nand NAND3 (N13312, N13298, N6671, N12871);
nand NAND2 (N13313, N13305, N4567);
or OR2 (N13314, N13306, N8701);
or OR2 (N13315, N13314, N790);
nor NOR2 (N13316, N13282, N11455);
nor NOR2 (N13317, N13302, N6086);
xor XOR2 (N13318, N13316, N12057);
nor NOR3 (N13319, N13315, N7386, N8509);
and AND2 (N13320, N13319, N6332);
nand NAND3 (N13321, N13317, N12541, N2812);
nand NAND3 (N13322, N13299, N12556, N3809);
nor NOR3 (N13323, N13310, N9593, N13144);
nand NAND4 (N13324, N13311, N4504, N5082, N9334);
buf BUF1 (N13325, N13320);
not NOT1 (N13326, N13312);
nor NOR4 (N13327, N13326, N9960, N1596, N3686);
and AND3 (N13328, N13322, N5676, N7475);
nand NAND3 (N13329, N13309, N12977, N13001);
buf BUF1 (N13330, N13318);
or OR4 (N13331, N13328, N4616, N12314, N9650);
buf BUF1 (N13332, N13324);
and AND2 (N13333, N13323, N343);
or OR3 (N13334, N13313, N10171, N12704);
or OR3 (N13335, N13334, N12905, N12709);
or OR2 (N13336, N13327, N8817);
nand NAND3 (N13337, N13330, N12382, N5608);
or OR2 (N13338, N13287, N10079);
buf BUF1 (N13339, N13333);
xor XOR2 (N13340, N13331, N1001);
nor NOR2 (N13341, N13339, N9662);
xor XOR2 (N13342, N13337, N12705);
or OR3 (N13343, N13329, N4116, N10408);
nand NAND3 (N13344, N13338, N8769, N2298);
not NOT1 (N13345, N13344);
xor XOR2 (N13346, N13343, N3214);
and AND3 (N13347, N13336, N7841, N12065);
buf BUF1 (N13348, N13342);
buf BUF1 (N13349, N13347);
nor NOR4 (N13350, N13335, N7527, N5544, N7457);
not NOT1 (N13351, N13332);
nand NAND2 (N13352, N13351, N4882);
buf BUF1 (N13353, N13349);
buf BUF1 (N13354, N13345);
and AND3 (N13355, N13348, N766, N5893);
buf BUF1 (N13356, N13353);
and AND4 (N13357, N13356, N3527, N7555, N5530);
and AND4 (N13358, N13346, N5786, N10432, N1372);
nor NOR4 (N13359, N13350, N7151, N5926, N703);
and AND2 (N13360, N13354, N12136);
nor NOR2 (N13361, N13355, N9726);
nand NAND3 (N13362, N13321, N2117, N9983);
buf BUF1 (N13363, N13358);
and AND3 (N13364, N13363, N4566, N7838);
nor NOR4 (N13365, N13341, N11241, N10824, N2198);
or OR3 (N13366, N13325, N8141, N10166);
xor XOR2 (N13367, N13361, N3154);
xor XOR2 (N13368, N13352, N11451);
or OR3 (N13369, N13359, N1126, N9015);
nor NOR3 (N13370, N13367, N12527, N5139);
nand NAND3 (N13371, N13357, N12880, N5595);
not NOT1 (N13372, N13340);
not NOT1 (N13373, N13369);
buf BUF1 (N13374, N13364);
buf BUF1 (N13375, N13370);
or OR3 (N13376, N13374, N993, N929);
not NOT1 (N13377, N13362);
and AND2 (N13378, N13372, N9251);
and AND2 (N13379, N13375, N1631);
xor XOR2 (N13380, N13365, N2791);
buf BUF1 (N13381, N13377);
and AND4 (N13382, N13360, N12659, N2317, N6756);
nor NOR3 (N13383, N13378, N13060, N6915);
or OR3 (N13384, N13381, N5148, N6408);
buf BUF1 (N13385, N13380);
and AND4 (N13386, N13384, N6985, N1830, N13136);
xor XOR2 (N13387, N13373, N8284);
not NOT1 (N13388, N13387);
nand NAND3 (N13389, N13366, N358, N12037);
xor XOR2 (N13390, N13385, N4955);
nor NOR2 (N13391, N13390, N8971);
or OR3 (N13392, N13383, N12170, N8645);
nand NAND3 (N13393, N13379, N3301, N13290);
not NOT1 (N13394, N13382);
buf BUF1 (N13395, N13376);
xor XOR2 (N13396, N13386, N7201);
xor XOR2 (N13397, N13395, N6455);
not NOT1 (N13398, N13397);
or OR2 (N13399, N13393, N5630);
not NOT1 (N13400, N13396);
buf BUF1 (N13401, N13388);
buf BUF1 (N13402, N13401);
nor NOR2 (N13403, N13392, N1754);
xor XOR2 (N13404, N13399, N6001);
not NOT1 (N13405, N13400);
not NOT1 (N13406, N13398);
not NOT1 (N13407, N13403);
nand NAND4 (N13408, N13394, N4860, N7420, N13406);
xor XOR2 (N13409, N12502, N516);
xor XOR2 (N13410, N13404, N2324);
buf BUF1 (N13411, N13402);
or OR3 (N13412, N13389, N6216, N9822);
xor XOR2 (N13413, N13412, N8407);
not NOT1 (N13414, N13409);
buf BUF1 (N13415, N13411);
or OR3 (N13416, N13368, N12790, N8671);
and AND3 (N13417, N13407, N9853, N8772);
nor NOR3 (N13418, N13415, N11518, N1199);
nor NOR3 (N13419, N13408, N7173, N2598);
not NOT1 (N13420, N13418);
xor XOR2 (N13421, N13391, N3183);
or OR4 (N13422, N13414, N5479, N5274, N9537);
not NOT1 (N13423, N13421);
nor NOR2 (N13424, N13419, N9119);
buf BUF1 (N13425, N13423);
buf BUF1 (N13426, N13410);
and AND3 (N13427, N13426, N1793, N6061);
xor XOR2 (N13428, N13427, N13114);
nand NAND3 (N13429, N13422, N5269, N9935);
nor NOR3 (N13430, N13417, N8311, N9826);
not NOT1 (N13431, N13428);
not NOT1 (N13432, N13413);
xor XOR2 (N13433, N13429, N6937);
buf BUF1 (N13434, N13424);
or OR3 (N13435, N13405, N8525, N860);
or OR4 (N13436, N13416, N11551, N7463, N12550);
buf BUF1 (N13437, N13436);
nor NOR2 (N13438, N13437, N11490);
buf BUF1 (N13439, N13434);
and AND2 (N13440, N13371, N4948);
nor NOR2 (N13441, N13430, N5705);
and AND3 (N13442, N13425, N1950, N9586);
not NOT1 (N13443, N13441);
xor XOR2 (N13444, N13435, N9359);
nor NOR4 (N13445, N13420, N8410, N1112, N12743);
not NOT1 (N13446, N13440);
nand NAND3 (N13447, N13445, N11196, N1387);
not NOT1 (N13448, N13433);
buf BUF1 (N13449, N13448);
xor XOR2 (N13450, N13438, N4440);
not NOT1 (N13451, N13431);
xor XOR2 (N13452, N13446, N4174);
nor NOR2 (N13453, N13432, N618);
not NOT1 (N13454, N13439);
not NOT1 (N13455, N13449);
and AND3 (N13456, N13450, N10250, N3510);
xor XOR2 (N13457, N13444, N2497);
or OR4 (N13458, N13456, N5477, N11639, N405);
nand NAND3 (N13459, N13442, N10200, N1109);
and AND4 (N13460, N13455, N9956, N6685, N5189);
xor XOR2 (N13461, N13457, N7135);
not NOT1 (N13462, N13447);
nand NAND3 (N13463, N13443, N4663, N9274);
nor NOR4 (N13464, N13454, N9910, N10067, N6180);
nand NAND3 (N13465, N13459, N11552, N6015);
and AND4 (N13466, N13462, N6786, N6429, N8754);
not NOT1 (N13467, N13461);
or OR2 (N13468, N13465, N5424);
xor XOR2 (N13469, N13460, N10828);
and AND2 (N13470, N13467, N12157);
buf BUF1 (N13471, N13463);
nor NOR2 (N13472, N13469, N2137);
and AND2 (N13473, N13451, N12194);
xor XOR2 (N13474, N13470, N681);
xor XOR2 (N13475, N13464, N5079);
buf BUF1 (N13476, N13468);
or OR4 (N13477, N13475, N1490, N1085, N3364);
and AND3 (N13478, N13452, N2795, N3937);
xor XOR2 (N13479, N13473, N10212);
and AND2 (N13480, N13478, N6613);
buf BUF1 (N13481, N13479);
nor NOR3 (N13482, N13477, N6002, N11062);
buf BUF1 (N13483, N13482);
nand NAND3 (N13484, N13474, N2399, N13140);
nand NAND4 (N13485, N13472, N5446, N9020, N10004);
or OR2 (N13486, N13481, N10997);
buf BUF1 (N13487, N13471);
nand NAND2 (N13488, N13485, N10784);
nor NOR4 (N13489, N13453, N3922, N53, N815);
buf BUF1 (N13490, N13487);
nand NAND2 (N13491, N13488, N143);
nor NOR3 (N13492, N13483, N2970, N1696);
nor NOR2 (N13493, N13480, N4254);
nand NAND3 (N13494, N13458, N3725, N8310);
or OR4 (N13495, N13490, N7110, N3119, N1137);
xor XOR2 (N13496, N13493, N2293);
nand NAND4 (N13497, N13492, N654, N12244, N6456);
nand NAND4 (N13498, N13497, N11650, N6300, N11554);
nor NOR2 (N13499, N13498, N3522);
not NOT1 (N13500, N13476);
xor XOR2 (N13501, N13486, N4524);
nand NAND2 (N13502, N13499, N2282);
not NOT1 (N13503, N13496);
nand NAND4 (N13504, N13495, N4599, N8823, N11288);
and AND4 (N13505, N13491, N3988, N101, N3786);
buf BUF1 (N13506, N13489);
nor NOR2 (N13507, N13484, N694);
buf BUF1 (N13508, N13494);
xor XOR2 (N13509, N13507, N1787);
or OR4 (N13510, N13509, N1763, N5671, N1922);
xor XOR2 (N13511, N13510, N10947);
xor XOR2 (N13512, N13502, N6194);
and AND3 (N13513, N13505, N1366, N8124);
buf BUF1 (N13514, N13511);
buf BUF1 (N13515, N13513);
nand NAND2 (N13516, N13512, N1383);
xor XOR2 (N13517, N13516, N13204);
buf BUF1 (N13518, N13514);
not NOT1 (N13519, N13500);
nand NAND2 (N13520, N13466, N5310);
nor NOR3 (N13521, N13515, N11328, N3218);
buf BUF1 (N13522, N13521);
nor NOR2 (N13523, N13520, N10780);
nand NAND3 (N13524, N13506, N10738, N6558);
and AND4 (N13525, N13522, N6384, N13322, N10441);
buf BUF1 (N13526, N13525);
buf BUF1 (N13527, N13501);
not NOT1 (N13528, N13504);
not NOT1 (N13529, N13526);
buf BUF1 (N13530, N13508);
nand NAND4 (N13531, N13524, N3082, N4005, N10197);
buf BUF1 (N13532, N13503);
nand NAND2 (N13533, N13519, N4408);
buf BUF1 (N13534, N13517);
nand NAND2 (N13535, N13532, N10549);
xor XOR2 (N13536, N13531, N832);
nand NAND3 (N13537, N13518, N7159, N658);
and AND2 (N13538, N13533, N2746);
nor NOR4 (N13539, N13523, N7602, N11058, N7305);
or OR4 (N13540, N13536, N8043, N8751, N8597);
buf BUF1 (N13541, N13535);
and AND3 (N13542, N13537, N7627, N1191);
or OR2 (N13543, N13539, N3249);
xor XOR2 (N13544, N13540, N13358);
xor XOR2 (N13545, N13534, N9766);
nor NOR3 (N13546, N13542, N694, N12673);
buf BUF1 (N13547, N13543);
or OR2 (N13548, N13527, N632);
nand NAND3 (N13549, N13529, N13437, N4791);
or OR4 (N13550, N13545, N6914, N5836, N11126);
nand NAND2 (N13551, N13528, N11403);
and AND4 (N13552, N13544, N4695, N2037, N12726);
xor XOR2 (N13553, N13548, N1485);
not NOT1 (N13554, N13553);
xor XOR2 (N13555, N13549, N10496);
or OR3 (N13556, N13552, N3717, N4421);
xor XOR2 (N13557, N13554, N1518);
buf BUF1 (N13558, N13551);
and AND2 (N13559, N13547, N4902);
buf BUF1 (N13560, N13555);
buf BUF1 (N13561, N13560);
xor XOR2 (N13562, N13557, N2742);
buf BUF1 (N13563, N13556);
buf BUF1 (N13564, N13559);
not NOT1 (N13565, N13538);
buf BUF1 (N13566, N13558);
and AND4 (N13567, N13550, N7341, N4180, N5231);
nor NOR4 (N13568, N13541, N52, N3959, N12486);
and AND3 (N13569, N13546, N4591, N12803);
nor NOR2 (N13570, N13567, N6126);
not NOT1 (N13571, N13563);
not NOT1 (N13572, N13571);
not NOT1 (N13573, N13530);
buf BUF1 (N13574, N13561);
nor NOR3 (N13575, N13572, N11349, N8103);
buf BUF1 (N13576, N13568);
buf BUF1 (N13577, N13564);
xor XOR2 (N13578, N13576, N9094);
buf BUF1 (N13579, N13573);
nand NAND4 (N13580, N13566, N3647, N57, N6836);
or OR4 (N13581, N13569, N12706, N7584, N2374);
and AND2 (N13582, N13577, N8350);
and AND2 (N13583, N13562, N8317);
xor XOR2 (N13584, N13578, N10473);
and AND2 (N13585, N13570, N10752);
nand NAND4 (N13586, N13565, N6722, N3978, N1169);
nand NAND4 (N13587, N13579, N10802, N2311, N3034);
and AND4 (N13588, N13587, N6873, N7383, N3067);
not NOT1 (N13589, N13580);
and AND2 (N13590, N13581, N154);
or OR4 (N13591, N13588, N1779, N13479, N10367);
buf BUF1 (N13592, N13583);
and AND2 (N13593, N13582, N11836);
buf BUF1 (N13594, N13585);
xor XOR2 (N13595, N13575, N699);
nand NAND4 (N13596, N13574, N1091, N9333, N4621);
nor NOR3 (N13597, N13593, N9385, N10980);
nand NAND4 (N13598, N13590, N9477, N13307, N3110);
nor NOR3 (N13599, N13595, N2250, N3881);
or OR4 (N13600, N13589, N9222, N6935, N9373);
not NOT1 (N13601, N13592);
not NOT1 (N13602, N13597);
nand NAND2 (N13603, N13600, N7139);
xor XOR2 (N13604, N13598, N8447);
or OR3 (N13605, N13604, N6525, N1804);
or OR2 (N13606, N13605, N8000);
and AND3 (N13607, N13591, N1162, N7849);
nor NOR3 (N13608, N13586, N11768, N8474);
xor XOR2 (N13609, N13607, N11416);
nand NAND3 (N13610, N13584, N11321, N12278);
nor NOR2 (N13611, N13599, N12066);
and AND4 (N13612, N13596, N10519, N3098, N10736);
and AND4 (N13613, N13594, N12852, N9010, N1034);
and AND3 (N13614, N13612, N7907, N1083);
or OR4 (N13615, N13603, N5334, N9589, N670);
and AND3 (N13616, N13608, N454, N8055);
xor XOR2 (N13617, N13609, N1844);
not NOT1 (N13618, N13606);
buf BUF1 (N13619, N13616);
not NOT1 (N13620, N13613);
nor NOR2 (N13621, N13610, N2573);
buf BUF1 (N13622, N13618);
or OR2 (N13623, N13622, N5012);
buf BUF1 (N13624, N13621);
or OR2 (N13625, N13614, N6359);
buf BUF1 (N13626, N13625);
and AND4 (N13627, N13623, N6478, N5863, N8971);
not NOT1 (N13628, N13611);
or OR4 (N13629, N13627, N5422, N12687, N6531);
and AND3 (N13630, N13619, N5718, N3332);
or OR2 (N13631, N13620, N12122);
or OR3 (N13632, N13628, N8279, N10929);
buf BUF1 (N13633, N13617);
and AND4 (N13634, N13633, N9935, N5834, N4445);
and AND2 (N13635, N13630, N4413);
nand NAND2 (N13636, N13626, N12767);
xor XOR2 (N13637, N13624, N11359);
not NOT1 (N13638, N13601);
nand NAND3 (N13639, N13635, N11264, N13285);
xor XOR2 (N13640, N13634, N6068);
not NOT1 (N13641, N13631);
nor NOR4 (N13642, N13640, N421, N10053, N4826);
and AND2 (N13643, N13638, N5942);
nand NAND2 (N13644, N13632, N8571);
nand NAND4 (N13645, N13643, N11382, N1767, N12117);
or OR3 (N13646, N13637, N4791, N7767);
nor NOR2 (N13647, N13636, N13373);
nor NOR2 (N13648, N13647, N4269);
not NOT1 (N13649, N13639);
and AND4 (N13650, N13642, N7423, N3387, N5393);
xor XOR2 (N13651, N13649, N200);
xor XOR2 (N13652, N13641, N9012);
or OR3 (N13653, N13650, N4737, N6317);
and AND4 (N13654, N13644, N5094, N9870, N6414);
nor NOR2 (N13655, N13653, N11017);
nand NAND2 (N13656, N13602, N1920);
buf BUF1 (N13657, N13656);
nor NOR4 (N13658, N13654, N3158, N3378, N7659);
nor NOR3 (N13659, N13655, N11928, N11974);
xor XOR2 (N13660, N13615, N4962);
not NOT1 (N13661, N13660);
and AND4 (N13662, N13661, N5673, N10771, N12277);
buf BUF1 (N13663, N13645);
nand NAND3 (N13664, N13658, N8437, N6696);
not NOT1 (N13665, N13652);
nand NAND4 (N13666, N13665, N11270, N3443, N8055);
nand NAND4 (N13667, N13648, N4545, N2175, N12084);
or OR2 (N13668, N13646, N12239);
xor XOR2 (N13669, N13659, N9263);
and AND4 (N13670, N13657, N3138, N1176, N12545);
and AND2 (N13671, N13651, N8930);
nor NOR4 (N13672, N13667, N3821, N1213, N4649);
not NOT1 (N13673, N13629);
and AND4 (N13674, N13673, N6704, N957, N6476);
xor XOR2 (N13675, N13671, N8317);
nor NOR3 (N13676, N13666, N8337, N5941);
xor XOR2 (N13677, N13662, N1638);
nand NAND3 (N13678, N13664, N892, N10134);
nand NAND4 (N13679, N13669, N8925, N9814, N8986);
or OR3 (N13680, N13676, N1438, N8476);
xor XOR2 (N13681, N13674, N5470);
and AND2 (N13682, N13672, N3966);
or OR2 (N13683, N13682, N13219);
or OR4 (N13684, N13681, N6756, N97, N12372);
and AND2 (N13685, N13670, N1417);
buf BUF1 (N13686, N13683);
buf BUF1 (N13687, N13668);
or OR3 (N13688, N13685, N9101, N7921);
or OR3 (N13689, N13684, N4314, N1632);
xor XOR2 (N13690, N13687, N12354);
not NOT1 (N13691, N13690);
xor XOR2 (N13692, N13686, N9355);
xor XOR2 (N13693, N13677, N13043);
nor NOR3 (N13694, N13691, N9240, N8251);
nand NAND2 (N13695, N13693, N7074);
buf BUF1 (N13696, N13680);
nand NAND4 (N13697, N13688, N12989, N10817, N9839);
xor XOR2 (N13698, N13675, N8981);
or OR4 (N13699, N13696, N5419, N2586, N9118);
nor NOR3 (N13700, N13689, N1015, N13107);
nor NOR3 (N13701, N13692, N5606, N9617);
xor XOR2 (N13702, N13678, N11535);
not NOT1 (N13703, N13697);
and AND4 (N13704, N13679, N10583, N874, N13100);
or OR3 (N13705, N13704, N2720, N9413);
nor NOR3 (N13706, N13694, N7234, N10849);
nor NOR3 (N13707, N13698, N1004, N6466);
and AND2 (N13708, N13699, N12293);
buf BUF1 (N13709, N13701);
nand NAND2 (N13710, N13707, N4304);
nor NOR2 (N13711, N13708, N10088);
not NOT1 (N13712, N13706);
xor XOR2 (N13713, N13700, N3110);
buf BUF1 (N13714, N13663);
buf BUF1 (N13715, N13713);
nand NAND2 (N13716, N13705, N9225);
xor XOR2 (N13717, N13716, N6696);
nor NOR4 (N13718, N13702, N1418, N3108, N8036);
not NOT1 (N13719, N13703);
not NOT1 (N13720, N13714);
nand NAND3 (N13721, N13715, N4480, N7339);
and AND2 (N13722, N13710, N6895);
nor NOR3 (N13723, N13721, N10402, N6673);
buf BUF1 (N13724, N13712);
buf BUF1 (N13725, N13711);
nor NOR2 (N13726, N13717, N9447);
nor NOR2 (N13727, N13719, N264);
or OR2 (N13728, N13726, N5144);
nor NOR3 (N13729, N13722, N2672, N13395);
xor XOR2 (N13730, N13718, N11312);
nor NOR2 (N13731, N13729, N9463);
nor NOR4 (N13732, N13720, N2111, N12292, N2042);
xor XOR2 (N13733, N13730, N2467);
or OR3 (N13734, N13709, N10319, N11458);
or OR3 (N13735, N13723, N1971, N1330);
nand NAND2 (N13736, N13727, N3618);
nor NOR4 (N13737, N13735, N2913, N849, N7519);
nand NAND2 (N13738, N13728, N10656);
and AND4 (N13739, N13733, N205, N12904, N12917);
or OR4 (N13740, N13736, N13191, N3789, N7828);
and AND3 (N13741, N13739, N8845, N4852);
not NOT1 (N13742, N13732);
buf BUF1 (N13743, N13738);
or OR4 (N13744, N13743, N7159, N12519, N10778);
and AND3 (N13745, N13724, N303, N8528);
xor XOR2 (N13746, N13744, N13535);
and AND4 (N13747, N13740, N8989, N8831, N5143);
not NOT1 (N13748, N13731);
or OR2 (N13749, N13747, N10992);
not NOT1 (N13750, N13737);
nor NOR3 (N13751, N13734, N8328, N1022);
not NOT1 (N13752, N13745);
nand NAND3 (N13753, N13746, N821, N11997);
nand NAND4 (N13754, N13752, N7048, N8582, N11594);
and AND3 (N13755, N13748, N13365, N2019);
nand NAND3 (N13756, N13751, N5671, N1508);
or OR4 (N13757, N13754, N4832, N10728, N10976);
or OR4 (N13758, N13755, N12596, N5684, N10390);
not NOT1 (N13759, N13756);
and AND4 (N13760, N13753, N10897, N8961, N2810);
nor NOR4 (N13761, N13695, N9885, N7371, N7750);
buf BUF1 (N13762, N13750);
xor XOR2 (N13763, N13760, N4921);
not NOT1 (N13764, N13741);
buf BUF1 (N13765, N13761);
not NOT1 (N13766, N13758);
not NOT1 (N13767, N13759);
nor NOR3 (N13768, N13742, N1870, N7675);
not NOT1 (N13769, N13749);
or OR2 (N13770, N13765, N13696);
buf BUF1 (N13771, N13762);
not NOT1 (N13772, N13766);
or OR2 (N13773, N13770, N10176);
buf BUF1 (N13774, N13725);
not NOT1 (N13775, N13757);
not NOT1 (N13776, N13774);
and AND2 (N13777, N13775, N1950);
or OR2 (N13778, N13772, N9147);
xor XOR2 (N13779, N13763, N7879);
nand NAND2 (N13780, N13771, N1805);
buf BUF1 (N13781, N13777);
xor XOR2 (N13782, N13780, N8140);
not NOT1 (N13783, N13764);
and AND4 (N13784, N13776, N1566, N10347, N144);
not NOT1 (N13785, N13779);
or OR3 (N13786, N13767, N8927, N2792);
nor NOR4 (N13787, N13769, N6812, N12649, N1991);
not NOT1 (N13788, N13787);
nor NOR2 (N13789, N13778, N957);
nor NOR3 (N13790, N13773, N10442, N11836);
or OR2 (N13791, N13768, N458);
xor XOR2 (N13792, N13783, N11170);
xor XOR2 (N13793, N13791, N8);
nor NOR3 (N13794, N13790, N5713, N13478);
and AND3 (N13795, N13789, N8533, N12740);
or OR2 (N13796, N13792, N11465);
or OR3 (N13797, N13795, N13032, N5309);
xor XOR2 (N13798, N13782, N2895);
or OR2 (N13799, N13786, N10515);
nand NAND4 (N13800, N13797, N7391, N8114, N8955);
not NOT1 (N13801, N13781);
not NOT1 (N13802, N13793);
xor XOR2 (N13803, N13785, N6411);
nand NAND3 (N13804, N13794, N12378, N10452);
or OR2 (N13805, N13796, N1067);
or OR2 (N13806, N13804, N12083);
nand NAND3 (N13807, N13803, N2082, N13406);
nand NAND3 (N13808, N13806, N7240, N862);
xor XOR2 (N13809, N13798, N8701);
and AND4 (N13810, N13807, N10745, N927, N4348);
and AND3 (N13811, N13809, N6147, N612);
or OR2 (N13812, N13800, N7611);
not NOT1 (N13813, N13812);
nand NAND3 (N13814, N13810, N9024, N7098);
nor NOR3 (N13815, N13805, N2975, N9325);
or OR4 (N13816, N13815, N13575, N6583, N6087);
and AND4 (N13817, N13799, N5325, N3911, N4899);
xor XOR2 (N13818, N13811, N11880);
nand NAND3 (N13819, N13801, N9404, N2167);
xor XOR2 (N13820, N13814, N1412);
xor XOR2 (N13821, N13784, N13814);
or OR3 (N13822, N13821, N2083, N1982);
buf BUF1 (N13823, N13813);
xor XOR2 (N13824, N13818, N10251);
xor XOR2 (N13825, N13820, N9803);
nor NOR4 (N13826, N13802, N10084, N9283, N6090);
nand NAND2 (N13827, N13823, N4984);
xor XOR2 (N13828, N13816, N177);
or OR4 (N13829, N13822, N12790, N9758, N2278);
or OR4 (N13830, N13808, N6408, N9809, N9474);
buf BUF1 (N13831, N13829);
xor XOR2 (N13832, N13825, N1455);
or OR4 (N13833, N13826, N4357, N9803, N2427);
nor NOR4 (N13834, N13824, N3473, N12944, N408);
nand NAND2 (N13835, N13834, N467);
and AND3 (N13836, N13828, N9596, N13179);
not NOT1 (N13837, N13819);
nand NAND4 (N13838, N13837, N6179, N5661, N9192);
nor NOR3 (N13839, N13817, N13148, N6957);
or OR4 (N13840, N13831, N6943, N6952, N8636);
xor XOR2 (N13841, N13838, N7292);
or OR2 (N13842, N13835, N11648);
or OR4 (N13843, N13830, N11510, N3137, N3671);
xor XOR2 (N13844, N13843, N8356);
xor XOR2 (N13845, N13842, N5251);
and AND2 (N13846, N13833, N2381);
xor XOR2 (N13847, N13832, N5174);
buf BUF1 (N13848, N13847);
buf BUF1 (N13849, N13839);
or OR4 (N13850, N13849, N3262, N8362, N5943);
xor XOR2 (N13851, N13848, N9584);
or OR3 (N13852, N13850, N3200, N10644);
or OR3 (N13853, N13836, N815, N682);
nor NOR3 (N13854, N13827, N6312, N9372);
nand NAND2 (N13855, N13840, N12378);
not NOT1 (N13856, N13851);
nand NAND3 (N13857, N13844, N917, N3131);
buf BUF1 (N13858, N13853);
xor XOR2 (N13859, N13852, N4595);
buf BUF1 (N13860, N13846);
nor NOR3 (N13861, N13860, N3988, N12231);
not NOT1 (N13862, N13788);
nand NAND2 (N13863, N13861, N12186);
and AND4 (N13864, N13856, N4231, N7454, N6109);
not NOT1 (N13865, N13864);
xor XOR2 (N13866, N13863, N13244);
or OR3 (N13867, N13858, N8884, N3366);
xor XOR2 (N13868, N13854, N1874);
and AND3 (N13869, N13867, N4671, N7093);
xor XOR2 (N13870, N13841, N9480);
and AND4 (N13871, N13862, N3158, N5154, N6240);
or OR4 (N13872, N13855, N9337, N13703, N10542);
nand NAND2 (N13873, N13865, N10268);
and AND2 (N13874, N13872, N441);
nor NOR2 (N13875, N13870, N4021);
xor XOR2 (N13876, N13857, N2404);
xor XOR2 (N13877, N13876, N4089);
buf BUF1 (N13878, N13868);
xor XOR2 (N13879, N13877, N8086);
buf BUF1 (N13880, N13878);
nand NAND3 (N13881, N13845, N6901, N2754);
nor NOR4 (N13882, N13866, N6837, N84, N2100);
not NOT1 (N13883, N13879);
buf BUF1 (N13884, N13882);
buf BUF1 (N13885, N13859);
nor NOR2 (N13886, N13873, N5985);
and AND4 (N13887, N13883, N1082, N3408, N10661);
not NOT1 (N13888, N13881);
xor XOR2 (N13889, N13869, N13360);
not NOT1 (N13890, N13880);
xor XOR2 (N13891, N13890, N13174);
and AND2 (N13892, N13884, N7232);
nand NAND4 (N13893, N13886, N6905, N574, N3420);
or OR3 (N13894, N13889, N7814, N12747);
or OR4 (N13895, N13894, N12709, N4197, N12316);
nand NAND2 (N13896, N13895, N5808);
xor XOR2 (N13897, N13887, N7534);
and AND3 (N13898, N13897, N4296, N13165);
not NOT1 (N13899, N13875);
xor XOR2 (N13900, N13893, N5896);
nor NOR3 (N13901, N13874, N10653, N12248);
xor XOR2 (N13902, N13892, N2979);
xor XOR2 (N13903, N13899, N6753);
xor XOR2 (N13904, N13888, N10225);
buf BUF1 (N13905, N13904);
and AND3 (N13906, N13903, N13607, N4117);
nor NOR3 (N13907, N13885, N9405, N11545);
and AND4 (N13908, N13898, N7777, N5386, N13450);
not NOT1 (N13909, N13891);
and AND2 (N13910, N13902, N11127);
xor XOR2 (N13911, N13907, N12046);
buf BUF1 (N13912, N13910);
and AND3 (N13913, N13896, N8642, N1265);
xor XOR2 (N13914, N13905, N5125);
nand NAND3 (N13915, N13913, N3904, N1740);
buf BUF1 (N13916, N13906);
or OR4 (N13917, N13908, N12741, N1685, N6773);
buf BUF1 (N13918, N13915);
or OR4 (N13919, N13914, N6282, N10531, N11745);
not NOT1 (N13920, N13917);
and AND4 (N13921, N13916, N8875, N2679, N1943);
nor NOR3 (N13922, N13901, N3792, N9529);
nor NOR2 (N13923, N13918, N3399);
or OR4 (N13924, N13909, N9376, N4342, N5818);
xor XOR2 (N13925, N13920, N13888);
and AND4 (N13926, N13919, N5799, N1545, N1494);
xor XOR2 (N13927, N13921, N6324);
nor NOR2 (N13928, N13923, N7029);
and AND3 (N13929, N13925, N12916, N11387);
not NOT1 (N13930, N13871);
xor XOR2 (N13931, N13930, N13878);
and AND4 (N13932, N13926, N7626, N10073, N9170);
buf BUF1 (N13933, N13927);
buf BUF1 (N13934, N13924);
buf BUF1 (N13935, N13934);
nor NOR4 (N13936, N13933, N4546, N11168, N10199);
or OR3 (N13937, N13900, N3143, N8302);
buf BUF1 (N13938, N13936);
not NOT1 (N13939, N13937);
or OR2 (N13940, N13938, N4379);
nand NAND4 (N13941, N13911, N10227, N465, N358);
and AND4 (N13942, N13932, N13398, N249, N2417);
and AND3 (N13943, N13942, N1939, N385);
or OR2 (N13944, N13931, N13806);
and AND2 (N13945, N13944, N3983);
nor NOR4 (N13946, N13929, N1135, N10773, N8437);
xor XOR2 (N13947, N13941, N13001);
nor NOR4 (N13948, N13940, N687, N1356, N388);
and AND2 (N13949, N13943, N4611);
and AND2 (N13950, N13945, N9497);
buf BUF1 (N13951, N13912);
and AND2 (N13952, N13948, N862);
nor NOR2 (N13953, N13946, N12999);
xor XOR2 (N13954, N13952, N13682);
nand NAND4 (N13955, N13939, N1851, N11447, N7325);
and AND2 (N13956, N13954, N12269);
nand NAND4 (N13957, N13922, N3792, N5039, N6609);
and AND3 (N13958, N13928, N3226, N7023);
or OR3 (N13959, N13935, N2268, N8917);
or OR4 (N13960, N13956, N7445, N2692, N7550);
nor NOR2 (N13961, N13955, N3938);
buf BUF1 (N13962, N13949);
or OR3 (N13963, N13958, N4076, N9144);
or OR4 (N13964, N13959, N1673, N528, N2893);
xor XOR2 (N13965, N13950, N11407);
and AND2 (N13966, N13951, N13898);
or OR2 (N13967, N13947, N3489);
or OR4 (N13968, N13962, N13414, N13559, N7015);
or OR3 (N13969, N13960, N7928, N633);
nor NOR2 (N13970, N13966, N11603);
nand NAND4 (N13971, N13961, N12204, N8762, N7494);
nor NOR4 (N13972, N13965, N8819, N13254, N1277);
xor XOR2 (N13973, N13953, N8547);
buf BUF1 (N13974, N13970);
buf BUF1 (N13975, N13972);
and AND2 (N13976, N13974, N6749);
not NOT1 (N13977, N13976);
not NOT1 (N13978, N13963);
or OR3 (N13979, N13971, N9494, N10688);
nor NOR3 (N13980, N13977, N13792, N2391);
and AND4 (N13981, N13957, N5605, N10718, N4586);
not NOT1 (N13982, N13964);
buf BUF1 (N13983, N13979);
or OR4 (N13984, N13983, N88, N1224, N5394);
or OR2 (N13985, N13973, N6014);
or OR4 (N13986, N13984, N8904, N12312, N6382);
or OR2 (N13987, N13985, N12263);
xor XOR2 (N13988, N13968, N8838);
nor NOR4 (N13989, N13967, N4988, N3417, N8922);
nor NOR4 (N13990, N13981, N4384, N11109, N7467);
buf BUF1 (N13991, N13986);
nor NOR4 (N13992, N13988, N9587, N6614, N5179);
or OR3 (N13993, N13969, N3920, N3301);
buf BUF1 (N13994, N13991);
not NOT1 (N13995, N13989);
or OR4 (N13996, N13980, N7820, N10187, N1777);
or OR4 (N13997, N13995, N6723, N3707, N13670);
xor XOR2 (N13998, N13982, N3366);
buf BUF1 (N13999, N13996);
and AND3 (N14000, N13978, N2706, N13540);
and AND2 (N14001, N13997, N2172);
and AND2 (N14002, N13998, N324);
and AND2 (N14003, N13975, N13842);
or OR2 (N14004, N13992, N13434);
nor NOR4 (N14005, N13994, N7586, N10811, N9329);
and AND3 (N14006, N13987, N11525, N13821);
nor NOR2 (N14007, N13990, N11963);
nand NAND4 (N14008, N14006, N5209, N9647, N13061);
xor XOR2 (N14009, N14008, N10292);
nand NAND2 (N14010, N14007, N3482);
nand NAND3 (N14011, N14004, N2380, N12586);
not NOT1 (N14012, N14001);
nand NAND3 (N14013, N13993, N8218, N9731);
buf BUF1 (N14014, N14009);
not NOT1 (N14015, N13999);
xor XOR2 (N14016, N14013, N949);
not NOT1 (N14017, N14012);
xor XOR2 (N14018, N14002, N530);
nor NOR2 (N14019, N14005, N987);
nor NOR2 (N14020, N14017, N3556);
buf BUF1 (N14021, N14000);
nand NAND4 (N14022, N14014, N9472, N5893, N5922);
and AND2 (N14023, N14020, N6790);
xor XOR2 (N14024, N14023, N5882);
buf BUF1 (N14025, N14021);
or OR4 (N14026, N14016, N9123, N3230, N4370);
and AND3 (N14027, N14003, N8703, N10854);
nand NAND4 (N14028, N14027, N1761, N10380, N1472);
not NOT1 (N14029, N14026);
xor XOR2 (N14030, N14025, N8992);
nor NOR3 (N14031, N14018, N12431, N11661);
and AND2 (N14032, N14031, N11788);
nand NAND2 (N14033, N14029, N12131);
nand NAND3 (N14034, N14015, N11561, N7440);
xor XOR2 (N14035, N14011, N5784);
and AND3 (N14036, N14019, N7267, N10666);
and AND2 (N14037, N14033, N8324);
nor NOR3 (N14038, N14034, N9770, N10754);
and AND2 (N14039, N14028, N4408);
not NOT1 (N14040, N14024);
not NOT1 (N14041, N14039);
nand NAND4 (N14042, N14038, N10246, N9447, N10766);
xor XOR2 (N14043, N14037, N835);
nand NAND3 (N14044, N14035, N7204, N10382);
nor NOR2 (N14045, N14030, N6992);
or OR3 (N14046, N14032, N10173, N13373);
nor NOR3 (N14047, N14041, N12247, N10296);
xor XOR2 (N14048, N14047, N3393);
not NOT1 (N14049, N14048);
and AND4 (N14050, N14044, N7704, N13745, N5651);
buf BUF1 (N14051, N14046);
or OR3 (N14052, N14045, N9460, N4601);
not NOT1 (N14053, N14036);
not NOT1 (N14054, N14022);
buf BUF1 (N14055, N14050);
nor NOR3 (N14056, N14055, N11814, N3000);
and AND2 (N14057, N14043, N4715);
not NOT1 (N14058, N14049);
and AND4 (N14059, N14040, N6705, N10604, N8338);
xor XOR2 (N14060, N14010, N739);
buf BUF1 (N14061, N14059);
nand NAND3 (N14062, N14042, N5908, N11712);
buf BUF1 (N14063, N14060);
or OR3 (N14064, N14056, N271, N4228);
buf BUF1 (N14065, N14054);
buf BUF1 (N14066, N14061);
not NOT1 (N14067, N14053);
and AND2 (N14068, N14052, N455);
nand NAND3 (N14069, N14066, N3606, N8108);
and AND2 (N14070, N14064, N10559);
not NOT1 (N14071, N14062);
xor XOR2 (N14072, N14068, N9314);
xor XOR2 (N14073, N14071, N5456);
nand NAND2 (N14074, N14051, N1036);
nand NAND4 (N14075, N14058, N1736, N3674, N7074);
nand NAND3 (N14076, N14073, N3811, N11497);
and AND3 (N14077, N14067, N10855, N2900);
xor XOR2 (N14078, N14070, N8589);
xor XOR2 (N14079, N14074, N7377);
and AND4 (N14080, N14065, N1394, N3399, N425);
xor XOR2 (N14081, N14057, N286);
xor XOR2 (N14082, N14076, N5210);
xor XOR2 (N14083, N14072, N9565);
nor NOR4 (N14084, N14083, N835, N1799, N8446);
nor NOR3 (N14085, N14075, N9786, N6286);
nand NAND4 (N14086, N14078, N640, N12800, N8825);
xor XOR2 (N14087, N14084, N12450);
not NOT1 (N14088, N14069);
nand NAND4 (N14089, N14086, N9599, N11051, N11771);
xor XOR2 (N14090, N14087, N931);
xor XOR2 (N14091, N14082, N4549);
nand NAND4 (N14092, N14081, N4200, N8101, N3456);
buf BUF1 (N14093, N14080);
or OR4 (N14094, N14093, N7375, N1903, N3331);
xor XOR2 (N14095, N14094, N12894);
not NOT1 (N14096, N14063);
or OR4 (N14097, N14088, N9916, N9954, N2847);
nor NOR4 (N14098, N14085, N11606, N2914, N3578);
nor NOR3 (N14099, N14079, N2656, N5429);
xor XOR2 (N14100, N14095, N3259);
buf BUF1 (N14101, N14098);
or OR3 (N14102, N14099, N6601, N14025);
or OR3 (N14103, N14102, N8205, N5954);
buf BUF1 (N14104, N14097);
nand NAND2 (N14105, N14096, N3503);
buf BUF1 (N14106, N14105);
nor NOR3 (N14107, N14092, N1433, N3406);
buf BUF1 (N14108, N14101);
not NOT1 (N14109, N14106);
and AND3 (N14110, N14091, N6401, N12383);
buf BUF1 (N14111, N14109);
xor XOR2 (N14112, N14110, N10132);
nor NOR3 (N14113, N14103, N9056, N8843);
buf BUF1 (N14114, N14089);
xor XOR2 (N14115, N14100, N12251);
not NOT1 (N14116, N14113);
nand NAND2 (N14117, N14114, N2899);
nand NAND3 (N14118, N14115, N11134, N12293);
nand NAND4 (N14119, N14117, N13116, N11685, N12449);
not NOT1 (N14120, N14119);
xor XOR2 (N14121, N14118, N6691);
nor NOR2 (N14122, N14107, N1254);
nor NOR2 (N14123, N14116, N6594);
nand NAND3 (N14124, N14111, N11152, N14009);
or OR3 (N14125, N14122, N3169, N11145);
buf BUF1 (N14126, N14120);
nor NOR4 (N14127, N14121, N9873, N2568, N1193);
buf BUF1 (N14128, N14077);
nand NAND2 (N14129, N14126, N6493);
buf BUF1 (N14130, N14090);
and AND2 (N14131, N14108, N544);
xor XOR2 (N14132, N14104, N8310);
or OR3 (N14133, N14132, N12593, N4503);
buf BUF1 (N14134, N14128);
and AND3 (N14135, N14129, N6180, N1724);
buf BUF1 (N14136, N14134);
not NOT1 (N14137, N14135);
nand NAND4 (N14138, N14127, N14078, N6838, N11992);
buf BUF1 (N14139, N14137);
buf BUF1 (N14140, N14133);
xor XOR2 (N14141, N14131, N5995);
not NOT1 (N14142, N14130);
or OR3 (N14143, N14139, N515, N9156);
buf BUF1 (N14144, N14141);
or OR3 (N14145, N14123, N8770, N3344);
buf BUF1 (N14146, N14143);
buf BUF1 (N14147, N14145);
nand NAND3 (N14148, N14146, N7064, N10159);
or OR2 (N14149, N14140, N5779);
and AND2 (N14150, N14149, N1657);
nand NAND3 (N14151, N14147, N12128, N8909);
and AND4 (N14152, N14150, N1444, N5448, N13241);
nand NAND4 (N14153, N14151, N13752, N5633, N2606);
and AND3 (N14154, N14124, N7029, N13510);
not NOT1 (N14155, N14144);
buf BUF1 (N14156, N14136);
and AND2 (N14157, N14142, N1283);
not NOT1 (N14158, N14157);
not NOT1 (N14159, N14154);
or OR3 (N14160, N14155, N3069, N3884);
or OR3 (N14161, N14125, N12503, N3942);
buf BUF1 (N14162, N14152);
and AND3 (N14163, N14160, N10156, N12457);
buf BUF1 (N14164, N14161);
nor NOR4 (N14165, N14138, N4512, N12169, N13205);
and AND2 (N14166, N14163, N9161);
not NOT1 (N14167, N14162);
nor NOR3 (N14168, N14112, N710, N8840);
nor NOR2 (N14169, N14168, N12599);
nor NOR3 (N14170, N14164, N4851, N11611);
and AND2 (N14171, N14170, N10415);
buf BUF1 (N14172, N14167);
buf BUF1 (N14173, N14159);
or OR3 (N14174, N14171, N10318, N6780);
nor NOR3 (N14175, N14148, N239, N2928);
nand NAND4 (N14176, N14153, N7419, N1446, N14085);
nand NAND4 (N14177, N14173, N687, N6233, N2611);
not NOT1 (N14178, N14169);
or OR4 (N14179, N14176, N8612, N13656, N6575);
xor XOR2 (N14180, N14165, N2903);
xor XOR2 (N14181, N14158, N10559);
not NOT1 (N14182, N14166);
nor NOR3 (N14183, N14175, N479, N12840);
xor XOR2 (N14184, N14174, N3223);
and AND3 (N14185, N14183, N6400, N323);
nor NOR2 (N14186, N14172, N8250);
nand NAND4 (N14187, N14177, N5033, N11728, N9530);
or OR2 (N14188, N14179, N10625);
and AND2 (N14189, N14184, N2224);
and AND4 (N14190, N14182, N10647, N2953, N12717);
nor NOR3 (N14191, N14189, N10158, N5074);
and AND3 (N14192, N14191, N1627, N2638);
nand NAND4 (N14193, N14190, N12943, N953, N3616);
xor XOR2 (N14194, N14156, N8723);
nor NOR3 (N14195, N14185, N8243, N6471);
buf BUF1 (N14196, N14193);
nor NOR4 (N14197, N14178, N6961, N7662, N7531);
nor NOR3 (N14198, N14186, N3676, N10691);
nor NOR3 (N14199, N14180, N5334, N1661);
not NOT1 (N14200, N14188);
buf BUF1 (N14201, N14199);
nand NAND4 (N14202, N14181, N8758, N10580, N6855);
or OR3 (N14203, N14195, N8115, N2526);
or OR4 (N14204, N14192, N14093, N1143, N11372);
not NOT1 (N14205, N14204);
or OR3 (N14206, N14194, N4397, N3901);
buf BUF1 (N14207, N14205);
buf BUF1 (N14208, N14198);
xor XOR2 (N14209, N14207, N6241);
and AND4 (N14210, N14200, N12725, N725, N8029);
nor NOR3 (N14211, N14206, N9553, N5018);
nor NOR3 (N14212, N14187, N7024, N4877);
buf BUF1 (N14213, N14211);
nand NAND4 (N14214, N14201, N9082, N88, N9110);
or OR2 (N14215, N14202, N9072);
xor XOR2 (N14216, N14209, N10678);
buf BUF1 (N14217, N14196);
and AND2 (N14218, N14212, N6315);
not NOT1 (N14219, N14215);
or OR2 (N14220, N14219, N868);
and AND2 (N14221, N14214, N11350);
and AND2 (N14222, N14220, N8965);
nor NOR4 (N14223, N14197, N3991, N7826, N4924);
nor NOR3 (N14224, N14221, N4453, N3258);
and AND3 (N14225, N14217, N13269, N117);
xor XOR2 (N14226, N14225, N6109);
nand NAND2 (N14227, N14218, N1306);
xor XOR2 (N14228, N14203, N7364);
or OR4 (N14229, N14222, N8833, N8322, N11570);
not NOT1 (N14230, N14213);
buf BUF1 (N14231, N14226);
not NOT1 (N14232, N14229);
or OR3 (N14233, N14230, N5202, N10170);
and AND2 (N14234, N14210, N347);
not NOT1 (N14235, N14233);
buf BUF1 (N14236, N14228);
and AND2 (N14237, N14234, N4369);
nor NOR4 (N14238, N14231, N7200, N12274, N5451);
xor XOR2 (N14239, N14208, N1493);
and AND3 (N14240, N14227, N5391, N5546);
and AND2 (N14241, N14216, N10207);
xor XOR2 (N14242, N14235, N11536);
nor NOR4 (N14243, N14224, N9835, N8049, N8944);
nor NOR3 (N14244, N14223, N9829, N9282);
and AND2 (N14245, N14244, N4440);
not NOT1 (N14246, N14245);
buf BUF1 (N14247, N14237);
nor NOR2 (N14248, N14243, N6889);
nand NAND2 (N14249, N14238, N5782);
and AND3 (N14250, N14232, N1926, N6636);
not NOT1 (N14251, N14239);
xor XOR2 (N14252, N14249, N4135);
nand NAND3 (N14253, N14240, N13842, N9030);
and AND2 (N14254, N14236, N12727);
and AND3 (N14255, N14252, N13757, N11684);
nand NAND4 (N14256, N14246, N971, N2865, N11536);
not NOT1 (N14257, N14241);
and AND3 (N14258, N14251, N1955, N14127);
or OR3 (N14259, N14255, N3925, N8846);
buf BUF1 (N14260, N14247);
nor NOR2 (N14261, N14242, N8394);
xor XOR2 (N14262, N14260, N3769);
or OR3 (N14263, N14250, N7360, N2805);
not NOT1 (N14264, N14261);
and AND2 (N14265, N14254, N10974);
xor XOR2 (N14266, N14256, N9067);
xor XOR2 (N14267, N14248, N5275);
not NOT1 (N14268, N14263);
not NOT1 (N14269, N14253);
buf BUF1 (N14270, N14265);
nor NOR3 (N14271, N14264, N4374, N13247);
not NOT1 (N14272, N14269);
buf BUF1 (N14273, N14266);
or OR2 (N14274, N14270, N1191);
nand NAND2 (N14275, N14272, N799);
buf BUF1 (N14276, N14275);
or OR3 (N14277, N14271, N14167, N831);
nor NOR4 (N14278, N14268, N6022, N867, N10211);
and AND4 (N14279, N14267, N4191, N7956, N11385);
and AND4 (N14280, N14277, N5818, N7799, N10777);
and AND4 (N14281, N14257, N9254, N8554, N2313);
not NOT1 (N14282, N14281);
nand NAND4 (N14283, N14278, N9718, N13207, N2914);
buf BUF1 (N14284, N14259);
xor XOR2 (N14285, N14258, N4485);
and AND2 (N14286, N14285, N8765);
xor XOR2 (N14287, N14276, N4791);
xor XOR2 (N14288, N14286, N4124);
not NOT1 (N14289, N14284);
not NOT1 (N14290, N14274);
and AND4 (N14291, N14288, N4919, N9802, N2427);
or OR4 (N14292, N14289, N6395, N13492, N6789);
nand NAND2 (N14293, N14282, N5349);
or OR2 (N14294, N14292, N3238);
xor XOR2 (N14295, N14294, N3497);
not NOT1 (N14296, N14283);
buf BUF1 (N14297, N14287);
nand NAND2 (N14298, N14273, N8203);
nand NAND3 (N14299, N14279, N801, N5727);
not NOT1 (N14300, N14298);
xor XOR2 (N14301, N14293, N4397);
buf BUF1 (N14302, N14291);
buf BUF1 (N14303, N14295);
xor XOR2 (N14304, N14302, N7193);
or OR3 (N14305, N14300, N13153, N9300);
not NOT1 (N14306, N14305);
buf BUF1 (N14307, N14304);
xor XOR2 (N14308, N14296, N8016);
or OR3 (N14309, N14307, N9646, N3736);
or OR3 (N14310, N14301, N12178, N12557);
xor XOR2 (N14311, N14303, N4698);
buf BUF1 (N14312, N14311);
nand NAND2 (N14313, N14290, N10492);
nor NOR2 (N14314, N14312, N899);
nor NOR2 (N14315, N14297, N3590);
nor NOR2 (N14316, N14308, N673);
not NOT1 (N14317, N14315);
nor NOR3 (N14318, N14317, N5168, N8397);
or OR4 (N14319, N14309, N6097, N3196, N8800);
not NOT1 (N14320, N14280);
and AND4 (N14321, N14299, N6712, N8744, N9564);
nor NOR4 (N14322, N14316, N1617, N6942, N3262);
nand NAND4 (N14323, N14322, N712, N12762, N3266);
and AND3 (N14324, N14323, N14105, N10627);
buf BUF1 (N14325, N14310);
and AND2 (N14326, N14319, N8632);
nor NOR4 (N14327, N14321, N4013, N12723, N2774);
nand NAND4 (N14328, N14325, N8328, N9882, N2213);
nand NAND4 (N14329, N14320, N10955, N1342, N7306);
buf BUF1 (N14330, N14306);
xor XOR2 (N14331, N14318, N699);
buf BUF1 (N14332, N14328);
and AND3 (N14333, N14314, N2066, N2744);
not NOT1 (N14334, N14326);
buf BUF1 (N14335, N14332);
or OR3 (N14336, N14324, N4864, N559);
and AND2 (N14337, N14335, N2622);
nand NAND3 (N14338, N14330, N4896, N7679);
xor XOR2 (N14339, N14337, N3029);
xor XOR2 (N14340, N14336, N1855);
buf BUF1 (N14341, N14329);
nand NAND2 (N14342, N14333, N11414);
or OR4 (N14343, N14338, N5905, N5065, N7452);
or OR4 (N14344, N14339, N7868, N10570, N3535);
buf BUF1 (N14345, N14344);
buf BUF1 (N14346, N14345);
or OR3 (N14347, N14331, N11870, N14018);
and AND4 (N14348, N14346, N11669, N7943, N6205);
not NOT1 (N14349, N14347);
xor XOR2 (N14350, N14349, N3923);
buf BUF1 (N14351, N14327);
not NOT1 (N14352, N14334);
and AND2 (N14353, N14342, N9430);
buf BUF1 (N14354, N14341);
buf BUF1 (N14355, N14348);
not NOT1 (N14356, N14340);
nor NOR2 (N14357, N14353, N10239);
or OR2 (N14358, N14356, N5815);
nand NAND4 (N14359, N14357, N10474, N11606, N4867);
and AND3 (N14360, N14354, N7459, N9369);
xor XOR2 (N14361, N14355, N7446);
buf BUF1 (N14362, N14262);
xor XOR2 (N14363, N14352, N11343);
xor XOR2 (N14364, N14362, N14291);
buf BUF1 (N14365, N14363);
not NOT1 (N14366, N14365);
not NOT1 (N14367, N14361);
not NOT1 (N14368, N14367);
xor XOR2 (N14369, N14360, N5042);
and AND4 (N14370, N14350, N2632, N4702, N14226);
buf BUF1 (N14371, N14359);
or OR3 (N14372, N14351, N11823, N13289);
nor NOR4 (N14373, N14313, N9488, N11047, N1783);
nand NAND2 (N14374, N14358, N3233);
buf BUF1 (N14375, N14368);
or OR2 (N14376, N14369, N2265);
xor XOR2 (N14377, N14370, N10516);
buf BUF1 (N14378, N14373);
and AND2 (N14379, N14377, N10789);
nor NOR4 (N14380, N14376, N13069, N13678, N7761);
or OR3 (N14381, N14378, N8345, N3132);
nand NAND2 (N14382, N14372, N8907);
not NOT1 (N14383, N14364);
not NOT1 (N14384, N14375);
buf BUF1 (N14385, N14366);
xor XOR2 (N14386, N14374, N12443);
and AND3 (N14387, N14343, N10291, N12076);
xor XOR2 (N14388, N14386, N3650);
nand NAND2 (N14389, N14381, N11508);
and AND2 (N14390, N14379, N10701);
nand NAND4 (N14391, N14371, N5947, N13316, N6603);
xor XOR2 (N14392, N14387, N1503);
and AND4 (N14393, N14380, N13645, N4271, N2952);
buf BUF1 (N14394, N14388);
and AND2 (N14395, N14393, N1935);
not NOT1 (N14396, N14382);
xor XOR2 (N14397, N14385, N2772);
nor NOR2 (N14398, N14383, N9563);
nand NAND4 (N14399, N14390, N1182, N6856, N7420);
xor XOR2 (N14400, N14391, N12850);
buf BUF1 (N14401, N14389);
buf BUF1 (N14402, N14401);
buf BUF1 (N14403, N14384);
and AND4 (N14404, N14403, N161, N3678, N5491);
nor NOR2 (N14405, N14394, N14001);
xor XOR2 (N14406, N14405, N2140);
nand NAND2 (N14407, N14404, N8868);
nand NAND4 (N14408, N14406, N2543, N10168, N11339);
and AND3 (N14409, N14398, N8260, N8873);
not NOT1 (N14410, N14392);
buf BUF1 (N14411, N14402);
buf BUF1 (N14412, N14409);
or OR2 (N14413, N14408, N11766);
buf BUF1 (N14414, N14407);
and AND2 (N14415, N14397, N9051);
nand NAND3 (N14416, N14415, N6714, N7410);
nand NAND3 (N14417, N14413, N15, N4862);
not NOT1 (N14418, N14412);
nor NOR4 (N14419, N14417, N6942, N1380, N10028);
not NOT1 (N14420, N14416);
or OR3 (N14421, N14419, N5904, N10691);
nor NOR3 (N14422, N14420, N7709, N1111);
not NOT1 (N14423, N14414);
nand NAND3 (N14424, N14400, N10525, N6444);
buf BUF1 (N14425, N14423);
nand NAND2 (N14426, N14425, N10810);
and AND3 (N14427, N14421, N12841, N14405);
xor XOR2 (N14428, N14427, N8843);
buf BUF1 (N14429, N14410);
xor XOR2 (N14430, N14411, N14171);
nor NOR4 (N14431, N14428, N6492, N1349, N10704);
buf BUF1 (N14432, N14424);
not NOT1 (N14433, N14396);
nor NOR4 (N14434, N14432, N6199, N9101, N8177);
nand NAND3 (N14435, N14422, N5474, N81);
nor NOR4 (N14436, N14431, N9540, N2379, N6595);
buf BUF1 (N14437, N14434);
nor NOR2 (N14438, N14399, N49);
nand NAND4 (N14439, N14418, N2594, N12624, N5196);
and AND2 (N14440, N14433, N5324);
or OR4 (N14441, N14395, N13169, N9549, N4295);
buf BUF1 (N14442, N14437);
buf BUF1 (N14443, N14429);
and AND3 (N14444, N14435, N12926, N13414);
nor NOR4 (N14445, N14443, N12564, N4561, N6223);
xor XOR2 (N14446, N14426, N2631);
xor XOR2 (N14447, N14444, N13007);
and AND2 (N14448, N14445, N8976);
or OR2 (N14449, N14442, N12608);
not NOT1 (N14450, N14430);
nor NOR2 (N14451, N14450, N9879);
not NOT1 (N14452, N14449);
or OR3 (N14453, N14452, N12903, N7761);
or OR4 (N14454, N14446, N2071, N11381, N14297);
and AND4 (N14455, N14451, N7440, N12562, N11169);
and AND3 (N14456, N14436, N9704, N11956);
xor XOR2 (N14457, N14456, N7021);
buf BUF1 (N14458, N14447);
and AND2 (N14459, N14454, N1126);
or OR4 (N14460, N14453, N12579, N7659, N4594);
not NOT1 (N14461, N14448);
or OR4 (N14462, N14438, N12281, N6016, N3501);
and AND3 (N14463, N14440, N9310, N4786);
and AND2 (N14464, N14462, N8090);
or OR2 (N14465, N14461, N7244);
nor NOR4 (N14466, N14441, N1322, N9233, N10691);
or OR2 (N14467, N14465, N13719);
not NOT1 (N14468, N14464);
xor XOR2 (N14469, N14455, N258);
nand NAND2 (N14470, N14467, N10848);
nor NOR2 (N14471, N14460, N10735);
or OR3 (N14472, N14470, N5591, N4934);
nand NAND3 (N14473, N14468, N231, N3130);
xor XOR2 (N14474, N14472, N9561);
xor XOR2 (N14475, N14459, N13109);
not NOT1 (N14476, N14466);
and AND3 (N14477, N14475, N7895, N5677);
not NOT1 (N14478, N14439);
nor NOR4 (N14479, N14476, N3055, N7626, N664);
not NOT1 (N14480, N14473);
not NOT1 (N14481, N14471);
buf BUF1 (N14482, N14480);
nor NOR2 (N14483, N14457, N8868);
not NOT1 (N14484, N14481);
nand NAND2 (N14485, N14484, N2000);
not NOT1 (N14486, N14482);
or OR2 (N14487, N14469, N486);
buf BUF1 (N14488, N14483);
and AND2 (N14489, N14488, N10999);
nand NAND3 (N14490, N14485, N7366, N4040);
or OR4 (N14491, N14489, N424, N6, N10386);
xor XOR2 (N14492, N14487, N4400);
or OR3 (N14493, N14458, N5320, N6659);
or OR4 (N14494, N14486, N12148, N6683, N10396);
nor NOR4 (N14495, N14494, N6014, N12997, N3996);
buf BUF1 (N14496, N14490);
or OR3 (N14497, N14479, N12072, N7981);
not NOT1 (N14498, N14478);
or OR4 (N14499, N14463, N5700, N9980, N8451);
buf BUF1 (N14500, N14493);
nor NOR3 (N14501, N14491, N9675, N2366);
and AND3 (N14502, N14497, N46, N12308);
not NOT1 (N14503, N14496);
not NOT1 (N14504, N14500);
xor XOR2 (N14505, N14502, N2608);
and AND2 (N14506, N14505, N11904);
not NOT1 (N14507, N14477);
xor XOR2 (N14508, N14501, N2009);
buf BUF1 (N14509, N14492);
xor XOR2 (N14510, N14503, N13575);
xor XOR2 (N14511, N14508, N804);
xor XOR2 (N14512, N14504, N8994);
xor XOR2 (N14513, N14507, N1227);
and AND4 (N14514, N14509, N14359, N5336, N1252);
and AND4 (N14515, N14506, N142, N67, N5059);
nand NAND2 (N14516, N14514, N2315);
not NOT1 (N14517, N14516);
xor XOR2 (N14518, N14510, N6319);
buf BUF1 (N14519, N14495);
buf BUF1 (N14520, N14511);
not NOT1 (N14521, N14519);
buf BUF1 (N14522, N14521);
buf BUF1 (N14523, N14522);
nor NOR4 (N14524, N14498, N4930, N8949, N5577);
xor XOR2 (N14525, N14524, N4100);
or OR2 (N14526, N14525, N5414);
nor NOR2 (N14527, N14518, N1741);
or OR2 (N14528, N14523, N8284);
xor XOR2 (N14529, N14513, N7406);
nand NAND3 (N14530, N14517, N4625, N2973);
buf BUF1 (N14531, N14530);
xor XOR2 (N14532, N14527, N464);
or OR2 (N14533, N14512, N9254);
and AND2 (N14534, N14520, N11237);
xor XOR2 (N14535, N14529, N8850);
nand NAND2 (N14536, N14531, N12371);
not NOT1 (N14537, N14526);
not NOT1 (N14538, N14528);
and AND3 (N14539, N14534, N860, N9091);
or OR3 (N14540, N14533, N14369, N6293);
buf BUF1 (N14541, N14540);
or OR3 (N14542, N14538, N11551, N3810);
not NOT1 (N14543, N14532);
or OR4 (N14544, N14542, N695, N1712, N3740);
nor NOR4 (N14545, N14499, N5552, N13301, N3661);
or OR4 (N14546, N14535, N2106, N6918, N12278);
nor NOR2 (N14547, N14545, N8217);
xor XOR2 (N14548, N14543, N5076);
buf BUF1 (N14549, N14537);
not NOT1 (N14550, N14544);
xor XOR2 (N14551, N14539, N2438);
nor NOR3 (N14552, N14515, N5643, N38);
and AND3 (N14553, N14474, N1459, N13844);
xor XOR2 (N14554, N14546, N14207);
or OR2 (N14555, N14552, N9946);
xor XOR2 (N14556, N14555, N325);
nor NOR3 (N14557, N14541, N11971, N13159);
not NOT1 (N14558, N14551);
buf BUF1 (N14559, N14549);
or OR3 (N14560, N14547, N5632, N6139);
nor NOR4 (N14561, N14553, N3766, N8027, N7204);
nand NAND2 (N14562, N14557, N8510);
or OR3 (N14563, N14558, N1949, N329);
and AND3 (N14564, N14563, N12374, N9590);
nor NOR2 (N14565, N14561, N9412);
buf BUF1 (N14566, N14564);
not NOT1 (N14567, N14556);
nand NAND3 (N14568, N14554, N3347, N7284);
and AND3 (N14569, N14565, N11685, N9599);
not NOT1 (N14570, N14536);
nand NAND3 (N14571, N14569, N3887, N10854);
nand NAND3 (N14572, N14560, N7950, N3926);
nor NOR2 (N14573, N14567, N7805);
not NOT1 (N14574, N14568);
buf BUF1 (N14575, N14570);
not NOT1 (N14576, N14575);
nand NAND2 (N14577, N14559, N11093);
nor NOR3 (N14578, N14566, N7172, N3894);
nor NOR4 (N14579, N14573, N3040, N1133, N635);
nand NAND4 (N14580, N14576, N13166, N8017, N12883);
or OR4 (N14581, N14579, N8578, N6924, N8067);
or OR3 (N14582, N14581, N1119, N846);
nand NAND2 (N14583, N14550, N7927);
xor XOR2 (N14584, N14582, N11854);
xor XOR2 (N14585, N14562, N4820);
nand NAND2 (N14586, N14585, N5549);
nor NOR4 (N14587, N14572, N4200, N7946, N7259);
and AND2 (N14588, N14574, N7978);
buf BUF1 (N14589, N14577);
xor XOR2 (N14590, N14588, N12322);
or OR4 (N14591, N14586, N13850, N13332, N14485);
or OR3 (N14592, N14578, N9774, N10887);
xor XOR2 (N14593, N14548, N6552);
xor XOR2 (N14594, N14571, N6346);
or OR4 (N14595, N14583, N2355, N363, N6799);
nor NOR3 (N14596, N14595, N3793, N12030);
or OR4 (N14597, N14584, N7225, N12684, N13165);
not NOT1 (N14598, N14589);
xor XOR2 (N14599, N14580, N12837);
nand NAND3 (N14600, N14599, N7722, N9072);
not NOT1 (N14601, N14592);
or OR3 (N14602, N14601, N4461, N6484);
nand NAND2 (N14603, N14590, N6134);
not NOT1 (N14604, N14597);
buf BUF1 (N14605, N14591);
or OR2 (N14606, N14593, N2466);
or OR2 (N14607, N14596, N9223);
buf BUF1 (N14608, N14600);
and AND4 (N14609, N14605, N7321, N10558, N13948);
not NOT1 (N14610, N14594);
nand NAND3 (N14611, N14604, N3691, N8382);
nor NOR3 (N14612, N14609, N6329, N5926);
and AND3 (N14613, N14608, N10937, N7348);
buf BUF1 (N14614, N14607);
or OR2 (N14615, N14606, N2488);
buf BUF1 (N14616, N14615);
not NOT1 (N14617, N14587);
nand NAND4 (N14618, N14617, N6803, N47, N12220);
nor NOR4 (N14619, N14612, N1670, N3120, N304);
nor NOR3 (N14620, N14616, N14179, N8331);
xor XOR2 (N14621, N14603, N3974);
not NOT1 (N14622, N14614);
not NOT1 (N14623, N14613);
or OR2 (N14624, N14618, N13217);
nor NOR3 (N14625, N14620, N1843, N8770);
nand NAND2 (N14626, N14598, N14232);
nor NOR2 (N14627, N14611, N1761);
or OR2 (N14628, N14627, N12137);
or OR3 (N14629, N14602, N10743, N6530);
nor NOR3 (N14630, N14623, N1825, N13410);
buf BUF1 (N14631, N14610);
or OR2 (N14632, N14629, N12483);
or OR2 (N14633, N14621, N13627);
and AND4 (N14634, N14626, N2281, N11595, N11178);
or OR4 (N14635, N14622, N12566, N13460, N1751);
not NOT1 (N14636, N14628);
nor NOR3 (N14637, N14619, N7226, N1737);
xor XOR2 (N14638, N14636, N9693);
xor XOR2 (N14639, N14630, N622);
nand NAND4 (N14640, N14625, N12607, N3267, N2635);
buf BUF1 (N14641, N14639);
nand NAND4 (N14642, N14637, N10212, N9807, N5049);
or OR3 (N14643, N14642, N9844, N5479);
nand NAND3 (N14644, N14638, N12518, N11682);
xor XOR2 (N14645, N14632, N5551);
xor XOR2 (N14646, N14635, N3171);
and AND2 (N14647, N14643, N8205);
or OR2 (N14648, N14634, N6213);
nor NOR4 (N14649, N14631, N9496, N5057, N3447);
xor XOR2 (N14650, N14640, N9018);
not NOT1 (N14651, N14644);
xor XOR2 (N14652, N14649, N12334);
not NOT1 (N14653, N14624);
buf BUF1 (N14654, N14648);
or OR2 (N14655, N14650, N2749);
or OR3 (N14656, N14641, N13625, N402);
or OR3 (N14657, N14651, N4553, N9615);
nand NAND4 (N14658, N14647, N14071, N5075, N6664);
not NOT1 (N14659, N14646);
buf BUF1 (N14660, N14659);
or OR4 (N14661, N14657, N1645, N10044, N6319);
not NOT1 (N14662, N14661);
or OR4 (N14663, N14653, N1208, N3415, N4665);
xor XOR2 (N14664, N14655, N11553);
and AND2 (N14665, N14664, N14182);
not NOT1 (N14666, N14633);
not NOT1 (N14667, N14660);
buf BUF1 (N14668, N14662);
xor XOR2 (N14669, N14652, N2522);
buf BUF1 (N14670, N14663);
and AND2 (N14671, N14668, N2450);
or OR4 (N14672, N14656, N540, N6911, N12983);
and AND2 (N14673, N14669, N8506);
not NOT1 (N14674, N14665);
not NOT1 (N14675, N14658);
and AND3 (N14676, N14671, N516, N13795);
xor XOR2 (N14677, N14675, N4606);
and AND4 (N14678, N14666, N9553, N2388, N10799);
nor NOR2 (N14679, N14678, N5184);
and AND3 (N14680, N14676, N10047, N8338);
or OR3 (N14681, N14672, N2568, N3742);
or OR2 (N14682, N14674, N2004);
not NOT1 (N14683, N14673);
xor XOR2 (N14684, N14679, N271);
or OR3 (N14685, N14670, N7024, N5154);
buf BUF1 (N14686, N14680);
xor XOR2 (N14687, N14682, N2897);
not NOT1 (N14688, N14681);
not NOT1 (N14689, N14667);
nand NAND4 (N14690, N14684, N12587, N14385, N13820);
nand NAND4 (N14691, N14687, N11433, N2738, N11173);
not NOT1 (N14692, N14689);
nor NOR2 (N14693, N14691, N1588);
buf BUF1 (N14694, N14683);
nor NOR3 (N14695, N14688, N4679, N1188);
or OR4 (N14696, N14692, N9448, N5024, N6415);
or OR2 (N14697, N14694, N14426);
nand NAND3 (N14698, N14686, N10080, N9131);
xor XOR2 (N14699, N14690, N6196);
or OR2 (N14700, N14696, N12895);
not NOT1 (N14701, N14699);
nor NOR4 (N14702, N14645, N9509, N12532, N6922);
or OR2 (N14703, N14701, N7552);
and AND2 (N14704, N14702, N13389);
not NOT1 (N14705, N14698);
and AND3 (N14706, N14693, N4979, N9513);
buf BUF1 (N14707, N14703);
buf BUF1 (N14708, N14677);
not NOT1 (N14709, N14654);
and AND2 (N14710, N14695, N6565);
buf BUF1 (N14711, N14705);
xor XOR2 (N14712, N14704, N11375);
nand NAND2 (N14713, N14708, N11870);
or OR2 (N14714, N14700, N5313);
nor NOR2 (N14715, N14697, N7907);
and AND3 (N14716, N14715, N836, N7200);
or OR4 (N14717, N14707, N5561, N2302, N9190);
and AND4 (N14718, N14710, N8352, N14300, N7799);
and AND2 (N14719, N14709, N1267);
xor XOR2 (N14720, N14714, N10706);
nand NAND3 (N14721, N14712, N350, N7176);
or OR4 (N14722, N14720, N3182, N11645, N14251);
and AND3 (N14723, N14716, N11868, N2746);
buf BUF1 (N14724, N14722);
buf BUF1 (N14725, N14711);
and AND4 (N14726, N14685, N254, N4770, N8973);
not NOT1 (N14727, N14706);
nor NOR2 (N14728, N14727, N8061);
buf BUF1 (N14729, N14726);
or OR3 (N14730, N14728, N11834, N11812);
xor XOR2 (N14731, N14721, N5379);
or OR2 (N14732, N14718, N5822);
buf BUF1 (N14733, N14729);
not NOT1 (N14734, N14725);
nand NAND4 (N14735, N14731, N12039, N3361, N12541);
nand NAND2 (N14736, N14713, N11663);
and AND4 (N14737, N14719, N7810, N11609, N5218);
nor NOR4 (N14738, N14733, N6256, N6470, N9925);
nand NAND4 (N14739, N14724, N5560, N11375, N5177);
nor NOR4 (N14740, N14732, N7036, N10500, N3497);
not NOT1 (N14741, N14736);
or OR3 (N14742, N14730, N189, N14631);
not NOT1 (N14743, N14741);
or OR4 (N14744, N14743, N5113, N7329, N3600);
not NOT1 (N14745, N14739);
not NOT1 (N14746, N14737);
buf BUF1 (N14747, N14744);
nor NOR4 (N14748, N14742, N10252, N2739, N1067);
or OR2 (N14749, N14747, N3900);
nor NOR2 (N14750, N14738, N5372);
not NOT1 (N14751, N14745);
buf BUF1 (N14752, N14723);
and AND2 (N14753, N14740, N9847);
xor XOR2 (N14754, N14749, N2973);
not NOT1 (N14755, N14717);
and AND4 (N14756, N14734, N2812, N13323, N2583);
not NOT1 (N14757, N14748);
xor XOR2 (N14758, N14746, N11961);
nand NAND3 (N14759, N14735, N3308, N1442);
or OR4 (N14760, N14752, N2199, N4724, N10033);
buf BUF1 (N14761, N14755);
nand NAND2 (N14762, N14760, N5890);
nand NAND2 (N14763, N14761, N11129);
xor XOR2 (N14764, N14763, N12871);
buf BUF1 (N14765, N14754);
and AND4 (N14766, N14756, N1831, N13425, N3364);
or OR3 (N14767, N14758, N2675, N890);
nor NOR2 (N14768, N14766, N8801);
nand NAND4 (N14769, N14757, N14262, N7718, N11338);
buf BUF1 (N14770, N14762);
not NOT1 (N14771, N14759);
xor XOR2 (N14772, N14753, N11520);
or OR4 (N14773, N14765, N6488, N6992, N8665);
and AND3 (N14774, N14769, N11348, N6894);
nor NOR3 (N14775, N14767, N1326, N572);
xor XOR2 (N14776, N14771, N11197);
nor NOR2 (N14777, N14776, N14710);
buf BUF1 (N14778, N14764);
nand NAND3 (N14779, N14772, N12725, N8588);
and AND3 (N14780, N14773, N13557, N3485);
and AND3 (N14781, N14751, N4043, N9506);
not NOT1 (N14782, N14781);
or OR3 (N14783, N14768, N821, N8290);
buf BUF1 (N14784, N14774);
and AND2 (N14785, N14770, N11247);
nor NOR2 (N14786, N14785, N4189);
or OR3 (N14787, N14783, N9836, N6026);
and AND2 (N14788, N14750, N4099);
xor XOR2 (N14789, N14786, N6514);
nor NOR2 (N14790, N14778, N4401);
and AND3 (N14791, N14784, N7257, N6783);
xor XOR2 (N14792, N14780, N7404);
and AND2 (N14793, N14782, N7786);
or OR4 (N14794, N14779, N3686, N3370, N9827);
nand NAND4 (N14795, N14794, N8996, N11787, N6613);
nand NAND3 (N14796, N14777, N6227, N7871);
buf BUF1 (N14797, N14792);
or OR3 (N14798, N14788, N7608, N13769);
buf BUF1 (N14799, N14798);
xor XOR2 (N14800, N14787, N6701);
nor NOR2 (N14801, N14796, N3225);
and AND4 (N14802, N14800, N2775, N11259, N2504);
xor XOR2 (N14803, N14793, N8425);
nor NOR3 (N14804, N14801, N14127, N13336);
and AND3 (N14805, N14804, N7296, N3005);
nor NOR4 (N14806, N14795, N2299, N13193, N7584);
buf BUF1 (N14807, N14791);
buf BUF1 (N14808, N14775);
xor XOR2 (N14809, N14797, N3547);
and AND3 (N14810, N14809, N12011, N2436);
nand NAND2 (N14811, N14808, N1849);
not NOT1 (N14812, N14805);
xor XOR2 (N14813, N14803, N3519);
and AND2 (N14814, N14790, N3357);
and AND3 (N14815, N14811, N2348, N12452);
xor XOR2 (N14816, N14812, N10421);
xor XOR2 (N14817, N14789, N3002);
and AND3 (N14818, N14802, N9945, N10817);
and AND3 (N14819, N14816, N9294, N7306);
xor XOR2 (N14820, N14817, N5997);
nor NOR4 (N14821, N14820, N10578, N12481, N12289);
nand NAND3 (N14822, N14799, N9027, N8077);
and AND3 (N14823, N14813, N4883, N3873);
buf BUF1 (N14824, N14823);
xor XOR2 (N14825, N14810, N2172);
or OR4 (N14826, N14819, N11760, N3357, N3151);
xor XOR2 (N14827, N14821, N145);
xor XOR2 (N14828, N14826, N1354);
nand NAND2 (N14829, N14806, N8764);
and AND2 (N14830, N14818, N10035);
nand NAND3 (N14831, N14829, N3409, N11822);
xor XOR2 (N14832, N14815, N13506);
xor XOR2 (N14833, N14824, N8430);
or OR4 (N14834, N14827, N4121, N11217, N7388);
or OR3 (N14835, N14814, N13718, N11209);
nand NAND4 (N14836, N14807, N7983, N457, N5251);
not NOT1 (N14837, N14834);
xor XOR2 (N14838, N14828, N5420);
buf BUF1 (N14839, N14832);
and AND4 (N14840, N14822, N12537, N3948, N4029);
and AND4 (N14841, N14839, N10737, N12844, N10290);
nand NAND3 (N14842, N14837, N11079, N3312);
xor XOR2 (N14843, N14842, N4878);
buf BUF1 (N14844, N14843);
not NOT1 (N14845, N14840);
not NOT1 (N14846, N14841);
nand NAND2 (N14847, N14845, N5853);
not NOT1 (N14848, N14844);
not NOT1 (N14849, N14847);
and AND3 (N14850, N14831, N3306, N14251);
nor NOR2 (N14851, N14833, N7661);
or OR4 (N14852, N14848, N6578, N5515, N4423);
xor XOR2 (N14853, N14838, N13175);
nor NOR3 (N14854, N14836, N5518, N14762);
nor NOR3 (N14855, N14852, N3278, N9298);
xor XOR2 (N14856, N14849, N4542);
xor XOR2 (N14857, N14846, N11067);
nor NOR3 (N14858, N14835, N12605, N5243);
and AND2 (N14859, N14851, N11238);
not NOT1 (N14860, N14859);
buf BUF1 (N14861, N14850);
not NOT1 (N14862, N14825);
nor NOR4 (N14863, N14857, N121, N3978, N11911);
nand NAND2 (N14864, N14860, N6898);
and AND4 (N14865, N14863, N12650, N776, N11438);
nand NAND4 (N14866, N14862, N3002, N14324, N525);
xor XOR2 (N14867, N14856, N7488);
xor XOR2 (N14868, N14864, N7161);
xor XOR2 (N14869, N14866, N11985);
nand NAND3 (N14870, N14858, N4105, N3724);
xor XOR2 (N14871, N14868, N8540);
not NOT1 (N14872, N14853);
buf BUF1 (N14873, N14867);
nor NOR4 (N14874, N14872, N2789, N9410, N3769);
xor XOR2 (N14875, N14855, N3516);
not NOT1 (N14876, N14874);
nand NAND3 (N14877, N14870, N11864, N13808);
xor XOR2 (N14878, N14875, N13517);
nand NAND4 (N14879, N14865, N2824, N6731, N11213);
not NOT1 (N14880, N14876);
not NOT1 (N14881, N14877);
nand NAND2 (N14882, N14871, N6032);
buf BUF1 (N14883, N14873);
nor NOR2 (N14884, N14882, N9657);
and AND4 (N14885, N14878, N11174, N508, N7704);
not NOT1 (N14886, N14879);
buf BUF1 (N14887, N14861);
or OR3 (N14888, N14887, N6171, N11220);
and AND2 (N14889, N14886, N3439);
xor XOR2 (N14890, N14884, N5357);
or OR2 (N14891, N14830, N12240);
buf BUF1 (N14892, N14880);
buf BUF1 (N14893, N14890);
or OR3 (N14894, N14892, N2603, N3380);
or OR3 (N14895, N14893, N2949, N7070);
nand NAND3 (N14896, N14891, N2315, N14149);
or OR3 (N14897, N14885, N3733, N10629);
and AND3 (N14898, N14896, N7805, N4738);
not NOT1 (N14899, N14895);
xor XOR2 (N14900, N14889, N6543);
nand NAND4 (N14901, N14894, N14682, N12856, N9113);
nand NAND3 (N14902, N14901, N664, N337);
and AND3 (N14903, N14869, N14523, N4000);
nand NAND2 (N14904, N14854, N8576);
xor XOR2 (N14905, N14898, N12953);
nor NOR2 (N14906, N14904, N13631);
buf BUF1 (N14907, N14903);
not NOT1 (N14908, N14902);
xor XOR2 (N14909, N14899, N3078);
or OR2 (N14910, N14908, N8528);
buf BUF1 (N14911, N14910);
buf BUF1 (N14912, N14881);
buf BUF1 (N14913, N14906);
xor XOR2 (N14914, N14913, N3926);
not NOT1 (N14915, N14883);
buf BUF1 (N14916, N14911);
not NOT1 (N14917, N14905);
and AND4 (N14918, N14897, N11870, N2647, N12007);
buf BUF1 (N14919, N14917);
nand NAND2 (N14920, N14915, N8696);
nor NOR2 (N14921, N14916, N8631);
buf BUF1 (N14922, N14914);
or OR3 (N14923, N14918, N3067, N957);
nand NAND2 (N14924, N14921, N13389);
and AND2 (N14925, N14924, N1329);
nand NAND3 (N14926, N14909, N3413, N10926);
buf BUF1 (N14927, N14900);
nor NOR3 (N14928, N14927, N4851, N816);
and AND3 (N14929, N14919, N3663, N6728);
nand NAND4 (N14930, N14888, N6470, N6164, N10898);
nor NOR3 (N14931, N14912, N9330, N6922);
nand NAND4 (N14932, N14907, N4461, N3470, N13176);
or OR2 (N14933, N14925, N760);
not NOT1 (N14934, N14929);
or OR4 (N14935, N14933, N10971, N13756, N7229);
or OR2 (N14936, N14935, N13406);
nand NAND3 (N14937, N14923, N5949, N12947);
nor NOR2 (N14938, N14926, N9343);
nand NAND3 (N14939, N14938, N5517, N13526);
or OR4 (N14940, N14928, N7861, N14629, N9175);
or OR3 (N14941, N14932, N8409, N11185);
nand NAND2 (N14942, N14940, N9556);
xor XOR2 (N14943, N14941, N10440);
xor XOR2 (N14944, N14934, N1473);
and AND4 (N14945, N14922, N11371, N10648, N6394);
and AND3 (N14946, N14942, N5730, N544);
nand NAND2 (N14947, N14931, N8765);
buf BUF1 (N14948, N14937);
not NOT1 (N14949, N14943);
not NOT1 (N14950, N14947);
xor XOR2 (N14951, N14946, N7645);
buf BUF1 (N14952, N14950);
buf BUF1 (N14953, N14944);
or OR4 (N14954, N14949, N7504, N14285, N9416);
and AND4 (N14955, N14936, N3195, N11432, N3402);
nor NOR4 (N14956, N14955, N13961, N6871, N7185);
or OR4 (N14957, N14948, N855, N1898, N5524);
or OR2 (N14958, N14953, N11297);
not NOT1 (N14959, N14956);
buf BUF1 (N14960, N14920);
and AND4 (N14961, N14952, N11372, N6617, N3492);
not NOT1 (N14962, N14958);
nand NAND4 (N14963, N14945, N13237, N4743, N2282);
nand NAND4 (N14964, N14930, N11020, N3618, N13336);
not NOT1 (N14965, N14961);
nor NOR4 (N14966, N14951, N867, N12992, N9998);
nor NOR3 (N14967, N14939, N5703, N10645);
and AND4 (N14968, N14954, N11594, N14247, N2320);
not NOT1 (N14969, N14966);
not NOT1 (N14970, N14968);
nand NAND2 (N14971, N14969, N13067);
buf BUF1 (N14972, N14967);
nand NAND3 (N14973, N14957, N9458, N112);
or OR2 (N14974, N14970, N14785);
xor XOR2 (N14975, N14972, N2359);
xor XOR2 (N14976, N14971, N9591);
or OR2 (N14977, N14976, N7875);
not NOT1 (N14978, N14977);
buf BUF1 (N14979, N14973);
xor XOR2 (N14980, N14974, N5073);
not NOT1 (N14981, N14964);
nor NOR4 (N14982, N14979, N923, N11454, N4988);
and AND3 (N14983, N14978, N8745, N7922);
nor NOR2 (N14984, N14983, N11193);
buf BUF1 (N14985, N14959);
not NOT1 (N14986, N14980);
nand NAND3 (N14987, N14965, N12975, N13511);
nor NOR2 (N14988, N14975, N1627);
xor XOR2 (N14989, N14988, N1529);
and AND2 (N14990, N14960, N9910);
xor XOR2 (N14991, N14987, N11694);
xor XOR2 (N14992, N14981, N6356);
not NOT1 (N14993, N14984);
xor XOR2 (N14994, N14982, N10620);
xor XOR2 (N14995, N14989, N10709);
and AND2 (N14996, N14962, N9651);
or OR3 (N14997, N14992, N918, N337);
not NOT1 (N14998, N14985);
not NOT1 (N14999, N14993);
or OR2 (N15000, N14991, N7753);
or OR4 (N15001, N14986, N11616, N8862, N10701);
not NOT1 (N15002, N14963);
buf BUF1 (N15003, N14990);
xor XOR2 (N15004, N14998, N4671);
and AND3 (N15005, N14994, N6192, N5642);
or OR4 (N15006, N14995, N1273, N8403, N8325);
buf BUF1 (N15007, N15001);
nor NOR4 (N15008, N15003, N3686, N13750, N9928);
not NOT1 (N15009, N15002);
buf BUF1 (N15010, N15009);
nor NOR4 (N15011, N15006, N4460, N14156, N11849);
not NOT1 (N15012, N15008);
buf BUF1 (N15013, N15010);
not NOT1 (N15014, N15012);
nand NAND4 (N15015, N15007, N8012, N213, N5728);
nand NAND2 (N15016, N15004, N41);
and AND3 (N15017, N15016, N5834, N5877);
buf BUF1 (N15018, N15011);
not NOT1 (N15019, N14999);
not NOT1 (N15020, N14996);
buf BUF1 (N15021, N15000);
nor NOR3 (N15022, N15019, N5005, N8295);
not NOT1 (N15023, N15017);
or OR3 (N15024, N15005, N7749, N276);
and AND3 (N15025, N15013, N4657, N12987);
nor NOR3 (N15026, N15024, N9338, N13425);
and AND3 (N15027, N15026, N1134, N3593);
and AND4 (N15028, N15021, N5488, N4570, N7368);
or OR4 (N15029, N15018, N10026, N3020, N7544);
or OR4 (N15030, N15022, N7630, N4881, N14951);
buf BUF1 (N15031, N15014);
nor NOR3 (N15032, N15028, N11742, N695);
or OR2 (N15033, N15025, N8401);
nor NOR2 (N15034, N15031, N8143);
xor XOR2 (N15035, N15034, N14726);
not NOT1 (N15036, N15020);
and AND4 (N15037, N15035, N9829, N12233, N3925);
nor NOR2 (N15038, N14997, N7746);
nand NAND4 (N15039, N15030, N218, N1148, N13844);
nand NAND3 (N15040, N15029, N1385, N12773);
xor XOR2 (N15041, N15038, N3395);
or OR3 (N15042, N15036, N14485, N3823);
xor XOR2 (N15043, N15023, N5224);
not NOT1 (N15044, N15039);
and AND2 (N15045, N15033, N8441);
xor XOR2 (N15046, N15045, N202);
or OR4 (N15047, N15042, N11087, N9045, N10706);
buf BUF1 (N15048, N15046);
buf BUF1 (N15049, N15015);
nand NAND4 (N15050, N15044, N7020, N9456, N4887);
xor XOR2 (N15051, N15037, N11582);
buf BUF1 (N15052, N15027);
buf BUF1 (N15053, N15052);
xor XOR2 (N15054, N15041, N14390);
or OR3 (N15055, N15051, N5214, N13693);
or OR4 (N15056, N15054, N10775, N14102, N58);
nor NOR3 (N15057, N15056, N6946, N2778);
not NOT1 (N15058, N15055);
not NOT1 (N15059, N15050);
nand NAND2 (N15060, N15048, N10244);
xor XOR2 (N15061, N15060, N11195);
buf BUF1 (N15062, N15053);
buf BUF1 (N15063, N15058);
nor NOR4 (N15064, N15057, N14679, N10098, N1774);
nand NAND3 (N15065, N15040, N1352, N4257);
xor XOR2 (N15066, N15062, N6532);
buf BUF1 (N15067, N15063);
buf BUF1 (N15068, N15065);
nor NOR2 (N15069, N15064, N2438);
nand NAND2 (N15070, N15066, N12511);
xor XOR2 (N15071, N15032, N5832);
or OR4 (N15072, N15043, N8908, N3454, N1438);
not NOT1 (N15073, N15070);
not NOT1 (N15074, N15073);
xor XOR2 (N15075, N15074, N13436);
nor NOR2 (N15076, N15072, N1832);
nor NOR4 (N15077, N15047, N11807, N9309, N939);
not NOT1 (N15078, N15076);
buf BUF1 (N15079, N15077);
or OR3 (N15080, N15071, N8993, N2304);
buf BUF1 (N15081, N15067);
nand NAND2 (N15082, N15069, N6160);
or OR4 (N15083, N15059, N14117, N10152, N5474);
buf BUF1 (N15084, N15061);
or OR3 (N15085, N15075, N2626, N9206);
or OR4 (N15086, N15084, N13012, N13074, N14948);
or OR2 (N15087, N15078, N2783);
or OR3 (N15088, N15079, N15081, N5693);
not NOT1 (N15089, N7379);
xor XOR2 (N15090, N15068, N603);
and AND4 (N15091, N15049, N2882, N12521, N13000);
buf BUF1 (N15092, N15088);
or OR3 (N15093, N15091, N7925, N13160);
xor XOR2 (N15094, N15080, N6305);
xor XOR2 (N15095, N15094, N3);
nor NOR2 (N15096, N15086, N8447);
and AND3 (N15097, N15092, N646, N8591);
and AND4 (N15098, N15089, N2745, N3970, N581);
buf BUF1 (N15099, N15087);
nor NOR4 (N15100, N15083, N3565, N11572, N1992);
not NOT1 (N15101, N15100);
not NOT1 (N15102, N15098);
not NOT1 (N15103, N15082);
buf BUF1 (N15104, N15085);
buf BUF1 (N15105, N15101);
buf BUF1 (N15106, N15099);
not NOT1 (N15107, N15095);
not NOT1 (N15108, N15103);
or OR3 (N15109, N15104, N11678, N14998);
not NOT1 (N15110, N15097);
nand NAND4 (N15111, N15096, N13944, N5467, N2121);
nor NOR2 (N15112, N15111, N9878);
or OR2 (N15113, N15105, N12368);
or OR4 (N15114, N15102, N5564, N7544, N11930);
buf BUF1 (N15115, N15108);
xor XOR2 (N15116, N15110, N11245);
buf BUF1 (N15117, N15109);
and AND2 (N15118, N15107, N1244);
buf BUF1 (N15119, N15116);
nand NAND4 (N15120, N15114, N12212, N10222, N11879);
nand NAND2 (N15121, N15106, N1654);
buf BUF1 (N15122, N15113);
nand NAND2 (N15123, N15118, N3949);
buf BUF1 (N15124, N15112);
buf BUF1 (N15125, N15120);
nand NAND4 (N15126, N15115, N3689, N8467, N8260);
nor NOR4 (N15127, N15090, N1880, N947, N7555);
not NOT1 (N15128, N15117);
nand NAND4 (N15129, N15124, N11201, N4968, N14885);
or OR2 (N15130, N15121, N3885);
xor XOR2 (N15131, N15126, N12214);
buf BUF1 (N15132, N15119);
nor NOR2 (N15133, N15129, N10134);
and AND4 (N15134, N15093, N9174, N12492, N11369);
or OR2 (N15135, N15131, N11876);
xor XOR2 (N15136, N15128, N12462);
xor XOR2 (N15137, N15133, N10146);
nor NOR3 (N15138, N15134, N9351, N1789);
not NOT1 (N15139, N15135);
xor XOR2 (N15140, N15123, N7268);
not NOT1 (N15141, N15139);
nor NOR4 (N15142, N15122, N12805, N3271, N11124);
and AND3 (N15143, N15132, N8015, N14335);
buf BUF1 (N15144, N15127);
or OR3 (N15145, N15136, N3825, N916);
not NOT1 (N15146, N15140);
nor NOR2 (N15147, N15145, N4041);
buf BUF1 (N15148, N15147);
nand NAND2 (N15149, N15130, N11524);
nor NOR3 (N15150, N15148, N5631, N12088);
or OR4 (N15151, N15149, N8053, N10454, N9489);
not NOT1 (N15152, N15151);
nand NAND2 (N15153, N15137, N7947);
buf BUF1 (N15154, N15142);
and AND2 (N15155, N15150, N11409);
buf BUF1 (N15156, N15144);
xor XOR2 (N15157, N15138, N10483);
and AND3 (N15158, N15153, N12391, N13800);
buf BUF1 (N15159, N15157);
or OR2 (N15160, N15146, N12605);
buf BUF1 (N15161, N15154);
nand NAND4 (N15162, N15141, N3342, N14740, N4566);
buf BUF1 (N15163, N15143);
nor NOR2 (N15164, N15156, N4536);
and AND3 (N15165, N15162, N6191, N11860);
not NOT1 (N15166, N15152);
or OR3 (N15167, N15165, N11790, N9701);
nor NOR4 (N15168, N15163, N5846, N8100, N3361);
nor NOR2 (N15169, N15160, N5885);
xor XOR2 (N15170, N15158, N9927);
nand NAND4 (N15171, N15155, N11880, N4601, N14952);
nand NAND3 (N15172, N15170, N11616, N7754);
nand NAND2 (N15173, N15166, N4363);
not NOT1 (N15174, N15159);
and AND2 (N15175, N15171, N1297);
xor XOR2 (N15176, N15172, N13586);
nor NOR3 (N15177, N15175, N8270, N9311);
or OR4 (N15178, N15168, N10075, N13525, N12859);
buf BUF1 (N15179, N15176);
or OR3 (N15180, N15161, N9986, N3059);
buf BUF1 (N15181, N15167);
xor XOR2 (N15182, N15179, N10047);
xor XOR2 (N15183, N15125, N1656);
not NOT1 (N15184, N15178);
buf BUF1 (N15185, N15169);
nor NOR3 (N15186, N15180, N8639, N4746);
xor XOR2 (N15187, N15185, N14580);
buf BUF1 (N15188, N15164);
or OR3 (N15189, N15174, N6872, N7947);
and AND3 (N15190, N15187, N133, N14681);
buf BUF1 (N15191, N15188);
nand NAND3 (N15192, N15186, N4542, N3929);
buf BUF1 (N15193, N15191);
and AND4 (N15194, N15189, N4373, N14562, N4400);
nand NAND2 (N15195, N15173, N102);
not NOT1 (N15196, N15181);
not NOT1 (N15197, N15194);
not NOT1 (N15198, N15193);
xor XOR2 (N15199, N15196, N5493);
or OR2 (N15200, N15199, N273);
nor NOR2 (N15201, N15192, N3932);
and AND4 (N15202, N15184, N9599, N13144, N6656);
nor NOR2 (N15203, N15202, N12587);
buf BUF1 (N15204, N15182);
xor XOR2 (N15205, N15201, N13284);
not NOT1 (N15206, N15195);
and AND2 (N15207, N15204, N3524);
buf BUF1 (N15208, N15207);
nand NAND3 (N15209, N15203, N8843, N5682);
not NOT1 (N15210, N15190);
not NOT1 (N15211, N15198);
nand NAND2 (N15212, N15177, N12289);
xor XOR2 (N15213, N15206, N9955);
buf BUF1 (N15214, N15209);
nand NAND2 (N15215, N15200, N5651);
or OR2 (N15216, N15208, N1183);
buf BUF1 (N15217, N15216);
xor XOR2 (N15218, N15197, N487);
and AND4 (N15219, N15215, N13344, N11976, N9655);
xor XOR2 (N15220, N15212, N6357);
and AND4 (N15221, N15220, N5600, N12429, N7022);
buf BUF1 (N15222, N15213);
or OR4 (N15223, N15183, N12880, N13244, N11868);
and AND2 (N15224, N15205, N4262);
and AND4 (N15225, N15211, N14602, N14667, N2467);
xor XOR2 (N15226, N15217, N14657);
nand NAND2 (N15227, N15221, N8494);
xor XOR2 (N15228, N15223, N3277);
not NOT1 (N15229, N15210);
nand NAND2 (N15230, N15222, N4562);
or OR3 (N15231, N15228, N14778, N3686);
not NOT1 (N15232, N15225);
not NOT1 (N15233, N15227);
nor NOR2 (N15234, N15214, N13171);
buf BUF1 (N15235, N15231);
xor XOR2 (N15236, N15234, N1276);
and AND2 (N15237, N15218, N6636);
or OR2 (N15238, N15237, N8274);
and AND2 (N15239, N15224, N3824);
buf BUF1 (N15240, N15229);
buf BUF1 (N15241, N15238);
nand NAND2 (N15242, N15232, N5691);
or OR3 (N15243, N15219, N9296, N8804);
xor XOR2 (N15244, N15241, N394);
nand NAND4 (N15245, N15230, N11774, N11462, N4439);
xor XOR2 (N15246, N15239, N4180);
not NOT1 (N15247, N15233);
or OR3 (N15248, N15246, N4694, N2216);
nand NAND3 (N15249, N15243, N2401, N8429);
or OR4 (N15250, N15236, N8835, N351, N14907);
and AND2 (N15251, N15244, N8067);
or OR3 (N15252, N15242, N7817, N10803);
not NOT1 (N15253, N15250);
buf BUF1 (N15254, N15245);
xor XOR2 (N15255, N15235, N12053);
not NOT1 (N15256, N15249);
nor NOR3 (N15257, N15251, N12803, N13081);
nor NOR2 (N15258, N15256, N2721);
buf BUF1 (N15259, N15258);
or OR4 (N15260, N15259, N1930, N10289, N10616);
nand NAND2 (N15261, N15253, N8360);
nor NOR2 (N15262, N15261, N10410);
and AND2 (N15263, N15260, N3389);
not NOT1 (N15264, N15247);
not NOT1 (N15265, N15264);
and AND4 (N15266, N15265, N3977, N10184, N6362);
nor NOR3 (N15267, N15255, N4752, N7900);
not NOT1 (N15268, N15248);
or OR4 (N15269, N15226, N5768, N10953, N8671);
buf BUF1 (N15270, N15257);
xor XOR2 (N15271, N15263, N11959);
and AND4 (N15272, N15268, N13127, N7470, N9807);
nor NOR3 (N15273, N15252, N6849, N9904);
buf BUF1 (N15274, N15272);
xor XOR2 (N15275, N15240, N7991);
buf BUF1 (N15276, N15266);
nand NAND3 (N15277, N15262, N923, N4525);
nor NOR2 (N15278, N15273, N8622);
nor NOR3 (N15279, N15267, N9012, N4007);
xor XOR2 (N15280, N15269, N13035);
not NOT1 (N15281, N15270);
not NOT1 (N15282, N15279);
nand NAND2 (N15283, N15277, N13782);
xor XOR2 (N15284, N15276, N13378);
and AND4 (N15285, N15278, N11634, N11733, N8112);
or OR3 (N15286, N15283, N13801, N5383);
nor NOR3 (N15287, N15280, N14503, N7793);
xor XOR2 (N15288, N15282, N9259);
xor XOR2 (N15289, N15275, N6036);
nor NOR4 (N15290, N15285, N11689, N9056, N13948);
xor XOR2 (N15291, N15288, N12523);
nand NAND3 (N15292, N15271, N11980, N8662);
nand NAND3 (N15293, N15291, N7383, N3516);
buf BUF1 (N15294, N15289);
and AND3 (N15295, N15292, N2176, N6415);
buf BUF1 (N15296, N15284);
and AND4 (N15297, N15294, N6082, N4332, N8567);
xor XOR2 (N15298, N15295, N3096);
not NOT1 (N15299, N15293);
buf BUF1 (N15300, N15296);
or OR2 (N15301, N15298, N7691);
nor NOR2 (N15302, N15301, N3474);
buf BUF1 (N15303, N15302);
not NOT1 (N15304, N15297);
or OR2 (N15305, N15286, N748);
or OR2 (N15306, N15300, N826);
nand NAND4 (N15307, N15305, N14312, N13174, N15290);
not NOT1 (N15308, N7016);
xor XOR2 (N15309, N15304, N6584);
buf BUF1 (N15310, N15281);
buf BUF1 (N15311, N15308);
buf BUF1 (N15312, N15274);
buf BUF1 (N15313, N15310);
not NOT1 (N15314, N15313);
nand NAND4 (N15315, N15314, N2885, N9076, N6057);
and AND4 (N15316, N15312, N1552, N9195, N2947);
buf BUF1 (N15317, N15287);
xor XOR2 (N15318, N15303, N3101);
xor XOR2 (N15319, N15254, N791);
nand NAND3 (N15320, N15315, N7281, N9623);
buf BUF1 (N15321, N15306);
not NOT1 (N15322, N15316);
nand NAND4 (N15323, N15319, N4541, N12733, N410);
not NOT1 (N15324, N15317);
xor XOR2 (N15325, N15320, N13623);
nand NAND3 (N15326, N15323, N13882, N15309);
or OR3 (N15327, N2934, N4120, N6357);
xor XOR2 (N15328, N15322, N9256);
nor NOR4 (N15329, N15326, N7113, N11138, N11606);
or OR2 (N15330, N15311, N14019);
or OR2 (N15331, N15330, N702);
xor XOR2 (N15332, N15324, N11425);
or OR3 (N15333, N15331, N4538, N5567);
or OR4 (N15334, N15307, N10338, N458, N9004);
and AND4 (N15335, N15333, N8221, N13982, N10178);
or OR4 (N15336, N15318, N1173, N191, N1772);
or OR4 (N15337, N15328, N8513, N4770, N2355);
nand NAND3 (N15338, N15336, N13378, N333);
nor NOR3 (N15339, N15321, N8307, N2152);
or OR4 (N15340, N15327, N14743, N2035, N14353);
and AND4 (N15341, N15299, N6868, N8863, N7713);
buf BUF1 (N15342, N15332);
xor XOR2 (N15343, N15342, N3550);
nor NOR2 (N15344, N15338, N1847);
xor XOR2 (N15345, N15341, N4676);
buf BUF1 (N15346, N15325);
not NOT1 (N15347, N15345);
nand NAND4 (N15348, N15347, N8731, N7223, N6109);
buf BUF1 (N15349, N15334);
buf BUF1 (N15350, N15340);
buf BUF1 (N15351, N15335);
xor XOR2 (N15352, N15349, N2470);
buf BUF1 (N15353, N15352);
xor XOR2 (N15354, N15339, N194);
buf BUF1 (N15355, N15329);
and AND2 (N15356, N15350, N368);
xor XOR2 (N15357, N15344, N662);
buf BUF1 (N15358, N15357);
nor NOR3 (N15359, N15346, N426, N2940);
buf BUF1 (N15360, N15348);
nand NAND4 (N15361, N15351, N6885, N6016, N6449);
or OR2 (N15362, N15354, N1837);
or OR4 (N15363, N15361, N4548, N10789, N9108);
nor NOR2 (N15364, N15359, N1608);
not NOT1 (N15365, N15362);
not NOT1 (N15366, N15343);
nand NAND4 (N15367, N15360, N9396, N286, N10178);
buf BUF1 (N15368, N15355);
or OR3 (N15369, N15358, N11247, N8814);
or OR4 (N15370, N15367, N6386, N4069, N6792);
nor NOR2 (N15371, N15363, N10472);
nor NOR4 (N15372, N15366, N3640, N4512, N13827);
and AND2 (N15373, N15370, N13956);
buf BUF1 (N15374, N15337);
buf BUF1 (N15375, N15369);
and AND4 (N15376, N15374, N5697, N1655, N4985);
and AND2 (N15377, N15376, N3524);
nor NOR2 (N15378, N15356, N773);
xor XOR2 (N15379, N15372, N8511);
or OR3 (N15380, N15379, N1380, N927);
buf BUF1 (N15381, N15364);
not NOT1 (N15382, N15381);
and AND4 (N15383, N15380, N9157, N7831, N13592);
and AND2 (N15384, N15375, N13259);
nor NOR2 (N15385, N15373, N4219);
nand NAND3 (N15386, N15365, N15152, N4606);
not NOT1 (N15387, N15371);
nand NAND4 (N15388, N15387, N2110, N6243, N1782);
or OR2 (N15389, N15353, N4269);
or OR4 (N15390, N15384, N9212, N9642, N6312);
nand NAND3 (N15391, N15385, N4588, N5719);
and AND2 (N15392, N15383, N5109);
and AND3 (N15393, N15391, N3052, N15074);
nor NOR3 (N15394, N15377, N1825, N9232);
nand NAND3 (N15395, N15388, N446, N11387);
xor XOR2 (N15396, N15378, N3624);
not NOT1 (N15397, N15368);
not NOT1 (N15398, N15390);
nand NAND3 (N15399, N15382, N4234, N9796);
nand NAND3 (N15400, N15396, N10931, N4341);
not NOT1 (N15401, N15398);
nand NAND4 (N15402, N15395, N3064, N1270, N4925);
buf BUF1 (N15403, N15392);
and AND2 (N15404, N15401, N13789);
not NOT1 (N15405, N15389);
not NOT1 (N15406, N15404);
or OR3 (N15407, N15393, N3307, N12141);
or OR2 (N15408, N15402, N9190);
nor NOR2 (N15409, N15403, N7657);
xor XOR2 (N15410, N15405, N13125);
not NOT1 (N15411, N15386);
nand NAND4 (N15412, N15406, N8195, N2740, N10710);
nor NOR2 (N15413, N15394, N3484);
nand NAND2 (N15414, N15397, N12159);
not NOT1 (N15415, N15413);
nor NOR3 (N15416, N15412, N12034, N11956);
xor XOR2 (N15417, N15399, N7291);
nand NAND4 (N15418, N15411, N13477, N182, N12568);
xor XOR2 (N15419, N15414, N4193);
nand NAND3 (N15420, N15416, N8438, N12834);
xor XOR2 (N15421, N15420, N9657);
or OR4 (N15422, N15410, N5571, N7963, N1451);
nor NOR2 (N15423, N15408, N6352);
and AND2 (N15424, N15417, N11127);
or OR3 (N15425, N15421, N12153, N1888);
not NOT1 (N15426, N15409);
and AND2 (N15427, N15419, N10034);
or OR2 (N15428, N15422, N5933);
not NOT1 (N15429, N15424);
xor XOR2 (N15430, N15427, N5730);
nor NOR2 (N15431, N15407, N4717);
or OR4 (N15432, N15430, N3409, N2497, N11969);
not NOT1 (N15433, N15425);
nand NAND3 (N15434, N15426, N8149, N85);
xor XOR2 (N15435, N15434, N58);
xor XOR2 (N15436, N15432, N1464);
nand NAND3 (N15437, N15435, N7970, N5294);
nand NAND2 (N15438, N15429, N7884);
and AND2 (N15439, N15431, N706);
buf BUF1 (N15440, N15418);
xor XOR2 (N15441, N15400, N2884);
nand NAND4 (N15442, N15440, N3192, N4719, N15318);
not NOT1 (N15443, N15433);
nand NAND3 (N15444, N15428, N12434, N10874);
and AND3 (N15445, N15423, N5540, N14383);
not NOT1 (N15446, N15444);
and AND3 (N15447, N15443, N5736, N14055);
or OR4 (N15448, N15442, N478, N14344, N2735);
xor XOR2 (N15449, N15415, N5597);
nor NOR2 (N15450, N15441, N10722);
and AND3 (N15451, N15437, N3471, N559);
xor XOR2 (N15452, N15447, N5338);
not NOT1 (N15453, N15438);
nor NOR4 (N15454, N15448, N5264, N3804, N12879);
buf BUF1 (N15455, N15450);
buf BUF1 (N15456, N15445);
not NOT1 (N15457, N15446);
xor XOR2 (N15458, N15449, N7277);
xor XOR2 (N15459, N15456, N12476);
not NOT1 (N15460, N15455);
buf BUF1 (N15461, N15452);
nand NAND3 (N15462, N15459, N5758, N2743);
buf BUF1 (N15463, N15460);
or OR3 (N15464, N15454, N3574, N2796);
and AND2 (N15465, N15453, N5434);
nor NOR4 (N15466, N15458, N3777, N852, N4943);
nand NAND2 (N15467, N15462, N4535);
nand NAND4 (N15468, N15465, N9274, N9753, N6478);
buf BUF1 (N15469, N15464);
and AND4 (N15470, N15451, N13454, N7496, N12943);
buf BUF1 (N15471, N15469);
nand NAND3 (N15472, N15461, N10204, N5025);
xor XOR2 (N15473, N15472, N13175);
and AND4 (N15474, N15463, N14409, N9456, N7970);
or OR3 (N15475, N15468, N14828, N10885);
buf BUF1 (N15476, N15471);
or OR2 (N15477, N15476, N5369);
buf BUF1 (N15478, N15477);
or OR2 (N15479, N15474, N12819);
nor NOR3 (N15480, N15466, N14663, N592);
nand NAND3 (N15481, N15470, N4566, N14216);
buf BUF1 (N15482, N15467);
not NOT1 (N15483, N15480);
nand NAND3 (N15484, N15481, N5570, N8486);
buf BUF1 (N15485, N15478);
xor XOR2 (N15486, N15475, N540);
not NOT1 (N15487, N15484);
xor XOR2 (N15488, N15483, N12252);
or OR3 (N15489, N15479, N4076, N15181);
and AND2 (N15490, N15457, N9184);
buf BUF1 (N15491, N15489);
buf BUF1 (N15492, N15491);
buf BUF1 (N15493, N15492);
xor XOR2 (N15494, N15482, N1960);
xor XOR2 (N15495, N15494, N7007);
not NOT1 (N15496, N15436);
nand NAND3 (N15497, N15473, N9816, N8490);
not NOT1 (N15498, N15487);
or OR4 (N15499, N15493, N3381, N10843, N3437);
nand NAND2 (N15500, N15495, N4428);
buf BUF1 (N15501, N15485);
and AND2 (N15502, N15501, N14865);
not NOT1 (N15503, N15439);
not NOT1 (N15504, N15497);
and AND3 (N15505, N15496, N4942, N5478);
nor NOR2 (N15506, N15505, N5137);
nor NOR2 (N15507, N15499, N4280);
or OR2 (N15508, N15486, N9386);
nand NAND4 (N15509, N15504, N11981, N736, N10423);
and AND3 (N15510, N15506, N14751, N14697);
xor XOR2 (N15511, N15509, N1525);
nand NAND2 (N15512, N15500, N12386);
nor NOR2 (N15513, N15503, N3794);
or OR4 (N15514, N15488, N2308, N7594, N15375);
xor XOR2 (N15515, N15514, N1908);
buf BUF1 (N15516, N15515);
or OR2 (N15517, N15508, N3457);
nand NAND2 (N15518, N15510, N12655);
not NOT1 (N15519, N15511);
xor XOR2 (N15520, N15512, N14915);
xor XOR2 (N15521, N15520, N3175);
not NOT1 (N15522, N15507);
not NOT1 (N15523, N15518);
buf BUF1 (N15524, N15517);
xor XOR2 (N15525, N15498, N7615);
and AND4 (N15526, N15490, N14798, N14476, N4623);
buf BUF1 (N15527, N15522);
buf BUF1 (N15528, N15519);
not NOT1 (N15529, N15513);
xor XOR2 (N15530, N15526, N3861);
and AND3 (N15531, N15528, N15320, N13710);
and AND4 (N15532, N15523, N6711, N11908, N6063);
nor NOR4 (N15533, N15502, N7515, N14523, N7993);
nor NOR4 (N15534, N15533, N8028, N1850, N11074);
nor NOR2 (N15535, N15532, N5045);
not NOT1 (N15536, N15521);
nor NOR2 (N15537, N15527, N5291);
or OR3 (N15538, N15530, N14482, N15191);
nor NOR4 (N15539, N15531, N7340, N1529, N276);
not NOT1 (N15540, N15535);
not NOT1 (N15541, N15537);
nand NAND4 (N15542, N15540, N14330, N15234, N8167);
or OR2 (N15543, N15542, N11884);
not NOT1 (N15544, N15529);
buf BUF1 (N15545, N15534);
and AND3 (N15546, N15538, N13063, N2156);
buf BUF1 (N15547, N15545);
nor NOR4 (N15548, N15547, N11644, N6880, N10859);
or OR2 (N15549, N15525, N11111);
and AND3 (N15550, N15546, N4511, N1408);
nor NOR2 (N15551, N15543, N7791);
nand NAND3 (N15552, N15544, N7412, N6024);
not NOT1 (N15553, N15548);
or OR3 (N15554, N15550, N453, N8744);
nand NAND4 (N15555, N15516, N12089, N2615, N12006);
or OR3 (N15556, N15541, N14246, N10721);
or OR3 (N15557, N15524, N9590, N5868);
xor XOR2 (N15558, N15549, N5217);
buf BUF1 (N15559, N15536);
not NOT1 (N15560, N15555);
or OR4 (N15561, N15539, N12652, N15264, N13845);
xor XOR2 (N15562, N15559, N10824);
not NOT1 (N15563, N15560);
xor XOR2 (N15564, N15556, N1842);
nor NOR2 (N15565, N15557, N7331);
nor NOR4 (N15566, N15562, N278, N849, N15327);
xor XOR2 (N15567, N15551, N13023);
and AND3 (N15568, N15553, N3397, N9656);
and AND3 (N15569, N15554, N13695, N5777);
or OR2 (N15570, N15565, N12163);
or OR3 (N15571, N15552, N13925, N14619);
or OR3 (N15572, N15566, N965, N1470);
not NOT1 (N15573, N15564);
and AND2 (N15574, N15568, N469);
and AND4 (N15575, N15573, N6881, N5379, N13266);
nand NAND2 (N15576, N15570, N8638);
xor XOR2 (N15577, N15574, N3113);
nand NAND4 (N15578, N15576, N9068, N7750, N9347);
or OR2 (N15579, N15567, N14231);
or OR2 (N15580, N15572, N14292);
nor NOR3 (N15581, N15579, N5323, N8116);
nand NAND4 (N15582, N15581, N13689, N12228, N6193);
or OR4 (N15583, N15582, N6250, N7091, N8238);
or OR2 (N15584, N15583, N15047);
not NOT1 (N15585, N15558);
nand NAND4 (N15586, N15585, N2789, N9399, N13146);
or OR3 (N15587, N15586, N3025, N7931);
xor XOR2 (N15588, N15577, N7381);
xor XOR2 (N15589, N15561, N980);
and AND2 (N15590, N15587, N12982);
and AND4 (N15591, N15569, N11246, N13683, N3765);
or OR2 (N15592, N15563, N1709);
not NOT1 (N15593, N15591);
nor NOR4 (N15594, N15580, N13494, N11016, N12803);
not NOT1 (N15595, N15589);
xor XOR2 (N15596, N15578, N8449);
or OR3 (N15597, N15590, N3040, N10994);
or OR2 (N15598, N15595, N11705);
or OR3 (N15599, N15597, N12584, N13213);
nor NOR3 (N15600, N15588, N15351, N3762);
buf BUF1 (N15601, N15584);
and AND3 (N15602, N15594, N1632, N13612);
nand NAND3 (N15603, N15596, N6172, N6164);
and AND3 (N15604, N15602, N3638, N9802);
buf BUF1 (N15605, N15571);
nand NAND2 (N15606, N15605, N11513);
buf BUF1 (N15607, N15599);
nor NOR4 (N15608, N15601, N930, N14031, N120);
nand NAND3 (N15609, N15604, N1574, N8256);
nand NAND4 (N15610, N15575, N594, N13704, N659);
nor NOR3 (N15611, N15606, N6157, N10926);
nor NOR3 (N15612, N15609, N9522, N10025);
nand NAND4 (N15613, N15607, N957, N13772, N8173);
buf BUF1 (N15614, N15612);
nor NOR2 (N15615, N15611, N7020);
or OR4 (N15616, N15600, N3500, N9369, N3489);
nand NAND3 (N15617, N15616, N3245, N13707);
xor XOR2 (N15618, N15593, N4716);
not NOT1 (N15619, N15610);
buf BUF1 (N15620, N15619);
nand NAND3 (N15621, N15603, N9046, N5602);
nand NAND4 (N15622, N15613, N10447, N6617, N7622);
and AND4 (N15623, N15592, N14477, N14597, N8126);
nand NAND2 (N15624, N15620, N7130);
not NOT1 (N15625, N15622);
not NOT1 (N15626, N15614);
or OR3 (N15627, N15624, N8510, N12092);
and AND4 (N15628, N15608, N2115, N9019, N972);
nand NAND3 (N15629, N15617, N11894, N13500);
and AND3 (N15630, N15626, N619, N4335);
not NOT1 (N15631, N15615);
buf BUF1 (N15632, N15627);
or OR3 (N15633, N15632, N1125, N8607);
buf BUF1 (N15634, N15628);
nand NAND4 (N15635, N15623, N13137, N7693, N10114);
nor NOR4 (N15636, N15625, N12450, N4197, N14914);
nor NOR3 (N15637, N15631, N15214, N2742);
buf BUF1 (N15638, N15637);
or OR4 (N15639, N15638, N1797, N6635, N2391);
or OR4 (N15640, N15618, N8251, N10206, N8226);
nor NOR3 (N15641, N15630, N7664, N14994);
nor NOR4 (N15642, N15633, N1907, N7735, N6057);
xor XOR2 (N15643, N15636, N3609);
buf BUF1 (N15644, N15629);
nor NOR3 (N15645, N15639, N7818, N14630);
nor NOR4 (N15646, N15645, N3511, N46, N5486);
xor XOR2 (N15647, N15634, N2555);
nand NAND2 (N15648, N15621, N9451);
xor XOR2 (N15649, N15641, N4290);
nand NAND4 (N15650, N15642, N705, N1682, N2486);
buf BUF1 (N15651, N15647);
nand NAND4 (N15652, N15644, N15175, N9679, N1108);
xor XOR2 (N15653, N15635, N11520);
nand NAND3 (N15654, N15598, N1482, N3210);
not NOT1 (N15655, N15640);
and AND4 (N15656, N15646, N3729, N11813, N15295);
or OR2 (N15657, N15648, N3525);
buf BUF1 (N15658, N15654);
not NOT1 (N15659, N15649);
xor XOR2 (N15660, N15657, N14178);
and AND4 (N15661, N15651, N2861, N14257, N10566);
or OR2 (N15662, N15661, N1635);
nand NAND3 (N15663, N15653, N6566, N6286);
or OR3 (N15664, N15660, N11557, N737);
not NOT1 (N15665, N15655);
xor XOR2 (N15666, N15665, N156);
nor NOR3 (N15667, N15664, N12767, N2936);
nand NAND4 (N15668, N15666, N2643, N6226, N9466);
nand NAND3 (N15669, N15656, N1930, N3253);
and AND4 (N15670, N15669, N2501, N2677, N12885);
and AND3 (N15671, N15659, N6600, N12565);
not NOT1 (N15672, N15663);
buf BUF1 (N15673, N15671);
nand NAND4 (N15674, N15667, N10664, N15668, N1715);
or OR4 (N15675, N14893, N3429, N10959, N10229);
and AND3 (N15676, N15650, N9605, N7223);
xor XOR2 (N15677, N15674, N11947);
nand NAND4 (N15678, N15672, N6203, N8645, N2934);
not NOT1 (N15679, N15675);
not NOT1 (N15680, N15652);
xor XOR2 (N15681, N15680, N5639);
and AND3 (N15682, N15676, N7599, N12438);
or OR4 (N15683, N15670, N3373, N12240, N13168);
xor XOR2 (N15684, N15679, N4637);
xor XOR2 (N15685, N15681, N10519);
nand NAND4 (N15686, N15685, N14678, N6593, N11431);
xor XOR2 (N15687, N15682, N1281);
or OR2 (N15688, N15662, N5589);
not NOT1 (N15689, N15688);
or OR2 (N15690, N15678, N6531);
not NOT1 (N15691, N15658);
nand NAND2 (N15692, N15673, N4788);
not NOT1 (N15693, N15687);
nand NAND4 (N15694, N15684, N1490, N13285, N14969);
buf BUF1 (N15695, N15683);
and AND4 (N15696, N15694, N2431, N11777, N7052);
nor NOR4 (N15697, N15696, N10367, N4140, N11660);
xor XOR2 (N15698, N15643, N3195);
and AND4 (N15699, N15677, N1991, N5293, N12303);
and AND2 (N15700, N15697, N7443);
and AND2 (N15701, N15698, N13972);
or OR2 (N15702, N15695, N2);
and AND3 (N15703, N15701, N4916, N1989);
not NOT1 (N15704, N15691);
nand NAND2 (N15705, N15702, N11956);
or OR2 (N15706, N15699, N14022);
nand NAND2 (N15707, N15704, N1158);
and AND4 (N15708, N15692, N7072, N15671, N8246);
nor NOR2 (N15709, N15703, N5906);
not NOT1 (N15710, N15705);
buf BUF1 (N15711, N15693);
buf BUF1 (N15712, N15708);
not NOT1 (N15713, N15712);
not NOT1 (N15714, N15711);
buf BUF1 (N15715, N15706);
or OR4 (N15716, N15707, N1306, N5003, N8133);
and AND4 (N15717, N15714, N5595, N2837, N4943);
buf BUF1 (N15718, N15710);
or OR3 (N15719, N15713, N13871, N243);
nor NOR2 (N15720, N15716, N7986);
or OR3 (N15721, N15689, N5013, N1243);
buf BUF1 (N15722, N15715);
buf BUF1 (N15723, N15719);
and AND4 (N15724, N15720, N8787, N4388, N8630);
nor NOR4 (N15725, N15700, N4652, N5055, N169);
and AND4 (N15726, N15721, N4441, N15483, N8484);
xor XOR2 (N15727, N15718, N1292);
nand NAND3 (N15728, N15690, N6490, N5510);
not NOT1 (N15729, N15723);
buf BUF1 (N15730, N15729);
or OR3 (N15731, N15725, N2192, N15100);
nand NAND2 (N15732, N15731, N14673);
not NOT1 (N15733, N15686);
nor NOR3 (N15734, N15722, N13194, N9987);
or OR2 (N15735, N15733, N10675);
nand NAND3 (N15736, N15732, N9383, N10671);
and AND3 (N15737, N15727, N379, N11764);
or OR4 (N15738, N15717, N11663, N6501, N1927);
and AND3 (N15739, N15737, N6067, N9465);
buf BUF1 (N15740, N15726);
buf BUF1 (N15741, N15736);
not NOT1 (N15742, N15709);
buf BUF1 (N15743, N15735);
not NOT1 (N15744, N15724);
and AND3 (N15745, N15743, N14611, N13207);
xor XOR2 (N15746, N15728, N14375);
and AND4 (N15747, N15734, N6132, N12652, N5025);
xor XOR2 (N15748, N15740, N1628);
nand NAND2 (N15749, N15730, N8188);
nor NOR3 (N15750, N15744, N13865, N8019);
xor XOR2 (N15751, N15738, N1076);
nand NAND3 (N15752, N15749, N7156, N14650);
and AND2 (N15753, N15747, N15696);
and AND2 (N15754, N15750, N12430);
nand NAND3 (N15755, N15739, N7094, N8867);
nor NOR4 (N15756, N15754, N6243, N6048, N1056);
nor NOR2 (N15757, N15753, N10971);
nor NOR4 (N15758, N15748, N12637, N13826, N3461);
nor NOR4 (N15759, N15751, N14155, N2940, N123);
nor NOR4 (N15760, N15752, N5730, N13964, N13293);
xor XOR2 (N15761, N15756, N11186);
nand NAND4 (N15762, N15757, N12429, N12674, N15729);
nor NOR3 (N15763, N15762, N8492, N11330);
or OR4 (N15764, N15745, N15147, N12705, N13000);
nand NAND2 (N15765, N15760, N6581);
nor NOR4 (N15766, N15763, N7432, N9366, N14830);
nand NAND2 (N15767, N15742, N1022);
nor NOR2 (N15768, N15755, N6620);
nor NOR4 (N15769, N15764, N3245, N6597, N10287);
nand NAND2 (N15770, N15759, N14292);
nand NAND4 (N15771, N15765, N799, N2407, N533);
buf BUF1 (N15772, N15746);
or OR2 (N15773, N15768, N14958);
nand NAND2 (N15774, N15741, N9445);
nand NAND3 (N15775, N15758, N1381, N15707);
or OR3 (N15776, N15770, N8748, N8784);
nor NOR2 (N15777, N15766, N12758);
xor XOR2 (N15778, N15772, N8006);
xor XOR2 (N15779, N15778, N1755);
or OR2 (N15780, N15774, N5590);
xor XOR2 (N15781, N15775, N7323);
not NOT1 (N15782, N15781);
or OR3 (N15783, N15777, N14076, N12030);
and AND2 (N15784, N15761, N2646);
xor XOR2 (N15785, N15769, N5070);
and AND3 (N15786, N15783, N12811, N524);
nand NAND3 (N15787, N15784, N13184, N9736);
buf BUF1 (N15788, N15780);
nand NAND2 (N15789, N15788, N10259);
and AND2 (N15790, N15767, N15442);
buf BUF1 (N15791, N15789);
or OR3 (N15792, N15785, N13286, N14629);
and AND2 (N15793, N15790, N13033);
nand NAND4 (N15794, N15792, N3875, N11789, N1515);
nand NAND4 (N15795, N15794, N13712, N12748, N6029);
buf BUF1 (N15796, N15786);
nor NOR4 (N15797, N15796, N1986, N18, N367);
nor NOR3 (N15798, N15791, N7348, N11270);
or OR3 (N15799, N15779, N5510, N2463);
buf BUF1 (N15800, N15795);
xor XOR2 (N15801, N15776, N880);
and AND2 (N15802, N15782, N2866);
or OR2 (N15803, N15800, N13600);
not NOT1 (N15804, N15803);
nor NOR2 (N15805, N15793, N6316);
or OR2 (N15806, N15797, N2298);
buf BUF1 (N15807, N15787);
nand NAND3 (N15808, N15807, N10280, N316);
nand NAND4 (N15809, N15806, N9830, N5676, N5425);
buf BUF1 (N15810, N15773);
and AND4 (N15811, N15801, N10094, N15590, N10744);
xor XOR2 (N15812, N15798, N14164);
nand NAND4 (N15813, N15771, N10090, N11223, N13738);
buf BUF1 (N15814, N15812);
nor NOR3 (N15815, N15814, N13510, N5596);
or OR2 (N15816, N15809, N2598);
and AND4 (N15817, N15810, N155, N10989, N2745);
and AND2 (N15818, N15799, N1623);
nand NAND3 (N15819, N15805, N3696, N5025);
buf BUF1 (N15820, N15813);
xor XOR2 (N15821, N15808, N7445);
not NOT1 (N15822, N15816);
or OR2 (N15823, N15804, N13941);
not NOT1 (N15824, N15817);
xor XOR2 (N15825, N15822, N7581);
nand NAND4 (N15826, N15823, N1406, N2698, N2627);
nor NOR2 (N15827, N15826, N2269);
nor NOR4 (N15828, N15818, N8484, N1358, N13067);
or OR2 (N15829, N15825, N7663);
and AND2 (N15830, N15821, N7499);
not NOT1 (N15831, N15828);
or OR4 (N15832, N15824, N2634, N15404, N6824);
xor XOR2 (N15833, N15802, N13165);
buf BUF1 (N15834, N15827);
xor XOR2 (N15835, N15820, N11113);
xor XOR2 (N15836, N15832, N5817);
nand NAND2 (N15837, N15811, N11690);
buf BUF1 (N15838, N15815);
buf BUF1 (N15839, N15837);
or OR3 (N15840, N15839, N5402, N10675);
and AND3 (N15841, N15819, N12762, N8089);
nand NAND2 (N15842, N15833, N11819);
buf BUF1 (N15843, N15842);
and AND3 (N15844, N15835, N13348, N14354);
nor NOR3 (N15845, N15836, N9810, N6559);
xor XOR2 (N15846, N15834, N1775);
buf BUF1 (N15847, N15845);
and AND2 (N15848, N15830, N6658);
and AND4 (N15849, N15838, N3087, N1170, N12377);
nand NAND4 (N15850, N15848, N7349, N8632, N7843);
or OR4 (N15851, N15831, N9757, N15689, N10446);
and AND3 (N15852, N15840, N3574, N12133);
or OR4 (N15853, N15850, N7781, N10404, N2588);
nor NOR2 (N15854, N15851, N3460);
buf BUF1 (N15855, N15847);
xor XOR2 (N15856, N15843, N3845);
xor XOR2 (N15857, N15846, N2571);
not NOT1 (N15858, N15855);
buf BUF1 (N15859, N15856);
xor XOR2 (N15860, N15841, N14609);
nand NAND3 (N15861, N15853, N341, N11758);
nor NOR3 (N15862, N15861, N2305, N2742);
nand NAND2 (N15863, N15854, N13874);
buf BUF1 (N15864, N15860);
nor NOR4 (N15865, N15849, N8289, N11289, N14053);
nand NAND2 (N15866, N15858, N15277);
or OR2 (N15867, N15859, N338);
xor XOR2 (N15868, N15866, N11915);
not NOT1 (N15869, N15852);
nor NOR4 (N15870, N15869, N9809, N13514, N4606);
or OR4 (N15871, N15867, N9646, N13408, N6180);
buf BUF1 (N15872, N15829);
nand NAND3 (N15873, N15857, N6023, N14643);
buf BUF1 (N15874, N15844);
xor XOR2 (N15875, N15865, N6581);
buf BUF1 (N15876, N15868);
and AND4 (N15877, N15873, N11429, N1995, N10506);
not NOT1 (N15878, N15875);
nand NAND2 (N15879, N15874, N10664);
xor XOR2 (N15880, N15863, N5368);
buf BUF1 (N15881, N15864);
nand NAND2 (N15882, N15870, N7721);
and AND2 (N15883, N15877, N15716);
and AND4 (N15884, N15862, N8672, N6570, N10976);
and AND4 (N15885, N15876, N6621, N15335, N9);
and AND4 (N15886, N15882, N10935, N12994, N116);
xor XOR2 (N15887, N15885, N3011);
nand NAND4 (N15888, N15872, N1545, N13341, N6379);
nor NOR3 (N15889, N15879, N15073, N7460);
and AND2 (N15890, N15878, N10779);
nand NAND4 (N15891, N15881, N1190, N5008, N8068);
nor NOR3 (N15892, N15891, N194, N6226);
and AND2 (N15893, N15883, N12237);
xor XOR2 (N15894, N15890, N12035);
xor XOR2 (N15895, N15884, N5397);
or OR4 (N15896, N15894, N2310, N15641, N6431);
and AND3 (N15897, N15896, N15471, N15852);
nor NOR2 (N15898, N15886, N3121);
or OR2 (N15899, N15897, N6081);
nor NOR3 (N15900, N15889, N8298, N13968);
and AND4 (N15901, N15899, N13658, N5053, N11739);
xor XOR2 (N15902, N15871, N3733);
nand NAND3 (N15903, N15892, N158, N15028);
nor NOR4 (N15904, N15901, N12924, N9899, N12387);
nor NOR3 (N15905, N15898, N10986, N10084);
nand NAND4 (N15906, N15903, N767, N12444, N3993);
nand NAND2 (N15907, N15904, N14892);
nand NAND3 (N15908, N15888, N12489, N6968);
nand NAND2 (N15909, N15887, N15607);
and AND2 (N15910, N15905, N5751);
nand NAND2 (N15911, N15908, N15531);
buf BUF1 (N15912, N15907);
nor NOR3 (N15913, N15900, N14048, N1214);
not NOT1 (N15914, N15906);
and AND2 (N15915, N15902, N3723);
or OR3 (N15916, N15895, N1512, N4195);
xor XOR2 (N15917, N15912, N8901);
and AND4 (N15918, N15915, N4571, N14287, N11195);
or OR2 (N15919, N15917, N15615);
xor XOR2 (N15920, N15913, N5974);
xor XOR2 (N15921, N15880, N10721);
nand NAND4 (N15922, N15918, N12964, N8047, N11314);
not NOT1 (N15923, N15916);
not NOT1 (N15924, N15909);
not NOT1 (N15925, N15921);
buf BUF1 (N15926, N15922);
buf BUF1 (N15927, N15910);
and AND2 (N15928, N15924, N1465);
or OR4 (N15929, N15914, N4908, N7648, N2595);
buf BUF1 (N15930, N15920);
xor XOR2 (N15931, N15926, N4233);
and AND2 (N15932, N15925, N381);
nand NAND2 (N15933, N15927, N8944);
or OR4 (N15934, N15928, N5793, N3594, N1598);
and AND2 (N15935, N15932, N6690);
or OR3 (N15936, N15933, N2325, N11206);
nand NAND4 (N15937, N15929, N11432, N3032, N3169);
nand NAND4 (N15938, N15911, N13135, N5931, N1311);
and AND2 (N15939, N15919, N13528);
or OR2 (N15940, N15923, N8486);
nand NAND4 (N15941, N15893, N15805, N11107, N2055);
not NOT1 (N15942, N15938);
nor NOR4 (N15943, N15942, N10195, N6225, N9199);
nor NOR4 (N15944, N15940, N15331, N11964, N12893);
nand NAND4 (N15945, N15931, N14251, N13378, N14792);
nor NOR4 (N15946, N15939, N12561, N3291, N229);
nor NOR4 (N15947, N15935, N7344, N6730, N1420);
nor NOR2 (N15948, N15944, N3437);
and AND4 (N15949, N15947, N2101, N4192, N12189);
or OR3 (N15950, N15934, N5704, N5947);
or OR2 (N15951, N15937, N4444);
xor XOR2 (N15952, N15949, N12190);
nand NAND2 (N15953, N15948, N11111);
nor NOR2 (N15954, N15951, N4018);
xor XOR2 (N15955, N15950, N1049);
nor NOR3 (N15956, N15955, N12291, N15021);
and AND4 (N15957, N15930, N14807, N11469, N6087);
buf BUF1 (N15958, N15936);
not NOT1 (N15959, N15958);
and AND2 (N15960, N15954, N9919);
and AND2 (N15961, N15957, N12746);
or OR4 (N15962, N15961, N1258, N15237, N5159);
xor XOR2 (N15963, N15959, N15069);
or OR4 (N15964, N15953, N1296, N13330, N7362);
or OR3 (N15965, N15960, N4832, N14487);
not NOT1 (N15966, N15962);
nor NOR3 (N15967, N15946, N1913, N12499);
nand NAND4 (N15968, N15945, N15006, N4732, N4724);
nor NOR4 (N15969, N15968, N7827, N5849, N15759);
nand NAND4 (N15970, N15967, N15301, N14712, N5184);
buf BUF1 (N15971, N15966);
buf BUF1 (N15972, N15971);
and AND4 (N15973, N15965, N5620, N8204, N10076);
not NOT1 (N15974, N15943);
not NOT1 (N15975, N15973);
or OR2 (N15976, N15969, N3306);
not NOT1 (N15977, N15963);
or OR2 (N15978, N15974, N3895);
or OR2 (N15979, N15975, N1254);
not NOT1 (N15980, N15977);
nor NOR3 (N15981, N15952, N12751, N8164);
and AND4 (N15982, N15970, N14663, N12788, N12987);
nor NOR2 (N15983, N15964, N3640);
nor NOR2 (N15984, N15976, N2894);
nand NAND3 (N15985, N15980, N4299, N7713);
xor XOR2 (N15986, N15984, N4410);
not NOT1 (N15987, N15978);
buf BUF1 (N15988, N15985);
or OR4 (N15989, N15956, N9155, N4059, N3712);
nor NOR4 (N15990, N15983, N14215, N5597, N11001);
or OR3 (N15991, N15989, N11757, N6261);
xor XOR2 (N15992, N15972, N920);
or OR2 (N15993, N15990, N14144);
and AND4 (N15994, N15988, N8666, N4119, N9893);
buf BUF1 (N15995, N15991);
nand NAND3 (N15996, N15987, N9500, N6945);
not NOT1 (N15997, N15941);
xor XOR2 (N15998, N15994, N10930);
xor XOR2 (N15999, N15995, N3232);
not NOT1 (N16000, N15986);
nand NAND2 (N16001, N15999, N15481);
nand NAND2 (N16002, N16000, N14443);
nor NOR2 (N16003, N15993, N2101);
or OR3 (N16004, N15979, N6393, N11786);
and AND2 (N16005, N15997, N6896);
or OR3 (N16006, N15992, N893, N1524);
xor XOR2 (N16007, N16001, N14746);
nand NAND2 (N16008, N16004, N4777);
not NOT1 (N16009, N15996);
or OR4 (N16010, N15998, N8924, N9101, N9347);
nand NAND3 (N16011, N15981, N933, N15853);
and AND4 (N16012, N16008, N15804, N4933, N8513);
and AND2 (N16013, N16010, N6930);
or OR2 (N16014, N16002, N7152);
and AND2 (N16015, N16013, N8471);
or OR3 (N16016, N16012, N11043, N11421);
or OR3 (N16017, N16005, N1989, N5502);
endmodule