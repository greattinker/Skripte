// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11;

output N509,N492,N504,N505,N510,N506,N495,N508,N507,N511;

buf BUF1 (N12, N10);
and AND3 (N13, N8, N11, N3);
not NOT1 (N14, N11);
nor NOR2 (N15, N12, N14);
not NOT1 (N16, N7);
nand NAND3 (N17, N12, N13, N5);
or OR2 (N18, N12, N11);
or OR3 (N19, N7, N10, N18);
and AND2 (N20, N2, N16);
not NOT1 (N21, N20);
not NOT1 (N22, N21);
buf BUF1 (N23, N10);
nand NAND2 (N24, N16, N21);
and AND2 (N25, N13, N21);
nand NAND3 (N26, N15, N13, N1);
or OR3 (N27, N24, N5, N14);
and AND4 (N28, N21, N18, N22, N23);
and AND2 (N29, N10, N2);
buf BUF1 (N30, N20);
or OR3 (N31, N2, N25, N11);
not NOT1 (N32, N7);
nand NAND4 (N33, N24, N7, N20, N1);
nand NAND4 (N34, N33, N12, N13, N23);
nor NOR2 (N35, N17, N16);
nand NAND2 (N36, N30, N14);
nand NAND3 (N37, N26, N12, N32);
nor NOR3 (N38, N19, N8, N32);
not NOT1 (N39, N14);
nor NOR3 (N40, N36, N21, N6);
and AND2 (N41, N31, N4);
nand NAND3 (N42, N29, N21, N34);
not NOT1 (N43, N9);
or OR3 (N44, N42, N6, N33);
and AND3 (N45, N27, N5, N13);
nor NOR4 (N46, N40, N3, N35, N13);
buf BUF1 (N47, N38);
xor XOR2 (N48, N39, N2);
or OR4 (N49, N14, N21, N26, N24);
not NOT1 (N50, N44);
buf BUF1 (N51, N49);
and AND2 (N52, N50, N49);
and AND3 (N53, N48, N30, N13);
nand NAND2 (N54, N53, N12);
and AND2 (N55, N37, N25);
xor XOR2 (N56, N43, N37);
or OR2 (N57, N41, N34);
nor NOR2 (N58, N52, N31);
or OR2 (N59, N57, N27);
nand NAND4 (N60, N59, N6, N43, N59);
buf BUF1 (N61, N28);
not NOT1 (N62, N51);
and AND3 (N63, N55, N47, N31);
not NOT1 (N64, N51);
xor XOR2 (N65, N54, N48);
or OR3 (N66, N64, N34, N24);
nor NOR4 (N67, N58, N52, N13, N2);
xor XOR2 (N68, N67, N47);
and AND4 (N69, N45, N50, N2, N27);
or OR3 (N70, N68, N25, N22);
nand NAND2 (N71, N65, N45);
or OR4 (N72, N63, N59, N40, N14);
xor XOR2 (N73, N69, N35);
nor NOR4 (N74, N70, N48, N58, N19);
or OR2 (N75, N46, N21);
nand NAND2 (N76, N71, N24);
or OR3 (N77, N76, N41, N33);
or OR3 (N78, N73, N6, N9);
buf BUF1 (N79, N66);
nor NOR2 (N80, N61, N45);
and AND2 (N81, N80, N70);
nor NOR4 (N82, N72, N74, N66, N6);
nand NAND3 (N83, N10, N40, N80);
not NOT1 (N84, N77);
nor NOR2 (N85, N78, N81);
or OR3 (N86, N44, N14, N12);
nor NOR4 (N87, N85, N2, N61, N20);
nor NOR2 (N88, N82, N8);
nor NOR4 (N89, N56, N80, N59, N83);
or OR4 (N90, N89, N5, N60, N44);
buf BUF1 (N91, N20);
and AND3 (N92, N31, N23, N76);
not NOT1 (N93, N86);
buf BUF1 (N94, N92);
and AND2 (N95, N87, N77);
nand NAND4 (N96, N79, N81, N18, N95);
not NOT1 (N97, N96);
nor NOR4 (N98, N66, N91, N22, N67);
or OR4 (N99, N23, N58, N18, N25);
nand NAND3 (N100, N93, N8, N63);
buf BUF1 (N101, N84);
not NOT1 (N102, N99);
not NOT1 (N103, N100);
nor NOR3 (N104, N97, N80, N16);
nor NOR3 (N105, N102, N16, N52);
nor NOR4 (N106, N103, N68, N16, N66);
or OR2 (N107, N88, N35);
nand NAND4 (N108, N62, N76, N101, N41);
buf BUF1 (N109, N54);
or OR2 (N110, N105, N1);
nor NOR2 (N111, N90, N84);
not NOT1 (N112, N106);
buf BUF1 (N113, N110);
buf BUF1 (N114, N112);
buf BUF1 (N115, N104);
not NOT1 (N116, N109);
and AND3 (N117, N108, N110, N3);
or OR4 (N118, N107, N76, N91, N104);
nand NAND4 (N119, N115, N86, N118, N16);
nor NOR3 (N120, N6, N111, N49);
not NOT1 (N121, N30);
nand NAND2 (N122, N119, N22);
or OR2 (N123, N113, N100);
nor NOR4 (N124, N114, N43, N69, N9);
not NOT1 (N125, N117);
buf BUF1 (N126, N122);
or OR3 (N127, N124, N113, N50);
nor NOR2 (N128, N116, N81);
or OR3 (N129, N121, N98, N102);
buf BUF1 (N130, N36);
buf BUF1 (N131, N125);
or OR3 (N132, N130, N94, N8);
or OR4 (N133, N132, N69, N81, N12);
and AND3 (N134, N40, N92, N36);
nor NOR2 (N135, N126, N126);
or OR2 (N136, N133, N15);
and AND4 (N137, N75, N119, N106, N5);
and AND2 (N138, N128, N6);
buf BUF1 (N139, N123);
buf BUF1 (N140, N139);
nor NOR4 (N141, N129, N132, N122, N100);
nand NAND2 (N142, N138, N6);
or OR4 (N143, N135, N88, N112, N137);
and AND2 (N144, N28, N138);
and AND2 (N145, N136, N43);
xor XOR2 (N146, N145, N17);
xor XOR2 (N147, N127, N42);
buf BUF1 (N148, N143);
not NOT1 (N149, N131);
nand NAND2 (N150, N146, N121);
nand NAND4 (N151, N144, N146, N118, N89);
not NOT1 (N152, N150);
xor XOR2 (N153, N141, N63);
nor NOR4 (N154, N149, N133, N40, N55);
xor XOR2 (N155, N152, N4);
nor NOR4 (N156, N155, N78, N22, N60);
nand NAND2 (N157, N142, N71);
buf BUF1 (N158, N151);
nor NOR3 (N159, N134, N101, N94);
xor XOR2 (N160, N158, N72);
nand NAND4 (N161, N140, N87, N92, N25);
nor NOR3 (N162, N161, N87, N34);
or OR3 (N163, N147, N51, N71);
buf BUF1 (N164, N154);
nand NAND2 (N165, N162, N151);
nor NOR2 (N166, N159, N17);
or OR4 (N167, N166, N19, N42, N2);
or OR4 (N168, N164, N147, N95, N118);
or OR4 (N169, N167, N62, N161, N164);
xor XOR2 (N170, N157, N19);
not NOT1 (N171, N168);
nor NOR2 (N172, N148, N160);
xor XOR2 (N173, N135, N54);
nand NAND3 (N174, N163, N166, N155);
nand NAND3 (N175, N165, N65, N67);
or OR3 (N176, N174, N102, N114);
not NOT1 (N177, N172);
or OR4 (N178, N170, N123, N97, N30);
or OR2 (N179, N173, N100);
buf BUF1 (N180, N179);
or OR4 (N181, N177, N123, N180, N177);
buf BUF1 (N182, N68);
nand NAND2 (N183, N176, N132);
or OR2 (N184, N153, N76);
not NOT1 (N185, N184);
and AND4 (N186, N178, N167, N113, N122);
buf BUF1 (N187, N181);
and AND4 (N188, N183, N28, N123, N54);
and AND3 (N189, N175, N30, N45);
xor XOR2 (N190, N187, N49);
xor XOR2 (N191, N156, N145);
nand NAND3 (N192, N189, N155, N111);
buf BUF1 (N193, N190);
or OR2 (N194, N182, N40);
buf BUF1 (N195, N186);
or OR4 (N196, N194, N8, N105, N185);
nand NAND3 (N197, N136, N23, N22);
not NOT1 (N198, N193);
buf BUF1 (N199, N171);
not NOT1 (N200, N120);
xor XOR2 (N201, N192, N68);
nand NAND4 (N202, N197, N100, N110, N175);
not NOT1 (N203, N169);
buf BUF1 (N204, N201);
xor XOR2 (N205, N204, N110);
not NOT1 (N206, N200);
xor XOR2 (N207, N202, N101);
nand NAND4 (N208, N188, N155, N58, N79);
xor XOR2 (N209, N198, N80);
and AND4 (N210, N199, N64, N48, N52);
nor NOR3 (N211, N205, N51, N119);
buf BUF1 (N212, N196);
and AND3 (N213, N208, N21, N105);
not NOT1 (N214, N195);
and AND2 (N215, N213, N152);
and AND4 (N216, N214, N205, N22, N82);
buf BUF1 (N217, N211);
nor NOR4 (N218, N203, N73, N146, N170);
not NOT1 (N219, N215);
not NOT1 (N220, N207);
and AND2 (N221, N219, N181);
buf BUF1 (N222, N210);
or OR4 (N223, N218, N211, N128, N115);
nor NOR3 (N224, N222, N194, N217);
and AND2 (N225, N213, N52);
or OR4 (N226, N220, N204, N35, N97);
and AND3 (N227, N191, N169, N204);
or OR3 (N228, N227, N79, N175);
or OR2 (N229, N228, N164);
and AND2 (N230, N212, N46);
nand NAND2 (N231, N226, N199);
and AND4 (N232, N229, N92, N203, N122);
nand NAND3 (N233, N232, N27, N216);
xor XOR2 (N234, N63, N66);
not NOT1 (N235, N230);
xor XOR2 (N236, N209, N146);
nand NAND3 (N237, N224, N65, N191);
not NOT1 (N238, N206);
or OR4 (N239, N235, N13, N177, N226);
buf BUF1 (N240, N223);
not NOT1 (N241, N231);
not NOT1 (N242, N225);
nand NAND4 (N243, N221, N65, N126, N95);
nand NAND2 (N244, N238, N157);
or OR2 (N245, N239, N197);
xor XOR2 (N246, N241, N67);
xor XOR2 (N247, N244, N87);
or OR2 (N248, N240, N116);
xor XOR2 (N249, N237, N12);
not NOT1 (N250, N242);
nand NAND4 (N251, N246, N244, N250, N24);
buf BUF1 (N252, N6);
or OR3 (N253, N249, N104, N60);
or OR2 (N254, N251, N48);
not NOT1 (N255, N253);
nor NOR4 (N256, N233, N49, N44, N88);
xor XOR2 (N257, N236, N202);
nand NAND3 (N258, N247, N109, N45);
nor NOR4 (N259, N254, N221, N243, N100);
nor NOR2 (N260, N102, N43);
and AND4 (N261, N258, N134, N42, N30);
and AND4 (N262, N256, N203, N245, N22);
or OR4 (N263, N251, N192, N149, N205);
not NOT1 (N264, N252);
xor XOR2 (N265, N264, N42);
and AND4 (N266, N262, N115, N237, N214);
nand NAND2 (N267, N266, N80);
nand NAND4 (N268, N263, N96, N98, N80);
xor XOR2 (N269, N260, N159);
nand NAND4 (N270, N255, N89, N73, N65);
nor NOR4 (N271, N257, N223, N98, N67);
buf BUF1 (N272, N261);
and AND4 (N273, N271, N237, N75, N186);
buf BUF1 (N274, N267);
nand NAND3 (N275, N268, N79, N200);
xor XOR2 (N276, N269, N270);
nor NOR2 (N277, N55, N184);
not NOT1 (N278, N259);
not NOT1 (N279, N276);
not NOT1 (N280, N278);
xor XOR2 (N281, N275, N216);
or OR3 (N282, N248, N24, N140);
not NOT1 (N283, N281);
nand NAND3 (N284, N272, N194, N206);
buf BUF1 (N285, N265);
and AND3 (N286, N279, N245, N250);
or OR4 (N287, N282, N27, N258, N87);
and AND4 (N288, N273, N253, N245, N248);
buf BUF1 (N289, N285);
buf BUF1 (N290, N274);
and AND2 (N291, N286, N197);
or OR4 (N292, N283, N68, N99, N275);
buf BUF1 (N293, N287);
nor NOR3 (N294, N291, N49, N202);
and AND3 (N295, N294, N88, N65);
xor XOR2 (N296, N292, N40);
xor XOR2 (N297, N280, N266);
nor NOR4 (N298, N284, N281, N87, N44);
xor XOR2 (N299, N297, N218);
nand NAND3 (N300, N295, N1, N4);
nor NOR3 (N301, N234, N122, N7);
or OR4 (N302, N296, N77, N275, N115);
and AND3 (N303, N301, N233, N187);
not NOT1 (N304, N288);
buf BUF1 (N305, N289);
not NOT1 (N306, N304);
xor XOR2 (N307, N306, N141);
and AND4 (N308, N302, N56, N227, N93);
xor XOR2 (N309, N305, N15);
xor XOR2 (N310, N293, N185);
buf BUF1 (N311, N299);
or OR3 (N312, N309, N68, N50);
xor XOR2 (N313, N298, N125);
nor NOR2 (N314, N303, N280);
nand NAND4 (N315, N310, N293, N274, N171);
nor NOR4 (N316, N277, N44, N179, N192);
nor NOR2 (N317, N316, N285);
nor NOR4 (N318, N290, N245, N69, N88);
or OR4 (N319, N308, N296, N135, N213);
and AND2 (N320, N318, N8);
xor XOR2 (N321, N312, N310);
or OR4 (N322, N317, N252, N105, N213);
or OR4 (N323, N311, N140, N184, N65);
or OR4 (N324, N320, N231, N277, N141);
nor NOR4 (N325, N324, N261, N322, N83);
xor XOR2 (N326, N129, N56);
or OR2 (N327, N300, N223);
xor XOR2 (N328, N326, N118);
nor NOR3 (N329, N314, N253, N217);
nor NOR2 (N330, N323, N59);
xor XOR2 (N331, N328, N168);
or OR4 (N332, N315, N201, N122, N45);
xor XOR2 (N333, N329, N101);
xor XOR2 (N334, N307, N266);
or OR4 (N335, N313, N153, N288, N230);
nor NOR3 (N336, N327, N155, N323);
nor NOR3 (N337, N336, N310, N2);
and AND3 (N338, N325, N283, N44);
xor XOR2 (N339, N332, N96);
nor NOR4 (N340, N330, N98, N123, N235);
or OR3 (N341, N319, N14, N10);
nand NAND4 (N342, N337, N256, N90, N239);
or OR4 (N343, N331, N115, N170, N108);
nor NOR3 (N344, N321, N298, N211);
nand NAND4 (N345, N339, N192, N220, N122);
xor XOR2 (N346, N345, N291);
buf BUF1 (N347, N341);
or OR4 (N348, N346, N268, N70, N258);
nor NOR3 (N349, N335, N67, N125);
nor NOR4 (N350, N334, N266, N235, N163);
or OR3 (N351, N342, N84, N116);
nor NOR4 (N352, N333, N82, N250, N316);
buf BUF1 (N353, N349);
xor XOR2 (N354, N353, N176);
buf BUF1 (N355, N344);
and AND3 (N356, N348, N50, N191);
nor NOR3 (N357, N347, N274, N8);
nand NAND4 (N358, N351, N297, N199, N43);
nand NAND4 (N359, N355, N59, N245, N247);
and AND4 (N360, N356, N16, N281, N115);
buf BUF1 (N361, N352);
buf BUF1 (N362, N357);
xor XOR2 (N363, N354, N141);
xor XOR2 (N364, N360, N85);
nand NAND4 (N365, N340, N204, N195, N54);
nor NOR2 (N366, N363, N72);
nand NAND4 (N367, N362, N290, N211, N276);
and AND2 (N368, N366, N119);
nor NOR4 (N369, N365, N162, N176, N159);
xor XOR2 (N370, N359, N3);
or OR2 (N371, N343, N191);
not NOT1 (N372, N364);
and AND4 (N373, N358, N368, N184, N308);
nand NAND4 (N374, N24, N285, N97, N274);
or OR4 (N375, N367, N93, N207, N126);
nor NOR4 (N376, N372, N17, N98, N103);
not NOT1 (N377, N338);
not NOT1 (N378, N361);
nand NAND3 (N379, N371, N129, N87);
xor XOR2 (N380, N377, N15);
buf BUF1 (N381, N375);
and AND4 (N382, N373, N216, N280, N353);
buf BUF1 (N383, N370);
buf BUF1 (N384, N379);
and AND2 (N385, N380, N328);
nor NOR4 (N386, N384, N18, N160, N270);
not NOT1 (N387, N381);
and AND3 (N388, N387, N375, N154);
xor XOR2 (N389, N386, N182);
not NOT1 (N390, N369);
not NOT1 (N391, N385);
nand NAND4 (N392, N382, N2, N115, N93);
not NOT1 (N393, N383);
not NOT1 (N394, N392);
not NOT1 (N395, N378);
xor XOR2 (N396, N350, N84);
and AND4 (N397, N395, N52, N42, N42);
and AND3 (N398, N397, N393, N66);
nand NAND2 (N399, N398, N301);
xor XOR2 (N400, N130, N37);
and AND3 (N401, N396, N398, N202);
nand NAND2 (N402, N401, N286);
nor NOR4 (N403, N389, N72, N53, N158);
nand NAND4 (N404, N403, N96, N75, N193);
or OR4 (N405, N399, N203, N403, N44);
or OR3 (N406, N391, N33, N131);
or OR3 (N407, N388, N341, N14);
not NOT1 (N408, N402);
or OR4 (N409, N390, N105, N381, N373);
nor NOR3 (N410, N394, N16, N187);
or OR2 (N411, N376, N117);
not NOT1 (N412, N406);
or OR4 (N413, N412, N112, N119, N190);
nand NAND3 (N414, N409, N94, N320);
nor NOR3 (N415, N407, N288, N62);
buf BUF1 (N416, N405);
buf BUF1 (N417, N411);
xor XOR2 (N418, N417, N66);
and AND3 (N419, N414, N79, N219);
buf BUF1 (N420, N408);
and AND4 (N421, N374, N411, N69, N402);
nor NOR4 (N422, N421, N37, N185, N101);
nor NOR4 (N423, N415, N398, N93, N14);
buf BUF1 (N424, N416);
nor NOR2 (N425, N413, N351);
not NOT1 (N426, N419);
xor XOR2 (N427, N400, N153);
nor NOR3 (N428, N404, N388, N158);
or OR4 (N429, N424, N246, N305, N237);
xor XOR2 (N430, N428, N138);
or OR3 (N431, N422, N141, N387);
buf BUF1 (N432, N420);
nor NOR4 (N433, N429, N312, N72, N365);
nor NOR3 (N434, N433, N380, N149);
xor XOR2 (N435, N410, N393);
xor XOR2 (N436, N423, N136);
nor NOR3 (N437, N427, N268, N318);
not NOT1 (N438, N426);
and AND3 (N439, N431, N274, N343);
or OR3 (N440, N418, N377, N146);
nand NAND3 (N441, N432, N220, N342);
nor NOR3 (N442, N430, N255, N390);
buf BUF1 (N443, N437);
nand NAND3 (N444, N436, N99, N317);
buf BUF1 (N445, N439);
and AND2 (N446, N445, N196);
and AND4 (N447, N443, N22, N181, N106);
nor NOR2 (N448, N441, N258);
and AND3 (N449, N438, N185, N27);
nand NAND3 (N450, N449, N180, N115);
nand NAND3 (N451, N446, N357, N347);
not NOT1 (N452, N451);
buf BUF1 (N453, N448);
xor XOR2 (N454, N435, N246);
xor XOR2 (N455, N440, N362);
xor XOR2 (N456, N453, N40);
nor NOR2 (N457, N447, N17);
or OR2 (N458, N425, N254);
nor NOR2 (N459, N456, N6);
nand NAND2 (N460, N454, N329);
or OR4 (N461, N459, N256, N436, N56);
not NOT1 (N462, N434);
and AND3 (N463, N452, N322, N366);
nand NAND3 (N464, N458, N216, N38);
nand NAND4 (N465, N463, N126, N186, N31);
buf BUF1 (N466, N460);
nor NOR2 (N467, N466, N92);
buf BUF1 (N468, N461);
nor NOR4 (N469, N444, N271, N184, N389);
xor XOR2 (N470, N467, N229);
buf BUF1 (N471, N465);
xor XOR2 (N472, N464, N288);
xor XOR2 (N473, N442, N258);
or OR2 (N474, N450, N447);
nor NOR3 (N475, N455, N134, N164);
or OR4 (N476, N474, N372, N393, N62);
xor XOR2 (N477, N471, N268);
buf BUF1 (N478, N469);
buf BUF1 (N479, N475);
nor NOR3 (N480, N479, N67, N48);
xor XOR2 (N481, N472, N196);
nand NAND4 (N482, N462, N157, N333, N92);
nand NAND4 (N483, N478, N323, N376, N159);
nand NAND3 (N484, N468, N90, N170);
not NOT1 (N485, N476);
not NOT1 (N486, N470);
or OR2 (N487, N481, N335);
buf BUF1 (N488, N484);
and AND2 (N489, N483, N438);
nand NAND2 (N490, N489, N337);
nor NOR2 (N491, N482, N162);
not NOT1 (N492, N457);
not NOT1 (N493, N480);
nand NAND4 (N494, N493, N249, N338, N33);
buf BUF1 (N495, N490);
buf BUF1 (N496, N491);
and AND3 (N497, N496, N212, N478);
buf BUF1 (N498, N485);
buf BUF1 (N499, N477);
and AND3 (N500, N497, N30, N295);
nand NAND2 (N501, N499, N68);
and AND3 (N502, N494, N149, N417);
or OR3 (N503, N501, N243, N126);
nor NOR4 (N504, N503, N450, N117, N340);
buf BUF1 (N505, N488);
or OR4 (N506, N473, N111, N431, N206);
xor XOR2 (N507, N502, N309);
or OR4 (N508, N500, N252, N347, N490);
and AND4 (N509, N487, N316, N158, N59);
nor NOR4 (N510, N498, N243, N76, N219);
xor XOR2 (N511, N486, N134);
endmodule