// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22;

output N12811,N12792,N12801,N12820,N12818,N12809,N12821,N12816,N12810,N12822;

not NOT1 (N23, N17);
buf BUF1 (N24, N2);
or OR2 (N25, N16, N11);
nor NOR4 (N26, N19, N23, N19, N1);
not NOT1 (N27, N11);
nor NOR3 (N28, N8, N18, N24);
nor NOR2 (N29, N6, N2);
buf BUF1 (N30, N9);
and AND3 (N31, N9, N14, N7);
nand NAND4 (N32, N26, N17, N30, N16);
nand NAND4 (N33, N27, N11, N13, N29);
and AND2 (N34, N17, N20);
nand NAND2 (N35, N20, N29);
xor XOR2 (N36, N17, N5);
not NOT1 (N37, N34);
xor XOR2 (N38, N6, N27);
buf BUF1 (N39, N4);
xor XOR2 (N40, N38, N17);
xor XOR2 (N41, N39, N30);
and AND2 (N42, N31, N40);
and AND2 (N43, N40, N33);
or OR4 (N44, N35, N11, N26, N14);
xor XOR2 (N45, N24, N18);
buf BUF1 (N46, N36);
xor XOR2 (N47, N37, N4);
xor XOR2 (N48, N42, N5);
or OR2 (N49, N44, N27);
xor XOR2 (N50, N41, N6);
or OR4 (N51, N49, N20, N35, N10);
nor NOR2 (N52, N28, N26);
nand NAND2 (N53, N48, N2);
not NOT1 (N54, N50);
buf BUF1 (N55, N51);
xor XOR2 (N56, N25, N21);
not NOT1 (N57, N54);
and AND3 (N58, N46, N19, N50);
nand NAND3 (N59, N47, N30, N56);
xor XOR2 (N60, N34, N53);
buf BUF1 (N61, N4);
xor XOR2 (N62, N60, N46);
and AND3 (N63, N32, N30, N45);
and AND4 (N64, N22, N63, N34, N29);
xor XOR2 (N65, N34, N29);
and AND4 (N66, N52, N56, N16, N55);
xor XOR2 (N67, N35, N1);
and AND2 (N68, N66, N33);
and AND3 (N69, N64, N59, N59);
buf BUF1 (N70, N23);
or OR3 (N71, N57, N17, N54);
nor NOR4 (N72, N70, N14, N2, N71);
xor XOR2 (N73, N41, N44);
not NOT1 (N74, N61);
xor XOR2 (N75, N62, N31);
not NOT1 (N76, N68);
not NOT1 (N77, N73);
nor NOR2 (N78, N67, N61);
or OR3 (N79, N77, N30, N29);
not NOT1 (N80, N78);
nor NOR3 (N81, N75, N67, N70);
nand NAND3 (N82, N69, N19, N73);
nand NAND3 (N83, N76, N48, N34);
not NOT1 (N84, N58);
and AND4 (N85, N72, N13, N62, N35);
and AND3 (N86, N80, N47, N39);
or OR4 (N87, N84, N70, N56, N5);
nor NOR4 (N88, N85, N60, N66, N76);
xor XOR2 (N89, N43, N58);
xor XOR2 (N90, N82, N56);
and AND3 (N91, N87, N53, N4);
not NOT1 (N92, N89);
nor NOR3 (N93, N79, N55, N65);
or OR4 (N94, N23, N77, N67, N64);
buf BUF1 (N95, N92);
not NOT1 (N96, N88);
not NOT1 (N97, N83);
nor NOR4 (N98, N96, N39, N26, N49);
nand NAND3 (N99, N93, N27, N95);
not NOT1 (N100, N74);
nor NOR2 (N101, N58, N45);
or OR4 (N102, N98, N26, N28, N70);
or OR2 (N103, N102, N11);
not NOT1 (N104, N99);
not NOT1 (N105, N103);
not NOT1 (N106, N105);
xor XOR2 (N107, N90, N58);
and AND2 (N108, N107, N58);
not NOT1 (N109, N108);
buf BUF1 (N110, N106);
buf BUF1 (N111, N91);
not NOT1 (N112, N81);
or OR2 (N113, N104, N7);
buf BUF1 (N114, N94);
not NOT1 (N115, N100);
or OR2 (N116, N110, N53);
buf BUF1 (N117, N86);
nor NOR2 (N118, N101, N76);
nor NOR2 (N119, N113, N113);
nand NAND3 (N120, N118, N112, N76);
or OR4 (N121, N40, N52, N89, N63);
nor NOR3 (N122, N111, N61, N41);
nand NAND2 (N123, N116, N120);
or OR4 (N124, N59, N63, N62, N82);
not NOT1 (N125, N115);
nor NOR3 (N126, N97, N15, N56);
xor XOR2 (N127, N123, N27);
and AND3 (N128, N121, N87, N86);
nand NAND4 (N129, N126, N69, N124, N18);
or OR2 (N130, N35, N66);
not NOT1 (N131, N122);
nor NOR2 (N132, N131, N81);
buf BUF1 (N133, N119);
and AND2 (N134, N129, N105);
or OR2 (N135, N134, N1);
nor NOR3 (N136, N117, N21, N32);
buf BUF1 (N137, N135);
xor XOR2 (N138, N114, N39);
xor XOR2 (N139, N127, N128);
not NOT1 (N140, N91);
or OR2 (N141, N125, N119);
or OR2 (N142, N140, N32);
buf BUF1 (N143, N138);
and AND3 (N144, N136, N82, N47);
or OR2 (N145, N142, N13);
or OR3 (N146, N145, N128, N41);
xor XOR2 (N147, N109, N77);
and AND4 (N148, N144, N20, N46, N96);
nor NOR3 (N149, N139, N21, N140);
nor NOR4 (N150, N132, N18, N81, N136);
nand NAND3 (N151, N146, N141, N15);
nor NOR4 (N152, N12, N149, N15, N131);
not NOT1 (N153, N81);
buf BUF1 (N154, N130);
buf BUF1 (N155, N153);
xor XOR2 (N156, N151, N39);
not NOT1 (N157, N143);
or OR3 (N158, N155, N7, N19);
and AND2 (N159, N137, N146);
nand NAND4 (N160, N148, N23, N128, N119);
and AND2 (N161, N156, N1);
xor XOR2 (N162, N150, N19);
not NOT1 (N163, N158);
nand NAND4 (N164, N160, N73, N54, N19);
nor NOR3 (N165, N154, N134, N134);
nand NAND4 (N166, N163, N7, N160, N104);
nand NAND2 (N167, N147, N149);
nor NOR2 (N168, N157, N83);
not NOT1 (N169, N162);
xor XOR2 (N170, N159, N84);
and AND3 (N171, N170, N124, N13);
or OR2 (N172, N168, N49);
or OR4 (N173, N133, N100, N84, N28);
nor NOR4 (N174, N172, N118, N148, N43);
and AND4 (N175, N174, N85, N98, N55);
xor XOR2 (N176, N166, N73);
xor XOR2 (N177, N173, N41);
nor NOR4 (N178, N164, N113, N65, N4);
nor NOR3 (N179, N165, N39, N54);
xor XOR2 (N180, N152, N162);
and AND4 (N181, N179, N69, N52, N14);
and AND4 (N182, N181, N144, N14, N71);
not NOT1 (N183, N178);
or OR4 (N184, N171, N142, N149, N163);
not NOT1 (N185, N169);
nor NOR4 (N186, N177, N144, N171, N114);
nor NOR4 (N187, N167, N83, N74, N64);
or OR2 (N188, N180, N25);
or OR4 (N189, N185, N140, N129, N97);
not NOT1 (N190, N183);
and AND4 (N191, N188, N129, N9, N52);
nor NOR3 (N192, N161, N86, N149);
buf BUF1 (N193, N190);
or OR3 (N194, N175, N43, N177);
nand NAND2 (N195, N194, N64);
or OR3 (N196, N195, N170, N100);
nand NAND4 (N197, N192, N157, N173, N172);
not NOT1 (N198, N176);
or OR4 (N199, N186, N177, N147, N42);
nand NAND2 (N200, N197, N2);
nand NAND3 (N201, N182, N200, N5);
buf BUF1 (N202, N170);
and AND4 (N203, N196, N6, N119, N145);
not NOT1 (N204, N189);
xor XOR2 (N205, N184, N93);
xor XOR2 (N206, N204, N87);
nand NAND2 (N207, N198, N116);
buf BUF1 (N208, N203);
and AND4 (N209, N201, N150, N187, N32);
and AND4 (N210, N97, N171, N139, N65);
nor NOR4 (N211, N202, N45, N10, N23);
nand NAND2 (N212, N199, N200);
and AND2 (N213, N209, N81);
xor XOR2 (N214, N208, N170);
or OR2 (N215, N212, N198);
xor XOR2 (N216, N205, N202);
not NOT1 (N217, N214);
or OR4 (N218, N191, N200, N144, N96);
not NOT1 (N219, N218);
nor NOR2 (N220, N219, N191);
buf BUF1 (N221, N215);
nand NAND4 (N222, N213, N99, N83, N30);
buf BUF1 (N223, N217);
buf BUF1 (N224, N223);
buf BUF1 (N225, N206);
not NOT1 (N226, N224);
nor NOR3 (N227, N226, N206, N31);
buf BUF1 (N228, N227);
not NOT1 (N229, N210);
nand NAND3 (N230, N211, N162, N17);
buf BUF1 (N231, N216);
not NOT1 (N232, N221);
nand NAND2 (N233, N232, N69);
xor XOR2 (N234, N225, N39);
xor XOR2 (N235, N231, N71);
nand NAND2 (N236, N235, N93);
nor NOR2 (N237, N220, N143);
nand NAND2 (N238, N234, N200);
nor NOR2 (N239, N222, N2);
nor NOR2 (N240, N236, N119);
buf BUF1 (N241, N193);
xor XOR2 (N242, N233, N229);
xor XOR2 (N243, N30, N225);
nor NOR3 (N244, N228, N81, N55);
nor NOR2 (N245, N240, N211);
not NOT1 (N246, N242);
buf BUF1 (N247, N207);
nor NOR3 (N248, N244, N76, N128);
xor XOR2 (N249, N239, N242);
and AND4 (N250, N246, N202, N143, N137);
not NOT1 (N251, N230);
not NOT1 (N252, N238);
not NOT1 (N253, N243);
xor XOR2 (N254, N247, N107);
nand NAND4 (N255, N252, N79, N138, N212);
nand NAND4 (N256, N254, N150, N178, N201);
nor NOR4 (N257, N256, N50, N82, N247);
buf BUF1 (N258, N248);
xor XOR2 (N259, N249, N36);
and AND4 (N260, N245, N235, N240, N102);
not NOT1 (N261, N257);
not NOT1 (N262, N241);
buf BUF1 (N263, N262);
buf BUF1 (N264, N260);
not NOT1 (N265, N255);
buf BUF1 (N266, N250);
not NOT1 (N267, N258);
or OR2 (N268, N259, N216);
xor XOR2 (N269, N267, N143);
xor XOR2 (N270, N266, N88);
and AND2 (N271, N269, N178);
or OR4 (N272, N263, N231, N49, N259);
not NOT1 (N273, N272);
and AND2 (N274, N253, N73);
buf BUF1 (N275, N271);
not NOT1 (N276, N265);
nand NAND2 (N277, N251, N237);
nand NAND2 (N278, N157, N258);
nor NOR3 (N279, N268, N35, N257);
and AND3 (N280, N261, N124, N17);
or OR2 (N281, N276, N129);
nor NOR2 (N282, N281, N2);
or OR4 (N283, N270, N30, N132, N100);
and AND4 (N284, N278, N198, N211, N129);
and AND3 (N285, N275, N121, N154);
and AND2 (N286, N279, N243);
buf BUF1 (N287, N273);
xor XOR2 (N288, N284, N122);
or OR2 (N289, N274, N28);
xor XOR2 (N290, N282, N271);
buf BUF1 (N291, N289);
and AND2 (N292, N286, N245);
nor NOR4 (N293, N264, N131, N201, N162);
nand NAND3 (N294, N285, N269, N95);
nand NAND3 (N295, N293, N244, N287);
nand NAND3 (N296, N7, N29, N46);
and AND2 (N297, N290, N3);
and AND3 (N298, N277, N222, N65);
xor XOR2 (N299, N291, N142);
not NOT1 (N300, N294);
buf BUF1 (N301, N295);
nor NOR2 (N302, N297, N197);
or OR2 (N303, N302, N85);
nor NOR3 (N304, N283, N226, N12);
or OR2 (N305, N292, N227);
and AND2 (N306, N298, N243);
and AND4 (N307, N306, N119, N202, N284);
xor XOR2 (N308, N301, N80);
and AND2 (N309, N296, N102);
buf BUF1 (N310, N303);
not NOT1 (N311, N304);
nand NAND3 (N312, N288, N3, N77);
nor NOR3 (N313, N309, N201, N174);
buf BUF1 (N314, N313);
nand NAND3 (N315, N312, N283, N13);
not NOT1 (N316, N315);
xor XOR2 (N317, N299, N73);
buf BUF1 (N318, N308);
and AND3 (N319, N311, N88, N317);
nor NOR2 (N320, N127, N184);
not NOT1 (N321, N318);
nand NAND4 (N322, N319, N305, N55, N251);
nand NAND4 (N323, N222, N240, N280, N103);
nand NAND2 (N324, N72, N108);
not NOT1 (N325, N323);
not NOT1 (N326, N324);
buf BUF1 (N327, N326);
or OR4 (N328, N310, N279, N15, N287);
buf BUF1 (N329, N325);
nand NAND3 (N330, N316, N285, N231);
buf BUF1 (N331, N321);
or OR2 (N332, N327, N182);
not NOT1 (N333, N329);
and AND2 (N334, N307, N315);
not NOT1 (N335, N331);
xor XOR2 (N336, N333, N165);
nand NAND3 (N337, N330, N324, N152);
or OR2 (N338, N334, N215);
nand NAND2 (N339, N314, N16);
nor NOR3 (N340, N322, N8, N95);
xor XOR2 (N341, N337, N34);
and AND3 (N342, N341, N279, N279);
nand NAND4 (N343, N335, N111, N309, N245);
nor NOR4 (N344, N339, N269, N241, N7);
nor NOR3 (N345, N332, N127, N164);
and AND3 (N346, N340, N66, N124);
not NOT1 (N347, N345);
xor XOR2 (N348, N336, N208);
xor XOR2 (N349, N338, N96);
nor NOR4 (N350, N342, N304, N89, N177);
xor XOR2 (N351, N320, N191);
buf BUF1 (N352, N348);
or OR4 (N353, N328, N145, N188, N292);
buf BUF1 (N354, N352);
not NOT1 (N355, N347);
and AND4 (N356, N344, N231, N157, N7);
xor XOR2 (N357, N356, N264);
or OR3 (N358, N300, N69, N319);
nor NOR4 (N359, N350, N169, N255, N262);
nand NAND4 (N360, N351, N74, N1, N235);
not NOT1 (N361, N353);
nor NOR2 (N362, N349, N39);
and AND3 (N363, N343, N164, N352);
not NOT1 (N364, N354);
not NOT1 (N365, N362);
not NOT1 (N366, N359);
buf BUF1 (N367, N357);
nor NOR3 (N368, N346, N251, N340);
not NOT1 (N369, N366);
xor XOR2 (N370, N358, N57);
nor NOR3 (N371, N364, N274, N159);
not NOT1 (N372, N369);
or OR2 (N373, N363, N252);
not NOT1 (N374, N368);
buf BUF1 (N375, N365);
not NOT1 (N376, N355);
not NOT1 (N377, N374);
xor XOR2 (N378, N376, N354);
nor NOR2 (N379, N370, N286);
not NOT1 (N380, N375);
nor NOR4 (N381, N372, N268, N298, N218);
buf BUF1 (N382, N380);
xor XOR2 (N383, N378, N373);
not NOT1 (N384, N93);
buf BUF1 (N385, N377);
or OR4 (N386, N367, N200, N15, N84);
not NOT1 (N387, N385);
nor NOR4 (N388, N371, N269, N123, N148);
buf BUF1 (N389, N388);
xor XOR2 (N390, N361, N20);
and AND3 (N391, N381, N199, N342);
buf BUF1 (N392, N386);
buf BUF1 (N393, N360);
nor NOR2 (N394, N384, N351);
or OR4 (N395, N390, N329, N130, N292);
and AND2 (N396, N395, N13);
nor NOR3 (N397, N391, N271, N247);
not NOT1 (N398, N387);
or OR3 (N399, N397, N279, N101);
buf BUF1 (N400, N398);
or OR2 (N401, N399, N116);
buf BUF1 (N402, N383);
nand NAND3 (N403, N400, N169, N111);
nand NAND2 (N404, N394, N258);
buf BUF1 (N405, N403);
not NOT1 (N406, N405);
buf BUF1 (N407, N406);
nand NAND2 (N408, N393, N304);
not NOT1 (N409, N392);
and AND3 (N410, N379, N46, N398);
xor XOR2 (N411, N407, N180);
or OR4 (N412, N411, N2, N84, N198);
not NOT1 (N413, N409);
not NOT1 (N414, N410);
nor NOR3 (N415, N401, N292, N58);
nand NAND2 (N416, N404, N325);
and AND2 (N417, N389, N294);
and AND3 (N418, N417, N231, N58);
buf BUF1 (N419, N408);
nand NAND3 (N420, N415, N84, N222);
xor XOR2 (N421, N418, N367);
not NOT1 (N422, N414);
not NOT1 (N423, N412);
nor NOR3 (N424, N402, N23, N275);
and AND2 (N425, N420, N351);
nor NOR4 (N426, N416, N359, N107, N379);
and AND3 (N427, N422, N102, N372);
and AND2 (N428, N396, N374);
nor NOR4 (N429, N428, N32, N40, N428);
xor XOR2 (N430, N426, N42);
nand NAND2 (N431, N423, N37);
buf BUF1 (N432, N425);
and AND4 (N433, N431, N75, N424, N255);
nand NAND2 (N434, N349, N420);
not NOT1 (N435, N413);
nor NOR3 (N436, N429, N166, N145);
nor NOR2 (N437, N436, N123);
or OR3 (N438, N433, N137, N45);
buf BUF1 (N439, N382);
nor NOR4 (N440, N438, N175, N307, N202);
not NOT1 (N441, N434);
nand NAND3 (N442, N421, N30, N128);
nor NOR3 (N443, N441, N79, N264);
buf BUF1 (N444, N440);
or OR2 (N445, N437, N97);
and AND3 (N446, N427, N346, N416);
or OR2 (N447, N430, N400);
nand NAND3 (N448, N446, N385, N251);
buf BUF1 (N449, N432);
or OR2 (N450, N444, N22);
not NOT1 (N451, N443);
or OR2 (N452, N450, N116);
nand NAND3 (N453, N435, N293, N44);
or OR3 (N454, N419, N114, N325);
xor XOR2 (N455, N448, N4);
not NOT1 (N456, N452);
not NOT1 (N457, N447);
and AND2 (N458, N442, N116);
xor XOR2 (N459, N454, N364);
buf BUF1 (N460, N459);
or OR3 (N461, N445, N167, N24);
not NOT1 (N462, N449);
nand NAND2 (N463, N456, N319);
and AND2 (N464, N439, N47);
and AND2 (N465, N461, N125);
buf BUF1 (N466, N453);
buf BUF1 (N467, N465);
xor XOR2 (N468, N463, N347);
buf BUF1 (N469, N462);
nand NAND3 (N470, N460, N388, N455);
xor XOR2 (N471, N91, N431);
not NOT1 (N472, N470);
or OR3 (N473, N467, N445, N63);
and AND3 (N474, N472, N324, N238);
xor XOR2 (N475, N473, N124);
not NOT1 (N476, N475);
and AND4 (N477, N469, N142, N421, N368);
xor XOR2 (N478, N457, N446);
nand NAND4 (N479, N451, N119, N227, N36);
nor NOR2 (N480, N477, N166);
nand NAND4 (N481, N464, N44, N110, N11);
and AND3 (N482, N458, N139, N214);
nor NOR4 (N483, N476, N328, N37, N298);
and AND2 (N484, N480, N78);
nand NAND3 (N485, N483, N378, N20);
nor NOR4 (N486, N484, N174, N154, N420);
not NOT1 (N487, N485);
nand NAND2 (N488, N482, N16);
or OR2 (N489, N488, N466);
xor XOR2 (N490, N368, N353);
nor NOR3 (N491, N479, N488, N311);
xor XOR2 (N492, N481, N393);
buf BUF1 (N493, N471);
buf BUF1 (N494, N489);
xor XOR2 (N495, N492, N189);
nand NAND2 (N496, N491, N344);
or OR3 (N497, N487, N128, N222);
buf BUF1 (N498, N496);
and AND2 (N499, N494, N34);
not NOT1 (N500, N490);
xor XOR2 (N501, N500, N272);
not NOT1 (N502, N498);
nand NAND4 (N503, N493, N235, N159, N55);
buf BUF1 (N504, N486);
nand NAND2 (N505, N499, N366);
buf BUF1 (N506, N504);
buf BUF1 (N507, N505);
xor XOR2 (N508, N497, N184);
nor NOR2 (N509, N468, N27);
not NOT1 (N510, N501);
xor XOR2 (N511, N478, N264);
not NOT1 (N512, N506);
nand NAND2 (N513, N508, N353);
and AND4 (N514, N509, N123, N393, N269);
nor NOR3 (N515, N502, N464, N493);
nand NAND4 (N516, N474, N293, N364, N404);
or OR3 (N517, N514, N443, N352);
or OR2 (N518, N516, N66);
nor NOR4 (N519, N511, N231, N241, N318);
buf BUF1 (N520, N518);
buf BUF1 (N521, N510);
not NOT1 (N522, N517);
nor NOR2 (N523, N519, N280);
or OR3 (N524, N515, N514, N479);
or OR2 (N525, N520, N364);
not NOT1 (N526, N507);
and AND3 (N527, N524, N405, N256);
or OR4 (N528, N526, N453, N443, N311);
nand NAND4 (N529, N523, N229, N423, N297);
and AND3 (N530, N525, N449, N180);
and AND3 (N531, N529, N399, N254);
or OR3 (N532, N527, N310, N260);
or OR2 (N533, N512, N141);
buf BUF1 (N534, N533);
or OR4 (N535, N513, N450, N489, N10);
nor NOR4 (N536, N535, N28, N485, N388);
or OR3 (N537, N536, N377, N360);
or OR2 (N538, N528, N529);
nor NOR2 (N539, N531, N442);
not NOT1 (N540, N532);
and AND3 (N541, N521, N46, N1);
buf BUF1 (N542, N534);
nor NOR3 (N543, N503, N309, N50);
and AND4 (N544, N495, N284, N378, N315);
nand NAND4 (N545, N541, N429, N183, N43);
nor NOR2 (N546, N539, N503);
not NOT1 (N547, N530);
not NOT1 (N548, N542);
buf BUF1 (N549, N543);
or OR3 (N550, N538, N176, N265);
nor NOR4 (N551, N546, N27, N314, N150);
xor XOR2 (N552, N551, N351);
buf BUF1 (N553, N537);
not NOT1 (N554, N552);
and AND3 (N555, N550, N286, N496);
xor XOR2 (N556, N548, N342);
and AND2 (N557, N522, N184);
not NOT1 (N558, N554);
buf BUF1 (N559, N540);
or OR4 (N560, N557, N452, N96, N428);
xor XOR2 (N561, N547, N267);
buf BUF1 (N562, N560);
not NOT1 (N563, N562);
not NOT1 (N564, N556);
nand NAND2 (N565, N544, N73);
xor XOR2 (N566, N549, N29);
nand NAND3 (N567, N553, N492, N268);
and AND3 (N568, N559, N562, N29);
not NOT1 (N569, N566);
nand NAND4 (N570, N565, N552, N374, N440);
nand NAND3 (N571, N567, N83, N321);
nor NOR2 (N572, N570, N97);
nand NAND4 (N573, N545, N72, N198, N129);
not NOT1 (N574, N573);
nor NOR4 (N575, N555, N297, N240, N548);
or OR2 (N576, N563, N388);
nor NOR2 (N577, N575, N352);
xor XOR2 (N578, N568, N316);
buf BUF1 (N579, N561);
not NOT1 (N580, N577);
or OR3 (N581, N576, N118, N491);
and AND2 (N582, N581, N64);
or OR2 (N583, N574, N303);
and AND4 (N584, N578, N405, N84, N254);
xor XOR2 (N585, N579, N226);
xor XOR2 (N586, N558, N348);
or OR2 (N587, N586, N358);
nor NOR3 (N588, N572, N459, N546);
not NOT1 (N589, N564);
or OR3 (N590, N588, N362, N485);
buf BUF1 (N591, N585);
nor NOR4 (N592, N589, N586, N449, N166);
or OR2 (N593, N571, N275);
not NOT1 (N594, N582);
buf BUF1 (N595, N569);
xor XOR2 (N596, N583, N237);
or OR3 (N597, N590, N419, N442);
buf BUF1 (N598, N584);
not NOT1 (N599, N596);
nor NOR2 (N600, N598, N524);
nor NOR2 (N601, N595, N386);
and AND3 (N602, N592, N89, N25);
xor XOR2 (N603, N599, N349);
or OR2 (N604, N591, N193);
buf BUF1 (N605, N600);
and AND2 (N606, N605, N88);
and AND2 (N607, N603, N26);
nand NAND3 (N608, N604, N328, N349);
nor NOR3 (N609, N607, N167, N304);
not NOT1 (N610, N597);
or OR4 (N611, N610, N220, N86, N255);
or OR3 (N612, N594, N205, N120);
nand NAND3 (N613, N611, N41, N265);
buf BUF1 (N614, N602);
and AND4 (N615, N609, N445, N183, N78);
nand NAND2 (N616, N587, N582);
buf BUF1 (N617, N593);
and AND4 (N618, N617, N213, N91, N399);
and AND3 (N619, N608, N221, N226);
nand NAND4 (N620, N580, N7, N169, N375);
and AND3 (N621, N616, N526, N48);
and AND2 (N622, N613, N464);
and AND3 (N623, N621, N482, N595);
nand NAND2 (N624, N618, N259);
or OR4 (N625, N624, N464, N413, N86);
nand NAND2 (N626, N614, N322);
not NOT1 (N627, N612);
not NOT1 (N628, N627);
or OR4 (N629, N622, N134, N437, N4);
nand NAND4 (N630, N628, N462, N71, N154);
xor XOR2 (N631, N626, N45);
nand NAND3 (N632, N620, N244, N392);
nand NAND3 (N633, N606, N6, N79);
nor NOR2 (N634, N629, N559);
xor XOR2 (N635, N625, N103);
or OR2 (N636, N634, N162);
xor XOR2 (N637, N633, N177);
nand NAND2 (N638, N631, N328);
and AND2 (N639, N632, N94);
and AND3 (N640, N638, N405, N554);
and AND4 (N641, N601, N149, N390, N414);
and AND3 (N642, N640, N185, N592);
or OR2 (N643, N615, N29);
and AND2 (N644, N643, N143);
buf BUF1 (N645, N644);
or OR4 (N646, N623, N342, N122, N410);
not NOT1 (N647, N646);
nor NOR3 (N648, N641, N96, N232);
and AND4 (N649, N619, N586, N256, N573);
xor XOR2 (N650, N647, N155);
not NOT1 (N651, N630);
nor NOR4 (N652, N645, N90, N498, N304);
buf BUF1 (N653, N651);
buf BUF1 (N654, N635);
buf BUF1 (N655, N648);
or OR3 (N656, N636, N36, N131);
buf BUF1 (N657, N639);
and AND2 (N658, N642, N42);
and AND4 (N659, N652, N2, N88, N216);
nor NOR2 (N660, N659, N403);
nor NOR3 (N661, N660, N275, N561);
not NOT1 (N662, N637);
nand NAND4 (N663, N650, N406, N579, N579);
nor NOR4 (N664, N663, N460, N657, N461);
nand NAND2 (N665, N252, N409);
xor XOR2 (N666, N662, N216);
nand NAND2 (N667, N656, N216);
nor NOR2 (N668, N667, N345);
buf BUF1 (N669, N661);
or OR3 (N670, N668, N329, N485);
not NOT1 (N671, N649);
xor XOR2 (N672, N669, N216);
nor NOR4 (N673, N664, N614, N524, N451);
xor XOR2 (N674, N653, N438);
nor NOR2 (N675, N666, N266);
xor XOR2 (N676, N673, N532);
and AND4 (N677, N674, N148, N76, N377);
nand NAND4 (N678, N655, N591, N82, N653);
buf BUF1 (N679, N675);
xor XOR2 (N680, N679, N225);
buf BUF1 (N681, N671);
buf BUF1 (N682, N676);
nand NAND4 (N683, N672, N141, N481, N420);
not NOT1 (N684, N677);
buf BUF1 (N685, N684);
not NOT1 (N686, N680);
or OR2 (N687, N681, N647);
buf BUF1 (N688, N670);
buf BUF1 (N689, N682);
nor NOR4 (N690, N686, N114, N568, N584);
buf BUF1 (N691, N658);
nor NOR2 (N692, N690, N124);
xor XOR2 (N693, N678, N510);
or OR2 (N694, N683, N606);
buf BUF1 (N695, N692);
xor XOR2 (N696, N654, N373);
not NOT1 (N697, N685);
and AND3 (N698, N693, N116, N115);
or OR4 (N699, N689, N185, N42, N238);
and AND4 (N700, N699, N247, N473, N406);
nand NAND3 (N701, N694, N270, N176);
nand NAND2 (N702, N698, N615);
nand NAND4 (N703, N697, N696, N310, N104);
or OR3 (N704, N254, N617, N252);
buf BUF1 (N705, N688);
or OR3 (N706, N691, N347, N9);
xor XOR2 (N707, N706, N317);
and AND2 (N708, N702, N98);
not NOT1 (N709, N701);
not NOT1 (N710, N695);
and AND3 (N711, N705, N181, N477);
xor XOR2 (N712, N704, N641);
nor NOR4 (N713, N665, N381, N514, N477);
not NOT1 (N714, N687);
xor XOR2 (N715, N713, N441);
and AND4 (N716, N711, N353, N16, N240);
buf BUF1 (N717, N714);
nand NAND4 (N718, N715, N518, N204, N435);
nand NAND4 (N719, N717, N642, N370, N473);
nor NOR3 (N720, N710, N639, N317);
and AND3 (N721, N707, N635, N534);
nor NOR4 (N722, N720, N397, N455, N514);
not NOT1 (N723, N722);
buf BUF1 (N724, N716);
nor NOR2 (N725, N721, N141);
not NOT1 (N726, N719);
nor NOR4 (N727, N723, N206, N636, N693);
buf BUF1 (N728, N727);
nand NAND4 (N729, N712, N33, N621, N676);
xor XOR2 (N730, N703, N303);
nor NOR2 (N731, N729, N160);
not NOT1 (N732, N708);
xor XOR2 (N733, N730, N349);
nor NOR3 (N734, N724, N648, N77);
nor NOR3 (N735, N700, N493, N465);
xor XOR2 (N736, N731, N734);
nor NOR3 (N737, N494, N36, N225);
not NOT1 (N738, N737);
nor NOR4 (N739, N725, N213, N654, N589);
xor XOR2 (N740, N726, N23);
xor XOR2 (N741, N739, N493);
or OR2 (N742, N740, N174);
xor XOR2 (N743, N718, N377);
nand NAND3 (N744, N733, N75, N730);
or OR4 (N745, N735, N143, N550, N515);
nor NOR3 (N746, N742, N561, N316);
buf BUF1 (N747, N728);
and AND4 (N748, N745, N549, N673, N407);
nor NOR4 (N749, N744, N436, N367, N687);
not NOT1 (N750, N736);
nor NOR4 (N751, N743, N522, N686, N729);
xor XOR2 (N752, N709, N19);
nor NOR2 (N753, N750, N373);
nand NAND2 (N754, N751, N414);
nor NOR2 (N755, N732, N438);
buf BUF1 (N756, N741);
and AND2 (N757, N754, N103);
nor NOR3 (N758, N749, N621, N574);
buf BUF1 (N759, N748);
nor NOR2 (N760, N757, N602);
not NOT1 (N761, N760);
nor NOR2 (N762, N758, N126);
not NOT1 (N763, N746);
nand NAND2 (N764, N763, N2);
xor XOR2 (N765, N755, N711);
buf BUF1 (N766, N747);
not NOT1 (N767, N766);
or OR4 (N768, N765, N264, N129, N718);
xor XOR2 (N769, N738, N441);
and AND3 (N770, N767, N14, N534);
and AND3 (N771, N756, N268, N50);
and AND4 (N772, N768, N767, N490, N187);
nand NAND2 (N773, N752, N528);
or OR2 (N774, N773, N394);
not NOT1 (N775, N769);
buf BUF1 (N776, N759);
nor NOR2 (N777, N772, N54);
nand NAND4 (N778, N771, N290, N623, N213);
nand NAND3 (N779, N776, N644, N560);
buf BUF1 (N780, N778);
not NOT1 (N781, N775);
and AND4 (N782, N753, N392, N6, N310);
not NOT1 (N783, N764);
nand NAND4 (N784, N761, N350, N731, N24);
buf BUF1 (N785, N774);
buf BUF1 (N786, N785);
nor NOR4 (N787, N784, N533, N110, N418);
or OR3 (N788, N770, N785, N373);
not NOT1 (N789, N783);
buf BUF1 (N790, N781);
buf BUF1 (N791, N762);
nor NOR2 (N792, N789, N88);
xor XOR2 (N793, N792, N776);
or OR3 (N794, N788, N126, N445);
xor XOR2 (N795, N777, N438);
and AND4 (N796, N794, N406, N536, N794);
and AND4 (N797, N780, N598, N402, N60);
nand NAND2 (N798, N790, N187);
not NOT1 (N799, N795);
nand NAND3 (N800, N782, N135, N444);
buf BUF1 (N801, N793);
nand NAND3 (N802, N779, N534, N297);
and AND3 (N803, N791, N5, N6);
xor XOR2 (N804, N799, N553);
buf BUF1 (N805, N801);
buf BUF1 (N806, N804);
and AND3 (N807, N797, N187, N655);
or OR3 (N808, N806, N666, N372);
not NOT1 (N809, N787);
xor XOR2 (N810, N786, N110);
not NOT1 (N811, N796);
not NOT1 (N812, N798);
nor NOR2 (N813, N802, N143);
not NOT1 (N814, N808);
buf BUF1 (N815, N803);
xor XOR2 (N816, N809, N101);
or OR4 (N817, N811, N180, N721, N750);
xor XOR2 (N818, N805, N579);
or OR4 (N819, N818, N454, N480, N487);
xor XOR2 (N820, N814, N17);
nor NOR3 (N821, N820, N561, N379);
nor NOR2 (N822, N800, N92);
or OR2 (N823, N817, N55);
not NOT1 (N824, N815);
buf BUF1 (N825, N812);
nor NOR4 (N826, N810, N394, N550, N103);
buf BUF1 (N827, N822);
or OR3 (N828, N824, N194, N517);
buf BUF1 (N829, N825);
and AND2 (N830, N813, N463);
and AND2 (N831, N819, N625);
xor XOR2 (N832, N827, N726);
buf BUF1 (N833, N823);
not NOT1 (N834, N826);
nor NOR2 (N835, N828, N203);
xor XOR2 (N836, N829, N289);
and AND3 (N837, N832, N606, N223);
buf BUF1 (N838, N835);
xor XOR2 (N839, N833, N699);
nor NOR3 (N840, N837, N104, N835);
buf BUF1 (N841, N807);
and AND2 (N842, N834, N560);
not NOT1 (N843, N821);
nor NOR2 (N844, N841, N574);
nand NAND4 (N845, N843, N367, N824, N233);
nor NOR4 (N846, N816, N586, N316, N570);
or OR3 (N847, N836, N307, N171);
xor XOR2 (N848, N840, N168);
or OR3 (N849, N844, N84, N692);
xor XOR2 (N850, N846, N387);
buf BUF1 (N851, N831);
nor NOR4 (N852, N847, N548, N517, N452);
not NOT1 (N853, N850);
or OR2 (N854, N838, N382);
nor NOR4 (N855, N852, N227, N396, N745);
not NOT1 (N856, N845);
nor NOR4 (N857, N856, N709, N419, N697);
and AND2 (N858, N842, N69);
and AND3 (N859, N858, N780, N301);
and AND2 (N860, N851, N148);
nand NAND3 (N861, N830, N170, N335);
or OR2 (N862, N857, N504);
not NOT1 (N863, N861);
nand NAND4 (N864, N839, N264, N304, N422);
nand NAND4 (N865, N859, N320, N12, N550);
nand NAND4 (N866, N864, N306, N384, N5);
or OR3 (N867, N865, N198, N522);
nand NAND2 (N868, N853, N39);
buf BUF1 (N869, N868);
not NOT1 (N870, N848);
not NOT1 (N871, N863);
or OR3 (N872, N860, N210, N218);
buf BUF1 (N873, N866);
nor NOR4 (N874, N862, N339, N146, N415);
nor NOR4 (N875, N869, N676, N67, N171);
not NOT1 (N876, N855);
and AND2 (N877, N871, N761);
buf BUF1 (N878, N873);
nand NAND4 (N879, N874, N822, N213, N114);
buf BUF1 (N880, N878);
nor NOR2 (N881, N872, N834);
buf BUF1 (N882, N854);
nor NOR4 (N883, N882, N581, N828, N18);
nor NOR4 (N884, N875, N357, N788, N336);
xor XOR2 (N885, N879, N264);
or OR2 (N886, N880, N375);
nor NOR2 (N887, N876, N211);
nor NOR2 (N888, N884, N461);
nor NOR2 (N889, N877, N472);
nand NAND3 (N890, N870, N716, N271);
xor XOR2 (N891, N867, N702);
nand NAND2 (N892, N887, N61);
xor XOR2 (N893, N888, N239);
xor XOR2 (N894, N883, N753);
or OR3 (N895, N889, N126, N248);
xor XOR2 (N896, N886, N715);
nor NOR3 (N897, N892, N61, N276);
nor NOR2 (N898, N897, N468);
or OR2 (N899, N894, N350);
not NOT1 (N900, N891);
xor XOR2 (N901, N890, N191);
not NOT1 (N902, N895);
or OR3 (N903, N900, N838, N113);
buf BUF1 (N904, N849);
nor NOR4 (N905, N899, N894, N53, N641);
and AND2 (N906, N901, N828);
nand NAND2 (N907, N905, N379);
xor XOR2 (N908, N903, N569);
or OR2 (N909, N904, N113);
or OR4 (N910, N908, N872, N674, N280);
xor XOR2 (N911, N910, N900);
nor NOR4 (N912, N893, N782, N771, N847);
xor XOR2 (N913, N912, N509);
buf BUF1 (N914, N896);
not NOT1 (N915, N909);
nand NAND4 (N916, N902, N467, N349, N19);
buf BUF1 (N917, N911);
nor NOR3 (N918, N914, N433, N358);
nand NAND4 (N919, N881, N551, N537, N910);
not NOT1 (N920, N917);
and AND3 (N921, N885, N881, N563);
not NOT1 (N922, N921);
xor XOR2 (N923, N919, N11);
xor XOR2 (N924, N907, N882);
not NOT1 (N925, N920);
nor NOR4 (N926, N918, N359, N294, N345);
and AND3 (N927, N922, N783, N193);
xor XOR2 (N928, N898, N408);
nor NOR2 (N929, N915, N272);
and AND4 (N930, N924, N433, N190, N471);
buf BUF1 (N931, N925);
or OR2 (N932, N926, N230);
nor NOR2 (N933, N927, N594);
and AND4 (N934, N931, N96, N803, N187);
not NOT1 (N935, N929);
buf BUF1 (N936, N932);
xor XOR2 (N937, N936, N319);
not NOT1 (N938, N928);
nor NOR4 (N939, N934, N392, N929, N467);
xor XOR2 (N940, N906, N873);
nand NAND3 (N941, N938, N596, N365);
buf BUF1 (N942, N916);
or OR3 (N943, N930, N737, N558);
xor XOR2 (N944, N935, N883);
or OR2 (N945, N942, N548);
or OR2 (N946, N945, N207);
not NOT1 (N947, N940);
nand NAND3 (N948, N941, N223, N400);
buf BUF1 (N949, N937);
buf BUF1 (N950, N943);
buf BUF1 (N951, N939);
buf BUF1 (N952, N933);
nand NAND3 (N953, N948, N632, N87);
not NOT1 (N954, N944);
buf BUF1 (N955, N913);
nand NAND3 (N956, N950, N438, N32);
or OR3 (N957, N955, N646, N899);
and AND3 (N958, N957, N504, N758);
buf BUF1 (N959, N923);
buf BUF1 (N960, N953);
nand NAND3 (N961, N959, N293, N685);
buf BUF1 (N962, N951);
and AND2 (N963, N960, N869);
buf BUF1 (N964, N956);
not NOT1 (N965, N949);
not NOT1 (N966, N962);
not NOT1 (N967, N952);
not NOT1 (N968, N964);
xor XOR2 (N969, N963, N444);
and AND2 (N970, N966, N708);
or OR2 (N971, N961, N526);
or OR2 (N972, N971, N687);
xor XOR2 (N973, N946, N583);
not NOT1 (N974, N958);
and AND3 (N975, N972, N164, N952);
nand NAND4 (N976, N975, N949, N244, N816);
buf BUF1 (N977, N970);
buf BUF1 (N978, N974);
not NOT1 (N979, N947);
nor NOR2 (N980, N969, N918);
nand NAND2 (N981, N977, N597);
or OR2 (N982, N981, N840);
buf BUF1 (N983, N979);
nor NOR4 (N984, N965, N763, N277, N778);
not NOT1 (N985, N954);
nor NOR3 (N986, N983, N633, N761);
and AND4 (N987, N973, N397, N468, N343);
xor XOR2 (N988, N976, N507);
xor XOR2 (N989, N980, N45);
not NOT1 (N990, N984);
not NOT1 (N991, N990);
nand NAND2 (N992, N987, N603);
and AND2 (N993, N968, N984);
or OR2 (N994, N989, N600);
nand NAND2 (N995, N986, N886);
or OR2 (N996, N985, N211);
nor NOR3 (N997, N988, N859, N701);
not NOT1 (N998, N982);
not NOT1 (N999, N993);
or OR3 (N1000, N978, N699, N947);
nor NOR4 (N1001, N994, N46, N823, N240);
nand NAND4 (N1002, N967, N999, N366, N726);
not NOT1 (N1003, N64);
or OR4 (N1004, N997, N645, N55, N538);
not NOT1 (N1005, N1001);
buf BUF1 (N1006, N1002);
or OR2 (N1007, N1003, N633);
xor XOR2 (N1008, N1007, N123);
nor NOR4 (N1009, N1005, N806, N861, N527);
nand NAND2 (N1010, N998, N740);
xor XOR2 (N1011, N1008, N350);
nand NAND2 (N1012, N995, N617);
xor XOR2 (N1013, N1012, N303);
nor NOR4 (N1014, N1009, N787, N287, N359);
nand NAND2 (N1015, N1011, N204);
nor NOR2 (N1016, N1000, N61);
buf BUF1 (N1017, N1006);
and AND4 (N1018, N1015, N723, N159, N844);
or OR3 (N1019, N991, N261, N391);
not NOT1 (N1020, N1018);
not NOT1 (N1021, N996);
xor XOR2 (N1022, N1010, N651);
xor XOR2 (N1023, N1014, N706);
buf BUF1 (N1024, N1020);
nor NOR2 (N1025, N1023, N743);
nor NOR3 (N1026, N1021, N680, N729);
and AND4 (N1027, N1024, N949, N478, N636);
buf BUF1 (N1028, N1004);
or OR3 (N1029, N1019, N314, N15);
xor XOR2 (N1030, N992, N5);
buf BUF1 (N1031, N1029);
or OR3 (N1032, N1016, N488, N841);
nor NOR3 (N1033, N1026, N47, N26);
xor XOR2 (N1034, N1028, N932);
buf BUF1 (N1035, N1031);
and AND4 (N1036, N1033, N395, N401, N338);
buf BUF1 (N1037, N1034);
and AND2 (N1038, N1035, N136);
nor NOR3 (N1039, N1038, N898, N805);
not NOT1 (N1040, N1030);
nor NOR2 (N1041, N1022, N599);
buf BUF1 (N1042, N1025);
and AND4 (N1043, N1039, N874, N121, N755);
nor NOR2 (N1044, N1037, N805);
nand NAND4 (N1045, N1027, N509, N84, N990);
and AND4 (N1046, N1032, N392, N750, N1026);
or OR3 (N1047, N1046, N773, N21);
xor XOR2 (N1048, N1041, N755);
nor NOR4 (N1049, N1042, N505, N347, N231);
and AND3 (N1050, N1049, N232, N133);
xor XOR2 (N1051, N1047, N621);
buf BUF1 (N1052, N1051);
xor XOR2 (N1053, N1052, N617);
nor NOR2 (N1054, N1050, N769);
nor NOR2 (N1055, N1043, N555);
not NOT1 (N1056, N1017);
or OR4 (N1057, N1056, N590, N210, N794);
or OR4 (N1058, N1044, N154, N856, N564);
and AND3 (N1059, N1057, N370, N199);
buf BUF1 (N1060, N1054);
or OR3 (N1061, N1036, N691, N907);
and AND4 (N1062, N1045, N793, N77, N660);
not NOT1 (N1063, N1061);
xor XOR2 (N1064, N1059, N606);
nand NAND2 (N1065, N1013, N408);
not NOT1 (N1066, N1040);
buf BUF1 (N1067, N1048);
nand NAND4 (N1068, N1066, N937, N975, N866);
not NOT1 (N1069, N1060);
not NOT1 (N1070, N1062);
nand NAND3 (N1071, N1058, N231, N729);
nand NAND2 (N1072, N1055, N428);
buf BUF1 (N1073, N1064);
not NOT1 (N1074, N1071);
and AND2 (N1075, N1070, N493);
and AND2 (N1076, N1075, N346);
buf BUF1 (N1077, N1067);
nand NAND3 (N1078, N1069, N822, N214);
and AND4 (N1079, N1053, N789, N403, N800);
xor XOR2 (N1080, N1076, N867);
nor NOR2 (N1081, N1077, N279);
and AND4 (N1082, N1072, N1019, N155, N167);
or OR3 (N1083, N1078, N271, N281);
or OR2 (N1084, N1074, N825);
or OR3 (N1085, N1063, N793, N481);
buf BUF1 (N1086, N1085);
nand NAND4 (N1087, N1081, N138, N976, N735);
and AND3 (N1088, N1065, N840, N561);
not NOT1 (N1089, N1073);
buf BUF1 (N1090, N1080);
nor NOR4 (N1091, N1088, N548, N140, N201);
nor NOR2 (N1092, N1089, N560);
not NOT1 (N1093, N1087);
not NOT1 (N1094, N1083);
xor XOR2 (N1095, N1082, N1015);
xor XOR2 (N1096, N1068, N1063);
and AND3 (N1097, N1094, N635, N1053);
buf BUF1 (N1098, N1091);
nand NAND4 (N1099, N1097, N871, N906, N1024);
and AND3 (N1100, N1095, N983, N661);
nand NAND2 (N1101, N1090, N1002);
and AND4 (N1102, N1079, N218, N798, N118);
xor XOR2 (N1103, N1084, N257);
not NOT1 (N1104, N1103);
nand NAND2 (N1105, N1104, N92);
nand NAND2 (N1106, N1100, N111);
and AND2 (N1107, N1105, N983);
xor XOR2 (N1108, N1102, N117);
buf BUF1 (N1109, N1086);
xor XOR2 (N1110, N1107, N76);
xor XOR2 (N1111, N1106, N140);
not NOT1 (N1112, N1092);
nand NAND4 (N1113, N1109, N237, N1045, N218);
nand NAND3 (N1114, N1113, N1088, N778);
or OR2 (N1115, N1098, N71);
xor XOR2 (N1116, N1101, N372);
and AND4 (N1117, N1115, N156, N492, N606);
buf BUF1 (N1118, N1093);
buf BUF1 (N1119, N1099);
or OR4 (N1120, N1119, N1079, N1006, N531);
not NOT1 (N1121, N1118);
or OR3 (N1122, N1120, N69, N809);
nand NAND2 (N1123, N1108, N150);
not NOT1 (N1124, N1110);
not NOT1 (N1125, N1116);
xor XOR2 (N1126, N1122, N721);
nor NOR2 (N1127, N1123, N721);
not NOT1 (N1128, N1112);
xor XOR2 (N1129, N1128, N1035);
not NOT1 (N1130, N1111);
nand NAND4 (N1131, N1126, N506, N414, N610);
not NOT1 (N1132, N1125);
nand NAND2 (N1133, N1124, N756);
nor NOR3 (N1134, N1132, N167, N484);
xor XOR2 (N1135, N1096, N1000);
and AND4 (N1136, N1134, N816, N188, N235);
nor NOR4 (N1137, N1130, N212, N418, N409);
or OR3 (N1138, N1131, N954, N111);
and AND2 (N1139, N1117, N157);
or OR3 (N1140, N1127, N273, N907);
xor XOR2 (N1141, N1137, N903);
xor XOR2 (N1142, N1114, N122);
buf BUF1 (N1143, N1133);
nor NOR2 (N1144, N1129, N663);
xor XOR2 (N1145, N1144, N816);
not NOT1 (N1146, N1140);
xor XOR2 (N1147, N1142, N297);
xor XOR2 (N1148, N1121, N419);
nor NOR4 (N1149, N1143, N1088, N483, N26);
xor XOR2 (N1150, N1147, N228);
nand NAND2 (N1151, N1150, N77);
buf BUF1 (N1152, N1141);
and AND2 (N1153, N1148, N267);
xor XOR2 (N1154, N1136, N347);
not NOT1 (N1155, N1145);
nand NAND2 (N1156, N1146, N703);
not NOT1 (N1157, N1155);
xor XOR2 (N1158, N1151, N559);
nor NOR2 (N1159, N1157, N952);
xor XOR2 (N1160, N1152, N388);
nor NOR3 (N1161, N1138, N342, N177);
or OR3 (N1162, N1154, N780, N687);
not NOT1 (N1163, N1161);
or OR3 (N1164, N1156, N1065, N306);
buf BUF1 (N1165, N1164);
and AND2 (N1166, N1158, N1022);
and AND3 (N1167, N1162, N267, N71);
or OR3 (N1168, N1165, N140, N25);
nand NAND2 (N1169, N1135, N848);
xor XOR2 (N1170, N1159, N380);
nor NOR2 (N1171, N1163, N623);
or OR3 (N1172, N1160, N654, N266);
not NOT1 (N1173, N1167);
xor XOR2 (N1174, N1172, N274);
and AND2 (N1175, N1170, N845);
not NOT1 (N1176, N1166);
nand NAND4 (N1177, N1176, N521, N363, N546);
nor NOR4 (N1178, N1173, N219, N913, N985);
and AND2 (N1179, N1149, N975);
or OR3 (N1180, N1169, N1123, N382);
xor XOR2 (N1181, N1139, N254);
nand NAND4 (N1182, N1153, N1002, N966, N519);
or OR2 (N1183, N1178, N688);
not NOT1 (N1184, N1183);
and AND2 (N1185, N1177, N326);
nor NOR2 (N1186, N1175, N252);
and AND2 (N1187, N1171, N370);
not NOT1 (N1188, N1186);
buf BUF1 (N1189, N1184);
buf BUF1 (N1190, N1189);
or OR3 (N1191, N1187, N634, N1173);
nand NAND4 (N1192, N1180, N224, N1085, N798);
and AND3 (N1193, N1182, N691, N249);
not NOT1 (N1194, N1174);
buf BUF1 (N1195, N1181);
and AND2 (N1196, N1192, N356);
or OR4 (N1197, N1185, N128, N174, N473);
or OR4 (N1198, N1168, N109, N545, N595);
nand NAND2 (N1199, N1194, N749);
nand NAND3 (N1200, N1179, N454, N542);
not NOT1 (N1201, N1193);
not NOT1 (N1202, N1197);
not NOT1 (N1203, N1200);
not NOT1 (N1204, N1203);
not NOT1 (N1205, N1198);
or OR4 (N1206, N1188, N528, N943, N299);
not NOT1 (N1207, N1195);
buf BUF1 (N1208, N1191);
xor XOR2 (N1209, N1204, N257);
not NOT1 (N1210, N1209);
or OR3 (N1211, N1199, N336, N700);
nor NOR2 (N1212, N1210, N641);
xor XOR2 (N1213, N1211, N384);
nand NAND2 (N1214, N1208, N708);
or OR2 (N1215, N1207, N398);
nand NAND2 (N1216, N1202, N30);
buf BUF1 (N1217, N1216);
nand NAND3 (N1218, N1215, N471, N485);
xor XOR2 (N1219, N1201, N724);
and AND4 (N1220, N1214, N339, N492, N311);
xor XOR2 (N1221, N1196, N65);
buf BUF1 (N1222, N1205);
buf BUF1 (N1223, N1219);
xor XOR2 (N1224, N1213, N663);
buf BUF1 (N1225, N1224);
not NOT1 (N1226, N1212);
buf BUF1 (N1227, N1222);
and AND3 (N1228, N1190, N323, N428);
nor NOR3 (N1229, N1225, N1032, N687);
and AND3 (N1230, N1227, N67, N135);
and AND4 (N1231, N1217, N524, N1213, N136);
xor XOR2 (N1232, N1226, N7);
nor NOR4 (N1233, N1218, N808, N1122, N1047);
buf BUF1 (N1234, N1223);
buf BUF1 (N1235, N1221);
nand NAND2 (N1236, N1230, N1069);
not NOT1 (N1237, N1206);
or OR2 (N1238, N1220, N683);
or OR4 (N1239, N1231, N210, N1059, N1134);
buf BUF1 (N1240, N1233);
nor NOR3 (N1241, N1234, N112, N541);
nor NOR4 (N1242, N1240, N978, N948, N856);
nand NAND3 (N1243, N1235, N95, N334);
not NOT1 (N1244, N1232);
not NOT1 (N1245, N1243);
or OR3 (N1246, N1239, N1236, N986);
buf BUF1 (N1247, N316);
nor NOR2 (N1248, N1241, N238);
nand NAND4 (N1249, N1244, N1104, N73, N494);
nor NOR3 (N1250, N1245, N558, N644);
nand NAND3 (N1251, N1229, N1186, N247);
and AND2 (N1252, N1248, N81);
not NOT1 (N1253, N1250);
or OR3 (N1254, N1251, N1223, N170);
buf BUF1 (N1255, N1228);
not NOT1 (N1256, N1255);
buf BUF1 (N1257, N1237);
not NOT1 (N1258, N1238);
not NOT1 (N1259, N1252);
nand NAND4 (N1260, N1249, N187, N1175, N1018);
nand NAND2 (N1261, N1246, N833);
and AND3 (N1262, N1253, N552, N385);
buf BUF1 (N1263, N1258);
nor NOR2 (N1264, N1260, N615);
buf BUF1 (N1265, N1247);
buf BUF1 (N1266, N1263);
or OR2 (N1267, N1262, N1054);
or OR3 (N1268, N1261, N726, N1043);
and AND4 (N1269, N1265, N257, N1010, N964);
and AND3 (N1270, N1257, N1220, N687);
nor NOR3 (N1271, N1266, N144, N486);
nand NAND4 (N1272, N1256, N423, N203, N722);
nor NOR4 (N1273, N1271, N3, N597, N728);
not NOT1 (N1274, N1259);
not NOT1 (N1275, N1264);
buf BUF1 (N1276, N1273);
and AND4 (N1277, N1275, N743, N663, N646);
buf BUF1 (N1278, N1277);
not NOT1 (N1279, N1278);
nor NOR3 (N1280, N1274, N580, N890);
nor NOR4 (N1281, N1242, N907, N274, N245);
xor XOR2 (N1282, N1281, N425);
or OR2 (N1283, N1279, N1155);
nand NAND4 (N1284, N1283, N1196, N1219, N792);
nor NOR2 (N1285, N1270, N614);
xor XOR2 (N1286, N1276, N652);
and AND3 (N1287, N1282, N901, N1168);
xor XOR2 (N1288, N1285, N698);
or OR2 (N1289, N1284, N1131);
and AND4 (N1290, N1286, N1051, N76, N588);
and AND2 (N1291, N1287, N637);
not NOT1 (N1292, N1269);
nor NOR4 (N1293, N1272, N1060, N1277, N600);
nand NAND4 (N1294, N1291, N56, N332, N744);
buf BUF1 (N1295, N1280);
and AND2 (N1296, N1288, N841);
or OR4 (N1297, N1254, N98, N152, N938);
or OR2 (N1298, N1292, N1221);
and AND4 (N1299, N1298, N1078, N386, N87);
and AND2 (N1300, N1299, N465);
xor XOR2 (N1301, N1289, N1100);
xor XOR2 (N1302, N1297, N1259);
nand NAND4 (N1303, N1300, N950, N661, N781);
nor NOR2 (N1304, N1268, N695);
not NOT1 (N1305, N1304);
not NOT1 (N1306, N1290);
not NOT1 (N1307, N1301);
and AND4 (N1308, N1307, N713, N456, N542);
and AND4 (N1309, N1267, N641, N952, N858);
xor XOR2 (N1310, N1303, N69);
nor NOR3 (N1311, N1296, N752, N908);
nor NOR3 (N1312, N1308, N19, N743);
buf BUF1 (N1313, N1310);
buf BUF1 (N1314, N1312);
buf BUF1 (N1315, N1305);
or OR3 (N1316, N1309, N1094, N255);
and AND2 (N1317, N1302, N379);
and AND3 (N1318, N1315, N15, N280);
buf BUF1 (N1319, N1295);
xor XOR2 (N1320, N1306, N115);
and AND2 (N1321, N1314, N158);
xor XOR2 (N1322, N1313, N300);
nand NAND3 (N1323, N1318, N291, N481);
nor NOR4 (N1324, N1294, N252, N745, N547);
buf BUF1 (N1325, N1321);
nand NAND4 (N1326, N1323, N1186, N668, N35);
or OR4 (N1327, N1324, N332, N797, N282);
xor XOR2 (N1328, N1319, N662);
buf BUF1 (N1329, N1325);
not NOT1 (N1330, N1327);
nor NOR4 (N1331, N1330, N951, N479, N1201);
not NOT1 (N1332, N1322);
or OR2 (N1333, N1317, N539);
buf BUF1 (N1334, N1333);
nand NAND2 (N1335, N1311, N442);
nor NOR4 (N1336, N1335, N1149, N750, N1068);
nand NAND2 (N1337, N1293, N125);
and AND4 (N1338, N1326, N517, N101, N645);
buf BUF1 (N1339, N1329);
not NOT1 (N1340, N1328);
xor XOR2 (N1341, N1331, N1137);
buf BUF1 (N1342, N1316);
nand NAND4 (N1343, N1337, N556, N1326, N1193);
buf BUF1 (N1344, N1336);
buf BUF1 (N1345, N1332);
or OR2 (N1346, N1320, N1215);
nand NAND2 (N1347, N1344, N512);
or OR4 (N1348, N1339, N450, N938, N584);
and AND2 (N1349, N1338, N968);
or OR3 (N1350, N1348, N1131, N905);
buf BUF1 (N1351, N1340);
xor XOR2 (N1352, N1343, N1027);
xor XOR2 (N1353, N1341, N415);
xor XOR2 (N1354, N1351, N938);
and AND4 (N1355, N1349, N579, N756, N1167);
nand NAND3 (N1356, N1352, N778, N197);
and AND3 (N1357, N1334, N644, N231);
xor XOR2 (N1358, N1357, N76);
xor XOR2 (N1359, N1355, N860);
or OR3 (N1360, N1354, N810, N1129);
buf BUF1 (N1361, N1345);
and AND4 (N1362, N1359, N1308, N648, N915);
nor NOR4 (N1363, N1362, N832, N413, N984);
nor NOR3 (N1364, N1342, N1301, N430);
buf BUF1 (N1365, N1350);
nand NAND4 (N1366, N1360, N1005, N870, N692);
not NOT1 (N1367, N1366);
nand NAND4 (N1368, N1361, N641, N590, N413);
and AND2 (N1369, N1356, N1142);
xor XOR2 (N1370, N1353, N932);
and AND2 (N1371, N1358, N1251);
and AND2 (N1372, N1370, N853);
buf BUF1 (N1373, N1365);
and AND2 (N1374, N1369, N1350);
and AND3 (N1375, N1371, N968, N1119);
nor NOR4 (N1376, N1372, N151, N376, N247);
xor XOR2 (N1377, N1367, N586);
and AND3 (N1378, N1368, N136, N392);
xor XOR2 (N1379, N1347, N850);
nand NAND3 (N1380, N1377, N856, N816);
nor NOR4 (N1381, N1374, N673, N264, N265);
xor XOR2 (N1382, N1375, N359);
or OR2 (N1383, N1346, N663);
nand NAND2 (N1384, N1363, N1231);
nand NAND3 (N1385, N1384, N958, N1180);
and AND2 (N1386, N1383, N313);
not NOT1 (N1387, N1381);
xor XOR2 (N1388, N1379, N1149);
buf BUF1 (N1389, N1388);
and AND4 (N1390, N1386, N1170, N1135, N725);
or OR4 (N1391, N1389, N801, N1066, N1019);
or OR2 (N1392, N1376, N139);
xor XOR2 (N1393, N1390, N437);
or OR2 (N1394, N1385, N1269);
xor XOR2 (N1395, N1382, N574);
nor NOR3 (N1396, N1378, N428, N382);
not NOT1 (N1397, N1392);
nor NOR3 (N1398, N1394, N610, N1382);
nor NOR3 (N1399, N1364, N994, N1376);
xor XOR2 (N1400, N1387, N382);
and AND2 (N1401, N1391, N325);
not NOT1 (N1402, N1397);
and AND2 (N1403, N1398, N1384);
buf BUF1 (N1404, N1393);
nor NOR4 (N1405, N1401, N414, N1228, N340);
nor NOR4 (N1406, N1380, N1196, N1248, N867);
nor NOR4 (N1407, N1396, N1016, N101, N75);
nor NOR4 (N1408, N1402, N1046, N175, N1276);
buf BUF1 (N1409, N1405);
nor NOR2 (N1410, N1406, N171);
nor NOR2 (N1411, N1373, N940);
or OR4 (N1412, N1403, N971, N639, N966);
nand NAND4 (N1413, N1411, N782, N412, N692);
buf BUF1 (N1414, N1404);
buf BUF1 (N1415, N1395);
nor NOR2 (N1416, N1414, N75);
buf BUF1 (N1417, N1400);
and AND4 (N1418, N1413, N593, N988, N748);
nor NOR4 (N1419, N1418, N314, N57, N704);
and AND4 (N1420, N1416, N872, N1139, N481);
or OR2 (N1421, N1412, N402);
nor NOR3 (N1422, N1415, N476, N690);
nand NAND4 (N1423, N1417, N833, N1398, N985);
nand NAND4 (N1424, N1399, N1066, N955, N938);
xor XOR2 (N1425, N1409, N187);
nand NAND4 (N1426, N1407, N1114, N1332, N919);
nand NAND2 (N1427, N1408, N625);
xor XOR2 (N1428, N1410, N85);
xor XOR2 (N1429, N1421, N700);
and AND3 (N1430, N1425, N1109, N660);
and AND2 (N1431, N1429, N971);
or OR3 (N1432, N1431, N824, N358);
and AND2 (N1433, N1430, N619);
nand NAND2 (N1434, N1420, N127);
or OR4 (N1435, N1427, N913, N295, N483);
nand NAND2 (N1436, N1419, N12);
nor NOR2 (N1437, N1433, N72);
xor XOR2 (N1438, N1423, N1391);
not NOT1 (N1439, N1432);
xor XOR2 (N1440, N1435, N670);
not NOT1 (N1441, N1428);
nor NOR2 (N1442, N1434, N1053);
and AND4 (N1443, N1436, N504, N539, N559);
not NOT1 (N1444, N1422);
nor NOR4 (N1445, N1424, N656, N1096, N453);
xor XOR2 (N1446, N1444, N1441);
nor NOR3 (N1447, N1034, N813, N349);
not NOT1 (N1448, N1442);
buf BUF1 (N1449, N1439);
nor NOR3 (N1450, N1445, N625, N722);
xor XOR2 (N1451, N1447, N1153);
nor NOR2 (N1452, N1451, N182);
nor NOR2 (N1453, N1449, N433);
xor XOR2 (N1454, N1438, N1084);
xor XOR2 (N1455, N1446, N922);
xor XOR2 (N1456, N1426, N699);
not NOT1 (N1457, N1443);
nand NAND2 (N1458, N1437, N1254);
nand NAND4 (N1459, N1448, N1025, N1390, N1006);
buf BUF1 (N1460, N1454);
buf BUF1 (N1461, N1452);
nand NAND4 (N1462, N1450, N951, N522, N719);
nand NAND3 (N1463, N1459, N394, N303);
or OR4 (N1464, N1455, N563, N545, N1210);
nand NAND2 (N1465, N1453, N405);
nor NOR3 (N1466, N1458, N245, N1339);
nand NAND2 (N1467, N1463, N457);
nor NOR4 (N1468, N1464, N1109, N217, N627);
nor NOR4 (N1469, N1465, N1099, N1172, N925);
nand NAND4 (N1470, N1468, N790, N699, N1313);
nor NOR2 (N1471, N1469, N585);
nor NOR4 (N1472, N1462, N977, N1331, N1289);
or OR4 (N1473, N1456, N213, N400, N329);
nor NOR3 (N1474, N1471, N535, N316);
not NOT1 (N1475, N1457);
nand NAND3 (N1476, N1460, N1349, N229);
nand NAND2 (N1477, N1472, N29);
xor XOR2 (N1478, N1475, N271);
nand NAND3 (N1479, N1474, N521, N555);
not NOT1 (N1480, N1467);
nor NOR2 (N1481, N1470, N291);
or OR4 (N1482, N1466, N697, N606, N103);
not NOT1 (N1483, N1479);
not NOT1 (N1484, N1477);
buf BUF1 (N1485, N1478);
nor NOR3 (N1486, N1481, N16, N1222);
and AND2 (N1487, N1473, N166);
nor NOR3 (N1488, N1461, N660, N627);
nor NOR2 (N1489, N1440, N1374);
and AND4 (N1490, N1482, N1395, N655, N1244);
or OR3 (N1491, N1483, N1450, N251);
nand NAND2 (N1492, N1484, N45);
nand NAND3 (N1493, N1489, N542, N142);
nor NOR3 (N1494, N1491, N1190, N913);
not NOT1 (N1495, N1488);
nor NOR2 (N1496, N1495, N562);
not NOT1 (N1497, N1486);
not NOT1 (N1498, N1496);
not NOT1 (N1499, N1487);
or OR4 (N1500, N1480, N215, N354, N654);
nor NOR4 (N1501, N1490, N383, N1011, N268);
or OR2 (N1502, N1492, N1364);
not NOT1 (N1503, N1493);
and AND3 (N1504, N1500, N1456, N192);
and AND4 (N1505, N1501, N110, N1370, N1417);
xor XOR2 (N1506, N1494, N384);
and AND3 (N1507, N1502, N461, N1184);
or OR3 (N1508, N1507, N704, N963);
xor XOR2 (N1509, N1506, N1285);
nor NOR2 (N1510, N1508, N466);
and AND4 (N1511, N1509, N724, N878, N411);
and AND4 (N1512, N1499, N232, N1498, N1215);
and AND2 (N1513, N847, N526);
or OR4 (N1514, N1505, N1304, N620, N1017);
and AND3 (N1515, N1510, N1458, N1383);
buf BUF1 (N1516, N1476);
nand NAND3 (N1517, N1503, N908, N265);
buf BUF1 (N1518, N1515);
nor NOR4 (N1519, N1517, N785, N1198, N1033);
xor XOR2 (N1520, N1511, N835);
xor XOR2 (N1521, N1514, N492);
xor XOR2 (N1522, N1521, N518);
nor NOR3 (N1523, N1522, N669, N1370);
xor XOR2 (N1524, N1520, N623);
and AND3 (N1525, N1523, N893, N254);
nand NAND3 (N1526, N1518, N372, N781);
xor XOR2 (N1527, N1516, N236);
or OR4 (N1528, N1527, N85, N96, N1432);
buf BUF1 (N1529, N1519);
nor NOR2 (N1530, N1512, N1115);
or OR2 (N1531, N1524, N1491);
or OR2 (N1532, N1513, N1275);
not NOT1 (N1533, N1497);
not NOT1 (N1534, N1532);
or OR2 (N1535, N1525, N1060);
nor NOR2 (N1536, N1528, N676);
or OR3 (N1537, N1535, N1207, N1018);
and AND3 (N1538, N1530, N567, N1014);
nor NOR3 (N1539, N1531, N1190, N1461);
or OR4 (N1540, N1537, N773, N250, N939);
and AND2 (N1541, N1529, N1130);
not NOT1 (N1542, N1536);
not NOT1 (N1543, N1540);
nand NAND4 (N1544, N1504, N1035, N933, N909);
nand NAND2 (N1545, N1539, N113);
not NOT1 (N1546, N1544);
xor XOR2 (N1547, N1541, N750);
xor XOR2 (N1548, N1542, N229);
xor XOR2 (N1549, N1485, N221);
or OR3 (N1550, N1533, N1246, N1031);
not NOT1 (N1551, N1548);
nor NOR2 (N1552, N1546, N609);
xor XOR2 (N1553, N1545, N953);
or OR3 (N1554, N1550, N1374, N902);
buf BUF1 (N1555, N1551);
nor NOR2 (N1556, N1538, N437);
xor XOR2 (N1557, N1526, N1152);
nor NOR4 (N1558, N1553, N758, N683, N1283);
and AND3 (N1559, N1543, N971, N1179);
buf BUF1 (N1560, N1547);
or OR4 (N1561, N1554, N1405, N427, N1521);
or OR4 (N1562, N1557, N700, N160, N206);
nor NOR2 (N1563, N1561, N1239);
xor XOR2 (N1564, N1558, N731);
or OR4 (N1565, N1555, N115, N1552, N161);
nor NOR2 (N1566, N895, N261);
nor NOR3 (N1567, N1564, N1341, N54);
nor NOR2 (N1568, N1567, N1225);
xor XOR2 (N1569, N1560, N811);
or OR4 (N1570, N1568, N1328, N1545, N103);
nor NOR3 (N1571, N1549, N497, N893);
and AND2 (N1572, N1570, N673);
or OR4 (N1573, N1534, N789, N474, N1041);
or OR3 (N1574, N1556, N1315, N1210);
nand NAND3 (N1575, N1572, N708, N1029);
or OR4 (N1576, N1566, N530, N1266, N223);
nand NAND3 (N1577, N1574, N1146, N236);
not NOT1 (N1578, N1565);
buf BUF1 (N1579, N1577);
nor NOR2 (N1580, N1563, N1148);
nand NAND4 (N1581, N1569, N900, N220, N1573);
buf BUF1 (N1582, N784);
or OR4 (N1583, N1559, N12, N1374, N1496);
buf BUF1 (N1584, N1576);
nand NAND4 (N1585, N1562, N1109, N648, N487);
buf BUF1 (N1586, N1578);
not NOT1 (N1587, N1583);
not NOT1 (N1588, N1571);
nand NAND3 (N1589, N1584, N231, N1423);
nor NOR2 (N1590, N1579, N1112);
buf BUF1 (N1591, N1582);
not NOT1 (N1592, N1586);
buf BUF1 (N1593, N1592);
or OR3 (N1594, N1590, N694, N181);
or OR3 (N1595, N1593, N977, N671);
and AND3 (N1596, N1591, N684, N434);
xor XOR2 (N1597, N1585, N707);
nand NAND3 (N1598, N1594, N1551, N1005);
nor NOR2 (N1599, N1580, N1333);
and AND2 (N1600, N1589, N409);
buf BUF1 (N1601, N1600);
nor NOR4 (N1602, N1581, N831, N192, N812);
xor XOR2 (N1603, N1601, N1343);
not NOT1 (N1604, N1599);
xor XOR2 (N1605, N1603, N849);
xor XOR2 (N1606, N1605, N229);
and AND3 (N1607, N1606, N208, N1311);
nor NOR4 (N1608, N1602, N1453, N1379, N439);
not NOT1 (N1609, N1597);
or OR4 (N1610, N1595, N805, N1406, N903);
buf BUF1 (N1611, N1596);
xor XOR2 (N1612, N1611, N1193);
xor XOR2 (N1613, N1604, N550);
not NOT1 (N1614, N1575);
or OR2 (N1615, N1588, N638);
xor XOR2 (N1616, N1610, N905);
nand NAND4 (N1617, N1616, N1061, N1129, N167);
nor NOR3 (N1618, N1617, N265, N636);
not NOT1 (N1619, N1612);
buf BUF1 (N1620, N1614);
and AND3 (N1621, N1587, N881, N1288);
nand NAND2 (N1622, N1609, N1455);
and AND2 (N1623, N1620, N183);
nand NAND3 (N1624, N1598, N383, N1207);
nor NOR2 (N1625, N1619, N873);
buf BUF1 (N1626, N1608);
not NOT1 (N1627, N1607);
or OR3 (N1628, N1613, N23, N215);
and AND4 (N1629, N1618, N219, N972, N1191);
buf BUF1 (N1630, N1622);
nand NAND2 (N1631, N1629, N918);
buf BUF1 (N1632, N1626);
and AND2 (N1633, N1627, N973);
not NOT1 (N1634, N1633);
or OR4 (N1635, N1634, N1444, N1205, N304);
or OR3 (N1636, N1632, N990, N1200);
buf BUF1 (N1637, N1631);
and AND3 (N1638, N1625, N478, N349);
or OR2 (N1639, N1624, N1620);
or OR3 (N1640, N1615, N1175, N1070);
buf BUF1 (N1641, N1623);
and AND4 (N1642, N1635, N764, N335, N1379);
xor XOR2 (N1643, N1628, N1505);
xor XOR2 (N1644, N1641, N1593);
xor XOR2 (N1645, N1621, N387);
or OR3 (N1646, N1630, N1444, N1044);
or OR3 (N1647, N1637, N1466, N490);
xor XOR2 (N1648, N1638, N1242);
and AND4 (N1649, N1640, N1552, N407, N1067);
not NOT1 (N1650, N1644);
or OR4 (N1651, N1647, N192, N577, N980);
and AND2 (N1652, N1643, N729);
not NOT1 (N1653, N1650);
nand NAND3 (N1654, N1645, N893, N1235);
or OR3 (N1655, N1639, N987, N680);
nand NAND2 (N1656, N1648, N883);
buf BUF1 (N1657, N1656);
nor NOR4 (N1658, N1653, N422, N744, N31);
or OR2 (N1659, N1649, N639);
and AND3 (N1660, N1646, N1605, N1306);
xor XOR2 (N1661, N1636, N1030);
not NOT1 (N1662, N1658);
and AND2 (N1663, N1654, N668);
nor NOR4 (N1664, N1662, N1407, N388, N1655);
nor NOR3 (N1665, N182, N1109, N623);
nand NAND3 (N1666, N1652, N640, N1510);
buf BUF1 (N1667, N1659);
not NOT1 (N1668, N1663);
xor XOR2 (N1669, N1660, N821);
or OR2 (N1670, N1669, N673);
nand NAND2 (N1671, N1670, N964);
and AND2 (N1672, N1661, N980);
buf BUF1 (N1673, N1671);
buf BUF1 (N1674, N1672);
and AND3 (N1675, N1667, N244, N603);
nand NAND4 (N1676, N1666, N1351, N675, N1623);
and AND2 (N1677, N1674, N902);
not NOT1 (N1678, N1651);
nor NOR3 (N1679, N1665, N1079, N246);
nor NOR2 (N1680, N1664, N352);
or OR4 (N1681, N1676, N221, N324, N1180);
nand NAND2 (N1682, N1668, N717);
or OR2 (N1683, N1682, N647);
buf BUF1 (N1684, N1678);
nor NOR3 (N1685, N1679, N961, N834);
xor XOR2 (N1686, N1680, N116);
and AND4 (N1687, N1686, N954, N1208, N1626);
buf BUF1 (N1688, N1687);
xor XOR2 (N1689, N1681, N215);
and AND4 (N1690, N1673, N1113, N1632, N1119);
not NOT1 (N1691, N1675);
or OR3 (N1692, N1677, N186, N1438);
and AND3 (N1693, N1692, N398, N35);
nor NOR4 (N1694, N1688, N104, N940, N1673);
buf BUF1 (N1695, N1690);
nor NOR2 (N1696, N1689, N323);
or OR3 (N1697, N1683, N886, N1467);
nor NOR3 (N1698, N1697, N572, N1467);
nor NOR2 (N1699, N1684, N290);
nand NAND4 (N1700, N1691, N825, N1060, N141);
or OR4 (N1701, N1698, N1019, N717, N977);
xor XOR2 (N1702, N1657, N521);
not NOT1 (N1703, N1694);
nor NOR4 (N1704, N1695, N1547, N1211, N856);
nor NOR4 (N1705, N1685, N923, N170, N878);
and AND4 (N1706, N1693, N1635, N466, N265);
not NOT1 (N1707, N1703);
nand NAND4 (N1708, N1700, N1012, N650, N39);
xor XOR2 (N1709, N1701, N1661);
or OR4 (N1710, N1642, N559, N1472, N461);
xor XOR2 (N1711, N1704, N1381);
xor XOR2 (N1712, N1702, N235);
nor NOR4 (N1713, N1709, N1044, N1297, N611);
and AND4 (N1714, N1713, N1507, N39, N314);
nand NAND4 (N1715, N1708, N306, N86, N935);
not NOT1 (N1716, N1715);
not NOT1 (N1717, N1707);
nand NAND4 (N1718, N1717, N556, N917, N105);
nand NAND3 (N1719, N1714, N97, N668);
nand NAND4 (N1720, N1712, N1207, N192, N804);
or OR2 (N1721, N1706, N1186);
or OR3 (N1722, N1719, N62, N686);
nor NOR3 (N1723, N1722, N611, N1366);
and AND2 (N1724, N1710, N555);
xor XOR2 (N1725, N1699, N1234);
xor XOR2 (N1726, N1721, N1259);
nor NOR4 (N1727, N1716, N468, N471, N1589);
and AND4 (N1728, N1718, N629, N1111, N775);
not NOT1 (N1729, N1724);
xor XOR2 (N1730, N1720, N1256);
not NOT1 (N1731, N1723);
buf BUF1 (N1732, N1731);
xor XOR2 (N1733, N1727, N150);
and AND4 (N1734, N1696, N949, N1299, N844);
nor NOR2 (N1735, N1733, N1613);
buf BUF1 (N1736, N1725);
buf BUF1 (N1737, N1732);
xor XOR2 (N1738, N1734, N1724);
not NOT1 (N1739, N1736);
or OR2 (N1740, N1738, N867);
and AND4 (N1741, N1729, N335, N1344, N1077);
or OR4 (N1742, N1730, N677, N48, N1558);
xor XOR2 (N1743, N1739, N1700);
xor XOR2 (N1744, N1742, N984);
and AND3 (N1745, N1711, N122, N119);
or OR2 (N1746, N1705, N386);
xor XOR2 (N1747, N1746, N846);
xor XOR2 (N1748, N1741, N856);
nor NOR3 (N1749, N1745, N855, N1558);
buf BUF1 (N1750, N1728);
xor XOR2 (N1751, N1747, N1659);
or OR3 (N1752, N1751, N1216, N1131);
or OR3 (N1753, N1740, N139, N337);
and AND3 (N1754, N1752, N788, N664);
xor XOR2 (N1755, N1744, N135);
nand NAND4 (N1756, N1726, N563, N803, N165);
and AND2 (N1757, N1748, N1449);
nand NAND3 (N1758, N1754, N8, N5);
not NOT1 (N1759, N1737);
or OR2 (N1760, N1735, N931);
and AND3 (N1761, N1753, N1172, N548);
or OR3 (N1762, N1757, N606, N1021);
and AND4 (N1763, N1762, N415, N827, N254);
not NOT1 (N1764, N1750);
nor NOR2 (N1765, N1755, N728);
not NOT1 (N1766, N1760);
or OR2 (N1767, N1758, N1759);
nor NOR2 (N1768, N391, N155);
nand NAND3 (N1769, N1764, N494, N1209);
nand NAND4 (N1770, N1768, N372, N1472, N1305);
xor XOR2 (N1771, N1769, N440);
not NOT1 (N1772, N1756);
or OR4 (N1773, N1763, N109, N1503, N1083);
nor NOR4 (N1774, N1767, N98, N735, N129);
buf BUF1 (N1775, N1772);
not NOT1 (N1776, N1770);
not NOT1 (N1777, N1761);
or OR2 (N1778, N1776, N108);
xor XOR2 (N1779, N1771, N464);
nand NAND2 (N1780, N1777, N148);
buf BUF1 (N1781, N1774);
nand NAND3 (N1782, N1779, N1604, N1494);
and AND3 (N1783, N1782, N320, N565);
not NOT1 (N1784, N1766);
and AND4 (N1785, N1783, N106, N668, N21);
and AND2 (N1786, N1773, N502);
buf BUF1 (N1787, N1749);
and AND2 (N1788, N1786, N534);
nand NAND2 (N1789, N1784, N456);
not NOT1 (N1790, N1787);
not NOT1 (N1791, N1778);
buf BUF1 (N1792, N1781);
xor XOR2 (N1793, N1765, N1354);
not NOT1 (N1794, N1788);
and AND3 (N1795, N1789, N72, N155);
or OR2 (N1796, N1794, N1460);
not NOT1 (N1797, N1780);
or OR4 (N1798, N1775, N1289, N1773, N1613);
xor XOR2 (N1799, N1785, N91);
and AND4 (N1800, N1796, N300, N1464, N386);
buf BUF1 (N1801, N1798);
xor XOR2 (N1802, N1800, N230);
and AND3 (N1803, N1797, N1239, N559);
xor XOR2 (N1804, N1795, N857);
xor XOR2 (N1805, N1801, N5);
and AND3 (N1806, N1802, N1380, N1470);
xor XOR2 (N1807, N1806, N226);
xor XOR2 (N1808, N1805, N1766);
nand NAND3 (N1809, N1792, N1000, N1462);
xor XOR2 (N1810, N1804, N1569);
nand NAND3 (N1811, N1807, N1738, N199);
or OR3 (N1812, N1791, N109, N1242);
not NOT1 (N1813, N1809);
or OR4 (N1814, N1743, N208, N1642, N1666);
nor NOR3 (N1815, N1808, N1104, N318);
and AND4 (N1816, N1799, N1766, N1460, N1100);
or OR4 (N1817, N1816, N580, N458, N1478);
not NOT1 (N1818, N1812);
not NOT1 (N1819, N1810);
nand NAND2 (N1820, N1790, N1761);
nand NAND4 (N1821, N1814, N550, N475, N1442);
not NOT1 (N1822, N1803);
not NOT1 (N1823, N1820);
buf BUF1 (N1824, N1821);
or OR3 (N1825, N1818, N1011, N459);
or OR2 (N1826, N1813, N374);
nor NOR3 (N1827, N1815, N1637, N316);
not NOT1 (N1828, N1811);
or OR4 (N1829, N1793, N1640, N127, N1378);
and AND3 (N1830, N1823, N789, N735);
buf BUF1 (N1831, N1819);
not NOT1 (N1832, N1824);
nor NOR2 (N1833, N1830, N1258);
buf BUF1 (N1834, N1829);
nand NAND3 (N1835, N1832, N1366, N1638);
nor NOR2 (N1836, N1833, N1539);
buf BUF1 (N1837, N1828);
nand NAND4 (N1838, N1837, N1132, N1180, N1);
and AND3 (N1839, N1825, N1161, N510);
or OR3 (N1840, N1827, N175, N1491);
or OR3 (N1841, N1831, N920, N1834);
buf BUF1 (N1842, N1566);
or OR2 (N1843, N1817, N314);
buf BUF1 (N1844, N1822);
nor NOR2 (N1845, N1838, N795);
not NOT1 (N1846, N1840);
nand NAND2 (N1847, N1841, N1092);
nor NOR3 (N1848, N1844, N387, N293);
or OR3 (N1849, N1842, N77, N1099);
nor NOR3 (N1850, N1845, N125, N949);
or OR4 (N1851, N1839, N1032, N1651, N1222);
nand NAND4 (N1852, N1835, N1380, N516, N1589);
nor NOR2 (N1853, N1848, N1465);
buf BUF1 (N1854, N1849);
and AND3 (N1855, N1846, N1404, N894);
xor XOR2 (N1856, N1843, N187);
nand NAND3 (N1857, N1847, N728, N1191);
or OR4 (N1858, N1853, N234, N563, N1386);
and AND4 (N1859, N1826, N858, N71, N1525);
xor XOR2 (N1860, N1854, N1032);
not NOT1 (N1861, N1855);
buf BUF1 (N1862, N1856);
nand NAND3 (N1863, N1857, N1552, N343);
not NOT1 (N1864, N1860);
not NOT1 (N1865, N1858);
buf BUF1 (N1866, N1862);
or OR4 (N1867, N1859, N157, N1201, N1339);
nand NAND4 (N1868, N1863, N954, N1247, N449);
and AND2 (N1869, N1861, N517);
nand NAND3 (N1870, N1836, N1698, N1699);
and AND2 (N1871, N1866, N1139);
not NOT1 (N1872, N1851);
and AND2 (N1873, N1865, N298);
nor NOR4 (N1874, N1852, N716, N1580, N1808);
or OR3 (N1875, N1868, N581, N1440);
nor NOR2 (N1876, N1850, N1873);
buf BUF1 (N1877, N406);
nor NOR3 (N1878, N1872, N21, N549);
xor XOR2 (N1879, N1870, N367);
not NOT1 (N1880, N1875);
nand NAND4 (N1881, N1871, N267, N1483, N852);
not NOT1 (N1882, N1877);
xor XOR2 (N1883, N1869, N1446);
not NOT1 (N1884, N1881);
nand NAND2 (N1885, N1874, N576);
xor XOR2 (N1886, N1867, N1694);
nor NOR2 (N1887, N1882, N1442);
buf BUF1 (N1888, N1879);
or OR3 (N1889, N1885, N1690, N1144);
and AND2 (N1890, N1889, N792);
xor XOR2 (N1891, N1880, N1092);
nor NOR3 (N1892, N1888, N31, N343);
buf BUF1 (N1893, N1890);
or OR2 (N1894, N1883, N61);
nand NAND3 (N1895, N1886, N795, N1844);
or OR2 (N1896, N1876, N1583);
buf BUF1 (N1897, N1891);
buf BUF1 (N1898, N1896);
and AND4 (N1899, N1884, N716, N1704, N479);
xor XOR2 (N1900, N1887, N534);
nand NAND4 (N1901, N1899, N334, N1097, N1142);
not NOT1 (N1902, N1892);
not NOT1 (N1903, N1894);
not NOT1 (N1904, N1901);
nor NOR2 (N1905, N1897, N548);
or OR2 (N1906, N1902, N1834);
nand NAND2 (N1907, N1903, N638);
not NOT1 (N1908, N1893);
not NOT1 (N1909, N1900);
buf BUF1 (N1910, N1905);
or OR2 (N1911, N1909, N482);
xor XOR2 (N1912, N1898, N560);
xor XOR2 (N1913, N1908, N31);
buf BUF1 (N1914, N1864);
or OR3 (N1915, N1895, N1339, N1880);
xor XOR2 (N1916, N1911, N235);
buf BUF1 (N1917, N1913);
buf BUF1 (N1918, N1915);
not NOT1 (N1919, N1878);
nor NOR2 (N1920, N1912, N1429);
xor XOR2 (N1921, N1907, N1016);
or OR2 (N1922, N1904, N1190);
xor XOR2 (N1923, N1906, N369);
nor NOR4 (N1924, N1910, N519, N218, N946);
nor NOR2 (N1925, N1914, N1534);
nor NOR3 (N1926, N1921, N95, N1840);
and AND3 (N1927, N1920, N1242, N1842);
or OR3 (N1928, N1918, N1730, N1692);
and AND3 (N1929, N1916, N1251, N1464);
or OR4 (N1930, N1917, N783, N277, N296);
xor XOR2 (N1931, N1929, N731);
or OR2 (N1932, N1928, N550);
or OR4 (N1933, N1926, N1253, N1898, N1150);
nand NAND3 (N1934, N1924, N1091, N537);
buf BUF1 (N1935, N1922);
nor NOR3 (N1936, N1935, N877, N624);
and AND3 (N1937, N1933, N1592, N1659);
nand NAND2 (N1938, N1934, N701);
or OR3 (N1939, N1938, N545, N1254);
nand NAND3 (N1940, N1927, N240, N1367);
or OR4 (N1941, N1930, N215, N566, N1839);
not NOT1 (N1942, N1932);
not NOT1 (N1943, N1939);
or OR2 (N1944, N1937, N1359);
or OR2 (N1945, N1944, N1278);
nor NOR3 (N1946, N1936, N585, N1878);
xor XOR2 (N1947, N1946, N1766);
and AND2 (N1948, N1943, N1755);
buf BUF1 (N1949, N1947);
nor NOR4 (N1950, N1945, N1117, N1709, N908);
nand NAND2 (N1951, N1931, N287);
xor XOR2 (N1952, N1942, N1828);
and AND2 (N1953, N1925, N10);
nand NAND4 (N1954, N1941, N1392, N1907, N526);
or OR3 (N1955, N1949, N1723, N393);
xor XOR2 (N1956, N1948, N1892);
xor XOR2 (N1957, N1923, N768);
not NOT1 (N1958, N1957);
nand NAND4 (N1959, N1951, N634, N228, N1463);
xor XOR2 (N1960, N1956, N111);
nor NOR4 (N1961, N1919, N1057, N402, N1081);
nor NOR4 (N1962, N1954, N1773, N1833, N1430);
buf BUF1 (N1963, N1959);
nor NOR4 (N1964, N1958, N24, N964, N844);
not NOT1 (N1965, N1955);
or OR3 (N1966, N1963, N1086, N1108);
nand NAND4 (N1967, N1962, N149, N1229, N1749);
buf BUF1 (N1968, N1964);
buf BUF1 (N1969, N1965);
buf BUF1 (N1970, N1967);
not NOT1 (N1971, N1966);
or OR2 (N1972, N1971, N1257);
or OR3 (N1973, N1960, N1206, N25);
and AND3 (N1974, N1953, N608, N174);
xor XOR2 (N1975, N1961, N579);
nand NAND3 (N1976, N1972, N1255, N1485);
nand NAND2 (N1977, N1975, N1308);
or OR2 (N1978, N1970, N1790);
nor NOR4 (N1979, N1969, N695, N1767, N1115);
nor NOR4 (N1980, N1940, N1944, N1946, N301);
buf BUF1 (N1981, N1977);
not NOT1 (N1982, N1981);
nand NAND4 (N1983, N1973, N1963, N1363, N1657);
nand NAND2 (N1984, N1983, N1730);
and AND2 (N1985, N1978, N520);
not NOT1 (N1986, N1968);
nand NAND2 (N1987, N1974, N438);
not NOT1 (N1988, N1979);
and AND2 (N1989, N1988, N17);
and AND2 (N1990, N1950, N1484);
and AND4 (N1991, N1986, N1428, N19, N1467);
buf BUF1 (N1992, N1987);
or OR2 (N1993, N1991, N1076);
not NOT1 (N1994, N1976);
nand NAND3 (N1995, N1994, N142, N1522);
nor NOR3 (N1996, N1990, N996, N1041);
xor XOR2 (N1997, N1995, N1643);
buf BUF1 (N1998, N1996);
or OR3 (N1999, N1980, N1485, N1803);
nand NAND3 (N2000, N1984, N1663, N1425);
and AND4 (N2001, N1985, N1683, N928, N923);
nand NAND4 (N2002, N1989, N1504, N953, N579);
or OR3 (N2003, N2000, N1824, N1469);
and AND2 (N2004, N1999, N1515);
xor XOR2 (N2005, N1982, N161);
and AND3 (N2006, N1992, N925, N58);
buf BUF1 (N2007, N1998);
nand NAND4 (N2008, N2001, N1238, N985, N228);
not NOT1 (N2009, N1952);
nand NAND3 (N2010, N2003, N2003, N52);
xor XOR2 (N2011, N2006, N1604);
xor XOR2 (N2012, N2002, N1477);
nor NOR3 (N2013, N2007, N90, N488);
or OR4 (N2014, N1997, N1386, N184, N1827);
or OR4 (N2015, N2005, N855, N1005, N1009);
not NOT1 (N2016, N2011);
nand NAND4 (N2017, N2015, N1529, N1282, N295);
and AND2 (N2018, N2012, N1751);
nor NOR4 (N2019, N2014, N1628, N2013, N738);
or OR2 (N2020, N31, N1354);
xor XOR2 (N2021, N2016, N479);
buf BUF1 (N2022, N2008);
or OR4 (N2023, N2009, N1551, N532, N642);
or OR4 (N2024, N2017, N1436, N599, N686);
and AND4 (N2025, N2024, N741, N676, N1954);
nand NAND3 (N2026, N1993, N1585, N2006);
and AND3 (N2027, N2021, N835, N1236);
nor NOR4 (N2028, N2027, N874, N139, N1357);
or OR4 (N2029, N2004, N1878, N1611, N685);
buf BUF1 (N2030, N2010);
or OR3 (N2031, N2025, N1262, N1886);
nor NOR4 (N2032, N2019, N986, N1640, N1974);
nor NOR3 (N2033, N2032, N369, N1351);
nand NAND3 (N2034, N2028, N1276, N1874);
nor NOR2 (N2035, N2020, N798);
nor NOR4 (N2036, N2030, N1310, N1467, N859);
xor XOR2 (N2037, N2023, N1533);
and AND4 (N2038, N2026, N161, N1525, N1947);
buf BUF1 (N2039, N2031);
not NOT1 (N2040, N2022);
or OR3 (N2041, N2034, N1465, N861);
not NOT1 (N2042, N2037);
nand NAND3 (N2043, N2035, N2026, N1597);
not NOT1 (N2044, N2029);
nor NOR4 (N2045, N2038, N486, N1224, N1486);
nor NOR2 (N2046, N2044, N868);
not NOT1 (N2047, N2041);
and AND4 (N2048, N2042, N640, N1240, N412);
nand NAND3 (N2049, N2036, N1127, N1924);
xor XOR2 (N2050, N2049, N504);
nor NOR4 (N2051, N2050, N977, N267, N189);
nand NAND2 (N2052, N2018, N257);
xor XOR2 (N2053, N2052, N701);
nor NOR4 (N2054, N2039, N448, N445, N1491);
or OR3 (N2055, N2045, N583, N636);
xor XOR2 (N2056, N2054, N1102);
nor NOR3 (N2057, N2051, N167, N582);
nand NAND3 (N2058, N2040, N1250, N557);
or OR3 (N2059, N2047, N625, N1268);
or OR4 (N2060, N2058, N487, N1333, N731);
and AND2 (N2061, N2057, N1695);
nor NOR4 (N2062, N2056, N1635, N905, N71);
xor XOR2 (N2063, N2062, N8);
buf BUF1 (N2064, N2059);
xor XOR2 (N2065, N2055, N925);
not NOT1 (N2066, N2048);
buf BUF1 (N2067, N2043);
and AND2 (N2068, N2063, N656);
and AND4 (N2069, N2064, N519, N867, N515);
xor XOR2 (N2070, N2046, N500);
nand NAND4 (N2071, N2067, N1576, N1886, N1718);
and AND2 (N2072, N2066, N549);
nor NOR3 (N2073, N2070, N621, N1421);
xor XOR2 (N2074, N2072, N1693);
or OR3 (N2075, N2033, N964, N199);
buf BUF1 (N2076, N2071);
or OR3 (N2077, N2074, N473, N974);
nand NAND2 (N2078, N2073, N782);
xor XOR2 (N2079, N2069, N1958);
or OR3 (N2080, N2078, N1317, N1794);
xor XOR2 (N2081, N2065, N1538);
xor XOR2 (N2082, N2068, N722);
nand NAND3 (N2083, N2076, N1805, N948);
buf BUF1 (N2084, N2083);
not NOT1 (N2085, N2060);
buf BUF1 (N2086, N2079);
nand NAND3 (N2087, N2077, N1428, N588);
or OR2 (N2088, N2075, N886);
or OR4 (N2089, N2087, N2064, N97, N251);
or OR4 (N2090, N2086, N1078, N1436, N740);
nor NOR2 (N2091, N2090, N1828);
xor XOR2 (N2092, N2085, N131);
xor XOR2 (N2093, N2082, N126);
nand NAND3 (N2094, N2091, N251, N10);
and AND3 (N2095, N2089, N290, N87);
not NOT1 (N2096, N2094);
and AND2 (N2097, N2092, N1947);
xor XOR2 (N2098, N2080, N1144);
or OR3 (N2099, N2093, N1002, N1445);
or OR3 (N2100, N2098, N1420, N1205);
and AND2 (N2101, N2100, N737);
buf BUF1 (N2102, N2099);
not NOT1 (N2103, N2084);
or OR3 (N2104, N2103, N549, N898);
not NOT1 (N2105, N2081);
or OR2 (N2106, N2096, N955);
not NOT1 (N2107, N2061);
or OR4 (N2108, N2104, N1782, N797, N818);
nor NOR4 (N2109, N2105, N1329, N1298, N1938);
nor NOR4 (N2110, N2088, N1600, N647, N340);
nor NOR3 (N2111, N2097, N1571, N1954);
not NOT1 (N2112, N2109);
xor XOR2 (N2113, N2095, N1944);
not NOT1 (N2114, N2102);
buf BUF1 (N2115, N2053);
nor NOR4 (N2116, N2110, N2058, N769, N1085);
nand NAND2 (N2117, N2111, N1000);
or OR2 (N2118, N2115, N1803);
and AND2 (N2119, N2113, N1335);
nor NOR3 (N2120, N2101, N1109, N1040);
nand NAND4 (N2121, N2114, N1608, N35, N981);
nand NAND3 (N2122, N2119, N640, N2038);
buf BUF1 (N2123, N2118);
and AND3 (N2124, N2117, N2110, N1474);
buf BUF1 (N2125, N2108);
not NOT1 (N2126, N2112);
xor XOR2 (N2127, N2106, N1540);
nand NAND4 (N2128, N2107, N33, N1736, N1800);
nand NAND3 (N2129, N2116, N399, N1038);
or OR4 (N2130, N2127, N1509, N575, N730);
not NOT1 (N2131, N2124);
nor NOR3 (N2132, N2129, N1977, N319);
xor XOR2 (N2133, N2122, N631);
not NOT1 (N2134, N2131);
xor XOR2 (N2135, N2133, N335);
not NOT1 (N2136, N2135);
and AND3 (N2137, N2121, N7, N2017);
buf BUF1 (N2138, N2137);
not NOT1 (N2139, N2123);
not NOT1 (N2140, N2128);
xor XOR2 (N2141, N2132, N1444);
not NOT1 (N2142, N2126);
or OR4 (N2143, N2141, N1813, N993, N888);
nor NOR4 (N2144, N2140, N51, N26, N1609);
xor XOR2 (N2145, N2142, N639);
xor XOR2 (N2146, N2134, N1587);
xor XOR2 (N2147, N2130, N1546);
buf BUF1 (N2148, N2136);
buf BUF1 (N2149, N2125);
nor NOR3 (N2150, N2143, N244, N1720);
nand NAND3 (N2151, N2144, N399, N63);
nor NOR2 (N2152, N2120, N249);
xor XOR2 (N2153, N2152, N474);
and AND2 (N2154, N2150, N77);
and AND4 (N2155, N2153, N1637, N1352, N539);
not NOT1 (N2156, N2138);
xor XOR2 (N2157, N2155, N1987);
not NOT1 (N2158, N2157);
buf BUF1 (N2159, N2154);
buf BUF1 (N2160, N2151);
and AND4 (N2161, N2159, N1241, N150, N31);
buf BUF1 (N2162, N2147);
not NOT1 (N2163, N2160);
xor XOR2 (N2164, N2149, N1365);
nor NOR2 (N2165, N2163, N1707);
and AND4 (N2166, N2139, N1746, N1516, N1245);
not NOT1 (N2167, N2148);
nand NAND3 (N2168, N2167, N1060, N2053);
xor XOR2 (N2169, N2161, N1600);
xor XOR2 (N2170, N2145, N1193);
not NOT1 (N2171, N2169);
nand NAND3 (N2172, N2171, N1781, N1185);
nand NAND2 (N2173, N2166, N768);
xor XOR2 (N2174, N2170, N106);
xor XOR2 (N2175, N2164, N1430);
not NOT1 (N2176, N2162);
nor NOR2 (N2177, N2174, N2171);
nand NAND2 (N2178, N2176, N665);
xor XOR2 (N2179, N2146, N1379);
nor NOR2 (N2180, N2172, N133);
or OR2 (N2181, N2179, N2116);
or OR4 (N2182, N2175, N2134, N517, N290);
and AND2 (N2183, N2168, N1807);
not NOT1 (N2184, N2182);
xor XOR2 (N2185, N2183, N1868);
nand NAND4 (N2186, N2185, N1927, N1948, N952);
or OR4 (N2187, N2178, N87, N470, N1009);
buf BUF1 (N2188, N2165);
or OR4 (N2189, N2184, N1904, N983, N1817);
nand NAND2 (N2190, N2177, N788);
and AND3 (N2191, N2156, N537, N1765);
xor XOR2 (N2192, N2188, N2090);
nand NAND3 (N2193, N2187, N1295, N1158);
not NOT1 (N2194, N2192);
and AND4 (N2195, N2158, N2098, N978, N1295);
nor NOR3 (N2196, N2181, N1925, N266);
or OR4 (N2197, N2180, N200, N200, N1656);
nor NOR2 (N2198, N2196, N511);
xor XOR2 (N2199, N2189, N912);
or OR4 (N2200, N2194, N1627, N1714, N1182);
and AND2 (N2201, N2195, N2046);
nor NOR4 (N2202, N2186, N1726, N177, N1353);
and AND4 (N2203, N2197, N1217, N397, N1214);
and AND2 (N2204, N2193, N2065);
nor NOR4 (N2205, N2173, N1038, N368, N171);
or OR4 (N2206, N2199, N2115, N1431, N621);
nor NOR2 (N2207, N2190, N1086);
and AND4 (N2208, N2207, N1080, N1330, N523);
xor XOR2 (N2209, N2203, N1706);
and AND3 (N2210, N2209, N603, N485);
nand NAND3 (N2211, N2204, N2004, N1772);
and AND2 (N2212, N2201, N1336);
or OR3 (N2213, N2205, N628, N1820);
not NOT1 (N2214, N2211);
nand NAND4 (N2215, N2206, N1315, N160, N1829);
nand NAND3 (N2216, N2212, N888, N1379);
nor NOR3 (N2217, N2216, N2141, N1316);
buf BUF1 (N2218, N2213);
not NOT1 (N2219, N2217);
nand NAND4 (N2220, N2218, N1388, N1504, N1562);
or OR4 (N2221, N2202, N232, N242, N196);
nor NOR3 (N2222, N2221, N718, N168);
or OR2 (N2223, N2191, N1091);
nand NAND2 (N2224, N2208, N517);
or OR2 (N2225, N2219, N1383);
buf BUF1 (N2226, N2198);
nand NAND2 (N2227, N2223, N736);
or OR4 (N2228, N2226, N1833, N228, N1856);
xor XOR2 (N2229, N2228, N1267);
not NOT1 (N2230, N2227);
xor XOR2 (N2231, N2224, N2113);
and AND3 (N2232, N2229, N1216, N836);
or OR4 (N2233, N2210, N1762, N1022, N1152);
nand NAND2 (N2234, N2200, N1032);
or OR4 (N2235, N2233, N629, N1404, N1127);
buf BUF1 (N2236, N2232);
buf BUF1 (N2237, N2214);
nor NOR3 (N2238, N2222, N1030, N560);
and AND3 (N2239, N2237, N737, N88);
nor NOR2 (N2240, N2239, N1880);
and AND4 (N2241, N2230, N316, N2079, N428);
nor NOR2 (N2242, N2241, N549);
xor XOR2 (N2243, N2215, N1338);
and AND2 (N2244, N2220, N781);
buf BUF1 (N2245, N2240);
nand NAND3 (N2246, N2238, N30, N155);
nand NAND3 (N2247, N2236, N1331, N1964);
not NOT1 (N2248, N2235);
not NOT1 (N2249, N2247);
nand NAND2 (N2250, N2249, N350);
nor NOR2 (N2251, N2243, N747);
or OR4 (N2252, N2244, N1422, N1363, N638);
nand NAND3 (N2253, N2252, N1402, N532);
or OR4 (N2254, N2234, N767, N273, N1583);
buf BUF1 (N2255, N2245);
xor XOR2 (N2256, N2253, N1282);
nor NOR3 (N2257, N2242, N984, N740);
nand NAND4 (N2258, N2257, N711, N2034, N1756);
nand NAND3 (N2259, N2256, N1519, N2009);
not NOT1 (N2260, N2225);
and AND3 (N2261, N2246, N489, N1256);
xor XOR2 (N2262, N2261, N1969);
nand NAND2 (N2263, N2250, N1614);
or OR3 (N2264, N2231, N764, N1047);
buf BUF1 (N2265, N2264);
buf BUF1 (N2266, N2258);
nor NOR2 (N2267, N2266, N2034);
and AND3 (N2268, N2251, N1755, N1236);
and AND4 (N2269, N2267, N755, N739, N1135);
nor NOR3 (N2270, N2259, N1179, N627);
xor XOR2 (N2271, N2248, N1283);
or OR2 (N2272, N2271, N710);
or OR4 (N2273, N2255, N2186, N2165, N1261);
not NOT1 (N2274, N2268);
nor NOR4 (N2275, N2274, N2252, N1305, N1883);
and AND2 (N2276, N2272, N1024);
nor NOR2 (N2277, N2262, N562);
xor XOR2 (N2278, N2273, N560);
xor XOR2 (N2279, N2276, N758);
nand NAND4 (N2280, N2270, N2148, N1881, N834);
buf BUF1 (N2281, N2265);
not NOT1 (N2282, N2278);
not NOT1 (N2283, N2277);
xor XOR2 (N2284, N2269, N188);
and AND3 (N2285, N2281, N241, N137);
and AND2 (N2286, N2284, N353);
and AND3 (N2287, N2263, N2152, N801);
nand NAND3 (N2288, N2285, N1814, N1782);
not NOT1 (N2289, N2283);
or OR3 (N2290, N2286, N1537, N571);
nand NAND2 (N2291, N2260, N640);
and AND4 (N2292, N2288, N425, N1133, N965);
nor NOR4 (N2293, N2282, N484, N1047, N832);
not NOT1 (N2294, N2279);
or OR2 (N2295, N2291, N2018);
buf BUF1 (N2296, N2292);
nor NOR3 (N2297, N2275, N1103, N231);
nor NOR2 (N2298, N2297, N1099);
and AND3 (N2299, N2296, N1973, N1907);
not NOT1 (N2300, N2254);
not NOT1 (N2301, N2293);
buf BUF1 (N2302, N2298);
xor XOR2 (N2303, N2295, N1396);
nand NAND2 (N2304, N2294, N169);
or OR4 (N2305, N2290, N1738, N1403, N622);
nand NAND4 (N2306, N2303, N1990, N943, N1048);
xor XOR2 (N2307, N2304, N339);
not NOT1 (N2308, N2289);
nand NAND2 (N2309, N2299, N1044);
xor XOR2 (N2310, N2302, N1716);
nor NOR2 (N2311, N2307, N176);
or OR4 (N2312, N2310, N1166, N1412, N451);
nor NOR4 (N2313, N2308, N1905, N166, N2102);
and AND4 (N2314, N2287, N30, N567, N562);
nor NOR4 (N2315, N2314, N136, N752, N2019);
not NOT1 (N2316, N2280);
nand NAND2 (N2317, N2313, N1775);
xor XOR2 (N2318, N2311, N345);
or OR4 (N2319, N2312, N115, N395, N1234);
nand NAND2 (N2320, N2318, N1417);
buf BUF1 (N2321, N2305);
xor XOR2 (N2322, N2315, N897);
not NOT1 (N2323, N2321);
buf BUF1 (N2324, N2322);
not NOT1 (N2325, N2323);
not NOT1 (N2326, N2319);
and AND4 (N2327, N2316, N913, N1542, N1304);
nor NOR4 (N2328, N2320, N49, N1016, N1701);
and AND4 (N2329, N2328, N889, N1653, N1731);
and AND4 (N2330, N2327, N726, N1999, N576);
nor NOR4 (N2331, N2306, N1006, N1389, N1190);
or OR3 (N2332, N2330, N324, N295);
nor NOR2 (N2333, N2317, N1678);
buf BUF1 (N2334, N2324);
and AND3 (N2335, N2300, N1584, N10);
buf BUF1 (N2336, N2325);
not NOT1 (N2337, N2329);
nand NAND4 (N2338, N2336, N2234, N513, N1021);
buf BUF1 (N2339, N2326);
or OR3 (N2340, N2338, N2322, N540);
nor NOR4 (N2341, N2339, N1994, N48, N1515);
nor NOR2 (N2342, N2309, N1698);
not NOT1 (N2343, N2340);
and AND4 (N2344, N2333, N1146, N523, N72);
nor NOR3 (N2345, N2341, N2008, N2286);
and AND4 (N2346, N2335, N724, N144, N1649);
xor XOR2 (N2347, N2345, N625);
xor XOR2 (N2348, N2347, N2300);
nand NAND3 (N2349, N2346, N918, N1582);
not NOT1 (N2350, N2337);
nand NAND3 (N2351, N2349, N1413, N1961);
and AND2 (N2352, N2331, N371);
buf BUF1 (N2353, N2350);
and AND2 (N2354, N2301, N2350);
or OR2 (N2355, N2343, N2322);
buf BUF1 (N2356, N2342);
nor NOR4 (N2357, N2356, N80, N533, N1125);
nor NOR2 (N2358, N2354, N2230);
not NOT1 (N2359, N2351);
xor XOR2 (N2360, N2353, N811);
xor XOR2 (N2361, N2352, N2245);
nor NOR4 (N2362, N2355, N1138, N818, N2313);
nand NAND2 (N2363, N2334, N1959);
or OR3 (N2364, N2362, N777, N403);
xor XOR2 (N2365, N2361, N917);
nand NAND4 (N2366, N2332, N634, N110, N1357);
nor NOR3 (N2367, N2357, N2293, N1396);
or OR2 (N2368, N2359, N1866);
xor XOR2 (N2369, N2360, N1470);
nor NOR2 (N2370, N2344, N217);
or OR4 (N2371, N2348, N2019, N2066, N418);
nand NAND2 (N2372, N2371, N784);
or OR4 (N2373, N2365, N1820, N995, N240);
nor NOR4 (N2374, N2363, N1272, N1776, N1868);
buf BUF1 (N2375, N2368);
buf BUF1 (N2376, N2358);
and AND3 (N2377, N2373, N2146, N164);
nand NAND3 (N2378, N2364, N40, N598);
not NOT1 (N2379, N2376);
and AND2 (N2380, N2366, N2052);
nand NAND3 (N2381, N2375, N308, N1218);
buf BUF1 (N2382, N2379);
nor NOR4 (N2383, N2367, N1811, N1666, N679);
not NOT1 (N2384, N2377);
not NOT1 (N2385, N2383);
xor XOR2 (N2386, N2385, N2087);
and AND3 (N2387, N2378, N1652, N2090);
or OR2 (N2388, N2372, N132);
nand NAND2 (N2389, N2374, N937);
not NOT1 (N2390, N2386);
xor XOR2 (N2391, N2390, N63);
nor NOR2 (N2392, N2380, N239);
or OR2 (N2393, N2389, N620);
xor XOR2 (N2394, N2369, N1892);
and AND4 (N2395, N2393, N477, N319, N1363);
not NOT1 (N2396, N2387);
nand NAND4 (N2397, N2381, N1480, N1437, N1113);
and AND4 (N2398, N2384, N1050, N696, N1616);
not NOT1 (N2399, N2394);
nor NOR2 (N2400, N2382, N1920);
xor XOR2 (N2401, N2388, N1968);
xor XOR2 (N2402, N2370, N868);
nand NAND3 (N2403, N2400, N2249, N564);
or OR4 (N2404, N2396, N1041, N444, N341);
buf BUF1 (N2405, N2392);
not NOT1 (N2406, N2395);
not NOT1 (N2407, N2401);
or OR3 (N2408, N2404, N781, N738);
nand NAND3 (N2409, N2406, N700, N1521);
not NOT1 (N2410, N2391);
xor XOR2 (N2411, N2409, N761);
not NOT1 (N2412, N2397);
or OR2 (N2413, N2410, N1542);
and AND2 (N2414, N2402, N509);
xor XOR2 (N2415, N2412, N1683);
and AND2 (N2416, N2399, N1876);
nor NOR2 (N2417, N2415, N984);
xor XOR2 (N2418, N2403, N469);
xor XOR2 (N2419, N2407, N956);
and AND2 (N2420, N2405, N831);
or OR4 (N2421, N2420, N886, N2309, N635);
or OR2 (N2422, N2411, N1845);
or OR3 (N2423, N2422, N589, N1321);
buf BUF1 (N2424, N2423);
not NOT1 (N2425, N2418);
nand NAND3 (N2426, N2413, N1932, N1798);
or OR2 (N2427, N2398, N1892);
nand NAND3 (N2428, N2408, N1579, N1770);
nor NOR3 (N2429, N2426, N1333, N59);
and AND3 (N2430, N2421, N202, N484);
nor NOR3 (N2431, N2424, N788, N945);
nor NOR2 (N2432, N2419, N1402);
not NOT1 (N2433, N2432);
not NOT1 (N2434, N2425);
or OR4 (N2435, N2429, N1979, N1191, N2415);
buf BUF1 (N2436, N2417);
nor NOR2 (N2437, N2427, N1876);
buf BUF1 (N2438, N2428);
xor XOR2 (N2439, N2431, N286);
and AND3 (N2440, N2414, N1785, N1614);
xor XOR2 (N2441, N2416, N1943);
xor XOR2 (N2442, N2436, N799);
buf BUF1 (N2443, N2435);
and AND3 (N2444, N2443, N755, N1000);
nand NAND2 (N2445, N2433, N616);
not NOT1 (N2446, N2434);
or OR2 (N2447, N2437, N330);
buf BUF1 (N2448, N2441);
xor XOR2 (N2449, N2444, N419);
not NOT1 (N2450, N2449);
or OR4 (N2451, N2450, N1130, N293, N1307);
nor NOR2 (N2452, N2445, N1538);
nor NOR2 (N2453, N2440, N189);
and AND2 (N2454, N2452, N1327);
not NOT1 (N2455, N2451);
not NOT1 (N2456, N2453);
nand NAND2 (N2457, N2454, N1749);
nor NOR3 (N2458, N2457, N436, N1430);
xor XOR2 (N2459, N2442, N541);
nand NAND2 (N2460, N2456, N627);
buf BUF1 (N2461, N2447);
nor NOR4 (N2462, N2455, N909, N347, N55);
buf BUF1 (N2463, N2460);
nand NAND2 (N2464, N2463, N1948);
nor NOR2 (N2465, N2458, N609);
or OR3 (N2466, N2439, N2007, N2175);
or OR2 (N2467, N2464, N416);
nor NOR2 (N2468, N2438, N284);
xor XOR2 (N2469, N2461, N656);
buf BUF1 (N2470, N2469);
nor NOR3 (N2471, N2467, N510, N1020);
nand NAND3 (N2472, N2470, N868, N139);
or OR3 (N2473, N2430, N2456, N1392);
and AND2 (N2474, N2459, N41);
xor XOR2 (N2475, N2465, N1101);
buf BUF1 (N2476, N2472);
and AND2 (N2477, N2473, N135);
buf BUF1 (N2478, N2462);
not NOT1 (N2479, N2468);
nand NAND3 (N2480, N2479, N2351, N445);
xor XOR2 (N2481, N2466, N2005);
nand NAND4 (N2482, N2446, N1992, N413, N1421);
nand NAND4 (N2483, N2475, N646, N2359, N1867);
and AND3 (N2484, N2482, N1630, N2339);
nor NOR4 (N2485, N2471, N635, N2436, N1719);
xor XOR2 (N2486, N2477, N1143);
and AND3 (N2487, N2448, N780, N456);
and AND3 (N2488, N2485, N2174, N1695);
nand NAND3 (N2489, N2484, N34, N654);
and AND4 (N2490, N2487, N858, N142, N548);
xor XOR2 (N2491, N2489, N1619);
and AND2 (N2492, N2486, N723);
nor NOR4 (N2493, N2476, N99, N1116, N477);
buf BUF1 (N2494, N2490);
not NOT1 (N2495, N2491);
xor XOR2 (N2496, N2488, N1551);
nand NAND4 (N2497, N2483, N2368, N593, N2123);
or OR3 (N2498, N2496, N1012, N69);
not NOT1 (N2499, N2493);
or OR2 (N2500, N2497, N2139);
buf BUF1 (N2501, N2474);
and AND2 (N2502, N2494, N1934);
nor NOR2 (N2503, N2478, N2496);
xor XOR2 (N2504, N2501, N1511);
not NOT1 (N2505, N2502);
or OR4 (N2506, N2505, N2059, N1858, N107);
buf BUF1 (N2507, N2499);
not NOT1 (N2508, N2498);
or OR4 (N2509, N2508, N392, N509, N1041);
nand NAND4 (N2510, N2495, N1072, N1178, N2041);
not NOT1 (N2511, N2506);
or OR3 (N2512, N2480, N161, N1765);
buf BUF1 (N2513, N2512);
nand NAND4 (N2514, N2500, N123, N1724, N479);
nor NOR3 (N2515, N2510, N1207, N2439);
nor NOR4 (N2516, N2511, N1749, N320, N103);
xor XOR2 (N2517, N2516, N1135);
xor XOR2 (N2518, N2507, N2350);
not NOT1 (N2519, N2504);
nand NAND4 (N2520, N2492, N109, N782, N22);
nor NOR3 (N2521, N2509, N1564, N225);
or OR4 (N2522, N2520, N1893, N1977, N108);
not NOT1 (N2523, N2481);
xor XOR2 (N2524, N2518, N845);
and AND3 (N2525, N2515, N2128, N1710);
buf BUF1 (N2526, N2517);
xor XOR2 (N2527, N2514, N1899);
or OR2 (N2528, N2523, N472);
or OR3 (N2529, N2519, N2491, N1556);
nor NOR4 (N2530, N2503, N2036, N1732, N4);
or OR2 (N2531, N2527, N303);
nor NOR3 (N2532, N2531, N297, N1053);
nand NAND4 (N2533, N2521, N1220, N469, N664);
buf BUF1 (N2534, N2522);
xor XOR2 (N2535, N2528, N1110);
buf BUF1 (N2536, N2532);
not NOT1 (N2537, N2534);
nand NAND3 (N2538, N2530, N1397, N2397);
buf BUF1 (N2539, N2533);
buf BUF1 (N2540, N2537);
nand NAND2 (N2541, N2539, N1089);
and AND4 (N2542, N2535, N1509, N1819, N1779);
nor NOR2 (N2543, N2538, N1732);
not NOT1 (N2544, N2524);
nand NAND2 (N2545, N2529, N1503);
and AND2 (N2546, N2544, N1235);
nand NAND3 (N2547, N2540, N1365, N549);
and AND3 (N2548, N2525, N170, N104);
nand NAND2 (N2549, N2545, N1288);
xor XOR2 (N2550, N2526, N1778);
xor XOR2 (N2551, N2549, N1920);
not NOT1 (N2552, N2550);
nand NAND4 (N2553, N2551, N298, N843, N679);
nand NAND4 (N2554, N2536, N567, N2241, N834);
or OR4 (N2555, N2543, N909, N1478, N1583);
or OR4 (N2556, N2541, N349, N2177, N2046);
or OR2 (N2557, N2542, N29);
and AND3 (N2558, N2546, N181, N1626);
nor NOR2 (N2559, N2558, N1342);
buf BUF1 (N2560, N2559);
not NOT1 (N2561, N2554);
and AND3 (N2562, N2547, N1642, N904);
buf BUF1 (N2563, N2557);
not NOT1 (N2564, N2562);
nor NOR4 (N2565, N2564, N881, N264, N175);
nor NOR3 (N2566, N2548, N2403, N2466);
and AND3 (N2567, N2563, N1109, N279);
xor XOR2 (N2568, N2565, N620);
not NOT1 (N2569, N2561);
not NOT1 (N2570, N2566);
nor NOR3 (N2571, N2567, N1129, N662);
nand NAND3 (N2572, N2568, N1452, N222);
or OR4 (N2573, N2571, N1476, N2042, N2092);
xor XOR2 (N2574, N2555, N1587);
nand NAND2 (N2575, N2569, N1864);
nor NOR4 (N2576, N2553, N1042, N108, N458);
not NOT1 (N2577, N2513);
nand NAND4 (N2578, N2573, N1751, N990, N1426);
nor NOR2 (N2579, N2560, N1124);
and AND3 (N2580, N2576, N455, N390);
or OR2 (N2581, N2575, N2071);
not NOT1 (N2582, N2577);
and AND4 (N2583, N2582, N1333, N1901, N1227);
or OR3 (N2584, N2580, N50, N1958);
or OR3 (N2585, N2556, N1527, N1935);
xor XOR2 (N2586, N2572, N1611);
nand NAND2 (N2587, N2585, N480);
nand NAND3 (N2588, N2581, N1929, N1224);
nor NOR3 (N2589, N2587, N1671, N948);
nand NAND4 (N2590, N2579, N1371, N1382, N1109);
nand NAND3 (N2591, N2570, N1976, N532);
buf BUF1 (N2592, N2583);
not NOT1 (N2593, N2592);
buf BUF1 (N2594, N2574);
xor XOR2 (N2595, N2591, N67);
buf BUF1 (N2596, N2584);
buf BUF1 (N2597, N2590);
and AND2 (N2598, N2597, N880);
or OR3 (N2599, N2594, N2458, N1912);
or OR4 (N2600, N2588, N94, N237, N1604);
or OR3 (N2601, N2552, N2188, N2211);
buf BUF1 (N2602, N2600);
xor XOR2 (N2603, N2596, N2233);
xor XOR2 (N2604, N2601, N239);
nand NAND3 (N2605, N2586, N235, N1204);
and AND3 (N2606, N2595, N148, N767);
not NOT1 (N2607, N2602);
and AND2 (N2608, N2589, N2528);
xor XOR2 (N2609, N2599, N1416);
nor NOR4 (N2610, N2607, N1236, N965, N522);
or OR3 (N2611, N2606, N2543, N1910);
nor NOR4 (N2612, N2578, N717, N525, N182);
nand NAND4 (N2613, N2598, N1334, N2580, N1474);
nand NAND3 (N2614, N2609, N836, N402);
nor NOR3 (N2615, N2614, N628, N1240);
or OR2 (N2616, N2604, N899);
nand NAND3 (N2617, N2615, N1080, N2233);
or OR4 (N2618, N2613, N353, N976, N1854);
nand NAND3 (N2619, N2608, N817, N729);
nand NAND3 (N2620, N2593, N1316, N1392);
not NOT1 (N2621, N2611);
or OR4 (N2622, N2619, N1180, N1972, N2103);
buf BUF1 (N2623, N2610);
not NOT1 (N2624, N2620);
and AND3 (N2625, N2605, N2033, N1634);
buf BUF1 (N2626, N2603);
xor XOR2 (N2627, N2623, N176);
or OR4 (N2628, N2625, N2067, N1781, N1476);
nor NOR2 (N2629, N2621, N2586);
and AND2 (N2630, N2616, N2104);
not NOT1 (N2631, N2628);
buf BUF1 (N2632, N2624);
or OR4 (N2633, N2632, N373, N1747, N1358);
and AND2 (N2634, N2633, N1039);
and AND3 (N2635, N2622, N643, N1966);
nand NAND4 (N2636, N2634, N838, N914, N1807);
buf BUF1 (N2637, N2612);
nor NOR3 (N2638, N2630, N1883, N522);
and AND4 (N2639, N2635, N1777, N520, N2010);
and AND4 (N2640, N2627, N2344, N2365, N1454);
nand NAND2 (N2641, N2638, N2430);
nor NOR4 (N2642, N2636, N538, N247, N2151);
buf BUF1 (N2643, N2629);
buf BUF1 (N2644, N2631);
nor NOR2 (N2645, N2617, N823);
not NOT1 (N2646, N2626);
and AND2 (N2647, N2644, N1794);
and AND4 (N2648, N2645, N2227, N1191, N948);
and AND3 (N2649, N2640, N1550, N296);
buf BUF1 (N2650, N2647);
or OR3 (N2651, N2649, N2635, N855);
not NOT1 (N2652, N2643);
nor NOR3 (N2653, N2650, N1567, N69);
nand NAND3 (N2654, N2651, N661, N1776);
or OR4 (N2655, N2637, N905, N2621, N1194);
nand NAND4 (N2656, N2642, N2448, N58, N1582);
or OR4 (N2657, N2656, N1109, N1859, N497);
not NOT1 (N2658, N2646);
and AND3 (N2659, N2639, N2353, N1481);
and AND2 (N2660, N2654, N1882);
or OR2 (N2661, N2653, N2621);
xor XOR2 (N2662, N2661, N18);
xor XOR2 (N2663, N2657, N671);
nor NOR4 (N2664, N2618, N1205, N1538, N946);
nor NOR3 (N2665, N2655, N854, N1558);
nor NOR2 (N2666, N2660, N2634);
nand NAND4 (N2667, N2648, N2244, N1226, N2535);
xor XOR2 (N2668, N2665, N2195);
not NOT1 (N2669, N2667);
not NOT1 (N2670, N2664);
xor XOR2 (N2671, N2666, N2207);
not NOT1 (N2672, N2668);
and AND3 (N2673, N2652, N1870, N1762);
and AND2 (N2674, N2670, N747);
nor NOR2 (N2675, N2663, N1048);
nor NOR2 (N2676, N2672, N164);
xor XOR2 (N2677, N2669, N108);
not NOT1 (N2678, N2641);
buf BUF1 (N2679, N2658);
or OR2 (N2680, N2679, N862);
buf BUF1 (N2681, N2659);
xor XOR2 (N2682, N2673, N357);
not NOT1 (N2683, N2681);
not NOT1 (N2684, N2683);
nand NAND4 (N2685, N2675, N129, N351, N1953);
buf BUF1 (N2686, N2685);
not NOT1 (N2687, N2686);
nor NOR3 (N2688, N2682, N2383, N595);
buf BUF1 (N2689, N2678);
xor XOR2 (N2690, N2688, N1624);
xor XOR2 (N2691, N2687, N1959);
nor NOR4 (N2692, N2677, N2032, N1944, N2157);
or OR3 (N2693, N2689, N1281, N1988);
and AND2 (N2694, N2671, N2230);
and AND2 (N2695, N2693, N2461);
nand NAND4 (N2696, N2690, N2035, N352, N203);
nor NOR3 (N2697, N2691, N179, N789);
xor XOR2 (N2698, N2697, N1113);
nor NOR3 (N2699, N2698, N1887, N2428);
nand NAND2 (N2700, N2696, N454);
not NOT1 (N2701, N2695);
nand NAND3 (N2702, N2674, N1001, N487);
nand NAND3 (N2703, N2680, N887, N1014);
and AND2 (N2704, N2662, N2177);
nor NOR4 (N2705, N2700, N1259, N2052, N2684);
and AND3 (N2706, N1420, N79, N2455);
or OR2 (N2707, N2702, N2546);
xor XOR2 (N2708, N2676, N1695);
nor NOR2 (N2709, N2706, N1155);
xor XOR2 (N2710, N2703, N944);
not NOT1 (N2711, N2692);
xor XOR2 (N2712, N2708, N639);
xor XOR2 (N2713, N2705, N583);
or OR3 (N2714, N2694, N1618, N1534);
buf BUF1 (N2715, N2699);
nor NOR2 (N2716, N2710, N919);
nand NAND2 (N2717, N2715, N2030);
or OR2 (N2718, N2709, N1866);
xor XOR2 (N2719, N2711, N1323);
nor NOR4 (N2720, N2717, N1213, N323, N2414);
buf BUF1 (N2721, N2712);
not NOT1 (N2722, N2721);
not NOT1 (N2723, N2720);
nor NOR3 (N2724, N2714, N2640, N1581);
not NOT1 (N2725, N2701);
not NOT1 (N2726, N2704);
nor NOR4 (N2727, N2723, N643, N794, N313);
nor NOR3 (N2728, N2727, N1318, N1424);
not NOT1 (N2729, N2719);
buf BUF1 (N2730, N2724);
or OR2 (N2731, N2729, N1127);
and AND4 (N2732, N2730, N1832, N1903, N1420);
or OR4 (N2733, N2732, N729, N537, N834);
buf BUF1 (N2734, N2733);
or OR3 (N2735, N2726, N2059, N2528);
nand NAND4 (N2736, N2735, N1489, N1666, N1534);
or OR4 (N2737, N2713, N2466, N1018, N731);
xor XOR2 (N2738, N2734, N893);
nor NOR3 (N2739, N2737, N1465, N2522);
not NOT1 (N2740, N2731);
or OR4 (N2741, N2738, N1938, N1217, N2455);
nor NOR3 (N2742, N2718, N945, N1137);
not NOT1 (N2743, N2740);
and AND3 (N2744, N2722, N2540, N764);
xor XOR2 (N2745, N2744, N886);
buf BUF1 (N2746, N2739);
or OR2 (N2747, N2716, N2338);
not NOT1 (N2748, N2743);
or OR3 (N2749, N2725, N695, N1516);
xor XOR2 (N2750, N2707, N2659);
nor NOR3 (N2751, N2736, N628, N535);
xor XOR2 (N2752, N2746, N1628);
nor NOR4 (N2753, N2741, N716, N1358, N1580);
nand NAND3 (N2754, N2753, N2688, N295);
buf BUF1 (N2755, N2754);
nor NOR4 (N2756, N2751, N2267, N1214, N849);
not NOT1 (N2757, N2749);
nor NOR3 (N2758, N2742, N1294, N1571);
xor XOR2 (N2759, N2758, N2241);
nand NAND3 (N2760, N2745, N522, N1192);
nand NAND4 (N2761, N2747, N2163, N540, N2458);
or OR4 (N2762, N2752, N974, N1255, N1634);
not NOT1 (N2763, N2759);
xor XOR2 (N2764, N2756, N293);
nor NOR2 (N2765, N2764, N2670);
buf BUF1 (N2766, N2761);
nor NOR4 (N2767, N2763, N2595, N1648, N1389);
xor XOR2 (N2768, N2755, N2534);
buf BUF1 (N2769, N2767);
buf BUF1 (N2770, N2766);
or OR4 (N2771, N2765, N908, N1724, N2658);
or OR2 (N2772, N2728, N2073);
not NOT1 (N2773, N2760);
nor NOR2 (N2774, N2750, N286);
and AND4 (N2775, N2769, N2581, N31, N1184);
not NOT1 (N2776, N2770);
and AND3 (N2777, N2768, N2585, N1811);
not NOT1 (N2778, N2774);
not NOT1 (N2779, N2762);
or OR2 (N2780, N2777, N1832);
buf BUF1 (N2781, N2757);
or OR2 (N2782, N2780, N62);
not NOT1 (N2783, N2772);
and AND4 (N2784, N2775, N2478, N1938, N1742);
buf BUF1 (N2785, N2784);
xor XOR2 (N2786, N2779, N2528);
nand NAND4 (N2787, N2785, N204, N223, N1809);
xor XOR2 (N2788, N2748, N644);
or OR4 (N2789, N2778, N2349, N1384, N1764);
xor XOR2 (N2790, N2786, N2334);
and AND2 (N2791, N2782, N1565);
nand NAND4 (N2792, N2791, N866, N2760, N446);
nor NOR2 (N2793, N2790, N1309);
or OR4 (N2794, N2787, N204, N70, N1944);
buf BUF1 (N2795, N2789);
or OR3 (N2796, N2783, N124, N1047);
or OR2 (N2797, N2794, N2630);
buf BUF1 (N2798, N2771);
nand NAND2 (N2799, N2773, N2459);
not NOT1 (N2800, N2795);
nor NOR3 (N2801, N2800, N1540, N2370);
or OR3 (N2802, N2776, N503, N384);
xor XOR2 (N2803, N2798, N2187);
or OR4 (N2804, N2793, N155, N2308, N638);
and AND3 (N2805, N2788, N2142, N227);
or OR3 (N2806, N2796, N648, N1536);
nand NAND4 (N2807, N2781, N632, N1330, N288);
and AND2 (N2808, N2792, N1095);
not NOT1 (N2809, N2808);
and AND3 (N2810, N2807, N745, N2792);
buf BUF1 (N2811, N2804);
nand NAND2 (N2812, N2803, N1784);
buf BUF1 (N2813, N2810);
nand NAND2 (N2814, N2802, N644);
nand NAND2 (N2815, N2799, N2038);
buf BUF1 (N2816, N2811);
not NOT1 (N2817, N2797);
nand NAND4 (N2818, N2815, N1318, N1116, N838);
buf BUF1 (N2819, N2805);
or OR4 (N2820, N2816, N656, N2231, N19);
or OR2 (N2821, N2814, N775);
xor XOR2 (N2822, N2821, N1042);
xor XOR2 (N2823, N2809, N1776);
and AND2 (N2824, N2822, N909);
or OR4 (N2825, N2824, N1045, N1333, N186);
not NOT1 (N2826, N2806);
and AND3 (N2827, N2825, N2438, N918);
not NOT1 (N2828, N2817);
xor XOR2 (N2829, N2813, N821);
buf BUF1 (N2830, N2818);
nor NOR2 (N2831, N2823, N974);
nand NAND4 (N2832, N2828, N957, N2455, N2411);
or OR2 (N2833, N2830, N2103);
buf BUF1 (N2834, N2801);
nand NAND4 (N2835, N2819, N1123, N1707, N1704);
nand NAND4 (N2836, N2829, N821, N1290, N1974);
nor NOR3 (N2837, N2833, N2598, N2708);
nand NAND2 (N2838, N2812, N2304);
nor NOR3 (N2839, N2832, N1136, N2108);
or OR4 (N2840, N2834, N346, N259, N1642);
nor NOR3 (N2841, N2837, N239, N550);
and AND2 (N2842, N2836, N995);
and AND3 (N2843, N2826, N1049, N127);
and AND4 (N2844, N2840, N743, N2435, N1229);
or OR4 (N2845, N2831, N526, N209, N948);
xor XOR2 (N2846, N2839, N1971);
and AND3 (N2847, N2844, N443, N2362);
buf BUF1 (N2848, N2845);
nor NOR3 (N2849, N2835, N386, N213);
buf BUF1 (N2850, N2849);
and AND4 (N2851, N2841, N2261, N285, N1637);
and AND3 (N2852, N2850, N65, N1677);
or OR2 (N2853, N2846, N2703);
or OR3 (N2854, N2847, N1347, N2646);
not NOT1 (N2855, N2842);
not NOT1 (N2856, N2852);
nand NAND3 (N2857, N2855, N1750, N1601);
and AND4 (N2858, N2843, N1272, N2496, N1342);
and AND4 (N2859, N2827, N233, N1023, N102);
not NOT1 (N2860, N2857);
not NOT1 (N2861, N2859);
or OR4 (N2862, N2861, N855, N1244, N2350);
xor XOR2 (N2863, N2858, N636);
or OR3 (N2864, N2856, N1860, N1168);
xor XOR2 (N2865, N2862, N83);
nand NAND2 (N2866, N2851, N720);
nor NOR2 (N2867, N2866, N1107);
buf BUF1 (N2868, N2865);
and AND3 (N2869, N2864, N2425, N1186);
or OR2 (N2870, N2860, N288);
not NOT1 (N2871, N2854);
and AND2 (N2872, N2869, N1775);
nor NOR4 (N2873, N2867, N810, N1290, N602);
not NOT1 (N2874, N2870);
nor NOR4 (N2875, N2868, N790, N994, N1494);
nor NOR4 (N2876, N2875, N2792, N2048, N1968);
nand NAND2 (N2877, N2820, N869);
and AND2 (N2878, N2863, N638);
buf BUF1 (N2879, N2874);
nor NOR4 (N2880, N2879, N1456, N2861, N144);
nand NAND2 (N2881, N2878, N113);
nand NAND4 (N2882, N2873, N1228, N1409, N1766);
nor NOR4 (N2883, N2880, N1627, N1785, N2074);
xor XOR2 (N2884, N2853, N995);
not NOT1 (N2885, N2883);
buf BUF1 (N2886, N2885);
nand NAND3 (N2887, N2838, N920, N1795);
nand NAND2 (N2888, N2871, N2777);
xor XOR2 (N2889, N2881, N2829);
not NOT1 (N2890, N2887);
nor NOR3 (N2891, N2888, N1075, N2526);
and AND2 (N2892, N2884, N1419);
and AND4 (N2893, N2882, N2436, N1327, N1574);
nand NAND3 (N2894, N2891, N2583, N2659);
nor NOR2 (N2895, N2893, N678);
xor XOR2 (N2896, N2889, N1070);
or OR3 (N2897, N2877, N729, N1673);
buf BUF1 (N2898, N2892);
nand NAND3 (N2899, N2894, N1513, N2572);
and AND3 (N2900, N2890, N2474, N1557);
or OR4 (N2901, N2899, N618, N375, N2257);
nor NOR3 (N2902, N2901, N1, N2268);
and AND4 (N2903, N2876, N738, N2076, N2881);
and AND3 (N2904, N2872, N1357, N1422);
not NOT1 (N2905, N2898);
and AND2 (N2906, N2902, N1640);
nor NOR2 (N2907, N2905, N1921);
not NOT1 (N2908, N2897);
and AND4 (N2909, N2895, N1474, N2315, N446);
and AND3 (N2910, N2848, N2400, N2650);
not NOT1 (N2911, N2906);
or OR2 (N2912, N2900, N986);
xor XOR2 (N2913, N2908, N543);
nand NAND3 (N2914, N2909, N1981, N2620);
and AND4 (N2915, N2896, N2838, N451, N399);
nand NAND3 (N2916, N2904, N2413, N2303);
nand NAND3 (N2917, N2886, N2583, N1991);
xor XOR2 (N2918, N2903, N2232);
buf BUF1 (N2919, N2915);
xor XOR2 (N2920, N2913, N636);
buf BUF1 (N2921, N2907);
and AND3 (N2922, N2918, N312, N2120);
and AND4 (N2923, N2910, N894, N2250, N1985);
xor XOR2 (N2924, N2914, N1386);
nand NAND4 (N2925, N2922, N2474, N1237, N1476);
buf BUF1 (N2926, N2920);
xor XOR2 (N2927, N2924, N903);
xor XOR2 (N2928, N2912, N1133);
nand NAND4 (N2929, N2926, N1293, N2567, N1271);
nor NOR4 (N2930, N2928, N2916, N1156, N1914);
not NOT1 (N2931, N838);
nand NAND4 (N2932, N2911, N1597, N2244, N802);
buf BUF1 (N2933, N2930);
or OR2 (N2934, N2931, N1621);
xor XOR2 (N2935, N2923, N111);
or OR3 (N2936, N2927, N1853, N155);
not NOT1 (N2937, N2932);
and AND3 (N2938, N2934, N2192, N1397);
nor NOR4 (N2939, N2925, N123, N2728, N1861);
not NOT1 (N2940, N2919);
nor NOR3 (N2941, N2917, N1677, N2635);
nor NOR2 (N2942, N2933, N2431);
buf BUF1 (N2943, N2937);
and AND3 (N2944, N2921, N2807, N629);
nor NOR3 (N2945, N2936, N1088, N2820);
not NOT1 (N2946, N2940);
or OR4 (N2947, N2939, N467, N227, N2651);
and AND3 (N2948, N2942, N2410, N339);
buf BUF1 (N2949, N2944);
xor XOR2 (N2950, N2947, N2733);
and AND2 (N2951, N2935, N2480);
nand NAND2 (N2952, N2949, N440);
nor NOR4 (N2953, N2929, N10, N2184, N1462);
nor NOR3 (N2954, N2941, N2335, N2336);
and AND2 (N2955, N2938, N203);
and AND2 (N2956, N2955, N982);
or OR3 (N2957, N2943, N2441, N1616);
and AND3 (N2958, N2946, N213, N1658);
xor XOR2 (N2959, N2956, N1471);
xor XOR2 (N2960, N2954, N79);
xor XOR2 (N2961, N2959, N2786);
buf BUF1 (N2962, N2950);
not NOT1 (N2963, N2957);
not NOT1 (N2964, N2948);
nor NOR3 (N2965, N2963, N2317, N792);
or OR2 (N2966, N2960, N959);
or OR2 (N2967, N2952, N1762);
or OR4 (N2968, N2967, N228, N342, N905);
not NOT1 (N2969, N2951);
nand NAND4 (N2970, N2965, N1943, N28, N2253);
nand NAND3 (N2971, N2953, N1969, N2863);
not NOT1 (N2972, N2962);
nand NAND2 (N2973, N2964, N402);
buf BUF1 (N2974, N2958);
nor NOR2 (N2975, N2970, N2193);
nand NAND2 (N2976, N2945, N1323);
buf BUF1 (N2977, N2976);
or OR2 (N2978, N2975, N1621);
or OR2 (N2979, N2961, N374);
and AND2 (N2980, N2966, N2265);
not NOT1 (N2981, N2977);
nand NAND4 (N2982, N2980, N300, N2081, N2011);
and AND4 (N2983, N2978, N363, N1609, N2031);
nor NOR4 (N2984, N2972, N1104, N367, N1889);
nand NAND4 (N2985, N2984, N2559, N1150, N2597);
nand NAND4 (N2986, N2974, N372, N1895, N1373);
buf BUF1 (N2987, N2973);
or OR3 (N2988, N2985, N346, N2986);
not NOT1 (N2989, N359);
xor XOR2 (N2990, N2981, N1091);
or OR3 (N2991, N2968, N29, N702);
and AND3 (N2992, N2983, N843, N2287);
or OR2 (N2993, N2991, N1318);
and AND3 (N2994, N2988, N31, N113);
and AND3 (N2995, N2992, N2052, N686);
or OR4 (N2996, N2995, N2225, N273, N2898);
nor NOR4 (N2997, N2971, N1145, N1561, N2275);
xor XOR2 (N2998, N2993, N1825);
or OR2 (N2999, N2996, N2786);
xor XOR2 (N3000, N2990, N1099);
or OR3 (N3001, N2998, N99, N2407);
and AND3 (N3002, N2999, N1069, N433);
or OR2 (N3003, N2969, N2510);
and AND4 (N3004, N3002, N2828, N1218, N101);
xor XOR2 (N3005, N3004, N508);
not NOT1 (N3006, N3005);
buf BUF1 (N3007, N3003);
xor XOR2 (N3008, N3006, N1355);
buf BUF1 (N3009, N2982);
not NOT1 (N3010, N3009);
and AND2 (N3011, N3000, N1378);
nor NOR4 (N3012, N2987, N1765, N747, N2341);
not NOT1 (N3013, N2989);
or OR2 (N3014, N3007, N2085);
or OR2 (N3015, N2979, N715);
or OR4 (N3016, N3010, N1821, N198, N1567);
nand NAND4 (N3017, N3016, N1718, N1274, N1226);
xor XOR2 (N3018, N2994, N938);
xor XOR2 (N3019, N3018, N1319);
buf BUF1 (N3020, N3017);
or OR4 (N3021, N3001, N55, N1492, N2047);
nand NAND4 (N3022, N3015, N1764, N508, N1128);
nor NOR2 (N3023, N3022, N2072);
buf BUF1 (N3024, N3021);
buf BUF1 (N3025, N3012);
buf BUF1 (N3026, N3023);
xor XOR2 (N3027, N2997, N743);
not NOT1 (N3028, N3020);
or OR3 (N3029, N3008, N1480, N2592);
nor NOR4 (N3030, N3028, N1811, N656, N1894);
buf BUF1 (N3031, N3027);
nand NAND3 (N3032, N3014, N3022, N1267);
buf BUF1 (N3033, N3024);
or OR2 (N3034, N3029, N1097);
buf BUF1 (N3035, N3031);
not NOT1 (N3036, N3026);
not NOT1 (N3037, N3011);
buf BUF1 (N3038, N3032);
xor XOR2 (N3039, N3013, N1974);
nor NOR3 (N3040, N3033, N1696, N1898);
buf BUF1 (N3041, N3039);
not NOT1 (N3042, N3040);
buf BUF1 (N3043, N3035);
xor XOR2 (N3044, N3037, N2193);
xor XOR2 (N3045, N3044, N2456);
and AND3 (N3046, N3042, N1270, N2025);
nand NAND4 (N3047, N3025, N1411, N882, N1992);
and AND2 (N3048, N3036, N2193);
xor XOR2 (N3049, N3019, N1907);
and AND3 (N3050, N3041, N746, N98);
or OR3 (N3051, N3034, N2338, N1381);
or OR3 (N3052, N3047, N2210, N164);
not NOT1 (N3053, N3030);
xor XOR2 (N3054, N3046, N2142);
buf BUF1 (N3055, N3051);
or OR4 (N3056, N3048, N2101, N849, N1479);
not NOT1 (N3057, N3055);
buf BUF1 (N3058, N3045);
nand NAND4 (N3059, N3049, N372, N2465, N679);
xor XOR2 (N3060, N3038, N320);
xor XOR2 (N3061, N3057, N1420);
nand NAND2 (N3062, N3050, N2145);
buf BUF1 (N3063, N3058);
nand NAND2 (N3064, N3060, N820);
and AND3 (N3065, N3059, N1611, N2002);
and AND2 (N3066, N3052, N1124);
or OR3 (N3067, N3053, N3016, N2655);
nor NOR4 (N3068, N3056, N1905, N1497, N288);
xor XOR2 (N3069, N3068, N203);
and AND2 (N3070, N3063, N2233);
and AND4 (N3071, N3065, N492, N654, N261);
xor XOR2 (N3072, N3062, N1901);
nand NAND4 (N3073, N3066, N664, N1362, N114);
or OR2 (N3074, N3061, N2760);
nor NOR3 (N3075, N3054, N2768, N1271);
buf BUF1 (N3076, N3072);
nand NAND4 (N3077, N3071, N2058, N293, N352);
xor XOR2 (N3078, N3077, N1334);
buf BUF1 (N3079, N3075);
xor XOR2 (N3080, N3069, N745);
not NOT1 (N3081, N3076);
not NOT1 (N3082, N3081);
not NOT1 (N3083, N3064);
nand NAND3 (N3084, N3067, N2941, N1134);
nor NOR4 (N3085, N3073, N142, N1801, N823);
nand NAND2 (N3086, N3043, N169);
buf BUF1 (N3087, N3083);
buf BUF1 (N3088, N3080);
and AND4 (N3089, N3078, N1680, N1877, N1705);
and AND4 (N3090, N3074, N3020, N1502, N2428);
nand NAND4 (N3091, N3085, N2902, N473, N1125);
buf BUF1 (N3092, N3070);
xor XOR2 (N3093, N3089, N2237);
nand NAND2 (N3094, N3093, N2683);
and AND2 (N3095, N3086, N1034);
not NOT1 (N3096, N3088);
and AND4 (N3097, N3090, N2635, N396, N1050);
nor NOR4 (N3098, N3079, N1662, N249, N2730);
nor NOR2 (N3099, N3082, N2240);
nand NAND2 (N3100, N3084, N2381);
buf BUF1 (N3101, N3097);
nand NAND3 (N3102, N3101, N596, N629);
not NOT1 (N3103, N3087);
nand NAND2 (N3104, N3102, N1940);
nand NAND3 (N3105, N3099, N761, N2420);
nor NOR2 (N3106, N3105, N475);
or OR4 (N3107, N3091, N1704, N2431, N118);
not NOT1 (N3108, N3096);
nand NAND4 (N3109, N3092, N57, N2408, N482);
and AND4 (N3110, N3106, N1012, N2214, N1482);
buf BUF1 (N3111, N3110);
not NOT1 (N3112, N3100);
nor NOR4 (N3113, N3112, N965, N1810, N143);
nor NOR4 (N3114, N3095, N1502, N242, N2443);
nand NAND3 (N3115, N3103, N2276, N2367);
nor NOR4 (N3116, N3094, N2180, N82, N2286);
xor XOR2 (N3117, N3109, N2673);
nand NAND4 (N3118, N3113, N2069, N2827, N1624);
xor XOR2 (N3119, N3117, N1960);
xor XOR2 (N3120, N3116, N2795);
nand NAND3 (N3121, N3115, N2467, N2880);
or OR3 (N3122, N3098, N173, N1246);
and AND2 (N3123, N3108, N1981);
or OR2 (N3124, N3114, N60);
or OR4 (N3125, N3123, N516, N769, N2740);
nor NOR3 (N3126, N3119, N246, N127);
nor NOR4 (N3127, N3104, N1829, N1661, N876);
or OR3 (N3128, N3127, N1923, N1432);
buf BUF1 (N3129, N3128);
buf BUF1 (N3130, N3111);
not NOT1 (N3131, N3124);
nor NOR3 (N3132, N3130, N2145, N385);
nand NAND4 (N3133, N3107, N1862, N2787, N1644);
xor XOR2 (N3134, N3120, N189);
and AND4 (N3135, N3125, N1833, N676, N535);
xor XOR2 (N3136, N3129, N3122);
and AND2 (N3137, N2152, N862);
nand NAND2 (N3138, N3137, N1759);
buf BUF1 (N3139, N3118);
not NOT1 (N3140, N3138);
nor NOR4 (N3141, N3121, N2040, N2829, N86);
nor NOR3 (N3142, N3133, N1653, N548);
and AND4 (N3143, N3131, N1284, N2808, N3019);
or OR3 (N3144, N3134, N2410, N1869);
not NOT1 (N3145, N3142);
nor NOR3 (N3146, N3145, N927, N1561);
not NOT1 (N3147, N3141);
nor NOR4 (N3148, N3136, N1028, N2645, N981);
and AND2 (N3149, N3132, N1611);
and AND2 (N3150, N3143, N3134);
or OR3 (N3151, N3135, N1713, N2598);
buf BUF1 (N3152, N3139);
nor NOR4 (N3153, N3152, N2433, N3, N1868);
or OR2 (N3154, N3150, N1983);
nand NAND2 (N3155, N3154, N1431);
nor NOR3 (N3156, N3146, N2049, N432);
or OR2 (N3157, N3148, N2523);
or OR2 (N3158, N3147, N2277);
nor NOR3 (N3159, N3144, N2166, N1519);
xor XOR2 (N3160, N3149, N81);
and AND4 (N3161, N3153, N2203, N260, N2041);
nand NAND3 (N3162, N3159, N1756, N1876);
not NOT1 (N3163, N3126);
not NOT1 (N3164, N3162);
or OR4 (N3165, N3163, N1533, N2279, N874);
or OR4 (N3166, N3157, N184, N1043, N1582);
nand NAND4 (N3167, N3151, N1514, N1733, N3160);
nand NAND3 (N3168, N2625, N1498, N2710);
and AND3 (N3169, N3165, N611, N425);
nor NOR4 (N3170, N3158, N2278, N634, N1559);
not NOT1 (N3171, N3169);
nand NAND4 (N3172, N3168, N3083, N1060, N1850);
not NOT1 (N3173, N3170);
or OR2 (N3174, N3140, N107);
and AND3 (N3175, N3166, N463, N2034);
or OR3 (N3176, N3164, N2500, N1359);
xor XOR2 (N3177, N3173, N1246);
not NOT1 (N3178, N3171);
xor XOR2 (N3179, N3167, N61);
and AND4 (N3180, N3178, N1676, N1435, N1958);
nor NOR3 (N3181, N3161, N379, N2742);
not NOT1 (N3182, N3175);
nand NAND2 (N3183, N3176, N2890);
nand NAND3 (N3184, N3180, N455, N1760);
buf BUF1 (N3185, N3172);
or OR2 (N3186, N3183, N2569);
or OR4 (N3187, N3181, N711, N2409, N136);
and AND4 (N3188, N3187, N2212, N2972, N1215);
not NOT1 (N3189, N3186);
nor NOR3 (N3190, N3189, N2279, N580);
or OR3 (N3191, N3182, N1756, N58);
buf BUF1 (N3192, N3191);
nor NOR2 (N3193, N3184, N1243);
buf BUF1 (N3194, N3155);
nand NAND4 (N3195, N3156, N587, N1908, N1059);
nand NAND3 (N3196, N3192, N273, N1945);
not NOT1 (N3197, N3179);
xor XOR2 (N3198, N3197, N3075);
buf BUF1 (N3199, N3174);
nand NAND3 (N3200, N3196, N849, N1643);
nor NOR2 (N3201, N3199, N3062);
nor NOR2 (N3202, N3177, N1047);
xor XOR2 (N3203, N3193, N400);
xor XOR2 (N3204, N3188, N218);
nand NAND4 (N3205, N3202, N249, N2375, N402);
buf BUF1 (N3206, N3204);
xor XOR2 (N3207, N3200, N3167);
buf BUF1 (N3208, N3206);
nand NAND4 (N3209, N3205, N2054, N148, N709);
xor XOR2 (N3210, N3201, N1712);
xor XOR2 (N3211, N3207, N1844);
not NOT1 (N3212, N3209);
xor XOR2 (N3213, N3211, N2100);
xor XOR2 (N3214, N3198, N725);
nor NOR4 (N3215, N3203, N100, N2007, N1621);
nand NAND4 (N3216, N3212, N1759, N2286, N1967);
xor XOR2 (N3217, N3216, N1243);
and AND3 (N3218, N3195, N1984, N1421);
nor NOR2 (N3219, N3217, N2423);
or OR4 (N3220, N3194, N2746, N1351, N1115);
or OR4 (N3221, N3215, N2427, N1180, N2531);
or OR3 (N3222, N3208, N1807, N441);
not NOT1 (N3223, N3214);
not NOT1 (N3224, N3219);
or OR2 (N3225, N3213, N2328);
or OR4 (N3226, N3220, N1460, N726, N2346);
xor XOR2 (N3227, N3226, N1933);
nor NOR3 (N3228, N3210, N768, N384);
or OR2 (N3229, N3225, N2835);
buf BUF1 (N3230, N3185);
or OR4 (N3231, N3228, N3017, N1397, N2171);
nand NAND3 (N3232, N3231, N783, N2959);
nor NOR3 (N3233, N3218, N953, N726);
not NOT1 (N3234, N3221);
or OR4 (N3235, N3234, N30, N1102, N1454);
not NOT1 (N3236, N3222);
or OR3 (N3237, N3232, N3092, N3107);
or OR2 (N3238, N3229, N496);
xor XOR2 (N3239, N3190, N1777);
buf BUF1 (N3240, N3227);
nor NOR2 (N3241, N3240, N1241);
xor XOR2 (N3242, N3230, N1891);
or OR3 (N3243, N3224, N2470, N1147);
xor XOR2 (N3244, N3233, N876);
and AND2 (N3245, N3235, N454);
or OR4 (N3246, N3241, N1798, N1680, N2925);
xor XOR2 (N3247, N3244, N105);
not NOT1 (N3248, N3238);
xor XOR2 (N3249, N3245, N206);
nand NAND3 (N3250, N3242, N1366, N2206);
nor NOR4 (N3251, N3250, N2189, N25, N63);
or OR3 (N3252, N3239, N327, N1700);
buf BUF1 (N3253, N3236);
and AND2 (N3254, N3248, N732);
xor XOR2 (N3255, N3251, N1351);
xor XOR2 (N3256, N3237, N2268);
xor XOR2 (N3257, N3243, N2174);
not NOT1 (N3258, N3255);
not NOT1 (N3259, N3253);
nand NAND4 (N3260, N3247, N1883, N3068, N563);
xor XOR2 (N3261, N3257, N578);
not NOT1 (N3262, N3246);
or OR3 (N3263, N3256, N1604, N1696);
not NOT1 (N3264, N3261);
not NOT1 (N3265, N3254);
and AND4 (N3266, N3252, N2802, N1641, N1939);
nand NAND4 (N3267, N3264, N2235, N1932, N83);
not NOT1 (N3268, N3267);
and AND4 (N3269, N3265, N3194, N229, N1646);
not NOT1 (N3270, N3262);
or OR3 (N3271, N3266, N3251, N352);
and AND3 (N3272, N3249, N1436, N2485);
or OR4 (N3273, N3223, N2780, N2001, N983);
xor XOR2 (N3274, N3273, N3201);
nor NOR3 (N3275, N3269, N637, N3165);
xor XOR2 (N3276, N3274, N2873);
buf BUF1 (N3277, N3268);
xor XOR2 (N3278, N3276, N2872);
buf BUF1 (N3279, N3275);
buf BUF1 (N3280, N3258);
nand NAND3 (N3281, N3270, N477, N1877);
not NOT1 (N3282, N3263);
xor XOR2 (N3283, N3279, N3192);
and AND3 (N3284, N3259, N3130, N2825);
or OR3 (N3285, N3283, N2676, N452);
buf BUF1 (N3286, N3277);
nor NOR2 (N3287, N3271, N1449);
nor NOR3 (N3288, N3272, N939, N1275);
or OR4 (N3289, N3278, N2829, N322, N378);
nor NOR4 (N3290, N3281, N1763, N574, N801);
xor XOR2 (N3291, N3285, N2395);
or OR3 (N3292, N3290, N1596, N3026);
nor NOR3 (N3293, N3287, N760, N1648);
and AND4 (N3294, N3286, N2850, N1009, N2650);
buf BUF1 (N3295, N3284);
or OR4 (N3296, N3291, N2396, N464, N1862);
nor NOR2 (N3297, N3293, N1477);
nand NAND4 (N3298, N3280, N1042, N3161, N732);
and AND2 (N3299, N3260, N1540);
xor XOR2 (N3300, N3299, N1542);
nor NOR2 (N3301, N3292, N2690);
xor XOR2 (N3302, N3298, N2633);
not NOT1 (N3303, N3297);
xor XOR2 (N3304, N3303, N1023);
xor XOR2 (N3305, N3302, N2449);
xor XOR2 (N3306, N3305, N2530);
and AND4 (N3307, N3300, N2973, N636, N1755);
nand NAND2 (N3308, N3288, N770);
nor NOR2 (N3309, N3308, N648);
nand NAND3 (N3310, N3295, N1204, N1505);
or OR3 (N3311, N3306, N2724, N1160);
nor NOR2 (N3312, N3289, N1818);
and AND3 (N3313, N3310, N1177, N1662);
not NOT1 (N3314, N3301);
or OR3 (N3315, N3309, N558, N3227);
or OR3 (N3316, N3314, N1520, N2991);
and AND4 (N3317, N3316, N1550, N3048, N503);
not NOT1 (N3318, N3282);
nand NAND2 (N3319, N3318, N452);
buf BUF1 (N3320, N3294);
xor XOR2 (N3321, N3296, N1505);
or OR4 (N3322, N3307, N176, N660, N2035);
xor XOR2 (N3323, N3311, N145);
or OR4 (N3324, N3312, N2821, N2026, N3246);
xor XOR2 (N3325, N3313, N1847);
buf BUF1 (N3326, N3304);
and AND2 (N3327, N3325, N2448);
not NOT1 (N3328, N3322);
or OR3 (N3329, N3324, N2286, N2425);
xor XOR2 (N3330, N3317, N107);
not NOT1 (N3331, N3319);
buf BUF1 (N3332, N3315);
and AND4 (N3333, N3332, N1863, N410, N1275);
or OR3 (N3334, N3331, N447, N1747);
buf BUF1 (N3335, N3329);
not NOT1 (N3336, N3323);
or OR3 (N3337, N3336, N47, N780);
not NOT1 (N3338, N3326);
and AND4 (N3339, N3327, N366, N345, N2972);
and AND4 (N3340, N3321, N76, N2958, N765);
not NOT1 (N3341, N3334);
or OR2 (N3342, N3320, N3241);
not NOT1 (N3343, N3333);
xor XOR2 (N3344, N3330, N851);
or OR2 (N3345, N3342, N2364);
xor XOR2 (N3346, N3340, N2608);
nor NOR2 (N3347, N3345, N3015);
nor NOR4 (N3348, N3344, N2725, N2003, N1039);
buf BUF1 (N3349, N3341);
nand NAND2 (N3350, N3338, N1278);
buf BUF1 (N3351, N3349);
and AND2 (N3352, N3328, N2416);
nor NOR4 (N3353, N3351, N829, N679, N1137);
or OR4 (N3354, N3343, N162, N1529, N1212);
buf BUF1 (N3355, N3350);
not NOT1 (N3356, N3346);
and AND3 (N3357, N3348, N1203, N1756);
nand NAND4 (N3358, N3352, N2369, N1888, N2956);
not NOT1 (N3359, N3354);
or OR2 (N3360, N3356, N2743);
not NOT1 (N3361, N3358);
nor NOR2 (N3362, N3339, N2423);
and AND2 (N3363, N3361, N3321);
nor NOR3 (N3364, N3347, N3160, N2212);
nor NOR3 (N3365, N3337, N1001, N2078);
nor NOR3 (N3366, N3357, N1512, N1694);
xor XOR2 (N3367, N3362, N2387);
buf BUF1 (N3368, N3360);
and AND3 (N3369, N3366, N2010, N1676);
nand NAND4 (N3370, N3363, N2259, N1011, N741);
or OR3 (N3371, N3369, N2888, N3082);
buf BUF1 (N3372, N3365);
not NOT1 (N3373, N3355);
nand NAND3 (N3374, N3373, N667, N1419);
xor XOR2 (N3375, N3374, N1045);
not NOT1 (N3376, N3353);
buf BUF1 (N3377, N3372);
nand NAND2 (N3378, N3371, N2387);
not NOT1 (N3379, N3364);
and AND2 (N3380, N3368, N3023);
or OR4 (N3381, N3377, N2505, N145, N562);
not NOT1 (N3382, N3380);
buf BUF1 (N3383, N3381);
nand NAND2 (N3384, N3382, N3000);
or OR3 (N3385, N3379, N2649, N3100);
xor XOR2 (N3386, N3359, N1136);
not NOT1 (N3387, N3386);
not NOT1 (N3388, N3370);
xor XOR2 (N3389, N3378, N906);
or OR2 (N3390, N3385, N2133);
xor XOR2 (N3391, N3376, N578);
or OR2 (N3392, N3391, N386);
nor NOR3 (N3393, N3388, N639, N316);
or OR4 (N3394, N3383, N535, N37, N2388);
or OR3 (N3395, N3375, N2264, N3114);
not NOT1 (N3396, N3389);
xor XOR2 (N3397, N3394, N2562);
and AND2 (N3398, N3384, N2094);
xor XOR2 (N3399, N3398, N847);
not NOT1 (N3400, N3335);
buf BUF1 (N3401, N3399);
not NOT1 (N3402, N3392);
nand NAND4 (N3403, N3402, N1022, N2720, N1299);
or OR4 (N3404, N3401, N553, N59, N1329);
and AND3 (N3405, N3367, N2770, N3007);
xor XOR2 (N3406, N3404, N792);
xor XOR2 (N3407, N3396, N1342);
nor NOR2 (N3408, N3387, N100);
xor XOR2 (N3409, N3406, N633);
nand NAND4 (N3410, N3409, N2871, N2248, N241);
buf BUF1 (N3411, N3390);
xor XOR2 (N3412, N3393, N2827);
nand NAND2 (N3413, N3410, N3016);
nand NAND2 (N3414, N3403, N2271);
nor NOR4 (N3415, N3395, N1267, N193, N914);
nand NAND4 (N3416, N3397, N2896, N30, N2407);
nor NOR4 (N3417, N3415, N3318, N927, N2774);
nand NAND2 (N3418, N3414, N2771);
not NOT1 (N3419, N3405);
buf BUF1 (N3420, N3418);
not NOT1 (N3421, N3400);
not NOT1 (N3422, N3416);
nor NOR3 (N3423, N3422, N1787, N2694);
nand NAND3 (N3424, N3412, N921, N2361);
not NOT1 (N3425, N3413);
and AND3 (N3426, N3419, N2815, N2706);
xor XOR2 (N3427, N3424, N2821);
nor NOR3 (N3428, N3420, N2359, N1770);
nor NOR2 (N3429, N3407, N2217);
and AND2 (N3430, N3408, N943);
xor XOR2 (N3431, N3425, N1449);
buf BUF1 (N3432, N3426);
not NOT1 (N3433, N3411);
xor XOR2 (N3434, N3417, N1058);
and AND3 (N3435, N3431, N1670, N361);
nand NAND2 (N3436, N3423, N2643);
or OR3 (N3437, N3436, N1897, N2716);
not NOT1 (N3438, N3432);
xor XOR2 (N3439, N3433, N3398);
nor NOR4 (N3440, N3421, N2539, N2828, N2885);
and AND2 (N3441, N3440, N1025);
and AND4 (N3442, N3441, N1342, N1988, N1778);
not NOT1 (N3443, N3437);
nand NAND4 (N3444, N3442, N317, N1733, N2315);
and AND2 (N3445, N3430, N2297);
nor NOR4 (N3446, N3429, N1734, N2575, N3251);
xor XOR2 (N3447, N3434, N2612);
or OR4 (N3448, N3435, N8, N2790, N729);
or OR2 (N3449, N3439, N837);
and AND3 (N3450, N3428, N2314, N1315);
nand NAND2 (N3451, N3447, N1856);
xor XOR2 (N3452, N3450, N2917);
buf BUF1 (N3453, N3451);
buf BUF1 (N3454, N3448);
not NOT1 (N3455, N3427);
nor NOR4 (N3456, N3449, N2487, N102, N2548);
or OR3 (N3457, N3454, N2061, N814);
not NOT1 (N3458, N3456);
buf BUF1 (N3459, N3443);
and AND4 (N3460, N3444, N2183, N2473, N3259);
not NOT1 (N3461, N3457);
xor XOR2 (N3462, N3459, N3289);
or OR3 (N3463, N3460, N317, N1422);
or OR3 (N3464, N3446, N3278, N3104);
buf BUF1 (N3465, N3458);
or OR4 (N3466, N3455, N3177, N2016, N2662);
not NOT1 (N3467, N3438);
or OR2 (N3468, N3467, N1313);
not NOT1 (N3469, N3463);
not NOT1 (N3470, N3453);
not NOT1 (N3471, N3464);
not NOT1 (N3472, N3462);
nor NOR3 (N3473, N3445, N220, N932);
and AND3 (N3474, N3465, N881, N305);
xor XOR2 (N3475, N3466, N193);
not NOT1 (N3476, N3475);
or OR3 (N3477, N3468, N3009, N1426);
xor XOR2 (N3478, N3477, N2872);
nor NOR2 (N3479, N3472, N1046);
xor XOR2 (N3480, N3461, N3132);
buf BUF1 (N3481, N3476);
or OR4 (N3482, N3470, N2235, N2193, N1799);
buf BUF1 (N3483, N3479);
and AND2 (N3484, N3481, N2465);
nor NOR3 (N3485, N3471, N790, N516);
nor NOR2 (N3486, N3452, N2444);
nor NOR3 (N3487, N3469, N2702, N2656);
nand NAND4 (N3488, N3483, N3194, N1558, N2878);
nor NOR4 (N3489, N3474, N2506, N745, N3300);
buf BUF1 (N3490, N3485);
not NOT1 (N3491, N3480);
and AND3 (N3492, N3488, N2801, N2237);
or OR3 (N3493, N3482, N1799, N1583);
xor XOR2 (N3494, N3492, N36);
xor XOR2 (N3495, N3478, N603);
or OR4 (N3496, N3473, N3052, N1446, N2023);
nand NAND2 (N3497, N3486, N3343);
nor NOR2 (N3498, N3496, N3109);
nor NOR4 (N3499, N3490, N1433, N2359, N1875);
nor NOR4 (N3500, N3495, N1144, N3462, N838);
buf BUF1 (N3501, N3484);
nor NOR2 (N3502, N3499, N1641);
nor NOR3 (N3503, N3489, N1742, N3027);
buf BUF1 (N3504, N3500);
nor NOR3 (N3505, N3494, N1761, N2209);
not NOT1 (N3506, N3501);
not NOT1 (N3507, N3505);
or OR4 (N3508, N3487, N1777, N1751, N429);
xor XOR2 (N3509, N3504, N732);
nand NAND2 (N3510, N3506, N3045);
buf BUF1 (N3511, N3509);
buf BUF1 (N3512, N3497);
nor NOR4 (N3513, N3491, N615, N125, N3085);
buf BUF1 (N3514, N3510);
nor NOR4 (N3515, N3493, N3352, N1869, N1946);
not NOT1 (N3516, N3503);
and AND3 (N3517, N3514, N619, N3049);
nand NAND2 (N3518, N3512, N30);
nand NAND4 (N3519, N3516, N714, N3295, N1433);
nor NOR3 (N3520, N3498, N1668, N3188);
nand NAND4 (N3521, N3513, N791, N1465, N206);
nand NAND2 (N3522, N3520, N278);
and AND2 (N3523, N3518, N3075);
nor NOR2 (N3524, N3517, N830);
buf BUF1 (N3525, N3522);
nand NAND3 (N3526, N3525, N2220, N872);
not NOT1 (N3527, N3511);
and AND2 (N3528, N3502, N660);
not NOT1 (N3529, N3515);
buf BUF1 (N3530, N3527);
nor NOR3 (N3531, N3526, N603, N2922);
buf BUF1 (N3532, N3523);
not NOT1 (N3533, N3532);
xor XOR2 (N3534, N3531, N432);
or OR2 (N3535, N3534, N880);
and AND2 (N3536, N3528, N2282);
buf BUF1 (N3537, N3529);
nand NAND2 (N3538, N3537, N318);
or OR4 (N3539, N3533, N3104, N3270, N97);
nand NAND4 (N3540, N3519, N1835, N318, N1832);
nor NOR4 (N3541, N3521, N2383, N856, N1598);
nor NOR3 (N3542, N3508, N1739, N3470);
not NOT1 (N3543, N3530);
nor NOR2 (N3544, N3535, N2043);
not NOT1 (N3545, N3544);
buf BUF1 (N3546, N3539);
or OR2 (N3547, N3538, N3028);
nor NOR2 (N3548, N3536, N2724);
or OR2 (N3549, N3543, N2015);
buf BUF1 (N3550, N3547);
and AND2 (N3551, N3507, N467);
xor XOR2 (N3552, N3545, N2305);
or OR4 (N3553, N3552, N2123, N2877, N438);
buf BUF1 (N3554, N3553);
and AND2 (N3555, N3551, N3041);
not NOT1 (N3556, N3554);
not NOT1 (N3557, N3524);
xor XOR2 (N3558, N3550, N3508);
not NOT1 (N3559, N3556);
not NOT1 (N3560, N3541);
and AND4 (N3561, N3560, N885, N2754, N3398);
nand NAND2 (N3562, N3559, N1616);
or OR4 (N3563, N3558, N488, N2122, N3061);
or OR3 (N3564, N3561, N2076, N720);
buf BUF1 (N3565, N3563);
buf BUF1 (N3566, N3549);
not NOT1 (N3567, N3546);
or OR3 (N3568, N3540, N1270, N1109);
buf BUF1 (N3569, N3564);
xor XOR2 (N3570, N3557, N1128);
or OR3 (N3571, N3566, N3061, N178);
xor XOR2 (N3572, N3569, N2133);
not NOT1 (N3573, N3570);
buf BUF1 (N3574, N3573);
or OR3 (N3575, N3571, N2798, N1056);
xor XOR2 (N3576, N3575, N183);
and AND2 (N3577, N3555, N1192);
and AND2 (N3578, N3568, N3024);
not NOT1 (N3579, N3565);
and AND2 (N3580, N3577, N2346);
not NOT1 (N3581, N3572);
buf BUF1 (N3582, N3578);
nand NAND2 (N3583, N3574, N771);
xor XOR2 (N3584, N3580, N1729);
nor NOR2 (N3585, N3579, N2573);
and AND4 (N3586, N3548, N3101, N3087, N3207);
and AND4 (N3587, N3582, N3399, N1084, N1573);
nor NOR2 (N3588, N3576, N322);
buf BUF1 (N3589, N3585);
or OR3 (N3590, N3589, N1909, N2121);
nor NOR3 (N3591, N3583, N848, N3252);
not NOT1 (N3592, N3562);
xor XOR2 (N3593, N3592, N1990);
buf BUF1 (N3594, N3586);
buf BUF1 (N3595, N3591);
not NOT1 (N3596, N3567);
nor NOR3 (N3597, N3587, N1084, N3274);
nand NAND2 (N3598, N3588, N1416);
and AND3 (N3599, N3595, N3320, N3152);
or OR3 (N3600, N3593, N2017, N1051);
nand NAND4 (N3601, N3542, N2067, N2665, N678);
nand NAND3 (N3602, N3598, N1836, N2269);
nor NOR2 (N3603, N3590, N663);
nor NOR3 (N3604, N3581, N3313, N624);
nor NOR4 (N3605, N3600, N278, N3230, N2548);
or OR2 (N3606, N3601, N1550);
and AND3 (N3607, N3594, N3147, N2106);
and AND3 (N3608, N3607, N1488, N1365);
and AND3 (N3609, N3599, N2069, N154);
xor XOR2 (N3610, N3605, N1729);
nor NOR3 (N3611, N3597, N472, N2006);
xor XOR2 (N3612, N3610, N2126);
or OR4 (N3613, N3602, N2562, N2886, N2212);
xor XOR2 (N3614, N3611, N2576);
buf BUF1 (N3615, N3612);
nand NAND4 (N3616, N3606, N311, N3134, N2812);
xor XOR2 (N3617, N3615, N1624);
nor NOR3 (N3618, N3604, N2657, N1571);
and AND2 (N3619, N3617, N1180);
not NOT1 (N3620, N3584);
nor NOR2 (N3621, N3603, N2200);
buf BUF1 (N3622, N3613);
nor NOR3 (N3623, N3616, N1899, N3372);
and AND2 (N3624, N3596, N2903);
and AND3 (N3625, N3624, N3261, N3350);
nor NOR3 (N3626, N3623, N2435, N1606);
nor NOR3 (N3627, N3626, N2965, N328);
not NOT1 (N3628, N3621);
not NOT1 (N3629, N3627);
or OR3 (N3630, N3622, N219, N3558);
not NOT1 (N3631, N3614);
and AND3 (N3632, N3620, N469, N3578);
and AND2 (N3633, N3618, N2317);
buf BUF1 (N3634, N3609);
xor XOR2 (N3635, N3633, N2513);
nor NOR4 (N3636, N3625, N1121, N15, N2831);
buf BUF1 (N3637, N3628);
buf BUF1 (N3638, N3632);
not NOT1 (N3639, N3608);
or OR3 (N3640, N3637, N686, N2197);
buf BUF1 (N3641, N3635);
not NOT1 (N3642, N3629);
xor XOR2 (N3643, N3642, N1947);
not NOT1 (N3644, N3619);
nor NOR2 (N3645, N3631, N959);
or OR3 (N3646, N3636, N1152, N1736);
xor XOR2 (N3647, N3643, N742);
nand NAND4 (N3648, N3641, N968, N3106, N1601);
not NOT1 (N3649, N3634);
or OR3 (N3650, N3649, N2424, N246);
and AND3 (N3651, N3640, N2850, N1220);
buf BUF1 (N3652, N3645);
xor XOR2 (N3653, N3639, N1531);
and AND3 (N3654, N3630, N2403, N681);
not NOT1 (N3655, N3651);
not NOT1 (N3656, N3653);
buf BUF1 (N3657, N3648);
nor NOR4 (N3658, N3656, N1142, N646, N1937);
and AND2 (N3659, N3650, N2520);
or OR4 (N3660, N3647, N1409, N3402, N3520);
not NOT1 (N3661, N3638);
xor XOR2 (N3662, N3646, N2876);
nor NOR3 (N3663, N3654, N425, N2619);
buf BUF1 (N3664, N3655);
and AND2 (N3665, N3662, N2921);
nor NOR2 (N3666, N3661, N865);
xor XOR2 (N3667, N3660, N3217);
and AND2 (N3668, N3667, N3625);
and AND4 (N3669, N3652, N1757, N2171, N1969);
or OR2 (N3670, N3669, N3436);
buf BUF1 (N3671, N3665);
or OR3 (N3672, N3644, N1895, N1063);
and AND4 (N3673, N3670, N2084, N3070, N168);
nand NAND4 (N3674, N3663, N1945, N2181, N1550);
buf BUF1 (N3675, N3666);
or OR2 (N3676, N3671, N3331);
buf BUF1 (N3677, N3657);
buf BUF1 (N3678, N3658);
or OR3 (N3679, N3668, N2741, N2905);
or OR2 (N3680, N3673, N2062);
xor XOR2 (N3681, N3659, N2707);
and AND3 (N3682, N3678, N3311, N55);
buf BUF1 (N3683, N3682);
xor XOR2 (N3684, N3679, N990);
and AND2 (N3685, N3683, N3509);
or OR4 (N3686, N3677, N1246, N3471, N1384);
nand NAND2 (N3687, N3672, N3183);
and AND3 (N3688, N3681, N2474, N514);
not NOT1 (N3689, N3664);
xor XOR2 (N3690, N3674, N1581);
nor NOR3 (N3691, N3685, N1278, N2934);
nor NOR4 (N3692, N3689, N3167, N2332, N1171);
and AND3 (N3693, N3675, N1180, N2066);
or OR2 (N3694, N3690, N2244);
nor NOR3 (N3695, N3676, N2456, N3142);
or OR2 (N3696, N3694, N2952);
not NOT1 (N3697, N3696);
and AND4 (N3698, N3697, N41, N1977, N2229);
or OR3 (N3699, N3692, N2949, N3438);
and AND3 (N3700, N3687, N3382, N5);
xor XOR2 (N3701, N3699, N2025);
or OR3 (N3702, N3695, N1117, N1699);
nor NOR2 (N3703, N3698, N2125);
not NOT1 (N3704, N3691);
or OR2 (N3705, N3693, N3112);
nand NAND3 (N3706, N3701, N1169, N3572);
nand NAND4 (N3707, N3684, N523, N1415, N2102);
not NOT1 (N3708, N3707);
not NOT1 (N3709, N3686);
buf BUF1 (N3710, N3680);
or OR4 (N3711, N3705, N2154, N756, N1147);
or OR2 (N3712, N3710, N2475);
buf BUF1 (N3713, N3709);
or OR2 (N3714, N3704, N2392);
nor NOR3 (N3715, N3688, N507, N2017);
or OR3 (N3716, N3700, N2735, N3574);
or OR3 (N3717, N3715, N681, N2136);
nand NAND2 (N3718, N3708, N2692);
nor NOR4 (N3719, N3702, N1534, N2099, N1657);
or OR4 (N3720, N3714, N69, N1500, N1337);
nand NAND3 (N3721, N3716, N640, N832);
xor XOR2 (N3722, N3711, N665);
nor NOR2 (N3723, N3719, N3384);
buf BUF1 (N3724, N3703);
nand NAND2 (N3725, N3712, N3043);
nor NOR4 (N3726, N3722, N725, N2894, N3020);
and AND4 (N3727, N3723, N2168, N3385, N1937);
xor XOR2 (N3728, N3718, N2462);
nor NOR4 (N3729, N3724, N3507, N2899, N229);
not NOT1 (N3730, N3706);
and AND3 (N3731, N3730, N1329, N474);
or OR3 (N3732, N3721, N1120, N346);
and AND3 (N3733, N3726, N1625, N2048);
or OR4 (N3734, N3717, N809, N1357, N750);
and AND2 (N3735, N3728, N3709);
or OR4 (N3736, N3729, N776, N1987, N2006);
not NOT1 (N3737, N3732);
nor NOR2 (N3738, N3725, N971);
not NOT1 (N3739, N3738);
nand NAND2 (N3740, N3739, N756);
and AND2 (N3741, N3713, N1613);
and AND3 (N3742, N3740, N2468, N467);
nor NOR2 (N3743, N3733, N1392);
not NOT1 (N3744, N3737);
xor XOR2 (N3745, N3720, N716);
or OR4 (N3746, N3743, N2255, N2862, N2345);
nor NOR3 (N3747, N3742, N77, N764);
nor NOR4 (N3748, N3741, N956, N2252, N1241);
and AND3 (N3749, N3727, N2859, N693);
buf BUF1 (N3750, N3731);
nor NOR4 (N3751, N3744, N1948, N1757, N2193);
nand NAND2 (N3752, N3747, N2134);
and AND4 (N3753, N3750, N475, N2234, N1856);
not NOT1 (N3754, N3734);
nand NAND2 (N3755, N3746, N169);
or OR3 (N3756, N3745, N740, N1645);
buf BUF1 (N3757, N3751);
nor NOR3 (N3758, N3736, N1445, N3118);
xor XOR2 (N3759, N3749, N1019);
not NOT1 (N3760, N3759);
or OR2 (N3761, N3755, N1434);
buf BUF1 (N3762, N3748);
xor XOR2 (N3763, N3760, N2780);
nand NAND3 (N3764, N3756, N2986, N673);
nor NOR2 (N3765, N3764, N2295);
nor NOR3 (N3766, N3757, N1720, N2211);
nand NAND2 (N3767, N3765, N2233);
buf BUF1 (N3768, N3766);
xor XOR2 (N3769, N3763, N3069);
nor NOR4 (N3770, N3758, N1537, N2867, N1327);
xor XOR2 (N3771, N3753, N3185);
or OR3 (N3772, N3768, N2816, N2230);
buf BUF1 (N3773, N3772);
buf BUF1 (N3774, N3754);
not NOT1 (N3775, N3761);
or OR4 (N3776, N3752, N815, N1937, N535);
buf BUF1 (N3777, N3767);
or OR3 (N3778, N3769, N3623, N667);
or OR4 (N3779, N3776, N3063, N1787, N2812);
not NOT1 (N3780, N3778);
buf BUF1 (N3781, N3775);
nand NAND4 (N3782, N3780, N738, N3451, N3408);
buf BUF1 (N3783, N3782);
nor NOR4 (N3784, N3781, N2928, N1028, N277);
and AND3 (N3785, N3735, N3671, N2688);
not NOT1 (N3786, N3773);
or OR3 (N3787, N3785, N3433, N3521);
or OR3 (N3788, N3787, N2607, N2289);
buf BUF1 (N3789, N3788);
nor NOR4 (N3790, N3789, N2187, N2040, N2644);
nand NAND2 (N3791, N3771, N3123);
buf BUF1 (N3792, N3786);
or OR2 (N3793, N3779, N3772);
xor XOR2 (N3794, N3792, N2995);
xor XOR2 (N3795, N3762, N2945);
xor XOR2 (N3796, N3795, N3732);
nand NAND2 (N3797, N3784, N1817);
nand NAND2 (N3798, N3777, N1038);
nand NAND2 (N3799, N3798, N1143);
nor NOR2 (N3800, N3793, N3329);
and AND4 (N3801, N3774, N2046, N2547, N310);
xor XOR2 (N3802, N3790, N3480);
nand NAND3 (N3803, N3770, N2273, N1099);
and AND2 (N3804, N3797, N624);
not NOT1 (N3805, N3791);
nand NAND4 (N3806, N3802, N2846, N630, N67);
or OR4 (N3807, N3801, N2467, N2958, N2150);
nand NAND3 (N3808, N3803, N1288, N1607);
or OR2 (N3809, N3806, N2353);
not NOT1 (N3810, N3783);
or OR2 (N3811, N3810, N2271);
and AND3 (N3812, N3799, N1724, N3219);
and AND4 (N3813, N3809, N81, N890, N3013);
not NOT1 (N3814, N3800);
xor XOR2 (N3815, N3796, N1405);
nand NAND4 (N3816, N3814, N2183, N2362, N2727);
not NOT1 (N3817, N3804);
and AND2 (N3818, N3813, N2947);
not NOT1 (N3819, N3818);
buf BUF1 (N3820, N3808);
not NOT1 (N3821, N3815);
nor NOR3 (N3822, N3811, N2191, N1626);
not NOT1 (N3823, N3812);
not NOT1 (N3824, N3823);
and AND2 (N3825, N3819, N210);
not NOT1 (N3826, N3817);
not NOT1 (N3827, N3794);
xor XOR2 (N3828, N3827, N978);
xor XOR2 (N3829, N3824, N1605);
nor NOR2 (N3830, N3820, N1301);
buf BUF1 (N3831, N3829);
xor XOR2 (N3832, N3805, N489);
xor XOR2 (N3833, N3807, N835);
nor NOR3 (N3834, N3832, N33, N2986);
nand NAND3 (N3835, N3834, N3637, N2441);
buf BUF1 (N3836, N3822);
buf BUF1 (N3837, N3836);
not NOT1 (N3838, N3821);
xor XOR2 (N3839, N3816, N3794);
nand NAND3 (N3840, N3830, N3484, N2183);
or OR2 (N3841, N3825, N2201);
or OR2 (N3842, N3835, N2347);
nor NOR4 (N3843, N3842, N50, N1959, N1452);
not NOT1 (N3844, N3838);
nor NOR2 (N3845, N3839, N2080);
nor NOR4 (N3846, N3837, N182, N1915, N30);
xor XOR2 (N3847, N3841, N1200);
buf BUF1 (N3848, N3847);
nand NAND2 (N3849, N3844, N2023);
nor NOR4 (N3850, N3848, N3345, N990, N2087);
and AND3 (N3851, N3849, N2425, N3842);
nor NOR4 (N3852, N3833, N1923, N1014, N2977);
nand NAND2 (N3853, N3852, N644);
buf BUF1 (N3854, N3853);
xor XOR2 (N3855, N3826, N2206);
not NOT1 (N3856, N3854);
or OR3 (N3857, N3840, N1090, N665);
or OR4 (N3858, N3851, N1896, N1882, N3038);
nand NAND4 (N3859, N3856, N791, N3147, N1295);
and AND3 (N3860, N3859, N2297, N369);
not NOT1 (N3861, N3831);
nor NOR4 (N3862, N3860, N1706, N1154, N1792);
or OR2 (N3863, N3828, N2048);
or OR3 (N3864, N3858, N3740, N1518);
nand NAND3 (N3865, N3861, N3756, N2988);
nor NOR2 (N3866, N3857, N3262);
nand NAND2 (N3867, N3845, N390);
nor NOR2 (N3868, N3855, N3579);
buf BUF1 (N3869, N3843);
or OR3 (N3870, N3869, N2966, N2663);
xor XOR2 (N3871, N3865, N311);
or OR2 (N3872, N3868, N580);
nand NAND3 (N3873, N3850, N2913, N3299);
or OR4 (N3874, N3846, N3322, N775, N3528);
xor XOR2 (N3875, N3871, N1585);
nor NOR2 (N3876, N3866, N3254);
nand NAND2 (N3877, N3872, N1514);
xor XOR2 (N3878, N3876, N1384);
nand NAND4 (N3879, N3875, N54, N2987, N778);
or OR2 (N3880, N3862, N3773);
nand NAND3 (N3881, N3863, N3045, N3846);
or OR2 (N3882, N3874, N3657);
nor NOR3 (N3883, N3864, N1288, N1308);
nand NAND4 (N3884, N3867, N1250, N1983, N272);
nor NOR3 (N3885, N3882, N92, N3523);
not NOT1 (N3886, N3873);
xor XOR2 (N3887, N3885, N1030);
nand NAND4 (N3888, N3887, N1390, N2435, N303);
not NOT1 (N3889, N3879);
not NOT1 (N3890, N3870);
and AND4 (N3891, N3888, N2731, N2987, N1494);
nand NAND2 (N3892, N3886, N3746);
xor XOR2 (N3893, N3889, N2594);
and AND2 (N3894, N3880, N919);
or OR2 (N3895, N3890, N3100);
nor NOR3 (N3896, N3895, N3459, N1788);
xor XOR2 (N3897, N3878, N391);
nor NOR2 (N3898, N3891, N2737);
nor NOR4 (N3899, N3883, N3461, N1087, N3808);
and AND2 (N3900, N3881, N2509);
buf BUF1 (N3901, N3900);
and AND2 (N3902, N3899, N2187);
buf BUF1 (N3903, N3894);
xor XOR2 (N3904, N3877, N657);
buf BUF1 (N3905, N3902);
buf BUF1 (N3906, N3898);
buf BUF1 (N3907, N3893);
nand NAND2 (N3908, N3897, N1314);
or OR4 (N3909, N3905, N104, N2019, N1547);
nand NAND4 (N3910, N3892, N2099, N862, N789);
not NOT1 (N3911, N3896);
or OR4 (N3912, N3910, N3376, N2114, N1998);
nand NAND4 (N3913, N3909, N2073, N2983, N3123);
xor XOR2 (N3914, N3907, N499);
nor NOR3 (N3915, N3913, N243, N2659);
nor NOR3 (N3916, N3901, N1842, N1794);
buf BUF1 (N3917, N3916);
xor XOR2 (N3918, N3908, N1186);
and AND2 (N3919, N3915, N2909);
not NOT1 (N3920, N3911);
nand NAND3 (N3921, N3912, N194, N2265);
nand NAND4 (N3922, N3921, N3775, N2992, N2284);
and AND2 (N3923, N3884, N3649);
nand NAND3 (N3924, N3919, N1556, N2526);
and AND2 (N3925, N3906, N2974);
not NOT1 (N3926, N3914);
nand NAND3 (N3927, N3925, N2359, N3651);
nand NAND4 (N3928, N3922, N1231, N1620, N2861);
nor NOR4 (N3929, N3904, N272, N2061, N2354);
or OR3 (N3930, N3929, N626, N3800);
nand NAND3 (N3931, N3928, N896, N1485);
nand NAND3 (N3932, N3903, N2297, N1523);
and AND2 (N3933, N3920, N3256);
nand NAND3 (N3934, N3918, N3174, N2684);
xor XOR2 (N3935, N3934, N1985);
or OR4 (N3936, N3935, N2921, N1997, N335);
buf BUF1 (N3937, N3936);
and AND2 (N3938, N3917, N2048);
nand NAND2 (N3939, N3924, N1106);
not NOT1 (N3940, N3938);
or OR2 (N3941, N3940, N1744);
nor NOR2 (N3942, N3931, N2520);
buf BUF1 (N3943, N3927);
buf BUF1 (N3944, N3937);
or OR2 (N3945, N3926, N270);
and AND2 (N3946, N3939, N1597);
buf BUF1 (N3947, N3943);
xor XOR2 (N3948, N3946, N3516);
nand NAND3 (N3949, N3932, N1182, N3362);
nand NAND3 (N3950, N3942, N1822, N964);
nor NOR4 (N3951, N3949, N2173, N3022, N3052);
or OR2 (N3952, N3930, N1903);
not NOT1 (N3953, N3952);
and AND4 (N3954, N3941, N2920, N2386, N3236);
buf BUF1 (N3955, N3923);
or OR2 (N3956, N3948, N870);
xor XOR2 (N3957, N3947, N2652);
and AND4 (N3958, N3957, N2548, N3221, N3950);
nand NAND4 (N3959, N3527, N26, N2754, N2868);
nor NOR3 (N3960, N3945, N3290, N3438);
nand NAND3 (N3961, N3933, N2832, N3725);
nand NAND4 (N3962, N3961, N3614, N2940, N878);
nand NAND2 (N3963, N3944, N2196);
and AND4 (N3964, N3963, N2449, N1093, N3338);
buf BUF1 (N3965, N3958);
buf BUF1 (N3966, N3962);
nand NAND2 (N3967, N3955, N3331);
and AND4 (N3968, N3956, N3658, N1444, N492);
or OR3 (N3969, N3953, N3406, N821);
and AND4 (N3970, N3951, N1790, N3494, N1064);
nand NAND2 (N3971, N3970, N3719);
nor NOR3 (N3972, N3960, N563, N1155);
buf BUF1 (N3973, N3964);
xor XOR2 (N3974, N3971, N1527);
and AND2 (N3975, N3972, N2699);
or OR2 (N3976, N3966, N3507);
nand NAND3 (N3977, N3974, N882, N927);
xor XOR2 (N3978, N3976, N2743);
or OR4 (N3979, N3977, N3341, N1953, N1215);
not NOT1 (N3980, N3975);
nor NOR3 (N3981, N3954, N2378, N1595);
not NOT1 (N3982, N3978);
buf BUF1 (N3983, N3979);
nand NAND4 (N3984, N3959, N1549, N1246, N3561);
nand NAND4 (N3985, N3983, N2437, N497, N1803);
nor NOR3 (N3986, N3984, N3070, N3621);
nand NAND3 (N3987, N3965, N3931, N2270);
or OR2 (N3988, N3982, N855);
nand NAND2 (N3989, N3987, N1621);
or OR2 (N3990, N3981, N3083);
buf BUF1 (N3991, N3985);
nor NOR3 (N3992, N3969, N2069, N867);
nor NOR2 (N3993, N3980, N2295);
buf BUF1 (N3994, N3991);
nor NOR4 (N3995, N3988, N1473, N2559, N2238);
not NOT1 (N3996, N3973);
nand NAND4 (N3997, N3989, N3035, N765, N749);
and AND3 (N3998, N3996, N1450, N2884);
nand NAND4 (N3999, N3994, N1528, N2313, N1549);
nand NAND2 (N4000, N3998, N558);
xor XOR2 (N4001, N3995, N959);
nand NAND4 (N4002, N3986, N1223, N843, N2656);
and AND4 (N4003, N3993, N1216, N33, N1854);
or OR3 (N4004, N4002, N628, N2459);
buf BUF1 (N4005, N3992);
not NOT1 (N4006, N3968);
nand NAND4 (N4007, N4004, N704, N1094, N2197);
and AND4 (N4008, N4003, N598, N3455, N1865);
xor XOR2 (N4009, N4005, N3914);
xor XOR2 (N4010, N3997, N917);
or OR4 (N4011, N4006, N3789, N513, N1935);
xor XOR2 (N4012, N4010, N99);
and AND2 (N4013, N4009, N3142);
buf BUF1 (N4014, N4013);
nor NOR2 (N4015, N4008, N3772);
and AND4 (N4016, N4014, N1926, N3580, N3988);
not NOT1 (N4017, N3990);
nor NOR4 (N4018, N3967, N3182, N1598, N2778);
nor NOR4 (N4019, N4017, N320, N2010, N2518);
not NOT1 (N4020, N4019);
nand NAND3 (N4021, N4016, N2603, N2799);
buf BUF1 (N4022, N4018);
buf BUF1 (N4023, N4022);
nand NAND3 (N4024, N4021, N1925, N1974);
not NOT1 (N4025, N3999);
nand NAND3 (N4026, N4025, N1122, N1497);
nand NAND2 (N4027, N4011, N1861);
not NOT1 (N4028, N4020);
and AND4 (N4029, N4026, N3351, N926, N3966);
buf BUF1 (N4030, N4012);
not NOT1 (N4031, N4000);
and AND4 (N4032, N4031, N3583, N485, N2021);
nor NOR2 (N4033, N4027, N451);
nor NOR3 (N4034, N4001, N216, N669);
buf BUF1 (N4035, N4028);
not NOT1 (N4036, N4029);
not NOT1 (N4037, N4036);
nor NOR3 (N4038, N4030, N576, N3345);
buf BUF1 (N4039, N4032);
nor NOR4 (N4040, N4037, N7, N3885, N1623);
or OR2 (N4041, N4034, N2828);
or OR3 (N4042, N4023, N1316, N1886);
buf BUF1 (N4043, N4040);
nor NOR3 (N4044, N4007, N2918, N1275);
not NOT1 (N4045, N4044);
xor XOR2 (N4046, N4038, N4031);
and AND4 (N4047, N4046, N687, N2065, N3408);
xor XOR2 (N4048, N4039, N2097);
and AND2 (N4049, N4043, N333);
and AND4 (N4050, N4015, N3678, N1550, N1364);
not NOT1 (N4051, N4033);
and AND2 (N4052, N4049, N3465);
buf BUF1 (N4053, N4042);
nor NOR2 (N4054, N4035, N2500);
buf BUF1 (N4055, N4053);
not NOT1 (N4056, N4054);
nor NOR2 (N4057, N4041, N3266);
or OR4 (N4058, N4048, N33, N2528, N3896);
buf BUF1 (N4059, N4045);
xor XOR2 (N4060, N4055, N2528);
or OR2 (N4061, N4058, N2678);
not NOT1 (N4062, N4060);
buf BUF1 (N4063, N4050);
and AND4 (N4064, N4063, N2165, N235, N274);
or OR2 (N4065, N4056, N3767);
buf BUF1 (N4066, N4065);
xor XOR2 (N4067, N4059, N2086);
nand NAND3 (N4068, N4061, N1370, N3430);
and AND2 (N4069, N4047, N382);
xor XOR2 (N4070, N4062, N326);
xor XOR2 (N4071, N4068, N3901);
nand NAND2 (N4072, N4064, N2186);
or OR3 (N4073, N4071, N2218, N2686);
xor XOR2 (N4074, N4069, N4007);
nand NAND3 (N4075, N4052, N3954, N814);
xor XOR2 (N4076, N4074, N2877);
not NOT1 (N4077, N4024);
not NOT1 (N4078, N4072);
xor XOR2 (N4079, N4051, N2418);
not NOT1 (N4080, N4077);
xor XOR2 (N4081, N4079, N1158);
and AND4 (N4082, N4070, N3313, N2596, N1520);
not NOT1 (N4083, N4080);
buf BUF1 (N4084, N4081);
nand NAND4 (N4085, N4067, N823, N739, N1038);
and AND3 (N4086, N4057, N1554, N1166);
buf BUF1 (N4087, N4083);
nor NOR2 (N4088, N4085, N140);
or OR2 (N4089, N4078, N3563);
buf BUF1 (N4090, N4073);
nor NOR2 (N4091, N4076, N652);
or OR3 (N4092, N4066, N526, N2890);
xor XOR2 (N4093, N4086, N2620);
xor XOR2 (N4094, N4082, N3555);
not NOT1 (N4095, N4087);
or OR4 (N4096, N4091, N569, N3404, N922);
nand NAND3 (N4097, N4089, N2175, N661);
nand NAND3 (N4098, N4093, N3213, N3176);
nor NOR4 (N4099, N4090, N1687, N2545, N2706);
nand NAND3 (N4100, N4099, N1660, N2142);
buf BUF1 (N4101, N4088);
or OR4 (N4102, N4094, N1765, N3979, N2437);
and AND4 (N4103, N4075, N1104, N3369, N2330);
buf BUF1 (N4104, N4101);
nand NAND3 (N4105, N4103, N1909, N179);
or OR2 (N4106, N4096, N2311);
not NOT1 (N4107, N4104);
nor NOR4 (N4108, N4084, N1157, N1471, N1270);
nand NAND2 (N4109, N4106, N1445);
or OR3 (N4110, N4107, N2389, N583);
buf BUF1 (N4111, N4097);
buf BUF1 (N4112, N4110);
and AND3 (N4113, N4095, N3121, N327);
xor XOR2 (N4114, N4098, N1904);
nor NOR2 (N4115, N4109, N1354);
buf BUF1 (N4116, N4102);
not NOT1 (N4117, N4105);
or OR3 (N4118, N4108, N2437, N386);
not NOT1 (N4119, N4115);
nor NOR3 (N4120, N4116, N3228, N2007);
xor XOR2 (N4121, N4117, N769);
xor XOR2 (N4122, N4111, N4029);
or OR4 (N4123, N4119, N2659, N575, N639);
or OR2 (N4124, N4122, N3835);
and AND4 (N4125, N4112, N3539, N1612, N1948);
xor XOR2 (N4126, N4092, N841);
nor NOR3 (N4127, N4124, N3023, N1242);
not NOT1 (N4128, N4121);
nand NAND3 (N4129, N4125, N2519, N4051);
not NOT1 (N4130, N4128);
nand NAND4 (N4131, N4118, N1330, N2613, N1704);
xor XOR2 (N4132, N4123, N1008);
and AND4 (N4133, N4131, N2679, N4061, N3392);
xor XOR2 (N4134, N4129, N454);
buf BUF1 (N4135, N4113);
and AND4 (N4136, N4126, N754, N3150, N1564);
nor NOR3 (N4137, N4135, N1773, N2270);
nand NAND3 (N4138, N4100, N1191, N1152);
and AND4 (N4139, N4134, N2436, N2803, N2890);
buf BUF1 (N4140, N4114);
or OR3 (N4141, N4133, N3943, N3952);
xor XOR2 (N4142, N4141, N2879);
buf BUF1 (N4143, N4139);
nor NOR3 (N4144, N4143, N1155, N192);
not NOT1 (N4145, N4138);
nand NAND4 (N4146, N4127, N3143, N2307, N2174);
nor NOR4 (N4147, N4120, N3974, N989, N1958);
buf BUF1 (N4148, N4144);
or OR2 (N4149, N4132, N771);
buf BUF1 (N4150, N4140);
not NOT1 (N4151, N4142);
nand NAND3 (N4152, N4147, N2466, N3557);
buf BUF1 (N4153, N4152);
or OR2 (N4154, N4130, N1135);
and AND3 (N4155, N4153, N3894, N2725);
and AND4 (N4156, N4151, N346, N2722, N2156);
or OR3 (N4157, N4136, N3558, N708);
and AND3 (N4158, N4157, N3304, N433);
not NOT1 (N4159, N4154);
or OR4 (N4160, N4148, N2912, N1538, N3610);
buf BUF1 (N4161, N4155);
and AND4 (N4162, N4150, N54, N2724, N2003);
and AND3 (N4163, N4161, N3084, N2874);
xor XOR2 (N4164, N4149, N810);
and AND4 (N4165, N4163, N3301, N2224, N2413);
nor NOR4 (N4166, N4164, N40, N2242, N3743);
nor NOR2 (N4167, N4158, N2567);
or OR2 (N4168, N4159, N2695);
nor NOR3 (N4169, N4166, N1906, N2266);
buf BUF1 (N4170, N4165);
not NOT1 (N4171, N4137);
not NOT1 (N4172, N4168);
and AND2 (N4173, N4167, N3364);
or OR4 (N4174, N4146, N3095, N1063, N2613);
nand NAND2 (N4175, N4160, N400);
xor XOR2 (N4176, N4162, N2201);
or OR4 (N4177, N4145, N1407, N1478, N1099);
buf BUF1 (N4178, N4173);
or OR2 (N4179, N4170, N4100);
or OR2 (N4180, N4176, N2944);
nand NAND3 (N4181, N4180, N1974, N4095);
nand NAND2 (N4182, N4181, N3760);
nand NAND3 (N4183, N4169, N3838, N1197);
and AND4 (N4184, N4178, N1619, N1325, N2016);
and AND4 (N4185, N4175, N2048, N1639, N487);
nand NAND4 (N4186, N4156, N3363, N3152, N2112);
nand NAND4 (N4187, N4186, N1955, N2770, N25);
or OR4 (N4188, N4174, N490, N2838, N2158);
xor XOR2 (N4189, N4172, N3564);
and AND2 (N4190, N4179, N3372);
not NOT1 (N4191, N4182);
xor XOR2 (N4192, N4185, N2620);
not NOT1 (N4193, N4171);
and AND4 (N4194, N4188, N3773, N1065, N4168);
buf BUF1 (N4195, N4184);
buf BUF1 (N4196, N4189);
and AND3 (N4197, N4192, N1075, N287);
or OR2 (N4198, N4197, N3702);
not NOT1 (N4199, N4177);
or OR4 (N4200, N4194, N2166, N2330, N3814);
or OR3 (N4201, N4191, N4063, N2473);
nand NAND3 (N4202, N4196, N2535, N3335);
and AND3 (N4203, N4201, N3568, N3592);
nor NOR4 (N4204, N4187, N3411, N2623, N901);
buf BUF1 (N4205, N4199);
nand NAND4 (N4206, N4195, N3532, N2415, N2595);
xor XOR2 (N4207, N4183, N2148);
buf BUF1 (N4208, N4207);
or OR4 (N4209, N4204, N3439, N2925, N1397);
xor XOR2 (N4210, N4205, N2534);
xor XOR2 (N4211, N4190, N2552);
buf BUF1 (N4212, N4208);
xor XOR2 (N4213, N4193, N2748);
not NOT1 (N4214, N4209);
not NOT1 (N4215, N4211);
not NOT1 (N4216, N4200);
buf BUF1 (N4217, N4210);
or OR4 (N4218, N4216, N3388, N4111, N1767);
or OR3 (N4219, N4213, N3910, N3413);
buf BUF1 (N4220, N4219);
not NOT1 (N4221, N4206);
nor NOR3 (N4222, N4214, N3781, N2246);
buf BUF1 (N4223, N4222);
xor XOR2 (N4224, N4217, N1967);
xor XOR2 (N4225, N4198, N102);
not NOT1 (N4226, N4218);
nand NAND3 (N4227, N4220, N1222, N3248);
and AND2 (N4228, N4215, N2759);
nand NAND2 (N4229, N4203, N4047);
nand NAND4 (N4230, N4226, N1434, N2482, N3188);
xor XOR2 (N4231, N4223, N2677);
buf BUF1 (N4232, N4224);
nand NAND2 (N4233, N4229, N3195);
nor NOR4 (N4234, N4233, N4054, N195, N2116);
and AND3 (N4235, N4228, N1279, N1849);
nand NAND2 (N4236, N4225, N2236);
xor XOR2 (N4237, N4231, N1801);
xor XOR2 (N4238, N4236, N3808);
not NOT1 (N4239, N4221);
nand NAND2 (N4240, N4239, N2394);
or OR3 (N4241, N4235, N2833, N2698);
nand NAND3 (N4242, N4232, N128, N1705);
nand NAND2 (N4243, N4212, N3865);
nand NAND3 (N4244, N4241, N1905, N2501);
not NOT1 (N4245, N4234);
buf BUF1 (N4246, N4237);
nand NAND2 (N4247, N4230, N2179);
nor NOR2 (N4248, N4240, N2431);
nor NOR2 (N4249, N4248, N2767);
not NOT1 (N4250, N4249);
buf BUF1 (N4251, N4227);
buf BUF1 (N4252, N4250);
not NOT1 (N4253, N4238);
nand NAND3 (N4254, N4243, N2778, N2538);
nand NAND3 (N4255, N4246, N393, N786);
nor NOR2 (N4256, N4254, N3888);
nor NOR2 (N4257, N4252, N1126);
not NOT1 (N4258, N4253);
and AND3 (N4259, N4242, N2728, N356);
not NOT1 (N4260, N4255);
or OR4 (N4261, N4260, N2711, N3458, N3085);
buf BUF1 (N4262, N4257);
or OR4 (N4263, N4244, N4020, N2759, N2129);
and AND4 (N4264, N4202, N1068, N981, N3184);
not NOT1 (N4265, N4261);
xor XOR2 (N4266, N4259, N2648);
nor NOR2 (N4267, N4266, N3300);
not NOT1 (N4268, N4264);
not NOT1 (N4269, N4258);
nand NAND4 (N4270, N4245, N4248, N2357, N1566);
not NOT1 (N4271, N4267);
or OR2 (N4272, N4269, N790);
nor NOR4 (N4273, N4268, N1364, N1965, N292);
buf BUF1 (N4274, N4271);
nor NOR4 (N4275, N4263, N1869, N1657, N1645);
or OR2 (N4276, N4274, N407);
nand NAND4 (N4277, N4256, N1866, N3309, N2574);
and AND4 (N4278, N4275, N2630, N3989, N3689);
xor XOR2 (N4279, N4262, N3147);
xor XOR2 (N4280, N4272, N1440);
not NOT1 (N4281, N4265);
xor XOR2 (N4282, N4247, N3925);
or OR3 (N4283, N4277, N1663, N1571);
or OR2 (N4284, N4281, N625);
or OR2 (N4285, N4278, N1963);
xor XOR2 (N4286, N4283, N1449);
and AND2 (N4287, N4273, N2610);
nor NOR2 (N4288, N4280, N3804);
not NOT1 (N4289, N4286);
nor NOR3 (N4290, N4270, N2260, N3832);
nand NAND3 (N4291, N4276, N3411, N2298);
nand NAND3 (N4292, N4291, N2348, N3106);
nand NAND2 (N4293, N4251, N2435);
or OR2 (N4294, N4279, N3712);
buf BUF1 (N4295, N4290);
and AND2 (N4296, N4282, N403);
and AND2 (N4297, N4294, N341);
xor XOR2 (N4298, N4296, N124);
xor XOR2 (N4299, N4293, N2550);
xor XOR2 (N4300, N4289, N604);
not NOT1 (N4301, N4285);
buf BUF1 (N4302, N4299);
or OR3 (N4303, N4292, N3688, N2848);
or OR3 (N4304, N4287, N1287, N2817);
xor XOR2 (N4305, N4298, N3587);
xor XOR2 (N4306, N4305, N1471);
and AND4 (N4307, N4284, N2986, N230, N4275);
nor NOR4 (N4308, N4304, N3966, N3544, N3306);
or OR2 (N4309, N4297, N2439);
or OR3 (N4310, N4307, N2480, N1681);
nand NAND3 (N4311, N4309, N2047, N126);
and AND2 (N4312, N4308, N2502);
nor NOR3 (N4313, N4306, N793, N1769);
nand NAND2 (N4314, N4301, N2837);
and AND4 (N4315, N4311, N2497, N2293, N275);
nor NOR4 (N4316, N4302, N2982, N575, N3215);
nor NOR2 (N4317, N4303, N2451);
and AND3 (N4318, N4312, N3449, N227);
nand NAND2 (N4319, N4316, N1467);
or OR2 (N4320, N4315, N2019);
and AND2 (N4321, N4317, N3705);
nand NAND3 (N4322, N4295, N956, N228);
not NOT1 (N4323, N4320);
xor XOR2 (N4324, N4310, N359);
or OR2 (N4325, N4318, N1961);
and AND4 (N4326, N4319, N3762, N3210, N2777);
nand NAND3 (N4327, N4321, N694, N1245);
not NOT1 (N4328, N4327);
xor XOR2 (N4329, N4300, N2529);
nor NOR2 (N4330, N4288, N3769);
buf BUF1 (N4331, N4324);
nand NAND4 (N4332, N4322, N2237, N818, N321);
nor NOR3 (N4333, N4326, N199, N3612);
xor XOR2 (N4334, N4313, N2469);
xor XOR2 (N4335, N4330, N2902);
or OR4 (N4336, N4333, N3830, N3218, N2195);
and AND2 (N4337, N4334, N902);
xor XOR2 (N4338, N4331, N547);
xor XOR2 (N4339, N4332, N4282);
nand NAND2 (N4340, N4339, N2484);
and AND3 (N4341, N4325, N366, N1956);
nand NAND3 (N4342, N4336, N1639, N2301);
nor NOR4 (N4343, N4340, N1493, N3520, N1312);
or OR4 (N4344, N4323, N248, N1517, N2419);
or OR4 (N4345, N4329, N1539, N3885, N3880);
nand NAND4 (N4346, N4314, N2878, N1106, N692);
nand NAND3 (N4347, N4344, N3271, N202);
or OR4 (N4348, N4341, N4152, N1248, N725);
and AND4 (N4349, N4342, N164, N69, N619);
or OR4 (N4350, N4348, N1303, N1105, N97);
buf BUF1 (N4351, N4349);
buf BUF1 (N4352, N4335);
xor XOR2 (N4353, N4345, N14);
nand NAND3 (N4354, N4338, N4213, N1694);
or OR4 (N4355, N4343, N1641, N2436, N1114);
and AND4 (N4356, N4351, N2422, N1052, N2894);
not NOT1 (N4357, N4356);
or OR3 (N4358, N4353, N564, N2560);
nand NAND4 (N4359, N4347, N1568, N2095, N4205);
nand NAND4 (N4360, N4350, N2185, N3782, N3985);
and AND2 (N4361, N4354, N1624);
buf BUF1 (N4362, N4361);
nor NOR2 (N4363, N4359, N620);
and AND3 (N4364, N4346, N2422, N921);
or OR4 (N4365, N4364, N3384, N31, N462);
xor XOR2 (N4366, N4358, N3502);
and AND3 (N4367, N4363, N2074, N3840);
buf BUF1 (N4368, N4365);
nand NAND2 (N4369, N4362, N1617);
nor NOR3 (N4370, N4368, N2901, N3208);
and AND3 (N4371, N4328, N3162, N325);
nand NAND2 (N4372, N4366, N3910);
buf BUF1 (N4373, N4371);
buf BUF1 (N4374, N4370);
xor XOR2 (N4375, N4352, N349);
not NOT1 (N4376, N4375);
or OR2 (N4377, N4374, N3621);
or OR2 (N4378, N4355, N534);
xor XOR2 (N4379, N4367, N2471);
not NOT1 (N4380, N4357);
buf BUF1 (N4381, N4369);
or OR2 (N4382, N4381, N4027);
and AND4 (N4383, N4373, N3402, N212, N1134);
not NOT1 (N4384, N4337);
not NOT1 (N4385, N4383);
nor NOR3 (N4386, N4379, N4067, N2713);
and AND2 (N4387, N4372, N4129);
or OR3 (N4388, N4384, N1742, N1559);
not NOT1 (N4389, N4376);
nor NOR3 (N4390, N4386, N2657, N3809);
or OR3 (N4391, N4385, N843, N3517);
nor NOR3 (N4392, N4378, N575, N998);
buf BUF1 (N4393, N4389);
nand NAND4 (N4394, N4360, N1690, N3960, N2492);
nor NOR3 (N4395, N4380, N1300, N3514);
buf BUF1 (N4396, N4388);
buf BUF1 (N4397, N4393);
xor XOR2 (N4398, N4390, N3683);
or OR2 (N4399, N4392, N2663);
buf BUF1 (N4400, N4387);
xor XOR2 (N4401, N4391, N591);
nor NOR3 (N4402, N4382, N1973, N3753);
and AND4 (N4403, N4399, N401, N3183, N147);
and AND2 (N4404, N4403, N2352);
nand NAND2 (N4405, N4377, N2660);
nor NOR3 (N4406, N4400, N3972, N2548);
nor NOR4 (N4407, N4405, N2172, N256, N1847);
nand NAND4 (N4408, N4402, N4015, N3172, N2518);
nand NAND3 (N4409, N4395, N3320, N774);
nor NOR2 (N4410, N4401, N3698);
not NOT1 (N4411, N4394);
xor XOR2 (N4412, N4396, N1445);
xor XOR2 (N4413, N4398, N2166);
not NOT1 (N4414, N4412);
or OR4 (N4415, N4414, N3610, N2288, N1969);
and AND3 (N4416, N4407, N4213, N3769);
buf BUF1 (N4417, N4408);
buf BUF1 (N4418, N4411);
and AND4 (N4419, N4397, N4227, N1187, N2033);
xor XOR2 (N4420, N4416, N2063);
or OR3 (N4421, N4413, N995, N2782);
xor XOR2 (N4422, N4417, N4141);
nor NOR4 (N4423, N4415, N472, N4236, N2402);
nand NAND2 (N4424, N4420, N4256);
buf BUF1 (N4425, N4409);
not NOT1 (N4426, N4410);
or OR2 (N4427, N4406, N1159);
not NOT1 (N4428, N4426);
buf BUF1 (N4429, N4404);
buf BUF1 (N4430, N4428);
nor NOR2 (N4431, N4429, N3654);
not NOT1 (N4432, N4427);
xor XOR2 (N4433, N4430, N296);
nand NAND2 (N4434, N4431, N604);
or OR2 (N4435, N4419, N3630);
nand NAND2 (N4436, N4418, N3563);
nor NOR4 (N4437, N4434, N3545, N2604, N397);
or OR3 (N4438, N4436, N717, N1963);
xor XOR2 (N4439, N4424, N2434);
nor NOR3 (N4440, N4425, N2577, N227);
nand NAND4 (N4441, N4432, N4033, N3152, N3733);
nor NOR2 (N4442, N4423, N2276);
and AND3 (N4443, N4442, N2357, N355);
nor NOR2 (N4444, N4440, N2911);
xor XOR2 (N4445, N4435, N576);
nand NAND3 (N4446, N4444, N4211, N2427);
or OR4 (N4447, N4437, N705, N4036, N3653);
nand NAND4 (N4448, N4438, N2859, N1729, N801);
not NOT1 (N4449, N4439);
xor XOR2 (N4450, N4443, N1110);
xor XOR2 (N4451, N4446, N3723);
not NOT1 (N4452, N4449);
nand NAND2 (N4453, N4433, N2101);
xor XOR2 (N4454, N4447, N130);
and AND2 (N4455, N4448, N3020);
nand NAND3 (N4456, N4455, N2465, N791);
buf BUF1 (N4457, N4445);
or OR3 (N4458, N4451, N2205, N3096);
or OR2 (N4459, N4453, N288);
nor NOR2 (N4460, N4450, N3527);
not NOT1 (N4461, N4441);
and AND3 (N4462, N4422, N590, N647);
buf BUF1 (N4463, N4458);
nor NOR4 (N4464, N4462, N2376, N2016, N4434);
or OR4 (N4465, N4421, N4196, N4025, N1283);
nor NOR2 (N4466, N4457, N4356);
buf BUF1 (N4467, N4460);
or OR2 (N4468, N4461, N3228);
or OR3 (N4469, N4452, N467, N355);
not NOT1 (N4470, N4469);
buf BUF1 (N4471, N4456);
and AND3 (N4472, N4471, N1936, N613);
and AND4 (N4473, N4467, N1684, N2331, N973);
buf BUF1 (N4474, N4464);
and AND3 (N4475, N4465, N1918, N4127);
nand NAND4 (N4476, N4468, N176, N239, N2574);
nor NOR3 (N4477, N4454, N4179, N1877);
or OR3 (N4478, N4474, N2914, N3460);
or OR2 (N4479, N4463, N2292);
nand NAND4 (N4480, N4473, N2666, N3575, N51);
nor NOR4 (N4481, N4477, N4464, N2220, N3734);
or OR4 (N4482, N4478, N3657, N3438, N4215);
xor XOR2 (N4483, N4481, N2310);
not NOT1 (N4484, N4475);
and AND2 (N4485, N4459, N1194);
and AND3 (N4486, N4476, N2789, N3989);
or OR2 (N4487, N4479, N1683);
nor NOR2 (N4488, N4472, N2621);
or OR4 (N4489, N4486, N3260, N1490, N217);
or OR4 (N4490, N4489, N2474, N474, N3344);
nand NAND2 (N4491, N4490, N4142);
buf BUF1 (N4492, N4482);
buf BUF1 (N4493, N4492);
xor XOR2 (N4494, N4493, N1920);
or OR2 (N4495, N4470, N1332);
or OR2 (N4496, N4484, N2911);
or OR2 (N4497, N4480, N2241);
and AND3 (N4498, N4497, N2585, N3643);
not NOT1 (N4499, N4495);
or OR4 (N4500, N4496, N3448, N2532, N2273);
nand NAND4 (N4501, N4483, N1129, N1539, N1315);
nand NAND2 (N4502, N4488, N1707);
or OR4 (N4503, N4487, N4010, N2287, N2655);
and AND4 (N4504, N4501, N1695, N2158, N4039);
buf BUF1 (N4505, N4494);
and AND2 (N4506, N4498, N3866);
and AND2 (N4507, N4466, N87);
and AND2 (N4508, N4504, N2115);
not NOT1 (N4509, N4506);
nor NOR4 (N4510, N4503, N1405, N4400, N1250);
buf BUF1 (N4511, N4485);
xor XOR2 (N4512, N4499, N4510);
nor NOR3 (N4513, N1216, N4204, N921);
xor XOR2 (N4514, N4507, N2325);
or OR4 (N4515, N4502, N4338, N1124, N2902);
buf BUF1 (N4516, N4508);
not NOT1 (N4517, N4512);
buf BUF1 (N4518, N4491);
nor NOR4 (N4519, N4515, N4454, N3375, N3973);
xor XOR2 (N4520, N4518, N76);
nand NAND3 (N4521, N4500, N3277, N2795);
or OR2 (N4522, N4519, N4155);
xor XOR2 (N4523, N4505, N2911);
not NOT1 (N4524, N4523);
nor NOR4 (N4525, N4509, N2213, N239, N3647);
xor XOR2 (N4526, N4520, N709);
and AND3 (N4527, N4516, N3319, N145);
not NOT1 (N4528, N4511);
not NOT1 (N4529, N4525);
and AND4 (N4530, N4524, N3808, N4352, N2384);
nand NAND2 (N4531, N4517, N3769);
xor XOR2 (N4532, N4531, N310);
xor XOR2 (N4533, N4527, N2406);
nand NAND4 (N4534, N4513, N353, N4510, N4424);
or OR4 (N4535, N4526, N359, N168, N1074);
not NOT1 (N4536, N4530);
buf BUF1 (N4537, N4535);
nor NOR3 (N4538, N4522, N310, N3493);
nand NAND2 (N4539, N4537, N2927);
or OR2 (N4540, N4528, N1237);
not NOT1 (N4541, N4529);
xor XOR2 (N4542, N4540, N1235);
or OR4 (N4543, N4514, N3737, N1964, N3789);
nor NOR4 (N4544, N4538, N246, N1602, N4268);
xor XOR2 (N4545, N4539, N2597);
xor XOR2 (N4546, N4542, N4360);
nand NAND3 (N4547, N4534, N2987, N2794);
nand NAND2 (N4548, N4546, N3116);
xor XOR2 (N4549, N4543, N3757);
not NOT1 (N4550, N4536);
nor NOR2 (N4551, N4521, N2308);
and AND2 (N4552, N4544, N3);
or OR2 (N4553, N4532, N3123);
xor XOR2 (N4554, N4545, N168);
buf BUF1 (N4555, N4551);
and AND2 (N4556, N4550, N4277);
nor NOR4 (N4557, N4556, N3620, N2436, N3155);
nor NOR3 (N4558, N4547, N214, N3682);
xor XOR2 (N4559, N4549, N726);
buf BUF1 (N4560, N4557);
not NOT1 (N4561, N4558);
nor NOR2 (N4562, N4553, N4010);
or OR4 (N4563, N4561, N3040, N3959, N7);
and AND4 (N4564, N4548, N1599, N1117, N3865);
nand NAND4 (N4565, N4564, N2619, N492, N2277);
and AND2 (N4566, N4565, N1948);
xor XOR2 (N4567, N4533, N3771);
or OR3 (N4568, N4559, N538, N4539);
buf BUF1 (N4569, N4567);
or OR2 (N4570, N4562, N3529);
buf BUF1 (N4571, N4552);
or OR3 (N4572, N4566, N402, N1975);
nor NOR2 (N4573, N4572, N3718);
not NOT1 (N4574, N4573);
nand NAND4 (N4575, N4554, N2188, N181, N4394);
buf BUF1 (N4576, N4574);
buf BUF1 (N4577, N4569);
not NOT1 (N4578, N4560);
nand NAND4 (N4579, N4568, N120, N2824, N3348);
nor NOR4 (N4580, N4541, N2964, N2541, N411);
nor NOR3 (N4581, N4570, N806, N1555);
xor XOR2 (N4582, N4580, N1733);
nor NOR2 (N4583, N4578, N696);
or OR2 (N4584, N4579, N3813);
and AND2 (N4585, N4577, N2600);
or OR2 (N4586, N4585, N4557);
not NOT1 (N4587, N4583);
or OR3 (N4588, N4587, N1014, N2778);
nor NOR2 (N4589, N4584, N3360);
buf BUF1 (N4590, N4588);
buf BUF1 (N4591, N4586);
not NOT1 (N4592, N4571);
buf BUF1 (N4593, N4582);
and AND3 (N4594, N4592, N2332, N3206);
not NOT1 (N4595, N4590);
nand NAND2 (N4596, N4581, N1263);
nand NAND4 (N4597, N4589, N1217, N2095, N2322);
not NOT1 (N4598, N4575);
or OR2 (N4599, N4576, N2167);
or OR3 (N4600, N4594, N3320, N2059);
buf BUF1 (N4601, N4600);
nand NAND4 (N4602, N4598, N822, N547, N412);
or OR2 (N4603, N4601, N2548);
not NOT1 (N4604, N4563);
nand NAND4 (N4605, N4604, N1602, N113, N2455);
xor XOR2 (N4606, N4603, N875);
buf BUF1 (N4607, N4606);
buf BUF1 (N4608, N4599);
not NOT1 (N4609, N4602);
xor XOR2 (N4610, N4609, N4183);
and AND3 (N4611, N4593, N3137, N370);
nor NOR3 (N4612, N4597, N2671, N3262);
not NOT1 (N4613, N4611);
nor NOR4 (N4614, N4605, N4527, N248, N313);
buf BUF1 (N4615, N4607);
not NOT1 (N4616, N4612);
nor NOR4 (N4617, N4615, N4499, N2460, N4422);
buf BUF1 (N4618, N4617);
buf BUF1 (N4619, N4591);
and AND4 (N4620, N4613, N4547, N1075, N156);
buf BUF1 (N4621, N4610);
not NOT1 (N4622, N4555);
or OR4 (N4623, N4622, N4376, N3363, N1436);
or OR4 (N4624, N4621, N851, N3062, N607);
nor NOR4 (N4625, N4624, N4357, N244, N3453);
and AND2 (N4626, N4614, N4466);
or OR3 (N4627, N4618, N1207, N2030);
and AND4 (N4628, N4625, N1354, N2898, N2325);
nand NAND2 (N4629, N4623, N567);
nor NOR4 (N4630, N4596, N4094, N2857, N195);
nand NAND3 (N4631, N4616, N4563, N1995);
nand NAND3 (N4632, N4630, N3625, N2730);
nor NOR2 (N4633, N4619, N4228);
xor XOR2 (N4634, N4608, N3143);
not NOT1 (N4635, N4626);
xor XOR2 (N4636, N4595, N3523);
xor XOR2 (N4637, N4627, N2043);
nor NOR3 (N4638, N4632, N296, N117);
nor NOR4 (N4639, N4634, N1997, N3467, N3106);
buf BUF1 (N4640, N4633);
nand NAND2 (N4641, N4620, N4303);
or OR4 (N4642, N4641, N2135, N3163, N4037);
and AND2 (N4643, N4639, N2458);
and AND4 (N4644, N4629, N1447, N1643, N4419);
or OR2 (N4645, N4638, N94);
nand NAND3 (N4646, N4635, N3948, N193);
nor NOR2 (N4647, N4628, N1578);
xor XOR2 (N4648, N4643, N1875);
nand NAND3 (N4649, N4637, N1468, N5);
nand NAND3 (N4650, N4646, N3258, N299);
and AND4 (N4651, N4642, N3878, N4120, N1001);
not NOT1 (N4652, N4644);
nand NAND4 (N4653, N4640, N3877, N4221, N2680);
nand NAND4 (N4654, N4649, N4612, N2899, N1658);
xor XOR2 (N4655, N4650, N2394);
buf BUF1 (N4656, N4645);
or OR3 (N4657, N4651, N4526, N438);
not NOT1 (N4658, N4652);
and AND3 (N4659, N4654, N2907, N2730);
buf BUF1 (N4660, N4648);
buf BUF1 (N4661, N4647);
not NOT1 (N4662, N4655);
and AND3 (N4663, N4657, N3186, N3972);
or OR4 (N4664, N4663, N3442, N2038, N3333);
buf BUF1 (N4665, N4656);
nand NAND4 (N4666, N4661, N3229, N1385, N1267);
or OR4 (N4667, N4636, N2570, N4260, N1870);
and AND2 (N4668, N4662, N2273);
or OR4 (N4669, N4664, N47, N3001, N365);
buf BUF1 (N4670, N4669);
nand NAND4 (N4671, N4659, N4001, N3137, N1264);
xor XOR2 (N4672, N4666, N3120);
nor NOR4 (N4673, N4653, N812, N3663, N203);
and AND2 (N4674, N4665, N257);
xor XOR2 (N4675, N4672, N3228);
not NOT1 (N4676, N4658);
nand NAND3 (N4677, N4667, N3865, N2130);
and AND4 (N4678, N4660, N3409, N2162, N2391);
and AND3 (N4679, N4631, N345, N428);
nor NOR4 (N4680, N4675, N3682, N4136, N733);
and AND4 (N4681, N4680, N4121, N1676, N2857);
xor XOR2 (N4682, N4674, N258);
buf BUF1 (N4683, N4682);
xor XOR2 (N4684, N4671, N2816);
or OR3 (N4685, N4681, N3958, N2936);
or OR4 (N4686, N4685, N3048, N3176, N1132);
xor XOR2 (N4687, N4673, N3408);
buf BUF1 (N4688, N4686);
buf BUF1 (N4689, N4688);
not NOT1 (N4690, N4683);
or OR4 (N4691, N4678, N3032, N3599, N2596);
xor XOR2 (N4692, N4684, N4188);
or OR2 (N4693, N4670, N2950);
buf BUF1 (N4694, N4692);
nand NAND2 (N4695, N4694, N112);
nor NOR4 (N4696, N4690, N3012, N15, N809);
or OR3 (N4697, N4695, N1059, N2153);
and AND2 (N4698, N4677, N4564);
or OR4 (N4699, N4676, N2348, N1625, N297);
and AND3 (N4700, N4668, N1284, N2584);
and AND4 (N4701, N4696, N1855, N168, N2390);
nand NAND4 (N4702, N4687, N2124, N2041, N3496);
and AND3 (N4703, N4697, N1324, N1702);
nand NAND2 (N4704, N4689, N1502);
buf BUF1 (N4705, N4698);
not NOT1 (N4706, N4703);
buf BUF1 (N4707, N4704);
buf BUF1 (N4708, N4705);
or OR2 (N4709, N4699, N2930);
and AND3 (N4710, N4679, N1470, N3979);
and AND3 (N4711, N4708, N2775, N471);
nand NAND2 (N4712, N4702, N2338);
not NOT1 (N4713, N4709);
nor NOR3 (N4714, N4711, N1102, N3201);
and AND3 (N4715, N4706, N4223, N3914);
and AND2 (N4716, N4691, N2469);
not NOT1 (N4717, N4715);
and AND3 (N4718, N4714, N2150, N4358);
not NOT1 (N4719, N4717);
nor NOR3 (N4720, N4700, N3428, N69);
not NOT1 (N4721, N4710);
xor XOR2 (N4722, N4719, N2550);
nor NOR2 (N4723, N4707, N945);
nor NOR4 (N4724, N4716, N1616, N1041, N1146);
buf BUF1 (N4725, N4720);
buf BUF1 (N4726, N4712);
and AND2 (N4727, N4724, N2096);
nand NAND4 (N4728, N4726, N2563, N3184, N237);
or OR4 (N4729, N4722, N744, N3566, N2466);
nand NAND4 (N4730, N4721, N4269, N4206, N2746);
xor XOR2 (N4731, N4718, N4686);
not NOT1 (N4732, N4727);
nor NOR2 (N4733, N4729, N3368);
or OR3 (N4734, N4733, N2178, N3830);
xor XOR2 (N4735, N4734, N3987);
and AND3 (N4736, N4730, N3354, N3102);
xor XOR2 (N4737, N4732, N1123);
nor NOR2 (N4738, N4693, N1612);
not NOT1 (N4739, N4728);
buf BUF1 (N4740, N4739);
or OR4 (N4741, N4701, N3328, N3696, N4432);
not NOT1 (N4742, N4741);
nor NOR3 (N4743, N4742, N153, N2837);
and AND4 (N4744, N4735, N3861, N3494, N3934);
nand NAND2 (N4745, N4723, N3090);
not NOT1 (N4746, N4736);
nor NOR4 (N4747, N4740, N237, N3731, N2402);
nor NOR4 (N4748, N4731, N4006, N992, N1623);
not NOT1 (N4749, N4745);
not NOT1 (N4750, N4747);
nor NOR3 (N4751, N4713, N399, N1358);
not NOT1 (N4752, N4738);
xor XOR2 (N4753, N4737, N2965);
or OR2 (N4754, N4743, N2910);
and AND3 (N4755, N4754, N2375, N148);
nand NAND3 (N4756, N4744, N4152, N3796);
or OR4 (N4757, N4756, N2127, N1551, N107);
nor NOR4 (N4758, N4746, N3864, N2209, N4421);
nor NOR4 (N4759, N4758, N2199, N3456, N4577);
or OR4 (N4760, N4725, N3919, N1470, N3673);
nor NOR4 (N4761, N4759, N2238, N3699, N2526);
nor NOR2 (N4762, N4753, N3618);
buf BUF1 (N4763, N4757);
buf BUF1 (N4764, N4755);
buf BUF1 (N4765, N4760);
buf BUF1 (N4766, N4765);
nor NOR3 (N4767, N4749, N2203, N3524);
not NOT1 (N4768, N4764);
xor XOR2 (N4769, N4763, N3989);
nand NAND4 (N4770, N4751, N1794, N566, N3664);
nor NOR3 (N4771, N4761, N3016, N4369);
nand NAND4 (N4772, N4766, N3518, N1227, N3428);
not NOT1 (N4773, N4770);
nor NOR2 (N4774, N4767, N1998);
and AND4 (N4775, N4773, N629, N1252, N93);
and AND4 (N4776, N4775, N3804, N4103, N4355);
or OR4 (N4777, N4771, N3394, N2024, N3942);
nand NAND3 (N4778, N4772, N1514, N436);
buf BUF1 (N4779, N4750);
buf BUF1 (N4780, N4776);
buf BUF1 (N4781, N4748);
and AND3 (N4782, N4780, N4165, N3018);
xor XOR2 (N4783, N4782, N4061);
nand NAND3 (N4784, N4779, N2083, N3833);
and AND2 (N4785, N4781, N1656);
nand NAND4 (N4786, N4774, N2864, N1154, N2795);
not NOT1 (N4787, N4777);
or OR2 (N4788, N4786, N3032);
nor NOR4 (N4789, N4762, N58, N2863, N3007);
buf BUF1 (N4790, N4768);
nand NAND2 (N4791, N4789, N764);
buf BUF1 (N4792, N4752);
buf BUF1 (N4793, N4783);
not NOT1 (N4794, N4790);
not NOT1 (N4795, N4794);
and AND3 (N4796, N4778, N1011, N2674);
buf BUF1 (N4797, N4793);
xor XOR2 (N4798, N4795, N2588);
buf BUF1 (N4799, N4788);
and AND2 (N4800, N4799, N1442);
xor XOR2 (N4801, N4787, N2073);
and AND2 (N4802, N4792, N1109);
or OR2 (N4803, N4796, N2755);
nand NAND3 (N4804, N4803, N3454, N4774);
and AND3 (N4805, N4804, N1308, N2003);
or OR2 (N4806, N4785, N2988);
nand NAND3 (N4807, N4800, N3234, N4443);
or OR4 (N4808, N4802, N1292, N4523, N3896);
and AND4 (N4809, N4808, N3558, N1552, N613);
or OR4 (N4810, N4806, N629, N3756, N4528);
and AND3 (N4811, N4809, N238, N103);
nor NOR4 (N4812, N4798, N241, N2198, N1569);
or OR3 (N4813, N4810, N4001, N4130);
nand NAND3 (N4814, N4813, N2450, N4600);
buf BUF1 (N4815, N4807);
buf BUF1 (N4816, N4812);
buf BUF1 (N4817, N4791);
and AND2 (N4818, N4801, N159);
and AND2 (N4819, N4797, N1370);
nand NAND3 (N4820, N4814, N675, N4274);
buf BUF1 (N4821, N4769);
nand NAND4 (N4822, N4821, N88, N1014, N466);
xor XOR2 (N4823, N4817, N1167);
and AND3 (N4824, N4823, N4092, N1005);
not NOT1 (N4825, N4822);
buf BUF1 (N4826, N4811);
and AND2 (N4827, N4826, N2924);
nand NAND3 (N4828, N4815, N1043, N3374);
or OR3 (N4829, N4820, N397, N2381);
nor NOR3 (N4830, N4824, N2563, N1037);
or OR3 (N4831, N4818, N4007, N2858);
xor XOR2 (N4832, N4784, N1832);
not NOT1 (N4833, N4830);
and AND3 (N4834, N4825, N729, N3229);
nor NOR3 (N4835, N4805, N4421, N3358);
not NOT1 (N4836, N4829);
xor XOR2 (N4837, N4835, N947);
xor XOR2 (N4838, N4836, N4439);
xor XOR2 (N4839, N4816, N358);
xor XOR2 (N4840, N4831, N451);
not NOT1 (N4841, N4840);
nor NOR2 (N4842, N4832, N1180);
xor XOR2 (N4843, N4842, N3307);
not NOT1 (N4844, N4834);
xor XOR2 (N4845, N4827, N1632);
xor XOR2 (N4846, N4844, N565);
buf BUF1 (N4847, N4843);
and AND2 (N4848, N4833, N2710);
buf BUF1 (N4849, N4845);
not NOT1 (N4850, N4839);
nor NOR4 (N4851, N4847, N1652, N1450, N827);
nor NOR2 (N4852, N4851, N3830);
not NOT1 (N4853, N4848);
xor XOR2 (N4854, N4819, N2825);
nor NOR3 (N4855, N4850, N4222, N2612);
nor NOR3 (N4856, N4852, N787, N2226);
or OR3 (N4857, N4841, N1430, N1024);
and AND2 (N4858, N4857, N560);
xor XOR2 (N4859, N4846, N615);
nand NAND2 (N4860, N4837, N1499);
nor NOR3 (N4861, N4855, N4252, N3679);
and AND3 (N4862, N4860, N935, N978);
or OR3 (N4863, N4854, N2609, N432);
nor NOR4 (N4864, N4858, N884, N1061, N1590);
or OR2 (N4865, N4864, N4271);
buf BUF1 (N4866, N4856);
and AND4 (N4867, N4828, N3385, N4517, N3325);
buf BUF1 (N4868, N4866);
nand NAND3 (N4869, N4838, N534, N3355);
nor NOR4 (N4870, N4862, N3843, N4246, N1260);
not NOT1 (N4871, N4863);
xor XOR2 (N4872, N4868, N175);
and AND4 (N4873, N4859, N2890, N211, N4854);
nor NOR2 (N4874, N4871, N3810);
nor NOR3 (N4875, N4869, N17, N4270);
buf BUF1 (N4876, N4870);
nor NOR4 (N4877, N4861, N3400, N65, N4492);
buf BUF1 (N4878, N4876);
and AND4 (N4879, N4873, N1911, N2121, N2158);
or OR2 (N4880, N4853, N2706);
not NOT1 (N4881, N4849);
or OR3 (N4882, N4867, N534, N349);
and AND3 (N4883, N4872, N4458, N1313);
nor NOR4 (N4884, N4874, N714, N4836, N1323);
not NOT1 (N4885, N4865);
nand NAND4 (N4886, N4884, N4185, N3311, N4482);
not NOT1 (N4887, N4877);
buf BUF1 (N4888, N4875);
nor NOR2 (N4889, N4879, N2464);
nand NAND4 (N4890, N4886, N2105, N3467, N426);
not NOT1 (N4891, N4883);
buf BUF1 (N4892, N4889);
or OR4 (N4893, N4885, N1165, N76, N2052);
buf BUF1 (N4894, N4878);
not NOT1 (N4895, N4880);
not NOT1 (N4896, N4895);
nand NAND3 (N4897, N4887, N1278, N2244);
buf BUF1 (N4898, N4893);
nor NOR4 (N4899, N4890, N1028, N2718, N2846);
nand NAND3 (N4900, N4899, N1912, N466);
nand NAND2 (N4901, N4897, N2932);
not NOT1 (N4902, N4901);
buf BUF1 (N4903, N4888);
nor NOR4 (N4904, N4896, N163, N3670, N2561);
or OR2 (N4905, N4903, N1866);
nor NOR4 (N4906, N4902, N4266, N136, N4626);
xor XOR2 (N4907, N4891, N2484);
or OR3 (N4908, N4907, N4597, N3777);
and AND2 (N4909, N4881, N3376);
nor NOR2 (N4910, N4892, N531);
nand NAND4 (N4911, N4900, N3856, N2792, N2188);
nor NOR4 (N4912, N4911, N2497, N3222, N1165);
not NOT1 (N4913, N4910);
nor NOR4 (N4914, N4906, N3884, N4037, N536);
nand NAND4 (N4915, N4913, N4721, N3569, N1998);
buf BUF1 (N4916, N4904);
xor XOR2 (N4917, N4909, N2091);
not NOT1 (N4918, N4915);
nand NAND4 (N4919, N4917, N1083, N592, N320);
not NOT1 (N4920, N4918);
nand NAND4 (N4921, N4914, N3888, N2132, N3499);
and AND2 (N4922, N4898, N3345);
and AND3 (N4923, N4921, N3213, N2722);
buf BUF1 (N4924, N4905);
buf BUF1 (N4925, N4894);
nor NOR4 (N4926, N4919, N2342, N3295, N1254);
nand NAND3 (N4927, N4923, N274, N3374);
and AND2 (N4928, N4916, N4230);
buf BUF1 (N4929, N4926);
and AND3 (N4930, N4924, N2992, N1815);
nor NOR4 (N4931, N4882, N4523, N3531, N2177);
nand NAND3 (N4932, N4925, N1107, N133);
xor XOR2 (N4933, N4922, N394);
nand NAND2 (N4934, N4928, N4740);
and AND4 (N4935, N4934, N2885, N1617, N4356);
buf BUF1 (N4936, N4930);
not NOT1 (N4937, N4936);
nor NOR3 (N4938, N4935, N4658, N4935);
or OR4 (N4939, N4920, N1071, N3777, N1820);
or OR3 (N4940, N4938, N4020, N3307);
nor NOR2 (N4941, N4912, N2321);
xor XOR2 (N4942, N4932, N4137);
buf BUF1 (N4943, N4927);
nand NAND3 (N4944, N4942, N3388, N4916);
or OR2 (N4945, N4929, N2306);
buf BUF1 (N4946, N4908);
not NOT1 (N4947, N4943);
and AND3 (N4948, N4944, N1682, N649);
not NOT1 (N4949, N4939);
or OR2 (N4950, N4937, N3012);
buf BUF1 (N4951, N4946);
nand NAND4 (N4952, N4951, N2025, N2773, N3586);
xor XOR2 (N4953, N4952, N3046);
nand NAND4 (N4954, N4949, N1906, N109, N590);
or OR4 (N4955, N4945, N3661, N1429, N1161);
nand NAND4 (N4956, N4950, N4070, N3047, N2763);
or OR4 (N4957, N4940, N4539, N2916, N3848);
or OR3 (N4958, N4956, N2115, N2003);
and AND3 (N4959, N4931, N2978, N53);
and AND4 (N4960, N4933, N4876, N3175, N78);
nand NAND3 (N4961, N4959, N1956, N389);
xor XOR2 (N4962, N4953, N3424);
and AND2 (N4963, N4955, N3433);
and AND2 (N4964, N4941, N3421);
or OR3 (N4965, N4958, N775, N699);
xor XOR2 (N4966, N4954, N1771);
not NOT1 (N4967, N4966);
xor XOR2 (N4968, N4964, N2397);
nand NAND4 (N4969, N4947, N4829, N2148, N3805);
nand NAND3 (N4970, N4962, N4376, N3145);
buf BUF1 (N4971, N4970);
xor XOR2 (N4972, N4948, N4356);
nand NAND4 (N4973, N4969, N2575, N1669, N4678);
and AND2 (N4974, N4961, N355);
buf BUF1 (N4975, N4960);
buf BUF1 (N4976, N4973);
nand NAND2 (N4977, N4976, N4513);
or OR2 (N4978, N4963, N2955);
nand NAND3 (N4979, N4971, N2663, N2628);
nand NAND4 (N4980, N4974, N530, N14, N4140);
nand NAND4 (N4981, N4978, N3273, N3568, N3321);
and AND4 (N4982, N4979, N655, N914, N388);
or OR2 (N4983, N4980, N1333);
nand NAND4 (N4984, N4957, N919, N3198, N4244);
nor NOR4 (N4985, N4975, N1349, N898, N4206);
not NOT1 (N4986, N4965);
nor NOR3 (N4987, N4981, N3862, N4744);
or OR4 (N4988, N4982, N2654, N3058, N624);
and AND4 (N4989, N4968, N2817, N289, N4585);
and AND2 (N4990, N4986, N2602);
xor XOR2 (N4991, N4988, N3223);
and AND2 (N4992, N4967, N2162);
or OR2 (N4993, N4991, N180);
xor XOR2 (N4994, N4972, N3116);
and AND4 (N4995, N4993, N1923, N1616, N3059);
xor XOR2 (N4996, N4987, N3233);
and AND2 (N4997, N4994, N3883);
nand NAND4 (N4998, N4992, N983, N4865, N4871);
nor NOR2 (N4999, N4990, N4633);
nand NAND3 (N5000, N4999, N1391, N4816);
buf BUF1 (N5001, N4997);
nor NOR3 (N5002, N4989, N4286, N1661);
not NOT1 (N5003, N4977);
not NOT1 (N5004, N5000);
nor NOR3 (N5005, N5001, N3790, N1126);
nor NOR3 (N5006, N4985, N4235, N2443);
and AND2 (N5007, N4995, N1349);
nand NAND3 (N5008, N4998, N531, N1631);
and AND3 (N5009, N5007, N254, N1070);
nor NOR3 (N5010, N5004, N4203, N2891);
buf BUF1 (N5011, N5008);
buf BUF1 (N5012, N4983);
not NOT1 (N5013, N4996);
or OR4 (N5014, N5009, N2190, N3945, N2857);
nor NOR2 (N5015, N5014, N1885);
not NOT1 (N5016, N5002);
nand NAND4 (N5017, N5013, N3081, N4678, N831);
nand NAND2 (N5018, N5015, N618);
and AND4 (N5019, N5018, N4327, N1117, N2574);
buf BUF1 (N5020, N5010);
nor NOR2 (N5021, N5017, N3371);
buf BUF1 (N5022, N5016);
or OR3 (N5023, N5012, N3779, N3499);
xor XOR2 (N5024, N5011, N1368);
not NOT1 (N5025, N4984);
or OR3 (N5026, N5006, N3711, N4879);
xor XOR2 (N5027, N5005, N3666);
not NOT1 (N5028, N5019);
and AND2 (N5029, N5022, N493);
not NOT1 (N5030, N5025);
nand NAND4 (N5031, N5021, N4960, N4494, N2224);
or OR3 (N5032, N5031, N732, N311);
buf BUF1 (N5033, N5003);
buf BUF1 (N5034, N5033);
nand NAND3 (N5035, N5024, N3758, N4184);
nand NAND3 (N5036, N5028, N2083, N587);
and AND2 (N5037, N5032, N1192);
or OR3 (N5038, N5023, N1842, N2360);
and AND3 (N5039, N5036, N2395, N677);
xor XOR2 (N5040, N5026, N2277);
or OR3 (N5041, N5027, N2296, N2787);
nand NAND2 (N5042, N5039, N4715);
xor XOR2 (N5043, N5035, N2823);
nand NAND3 (N5044, N5043, N3763, N4054);
not NOT1 (N5045, N5034);
nand NAND2 (N5046, N5044, N1605);
buf BUF1 (N5047, N5020);
nor NOR4 (N5048, N5046, N3129, N3707, N3317);
nor NOR2 (N5049, N5045, N1664);
xor XOR2 (N5050, N5041, N1140);
and AND3 (N5051, N5029, N4891, N2152);
buf BUF1 (N5052, N5051);
and AND4 (N5053, N5049, N939, N1296, N678);
or OR3 (N5054, N5047, N552, N1303);
and AND2 (N5055, N5040, N2536);
xor XOR2 (N5056, N5048, N2513);
nand NAND3 (N5057, N5053, N1586, N3097);
buf BUF1 (N5058, N5042);
nand NAND3 (N5059, N5054, N2012, N689);
and AND4 (N5060, N5038, N3271, N2863, N2479);
nand NAND4 (N5061, N5052, N1765, N1443, N2741);
and AND2 (N5062, N5055, N3051);
buf BUF1 (N5063, N5060);
or OR2 (N5064, N5057, N2538);
or OR2 (N5065, N5063, N2362);
xor XOR2 (N5066, N5061, N3022);
buf BUF1 (N5067, N5056);
nor NOR4 (N5068, N5050, N4163, N480, N962);
or OR2 (N5069, N5068, N3494);
xor XOR2 (N5070, N5062, N3955);
and AND4 (N5071, N5059, N3440, N4619, N3663);
nor NOR3 (N5072, N5030, N2610, N3962);
or OR3 (N5073, N5070, N3988, N4294);
nand NAND2 (N5074, N5073, N3070);
or OR2 (N5075, N5072, N4231);
nor NOR2 (N5076, N5071, N598);
nand NAND2 (N5077, N5066, N105);
or OR3 (N5078, N5075, N3991, N2966);
not NOT1 (N5079, N5077);
xor XOR2 (N5080, N5079, N4505);
or OR4 (N5081, N5067, N520, N2322, N2189);
or OR3 (N5082, N5076, N1837, N2961);
nor NOR3 (N5083, N5064, N1921, N3468);
or OR2 (N5084, N5078, N2998);
not NOT1 (N5085, N5069);
nand NAND4 (N5086, N5081, N4813, N4398, N178);
nand NAND4 (N5087, N5080, N4839, N4052, N3940);
buf BUF1 (N5088, N5058);
nor NOR2 (N5089, N5082, N2545);
nor NOR3 (N5090, N5065, N2021, N4236);
buf BUF1 (N5091, N5090);
nand NAND3 (N5092, N5089, N3248, N4285);
not NOT1 (N5093, N5088);
buf BUF1 (N5094, N5083);
buf BUF1 (N5095, N5087);
or OR2 (N5096, N5094, N1226);
nor NOR4 (N5097, N5086, N2370, N4986, N1673);
buf BUF1 (N5098, N5096);
and AND3 (N5099, N5095, N2086, N5003);
nor NOR2 (N5100, N5037, N4118);
xor XOR2 (N5101, N5092, N949);
xor XOR2 (N5102, N5100, N2788);
buf BUF1 (N5103, N5101);
or OR3 (N5104, N5085, N3154, N791);
nand NAND3 (N5105, N5099, N1690, N2540);
not NOT1 (N5106, N5103);
not NOT1 (N5107, N5106);
not NOT1 (N5108, N5105);
xor XOR2 (N5109, N5074, N2742);
not NOT1 (N5110, N5098);
nand NAND2 (N5111, N5102, N1116);
not NOT1 (N5112, N5108);
nor NOR4 (N5113, N5111, N424, N2729, N394);
nor NOR2 (N5114, N5112, N944);
xor XOR2 (N5115, N5107, N1439);
nand NAND2 (N5116, N5113, N94);
buf BUF1 (N5117, N5110);
buf BUF1 (N5118, N5097);
nor NOR3 (N5119, N5109, N1529, N4582);
buf BUF1 (N5120, N5104);
not NOT1 (N5121, N5119);
and AND3 (N5122, N5117, N3874, N4001);
nand NAND3 (N5123, N5114, N809, N1324);
nor NOR3 (N5124, N5120, N4857, N3780);
xor XOR2 (N5125, N5121, N1015);
nor NOR3 (N5126, N5115, N1610, N245);
or OR4 (N5127, N5084, N2729, N3994, N3134);
and AND3 (N5128, N5091, N1578, N3260);
buf BUF1 (N5129, N5122);
and AND4 (N5130, N5126, N3128, N2459, N4164);
buf BUF1 (N5131, N5130);
xor XOR2 (N5132, N5128, N460);
buf BUF1 (N5133, N5125);
not NOT1 (N5134, N5093);
nor NOR2 (N5135, N5132, N2732);
xor XOR2 (N5136, N5129, N3072);
and AND3 (N5137, N5127, N3458, N2752);
xor XOR2 (N5138, N5135, N1698);
or OR4 (N5139, N5136, N1899, N4134, N1115);
xor XOR2 (N5140, N5124, N3242);
or OR3 (N5141, N5137, N4751, N2891);
nor NOR3 (N5142, N5139, N1925, N68);
buf BUF1 (N5143, N5134);
nor NOR4 (N5144, N5143, N307, N783, N415);
and AND3 (N5145, N5141, N336, N2497);
and AND3 (N5146, N5133, N1484, N89);
or OR4 (N5147, N5144, N529, N2896, N4113);
not NOT1 (N5148, N5118);
not NOT1 (N5149, N5116);
not NOT1 (N5150, N5146);
nand NAND3 (N5151, N5142, N1889, N4862);
or OR3 (N5152, N5151, N4199, N861);
xor XOR2 (N5153, N5149, N4898);
and AND3 (N5154, N5148, N1877, N458);
xor XOR2 (N5155, N5150, N2953);
not NOT1 (N5156, N5145);
and AND4 (N5157, N5131, N1703, N3691, N1430);
nand NAND2 (N5158, N5147, N3561);
and AND3 (N5159, N5157, N1856, N479);
and AND2 (N5160, N5158, N2483);
xor XOR2 (N5161, N5156, N1855);
nand NAND2 (N5162, N5155, N3319);
or OR2 (N5163, N5159, N452);
and AND4 (N5164, N5162, N280, N3816, N2775);
nor NOR4 (N5165, N5138, N497, N4253, N4223);
or OR4 (N5166, N5140, N4545, N3234, N967);
nor NOR2 (N5167, N5153, N1766);
and AND3 (N5168, N5160, N2984, N1535);
nand NAND4 (N5169, N5154, N2288, N1275, N1109);
and AND4 (N5170, N5166, N1998, N1047, N4833);
nor NOR4 (N5171, N5123, N351, N2687, N4831);
nand NAND4 (N5172, N5164, N197, N4714, N1668);
and AND4 (N5173, N5169, N2290, N237, N1790);
and AND2 (N5174, N5161, N3711);
nor NOR3 (N5175, N5170, N1339, N2132);
nand NAND4 (N5176, N5173, N3073, N1156, N1268);
and AND2 (N5177, N5175, N3265);
and AND3 (N5178, N5167, N1453, N76);
or OR3 (N5179, N5178, N530, N5037);
or OR2 (N5180, N5152, N2230);
or OR3 (N5181, N5171, N677, N2817);
xor XOR2 (N5182, N5180, N1087);
nor NOR2 (N5183, N5179, N4710);
buf BUF1 (N5184, N5174);
xor XOR2 (N5185, N5181, N3915);
or OR4 (N5186, N5172, N3857, N1342, N3292);
or OR3 (N5187, N5182, N2414, N214);
and AND3 (N5188, N5187, N3371, N1022);
nand NAND3 (N5189, N5188, N1489, N2591);
not NOT1 (N5190, N5165);
and AND4 (N5191, N5189, N28, N3025, N5175);
not NOT1 (N5192, N5168);
nand NAND2 (N5193, N5192, N622);
and AND2 (N5194, N5184, N1917);
nand NAND2 (N5195, N5191, N2529);
buf BUF1 (N5196, N5163);
nor NOR4 (N5197, N5195, N3983, N375, N3277);
buf BUF1 (N5198, N5194);
nor NOR2 (N5199, N5176, N2119);
nand NAND2 (N5200, N5185, N2818);
xor XOR2 (N5201, N5193, N728);
nor NOR2 (N5202, N5186, N4131);
nor NOR3 (N5203, N5202, N4133, N627);
nor NOR4 (N5204, N5183, N1235, N4614, N524);
xor XOR2 (N5205, N5204, N1720);
xor XOR2 (N5206, N5177, N248);
not NOT1 (N5207, N5196);
buf BUF1 (N5208, N5199);
xor XOR2 (N5209, N5201, N3544);
buf BUF1 (N5210, N5190);
xor XOR2 (N5211, N5207, N3126);
and AND4 (N5212, N5211, N1091, N1848, N3435);
buf BUF1 (N5213, N5197);
nor NOR2 (N5214, N5212, N1314);
buf BUF1 (N5215, N5214);
xor XOR2 (N5216, N5209, N630);
nor NOR4 (N5217, N5200, N1653, N890, N3654);
buf BUF1 (N5218, N5203);
not NOT1 (N5219, N5208);
and AND4 (N5220, N5215, N2199, N4128, N3076);
xor XOR2 (N5221, N5198, N4256);
xor XOR2 (N5222, N5219, N217);
and AND3 (N5223, N5216, N4702, N3933);
nor NOR2 (N5224, N5223, N1048);
nor NOR3 (N5225, N5220, N2840, N4213);
nor NOR4 (N5226, N5213, N496, N3328, N1405);
nor NOR4 (N5227, N5206, N663, N2750, N4070);
nor NOR3 (N5228, N5217, N1439, N2226);
nand NAND3 (N5229, N5218, N4823, N4189);
and AND4 (N5230, N5222, N4706, N2703, N3580);
nor NOR2 (N5231, N5225, N2385);
nand NAND4 (N5232, N5226, N2104, N709, N3368);
and AND3 (N5233, N5224, N4328, N3113);
buf BUF1 (N5234, N5228);
and AND2 (N5235, N5210, N3278);
xor XOR2 (N5236, N5232, N1785);
or OR2 (N5237, N5236, N2493);
and AND2 (N5238, N5230, N3883);
nand NAND4 (N5239, N5229, N701, N2175, N3526);
or OR3 (N5240, N5234, N1280, N3137);
nor NOR3 (N5241, N5238, N2345, N3132);
xor XOR2 (N5242, N5231, N3491);
nor NOR3 (N5243, N5237, N4173, N3794);
and AND3 (N5244, N5241, N383, N539);
not NOT1 (N5245, N5242);
nand NAND3 (N5246, N5227, N1987, N2220);
not NOT1 (N5247, N5233);
nand NAND3 (N5248, N5240, N1147, N4300);
and AND3 (N5249, N5235, N640, N2282);
not NOT1 (N5250, N5248);
not NOT1 (N5251, N5246);
or OR2 (N5252, N5221, N4422);
xor XOR2 (N5253, N5205, N386);
nand NAND2 (N5254, N5251, N2990);
nand NAND4 (N5255, N5244, N5099, N1924, N5013);
and AND3 (N5256, N5243, N1780, N5245);
not NOT1 (N5257, N2735);
or OR3 (N5258, N5257, N4847, N2865);
nand NAND4 (N5259, N5258, N1501, N2087, N3583);
buf BUF1 (N5260, N5239);
xor XOR2 (N5261, N5250, N1910);
not NOT1 (N5262, N5247);
nor NOR4 (N5263, N5252, N212, N1310, N4728);
not NOT1 (N5264, N5255);
not NOT1 (N5265, N5260);
buf BUF1 (N5266, N5259);
and AND3 (N5267, N5261, N3919, N2123);
not NOT1 (N5268, N5263);
not NOT1 (N5269, N5249);
xor XOR2 (N5270, N5265, N3064);
xor XOR2 (N5271, N5267, N4202);
and AND4 (N5272, N5253, N618, N4293, N1780);
not NOT1 (N5273, N5256);
not NOT1 (N5274, N5266);
nand NAND4 (N5275, N5262, N4502, N2155, N932);
nand NAND3 (N5276, N5273, N2875, N931);
and AND2 (N5277, N5274, N1933);
xor XOR2 (N5278, N5275, N1435);
nor NOR4 (N5279, N5270, N3604, N2722, N333);
or OR2 (N5280, N5264, N1610);
xor XOR2 (N5281, N5278, N4061);
nand NAND3 (N5282, N5254, N260, N3376);
and AND4 (N5283, N5268, N2015, N2322, N727);
or OR3 (N5284, N5283, N4805, N4525);
nand NAND3 (N5285, N5284, N1747, N3837);
not NOT1 (N5286, N5281);
or OR4 (N5287, N5286, N1179, N1344, N3581);
nand NAND4 (N5288, N5287, N3954, N1668, N638);
nor NOR4 (N5289, N5269, N4957, N3493, N1329);
xor XOR2 (N5290, N5285, N4878);
xor XOR2 (N5291, N5289, N3531);
buf BUF1 (N5292, N5279);
and AND4 (N5293, N5288, N1505, N1838, N4716);
not NOT1 (N5294, N5290);
xor XOR2 (N5295, N5280, N4760);
nor NOR2 (N5296, N5276, N2193);
not NOT1 (N5297, N5282);
not NOT1 (N5298, N5295);
and AND2 (N5299, N5271, N3962);
nand NAND2 (N5300, N5292, N1192);
nor NOR3 (N5301, N5272, N3316, N4219);
buf BUF1 (N5302, N5293);
nor NOR2 (N5303, N5291, N3078);
nor NOR2 (N5304, N5301, N1704);
xor XOR2 (N5305, N5277, N817);
buf BUF1 (N5306, N5300);
not NOT1 (N5307, N5304);
nor NOR4 (N5308, N5305, N1083, N4897, N2612);
and AND3 (N5309, N5298, N3684, N4872);
or OR2 (N5310, N5294, N2395);
not NOT1 (N5311, N5297);
and AND4 (N5312, N5311, N2247, N2251, N2399);
or OR2 (N5313, N5299, N2418);
nor NOR2 (N5314, N5303, N1187);
not NOT1 (N5315, N5302);
nand NAND4 (N5316, N5310, N2092, N5042, N302);
and AND2 (N5317, N5296, N2055);
and AND4 (N5318, N5314, N419, N3829, N976);
or OR3 (N5319, N5312, N4297, N2264);
nand NAND2 (N5320, N5307, N2991);
or OR4 (N5321, N5308, N4521, N2121, N5018);
not NOT1 (N5322, N5306);
xor XOR2 (N5323, N5313, N3633);
and AND2 (N5324, N5316, N1786);
xor XOR2 (N5325, N5317, N2330);
xor XOR2 (N5326, N5321, N3090);
not NOT1 (N5327, N5319);
or OR2 (N5328, N5318, N4059);
not NOT1 (N5329, N5328);
nor NOR2 (N5330, N5329, N3013);
xor XOR2 (N5331, N5324, N3455);
nand NAND2 (N5332, N5320, N912);
and AND2 (N5333, N5326, N3837);
nor NOR3 (N5334, N5322, N637, N2625);
and AND2 (N5335, N5331, N1083);
nand NAND2 (N5336, N5330, N1200);
nand NAND4 (N5337, N5336, N4482, N2800, N5067);
nor NOR4 (N5338, N5334, N2413, N3821, N5046);
or OR3 (N5339, N5335, N2110, N2971);
or OR4 (N5340, N5325, N1257, N2334, N794);
nand NAND3 (N5341, N5315, N980, N2025);
and AND3 (N5342, N5340, N1725, N1123);
buf BUF1 (N5343, N5339);
xor XOR2 (N5344, N5309, N599);
xor XOR2 (N5345, N5333, N4543);
not NOT1 (N5346, N5327);
or OR3 (N5347, N5341, N3613, N1322);
xor XOR2 (N5348, N5323, N4224);
or OR4 (N5349, N5332, N2750, N483, N3920);
xor XOR2 (N5350, N5349, N1076);
xor XOR2 (N5351, N5338, N3746);
nor NOR3 (N5352, N5344, N2007, N1775);
or OR3 (N5353, N5342, N3864, N4567);
not NOT1 (N5354, N5353);
nand NAND3 (N5355, N5348, N1638, N2597);
or OR4 (N5356, N5351, N4131, N4972, N1723);
buf BUF1 (N5357, N5352);
and AND2 (N5358, N5347, N4854);
xor XOR2 (N5359, N5343, N2910);
or OR4 (N5360, N5359, N3027, N596, N2687);
and AND2 (N5361, N5355, N2343);
xor XOR2 (N5362, N5357, N3759);
xor XOR2 (N5363, N5362, N2844);
xor XOR2 (N5364, N5354, N650);
buf BUF1 (N5365, N5346);
and AND3 (N5366, N5350, N5148, N5012);
nand NAND3 (N5367, N5363, N5000, N2685);
nand NAND4 (N5368, N5367, N3384, N1401, N4210);
not NOT1 (N5369, N5356);
nor NOR4 (N5370, N5365, N4995, N3298, N1583);
not NOT1 (N5371, N5337);
and AND2 (N5372, N5364, N979);
not NOT1 (N5373, N5368);
nor NOR4 (N5374, N5372, N3576, N4660, N3334);
and AND3 (N5375, N5373, N106, N207);
or OR3 (N5376, N5360, N2606, N1400);
buf BUF1 (N5377, N5371);
buf BUF1 (N5378, N5377);
xor XOR2 (N5379, N5376, N3857);
nand NAND3 (N5380, N5370, N3071, N1134);
or OR2 (N5381, N5380, N2332);
and AND3 (N5382, N5374, N2601, N954);
xor XOR2 (N5383, N5358, N129);
buf BUF1 (N5384, N5382);
not NOT1 (N5385, N5384);
and AND3 (N5386, N5375, N5182, N3430);
or OR2 (N5387, N5345, N2185);
buf BUF1 (N5388, N5383);
or OR3 (N5389, N5366, N5362, N738);
not NOT1 (N5390, N5386);
nor NOR3 (N5391, N5389, N3149, N4474);
or OR2 (N5392, N5391, N2011);
nand NAND3 (N5393, N5387, N1057, N693);
or OR3 (N5394, N5388, N1581, N3224);
nand NAND4 (N5395, N5394, N4935, N3407, N3273);
nand NAND4 (N5396, N5392, N968, N2454, N4233);
not NOT1 (N5397, N5379);
xor XOR2 (N5398, N5397, N3964);
xor XOR2 (N5399, N5398, N2467);
nor NOR4 (N5400, N5399, N1534, N1678, N1217);
and AND3 (N5401, N5395, N2162, N2710);
xor XOR2 (N5402, N5378, N4497);
and AND4 (N5403, N5369, N4433, N1521, N2018);
buf BUF1 (N5404, N5396);
nor NOR3 (N5405, N5401, N3726, N4159);
buf BUF1 (N5406, N5405);
and AND3 (N5407, N5403, N2001, N908);
nand NAND3 (N5408, N5402, N649, N1192);
or OR3 (N5409, N5393, N520, N1802);
buf BUF1 (N5410, N5385);
not NOT1 (N5411, N5361);
buf BUF1 (N5412, N5381);
and AND3 (N5413, N5409, N3583, N4108);
and AND4 (N5414, N5406, N2065, N4918, N5385);
and AND4 (N5415, N5407, N2485, N430, N4249);
xor XOR2 (N5416, N5414, N3483);
xor XOR2 (N5417, N5404, N4224);
xor XOR2 (N5418, N5412, N2572);
not NOT1 (N5419, N5408);
nor NOR3 (N5420, N5415, N2823, N1419);
nor NOR3 (N5421, N5390, N111, N3797);
or OR4 (N5422, N5400, N3884, N3273, N927);
and AND3 (N5423, N5416, N1161, N2920);
nor NOR3 (N5424, N5413, N1568, N484);
nor NOR3 (N5425, N5422, N1633, N3241);
buf BUF1 (N5426, N5424);
buf BUF1 (N5427, N5410);
buf BUF1 (N5428, N5418);
nand NAND4 (N5429, N5428, N1980, N3911, N1869);
nor NOR2 (N5430, N5417, N2373);
and AND2 (N5431, N5425, N3983);
and AND3 (N5432, N5411, N3545, N4131);
xor XOR2 (N5433, N5421, N3918);
nor NOR2 (N5434, N5427, N43);
and AND2 (N5435, N5432, N1683);
nand NAND4 (N5436, N5426, N1207, N484, N3973);
buf BUF1 (N5437, N5433);
buf BUF1 (N5438, N5429);
nor NOR3 (N5439, N5430, N5323, N1932);
buf BUF1 (N5440, N5431);
xor XOR2 (N5441, N5419, N4780);
xor XOR2 (N5442, N5438, N3116);
or OR2 (N5443, N5442, N1408);
nand NAND3 (N5444, N5436, N5238, N3294);
and AND4 (N5445, N5434, N2696, N3082, N1221);
xor XOR2 (N5446, N5435, N5183);
or OR2 (N5447, N5423, N197);
buf BUF1 (N5448, N5443);
nand NAND2 (N5449, N5446, N4390);
not NOT1 (N5450, N5437);
and AND4 (N5451, N5439, N1069, N1460, N5309);
and AND2 (N5452, N5449, N4582);
and AND4 (N5453, N5444, N1835, N3521, N197);
or OR4 (N5454, N5453, N3044, N1016, N3933);
and AND3 (N5455, N5448, N949, N342);
and AND4 (N5456, N5454, N2817, N3760, N1854);
buf BUF1 (N5457, N5440);
and AND3 (N5458, N5441, N603, N4404);
nor NOR4 (N5459, N5452, N3898, N3571, N5019);
xor XOR2 (N5460, N5445, N2635);
nand NAND3 (N5461, N5460, N2576, N2271);
nor NOR3 (N5462, N5447, N4524, N3914);
or OR2 (N5463, N5420, N4879);
xor XOR2 (N5464, N5462, N370);
nor NOR3 (N5465, N5461, N4527, N42);
nand NAND4 (N5466, N5455, N1249, N4149, N2223);
not NOT1 (N5467, N5464);
nor NOR4 (N5468, N5458, N3655, N3694, N4612);
or OR3 (N5469, N5459, N11, N5058);
and AND2 (N5470, N5456, N4156);
buf BUF1 (N5471, N5451);
nand NAND2 (N5472, N5467, N2513);
and AND4 (N5473, N5469, N2436, N1366, N4678);
and AND2 (N5474, N5473, N5360);
buf BUF1 (N5475, N5465);
nand NAND4 (N5476, N5468, N2192, N2615, N170);
and AND2 (N5477, N5457, N765);
and AND3 (N5478, N5470, N174, N885);
and AND3 (N5479, N5477, N1166, N4549);
nor NOR4 (N5480, N5479, N3951, N2179, N5219);
nand NAND2 (N5481, N5450, N4085);
or OR2 (N5482, N5472, N3768);
or OR2 (N5483, N5463, N5064);
xor XOR2 (N5484, N5481, N1584);
buf BUF1 (N5485, N5474);
xor XOR2 (N5486, N5480, N3576);
xor XOR2 (N5487, N5483, N1239);
or OR4 (N5488, N5484, N27, N2581, N4303);
nor NOR3 (N5489, N5478, N920, N2622);
and AND2 (N5490, N5489, N5268);
nor NOR4 (N5491, N5476, N5081, N2040, N5262);
buf BUF1 (N5492, N5475);
nor NOR2 (N5493, N5490, N2925);
or OR4 (N5494, N5493, N3521, N3748, N983);
xor XOR2 (N5495, N5491, N5295);
nor NOR4 (N5496, N5487, N4755, N4396, N4135);
or OR4 (N5497, N5482, N3116, N5039, N4816);
nor NOR2 (N5498, N5495, N1834);
nand NAND3 (N5499, N5485, N1076, N2027);
nand NAND3 (N5500, N5496, N1514, N4293);
or OR3 (N5501, N5486, N4219, N2044);
nor NOR2 (N5502, N5492, N208);
nor NOR3 (N5503, N5499, N3295, N4637);
nor NOR3 (N5504, N5500, N3546, N1081);
or OR4 (N5505, N5498, N5100, N3634, N2444);
nand NAND4 (N5506, N5504, N1656, N602, N156);
nor NOR3 (N5507, N5502, N4166, N4042);
nor NOR4 (N5508, N5503, N662, N1671, N1046);
nor NOR4 (N5509, N5508, N4027, N3517, N314);
nand NAND4 (N5510, N5466, N1766, N5142, N4116);
xor XOR2 (N5511, N5506, N4289);
or OR4 (N5512, N5494, N5015, N3467, N3514);
nor NOR2 (N5513, N5505, N4907);
nand NAND4 (N5514, N5507, N1211, N300, N2515);
and AND2 (N5515, N5512, N660);
and AND4 (N5516, N5488, N5195, N4960, N3932);
and AND4 (N5517, N5513, N895, N3382, N1350);
xor XOR2 (N5518, N5514, N5110);
nand NAND3 (N5519, N5517, N2073, N1523);
not NOT1 (N5520, N5519);
not NOT1 (N5521, N5501);
buf BUF1 (N5522, N5497);
xor XOR2 (N5523, N5521, N4207);
buf BUF1 (N5524, N5522);
buf BUF1 (N5525, N5511);
nand NAND4 (N5526, N5525, N4428, N1327, N1809);
nor NOR4 (N5527, N5520, N2402, N3375, N1780);
not NOT1 (N5528, N5516);
not NOT1 (N5529, N5509);
nor NOR3 (N5530, N5527, N3900, N640);
xor XOR2 (N5531, N5530, N994);
and AND2 (N5532, N5518, N3788);
nor NOR3 (N5533, N5524, N909, N4683);
xor XOR2 (N5534, N5533, N2179);
buf BUF1 (N5535, N5526);
and AND3 (N5536, N5523, N3617, N1724);
or OR2 (N5537, N5532, N4193);
nand NAND4 (N5538, N5510, N4146, N89, N2473);
or OR4 (N5539, N5536, N4125, N3124, N4101);
buf BUF1 (N5540, N5515);
nor NOR3 (N5541, N5539, N325, N3731);
not NOT1 (N5542, N5541);
or OR4 (N5543, N5471, N991, N1593, N325);
not NOT1 (N5544, N5543);
and AND4 (N5545, N5531, N1708, N2649, N2937);
nor NOR3 (N5546, N5542, N1800, N3195);
or OR4 (N5547, N5535, N4836, N2583, N3664);
nor NOR4 (N5548, N5528, N4457, N1666, N4402);
or OR2 (N5549, N5540, N4861);
xor XOR2 (N5550, N5545, N2043);
buf BUF1 (N5551, N5546);
nor NOR3 (N5552, N5529, N2032, N1482);
buf BUF1 (N5553, N5551);
nor NOR2 (N5554, N5537, N4460);
not NOT1 (N5555, N5550);
not NOT1 (N5556, N5538);
nor NOR2 (N5557, N5534, N4818);
buf BUF1 (N5558, N5549);
nand NAND4 (N5559, N5553, N2737, N3533, N158);
nor NOR4 (N5560, N5544, N2965, N5221, N4918);
xor XOR2 (N5561, N5556, N3764);
or OR4 (N5562, N5557, N4420, N4212, N673);
and AND2 (N5563, N5558, N1092);
nand NAND2 (N5564, N5554, N5008);
or OR2 (N5565, N5555, N2405);
nand NAND4 (N5566, N5564, N1321, N5333, N1034);
not NOT1 (N5567, N5562);
not NOT1 (N5568, N5548);
nand NAND2 (N5569, N5547, N3193);
or OR3 (N5570, N5559, N41, N4151);
xor XOR2 (N5571, N5560, N147);
not NOT1 (N5572, N5569);
buf BUF1 (N5573, N5561);
nor NOR3 (N5574, N5565, N2192, N175);
not NOT1 (N5575, N5563);
nor NOR3 (N5576, N5572, N5496, N872);
or OR2 (N5577, N5552, N5570);
and AND4 (N5578, N4785, N2405, N4569, N3771);
not NOT1 (N5579, N5577);
and AND4 (N5580, N5574, N1354, N2604, N4295);
xor XOR2 (N5581, N5573, N4654);
nand NAND4 (N5582, N5579, N2189, N2434, N5517);
nor NOR2 (N5583, N5576, N1073);
and AND4 (N5584, N5575, N1970, N1856, N1417);
buf BUF1 (N5585, N5582);
not NOT1 (N5586, N5584);
nand NAND3 (N5587, N5567, N692, N2799);
nor NOR3 (N5588, N5578, N2516, N2268);
xor XOR2 (N5589, N5568, N5495);
nor NOR3 (N5590, N5586, N1577, N2601);
xor XOR2 (N5591, N5588, N1173);
or OR4 (N5592, N5571, N4072, N2225, N5096);
buf BUF1 (N5593, N5589);
or OR3 (N5594, N5583, N3048, N3445);
and AND3 (N5595, N5592, N2064, N2190);
nor NOR4 (N5596, N5587, N1047, N1598, N424);
xor XOR2 (N5597, N5581, N208);
xor XOR2 (N5598, N5595, N92);
xor XOR2 (N5599, N5591, N3317);
nand NAND4 (N5600, N5596, N289, N5102, N2999);
nand NAND2 (N5601, N5598, N2182);
and AND2 (N5602, N5594, N2570);
or OR2 (N5603, N5590, N3521);
nor NOR3 (N5604, N5601, N1300, N1059);
nor NOR2 (N5605, N5593, N3224);
nor NOR3 (N5606, N5605, N3608, N765);
buf BUF1 (N5607, N5600);
and AND2 (N5608, N5597, N4427);
nand NAND4 (N5609, N5599, N5406, N3939, N2960);
not NOT1 (N5610, N5602);
nor NOR3 (N5611, N5610, N1820, N4435);
and AND2 (N5612, N5607, N4233);
xor XOR2 (N5613, N5566, N3251);
or OR2 (N5614, N5580, N1714);
buf BUF1 (N5615, N5613);
or OR4 (N5616, N5585, N4267, N3442, N257);
and AND3 (N5617, N5608, N746, N2896);
buf BUF1 (N5618, N5615);
nor NOR3 (N5619, N5609, N3216, N1301);
nand NAND3 (N5620, N5619, N1430, N498);
nor NOR3 (N5621, N5620, N1552, N1201);
nand NAND2 (N5622, N5616, N1293);
xor XOR2 (N5623, N5603, N1485);
buf BUF1 (N5624, N5621);
and AND2 (N5625, N5604, N1492);
not NOT1 (N5626, N5625);
nand NAND3 (N5627, N5612, N1327, N2015);
not NOT1 (N5628, N5614);
or OR4 (N5629, N5628, N3485, N1566, N3241);
not NOT1 (N5630, N5623);
and AND2 (N5631, N5611, N1143);
nand NAND4 (N5632, N5618, N2843, N3305, N748);
or OR3 (N5633, N5626, N4020, N3483);
or OR4 (N5634, N5606, N3541, N501, N3301);
nor NOR2 (N5635, N5632, N4837);
nand NAND3 (N5636, N5633, N2350, N3227);
or OR2 (N5637, N5622, N3894);
nor NOR4 (N5638, N5630, N334, N2960, N1616);
not NOT1 (N5639, N5627);
not NOT1 (N5640, N5617);
not NOT1 (N5641, N5637);
not NOT1 (N5642, N5640);
or OR4 (N5643, N5638, N2405, N279, N3247);
or OR2 (N5644, N5641, N1068);
and AND4 (N5645, N5631, N1808, N352, N4934);
not NOT1 (N5646, N5644);
xor XOR2 (N5647, N5642, N4198);
xor XOR2 (N5648, N5643, N4107);
buf BUF1 (N5649, N5629);
buf BUF1 (N5650, N5624);
nor NOR3 (N5651, N5650, N248, N894);
not NOT1 (N5652, N5639);
xor XOR2 (N5653, N5636, N5406);
nor NOR3 (N5654, N5653, N1465, N4490);
xor XOR2 (N5655, N5654, N448);
xor XOR2 (N5656, N5647, N3077);
not NOT1 (N5657, N5646);
or OR3 (N5658, N5651, N4178, N5608);
and AND3 (N5659, N5658, N3940, N443);
and AND4 (N5660, N5634, N2683, N1485, N1043);
nand NAND3 (N5661, N5645, N2592, N4391);
not NOT1 (N5662, N5655);
and AND3 (N5663, N5661, N5548, N4346);
not NOT1 (N5664, N5659);
nor NOR2 (N5665, N5663, N5488);
nand NAND3 (N5666, N5649, N1585, N602);
nand NAND3 (N5667, N5666, N1814, N208);
nor NOR2 (N5668, N5665, N2356);
not NOT1 (N5669, N5667);
not NOT1 (N5670, N5657);
or OR2 (N5671, N5652, N1707);
nand NAND3 (N5672, N5670, N1529, N2580);
xor XOR2 (N5673, N5664, N2902);
buf BUF1 (N5674, N5668);
xor XOR2 (N5675, N5669, N2099);
xor XOR2 (N5676, N5648, N1424);
nand NAND4 (N5677, N5673, N2042, N4030, N5487);
buf BUF1 (N5678, N5660);
nor NOR4 (N5679, N5635, N4392, N877, N5321);
nor NOR2 (N5680, N5679, N903);
buf BUF1 (N5681, N5662);
or OR4 (N5682, N5680, N5348, N2689, N41);
and AND4 (N5683, N5656, N5639, N3535, N5183);
or OR2 (N5684, N5671, N967);
nand NAND3 (N5685, N5684, N5414, N2072);
not NOT1 (N5686, N5675);
nor NOR3 (N5687, N5674, N1066, N641);
xor XOR2 (N5688, N5681, N2477);
and AND2 (N5689, N5688, N3257);
buf BUF1 (N5690, N5687);
xor XOR2 (N5691, N5685, N4611);
nand NAND4 (N5692, N5678, N5145, N900, N1299);
nor NOR3 (N5693, N5672, N553, N3010);
nor NOR4 (N5694, N5689, N4471, N702, N3658);
nor NOR2 (N5695, N5686, N800);
and AND4 (N5696, N5692, N1237, N4201, N1591);
and AND2 (N5697, N5695, N4003);
nor NOR3 (N5698, N5682, N3239, N5191);
or OR3 (N5699, N5696, N3477, N54);
nand NAND4 (N5700, N5691, N5096, N3435, N4646);
xor XOR2 (N5701, N5690, N4508);
and AND2 (N5702, N5676, N3521);
xor XOR2 (N5703, N5698, N3897);
nor NOR2 (N5704, N5701, N2907);
nor NOR4 (N5705, N5704, N3895, N406, N4446);
buf BUF1 (N5706, N5694);
not NOT1 (N5707, N5683);
nor NOR2 (N5708, N5705, N4441);
buf BUF1 (N5709, N5677);
nor NOR2 (N5710, N5707, N3250);
and AND3 (N5711, N5693, N3227, N3937);
nand NAND4 (N5712, N5700, N1416, N3828, N664);
buf BUF1 (N5713, N5708);
or OR4 (N5714, N5712, N3600, N2672, N5568);
not NOT1 (N5715, N5710);
and AND3 (N5716, N5702, N2145, N669);
nor NOR3 (N5717, N5716, N2347, N1841);
buf BUF1 (N5718, N5717);
buf BUF1 (N5719, N5697);
and AND4 (N5720, N5715, N3744, N4960, N1756);
or OR2 (N5721, N5713, N4912);
buf BUF1 (N5722, N5721);
and AND4 (N5723, N5714, N1440, N5392, N2644);
or OR3 (N5724, N5719, N1310, N1181);
nor NOR2 (N5725, N5723, N3206);
xor XOR2 (N5726, N5722, N4701);
buf BUF1 (N5727, N5703);
nand NAND2 (N5728, N5726, N102);
nor NOR4 (N5729, N5711, N4224, N1768, N1814);
nor NOR2 (N5730, N5706, N2596);
buf BUF1 (N5731, N5727);
xor XOR2 (N5732, N5729, N1182);
and AND4 (N5733, N5699, N3360, N1156, N4647);
and AND2 (N5734, N5709, N3188);
buf BUF1 (N5735, N5725);
buf BUF1 (N5736, N5720);
not NOT1 (N5737, N5728);
xor XOR2 (N5738, N5730, N14);
nand NAND3 (N5739, N5731, N5525, N3945);
not NOT1 (N5740, N5718);
not NOT1 (N5741, N5736);
or OR4 (N5742, N5739, N4103, N3715, N2076);
not NOT1 (N5743, N5738);
buf BUF1 (N5744, N5734);
and AND4 (N5745, N5743, N5650, N1918, N259);
nand NAND3 (N5746, N5737, N1362, N692);
and AND3 (N5747, N5746, N3390, N2617);
or OR4 (N5748, N5745, N3326, N457, N2257);
or OR4 (N5749, N5748, N5053, N5092, N4423);
and AND3 (N5750, N5733, N2769, N5115);
not NOT1 (N5751, N5749);
or OR3 (N5752, N5732, N3132, N4192);
and AND3 (N5753, N5744, N5658, N2205);
and AND2 (N5754, N5741, N4472);
or OR2 (N5755, N5747, N179);
not NOT1 (N5756, N5751);
buf BUF1 (N5757, N5755);
xor XOR2 (N5758, N5753, N5012);
and AND3 (N5759, N5742, N2410, N1131);
xor XOR2 (N5760, N5758, N3103);
nor NOR3 (N5761, N5756, N3102, N1836);
not NOT1 (N5762, N5754);
xor XOR2 (N5763, N5762, N2513);
nand NAND2 (N5764, N5752, N2522);
nor NOR4 (N5765, N5763, N2106, N939, N4621);
buf BUF1 (N5766, N5735);
xor XOR2 (N5767, N5761, N229);
or OR3 (N5768, N5724, N3347, N1667);
buf BUF1 (N5769, N5767);
and AND2 (N5770, N5764, N4639);
or OR3 (N5771, N5750, N5408, N5649);
buf BUF1 (N5772, N5770);
nor NOR2 (N5773, N5766, N2470);
or OR3 (N5774, N5760, N5592, N2492);
nor NOR3 (N5775, N5740, N3653, N3644);
not NOT1 (N5776, N5765);
not NOT1 (N5777, N5757);
nor NOR2 (N5778, N5771, N4374);
nand NAND4 (N5779, N5769, N3297, N3905, N4120);
or OR4 (N5780, N5777, N5209, N1857, N5185);
not NOT1 (N5781, N5773);
or OR3 (N5782, N5781, N5301, N1675);
nor NOR2 (N5783, N5774, N5184);
and AND2 (N5784, N5772, N2821);
xor XOR2 (N5785, N5768, N4106);
nor NOR4 (N5786, N5782, N1022, N738, N4419);
nor NOR2 (N5787, N5779, N5437);
nand NAND2 (N5788, N5759, N2293);
nand NAND2 (N5789, N5788, N457);
buf BUF1 (N5790, N5783);
or OR3 (N5791, N5785, N870, N3281);
and AND3 (N5792, N5776, N4920, N3345);
nor NOR2 (N5793, N5789, N935);
nand NAND3 (N5794, N5787, N4613, N3465);
xor XOR2 (N5795, N5791, N2493);
or OR2 (N5796, N5794, N4860);
xor XOR2 (N5797, N5775, N2952);
nand NAND4 (N5798, N5778, N5777, N5257, N2639);
nand NAND2 (N5799, N5798, N4622);
and AND4 (N5800, N5790, N1109, N621, N5127);
or OR3 (N5801, N5796, N2439, N3554);
and AND2 (N5802, N5786, N2430);
nand NAND2 (N5803, N5780, N2300);
and AND4 (N5804, N5793, N5685, N1108, N4144);
and AND3 (N5805, N5801, N3826, N4675);
nor NOR4 (N5806, N5784, N1997, N648, N5518);
xor XOR2 (N5807, N5806, N3640);
xor XOR2 (N5808, N5802, N4719);
or OR3 (N5809, N5803, N1927, N291);
nor NOR4 (N5810, N5797, N4789, N2369, N2943);
or OR3 (N5811, N5792, N5297, N2744);
or OR4 (N5812, N5807, N2412, N1756, N3838);
and AND3 (N5813, N5811, N3776, N3398);
and AND2 (N5814, N5804, N3607);
not NOT1 (N5815, N5812);
nand NAND3 (N5816, N5813, N3012, N7);
xor XOR2 (N5817, N5795, N4250);
xor XOR2 (N5818, N5816, N1724);
nand NAND4 (N5819, N5800, N3976, N408, N5304);
nor NOR3 (N5820, N5814, N4536, N723);
nor NOR3 (N5821, N5799, N622, N4063);
xor XOR2 (N5822, N5805, N4168);
nand NAND3 (N5823, N5821, N3718, N5764);
and AND4 (N5824, N5822, N4443, N814, N3349);
buf BUF1 (N5825, N5820);
or OR2 (N5826, N5815, N2632);
and AND2 (N5827, N5824, N2552);
nand NAND3 (N5828, N5808, N870, N4224);
nand NAND2 (N5829, N5818, N4538);
nand NAND3 (N5830, N5826, N1232, N3185);
or OR3 (N5831, N5825, N5419, N2288);
nand NAND4 (N5832, N5830, N2134, N3299, N27);
buf BUF1 (N5833, N5832);
or OR4 (N5834, N5817, N3834, N5448, N93);
nand NAND4 (N5835, N5834, N5646, N2553, N189);
xor XOR2 (N5836, N5810, N5053);
or OR2 (N5837, N5835, N5260);
buf BUF1 (N5838, N5831);
buf BUF1 (N5839, N5823);
nor NOR2 (N5840, N5838, N3645);
not NOT1 (N5841, N5837);
xor XOR2 (N5842, N5819, N2507);
xor XOR2 (N5843, N5842, N4655);
nor NOR4 (N5844, N5840, N5626, N1013, N1757);
not NOT1 (N5845, N5829);
not NOT1 (N5846, N5844);
nor NOR3 (N5847, N5833, N4919, N5087);
xor XOR2 (N5848, N5827, N4851);
xor XOR2 (N5849, N5845, N549);
not NOT1 (N5850, N5839);
xor XOR2 (N5851, N5841, N3991);
and AND3 (N5852, N5848, N582, N2744);
and AND2 (N5853, N5850, N2023);
buf BUF1 (N5854, N5809);
buf BUF1 (N5855, N5836);
xor XOR2 (N5856, N5855, N3511);
or OR2 (N5857, N5856, N2256);
not NOT1 (N5858, N5854);
nor NOR2 (N5859, N5858, N1323);
and AND3 (N5860, N5857, N4581, N1977);
or OR3 (N5861, N5828, N5277, N2904);
buf BUF1 (N5862, N5852);
nor NOR2 (N5863, N5849, N5321);
xor XOR2 (N5864, N5860, N5438);
buf BUF1 (N5865, N5846);
not NOT1 (N5866, N5859);
or OR3 (N5867, N5853, N2806, N311);
and AND4 (N5868, N5861, N3957, N1772, N1756);
buf BUF1 (N5869, N5862);
or OR2 (N5870, N5847, N1755);
nand NAND3 (N5871, N5870, N2453, N1353);
or OR3 (N5872, N5868, N861, N1080);
or OR2 (N5873, N5863, N1640);
xor XOR2 (N5874, N5871, N201);
xor XOR2 (N5875, N5869, N4189);
not NOT1 (N5876, N5864);
and AND3 (N5877, N5865, N5317, N5260);
xor XOR2 (N5878, N5873, N4154);
not NOT1 (N5879, N5867);
xor XOR2 (N5880, N5874, N1804);
nand NAND2 (N5881, N5843, N622);
not NOT1 (N5882, N5875);
nand NAND3 (N5883, N5851, N3212, N2079);
buf BUF1 (N5884, N5883);
xor XOR2 (N5885, N5872, N3592);
nand NAND3 (N5886, N5882, N1132, N1336);
and AND4 (N5887, N5880, N5586, N4891, N2625);
buf BUF1 (N5888, N5878);
xor XOR2 (N5889, N5866, N1299);
or OR4 (N5890, N5889, N340, N4391, N16);
buf BUF1 (N5891, N5888);
buf BUF1 (N5892, N5887);
and AND4 (N5893, N5892, N2740, N3629, N618);
xor XOR2 (N5894, N5884, N4380);
not NOT1 (N5895, N5893);
buf BUF1 (N5896, N5876);
nand NAND4 (N5897, N5877, N3692, N402, N4924);
or OR2 (N5898, N5891, N2166);
nand NAND2 (N5899, N5886, N4056);
buf BUF1 (N5900, N5896);
or OR4 (N5901, N5897, N860, N5578, N3975);
nand NAND3 (N5902, N5894, N4726, N3269);
nand NAND2 (N5903, N5899, N3288);
or OR4 (N5904, N5881, N5609, N4890, N418);
buf BUF1 (N5905, N5901);
buf BUF1 (N5906, N5898);
xor XOR2 (N5907, N5890, N2056);
or OR4 (N5908, N5895, N5415, N2999, N55);
nand NAND2 (N5909, N5885, N4368);
xor XOR2 (N5910, N5904, N1541);
nor NOR4 (N5911, N5879, N4080, N139, N1313);
not NOT1 (N5912, N5908);
buf BUF1 (N5913, N5912);
and AND2 (N5914, N5910, N2532);
buf BUF1 (N5915, N5909);
nand NAND4 (N5916, N5905, N1867, N3360, N514);
nor NOR3 (N5917, N5907, N1138, N3198);
nor NOR4 (N5918, N5902, N1472, N5429, N862);
and AND3 (N5919, N5906, N1940, N700);
nor NOR2 (N5920, N5918, N3364);
buf BUF1 (N5921, N5917);
buf BUF1 (N5922, N5915);
nand NAND3 (N5923, N5920, N2885, N550);
nand NAND4 (N5924, N5922, N2717, N5054, N1811);
or OR3 (N5925, N5916, N1075, N2931);
not NOT1 (N5926, N5921);
or OR4 (N5927, N5913, N3433, N4907, N2199);
nand NAND3 (N5928, N5903, N4415, N4323);
not NOT1 (N5929, N5919);
buf BUF1 (N5930, N5923);
nor NOR4 (N5931, N5911, N5912, N1878, N4220);
and AND4 (N5932, N5924, N1880, N2756, N5081);
or OR2 (N5933, N5929, N4892);
not NOT1 (N5934, N5932);
not NOT1 (N5935, N5931);
not NOT1 (N5936, N5935);
buf BUF1 (N5937, N5933);
not NOT1 (N5938, N5930);
not NOT1 (N5939, N5926);
buf BUF1 (N5940, N5936);
buf BUF1 (N5941, N5928);
and AND2 (N5942, N5934, N3122);
or OR2 (N5943, N5925, N2174);
not NOT1 (N5944, N5942);
or OR2 (N5945, N5944, N3202);
or OR4 (N5946, N5937, N3481, N2995, N2951);
nor NOR3 (N5947, N5939, N546, N1603);
nor NOR4 (N5948, N5914, N4577, N4462, N47);
buf BUF1 (N5949, N5938);
or OR4 (N5950, N5900, N2847, N5938, N213);
not NOT1 (N5951, N5946);
and AND4 (N5952, N5951, N1927, N3516, N2967);
and AND2 (N5953, N5927, N2942);
buf BUF1 (N5954, N5945);
xor XOR2 (N5955, N5948, N225);
nand NAND2 (N5956, N5943, N4287);
buf BUF1 (N5957, N5952);
nand NAND3 (N5958, N5947, N1113, N2777);
not NOT1 (N5959, N5950);
buf BUF1 (N5960, N5949);
or OR4 (N5961, N5958, N5087, N5333, N4699);
buf BUF1 (N5962, N5956);
nor NOR4 (N5963, N5940, N18, N5403, N2340);
xor XOR2 (N5964, N5955, N1391);
not NOT1 (N5965, N5953);
nor NOR4 (N5966, N5962, N2450, N2593, N1009);
not NOT1 (N5967, N5961);
xor XOR2 (N5968, N5964, N3198);
not NOT1 (N5969, N5963);
buf BUF1 (N5970, N5959);
nand NAND3 (N5971, N5965, N4727, N4381);
nor NOR2 (N5972, N5966, N1838);
nand NAND4 (N5973, N5971, N5931, N1116, N1875);
or OR3 (N5974, N5954, N4047, N116);
nand NAND4 (N5975, N5970, N2790, N837, N5211);
nand NAND3 (N5976, N5969, N4624, N4936);
or OR2 (N5977, N5941, N3863);
and AND3 (N5978, N5972, N5380, N3275);
xor XOR2 (N5979, N5960, N3805);
nor NOR2 (N5980, N5968, N1545);
nand NAND4 (N5981, N5967, N5287, N3147, N1884);
xor XOR2 (N5982, N5977, N2925);
not NOT1 (N5983, N5974);
nor NOR3 (N5984, N5980, N522, N1900);
and AND4 (N5985, N5981, N5624, N3237, N1834);
or OR2 (N5986, N5957, N5474);
and AND4 (N5987, N5985, N5644, N1003, N870);
xor XOR2 (N5988, N5975, N1353);
xor XOR2 (N5989, N5976, N3756);
not NOT1 (N5990, N5984);
not NOT1 (N5991, N5989);
nand NAND3 (N5992, N5983, N3285, N4004);
nand NAND4 (N5993, N5991, N3672, N56, N3724);
buf BUF1 (N5994, N5986);
nand NAND3 (N5995, N5988, N2780, N4696);
xor XOR2 (N5996, N5994, N5133);
xor XOR2 (N5997, N5987, N187);
xor XOR2 (N5998, N5990, N2158);
nand NAND4 (N5999, N5992, N2511, N616, N2637);
buf BUF1 (N6000, N5973);
xor XOR2 (N6001, N6000, N1961);
buf BUF1 (N6002, N5996);
nor NOR3 (N6003, N5978, N2085, N4848);
nor NOR3 (N6004, N5999, N3400, N224);
xor XOR2 (N6005, N6002, N5632);
or OR3 (N6006, N5997, N5704, N1055);
xor XOR2 (N6007, N6005, N3413);
or OR3 (N6008, N5993, N1662, N5411);
buf BUF1 (N6009, N6001);
buf BUF1 (N6010, N6004);
xor XOR2 (N6011, N5995, N465);
xor XOR2 (N6012, N6003, N3381);
nor NOR2 (N6013, N6009, N371);
nor NOR2 (N6014, N5982, N1134);
or OR4 (N6015, N6008, N5726, N5279, N5442);
buf BUF1 (N6016, N6007);
xor XOR2 (N6017, N6016, N3127);
buf BUF1 (N6018, N6006);
and AND4 (N6019, N6011, N3552, N5989, N568);
nand NAND4 (N6020, N5979, N4868, N2429, N1407);
buf BUF1 (N6021, N6020);
not NOT1 (N6022, N6015);
and AND3 (N6023, N6017, N521, N1474);
not NOT1 (N6024, N6018);
xor XOR2 (N6025, N6023, N3633);
nor NOR3 (N6026, N6014, N5978, N3772);
nor NOR2 (N6027, N6021, N5272);
xor XOR2 (N6028, N6010, N4250);
nor NOR3 (N6029, N6028, N693, N627);
nand NAND2 (N6030, N6026, N2735);
nand NAND2 (N6031, N6012, N484);
not NOT1 (N6032, N6022);
xor XOR2 (N6033, N6030, N228);
or OR4 (N6034, N6029, N4185, N1095, N4984);
or OR3 (N6035, N6024, N4034, N3526);
and AND2 (N6036, N6032, N51);
xor XOR2 (N6037, N6035, N990);
nor NOR2 (N6038, N6027, N823);
nand NAND2 (N6039, N6034, N1078);
nor NOR3 (N6040, N5998, N2005, N5299);
not NOT1 (N6041, N6038);
nor NOR2 (N6042, N6025, N1064);
and AND4 (N6043, N6041, N4030, N1948, N3887);
nand NAND4 (N6044, N6019, N3400, N2068, N3069);
buf BUF1 (N6045, N6039);
nand NAND3 (N6046, N6036, N4772, N3259);
and AND4 (N6047, N6043, N5130, N1668, N936);
nor NOR4 (N6048, N6044, N1272, N4188, N3488);
xor XOR2 (N6049, N6047, N5584);
buf BUF1 (N6050, N6042);
and AND2 (N6051, N6033, N731);
buf BUF1 (N6052, N6046);
xor XOR2 (N6053, N6052, N1404);
xor XOR2 (N6054, N6051, N4756);
or OR4 (N6055, N6050, N4798, N5646, N4339);
or OR2 (N6056, N6048, N4515);
nor NOR3 (N6057, N6031, N4038, N594);
nand NAND4 (N6058, N6055, N4691, N2590, N496);
not NOT1 (N6059, N6049);
and AND3 (N6060, N6058, N491, N2005);
xor XOR2 (N6061, N6057, N4855);
nand NAND2 (N6062, N6013, N5634);
nand NAND4 (N6063, N6062, N4873, N553, N2054);
xor XOR2 (N6064, N6040, N2604);
not NOT1 (N6065, N6059);
nor NOR2 (N6066, N6060, N3476);
and AND4 (N6067, N6063, N3059, N4408, N1667);
and AND4 (N6068, N6053, N3047, N3783, N5665);
or OR3 (N6069, N6037, N2081, N3344);
nor NOR4 (N6070, N6066, N3989, N3307, N3858);
nor NOR3 (N6071, N6061, N3415, N608);
or OR4 (N6072, N6067, N4195, N3405, N2362);
buf BUF1 (N6073, N6064);
or OR4 (N6074, N6070, N4278, N3120, N3812);
buf BUF1 (N6075, N6069);
and AND4 (N6076, N6054, N2000, N5011, N5004);
nand NAND2 (N6077, N6075, N2142);
nand NAND2 (N6078, N6076, N957);
nor NOR2 (N6079, N6074, N3074);
and AND3 (N6080, N6056, N5749, N1800);
or OR4 (N6081, N6080, N3559, N5641, N3144);
nand NAND3 (N6082, N6077, N5506, N4043);
nor NOR2 (N6083, N6082, N3842);
nor NOR2 (N6084, N6083, N69);
nand NAND4 (N6085, N6081, N1831, N4597, N1260);
or OR4 (N6086, N6073, N86, N431, N3923);
nor NOR4 (N6087, N6071, N4149, N3338, N140);
nand NAND4 (N6088, N6078, N5969, N2511, N5178);
nand NAND4 (N6089, N6086, N3144, N1080, N5318);
xor XOR2 (N6090, N6079, N3595);
and AND2 (N6091, N6088, N4996);
nor NOR3 (N6092, N6091, N5091, N1448);
and AND4 (N6093, N6090, N4150, N2525, N4539);
not NOT1 (N6094, N6068);
nand NAND4 (N6095, N6094, N2025, N4926, N412);
or OR2 (N6096, N6089, N221);
nand NAND2 (N6097, N6084, N5887);
xor XOR2 (N6098, N6087, N3403);
and AND4 (N6099, N6098, N4318, N4637, N323);
and AND4 (N6100, N6085, N1665, N40, N5139);
or OR3 (N6101, N6096, N3652, N1952);
buf BUF1 (N6102, N6065);
and AND4 (N6103, N6093, N1358, N4467, N2265);
nand NAND2 (N6104, N6045, N3182);
nor NOR3 (N6105, N6095, N54, N4186);
xor XOR2 (N6106, N6099, N1116);
not NOT1 (N6107, N6104);
nor NOR2 (N6108, N6102, N800);
xor XOR2 (N6109, N6097, N4912);
and AND2 (N6110, N6103, N2847);
not NOT1 (N6111, N6072);
nand NAND3 (N6112, N6106, N2248, N3742);
or OR2 (N6113, N6112, N2556);
or OR3 (N6114, N6111, N5602, N1287);
nor NOR2 (N6115, N6092, N2794);
and AND2 (N6116, N6108, N2104);
or OR4 (N6117, N6113, N5869, N4700, N191);
buf BUF1 (N6118, N6117);
nand NAND2 (N6119, N6107, N4610);
nand NAND4 (N6120, N6100, N1061, N875, N1649);
nand NAND3 (N6121, N6101, N2489, N1220);
and AND4 (N6122, N6120, N1742, N5955, N5835);
nand NAND4 (N6123, N6116, N3857, N28, N762);
xor XOR2 (N6124, N6109, N3911);
and AND4 (N6125, N6105, N1843, N576, N1689);
nor NOR3 (N6126, N6125, N5005, N1221);
or OR4 (N6127, N6124, N4460, N2692, N675);
nor NOR2 (N6128, N6127, N308);
and AND4 (N6129, N6115, N765, N1273, N370);
buf BUF1 (N6130, N6114);
or OR2 (N6131, N6122, N5722);
xor XOR2 (N6132, N6121, N1691);
nor NOR2 (N6133, N6132, N4489);
and AND2 (N6134, N6123, N507);
buf BUF1 (N6135, N6128);
buf BUF1 (N6136, N6126);
nand NAND4 (N6137, N6119, N4484, N1411, N1032);
nand NAND3 (N6138, N6131, N411, N1723);
nor NOR4 (N6139, N6136, N383, N289, N4579);
or OR2 (N6140, N6135, N699);
nand NAND3 (N6141, N6118, N4694, N6059);
and AND3 (N6142, N6140, N5622, N4722);
and AND3 (N6143, N6134, N6093, N4927);
buf BUF1 (N6144, N6139);
and AND2 (N6145, N6110, N4466);
not NOT1 (N6146, N6144);
not NOT1 (N6147, N6129);
or OR2 (N6148, N6141, N5991);
nor NOR4 (N6149, N6142, N4467, N2700, N6103);
buf BUF1 (N6150, N6138);
not NOT1 (N6151, N6148);
nor NOR3 (N6152, N6130, N344, N5817);
and AND3 (N6153, N6151, N5110, N2233);
nor NOR2 (N6154, N6146, N1551);
or OR2 (N6155, N6150, N1988);
and AND4 (N6156, N6154, N878, N5700, N2527);
nand NAND4 (N6157, N6156, N4736, N2531, N1161);
nor NOR2 (N6158, N6147, N2419);
or OR2 (N6159, N6152, N5766);
not NOT1 (N6160, N6158);
xor XOR2 (N6161, N6133, N5402);
nor NOR4 (N6162, N6155, N5388, N5087, N5341);
or OR4 (N6163, N6157, N3132, N3362, N2334);
xor XOR2 (N6164, N6143, N4029);
or OR4 (N6165, N6137, N467, N3073, N5837);
and AND2 (N6166, N6163, N2296);
and AND2 (N6167, N6145, N4638);
and AND3 (N6168, N6153, N2031, N2679);
nand NAND3 (N6169, N6166, N5579, N4048);
nor NOR4 (N6170, N6162, N1366, N5356, N1384);
nand NAND2 (N6171, N6169, N1561);
not NOT1 (N6172, N6159);
buf BUF1 (N6173, N6149);
not NOT1 (N6174, N6167);
and AND3 (N6175, N6170, N173, N3698);
buf BUF1 (N6176, N6168);
buf BUF1 (N6177, N6173);
xor XOR2 (N6178, N6174, N483);
nand NAND3 (N6179, N6160, N505, N5849);
and AND3 (N6180, N6175, N3470, N3982);
and AND4 (N6181, N6177, N3604, N5878, N6024);
not NOT1 (N6182, N6176);
not NOT1 (N6183, N6164);
nand NAND2 (N6184, N6165, N2112);
nand NAND2 (N6185, N6161, N1732);
xor XOR2 (N6186, N6181, N3367);
xor XOR2 (N6187, N6184, N5159);
or OR2 (N6188, N6182, N931);
nand NAND2 (N6189, N6179, N3402);
nor NOR2 (N6190, N6172, N2188);
and AND2 (N6191, N6188, N1879);
buf BUF1 (N6192, N6171);
buf BUF1 (N6193, N6187);
nor NOR4 (N6194, N6192, N244, N460, N4420);
not NOT1 (N6195, N6183);
and AND2 (N6196, N6191, N4521);
xor XOR2 (N6197, N6189, N3621);
nor NOR2 (N6198, N6180, N5177);
or OR4 (N6199, N6186, N2130, N4869, N4812);
buf BUF1 (N6200, N6193);
or OR2 (N6201, N6178, N5884);
not NOT1 (N6202, N6199);
or OR3 (N6203, N6195, N5462, N432);
nand NAND2 (N6204, N6202, N3413);
xor XOR2 (N6205, N6197, N4792);
or OR2 (N6206, N6198, N4679);
xor XOR2 (N6207, N6201, N4999);
or OR4 (N6208, N6200, N4021, N2125, N4692);
not NOT1 (N6209, N6204);
or OR2 (N6210, N6208, N286);
not NOT1 (N6211, N6207);
nand NAND3 (N6212, N6209, N3768, N1648);
buf BUF1 (N6213, N6205);
buf BUF1 (N6214, N6194);
nand NAND2 (N6215, N6203, N3013);
or OR4 (N6216, N6214, N924, N5662, N3507);
or OR3 (N6217, N6185, N1365, N3211);
not NOT1 (N6218, N6217);
nor NOR3 (N6219, N6210, N2740, N3455);
nand NAND4 (N6220, N6190, N3008, N3792, N3441);
not NOT1 (N6221, N6218);
buf BUF1 (N6222, N6216);
not NOT1 (N6223, N6221);
xor XOR2 (N6224, N6220, N658);
or OR4 (N6225, N6213, N5381, N4707, N5026);
buf BUF1 (N6226, N6223);
and AND4 (N6227, N6196, N286, N5194, N6152);
xor XOR2 (N6228, N6222, N5467);
or OR4 (N6229, N6219, N42, N3498, N4756);
buf BUF1 (N6230, N6224);
nor NOR3 (N6231, N6211, N3639, N3829);
and AND3 (N6232, N6226, N3099, N5050);
not NOT1 (N6233, N6206);
nand NAND4 (N6234, N6228, N122, N541, N2613);
or OR3 (N6235, N6234, N3322, N958);
buf BUF1 (N6236, N6212);
buf BUF1 (N6237, N6230);
not NOT1 (N6238, N6236);
nand NAND4 (N6239, N6231, N5686, N1818, N4734);
and AND3 (N6240, N6215, N5129, N2640);
nor NOR3 (N6241, N6229, N4262, N4238);
buf BUF1 (N6242, N6227);
nor NOR4 (N6243, N6235, N3010, N3966, N3404);
and AND3 (N6244, N6233, N2116, N1762);
nand NAND2 (N6245, N6242, N5689);
nand NAND2 (N6246, N6240, N1059);
nand NAND3 (N6247, N6244, N5787, N5317);
buf BUF1 (N6248, N6232);
nor NOR4 (N6249, N6246, N2918, N3202, N4298);
xor XOR2 (N6250, N6249, N4277);
buf BUF1 (N6251, N6239);
nand NAND3 (N6252, N6241, N393, N4487);
nor NOR3 (N6253, N6251, N439, N5503);
nand NAND4 (N6254, N6247, N5047, N2510, N5537);
buf BUF1 (N6255, N6250);
buf BUF1 (N6256, N6254);
nand NAND3 (N6257, N6245, N4108, N2723);
and AND2 (N6258, N6248, N5894);
nor NOR2 (N6259, N6238, N5253);
nand NAND4 (N6260, N6253, N2545, N3694, N4169);
nor NOR4 (N6261, N6252, N4581, N997, N5513);
xor XOR2 (N6262, N6259, N1860);
not NOT1 (N6263, N6237);
nand NAND4 (N6264, N6260, N2117, N4333, N1202);
nor NOR2 (N6265, N6225, N415);
nor NOR2 (N6266, N6263, N4261);
or OR4 (N6267, N6256, N534, N661, N3185);
xor XOR2 (N6268, N6265, N3479);
not NOT1 (N6269, N6267);
or OR3 (N6270, N6262, N3936, N4638);
and AND3 (N6271, N6243, N3591, N5685);
buf BUF1 (N6272, N6269);
or OR3 (N6273, N6271, N4321, N1178);
nor NOR2 (N6274, N6270, N295);
xor XOR2 (N6275, N6273, N5968);
and AND4 (N6276, N6264, N1792, N3200, N3116);
xor XOR2 (N6277, N6258, N5384);
nand NAND4 (N6278, N6272, N5447, N4651, N2428);
nand NAND3 (N6279, N6266, N5944, N2646);
buf BUF1 (N6280, N6261);
not NOT1 (N6281, N6257);
or OR2 (N6282, N6276, N104);
nand NAND3 (N6283, N6274, N3423, N2143);
buf BUF1 (N6284, N6281);
and AND2 (N6285, N6255, N3814);
xor XOR2 (N6286, N6275, N2318);
not NOT1 (N6287, N6280);
not NOT1 (N6288, N6282);
nor NOR2 (N6289, N6279, N2940);
nor NOR2 (N6290, N6284, N617);
nor NOR3 (N6291, N6283, N5982, N3208);
nand NAND3 (N6292, N6278, N4271, N423);
nor NOR2 (N6293, N6288, N4043);
or OR2 (N6294, N6285, N2339);
nor NOR3 (N6295, N6291, N6053, N1481);
xor XOR2 (N6296, N6286, N1008);
or OR3 (N6297, N6277, N5917, N2335);
not NOT1 (N6298, N6268);
or OR3 (N6299, N6297, N3158, N2126);
or OR3 (N6300, N6292, N3658, N1749);
or OR4 (N6301, N6289, N5235, N1175, N2682);
buf BUF1 (N6302, N6301);
nand NAND3 (N6303, N6300, N2304, N4108);
nor NOR3 (N6304, N6303, N4135, N1126);
or OR4 (N6305, N6298, N5210, N2876, N5609);
xor XOR2 (N6306, N6290, N4136);
and AND4 (N6307, N6293, N3593, N1749, N727);
buf BUF1 (N6308, N6287);
nand NAND3 (N6309, N6305, N3663, N3063);
xor XOR2 (N6310, N6304, N4217);
nand NAND4 (N6311, N6306, N3129, N4337, N2151);
not NOT1 (N6312, N6308);
not NOT1 (N6313, N6302);
nand NAND4 (N6314, N6307, N3972, N892, N4338);
and AND3 (N6315, N6310, N2444, N1065);
not NOT1 (N6316, N6309);
nand NAND3 (N6317, N6294, N410, N4256);
and AND4 (N6318, N6314, N89, N5267, N2216);
nand NAND2 (N6319, N6317, N4620);
and AND2 (N6320, N6312, N1931);
and AND4 (N6321, N6311, N1488, N4707, N5375);
nand NAND2 (N6322, N6315, N1224);
buf BUF1 (N6323, N6299);
nor NOR2 (N6324, N6321, N5428);
or OR4 (N6325, N6323, N2062, N3589, N3968);
xor XOR2 (N6326, N6318, N5240);
nor NOR4 (N6327, N6313, N5684, N2355, N4843);
nand NAND2 (N6328, N6326, N4535);
nor NOR2 (N6329, N6320, N1623);
nand NAND3 (N6330, N6319, N4354, N3092);
xor XOR2 (N6331, N6322, N5540);
and AND4 (N6332, N6330, N4331, N1759, N3169);
nand NAND4 (N6333, N6329, N5693, N4370, N3602);
nor NOR3 (N6334, N6327, N4552, N355);
or OR3 (N6335, N6325, N781, N3366);
or OR4 (N6336, N6316, N1861, N2850, N1882);
xor XOR2 (N6337, N6331, N2771);
xor XOR2 (N6338, N6332, N3771);
xor XOR2 (N6339, N6333, N5596);
nand NAND2 (N6340, N6337, N3407);
or OR3 (N6341, N6324, N2338, N4835);
not NOT1 (N6342, N6334);
nor NOR4 (N6343, N6338, N1582, N1266, N6028);
nor NOR3 (N6344, N6339, N2980, N686);
nor NOR3 (N6345, N6341, N2336, N3965);
nand NAND4 (N6346, N6335, N6139, N4684, N915);
or OR4 (N6347, N6346, N821, N4734, N287);
xor XOR2 (N6348, N6344, N5634);
or OR3 (N6349, N6340, N5214, N610);
xor XOR2 (N6350, N6349, N8);
nand NAND4 (N6351, N6345, N4505, N1606, N6241);
not NOT1 (N6352, N6347);
or OR4 (N6353, N6336, N4987, N6057, N161);
xor XOR2 (N6354, N6348, N6150);
xor XOR2 (N6355, N6353, N4768);
buf BUF1 (N6356, N6352);
and AND2 (N6357, N6355, N6093);
nor NOR4 (N6358, N6342, N4979, N2781, N1648);
or OR3 (N6359, N6328, N6122, N2086);
or OR4 (N6360, N6357, N532, N3664, N4039);
buf BUF1 (N6361, N6360);
and AND3 (N6362, N6351, N1495, N3287);
buf BUF1 (N6363, N6362);
xor XOR2 (N6364, N6356, N6257);
xor XOR2 (N6365, N6358, N3055);
not NOT1 (N6366, N6361);
buf BUF1 (N6367, N6359);
nand NAND4 (N6368, N6365, N2894, N264, N1586);
or OR2 (N6369, N6367, N4722);
nand NAND4 (N6370, N6295, N5669, N3843, N3534);
and AND4 (N6371, N6363, N4950, N1142, N1967);
and AND3 (N6372, N6368, N2507, N5313);
nor NOR3 (N6373, N6370, N3668, N5735);
xor XOR2 (N6374, N6343, N2877);
buf BUF1 (N6375, N6374);
and AND3 (N6376, N6371, N4256, N2133);
or OR4 (N6377, N6373, N4653, N712, N1633);
xor XOR2 (N6378, N6369, N4238);
nor NOR2 (N6379, N6372, N1072);
or OR4 (N6380, N6375, N2429, N4875, N564);
xor XOR2 (N6381, N6354, N4776);
buf BUF1 (N6382, N6366);
not NOT1 (N6383, N6350);
nor NOR2 (N6384, N6364, N5395);
or OR4 (N6385, N6379, N6320, N3648, N2690);
xor XOR2 (N6386, N6296, N1782);
and AND3 (N6387, N6384, N468, N6167);
not NOT1 (N6388, N6383);
buf BUF1 (N6389, N6386);
nand NAND2 (N6390, N6389, N1515);
nor NOR4 (N6391, N6380, N947, N3708, N37);
not NOT1 (N6392, N6388);
buf BUF1 (N6393, N6382);
buf BUF1 (N6394, N6378);
buf BUF1 (N6395, N6393);
buf BUF1 (N6396, N6376);
not NOT1 (N6397, N6387);
buf BUF1 (N6398, N6377);
nand NAND3 (N6399, N6391, N3963, N4521);
nor NOR4 (N6400, N6397, N5843, N4752, N720);
xor XOR2 (N6401, N6394, N1012);
nand NAND3 (N6402, N6396, N3892, N4038);
nand NAND2 (N6403, N6395, N1312);
not NOT1 (N6404, N6401);
xor XOR2 (N6405, N6404, N39);
xor XOR2 (N6406, N6400, N1556);
nand NAND4 (N6407, N6390, N1277, N2547, N5217);
nor NOR4 (N6408, N6403, N531, N6352, N2897);
not NOT1 (N6409, N6399);
nor NOR4 (N6410, N6381, N354, N5391, N1429);
buf BUF1 (N6411, N6398);
buf BUF1 (N6412, N6392);
nor NOR4 (N6413, N6410, N3850, N2015, N3934);
buf BUF1 (N6414, N6406);
nor NOR4 (N6415, N6414, N4646, N633, N1876);
nor NOR4 (N6416, N6412, N5595, N3603, N6357);
buf BUF1 (N6417, N6402);
xor XOR2 (N6418, N6416, N3808);
or OR2 (N6419, N6418, N5315);
buf BUF1 (N6420, N6408);
or OR3 (N6421, N6411, N709, N5713);
and AND4 (N6422, N6413, N980, N2535, N4441);
or OR4 (N6423, N6417, N1951, N300, N5870);
and AND2 (N6424, N6385, N2444);
or OR4 (N6425, N6420, N4865, N3078, N1316);
nand NAND4 (N6426, N6419, N1193, N1277, N649);
nor NOR4 (N6427, N6405, N1754, N4057, N3536);
or OR2 (N6428, N6422, N1341);
not NOT1 (N6429, N6421);
buf BUF1 (N6430, N6429);
and AND4 (N6431, N6430, N5244, N2331, N4434);
nor NOR3 (N6432, N6415, N1185, N2400);
nor NOR4 (N6433, N6427, N222, N2308, N4906);
buf BUF1 (N6434, N6407);
buf BUF1 (N6435, N6431);
or OR2 (N6436, N6425, N4164);
nand NAND4 (N6437, N6432, N4092, N1500, N2036);
and AND2 (N6438, N6409, N3089);
xor XOR2 (N6439, N6438, N2937);
nor NOR3 (N6440, N6434, N4501, N4776);
buf BUF1 (N6441, N6423);
nand NAND4 (N6442, N6433, N4040, N2374, N2566);
nand NAND2 (N6443, N6441, N3725);
nand NAND4 (N6444, N6443, N4702, N1786, N3143);
xor XOR2 (N6445, N6428, N4236);
nor NOR4 (N6446, N6437, N2930, N2260, N4777);
buf BUF1 (N6447, N6436);
and AND2 (N6448, N6444, N473);
buf BUF1 (N6449, N6435);
nor NOR3 (N6450, N6442, N1228, N4921);
and AND4 (N6451, N6440, N2562, N158, N136);
not NOT1 (N6452, N6424);
and AND3 (N6453, N6426, N4671, N4256);
xor XOR2 (N6454, N6448, N3386);
buf BUF1 (N6455, N6446);
nor NOR3 (N6456, N6452, N1570, N974);
and AND3 (N6457, N6455, N3474, N1618);
xor XOR2 (N6458, N6439, N3323);
and AND2 (N6459, N6458, N1225);
and AND4 (N6460, N6459, N3028, N1362, N3578);
buf BUF1 (N6461, N6457);
nor NOR2 (N6462, N6453, N2593);
or OR3 (N6463, N6445, N2018, N2746);
not NOT1 (N6464, N6463);
nand NAND3 (N6465, N6456, N2081, N1511);
buf BUF1 (N6466, N6461);
xor XOR2 (N6467, N6454, N2447);
or OR3 (N6468, N6451, N4658, N1188);
nand NAND4 (N6469, N6464, N3569, N3742, N2730);
and AND2 (N6470, N6468, N3388);
not NOT1 (N6471, N6467);
xor XOR2 (N6472, N6447, N5489);
nor NOR2 (N6473, N6462, N5062);
not NOT1 (N6474, N6450);
and AND2 (N6475, N6466, N5196);
and AND2 (N6476, N6470, N259);
and AND3 (N6477, N6473, N4390, N3083);
nand NAND2 (N6478, N6476, N6344);
nand NAND3 (N6479, N6475, N3520, N3184);
not NOT1 (N6480, N6460);
not NOT1 (N6481, N6479);
buf BUF1 (N6482, N6481);
xor XOR2 (N6483, N6471, N3351);
and AND2 (N6484, N6478, N4144);
nor NOR4 (N6485, N6477, N5297, N218, N5346);
not NOT1 (N6486, N6484);
nor NOR4 (N6487, N6483, N404, N470, N2299);
not NOT1 (N6488, N6474);
nor NOR3 (N6489, N6487, N5046, N3208);
xor XOR2 (N6490, N6482, N5764);
and AND2 (N6491, N6490, N2549);
xor XOR2 (N6492, N6486, N5599);
or OR3 (N6493, N6465, N1603, N4119);
xor XOR2 (N6494, N6469, N5969);
and AND2 (N6495, N6493, N4903);
and AND4 (N6496, N6488, N608, N112, N484);
xor XOR2 (N6497, N6480, N520);
buf BUF1 (N6498, N6495);
and AND3 (N6499, N6485, N1195, N1855);
xor XOR2 (N6500, N6491, N3099);
xor XOR2 (N6501, N6498, N3852);
xor XOR2 (N6502, N6497, N4427);
and AND3 (N6503, N6449, N1817, N2005);
not NOT1 (N6504, N6502);
or OR4 (N6505, N6499, N1384, N6462, N121);
nor NOR3 (N6506, N6503, N1316, N504);
or OR2 (N6507, N6505, N5376);
buf BUF1 (N6508, N6496);
not NOT1 (N6509, N6489);
buf BUF1 (N6510, N6507);
buf BUF1 (N6511, N6510);
not NOT1 (N6512, N6509);
nand NAND4 (N6513, N6508, N3806, N3477, N6084);
xor XOR2 (N6514, N6511, N2160);
or OR3 (N6515, N6492, N6362, N2214);
not NOT1 (N6516, N6494);
and AND3 (N6517, N6514, N1875, N3717);
and AND2 (N6518, N6506, N41);
and AND3 (N6519, N6516, N1069, N3926);
not NOT1 (N6520, N6519);
and AND2 (N6521, N6517, N6087);
nand NAND2 (N6522, N6501, N1492);
or OR4 (N6523, N6515, N51, N3821, N2839);
buf BUF1 (N6524, N6472);
and AND3 (N6525, N6513, N1848, N6476);
buf BUF1 (N6526, N6504);
or OR2 (N6527, N6522, N5613);
nor NOR2 (N6528, N6523, N4862);
xor XOR2 (N6529, N6520, N2765);
xor XOR2 (N6530, N6524, N1391);
nor NOR2 (N6531, N6525, N927);
and AND4 (N6532, N6531, N5771, N4858, N3442);
xor XOR2 (N6533, N6521, N517);
and AND3 (N6534, N6500, N4689, N439);
not NOT1 (N6535, N6527);
and AND2 (N6536, N6518, N4661);
not NOT1 (N6537, N6512);
not NOT1 (N6538, N6529);
nor NOR3 (N6539, N6533, N5305, N3469);
and AND2 (N6540, N6528, N5756);
xor XOR2 (N6541, N6540, N3245);
nor NOR2 (N6542, N6526, N1467);
xor XOR2 (N6543, N6539, N5942);
or OR2 (N6544, N6542, N4717);
nor NOR3 (N6545, N6544, N485, N2743);
buf BUF1 (N6546, N6535);
not NOT1 (N6547, N6543);
nor NOR4 (N6548, N6530, N2572, N90, N3456);
xor XOR2 (N6549, N6541, N4831);
and AND3 (N6550, N6536, N3150, N691);
nand NAND4 (N6551, N6532, N1147, N2040, N6488);
nand NAND4 (N6552, N6547, N4722, N1203, N348);
not NOT1 (N6553, N6545);
nor NOR4 (N6554, N6552, N3262, N2921, N485);
nor NOR3 (N6555, N6548, N6391, N1768);
nor NOR2 (N6556, N6555, N112);
buf BUF1 (N6557, N6556);
xor XOR2 (N6558, N6537, N3598);
not NOT1 (N6559, N6534);
or OR3 (N6560, N6538, N2754, N1842);
buf BUF1 (N6561, N6554);
nand NAND2 (N6562, N6557, N4240);
xor XOR2 (N6563, N6551, N3331);
not NOT1 (N6564, N6561);
buf BUF1 (N6565, N6558);
not NOT1 (N6566, N6549);
buf BUF1 (N6567, N6559);
and AND4 (N6568, N6567, N3250, N1397, N4626);
buf BUF1 (N6569, N6550);
nor NOR4 (N6570, N6546, N5829, N4310, N2771);
or OR2 (N6571, N6560, N3951);
xor XOR2 (N6572, N6566, N4594);
nor NOR3 (N6573, N6553, N1995, N5683);
and AND4 (N6574, N6565, N397, N2407, N2913);
not NOT1 (N6575, N6562);
or OR2 (N6576, N6572, N542);
nor NOR2 (N6577, N6576, N5055);
and AND3 (N6578, N6573, N427, N5819);
nor NOR2 (N6579, N6571, N67);
not NOT1 (N6580, N6563);
and AND2 (N6581, N6578, N5908);
or OR3 (N6582, N6577, N6515, N33);
and AND2 (N6583, N6568, N1659);
buf BUF1 (N6584, N6564);
and AND2 (N6585, N6580, N2495);
nor NOR2 (N6586, N6574, N5272);
buf BUF1 (N6587, N6570);
or OR3 (N6588, N6584, N4601, N6031);
buf BUF1 (N6589, N6579);
nor NOR4 (N6590, N6575, N2490, N3322, N3090);
xor XOR2 (N6591, N6582, N1078);
or OR4 (N6592, N6590, N5989, N6194, N2170);
nand NAND4 (N6593, N6583, N818, N698, N4582);
or OR2 (N6594, N6589, N2531);
or OR4 (N6595, N6587, N2650, N2104, N6282);
nand NAND4 (N6596, N6592, N3966, N688, N5974);
nand NAND4 (N6597, N6585, N5321, N3313, N3207);
nor NOR2 (N6598, N6569, N4218);
nor NOR2 (N6599, N6597, N2561);
not NOT1 (N6600, N6588);
not NOT1 (N6601, N6599);
not NOT1 (N6602, N6581);
or OR2 (N6603, N6602, N2952);
and AND4 (N6604, N6600, N4191, N1744, N684);
and AND3 (N6605, N6596, N3573, N4973);
not NOT1 (N6606, N6605);
nand NAND4 (N6607, N6595, N3617, N6459, N4664);
nor NOR3 (N6608, N6606, N5294, N1654);
xor XOR2 (N6609, N6586, N1305);
xor XOR2 (N6610, N6603, N4580);
nor NOR2 (N6611, N6601, N2044);
xor XOR2 (N6612, N6608, N5852);
not NOT1 (N6613, N6611);
not NOT1 (N6614, N6613);
and AND3 (N6615, N6604, N238, N1962);
xor XOR2 (N6616, N6610, N2089);
nor NOR4 (N6617, N6612, N1896, N6493, N3540);
and AND3 (N6618, N6616, N2032, N6524);
and AND2 (N6619, N6591, N180);
buf BUF1 (N6620, N6609);
nor NOR3 (N6621, N6598, N4121, N683);
not NOT1 (N6622, N6617);
nor NOR3 (N6623, N6620, N2545, N5856);
nand NAND4 (N6624, N6594, N3227, N775, N6570);
and AND3 (N6625, N6614, N3226, N1517);
and AND2 (N6626, N6625, N3466);
and AND3 (N6627, N6622, N6268, N2432);
buf BUF1 (N6628, N6624);
nor NOR3 (N6629, N6615, N6019, N4752);
or OR3 (N6630, N6593, N82, N4971);
nor NOR2 (N6631, N6629, N6314);
buf BUF1 (N6632, N6628);
or OR4 (N6633, N6631, N3988, N2195, N6174);
buf BUF1 (N6634, N6623);
not NOT1 (N6635, N6607);
nand NAND3 (N6636, N6621, N5269, N3201);
nor NOR4 (N6637, N6634, N2035, N5256, N6221);
and AND3 (N6638, N6630, N4269, N1101);
not NOT1 (N6639, N6635);
or OR4 (N6640, N6633, N1155, N5984, N5500);
and AND4 (N6641, N6637, N448, N5242, N1084);
nor NOR2 (N6642, N6619, N596);
not NOT1 (N6643, N6642);
or OR4 (N6644, N6641, N129, N863, N5758);
xor XOR2 (N6645, N6626, N899);
or OR3 (N6646, N6618, N5478, N1623);
xor XOR2 (N6647, N6644, N4703);
nor NOR3 (N6648, N6627, N3934, N3986);
buf BUF1 (N6649, N6636);
nor NOR2 (N6650, N6646, N3047);
xor XOR2 (N6651, N6638, N2654);
and AND4 (N6652, N6632, N1141, N3062, N1691);
or OR4 (N6653, N6640, N2648, N4999, N3634);
and AND3 (N6654, N6653, N6305, N4460);
nand NAND3 (N6655, N6651, N1259, N397);
xor XOR2 (N6656, N6645, N5517);
buf BUF1 (N6657, N6650);
xor XOR2 (N6658, N6657, N3444);
and AND2 (N6659, N6658, N6463);
buf BUF1 (N6660, N6655);
nand NAND2 (N6661, N6652, N5885);
nor NOR2 (N6662, N6660, N3060);
or OR3 (N6663, N6656, N3013, N1856);
not NOT1 (N6664, N6663);
not NOT1 (N6665, N6643);
and AND2 (N6666, N6639, N3203);
buf BUF1 (N6667, N6664);
xor XOR2 (N6668, N6661, N6387);
xor XOR2 (N6669, N6668, N4517);
xor XOR2 (N6670, N6669, N5944);
buf BUF1 (N6671, N6665);
nor NOR2 (N6672, N6662, N5345);
not NOT1 (N6673, N6654);
or OR3 (N6674, N6649, N5375, N2112);
xor XOR2 (N6675, N6674, N3817);
or OR3 (N6676, N6667, N6046, N1792);
buf BUF1 (N6677, N6672);
xor XOR2 (N6678, N6659, N288);
and AND4 (N6679, N6678, N119, N3847, N4191);
not NOT1 (N6680, N6648);
nand NAND3 (N6681, N6679, N328, N2588);
nor NOR4 (N6682, N6647, N2253, N4634, N451);
nor NOR2 (N6683, N6681, N733);
buf BUF1 (N6684, N6670);
and AND4 (N6685, N6680, N1393, N5259, N4407);
not NOT1 (N6686, N6685);
or OR2 (N6687, N6683, N2603);
not NOT1 (N6688, N6673);
buf BUF1 (N6689, N6675);
nand NAND4 (N6690, N6677, N2177, N1822, N5033);
not NOT1 (N6691, N6671);
nor NOR2 (N6692, N6690, N763);
xor XOR2 (N6693, N6687, N2900);
not NOT1 (N6694, N6693);
not NOT1 (N6695, N6689);
buf BUF1 (N6696, N6676);
buf BUF1 (N6697, N6684);
or OR4 (N6698, N6696, N5205, N3945, N1176);
xor XOR2 (N6699, N6697, N1530);
nor NOR3 (N6700, N6691, N4434, N2893);
or OR3 (N6701, N6695, N2238, N387);
and AND2 (N6702, N6701, N2466);
and AND4 (N6703, N6700, N526, N4677, N6041);
not NOT1 (N6704, N6694);
and AND4 (N6705, N6688, N3437, N5286, N28);
not NOT1 (N6706, N6686);
or OR3 (N6707, N6692, N5565, N1178);
or OR3 (N6708, N6666, N655, N5180);
nor NOR2 (N6709, N6708, N161);
and AND2 (N6710, N6707, N5655);
and AND3 (N6711, N6698, N4368, N2731);
xor XOR2 (N6712, N6702, N4267);
not NOT1 (N6713, N6709);
xor XOR2 (N6714, N6682, N2250);
and AND2 (N6715, N6710, N6534);
nor NOR2 (N6716, N6706, N4721);
buf BUF1 (N6717, N6716);
xor XOR2 (N6718, N6717, N1758);
and AND4 (N6719, N6699, N3730, N3966, N4902);
or OR4 (N6720, N6704, N4821, N5280, N3806);
nor NOR2 (N6721, N6711, N408);
xor XOR2 (N6722, N6712, N1650);
xor XOR2 (N6723, N6721, N3849);
nor NOR4 (N6724, N6705, N2316, N4325, N3930);
xor XOR2 (N6725, N6713, N920);
nand NAND3 (N6726, N6723, N3079, N5028);
and AND3 (N6727, N6725, N4622, N1304);
or OR3 (N6728, N6724, N1475, N1970);
buf BUF1 (N6729, N6722);
not NOT1 (N6730, N6703);
nor NOR2 (N6731, N6714, N5470);
or OR2 (N6732, N6730, N3114);
xor XOR2 (N6733, N6727, N6103);
or OR3 (N6734, N6720, N2208, N5727);
nor NOR3 (N6735, N6731, N3803, N5447);
nor NOR4 (N6736, N6732, N157, N443, N1377);
nor NOR3 (N6737, N6719, N6449, N648);
not NOT1 (N6738, N6728);
xor XOR2 (N6739, N6735, N3378);
not NOT1 (N6740, N6736);
not NOT1 (N6741, N6729);
nor NOR3 (N6742, N6718, N1157, N6093);
and AND3 (N6743, N6733, N73, N5812);
nand NAND4 (N6744, N6738, N3571, N4205, N2588);
and AND3 (N6745, N6739, N5010, N4415);
or OR3 (N6746, N6740, N3580, N1328);
buf BUF1 (N6747, N6746);
not NOT1 (N6748, N6734);
buf BUF1 (N6749, N6748);
buf BUF1 (N6750, N6726);
xor XOR2 (N6751, N6715, N783);
not NOT1 (N6752, N6743);
xor XOR2 (N6753, N6742, N4927);
buf BUF1 (N6754, N6744);
not NOT1 (N6755, N6754);
nand NAND2 (N6756, N6751, N4544);
nand NAND4 (N6757, N6755, N1299, N4018, N1360);
or OR3 (N6758, N6753, N126, N4910);
or OR2 (N6759, N6741, N6665);
nor NOR2 (N6760, N6749, N2138);
nor NOR3 (N6761, N6760, N5479, N3628);
or OR4 (N6762, N6761, N2811, N5790, N3261);
nor NOR3 (N6763, N6756, N2463, N6046);
nand NAND2 (N6764, N6763, N6130);
and AND2 (N6765, N6737, N1123);
not NOT1 (N6766, N6758);
xor XOR2 (N6767, N6762, N2466);
or OR4 (N6768, N6764, N1538, N1065, N5604);
or OR2 (N6769, N6745, N2914);
nand NAND4 (N6770, N6750, N1526, N3696, N4421);
not NOT1 (N6771, N6768);
not NOT1 (N6772, N6770);
nand NAND3 (N6773, N6757, N2554, N4274);
and AND3 (N6774, N6769, N5238, N3967);
not NOT1 (N6775, N6774);
not NOT1 (N6776, N6767);
and AND4 (N6777, N6775, N1898, N4810, N4430);
not NOT1 (N6778, N6776);
xor XOR2 (N6779, N6772, N5576);
and AND2 (N6780, N6766, N6505);
nor NOR4 (N6781, N6773, N4777, N3778, N6006);
nor NOR3 (N6782, N6779, N1080, N6661);
not NOT1 (N6783, N6782);
not NOT1 (N6784, N6781);
buf BUF1 (N6785, N6778);
nand NAND3 (N6786, N6765, N2801, N5916);
not NOT1 (N6787, N6786);
not NOT1 (N6788, N6783);
or OR2 (N6789, N6780, N200);
nor NOR3 (N6790, N6788, N1005, N694);
nand NAND3 (N6791, N6759, N3807, N4470);
nand NAND3 (N6792, N6789, N6113, N4864);
not NOT1 (N6793, N6771);
nor NOR4 (N6794, N6752, N4953, N6436, N3775);
or OR4 (N6795, N6791, N2505, N6544, N1988);
nor NOR3 (N6796, N6784, N2902, N780);
buf BUF1 (N6797, N6792);
or OR2 (N6798, N6794, N642);
nand NAND4 (N6799, N6777, N6107, N4589, N5919);
or OR3 (N6800, N6787, N3234, N6120);
buf BUF1 (N6801, N6793);
nor NOR2 (N6802, N6800, N2303);
xor XOR2 (N6803, N6795, N6120);
and AND4 (N6804, N6801, N4786, N4132, N1075);
or OR4 (N6805, N6799, N5079, N227, N2361);
nand NAND3 (N6806, N6798, N4576, N2109);
nor NOR3 (N6807, N6790, N6492, N5749);
nor NOR3 (N6808, N6796, N3574, N6347);
nand NAND3 (N6809, N6807, N4016, N1798);
nand NAND3 (N6810, N6802, N3790, N4964);
and AND2 (N6811, N6804, N3785);
nor NOR2 (N6812, N6785, N1283);
nor NOR4 (N6813, N6808, N1815, N4170, N64);
nor NOR2 (N6814, N6809, N4008);
or OR4 (N6815, N6805, N1063, N147, N3744);
xor XOR2 (N6816, N6806, N1818);
or OR3 (N6817, N6747, N582, N2921);
xor XOR2 (N6818, N6810, N3208);
or OR2 (N6819, N6817, N5665);
buf BUF1 (N6820, N6812);
buf BUF1 (N6821, N6813);
buf BUF1 (N6822, N6820);
xor XOR2 (N6823, N6814, N4734);
buf BUF1 (N6824, N6816);
xor XOR2 (N6825, N6821, N6726);
or OR2 (N6826, N6823, N1517);
and AND4 (N6827, N6825, N57, N156, N3249);
nand NAND4 (N6828, N6811, N5787, N5238, N5731);
not NOT1 (N6829, N6827);
nor NOR3 (N6830, N6824, N163, N5120);
nand NAND2 (N6831, N6815, N3488);
nand NAND2 (N6832, N6830, N4633);
nor NOR2 (N6833, N6818, N6199);
or OR4 (N6834, N6822, N470, N3709, N3081);
buf BUF1 (N6835, N6803);
and AND4 (N6836, N6832, N2510, N5249, N688);
nor NOR3 (N6837, N6797, N4231, N5970);
xor XOR2 (N6838, N6829, N3690);
nand NAND2 (N6839, N6837, N2621);
not NOT1 (N6840, N6836);
or OR3 (N6841, N6834, N3331, N2103);
xor XOR2 (N6842, N6835, N4195);
nand NAND4 (N6843, N6838, N5681, N3874, N563);
xor XOR2 (N6844, N6819, N4427);
not NOT1 (N6845, N6826);
xor XOR2 (N6846, N6840, N4379);
buf BUF1 (N6847, N6833);
and AND2 (N6848, N6847, N1865);
nor NOR4 (N6849, N6842, N1147, N1731, N2950);
and AND3 (N6850, N6828, N3436, N1612);
and AND3 (N6851, N6849, N3205, N4790);
or OR3 (N6852, N6848, N5939, N5246);
or OR3 (N6853, N6846, N812, N3273);
buf BUF1 (N6854, N6853);
buf BUF1 (N6855, N6851);
buf BUF1 (N6856, N6845);
buf BUF1 (N6857, N6850);
nor NOR3 (N6858, N6841, N932, N249);
xor XOR2 (N6859, N6854, N2777);
not NOT1 (N6860, N6839);
and AND3 (N6861, N6857, N3084, N2623);
or OR3 (N6862, N6843, N5454, N4450);
not NOT1 (N6863, N6852);
and AND2 (N6864, N6861, N6537);
nor NOR4 (N6865, N6863, N6707, N5791, N5810);
not NOT1 (N6866, N6858);
buf BUF1 (N6867, N6844);
nand NAND4 (N6868, N6855, N2764, N5228, N2755);
not NOT1 (N6869, N6866);
xor XOR2 (N6870, N6856, N4873);
or OR4 (N6871, N6864, N3679, N4361, N5379);
buf BUF1 (N6872, N6871);
not NOT1 (N6873, N6862);
and AND2 (N6874, N6860, N4254);
and AND3 (N6875, N6874, N4072, N5562);
xor XOR2 (N6876, N6865, N2285);
and AND4 (N6877, N6831, N5903, N1195, N281);
nor NOR2 (N6878, N6873, N5035);
buf BUF1 (N6879, N6867);
nor NOR2 (N6880, N6872, N3305);
and AND2 (N6881, N6869, N1404);
not NOT1 (N6882, N6881);
xor XOR2 (N6883, N6875, N875);
buf BUF1 (N6884, N6868);
or OR3 (N6885, N6883, N2283, N758);
not NOT1 (N6886, N6884);
not NOT1 (N6887, N6886);
or OR4 (N6888, N6882, N3253, N2129, N1688);
nand NAND2 (N6889, N6880, N1300);
nor NOR2 (N6890, N6876, N6889);
nor NOR4 (N6891, N4349, N5789, N1246, N3169);
or OR3 (N6892, N6888, N4184, N4490);
xor XOR2 (N6893, N6878, N3425);
or OR4 (N6894, N6887, N1050, N1234, N3624);
and AND3 (N6895, N6885, N5791, N2702);
buf BUF1 (N6896, N6890);
and AND2 (N6897, N6895, N3427);
xor XOR2 (N6898, N6870, N1447);
nand NAND4 (N6899, N6893, N5072, N5076, N2621);
xor XOR2 (N6900, N6896, N4952);
not NOT1 (N6901, N6894);
nor NOR4 (N6902, N6891, N5630, N2270, N6660);
buf BUF1 (N6903, N6902);
nand NAND2 (N6904, N6898, N6424);
not NOT1 (N6905, N6877);
buf BUF1 (N6906, N6904);
and AND2 (N6907, N6901, N5849);
xor XOR2 (N6908, N6900, N3414);
nand NAND2 (N6909, N6879, N761);
nand NAND3 (N6910, N6897, N883, N668);
or OR4 (N6911, N6903, N3669, N1317, N5270);
not NOT1 (N6912, N6909);
xor XOR2 (N6913, N6908, N5289);
xor XOR2 (N6914, N6859, N6144);
or OR3 (N6915, N6910, N4141, N3575);
and AND3 (N6916, N6905, N2438, N4795);
nand NAND4 (N6917, N6913, N119, N1108, N4906);
nor NOR4 (N6918, N6911, N2733, N1112, N1465);
xor XOR2 (N6919, N6918, N5893);
nor NOR4 (N6920, N6892, N6764, N6009, N4726);
or OR4 (N6921, N6915, N668, N2054, N3184);
and AND4 (N6922, N6899, N4017, N2176, N1245);
xor XOR2 (N6923, N6914, N6001);
buf BUF1 (N6924, N6919);
not NOT1 (N6925, N6921);
nor NOR4 (N6926, N6923, N1286, N343, N6300);
or OR3 (N6927, N6907, N4710, N6509);
xor XOR2 (N6928, N6906, N1185);
buf BUF1 (N6929, N6922);
and AND4 (N6930, N6917, N5284, N5075, N5058);
xor XOR2 (N6931, N6927, N3551);
nor NOR2 (N6932, N6928, N5220);
or OR3 (N6933, N6930, N3428, N376);
not NOT1 (N6934, N6933);
not NOT1 (N6935, N6929);
not NOT1 (N6936, N6912);
and AND4 (N6937, N6932, N4700, N1376, N5294);
and AND4 (N6938, N6937, N3591, N5444, N2715);
or OR3 (N6939, N6935, N904, N2343);
nor NOR2 (N6940, N6939, N6414);
and AND2 (N6941, N6925, N934);
nand NAND3 (N6942, N6916, N5053, N5358);
not NOT1 (N6943, N6926);
and AND3 (N6944, N6924, N1249, N3887);
nand NAND3 (N6945, N6941, N1999, N1182);
buf BUF1 (N6946, N6940);
not NOT1 (N6947, N6920);
nand NAND2 (N6948, N6944, N5321);
not NOT1 (N6949, N6943);
or OR4 (N6950, N6947, N3055, N766, N3870);
not NOT1 (N6951, N6948);
buf BUF1 (N6952, N6934);
buf BUF1 (N6953, N6951);
nor NOR2 (N6954, N6952, N3045);
nor NOR3 (N6955, N6949, N3521, N2359);
xor XOR2 (N6956, N6942, N542);
and AND2 (N6957, N6950, N3260);
not NOT1 (N6958, N6946);
nor NOR4 (N6959, N6957, N5090, N154, N1609);
nor NOR2 (N6960, N6959, N5160);
nor NOR4 (N6961, N6960, N5485, N6382, N6864);
or OR3 (N6962, N6955, N3131, N636);
nor NOR2 (N6963, N6945, N3006);
nand NAND3 (N6964, N6938, N2315, N635);
nor NOR3 (N6965, N6956, N6543, N1364);
not NOT1 (N6966, N6931);
nand NAND2 (N6967, N6965, N3628);
or OR4 (N6968, N6954, N4222, N5398, N3161);
buf BUF1 (N6969, N6962);
buf BUF1 (N6970, N6967);
and AND3 (N6971, N6964, N2209, N994);
buf BUF1 (N6972, N6953);
nand NAND2 (N6973, N6970, N6906);
nor NOR2 (N6974, N6969, N3736);
nor NOR3 (N6975, N6973, N5409, N1930);
not NOT1 (N6976, N6975);
nor NOR4 (N6977, N6958, N6366, N3463, N4096);
buf BUF1 (N6978, N6976);
and AND3 (N6979, N6974, N1441, N3459);
nand NAND4 (N6980, N6979, N2874, N555, N5886);
or OR2 (N6981, N6936, N5275);
xor XOR2 (N6982, N6971, N1879);
or OR2 (N6983, N6980, N3594);
nor NOR4 (N6984, N6968, N3712, N3945, N6449);
xor XOR2 (N6985, N6983, N3985);
and AND4 (N6986, N6963, N4540, N1412, N4927);
or OR3 (N6987, N6982, N5413, N4136);
or OR4 (N6988, N6987, N6836, N2023, N2003);
xor XOR2 (N6989, N6986, N830);
or OR2 (N6990, N6961, N2145);
xor XOR2 (N6991, N6985, N1081);
nand NAND2 (N6992, N6988, N4040);
buf BUF1 (N6993, N6990);
xor XOR2 (N6994, N6991, N3086);
nand NAND3 (N6995, N6989, N6954, N194);
xor XOR2 (N6996, N6972, N2683);
and AND3 (N6997, N6981, N4305, N2763);
buf BUF1 (N6998, N6977);
not NOT1 (N6999, N6997);
or OR3 (N7000, N6993, N1978, N2078);
nor NOR4 (N7001, N6992, N1475, N2503, N643);
xor XOR2 (N7002, N6996, N2271);
buf BUF1 (N7003, N6994);
nor NOR3 (N7004, N6995, N6636, N2923);
buf BUF1 (N7005, N6998);
xor XOR2 (N7006, N6999, N4120);
nor NOR2 (N7007, N6978, N6741);
nor NOR2 (N7008, N7005, N4503);
nand NAND4 (N7009, N6966, N2751, N3047, N6076);
xor XOR2 (N7010, N7004, N4932);
buf BUF1 (N7011, N7010);
buf BUF1 (N7012, N7001);
buf BUF1 (N7013, N7012);
and AND2 (N7014, N7013, N3147);
xor XOR2 (N7015, N7009, N3458);
nand NAND4 (N7016, N7002, N6428, N1625, N6713);
nor NOR2 (N7017, N6984, N6821);
nor NOR2 (N7018, N7007, N803);
nor NOR3 (N7019, N7006, N4480, N1023);
buf BUF1 (N7020, N7018);
nand NAND2 (N7021, N7016, N1085);
and AND3 (N7022, N7000, N17, N2456);
and AND2 (N7023, N7015, N3351);
or OR4 (N7024, N7003, N2894, N2653, N5089);
nand NAND3 (N7025, N7023, N2615, N3675);
xor XOR2 (N7026, N7021, N5951);
buf BUF1 (N7027, N7020);
and AND3 (N7028, N7011, N4416, N2894);
xor XOR2 (N7029, N7025, N4457);
xor XOR2 (N7030, N7027, N1699);
xor XOR2 (N7031, N7026, N1495);
or OR3 (N7032, N7022, N2217, N5549);
nand NAND3 (N7033, N7028, N2377, N3307);
and AND2 (N7034, N7031, N1587);
and AND4 (N7035, N7019, N778, N3431, N6674);
or OR4 (N7036, N7034, N945, N3586, N6090);
not NOT1 (N7037, N7032);
nor NOR3 (N7038, N7008, N2897, N4579);
xor XOR2 (N7039, N7037, N2959);
nand NAND2 (N7040, N7035, N4084);
or OR4 (N7041, N7033, N2144, N1552, N4590);
or OR3 (N7042, N7030, N5814, N782);
nand NAND2 (N7043, N7029, N5720);
or OR3 (N7044, N7043, N2451, N6115);
not NOT1 (N7045, N7044);
xor XOR2 (N7046, N7024, N1086);
nand NAND4 (N7047, N7017, N5555, N4859, N3421);
nor NOR3 (N7048, N7038, N2567, N5466);
and AND4 (N7049, N7039, N3974, N5699, N2744);
xor XOR2 (N7050, N7047, N6170);
not NOT1 (N7051, N7050);
buf BUF1 (N7052, N7041);
and AND4 (N7053, N7046, N5504, N929, N89);
not NOT1 (N7054, N7053);
or OR4 (N7055, N7054, N6846, N6964, N6514);
nand NAND2 (N7056, N7049, N1321);
and AND2 (N7057, N7056, N4904);
or OR2 (N7058, N7040, N6262);
and AND2 (N7059, N7036, N2645);
and AND3 (N7060, N7055, N4782, N2701);
or OR4 (N7061, N7059, N4993, N3959, N4154);
not NOT1 (N7062, N7042);
and AND2 (N7063, N7060, N4729);
nand NAND2 (N7064, N7045, N811);
not NOT1 (N7065, N7048);
nand NAND4 (N7066, N7057, N6003, N4867, N3297);
nand NAND4 (N7067, N7051, N3988, N3779, N395);
nor NOR2 (N7068, N7063, N676);
nand NAND4 (N7069, N7065, N4668, N1301, N3256);
and AND4 (N7070, N7069, N2500, N3136, N1668);
not NOT1 (N7071, N7052);
nor NOR4 (N7072, N7058, N4299, N2183, N3924);
or OR4 (N7073, N7072, N2939, N4522, N4169);
or OR4 (N7074, N7071, N4292, N3814, N1133);
nand NAND3 (N7075, N7014, N6416, N5674);
or OR3 (N7076, N7064, N1982, N1878);
xor XOR2 (N7077, N7068, N1170);
not NOT1 (N7078, N7066);
buf BUF1 (N7079, N7073);
nand NAND3 (N7080, N7074, N3121, N3138);
xor XOR2 (N7081, N7061, N1515);
nor NOR2 (N7082, N7079, N6305);
nor NOR4 (N7083, N7076, N688, N473, N820);
nand NAND3 (N7084, N7082, N6551, N1702);
nor NOR2 (N7085, N7078, N6362);
or OR4 (N7086, N7085, N1909, N61, N449);
nor NOR2 (N7087, N7086, N5326);
not NOT1 (N7088, N7075);
buf BUF1 (N7089, N7084);
nand NAND3 (N7090, N7081, N5018, N4448);
nand NAND3 (N7091, N7062, N3508, N2525);
buf BUF1 (N7092, N7070);
nor NOR4 (N7093, N7090, N581, N6681, N1264);
and AND4 (N7094, N7083, N3675, N4705, N4625);
buf BUF1 (N7095, N7088);
buf BUF1 (N7096, N7092);
and AND2 (N7097, N7091, N5134);
not NOT1 (N7098, N7096);
or OR3 (N7099, N7097, N1139, N5193);
or OR2 (N7100, N7098, N6235);
nor NOR4 (N7101, N7089, N7080, N1279, N3500);
buf BUF1 (N7102, N5084);
nand NAND3 (N7103, N7100, N2842, N2615);
xor XOR2 (N7104, N7099, N6986);
xor XOR2 (N7105, N7101, N382);
buf BUF1 (N7106, N7102);
not NOT1 (N7107, N7103);
nand NAND4 (N7108, N7107, N6418, N5418, N876);
nor NOR2 (N7109, N7104, N2773);
xor XOR2 (N7110, N7109, N5304);
not NOT1 (N7111, N7087);
and AND3 (N7112, N7077, N5766, N4952);
not NOT1 (N7113, N7095);
nand NAND4 (N7114, N7112, N626, N3732, N218);
nor NOR3 (N7115, N7106, N5680, N4263);
or OR3 (N7116, N7105, N45, N2312);
xor XOR2 (N7117, N7111, N6524);
or OR3 (N7118, N7108, N4451, N6279);
or OR3 (N7119, N7093, N4065, N6209);
xor XOR2 (N7120, N7118, N5125);
buf BUF1 (N7121, N7110);
or OR4 (N7122, N7094, N4967, N2089, N3060);
not NOT1 (N7123, N7119);
not NOT1 (N7124, N7115);
xor XOR2 (N7125, N7117, N5909);
buf BUF1 (N7126, N7124);
and AND3 (N7127, N7123, N5902, N5854);
nand NAND3 (N7128, N7116, N5842, N6622);
or OR4 (N7129, N7067, N5508, N3770, N5813);
or OR2 (N7130, N7114, N5569);
and AND3 (N7131, N7122, N3265, N5892);
or OR3 (N7132, N7128, N5299, N2301);
buf BUF1 (N7133, N7113);
not NOT1 (N7134, N7129);
buf BUF1 (N7135, N7126);
xor XOR2 (N7136, N7130, N5093);
xor XOR2 (N7137, N7134, N1475);
and AND4 (N7138, N7135, N3320, N4692, N5431);
nor NOR4 (N7139, N7125, N4401, N6096, N2437);
not NOT1 (N7140, N7139);
xor XOR2 (N7141, N7132, N1753);
xor XOR2 (N7142, N7133, N710);
buf BUF1 (N7143, N7127);
and AND2 (N7144, N7140, N3292);
or OR3 (N7145, N7120, N5025, N499);
and AND4 (N7146, N7136, N5694, N6726, N4130);
xor XOR2 (N7147, N7131, N5452);
or OR4 (N7148, N7137, N3007, N3449, N1180);
or OR4 (N7149, N7148, N1466, N3879, N5819);
nand NAND3 (N7150, N7149, N4569, N6708);
not NOT1 (N7151, N7138);
or OR3 (N7152, N7121, N135, N2350);
nor NOR3 (N7153, N7152, N665, N96);
and AND2 (N7154, N7146, N2312);
and AND4 (N7155, N7144, N2828, N530, N3934);
xor XOR2 (N7156, N7145, N4769);
nand NAND4 (N7157, N7155, N3770, N5331, N2313);
or OR4 (N7158, N7147, N3724, N6905, N7127);
and AND2 (N7159, N7143, N4487);
not NOT1 (N7160, N7151);
buf BUF1 (N7161, N7153);
nand NAND4 (N7162, N7161, N3293, N6680, N1280);
nor NOR3 (N7163, N7156, N1779, N733);
xor XOR2 (N7164, N7158, N5705);
nor NOR2 (N7165, N7150, N3745);
and AND2 (N7166, N7162, N6817);
xor XOR2 (N7167, N7165, N3633);
buf BUF1 (N7168, N7154);
and AND4 (N7169, N7168, N1742, N3504, N6233);
buf BUF1 (N7170, N7163);
xor XOR2 (N7171, N7164, N612);
buf BUF1 (N7172, N7159);
nand NAND4 (N7173, N7166, N952, N5993, N673);
nor NOR2 (N7174, N7172, N4916);
nor NOR3 (N7175, N7141, N5107, N6613);
xor XOR2 (N7176, N7160, N3985);
or OR2 (N7177, N7170, N1514);
or OR2 (N7178, N7175, N3061);
not NOT1 (N7179, N7173);
nand NAND3 (N7180, N7177, N5909, N6787);
xor XOR2 (N7181, N7174, N4267);
and AND4 (N7182, N7169, N6745, N4659, N2763);
or OR2 (N7183, N7180, N3800);
and AND2 (N7184, N7183, N6638);
and AND4 (N7185, N7142, N6269, N2843, N2932);
buf BUF1 (N7186, N7185);
nand NAND3 (N7187, N7178, N6541, N3732);
xor XOR2 (N7188, N7171, N1950);
and AND3 (N7189, N7179, N1296, N3100);
and AND3 (N7190, N7189, N924, N7054);
buf BUF1 (N7191, N7181);
xor XOR2 (N7192, N7186, N5600);
and AND2 (N7193, N7184, N4736);
nand NAND4 (N7194, N7191, N3778, N2281, N263);
buf BUF1 (N7195, N7176);
nor NOR4 (N7196, N7195, N2770, N2030, N6659);
buf BUF1 (N7197, N7192);
nand NAND3 (N7198, N7188, N1443, N1161);
nor NOR3 (N7199, N7182, N2625, N4083);
and AND4 (N7200, N7194, N1550, N6973, N3709);
or OR4 (N7201, N7193, N5305, N6492, N290);
nand NAND3 (N7202, N7157, N6310, N6636);
buf BUF1 (N7203, N7190);
or OR3 (N7204, N7196, N2512, N5859);
or OR3 (N7205, N7197, N6007, N1837);
xor XOR2 (N7206, N7200, N2312);
nand NAND4 (N7207, N7198, N1982, N6806, N2347);
or OR3 (N7208, N7205, N4136, N2600);
nor NOR2 (N7209, N7206, N5012);
not NOT1 (N7210, N7167);
nor NOR2 (N7211, N7187, N3248);
or OR4 (N7212, N7207, N1207, N5708, N293);
xor XOR2 (N7213, N7203, N5926);
or OR2 (N7214, N7201, N709);
nor NOR3 (N7215, N7214, N1700, N1488);
or OR4 (N7216, N7211, N6682, N777, N3455);
nand NAND4 (N7217, N7212, N6652, N2550, N5672);
nand NAND2 (N7218, N7199, N1571);
and AND4 (N7219, N7217, N692, N1538, N4734);
and AND4 (N7220, N7208, N4530, N1333, N976);
buf BUF1 (N7221, N7218);
not NOT1 (N7222, N7216);
buf BUF1 (N7223, N7220);
nand NAND3 (N7224, N7202, N5291, N2560);
xor XOR2 (N7225, N7223, N2355);
nand NAND3 (N7226, N7209, N2685, N1196);
xor XOR2 (N7227, N7224, N1548);
buf BUF1 (N7228, N7204);
buf BUF1 (N7229, N7227);
or OR4 (N7230, N7221, N1479, N737, N4281);
nor NOR4 (N7231, N7215, N2412, N557, N4630);
nor NOR3 (N7232, N7225, N6308, N6707);
nor NOR2 (N7233, N7222, N5593);
nand NAND4 (N7234, N7233, N6983, N5621, N5300);
buf BUF1 (N7235, N7231);
and AND3 (N7236, N7213, N5532, N913);
nand NAND3 (N7237, N7232, N35, N1909);
nor NOR3 (N7238, N7235, N635, N4236);
xor XOR2 (N7239, N7230, N1010);
not NOT1 (N7240, N7239);
nand NAND4 (N7241, N7237, N1241, N3896, N3252);
or OR3 (N7242, N7219, N5320, N696);
buf BUF1 (N7243, N7242);
nand NAND3 (N7244, N7234, N6294, N2129);
xor XOR2 (N7245, N7229, N2410);
buf BUF1 (N7246, N7238);
buf BUF1 (N7247, N7244);
nand NAND3 (N7248, N7236, N1858, N3392);
not NOT1 (N7249, N7246);
xor XOR2 (N7250, N7228, N7039);
not NOT1 (N7251, N7250);
not NOT1 (N7252, N7249);
and AND3 (N7253, N7210, N2271, N7176);
not NOT1 (N7254, N7251);
buf BUF1 (N7255, N7253);
nand NAND4 (N7256, N7254, N4273, N5294, N6996);
nand NAND3 (N7257, N7241, N3677, N6746);
not NOT1 (N7258, N7255);
buf BUF1 (N7259, N7240);
nor NOR2 (N7260, N7248, N1625);
buf BUF1 (N7261, N7247);
or OR3 (N7262, N7252, N2422, N4771);
nor NOR2 (N7263, N7258, N1502);
buf BUF1 (N7264, N7260);
xor XOR2 (N7265, N7257, N739);
nand NAND4 (N7266, N7245, N2722, N4294, N6597);
nor NOR3 (N7267, N7259, N5783, N2773);
nand NAND3 (N7268, N7264, N5746, N6507);
or OR2 (N7269, N7256, N4890);
and AND4 (N7270, N7267, N6747, N1265, N3513);
xor XOR2 (N7271, N7265, N3050);
not NOT1 (N7272, N7268);
buf BUF1 (N7273, N7226);
nor NOR3 (N7274, N7261, N3895, N3061);
and AND2 (N7275, N7271, N5399);
xor XOR2 (N7276, N7273, N3017);
xor XOR2 (N7277, N7269, N4791);
or OR2 (N7278, N7276, N3334);
nor NOR4 (N7279, N7270, N4890, N1940, N1692);
xor XOR2 (N7280, N7263, N4994);
xor XOR2 (N7281, N7278, N5712);
not NOT1 (N7282, N7272);
not NOT1 (N7283, N7279);
or OR3 (N7284, N7275, N5533, N5186);
or OR3 (N7285, N7243, N5852, N3487);
xor XOR2 (N7286, N7266, N5226);
or OR2 (N7287, N7286, N3839);
not NOT1 (N7288, N7277);
xor XOR2 (N7289, N7282, N582);
nand NAND2 (N7290, N7283, N6594);
or OR2 (N7291, N7287, N1507);
xor XOR2 (N7292, N7284, N716);
nand NAND2 (N7293, N7281, N6373);
xor XOR2 (N7294, N7289, N2842);
or OR2 (N7295, N7262, N5133);
not NOT1 (N7296, N7274);
nand NAND3 (N7297, N7296, N6614, N3566);
and AND3 (N7298, N7290, N4034, N2700);
and AND4 (N7299, N7285, N3817, N4281, N5802);
or OR4 (N7300, N7299, N715, N6961, N657);
nand NAND2 (N7301, N7292, N6408);
not NOT1 (N7302, N7291);
buf BUF1 (N7303, N7297);
buf BUF1 (N7304, N7300);
nor NOR4 (N7305, N7298, N4196, N6973, N6321);
not NOT1 (N7306, N7303);
and AND4 (N7307, N7280, N740, N961, N4742);
and AND2 (N7308, N7294, N5628);
buf BUF1 (N7309, N7295);
buf BUF1 (N7310, N7309);
buf BUF1 (N7311, N7308);
and AND2 (N7312, N7311, N1049);
or OR2 (N7313, N7302, N4496);
nor NOR2 (N7314, N7312, N3036);
not NOT1 (N7315, N7293);
nand NAND3 (N7316, N7288, N1489, N7095);
nand NAND2 (N7317, N7315, N2788);
buf BUF1 (N7318, N7313);
nand NAND4 (N7319, N7314, N6657, N2750, N5087);
not NOT1 (N7320, N7301);
nand NAND3 (N7321, N7310, N6525, N2922);
or OR2 (N7322, N7305, N5228);
nand NAND4 (N7323, N7304, N958, N87, N1009);
xor XOR2 (N7324, N7318, N7104);
or OR2 (N7325, N7317, N1828);
not NOT1 (N7326, N7307);
xor XOR2 (N7327, N7326, N4695);
xor XOR2 (N7328, N7327, N1676);
or OR2 (N7329, N7325, N3431);
buf BUF1 (N7330, N7322);
or OR2 (N7331, N7324, N5469);
nor NOR2 (N7332, N7316, N1803);
buf BUF1 (N7333, N7328);
or OR2 (N7334, N7321, N5745);
not NOT1 (N7335, N7330);
nand NAND4 (N7336, N7319, N6246, N765, N2390);
nand NAND3 (N7337, N7306, N6004, N6066);
nand NAND4 (N7338, N7331, N3809, N6957, N2401);
not NOT1 (N7339, N7320);
or OR4 (N7340, N7335, N89, N6497, N3202);
nand NAND4 (N7341, N7340, N3030, N779, N4456);
not NOT1 (N7342, N7329);
nand NAND3 (N7343, N7339, N5554, N5069);
xor XOR2 (N7344, N7342, N7082);
nand NAND3 (N7345, N7344, N6746, N1872);
buf BUF1 (N7346, N7333);
nand NAND3 (N7347, N7332, N696, N1546);
or OR4 (N7348, N7346, N3165, N686, N1728);
nand NAND3 (N7349, N7347, N1580, N3090);
xor XOR2 (N7350, N7336, N4140);
xor XOR2 (N7351, N7349, N2748);
and AND2 (N7352, N7323, N5142);
or OR3 (N7353, N7351, N5112, N3172);
and AND3 (N7354, N7352, N815, N3066);
buf BUF1 (N7355, N7353);
buf BUF1 (N7356, N7341);
buf BUF1 (N7357, N7348);
nor NOR3 (N7358, N7337, N2240, N4648);
buf BUF1 (N7359, N7338);
nor NOR4 (N7360, N7355, N715, N3722, N5174);
xor XOR2 (N7361, N7334, N3553);
nor NOR4 (N7362, N7345, N3608, N344, N4316);
nand NAND2 (N7363, N7356, N2449);
or OR4 (N7364, N7363, N3153, N3806, N6588);
nand NAND4 (N7365, N7357, N2067, N81, N3590);
xor XOR2 (N7366, N7361, N4336);
nand NAND2 (N7367, N7350, N6501);
buf BUF1 (N7368, N7360);
buf BUF1 (N7369, N7367);
nor NOR4 (N7370, N7364, N2424, N5815, N3625);
and AND3 (N7371, N7358, N6685, N4794);
and AND4 (N7372, N7368, N175, N3584, N3627);
not NOT1 (N7373, N7366);
nand NAND3 (N7374, N7370, N3999, N6281);
buf BUF1 (N7375, N7372);
or OR4 (N7376, N7359, N2606, N6896, N298);
nor NOR4 (N7377, N7362, N37, N2694, N3569);
and AND2 (N7378, N7371, N2117);
buf BUF1 (N7379, N7369);
and AND3 (N7380, N7343, N6850, N1720);
buf BUF1 (N7381, N7380);
not NOT1 (N7382, N7381);
nor NOR4 (N7383, N7376, N5149, N2164, N1267);
not NOT1 (N7384, N7373);
or OR4 (N7385, N7384, N2878, N5911, N1594);
or OR3 (N7386, N7382, N1040, N3021);
buf BUF1 (N7387, N7379);
nand NAND3 (N7388, N7365, N7006, N3111);
and AND4 (N7389, N7354, N4880, N6227, N5529);
nor NOR2 (N7390, N7385, N6428);
not NOT1 (N7391, N7386);
buf BUF1 (N7392, N7383);
nand NAND3 (N7393, N7389, N3222, N3535);
not NOT1 (N7394, N7388);
or OR4 (N7395, N7392, N2157, N5956, N3403);
xor XOR2 (N7396, N7390, N3849);
or OR2 (N7397, N7387, N5142);
nand NAND2 (N7398, N7393, N5271);
nor NOR3 (N7399, N7391, N1198, N6871);
or OR4 (N7400, N7398, N4570, N3804, N5412);
buf BUF1 (N7401, N7397);
or OR2 (N7402, N7401, N996);
not NOT1 (N7403, N7378);
nor NOR3 (N7404, N7402, N4321, N3874);
xor XOR2 (N7405, N7400, N4399);
nand NAND4 (N7406, N7396, N5910, N3478, N4172);
nor NOR3 (N7407, N7403, N6239, N2536);
or OR2 (N7408, N7394, N6277);
nand NAND3 (N7409, N7404, N1019, N1545);
nor NOR3 (N7410, N7406, N3472, N2080);
and AND2 (N7411, N7405, N3232);
or OR2 (N7412, N7407, N3648);
nor NOR4 (N7413, N7395, N5903, N3019, N4361);
or OR3 (N7414, N7408, N2145, N6152);
and AND4 (N7415, N7377, N5794, N1700, N1511);
not NOT1 (N7416, N7409);
nand NAND2 (N7417, N7415, N1582);
buf BUF1 (N7418, N7410);
and AND4 (N7419, N7374, N1380, N6687, N5998);
buf BUF1 (N7420, N7419);
and AND3 (N7421, N7411, N468, N2753);
nand NAND2 (N7422, N7412, N6838);
not NOT1 (N7423, N7414);
xor XOR2 (N7424, N7418, N3084);
nor NOR3 (N7425, N7423, N2441, N978);
buf BUF1 (N7426, N7422);
not NOT1 (N7427, N7375);
nand NAND3 (N7428, N7421, N2624, N3300);
and AND4 (N7429, N7413, N3922, N4417, N6167);
not NOT1 (N7430, N7426);
nand NAND3 (N7431, N7425, N7312, N6339);
and AND2 (N7432, N7428, N6443);
buf BUF1 (N7433, N7427);
nor NOR4 (N7434, N7399, N963, N2010, N1468);
not NOT1 (N7435, N7420);
xor XOR2 (N7436, N7430, N4524);
nand NAND3 (N7437, N7417, N6160, N1654);
buf BUF1 (N7438, N7431);
not NOT1 (N7439, N7433);
xor XOR2 (N7440, N7424, N7212);
or OR4 (N7441, N7432, N2260, N1791, N2242);
nor NOR4 (N7442, N7441, N289, N5152, N6305);
or OR4 (N7443, N7434, N622, N1481, N480);
nand NAND2 (N7444, N7440, N2621);
nor NOR3 (N7445, N7437, N5190, N2457);
and AND4 (N7446, N7416, N3159, N269, N5746);
buf BUF1 (N7447, N7435);
or OR4 (N7448, N7429, N1782, N6357, N3442);
buf BUF1 (N7449, N7443);
nand NAND4 (N7450, N7436, N354, N869, N2487);
or OR3 (N7451, N7448, N74, N7122);
not NOT1 (N7452, N7449);
or OR4 (N7453, N7444, N5937, N6344, N7385);
xor XOR2 (N7454, N7445, N5923);
nand NAND2 (N7455, N7453, N4763);
or OR2 (N7456, N7451, N5642);
nor NOR2 (N7457, N7456, N5002);
or OR3 (N7458, N7452, N4354, N1373);
nor NOR2 (N7459, N7446, N2195);
and AND2 (N7460, N7458, N5416);
buf BUF1 (N7461, N7460);
or OR4 (N7462, N7461, N226, N5661, N4524);
and AND2 (N7463, N7442, N4046);
not NOT1 (N7464, N7462);
nand NAND2 (N7465, N7447, N3237);
nand NAND3 (N7466, N7457, N938, N4858);
xor XOR2 (N7467, N7439, N1123);
nor NOR3 (N7468, N7455, N5404, N2756);
xor XOR2 (N7469, N7465, N6346);
nor NOR2 (N7470, N7464, N6964);
nand NAND2 (N7471, N7467, N2229);
nor NOR2 (N7472, N7463, N6256);
nand NAND3 (N7473, N7470, N1287, N6674);
nor NOR3 (N7474, N7466, N391, N3068);
buf BUF1 (N7475, N7469);
xor XOR2 (N7476, N7468, N5229);
or OR3 (N7477, N7474, N3679, N6715);
nor NOR4 (N7478, N7477, N6394, N1974, N1206);
nor NOR4 (N7479, N7473, N3058, N3932, N4965);
xor XOR2 (N7480, N7472, N4347);
not NOT1 (N7481, N7471);
xor XOR2 (N7482, N7479, N1880);
nor NOR2 (N7483, N7478, N487);
nor NOR4 (N7484, N7481, N1678, N3628, N2877);
nor NOR4 (N7485, N7438, N7233, N2519, N2195);
buf BUF1 (N7486, N7480);
and AND2 (N7487, N7484, N753);
nand NAND4 (N7488, N7459, N3402, N2643, N6504);
nor NOR4 (N7489, N7482, N7097, N1872, N770);
buf BUF1 (N7490, N7475);
nand NAND3 (N7491, N7487, N4434, N3619);
or OR2 (N7492, N7485, N5777);
nand NAND3 (N7493, N7492, N6962, N6870);
xor XOR2 (N7494, N7493, N6694);
not NOT1 (N7495, N7490);
or OR4 (N7496, N7488, N226, N1361, N1027);
xor XOR2 (N7497, N7494, N553);
nor NOR4 (N7498, N7497, N4780, N3256, N3977);
xor XOR2 (N7499, N7496, N1071);
nand NAND3 (N7500, N7450, N2082, N7056);
nor NOR4 (N7501, N7491, N4969, N7424, N6655);
and AND4 (N7502, N7500, N6453, N1224, N6511);
and AND3 (N7503, N7454, N7494, N3001);
xor XOR2 (N7504, N7486, N5394);
nor NOR2 (N7505, N7495, N1061);
and AND2 (N7506, N7489, N4371);
nand NAND4 (N7507, N7499, N3359, N3946, N6131);
nor NOR4 (N7508, N7476, N228, N6868, N6503);
and AND2 (N7509, N7503, N788);
or OR4 (N7510, N7506, N1950, N6380, N1775);
and AND4 (N7511, N7507, N5119, N1143, N7178);
nor NOR2 (N7512, N7483, N4597);
nand NAND4 (N7513, N7511, N2788, N6746, N4202);
nor NOR3 (N7514, N7509, N92, N1775);
not NOT1 (N7515, N7508);
and AND4 (N7516, N7505, N5307, N4604, N5616);
nor NOR2 (N7517, N7502, N3235);
nor NOR4 (N7518, N7501, N3852, N7138, N2628);
nor NOR2 (N7519, N7498, N3288);
buf BUF1 (N7520, N7510);
nand NAND3 (N7521, N7513, N2668, N3409);
nand NAND2 (N7522, N7504, N4296);
nand NAND3 (N7523, N7522, N3805, N3510);
not NOT1 (N7524, N7520);
nor NOR4 (N7525, N7512, N4570, N2522, N643);
and AND3 (N7526, N7519, N2700, N461);
nor NOR2 (N7527, N7521, N5207);
nand NAND3 (N7528, N7517, N5202, N7482);
or OR2 (N7529, N7525, N11);
buf BUF1 (N7530, N7528);
nor NOR4 (N7531, N7524, N5778, N3104, N3516);
or OR4 (N7532, N7523, N49, N3073, N4493);
not NOT1 (N7533, N7518);
xor XOR2 (N7534, N7526, N4569);
not NOT1 (N7535, N7516);
nor NOR4 (N7536, N7532, N3634, N7030, N3699);
nand NAND3 (N7537, N7514, N6087, N2898);
xor XOR2 (N7538, N7534, N3034);
buf BUF1 (N7539, N7535);
xor XOR2 (N7540, N7538, N1817);
xor XOR2 (N7541, N7536, N7185);
or OR4 (N7542, N7533, N6819, N3954, N1780);
not NOT1 (N7543, N7529);
nor NOR3 (N7544, N7542, N3506, N1029);
nor NOR3 (N7545, N7541, N5519, N1728);
nor NOR4 (N7546, N7544, N1208, N1021, N1126);
not NOT1 (N7547, N7545);
nor NOR4 (N7548, N7539, N1752, N5134, N6577);
and AND3 (N7549, N7546, N5688, N5518);
not NOT1 (N7550, N7537);
and AND3 (N7551, N7540, N1747, N2085);
or OR3 (N7552, N7530, N2485, N3944);
nor NOR2 (N7553, N7515, N4426);
not NOT1 (N7554, N7531);
buf BUF1 (N7555, N7547);
nor NOR3 (N7556, N7527, N2621, N4083);
xor XOR2 (N7557, N7552, N5828);
buf BUF1 (N7558, N7554);
xor XOR2 (N7559, N7557, N2970);
buf BUF1 (N7560, N7553);
buf BUF1 (N7561, N7548);
or OR3 (N7562, N7543, N1972, N7315);
and AND2 (N7563, N7560, N1654);
nor NOR2 (N7564, N7561, N735);
nand NAND4 (N7565, N7551, N6316, N6578, N5727);
and AND4 (N7566, N7549, N3788, N4929, N2238);
buf BUF1 (N7567, N7563);
xor XOR2 (N7568, N7555, N186);
xor XOR2 (N7569, N7568, N4723);
nand NAND4 (N7570, N7556, N2716, N7188, N7073);
or OR3 (N7571, N7564, N4779, N5685);
nand NAND2 (N7572, N7571, N1101);
and AND3 (N7573, N7562, N232, N7255);
nand NAND4 (N7574, N7570, N6793, N1991, N3217);
xor XOR2 (N7575, N7573, N2879);
nor NOR4 (N7576, N7565, N2572, N6604, N528);
buf BUF1 (N7577, N7574);
xor XOR2 (N7578, N7567, N2598);
nor NOR3 (N7579, N7550, N6793, N1869);
buf BUF1 (N7580, N7569);
xor XOR2 (N7581, N7580, N950);
and AND4 (N7582, N7572, N1716, N1687, N3049);
xor XOR2 (N7583, N7578, N6654);
nand NAND4 (N7584, N7576, N5563, N661, N2249);
nand NAND4 (N7585, N7584, N4887, N3924, N5557);
nand NAND2 (N7586, N7579, N2561);
nand NAND3 (N7587, N7586, N2380, N6523);
not NOT1 (N7588, N7558);
xor XOR2 (N7589, N7577, N2987);
nand NAND3 (N7590, N7585, N1826, N7119);
xor XOR2 (N7591, N7575, N5480);
or OR4 (N7592, N7588, N3735, N6834, N4566);
not NOT1 (N7593, N7590);
and AND2 (N7594, N7581, N4635);
not NOT1 (N7595, N7594);
nand NAND4 (N7596, N7566, N7267, N6679, N1062);
xor XOR2 (N7597, N7596, N779);
or OR3 (N7598, N7593, N4926, N4614);
buf BUF1 (N7599, N7589);
nor NOR3 (N7600, N7592, N913, N6913);
nor NOR2 (N7601, N7591, N3658);
xor XOR2 (N7602, N7559, N6772);
and AND3 (N7603, N7583, N3995, N1095);
xor XOR2 (N7604, N7601, N5800);
xor XOR2 (N7605, N7604, N5555);
or OR4 (N7606, N7602, N7333, N6401, N5275);
xor XOR2 (N7607, N7606, N2963);
or OR2 (N7608, N7597, N6360);
xor XOR2 (N7609, N7607, N511);
nor NOR3 (N7610, N7603, N937, N7411);
xor XOR2 (N7611, N7608, N1189);
or OR3 (N7612, N7599, N5838, N4193);
xor XOR2 (N7613, N7612, N5162);
or OR2 (N7614, N7613, N7516);
not NOT1 (N7615, N7582);
not NOT1 (N7616, N7587);
or OR3 (N7617, N7609, N1277, N5592);
nand NAND4 (N7618, N7598, N6140, N4137, N6820);
nor NOR3 (N7619, N7616, N5191, N4887);
xor XOR2 (N7620, N7605, N3148);
xor XOR2 (N7621, N7618, N658);
not NOT1 (N7622, N7600);
nand NAND4 (N7623, N7611, N7138, N348, N7215);
buf BUF1 (N7624, N7619);
nand NAND2 (N7625, N7621, N6253);
buf BUF1 (N7626, N7625);
or OR4 (N7627, N7610, N7054, N2122, N707);
and AND4 (N7628, N7615, N1607, N4506, N6596);
xor XOR2 (N7629, N7623, N281);
xor XOR2 (N7630, N7628, N2904);
and AND3 (N7631, N7617, N609, N1637);
xor XOR2 (N7632, N7631, N5869);
buf BUF1 (N7633, N7632);
not NOT1 (N7634, N7595);
and AND2 (N7635, N7614, N3964);
and AND2 (N7636, N7622, N1989);
buf BUF1 (N7637, N7629);
not NOT1 (N7638, N7636);
nand NAND4 (N7639, N7630, N365, N1029, N6231);
nor NOR3 (N7640, N7637, N6878, N5742);
buf BUF1 (N7641, N7624);
buf BUF1 (N7642, N7627);
not NOT1 (N7643, N7620);
xor XOR2 (N7644, N7626, N3892);
and AND4 (N7645, N7643, N6910, N7183, N1109);
nor NOR3 (N7646, N7635, N7640, N4647);
nor NOR4 (N7647, N3299, N6860, N5290, N7612);
or OR2 (N7648, N7634, N4055);
not NOT1 (N7649, N7648);
nor NOR2 (N7650, N7644, N2993);
buf BUF1 (N7651, N7639);
nor NOR3 (N7652, N7642, N5829, N4863);
and AND3 (N7653, N7633, N5622, N2076);
nor NOR4 (N7654, N7638, N6335, N1683, N4057);
nor NOR3 (N7655, N7650, N542, N6987);
nand NAND4 (N7656, N7653, N2082, N5821, N5074);
xor XOR2 (N7657, N7651, N5098);
or OR3 (N7658, N7656, N7058, N6237);
xor XOR2 (N7659, N7645, N5724);
buf BUF1 (N7660, N7646);
nand NAND4 (N7661, N7654, N2181, N4306, N2152);
and AND4 (N7662, N7652, N6198, N2188, N5375);
nand NAND2 (N7663, N7647, N4315);
nor NOR4 (N7664, N7659, N7447, N520, N2165);
xor XOR2 (N7665, N7641, N6601);
buf BUF1 (N7666, N7657);
xor XOR2 (N7667, N7666, N5552);
not NOT1 (N7668, N7658);
not NOT1 (N7669, N7665);
xor XOR2 (N7670, N7649, N4594);
buf BUF1 (N7671, N7668);
buf BUF1 (N7672, N7670);
xor XOR2 (N7673, N7663, N4799);
buf BUF1 (N7674, N7655);
buf BUF1 (N7675, N7660);
xor XOR2 (N7676, N7672, N2921);
nand NAND4 (N7677, N7667, N2469, N3043, N81);
not NOT1 (N7678, N7662);
not NOT1 (N7679, N7675);
buf BUF1 (N7680, N7679);
nor NOR2 (N7681, N7677, N5927);
buf BUF1 (N7682, N7681);
xor XOR2 (N7683, N7676, N3916);
buf BUF1 (N7684, N7673);
not NOT1 (N7685, N7684);
xor XOR2 (N7686, N7678, N1741);
nor NOR2 (N7687, N7661, N1402);
buf BUF1 (N7688, N7669);
or OR3 (N7689, N7682, N5623, N7515);
and AND2 (N7690, N7685, N4349);
nor NOR3 (N7691, N7671, N3271, N2035);
not NOT1 (N7692, N7686);
nand NAND4 (N7693, N7692, N5675, N7636, N2697);
nor NOR3 (N7694, N7690, N728, N6371);
or OR2 (N7695, N7680, N6983);
nor NOR2 (N7696, N7693, N247);
buf BUF1 (N7697, N7674);
xor XOR2 (N7698, N7696, N2235);
xor XOR2 (N7699, N7698, N4865);
nand NAND4 (N7700, N7687, N1733, N6964, N2301);
not NOT1 (N7701, N7694);
xor XOR2 (N7702, N7699, N348);
buf BUF1 (N7703, N7683);
nor NOR4 (N7704, N7689, N5346, N5400, N5984);
nor NOR3 (N7705, N7697, N3433, N7497);
and AND2 (N7706, N7701, N4804);
xor XOR2 (N7707, N7703, N5480);
nand NAND4 (N7708, N7695, N6536, N641, N512);
not NOT1 (N7709, N7664);
nand NAND3 (N7710, N7691, N2008, N823);
nor NOR3 (N7711, N7702, N3731, N2045);
or OR4 (N7712, N7705, N2952, N3410, N1174);
buf BUF1 (N7713, N7707);
and AND3 (N7714, N7700, N4616, N1369);
xor XOR2 (N7715, N7714, N1950);
nand NAND3 (N7716, N7688, N6961, N6003);
nor NOR3 (N7717, N7709, N3172, N923);
and AND2 (N7718, N7706, N2429);
and AND2 (N7719, N7716, N5780);
nor NOR2 (N7720, N7704, N1017);
nand NAND3 (N7721, N7715, N5023, N6744);
nor NOR2 (N7722, N7720, N6459);
or OR2 (N7723, N7722, N2867);
xor XOR2 (N7724, N7723, N2155);
buf BUF1 (N7725, N7710);
and AND4 (N7726, N7718, N3409, N7549, N3037);
nand NAND4 (N7727, N7724, N517, N1840, N5004);
xor XOR2 (N7728, N7726, N2261);
nor NOR2 (N7729, N7725, N4349);
xor XOR2 (N7730, N7729, N3151);
and AND2 (N7731, N7728, N2533);
buf BUF1 (N7732, N7717);
not NOT1 (N7733, N7719);
not NOT1 (N7734, N7712);
nor NOR4 (N7735, N7727, N7706, N7416, N5632);
xor XOR2 (N7736, N7721, N1727);
xor XOR2 (N7737, N7733, N6613);
xor XOR2 (N7738, N7711, N4182);
buf BUF1 (N7739, N7713);
nor NOR3 (N7740, N7732, N7247, N1677);
nor NOR2 (N7741, N7738, N7683);
nand NAND2 (N7742, N7737, N5831);
or OR2 (N7743, N7739, N4515);
xor XOR2 (N7744, N7731, N6524);
and AND3 (N7745, N7740, N4005, N3950);
not NOT1 (N7746, N7743);
nand NAND2 (N7747, N7744, N3056);
or OR4 (N7748, N7745, N814, N4842, N226);
and AND3 (N7749, N7741, N3948, N569);
buf BUF1 (N7750, N7734);
xor XOR2 (N7751, N7736, N7593);
and AND2 (N7752, N7730, N3109);
nand NAND3 (N7753, N7751, N5857, N4583);
xor XOR2 (N7754, N7750, N3918);
buf BUF1 (N7755, N7708);
nor NOR2 (N7756, N7754, N341);
nor NOR3 (N7757, N7752, N1379, N5621);
nor NOR3 (N7758, N7742, N5963, N6609);
buf BUF1 (N7759, N7753);
or OR4 (N7760, N7758, N1737, N3371, N5118);
not NOT1 (N7761, N7757);
nand NAND2 (N7762, N7759, N5200);
nand NAND2 (N7763, N7762, N912);
not NOT1 (N7764, N7761);
nand NAND2 (N7765, N7746, N6071);
and AND2 (N7766, N7755, N5837);
and AND2 (N7767, N7760, N7116);
nor NOR4 (N7768, N7748, N7553, N6006, N7432);
xor XOR2 (N7769, N7764, N756);
xor XOR2 (N7770, N7767, N6666);
nand NAND4 (N7771, N7765, N1213, N5217, N7272);
nor NOR4 (N7772, N7749, N3669, N7199, N368);
xor XOR2 (N7773, N7763, N5169);
and AND4 (N7774, N7768, N942, N7273, N1109);
and AND3 (N7775, N7773, N961, N7504);
or OR3 (N7776, N7747, N7676, N1180);
not NOT1 (N7777, N7776);
xor XOR2 (N7778, N7766, N7744);
nand NAND3 (N7779, N7774, N6595, N5846);
nand NAND3 (N7780, N7770, N6589, N6097);
buf BUF1 (N7781, N7777);
not NOT1 (N7782, N7775);
not NOT1 (N7783, N7779);
nand NAND2 (N7784, N7756, N4090);
nand NAND3 (N7785, N7778, N3989, N4808);
not NOT1 (N7786, N7780);
xor XOR2 (N7787, N7785, N3829);
buf BUF1 (N7788, N7787);
nor NOR2 (N7789, N7772, N347);
nand NAND3 (N7790, N7786, N331, N7068);
or OR3 (N7791, N7735, N5412, N7390);
and AND3 (N7792, N7790, N2478, N5376);
nor NOR3 (N7793, N7792, N4442, N7481);
buf BUF1 (N7794, N7791);
xor XOR2 (N7795, N7784, N2558);
xor XOR2 (N7796, N7782, N2608);
buf BUF1 (N7797, N7796);
not NOT1 (N7798, N7771);
or OR4 (N7799, N7783, N6922, N2966, N7227);
nand NAND3 (N7800, N7781, N3319, N4708);
nor NOR3 (N7801, N7799, N3775, N3565);
not NOT1 (N7802, N7769);
and AND3 (N7803, N7801, N5628, N7152);
or OR4 (N7804, N7797, N5239, N6217, N6413);
and AND3 (N7805, N7798, N7359, N6902);
xor XOR2 (N7806, N7789, N7597);
nand NAND2 (N7807, N7803, N784);
not NOT1 (N7808, N7800);
not NOT1 (N7809, N7793);
not NOT1 (N7810, N7805);
or OR2 (N7811, N7809, N2878);
buf BUF1 (N7812, N7788);
not NOT1 (N7813, N7794);
not NOT1 (N7814, N7807);
and AND3 (N7815, N7811, N4153, N3621);
xor XOR2 (N7816, N7810, N3752);
nand NAND2 (N7817, N7816, N5631);
buf BUF1 (N7818, N7817);
or OR3 (N7819, N7808, N3405, N4017);
or OR3 (N7820, N7802, N6059, N5972);
nor NOR3 (N7821, N7820, N4174, N2664);
nand NAND4 (N7822, N7804, N7070, N3773, N4715);
and AND3 (N7823, N7815, N4267, N5714);
nand NAND4 (N7824, N7806, N979, N5541, N2676);
buf BUF1 (N7825, N7818);
nor NOR4 (N7826, N7795, N5840, N897, N7441);
buf BUF1 (N7827, N7821);
not NOT1 (N7828, N7813);
nand NAND2 (N7829, N7814, N4278);
not NOT1 (N7830, N7826);
nand NAND2 (N7831, N7823, N7072);
nand NAND3 (N7832, N7830, N6047, N4716);
xor XOR2 (N7833, N7831, N6913);
buf BUF1 (N7834, N7828);
xor XOR2 (N7835, N7822, N980);
buf BUF1 (N7836, N7825);
xor XOR2 (N7837, N7834, N2399);
not NOT1 (N7838, N7832);
nand NAND3 (N7839, N7835, N5889, N691);
nor NOR3 (N7840, N7812, N6202, N932);
nor NOR4 (N7841, N7840, N6870, N5282, N2395);
xor XOR2 (N7842, N7836, N5893);
nand NAND2 (N7843, N7838, N413);
xor XOR2 (N7844, N7837, N5382);
nand NAND3 (N7845, N7824, N2707, N7830);
or OR4 (N7846, N7843, N1414, N7451, N2793);
or OR3 (N7847, N7845, N7212, N3086);
nor NOR4 (N7848, N7844, N1495, N4156, N2251);
and AND3 (N7849, N7842, N1643, N1313);
and AND3 (N7850, N7827, N3685, N6841);
nand NAND4 (N7851, N7839, N3091, N1646, N5146);
and AND3 (N7852, N7848, N6978, N760);
nand NAND3 (N7853, N7849, N6388, N1771);
or OR3 (N7854, N7853, N3389, N3270);
nand NAND4 (N7855, N7841, N7829, N2792, N5501);
buf BUF1 (N7856, N2403);
buf BUF1 (N7857, N7851);
nand NAND2 (N7858, N7857, N874);
xor XOR2 (N7859, N7819, N5834);
and AND3 (N7860, N7833, N5045, N3707);
and AND3 (N7861, N7852, N2289, N4136);
nor NOR4 (N7862, N7860, N6498, N3845, N825);
and AND3 (N7863, N7858, N1829, N983);
nand NAND2 (N7864, N7859, N2715);
and AND2 (N7865, N7864, N2721);
buf BUF1 (N7866, N7847);
not NOT1 (N7867, N7862);
nand NAND4 (N7868, N7861, N1966, N810, N7028);
nor NOR4 (N7869, N7846, N2498, N602, N630);
not NOT1 (N7870, N7866);
not NOT1 (N7871, N7856);
not NOT1 (N7872, N7865);
nand NAND3 (N7873, N7863, N7672, N1264);
not NOT1 (N7874, N7854);
not NOT1 (N7875, N7872);
or OR3 (N7876, N7855, N1995, N7562);
nand NAND3 (N7877, N7850, N427, N7100);
buf BUF1 (N7878, N7871);
or OR2 (N7879, N7874, N40);
xor XOR2 (N7880, N7868, N4882);
buf BUF1 (N7881, N7878);
xor XOR2 (N7882, N7875, N7463);
nor NOR4 (N7883, N7880, N50, N3104, N2381);
nand NAND2 (N7884, N7876, N3458);
nor NOR4 (N7885, N7873, N2089, N7043, N6065);
xor XOR2 (N7886, N7884, N6486);
nand NAND3 (N7887, N7886, N3034, N2947);
nand NAND4 (N7888, N7885, N1652, N1514, N1511);
nor NOR3 (N7889, N7870, N3213, N227);
nand NAND3 (N7890, N7882, N7106, N1320);
or OR3 (N7891, N7881, N1304, N822);
xor XOR2 (N7892, N7888, N2943);
or OR4 (N7893, N7889, N891, N4825, N1172);
or OR2 (N7894, N7877, N2892);
buf BUF1 (N7895, N7869);
xor XOR2 (N7896, N7891, N2392);
and AND4 (N7897, N7887, N3389, N3018, N6266);
not NOT1 (N7898, N7897);
nor NOR4 (N7899, N7883, N3993, N1056, N534);
buf BUF1 (N7900, N7867);
nor NOR3 (N7901, N7899, N168, N762);
xor XOR2 (N7902, N7890, N3831);
not NOT1 (N7903, N7901);
not NOT1 (N7904, N7903);
xor XOR2 (N7905, N7894, N2070);
xor XOR2 (N7906, N7905, N326);
nand NAND2 (N7907, N7879, N2935);
xor XOR2 (N7908, N7902, N575);
xor XOR2 (N7909, N7900, N2438);
or OR2 (N7910, N7907, N1342);
buf BUF1 (N7911, N7910);
nand NAND2 (N7912, N7896, N6876);
nand NAND4 (N7913, N7895, N4043, N7621, N7380);
buf BUF1 (N7914, N7893);
or OR3 (N7915, N7906, N5400, N7783);
nor NOR3 (N7916, N7914, N5716, N1252);
nand NAND4 (N7917, N7915, N390, N7878, N4300);
nor NOR3 (N7918, N7917, N1018, N6002);
nand NAND4 (N7919, N7898, N3757, N3663, N954);
and AND2 (N7920, N7911, N1945);
or OR3 (N7921, N7904, N6609, N541);
and AND4 (N7922, N7908, N6503, N3822, N1298);
not NOT1 (N7923, N7916);
not NOT1 (N7924, N7923);
nand NAND3 (N7925, N7921, N1371, N4016);
nand NAND3 (N7926, N7892, N7338, N71);
not NOT1 (N7927, N7912);
or OR2 (N7928, N7925, N1980);
or OR3 (N7929, N7927, N4259, N6645);
nor NOR4 (N7930, N7928, N6363, N6477, N7622);
and AND3 (N7931, N7926, N7672, N1965);
and AND4 (N7932, N7913, N3721, N6908, N5070);
xor XOR2 (N7933, N7931, N4493);
nor NOR4 (N7934, N7909, N6220, N2589, N1745);
buf BUF1 (N7935, N7929);
nor NOR2 (N7936, N7935, N1362);
buf BUF1 (N7937, N7934);
and AND4 (N7938, N7933, N6092, N4223, N1290);
not NOT1 (N7939, N7920);
buf BUF1 (N7940, N7938);
nand NAND2 (N7941, N7939, N6758);
xor XOR2 (N7942, N7941, N880);
not NOT1 (N7943, N7922);
not NOT1 (N7944, N7932);
or OR3 (N7945, N7943, N3509, N478);
nor NOR4 (N7946, N7944, N4349, N3304, N1443);
nand NAND4 (N7947, N7924, N2954, N5239, N6514);
not NOT1 (N7948, N7937);
and AND4 (N7949, N7919, N2375, N3123, N3071);
or OR2 (N7950, N7945, N1902);
or OR3 (N7951, N7918, N7733, N3719);
nor NOR4 (N7952, N7930, N899, N3909, N2062);
nand NAND4 (N7953, N7948, N7013, N7095, N6707);
nand NAND2 (N7954, N7940, N20);
nand NAND3 (N7955, N7950, N7901, N5315);
or OR4 (N7956, N7949, N4260, N1576, N4706);
nor NOR2 (N7957, N7946, N1767);
and AND4 (N7958, N7956, N5410, N2624, N7932);
and AND2 (N7959, N7951, N984);
not NOT1 (N7960, N7952);
not NOT1 (N7961, N7955);
nand NAND4 (N7962, N7942, N1694, N5563, N2159);
nor NOR3 (N7963, N7954, N5071, N4996);
buf BUF1 (N7964, N7960);
not NOT1 (N7965, N7962);
buf BUF1 (N7966, N7963);
not NOT1 (N7967, N7947);
and AND3 (N7968, N7936, N5128, N6444);
not NOT1 (N7969, N7957);
xor XOR2 (N7970, N7969, N7908);
nand NAND2 (N7971, N7970, N38);
nor NOR3 (N7972, N7971, N4097, N4318);
xor XOR2 (N7973, N7972, N7903);
nand NAND2 (N7974, N7964, N7630);
not NOT1 (N7975, N7966);
nor NOR3 (N7976, N7965, N6449, N23);
nor NOR2 (N7977, N7959, N6183);
nor NOR4 (N7978, N7968, N4682, N3051, N1659);
nand NAND2 (N7979, N7958, N1982);
buf BUF1 (N7980, N7977);
and AND2 (N7981, N7979, N2547);
xor XOR2 (N7982, N7973, N7563);
xor XOR2 (N7983, N7975, N6472);
xor XOR2 (N7984, N7982, N6130);
nand NAND3 (N7985, N7976, N4690, N4947);
or OR2 (N7986, N7978, N5482);
buf BUF1 (N7987, N7984);
or OR2 (N7988, N7967, N3060);
buf BUF1 (N7989, N7980);
not NOT1 (N7990, N7985);
not NOT1 (N7991, N7961);
buf BUF1 (N7992, N7986);
buf BUF1 (N7993, N7988);
xor XOR2 (N7994, N7987, N3295);
or OR3 (N7995, N7991, N918, N2874);
buf BUF1 (N7996, N7990);
not NOT1 (N7997, N7974);
or OR3 (N7998, N7953, N1926, N6940);
buf BUF1 (N7999, N7994);
not NOT1 (N8000, N7998);
or OR3 (N8001, N7983, N6076, N318);
or OR4 (N8002, N8000, N2270, N2514, N1168);
or OR3 (N8003, N7999, N2267, N1059);
or OR4 (N8004, N8002, N4212, N2589, N1014);
nand NAND3 (N8005, N7996, N2954, N7141);
buf BUF1 (N8006, N7993);
not NOT1 (N8007, N7997);
nor NOR2 (N8008, N8004, N2866);
buf BUF1 (N8009, N8003);
xor XOR2 (N8010, N7989, N4120);
nand NAND2 (N8011, N8006, N69);
or OR3 (N8012, N7995, N2946, N4855);
or OR4 (N8013, N8009, N2004, N4432, N3441);
buf BUF1 (N8014, N8005);
xor XOR2 (N8015, N8010, N3344);
not NOT1 (N8016, N8014);
nor NOR4 (N8017, N8013, N7624, N574, N234);
buf BUF1 (N8018, N8008);
xor XOR2 (N8019, N8007, N1857);
and AND3 (N8020, N8019, N3708, N5993);
and AND4 (N8021, N8012, N2749, N1980, N7098);
and AND3 (N8022, N8011, N3455, N1310);
xor XOR2 (N8023, N7981, N4238);
nor NOR3 (N8024, N8020, N7504, N2837);
not NOT1 (N8025, N8001);
or OR2 (N8026, N8018, N1364);
and AND2 (N8027, N8022, N2217);
nor NOR2 (N8028, N8023, N1121);
nor NOR4 (N8029, N8028, N2850, N6598, N7771);
buf BUF1 (N8030, N8026);
not NOT1 (N8031, N8021);
xor XOR2 (N8032, N7992, N2678);
xor XOR2 (N8033, N8027, N4400);
and AND4 (N8034, N8015, N4328, N1735, N4914);
nor NOR3 (N8035, N8032, N7504, N2183);
buf BUF1 (N8036, N8031);
nor NOR2 (N8037, N8036, N1556);
nor NOR3 (N8038, N8030, N4108, N1577);
not NOT1 (N8039, N8038);
nand NAND3 (N8040, N8029, N7813, N7552);
nand NAND4 (N8041, N8025, N533, N1371, N5296);
not NOT1 (N8042, N8035);
nand NAND2 (N8043, N8017, N526);
nand NAND4 (N8044, N8034, N1532, N6350, N4620);
buf BUF1 (N8045, N8044);
and AND2 (N8046, N8040, N6171);
nor NOR3 (N8047, N8033, N7306, N2653);
and AND3 (N8048, N8047, N119, N2051);
xor XOR2 (N8049, N8024, N2933);
and AND3 (N8050, N8037, N4130, N7612);
nand NAND3 (N8051, N8050, N1873, N4744);
buf BUF1 (N8052, N8042);
nor NOR2 (N8053, N8039, N4641);
nor NOR3 (N8054, N8043, N4359, N1689);
and AND2 (N8055, N8049, N6216);
nand NAND3 (N8056, N8052, N5305, N6008);
nor NOR4 (N8057, N8055, N950, N3988, N3514);
xor XOR2 (N8058, N8057, N4284);
not NOT1 (N8059, N8058);
nor NOR4 (N8060, N8051, N6341, N6218, N7679);
buf BUF1 (N8061, N8059);
xor XOR2 (N8062, N8056, N3008);
nor NOR2 (N8063, N8045, N5277);
nand NAND2 (N8064, N8046, N3777);
nand NAND3 (N8065, N8054, N3739, N6455);
and AND4 (N8066, N8063, N4071, N5451, N7161);
and AND2 (N8067, N8061, N6027);
or OR2 (N8068, N8064, N3776);
or OR3 (N8069, N8016, N7830, N4882);
or OR2 (N8070, N8041, N1637);
or OR4 (N8071, N8060, N6067, N732, N5291);
or OR4 (N8072, N8053, N4707, N3394, N7265);
or OR3 (N8073, N8068, N923, N7417);
buf BUF1 (N8074, N8048);
xor XOR2 (N8075, N8070, N1170);
buf BUF1 (N8076, N8073);
not NOT1 (N8077, N8071);
not NOT1 (N8078, N8075);
not NOT1 (N8079, N8069);
xor XOR2 (N8080, N8076, N5939);
nand NAND2 (N8081, N8062, N8061);
not NOT1 (N8082, N8081);
nand NAND3 (N8083, N8078, N1244, N4170);
xor XOR2 (N8084, N8079, N35);
buf BUF1 (N8085, N8082);
or OR4 (N8086, N8065, N4953, N3095, N7981);
nand NAND3 (N8087, N8086, N2642, N7796);
nand NAND4 (N8088, N8084, N3244, N46, N2706);
or OR2 (N8089, N8085, N6580);
xor XOR2 (N8090, N8080, N1293);
or OR4 (N8091, N8066, N6742, N65, N6132);
or OR3 (N8092, N8090, N4511, N3814);
or OR4 (N8093, N8072, N7616, N3544, N3987);
not NOT1 (N8094, N8083);
nand NAND4 (N8095, N8094, N7894, N2608, N1092);
nor NOR4 (N8096, N8089, N774, N1369, N1929);
and AND3 (N8097, N8095, N5402, N5898);
nor NOR4 (N8098, N8091, N7515, N6263, N5111);
not NOT1 (N8099, N8077);
and AND2 (N8100, N8099, N3435);
nand NAND4 (N8101, N8097, N414, N1820, N1392);
and AND3 (N8102, N8088, N4638, N2445);
xor XOR2 (N8103, N8087, N7194);
xor XOR2 (N8104, N8098, N7037);
xor XOR2 (N8105, N8104, N6537);
nand NAND2 (N8106, N8100, N857);
and AND3 (N8107, N8101, N1227, N592);
and AND3 (N8108, N8105, N7657, N4134);
nor NOR4 (N8109, N8067, N7872, N6905, N5765);
and AND3 (N8110, N8109, N3178, N726);
or OR4 (N8111, N8108, N3295, N1240, N2721);
or OR4 (N8112, N8111, N5857, N2915, N6017);
not NOT1 (N8113, N8092);
nor NOR4 (N8114, N8103, N4127, N6544, N1049);
or OR3 (N8115, N8074, N5779, N5003);
xor XOR2 (N8116, N8096, N2687);
xor XOR2 (N8117, N8107, N5118);
buf BUF1 (N8118, N8102);
xor XOR2 (N8119, N8112, N6253);
xor XOR2 (N8120, N8093, N2281);
xor XOR2 (N8121, N8116, N1054);
nor NOR4 (N8122, N8115, N3003, N2785, N4185);
or OR3 (N8123, N8106, N2313, N2632);
and AND4 (N8124, N8113, N1511, N6315, N5264);
nor NOR4 (N8125, N8123, N6750, N2272, N4024);
or OR4 (N8126, N8110, N6439, N5483, N8022);
not NOT1 (N8127, N8124);
xor XOR2 (N8128, N8127, N2886);
or OR4 (N8129, N8120, N4450, N7950, N7745);
or OR2 (N8130, N8129, N1457);
nand NAND4 (N8131, N8119, N7183, N6397, N2724);
nor NOR3 (N8132, N8117, N6734, N7944);
nor NOR3 (N8133, N8130, N5069, N1932);
nor NOR4 (N8134, N8125, N2012, N947, N5138);
xor XOR2 (N8135, N8118, N583);
xor XOR2 (N8136, N8128, N2685);
xor XOR2 (N8137, N8136, N6844);
or OR3 (N8138, N8132, N3614, N6013);
or OR2 (N8139, N8114, N5063);
buf BUF1 (N8140, N8137);
and AND4 (N8141, N8131, N2707, N7036, N6681);
and AND3 (N8142, N8139, N109, N1017);
not NOT1 (N8143, N8140);
nor NOR2 (N8144, N8141, N7431);
buf BUF1 (N8145, N8121);
nand NAND3 (N8146, N8144, N4743, N5249);
and AND4 (N8147, N8133, N6258, N5154, N90);
xor XOR2 (N8148, N8122, N5179);
and AND4 (N8149, N8135, N5380, N2065, N6017);
buf BUF1 (N8150, N8134);
or OR3 (N8151, N8143, N1043, N664);
buf BUF1 (N8152, N8149);
or OR3 (N8153, N8142, N4988, N3470);
nor NOR4 (N8154, N8148, N7047, N2178, N1940);
nand NAND3 (N8155, N8126, N7871, N5331);
nand NAND3 (N8156, N8151, N2144, N5747);
nor NOR4 (N8157, N8155, N5253, N4911, N273);
buf BUF1 (N8158, N8152);
nor NOR3 (N8159, N8145, N5084, N5665);
buf BUF1 (N8160, N8158);
nand NAND4 (N8161, N8153, N4499, N4438, N4887);
nand NAND3 (N8162, N8146, N5653, N1612);
or OR3 (N8163, N8159, N5093, N7277);
not NOT1 (N8164, N8150);
nand NAND3 (N8165, N8161, N1313, N5471);
or OR4 (N8166, N8157, N574, N1807, N5354);
buf BUF1 (N8167, N8138);
nor NOR3 (N8168, N8156, N5699, N5599);
and AND3 (N8169, N8167, N706, N6791);
nand NAND2 (N8170, N8162, N7981);
nand NAND3 (N8171, N8166, N4206, N5555);
nand NAND3 (N8172, N8169, N5482, N2225);
nor NOR2 (N8173, N8171, N2932);
not NOT1 (N8174, N8147);
nor NOR4 (N8175, N8170, N779, N6823, N5870);
not NOT1 (N8176, N8174);
xor XOR2 (N8177, N8165, N6832);
buf BUF1 (N8178, N8175);
buf BUF1 (N8179, N8173);
buf BUF1 (N8180, N8160);
xor XOR2 (N8181, N8163, N3787);
nand NAND3 (N8182, N8180, N516, N7472);
nor NOR2 (N8183, N8177, N2035);
or OR4 (N8184, N8172, N6678, N3806, N5081);
xor XOR2 (N8185, N8182, N5628);
nor NOR3 (N8186, N8184, N5988, N348);
not NOT1 (N8187, N8185);
and AND4 (N8188, N8186, N5734, N6199, N2490);
xor XOR2 (N8189, N8181, N4999);
buf BUF1 (N8190, N8183);
nand NAND2 (N8191, N8168, N2309);
or OR2 (N8192, N8179, N202);
and AND3 (N8193, N8187, N914, N4748);
and AND4 (N8194, N8193, N2668, N6134, N1493);
buf BUF1 (N8195, N8188);
nand NAND3 (N8196, N8154, N186, N893);
nor NOR2 (N8197, N8195, N6810);
not NOT1 (N8198, N8197);
nand NAND3 (N8199, N8196, N5428, N5204);
nand NAND4 (N8200, N8176, N276, N4713, N2608);
and AND3 (N8201, N8199, N6720, N3113);
nand NAND3 (N8202, N8194, N2187, N4051);
not NOT1 (N8203, N8164);
xor XOR2 (N8204, N8192, N3557);
or OR2 (N8205, N8200, N6351);
and AND3 (N8206, N8190, N3130, N5349);
buf BUF1 (N8207, N8201);
nand NAND3 (N8208, N8207, N366, N7292);
buf BUF1 (N8209, N8202);
not NOT1 (N8210, N8178);
not NOT1 (N8211, N8198);
nand NAND4 (N8212, N8211, N5094, N1581, N2249);
nand NAND4 (N8213, N8209, N6177, N6332, N3955);
nand NAND4 (N8214, N8203, N5007, N367, N7669);
buf BUF1 (N8215, N8205);
or OR3 (N8216, N8204, N2816, N1535);
not NOT1 (N8217, N8189);
xor XOR2 (N8218, N8213, N2716);
nor NOR3 (N8219, N8215, N5285, N2438);
nand NAND3 (N8220, N8210, N5435, N6156);
xor XOR2 (N8221, N8219, N2637);
or OR4 (N8222, N8217, N7145, N530, N6754);
and AND4 (N8223, N8222, N565, N8197, N5413);
xor XOR2 (N8224, N8191, N702);
not NOT1 (N8225, N8214);
nor NOR3 (N8226, N8218, N224, N1633);
and AND3 (N8227, N8206, N4304, N8153);
nand NAND3 (N8228, N8224, N2575, N8047);
xor XOR2 (N8229, N8226, N4547);
or OR2 (N8230, N8208, N5642);
buf BUF1 (N8231, N8216);
nor NOR3 (N8232, N8225, N3550, N7499);
or OR2 (N8233, N8231, N7839);
or OR3 (N8234, N8223, N2197, N3645);
and AND3 (N8235, N8234, N6118, N6499);
xor XOR2 (N8236, N8232, N1772);
buf BUF1 (N8237, N8212);
xor XOR2 (N8238, N8221, N6101);
nand NAND4 (N8239, N8237, N6596, N3453, N2295);
nand NAND2 (N8240, N8229, N7433);
or OR3 (N8241, N8236, N5391, N4588);
and AND2 (N8242, N8239, N4282);
buf BUF1 (N8243, N8235);
and AND3 (N8244, N8238, N1037, N1087);
xor XOR2 (N8245, N8228, N1092);
not NOT1 (N8246, N8220);
nand NAND3 (N8247, N8244, N4864, N6258);
nor NOR4 (N8248, N8240, N5887, N2830, N3002);
or OR3 (N8249, N8242, N296, N2000);
and AND4 (N8250, N8230, N5313, N5998, N4264);
xor XOR2 (N8251, N8233, N1250);
nand NAND4 (N8252, N8250, N7798, N5309, N4020);
or OR2 (N8253, N8252, N912);
and AND3 (N8254, N8247, N7119, N5751);
nand NAND4 (N8255, N8251, N3488, N2311, N4703);
not NOT1 (N8256, N8249);
not NOT1 (N8257, N8255);
or OR4 (N8258, N8241, N1317, N7876, N5644);
not NOT1 (N8259, N8253);
not NOT1 (N8260, N8259);
and AND3 (N8261, N8260, N7523, N5484);
buf BUF1 (N8262, N8256);
nor NOR3 (N8263, N8257, N1704, N4804);
nand NAND3 (N8264, N8248, N7188, N2678);
buf BUF1 (N8265, N8227);
buf BUF1 (N8266, N8263);
nand NAND3 (N8267, N8258, N5924, N842);
or OR2 (N8268, N8262, N3620);
buf BUF1 (N8269, N8243);
and AND2 (N8270, N8264, N2700);
xor XOR2 (N8271, N8269, N40);
or OR2 (N8272, N8266, N1076);
and AND4 (N8273, N8267, N7448, N2097, N7473);
or OR2 (N8274, N8271, N5843);
not NOT1 (N8275, N8246);
not NOT1 (N8276, N8265);
or OR3 (N8277, N8272, N3144, N7750);
or OR4 (N8278, N8274, N7931, N7591, N1008);
xor XOR2 (N8279, N8261, N2137);
or OR4 (N8280, N8278, N5528, N1602, N1884);
nor NOR2 (N8281, N8280, N3401);
nor NOR3 (N8282, N8276, N2, N1901);
nand NAND4 (N8283, N8270, N3306, N6194, N3792);
nor NOR3 (N8284, N8281, N2527, N2684);
buf BUF1 (N8285, N8279);
nand NAND4 (N8286, N8285, N1314, N3309, N7033);
or OR2 (N8287, N8283, N5833);
nand NAND3 (N8288, N8245, N657, N2209);
buf BUF1 (N8289, N8277);
not NOT1 (N8290, N8289);
not NOT1 (N8291, N8254);
buf BUF1 (N8292, N8284);
or OR3 (N8293, N8268, N3611, N2371);
or OR3 (N8294, N8275, N7506, N8081);
and AND3 (N8295, N8287, N1069, N5196);
nor NOR3 (N8296, N8292, N2076, N7573);
xor XOR2 (N8297, N8288, N5483);
or OR3 (N8298, N8282, N2364, N2381);
buf BUF1 (N8299, N8294);
xor XOR2 (N8300, N8290, N1884);
nand NAND4 (N8301, N8297, N4113, N2425, N4249);
nor NOR2 (N8302, N8291, N6018);
not NOT1 (N8303, N8298);
or OR4 (N8304, N8299, N5664, N4239, N3582);
nand NAND2 (N8305, N8302, N1962);
nor NOR4 (N8306, N8304, N6613, N6672, N5242);
or OR4 (N8307, N8306, N1701, N6768, N6448);
xor XOR2 (N8308, N8300, N4608);
and AND2 (N8309, N8301, N2921);
or OR4 (N8310, N8309, N6698, N5709, N2946);
nor NOR2 (N8311, N8293, N335);
xor XOR2 (N8312, N8303, N481);
or OR3 (N8313, N8310, N2911, N1039);
buf BUF1 (N8314, N8305);
and AND4 (N8315, N8314, N262, N6911, N2712);
nand NAND2 (N8316, N8311, N1989);
xor XOR2 (N8317, N8308, N5420);
buf BUF1 (N8318, N8273);
nand NAND2 (N8319, N8307, N353);
xor XOR2 (N8320, N8315, N2356);
buf BUF1 (N8321, N8316);
xor XOR2 (N8322, N8313, N6389);
buf BUF1 (N8323, N8296);
xor XOR2 (N8324, N8319, N7173);
nor NOR3 (N8325, N8312, N959, N2140);
or OR4 (N8326, N8325, N1149, N6012, N1909);
nor NOR4 (N8327, N8323, N5417, N3341, N6789);
and AND4 (N8328, N8320, N4026, N7975, N5735);
nand NAND4 (N8329, N8328, N5671, N3429, N112);
not NOT1 (N8330, N8295);
or OR2 (N8331, N8327, N8220);
or OR3 (N8332, N8329, N948, N7008);
nand NAND2 (N8333, N8322, N6414);
buf BUF1 (N8334, N8321);
buf BUF1 (N8335, N8324);
buf BUF1 (N8336, N8330);
or OR2 (N8337, N8336, N128);
nand NAND2 (N8338, N8332, N2405);
or OR2 (N8339, N8326, N4993);
nor NOR4 (N8340, N8318, N2072, N1445, N2729);
buf BUF1 (N8341, N8338);
and AND3 (N8342, N8341, N3801, N1402);
and AND3 (N8343, N8334, N6881, N7977);
not NOT1 (N8344, N8317);
nor NOR3 (N8345, N8343, N2471, N991);
buf BUF1 (N8346, N8344);
nand NAND2 (N8347, N8345, N676);
or OR3 (N8348, N8339, N7789, N4584);
and AND3 (N8349, N8342, N4709, N2823);
xor XOR2 (N8350, N8337, N1423);
buf BUF1 (N8351, N8286);
nand NAND4 (N8352, N8347, N8289, N3202, N303);
nand NAND3 (N8353, N8348, N6036, N764);
nor NOR2 (N8354, N8346, N2821);
nand NAND3 (N8355, N8350, N592, N4858);
and AND2 (N8356, N8335, N3166);
or OR4 (N8357, N8353, N1677, N4508, N755);
and AND4 (N8358, N8333, N392, N6696, N3048);
nand NAND2 (N8359, N8351, N87);
xor XOR2 (N8360, N8340, N2710);
and AND2 (N8361, N8331, N853);
xor XOR2 (N8362, N8356, N7139);
and AND2 (N8363, N8352, N7077);
nand NAND2 (N8364, N8362, N7446);
or OR2 (N8365, N8358, N671);
or OR3 (N8366, N8363, N3687, N706);
and AND3 (N8367, N8366, N2877, N1268);
not NOT1 (N8368, N8367);
and AND4 (N8369, N8360, N700, N3725, N4199);
nand NAND2 (N8370, N8364, N3175);
xor XOR2 (N8371, N8355, N4103);
not NOT1 (N8372, N8354);
nand NAND4 (N8373, N8370, N7599, N1580, N4841);
not NOT1 (N8374, N8361);
xor XOR2 (N8375, N8357, N203);
nor NOR3 (N8376, N8372, N6905, N2723);
and AND2 (N8377, N8349, N5328);
not NOT1 (N8378, N8376);
xor XOR2 (N8379, N8359, N705);
buf BUF1 (N8380, N8375);
nor NOR3 (N8381, N8369, N6948, N1616);
xor XOR2 (N8382, N8381, N7072);
buf BUF1 (N8383, N8382);
and AND2 (N8384, N8368, N2114);
and AND3 (N8385, N8383, N4675, N6522);
nor NOR2 (N8386, N8380, N5286);
not NOT1 (N8387, N8371);
not NOT1 (N8388, N8384);
nand NAND2 (N8389, N8377, N5721);
nand NAND3 (N8390, N8389, N4043, N5008);
xor XOR2 (N8391, N8373, N7609);
and AND2 (N8392, N8365, N4268);
and AND4 (N8393, N8388, N404, N3067, N2068);
nand NAND3 (N8394, N8378, N3541, N3832);
or OR4 (N8395, N8390, N4023, N8175, N3984);
nor NOR3 (N8396, N8379, N7450, N563);
xor XOR2 (N8397, N8395, N3215);
not NOT1 (N8398, N8387);
and AND3 (N8399, N8392, N3355, N2146);
nand NAND3 (N8400, N8399, N7035, N7291);
xor XOR2 (N8401, N8386, N5592);
buf BUF1 (N8402, N8396);
buf BUF1 (N8403, N8398);
xor XOR2 (N8404, N8385, N4480);
nor NOR4 (N8405, N8391, N939, N1431, N6760);
xor XOR2 (N8406, N8374, N2506);
nand NAND2 (N8407, N8405, N90);
buf BUF1 (N8408, N8393);
and AND4 (N8409, N8394, N4577, N1032, N3278);
or OR4 (N8410, N8409, N7866, N3906, N73);
buf BUF1 (N8411, N8404);
nor NOR3 (N8412, N8408, N2574, N619);
or OR3 (N8413, N8402, N3739, N989);
nor NOR4 (N8414, N8412, N5046, N1844, N4688);
nand NAND4 (N8415, N8410, N4009, N1762, N6731);
nor NOR2 (N8416, N8415, N139);
xor XOR2 (N8417, N8414, N2070);
and AND2 (N8418, N8403, N6167);
or OR3 (N8419, N8406, N1693, N8363);
xor XOR2 (N8420, N8397, N381);
not NOT1 (N8421, N8401);
buf BUF1 (N8422, N8418);
xor XOR2 (N8423, N8421, N7196);
nand NAND2 (N8424, N8419, N2456);
nand NAND3 (N8425, N8424, N4508, N803);
not NOT1 (N8426, N8407);
or OR2 (N8427, N8416, N567);
nor NOR2 (N8428, N8425, N4391);
nand NAND4 (N8429, N8426, N4211, N3111, N4934);
and AND4 (N8430, N8422, N99, N7874, N2306);
nor NOR2 (N8431, N8423, N4954);
nand NAND4 (N8432, N8428, N3191, N790, N5835);
buf BUF1 (N8433, N8413);
nor NOR3 (N8434, N8430, N5803, N3762);
and AND2 (N8435, N8417, N5387);
or OR4 (N8436, N8420, N119, N5193, N665);
or OR3 (N8437, N8434, N1409, N2241);
nor NOR3 (N8438, N8437, N7899, N2295);
nand NAND3 (N8439, N8436, N8116, N3704);
xor XOR2 (N8440, N8435, N5973);
xor XOR2 (N8441, N8432, N3392);
nand NAND4 (N8442, N8440, N550, N8043, N6255);
xor XOR2 (N8443, N8433, N1611);
or OR4 (N8444, N8429, N7463, N2376, N4759);
xor XOR2 (N8445, N8442, N4553);
buf BUF1 (N8446, N8445);
xor XOR2 (N8447, N8444, N2660);
nand NAND3 (N8448, N8427, N6328, N5404);
buf BUF1 (N8449, N8411);
and AND3 (N8450, N8446, N339, N7662);
or OR4 (N8451, N8400, N2650, N6998, N6177);
not NOT1 (N8452, N8441);
buf BUF1 (N8453, N8438);
nor NOR4 (N8454, N8451, N5046, N5706, N3971);
xor XOR2 (N8455, N8449, N1376);
buf BUF1 (N8456, N8455);
buf BUF1 (N8457, N8443);
nor NOR3 (N8458, N8450, N508, N2253);
xor XOR2 (N8459, N8456, N2076);
nand NAND2 (N8460, N8431, N1822);
nand NAND2 (N8461, N8460, N5486);
nand NAND4 (N8462, N8461, N107, N987, N2991);
nor NOR2 (N8463, N8447, N2040);
xor XOR2 (N8464, N8448, N4737);
nor NOR2 (N8465, N8453, N1202);
xor XOR2 (N8466, N8464, N6496);
buf BUF1 (N8467, N8454);
not NOT1 (N8468, N8457);
and AND4 (N8469, N8465, N2861, N535, N2484);
or OR3 (N8470, N8466, N1189, N1989);
and AND2 (N8471, N8469, N2909);
nand NAND2 (N8472, N8458, N5587);
nor NOR3 (N8473, N8472, N1774, N2626);
nor NOR2 (N8474, N8468, N7654);
nand NAND2 (N8475, N8462, N4712);
xor XOR2 (N8476, N8439, N5821);
nand NAND2 (N8477, N8470, N1632);
nor NOR3 (N8478, N8474, N6085, N7574);
xor XOR2 (N8479, N8467, N4893);
nor NOR4 (N8480, N8477, N1493, N558, N798);
buf BUF1 (N8481, N8480);
buf BUF1 (N8482, N8459);
buf BUF1 (N8483, N8475);
or OR2 (N8484, N8452, N197);
nor NOR4 (N8485, N8476, N1058, N325, N979);
or OR2 (N8486, N8478, N8383);
xor XOR2 (N8487, N8471, N3909);
nor NOR4 (N8488, N8486, N5952, N3929, N1388);
nand NAND3 (N8489, N8481, N709, N5783);
nand NAND3 (N8490, N8483, N8255, N8124);
not NOT1 (N8491, N8488);
not NOT1 (N8492, N8484);
and AND4 (N8493, N8489, N2759, N1223, N2228);
not NOT1 (N8494, N8482);
buf BUF1 (N8495, N8492);
nor NOR3 (N8496, N8491, N6343, N4481);
not NOT1 (N8497, N8473);
nand NAND3 (N8498, N8493, N5149, N5108);
nand NAND2 (N8499, N8490, N7159);
nand NAND2 (N8500, N8496, N8296);
and AND3 (N8501, N8495, N6425, N5084);
nor NOR3 (N8502, N8494, N5407, N5163);
and AND4 (N8503, N8499, N2532, N1898, N1160);
buf BUF1 (N8504, N8503);
and AND3 (N8505, N8500, N3501, N2730);
nor NOR4 (N8506, N8498, N3902, N2481, N1168);
xor XOR2 (N8507, N8497, N4645);
not NOT1 (N8508, N8487);
buf BUF1 (N8509, N8507);
xor XOR2 (N8510, N8509, N593);
not NOT1 (N8511, N8505);
xor XOR2 (N8512, N8504, N3966);
and AND3 (N8513, N8501, N4727, N7457);
nand NAND4 (N8514, N8513, N1949, N4720, N5413);
and AND3 (N8515, N8479, N3552, N7900);
or OR4 (N8516, N8463, N8206, N6731, N4802);
nand NAND4 (N8517, N8510, N2062, N2051, N7575);
xor XOR2 (N8518, N8502, N897);
nand NAND3 (N8519, N8516, N8251, N6203);
xor XOR2 (N8520, N8519, N6858);
nand NAND4 (N8521, N8515, N1799, N8383, N1593);
nand NAND3 (N8522, N8517, N868, N2645);
buf BUF1 (N8523, N8514);
or OR4 (N8524, N8522, N3298, N4766, N6720);
nor NOR2 (N8525, N8521, N4767);
buf BUF1 (N8526, N8523);
xor XOR2 (N8527, N8520, N3536);
or OR4 (N8528, N8485, N2703, N3839, N4740);
nand NAND4 (N8529, N8525, N2022, N1158, N4387);
not NOT1 (N8530, N8529);
xor XOR2 (N8531, N8528, N3831);
buf BUF1 (N8532, N8530);
or OR3 (N8533, N8518, N717, N925);
and AND4 (N8534, N8512, N4341, N880, N3607);
not NOT1 (N8535, N8511);
or OR3 (N8536, N8526, N2368, N548);
nor NOR3 (N8537, N8532, N3220, N862);
not NOT1 (N8538, N8534);
or OR4 (N8539, N8535, N2430, N2012, N7016);
and AND4 (N8540, N8533, N751, N71, N2383);
buf BUF1 (N8541, N8508);
and AND3 (N8542, N8537, N4042, N4316);
not NOT1 (N8543, N8540);
nand NAND2 (N8544, N8524, N7703);
xor XOR2 (N8545, N8543, N4106);
buf BUF1 (N8546, N8541);
nand NAND4 (N8547, N8545, N5012, N7563, N745);
nand NAND4 (N8548, N8539, N5, N5580, N4649);
nand NAND3 (N8549, N8547, N4581, N2550);
and AND2 (N8550, N8544, N310);
or OR3 (N8551, N8548, N7169, N7897);
nand NAND2 (N8552, N8527, N979);
not NOT1 (N8553, N8546);
nor NOR3 (N8554, N8552, N4992, N4647);
or OR2 (N8555, N8538, N8291);
not NOT1 (N8556, N8551);
nand NAND4 (N8557, N8554, N5352, N2564, N3845);
buf BUF1 (N8558, N8557);
buf BUF1 (N8559, N8542);
nor NOR3 (N8560, N8536, N4661, N944);
xor XOR2 (N8561, N8555, N3625);
and AND4 (N8562, N8560, N3619, N5461, N1097);
or OR2 (N8563, N8558, N3164);
or OR2 (N8564, N8562, N2148);
not NOT1 (N8565, N8531);
nor NOR3 (N8566, N8564, N6055, N6135);
buf BUF1 (N8567, N8549);
and AND2 (N8568, N8567, N729);
nand NAND2 (N8569, N8563, N2085);
xor XOR2 (N8570, N8565, N6473);
buf BUF1 (N8571, N8569);
xor XOR2 (N8572, N8556, N5194);
and AND3 (N8573, N8572, N5606, N3939);
nand NAND3 (N8574, N8568, N4115, N1225);
xor XOR2 (N8575, N8553, N5343);
or OR3 (N8576, N8575, N2741, N6583);
nor NOR3 (N8577, N8566, N3089, N2955);
or OR2 (N8578, N8571, N2092);
not NOT1 (N8579, N8573);
nand NAND4 (N8580, N8550, N5809, N2973, N3624);
not NOT1 (N8581, N8579);
not NOT1 (N8582, N8581);
and AND2 (N8583, N8570, N1876);
or OR4 (N8584, N8577, N8355, N2398, N6179);
nor NOR4 (N8585, N8580, N6000, N8453, N4652);
and AND2 (N8586, N8561, N1024);
xor XOR2 (N8587, N8582, N2903);
nor NOR4 (N8588, N8578, N5526, N221, N7574);
buf BUF1 (N8589, N8588);
and AND3 (N8590, N8587, N5890, N5283);
not NOT1 (N8591, N8583);
or OR3 (N8592, N8590, N7493, N8511);
buf BUF1 (N8593, N8586);
not NOT1 (N8594, N8585);
nand NAND3 (N8595, N8559, N6856, N5418);
nor NOR2 (N8596, N8506, N3049);
not NOT1 (N8597, N8593);
not NOT1 (N8598, N8589);
buf BUF1 (N8599, N8597);
not NOT1 (N8600, N8591);
nand NAND2 (N8601, N8592, N6062);
buf BUF1 (N8602, N8576);
xor XOR2 (N8603, N8601, N3233);
nand NAND4 (N8604, N8596, N4657, N8251, N7987);
nand NAND3 (N8605, N8594, N5836, N7021);
or OR4 (N8606, N8574, N5266, N2439, N1405);
xor XOR2 (N8607, N8599, N6090);
not NOT1 (N8608, N8604);
nand NAND3 (N8609, N8605, N5878, N6722);
nor NOR4 (N8610, N8584, N8441, N7339, N8424);
nor NOR4 (N8611, N8607, N3852, N6268, N6677);
buf BUF1 (N8612, N8609);
nand NAND4 (N8613, N8595, N2118, N4729, N1371);
and AND2 (N8614, N8598, N4181);
nand NAND4 (N8615, N8603, N886, N3545, N3209);
nor NOR2 (N8616, N8611, N7820);
nor NOR4 (N8617, N8614, N1147, N4786, N8259);
not NOT1 (N8618, N8608);
buf BUF1 (N8619, N8612);
and AND4 (N8620, N8606, N5763, N2074, N1504);
nand NAND3 (N8621, N8610, N5543, N5215);
and AND4 (N8622, N8602, N3830, N4225, N6943);
nor NOR3 (N8623, N8613, N2846, N7302);
nand NAND4 (N8624, N8615, N2701, N4997, N4669);
and AND4 (N8625, N8623, N2027, N52, N8424);
buf BUF1 (N8626, N8619);
not NOT1 (N8627, N8620);
or OR3 (N8628, N8627, N1964, N7270);
nand NAND4 (N8629, N8626, N4017, N6458, N5225);
buf BUF1 (N8630, N8628);
and AND4 (N8631, N8625, N6126, N6338, N5284);
buf BUF1 (N8632, N8629);
buf BUF1 (N8633, N8621);
or OR3 (N8634, N8618, N6522, N3306);
not NOT1 (N8635, N8616);
not NOT1 (N8636, N8633);
nor NOR3 (N8637, N8634, N1119, N6375);
nor NOR3 (N8638, N8636, N1870, N5260);
not NOT1 (N8639, N8624);
xor XOR2 (N8640, N8622, N6777);
xor XOR2 (N8641, N8630, N351);
buf BUF1 (N8642, N8638);
nand NAND2 (N8643, N8642, N5491);
not NOT1 (N8644, N8617);
nand NAND4 (N8645, N8635, N6798, N8065, N8211);
nand NAND2 (N8646, N8631, N766);
not NOT1 (N8647, N8600);
not NOT1 (N8648, N8644);
and AND2 (N8649, N8647, N6031);
xor XOR2 (N8650, N8649, N47);
nor NOR4 (N8651, N8648, N5794, N1092, N5168);
nand NAND2 (N8652, N8651, N1591);
or OR4 (N8653, N8650, N3903, N5942, N7000);
nand NAND4 (N8654, N8639, N1390, N2276, N4100);
or OR2 (N8655, N8632, N767);
or OR4 (N8656, N8643, N6512, N6418, N8497);
and AND4 (N8657, N8652, N4787, N5916, N8615);
or OR3 (N8658, N8657, N4976, N3140);
buf BUF1 (N8659, N8646);
nand NAND3 (N8660, N8658, N4422, N4095);
xor XOR2 (N8661, N8640, N3007);
and AND4 (N8662, N8653, N6763, N3314, N6865);
buf BUF1 (N8663, N8645);
or OR3 (N8664, N8659, N1022, N7405);
nor NOR4 (N8665, N8641, N7606, N5394, N1980);
not NOT1 (N8666, N8656);
or OR4 (N8667, N8663, N4976, N5047, N846);
not NOT1 (N8668, N8665);
nand NAND4 (N8669, N8660, N4576, N7800, N4777);
nor NOR4 (N8670, N8637, N7642, N3270, N6389);
nand NAND3 (N8671, N8670, N6104, N2220);
not NOT1 (N8672, N8654);
or OR4 (N8673, N8661, N3013, N8648, N6806);
nand NAND3 (N8674, N8672, N4106, N5097);
or OR3 (N8675, N8673, N6831, N7717);
not NOT1 (N8676, N8668);
or OR3 (N8677, N8664, N1182, N1408);
nand NAND2 (N8678, N8666, N7979);
or OR2 (N8679, N8678, N8203);
xor XOR2 (N8680, N8679, N6790);
and AND2 (N8681, N8662, N340);
buf BUF1 (N8682, N8671);
not NOT1 (N8683, N8667);
and AND2 (N8684, N8683, N2271);
buf BUF1 (N8685, N8674);
nor NOR3 (N8686, N8677, N4220, N7725);
xor XOR2 (N8687, N8675, N2591);
or OR2 (N8688, N8684, N6926);
nor NOR2 (N8689, N8676, N5822);
xor XOR2 (N8690, N8682, N695);
nor NOR4 (N8691, N8689, N458, N1120, N5349);
nor NOR3 (N8692, N8691, N3141, N5741);
or OR3 (N8693, N8685, N133, N4824);
nor NOR2 (N8694, N8686, N5905);
and AND3 (N8695, N8687, N4661, N5467);
nor NOR2 (N8696, N8692, N529);
xor XOR2 (N8697, N8696, N6628);
buf BUF1 (N8698, N8681);
nor NOR2 (N8699, N8669, N2388);
and AND3 (N8700, N8688, N5521, N8379);
buf BUF1 (N8701, N8700);
nor NOR3 (N8702, N8697, N5477, N4242);
nor NOR2 (N8703, N8690, N6308);
buf BUF1 (N8704, N8703);
and AND3 (N8705, N8655, N3757, N1738);
nand NAND4 (N8706, N8699, N172, N116, N999);
nand NAND2 (N8707, N8680, N2198);
xor XOR2 (N8708, N8694, N182);
xor XOR2 (N8709, N8704, N1150);
xor XOR2 (N8710, N8709, N6123);
xor XOR2 (N8711, N8708, N6878);
buf BUF1 (N8712, N8695);
not NOT1 (N8713, N8701);
and AND3 (N8714, N8702, N4457, N949);
not NOT1 (N8715, N8693);
or OR2 (N8716, N8711, N229);
nand NAND3 (N8717, N8698, N1262, N448);
not NOT1 (N8718, N8706);
nor NOR3 (N8719, N8716, N3136, N1604);
not NOT1 (N8720, N8719);
nor NOR4 (N8721, N8717, N4995, N7848, N3871);
buf BUF1 (N8722, N8720);
xor XOR2 (N8723, N8722, N700);
nand NAND2 (N8724, N8721, N237);
buf BUF1 (N8725, N8723);
nand NAND4 (N8726, N8724, N1171, N184, N5415);
xor XOR2 (N8727, N8715, N3160);
or OR2 (N8728, N8705, N4980);
buf BUF1 (N8729, N8725);
and AND4 (N8730, N8710, N3284, N6343, N249);
or OR4 (N8731, N8726, N6249, N3512, N6484);
buf BUF1 (N8732, N8707);
nor NOR2 (N8733, N8731, N8384);
or OR2 (N8734, N8718, N3567);
nand NAND4 (N8735, N8728, N3065, N2287, N5627);
nor NOR4 (N8736, N8730, N4302, N5057, N1791);
nand NAND4 (N8737, N8727, N7661, N3319, N7103);
or OR4 (N8738, N8732, N8384, N3501, N7329);
xor XOR2 (N8739, N8729, N1660);
not NOT1 (N8740, N8735);
nor NOR4 (N8741, N8712, N2347, N3067, N1258);
not NOT1 (N8742, N8734);
nand NAND2 (N8743, N8740, N6332);
buf BUF1 (N8744, N8736);
nand NAND2 (N8745, N8743, N1866);
not NOT1 (N8746, N8741);
xor XOR2 (N8747, N8744, N958);
nor NOR4 (N8748, N8747, N8065, N3155, N862);
not NOT1 (N8749, N8739);
xor XOR2 (N8750, N8745, N626);
or OR3 (N8751, N8713, N8372, N4765);
not NOT1 (N8752, N8738);
or OR3 (N8753, N8752, N2797, N1780);
not NOT1 (N8754, N8751);
nor NOR2 (N8755, N8733, N2533);
nand NAND2 (N8756, N8755, N6300);
or OR2 (N8757, N8750, N2142);
not NOT1 (N8758, N8737);
xor XOR2 (N8759, N8753, N5843);
and AND4 (N8760, N8756, N3494, N5159, N3158);
buf BUF1 (N8761, N8757);
nor NOR2 (N8762, N8760, N8010);
xor XOR2 (N8763, N8714, N8604);
xor XOR2 (N8764, N8763, N8544);
xor XOR2 (N8765, N8761, N2623);
not NOT1 (N8766, N8762);
and AND4 (N8767, N8754, N5233, N6181, N4773);
nor NOR4 (N8768, N8758, N7615, N1459, N4421);
or OR2 (N8769, N8766, N7806);
buf BUF1 (N8770, N8748);
not NOT1 (N8771, N8764);
not NOT1 (N8772, N8765);
nand NAND4 (N8773, N8769, N2403, N2604, N7898);
xor XOR2 (N8774, N8759, N2878);
nand NAND3 (N8775, N8771, N6681, N1926);
xor XOR2 (N8776, N8773, N57);
and AND3 (N8777, N8749, N7980, N7205);
xor XOR2 (N8778, N8742, N1547);
not NOT1 (N8779, N8775);
and AND4 (N8780, N8770, N797, N3838, N1212);
or OR4 (N8781, N8776, N3664, N3058, N3009);
nor NOR4 (N8782, N8768, N8499, N2666, N1615);
nor NOR4 (N8783, N8774, N1474, N3584, N5653);
xor XOR2 (N8784, N8777, N549);
or OR3 (N8785, N8784, N7545, N5260);
buf BUF1 (N8786, N8783);
buf BUF1 (N8787, N8786);
nor NOR2 (N8788, N8772, N3515);
or OR4 (N8789, N8746, N7812, N6312, N6989);
or OR2 (N8790, N8779, N246);
nand NAND4 (N8791, N8782, N6978, N2408, N1538);
or OR2 (N8792, N8785, N7251);
and AND2 (N8793, N8790, N7879);
xor XOR2 (N8794, N8793, N7292);
nand NAND2 (N8795, N8781, N1256);
buf BUF1 (N8796, N8788);
not NOT1 (N8797, N8794);
xor XOR2 (N8798, N8796, N572);
and AND4 (N8799, N8778, N3165, N7775, N8608);
buf BUF1 (N8800, N8799);
not NOT1 (N8801, N8797);
nor NOR2 (N8802, N8801, N5146);
nor NOR3 (N8803, N8767, N1402, N4645);
not NOT1 (N8804, N8792);
buf BUF1 (N8805, N8791);
or OR2 (N8806, N8787, N3546);
or OR2 (N8807, N8805, N4973);
or OR2 (N8808, N8795, N7788);
not NOT1 (N8809, N8804);
not NOT1 (N8810, N8780);
xor XOR2 (N8811, N8800, N8705);
nor NOR2 (N8812, N8806, N6476);
nor NOR2 (N8813, N8808, N949);
buf BUF1 (N8814, N8813);
xor XOR2 (N8815, N8809, N6176);
and AND2 (N8816, N8811, N4262);
nor NOR4 (N8817, N8816, N541, N346, N1385);
or OR2 (N8818, N8815, N6924);
or OR4 (N8819, N8803, N6886, N4415, N2586);
xor XOR2 (N8820, N8814, N5913);
not NOT1 (N8821, N8818);
not NOT1 (N8822, N8810);
nor NOR3 (N8823, N8802, N162, N5194);
nand NAND4 (N8824, N8823, N1135, N7160, N241);
and AND3 (N8825, N8812, N4849, N3686);
nand NAND2 (N8826, N8825, N7274);
or OR3 (N8827, N8822, N2773, N4625);
or OR3 (N8828, N8817, N7700, N1295);
and AND4 (N8829, N8807, N7721, N3670, N6437);
buf BUF1 (N8830, N8789);
nand NAND4 (N8831, N8829, N472, N5039, N3791);
buf BUF1 (N8832, N8819);
nand NAND4 (N8833, N8827, N336, N3460, N1965);
and AND2 (N8834, N8832, N8492);
nor NOR3 (N8835, N8821, N7552, N1857);
and AND4 (N8836, N8826, N1348, N3000, N7616);
not NOT1 (N8837, N8831);
xor XOR2 (N8838, N8828, N1701);
nand NAND4 (N8839, N8834, N4667, N1573, N5041);
not NOT1 (N8840, N8836);
and AND2 (N8841, N8830, N5663);
buf BUF1 (N8842, N8824);
xor XOR2 (N8843, N8835, N7901);
not NOT1 (N8844, N8820);
and AND2 (N8845, N8833, N443);
nor NOR4 (N8846, N8838, N980, N5417, N3818);
nand NAND2 (N8847, N8843, N3907);
buf BUF1 (N8848, N8839);
and AND2 (N8849, N8848, N3515);
nand NAND3 (N8850, N8849, N2166, N8599);
buf BUF1 (N8851, N8840);
xor XOR2 (N8852, N8846, N243);
and AND4 (N8853, N8841, N121, N774, N5745);
not NOT1 (N8854, N8844);
and AND3 (N8855, N8798, N6827, N7521);
nor NOR4 (N8856, N8854, N5020, N6787, N7388);
xor XOR2 (N8857, N8855, N956);
buf BUF1 (N8858, N8851);
nor NOR3 (N8859, N8842, N2964, N5570);
buf BUF1 (N8860, N8845);
nor NOR3 (N8861, N8837, N3941, N6376);
not NOT1 (N8862, N8847);
and AND3 (N8863, N8853, N352, N6309);
buf BUF1 (N8864, N8861);
and AND4 (N8865, N8859, N658, N5907, N2496);
or OR4 (N8866, N8850, N430, N2744, N2734);
buf BUF1 (N8867, N8865);
or OR3 (N8868, N8860, N6326, N5773);
nand NAND3 (N8869, N8867, N1807, N1566);
xor XOR2 (N8870, N8857, N2770);
nand NAND3 (N8871, N8868, N623, N8217);
nand NAND4 (N8872, N8870, N2921, N6897, N7736);
xor XOR2 (N8873, N8852, N3860);
nor NOR2 (N8874, N8872, N5149);
and AND2 (N8875, N8874, N3357);
or OR2 (N8876, N8862, N8431);
not NOT1 (N8877, N8856);
not NOT1 (N8878, N8864);
or OR2 (N8879, N8858, N8723);
buf BUF1 (N8880, N8873);
buf BUF1 (N8881, N8866);
and AND2 (N8882, N8871, N7178);
nor NOR4 (N8883, N8881, N2007, N566, N7531);
not NOT1 (N8884, N8882);
nor NOR3 (N8885, N8879, N8443, N2417);
not NOT1 (N8886, N8884);
or OR3 (N8887, N8880, N6031, N2625);
nand NAND4 (N8888, N8886, N156, N4908, N6453);
xor XOR2 (N8889, N8875, N2314);
and AND3 (N8890, N8878, N1308, N5589);
or OR2 (N8891, N8890, N6395);
nor NOR2 (N8892, N8869, N803);
not NOT1 (N8893, N8876);
xor XOR2 (N8894, N8885, N6364);
not NOT1 (N8895, N8892);
buf BUF1 (N8896, N8888);
buf BUF1 (N8897, N8889);
and AND2 (N8898, N8887, N1917);
not NOT1 (N8899, N8891);
not NOT1 (N8900, N8877);
nor NOR4 (N8901, N8897, N8052, N1744, N7818);
buf BUF1 (N8902, N8893);
not NOT1 (N8903, N8894);
buf BUF1 (N8904, N8895);
not NOT1 (N8905, N8899);
and AND2 (N8906, N8863, N7445);
buf BUF1 (N8907, N8900);
or OR3 (N8908, N8901, N646, N7181);
not NOT1 (N8909, N8902);
xor XOR2 (N8910, N8906, N6583);
nand NAND2 (N8911, N8904, N3122);
buf BUF1 (N8912, N8896);
and AND4 (N8913, N8911, N2275, N254, N7654);
and AND2 (N8914, N8912, N3332);
not NOT1 (N8915, N8914);
buf BUF1 (N8916, N8910);
or OR3 (N8917, N8909, N7324, N6944);
not NOT1 (N8918, N8898);
nand NAND4 (N8919, N8917, N4332, N1309, N6247);
not NOT1 (N8920, N8907);
or OR4 (N8921, N8903, N7405, N1439, N7681);
not NOT1 (N8922, N8883);
nand NAND3 (N8923, N8916, N7895, N8057);
or OR2 (N8924, N8913, N548);
or OR4 (N8925, N8918, N8182, N7088, N153);
and AND3 (N8926, N8924, N6410, N2383);
or OR3 (N8927, N8920, N7406, N1497);
nand NAND2 (N8928, N8919, N1194);
and AND2 (N8929, N8923, N2070);
not NOT1 (N8930, N8926);
nand NAND2 (N8931, N8921, N7165);
and AND4 (N8932, N8928, N6323, N8115, N6938);
and AND2 (N8933, N8927, N2336);
buf BUF1 (N8934, N8915);
nor NOR3 (N8935, N8925, N3517, N4607);
not NOT1 (N8936, N8935);
xor XOR2 (N8937, N8933, N1326);
and AND3 (N8938, N8936, N8146, N5498);
not NOT1 (N8939, N8938);
not NOT1 (N8940, N8937);
buf BUF1 (N8941, N8908);
and AND4 (N8942, N8931, N2365, N3329, N2583);
or OR2 (N8943, N8932, N2448);
and AND3 (N8944, N8922, N8141, N3133);
nand NAND2 (N8945, N8943, N8086);
nor NOR2 (N8946, N8944, N963);
or OR2 (N8947, N8939, N4008);
not NOT1 (N8948, N8942);
not NOT1 (N8949, N8947);
nor NOR3 (N8950, N8941, N487, N263);
and AND3 (N8951, N8929, N6036, N7585);
nand NAND2 (N8952, N8934, N8584);
or OR4 (N8953, N8948, N175, N3087, N8320);
nand NAND2 (N8954, N8905, N5466);
and AND2 (N8955, N8951, N1711);
not NOT1 (N8956, N8954);
nor NOR4 (N8957, N8949, N7779, N5182, N4660);
or OR4 (N8958, N8945, N2178, N5247, N3775);
nor NOR4 (N8959, N8952, N5913, N2333, N257);
nand NAND4 (N8960, N8950, N7379, N2725, N8216);
not NOT1 (N8961, N8960);
xor XOR2 (N8962, N8953, N7998);
nand NAND2 (N8963, N8962, N2359);
or OR4 (N8964, N8963, N215, N8139, N5419);
not NOT1 (N8965, N8964);
buf BUF1 (N8966, N8961);
nand NAND2 (N8967, N8958, N477);
or OR3 (N8968, N8955, N8516, N7009);
and AND2 (N8969, N8965, N607);
nand NAND3 (N8970, N8940, N4421, N4949);
buf BUF1 (N8971, N8966);
not NOT1 (N8972, N8957);
or OR3 (N8973, N8969, N6944, N6878);
nor NOR2 (N8974, N8973, N742);
not NOT1 (N8975, N8972);
nand NAND4 (N8976, N8975, N7548, N5526, N5874);
and AND3 (N8977, N8976, N1000, N6198);
xor XOR2 (N8978, N8930, N8756);
and AND3 (N8979, N8959, N7110, N7783);
xor XOR2 (N8980, N8956, N645);
xor XOR2 (N8981, N8968, N3540);
nand NAND2 (N8982, N8977, N6022);
nor NOR2 (N8983, N8970, N3638);
buf BUF1 (N8984, N8981);
xor XOR2 (N8985, N8982, N1363);
buf BUF1 (N8986, N8979);
buf BUF1 (N8987, N8967);
xor XOR2 (N8988, N8984, N7236);
nor NOR3 (N8989, N8987, N7841, N7761);
xor XOR2 (N8990, N8983, N3057);
or OR4 (N8991, N8978, N7256, N3792, N1854);
not NOT1 (N8992, N8991);
not NOT1 (N8993, N8971);
nand NAND2 (N8994, N8974, N7318);
and AND4 (N8995, N8946, N2103, N2838, N7381);
buf BUF1 (N8996, N8990);
and AND2 (N8997, N8995, N5358);
or OR2 (N8998, N8986, N8368);
or OR3 (N8999, N8992, N7586, N2934);
xor XOR2 (N9000, N8998, N8223);
nor NOR4 (N9001, N8996, N6822, N6996, N45);
nand NAND2 (N9002, N8988, N1379);
and AND2 (N9003, N8994, N5202);
buf BUF1 (N9004, N9000);
not NOT1 (N9005, N8993);
buf BUF1 (N9006, N9001);
nand NAND4 (N9007, N8989, N170, N8356, N512);
xor XOR2 (N9008, N9002, N7502);
not NOT1 (N9009, N9006);
and AND2 (N9010, N9004, N2026);
nor NOR4 (N9011, N9005, N2418, N2358, N7519);
buf BUF1 (N9012, N8999);
buf BUF1 (N9013, N9003);
buf BUF1 (N9014, N8980);
xor XOR2 (N9015, N9010, N6379);
nor NOR2 (N9016, N8985, N6355);
xor XOR2 (N9017, N9007, N3010);
or OR2 (N9018, N9014, N6604);
nand NAND3 (N9019, N9013, N8328, N6517);
nand NAND4 (N9020, N9019, N4683, N347, N7495);
or OR3 (N9021, N9008, N2770, N7875);
nand NAND4 (N9022, N9017, N4768, N2731, N5980);
or OR3 (N9023, N9009, N285, N7523);
or OR2 (N9024, N9011, N3911);
nand NAND4 (N9025, N8997, N801, N4641, N7354);
xor XOR2 (N9026, N9023, N2697);
buf BUF1 (N9027, N9012);
nor NOR4 (N9028, N9027, N2301, N7293, N6027);
nor NOR3 (N9029, N9022, N4435, N4147);
nor NOR3 (N9030, N9021, N7049, N1618);
and AND2 (N9031, N9029, N3053);
not NOT1 (N9032, N9024);
not NOT1 (N9033, N9015);
buf BUF1 (N9034, N9020);
nor NOR3 (N9035, N9016, N6795, N6421);
not NOT1 (N9036, N9028);
nand NAND2 (N9037, N9025, N6731);
and AND2 (N9038, N9032, N2324);
nor NOR3 (N9039, N9035, N3410, N8093);
nand NAND4 (N9040, N9033, N1589, N5004, N254);
and AND2 (N9041, N9034, N7693);
nand NAND3 (N9042, N9018, N7800, N3652);
xor XOR2 (N9043, N9041, N8563);
or OR2 (N9044, N9030, N3199);
xor XOR2 (N9045, N9036, N2870);
xor XOR2 (N9046, N9043, N2567);
or OR2 (N9047, N9038, N3855);
nor NOR4 (N9048, N9045, N7781, N7843, N8565);
nand NAND4 (N9049, N9042, N3764, N46, N4648);
nor NOR4 (N9050, N9026, N8982, N7084, N3641);
xor XOR2 (N9051, N9039, N3984);
and AND4 (N9052, N9047, N4409, N1617, N4920);
xor XOR2 (N9053, N9052, N5374);
buf BUF1 (N9054, N9051);
nor NOR2 (N9055, N9048, N8541);
buf BUF1 (N9056, N9044);
not NOT1 (N9057, N9055);
xor XOR2 (N9058, N9057, N2212);
xor XOR2 (N9059, N9056, N8359);
nand NAND3 (N9060, N9031, N8787, N2057);
nand NAND2 (N9061, N9040, N9029);
nand NAND2 (N9062, N9049, N2030);
and AND2 (N9063, N9046, N1545);
nand NAND3 (N9064, N9037, N1201, N4339);
or OR2 (N9065, N9062, N5488);
nand NAND4 (N9066, N9053, N7036, N1044, N5702);
and AND3 (N9067, N9050, N3857, N5259);
buf BUF1 (N9068, N9060);
xor XOR2 (N9069, N9067, N8256);
not NOT1 (N9070, N9063);
buf BUF1 (N9071, N9054);
not NOT1 (N9072, N9059);
xor XOR2 (N9073, N9068, N813);
or OR4 (N9074, N9070, N7415, N8093, N4636);
xor XOR2 (N9075, N9073, N2622);
and AND2 (N9076, N9069, N423);
xor XOR2 (N9077, N9061, N680);
not NOT1 (N9078, N9074);
and AND3 (N9079, N9075, N8826, N2987);
and AND2 (N9080, N9077, N7812);
and AND4 (N9081, N9072, N2458, N285, N7166);
and AND4 (N9082, N9065, N2995, N1358, N4491);
xor XOR2 (N9083, N9066, N5537);
buf BUF1 (N9084, N9078);
buf BUF1 (N9085, N9079);
nand NAND2 (N9086, N9085, N959);
buf BUF1 (N9087, N9086);
and AND4 (N9088, N9071, N7994, N3336, N3383);
nand NAND3 (N9089, N9076, N1917, N1911);
not NOT1 (N9090, N9082);
buf BUF1 (N9091, N9081);
buf BUF1 (N9092, N9089);
nand NAND2 (N9093, N9090, N8480);
buf BUF1 (N9094, N9084);
or OR3 (N9095, N9080, N7239, N5589);
nand NAND4 (N9096, N9087, N7033, N5651, N556);
xor XOR2 (N9097, N9091, N7867);
or OR4 (N9098, N9093, N7422, N4708, N6284);
or OR3 (N9099, N9096, N7877, N6829);
xor XOR2 (N9100, N9099, N2183);
not NOT1 (N9101, N9058);
nand NAND4 (N9102, N9094, N2864, N8170, N8407);
or OR2 (N9103, N9102, N3229);
not NOT1 (N9104, N9083);
nand NAND2 (N9105, N9103, N7613);
not NOT1 (N9106, N9101);
buf BUF1 (N9107, N9097);
xor XOR2 (N9108, N9095, N4605);
xor XOR2 (N9109, N9092, N6042);
xor XOR2 (N9110, N9100, N373);
xor XOR2 (N9111, N9109, N6941);
nand NAND3 (N9112, N9106, N5062, N6998);
and AND3 (N9113, N9108, N2822, N5182);
nor NOR3 (N9114, N9104, N4169, N6352);
buf BUF1 (N9115, N9107);
nand NAND3 (N9116, N9111, N4935, N2772);
buf BUF1 (N9117, N9112);
nand NAND4 (N9118, N9114, N10, N2133, N8511);
buf BUF1 (N9119, N9098);
buf BUF1 (N9120, N9113);
and AND3 (N9121, N9118, N5212, N3131);
and AND3 (N9122, N9110, N4807, N6459);
not NOT1 (N9123, N9119);
nand NAND3 (N9124, N9064, N3600, N8798);
not NOT1 (N9125, N9123);
xor XOR2 (N9126, N9115, N6757);
xor XOR2 (N9127, N9121, N5721);
or OR3 (N9128, N9120, N2113, N5255);
nand NAND2 (N9129, N9125, N4499);
xor XOR2 (N9130, N9128, N4554);
xor XOR2 (N9131, N9116, N609);
or OR4 (N9132, N9124, N7342, N2955, N8831);
and AND3 (N9133, N9130, N4776, N3693);
not NOT1 (N9134, N9127);
buf BUF1 (N9135, N9131);
nor NOR4 (N9136, N9133, N2450, N6978, N3730);
xor XOR2 (N9137, N9129, N6413);
nor NOR2 (N9138, N9117, N3512);
nand NAND3 (N9139, N9122, N2090, N5154);
nor NOR2 (N9140, N9132, N2331);
nor NOR4 (N9141, N9126, N7997, N329, N3896);
nand NAND4 (N9142, N9134, N6512, N8035, N3564);
buf BUF1 (N9143, N9135);
or OR3 (N9144, N9139, N7529, N1861);
nand NAND2 (N9145, N9143, N4460);
and AND3 (N9146, N9137, N7718, N7291);
and AND2 (N9147, N9145, N4195);
not NOT1 (N9148, N9147);
xor XOR2 (N9149, N9105, N7080);
nor NOR3 (N9150, N9088, N6580, N8615);
or OR3 (N9151, N9141, N3653, N8465);
and AND3 (N9152, N9140, N8648, N5661);
nand NAND3 (N9153, N9151, N5193, N1522);
not NOT1 (N9154, N9149);
xor XOR2 (N9155, N9148, N5723);
nor NOR4 (N9156, N9146, N377, N4477, N6029);
or OR4 (N9157, N9156, N1202, N1099, N406);
and AND3 (N9158, N9136, N127, N3639);
or OR2 (N9159, N9154, N1276);
nand NAND3 (N9160, N9144, N3278, N1216);
buf BUF1 (N9161, N9160);
or OR4 (N9162, N9155, N8630, N7587, N9043);
or OR2 (N9163, N9152, N6309);
and AND3 (N9164, N9159, N5423, N4192);
buf BUF1 (N9165, N9161);
not NOT1 (N9166, N9142);
nor NOR4 (N9167, N9165, N43, N4908, N7559);
and AND4 (N9168, N9157, N2052, N3968, N542);
not NOT1 (N9169, N9164);
nand NAND2 (N9170, N9169, N7735);
nor NOR4 (N9171, N9150, N5414, N263, N8609);
nand NAND2 (N9172, N9171, N8925);
nand NAND3 (N9173, N9170, N5379, N8055);
and AND3 (N9174, N9138, N1100, N1518);
or OR2 (N9175, N9174, N5460);
or OR2 (N9176, N9158, N7544);
or OR4 (N9177, N9176, N7988, N7743, N4392);
nor NOR4 (N9178, N9163, N1644, N5756, N5694);
and AND4 (N9179, N9167, N5621, N7403, N6660);
nor NOR3 (N9180, N9178, N2213, N7413);
nor NOR4 (N9181, N9173, N3233, N3689, N5002);
buf BUF1 (N9182, N9166);
buf BUF1 (N9183, N9168);
nand NAND4 (N9184, N9183, N6432, N615, N147);
nor NOR4 (N9185, N9181, N3016, N1355, N9005);
xor XOR2 (N9186, N9177, N8279);
or OR3 (N9187, N9184, N8559, N6495);
buf BUF1 (N9188, N9185);
xor XOR2 (N9189, N9182, N831);
nor NOR4 (N9190, N9162, N4782, N7056, N2119);
buf BUF1 (N9191, N9189);
or OR3 (N9192, N9191, N3273, N845);
and AND4 (N9193, N9190, N7281, N8695, N611);
buf BUF1 (N9194, N9180);
xor XOR2 (N9195, N9187, N489);
xor XOR2 (N9196, N9195, N8673);
or OR4 (N9197, N9194, N2899, N1935, N8356);
nor NOR4 (N9198, N9179, N9004, N2306, N918);
or OR3 (N9199, N9172, N8369, N6842);
nor NOR4 (N9200, N9175, N4083, N7737, N6399);
xor XOR2 (N9201, N9188, N7233);
nand NAND3 (N9202, N9186, N4459, N6356);
and AND3 (N9203, N9153, N8276, N476);
buf BUF1 (N9204, N9198);
or OR2 (N9205, N9203, N8675);
and AND3 (N9206, N9204, N8842, N2889);
not NOT1 (N9207, N9193);
nor NOR3 (N9208, N9196, N2181, N4151);
or OR2 (N9209, N9192, N8586);
or OR4 (N9210, N9207, N2416, N2271, N7383);
not NOT1 (N9211, N9202);
nor NOR3 (N9212, N9209, N7961, N4827);
or OR3 (N9213, N9199, N8036, N1983);
xor XOR2 (N9214, N9210, N6975);
buf BUF1 (N9215, N9212);
or OR4 (N9216, N9211, N7373, N727, N7467);
and AND4 (N9217, N9214, N5272, N8521, N3161);
nand NAND3 (N9218, N9201, N585, N1877);
not NOT1 (N9219, N9208);
nor NOR4 (N9220, N9205, N7456, N7797, N4911);
and AND4 (N9221, N9200, N7791, N6218, N3929);
not NOT1 (N9222, N9219);
not NOT1 (N9223, N9221);
xor XOR2 (N9224, N9223, N7506);
and AND4 (N9225, N9213, N3733, N3280, N6587);
nor NOR4 (N9226, N9215, N5493, N4789, N5434);
and AND4 (N9227, N9224, N6732, N4602, N2234);
nand NAND4 (N9228, N9225, N1600, N1236, N3739);
buf BUF1 (N9229, N9222);
xor XOR2 (N9230, N9216, N7940);
and AND4 (N9231, N9206, N1847, N7918, N3111);
buf BUF1 (N9232, N9218);
nor NOR4 (N9233, N9217, N6149, N5422, N6352);
buf BUF1 (N9234, N9230);
nor NOR4 (N9235, N9197, N83, N7489, N1935);
not NOT1 (N9236, N9234);
and AND4 (N9237, N9235, N1965, N2082, N3946);
buf BUF1 (N9238, N9237);
nor NOR4 (N9239, N9232, N7713, N8927, N7225);
and AND2 (N9240, N9233, N1967);
nor NOR4 (N9241, N9236, N6044, N1659, N5824);
buf BUF1 (N9242, N9227);
or OR2 (N9243, N9238, N5064);
nor NOR4 (N9244, N9240, N8724, N7308, N2317);
buf BUF1 (N9245, N9220);
xor XOR2 (N9246, N9245, N1000);
or OR2 (N9247, N9231, N5932);
xor XOR2 (N9248, N9246, N1791);
not NOT1 (N9249, N9247);
not NOT1 (N9250, N9239);
or OR4 (N9251, N9226, N1283, N314, N6358);
buf BUF1 (N9252, N9244);
and AND3 (N9253, N9243, N5107, N5259);
xor XOR2 (N9254, N9248, N6571);
nand NAND3 (N9255, N9228, N691, N4132);
not NOT1 (N9256, N9250);
or OR2 (N9257, N9252, N3579);
xor XOR2 (N9258, N9256, N1020);
and AND3 (N9259, N9255, N7117, N5256);
buf BUF1 (N9260, N9249);
nor NOR2 (N9261, N9254, N6835);
or OR2 (N9262, N9251, N7396);
and AND2 (N9263, N9262, N7196);
and AND4 (N9264, N9257, N6655, N387, N9232);
and AND3 (N9265, N9253, N6498, N2989);
or OR4 (N9266, N9229, N4837, N8120, N3059);
nor NOR2 (N9267, N9266, N143);
or OR3 (N9268, N9242, N1895, N685);
and AND2 (N9269, N9258, N6121);
nand NAND2 (N9270, N9264, N3383);
xor XOR2 (N9271, N9268, N147);
buf BUF1 (N9272, N9260);
xor XOR2 (N9273, N9271, N1759);
and AND4 (N9274, N9241, N4698, N3816, N6505);
nor NOR4 (N9275, N9274, N4622, N6088, N7272);
xor XOR2 (N9276, N9270, N1742);
nor NOR2 (N9277, N9267, N3646);
or OR4 (N9278, N9273, N2953, N8712, N7020);
not NOT1 (N9279, N9263);
and AND4 (N9280, N9277, N4857, N7971, N656);
nand NAND4 (N9281, N9259, N4549, N5110, N7919);
and AND3 (N9282, N9265, N8108, N8762);
and AND4 (N9283, N9275, N4658, N5559, N5526);
nand NAND3 (N9284, N9276, N8857, N3649);
buf BUF1 (N9285, N9280);
and AND4 (N9286, N9261, N4920, N2545, N6334);
and AND4 (N9287, N9272, N3972, N5839, N3078);
or OR2 (N9288, N9282, N334);
or OR4 (N9289, N9283, N94, N8913, N4433);
and AND4 (N9290, N9288, N6713, N5558, N7277);
buf BUF1 (N9291, N9285);
nand NAND3 (N9292, N9269, N73, N7292);
nand NAND4 (N9293, N9278, N1257, N3763, N95);
nor NOR2 (N9294, N9284, N2120);
xor XOR2 (N9295, N9287, N952);
or OR2 (N9296, N9279, N612);
nand NAND3 (N9297, N9291, N5661, N4733);
nand NAND3 (N9298, N9296, N7178, N6021);
or OR4 (N9299, N9293, N3578, N1051, N5243);
xor XOR2 (N9300, N9299, N4399);
buf BUF1 (N9301, N9294);
nand NAND4 (N9302, N9300, N7531, N9156, N5584);
nand NAND2 (N9303, N9302, N8971);
nor NOR4 (N9304, N9303, N3886, N8374, N8657);
or OR2 (N9305, N9289, N265);
or OR4 (N9306, N9290, N88, N6878, N186);
nand NAND2 (N9307, N9286, N6784);
and AND2 (N9308, N9281, N6742);
not NOT1 (N9309, N9308);
and AND3 (N9310, N9304, N6445, N4869);
not NOT1 (N9311, N9309);
nand NAND2 (N9312, N9307, N809);
and AND3 (N9313, N9312, N6145, N4260);
nand NAND4 (N9314, N9292, N167, N4852, N8834);
and AND3 (N9315, N9298, N462, N5214);
not NOT1 (N9316, N9295);
nand NAND3 (N9317, N9316, N4771, N3425);
buf BUF1 (N9318, N9317);
buf BUF1 (N9319, N9314);
nand NAND2 (N9320, N9297, N7778);
xor XOR2 (N9321, N9306, N6326);
not NOT1 (N9322, N9321);
nor NOR2 (N9323, N9318, N1405);
and AND4 (N9324, N9311, N6573, N5866, N9040);
or OR2 (N9325, N9313, N4443);
nand NAND4 (N9326, N9323, N2666, N4983, N2385);
nor NOR2 (N9327, N9319, N992);
not NOT1 (N9328, N9305);
nand NAND4 (N9329, N9301, N5558, N6299, N1341);
not NOT1 (N9330, N9326);
buf BUF1 (N9331, N9329);
nand NAND2 (N9332, N9324, N3358);
xor XOR2 (N9333, N9331, N5333);
nor NOR3 (N9334, N9320, N7857, N5652);
or OR3 (N9335, N9310, N2812, N6774);
not NOT1 (N9336, N9332);
nand NAND3 (N9337, N9334, N2658, N7564);
or OR3 (N9338, N9336, N3101, N8993);
or OR3 (N9339, N9337, N5537, N704);
nor NOR3 (N9340, N9339, N7824, N4500);
not NOT1 (N9341, N9315);
nor NOR4 (N9342, N9330, N8600, N3813, N1391);
buf BUF1 (N9343, N9328);
nor NOR2 (N9344, N9343, N5564);
nor NOR2 (N9345, N9342, N5355);
not NOT1 (N9346, N9338);
nor NOR4 (N9347, N9335, N3758, N5254, N5889);
xor XOR2 (N9348, N9325, N7743);
buf BUF1 (N9349, N9333);
and AND2 (N9350, N9346, N4593);
nor NOR2 (N9351, N9340, N4469);
nor NOR2 (N9352, N9327, N1004);
not NOT1 (N9353, N9350);
xor XOR2 (N9354, N9349, N7250);
not NOT1 (N9355, N9344);
nor NOR2 (N9356, N9345, N5961);
xor XOR2 (N9357, N9322, N155);
and AND2 (N9358, N9357, N3501);
xor XOR2 (N9359, N9351, N7086);
not NOT1 (N9360, N9352);
nor NOR2 (N9361, N9341, N7836);
or OR2 (N9362, N9358, N1196);
or OR2 (N9363, N9347, N8645);
buf BUF1 (N9364, N9361);
nand NAND3 (N9365, N9354, N2574, N2626);
or OR3 (N9366, N9365, N5742, N7554);
or OR4 (N9367, N9363, N5169, N2288, N40);
xor XOR2 (N9368, N9348, N1361);
nand NAND2 (N9369, N9355, N8571);
nand NAND4 (N9370, N9367, N2378, N8267, N3124);
buf BUF1 (N9371, N9353);
nor NOR3 (N9372, N9359, N3189, N4940);
nor NOR2 (N9373, N9372, N7608);
and AND3 (N9374, N9364, N6010, N8915);
not NOT1 (N9375, N9368);
nor NOR4 (N9376, N9373, N1942, N5677, N8793);
buf BUF1 (N9377, N9374);
nor NOR4 (N9378, N9376, N2000, N3653, N1769);
or OR2 (N9379, N9371, N6714);
nor NOR4 (N9380, N9356, N4688, N9131, N3496);
and AND2 (N9381, N9360, N3419);
not NOT1 (N9382, N9369);
and AND2 (N9383, N9381, N4195);
not NOT1 (N9384, N9378);
or OR3 (N9385, N9362, N5657, N3825);
buf BUF1 (N9386, N9377);
or OR2 (N9387, N9384, N9340);
and AND2 (N9388, N9386, N4085);
nand NAND4 (N9389, N9385, N2730, N6267, N4991);
buf BUF1 (N9390, N9380);
nand NAND2 (N9391, N9370, N625);
not NOT1 (N9392, N9366);
or OR4 (N9393, N9389, N9369, N3315, N1054);
not NOT1 (N9394, N9387);
and AND4 (N9395, N9391, N6029, N4841, N8059);
and AND2 (N9396, N9393, N4249);
xor XOR2 (N9397, N9395, N5311);
not NOT1 (N9398, N9394);
and AND4 (N9399, N9375, N4371, N8012, N7422);
or OR3 (N9400, N9390, N4908, N3759);
xor XOR2 (N9401, N9383, N6043);
nor NOR3 (N9402, N9401, N6000, N8081);
not NOT1 (N9403, N9397);
or OR3 (N9404, N9382, N6903, N181);
buf BUF1 (N9405, N9399);
xor XOR2 (N9406, N9379, N1577);
nand NAND3 (N9407, N9402, N7166, N5963);
not NOT1 (N9408, N9392);
not NOT1 (N9409, N9403);
xor XOR2 (N9410, N9405, N2837);
buf BUF1 (N9411, N9410);
or OR4 (N9412, N9407, N1775, N5095, N3483);
or OR3 (N9413, N9400, N8055, N4609);
not NOT1 (N9414, N9408);
nand NAND3 (N9415, N9398, N7809, N3933);
not NOT1 (N9416, N9406);
buf BUF1 (N9417, N9409);
and AND4 (N9418, N9404, N8211, N488, N1195);
nand NAND4 (N9419, N9413, N7838, N4595, N3068);
or OR4 (N9420, N9412, N2046, N5324, N8376);
xor XOR2 (N9421, N9418, N3336);
xor XOR2 (N9422, N9414, N4154);
or OR4 (N9423, N9419, N1017, N1520, N76);
and AND4 (N9424, N9416, N2338, N7109, N1849);
nor NOR3 (N9425, N9411, N4505, N4150);
buf BUF1 (N9426, N9422);
not NOT1 (N9427, N9421);
and AND4 (N9428, N9426, N895, N5696, N5448);
not NOT1 (N9429, N9396);
nand NAND3 (N9430, N9428, N150, N616);
nand NAND3 (N9431, N9425, N9350, N4792);
and AND4 (N9432, N9430, N3188, N8863, N8529);
not NOT1 (N9433, N9432);
not NOT1 (N9434, N9433);
nor NOR2 (N9435, N9424, N1033);
and AND2 (N9436, N9427, N8316);
nand NAND2 (N9437, N9417, N7066);
not NOT1 (N9438, N9415);
xor XOR2 (N9439, N9420, N1214);
not NOT1 (N9440, N9436);
and AND2 (N9441, N9423, N9226);
buf BUF1 (N9442, N9388);
buf BUF1 (N9443, N9435);
nor NOR2 (N9444, N9438, N6286);
xor XOR2 (N9445, N9437, N4763);
and AND4 (N9446, N9434, N938, N9414, N3634);
or OR2 (N9447, N9444, N4719);
nand NAND2 (N9448, N9442, N862);
nor NOR3 (N9449, N9441, N2864, N5097);
nand NAND2 (N9450, N9429, N6667);
and AND2 (N9451, N9440, N7246);
xor XOR2 (N9452, N9447, N1297);
nand NAND4 (N9453, N9451, N475, N2897, N5777);
xor XOR2 (N9454, N9448, N1307);
not NOT1 (N9455, N9450);
buf BUF1 (N9456, N9455);
not NOT1 (N9457, N9453);
and AND2 (N9458, N9456, N3489);
and AND3 (N9459, N9439, N4598, N5594);
or OR4 (N9460, N9446, N5764, N6661, N5893);
not NOT1 (N9461, N9460);
buf BUF1 (N9462, N9431);
not NOT1 (N9463, N9461);
xor XOR2 (N9464, N9452, N1572);
buf BUF1 (N9465, N9457);
nand NAND4 (N9466, N9454, N4901, N3229, N8408);
nand NAND2 (N9467, N9466, N4552);
nor NOR3 (N9468, N9459, N5356, N4869);
xor XOR2 (N9469, N9463, N4348);
xor XOR2 (N9470, N9462, N2283);
and AND4 (N9471, N9445, N7268, N1723, N2828);
nor NOR4 (N9472, N9449, N3748, N9317, N2011);
xor XOR2 (N9473, N9458, N3660);
nor NOR3 (N9474, N9465, N1679, N5788);
nand NAND4 (N9475, N9468, N6531, N301, N7515);
nand NAND4 (N9476, N9467, N6595, N1580, N7401);
not NOT1 (N9477, N9470);
not NOT1 (N9478, N9473);
or OR3 (N9479, N9443, N5174, N6717);
not NOT1 (N9480, N9464);
xor XOR2 (N9481, N9477, N520);
and AND4 (N9482, N9469, N5074, N9176, N4025);
not NOT1 (N9483, N9482);
nor NOR3 (N9484, N9478, N530, N6398);
nand NAND2 (N9485, N9480, N7310);
xor XOR2 (N9486, N9475, N3528);
not NOT1 (N9487, N9484);
nand NAND2 (N9488, N9483, N3648);
or OR3 (N9489, N9488, N6046, N561);
and AND4 (N9490, N9489, N4223, N7293, N5913);
and AND4 (N9491, N9487, N4763, N1681, N2250);
nand NAND4 (N9492, N9485, N8866, N1775, N1077);
or OR3 (N9493, N9481, N6677, N6578);
xor XOR2 (N9494, N9479, N6190);
nor NOR4 (N9495, N9491, N5427, N830, N5367);
or OR4 (N9496, N9495, N7344, N4365, N8557);
buf BUF1 (N9497, N9474);
xor XOR2 (N9498, N9490, N3310);
buf BUF1 (N9499, N9471);
and AND4 (N9500, N9496, N5040, N6680, N8165);
nor NOR2 (N9501, N9494, N371);
nand NAND2 (N9502, N9492, N1887);
nor NOR4 (N9503, N9502, N2071, N1412, N4499);
and AND2 (N9504, N9499, N6361);
and AND3 (N9505, N9476, N9317, N8991);
buf BUF1 (N9506, N9498);
nor NOR3 (N9507, N9486, N5444, N6151);
buf BUF1 (N9508, N9500);
or OR4 (N9509, N9506, N490, N8100, N5874);
or OR2 (N9510, N9504, N5172);
and AND2 (N9511, N9505, N9026);
and AND3 (N9512, N9509, N969, N2897);
xor XOR2 (N9513, N9508, N6182);
nor NOR4 (N9514, N9513, N5983, N7883, N6835);
not NOT1 (N9515, N9472);
and AND4 (N9516, N9493, N794, N6862, N9092);
not NOT1 (N9517, N9511);
nor NOR4 (N9518, N9497, N6636, N2479, N7367);
nand NAND4 (N9519, N9517, N6212, N1014, N5155);
nor NOR3 (N9520, N9518, N2804, N6383);
nor NOR4 (N9521, N9512, N7782, N7865, N341);
and AND3 (N9522, N9514, N6145, N7829);
xor XOR2 (N9523, N9510, N4964);
xor XOR2 (N9524, N9519, N6489);
xor XOR2 (N9525, N9522, N3543);
not NOT1 (N9526, N9520);
nor NOR3 (N9527, N9503, N8374, N8114);
not NOT1 (N9528, N9527);
buf BUF1 (N9529, N9523);
and AND2 (N9530, N9524, N6555);
and AND4 (N9531, N9507, N9231, N7347, N3872);
buf BUF1 (N9532, N9529);
nand NAND2 (N9533, N9515, N5946);
and AND2 (N9534, N9532, N3586);
or OR3 (N9535, N9531, N4777, N140);
nand NAND3 (N9536, N9525, N9049, N7537);
and AND4 (N9537, N9535, N7642, N1514, N5684);
or OR3 (N9538, N9526, N8791, N3940);
nor NOR4 (N9539, N9528, N4800, N4439, N8804);
buf BUF1 (N9540, N9538);
not NOT1 (N9541, N9516);
and AND4 (N9542, N9533, N48, N4406, N2414);
and AND4 (N9543, N9521, N6939, N61, N4773);
and AND4 (N9544, N9501, N5695, N8110, N6196);
nor NOR3 (N9545, N9541, N5398, N364);
buf BUF1 (N9546, N9537);
or OR2 (N9547, N9542, N5482);
nor NOR3 (N9548, N9545, N578, N824);
and AND2 (N9549, N9546, N4707);
nand NAND4 (N9550, N9544, N4475, N2810, N2515);
not NOT1 (N9551, N9549);
or OR3 (N9552, N9530, N2823, N7268);
nor NOR4 (N9553, N9548, N971, N5085, N1432);
or OR4 (N9554, N9534, N1633, N4133, N320);
and AND3 (N9555, N9539, N1762, N1812);
nand NAND4 (N9556, N9551, N4152, N7880, N7419);
buf BUF1 (N9557, N9540);
and AND3 (N9558, N9557, N8472, N2316);
and AND3 (N9559, N9554, N8820, N2205);
xor XOR2 (N9560, N9536, N6447);
nor NOR2 (N9561, N9560, N40);
nor NOR3 (N9562, N9553, N3519, N2511);
and AND4 (N9563, N9556, N8766, N1776, N1129);
or OR2 (N9564, N9563, N846);
buf BUF1 (N9565, N9550);
nor NOR3 (N9566, N9561, N7594, N8680);
nand NAND2 (N9567, N9543, N5057);
or OR2 (N9568, N9562, N7824);
buf BUF1 (N9569, N9558);
not NOT1 (N9570, N9552);
nor NOR4 (N9571, N9547, N4129, N6629, N7252);
nand NAND2 (N9572, N9555, N1959);
and AND2 (N9573, N9565, N1605);
and AND4 (N9574, N9572, N4020, N3066, N4025);
not NOT1 (N9575, N9569);
xor XOR2 (N9576, N9567, N6893);
or OR4 (N9577, N9576, N133, N5308, N1819);
and AND3 (N9578, N9566, N9218, N9338);
not NOT1 (N9579, N9568);
nand NAND3 (N9580, N9579, N1879, N3610);
or OR3 (N9581, N9571, N7637, N84);
or OR4 (N9582, N9578, N5024, N3681, N6954);
not NOT1 (N9583, N9580);
not NOT1 (N9584, N9582);
nor NOR3 (N9585, N9583, N1914, N1842);
xor XOR2 (N9586, N9575, N2883);
not NOT1 (N9587, N9570);
xor XOR2 (N9588, N9577, N3350);
buf BUF1 (N9589, N9587);
or OR4 (N9590, N9581, N5612, N6793, N8276);
nand NAND3 (N9591, N9573, N3625, N2229);
or OR2 (N9592, N9589, N7419);
nand NAND4 (N9593, N9584, N6623, N99, N4867);
buf BUF1 (N9594, N9564);
or OR4 (N9595, N9586, N8564, N1197, N1996);
and AND2 (N9596, N9574, N7599);
and AND2 (N9597, N9585, N2260);
nor NOR4 (N9598, N9597, N4505, N9053, N8876);
and AND3 (N9599, N9590, N5567, N9101);
xor XOR2 (N9600, N9599, N6647);
nand NAND3 (N9601, N9593, N1053, N3615);
and AND2 (N9602, N9598, N9090);
or OR2 (N9603, N9594, N5554);
buf BUF1 (N9604, N9592);
not NOT1 (N9605, N9604);
not NOT1 (N9606, N9600);
xor XOR2 (N9607, N9602, N1068);
or OR4 (N9608, N9559, N6704, N1847, N4948);
not NOT1 (N9609, N9601);
and AND2 (N9610, N9588, N6962);
nand NAND2 (N9611, N9605, N541);
xor XOR2 (N9612, N9611, N1143);
not NOT1 (N9613, N9609);
and AND2 (N9614, N9613, N9116);
xor XOR2 (N9615, N9595, N8254);
and AND3 (N9616, N9614, N3872, N1683);
xor XOR2 (N9617, N9606, N1304);
xor XOR2 (N9618, N9591, N1989);
not NOT1 (N9619, N9607);
not NOT1 (N9620, N9615);
buf BUF1 (N9621, N9616);
xor XOR2 (N9622, N9618, N6769);
buf BUF1 (N9623, N9608);
and AND4 (N9624, N9610, N2992, N3429, N8468);
nor NOR4 (N9625, N9596, N7091, N7040, N4118);
and AND4 (N9626, N9624, N6268, N2987, N9316);
nand NAND4 (N9627, N9619, N7488, N2875, N4217);
xor XOR2 (N9628, N9621, N6882);
nand NAND2 (N9629, N9626, N3090);
not NOT1 (N9630, N9620);
not NOT1 (N9631, N9623);
and AND2 (N9632, N9622, N227);
buf BUF1 (N9633, N9629);
nor NOR2 (N9634, N9631, N4253);
or OR3 (N9635, N9625, N2565, N6158);
or OR3 (N9636, N9627, N420, N541);
buf BUF1 (N9637, N9630);
nand NAND3 (N9638, N9603, N4341, N8821);
or OR3 (N9639, N9636, N4443, N1607);
or OR4 (N9640, N9635, N8632, N2692, N682);
and AND2 (N9641, N9628, N5808);
or OR4 (N9642, N9632, N7188, N438, N6663);
not NOT1 (N9643, N9617);
and AND2 (N9644, N9634, N8066);
not NOT1 (N9645, N9637);
buf BUF1 (N9646, N9644);
buf BUF1 (N9647, N9643);
nor NOR4 (N9648, N9642, N4391, N2649, N7435);
and AND2 (N9649, N9647, N4854);
nand NAND3 (N9650, N9633, N8778, N6287);
and AND3 (N9651, N9612, N8555, N7174);
nand NAND3 (N9652, N9650, N8133, N9590);
nand NAND2 (N9653, N9651, N4350);
nand NAND4 (N9654, N9648, N7976, N2923, N8238);
and AND4 (N9655, N9641, N8430, N552, N4012);
or OR3 (N9656, N9638, N4736, N4212);
nand NAND3 (N9657, N9655, N6919, N3008);
buf BUF1 (N9658, N9653);
and AND2 (N9659, N9658, N2768);
nor NOR4 (N9660, N9659, N2289, N2109, N2987);
nor NOR4 (N9661, N9656, N3291, N5872, N8479);
not NOT1 (N9662, N9646);
nand NAND3 (N9663, N9660, N6727, N6349);
or OR4 (N9664, N9639, N6903, N3821, N1033);
nand NAND4 (N9665, N9649, N7602, N7031, N1297);
nand NAND2 (N9666, N9640, N4261);
nand NAND4 (N9667, N9662, N382, N3851, N1121);
and AND3 (N9668, N9663, N4642, N6262);
xor XOR2 (N9669, N9666, N4534);
not NOT1 (N9670, N9645);
not NOT1 (N9671, N9669);
nand NAND3 (N9672, N9664, N1808, N4597);
nand NAND4 (N9673, N9654, N5908, N6970, N8191);
or OR2 (N9674, N9667, N6378);
nor NOR4 (N9675, N9657, N775, N1751, N4753);
and AND2 (N9676, N9673, N7491);
not NOT1 (N9677, N9652);
xor XOR2 (N9678, N9672, N6980);
and AND3 (N9679, N9677, N9622, N9042);
buf BUF1 (N9680, N9678);
nand NAND2 (N9681, N9680, N2015);
xor XOR2 (N9682, N9668, N5392);
xor XOR2 (N9683, N9671, N6157);
buf BUF1 (N9684, N9675);
and AND2 (N9685, N9676, N6191);
not NOT1 (N9686, N9683);
xor XOR2 (N9687, N9674, N7941);
not NOT1 (N9688, N9670);
or OR3 (N9689, N9684, N7122, N4687);
nand NAND3 (N9690, N9689, N2336, N2133);
nand NAND2 (N9691, N9679, N2271);
nand NAND4 (N9692, N9682, N6070, N4298, N3163);
and AND2 (N9693, N9661, N2281);
nand NAND2 (N9694, N9687, N7066);
nor NOR4 (N9695, N9694, N8404, N6866, N4025);
not NOT1 (N9696, N9665);
and AND4 (N9697, N9686, N3569, N1228, N9383);
or OR4 (N9698, N9692, N1052, N1367, N4134);
nand NAND3 (N9699, N9693, N2727, N5878);
nand NAND4 (N9700, N9698, N9628, N465, N5944);
nor NOR4 (N9701, N9688, N6846, N2212, N894);
buf BUF1 (N9702, N9699);
nor NOR3 (N9703, N9701, N7291, N6177);
or OR2 (N9704, N9697, N5274);
nor NOR3 (N9705, N9702, N3447, N4040);
nand NAND3 (N9706, N9696, N6814, N8238);
xor XOR2 (N9707, N9703, N7908);
nor NOR2 (N9708, N9685, N7269);
nor NOR2 (N9709, N9705, N2339);
or OR2 (N9710, N9681, N4676);
and AND3 (N9711, N9708, N2535, N2240);
xor XOR2 (N9712, N9695, N8622);
or OR4 (N9713, N9706, N1906, N2356, N3656);
nand NAND3 (N9714, N9709, N7694, N1612);
buf BUF1 (N9715, N9711);
or OR3 (N9716, N9707, N3821, N1242);
nand NAND4 (N9717, N9710, N820, N9142, N3474);
and AND2 (N9718, N9704, N7236);
and AND3 (N9719, N9717, N1115, N2705);
buf BUF1 (N9720, N9712);
not NOT1 (N9721, N9690);
buf BUF1 (N9722, N9719);
and AND3 (N9723, N9700, N2746, N1934);
nor NOR3 (N9724, N9722, N8281, N9639);
or OR3 (N9725, N9691, N3882, N5915);
buf BUF1 (N9726, N9713);
nor NOR4 (N9727, N9716, N1217, N4480, N2242);
and AND4 (N9728, N9724, N7209, N8281, N8621);
or OR3 (N9729, N9725, N3277, N7663);
xor XOR2 (N9730, N9727, N8186);
xor XOR2 (N9731, N9723, N8825);
xor XOR2 (N9732, N9721, N9639);
nor NOR3 (N9733, N9714, N2239, N3443);
not NOT1 (N9734, N9718);
nor NOR3 (N9735, N9732, N1319, N3307);
or OR3 (N9736, N9720, N7155, N8823);
buf BUF1 (N9737, N9728);
xor XOR2 (N9738, N9729, N5998);
or OR3 (N9739, N9736, N509, N9155);
or OR4 (N9740, N9737, N3097, N9173, N2009);
and AND4 (N9741, N9738, N3985, N7573, N4568);
not NOT1 (N9742, N9741);
buf BUF1 (N9743, N9742);
nand NAND2 (N9744, N9730, N6018);
and AND4 (N9745, N9715, N1924, N8807, N601);
and AND3 (N9746, N9745, N8453, N9742);
or OR3 (N9747, N9740, N8044, N8627);
buf BUF1 (N9748, N9746);
nor NOR2 (N9749, N9733, N6147);
buf BUF1 (N9750, N9749);
nand NAND2 (N9751, N9747, N3645);
or OR2 (N9752, N9748, N1284);
nand NAND2 (N9753, N9731, N1474);
xor XOR2 (N9754, N9734, N2527);
or OR3 (N9755, N9744, N2969, N7468);
or OR4 (N9756, N9753, N5939, N5666, N9199);
and AND2 (N9757, N9726, N6633);
and AND3 (N9758, N9750, N999, N9153);
or OR3 (N9759, N9752, N1953, N5764);
and AND2 (N9760, N9758, N3885);
nor NOR2 (N9761, N9759, N3189);
or OR4 (N9762, N9735, N5981, N2407, N4953);
not NOT1 (N9763, N9743);
not NOT1 (N9764, N9754);
xor XOR2 (N9765, N9757, N5328);
and AND4 (N9766, N9762, N9534, N5353, N9269);
buf BUF1 (N9767, N9761);
xor XOR2 (N9768, N9765, N4878);
not NOT1 (N9769, N9760);
or OR3 (N9770, N9739, N7321, N5935);
xor XOR2 (N9771, N9769, N4486);
xor XOR2 (N9772, N9770, N7891);
nor NOR4 (N9773, N9763, N8868, N8455, N1171);
or OR4 (N9774, N9764, N8195, N6164, N2992);
nand NAND2 (N9775, N9766, N3187);
buf BUF1 (N9776, N9755);
nor NOR2 (N9777, N9771, N9096);
xor XOR2 (N9778, N9768, N4304);
buf BUF1 (N9779, N9756);
and AND2 (N9780, N9779, N9333);
xor XOR2 (N9781, N9778, N9440);
not NOT1 (N9782, N9776);
not NOT1 (N9783, N9780);
or OR2 (N9784, N9782, N7071);
or OR4 (N9785, N9783, N2766, N8392, N7772);
nand NAND4 (N9786, N9772, N5516, N6879, N7329);
buf BUF1 (N9787, N9775);
not NOT1 (N9788, N9774);
xor XOR2 (N9789, N9751, N8966);
buf BUF1 (N9790, N9788);
nor NOR2 (N9791, N9789, N514);
not NOT1 (N9792, N9781);
xor XOR2 (N9793, N9790, N9092);
or OR4 (N9794, N9777, N9644, N399, N3572);
xor XOR2 (N9795, N9784, N124);
and AND4 (N9796, N9794, N6602, N9396, N8422);
nor NOR4 (N9797, N9773, N6395, N7293, N278);
nand NAND3 (N9798, N9796, N6482, N6752);
and AND2 (N9799, N9792, N6144);
xor XOR2 (N9800, N9798, N5096);
nor NOR4 (N9801, N9793, N8334, N6767, N7328);
or OR3 (N9802, N9791, N6491, N6379);
nand NAND4 (N9803, N9795, N750, N6143, N2763);
nand NAND4 (N9804, N9801, N934, N8261, N819);
buf BUF1 (N9805, N9802);
or OR3 (N9806, N9805, N8148, N5330);
xor XOR2 (N9807, N9787, N3747);
nand NAND3 (N9808, N9767, N6037, N4112);
xor XOR2 (N9809, N9804, N2140);
buf BUF1 (N9810, N9786);
or OR3 (N9811, N9803, N3454, N2108);
xor XOR2 (N9812, N9808, N9012);
not NOT1 (N9813, N9809);
nand NAND4 (N9814, N9807, N2557, N9345, N4058);
nor NOR2 (N9815, N9814, N3588);
or OR4 (N9816, N9800, N4883, N8488, N2895);
nor NOR3 (N9817, N9806, N6355, N743);
and AND4 (N9818, N9797, N6884, N4728, N8860);
xor XOR2 (N9819, N9818, N7230);
and AND2 (N9820, N9815, N7101);
nand NAND2 (N9821, N9816, N5460);
xor XOR2 (N9822, N9810, N1491);
buf BUF1 (N9823, N9785);
or OR3 (N9824, N9820, N4303, N3897);
xor XOR2 (N9825, N9817, N3009);
not NOT1 (N9826, N9811);
buf BUF1 (N9827, N9799);
not NOT1 (N9828, N9822);
nand NAND3 (N9829, N9828, N5967, N4398);
nand NAND2 (N9830, N9826, N3572);
xor XOR2 (N9831, N9824, N601);
buf BUF1 (N9832, N9830);
or OR4 (N9833, N9831, N696, N511, N8760);
not NOT1 (N9834, N9823);
nor NOR3 (N9835, N9819, N3218, N2629);
buf BUF1 (N9836, N9812);
nor NOR2 (N9837, N9833, N9475);
or OR3 (N9838, N9835, N5286, N173);
not NOT1 (N9839, N9832);
xor XOR2 (N9840, N9839, N1415);
xor XOR2 (N9841, N9837, N4921);
and AND3 (N9842, N9827, N1189, N6283);
nor NOR4 (N9843, N9841, N5566, N2441, N1485);
or OR4 (N9844, N9838, N603, N3280, N4189);
nor NOR2 (N9845, N9843, N3);
nand NAND4 (N9846, N9825, N624, N3251, N7755);
not NOT1 (N9847, N9845);
xor XOR2 (N9848, N9844, N45);
buf BUF1 (N9849, N9834);
nand NAND2 (N9850, N9849, N8851);
nor NOR2 (N9851, N9847, N3969);
buf BUF1 (N9852, N9840);
xor XOR2 (N9853, N9836, N609);
nor NOR2 (N9854, N9829, N6177);
nand NAND4 (N9855, N9813, N1419, N262, N6868);
buf BUF1 (N9856, N9855);
xor XOR2 (N9857, N9846, N1277);
buf BUF1 (N9858, N9848);
and AND4 (N9859, N9857, N9358, N3264, N2672);
xor XOR2 (N9860, N9859, N5726);
nor NOR2 (N9861, N9842, N7937);
nor NOR4 (N9862, N9851, N8944, N9595, N2101);
or OR3 (N9863, N9858, N2113, N3379);
not NOT1 (N9864, N9850);
nor NOR3 (N9865, N9860, N4173, N6649);
or OR4 (N9866, N9864, N7461, N5158, N8661);
not NOT1 (N9867, N9866);
nand NAND4 (N9868, N9867, N2838, N7841, N578);
nand NAND2 (N9869, N9853, N3649);
or OR4 (N9870, N9863, N4126, N255, N8731);
buf BUF1 (N9871, N9870);
not NOT1 (N9872, N9821);
or OR2 (N9873, N9872, N4600);
buf BUF1 (N9874, N9854);
nor NOR2 (N9875, N9873, N1050);
xor XOR2 (N9876, N9868, N4944);
buf BUF1 (N9877, N9869);
or OR2 (N9878, N9862, N1305);
xor XOR2 (N9879, N9877, N8297);
and AND3 (N9880, N9874, N3768, N2844);
nand NAND2 (N9881, N9878, N821);
nand NAND3 (N9882, N9852, N9328, N9097);
nand NAND3 (N9883, N9881, N4249, N2681);
and AND4 (N9884, N9861, N2510, N2584, N4304);
buf BUF1 (N9885, N9871);
nor NOR2 (N9886, N9884, N4751);
or OR2 (N9887, N9886, N6746);
xor XOR2 (N9888, N9887, N191);
not NOT1 (N9889, N9875);
not NOT1 (N9890, N9879);
not NOT1 (N9891, N9883);
xor XOR2 (N9892, N9890, N6812);
or OR2 (N9893, N9891, N4602);
buf BUF1 (N9894, N9893);
xor XOR2 (N9895, N9889, N3526);
or OR2 (N9896, N9865, N7626);
or OR2 (N9897, N9888, N6999);
buf BUF1 (N9898, N9882);
buf BUF1 (N9899, N9885);
and AND4 (N9900, N9899, N8345, N2840, N4899);
xor XOR2 (N9901, N9897, N5674);
buf BUF1 (N9902, N9895);
xor XOR2 (N9903, N9892, N5278);
xor XOR2 (N9904, N9898, N3976);
buf BUF1 (N9905, N9876);
nand NAND3 (N9906, N9900, N148, N5067);
or OR4 (N9907, N9906, N9716, N6231, N1374);
nand NAND3 (N9908, N9901, N1509, N1211);
nor NOR3 (N9909, N9905, N566, N1256);
buf BUF1 (N9910, N9909);
buf BUF1 (N9911, N9902);
xor XOR2 (N9912, N9903, N8462);
not NOT1 (N9913, N9904);
not NOT1 (N9914, N9908);
and AND3 (N9915, N9907, N3002, N9545);
and AND2 (N9916, N9856, N4384);
nand NAND4 (N9917, N9894, N7066, N9187, N7158);
nor NOR4 (N9918, N9915, N333, N9304, N5301);
xor XOR2 (N9919, N9918, N5827);
xor XOR2 (N9920, N9911, N782);
not NOT1 (N9921, N9896);
xor XOR2 (N9922, N9921, N4232);
and AND4 (N9923, N9917, N9042, N6551, N2845);
buf BUF1 (N9924, N9913);
buf BUF1 (N9925, N9910);
xor XOR2 (N9926, N9925, N3837);
xor XOR2 (N9927, N9920, N8759);
xor XOR2 (N9928, N9924, N702);
not NOT1 (N9929, N9927);
xor XOR2 (N9930, N9916, N4908);
nor NOR4 (N9931, N9922, N9821, N4493, N2311);
and AND3 (N9932, N9880, N2882, N5953);
xor XOR2 (N9933, N9919, N3348);
not NOT1 (N9934, N9912);
nand NAND2 (N9935, N9923, N8525);
nand NAND3 (N9936, N9928, N7942, N2485);
nor NOR2 (N9937, N9930, N6497);
xor XOR2 (N9938, N9931, N573);
and AND3 (N9939, N9935, N1882, N4013);
buf BUF1 (N9940, N9914);
nor NOR4 (N9941, N9934, N9567, N7592, N6310);
nor NOR4 (N9942, N9926, N8801, N4058, N6533);
buf BUF1 (N9943, N9941);
or OR3 (N9944, N9938, N6304, N1695);
nand NAND3 (N9945, N9936, N428, N4169);
nand NAND2 (N9946, N9933, N9460);
nand NAND4 (N9947, N9946, N2314, N7519, N6191);
or OR3 (N9948, N9945, N5814, N8225);
and AND3 (N9949, N9944, N3234, N5874);
nor NOR3 (N9950, N9947, N3423, N8150);
not NOT1 (N9951, N9942);
nor NOR3 (N9952, N9948, N6280, N9298);
xor XOR2 (N9953, N9952, N953);
not NOT1 (N9954, N9949);
buf BUF1 (N9955, N9954);
nand NAND4 (N9956, N9940, N3282, N9598, N6663);
nand NAND4 (N9957, N9953, N4040, N2225, N6701);
nand NAND4 (N9958, N9943, N1591, N8621, N7845);
buf BUF1 (N9959, N9956);
nand NAND3 (N9960, N9950, N6609, N1929);
and AND2 (N9961, N9932, N7062);
and AND3 (N9962, N9957, N2541, N7593);
nand NAND3 (N9963, N9958, N2149, N6632);
xor XOR2 (N9964, N9962, N9054);
and AND4 (N9965, N9939, N8159, N7053, N9074);
xor XOR2 (N9966, N9960, N8020);
or OR2 (N9967, N9966, N4106);
buf BUF1 (N9968, N9964);
buf BUF1 (N9969, N9965);
xor XOR2 (N9970, N9968, N413);
nor NOR2 (N9971, N9937, N649);
not NOT1 (N9972, N9961);
or OR3 (N9973, N9929, N576, N2392);
xor XOR2 (N9974, N9967, N6403);
nand NAND2 (N9975, N9969, N8925);
nor NOR3 (N9976, N9975, N3118, N5334);
not NOT1 (N9977, N9959);
nand NAND2 (N9978, N9972, N9663);
and AND2 (N9979, N9976, N1920);
buf BUF1 (N9980, N9971);
xor XOR2 (N9981, N9980, N3467);
not NOT1 (N9982, N9978);
xor XOR2 (N9983, N9955, N8281);
buf BUF1 (N9984, N9963);
nor NOR4 (N9985, N9970, N2647, N3070, N6915);
buf BUF1 (N9986, N9984);
not NOT1 (N9987, N9985);
nor NOR4 (N9988, N9977, N2453, N8938, N5434);
not NOT1 (N9989, N9986);
buf BUF1 (N9990, N9951);
nor NOR3 (N9991, N9982, N6056, N540);
xor XOR2 (N9992, N9990, N7371);
nor NOR3 (N9993, N9991, N7589, N605);
buf BUF1 (N9994, N9987);
not NOT1 (N9995, N9974);
and AND2 (N9996, N9983, N7944);
nand NAND2 (N9997, N9995, N953);
or OR3 (N9998, N9994, N240, N3723);
nand NAND4 (N9999, N9993, N4809, N79, N4625);
nor NOR2 (N10000, N9981, N8426);
buf BUF1 (N10001, N10000);
not NOT1 (N10002, N9989);
buf BUF1 (N10003, N9979);
xor XOR2 (N10004, N10002, N9576);
nor NOR2 (N10005, N9999, N3918);
buf BUF1 (N10006, N10001);
or OR4 (N10007, N9992, N4486, N7369, N6939);
or OR2 (N10008, N10007, N3619);
xor XOR2 (N10009, N9998, N1572);
xor XOR2 (N10010, N10008, N8817);
and AND4 (N10011, N10005, N4668, N1755, N6998);
xor XOR2 (N10012, N9988, N6458);
or OR2 (N10013, N10006, N1860);
and AND4 (N10014, N10012, N7976, N8545, N315);
or OR2 (N10015, N9973, N6574);
and AND2 (N10016, N9997, N3709);
and AND4 (N10017, N10016, N8795, N2683, N4989);
and AND4 (N10018, N10003, N7163, N728, N8019);
xor XOR2 (N10019, N10015, N6860);
and AND3 (N10020, N10018, N3277, N8355);
nor NOR4 (N10021, N10013, N4149, N6067, N9724);
nor NOR4 (N10022, N10017, N5875, N1519, N3593);
not NOT1 (N10023, N9996);
nor NOR4 (N10024, N10019, N3136, N1730, N8264);
not NOT1 (N10025, N10020);
or OR4 (N10026, N10025, N534, N4481, N7120);
and AND2 (N10027, N10004, N7017);
buf BUF1 (N10028, N10023);
and AND4 (N10029, N10009, N4462, N2921, N2048);
buf BUF1 (N10030, N10010);
xor XOR2 (N10031, N10024, N3427);
not NOT1 (N10032, N10021);
nor NOR2 (N10033, N10028, N6809);
or OR4 (N10034, N10027, N8821, N160, N1767);
nand NAND2 (N10035, N10031, N2436);
nor NOR3 (N10036, N10035, N7430, N9636);
buf BUF1 (N10037, N10029);
buf BUF1 (N10038, N10037);
nor NOR4 (N10039, N10011, N7530, N180, N5707);
nand NAND4 (N10040, N10014, N3096, N2932, N1929);
buf BUF1 (N10041, N10039);
and AND4 (N10042, N10038, N8491, N4955, N4960);
or OR3 (N10043, N10042, N8150, N262);
and AND2 (N10044, N10022, N7883);
nand NAND4 (N10045, N10036, N6450, N8167, N5048);
not NOT1 (N10046, N10044);
buf BUF1 (N10047, N10033);
and AND3 (N10048, N10046, N7796, N4181);
not NOT1 (N10049, N10032);
nor NOR4 (N10050, N10026, N8481, N4990, N6703);
or OR4 (N10051, N10048, N9891, N8142, N232);
or OR3 (N10052, N10040, N1771, N233);
buf BUF1 (N10053, N10041);
nand NAND4 (N10054, N10030, N3294, N242, N9941);
or OR2 (N10055, N10034, N479);
xor XOR2 (N10056, N10055, N1684);
buf BUF1 (N10057, N10054);
or OR3 (N10058, N10053, N5927, N5537);
and AND2 (N10059, N10045, N7178);
and AND3 (N10060, N10050, N2286, N10008);
or OR2 (N10061, N10057, N7148);
nand NAND3 (N10062, N10060, N9135, N7656);
not NOT1 (N10063, N10056);
or OR3 (N10064, N10058, N4305, N6217);
buf BUF1 (N10065, N10063);
or OR2 (N10066, N10059, N8999);
nand NAND3 (N10067, N10049, N902, N8177);
buf BUF1 (N10068, N10052);
or OR4 (N10069, N10051, N9187, N6549, N3742);
buf BUF1 (N10070, N10043);
or OR4 (N10071, N10061, N4912, N2382, N5019);
and AND2 (N10072, N10068, N3946);
or OR2 (N10073, N10071, N4019);
nand NAND3 (N10074, N10065, N1370, N7891);
not NOT1 (N10075, N10073);
nand NAND2 (N10076, N10062, N6805);
nand NAND4 (N10077, N10072, N6134, N2925, N6233);
xor XOR2 (N10078, N10074, N3280);
buf BUF1 (N10079, N10076);
nand NAND4 (N10080, N10069, N8193, N6086, N69);
nand NAND3 (N10081, N10080, N7246, N9910);
or OR3 (N10082, N10064, N2912, N2047);
nor NOR2 (N10083, N10082, N4124);
nor NOR3 (N10084, N10067, N1074, N2882);
buf BUF1 (N10085, N10047);
xor XOR2 (N10086, N10077, N7361);
and AND4 (N10087, N10085, N1656, N3149, N427);
xor XOR2 (N10088, N10081, N1523);
not NOT1 (N10089, N10078);
or OR2 (N10090, N10079, N1405);
nor NOR3 (N10091, N10088, N8734, N542);
not NOT1 (N10092, N10087);
nand NAND4 (N10093, N10092, N7662, N8403, N9774);
not NOT1 (N10094, N10086);
and AND4 (N10095, N10089, N6190, N871, N7603);
buf BUF1 (N10096, N10084);
nor NOR2 (N10097, N10083, N2309);
and AND2 (N10098, N10091, N4442);
buf BUF1 (N10099, N10098);
nor NOR2 (N10100, N10075, N5106);
buf BUF1 (N10101, N10093);
buf BUF1 (N10102, N10066);
and AND4 (N10103, N10096, N2125, N9358, N7650);
nor NOR3 (N10104, N10103, N8518, N931);
and AND2 (N10105, N10099, N4458);
not NOT1 (N10106, N10104);
not NOT1 (N10107, N10101);
or OR2 (N10108, N10107, N5391);
buf BUF1 (N10109, N10095);
nand NAND3 (N10110, N10100, N6698, N6215);
nand NAND4 (N10111, N10109, N8309, N535, N5478);
nor NOR4 (N10112, N10105, N6754, N4697, N5531);
not NOT1 (N10113, N10094);
not NOT1 (N10114, N10090);
xor XOR2 (N10115, N10113, N3083);
or OR4 (N10116, N10070, N2851, N806, N10015);
nand NAND4 (N10117, N10108, N3655, N2314, N8143);
nor NOR2 (N10118, N10106, N5106);
nand NAND2 (N10119, N10111, N4621);
xor XOR2 (N10120, N10116, N6842);
and AND2 (N10121, N10119, N8683);
or OR2 (N10122, N10115, N7722);
or OR3 (N10123, N10097, N2431, N4007);
and AND2 (N10124, N10122, N3844);
nand NAND2 (N10125, N10118, N9535);
xor XOR2 (N10126, N10102, N229);
or OR4 (N10127, N10114, N10117, N4761, N8793);
nor NOR2 (N10128, N6998, N7200);
xor XOR2 (N10129, N10124, N9955);
not NOT1 (N10130, N10120);
not NOT1 (N10131, N10130);
not NOT1 (N10132, N10123);
nand NAND2 (N10133, N10126, N1861);
nand NAND4 (N10134, N10132, N218, N1665, N5849);
not NOT1 (N10135, N10129);
and AND2 (N10136, N10134, N7593);
buf BUF1 (N10137, N10112);
and AND4 (N10138, N10136, N7182, N6922, N2295);
nand NAND2 (N10139, N10131, N7767);
or OR2 (N10140, N10128, N3064);
nor NOR4 (N10141, N10137, N4642, N6313, N6226);
buf BUF1 (N10142, N10139);
xor XOR2 (N10143, N10135, N1776);
nor NOR4 (N10144, N10141, N8511, N7370, N9604);
or OR2 (N10145, N10125, N7602);
nor NOR4 (N10146, N10121, N10016, N3682, N421);
xor XOR2 (N10147, N10140, N9151);
nor NOR3 (N10148, N10146, N5754, N5075);
nand NAND3 (N10149, N10110, N1184, N2730);
nor NOR2 (N10150, N10127, N2361);
nand NAND3 (N10151, N10142, N4083, N4786);
and AND2 (N10152, N10133, N250);
and AND4 (N10153, N10152, N134, N6893, N1825);
nor NOR3 (N10154, N10151, N1144, N735);
nand NAND4 (N10155, N10145, N3931, N1671, N6197);
not NOT1 (N10156, N10148);
buf BUF1 (N10157, N10138);
or OR4 (N10158, N10155, N9126, N9028, N5100);
buf BUF1 (N10159, N10156);
xor XOR2 (N10160, N10144, N1089);
nor NOR3 (N10161, N10153, N6230, N9019);
not NOT1 (N10162, N10159);
and AND3 (N10163, N10160, N5267, N5968);
and AND4 (N10164, N10163, N7043, N202, N203);
nand NAND4 (N10165, N10164, N9963, N7879, N6163);
nor NOR4 (N10166, N10154, N5418, N3848, N5538);
or OR2 (N10167, N10150, N6155);
xor XOR2 (N10168, N10167, N1340);
xor XOR2 (N10169, N10158, N5391);
or OR2 (N10170, N10165, N4584);
buf BUF1 (N10171, N10162);
nand NAND3 (N10172, N10171, N3605, N521);
nor NOR3 (N10173, N10149, N3835, N7042);
nor NOR4 (N10174, N10166, N5794, N8422, N61);
or OR4 (N10175, N10173, N4184, N7201, N7237);
nor NOR4 (N10176, N10157, N2055, N857, N479);
xor XOR2 (N10177, N10161, N9727);
and AND2 (N10178, N10168, N855);
xor XOR2 (N10179, N10174, N4518);
nor NOR2 (N10180, N10172, N9160);
and AND3 (N10181, N10177, N2267, N457);
nand NAND2 (N10182, N10175, N5017);
nor NOR3 (N10183, N10178, N6952, N1523);
not NOT1 (N10184, N10180);
nand NAND3 (N10185, N10176, N6300, N4926);
not NOT1 (N10186, N10170);
not NOT1 (N10187, N10143);
or OR4 (N10188, N10187, N3078, N692, N7483);
nor NOR3 (N10189, N10186, N470, N646);
not NOT1 (N10190, N10185);
not NOT1 (N10191, N10190);
or OR4 (N10192, N10184, N4413, N9239, N5200);
and AND4 (N10193, N10147, N2143, N4200, N6372);
xor XOR2 (N10194, N10191, N4709);
and AND4 (N10195, N10193, N1623, N2277, N3518);
not NOT1 (N10196, N10179);
xor XOR2 (N10197, N10181, N8656);
and AND3 (N10198, N10196, N2466, N4943);
not NOT1 (N10199, N10192);
xor XOR2 (N10200, N10169, N3963);
and AND2 (N10201, N10194, N418);
nand NAND3 (N10202, N10182, N4840, N4376);
xor XOR2 (N10203, N10197, N9465);
or OR2 (N10204, N10183, N6363);
nor NOR2 (N10205, N10202, N83);
and AND3 (N10206, N10203, N4941, N8254);
not NOT1 (N10207, N10198);
nor NOR4 (N10208, N10204, N4787, N8427, N5203);
not NOT1 (N10209, N10195);
nand NAND3 (N10210, N10199, N343, N2586);
and AND4 (N10211, N10210, N10153, N4377, N6887);
xor XOR2 (N10212, N10188, N6085);
and AND4 (N10213, N10201, N4339, N3628, N9962);
nand NAND3 (N10214, N10211, N9271, N281);
nand NAND4 (N10215, N10212, N2026, N8324, N6269);
not NOT1 (N10216, N10200);
xor XOR2 (N10217, N10213, N1018);
and AND2 (N10218, N10205, N2982);
and AND3 (N10219, N10206, N9473, N3715);
not NOT1 (N10220, N10189);
buf BUF1 (N10221, N10209);
buf BUF1 (N10222, N10218);
nor NOR4 (N10223, N10214, N7398, N4629, N1626);
not NOT1 (N10224, N10208);
not NOT1 (N10225, N10222);
or OR4 (N10226, N10215, N3681, N436, N2035);
xor XOR2 (N10227, N10223, N9418);
nand NAND3 (N10228, N10225, N8835, N1152);
nand NAND2 (N10229, N10220, N8736);
or OR3 (N10230, N10229, N6487, N3987);
not NOT1 (N10231, N10227);
buf BUF1 (N10232, N10207);
and AND2 (N10233, N10221, N9285);
nand NAND2 (N10234, N10226, N362);
buf BUF1 (N10235, N10233);
buf BUF1 (N10236, N10234);
xor XOR2 (N10237, N10230, N5298);
and AND3 (N10238, N10236, N10045, N8976);
not NOT1 (N10239, N10232);
and AND4 (N10240, N10239, N1278, N3354, N5176);
nor NOR4 (N10241, N10216, N2269, N7157, N3555);
buf BUF1 (N10242, N10231);
or OR4 (N10243, N10228, N6321, N5241, N447);
or OR2 (N10244, N10217, N9148);
nand NAND4 (N10245, N10235, N1880, N7588, N7397);
buf BUF1 (N10246, N10241);
or OR2 (N10247, N10219, N1653);
or OR2 (N10248, N10245, N9271);
or OR3 (N10249, N10237, N2069, N7519);
buf BUF1 (N10250, N10246);
not NOT1 (N10251, N10242);
and AND3 (N10252, N10238, N5993, N5752);
buf BUF1 (N10253, N10251);
nor NOR3 (N10254, N10248, N798, N1573);
nor NOR4 (N10255, N10252, N127, N8354, N4578);
or OR4 (N10256, N10254, N914, N2527, N1917);
not NOT1 (N10257, N10255);
nor NOR3 (N10258, N10244, N4469, N8738);
xor XOR2 (N10259, N10224, N8314);
nand NAND4 (N10260, N10259, N1777, N4090, N2702);
nand NAND2 (N10261, N10250, N10095);
not NOT1 (N10262, N10249);
and AND3 (N10263, N10253, N5902, N7353);
nand NAND4 (N10264, N10261, N7450, N2553, N6511);
nor NOR2 (N10265, N10256, N4260);
and AND3 (N10266, N10258, N7312, N9150);
nor NOR2 (N10267, N10264, N3157);
nand NAND3 (N10268, N10266, N7812, N7375);
buf BUF1 (N10269, N10243);
nor NOR2 (N10270, N10269, N7606);
xor XOR2 (N10271, N10268, N2177);
not NOT1 (N10272, N10240);
xor XOR2 (N10273, N10267, N2072);
nand NAND4 (N10274, N10272, N9072, N7386, N1081);
buf BUF1 (N10275, N10271);
nand NAND3 (N10276, N10257, N4335, N2890);
xor XOR2 (N10277, N10270, N8627);
and AND3 (N10278, N10262, N7906, N1666);
or OR2 (N10279, N10247, N3961);
or OR2 (N10280, N10278, N9254);
xor XOR2 (N10281, N10276, N7719);
nand NAND4 (N10282, N10265, N4328, N6423, N4134);
not NOT1 (N10283, N10260);
and AND3 (N10284, N10280, N2626, N5308);
xor XOR2 (N10285, N10281, N1154);
buf BUF1 (N10286, N10263);
buf BUF1 (N10287, N10274);
or OR4 (N10288, N10283, N7878, N4889, N1724);
not NOT1 (N10289, N10288);
and AND2 (N10290, N10287, N842);
nand NAND3 (N10291, N10289, N1569, N3062);
not NOT1 (N10292, N10275);
not NOT1 (N10293, N10286);
or OR4 (N10294, N10290, N7867, N279, N532);
xor XOR2 (N10295, N10291, N4667);
buf BUF1 (N10296, N10277);
not NOT1 (N10297, N10293);
buf BUF1 (N10298, N10282);
and AND3 (N10299, N10295, N2514, N4221);
or OR4 (N10300, N10284, N1151, N3628, N4952);
and AND2 (N10301, N10279, N4398);
nor NOR3 (N10302, N10297, N2060, N3379);
nand NAND4 (N10303, N10301, N3515, N8876, N997);
nor NOR4 (N10304, N10298, N738, N256, N3759);
and AND4 (N10305, N10299, N4730, N4575, N7470);
nand NAND2 (N10306, N10296, N1816);
nand NAND3 (N10307, N10305, N2624, N7332);
and AND3 (N10308, N10302, N7878, N9587);
xor XOR2 (N10309, N10294, N3484);
or OR3 (N10310, N10304, N828, N8262);
nand NAND2 (N10311, N10292, N1791);
nor NOR3 (N10312, N10307, N4302, N9258);
buf BUF1 (N10313, N10309);
and AND2 (N10314, N10300, N3317);
buf BUF1 (N10315, N10311);
xor XOR2 (N10316, N10310, N9475);
xor XOR2 (N10317, N10315, N3853);
nor NOR2 (N10318, N10312, N8868);
nor NOR4 (N10319, N10306, N2206, N5973, N9816);
buf BUF1 (N10320, N10316);
xor XOR2 (N10321, N10317, N2206);
nand NAND2 (N10322, N10313, N4167);
and AND2 (N10323, N10308, N7258);
nor NOR3 (N10324, N10318, N7190, N9781);
nand NAND3 (N10325, N10323, N4794, N4517);
nor NOR2 (N10326, N10321, N6782);
not NOT1 (N10327, N10325);
nor NOR2 (N10328, N10326, N397);
nor NOR4 (N10329, N10314, N6314, N3982, N3204);
and AND4 (N10330, N10328, N6523, N3242, N9982);
xor XOR2 (N10331, N10327, N6545);
nor NOR4 (N10332, N10273, N4293, N5125, N6943);
and AND2 (N10333, N10319, N8161);
not NOT1 (N10334, N10330);
xor XOR2 (N10335, N10333, N620);
nand NAND4 (N10336, N10335, N1609, N7609, N10038);
nor NOR4 (N10337, N10336, N4011, N5107, N6377);
nand NAND3 (N10338, N10285, N871, N2327);
xor XOR2 (N10339, N10331, N1278);
and AND4 (N10340, N10329, N1123, N8288, N4847);
or OR4 (N10341, N10340, N2320, N5472, N5978);
nand NAND3 (N10342, N10341, N8455, N3792);
and AND2 (N10343, N10320, N7098);
nand NAND4 (N10344, N10332, N5856, N3570, N5551);
not NOT1 (N10345, N10324);
nand NAND3 (N10346, N10344, N4118, N1362);
buf BUF1 (N10347, N10342);
xor XOR2 (N10348, N10334, N1549);
or OR2 (N10349, N10338, N2009);
or OR3 (N10350, N10348, N7803, N2769);
nand NAND2 (N10351, N10343, N6368);
xor XOR2 (N10352, N10350, N4003);
and AND2 (N10353, N10347, N856);
buf BUF1 (N10354, N10337);
buf BUF1 (N10355, N10354);
not NOT1 (N10356, N10351);
nand NAND4 (N10357, N10339, N2664, N7887, N1201);
buf BUF1 (N10358, N10346);
or OR2 (N10359, N10303, N3506);
and AND4 (N10360, N10357, N645, N6084, N8269);
or OR4 (N10361, N10345, N3187, N9511, N2636);
or OR4 (N10362, N10353, N8117, N880, N1926);
nor NOR4 (N10363, N10349, N1039, N1524, N277);
nor NOR4 (N10364, N10360, N2875, N6768, N4869);
nor NOR2 (N10365, N10322, N8864);
or OR4 (N10366, N10364, N4735, N7175, N8888);
nand NAND3 (N10367, N10366, N506, N8082);
nor NOR3 (N10368, N10352, N632, N10119);
not NOT1 (N10369, N10365);
nor NOR4 (N10370, N10358, N8411, N3178, N4015);
xor XOR2 (N10371, N10359, N4089);
or OR3 (N10372, N10369, N4371, N10220);
buf BUF1 (N10373, N10363);
nand NAND3 (N10374, N10356, N6000, N4334);
nand NAND2 (N10375, N10374, N8316);
or OR3 (N10376, N10362, N8704, N4588);
nand NAND4 (N10377, N10361, N8058, N2772, N7121);
nand NAND3 (N10378, N10375, N360, N7129);
or OR4 (N10379, N10373, N7750, N1199, N8596);
nand NAND4 (N10380, N10372, N6406, N8393, N5735);
and AND4 (N10381, N10355, N7548, N2370, N3624);
buf BUF1 (N10382, N10379);
xor XOR2 (N10383, N10382, N3290);
or OR3 (N10384, N10367, N8283, N1345);
nor NOR4 (N10385, N10377, N5423, N7347, N9925);
nand NAND4 (N10386, N10370, N198, N91, N9018);
nand NAND2 (N10387, N10371, N8247);
not NOT1 (N10388, N10381);
and AND4 (N10389, N10387, N1287, N836, N7666);
and AND2 (N10390, N10378, N4916);
not NOT1 (N10391, N10380);
or OR3 (N10392, N10391, N5136, N881);
not NOT1 (N10393, N10389);
buf BUF1 (N10394, N10384);
buf BUF1 (N10395, N10388);
and AND2 (N10396, N10368, N409);
not NOT1 (N10397, N10396);
nand NAND3 (N10398, N10383, N10397, N1264);
buf BUF1 (N10399, N7148);
xor XOR2 (N10400, N10385, N9868);
nor NOR4 (N10401, N10393, N7792, N6898, N3344);
or OR4 (N10402, N10394, N7283, N4132, N1623);
nor NOR4 (N10403, N10392, N9104, N9450, N3247);
not NOT1 (N10404, N10386);
nand NAND2 (N10405, N10403, N5971);
buf BUF1 (N10406, N10395);
xor XOR2 (N10407, N10398, N5739);
and AND4 (N10408, N10404, N10043, N5340, N7451);
nand NAND4 (N10409, N10408, N7438, N5106, N8103);
nor NOR2 (N10410, N10409, N2193);
nor NOR3 (N10411, N10376, N2667, N3799);
or OR2 (N10412, N10402, N4883);
not NOT1 (N10413, N10410);
not NOT1 (N10414, N10406);
nor NOR4 (N10415, N10399, N3307, N2293, N7236);
xor XOR2 (N10416, N10390, N2616);
buf BUF1 (N10417, N10415);
not NOT1 (N10418, N10412);
nor NOR4 (N10419, N10414, N10299, N5085, N8080);
xor XOR2 (N10420, N10418, N5686);
not NOT1 (N10421, N10420);
and AND2 (N10422, N10407, N2059);
not NOT1 (N10423, N10413);
nand NAND2 (N10424, N10401, N5217);
and AND2 (N10425, N10417, N5160);
and AND2 (N10426, N10423, N2305);
or OR4 (N10427, N10424, N2957, N7083, N806);
buf BUF1 (N10428, N10422);
not NOT1 (N10429, N10425);
nor NOR2 (N10430, N10428, N3857);
nand NAND4 (N10431, N10427, N8544, N5255, N7549);
buf BUF1 (N10432, N10430);
and AND4 (N10433, N10432, N7577, N2394, N1182);
and AND3 (N10434, N10426, N7020, N2206);
xor XOR2 (N10435, N10411, N2803);
buf BUF1 (N10436, N10400);
nor NOR2 (N10437, N10435, N8791);
or OR4 (N10438, N10405, N8006, N1251, N760);
buf BUF1 (N10439, N10437);
xor XOR2 (N10440, N10416, N246);
not NOT1 (N10441, N10429);
or OR4 (N10442, N10419, N9933, N10241, N8169);
buf BUF1 (N10443, N10442);
nand NAND2 (N10444, N10434, N10172);
nor NOR2 (N10445, N10439, N4021);
not NOT1 (N10446, N10440);
buf BUF1 (N10447, N10443);
and AND3 (N10448, N10438, N5660, N7728);
nand NAND3 (N10449, N10431, N22, N6922);
and AND2 (N10450, N10446, N2754);
or OR3 (N10451, N10433, N7095, N1954);
xor XOR2 (N10452, N10441, N10315);
xor XOR2 (N10453, N10451, N6915);
xor XOR2 (N10454, N10452, N2969);
or OR3 (N10455, N10447, N9859, N4289);
buf BUF1 (N10456, N10448);
or OR4 (N10457, N10445, N10184, N9327, N2667);
nor NOR2 (N10458, N10457, N1683);
nor NOR3 (N10459, N10421, N8369, N2468);
and AND2 (N10460, N10436, N7153);
nor NOR2 (N10461, N10458, N3189);
nand NAND3 (N10462, N10459, N10157, N9928);
nand NAND4 (N10463, N10449, N2381, N2223, N9770);
xor XOR2 (N10464, N10463, N995);
and AND3 (N10465, N10455, N8569, N9336);
not NOT1 (N10466, N10444);
and AND4 (N10467, N10466, N467, N6191, N5847);
xor XOR2 (N10468, N10453, N2936);
xor XOR2 (N10469, N10454, N5752);
xor XOR2 (N10470, N10461, N7521);
nor NOR3 (N10471, N10470, N577, N8806);
xor XOR2 (N10472, N10468, N4034);
xor XOR2 (N10473, N10469, N6549);
nor NOR2 (N10474, N10450, N7119);
xor XOR2 (N10475, N10467, N4483);
buf BUF1 (N10476, N10465);
nor NOR3 (N10477, N10460, N5744, N675);
not NOT1 (N10478, N10462);
xor XOR2 (N10479, N10464, N3217);
nand NAND3 (N10480, N10473, N7559, N5514);
or OR2 (N10481, N10474, N6084);
and AND4 (N10482, N10471, N8896, N9893, N900);
nor NOR2 (N10483, N10472, N1201);
not NOT1 (N10484, N10456);
or OR4 (N10485, N10482, N3217, N1850, N5949);
xor XOR2 (N10486, N10475, N4415);
nand NAND2 (N10487, N10485, N2732);
and AND4 (N10488, N10480, N2763, N2612, N661);
nand NAND3 (N10489, N10478, N7217, N4917);
or OR4 (N10490, N10479, N9564, N281, N721);
nand NAND3 (N10491, N10487, N1174, N7195);
buf BUF1 (N10492, N10484);
and AND2 (N10493, N10483, N4929);
nor NOR2 (N10494, N10481, N3355);
not NOT1 (N10495, N10476);
not NOT1 (N10496, N10491);
or OR4 (N10497, N10493, N7890, N8860, N5554);
or OR2 (N10498, N10486, N4576);
and AND2 (N10499, N10494, N8065);
xor XOR2 (N10500, N10498, N270);
and AND2 (N10501, N10489, N2300);
buf BUF1 (N10502, N10501);
not NOT1 (N10503, N10495);
and AND4 (N10504, N10499, N647, N6683, N1978);
xor XOR2 (N10505, N10497, N8693);
and AND3 (N10506, N10503, N2175, N7395);
or OR3 (N10507, N10496, N3989, N7846);
nor NOR2 (N10508, N10502, N10175);
xor XOR2 (N10509, N10506, N3328);
or OR4 (N10510, N10509, N6419, N8278, N9263);
buf BUF1 (N10511, N10505);
buf BUF1 (N10512, N10511);
not NOT1 (N10513, N10492);
or OR4 (N10514, N10477, N5251, N6160, N6258);
or OR4 (N10515, N10500, N8009, N7613, N2160);
not NOT1 (N10516, N10514);
nand NAND2 (N10517, N10516, N583);
nor NOR2 (N10518, N10510, N3276);
buf BUF1 (N10519, N10507);
or OR3 (N10520, N10488, N10232, N6114);
and AND4 (N10521, N10517, N3065, N8196, N5549);
buf BUF1 (N10522, N10518);
buf BUF1 (N10523, N10512);
or OR4 (N10524, N10504, N9705, N4660, N5223);
or OR4 (N10525, N10523, N6969, N5416, N4140);
and AND2 (N10526, N10524, N7846);
not NOT1 (N10527, N10513);
buf BUF1 (N10528, N10522);
not NOT1 (N10529, N10527);
not NOT1 (N10530, N10515);
xor XOR2 (N10531, N10525, N5626);
and AND2 (N10532, N10528, N4005);
nand NAND2 (N10533, N10520, N2076);
buf BUF1 (N10534, N10508);
nand NAND2 (N10535, N10532, N6289);
nand NAND4 (N10536, N10521, N5141, N8251, N9121);
not NOT1 (N10537, N10490);
not NOT1 (N10538, N10535);
nand NAND4 (N10539, N10529, N8573, N681, N7641);
and AND3 (N10540, N10530, N9475, N4012);
or OR3 (N10541, N10540, N3831, N10426);
not NOT1 (N10542, N10519);
nand NAND4 (N10543, N10534, N9077, N6778, N747);
nand NAND2 (N10544, N10543, N8459);
and AND4 (N10545, N10541, N9467, N9862, N4141);
nand NAND3 (N10546, N10537, N9452, N8748);
xor XOR2 (N10547, N10545, N4385);
and AND4 (N10548, N10542, N9456, N1653, N5924);
nand NAND3 (N10549, N10544, N5172, N6614);
not NOT1 (N10550, N10533);
buf BUF1 (N10551, N10538);
and AND3 (N10552, N10546, N6181, N10255);
nand NAND3 (N10553, N10531, N185, N8426);
xor XOR2 (N10554, N10547, N3077);
not NOT1 (N10555, N10526);
buf BUF1 (N10556, N10549);
buf BUF1 (N10557, N10551);
xor XOR2 (N10558, N10556, N8369);
or OR4 (N10559, N10548, N1207, N2167, N1794);
or OR2 (N10560, N10539, N2923);
xor XOR2 (N10561, N10557, N6216);
or OR3 (N10562, N10561, N5545, N6132);
nor NOR4 (N10563, N10554, N579, N6840, N10351);
and AND2 (N10564, N10558, N3340);
buf BUF1 (N10565, N10560);
nand NAND2 (N10566, N10562, N7528);
buf BUF1 (N10567, N10559);
nand NAND2 (N10568, N10563, N5697);
xor XOR2 (N10569, N10566, N6252);
and AND2 (N10570, N10569, N6112);
not NOT1 (N10571, N10568);
nor NOR3 (N10572, N10564, N3967, N9311);
nand NAND2 (N10573, N10570, N8230);
or OR3 (N10574, N10552, N1329, N3420);
buf BUF1 (N10575, N10571);
not NOT1 (N10576, N10575);
and AND2 (N10577, N10555, N2423);
xor XOR2 (N10578, N10576, N3830);
or OR2 (N10579, N10574, N2487);
nor NOR4 (N10580, N10550, N8232, N7611, N7246);
not NOT1 (N10581, N10553);
not NOT1 (N10582, N10565);
xor XOR2 (N10583, N10577, N3135);
buf BUF1 (N10584, N10536);
nor NOR4 (N10585, N10579, N3061, N10045, N5804);
xor XOR2 (N10586, N10580, N9329);
not NOT1 (N10587, N10585);
xor XOR2 (N10588, N10578, N10530);
not NOT1 (N10589, N10587);
and AND4 (N10590, N10589, N1254, N5159, N175);
xor XOR2 (N10591, N10582, N9991);
not NOT1 (N10592, N10590);
not NOT1 (N10593, N10573);
and AND4 (N10594, N10584, N8883, N9045, N5618);
xor XOR2 (N10595, N10591, N4992);
nor NOR2 (N10596, N10567, N5934);
buf BUF1 (N10597, N10596);
nand NAND2 (N10598, N10588, N1021);
and AND2 (N10599, N10583, N10517);
nor NOR2 (N10600, N10593, N663);
buf BUF1 (N10601, N10572);
or OR3 (N10602, N10581, N8051, N7683);
and AND3 (N10603, N10601, N2668, N555);
not NOT1 (N10604, N10599);
or OR4 (N10605, N10602, N6678, N9541, N4596);
buf BUF1 (N10606, N10592);
nor NOR2 (N10607, N10598, N5856);
nor NOR3 (N10608, N10597, N5909, N6390);
not NOT1 (N10609, N10600);
not NOT1 (N10610, N10595);
and AND4 (N10611, N10608, N921, N7921, N1037);
nand NAND2 (N10612, N10611, N5506);
or OR4 (N10613, N10609, N1370, N6322, N6581);
nand NAND3 (N10614, N10610, N1429, N1361);
not NOT1 (N10615, N10612);
not NOT1 (N10616, N10614);
nand NAND4 (N10617, N10607, N6234, N4529, N3104);
nand NAND2 (N10618, N10604, N3241);
or OR3 (N10619, N10618, N5505, N2370);
and AND4 (N10620, N10594, N8754, N8786, N6396);
xor XOR2 (N10621, N10603, N8166);
or OR3 (N10622, N10613, N713, N9401);
buf BUF1 (N10623, N10620);
nor NOR2 (N10624, N10586, N3630);
or OR4 (N10625, N10619, N5199, N4110, N2802);
nor NOR4 (N10626, N10605, N1787, N7700, N1123);
or OR2 (N10627, N10623, N7985);
nand NAND3 (N10628, N10624, N5931, N9103);
or OR3 (N10629, N10606, N2460, N6597);
not NOT1 (N10630, N10625);
nor NOR3 (N10631, N10617, N7663, N8515);
and AND4 (N10632, N10616, N10359, N6337, N2793);
buf BUF1 (N10633, N10631);
nor NOR2 (N10634, N10632, N10016);
nand NAND3 (N10635, N10615, N1239, N2297);
or OR4 (N10636, N10627, N3253, N6380, N1194);
nor NOR2 (N10637, N10629, N1088);
nor NOR3 (N10638, N10628, N8630, N1376);
xor XOR2 (N10639, N10636, N9847);
or OR3 (N10640, N10637, N175, N1410);
not NOT1 (N10641, N10635);
xor XOR2 (N10642, N10639, N10521);
and AND2 (N10643, N10638, N1309);
or OR2 (N10644, N10641, N2260);
nand NAND2 (N10645, N10644, N3400);
and AND4 (N10646, N10622, N10339, N2159, N9191);
not NOT1 (N10647, N10626);
or OR4 (N10648, N10621, N3232, N3426, N2115);
nand NAND3 (N10649, N10630, N2141, N9279);
not NOT1 (N10650, N10647);
nor NOR4 (N10651, N10650, N1726, N9269, N3141);
nor NOR4 (N10652, N10643, N5412, N5834, N2398);
not NOT1 (N10653, N10645);
and AND2 (N10654, N10640, N8797);
nor NOR2 (N10655, N10654, N7972);
nand NAND3 (N10656, N10648, N8267, N6948);
nand NAND3 (N10657, N10634, N4684, N419);
buf BUF1 (N10658, N10646);
and AND4 (N10659, N10633, N8075, N4020, N6842);
nor NOR3 (N10660, N10657, N8365, N573);
or OR4 (N10661, N10649, N3327, N7428, N9465);
xor XOR2 (N10662, N10661, N6570);
buf BUF1 (N10663, N10659);
not NOT1 (N10664, N10656);
and AND2 (N10665, N10652, N8611);
nor NOR2 (N10666, N10664, N10337);
buf BUF1 (N10667, N10658);
and AND4 (N10668, N10665, N8551, N9096, N7000);
and AND3 (N10669, N10666, N8686, N3648);
nand NAND3 (N10670, N10660, N2152, N6360);
not NOT1 (N10671, N10651);
buf BUF1 (N10672, N10670);
nor NOR2 (N10673, N10671, N6619);
xor XOR2 (N10674, N10669, N7374);
xor XOR2 (N10675, N10663, N5432);
and AND3 (N10676, N10662, N3011, N4154);
nand NAND2 (N10677, N10668, N6607);
not NOT1 (N10678, N10676);
not NOT1 (N10679, N10655);
and AND2 (N10680, N10653, N1900);
buf BUF1 (N10681, N10678);
nand NAND3 (N10682, N10672, N3221, N7428);
xor XOR2 (N10683, N10667, N9034);
xor XOR2 (N10684, N10673, N4914);
xor XOR2 (N10685, N10677, N5876);
xor XOR2 (N10686, N10675, N10241);
xor XOR2 (N10687, N10679, N314);
nand NAND3 (N10688, N10686, N5960, N4029);
or OR4 (N10689, N10684, N5675, N9549, N7563);
or OR4 (N10690, N10687, N1983, N6461, N3950);
nand NAND4 (N10691, N10680, N7521, N3182, N4891);
or OR3 (N10692, N10689, N3921, N10619);
and AND3 (N10693, N10681, N3786, N2004);
xor XOR2 (N10694, N10682, N2822);
xor XOR2 (N10695, N10691, N1544);
nor NOR4 (N10696, N10693, N2778, N5659, N4222);
nor NOR2 (N10697, N10690, N1069);
nor NOR2 (N10698, N10697, N5948);
buf BUF1 (N10699, N10694);
nor NOR3 (N10700, N10699, N5821, N2809);
and AND4 (N10701, N10642, N10691, N825, N8846);
nand NAND3 (N10702, N10701, N3942, N6615);
xor XOR2 (N10703, N10696, N1929);
nand NAND3 (N10704, N10695, N7825, N9540);
and AND3 (N10705, N10692, N5986, N7679);
not NOT1 (N10706, N10705);
not NOT1 (N10707, N10706);
not NOT1 (N10708, N10674);
xor XOR2 (N10709, N10683, N1083);
not NOT1 (N10710, N10703);
nand NAND4 (N10711, N10707, N484, N10483, N655);
or OR4 (N10712, N10709, N18, N5134, N10310);
and AND4 (N10713, N10700, N256, N8562, N1021);
xor XOR2 (N10714, N10713, N883);
xor XOR2 (N10715, N10710, N219);
nand NAND2 (N10716, N10685, N9772);
not NOT1 (N10717, N10714);
not NOT1 (N10718, N10704);
nand NAND4 (N10719, N10711, N3449, N6235, N3934);
nor NOR2 (N10720, N10698, N2838);
and AND4 (N10721, N10708, N10283, N9335, N5408);
or OR4 (N10722, N10720, N3391, N3041, N2173);
nor NOR2 (N10723, N10688, N816);
nand NAND3 (N10724, N10716, N7247, N2097);
xor XOR2 (N10725, N10724, N6849);
or OR4 (N10726, N10718, N2305, N6451, N7039);
nor NOR3 (N10727, N10715, N2571, N10709);
buf BUF1 (N10728, N10722);
xor XOR2 (N10729, N10725, N3274);
nand NAND2 (N10730, N10726, N6822);
nand NAND3 (N10731, N10719, N5296, N1824);
nor NOR2 (N10732, N10712, N186);
or OR4 (N10733, N10721, N1950, N2773, N4438);
or OR4 (N10734, N10728, N8999, N4267, N3768);
buf BUF1 (N10735, N10727);
nand NAND2 (N10736, N10735, N10537);
nand NAND3 (N10737, N10731, N6863, N4244);
and AND3 (N10738, N10717, N5216, N10078);
xor XOR2 (N10739, N10738, N10245);
xor XOR2 (N10740, N10736, N3366);
and AND4 (N10741, N10740, N4951, N2290, N5849);
buf BUF1 (N10742, N10737);
and AND4 (N10743, N10732, N7883, N9792, N428);
nand NAND4 (N10744, N10723, N615, N5890, N6420);
buf BUF1 (N10745, N10742);
or OR4 (N10746, N10730, N10405, N4316, N7828);
nor NOR3 (N10747, N10729, N4538, N7860);
nor NOR2 (N10748, N10744, N9678);
buf BUF1 (N10749, N10734);
nand NAND3 (N10750, N10702, N10681, N9561);
buf BUF1 (N10751, N10749);
nor NOR2 (N10752, N10750, N10087);
buf BUF1 (N10753, N10748);
buf BUF1 (N10754, N10743);
nand NAND2 (N10755, N10753, N6152);
and AND3 (N10756, N10739, N3623, N7027);
not NOT1 (N10757, N10751);
nor NOR2 (N10758, N10741, N10651);
and AND2 (N10759, N10757, N2796);
nand NAND4 (N10760, N10733, N6121, N4857, N6370);
nor NOR4 (N10761, N10746, N9274, N8344, N5750);
or OR3 (N10762, N10756, N3601, N3274);
xor XOR2 (N10763, N10754, N1054);
or OR4 (N10764, N10747, N7983, N5858, N1585);
buf BUF1 (N10765, N10758);
and AND4 (N10766, N10764, N8261, N4022, N3325);
or OR4 (N10767, N10760, N10505, N5403, N9802);
and AND4 (N10768, N10752, N2308, N647, N5359);
and AND4 (N10769, N10765, N6693, N2780, N6053);
nand NAND4 (N10770, N10766, N9674, N882, N6924);
or OR3 (N10771, N10755, N2180, N5167);
or OR3 (N10772, N10759, N667, N5084);
nand NAND4 (N10773, N10763, N6689, N9651, N6424);
and AND4 (N10774, N10767, N9107, N1635, N8037);
nor NOR2 (N10775, N10769, N3629);
and AND3 (N10776, N10762, N9394, N7885);
not NOT1 (N10777, N10768);
and AND3 (N10778, N10771, N2840, N4931);
nand NAND4 (N10779, N10745, N10150, N2643, N4779);
not NOT1 (N10780, N10779);
xor XOR2 (N10781, N10775, N7857);
not NOT1 (N10782, N10781);
buf BUF1 (N10783, N10782);
or OR3 (N10784, N10777, N1334, N8624);
nand NAND2 (N10785, N10783, N5961);
or OR4 (N10786, N10780, N3945, N3465, N2091);
xor XOR2 (N10787, N10778, N9461);
and AND2 (N10788, N10784, N6246);
and AND2 (N10789, N10770, N7495);
buf BUF1 (N10790, N10785);
xor XOR2 (N10791, N10774, N9413);
and AND4 (N10792, N10786, N10123, N1027, N6867);
xor XOR2 (N10793, N10790, N4391);
nor NOR3 (N10794, N10776, N145, N9516);
and AND4 (N10795, N10761, N663, N964, N9084);
not NOT1 (N10796, N10795);
buf BUF1 (N10797, N10796);
nand NAND2 (N10798, N10794, N4993);
or OR4 (N10799, N10787, N8185, N5825, N7203);
buf BUF1 (N10800, N10797);
and AND2 (N10801, N10789, N7190);
nand NAND4 (N10802, N10792, N2595, N4761, N4478);
buf BUF1 (N10803, N10802);
nor NOR3 (N10804, N10803, N7873, N4259);
xor XOR2 (N10805, N10801, N9747);
and AND4 (N10806, N10800, N4922, N7632, N7841);
nand NAND4 (N10807, N10798, N4852, N10418, N7461);
or OR2 (N10808, N10799, N7370);
nand NAND3 (N10809, N10773, N10238, N3938);
not NOT1 (N10810, N10791);
xor XOR2 (N10811, N10793, N6789);
not NOT1 (N10812, N10805);
xor XOR2 (N10813, N10811, N7870);
nand NAND2 (N10814, N10788, N8075);
nand NAND3 (N10815, N10807, N2550, N10114);
not NOT1 (N10816, N10810);
xor XOR2 (N10817, N10772, N8655);
buf BUF1 (N10818, N10812);
xor XOR2 (N10819, N10816, N2139);
buf BUF1 (N10820, N10813);
nor NOR3 (N10821, N10817, N285, N9943);
or OR3 (N10822, N10820, N6483, N10259);
nand NAND2 (N10823, N10819, N7422);
buf BUF1 (N10824, N10815);
nand NAND4 (N10825, N10822, N8667, N1429, N10132);
xor XOR2 (N10826, N10809, N1130);
xor XOR2 (N10827, N10821, N5339);
and AND2 (N10828, N10814, N5437);
nand NAND4 (N10829, N10806, N1243, N4952, N2947);
nor NOR4 (N10830, N10829, N5490, N3786, N9483);
nor NOR3 (N10831, N10804, N5273, N627);
and AND4 (N10832, N10823, N6951, N6462, N10062);
or OR4 (N10833, N10831, N5114, N10518, N10016);
or OR2 (N10834, N10825, N6091);
nor NOR2 (N10835, N10833, N8676);
and AND3 (N10836, N10824, N10079, N3316);
buf BUF1 (N10837, N10828);
and AND4 (N10838, N10830, N9263, N8444, N6510);
or OR2 (N10839, N10818, N6149);
or OR3 (N10840, N10836, N9258, N8837);
nand NAND4 (N10841, N10808, N8937, N9098, N5632);
buf BUF1 (N10842, N10832);
nand NAND4 (N10843, N10842, N394, N4527, N5263);
not NOT1 (N10844, N10835);
buf BUF1 (N10845, N10841);
and AND4 (N10846, N10844, N3807, N5933, N10822);
xor XOR2 (N10847, N10839, N419);
nor NOR4 (N10848, N10845, N2419, N10528, N8831);
not NOT1 (N10849, N10837);
or OR2 (N10850, N10849, N4294);
nor NOR3 (N10851, N10840, N4517, N2101);
buf BUF1 (N10852, N10834);
buf BUF1 (N10853, N10850);
not NOT1 (N10854, N10846);
nor NOR3 (N10855, N10826, N2899, N6696);
nor NOR4 (N10856, N10847, N4436, N1665, N6499);
or OR4 (N10857, N10853, N3228, N142, N1943);
nand NAND4 (N10858, N10848, N1558, N1933, N4975);
and AND4 (N10859, N10857, N8559, N550, N7258);
nand NAND2 (N10860, N10852, N10302);
nor NOR3 (N10861, N10858, N1337, N10557);
buf BUF1 (N10862, N10854);
and AND4 (N10863, N10838, N4539, N6817, N10012);
or OR2 (N10864, N10861, N10633);
and AND4 (N10865, N10864, N3261, N4343, N4137);
nor NOR4 (N10866, N10862, N9141, N8430, N5550);
nor NOR3 (N10867, N10856, N10063, N1369);
and AND2 (N10868, N10863, N10050);
or OR4 (N10869, N10860, N509, N3025, N9006);
or OR4 (N10870, N10869, N8616, N5583, N3087);
xor XOR2 (N10871, N10859, N7028);
nand NAND4 (N10872, N10867, N1282, N2685, N865);
not NOT1 (N10873, N10855);
xor XOR2 (N10874, N10851, N1837);
xor XOR2 (N10875, N10868, N8182);
not NOT1 (N10876, N10870);
not NOT1 (N10877, N10875);
nand NAND2 (N10878, N10866, N979);
nor NOR3 (N10879, N10878, N10227, N3430);
nor NOR3 (N10880, N10874, N3916, N5511);
and AND2 (N10881, N10827, N1489);
not NOT1 (N10882, N10843);
not NOT1 (N10883, N10882);
buf BUF1 (N10884, N10876);
or OR2 (N10885, N10880, N10504);
nand NAND2 (N10886, N10872, N8928);
nand NAND2 (N10887, N10885, N7562);
not NOT1 (N10888, N10873);
not NOT1 (N10889, N10883);
nor NOR4 (N10890, N10879, N881, N2660, N6081);
buf BUF1 (N10891, N10888);
nor NOR4 (N10892, N10865, N10093, N2636, N5549);
nor NOR3 (N10893, N10890, N7297, N10765);
buf BUF1 (N10894, N10886);
xor XOR2 (N10895, N10881, N4677);
xor XOR2 (N10896, N10893, N3316);
and AND3 (N10897, N10877, N1001, N10605);
and AND3 (N10898, N10896, N8389, N9705);
not NOT1 (N10899, N10889);
nand NAND4 (N10900, N10892, N10216, N1516, N6145);
not NOT1 (N10901, N10884);
or OR3 (N10902, N10901, N5238, N4194);
buf BUF1 (N10903, N10894);
nor NOR2 (N10904, N10900, N1211);
and AND3 (N10905, N10898, N4043, N6213);
not NOT1 (N10906, N10897);
and AND2 (N10907, N10903, N10420);
xor XOR2 (N10908, N10905, N7858);
nand NAND3 (N10909, N10908, N172, N4847);
not NOT1 (N10910, N10899);
and AND3 (N10911, N10907, N9572, N10088);
nand NAND4 (N10912, N10904, N4939, N8381, N4912);
nor NOR3 (N10913, N10911, N2303, N2464);
nand NAND4 (N10914, N10887, N7926, N40, N7210);
nand NAND3 (N10915, N10913, N9027, N2579);
xor XOR2 (N10916, N10914, N4554);
buf BUF1 (N10917, N10912);
xor XOR2 (N10918, N10906, N2660);
buf BUF1 (N10919, N10915);
xor XOR2 (N10920, N10919, N1873);
nand NAND2 (N10921, N10895, N5284);
nor NOR4 (N10922, N10909, N8141, N6602, N4068);
nand NAND2 (N10923, N10920, N646);
xor XOR2 (N10924, N10871, N9955);
or OR4 (N10925, N10924, N9773, N7426, N10146);
not NOT1 (N10926, N10918);
not NOT1 (N10927, N10922);
nand NAND3 (N10928, N10927, N3935, N2635);
xor XOR2 (N10929, N10917, N674);
nor NOR2 (N10930, N10926, N7195);
or OR3 (N10931, N10921, N1645, N8713);
or OR2 (N10932, N10931, N7682);
buf BUF1 (N10933, N10923);
not NOT1 (N10934, N10925);
not NOT1 (N10935, N10902);
not NOT1 (N10936, N10934);
nor NOR4 (N10937, N10928, N9925, N9028, N1377);
nor NOR3 (N10938, N10937, N9933, N7777);
nand NAND4 (N10939, N10935, N4271, N6589, N9465);
not NOT1 (N10940, N10916);
or OR4 (N10941, N10930, N10467, N355, N10286);
or OR3 (N10942, N10941, N1891, N2293);
xor XOR2 (N10943, N10932, N28);
nand NAND2 (N10944, N10933, N4442);
nand NAND2 (N10945, N10940, N10529);
or OR2 (N10946, N10938, N639);
not NOT1 (N10947, N10910);
nor NOR4 (N10948, N10891, N2885, N9575, N9043);
buf BUF1 (N10949, N10936);
not NOT1 (N10950, N10942);
not NOT1 (N10951, N10948);
xor XOR2 (N10952, N10947, N2196);
xor XOR2 (N10953, N10952, N9720);
nor NOR4 (N10954, N10944, N4931, N10215, N9861);
nand NAND4 (N10955, N10946, N6097, N2916, N2054);
nand NAND4 (N10956, N10950, N4067, N68, N4955);
xor XOR2 (N10957, N10939, N6856);
xor XOR2 (N10958, N10943, N6222);
and AND3 (N10959, N10929, N7989, N4396);
or OR3 (N10960, N10954, N3772, N8416);
not NOT1 (N10961, N10957);
not NOT1 (N10962, N10958);
and AND3 (N10963, N10960, N19, N3931);
buf BUF1 (N10964, N10953);
nand NAND4 (N10965, N10951, N6080, N2459, N6419);
buf BUF1 (N10966, N10965);
buf BUF1 (N10967, N10955);
not NOT1 (N10968, N10961);
nand NAND4 (N10969, N10964, N3028, N6254, N4018);
and AND3 (N10970, N10966, N1840, N3609);
nor NOR3 (N10971, N10962, N1606, N5254);
xor XOR2 (N10972, N10949, N2313);
buf BUF1 (N10973, N10969);
and AND4 (N10974, N10973, N3020, N6317, N8323);
nand NAND2 (N10975, N10972, N6120);
nand NAND4 (N10976, N10974, N5029, N2755, N1903);
nand NAND2 (N10977, N10975, N7288);
nand NAND2 (N10978, N10956, N2701);
buf BUF1 (N10979, N10959);
nor NOR2 (N10980, N10967, N6016);
and AND4 (N10981, N10968, N5121, N6968, N9402);
nand NAND3 (N10982, N10976, N1813, N1135);
nand NAND4 (N10983, N10979, N10430, N1673, N8733);
and AND2 (N10984, N10982, N9832);
and AND3 (N10985, N10983, N6801, N7973);
nor NOR3 (N10986, N10978, N4863, N682);
and AND4 (N10987, N10970, N3154, N10724, N2338);
nand NAND2 (N10988, N10987, N4229);
nand NAND3 (N10989, N10985, N4278, N6887);
nor NOR3 (N10990, N10977, N4207, N9590);
buf BUF1 (N10991, N10986);
and AND4 (N10992, N10963, N8360, N6355, N2590);
nor NOR4 (N10993, N10980, N9427, N6603, N6776);
buf BUF1 (N10994, N10988);
nor NOR4 (N10995, N10994, N10820, N8308, N9129);
nand NAND4 (N10996, N10993, N8139, N9224, N652);
or OR3 (N10997, N10991, N31, N3752);
not NOT1 (N10998, N10989);
xor XOR2 (N10999, N10984, N308);
or OR4 (N11000, N10997, N10350, N9242, N4999);
nor NOR4 (N11001, N10995, N2637, N10204, N1242);
not NOT1 (N11002, N11001);
buf BUF1 (N11003, N10992);
not NOT1 (N11004, N10990);
and AND3 (N11005, N10998, N6887, N5143);
nand NAND4 (N11006, N11002, N5, N8843, N3495);
nor NOR4 (N11007, N11003, N10841, N3351, N7321);
buf BUF1 (N11008, N10996);
xor XOR2 (N11009, N11007, N3362);
nand NAND2 (N11010, N10945, N2358);
nand NAND3 (N11011, N11008, N10779, N7650);
nand NAND2 (N11012, N11005, N9144);
and AND4 (N11013, N11006, N3887, N6272, N10319);
or OR4 (N11014, N10981, N6335, N10639, N1669);
xor XOR2 (N11015, N10999, N8802);
or OR4 (N11016, N11010, N8306, N565, N4687);
buf BUF1 (N11017, N11011);
nor NOR2 (N11018, N11000, N2231);
not NOT1 (N11019, N11009);
or OR3 (N11020, N11017, N3380, N4348);
nand NAND4 (N11021, N11019, N3638, N3772, N773);
nor NOR2 (N11022, N11020, N5690);
xor XOR2 (N11023, N11013, N3788);
not NOT1 (N11024, N11014);
xor XOR2 (N11025, N11018, N9640);
not NOT1 (N11026, N11025);
not NOT1 (N11027, N11022);
xor XOR2 (N11028, N11004, N5309);
not NOT1 (N11029, N10971);
xor XOR2 (N11030, N11021, N7040);
nand NAND3 (N11031, N11023, N9245, N7902);
nor NOR4 (N11032, N11028, N5619, N5194, N6433);
buf BUF1 (N11033, N11012);
buf BUF1 (N11034, N11032);
nand NAND3 (N11035, N11031, N8156, N3082);
nand NAND4 (N11036, N11030, N6946, N8116, N5670);
nand NAND3 (N11037, N11024, N8359, N5497);
nor NOR2 (N11038, N11026, N31);
xor XOR2 (N11039, N11029, N5656);
or OR3 (N11040, N11039, N8505, N2027);
nor NOR2 (N11041, N11038, N4998);
not NOT1 (N11042, N11034);
not NOT1 (N11043, N11037);
and AND4 (N11044, N11040, N1577, N7321, N10542);
not NOT1 (N11045, N11015);
xor XOR2 (N11046, N11027, N3492);
not NOT1 (N11047, N11045);
nor NOR2 (N11048, N11047, N2115);
nand NAND3 (N11049, N11035, N9850, N856);
nor NOR4 (N11050, N11016, N3828, N6071, N7574);
buf BUF1 (N11051, N11042);
nand NAND4 (N11052, N11050, N8582, N769, N5719);
nor NOR3 (N11053, N11051, N9380, N367);
or OR4 (N11054, N11053, N5078, N6656, N7777);
xor XOR2 (N11055, N11036, N6085);
xor XOR2 (N11056, N11054, N5030);
or OR4 (N11057, N11052, N8304, N9191, N327);
or OR2 (N11058, N11046, N1771);
buf BUF1 (N11059, N11058);
and AND3 (N11060, N11044, N6422, N1967);
buf BUF1 (N11061, N11033);
xor XOR2 (N11062, N11061, N1734);
nor NOR4 (N11063, N11043, N2066, N6564, N6650);
buf BUF1 (N11064, N11059);
not NOT1 (N11065, N11057);
not NOT1 (N11066, N11041);
xor XOR2 (N11067, N11066, N10787);
or OR4 (N11068, N11064, N4320, N2991, N7973);
not NOT1 (N11069, N11060);
not NOT1 (N11070, N11063);
xor XOR2 (N11071, N11070, N3043);
buf BUF1 (N11072, N11065);
nor NOR4 (N11073, N11055, N9510, N3598, N8844);
nor NOR3 (N11074, N11067, N1449, N4807);
or OR4 (N11075, N11069, N7304, N4022, N9161);
and AND3 (N11076, N11075, N824, N4851);
buf BUF1 (N11077, N11074);
nor NOR4 (N11078, N11072, N7527, N9824, N10816);
and AND2 (N11079, N11071, N10395);
nor NOR4 (N11080, N11056, N2725, N4456, N5071);
nand NAND2 (N11081, N11068, N4643);
and AND4 (N11082, N11062, N3645, N9778, N10452);
and AND3 (N11083, N11082, N3149, N3190);
or OR2 (N11084, N11078, N7261);
or OR2 (N11085, N11084, N4240);
or OR4 (N11086, N11085, N10847, N10617, N6752);
and AND3 (N11087, N11077, N10105, N1509);
and AND4 (N11088, N11080, N7569, N176, N7257);
buf BUF1 (N11089, N11076);
buf BUF1 (N11090, N11049);
or OR3 (N11091, N11087, N1803, N6909);
and AND3 (N11092, N11081, N550, N9361);
nand NAND3 (N11093, N11091, N5059, N3316);
xor XOR2 (N11094, N11090, N10628);
or OR2 (N11095, N11086, N9115);
xor XOR2 (N11096, N11079, N3500);
or OR3 (N11097, N11088, N4979, N4696);
buf BUF1 (N11098, N11096);
nand NAND3 (N11099, N11083, N10151, N6944);
nor NOR4 (N11100, N11048, N10639, N10488, N9607);
and AND2 (N11101, N11095, N4348);
xor XOR2 (N11102, N11098, N9427);
xor XOR2 (N11103, N11102, N2080);
nand NAND2 (N11104, N11100, N10557);
or OR4 (N11105, N11099, N1990, N9632, N3249);
not NOT1 (N11106, N11105);
and AND4 (N11107, N11094, N6123, N7840, N665);
and AND3 (N11108, N11089, N4773, N3356);
nor NOR2 (N11109, N11101, N5149);
and AND4 (N11110, N11107, N8039, N2577, N5042);
nor NOR3 (N11111, N11110, N513, N629);
xor XOR2 (N11112, N11109, N5962);
and AND2 (N11113, N11111, N4763);
not NOT1 (N11114, N11073);
nor NOR4 (N11115, N11104, N9539, N9673, N5623);
and AND4 (N11116, N11113, N4802, N8588, N5773);
not NOT1 (N11117, N11116);
buf BUF1 (N11118, N11106);
nand NAND4 (N11119, N11112, N7920, N3387, N2312);
xor XOR2 (N11120, N11093, N1853);
nand NAND2 (N11121, N11120, N10713);
nor NOR3 (N11122, N11117, N9614, N658);
or OR2 (N11123, N11108, N10398);
not NOT1 (N11124, N11123);
buf BUF1 (N11125, N11124);
not NOT1 (N11126, N11092);
buf BUF1 (N11127, N11103);
and AND2 (N11128, N11121, N5600);
or OR2 (N11129, N11097, N7090);
or OR4 (N11130, N11129, N2356, N4527, N2915);
xor XOR2 (N11131, N11126, N6346);
nor NOR3 (N11132, N11122, N7630, N8046);
buf BUF1 (N11133, N11128);
xor XOR2 (N11134, N11125, N10329);
not NOT1 (N11135, N11131);
or OR3 (N11136, N11135, N9391, N6388);
buf BUF1 (N11137, N11127);
and AND3 (N11138, N11133, N2887, N10268);
not NOT1 (N11139, N11137);
nor NOR2 (N11140, N11119, N4896);
xor XOR2 (N11141, N11130, N10329);
or OR4 (N11142, N11132, N5961, N4098, N420);
xor XOR2 (N11143, N11115, N4545);
and AND4 (N11144, N11134, N7504, N8178, N6449);
nor NOR3 (N11145, N11114, N6166, N3170);
or OR4 (N11146, N11136, N3911, N744, N2589);
nand NAND2 (N11147, N11146, N8313);
not NOT1 (N11148, N11139);
nand NAND3 (N11149, N11141, N6151, N5104);
xor XOR2 (N11150, N11149, N2836);
nor NOR2 (N11151, N11147, N3784);
or OR3 (N11152, N11143, N10845, N4606);
and AND2 (N11153, N11150, N1964);
not NOT1 (N11154, N11144);
or OR3 (N11155, N11138, N4864, N8858);
buf BUF1 (N11156, N11148);
nor NOR2 (N11157, N11142, N7870);
or OR3 (N11158, N11157, N3376, N5022);
or OR3 (N11159, N11158, N2067, N6962);
nand NAND2 (N11160, N11145, N4738);
not NOT1 (N11161, N11140);
not NOT1 (N11162, N11156);
and AND2 (N11163, N11151, N10690);
or OR4 (N11164, N11155, N6501, N7486, N5540);
nand NAND2 (N11165, N11154, N10342);
nor NOR4 (N11166, N11161, N3733, N10882, N1377);
nand NAND2 (N11167, N11166, N8150);
or OR4 (N11168, N11162, N7144, N6412, N5356);
or OR4 (N11169, N11168, N10639, N1552, N7735);
nand NAND2 (N11170, N11169, N7692);
nand NAND4 (N11171, N11152, N3214, N2155, N7427);
nand NAND2 (N11172, N11160, N904);
and AND4 (N11173, N11172, N6691, N9519, N7534);
or OR4 (N11174, N11164, N3493, N254, N5991);
nand NAND4 (N11175, N11153, N7695, N5853, N5279);
xor XOR2 (N11176, N11173, N5105);
xor XOR2 (N11177, N11163, N2042);
xor XOR2 (N11178, N11176, N6461);
xor XOR2 (N11179, N11170, N9963);
nor NOR4 (N11180, N11179, N4523, N5290, N8327);
nor NOR3 (N11181, N11180, N9489, N2576);
or OR2 (N11182, N11159, N10542);
not NOT1 (N11183, N11165);
or OR3 (N11184, N11175, N4642, N2917);
or OR2 (N11185, N11183, N5162);
not NOT1 (N11186, N11174);
and AND4 (N11187, N11167, N3717, N7053, N1452);
nor NOR2 (N11188, N11187, N10914);
or OR4 (N11189, N11177, N2767, N3745, N1686);
and AND2 (N11190, N11171, N1840);
xor XOR2 (N11191, N11185, N3010);
or OR3 (N11192, N11188, N5419, N8480);
xor XOR2 (N11193, N11118, N1769);
nor NOR4 (N11194, N11181, N2733, N6412, N365);
and AND4 (N11195, N11182, N4698, N9882, N1371);
and AND2 (N11196, N11192, N10981);
and AND3 (N11197, N11178, N6830, N4315);
not NOT1 (N11198, N11194);
not NOT1 (N11199, N11189);
nor NOR4 (N11200, N11190, N1148, N330, N10708);
not NOT1 (N11201, N11195);
or OR4 (N11202, N11196, N5062, N7755, N1419);
buf BUF1 (N11203, N11191);
buf BUF1 (N11204, N11203);
xor XOR2 (N11205, N11198, N9502);
not NOT1 (N11206, N11200);
and AND2 (N11207, N11206, N4890);
xor XOR2 (N11208, N11202, N6697);
and AND3 (N11209, N11208, N9694, N4740);
nor NOR3 (N11210, N11197, N5669, N4955);
and AND2 (N11211, N11204, N2985);
nor NOR2 (N11212, N11207, N7018);
or OR3 (N11213, N11212, N6691, N9293);
nor NOR3 (N11214, N11211, N4783, N10022);
not NOT1 (N11215, N11193);
nand NAND3 (N11216, N11184, N123, N10558);
nor NOR2 (N11217, N11201, N1452);
xor XOR2 (N11218, N11214, N7190);
nor NOR4 (N11219, N11218, N2589, N7573, N4539);
and AND2 (N11220, N11219, N4666);
buf BUF1 (N11221, N11213);
nor NOR3 (N11222, N11216, N4656, N1003);
nand NAND4 (N11223, N11215, N6061, N6824, N10462);
xor XOR2 (N11224, N11220, N10569);
buf BUF1 (N11225, N11221);
buf BUF1 (N11226, N11217);
nand NAND2 (N11227, N11223, N690);
nor NOR4 (N11228, N11227, N215, N983, N3646);
xor XOR2 (N11229, N11210, N5839);
nand NAND2 (N11230, N11228, N8122);
and AND3 (N11231, N11224, N1285, N8429);
nor NOR2 (N11232, N11222, N9179);
not NOT1 (N11233, N11205);
nand NAND4 (N11234, N11186, N460, N4471, N6469);
and AND2 (N11235, N11229, N8275);
and AND2 (N11236, N11230, N7259);
buf BUF1 (N11237, N11209);
and AND2 (N11238, N11231, N5791);
buf BUF1 (N11239, N11232);
or OR3 (N11240, N11225, N8320, N192);
or OR3 (N11241, N11226, N8961, N6126);
and AND4 (N11242, N11199, N11069, N5030, N4505);
not NOT1 (N11243, N11233);
or OR3 (N11244, N11238, N2101, N7352);
and AND2 (N11245, N11235, N11020);
nor NOR3 (N11246, N11236, N3193, N8338);
buf BUF1 (N11247, N11237);
xor XOR2 (N11248, N11244, N5883);
and AND4 (N11249, N11242, N5249, N3412, N9618);
nor NOR3 (N11250, N11239, N5751, N1587);
nand NAND3 (N11251, N11234, N4643, N4538);
xor XOR2 (N11252, N11250, N2807);
xor XOR2 (N11253, N11240, N8741);
nor NOR4 (N11254, N11253, N4386, N5726, N290);
nand NAND3 (N11255, N11248, N5241, N8182);
nand NAND2 (N11256, N11252, N4990);
buf BUF1 (N11257, N11249);
and AND2 (N11258, N11246, N4746);
buf BUF1 (N11259, N11255);
nand NAND3 (N11260, N11259, N457, N9875);
not NOT1 (N11261, N11245);
nor NOR2 (N11262, N11254, N435);
nand NAND3 (N11263, N11262, N11220, N11032);
nor NOR2 (N11264, N11241, N10975);
nand NAND3 (N11265, N11247, N6723, N3477);
nand NAND3 (N11266, N11265, N1097, N7386);
buf BUF1 (N11267, N11256);
xor XOR2 (N11268, N11243, N9099);
or OR3 (N11269, N11264, N5168, N7600);
xor XOR2 (N11270, N11266, N7012);
buf BUF1 (N11271, N11268);
not NOT1 (N11272, N11257);
nor NOR4 (N11273, N11263, N4368, N9552, N1039);
not NOT1 (N11274, N11261);
nand NAND4 (N11275, N11270, N7388, N3194, N2909);
nor NOR2 (N11276, N11269, N1372);
xor XOR2 (N11277, N11271, N8680);
xor XOR2 (N11278, N11251, N5280);
or OR3 (N11279, N11273, N3629, N5944);
buf BUF1 (N11280, N11276);
buf BUF1 (N11281, N11278);
not NOT1 (N11282, N11275);
nor NOR2 (N11283, N11267, N8200);
nand NAND3 (N11284, N11274, N10023, N6249);
and AND3 (N11285, N11258, N9507, N2264);
nand NAND3 (N11286, N11280, N428, N4496);
not NOT1 (N11287, N11272);
buf BUF1 (N11288, N11283);
xor XOR2 (N11289, N11284, N10563);
nor NOR4 (N11290, N11260, N608, N1135, N10239);
nor NOR3 (N11291, N11281, N4881, N8168);
or OR2 (N11292, N11286, N7176);
and AND4 (N11293, N11292, N3070, N6064, N9334);
nand NAND2 (N11294, N11291, N822);
buf BUF1 (N11295, N11285);
xor XOR2 (N11296, N11279, N9886);
xor XOR2 (N11297, N11282, N4217);
xor XOR2 (N11298, N11294, N2594);
nor NOR4 (N11299, N11290, N5013, N10930, N3788);
nor NOR2 (N11300, N11289, N9829);
and AND3 (N11301, N11300, N7488, N1668);
not NOT1 (N11302, N11297);
buf BUF1 (N11303, N11287);
nor NOR2 (N11304, N11301, N5882);
or OR2 (N11305, N11302, N5118);
and AND2 (N11306, N11295, N10950);
xor XOR2 (N11307, N11303, N4483);
xor XOR2 (N11308, N11306, N2120);
not NOT1 (N11309, N11305);
nor NOR4 (N11310, N11309, N300, N7521, N3132);
nand NAND3 (N11311, N11296, N7962, N8326);
and AND3 (N11312, N11311, N4862, N1198);
and AND2 (N11313, N11293, N10224);
and AND2 (N11314, N11288, N7304);
nand NAND2 (N11315, N11299, N8814);
not NOT1 (N11316, N11304);
xor XOR2 (N11317, N11315, N8166);
xor XOR2 (N11318, N11313, N9485);
nand NAND2 (N11319, N11318, N3730);
and AND2 (N11320, N11317, N589);
not NOT1 (N11321, N11310);
nand NAND2 (N11322, N11312, N7156);
buf BUF1 (N11323, N11322);
or OR4 (N11324, N11323, N8544, N8907, N4831);
or OR2 (N11325, N11307, N4956);
and AND4 (N11326, N11314, N9364, N10689, N9266);
and AND4 (N11327, N11326, N8642, N10056, N4940);
xor XOR2 (N11328, N11308, N5382);
not NOT1 (N11329, N11328);
or OR3 (N11330, N11329, N1961, N7672);
nand NAND2 (N11331, N11330, N8793);
or OR4 (N11332, N11319, N9468, N2748, N5305);
or OR2 (N11333, N11320, N5746);
not NOT1 (N11334, N11277);
buf BUF1 (N11335, N11331);
buf BUF1 (N11336, N11333);
nand NAND4 (N11337, N11334, N3569, N8351, N8173);
nand NAND3 (N11338, N11298, N338, N2862);
nand NAND4 (N11339, N11316, N9527, N10993, N4108);
nand NAND4 (N11340, N11321, N11052, N6407, N3298);
not NOT1 (N11341, N11335);
nor NOR3 (N11342, N11337, N4227, N9394);
buf BUF1 (N11343, N11341);
buf BUF1 (N11344, N11327);
or OR4 (N11345, N11332, N7775, N7527, N8940);
or OR4 (N11346, N11325, N6418, N172, N1867);
nor NOR4 (N11347, N11324, N3924, N3037, N6132);
nand NAND2 (N11348, N11342, N7854);
and AND3 (N11349, N11339, N8142, N10352);
nor NOR4 (N11350, N11340, N7525, N8634, N7194);
nor NOR4 (N11351, N11345, N7097, N5028, N1572);
nand NAND2 (N11352, N11347, N2252);
buf BUF1 (N11353, N11351);
buf BUF1 (N11354, N11350);
buf BUF1 (N11355, N11336);
xor XOR2 (N11356, N11344, N9658);
buf BUF1 (N11357, N11338);
and AND4 (N11358, N11352, N6970, N10268, N4841);
not NOT1 (N11359, N11356);
or OR3 (N11360, N11349, N511, N8339);
nand NAND3 (N11361, N11343, N4854, N161);
xor XOR2 (N11362, N11359, N6137);
nand NAND3 (N11363, N11357, N8465, N849);
and AND4 (N11364, N11354, N6181, N3856, N4883);
or OR4 (N11365, N11363, N9172, N6902, N3685);
nor NOR2 (N11366, N11348, N6982);
not NOT1 (N11367, N11365);
xor XOR2 (N11368, N11355, N7207);
xor XOR2 (N11369, N11367, N8726);
xor XOR2 (N11370, N11368, N9779);
nand NAND2 (N11371, N11353, N9061);
buf BUF1 (N11372, N11370);
and AND3 (N11373, N11362, N10077, N5208);
or OR3 (N11374, N11372, N11189, N3449);
and AND2 (N11375, N11358, N5583);
xor XOR2 (N11376, N11375, N1641);
and AND3 (N11377, N11376, N7804, N2591);
xor XOR2 (N11378, N11369, N8229);
xor XOR2 (N11379, N11361, N4371);
buf BUF1 (N11380, N11364);
and AND3 (N11381, N11346, N157, N11379);
not NOT1 (N11382, N8143);
nand NAND4 (N11383, N11373, N5569, N5006, N4159);
nand NAND3 (N11384, N11382, N6091, N10934);
buf BUF1 (N11385, N11371);
not NOT1 (N11386, N11360);
nand NAND2 (N11387, N11381, N3973);
not NOT1 (N11388, N11374);
xor XOR2 (N11389, N11366, N107);
and AND2 (N11390, N11383, N6142);
and AND4 (N11391, N11389, N7122, N5112, N1747);
nor NOR3 (N11392, N11380, N9138, N3426);
and AND3 (N11393, N11391, N5884, N8114);
xor XOR2 (N11394, N11384, N6877);
buf BUF1 (N11395, N11392);
buf BUF1 (N11396, N11393);
xor XOR2 (N11397, N11395, N7405);
nand NAND4 (N11398, N11390, N3344, N3260, N9859);
not NOT1 (N11399, N11398);
buf BUF1 (N11400, N11396);
or OR2 (N11401, N11388, N8572);
nand NAND2 (N11402, N11401, N4081);
and AND2 (N11403, N11400, N3040);
buf BUF1 (N11404, N11387);
and AND3 (N11405, N11397, N6501, N3791);
buf BUF1 (N11406, N11405);
nor NOR4 (N11407, N11394, N7060, N5684, N4633);
and AND3 (N11408, N11406, N6621, N8290);
nor NOR4 (N11409, N11378, N10786, N4365, N1334);
and AND3 (N11410, N11385, N1660, N10517);
buf BUF1 (N11411, N11399);
nand NAND2 (N11412, N11411, N11206);
buf BUF1 (N11413, N11402);
or OR2 (N11414, N11403, N6652);
or OR3 (N11415, N11386, N9139, N2420);
nor NOR2 (N11416, N11410, N13);
xor XOR2 (N11417, N11412, N5503);
or OR4 (N11418, N11413, N6300, N9523, N1757);
and AND3 (N11419, N11416, N9949, N8899);
or OR3 (N11420, N11414, N5672, N6502);
xor XOR2 (N11421, N11415, N9793);
nand NAND3 (N11422, N11407, N8909, N10319);
not NOT1 (N11423, N11420);
not NOT1 (N11424, N11417);
nor NOR2 (N11425, N11421, N2916);
and AND3 (N11426, N11424, N1037, N2);
xor XOR2 (N11427, N11408, N5772);
nor NOR4 (N11428, N11426, N58, N6009, N2871);
and AND2 (N11429, N11428, N5666);
buf BUF1 (N11430, N11427);
xor XOR2 (N11431, N11419, N4158);
buf BUF1 (N11432, N11418);
buf BUF1 (N11433, N11430);
nand NAND3 (N11434, N11422, N4214, N4565);
nand NAND2 (N11435, N11425, N501);
nor NOR3 (N11436, N11429, N166, N9363);
nor NOR2 (N11437, N11409, N10630);
buf BUF1 (N11438, N11423);
not NOT1 (N11439, N11433);
xor XOR2 (N11440, N11431, N3647);
nor NOR4 (N11441, N11436, N7685, N1580, N7330);
nor NOR2 (N11442, N11432, N10393);
xor XOR2 (N11443, N11439, N8694);
not NOT1 (N11444, N11377);
and AND4 (N11445, N11443, N7830, N2574, N3421);
nor NOR3 (N11446, N11404, N4725, N6744);
or OR4 (N11447, N11440, N10614, N6879, N11411);
buf BUF1 (N11448, N11447);
buf BUF1 (N11449, N11434);
and AND2 (N11450, N11442, N4037);
nor NOR3 (N11451, N11446, N7878, N6977);
or OR4 (N11452, N11441, N7532, N3000, N3730);
not NOT1 (N11453, N11435);
not NOT1 (N11454, N11444);
buf BUF1 (N11455, N11438);
nand NAND2 (N11456, N11449, N904);
xor XOR2 (N11457, N11454, N4631);
buf BUF1 (N11458, N11437);
nand NAND2 (N11459, N11445, N1341);
not NOT1 (N11460, N11455);
not NOT1 (N11461, N11453);
and AND2 (N11462, N11456, N9392);
nor NOR4 (N11463, N11451, N601, N8795, N5020);
nor NOR2 (N11464, N11459, N3109);
not NOT1 (N11465, N11464);
not NOT1 (N11466, N11448);
and AND2 (N11467, N11466, N8119);
and AND2 (N11468, N11458, N9442);
xor XOR2 (N11469, N11450, N4086);
nand NAND3 (N11470, N11465, N4050, N7330);
and AND3 (N11471, N11469, N2619, N5673);
or OR3 (N11472, N11470, N1288, N5539);
nand NAND4 (N11473, N11471, N1317, N132, N11120);
buf BUF1 (N11474, N11461);
and AND4 (N11475, N11457, N3355, N3340, N3559);
buf BUF1 (N11476, N11460);
nand NAND4 (N11477, N11467, N7989, N8424, N276);
or OR3 (N11478, N11452, N5888, N9394);
or OR4 (N11479, N11478, N6003, N54, N8404);
and AND2 (N11480, N11472, N9795);
nor NOR3 (N11481, N11463, N7145, N10313);
or OR3 (N11482, N11475, N3261, N5335);
nor NOR3 (N11483, N11479, N5338, N9874);
buf BUF1 (N11484, N11483);
nor NOR3 (N11485, N11480, N571, N401);
xor XOR2 (N11486, N11468, N2425);
nor NOR2 (N11487, N11485, N7933);
and AND2 (N11488, N11476, N10359);
buf BUF1 (N11489, N11486);
buf BUF1 (N11490, N11481);
not NOT1 (N11491, N11473);
or OR2 (N11492, N11488, N7577);
nor NOR2 (N11493, N11491, N1176);
not NOT1 (N11494, N11484);
and AND3 (N11495, N11482, N5284, N317);
nor NOR2 (N11496, N11493, N2916);
xor XOR2 (N11497, N11494, N8451);
xor XOR2 (N11498, N11489, N213);
not NOT1 (N11499, N11496);
nor NOR3 (N11500, N11477, N4652, N661);
not NOT1 (N11501, N11500);
not NOT1 (N11502, N11462);
and AND3 (N11503, N11487, N9695, N8029);
buf BUF1 (N11504, N11474);
nor NOR3 (N11505, N11498, N4166, N5898);
not NOT1 (N11506, N11492);
buf BUF1 (N11507, N11495);
xor XOR2 (N11508, N11507, N2973);
nand NAND2 (N11509, N11497, N6350);
not NOT1 (N11510, N11509);
or OR3 (N11511, N11510, N910, N5307);
nor NOR4 (N11512, N11504, N847, N4067, N5718);
xor XOR2 (N11513, N11511, N8735);
not NOT1 (N11514, N11508);
and AND4 (N11515, N11512, N5233, N10667, N548);
nor NOR4 (N11516, N11501, N1092, N1503, N9205);
not NOT1 (N11517, N11499);
and AND2 (N11518, N11505, N6575);
and AND4 (N11519, N11502, N7401, N7883, N5294);
nand NAND4 (N11520, N11490, N9826, N11311, N2726);
nor NOR3 (N11521, N11514, N4464, N2838);
nand NAND2 (N11522, N11515, N4734);
nand NAND3 (N11523, N11518, N6176, N5768);
buf BUF1 (N11524, N11506);
nand NAND4 (N11525, N11513, N6318, N8767, N10935);
and AND3 (N11526, N11522, N4837, N1235);
buf BUF1 (N11527, N11517);
not NOT1 (N11528, N11526);
or OR3 (N11529, N11503, N913, N10063);
and AND3 (N11530, N11528, N800, N10047);
nor NOR2 (N11531, N11527, N4178);
xor XOR2 (N11532, N11529, N7083);
not NOT1 (N11533, N11521);
nor NOR3 (N11534, N11519, N3382, N9313);
and AND3 (N11535, N11530, N923, N10525);
nand NAND4 (N11536, N11531, N1035, N1124, N6222);
and AND4 (N11537, N11525, N9353, N4333, N6315);
not NOT1 (N11538, N11524);
nand NAND3 (N11539, N11538, N8182, N10953);
and AND3 (N11540, N11536, N2548, N10385);
not NOT1 (N11541, N11520);
buf BUF1 (N11542, N11540);
buf BUF1 (N11543, N11532);
nor NOR3 (N11544, N11533, N11211, N7753);
and AND3 (N11545, N11544, N2007, N5127);
nor NOR3 (N11546, N11534, N3281, N7365);
nand NAND4 (N11547, N11542, N7777, N9332, N10207);
xor XOR2 (N11548, N11537, N8333);
or OR4 (N11549, N11546, N758, N4248, N8923);
buf BUF1 (N11550, N11543);
not NOT1 (N11551, N11535);
or OR4 (N11552, N11523, N11550, N1144, N4478);
or OR4 (N11553, N7081, N6464, N604, N8983);
nor NOR2 (N11554, N11552, N11043);
buf BUF1 (N11555, N11547);
or OR4 (N11556, N11549, N7809, N9562, N9997);
not NOT1 (N11557, N11554);
xor XOR2 (N11558, N11516, N8856);
nor NOR2 (N11559, N11557, N8933);
or OR3 (N11560, N11559, N843, N8828);
nor NOR4 (N11561, N11541, N8078, N8368, N4807);
nand NAND2 (N11562, N11553, N2744);
not NOT1 (N11563, N11558);
nor NOR4 (N11564, N11548, N5406, N4483, N872);
buf BUF1 (N11565, N11561);
or OR3 (N11566, N11556, N2649, N8424);
xor XOR2 (N11567, N11551, N2852);
buf BUF1 (N11568, N11563);
and AND4 (N11569, N11555, N8127, N10878, N7821);
xor XOR2 (N11570, N11569, N5865);
nor NOR2 (N11571, N11560, N1743);
and AND2 (N11572, N11564, N8733);
nand NAND3 (N11573, N11539, N9142, N10842);
nor NOR4 (N11574, N11568, N848, N7584, N6677);
buf BUF1 (N11575, N11565);
not NOT1 (N11576, N11575);
xor XOR2 (N11577, N11566, N4484);
xor XOR2 (N11578, N11573, N9685);
nor NOR4 (N11579, N11578, N8997, N2832, N3703);
not NOT1 (N11580, N11574);
not NOT1 (N11581, N11571);
nor NOR3 (N11582, N11567, N4838, N3137);
xor XOR2 (N11583, N11577, N1662);
xor XOR2 (N11584, N11570, N5978);
and AND4 (N11585, N11579, N68, N9076, N7939);
nand NAND4 (N11586, N11584, N5136, N2115, N5018);
or OR2 (N11587, N11585, N403);
not NOT1 (N11588, N11583);
or OR4 (N11589, N11588, N11473, N9222, N6038);
nor NOR4 (N11590, N11562, N84, N1022, N4921);
or OR2 (N11591, N11590, N8475);
nor NOR3 (N11592, N11572, N10865, N8463);
and AND2 (N11593, N11581, N5026);
or OR2 (N11594, N11587, N683);
buf BUF1 (N11595, N11593);
nor NOR3 (N11596, N11595, N6313, N5911);
buf BUF1 (N11597, N11592);
buf BUF1 (N11598, N11586);
nand NAND4 (N11599, N11598, N11280, N9186, N4675);
nor NOR3 (N11600, N11545, N4391, N7796);
nor NOR2 (N11601, N11596, N60);
nand NAND3 (N11602, N11597, N3459, N8385);
nor NOR3 (N11603, N11594, N10881, N5671);
or OR4 (N11604, N11580, N10013, N560, N3227);
nor NOR2 (N11605, N11599, N4831);
not NOT1 (N11606, N11605);
or OR4 (N11607, N11591, N9196, N324, N9160);
and AND4 (N11608, N11582, N8658, N3326, N10640);
not NOT1 (N11609, N11601);
or OR2 (N11610, N11576, N7885);
xor XOR2 (N11611, N11600, N4618);
not NOT1 (N11612, N11602);
buf BUF1 (N11613, N11604);
and AND4 (N11614, N11609, N8459, N8900, N4016);
buf BUF1 (N11615, N11614);
not NOT1 (N11616, N11606);
and AND4 (N11617, N11616, N1870, N2369, N8717);
or OR3 (N11618, N11615, N7308, N6694);
xor XOR2 (N11619, N11607, N7464);
xor XOR2 (N11620, N11618, N6037);
nand NAND2 (N11621, N11589, N11318);
nand NAND3 (N11622, N11617, N4535, N5240);
or OR3 (N11623, N11612, N11405, N9299);
nor NOR2 (N11624, N11613, N3654);
nand NAND3 (N11625, N11611, N5688, N8902);
nor NOR4 (N11626, N11621, N2974, N3536, N2327);
or OR2 (N11627, N11625, N7896);
buf BUF1 (N11628, N11627);
not NOT1 (N11629, N11603);
not NOT1 (N11630, N11619);
buf BUF1 (N11631, N11628);
and AND4 (N11632, N11620, N5823, N3437, N1781);
nor NOR3 (N11633, N11626, N8672, N6272);
and AND2 (N11634, N11629, N7493);
xor XOR2 (N11635, N11610, N11397);
xor XOR2 (N11636, N11608, N4726);
nand NAND2 (N11637, N11632, N10994);
buf BUF1 (N11638, N11623);
buf BUF1 (N11639, N11633);
not NOT1 (N11640, N11634);
nand NAND3 (N11641, N11639, N2863, N10649);
nand NAND3 (N11642, N11624, N1384, N2065);
not NOT1 (N11643, N11631);
and AND2 (N11644, N11630, N10979);
not NOT1 (N11645, N11642);
xor XOR2 (N11646, N11645, N9045);
or OR4 (N11647, N11622, N10423, N9617, N7180);
or OR2 (N11648, N11641, N8688);
not NOT1 (N11649, N11640);
not NOT1 (N11650, N11648);
not NOT1 (N11651, N11649);
xor XOR2 (N11652, N11644, N11415);
not NOT1 (N11653, N11650);
buf BUF1 (N11654, N11651);
nor NOR4 (N11655, N11646, N3669, N4475, N5052);
not NOT1 (N11656, N11637);
nand NAND3 (N11657, N11655, N8193, N187);
xor XOR2 (N11658, N11656, N6871);
and AND4 (N11659, N11647, N10898, N10001, N293);
nor NOR2 (N11660, N11653, N10031);
buf BUF1 (N11661, N11659);
nand NAND2 (N11662, N11654, N6641);
xor XOR2 (N11663, N11658, N10401);
or OR2 (N11664, N11643, N2304);
and AND2 (N11665, N11636, N11555);
and AND3 (N11666, N11663, N8434, N4297);
nand NAND2 (N11667, N11660, N11015);
and AND2 (N11668, N11661, N9068);
not NOT1 (N11669, N11635);
nand NAND2 (N11670, N11669, N6222);
xor XOR2 (N11671, N11638, N8124);
not NOT1 (N11672, N11657);
or OR4 (N11673, N11670, N7083, N228, N7973);
nand NAND3 (N11674, N11666, N5209, N6340);
buf BUF1 (N11675, N11664);
nand NAND2 (N11676, N11674, N11291);
buf BUF1 (N11677, N11676);
and AND4 (N11678, N11671, N5575, N2535, N11078);
buf BUF1 (N11679, N11668);
not NOT1 (N11680, N11679);
or OR4 (N11681, N11667, N8992, N8372, N4379);
and AND4 (N11682, N11672, N619, N4469, N226);
xor XOR2 (N11683, N11678, N6853);
or OR2 (N11684, N11681, N6448);
nor NOR3 (N11685, N11677, N9280, N1378);
nand NAND3 (N11686, N11675, N10729, N6523);
or OR2 (N11687, N11682, N307);
nand NAND2 (N11688, N11680, N1049);
and AND4 (N11689, N11665, N1453, N3062, N9703);
nor NOR3 (N11690, N11684, N11169, N1245);
buf BUF1 (N11691, N11689);
or OR2 (N11692, N11686, N7955);
not NOT1 (N11693, N11692);
or OR3 (N11694, N11683, N298, N3496);
buf BUF1 (N11695, N11662);
not NOT1 (N11696, N11687);
buf BUF1 (N11697, N11691);
or OR3 (N11698, N11694, N3565, N2980);
not NOT1 (N11699, N11698);
and AND4 (N11700, N11685, N1566, N264, N980);
nand NAND3 (N11701, N11697, N7468, N3842);
nand NAND4 (N11702, N11690, N7646, N6920, N10747);
and AND2 (N11703, N11702, N5937);
xor XOR2 (N11704, N11673, N3593);
not NOT1 (N11705, N11688);
not NOT1 (N11706, N11703);
and AND2 (N11707, N11700, N2301);
or OR4 (N11708, N11696, N7841, N6711, N7568);
buf BUF1 (N11709, N11693);
not NOT1 (N11710, N11701);
xor XOR2 (N11711, N11704, N2574);
not NOT1 (N11712, N11699);
or OR2 (N11713, N11711, N3456);
buf BUF1 (N11714, N11709);
not NOT1 (N11715, N11706);
and AND4 (N11716, N11712, N8324, N2600, N1192);
not NOT1 (N11717, N11708);
not NOT1 (N11718, N11705);
buf BUF1 (N11719, N11717);
nor NOR3 (N11720, N11718, N3, N7707);
xor XOR2 (N11721, N11714, N10412);
and AND3 (N11722, N11715, N10631, N9058);
buf BUF1 (N11723, N11716);
nor NOR2 (N11724, N11710, N6015);
xor XOR2 (N11725, N11722, N3228);
buf BUF1 (N11726, N11721);
buf BUF1 (N11727, N11707);
xor XOR2 (N11728, N11723, N8345);
buf BUF1 (N11729, N11724);
or OR3 (N11730, N11726, N10238, N10682);
buf BUF1 (N11731, N11728);
nand NAND2 (N11732, N11731, N9600);
buf BUF1 (N11733, N11727);
nand NAND4 (N11734, N11713, N10670, N3173, N6792);
buf BUF1 (N11735, N11733);
and AND2 (N11736, N11729, N8786);
and AND2 (N11737, N11730, N8685);
or OR2 (N11738, N11695, N4999);
and AND2 (N11739, N11652, N7732);
nand NAND2 (N11740, N11732, N10434);
nor NOR3 (N11741, N11736, N5574, N5772);
or OR2 (N11742, N11741, N3263);
buf BUF1 (N11743, N11739);
xor XOR2 (N11744, N11735, N3224);
nor NOR4 (N11745, N11719, N6020, N7896, N5567);
nand NAND3 (N11746, N11737, N8267, N4092);
not NOT1 (N11747, N11725);
and AND3 (N11748, N11738, N9182, N4339);
and AND4 (N11749, N11734, N1766, N6845, N6067);
or OR3 (N11750, N11746, N7915, N3658);
xor XOR2 (N11751, N11748, N2626);
nor NOR4 (N11752, N11743, N6442, N11401, N5416);
nand NAND4 (N11753, N11745, N5572, N3426, N7820);
and AND4 (N11754, N11749, N7442, N11620, N6716);
nor NOR4 (N11755, N11754, N2623, N2061, N8891);
or OR2 (N11756, N11751, N1656);
buf BUF1 (N11757, N11740);
xor XOR2 (N11758, N11753, N9717);
xor XOR2 (N11759, N11747, N185);
and AND4 (N11760, N11757, N2456, N157, N5316);
xor XOR2 (N11761, N11750, N4940);
not NOT1 (N11762, N11755);
nor NOR3 (N11763, N11742, N10545, N11758);
or OR4 (N11764, N6093, N4311, N9325, N11448);
not NOT1 (N11765, N11752);
nand NAND3 (N11766, N11763, N8247, N399);
buf BUF1 (N11767, N11759);
and AND2 (N11768, N11765, N1771);
not NOT1 (N11769, N11762);
not NOT1 (N11770, N11769);
or OR4 (N11771, N11761, N11459, N6175, N10400);
nor NOR4 (N11772, N11771, N11736, N3678, N3375);
or OR4 (N11773, N11770, N10402, N8010, N5606);
nor NOR2 (N11774, N11744, N2485);
or OR4 (N11775, N11766, N1786, N8436, N6724);
buf BUF1 (N11776, N11774);
not NOT1 (N11777, N11760);
and AND2 (N11778, N11775, N7543);
xor XOR2 (N11779, N11720, N6812);
nor NOR3 (N11780, N11768, N10053, N11053);
xor XOR2 (N11781, N11777, N8346);
xor XOR2 (N11782, N11773, N6659);
nand NAND2 (N11783, N11767, N10550);
and AND4 (N11784, N11776, N398, N9043, N6015);
nand NAND2 (N11785, N11764, N11000);
nand NAND2 (N11786, N11779, N6012);
xor XOR2 (N11787, N11786, N5884);
and AND3 (N11788, N11778, N973, N842);
not NOT1 (N11789, N11787);
buf BUF1 (N11790, N11756);
and AND3 (N11791, N11790, N4928, N3059);
or OR2 (N11792, N11772, N2757);
nor NOR4 (N11793, N11788, N6224, N602, N10292);
not NOT1 (N11794, N11781);
not NOT1 (N11795, N11794);
buf BUF1 (N11796, N11782);
buf BUF1 (N11797, N11795);
and AND3 (N11798, N11783, N9064, N3377);
and AND2 (N11799, N11791, N10363);
nor NOR2 (N11800, N11793, N6765);
nand NAND3 (N11801, N11785, N4922, N8086);
or OR2 (N11802, N11789, N8735);
and AND2 (N11803, N11802, N2375);
xor XOR2 (N11804, N11800, N802);
nor NOR2 (N11805, N11804, N5625);
xor XOR2 (N11806, N11780, N4000);
buf BUF1 (N11807, N11806);
buf BUF1 (N11808, N11796);
xor XOR2 (N11809, N11808, N2003);
nor NOR3 (N11810, N11801, N3407, N6544);
or OR4 (N11811, N11799, N7115, N7893, N10221);
nor NOR2 (N11812, N11807, N3745);
and AND2 (N11813, N11797, N8359);
nor NOR2 (N11814, N11784, N751);
nor NOR3 (N11815, N11811, N955, N274);
buf BUF1 (N11816, N11803);
or OR2 (N11817, N11805, N6815);
nor NOR4 (N11818, N11816, N3792, N10049, N4562);
nand NAND3 (N11819, N11812, N2167, N10903);
buf BUF1 (N11820, N11819);
or OR3 (N11821, N11814, N3534, N4729);
xor XOR2 (N11822, N11817, N4903);
nor NOR4 (N11823, N11792, N7744, N5492, N9161);
and AND2 (N11824, N11815, N1420);
not NOT1 (N11825, N11810);
buf BUF1 (N11826, N11823);
xor XOR2 (N11827, N11821, N7084);
xor XOR2 (N11828, N11818, N6499);
not NOT1 (N11829, N11824);
xor XOR2 (N11830, N11825, N6175);
not NOT1 (N11831, N11826);
buf BUF1 (N11832, N11798);
nor NOR4 (N11833, N11809, N11752, N5690, N12);
and AND2 (N11834, N11820, N6410);
xor XOR2 (N11835, N11827, N2517);
not NOT1 (N11836, N11822);
and AND3 (N11837, N11830, N2585, N11791);
nand NAND3 (N11838, N11837, N10289, N10908);
buf BUF1 (N11839, N11835);
nor NOR4 (N11840, N11838, N2372, N1798, N9851);
nor NOR4 (N11841, N11829, N10899, N5441, N9381);
xor XOR2 (N11842, N11840, N7497);
nand NAND3 (N11843, N11831, N3120, N7759);
nand NAND2 (N11844, N11828, N9625);
not NOT1 (N11845, N11836);
nor NOR3 (N11846, N11833, N492, N10413);
and AND2 (N11847, N11846, N63);
not NOT1 (N11848, N11847);
nand NAND3 (N11849, N11813, N2286, N1829);
or OR3 (N11850, N11844, N5311, N11280);
or OR2 (N11851, N11843, N6006);
buf BUF1 (N11852, N11850);
nor NOR3 (N11853, N11851, N8559, N1294);
not NOT1 (N11854, N11852);
xor XOR2 (N11855, N11854, N7747);
and AND2 (N11856, N11832, N5759);
nor NOR3 (N11857, N11848, N3365, N11313);
and AND4 (N11858, N11841, N3789, N9595, N5366);
and AND2 (N11859, N11857, N6176);
and AND4 (N11860, N11849, N6456, N8030, N10154);
xor XOR2 (N11861, N11859, N6836);
nor NOR2 (N11862, N11842, N9951);
or OR4 (N11863, N11856, N9982, N3999, N1849);
buf BUF1 (N11864, N11853);
nor NOR3 (N11865, N11834, N885, N11256);
buf BUF1 (N11866, N11861);
nand NAND4 (N11867, N11860, N11284, N7900, N4016);
nor NOR4 (N11868, N11858, N1597, N2780, N3621);
nor NOR2 (N11869, N11865, N11682);
nand NAND3 (N11870, N11867, N100, N4131);
xor XOR2 (N11871, N11866, N8329);
xor XOR2 (N11872, N11871, N2517);
xor XOR2 (N11873, N11870, N9474);
or OR4 (N11874, N11862, N4687, N5575, N2892);
or OR3 (N11875, N11839, N6372, N1125);
and AND4 (N11876, N11869, N2151, N8537, N1913);
buf BUF1 (N11877, N11855);
nor NOR4 (N11878, N11864, N916, N2718, N10427);
nand NAND3 (N11879, N11875, N4264, N6018);
nand NAND2 (N11880, N11879, N10855);
and AND4 (N11881, N11873, N875, N2489, N3426);
and AND4 (N11882, N11845, N3224, N7126, N11759);
nand NAND4 (N11883, N11874, N2494, N6428, N2567);
nand NAND4 (N11884, N11881, N11153, N4038, N11729);
or OR4 (N11885, N11868, N861, N2943, N1836);
or OR3 (N11886, N11882, N376, N6490);
buf BUF1 (N11887, N11878);
buf BUF1 (N11888, N11876);
xor XOR2 (N11889, N11883, N10647);
xor XOR2 (N11890, N11880, N10075);
and AND3 (N11891, N11889, N10694, N9750);
and AND4 (N11892, N11887, N7506, N5924, N1444);
xor XOR2 (N11893, N11890, N9518);
buf BUF1 (N11894, N11877);
not NOT1 (N11895, N11891);
buf BUF1 (N11896, N11863);
buf BUF1 (N11897, N11888);
not NOT1 (N11898, N11896);
nand NAND3 (N11899, N11895, N11430, N3015);
nor NOR2 (N11900, N11893, N392);
or OR3 (N11901, N11897, N8658, N5239);
nand NAND4 (N11902, N11885, N3921, N6703, N6609);
and AND2 (N11903, N11892, N3828);
buf BUF1 (N11904, N11894);
not NOT1 (N11905, N11903);
buf BUF1 (N11906, N11905);
nand NAND4 (N11907, N11906, N10385, N9064, N9682);
or OR4 (N11908, N11907, N9619, N4612, N3223);
not NOT1 (N11909, N11886);
not NOT1 (N11910, N11908);
buf BUF1 (N11911, N11909);
nand NAND3 (N11912, N11900, N9270, N8373);
xor XOR2 (N11913, N11901, N6316);
nand NAND2 (N11914, N11899, N9635);
nand NAND4 (N11915, N11911, N11571, N4706, N6218);
xor XOR2 (N11916, N11898, N8041);
and AND4 (N11917, N11915, N2301, N2656, N3405);
nor NOR4 (N11918, N11902, N4244, N9247, N8563);
nor NOR4 (N11919, N11910, N7179, N1037, N6181);
and AND3 (N11920, N11913, N2894, N4028);
xor XOR2 (N11921, N11917, N9996);
xor XOR2 (N11922, N11920, N2848);
buf BUF1 (N11923, N11904);
buf BUF1 (N11924, N11919);
buf BUF1 (N11925, N11922);
xor XOR2 (N11926, N11912, N10439);
not NOT1 (N11927, N11914);
xor XOR2 (N11928, N11924, N1818);
or OR2 (N11929, N11872, N293);
not NOT1 (N11930, N11918);
xor XOR2 (N11931, N11926, N11155);
nand NAND2 (N11932, N11884, N10096);
buf BUF1 (N11933, N11932);
xor XOR2 (N11934, N11925, N9770);
buf BUF1 (N11935, N11929);
xor XOR2 (N11936, N11934, N9373);
buf BUF1 (N11937, N11921);
xor XOR2 (N11938, N11933, N11271);
not NOT1 (N11939, N11931);
or OR2 (N11940, N11935, N9319);
nor NOR4 (N11941, N11936, N1674, N8234, N10750);
buf BUF1 (N11942, N11940);
not NOT1 (N11943, N11930);
buf BUF1 (N11944, N11916);
xor XOR2 (N11945, N11927, N2631);
xor XOR2 (N11946, N11928, N977);
and AND2 (N11947, N11944, N11607);
xor XOR2 (N11948, N11941, N10030);
xor XOR2 (N11949, N11945, N853);
xor XOR2 (N11950, N11949, N10049);
xor XOR2 (N11951, N11950, N2048);
not NOT1 (N11952, N11943);
and AND3 (N11953, N11923, N7452, N6336);
and AND4 (N11954, N11947, N8412, N6117, N6628);
xor XOR2 (N11955, N11953, N1940);
nand NAND4 (N11956, N11948, N1586, N5497, N5257);
nor NOR2 (N11957, N11955, N11893);
buf BUF1 (N11958, N11938);
nand NAND2 (N11959, N11951, N6009);
and AND4 (N11960, N11956, N1807, N6394, N4892);
buf BUF1 (N11961, N11957);
buf BUF1 (N11962, N11942);
xor XOR2 (N11963, N11946, N6742);
nor NOR3 (N11964, N11952, N4584, N11792);
xor XOR2 (N11965, N11959, N250);
and AND2 (N11966, N11963, N9791);
nor NOR4 (N11967, N11965, N5438, N5180, N1880);
or OR3 (N11968, N11937, N2430, N8390);
buf BUF1 (N11969, N11964);
buf BUF1 (N11970, N11960);
nor NOR3 (N11971, N11970, N11926, N11168);
buf BUF1 (N11972, N11968);
or OR2 (N11973, N11972, N11200);
xor XOR2 (N11974, N11961, N3492);
nand NAND3 (N11975, N11969, N10225, N9082);
buf BUF1 (N11976, N11974);
buf BUF1 (N11977, N11971);
nor NOR4 (N11978, N11973, N6386, N4594, N1990);
not NOT1 (N11979, N11976);
buf BUF1 (N11980, N11962);
or OR4 (N11981, N11958, N9903, N3121, N7190);
and AND2 (N11982, N11981, N864);
nor NOR3 (N11983, N11980, N2127, N5524);
xor XOR2 (N11984, N11978, N9772);
buf BUF1 (N11985, N11977);
not NOT1 (N11986, N11966);
buf BUF1 (N11987, N11967);
and AND2 (N11988, N11954, N622);
not NOT1 (N11989, N11983);
buf BUF1 (N11990, N11939);
or OR4 (N11991, N11987, N399, N10902, N11761);
nor NOR3 (N11992, N11989, N10873, N5999);
buf BUF1 (N11993, N11975);
or OR4 (N11994, N11993, N639, N11132, N6356);
or OR2 (N11995, N11985, N6016);
or OR2 (N11996, N11988, N8332);
xor XOR2 (N11997, N11991, N5732);
and AND4 (N11998, N11995, N10294, N9200, N5788);
not NOT1 (N11999, N11997);
or OR3 (N12000, N11998, N9016, N8072);
xor XOR2 (N12001, N11994, N4500);
nor NOR2 (N12002, N12001, N5079);
or OR3 (N12003, N11990, N10084, N543);
nor NOR4 (N12004, N11996, N658, N5171, N7862);
nand NAND3 (N12005, N11986, N6732, N433);
nand NAND4 (N12006, N11984, N5409, N699, N146);
xor XOR2 (N12007, N12006, N10694);
nand NAND2 (N12008, N12002, N3687);
nor NOR2 (N12009, N11999, N3171);
nor NOR3 (N12010, N12004, N4652, N5841);
not NOT1 (N12011, N12005);
and AND2 (N12012, N12007, N11193);
or OR3 (N12013, N12010, N10840, N1868);
nand NAND4 (N12014, N11979, N8926, N4132, N8293);
nor NOR3 (N12015, N12000, N3780, N3042);
xor XOR2 (N12016, N12012, N620);
xor XOR2 (N12017, N12009, N9116);
not NOT1 (N12018, N12003);
buf BUF1 (N12019, N12016);
buf BUF1 (N12020, N11992);
nand NAND3 (N12021, N11982, N9396, N5305);
nor NOR4 (N12022, N12017, N11211, N11273, N5631);
or OR4 (N12023, N12011, N1081, N919, N286);
and AND2 (N12024, N12013, N11621);
or OR2 (N12025, N12022, N667);
nand NAND3 (N12026, N12014, N9147, N10171);
or OR4 (N12027, N12023, N5628, N7542, N5151);
xor XOR2 (N12028, N12019, N1293);
and AND4 (N12029, N12025, N2330, N5019, N6813);
nor NOR2 (N12030, N12024, N276);
or OR2 (N12031, N12008, N4259);
or OR4 (N12032, N12026, N3603, N11393, N9039);
nor NOR2 (N12033, N12027, N1229);
nor NOR2 (N12034, N12028, N580);
xor XOR2 (N12035, N12030, N1109);
or OR4 (N12036, N12018, N8811, N9771, N3257);
not NOT1 (N12037, N12032);
nand NAND2 (N12038, N12033, N3412);
xor XOR2 (N12039, N12031, N4844);
and AND2 (N12040, N12020, N250);
not NOT1 (N12041, N12038);
buf BUF1 (N12042, N12029);
not NOT1 (N12043, N12035);
and AND2 (N12044, N12040, N6864);
nor NOR4 (N12045, N12041, N5818, N8155, N3950);
nand NAND2 (N12046, N12037, N9116);
nand NAND4 (N12047, N12015, N6632, N4145, N2419);
or OR4 (N12048, N12047, N4001, N1387, N5999);
nand NAND4 (N12049, N12036, N10069, N7228, N8563);
buf BUF1 (N12050, N12048);
and AND3 (N12051, N12050, N10687, N11703);
nor NOR2 (N12052, N12042, N355);
and AND3 (N12053, N12046, N9459, N2123);
nor NOR4 (N12054, N12044, N7487, N6409, N2770);
or OR4 (N12055, N12039, N7333, N6783, N6926);
and AND4 (N12056, N12051, N4351, N2278, N6156);
nor NOR3 (N12057, N12056, N9889, N6758);
buf BUF1 (N12058, N12057);
or OR4 (N12059, N12049, N11624, N7682, N4132);
or OR3 (N12060, N12053, N3704, N8606);
xor XOR2 (N12061, N12034, N653);
and AND3 (N12062, N12043, N1352, N9284);
and AND2 (N12063, N12061, N10022);
buf BUF1 (N12064, N12055);
xor XOR2 (N12065, N12052, N7662);
not NOT1 (N12066, N12021);
and AND3 (N12067, N12062, N6941, N8409);
not NOT1 (N12068, N12054);
not NOT1 (N12069, N12063);
or OR3 (N12070, N12060, N5801, N9190);
and AND2 (N12071, N12070, N1869);
not NOT1 (N12072, N12045);
nand NAND2 (N12073, N12065, N2845);
not NOT1 (N12074, N12071);
buf BUF1 (N12075, N12064);
or OR4 (N12076, N12059, N6042, N5041, N2787);
not NOT1 (N12077, N12069);
xor XOR2 (N12078, N12076, N3623);
and AND4 (N12079, N12077, N4036, N1051, N242);
not NOT1 (N12080, N12066);
and AND3 (N12081, N12074, N10973, N1898);
buf BUF1 (N12082, N12073);
or OR3 (N12083, N12075, N1606, N4949);
and AND4 (N12084, N12080, N8692, N1515, N1661);
and AND3 (N12085, N12068, N8885, N3125);
buf BUF1 (N12086, N12083);
not NOT1 (N12087, N12067);
not NOT1 (N12088, N12087);
not NOT1 (N12089, N12081);
xor XOR2 (N12090, N12082, N10667);
or OR3 (N12091, N12084, N3586, N1673);
or OR3 (N12092, N12089, N11377, N9063);
and AND2 (N12093, N12072, N7668);
not NOT1 (N12094, N12088);
nand NAND2 (N12095, N12090, N11324);
nor NOR4 (N12096, N12093, N84, N8997, N11908);
not NOT1 (N12097, N12078);
not NOT1 (N12098, N12097);
xor XOR2 (N12099, N12091, N6026);
buf BUF1 (N12100, N12079);
xor XOR2 (N12101, N12085, N10652);
and AND3 (N12102, N12101, N3600, N118);
nand NAND2 (N12103, N12095, N8495);
and AND4 (N12104, N12102, N7056, N8243, N2226);
xor XOR2 (N12105, N12086, N4706);
or OR3 (N12106, N12105, N9626, N4353);
nand NAND2 (N12107, N12094, N3110);
or OR2 (N12108, N12103, N7516);
and AND4 (N12109, N12108, N1742, N8913, N9540);
xor XOR2 (N12110, N12100, N855);
nand NAND4 (N12111, N12058, N11504, N6259, N9143);
buf BUF1 (N12112, N12096);
nand NAND4 (N12113, N12109, N4252, N3597, N12000);
nand NAND3 (N12114, N12099, N10762, N9378);
nor NOR2 (N12115, N12104, N11267);
xor XOR2 (N12116, N12115, N1147);
buf BUF1 (N12117, N12114);
or OR4 (N12118, N12111, N11306, N10313, N514);
not NOT1 (N12119, N12113);
not NOT1 (N12120, N12117);
not NOT1 (N12121, N12092);
nor NOR4 (N12122, N12116, N8764, N11282, N2079);
and AND4 (N12123, N12118, N9571, N11113, N4668);
nand NAND2 (N12124, N12121, N6210);
not NOT1 (N12125, N12124);
buf BUF1 (N12126, N12122);
not NOT1 (N12127, N12110);
or OR3 (N12128, N12107, N7147, N1975);
or OR2 (N12129, N12098, N4825);
not NOT1 (N12130, N12123);
and AND4 (N12131, N12120, N3490, N8665, N4173);
nor NOR3 (N12132, N12125, N2032, N4237);
or OR3 (N12133, N12127, N9668, N7545);
and AND2 (N12134, N12130, N2172);
nor NOR3 (N12135, N12112, N11214, N4695);
xor XOR2 (N12136, N12134, N6348);
nand NAND3 (N12137, N12131, N606, N442);
buf BUF1 (N12138, N12133);
not NOT1 (N12139, N12137);
nand NAND2 (N12140, N12136, N6101);
and AND3 (N12141, N12126, N4483, N4170);
not NOT1 (N12142, N12132);
and AND4 (N12143, N12141, N517, N3031, N276);
not NOT1 (N12144, N12139);
and AND2 (N12145, N12135, N12062);
not NOT1 (N12146, N12138);
nor NOR3 (N12147, N12129, N2496, N10114);
not NOT1 (N12148, N12119);
nand NAND3 (N12149, N12142, N11160, N4257);
not NOT1 (N12150, N12147);
buf BUF1 (N12151, N12149);
buf BUF1 (N12152, N12128);
buf BUF1 (N12153, N12145);
buf BUF1 (N12154, N12150);
xor XOR2 (N12155, N12151, N6031);
or OR2 (N12156, N12148, N10255);
buf BUF1 (N12157, N12144);
nand NAND4 (N12158, N12152, N5012, N56, N7726);
nand NAND4 (N12159, N12143, N1693, N3622, N8740);
or OR4 (N12160, N12154, N2941, N4168, N1850);
nor NOR3 (N12161, N12140, N10510, N4740);
and AND3 (N12162, N12146, N7705, N3406);
and AND3 (N12163, N12161, N8932, N1017);
buf BUF1 (N12164, N12153);
buf BUF1 (N12165, N12160);
buf BUF1 (N12166, N12165);
nor NOR3 (N12167, N12156, N5733, N7844);
nand NAND4 (N12168, N12163, N6192, N3557, N2705);
xor XOR2 (N12169, N12158, N9366);
nor NOR2 (N12170, N12166, N4976);
xor XOR2 (N12171, N12167, N1003);
xor XOR2 (N12172, N12170, N7980);
not NOT1 (N12173, N12162);
nor NOR4 (N12174, N12157, N8112, N7251, N11545);
buf BUF1 (N12175, N12159);
not NOT1 (N12176, N12155);
and AND3 (N12177, N12164, N2723, N5776);
and AND3 (N12178, N12106, N2832, N7210);
xor XOR2 (N12179, N12168, N5097);
nor NOR4 (N12180, N12174, N9956, N11180, N9382);
nand NAND4 (N12181, N12175, N2497, N5208, N8054);
not NOT1 (N12182, N12171);
nand NAND3 (N12183, N12181, N6125, N1405);
nor NOR2 (N12184, N12178, N11875);
or OR3 (N12185, N12182, N7683, N12159);
nand NAND4 (N12186, N12169, N1410, N9831, N4329);
and AND4 (N12187, N12180, N5973, N8950, N2258);
nand NAND3 (N12188, N12177, N10174, N10653);
not NOT1 (N12189, N12185);
nor NOR3 (N12190, N12184, N2273, N4810);
nor NOR2 (N12191, N12183, N11703);
nor NOR2 (N12192, N12187, N10847);
nor NOR4 (N12193, N12190, N7911, N9720, N7630);
nand NAND3 (N12194, N12179, N7564, N5050);
not NOT1 (N12195, N12172);
buf BUF1 (N12196, N12195);
nand NAND2 (N12197, N12193, N2174);
not NOT1 (N12198, N12194);
buf BUF1 (N12199, N12197);
buf BUF1 (N12200, N12198);
buf BUF1 (N12201, N12188);
xor XOR2 (N12202, N12189, N4704);
not NOT1 (N12203, N12176);
and AND3 (N12204, N12186, N7854, N11749);
nor NOR2 (N12205, N12191, N1485);
or OR2 (N12206, N12201, N2265);
buf BUF1 (N12207, N12173);
or OR4 (N12208, N12205, N11473, N11569, N2912);
not NOT1 (N12209, N12204);
and AND3 (N12210, N12203, N1848, N2696);
buf BUF1 (N12211, N12206);
buf BUF1 (N12212, N12199);
or OR3 (N12213, N12192, N9062, N7824);
nor NOR2 (N12214, N12211, N4759);
xor XOR2 (N12215, N12213, N8284);
or OR3 (N12216, N12209, N9295, N9569);
and AND3 (N12217, N12196, N1925, N538);
nand NAND2 (N12218, N12214, N10384);
nand NAND2 (N12219, N12208, N2790);
and AND2 (N12220, N12215, N10167);
nor NOR4 (N12221, N12219, N10989, N2891, N9155);
or OR4 (N12222, N12207, N696, N7519, N7470);
nand NAND4 (N12223, N12221, N6646, N6132, N8756);
not NOT1 (N12224, N12200);
xor XOR2 (N12225, N12212, N11516);
not NOT1 (N12226, N12225);
nand NAND3 (N12227, N12220, N6489, N1044);
or OR4 (N12228, N12202, N7624, N4367, N6928);
nand NAND2 (N12229, N12226, N749);
xor XOR2 (N12230, N12228, N9492);
xor XOR2 (N12231, N12229, N6965);
or OR2 (N12232, N12223, N12151);
or OR3 (N12233, N12227, N7240, N4005);
nand NAND4 (N12234, N12217, N5907, N4454, N8750);
buf BUF1 (N12235, N12218);
nand NAND2 (N12236, N12233, N6588);
and AND2 (N12237, N12210, N3007);
nor NOR4 (N12238, N12237, N7882, N367, N10087);
or OR2 (N12239, N12235, N538);
not NOT1 (N12240, N12232);
buf BUF1 (N12241, N12234);
xor XOR2 (N12242, N12236, N4276);
not NOT1 (N12243, N12240);
nor NOR2 (N12244, N12241, N682);
not NOT1 (N12245, N12224);
not NOT1 (N12246, N12231);
xor XOR2 (N12247, N12222, N6765);
nor NOR4 (N12248, N12244, N7346, N517, N11961);
xor XOR2 (N12249, N12243, N1125);
nand NAND3 (N12250, N12245, N10978, N2575);
xor XOR2 (N12251, N12246, N6004);
nand NAND2 (N12252, N12216, N5454);
nor NOR3 (N12253, N12247, N8927, N295);
buf BUF1 (N12254, N12250);
not NOT1 (N12255, N12238);
nor NOR3 (N12256, N12253, N9007, N131);
or OR4 (N12257, N12254, N3129, N11189, N9837);
or OR2 (N12258, N12239, N381);
or OR4 (N12259, N12255, N1782, N7229, N11582);
nand NAND3 (N12260, N12256, N3015, N7169);
or OR3 (N12261, N12248, N233, N6369);
buf BUF1 (N12262, N12260);
not NOT1 (N12263, N12252);
xor XOR2 (N12264, N12242, N1970);
and AND4 (N12265, N12263, N9442, N12014, N7459);
buf BUF1 (N12266, N12264);
nand NAND4 (N12267, N12261, N4636, N12117, N180);
xor XOR2 (N12268, N12267, N8309);
xor XOR2 (N12269, N12230, N4991);
and AND4 (N12270, N12262, N610, N7784, N9049);
not NOT1 (N12271, N12265);
xor XOR2 (N12272, N12269, N4951);
and AND4 (N12273, N12266, N6808, N8716, N6199);
nor NOR4 (N12274, N12251, N4414, N12046, N7935);
xor XOR2 (N12275, N12271, N3724);
not NOT1 (N12276, N12272);
and AND2 (N12277, N12270, N36);
or OR4 (N12278, N12277, N7846, N2826, N1203);
nor NOR4 (N12279, N12274, N10464, N9927, N11693);
nor NOR4 (N12280, N12259, N9279, N11407, N6567);
or OR2 (N12281, N12268, N11274);
nor NOR4 (N12282, N12278, N7138, N5975, N7712);
and AND2 (N12283, N12276, N4566);
and AND4 (N12284, N12273, N7917, N4628, N2554);
xor XOR2 (N12285, N12284, N7015);
buf BUF1 (N12286, N12275);
nand NAND3 (N12287, N12281, N1907, N8080);
buf BUF1 (N12288, N12286);
nor NOR4 (N12289, N12279, N4442, N9937, N7133);
and AND3 (N12290, N12282, N2250, N5388);
and AND2 (N12291, N12249, N690);
or OR2 (N12292, N12257, N1766);
xor XOR2 (N12293, N12280, N1273);
and AND2 (N12294, N12290, N11713);
xor XOR2 (N12295, N12287, N6502);
or OR3 (N12296, N12292, N7864, N7579);
not NOT1 (N12297, N12288);
not NOT1 (N12298, N12295);
buf BUF1 (N12299, N12291);
xor XOR2 (N12300, N12283, N895);
not NOT1 (N12301, N12299);
buf BUF1 (N12302, N12294);
buf BUF1 (N12303, N12285);
not NOT1 (N12304, N12293);
not NOT1 (N12305, N12301);
xor XOR2 (N12306, N12303, N1995);
nor NOR2 (N12307, N12306, N9017);
nor NOR2 (N12308, N12305, N679);
nor NOR4 (N12309, N12289, N2578, N2474, N4876);
buf BUF1 (N12310, N12307);
nor NOR2 (N12311, N12302, N11527);
not NOT1 (N12312, N12300);
xor XOR2 (N12313, N12308, N3872);
buf BUF1 (N12314, N12297);
nor NOR3 (N12315, N12304, N2516, N8976);
buf BUF1 (N12316, N12314);
buf BUF1 (N12317, N12313);
nor NOR2 (N12318, N12315, N1731);
buf BUF1 (N12319, N12318);
buf BUF1 (N12320, N12319);
xor XOR2 (N12321, N12312, N528);
nand NAND2 (N12322, N12298, N11296);
xor XOR2 (N12323, N12258, N7726);
or OR4 (N12324, N12316, N10545, N6278, N8819);
xor XOR2 (N12325, N12317, N172);
nor NOR4 (N12326, N12310, N8430, N7916, N11140);
buf BUF1 (N12327, N12309);
xor XOR2 (N12328, N12320, N5534);
not NOT1 (N12329, N12325);
and AND2 (N12330, N12324, N5103);
not NOT1 (N12331, N12311);
buf BUF1 (N12332, N12330);
not NOT1 (N12333, N12328);
nand NAND3 (N12334, N12326, N10110, N7526);
not NOT1 (N12335, N12331);
and AND2 (N12336, N12323, N11677);
buf BUF1 (N12337, N12327);
or OR2 (N12338, N12322, N248);
or OR3 (N12339, N12296, N11658, N4389);
nand NAND2 (N12340, N12332, N5804);
buf BUF1 (N12341, N12336);
nor NOR3 (N12342, N12339, N3508, N431);
xor XOR2 (N12343, N12342, N11591);
nor NOR4 (N12344, N12340, N3001, N250, N10560);
nand NAND4 (N12345, N12335, N6599, N1047, N2374);
xor XOR2 (N12346, N12343, N1544);
nand NAND2 (N12347, N12345, N2940);
nand NAND2 (N12348, N12347, N8938);
nand NAND4 (N12349, N12329, N9412, N11435, N1986);
or OR3 (N12350, N12346, N5211, N3348);
and AND2 (N12351, N12333, N5556);
xor XOR2 (N12352, N12337, N5244);
nand NAND4 (N12353, N12349, N2057, N1136, N5327);
xor XOR2 (N12354, N12338, N9756);
not NOT1 (N12355, N12344);
xor XOR2 (N12356, N12354, N3810);
buf BUF1 (N12357, N12356);
nor NOR3 (N12358, N12341, N1744, N10003);
not NOT1 (N12359, N12348);
xor XOR2 (N12360, N12351, N9358);
nor NOR4 (N12361, N12350, N4031, N9511, N7715);
or OR2 (N12362, N12360, N1670);
buf BUF1 (N12363, N12321);
buf BUF1 (N12364, N12362);
buf BUF1 (N12365, N12352);
buf BUF1 (N12366, N12359);
xor XOR2 (N12367, N12353, N12088);
not NOT1 (N12368, N12363);
nor NOR2 (N12369, N12368, N6988);
and AND3 (N12370, N12365, N3887, N2410);
nor NOR4 (N12371, N12364, N10903, N11945, N9562);
or OR4 (N12372, N12369, N8557, N12169, N8174);
and AND3 (N12373, N12334, N11066, N4214);
nor NOR3 (N12374, N12361, N4266, N1904);
and AND4 (N12375, N12366, N539, N828, N11420);
nand NAND2 (N12376, N12357, N2457);
buf BUF1 (N12377, N12374);
xor XOR2 (N12378, N12373, N9613);
not NOT1 (N12379, N12375);
xor XOR2 (N12380, N12377, N1714);
buf BUF1 (N12381, N12378);
buf BUF1 (N12382, N12355);
or OR2 (N12383, N12371, N10860);
not NOT1 (N12384, N12367);
and AND3 (N12385, N12384, N1131, N7926);
and AND4 (N12386, N12382, N3339, N12110, N965);
and AND2 (N12387, N12372, N1200);
xor XOR2 (N12388, N12386, N6965);
nor NOR4 (N12389, N12370, N11010, N7597, N7573);
xor XOR2 (N12390, N12383, N3087);
or OR3 (N12391, N12376, N3490, N6340);
nand NAND4 (N12392, N12388, N3671, N9621, N12101);
and AND3 (N12393, N12381, N5475, N4959);
nor NOR3 (N12394, N12390, N7998, N10602);
nor NOR2 (N12395, N12391, N3676);
and AND3 (N12396, N12379, N4887, N4825);
nor NOR4 (N12397, N12387, N2098, N8317, N9728);
nor NOR4 (N12398, N12380, N10729, N3584, N9994);
buf BUF1 (N12399, N12398);
and AND2 (N12400, N12395, N2939);
not NOT1 (N12401, N12394);
nor NOR2 (N12402, N12397, N5693);
xor XOR2 (N12403, N12358, N8156);
or OR4 (N12404, N12393, N295, N2873, N11950);
and AND2 (N12405, N12399, N6473);
not NOT1 (N12406, N12404);
not NOT1 (N12407, N12385);
nand NAND3 (N12408, N12389, N5647, N10571);
nand NAND3 (N12409, N12408, N7523, N8015);
or OR3 (N12410, N12409, N2065, N3788);
nor NOR4 (N12411, N12410, N1380, N8600, N6476);
nand NAND3 (N12412, N12400, N5675, N4224);
xor XOR2 (N12413, N12406, N10215);
and AND4 (N12414, N12402, N8182, N8105, N2562);
buf BUF1 (N12415, N12401);
and AND2 (N12416, N12396, N6690);
not NOT1 (N12417, N12392);
or OR4 (N12418, N12414, N4471, N3958, N11505);
nor NOR3 (N12419, N12405, N5593, N6172);
not NOT1 (N12420, N12413);
xor XOR2 (N12421, N12412, N2210);
or OR2 (N12422, N12411, N5478);
nor NOR3 (N12423, N12415, N272, N4196);
nor NOR4 (N12424, N12416, N10312, N4975, N5160);
or OR3 (N12425, N12422, N3161, N3358);
nor NOR4 (N12426, N12418, N10160, N11488, N6701);
or OR4 (N12427, N12421, N1848, N1638, N8033);
or OR3 (N12428, N12427, N11384, N2436);
or OR4 (N12429, N12428, N10572, N8812, N4704);
nand NAND4 (N12430, N12426, N6818, N8236, N2597);
or OR4 (N12431, N12429, N8935, N2933, N1263);
nand NAND3 (N12432, N12419, N11062, N8919);
xor XOR2 (N12433, N12430, N1615);
nand NAND3 (N12434, N12423, N12348, N7012);
or OR2 (N12435, N12403, N3391);
or OR2 (N12436, N12425, N4609);
xor XOR2 (N12437, N12431, N3492);
not NOT1 (N12438, N12433);
buf BUF1 (N12439, N12434);
and AND4 (N12440, N12420, N4339, N11346, N9436);
or OR4 (N12441, N12438, N6935, N6212, N8532);
or OR2 (N12442, N12432, N11357);
not NOT1 (N12443, N12439);
and AND2 (N12444, N12442, N11622);
nor NOR2 (N12445, N12443, N4863);
not NOT1 (N12446, N12417);
buf BUF1 (N12447, N12445);
not NOT1 (N12448, N12447);
nor NOR2 (N12449, N12444, N3618);
and AND3 (N12450, N12446, N6673, N3610);
nand NAND2 (N12451, N12449, N8119);
nor NOR3 (N12452, N12448, N10554, N9269);
buf BUF1 (N12453, N12407);
nand NAND2 (N12454, N12424, N6868);
and AND3 (N12455, N12440, N10819, N10284);
not NOT1 (N12456, N12454);
and AND3 (N12457, N12436, N7494, N4447);
nor NOR4 (N12458, N12455, N1338, N9909, N4019);
nand NAND3 (N12459, N12437, N838, N2531);
nand NAND3 (N12460, N12456, N11716, N10613);
nor NOR2 (N12461, N12441, N7045);
or OR4 (N12462, N12458, N9158, N10431, N7284);
nor NOR2 (N12463, N12462, N8621);
nor NOR4 (N12464, N12457, N10797, N10807, N7754);
and AND4 (N12465, N12460, N4831, N8758, N3549);
not NOT1 (N12466, N12463);
and AND3 (N12467, N12451, N9581, N3729);
xor XOR2 (N12468, N12435, N2403);
buf BUF1 (N12469, N12466);
buf BUF1 (N12470, N12459);
xor XOR2 (N12471, N12450, N11352);
or OR2 (N12472, N12453, N5825);
not NOT1 (N12473, N12470);
not NOT1 (N12474, N12461);
nand NAND4 (N12475, N12473, N7533, N5302, N10456);
buf BUF1 (N12476, N12469);
or OR4 (N12477, N12467, N9384, N7750, N9085);
and AND4 (N12478, N12472, N9251, N390, N9777);
buf BUF1 (N12479, N12452);
buf BUF1 (N12480, N12476);
xor XOR2 (N12481, N12479, N8803);
buf BUF1 (N12482, N12464);
buf BUF1 (N12483, N12481);
or OR2 (N12484, N12477, N6017);
not NOT1 (N12485, N12468);
xor XOR2 (N12486, N12480, N11600);
not NOT1 (N12487, N12465);
or OR4 (N12488, N12483, N6766, N2558, N5926);
nand NAND4 (N12489, N12487, N2926, N2527, N10982);
nand NAND3 (N12490, N12474, N683, N447);
and AND3 (N12491, N12488, N2295, N5445);
xor XOR2 (N12492, N12471, N12126);
not NOT1 (N12493, N12478);
nor NOR2 (N12494, N12475, N9827);
nand NAND3 (N12495, N12484, N3475, N4683);
nand NAND3 (N12496, N12486, N11479, N8132);
or OR4 (N12497, N12490, N9822, N4971, N12002);
buf BUF1 (N12498, N12493);
nor NOR3 (N12499, N12492, N3518, N1929);
or OR2 (N12500, N12495, N6888);
buf BUF1 (N12501, N12491);
not NOT1 (N12502, N12482);
and AND2 (N12503, N12485, N10676);
buf BUF1 (N12504, N12498);
nor NOR3 (N12505, N12500, N12457, N3075);
nand NAND3 (N12506, N12505, N3306, N12496);
or OR2 (N12507, N2797, N3243);
not NOT1 (N12508, N12507);
nand NAND4 (N12509, N12503, N6896, N11302, N301);
nand NAND4 (N12510, N12494, N2180, N2823, N9821);
buf BUF1 (N12511, N12509);
or OR3 (N12512, N12501, N952, N3759);
nor NOR2 (N12513, N12506, N2653);
buf BUF1 (N12514, N12499);
not NOT1 (N12515, N12502);
or OR2 (N12516, N12489, N8738);
nand NAND3 (N12517, N12514, N3163, N1809);
nand NAND3 (N12518, N12515, N7275, N9264);
nor NOR3 (N12519, N12511, N4215, N7952);
nand NAND2 (N12520, N12516, N5126);
or OR4 (N12521, N12513, N842, N7392, N11681);
nand NAND4 (N12522, N12519, N11750, N3880, N10036);
nor NOR3 (N12523, N12510, N5812, N9823);
not NOT1 (N12524, N12518);
or OR3 (N12525, N12508, N4647, N10661);
and AND2 (N12526, N12525, N11329);
or OR4 (N12527, N12512, N10745, N4177, N12115);
nand NAND3 (N12528, N12523, N3069, N1693);
nor NOR2 (N12529, N12524, N49);
or OR4 (N12530, N12504, N10167, N1852, N5844);
not NOT1 (N12531, N12517);
or OR2 (N12532, N12497, N6919);
buf BUF1 (N12533, N12532);
nor NOR2 (N12534, N12521, N10781);
nor NOR3 (N12535, N12529, N4401, N11611);
and AND3 (N12536, N12527, N11132, N6740);
or OR3 (N12537, N12530, N10614, N8358);
or OR3 (N12538, N12533, N7735, N1448);
and AND4 (N12539, N12526, N5158, N10127, N1341);
nand NAND4 (N12540, N12534, N12080, N10871, N4955);
xor XOR2 (N12541, N12540, N12346);
xor XOR2 (N12542, N12536, N10139);
and AND3 (N12543, N12531, N6954, N12027);
xor XOR2 (N12544, N12543, N8003);
not NOT1 (N12545, N12539);
nor NOR3 (N12546, N12537, N7478, N7832);
buf BUF1 (N12547, N12541);
or OR4 (N12548, N12528, N4826, N6834, N182);
not NOT1 (N12549, N12544);
and AND3 (N12550, N12538, N9788, N10169);
not NOT1 (N12551, N12545);
nand NAND3 (N12552, N12520, N6285, N7795);
and AND2 (N12553, N12522, N5526);
buf BUF1 (N12554, N12549);
buf BUF1 (N12555, N12551);
not NOT1 (N12556, N12550);
nand NAND4 (N12557, N12548, N6499, N6655, N7379);
or OR2 (N12558, N12552, N11571);
nand NAND3 (N12559, N12553, N8350, N8067);
not NOT1 (N12560, N12558);
or OR2 (N12561, N12547, N1650);
not NOT1 (N12562, N12561);
xor XOR2 (N12563, N12535, N7716);
nor NOR4 (N12564, N12560, N6144, N11836, N7205);
nand NAND2 (N12565, N12559, N6152);
nand NAND2 (N12566, N12562, N1377);
xor XOR2 (N12567, N12554, N12555);
and AND4 (N12568, N2108, N2635, N5498, N4383);
xor XOR2 (N12569, N12563, N9004);
buf BUF1 (N12570, N12557);
buf BUF1 (N12571, N12556);
buf BUF1 (N12572, N12565);
or OR2 (N12573, N12564, N11475);
not NOT1 (N12574, N12573);
and AND3 (N12575, N12572, N3100, N3332);
buf BUF1 (N12576, N12542);
xor XOR2 (N12577, N12569, N4066);
or OR4 (N12578, N12567, N8512, N748, N5802);
xor XOR2 (N12579, N12566, N12534);
xor XOR2 (N12580, N12546, N1760);
and AND3 (N12581, N12571, N1781, N1326);
xor XOR2 (N12582, N12580, N481);
not NOT1 (N12583, N12576);
nand NAND2 (N12584, N12579, N1712);
nor NOR2 (N12585, N12578, N1976);
buf BUF1 (N12586, N12585);
nor NOR4 (N12587, N12583, N8917, N6244, N7549);
xor XOR2 (N12588, N12587, N9081);
and AND2 (N12589, N12570, N8064);
and AND4 (N12590, N12584, N8610, N2453, N4711);
nand NAND2 (N12591, N12589, N3596);
nand NAND4 (N12592, N12574, N3695, N9412, N8119);
nor NOR3 (N12593, N12581, N6746, N10542);
nor NOR4 (N12594, N12592, N4014, N10329, N11399);
buf BUF1 (N12595, N12586);
xor XOR2 (N12596, N12595, N10034);
nand NAND3 (N12597, N12591, N8917, N4256);
buf BUF1 (N12598, N12594);
or OR2 (N12599, N12575, N5802);
buf BUF1 (N12600, N12599);
nand NAND3 (N12601, N12577, N8342, N4102);
nand NAND3 (N12602, N12593, N7676, N647);
not NOT1 (N12603, N12582);
and AND3 (N12604, N12596, N18, N6518);
nand NAND4 (N12605, N12601, N4709, N5751, N11114);
and AND2 (N12606, N12604, N11386);
not NOT1 (N12607, N12603);
xor XOR2 (N12608, N12607, N9268);
or OR3 (N12609, N12600, N9640, N4665);
xor XOR2 (N12610, N12568, N12361);
and AND2 (N12611, N12610, N11455);
xor XOR2 (N12612, N12605, N9412);
xor XOR2 (N12613, N12597, N8253);
or OR2 (N12614, N12588, N2717);
buf BUF1 (N12615, N12598);
xor XOR2 (N12616, N12602, N7423);
nand NAND2 (N12617, N12611, N8173);
nand NAND4 (N12618, N12608, N6345, N8195, N12175);
or OR3 (N12619, N12615, N9391, N6499);
xor XOR2 (N12620, N12606, N2789);
or OR4 (N12621, N12619, N2211, N9077, N10539);
xor XOR2 (N12622, N12609, N1914);
not NOT1 (N12623, N12617);
buf BUF1 (N12624, N12622);
or OR3 (N12625, N12616, N2026, N10546);
nor NOR4 (N12626, N12621, N3864, N5437, N1435);
or OR2 (N12627, N12624, N8031);
or OR2 (N12628, N12614, N481);
or OR2 (N12629, N12613, N2789);
not NOT1 (N12630, N12612);
not NOT1 (N12631, N12625);
buf BUF1 (N12632, N12590);
and AND4 (N12633, N12627, N6624, N9419, N6752);
nand NAND2 (N12634, N12628, N6347);
nor NOR3 (N12635, N12631, N10863, N6046);
and AND4 (N12636, N12626, N7913, N6083, N8354);
not NOT1 (N12637, N12634);
or OR3 (N12638, N12636, N11986, N12456);
or OR2 (N12639, N12629, N11015);
nor NOR2 (N12640, N12618, N8467);
or OR2 (N12641, N12637, N5664);
not NOT1 (N12642, N12632);
buf BUF1 (N12643, N12641);
and AND3 (N12644, N12639, N6920, N8688);
xor XOR2 (N12645, N12633, N8753);
nand NAND2 (N12646, N12645, N11863);
buf BUF1 (N12647, N12623);
and AND2 (N12648, N12642, N11647);
nor NOR4 (N12649, N12630, N6503, N47, N11861);
buf BUF1 (N12650, N12646);
and AND4 (N12651, N12644, N4919, N3467, N10482);
nand NAND4 (N12652, N12620, N7860, N4768, N1746);
nand NAND4 (N12653, N12643, N5780, N9913, N12085);
nor NOR3 (N12654, N12640, N2836, N6721);
xor XOR2 (N12655, N12654, N8152);
or OR2 (N12656, N12648, N7286);
and AND2 (N12657, N12652, N9270);
xor XOR2 (N12658, N12638, N998);
buf BUF1 (N12659, N12647);
nand NAND4 (N12660, N12635, N8339, N7106, N10159);
and AND4 (N12661, N12657, N4109, N8782, N12103);
xor XOR2 (N12662, N12655, N5476);
xor XOR2 (N12663, N12649, N12174);
and AND3 (N12664, N12651, N6916, N2411);
and AND3 (N12665, N12659, N12038, N6328);
not NOT1 (N12666, N12658);
buf BUF1 (N12667, N12665);
or OR2 (N12668, N12650, N11876);
nand NAND4 (N12669, N12656, N9272, N5569, N3874);
buf BUF1 (N12670, N12666);
not NOT1 (N12671, N12668);
and AND2 (N12672, N12653, N10656);
nor NOR2 (N12673, N12667, N8221);
nor NOR3 (N12674, N12662, N3345, N8585);
nor NOR4 (N12675, N12670, N4939, N7390, N3626);
not NOT1 (N12676, N12672);
and AND4 (N12677, N12674, N7730, N652, N5600);
nor NOR3 (N12678, N12676, N5127, N7008);
not NOT1 (N12679, N12664);
not NOT1 (N12680, N12673);
or OR2 (N12681, N12671, N11742);
buf BUF1 (N12682, N12679);
or OR2 (N12683, N12682, N9512);
xor XOR2 (N12684, N12661, N10494);
nand NAND3 (N12685, N12683, N11386, N8849);
buf BUF1 (N12686, N12678);
not NOT1 (N12687, N12677);
xor XOR2 (N12688, N12675, N6794);
nor NOR3 (N12689, N12686, N11181, N1476);
nor NOR2 (N12690, N12663, N11231);
xor XOR2 (N12691, N12689, N6368);
nand NAND3 (N12692, N12688, N6187, N2630);
not NOT1 (N12693, N12680);
nand NAND4 (N12694, N12685, N8200, N2205, N4749);
not NOT1 (N12695, N12681);
not NOT1 (N12696, N12691);
or OR3 (N12697, N12693, N206, N244);
not NOT1 (N12698, N12660);
nor NOR3 (N12699, N12697, N8335, N3210);
buf BUF1 (N12700, N12669);
nor NOR2 (N12701, N12700, N12448);
nor NOR3 (N12702, N12698, N4983, N1887);
nand NAND4 (N12703, N12696, N1196, N5115, N850);
nand NAND2 (N12704, N12703, N1342);
nor NOR4 (N12705, N12687, N1138, N10407, N8831);
buf BUF1 (N12706, N12702);
or OR2 (N12707, N12694, N6379);
nor NOR4 (N12708, N12695, N6842, N5155, N7670);
or OR4 (N12709, N12708, N5230, N7045, N6782);
nand NAND3 (N12710, N12699, N166, N4086);
nand NAND2 (N12711, N12684, N238);
and AND2 (N12712, N12710, N5421);
xor XOR2 (N12713, N12690, N3419);
xor XOR2 (N12714, N12701, N10252);
nand NAND3 (N12715, N12713, N12659, N9053);
and AND4 (N12716, N12706, N9392, N9040, N6101);
nand NAND3 (N12717, N12715, N10248, N1865);
and AND4 (N12718, N12705, N7764, N3865, N1392);
not NOT1 (N12719, N12711);
or OR2 (N12720, N12716, N11073);
buf BUF1 (N12721, N12712);
or OR2 (N12722, N12707, N6527);
xor XOR2 (N12723, N12714, N3072);
or OR4 (N12724, N12692, N10893, N12445, N2452);
and AND4 (N12725, N12720, N5886, N2299, N8424);
nor NOR3 (N12726, N12723, N8230, N7542);
and AND4 (N12727, N12726, N1758, N7047, N2790);
xor XOR2 (N12728, N12718, N7279);
buf BUF1 (N12729, N12704);
nand NAND4 (N12730, N12729, N5713, N7708, N11327);
buf BUF1 (N12731, N12709);
not NOT1 (N12732, N12721);
nor NOR3 (N12733, N12724, N10483, N9610);
nand NAND2 (N12734, N12732, N8190);
nor NOR2 (N12735, N12728, N11843);
nand NAND2 (N12736, N12725, N447);
buf BUF1 (N12737, N12730);
not NOT1 (N12738, N12737);
not NOT1 (N12739, N12719);
or OR2 (N12740, N12738, N10686);
nor NOR4 (N12741, N12736, N11854, N6935, N7604);
nand NAND2 (N12742, N12739, N7650);
buf BUF1 (N12743, N12727);
nand NAND2 (N12744, N12741, N1283);
and AND4 (N12745, N12733, N6131, N3612, N8692);
nor NOR4 (N12746, N12744, N7739, N3170, N10268);
buf BUF1 (N12747, N12717);
buf BUF1 (N12748, N12734);
or OR3 (N12749, N12748, N3402, N7193);
buf BUF1 (N12750, N12747);
nor NOR3 (N12751, N12745, N540, N10339);
nor NOR4 (N12752, N12722, N2257, N671, N8216);
xor XOR2 (N12753, N12731, N12230);
and AND3 (N12754, N12746, N4822, N6844);
nor NOR4 (N12755, N12749, N5217, N11533, N2153);
not NOT1 (N12756, N12740);
or OR3 (N12757, N12755, N1439, N10580);
buf BUF1 (N12758, N12751);
nor NOR3 (N12759, N12752, N11760, N6670);
nor NOR4 (N12760, N12758, N10732, N11026, N12013);
buf BUF1 (N12761, N12754);
nor NOR3 (N12762, N12760, N4061, N5120);
or OR2 (N12763, N12756, N987);
buf BUF1 (N12764, N12750);
and AND4 (N12765, N12762, N4450, N9139, N2938);
buf BUF1 (N12766, N12757);
nor NOR2 (N12767, N12759, N1342);
xor XOR2 (N12768, N12766, N477);
and AND3 (N12769, N12743, N2389, N7206);
and AND4 (N12770, N12765, N5456, N7320, N510);
nand NAND2 (N12771, N12742, N1767);
or OR2 (N12772, N12768, N11501);
nand NAND3 (N12773, N12735, N7639, N9791);
xor XOR2 (N12774, N12753, N7797);
buf BUF1 (N12775, N12767);
buf BUF1 (N12776, N12772);
xor XOR2 (N12777, N12776, N3522);
not NOT1 (N12778, N12770);
nor NOR4 (N12779, N12773, N346, N4968, N3166);
and AND2 (N12780, N12778, N5356);
or OR3 (N12781, N12763, N761, N9944);
nand NAND4 (N12782, N12779, N8279, N11551, N2388);
nor NOR2 (N12783, N12761, N11458);
and AND4 (N12784, N12781, N4790, N9603, N5479);
not NOT1 (N12785, N12783);
nand NAND2 (N12786, N12774, N8262);
buf BUF1 (N12787, N12771);
and AND4 (N12788, N12775, N11601, N9854, N8368);
buf BUF1 (N12789, N12777);
nor NOR2 (N12790, N12784, N6799);
buf BUF1 (N12791, N12788);
and AND3 (N12792, N12785, N9504, N12458);
or OR4 (N12793, N12782, N6415, N12625, N8205);
buf BUF1 (N12794, N12791);
xor XOR2 (N12795, N12780, N1927);
buf BUF1 (N12796, N12795);
xor XOR2 (N12797, N12790, N6814);
or OR2 (N12798, N12787, N10429);
and AND2 (N12799, N12797, N8350);
not NOT1 (N12800, N12786);
nand NAND4 (N12801, N12793, N7386, N12446, N9666);
xor XOR2 (N12802, N12800, N11474);
xor XOR2 (N12803, N12802, N8427);
nand NAND3 (N12804, N12789, N10822, N9047);
not NOT1 (N12805, N12798);
nor NOR3 (N12806, N12803, N7832, N8867);
and AND3 (N12807, N12806, N12129, N9344);
and AND3 (N12808, N12805, N4571, N3018);
xor XOR2 (N12809, N12804, N3628);
nor NOR2 (N12810, N12769, N5014);
and AND3 (N12811, N12796, N7951, N1988);
xor XOR2 (N12812, N12807, N10216);
buf BUF1 (N12813, N12799);
buf BUF1 (N12814, N12812);
xor XOR2 (N12815, N12764, N11165);
not NOT1 (N12816, N12815);
nor NOR3 (N12817, N12813, N1942, N1282);
not NOT1 (N12818, N12794);
nor NOR3 (N12819, N12817, N10542, N8033);
nand NAND3 (N12820, N12814, N9730, N565);
or OR3 (N12821, N12808, N12199, N8287);
nand NAND4 (N12822, N12819, N791, N3690, N4712);
endmodule