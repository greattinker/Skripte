// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20;

output N2517,N2516,N2519,N2514,N2515,N2518,N2498,N2513,N2506,N2520;

and AND2 (N21, N9, N9);
buf BUF1 (N22, N18);
or OR4 (N23, N3, N10, N8, N13);
nor NOR2 (N24, N6, N18);
not NOT1 (N25, N3);
nand NAND2 (N26, N19, N5);
or OR3 (N27, N19, N19, N9);
nand NAND4 (N28, N23, N17, N16, N4);
not NOT1 (N29, N3);
and AND3 (N30, N13, N13, N8);
nor NOR2 (N31, N24, N24);
xor XOR2 (N32, N6, N17);
not NOT1 (N33, N27);
nor NOR3 (N34, N22, N4, N8);
nor NOR4 (N35, N21, N7, N22, N12);
xor XOR2 (N36, N29, N35);
nor NOR2 (N37, N21, N17);
not NOT1 (N38, N28);
nor NOR4 (N39, N34, N28, N10, N22);
buf BUF1 (N40, N25);
buf BUF1 (N41, N37);
buf BUF1 (N42, N32);
nor NOR2 (N43, N36, N8);
xor XOR2 (N44, N30, N43);
nor NOR3 (N45, N4, N10, N5);
xor XOR2 (N46, N45, N36);
nand NAND2 (N47, N26, N16);
and AND3 (N48, N33, N31, N30);
and AND4 (N49, N11, N18, N21, N45);
not NOT1 (N50, N48);
buf BUF1 (N51, N41);
not NOT1 (N52, N50);
buf BUF1 (N53, N44);
or OR2 (N54, N53, N53);
and AND2 (N55, N47, N15);
nor NOR2 (N56, N42, N42);
buf BUF1 (N57, N51);
buf BUF1 (N58, N38);
nand NAND2 (N59, N55, N55);
not NOT1 (N60, N46);
xor XOR2 (N61, N52, N22);
buf BUF1 (N62, N57);
nand NAND3 (N63, N40, N30, N48);
xor XOR2 (N64, N58, N3);
not NOT1 (N65, N63);
and AND2 (N66, N59, N64);
not NOT1 (N67, N53);
buf BUF1 (N68, N56);
or OR2 (N69, N54, N15);
not NOT1 (N70, N60);
or OR3 (N71, N68, N17, N15);
or OR3 (N72, N39, N10, N18);
nor NOR3 (N73, N49, N12, N26);
xor XOR2 (N74, N65, N52);
not NOT1 (N75, N70);
nand NAND2 (N76, N67, N71);
xor XOR2 (N77, N74, N32);
and AND3 (N78, N42, N38, N6);
nand NAND4 (N79, N69, N45, N45, N17);
not NOT1 (N80, N62);
and AND2 (N81, N72, N65);
or OR2 (N82, N76, N28);
and AND2 (N83, N81, N10);
nor NOR3 (N84, N80, N52, N18);
or OR3 (N85, N79, N38, N37);
or OR4 (N86, N73, N30, N15, N68);
not NOT1 (N87, N82);
xor XOR2 (N88, N86, N1);
and AND3 (N89, N77, N70, N53);
xor XOR2 (N90, N84, N7);
or OR4 (N91, N88, N83, N67, N59);
xor XOR2 (N92, N76, N70);
or OR4 (N93, N61, N46, N81, N1);
and AND4 (N94, N85, N83, N29, N51);
nor NOR3 (N95, N75, N9, N35);
and AND2 (N96, N87, N4);
not NOT1 (N97, N92);
xor XOR2 (N98, N96, N69);
xor XOR2 (N99, N78, N68);
nor NOR2 (N100, N94, N89);
or OR2 (N101, N38, N5);
not NOT1 (N102, N93);
not NOT1 (N103, N101);
or OR3 (N104, N100, N103, N93);
not NOT1 (N105, N5);
nor NOR2 (N106, N98, N78);
and AND4 (N107, N102, N101, N74, N4);
nand NAND4 (N108, N106, N4, N86, N78);
not NOT1 (N109, N99);
and AND4 (N110, N95, N86, N40, N72);
buf BUF1 (N111, N105);
buf BUF1 (N112, N66);
nor NOR2 (N113, N97, N76);
and AND4 (N114, N107, N73, N13, N110);
not NOT1 (N115, N93);
buf BUF1 (N116, N104);
and AND3 (N117, N113, N92, N83);
nor NOR4 (N118, N90, N102, N58, N67);
not NOT1 (N119, N109);
buf BUF1 (N120, N108);
buf BUF1 (N121, N120);
buf BUF1 (N122, N111);
and AND2 (N123, N116, N107);
and AND3 (N124, N123, N17, N13);
nand NAND4 (N125, N112, N93, N27, N111);
not NOT1 (N126, N124);
nor NOR3 (N127, N91, N77, N86);
xor XOR2 (N128, N118, N64);
xor XOR2 (N129, N122, N48);
or OR3 (N130, N128, N69, N63);
buf BUF1 (N131, N127);
and AND3 (N132, N121, N95, N50);
buf BUF1 (N133, N130);
not NOT1 (N134, N129);
not NOT1 (N135, N132);
and AND2 (N136, N135, N125);
or OR3 (N137, N71, N109, N22);
or OR3 (N138, N115, N41, N74);
and AND2 (N139, N134, N129);
not NOT1 (N140, N133);
not NOT1 (N141, N131);
nor NOR2 (N142, N137, N13);
and AND4 (N143, N126, N129, N80, N136);
nand NAND2 (N144, N82, N10);
nor NOR2 (N145, N117, N12);
not NOT1 (N146, N119);
xor XOR2 (N147, N138, N56);
and AND4 (N148, N141, N14, N87, N50);
nor NOR2 (N149, N140, N114);
and AND2 (N150, N18, N97);
nand NAND2 (N151, N150, N146);
xor XOR2 (N152, N38, N74);
buf BUF1 (N153, N139);
not NOT1 (N154, N147);
and AND2 (N155, N142, N142);
or OR4 (N156, N149, N27, N79, N104);
xor XOR2 (N157, N152, N38);
or OR3 (N158, N157, N147, N53);
buf BUF1 (N159, N151);
or OR3 (N160, N158, N107, N123);
not NOT1 (N161, N143);
nand NAND3 (N162, N156, N25, N23);
nor NOR2 (N163, N160, N118);
not NOT1 (N164, N155);
not NOT1 (N165, N163);
nand NAND3 (N166, N154, N66, N145);
and AND4 (N167, N129, N134, N33, N48);
nor NOR2 (N168, N162, N33);
nand NAND4 (N169, N148, N5, N134, N100);
xor XOR2 (N170, N165, N74);
and AND3 (N171, N166, N41, N50);
nand NAND4 (N172, N161, N98, N143, N92);
buf BUF1 (N173, N167);
and AND4 (N174, N164, N129, N137, N33);
nor NOR4 (N175, N169, N91, N23, N161);
and AND4 (N176, N175, N70, N140, N106);
not NOT1 (N177, N159);
xor XOR2 (N178, N176, N52);
xor XOR2 (N179, N178, N72);
nor NOR4 (N180, N173, N40, N13, N47);
and AND3 (N181, N177, N29, N159);
buf BUF1 (N182, N171);
nor NOR4 (N183, N182, N44, N47, N85);
and AND2 (N184, N170, N105);
and AND2 (N185, N168, N70);
buf BUF1 (N186, N183);
nand NAND4 (N187, N144, N96, N120, N11);
nor NOR4 (N188, N179, N74, N23, N91);
or OR3 (N189, N186, N97, N66);
not NOT1 (N190, N172);
and AND2 (N191, N187, N108);
buf BUF1 (N192, N184);
and AND3 (N193, N181, N64, N174);
or OR4 (N194, N84, N55, N57, N189);
buf BUF1 (N195, N10);
xor XOR2 (N196, N153, N14);
xor XOR2 (N197, N185, N156);
or OR3 (N198, N188, N99, N72);
nand NAND3 (N199, N191, N15, N78);
buf BUF1 (N200, N199);
and AND2 (N201, N190, N143);
buf BUF1 (N202, N194);
nand NAND4 (N203, N195, N189, N122, N181);
xor XOR2 (N204, N192, N37);
and AND3 (N205, N198, N81, N34);
buf BUF1 (N206, N196);
nor NOR3 (N207, N180, N3, N153);
nand NAND3 (N208, N193, N174, N53);
buf BUF1 (N209, N200);
xor XOR2 (N210, N203, N183);
and AND4 (N211, N205, N189, N68, N16);
nor NOR2 (N212, N208, N53);
buf BUF1 (N213, N211);
and AND2 (N214, N213, N45);
buf BUF1 (N215, N202);
not NOT1 (N216, N212);
nand NAND4 (N217, N209, N173, N200, N86);
xor XOR2 (N218, N201, N30);
buf BUF1 (N219, N197);
nor NOR4 (N220, N219, N107, N61, N107);
or OR3 (N221, N217, N197, N186);
and AND3 (N222, N215, N30, N195);
and AND2 (N223, N222, N178);
buf BUF1 (N224, N206);
or OR4 (N225, N221, N115, N117, N171);
or OR4 (N226, N210, N156, N43, N165);
or OR2 (N227, N204, N127);
buf BUF1 (N228, N227);
not NOT1 (N229, N226);
nand NAND4 (N230, N225, N150, N7, N33);
not NOT1 (N231, N229);
not NOT1 (N232, N224);
nor NOR2 (N233, N231, N36);
buf BUF1 (N234, N214);
not NOT1 (N235, N230);
nand NAND2 (N236, N235, N92);
xor XOR2 (N237, N218, N191);
nor NOR3 (N238, N223, N186, N71);
buf BUF1 (N239, N233);
nor NOR2 (N240, N207, N207);
nand NAND3 (N241, N239, N187, N204);
nor NOR4 (N242, N236, N217, N33, N64);
nand NAND3 (N243, N238, N154, N208);
nand NAND2 (N244, N216, N189);
buf BUF1 (N245, N244);
and AND2 (N246, N240, N151);
or OR4 (N247, N243, N53, N49, N246);
buf BUF1 (N248, N194);
not NOT1 (N249, N248);
nor NOR2 (N250, N242, N59);
and AND2 (N251, N250, N192);
and AND4 (N252, N249, N58, N208, N168);
xor XOR2 (N253, N252, N88);
nand NAND4 (N254, N220, N38, N120, N218);
and AND4 (N255, N254, N217, N6, N54);
buf BUF1 (N256, N237);
and AND4 (N257, N241, N56, N179, N105);
or OR4 (N258, N232, N249, N189, N74);
xor XOR2 (N259, N234, N2);
nor NOR2 (N260, N251, N65);
not NOT1 (N261, N256);
nor NOR3 (N262, N245, N212, N246);
and AND3 (N263, N253, N11, N10);
nand NAND4 (N264, N257, N197, N51, N204);
or OR3 (N265, N260, N213, N149);
nand NAND3 (N266, N258, N80, N132);
or OR3 (N267, N261, N157, N35);
or OR2 (N268, N263, N235);
not NOT1 (N269, N266);
and AND3 (N270, N259, N9, N189);
and AND4 (N271, N265, N115, N135, N158);
buf BUF1 (N272, N268);
nand NAND3 (N273, N272, N123, N4);
and AND3 (N274, N262, N187, N5);
buf BUF1 (N275, N247);
not NOT1 (N276, N273);
nor NOR4 (N277, N275, N66, N29, N55);
not NOT1 (N278, N264);
nand NAND3 (N279, N271, N260, N153);
not NOT1 (N280, N278);
or OR3 (N281, N280, N252, N236);
nand NAND3 (N282, N267, N237, N40);
nor NOR3 (N283, N279, N6, N219);
xor XOR2 (N284, N270, N146);
or OR4 (N285, N274, N227, N68, N146);
and AND3 (N286, N281, N37, N3);
and AND2 (N287, N255, N228);
and AND4 (N288, N129, N90, N92, N148);
not NOT1 (N289, N283);
buf BUF1 (N290, N284);
nand NAND2 (N291, N290, N177);
nand NAND3 (N292, N277, N243, N56);
xor XOR2 (N293, N289, N262);
nand NAND4 (N294, N292, N180, N175, N284);
nor NOR2 (N295, N276, N32);
xor XOR2 (N296, N285, N164);
nor NOR4 (N297, N291, N109, N203, N44);
xor XOR2 (N298, N297, N120);
or OR2 (N299, N288, N266);
buf BUF1 (N300, N298);
not NOT1 (N301, N269);
xor XOR2 (N302, N295, N49);
buf BUF1 (N303, N301);
nand NAND4 (N304, N287, N19, N170, N240);
nand NAND4 (N305, N303, N199, N48, N27);
buf BUF1 (N306, N293);
nor NOR3 (N307, N300, N95, N9);
buf BUF1 (N308, N306);
and AND2 (N309, N299, N82);
and AND2 (N310, N302, N211);
and AND2 (N311, N310, N93);
nand NAND4 (N312, N305, N109, N104, N31);
buf BUF1 (N313, N304);
xor XOR2 (N314, N308, N5);
not NOT1 (N315, N313);
and AND4 (N316, N309, N85, N298, N208);
xor XOR2 (N317, N282, N274);
or OR4 (N318, N315, N87, N146, N16);
buf BUF1 (N319, N314);
buf BUF1 (N320, N316);
not NOT1 (N321, N307);
not NOT1 (N322, N321);
or OR3 (N323, N320, N132, N83);
buf BUF1 (N324, N318);
nand NAND3 (N325, N324, N216, N239);
xor XOR2 (N326, N296, N211);
nand NAND4 (N327, N317, N91, N53, N289);
or OR3 (N328, N325, N252, N217);
xor XOR2 (N329, N312, N229);
nand NAND4 (N330, N319, N55, N93, N255);
or OR2 (N331, N330, N3);
xor XOR2 (N332, N329, N227);
xor XOR2 (N333, N331, N105);
nand NAND3 (N334, N323, N221, N63);
and AND4 (N335, N311, N178, N223, N16);
or OR4 (N336, N328, N174, N299, N233);
nor NOR2 (N337, N327, N217);
not NOT1 (N338, N336);
buf BUF1 (N339, N334);
nor NOR4 (N340, N294, N181, N144, N190);
not NOT1 (N341, N337);
nand NAND4 (N342, N335, N200, N151, N314);
and AND2 (N343, N338, N149);
nor NOR3 (N344, N322, N95, N129);
or OR4 (N345, N286, N157, N282, N57);
nand NAND3 (N346, N345, N74, N23);
nor NOR2 (N347, N340, N24);
not NOT1 (N348, N332);
nor NOR2 (N349, N346, N348);
xor XOR2 (N350, N7, N319);
xor XOR2 (N351, N333, N178);
xor XOR2 (N352, N344, N121);
nor NOR3 (N353, N349, N281, N234);
not NOT1 (N354, N341);
or OR3 (N355, N350, N306, N71);
and AND2 (N356, N343, N352);
nand NAND4 (N357, N356, N6, N244, N212);
and AND4 (N358, N187, N124, N234, N73);
not NOT1 (N359, N351);
nor NOR4 (N360, N358, N80, N67, N162);
xor XOR2 (N361, N342, N165);
nand NAND4 (N362, N339, N241, N77, N63);
nor NOR3 (N363, N357, N209, N275);
xor XOR2 (N364, N363, N216);
and AND2 (N365, N360, N82);
or OR2 (N366, N353, N310);
and AND2 (N367, N362, N161);
not NOT1 (N368, N365);
not NOT1 (N369, N361);
nor NOR2 (N370, N347, N62);
nor NOR3 (N371, N370, N142, N213);
or OR2 (N372, N368, N133);
not NOT1 (N373, N359);
buf BUF1 (N374, N364);
xor XOR2 (N375, N372, N287);
nor NOR3 (N376, N373, N354, N139);
and AND4 (N377, N12, N316, N357, N96);
not NOT1 (N378, N375);
buf BUF1 (N379, N377);
buf BUF1 (N380, N367);
not NOT1 (N381, N326);
or OR3 (N382, N371, N177, N339);
nor NOR4 (N383, N380, N351, N352, N281);
buf BUF1 (N384, N369);
not NOT1 (N385, N355);
nand NAND3 (N386, N384, N276, N68);
xor XOR2 (N387, N366, N299);
nor NOR3 (N388, N386, N205, N79);
nand NAND4 (N389, N378, N375, N318, N18);
nor NOR3 (N390, N382, N221, N249);
buf BUF1 (N391, N383);
not NOT1 (N392, N374);
xor XOR2 (N393, N388, N262);
and AND4 (N394, N392, N196, N220, N117);
and AND3 (N395, N379, N245, N297);
xor XOR2 (N396, N391, N45);
nor NOR3 (N397, N381, N257, N12);
xor XOR2 (N398, N390, N321);
buf BUF1 (N399, N394);
not NOT1 (N400, N398);
and AND2 (N401, N400, N307);
and AND2 (N402, N376, N118);
nand NAND4 (N403, N389, N277, N75, N176);
xor XOR2 (N404, N395, N319);
buf BUF1 (N405, N396);
xor XOR2 (N406, N393, N58);
buf BUF1 (N407, N387);
nand NAND3 (N408, N403, N407, N391);
xor XOR2 (N409, N153, N289);
xor XOR2 (N410, N404, N55);
nor NOR4 (N411, N409, N147, N199, N249);
or OR2 (N412, N410, N348);
nor NOR2 (N413, N411, N281);
nand NAND3 (N414, N399, N266, N388);
nand NAND3 (N415, N405, N70, N153);
buf BUF1 (N416, N406);
not NOT1 (N417, N402);
not NOT1 (N418, N416);
nand NAND4 (N419, N385, N301, N70, N128);
nor NOR3 (N420, N401, N52, N392);
nand NAND3 (N421, N413, N298, N14);
buf BUF1 (N422, N408);
xor XOR2 (N423, N418, N76);
not NOT1 (N424, N415);
and AND2 (N425, N414, N102);
and AND2 (N426, N420, N69);
buf BUF1 (N427, N425);
buf BUF1 (N428, N419);
nor NOR4 (N429, N421, N24, N195, N131);
not NOT1 (N430, N428);
nor NOR2 (N431, N429, N103);
or OR4 (N432, N430, N207, N404, N387);
or OR3 (N433, N397, N372, N45);
buf BUF1 (N434, N424);
not NOT1 (N435, N426);
nand NAND4 (N436, N431, N40, N256, N149);
not NOT1 (N437, N417);
nand NAND2 (N438, N433, N152);
nor NOR2 (N439, N423, N225);
or OR3 (N440, N436, N333, N323);
buf BUF1 (N441, N437);
nor NOR2 (N442, N412, N93);
xor XOR2 (N443, N432, N34);
buf BUF1 (N444, N422);
not NOT1 (N445, N427);
not NOT1 (N446, N441);
buf BUF1 (N447, N439);
or OR4 (N448, N435, N108, N411, N193);
buf BUF1 (N449, N446);
not NOT1 (N450, N443);
nand NAND2 (N451, N438, N406);
nor NOR3 (N452, N449, N349, N173);
or OR4 (N453, N447, N184, N73, N353);
nor NOR2 (N454, N451, N132);
and AND2 (N455, N445, N96);
buf BUF1 (N456, N448);
or OR4 (N457, N442, N33, N423, N320);
nor NOR3 (N458, N450, N296, N337);
xor XOR2 (N459, N452, N98);
buf BUF1 (N460, N457);
not NOT1 (N461, N444);
buf BUF1 (N462, N434);
or OR2 (N463, N458, N342);
buf BUF1 (N464, N440);
xor XOR2 (N465, N459, N296);
not NOT1 (N466, N463);
and AND2 (N467, N465, N156);
or OR4 (N468, N467, N443, N430, N299);
xor XOR2 (N469, N468, N241);
and AND4 (N470, N454, N85, N35, N451);
or OR4 (N471, N466, N124, N359, N233);
buf BUF1 (N472, N460);
or OR4 (N473, N469, N31, N431, N225);
xor XOR2 (N474, N461, N306);
nand NAND4 (N475, N470, N426, N459, N286);
not NOT1 (N476, N462);
buf BUF1 (N477, N456);
nor NOR2 (N478, N464, N310);
nor NOR4 (N479, N455, N371, N211, N88);
xor XOR2 (N480, N476, N168);
xor XOR2 (N481, N475, N202);
nand NAND4 (N482, N473, N233, N423, N325);
buf BUF1 (N483, N481);
nand NAND3 (N484, N471, N275, N342);
buf BUF1 (N485, N483);
xor XOR2 (N486, N482, N320);
or OR3 (N487, N472, N330, N274);
nor NOR3 (N488, N487, N458, N478);
buf BUF1 (N489, N285);
xor XOR2 (N490, N479, N469);
xor XOR2 (N491, N489, N81);
xor XOR2 (N492, N480, N89);
not NOT1 (N493, N488);
nor NOR2 (N494, N492, N330);
buf BUF1 (N495, N491);
xor XOR2 (N496, N495, N210);
nor NOR2 (N497, N490, N404);
buf BUF1 (N498, N477);
nand NAND2 (N499, N453, N459);
xor XOR2 (N500, N494, N189);
buf BUF1 (N501, N485);
xor XOR2 (N502, N501, N12);
not NOT1 (N503, N499);
and AND3 (N504, N484, N212, N360);
not NOT1 (N505, N504);
xor XOR2 (N506, N500, N248);
buf BUF1 (N507, N502);
xor XOR2 (N508, N493, N28);
or OR4 (N509, N497, N471, N203, N27);
nor NOR2 (N510, N506, N245);
and AND3 (N511, N486, N240, N46);
not NOT1 (N512, N508);
or OR2 (N513, N512, N505);
xor XOR2 (N514, N472, N124);
nand NAND2 (N515, N507, N438);
nor NOR3 (N516, N510, N395, N79);
nor NOR3 (N517, N511, N338, N96);
or OR3 (N518, N513, N348, N418);
or OR2 (N519, N474, N105);
buf BUF1 (N520, N514);
nand NAND4 (N521, N517, N195, N337, N435);
xor XOR2 (N522, N503, N23);
not NOT1 (N523, N498);
buf BUF1 (N524, N515);
nand NAND3 (N525, N518, N349, N252);
xor XOR2 (N526, N496, N90);
and AND2 (N527, N525, N309);
nand NAND3 (N528, N527, N451, N126);
not NOT1 (N529, N522);
nand NAND2 (N530, N526, N436);
or OR2 (N531, N520, N161);
nor NOR4 (N532, N528, N382, N505, N80);
buf BUF1 (N533, N523);
buf BUF1 (N534, N532);
or OR2 (N535, N529, N78);
buf BUF1 (N536, N519);
or OR2 (N537, N509, N463);
not NOT1 (N538, N533);
nand NAND3 (N539, N516, N405, N523);
nor NOR2 (N540, N521, N8);
not NOT1 (N541, N531);
nor NOR3 (N542, N540, N316, N101);
buf BUF1 (N543, N541);
xor XOR2 (N544, N537, N34);
not NOT1 (N545, N535);
nor NOR3 (N546, N545, N67, N22);
nor NOR3 (N547, N530, N84, N452);
and AND2 (N548, N538, N143);
nand NAND2 (N549, N542, N71);
and AND4 (N550, N524, N119, N228, N278);
buf BUF1 (N551, N543);
and AND2 (N552, N547, N475);
xor XOR2 (N553, N549, N511);
and AND3 (N554, N552, N439, N324);
nor NOR4 (N555, N548, N277, N437, N6);
buf BUF1 (N556, N536);
nor NOR2 (N557, N553, N146);
and AND3 (N558, N546, N46, N115);
or OR4 (N559, N544, N397, N48, N507);
or OR4 (N560, N539, N49, N525, N219);
nand NAND3 (N561, N556, N401, N291);
buf BUF1 (N562, N550);
nand NAND3 (N563, N560, N1, N120);
and AND3 (N564, N558, N257, N481);
nand NAND2 (N565, N564, N16);
or OR2 (N566, N565, N140);
not NOT1 (N567, N551);
and AND3 (N568, N559, N338, N301);
not NOT1 (N569, N563);
not NOT1 (N570, N566);
and AND3 (N571, N569, N8, N394);
nand NAND3 (N572, N534, N77, N394);
or OR4 (N573, N555, N527, N64, N370);
nor NOR4 (N574, N554, N149, N294, N318);
xor XOR2 (N575, N570, N343);
xor XOR2 (N576, N571, N435);
xor XOR2 (N577, N573, N226);
and AND3 (N578, N574, N460, N399);
buf BUF1 (N579, N567);
not NOT1 (N580, N561);
or OR3 (N581, N562, N130, N378);
or OR4 (N582, N557, N427, N114, N48);
or OR2 (N583, N582, N481);
and AND4 (N584, N572, N46, N215, N174);
not NOT1 (N585, N576);
xor XOR2 (N586, N584, N523);
nand NAND3 (N587, N568, N424, N418);
xor XOR2 (N588, N583, N189);
buf BUF1 (N589, N585);
nor NOR4 (N590, N578, N320, N253, N433);
or OR4 (N591, N577, N397, N140, N386);
nor NOR2 (N592, N581, N582);
nor NOR4 (N593, N587, N372, N523, N129);
buf BUF1 (N594, N591);
or OR4 (N595, N580, N75, N516, N463);
nand NAND3 (N596, N592, N522, N353);
or OR3 (N597, N575, N374, N51);
xor XOR2 (N598, N589, N505);
or OR2 (N599, N586, N549);
not NOT1 (N600, N579);
not NOT1 (N601, N593);
or OR3 (N602, N594, N62, N490);
buf BUF1 (N603, N599);
nand NAND2 (N604, N603, N130);
buf BUF1 (N605, N602);
not NOT1 (N606, N590);
buf BUF1 (N607, N588);
not NOT1 (N608, N606);
or OR3 (N609, N597, N296, N228);
buf BUF1 (N610, N600);
buf BUF1 (N611, N605);
nand NAND2 (N612, N596, N478);
nand NAND2 (N613, N598, N317);
or OR2 (N614, N610, N265);
buf BUF1 (N615, N601);
and AND4 (N616, N612, N218, N78, N325);
nor NOR2 (N617, N608, N199);
buf BUF1 (N618, N604);
or OR4 (N619, N614, N221, N433, N382);
not NOT1 (N620, N611);
and AND4 (N621, N619, N348, N215, N228);
buf BUF1 (N622, N607);
buf BUF1 (N623, N616);
buf BUF1 (N624, N595);
buf BUF1 (N625, N618);
or OR3 (N626, N620, N187, N196);
xor XOR2 (N627, N625, N453);
buf BUF1 (N628, N621);
buf BUF1 (N629, N627);
buf BUF1 (N630, N626);
not NOT1 (N631, N609);
buf BUF1 (N632, N622);
nand NAND3 (N633, N630, N36, N169);
not NOT1 (N634, N623);
buf BUF1 (N635, N624);
xor XOR2 (N636, N613, N391);
and AND2 (N637, N615, N490);
nand NAND2 (N638, N637, N321);
not NOT1 (N639, N628);
and AND4 (N640, N633, N197, N613, N415);
and AND2 (N641, N640, N367);
buf BUF1 (N642, N641);
buf BUF1 (N643, N629);
not NOT1 (N644, N617);
nor NOR4 (N645, N634, N459, N615, N120);
nand NAND4 (N646, N639, N427, N599, N15);
buf BUF1 (N647, N643);
buf BUF1 (N648, N635);
nor NOR2 (N649, N645, N13);
xor XOR2 (N650, N632, N591);
and AND2 (N651, N648, N301);
nor NOR3 (N652, N631, N530, N345);
and AND4 (N653, N651, N257, N647, N149);
buf BUF1 (N654, N467);
nor NOR2 (N655, N636, N366);
and AND3 (N656, N655, N176, N587);
nand NAND2 (N657, N644, N368);
and AND2 (N658, N654, N179);
nand NAND2 (N659, N653, N113);
buf BUF1 (N660, N649);
xor XOR2 (N661, N657, N324);
and AND3 (N662, N638, N611, N335);
nor NOR3 (N663, N660, N228, N448);
xor XOR2 (N664, N663, N565);
and AND2 (N665, N650, N557);
and AND4 (N666, N658, N17, N94, N367);
buf BUF1 (N667, N652);
and AND2 (N668, N642, N622);
nand NAND4 (N669, N668, N356, N285, N461);
or OR2 (N670, N666, N450);
not NOT1 (N671, N665);
xor XOR2 (N672, N670, N605);
nor NOR3 (N673, N669, N273, N267);
not NOT1 (N674, N646);
nor NOR3 (N675, N661, N456, N657);
not NOT1 (N676, N659);
xor XOR2 (N677, N667, N591);
xor XOR2 (N678, N677, N111);
nand NAND3 (N679, N664, N318, N486);
buf BUF1 (N680, N671);
or OR3 (N681, N674, N340, N408);
nor NOR4 (N682, N672, N498, N356, N56);
nand NAND3 (N683, N678, N498, N355);
nand NAND4 (N684, N656, N305, N20, N540);
nor NOR2 (N685, N682, N347);
xor XOR2 (N686, N675, N88);
nand NAND3 (N687, N681, N591, N587);
not NOT1 (N688, N685);
buf BUF1 (N689, N687);
or OR3 (N690, N662, N207, N602);
xor XOR2 (N691, N688, N665);
nand NAND2 (N692, N689, N104);
and AND2 (N693, N691, N189);
nand NAND4 (N694, N680, N674, N445, N196);
or OR4 (N695, N693, N158, N632, N415);
and AND4 (N696, N686, N141, N641, N601);
buf BUF1 (N697, N696);
nor NOR3 (N698, N694, N392, N181);
and AND2 (N699, N695, N341);
nand NAND4 (N700, N692, N38, N68, N458);
or OR2 (N701, N690, N143);
xor XOR2 (N702, N698, N151);
nor NOR3 (N703, N700, N474, N269);
buf BUF1 (N704, N683);
xor XOR2 (N705, N704, N377);
nand NAND2 (N706, N705, N373);
nand NAND4 (N707, N673, N223, N73, N566);
nand NAND3 (N708, N679, N258, N420);
nand NAND4 (N709, N699, N110, N83, N525);
and AND2 (N710, N676, N118);
nor NOR4 (N711, N709, N407, N527, N173);
xor XOR2 (N712, N697, N589);
nor NOR2 (N713, N706, N256);
nor NOR4 (N714, N702, N264, N324, N572);
nor NOR2 (N715, N714, N452);
and AND2 (N716, N712, N572);
buf BUF1 (N717, N701);
or OR3 (N718, N684, N342, N552);
nand NAND4 (N719, N717, N312, N574, N455);
buf BUF1 (N720, N703);
not NOT1 (N721, N710);
not NOT1 (N722, N708);
nor NOR3 (N723, N720, N141, N453);
and AND2 (N724, N718, N162);
buf BUF1 (N725, N713);
or OR2 (N726, N722, N46);
nand NAND4 (N727, N721, N408, N197, N615);
not NOT1 (N728, N707);
nor NOR4 (N729, N716, N89, N205, N120);
nor NOR4 (N730, N725, N408, N72, N714);
not NOT1 (N731, N730);
or OR2 (N732, N726, N444);
nand NAND2 (N733, N729, N318);
nand NAND4 (N734, N715, N399, N598, N382);
buf BUF1 (N735, N728);
xor XOR2 (N736, N719, N440);
and AND4 (N737, N723, N113, N669, N658);
xor XOR2 (N738, N724, N318);
xor XOR2 (N739, N727, N728);
buf BUF1 (N740, N733);
and AND3 (N741, N739, N156, N687);
not NOT1 (N742, N711);
nor NOR3 (N743, N732, N316, N319);
buf BUF1 (N744, N740);
xor XOR2 (N745, N735, N465);
nor NOR2 (N746, N731, N131);
and AND3 (N747, N741, N108, N545);
nor NOR2 (N748, N744, N16);
xor XOR2 (N749, N745, N86);
not NOT1 (N750, N737);
or OR3 (N751, N747, N608, N93);
buf BUF1 (N752, N748);
buf BUF1 (N753, N736);
buf BUF1 (N754, N743);
not NOT1 (N755, N751);
nand NAND3 (N756, N752, N76, N454);
buf BUF1 (N757, N750);
xor XOR2 (N758, N756, N212);
and AND4 (N759, N755, N55, N292, N704);
or OR4 (N760, N754, N289, N29, N332);
and AND4 (N761, N753, N627, N135, N309);
or OR2 (N762, N761, N500);
xor XOR2 (N763, N746, N607);
buf BUF1 (N764, N749);
not NOT1 (N765, N738);
and AND2 (N766, N760, N507);
buf BUF1 (N767, N765);
and AND3 (N768, N759, N190, N251);
buf BUF1 (N769, N734);
xor XOR2 (N770, N768, N597);
or OR3 (N771, N763, N757, N218);
buf BUF1 (N772, N575);
buf BUF1 (N773, N770);
buf BUF1 (N774, N773);
or OR4 (N775, N769, N87, N389, N292);
buf BUF1 (N776, N764);
or OR2 (N777, N775, N613);
buf BUF1 (N778, N742);
nand NAND4 (N779, N758, N78, N353, N82);
buf BUF1 (N780, N767);
not NOT1 (N781, N771);
not NOT1 (N782, N776);
nand NAND4 (N783, N777, N111, N106, N678);
or OR4 (N784, N778, N192, N647, N91);
not NOT1 (N785, N772);
not NOT1 (N786, N782);
xor XOR2 (N787, N783, N578);
or OR4 (N788, N784, N713, N486, N376);
nand NAND4 (N789, N766, N474, N114, N535);
buf BUF1 (N790, N788);
xor XOR2 (N791, N781, N118);
xor XOR2 (N792, N785, N277);
and AND3 (N793, N792, N489, N115);
xor XOR2 (N794, N793, N758);
buf BUF1 (N795, N787);
or OR2 (N796, N780, N36);
xor XOR2 (N797, N791, N763);
nand NAND4 (N798, N794, N253, N59, N671);
xor XOR2 (N799, N797, N153);
not NOT1 (N800, N798);
buf BUF1 (N801, N789);
xor XOR2 (N802, N790, N141);
not NOT1 (N803, N779);
buf BUF1 (N804, N786);
nand NAND3 (N805, N795, N344, N418);
or OR3 (N806, N804, N751, N182);
and AND4 (N807, N805, N661, N520, N604);
nor NOR4 (N808, N802, N452, N64, N359);
nand NAND4 (N809, N762, N794, N31, N639);
or OR4 (N810, N806, N629, N172, N746);
xor XOR2 (N811, N799, N469);
and AND4 (N812, N796, N171, N48, N360);
and AND3 (N813, N803, N643, N808);
and AND2 (N814, N94, N653);
or OR3 (N815, N812, N722, N176);
xor XOR2 (N816, N800, N530);
or OR4 (N817, N801, N794, N209, N640);
buf BUF1 (N818, N817);
or OR4 (N819, N774, N430, N396, N212);
xor XOR2 (N820, N818, N18);
buf BUF1 (N821, N809);
not NOT1 (N822, N820);
xor XOR2 (N823, N815, N811);
and AND4 (N824, N662, N57, N201, N144);
and AND3 (N825, N822, N369, N759);
not NOT1 (N826, N810);
and AND2 (N827, N825, N607);
or OR4 (N828, N824, N807, N227, N54);
and AND2 (N829, N567, N90);
xor XOR2 (N830, N821, N791);
not NOT1 (N831, N816);
buf BUF1 (N832, N827);
not NOT1 (N833, N814);
buf BUF1 (N834, N813);
nor NOR3 (N835, N823, N825, N439);
and AND3 (N836, N828, N309, N337);
nand NAND4 (N837, N830, N320, N414, N49);
and AND4 (N838, N831, N278, N746, N718);
or OR3 (N839, N829, N256, N805);
buf BUF1 (N840, N837);
not NOT1 (N841, N840);
or OR2 (N842, N819, N67);
buf BUF1 (N843, N834);
and AND4 (N844, N826, N480, N740, N264);
nor NOR3 (N845, N838, N721, N173);
or OR3 (N846, N835, N541, N795);
xor XOR2 (N847, N845, N106);
and AND3 (N848, N832, N334, N818);
nor NOR3 (N849, N836, N748, N522);
xor XOR2 (N850, N842, N461);
nand NAND4 (N851, N848, N216, N779, N276);
buf BUF1 (N852, N833);
not NOT1 (N853, N852);
not NOT1 (N854, N843);
or OR4 (N855, N841, N518, N19, N624);
xor XOR2 (N856, N846, N164);
not NOT1 (N857, N844);
xor XOR2 (N858, N854, N435);
or OR2 (N859, N857, N630);
not NOT1 (N860, N858);
xor XOR2 (N861, N860, N72);
not NOT1 (N862, N856);
xor XOR2 (N863, N849, N141);
nand NAND4 (N864, N839, N282, N118, N410);
buf BUF1 (N865, N850);
nand NAND3 (N866, N861, N405, N322);
xor XOR2 (N867, N862, N156);
nor NOR3 (N868, N865, N494, N586);
not NOT1 (N869, N853);
nor NOR4 (N870, N847, N809, N648, N605);
nor NOR3 (N871, N866, N423, N90);
buf BUF1 (N872, N855);
not NOT1 (N873, N867);
not NOT1 (N874, N871);
or OR4 (N875, N864, N335, N111, N356);
nor NOR4 (N876, N859, N301, N120, N268);
xor XOR2 (N877, N869, N369);
nand NAND4 (N878, N863, N123, N245, N45);
nand NAND4 (N879, N875, N422, N769, N650);
nand NAND2 (N880, N874, N419);
nand NAND2 (N881, N880, N283);
nor NOR3 (N882, N877, N821, N288);
xor XOR2 (N883, N870, N263);
nand NAND2 (N884, N878, N45);
not NOT1 (N885, N851);
not NOT1 (N886, N885);
not NOT1 (N887, N879);
buf BUF1 (N888, N876);
nand NAND3 (N889, N868, N581, N309);
buf BUF1 (N890, N883);
or OR3 (N891, N888, N85, N31);
nand NAND3 (N892, N873, N33, N15);
nand NAND3 (N893, N882, N880, N881);
and AND3 (N894, N324, N110, N568);
or OR2 (N895, N891, N100);
nand NAND4 (N896, N894, N604, N744, N155);
nand NAND3 (N897, N872, N226, N866);
nor NOR3 (N898, N886, N627, N617);
xor XOR2 (N899, N897, N405);
nand NAND2 (N900, N889, N569);
buf BUF1 (N901, N893);
nand NAND3 (N902, N898, N698, N875);
xor XOR2 (N903, N901, N567);
and AND2 (N904, N903, N840);
or OR4 (N905, N884, N792, N284, N44);
not NOT1 (N906, N904);
nor NOR4 (N907, N890, N416, N160, N392);
nand NAND2 (N908, N899, N281);
not NOT1 (N909, N906);
buf BUF1 (N910, N900);
buf BUF1 (N911, N905);
xor XOR2 (N912, N907, N111);
xor XOR2 (N913, N911, N759);
buf BUF1 (N914, N902);
nand NAND2 (N915, N908, N23);
buf BUF1 (N916, N914);
or OR3 (N917, N909, N370, N278);
buf BUF1 (N918, N912);
or OR4 (N919, N913, N138, N796, N916);
nor NOR3 (N920, N806, N77, N650);
nor NOR3 (N921, N887, N293, N484);
xor XOR2 (N922, N895, N72);
xor XOR2 (N923, N910, N441);
not NOT1 (N924, N915);
not NOT1 (N925, N896);
nand NAND2 (N926, N921, N201);
and AND2 (N927, N925, N396);
buf BUF1 (N928, N892);
not NOT1 (N929, N924);
and AND4 (N930, N920, N291, N854, N660);
buf BUF1 (N931, N918);
or OR4 (N932, N923, N466, N666, N58);
or OR2 (N933, N919, N83);
xor XOR2 (N934, N928, N139);
nand NAND2 (N935, N917, N811);
and AND2 (N936, N935, N130);
buf BUF1 (N937, N936);
nor NOR2 (N938, N922, N706);
nor NOR2 (N939, N938, N659);
xor XOR2 (N940, N934, N816);
not NOT1 (N941, N937);
nor NOR4 (N942, N927, N313, N470, N603);
and AND3 (N943, N939, N762, N134);
xor XOR2 (N944, N932, N451);
and AND3 (N945, N931, N429, N544);
and AND2 (N946, N944, N175);
and AND4 (N947, N933, N385, N561, N854);
and AND2 (N948, N930, N878);
nand NAND4 (N949, N940, N594, N410, N707);
buf BUF1 (N950, N943);
nor NOR2 (N951, N929, N645);
nor NOR2 (N952, N951, N920);
buf BUF1 (N953, N926);
xor XOR2 (N954, N948, N880);
nor NOR3 (N955, N950, N827, N500);
xor XOR2 (N956, N953, N916);
nand NAND4 (N957, N945, N722, N438, N636);
nand NAND4 (N958, N947, N54, N371, N527);
nand NAND4 (N959, N955, N725, N309, N829);
nor NOR2 (N960, N952, N447);
nor NOR3 (N961, N957, N727, N874);
xor XOR2 (N962, N946, N825);
and AND3 (N963, N958, N618, N383);
nand NAND4 (N964, N949, N471, N223, N198);
or OR2 (N965, N960, N804);
or OR2 (N966, N965, N145);
nor NOR4 (N967, N941, N172, N587, N203);
xor XOR2 (N968, N956, N656);
nor NOR4 (N969, N942, N297, N506, N225);
nand NAND3 (N970, N969, N218, N397);
not NOT1 (N971, N968);
nor NOR4 (N972, N964, N877, N468, N287);
buf BUF1 (N973, N954);
and AND4 (N974, N961, N157, N926, N522);
and AND2 (N975, N967, N612);
nand NAND3 (N976, N971, N79, N639);
and AND2 (N977, N973, N556);
or OR2 (N978, N970, N947);
buf BUF1 (N979, N959);
xor XOR2 (N980, N966, N657);
nor NOR4 (N981, N963, N486, N485, N115);
nor NOR4 (N982, N979, N441, N661, N88);
or OR3 (N983, N972, N212, N318);
nor NOR3 (N984, N977, N68, N194);
buf BUF1 (N985, N983);
xor XOR2 (N986, N982, N351);
buf BUF1 (N987, N974);
xor XOR2 (N988, N981, N540);
nand NAND4 (N989, N978, N894, N139, N263);
and AND2 (N990, N976, N44);
buf BUF1 (N991, N989);
xor XOR2 (N992, N962, N223);
and AND2 (N993, N980, N574);
or OR2 (N994, N984, N91);
buf BUF1 (N995, N993);
not NOT1 (N996, N987);
not NOT1 (N997, N992);
not NOT1 (N998, N986);
nor NOR3 (N999, N990, N889, N182);
buf BUF1 (N1000, N985);
nor NOR3 (N1001, N995, N342, N495);
nand NAND3 (N1002, N1001, N532, N969);
buf BUF1 (N1003, N1000);
nand NAND4 (N1004, N994, N544, N805, N708);
nor NOR4 (N1005, N975, N986, N318, N80);
not NOT1 (N1006, N1004);
buf BUF1 (N1007, N1002);
or OR2 (N1008, N999, N977);
xor XOR2 (N1009, N998, N640);
xor XOR2 (N1010, N996, N67);
buf BUF1 (N1011, N997);
and AND4 (N1012, N988, N148, N668, N262);
xor XOR2 (N1013, N1003, N370);
buf BUF1 (N1014, N1009);
and AND2 (N1015, N1010, N238);
nor NOR4 (N1016, N1014, N534, N472, N669);
nand NAND3 (N1017, N1007, N600, N427);
buf BUF1 (N1018, N1012);
or OR4 (N1019, N1018, N879, N590, N907);
or OR4 (N1020, N991, N1012, N550, N667);
or OR3 (N1021, N1006, N512, N803);
buf BUF1 (N1022, N1020);
nor NOR3 (N1023, N1015, N244, N889);
or OR3 (N1024, N1005, N323, N472);
buf BUF1 (N1025, N1008);
nand NAND4 (N1026, N1021, N879, N939, N888);
or OR3 (N1027, N1022, N960, N475);
and AND3 (N1028, N1027, N749, N665);
or OR4 (N1029, N1023, N384, N364, N907);
and AND2 (N1030, N1017, N476);
and AND2 (N1031, N1030, N999);
xor XOR2 (N1032, N1019, N714);
nand NAND2 (N1033, N1028, N760);
and AND3 (N1034, N1024, N21, N343);
or OR4 (N1035, N1026, N674, N437, N30);
buf BUF1 (N1036, N1032);
or OR2 (N1037, N1013, N894);
not NOT1 (N1038, N1035);
xor XOR2 (N1039, N1036, N246);
nor NOR2 (N1040, N1038, N424);
xor XOR2 (N1041, N1025, N563);
and AND2 (N1042, N1039, N504);
or OR3 (N1043, N1041, N872, N621);
nor NOR4 (N1044, N1011, N240, N831, N47);
nand NAND2 (N1045, N1016, N968);
nand NAND4 (N1046, N1031, N800, N413, N1012);
buf BUF1 (N1047, N1037);
xor XOR2 (N1048, N1042, N844);
buf BUF1 (N1049, N1033);
or OR3 (N1050, N1029, N665, N374);
not NOT1 (N1051, N1048);
xor XOR2 (N1052, N1034, N260);
not NOT1 (N1053, N1049);
nand NAND2 (N1054, N1050, N834);
nand NAND4 (N1055, N1046, N452, N3, N391);
and AND4 (N1056, N1055, N955, N503, N946);
or OR3 (N1057, N1051, N63, N774);
and AND4 (N1058, N1040, N483, N682, N297);
buf BUF1 (N1059, N1052);
xor XOR2 (N1060, N1057, N901);
xor XOR2 (N1061, N1045, N400);
nor NOR4 (N1062, N1061, N401, N134, N450);
nand NAND4 (N1063, N1056, N421, N193, N268);
buf BUF1 (N1064, N1054);
buf BUF1 (N1065, N1062);
nor NOR2 (N1066, N1053, N194);
and AND2 (N1067, N1065, N426);
buf BUF1 (N1068, N1058);
xor XOR2 (N1069, N1060, N1001);
not NOT1 (N1070, N1044);
not NOT1 (N1071, N1059);
nand NAND4 (N1072, N1063, N177, N160, N1047);
buf BUF1 (N1073, N96);
or OR2 (N1074, N1071, N74);
and AND2 (N1075, N1072, N583);
nand NAND2 (N1076, N1064, N407);
nand NAND4 (N1077, N1066, N416, N879, N725);
buf BUF1 (N1078, N1068);
nand NAND2 (N1079, N1073, N596);
or OR3 (N1080, N1043, N453, N429);
nor NOR2 (N1081, N1078, N265);
and AND2 (N1082, N1075, N412);
xor XOR2 (N1083, N1069, N838);
or OR4 (N1084, N1080, N47, N460, N318);
or OR2 (N1085, N1081, N50);
buf BUF1 (N1086, N1067);
and AND2 (N1087, N1084, N29);
nand NAND2 (N1088, N1070, N414);
not NOT1 (N1089, N1079);
nor NOR2 (N1090, N1087, N236);
and AND3 (N1091, N1076, N874, N388);
buf BUF1 (N1092, N1074);
nand NAND3 (N1093, N1086, N983, N435);
nor NOR4 (N1094, N1088, N357, N313, N1056);
nor NOR4 (N1095, N1082, N851, N516, N422);
buf BUF1 (N1096, N1095);
and AND3 (N1097, N1083, N219, N731);
buf BUF1 (N1098, N1089);
nand NAND4 (N1099, N1096, N1086, N141, N893);
buf BUF1 (N1100, N1094);
not NOT1 (N1101, N1090);
nand NAND4 (N1102, N1085, N671, N234, N344);
xor XOR2 (N1103, N1091, N1039);
not NOT1 (N1104, N1097);
and AND3 (N1105, N1098, N290, N416);
nor NOR4 (N1106, N1100, N584, N813, N202);
or OR2 (N1107, N1103, N841);
and AND3 (N1108, N1101, N637, N644);
or OR3 (N1109, N1092, N1107, N718);
buf BUF1 (N1110, N70);
not NOT1 (N1111, N1110);
nor NOR3 (N1112, N1108, N295, N937);
nand NAND2 (N1113, N1102, N1090);
buf BUF1 (N1114, N1106);
not NOT1 (N1115, N1093);
or OR4 (N1116, N1077, N82, N420, N830);
not NOT1 (N1117, N1113);
not NOT1 (N1118, N1112);
or OR3 (N1119, N1111, N775, N247);
xor XOR2 (N1120, N1115, N986);
xor XOR2 (N1121, N1105, N207);
nor NOR2 (N1122, N1121, N488);
nand NAND4 (N1123, N1119, N482, N627, N771);
nand NAND3 (N1124, N1123, N1084, N737);
not NOT1 (N1125, N1122);
not NOT1 (N1126, N1125);
not NOT1 (N1127, N1109);
nand NAND4 (N1128, N1104, N434, N621, N853);
not NOT1 (N1129, N1126);
not NOT1 (N1130, N1128);
and AND4 (N1131, N1127, N139, N928, N204);
and AND4 (N1132, N1118, N485, N154, N780);
nor NOR4 (N1133, N1131, N109, N176, N145);
nand NAND2 (N1134, N1130, N1059);
buf BUF1 (N1135, N1134);
and AND4 (N1136, N1116, N744, N944, N345);
nand NAND2 (N1137, N1133, N436);
nor NOR3 (N1138, N1132, N770, N1072);
or OR4 (N1139, N1099, N507, N1124, N646);
and AND4 (N1140, N668, N549, N847, N1028);
and AND4 (N1141, N1120, N637, N316, N1009);
or OR3 (N1142, N1138, N929, N189);
buf BUF1 (N1143, N1141);
or OR2 (N1144, N1117, N942);
nor NOR4 (N1145, N1136, N48, N701, N1020);
buf BUF1 (N1146, N1139);
nor NOR4 (N1147, N1137, N425, N742, N695);
not NOT1 (N1148, N1146);
or OR3 (N1149, N1148, N815, N1073);
and AND2 (N1150, N1144, N374);
or OR2 (N1151, N1143, N664);
not NOT1 (N1152, N1151);
not NOT1 (N1153, N1147);
and AND4 (N1154, N1153, N669, N933, N87);
not NOT1 (N1155, N1114);
not NOT1 (N1156, N1140);
buf BUF1 (N1157, N1156);
nor NOR3 (N1158, N1145, N233, N71);
xor XOR2 (N1159, N1129, N828);
and AND4 (N1160, N1158, N1051, N972, N1044);
or OR4 (N1161, N1160, N843, N988, N22);
or OR3 (N1162, N1155, N414, N588);
or OR4 (N1163, N1161, N360, N88, N806);
xor XOR2 (N1164, N1159, N1132);
xor XOR2 (N1165, N1149, N686);
xor XOR2 (N1166, N1157, N463);
xor XOR2 (N1167, N1142, N289);
and AND3 (N1168, N1150, N284, N80);
nor NOR4 (N1169, N1165, N718, N233, N1054);
and AND2 (N1170, N1162, N827);
nor NOR3 (N1171, N1164, N747, N1024);
and AND3 (N1172, N1168, N29, N9);
buf BUF1 (N1173, N1135);
xor XOR2 (N1174, N1173, N1094);
xor XOR2 (N1175, N1174, N893);
not NOT1 (N1176, N1170);
or OR2 (N1177, N1171, N545);
buf BUF1 (N1178, N1152);
or OR3 (N1179, N1154, N1123, N1015);
and AND4 (N1180, N1178, N1156, N578, N447);
nand NAND2 (N1181, N1167, N477);
buf BUF1 (N1182, N1169);
buf BUF1 (N1183, N1163);
and AND3 (N1184, N1182, N248, N675);
or OR3 (N1185, N1177, N835, N577);
or OR3 (N1186, N1183, N329, N880);
or OR2 (N1187, N1185, N986);
or OR4 (N1188, N1176, N1059, N457, N540);
buf BUF1 (N1189, N1172);
nor NOR3 (N1190, N1179, N851, N769);
nor NOR4 (N1191, N1184, N178, N1007, N722);
not NOT1 (N1192, N1166);
nor NOR3 (N1193, N1186, N844, N608);
xor XOR2 (N1194, N1189, N434);
or OR3 (N1195, N1192, N1089, N561);
xor XOR2 (N1196, N1191, N502);
xor XOR2 (N1197, N1188, N993);
and AND4 (N1198, N1194, N971, N587, N996);
nor NOR2 (N1199, N1195, N1161);
or OR2 (N1200, N1199, N983);
nand NAND3 (N1201, N1175, N1003, N1149);
and AND3 (N1202, N1201, N994, N178);
or OR3 (N1203, N1198, N730, N84);
or OR4 (N1204, N1196, N63, N298, N276);
not NOT1 (N1205, N1202);
not NOT1 (N1206, N1180);
or OR4 (N1207, N1197, N249, N734, N776);
nand NAND3 (N1208, N1205, N860, N46);
nand NAND3 (N1209, N1207, N1048, N661);
and AND2 (N1210, N1181, N801);
or OR2 (N1211, N1200, N601);
buf BUF1 (N1212, N1204);
and AND3 (N1213, N1187, N35, N1149);
not NOT1 (N1214, N1190);
xor XOR2 (N1215, N1206, N800);
buf BUF1 (N1216, N1214);
nor NOR3 (N1217, N1212, N456, N1105);
and AND4 (N1218, N1209, N63, N942, N599);
nor NOR4 (N1219, N1208, N60, N426, N1132);
and AND3 (N1220, N1211, N619, N295);
buf BUF1 (N1221, N1203);
nor NOR3 (N1222, N1210, N438, N125);
not NOT1 (N1223, N1213);
and AND4 (N1224, N1218, N224, N150, N886);
xor XOR2 (N1225, N1217, N458);
buf BUF1 (N1226, N1221);
buf BUF1 (N1227, N1226);
not NOT1 (N1228, N1223);
buf BUF1 (N1229, N1222);
xor XOR2 (N1230, N1227, N641);
and AND4 (N1231, N1228, N521, N182, N646);
and AND3 (N1232, N1193, N395, N1119);
xor XOR2 (N1233, N1215, N144);
nand NAND2 (N1234, N1229, N241);
or OR4 (N1235, N1234, N900, N978, N1187);
not NOT1 (N1236, N1232);
buf BUF1 (N1237, N1224);
or OR2 (N1238, N1231, N520);
or OR4 (N1239, N1219, N160, N776, N713);
not NOT1 (N1240, N1233);
nor NOR2 (N1241, N1237, N569);
nand NAND4 (N1242, N1240, N671, N623, N896);
or OR4 (N1243, N1230, N1112, N1205, N857);
nor NOR4 (N1244, N1243, N1051, N1006, N298);
xor XOR2 (N1245, N1216, N966);
nand NAND3 (N1246, N1239, N811, N33);
nand NAND2 (N1247, N1244, N245);
or OR4 (N1248, N1235, N77, N672, N1104);
nor NOR4 (N1249, N1247, N400, N576, N1075);
buf BUF1 (N1250, N1246);
xor XOR2 (N1251, N1238, N1171);
nor NOR3 (N1252, N1241, N255, N221);
nor NOR2 (N1253, N1220, N752);
not NOT1 (N1254, N1245);
nand NAND2 (N1255, N1252, N263);
nor NOR3 (N1256, N1255, N282, N920);
nand NAND2 (N1257, N1249, N300);
not NOT1 (N1258, N1254);
or OR4 (N1259, N1236, N1041, N1011, N979);
xor XOR2 (N1260, N1257, N472);
nor NOR4 (N1261, N1250, N420, N648, N833);
or OR2 (N1262, N1260, N882);
and AND2 (N1263, N1261, N678);
xor XOR2 (N1264, N1262, N370);
nand NAND4 (N1265, N1225, N425, N551, N706);
not NOT1 (N1266, N1258);
buf BUF1 (N1267, N1242);
not NOT1 (N1268, N1248);
buf BUF1 (N1269, N1256);
and AND3 (N1270, N1268, N325, N1047);
buf BUF1 (N1271, N1265);
nand NAND4 (N1272, N1259, N432, N791, N576);
not NOT1 (N1273, N1269);
nand NAND4 (N1274, N1271, N1065, N15, N191);
buf BUF1 (N1275, N1251);
nand NAND2 (N1276, N1273, N918);
xor XOR2 (N1277, N1274, N460);
xor XOR2 (N1278, N1276, N1118);
nand NAND2 (N1279, N1272, N636);
or OR2 (N1280, N1278, N875);
nor NOR2 (N1281, N1280, N483);
and AND4 (N1282, N1275, N269, N302, N437);
nand NAND3 (N1283, N1281, N1145, N1074);
buf BUF1 (N1284, N1279);
and AND4 (N1285, N1263, N394, N463, N278);
or OR2 (N1286, N1282, N810);
not NOT1 (N1287, N1266);
buf BUF1 (N1288, N1283);
nor NOR3 (N1289, N1253, N229, N767);
xor XOR2 (N1290, N1277, N115);
xor XOR2 (N1291, N1284, N436);
nand NAND4 (N1292, N1288, N45, N185, N19);
or OR2 (N1293, N1289, N322);
nand NAND2 (N1294, N1286, N540);
buf BUF1 (N1295, N1287);
nand NAND4 (N1296, N1290, N986, N133, N1279);
xor XOR2 (N1297, N1295, N913);
xor XOR2 (N1298, N1296, N186);
and AND2 (N1299, N1285, N211);
or OR3 (N1300, N1299, N312, N56);
nor NOR2 (N1301, N1264, N136);
nor NOR2 (N1302, N1270, N1293);
nor NOR2 (N1303, N20, N96);
and AND4 (N1304, N1300, N520, N1059, N1173);
nor NOR3 (N1305, N1302, N293, N110);
nor NOR4 (N1306, N1304, N40, N165, N475);
buf BUF1 (N1307, N1297);
not NOT1 (N1308, N1307);
nand NAND2 (N1309, N1292, N517);
buf BUF1 (N1310, N1306);
nand NAND2 (N1311, N1309, N304);
nor NOR3 (N1312, N1305, N841, N219);
nor NOR4 (N1313, N1310, N376, N689, N865);
or OR3 (N1314, N1308, N466, N715);
nand NAND3 (N1315, N1303, N787, N106);
nor NOR3 (N1316, N1267, N1239, N1193);
xor XOR2 (N1317, N1313, N892);
xor XOR2 (N1318, N1315, N526);
xor XOR2 (N1319, N1291, N483);
nand NAND2 (N1320, N1319, N954);
not NOT1 (N1321, N1317);
nand NAND4 (N1322, N1318, N147, N890, N549);
and AND2 (N1323, N1321, N1285);
buf BUF1 (N1324, N1323);
nor NOR2 (N1325, N1314, N1105);
nor NOR2 (N1326, N1301, N325);
not NOT1 (N1327, N1325);
nand NAND4 (N1328, N1312, N1202, N1157, N784);
xor XOR2 (N1329, N1320, N565);
nand NAND4 (N1330, N1316, N1283, N773, N41);
nor NOR4 (N1331, N1324, N873, N857, N983);
buf BUF1 (N1332, N1322);
xor XOR2 (N1333, N1332, N661);
not NOT1 (N1334, N1331);
and AND4 (N1335, N1333, N447, N871, N965);
or OR4 (N1336, N1311, N368, N957, N980);
and AND3 (N1337, N1294, N1109, N520);
xor XOR2 (N1338, N1328, N788);
nor NOR4 (N1339, N1334, N1146, N315, N1051);
or OR3 (N1340, N1338, N258, N458);
nor NOR4 (N1341, N1330, N149, N1274, N550);
buf BUF1 (N1342, N1339);
xor XOR2 (N1343, N1336, N420);
buf BUF1 (N1344, N1335);
or OR2 (N1345, N1329, N1025);
not NOT1 (N1346, N1342);
not NOT1 (N1347, N1343);
buf BUF1 (N1348, N1347);
or OR3 (N1349, N1344, N418, N295);
nor NOR4 (N1350, N1346, N460, N1266, N876);
or OR2 (N1351, N1341, N845);
buf BUF1 (N1352, N1340);
nor NOR4 (N1353, N1352, N96, N756, N446);
nor NOR4 (N1354, N1351, N194, N410, N529);
buf BUF1 (N1355, N1337);
xor XOR2 (N1356, N1326, N849);
buf BUF1 (N1357, N1354);
not NOT1 (N1358, N1348);
nor NOR4 (N1359, N1349, N956, N739, N289);
nor NOR4 (N1360, N1359, N298, N592, N1056);
or OR4 (N1361, N1355, N223, N883, N531);
xor XOR2 (N1362, N1360, N371);
nor NOR2 (N1363, N1356, N272);
or OR3 (N1364, N1361, N1315, N432);
nor NOR4 (N1365, N1357, N388, N924, N764);
not NOT1 (N1366, N1358);
nand NAND3 (N1367, N1298, N426, N241);
not NOT1 (N1368, N1350);
xor XOR2 (N1369, N1368, N768);
buf BUF1 (N1370, N1369);
and AND2 (N1371, N1370, N147);
or OR2 (N1372, N1363, N385);
nand NAND4 (N1373, N1367, N495, N805, N470);
buf BUF1 (N1374, N1364);
buf BUF1 (N1375, N1365);
or OR3 (N1376, N1362, N474, N1189);
not NOT1 (N1377, N1327);
or OR4 (N1378, N1371, N229, N967, N1369);
buf BUF1 (N1379, N1376);
not NOT1 (N1380, N1378);
and AND4 (N1381, N1345, N270, N77, N73);
and AND3 (N1382, N1374, N1048, N219);
buf BUF1 (N1383, N1380);
or OR3 (N1384, N1379, N496, N1110);
and AND2 (N1385, N1373, N1301);
xor XOR2 (N1386, N1385, N1229);
not NOT1 (N1387, N1377);
and AND3 (N1388, N1381, N1322, N295);
nor NOR4 (N1389, N1384, N276, N501, N1028);
buf BUF1 (N1390, N1366);
and AND3 (N1391, N1388, N286, N1239);
nor NOR3 (N1392, N1387, N5, N572);
and AND3 (N1393, N1392, N1114, N209);
nand NAND2 (N1394, N1390, N405);
not NOT1 (N1395, N1382);
not NOT1 (N1396, N1389);
and AND2 (N1397, N1395, N744);
nor NOR3 (N1398, N1396, N459, N347);
nand NAND2 (N1399, N1391, N1339);
and AND4 (N1400, N1383, N159, N204, N1101);
or OR2 (N1401, N1375, N721);
not NOT1 (N1402, N1394);
xor XOR2 (N1403, N1397, N751);
xor XOR2 (N1404, N1403, N304);
buf BUF1 (N1405, N1402);
buf BUF1 (N1406, N1401);
buf BUF1 (N1407, N1399);
xor XOR2 (N1408, N1372, N1225);
and AND3 (N1409, N1386, N1310, N1405);
buf BUF1 (N1410, N395);
or OR2 (N1411, N1407, N708);
or OR3 (N1412, N1409, N1003, N543);
and AND4 (N1413, N1411, N788, N993, N784);
buf BUF1 (N1414, N1398);
nand NAND2 (N1415, N1404, N194);
buf BUF1 (N1416, N1413);
not NOT1 (N1417, N1412);
nor NOR2 (N1418, N1415, N415);
not NOT1 (N1419, N1400);
nand NAND2 (N1420, N1418, N424);
xor XOR2 (N1421, N1408, N49);
nor NOR4 (N1422, N1420, N890, N803, N413);
xor XOR2 (N1423, N1414, N1107);
and AND3 (N1424, N1410, N485, N1002);
not NOT1 (N1425, N1424);
nor NOR4 (N1426, N1422, N1317, N778, N167);
or OR3 (N1427, N1353, N1087, N368);
xor XOR2 (N1428, N1417, N1080);
and AND4 (N1429, N1425, N1140, N259, N875);
or OR2 (N1430, N1416, N400);
nand NAND2 (N1431, N1406, N1061);
or OR3 (N1432, N1428, N1209, N989);
nand NAND3 (N1433, N1419, N1154, N795);
nand NAND3 (N1434, N1431, N1408, N464);
buf BUF1 (N1435, N1432);
buf BUF1 (N1436, N1427);
xor XOR2 (N1437, N1426, N345);
and AND2 (N1438, N1434, N912);
buf BUF1 (N1439, N1429);
nand NAND4 (N1440, N1437, N320, N824, N165);
not NOT1 (N1441, N1436);
not NOT1 (N1442, N1421);
or OR2 (N1443, N1435, N223);
not NOT1 (N1444, N1442);
buf BUF1 (N1445, N1443);
nand NAND3 (N1446, N1393, N1055, N1316);
nand NAND4 (N1447, N1446, N488, N673, N475);
buf BUF1 (N1448, N1447);
nand NAND2 (N1449, N1438, N700);
xor XOR2 (N1450, N1430, N1416);
and AND3 (N1451, N1423, N971, N356);
nand NAND4 (N1452, N1445, N686, N41, N1280);
or OR3 (N1453, N1439, N238, N1106);
buf BUF1 (N1454, N1453);
nand NAND4 (N1455, N1448, N1264, N135, N872);
or OR4 (N1456, N1452, N1275, N1326, N783);
xor XOR2 (N1457, N1441, N163);
nand NAND4 (N1458, N1454, N232, N566, N1421);
not NOT1 (N1459, N1455);
buf BUF1 (N1460, N1444);
and AND4 (N1461, N1460, N1008, N644, N685);
buf BUF1 (N1462, N1459);
nor NOR4 (N1463, N1451, N1410, N961, N975);
buf BUF1 (N1464, N1450);
buf BUF1 (N1465, N1464);
buf BUF1 (N1466, N1457);
not NOT1 (N1467, N1458);
not NOT1 (N1468, N1449);
and AND2 (N1469, N1466, N1190);
nor NOR2 (N1470, N1440, N1159);
buf BUF1 (N1471, N1456);
nor NOR4 (N1472, N1471, N1364, N630, N803);
not NOT1 (N1473, N1469);
not NOT1 (N1474, N1472);
nand NAND3 (N1475, N1470, N852, N1357);
and AND2 (N1476, N1461, N1418);
buf BUF1 (N1477, N1433);
or OR3 (N1478, N1462, N182, N1400);
nand NAND4 (N1479, N1476, N1243, N411, N605);
and AND3 (N1480, N1467, N1164, N358);
or OR2 (N1481, N1475, N543);
and AND2 (N1482, N1468, N7);
nand NAND4 (N1483, N1479, N512, N175, N1398);
and AND4 (N1484, N1480, N1043, N27, N878);
nor NOR3 (N1485, N1477, N242, N252);
xor XOR2 (N1486, N1482, N450);
or OR4 (N1487, N1473, N1443, N609, N761);
or OR4 (N1488, N1484, N1222, N201, N1050);
not NOT1 (N1489, N1485);
and AND2 (N1490, N1488, N853);
and AND3 (N1491, N1465, N1115, N455);
not NOT1 (N1492, N1487);
xor XOR2 (N1493, N1492, N310);
not NOT1 (N1494, N1474);
xor XOR2 (N1495, N1481, N963);
xor XOR2 (N1496, N1495, N955);
not NOT1 (N1497, N1478);
buf BUF1 (N1498, N1497);
nor NOR2 (N1499, N1489, N178);
nor NOR3 (N1500, N1483, N778, N99);
nor NOR4 (N1501, N1500, N632, N969, N413);
nand NAND2 (N1502, N1498, N1436);
xor XOR2 (N1503, N1496, N550);
or OR3 (N1504, N1501, N782, N288);
nor NOR4 (N1505, N1463, N62, N509, N518);
nand NAND2 (N1506, N1491, N89);
buf BUF1 (N1507, N1486);
not NOT1 (N1508, N1504);
not NOT1 (N1509, N1490);
or OR2 (N1510, N1506, N1337);
and AND3 (N1511, N1502, N802, N956);
not NOT1 (N1512, N1494);
nor NOR4 (N1513, N1505, N1279, N1359, N1026);
not NOT1 (N1514, N1509);
nand NAND4 (N1515, N1513, N1023, N541, N1393);
buf BUF1 (N1516, N1508);
xor XOR2 (N1517, N1511, N260);
not NOT1 (N1518, N1512);
nor NOR2 (N1519, N1510, N1066);
and AND3 (N1520, N1493, N1223, N1186);
buf BUF1 (N1521, N1518);
buf BUF1 (N1522, N1514);
xor XOR2 (N1523, N1520, N992);
xor XOR2 (N1524, N1523, N201);
buf BUF1 (N1525, N1515);
nor NOR3 (N1526, N1517, N621, N1491);
nor NOR3 (N1527, N1525, N883, N191);
xor XOR2 (N1528, N1519, N412);
xor XOR2 (N1529, N1528, N393);
or OR4 (N1530, N1516, N844, N500, N969);
and AND3 (N1531, N1499, N510, N932);
nand NAND4 (N1532, N1524, N514, N992, N1299);
or OR3 (N1533, N1522, N1338, N452);
not NOT1 (N1534, N1521);
buf BUF1 (N1535, N1533);
not NOT1 (N1536, N1527);
and AND2 (N1537, N1507, N1119);
buf BUF1 (N1538, N1534);
nand NAND4 (N1539, N1535, N546, N979, N1038);
and AND4 (N1540, N1532, N439, N1024, N732);
not NOT1 (N1541, N1536);
not NOT1 (N1542, N1526);
not NOT1 (N1543, N1537);
xor XOR2 (N1544, N1539, N228);
nor NOR3 (N1545, N1540, N148, N204);
xor XOR2 (N1546, N1541, N1533);
nor NOR3 (N1547, N1546, N1138, N29);
or OR3 (N1548, N1544, N356, N217);
xor XOR2 (N1549, N1503, N182);
not NOT1 (N1550, N1531);
or OR3 (N1551, N1538, N752, N844);
not NOT1 (N1552, N1547);
buf BUF1 (N1553, N1530);
or OR3 (N1554, N1550, N1033, N889);
or OR2 (N1555, N1551, N1482);
xor XOR2 (N1556, N1548, N892);
buf BUF1 (N1557, N1545);
or OR2 (N1558, N1556, N1524);
nand NAND3 (N1559, N1555, N836, N973);
and AND2 (N1560, N1549, N136);
or OR4 (N1561, N1553, N802, N1424, N1004);
nor NOR2 (N1562, N1552, N242);
nand NAND4 (N1563, N1557, N509, N1453, N1209);
nor NOR3 (N1564, N1558, N61, N908);
or OR3 (N1565, N1560, N167, N1445);
or OR2 (N1566, N1565, N146);
buf BUF1 (N1567, N1563);
nor NOR3 (N1568, N1543, N364, N848);
and AND3 (N1569, N1562, N365, N1154);
and AND3 (N1570, N1567, N978, N1283);
or OR3 (N1571, N1564, N891, N246);
nor NOR4 (N1572, N1542, N1142, N157, N1072);
buf BUF1 (N1573, N1568);
nor NOR2 (N1574, N1559, N799);
nor NOR2 (N1575, N1574, N245);
and AND4 (N1576, N1554, N266, N1223, N570);
not NOT1 (N1577, N1566);
and AND2 (N1578, N1575, N20);
nor NOR4 (N1579, N1576, N352, N1461, N1105);
nor NOR3 (N1580, N1571, N1135, N200);
nor NOR2 (N1581, N1573, N1164);
nor NOR2 (N1582, N1579, N1468);
and AND4 (N1583, N1580, N721, N334, N112);
or OR4 (N1584, N1561, N1299, N556, N1002);
or OR2 (N1585, N1529, N998);
and AND2 (N1586, N1583, N514);
or OR4 (N1587, N1586, N1420, N1338, N1486);
and AND3 (N1588, N1569, N495, N269);
and AND3 (N1589, N1582, N361, N790);
and AND4 (N1590, N1572, N138, N1562, N1355);
xor XOR2 (N1591, N1570, N681);
nand NAND2 (N1592, N1584, N1362);
not NOT1 (N1593, N1590);
xor XOR2 (N1594, N1592, N426);
or OR3 (N1595, N1594, N25, N1233);
not NOT1 (N1596, N1591);
not NOT1 (N1597, N1589);
buf BUF1 (N1598, N1593);
xor XOR2 (N1599, N1581, N1561);
xor XOR2 (N1600, N1596, N1106);
or OR3 (N1601, N1597, N1567, N73);
buf BUF1 (N1602, N1587);
and AND2 (N1603, N1577, N1547);
or OR3 (N1604, N1578, N870, N147);
buf BUF1 (N1605, N1600);
xor XOR2 (N1606, N1605, N1421);
or OR3 (N1607, N1585, N197, N1303);
nor NOR3 (N1608, N1602, N909, N201);
xor XOR2 (N1609, N1599, N1013);
nand NAND3 (N1610, N1588, N125, N1100);
or OR4 (N1611, N1610, N1342, N875, N816);
and AND2 (N1612, N1601, N1161);
and AND3 (N1613, N1604, N265, N266);
buf BUF1 (N1614, N1611);
or OR4 (N1615, N1612, N1249, N1346, N400);
and AND3 (N1616, N1595, N252, N898);
nand NAND2 (N1617, N1614, N1454);
or OR4 (N1618, N1609, N1597, N867, N262);
nand NAND2 (N1619, N1608, N1401);
nand NAND2 (N1620, N1607, N185);
nand NAND4 (N1621, N1617, N1558, N255, N1556);
or OR4 (N1622, N1598, N1576, N1365, N1232);
nand NAND4 (N1623, N1619, N362, N573, N1033);
nor NOR3 (N1624, N1615, N1313, N763);
xor XOR2 (N1625, N1613, N979);
xor XOR2 (N1626, N1620, N134);
nand NAND3 (N1627, N1621, N436, N41);
xor XOR2 (N1628, N1618, N868);
and AND3 (N1629, N1627, N335, N263);
or OR2 (N1630, N1606, N666);
not NOT1 (N1631, N1623);
nand NAND3 (N1632, N1631, N769, N466);
buf BUF1 (N1633, N1616);
xor XOR2 (N1634, N1628, N615);
buf BUF1 (N1635, N1622);
nand NAND3 (N1636, N1632, N540, N734);
nand NAND3 (N1637, N1635, N1163, N24);
nor NOR4 (N1638, N1624, N40, N1585, N693);
buf BUF1 (N1639, N1634);
nor NOR3 (N1640, N1629, N1096, N1250);
nand NAND4 (N1641, N1640, N1507, N610, N1482);
nand NAND4 (N1642, N1638, N7, N613, N689);
not NOT1 (N1643, N1625);
nor NOR4 (N1644, N1642, N106, N464, N537);
nor NOR2 (N1645, N1626, N1246);
nor NOR3 (N1646, N1639, N1185, N1100);
and AND3 (N1647, N1630, N1037, N800);
nor NOR2 (N1648, N1603, N963);
buf BUF1 (N1649, N1641);
xor XOR2 (N1650, N1648, N830);
xor XOR2 (N1651, N1637, N1461);
not NOT1 (N1652, N1643);
nand NAND3 (N1653, N1651, N1375, N791);
or OR3 (N1654, N1646, N897, N1327);
buf BUF1 (N1655, N1636);
or OR4 (N1656, N1649, N941, N49, N688);
buf BUF1 (N1657, N1633);
xor XOR2 (N1658, N1654, N1321);
and AND2 (N1659, N1650, N336);
nor NOR2 (N1660, N1656, N1405);
nand NAND4 (N1661, N1657, N215, N629, N850);
buf BUF1 (N1662, N1645);
buf BUF1 (N1663, N1660);
nor NOR3 (N1664, N1658, N946, N1372);
nand NAND3 (N1665, N1647, N650, N742);
not NOT1 (N1666, N1665);
or OR3 (N1667, N1644, N606, N692);
not NOT1 (N1668, N1664);
nor NOR4 (N1669, N1668, N1609, N1619, N1313);
and AND3 (N1670, N1655, N558, N710);
xor XOR2 (N1671, N1669, N61);
nor NOR3 (N1672, N1662, N275, N1216);
xor XOR2 (N1673, N1671, N1077);
nand NAND4 (N1674, N1652, N55, N33, N718);
buf BUF1 (N1675, N1667);
nor NOR2 (N1676, N1670, N1618);
xor XOR2 (N1677, N1663, N708);
or OR2 (N1678, N1659, N901);
or OR2 (N1679, N1672, N595);
not NOT1 (N1680, N1666);
and AND3 (N1681, N1653, N139, N476);
or OR4 (N1682, N1677, N1383, N948, N1604);
buf BUF1 (N1683, N1681);
or OR2 (N1684, N1682, N495);
buf BUF1 (N1685, N1679);
buf BUF1 (N1686, N1674);
buf BUF1 (N1687, N1673);
or OR4 (N1688, N1678, N354, N1512, N654);
and AND4 (N1689, N1684, N1003, N191, N682);
nor NOR2 (N1690, N1688, N1032);
nand NAND2 (N1691, N1689, N1061);
xor XOR2 (N1692, N1676, N572);
buf BUF1 (N1693, N1686);
nor NOR3 (N1694, N1675, N560, N1351);
or OR4 (N1695, N1687, N797, N1461, N427);
xor XOR2 (N1696, N1694, N1645);
not NOT1 (N1697, N1661);
buf BUF1 (N1698, N1685);
xor XOR2 (N1699, N1696, N445);
buf BUF1 (N1700, N1692);
and AND3 (N1701, N1695, N1630, N1359);
xor XOR2 (N1702, N1693, N360);
buf BUF1 (N1703, N1697);
xor XOR2 (N1704, N1699, N170);
and AND2 (N1705, N1690, N661);
nand NAND2 (N1706, N1698, N1670);
buf BUF1 (N1707, N1703);
xor XOR2 (N1708, N1701, N1509);
and AND4 (N1709, N1708, N1335, N1475, N928);
and AND2 (N1710, N1706, N280);
not NOT1 (N1711, N1710);
and AND2 (N1712, N1683, N1082);
and AND3 (N1713, N1705, N573, N1254);
and AND3 (N1714, N1704, N1490, N676);
nor NOR2 (N1715, N1714, N861);
nor NOR3 (N1716, N1680, N869, N1191);
buf BUF1 (N1717, N1712);
nor NOR4 (N1718, N1707, N915, N985, N1161);
not NOT1 (N1719, N1717);
not NOT1 (N1720, N1711);
not NOT1 (N1721, N1691);
or OR3 (N1722, N1716, N794, N1026);
or OR4 (N1723, N1719, N281, N596, N368);
or OR3 (N1724, N1721, N290, N475);
not NOT1 (N1725, N1713);
or OR2 (N1726, N1715, N673);
and AND2 (N1727, N1724, N1014);
nand NAND2 (N1728, N1720, N909);
buf BUF1 (N1729, N1718);
or OR4 (N1730, N1722, N60, N575, N1209);
or OR3 (N1731, N1709, N422, N329);
or OR2 (N1732, N1702, N1313);
nor NOR3 (N1733, N1730, N1087, N1464);
buf BUF1 (N1734, N1733);
and AND2 (N1735, N1728, N74);
or OR2 (N1736, N1700, N128);
xor XOR2 (N1737, N1727, N1642);
nand NAND2 (N1738, N1723, N923);
xor XOR2 (N1739, N1729, N1305);
nand NAND4 (N1740, N1735, N962, N1328, N555);
not NOT1 (N1741, N1740);
nor NOR4 (N1742, N1732, N392, N504, N108);
nor NOR2 (N1743, N1741, N820);
nand NAND2 (N1744, N1742, N439);
not NOT1 (N1745, N1743);
not NOT1 (N1746, N1739);
not NOT1 (N1747, N1731);
xor XOR2 (N1748, N1734, N1602);
not NOT1 (N1749, N1726);
buf BUF1 (N1750, N1736);
nor NOR2 (N1751, N1750, N928);
not NOT1 (N1752, N1737);
not NOT1 (N1753, N1749);
and AND3 (N1754, N1753, N545, N1313);
and AND4 (N1755, N1745, N903, N1591, N1162);
not NOT1 (N1756, N1746);
not NOT1 (N1757, N1744);
nand NAND3 (N1758, N1755, N289, N939);
and AND2 (N1759, N1756, N881);
nor NOR3 (N1760, N1758, N770, N1264);
not NOT1 (N1761, N1760);
buf BUF1 (N1762, N1752);
not NOT1 (N1763, N1757);
buf BUF1 (N1764, N1761);
and AND3 (N1765, N1762, N44, N92);
or OR4 (N1766, N1759, N1569, N423, N1514);
nor NOR4 (N1767, N1748, N1729, N1442, N757);
nor NOR4 (N1768, N1751, N315, N1747, N1299);
buf BUF1 (N1769, N1234);
nand NAND2 (N1770, N1765, N304);
buf BUF1 (N1771, N1725);
buf BUF1 (N1772, N1771);
or OR4 (N1773, N1763, N1230, N936, N708);
xor XOR2 (N1774, N1768, N989);
not NOT1 (N1775, N1764);
nand NAND3 (N1776, N1770, N1456, N487);
or OR4 (N1777, N1775, N804, N861, N474);
not NOT1 (N1778, N1769);
and AND3 (N1779, N1766, N1120, N1255);
not NOT1 (N1780, N1738);
or OR2 (N1781, N1773, N6);
buf BUF1 (N1782, N1777);
and AND3 (N1783, N1781, N272, N813);
xor XOR2 (N1784, N1782, N418);
not NOT1 (N1785, N1780);
xor XOR2 (N1786, N1785, N364);
and AND4 (N1787, N1786, N129, N946, N388);
nand NAND4 (N1788, N1772, N1663, N1372, N1264);
or OR4 (N1789, N1754, N693, N1516, N1744);
and AND3 (N1790, N1788, N715, N1096);
nor NOR2 (N1791, N1790, N1174);
buf BUF1 (N1792, N1776);
not NOT1 (N1793, N1784);
buf BUF1 (N1794, N1778);
and AND3 (N1795, N1792, N1668, N490);
or OR2 (N1796, N1794, N526);
or OR3 (N1797, N1791, N1499, N1460);
or OR3 (N1798, N1797, N1409, N1094);
nor NOR4 (N1799, N1793, N1344, N1056, N1249);
and AND3 (N1800, N1796, N1753, N310);
xor XOR2 (N1801, N1795, N1436);
and AND4 (N1802, N1779, N153, N339, N1029);
nand NAND2 (N1803, N1798, N1340);
nand NAND3 (N1804, N1799, N1422, N260);
or OR2 (N1805, N1804, N1438);
not NOT1 (N1806, N1767);
buf BUF1 (N1807, N1774);
or OR4 (N1808, N1803, N995, N1181, N316);
not NOT1 (N1809, N1807);
and AND3 (N1810, N1809, N1472, N1447);
or OR3 (N1811, N1801, N850, N970);
and AND2 (N1812, N1805, N967);
nor NOR3 (N1813, N1812, N34, N138);
or OR2 (N1814, N1806, N682);
not NOT1 (N1815, N1813);
not NOT1 (N1816, N1814);
buf BUF1 (N1817, N1811);
nand NAND2 (N1818, N1817, N667);
buf BUF1 (N1819, N1808);
xor XOR2 (N1820, N1818, N843);
buf BUF1 (N1821, N1800);
or OR2 (N1822, N1787, N533);
xor XOR2 (N1823, N1789, N1243);
not NOT1 (N1824, N1820);
nor NOR2 (N1825, N1822, N608);
xor XOR2 (N1826, N1802, N723);
buf BUF1 (N1827, N1824);
or OR2 (N1828, N1823, N1247);
buf BUF1 (N1829, N1783);
xor XOR2 (N1830, N1819, N1811);
xor XOR2 (N1831, N1830, N1085);
or OR4 (N1832, N1815, N1040, N1189, N817);
xor XOR2 (N1833, N1832, N1554);
xor XOR2 (N1834, N1816, N1832);
nor NOR4 (N1835, N1825, N1716, N415, N550);
nand NAND3 (N1836, N1833, N1288, N1185);
nor NOR4 (N1837, N1834, N1703, N220, N1209);
not NOT1 (N1838, N1837);
or OR2 (N1839, N1829, N308);
or OR4 (N1840, N1839, N1588, N208, N129);
nand NAND4 (N1841, N1838, N655, N964, N1617);
not NOT1 (N1842, N1835);
nor NOR2 (N1843, N1826, N641);
xor XOR2 (N1844, N1841, N1707);
xor XOR2 (N1845, N1840, N769);
and AND3 (N1846, N1821, N336, N85);
or OR2 (N1847, N1828, N495);
buf BUF1 (N1848, N1844);
buf BUF1 (N1849, N1846);
or OR2 (N1850, N1843, N368);
nor NOR2 (N1851, N1831, N204);
or OR2 (N1852, N1836, N1305);
and AND3 (N1853, N1810, N1323, N163);
nor NOR3 (N1854, N1845, N1230, N341);
not NOT1 (N1855, N1852);
or OR4 (N1856, N1854, N1575, N588, N869);
not NOT1 (N1857, N1856);
not NOT1 (N1858, N1853);
buf BUF1 (N1859, N1842);
nor NOR3 (N1860, N1827, N1384, N583);
nand NAND3 (N1861, N1848, N1500, N1003);
or OR2 (N1862, N1860, N1369);
or OR4 (N1863, N1858, N884, N335, N115);
nor NOR3 (N1864, N1851, N162, N1522);
nor NOR3 (N1865, N1859, N1236, N1836);
nand NAND3 (N1866, N1865, N1082, N887);
not NOT1 (N1867, N1849);
and AND2 (N1868, N1864, N339);
nor NOR3 (N1869, N1857, N774, N590);
or OR4 (N1870, N1868, N1114, N3, N1102);
or OR4 (N1871, N1850, N718, N1837, N762);
not NOT1 (N1872, N1867);
or OR4 (N1873, N1869, N1534, N465, N1602);
xor XOR2 (N1874, N1870, N396);
not NOT1 (N1875, N1863);
nand NAND2 (N1876, N1871, N953);
nor NOR3 (N1877, N1861, N456, N1449);
not NOT1 (N1878, N1876);
or OR2 (N1879, N1873, N677);
buf BUF1 (N1880, N1872);
nand NAND2 (N1881, N1847, N1858);
nand NAND3 (N1882, N1874, N1368, N1687);
buf BUF1 (N1883, N1879);
nand NAND2 (N1884, N1882, N1451);
and AND3 (N1885, N1875, N812, N1728);
buf BUF1 (N1886, N1880);
nor NOR2 (N1887, N1877, N14);
not NOT1 (N1888, N1862);
nor NOR4 (N1889, N1887, N1407, N346, N1128);
nand NAND3 (N1890, N1866, N1699, N1278);
and AND4 (N1891, N1855, N376, N941, N865);
or OR2 (N1892, N1886, N1396);
xor XOR2 (N1893, N1885, N880);
buf BUF1 (N1894, N1893);
or OR3 (N1895, N1881, N383, N1226);
nand NAND4 (N1896, N1891, N1621, N754, N967);
or OR4 (N1897, N1878, N1832, N1561, N1652);
buf BUF1 (N1898, N1897);
buf BUF1 (N1899, N1898);
or OR3 (N1900, N1895, N617, N1744);
nor NOR4 (N1901, N1888, N181, N1006, N1243);
not NOT1 (N1902, N1896);
xor XOR2 (N1903, N1884, N1364);
xor XOR2 (N1904, N1900, N1791);
nand NAND4 (N1905, N1904, N720, N1470, N442);
and AND4 (N1906, N1883, N8, N1685, N622);
nand NAND2 (N1907, N1902, N72);
or OR3 (N1908, N1890, N465, N924);
nand NAND3 (N1909, N1905, N1738, N530);
not NOT1 (N1910, N1909);
nand NAND4 (N1911, N1908, N1693, N1497, N1553);
nor NOR3 (N1912, N1894, N737, N1063);
nand NAND2 (N1913, N1892, N1390);
nand NAND4 (N1914, N1911, N1226, N566, N239);
nor NOR3 (N1915, N1910, N1776, N1193);
and AND3 (N1916, N1889, N797, N1239);
nor NOR2 (N1917, N1903, N1665);
not NOT1 (N1918, N1906);
nand NAND2 (N1919, N1918, N87);
or OR3 (N1920, N1915, N1663, N218);
or OR3 (N1921, N1913, N897, N1561);
buf BUF1 (N1922, N1899);
and AND4 (N1923, N1916, N506, N353, N1349);
nand NAND4 (N1924, N1907, N942, N507, N354);
nand NAND4 (N1925, N1901, N827, N1457, N1548);
nor NOR2 (N1926, N1921, N125);
not NOT1 (N1927, N1922);
or OR4 (N1928, N1925, N834, N566, N1058);
nor NOR2 (N1929, N1923, N1049);
not NOT1 (N1930, N1926);
not NOT1 (N1931, N1924);
buf BUF1 (N1932, N1929);
or OR4 (N1933, N1919, N1029, N138, N276);
buf BUF1 (N1934, N1917);
buf BUF1 (N1935, N1933);
or OR3 (N1936, N1928, N1690, N1921);
and AND4 (N1937, N1931, N60, N1067, N875);
not NOT1 (N1938, N1920);
or OR2 (N1939, N1936, N1446);
not NOT1 (N1940, N1930);
not NOT1 (N1941, N1938);
nand NAND3 (N1942, N1934, N253, N518);
and AND4 (N1943, N1935, N1648, N601, N1551);
and AND4 (N1944, N1940, N976, N82, N1116);
not NOT1 (N1945, N1942);
xor XOR2 (N1946, N1944, N1192);
xor XOR2 (N1947, N1927, N1252);
and AND2 (N1948, N1943, N1021);
or OR4 (N1949, N1947, N84, N184, N217);
buf BUF1 (N1950, N1912);
not NOT1 (N1951, N1946);
or OR4 (N1952, N1914, N1526, N1202, N988);
nand NAND4 (N1953, N1951, N1552, N731, N186);
and AND4 (N1954, N1937, N1576, N1473, N1269);
nand NAND4 (N1955, N1952, N698, N163, N218);
not NOT1 (N1956, N1945);
buf BUF1 (N1957, N1954);
and AND4 (N1958, N1955, N1419, N175, N1519);
buf BUF1 (N1959, N1932);
xor XOR2 (N1960, N1939, N1537);
buf BUF1 (N1961, N1949);
or OR2 (N1962, N1960, N533);
and AND3 (N1963, N1950, N73, N326);
nor NOR4 (N1964, N1957, N1564, N1957, N422);
buf BUF1 (N1965, N1948);
xor XOR2 (N1966, N1963, N1447);
not NOT1 (N1967, N1941);
xor XOR2 (N1968, N1956, N430);
not NOT1 (N1969, N1962);
xor XOR2 (N1970, N1958, N353);
nand NAND4 (N1971, N1968, N954, N1711, N87);
buf BUF1 (N1972, N1965);
nand NAND3 (N1973, N1964, N1647, N1645);
nor NOR3 (N1974, N1973, N854, N1300);
nor NOR4 (N1975, N1959, N515, N1001, N1384);
or OR4 (N1976, N1971, N182, N461, N379);
buf BUF1 (N1977, N1975);
nor NOR3 (N1978, N1967, N1353, N797);
and AND2 (N1979, N1977, N1289);
nand NAND4 (N1980, N1961, N985, N1544, N529);
nand NAND3 (N1981, N1976, N782, N1083);
xor XOR2 (N1982, N1978, N808);
not NOT1 (N1983, N1980);
nor NOR4 (N1984, N1970, N61, N166, N1930);
xor XOR2 (N1985, N1972, N651);
not NOT1 (N1986, N1969);
not NOT1 (N1987, N1981);
buf BUF1 (N1988, N1987);
buf BUF1 (N1989, N1986);
and AND3 (N1990, N1953, N1890, N923);
buf BUF1 (N1991, N1989);
not NOT1 (N1992, N1979);
nor NOR3 (N1993, N1988, N1940, N1736);
nor NOR3 (N1994, N1992, N648, N377);
and AND3 (N1995, N1994, N1829, N683);
not NOT1 (N1996, N1966);
buf BUF1 (N1997, N1996);
nor NOR4 (N1998, N1990, N1671, N372, N1823);
xor XOR2 (N1999, N1985, N725);
buf BUF1 (N2000, N1998);
nor NOR2 (N2001, N1991, N1012);
nand NAND3 (N2002, N1984, N404, N98);
nor NOR4 (N2003, N1982, N1755, N879, N1140);
not NOT1 (N2004, N1993);
nor NOR3 (N2005, N2004, N532, N875);
xor XOR2 (N2006, N1997, N1435);
or OR2 (N2007, N2003, N565);
nand NAND3 (N2008, N2005, N363, N1800);
or OR4 (N2009, N2001, N1976, N1188, N229);
and AND2 (N2010, N2008, N198);
or OR3 (N2011, N1995, N853, N1530);
not NOT1 (N2012, N2002);
nand NAND4 (N2013, N2006, N1876, N855, N768);
or OR4 (N2014, N2010, N966, N1339, N1761);
xor XOR2 (N2015, N1999, N1487);
and AND3 (N2016, N2009, N1901, N1191);
nor NOR3 (N2017, N2011, N95, N312);
and AND4 (N2018, N2000, N949, N471, N2);
or OR3 (N2019, N2015, N32, N449);
or OR4 (N2020, N2014, N102, N1129, N1061);
xor XOR2 (N2021, N2012, N533);
not NOT1 (N2022, N2016);
buf BUF1 (N2023, N2022);
or OR4 (N2024, N2021, N805, N913, N807);
nand NAND4 (N2025, N2013, N1751, N1210, N1896);
and AND4 (N2026, N1983, N816, N644, N1627);
and AND4 (N2027, N2025, N344, N896, N691);
nand NAND4 (N2028, N2020, N1157, N47, N1994);
and AND2 (N2029, N2017, N673);
buf BUF1 (N2030, N2027);
and AND4 (N2031, N2023, N1527, N1815, N1627);
or OR4 (N2032, N2024, N1145, N1600, N623);
and AND3 (N2033, N2026, N1900, N601);
nor NOR4 (N2034, N2007, N568, N1849, N1765);
xor XOR2 (N2035, N2018, N1565);
and AND4 (N2036, N2028, N1666, N1010, N996);
and AND4 (N2037, N2036, N1888, N1700, N662);
nor NOR4 (N2038, N2019, N468, N520, N1134);
xor XOR2 (N2039, N2032, N1450);
not NOT1 (N2040, N2034);
nand NAND2 (N2041, N2030, N370);
buf BUF1 (N2042, N1974);
and AND4 (N2043, N2038, N200, N149, N1062);
not NOT1 (N2044, N2039);
or OR4 (N2045, N2044, N1521, N1411, N522);
nand NAND3 (N2046, N2043, N338, N572);
and AND2 (N2047, N2042, N1043);
not NOT1 (N2048, N2040);
buf BUF1 (N2049, N2029);
not NOT1 (N2050, N2046);
not NOT1 (N2051, N2035);
or OR2 (N2052, N2050, N225);
not NOT1 (N2053, N2031);
xor XOR2 (N2054, N2037, N1716);
nor NOR2 (N2055, N2054, N288);
not NOT1 (N2056, N2033);
not NOT1 (N2057, N2052);
xor XOR2 (N2058, N2048, N872);
nand NAND4 (N2059, N2058, N321, N654, N815);
or OR2 (N2060, N2055, N205);
nand NAND3 (N2061, N2051, N965, N1735);
nand NAND4 (N2062, N2049, N1445, N1477, N321);
xor XOR2 (N2063, N2045, N1626);
nor NOR2 (N2064, N2041, N1682);
buf BUF1 (N2065, N2060);
and AND4 (N2066, N2061, N570, N1744, N506);
and AND4 (N2067, N2062, N1328, N845, N1758);
nand NAND3 (N2068, N2056, N1078, N188);
and AND4 (N2069, N2059, N824, N1799, N856);
not NOT1 (N2070, N2067);
nor NOR2 (N2071, N2068, N788);
nor NOR3 (N2072, N2066, N275, N1533);
buf BUF1 (N2073, N2053);
not NOT1 (N2074, N2064);
nor NOR3 (N2075, N2072, N311, N2);
nor NOR3 (N2076, N2057, N868, N723);
nor NOR4 (N2077, N2047, N154, N13, N1511);
or OR3 (N2078, N2073, N1877, N1711);
nand NAND3 (N2079, N2077, N1661, N798);
nor NOR4 (N2080, N2074, N1137, N1230, N1366);
buf BUF1 (N2081, N2076);
and AND3 (N2082, N2081, N2073, N1973);
buf BUF1 (N2083, N2070);
nand NAND4 (N2084, N2079, N1229, N1695, N1976);
or OR2 (N2085, N2080, N640);
buf BUF1 (N2086, N2078);
not NOT1 (N2087, N2085);
and AND3 (N2088, N2071, N1108, N1829);
or OR2 (N2089, N2063, N1711);
nor NOR4 (N2090, N2088, N1278, N1662, N1901);
not NOT1 (N2091, N2084);
and AND3 (N2092, N2086, N1998, N747);
or OR2 (N2093, N2089, N1292);
nor NOR4 (N2094, N2069, N1452, N378, N1704);
or OR2 (N2095, N2090, N1157);
nor NOR2 (N2096, N2093, N1688);
or OR3 (N2097, N2094, N739, N1273);
nor NOR2 (N2098, N2092, N1633);
xor XOR2 (N2099, N2087, N1073);
nor NOR3 (N2100, N2082, N1997, N1331);
not NOT1 (N2101, N2096);
buf BUF1 (N2102, N2095);
nand NAND2 (N2103, N2098, N1419);
or OR3 (N2104, N2083, N644, N1721);
xor XOR2 (N2105, N2101, N1654);
not NOT1 (N2106, N2097);
not NOT1 (N2107, N2075);
xor XOR2 (N2108, N2102, N761);
nand NAND4 (N2109, N2091, N1011, N1095, N2049);
xor XOR2 (N2110, N2106, N1470);
buf BUF1 (N2111, N2108);
nor NOR2 (N2112, N2099, N118);
not NOT1 (N2113, N2104);
nor NOR4 (N2114, N2111, N370, N481, N782);
xor XOR2 (N2115, N2105, N1239);
and AND4 (N2116, N2100, N685, N1376, N1332);
nor NOR2 (N2117, N2103, N1432);
and AND4 (N2118, N2112, N146, N1643, N829);
and AND3 (N2119, N2114, N207, N1887);
nand NAND2 (N2120, N2109, N749);
nand NAND3 (N2121, N2117, N1866, N504);
not NOT1 (N2122, N2115);
nor NOR2 (N2123, N2122, N1208);
and AND2 (N2124, N2116, N686);
not NOT1 (N2125, N2121);
or OR2 (N2126, N2124, N1000);
nand NAND2 (N2127, N2123, N1267);
and AND2 (N2128, N2065, N1091);
xor XOR2 (N2129, N2126, N609);
buf BUF1 (N2130, N2119);
not NOT1 (N2131, N2129);
xor XOR2 (N2132, N2113, N1686);
not NOT1 (N2133, N2132);
or OR2 (N2134, N2118, N844);
xor XOR2 (N2135, N2120, N28);
and AND4 (N2136, N2131, N105, N249, N168);
nand NAND2 (N2137, N2125, N1783);
not NOT1 (N2138, N2107);
and AND3 (N2139, N2130, N332, N809);
xor XOR2 (N2140, N2110, N1197);
not NOT1 (N2141, N2136);
nor NOR3 (N2142, N2133, N635, N189);
nand NAND4 (N2143, N2135, N847, N855, N728);
and AND3 (N2144, N2143, N1967, N1103);
buf BUF1 (N2145, N2144);
xor XOR2 (N2146, N2137, N1418);
or OR4 (N2147, N2146, N1338, N801, N2044);
xor XOR2 (N2148, N2142, N410);
buf BUF1 (N2149, N2147);
or OR3 (N2150, N2140, N1565, N1286);
not NOT1 (N2151, N2141);
not NOT1 (N2152, N2149);
xor XOR2 (N2153, N2127, N1215);
and AND2 (N2154, N2134, N324);
xor XOR2 (N2155, N2148, N813);
xor XOR2 (N2156, N2150, N845);
not NOT1 (N2157, N2152);
buf BUF1 (N2158, N2139);
nand NAND3 (N2159, N2158, N443, N233);
and AND4 (N2160, N2153, N800, N244, N128);
not NOT1 (N2161, N2157);
or OR4 (N2162, N2161, N688, N1912, N1205);
not NOT1 (N2163, N2155);
not NOT1 (N2164, N2159);
nor NOR3 (N2165, N2151, N603, N36);
nand NAND4 (N2166, N2164, N732, N280, N1225);
nand NAND4 (N2167, N2128, N255, N1249, N1709);
and AND2 (N2168, N2167, N725);
or OR2 (N2169, N2162, N867);
nand NAND2 (N2170, N2138, N1671);
nand NAND3 (N2171, N2156, N224, N2164);
nand NAND3 (N2172, N2163, N349, N68);
nand NAND3 (N2173, N2172, N533, N1578);
buf BUF1 (N2174, N2168);
and AND2 (N2175, N2160, N1582);
not NOT1 (N2176, N2165);
buf BUF1 (N2177, N2169);
or OR4 (N2178, N2176, N373, N1090, N1091);
or OR3 (N2179, N2178, N627, N1178);
and AND4 (N2180, N2175, N256, N537, N640);
nand NAND4 (N2181, N2154, N1823, N59, N1454);
or OR4 (N2182, N2177, N862, N36, N725);
buf BUF1 (N2183, N2145);
xor XOR2 (N2184, N2170, N1298);
nor NOR4 (N2185, N2183, N1128, N1177, N1670);
and AND2 (N2186, N2184, N301);
xor XOR2 (N2187, N2171, N355);
xor XOR2 (N2188, N2187, N1056);
nor NOR4 (N2189, N2173, N1978, N2043, N1028);
nand NAND4 (N2190, N2181, N2034, N653, N125);
nor NOR2 (N2191, N2190, N1662);
buf BUF1 (N2192, N2174);
xor XOR2 (N2193, N2191, N1024);
nand NAND4 (N2194, N2192, N1928, N1739, N1214);
and AND2 (N2195, N2179, N2067);
nor NOR4 (N2196, N2182, N1295, N560, N1311);
buf BUF1 (N2197, N2196);
nor NOR2 (N2198, N2180, N1142);
or OR3 (N2199, N2194, N46, N1613);
nand NAND4 (N2200, N2198, N1191, N878, N1542);
not NOT1 (N2201, N2197);
nor NOR3 (N2202, N2188, N789, N1731);
and AND2 (N2203, N2202, N336);
nand NAND3 (N2204, N2201, N1214, N926);
buf BUF1 (N2205, N2203);
nor NOR4 (N2206, N2193, N1128, N1529, N2167);
xor XOR2 (N2207, N2189, N2018);
not NOT1 (N2208, N2205);
buf BUF1 (N2209, N2199);
xor XOR2 (N2210, N2200, N1120);
or OR2 (N2211, N2206, N674);
nor NOR4 (N2212, N2211, N1988, N1806, N206);
buf BUF1 (N2213, N2186);
buf BUF1 (N2214, N2212);
buf BUF1 (N2215, N2209);
and AND2 (N2216, N2214, N1504);
nor NOR2 (N2217, N2213, N1117);
xor XOR2 (N2218, N2216, N1084);
and AND3 (N2219, N2208, N2199, N614);
not NOT1 (N2220, N2217);
nand NAND4 (N2221, N2210, N2127, N583, N422);
and AND2 (N2222, N2166, N560);
or OR4 (N2223, N2222, N1641, N1876, N1206);
nor NOR2 (N2224, N2215, N1256);
nand NAND3 (N2225, N2219, N1641, N1470);
and AND4 (N2226, N2223, N1286, N1620, N656);
and AND4 (N2227, N2221, N53, N25, N1271);
or OR4 (N2228, N2218, N110, N283, N1032);
xor XOR2 (N2229, N2228, N611);
buf BUF1 (N2230, N2227);
xor XOR2 (N2231, N2225, N1327);
buf BUF1 (N2232, N2185);
xor XOR2 (N2233, N2226, N1776);
nor NOR4 (N2234, N2207, N2208, N947, N38);
nor NOR3 (N2235, N2229, N1362, N953);
nand NAND3 (N2236, N2220, N1678, N1729);
nand NAND2 (N2237, N2235, N551);
not NOT1 (N2238, N2195);
and AND3 (N2239, N2237, N1135, N1172);
xor XOR2 (N2240, N2231, N2196);
nor NOR2 (N2241, N2233, N2015);
nand NAND2 (N2242, N2232, N1530);
xor XOR2 (N2243, N2224, N1384);
buf BUF1 (N2244, N2230);
buf BUF1 (N2245, N2242);
and AND4 (N2246, N2239, N1707, N1032, N1356);
and AND3 (N2247, N2204, N125, N2015);
nand NAND2 (N2248, N2244, N756);
and AND4 (N2249, N2236, N1381, N2095, N105);
or OR3 (N2250, N2234, N1043, N650);
or OR3 (N2251, N2243, N519, N300);
buf BUF1 (N2252, N2247);
buf BUF1 (N2253, N2246);
nor NOR4 (N2254, N2249, N1216, N2241, N445);
buf BUF1 (N2255, N1766);
nor NOR2 (N2256, N2248, N862);
xor XOR2 (N2257, N2250, N2038);
nor NOR3 (N2258, N2255, N965, N2045);
buf BUF1 (N2259, N2240);
nor NOR2 (N2260, N2256, N1008);
xor XOR2 (N2261, N2260, N609);
nand NAND2 (N2262, N2258, N1564);
xor XOR2 (N2263, N2262, N994);
xor XOR2 (N2264, N2263, N2241);
not NOT1 (N2265, N2252);
nor NOR4 (N2266, N2261, N473, N28, N1692);
nor NOR3 (N2267, N2264, N130, N1128);
buf BUF1 (N2268, N2253);
not NOT1 (N2269, N2254);
nor NOR4 (N2270, N2266, N586, N230, N1551);
buf BUF1 (N2271, N2238);
or OR3 (N2272, N2268, N2200, N689);
and AND3 (N2273, N2270, N1142, N929);
or OR2 (N2274, N2273, N1950);
xor XOR2 (N2275, N2265, N219);
xor XOR2 (N2276, N2269, N1884);
nand NAND2 (N2277, N2257, N1981);
and AND3 (N2278, N2275, N436, N1069);
and AND4 (N2279, N2267, N1521, N20, N805);
not NOT1 (N2280, N2259);
and AND4 (N2281, N2278, N998, N1220, N1716);
not NOT1 (N2282, N2277);
xor XOR2 (N2283, N2271, N493);
nand NAND4 (N2284, N2282, N1098, N589, N1726);
buf BUF1 (N2285, N2251);
nand NAND2 (N2286, N2279, N2191);
xor XOR2 (N2287, N2274, N1623);
and AND2 (N2288, N2245, N402);
nor NOR4 (N2289, N2287, N1133, N2126, N655);
nor NOR2 (N2290, N2288, N43);
buf BUF1 (N2291, N2281);
nand NAND4 (N2292, N2290, N1435, N311, N838);
or OR2 (N2293, N2283, N1175);
or OR4 (N2294, N2276, N1009, N809, N1251);
nor NOR2 (N2295, N2272, N1680);
not NOT1 (N2296, N2295);
xor XOR2 (N2297, N2286, N186);
nand NAND2 (N2298, N2285, N104);
not NOT1 (N2299, N2289);
or OR4 (N2300, N2284, N699, N1889, N1249);
nand NAND3 (N2301, N2280, N1891, N1211);
not NOT1 (N2302, N2301);
buf BUF1 (N2303, N2294);
xor XOR2 (N2304, N2298, N1888);
not NOT1 (N2305, N2291);
xor XOR2 (N2306, N2300, N1800);
xor XOR2 (N2307, N2297, N892);
buf BUF1 (N2308, N2305);
or OR2 (N2309, N2292, N2192);
buf BUF1 (N2310, N2302);
nand NAND2 (N2311, N2303, N2292);
nor NOR3 (N2312, N2311, N698, N1950);
not NOT1 (N2313, N2309);
not NOT1 (N2314, N2313);
buf BUF1 (N2315, N2304);
xor XOR2 (N2316, N2314, N408);
xor XOR2 (N2317, N2308, N1820);
nor NOR3 (N2318, N2312, N107, N2115);
or OR2 (N2319, N2306, N1526);
or OR4 (N2320, N2310, N1275, N678, N921);
nand NAND4 (N2321, N2318, N2278, N1606, N356);
or OR2 (N2322, N2316, N419);
nand NAND3 (N2323, N2320, N284, N83);
nor NOR4 (N2324, N2319, N422, N1765, N295);
buf BUF1 (N2325, N2323);
xor XOR2 (N2326, N2307, N1085);
nand NAND2 (N2327, N2293, N471);
buf BUF1 (N2328, N2325);
or OR2 (N2329, N2326, N1326);
not NOT1 (N2330, N2324);
or OR4 (N2331, N2296, N624, N1116, N51);
nand NAND3 (N2332, N2315, N1210, N102);
not NOT1 (N2333, N2331);
buf BUF1 (N2334, N2317);
nor NOR2 (N2335, N2329, N2188);
and AND3 (N2336, N2321, N839, N1373);
nand NAND3 (N2337, N2335, N465, N1072);
not NOT1 (N2338, N2330);
or OR4 (N2339, N2332, N2174, N866, N1276);
nor NOR4 (N2340, N2322, N1719, N462, N1620);
and AND3 (N2341, N2334, N1534, N25);
nor NOR3 (N2342, N2338, N1050, N1373);
or OR4 (N2343, N2340, N1649, N656, N1591);
buf BUF1 (N2344, N2327);
xor XOR2 (N2345, N2343, N985);
xor XOR2 (N2346, N2342, N164);
or OR2 (N2347, N2333, N837);
buf BUF1 (N2348, N2328);
nor NOR4 (N2349, N2344, N1549, N988, N1745);
nand NAND3 (N2350, N2341, N428, N2133);
nand NAND4 (N2351, N2348, N1660, N946, N1000);
buf BUF1 (N2352, N2349);
xor XOR2 (N2353, N2336, N2316);
xor XOR2 (N2354, N2347, N2334);
nand NAND2 (N2355, N2346, N1535);
xor XOR2 (N2356, N2354, N752);
nor NOR4 (N2357, N2299, N1389, N1218, N1229);
nand NAND3 (N2358, N2356, N1493, N323);
nor NOR3 (N2359, N2355, N1236, N2184);
buf BUF1 (N2360, N2357);
nand NAND3 (N2361, N2353, N2322, N2);
nor NOR3 (N2362, N2360, N1686, N2344);
and AND4 (N2363, N2337, N1265, N2007, N94);
nand NAND4 (N2364, N2362, N1657, N2092, N108);
nor NOR4 (N2365, N2339, N2361, N1358, N1888);
xor XOR2 (N2366, N2178, N283);
xor XOR2 (N2367, N2345, N1500);
or OR4 (N2368, N2358, N957, N1474, N2292);
nand NAND3 (N2369, N2365, N979, N1569);
or OR3 (N2370, N2366, N458, N1033);
and AND4 (N2371, N2370, N41, N1972, N635);
and AND3 (N2372, N2367, N1149, N740);
buf BUF1 (N2373, N2368);
not NOT1 (N2374, N2373);
nand NAND2 (N2375, N2350, N1183);
nand NAND4 (N2376, N2369, N256, N2268, N718);
buf BUF1 (N2377, N2351);
or OR3 (N2378, N2377, N507, N2081);
nand NAND4 (N2379, N2359, N360, N1742, N395);
and AND3 (N2380, N2376, N1099, N1670);
or OR4 (N2381, N2380, N1353, N838, N1248);
xor XOR2 (N2382, N2363, N522);
and AND4 (N2383, N2364, N1642, N2073, N2023);
and AND2 (N2384, N2379, N1989);
xor XOR2 (N2385, N2374, N2315);
or OR4 (N2386, N2371, N452, N2172, N595);
xor XOR2 (N2387, N2386, N1229);
nand NAND3 (N2388, N2372, N527, N796);
buf BUF1 (N2389, N2381);
nand NAND4 (N2390, N2385, N2016, N826, N1736);
or OR2 (N2391, N2382, N1210);
not NOT1 (N2392, N2389);
not NOT1 (N2393, N2352);
and AND4 (N2394, N2388, N573, N466, N1214);
nand NAND3 (N2395, N2394, N1017, N1514);
xor XOR2 (N2396, N2378, N1613);
nor NOR3 (N2397, N2387, N1964, N305);
and AND4 (N2398, N2375, N1026, N2126, N2208);
or OR3 (N2399, N2397, N1835, N1753);
nor NOR2 (N2400, N2399, N1388);
nor NOR3 (N2401, N2383, N52, N2354);
nand NAND4 (N2402, N2384, N1035, N1163, N2351);
nand NAND2 (N2403, N2392, N2122);
nand NAND2 (N2404, N2391, N2127);
and AND3 (N2405, N2402, N1416, N773);
nand NAND3 (N2406, N2396, N1433, N2152);
or OR2 (N2407, N2398, N1315);
xor XOR2 (N2408, N2403, N1976);
or OR2 (N2409, N2405, N842);
and AND3 (N2410, N2400, N355, N927);
not NOT1 (N2411, N2406);
nand NAND4 (N2412, N2410, N1834, N1872, N2262);
buf BUF1 (N2413, N2408);
or OR4 (N2414, N2411, N447, N1058, N2019);
nand NAND4 (N2415, N2390, N1934, N99, N552);
nor NOR3 (N2416, N2393, N778, N1907);
not NOT1 (N2417, N2404);
or OR4 (N2418, N2413, N422, N1062, N195);
buf BUF1 (N2419, N2407);
not NOT1 (N2420, N2401);
not NOT1 (N2421, N2416);
not NOT1 (N2422, N2415);
nand NAND3 (N2423, N2417, N277, N1112);
xor XOR2 (N2424, N2395, N172);
xor XOR2 (N2425, N2423, N1743);
or OR3 (N2426, N2412, N2031, N586);
nor NOR2 (N2427, N2424, N857);
buf BUF1 (N2428, N2414);
or OR4 (N2429, N2409, N1068, N1231, N1443);
nand NAND2 (N2430, N2418, N175);
and AND2 (N2431, N2428, N1182);
and AND4 (N2432, N2420, N19, N247, N279);
and AND4 (N2433, N2427, N1646, N971, N823);
not NOT1 (N2434, N2429);
or OR3 (N2435, N2421, N932, N781);
nand NAND4 (N2436, N2426, N1509, N2153, N740);
not NOT1 (N2437, N2430);
and AND2 (N2438, N2437, N948);
or OR2 (N2439, N2419, N424);
nor NOR2 (N2440, N2435, N48);
and AND3 (N2441, N2422, N511, N1659);
buf BUF1 (N2442, N2440);
nand NAND2 (N2443, N2425, N1615);
not NOT1 (N2444, N2441);
nand NAND4 (N2445, N2433, N537, N1543, N1087);
nand NAND4 (N2446, N2434, N1465, N231, N704);
nand NAND4 (N2447, N2442, N1294, N1194, N1763);
or OR3 (N2448, N2446, N534, N1110);
nor NOR2 (N2449, N2432, N1240);
and AND3 (N2450, N2444, N75, N1778);
buf BUF1 (N2451, N2449);
xor XOR2 (N2452, N2447, N1270);
nand NAND2 (N2453, N2450, N2147);
not NOT1 (N2454, N2439);
nor NOR3 (N2455, N2454, N1552, N2062);
and AND4 (N2456, N2431, N2303, N570, N96);
buf BUF1 (N2457, N2445);
xor XOR2 (N2458, N2455, N886);
and AND3 (N2459, N2443, N961, N498);
or OR4 (N2460, N2457, N229, N1881, N911);
not NOT1 (N2461, N2453);
nand NAND3 (N2462, N2459, N110, N1735);
not NOT1 (N2463, N2448);
nor NOR2 (N2464, N2451, N816);
not NOT1 (N2465, N2438);
xor XOR2 (N2466, N2463, N1806);
not NOT1 (N2467, N2436);
and AND3 (N2468, N2464, N2120, N563);
not NOT1 (N2469, N2460);
buf BUF1 (N2470, N2466);
not NOT1 (N2471, N2458);
nor NOR4 (N2472, N2470, N1217, N1487, N2048);
nor NOR4 (N2473, N2461, N1278, N2427, N589);
or OR4 (N2474, N2467, N38, N2181, N1420);
xor XOR2 (N2475, N2462, N1348);
or OR4 (N2476, N2469, N507, N336, N2318);
or OR2 (N2477, N2474, N82);
nor NOR2 (N2478, N2471, N2435);
and AND4 (N2479, N2452, N1642, N1506, N1806);
buf BUF1 (N2480, N2472);
nor NOR4 (N2481, N2465, N384, N2275, N2374);
buf BUF1 (N2482, N2479);
xor XOR2 (N2483, N2478, N931);
and AND3 (N2484, N2476, N686, N139);
xor XOR2 (N2485, N2482, N2332);
or OR2 (N2486, N2475, N2441);
not NOT1 (N2487, N2481);
or OR3 (N2488, N2487, N1210, N17);
xor XOR2 (N2489, N2456, N1910);
or OR2 (N2490, N2489, N58);
nand NAND4 (N2491, N2484, N848, N396, N870);
and AND4 (N2492, N2491, N306, N2343, N65);
xor XOR2 (N2493, N2490, N2017);
xor XOR2 (N2494, N2468, N1329);
nand NAND4 (N2495, N2480, N55, N403, N1558);
nor NOR4 (N2496, N2483, N1604, N1119, N488);
nand NAND3 (N2497, N2492, N1324, N1495);
and AND2 (N2498, N2473, N1634);
and AND3 (N2499, N2477, N1571, N1526);
nor NOR3 (N2500, N2485, N2303, N80);
and AND4 (N2501, N2494, N604, N1472, N229);
buf BUF1 (N2502, N2496);
nor NOR3 (N2503, N2495, N1623, N384);
and AND2 (N2504, N2499, N1882);
and AND2 (N2505, N2493, N1302);
nand NAND3 (N2506, N2497, N10, N366);
not NOT1 (N2507, N2500);
or OR3 (N2508, N2502, N1893, N1621);
or OR2 (N2509, N2488, N2220);
nand NAND3 (N2510, N2508, N698, N1296);
buf BUF1 (N2511, N2505);
nor NOR2 (N2512, N2510, N580);
buf BUF1 (N2513, N2504);
xor XOR2 (N2514, N2509, N1705);
buf BUF1 (N2515, N2512);
xor XOR2 (N2516, N2501, N103);
nor NOR4 (N2517, N2486, N222, N1494, N717);
and AND3 (N2518, N2511, N761, N1198);
xor XOR2 (N2519, N2507, N1355);
nor NOR3 (N2520, N2503, N1586, N2263);
endmodule