// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17;

output N811,N802,N800,N798,N812,N814,N816,N815,N810,N817;

nor NOR4 (N18, N17, N16, N12, N12);
or OR4 (N19, N12, N17, N6, N10);
buf BUF1 (N20, N14);
not NOT1 (N21, N16);
and AND3 (N22, N1, N13, N13);
nand NAND3 (N23, N19, N7, N11);
xor XOR2 (N24, N13, N17);
nor NOR4 (N25, N18, N20, N9, N6);
or OR2 (N26, N7, N2);
xor XOR2 (N27, N15, N25);
nand NAND2 (N28, N25, N10);
and AND2 (N29, N12, N2);
not NOT1 (N30, N24);
not NOT1 (N31, N2);
and AND3 (N32, N3, N23, N21);
nor NOR4 (N33, N29, N1, N25, N17);
and AND3 (N34, N1, N17, N18);
and AND4 (N35, N6, N27, N13, N4);
and AND2 (N36, N10, N30);
xor XOR2 (N37, N18, N13);
xor XOR2 (N38, N35, N9);
nand NAND4 (N39, N36, N6, N4, N7);
nor NOR3 (N40, N32, N1, N25);
not NOT1 (N41, N39);
and AND4 (N42, N37, N1, N3, N15);
nor NOR4 (N43, N28, N27, N19, N39);
xor XOR2 (N44, N43, N40);
nor NOR2 (N45, N6, N29);
xor XOR2 (N46, N41, N44);
xor XOR2 (N47, N13, N31);
nor NOR2 (N48, N14, N11);
nor NOR2 (N49, N48, N40);
xor XOR2 (N50, N22, N42);
or OR3 (N51, N5, N25, N46);
xor XOR2 (N52, N49, N49);
not NOT1 (N53, N7);
or OR3 (N54, N51, N37, N12);
buf BUF1 (N55, N53);
and AND2 (N56, N54, N21);
nand NAND3 (N57, N47, N35, N30);
nand NAND4 (N58, N33, N16, N10, N32);
buf BUF1 (N59, N38);
or OR4 (N60, N56, N30, N24, N4);
xor XOR2 (N61, N60, N26);
nand NAND4 (N62, N43, N14, N41, N39);
nand NAND4 (N63, N55, N31, N34, N13);
and AND4 (N64, N43, N58, N10, N59);
buf BUF1 (N65, N12);
or OR2 (N66, N40, N57);
buf BUF1 (N67, N41);
and AND4 (N68, N45, N9, N13, N47);
or OR4 (N69, N66, N48, N54, N33);
nand NAND4 (N70, N52, N18, N33, N8);
nand NAND2 (N71, N64, N11);
or OR2 (N72, N67, N8);
buf BUF1 (N73, N65);
nor NOR3 (N74, N68, N39, N29);
not NOT1 (N75, N72);
not NOT1 (N76, N71);
and AND4 (N77, N69, N23, N68, N54);
or OR3 (N78, N63, N54, N54);
not NOT1 (N79, N62);
nor NOR4 (N80, N76, N27, N9, N41);
buf BUF1 (N81, N79);
or OR3 (N82, N75, N50, N2);
and AND4 (N83, N17, N51, N63, N82);
buf BUF1 (N84, N34);
not NOT1 (N85, N83);
or OR4 (N86, N61, N4, N55, N26);
not NOT1 (N87, N81);
nor NOR4 (N88, N86, N79, N87, N64);
nor NOR4 (N89, N35, N16, N16, N6);
or OR3 (N90, N84, N89, N32);
nor NOR2 (N91, N10, N71);
nand NAND4 (N92, N70, N14, N23, N79);
and AND4 (N93, N74, N67, N19, N9);
nor NOR3 (N94, N85, N89, N36);
buf BUF1 (N95, N94);
not NOT1 (N96, N90);
buf BUF1 (N97, N77);
buf BUF1 (N98, N96);
and AND4 (N99, N97, N63, N42, N35);
not NOT1 (N100, N92);
nand NAND4 (N101, N93, N82, N13, N58);
buf BUF1 (N102, N80);
or OR3 (N103, N98, N23, N70);
xor XOR2 (N104, N91, N58);
nor NOR2 (N105, N78, N90);
not NOT1 (N106, N73);
nand NAND2 (N107, N99, N83);
and AND4 (N108, N104, N19, N2, N32);
xor XOR2 (N109, N103, N85);
nand NAND3 (N110, N107, N91, N93);
nor NOR4 (N111, N110, N42, N6, N11);
buf BUF1 (N112, N108);
xor XOR2 (N113, N112, N92);
xor XOR2 (N114, N113, N6);
nor NOR2 (N115, N101, N13);
nand NAND2 (N116, N111, N41);
not NOT1 (N117, N102);
nor NOR2 (N118, N115, N10);
xor XOR2 (N119, N114, N84);
not NOT1 (N120, N118);
nor NOR4 (N121, N88, N10, N46, N13);
or OR2 (N122, N121, N9);
or OR4 (N123, N105, N90, N5, N75);
nor NOR2 (N124, N95, N50);
buf BUF1 (N125, N119);
not NOT1 (N126, N123);
and AND3 (N127, N109, N96, N62);
and AND3 (N128, N124, N8, N8);
or OR2 (N129, N116, N69);
and AND4 (N130, N122, N72, N38, N76);
not NOT1 (N131, N126);
or OR3 (N132, N127, N97, N105);
nand NAND3 (N133, N128, N126, N58);
buf BUF1 (N134, N120);
not NOT1 (N135, N129);
nand NAND2 (N136, N117, N130);
or OR2 (N137, N126, N6);
not NOT1 (N138, N100);
nand NAND2 (N139, N125, N96);
not NOT1 (N140, N106);
nor NOR2 (N141, N133, N138);
or OR3 (N142, N117, N47, N107);
nor NOR4 (N143, N142, N54, N75, N122);
or OR4 (N144, N136, N107, N71, N72);
or OR4 (N145, N139, N25, N113, N16);
and AND2 (N146, N135, N86);
and AND4 (N147, N145, N30, N32, N87);
xor XOR2 (N148, N132, N106);
or OR2 (N149, N141, N142);
xor XOR2 (N150, N149, N129);
nand NAND4 (N151, N148, N18, N6, N81);
buf BUF1 (N152, N131);
and AND4 (N153, N137, N48, N13, N151);
xor XOR2 (N154, N128, N149);
not NOT1 (N155, N154);
nor NOR4 (N156, N140, N133, N118, N55);
not NOT1 (N157, N134);
xor XOR2 (N158, N143, N91);
xor XOR2 (N159, N150, N88);
xor XOR2 (N160, N158, N80);
not NOT1 (N161, N156);
xor XOR2 (N162, N161, N33);
not NOT1 (N163, N155);
xor XOR2 (N164, N160, N121);
nand NAND3 (N165, N162, N133, N116);
or OR2 (N166, N159, N139);
buf BUF1 (N167, N157);
nand NAND2 (N168, N163, N139);
xor XOR2 (N169, N144, N158);
nand NAND2 (N170, N167, N88);
xor XOR2 (N171, N168, N150);
and AND3 (N172, N169, N65, N154);
nor NOR2 (N173, N147, N24);
nor NOR2 (N174, N165, N171);
xor XOR2 (N175, N107, N60);
and AND4 (N176, N153, N171, N111, N16);
and AND4 (N177, N172, N64, N7, N132);
and AND3 (N178, N166, N139, N131);
nand NAND3 (N179, N146, N115, N40);
nor NOR3 (N180, N177, N82, N150);
xor XOR2 (N181, N170, N178);
not NOT1 (N182, N85);
nand NAND3 (N183, N164, N9, N155);
xor XOR2 (N184, N182, N127);
nor NOR4 (N185, N152, N115, N60, N183);
and AND3 (N186, N68, N43, N81);
nor NOR2 (N187, N173, N177);
not NOT1 (N188, N184);
buf BUF1 (N189, N175);
buf BUF1 (N190, N181);
not NOT1 (N191, N180);
or OR3 (N192, N187, N179, N135);
nand NAND3 (N193, N14, N88, N71);
and AND2 (N194, N189, N37);
or OR3 (N195, N194, N108, N78);
nor NOR4 (N196, N188, N62, N128, N139);
not NOT1 (N197, N186);
or OR2 (N198, N191, N99);
nor NOR3 (N199, N198, N63, N47);
or OR2 (N200, N192, N10);
xor XOR2 (N201, N196, N170);
nor NOR3 (N202, N174, N183, N11);
and AND2 (N203, N201, N122);
or OR3 (N204, N195, N102, N33);
and AND2 (N205, N197, N32);
or OR2 (N206, N205, N179);
buf BUF1 (N207, N185);
buf BUF1 (N208, N206);
xor XOR2 (N209, N199, N135);
nor NOR2 (N210, N207, N76);
buf BUF1 (N211, N200);
xor XOR2 (N212, N190, N185);
buf BUF1 (N213, N193);
buf BUF1 (N214, N212);
or OR4 (N215, N208, N25, N13, N187);
buf BUF1 (N216, N211);
or OR3 (N217, N209, N129, N136);
buf BUF1 (N218, N204);
or OR3 (N219, N202, N46, N175);
nand NAND4 (N220, N216, N124, N15, N88);
nand NAND4 (N221, N219, N75, N184, N219);
nor NOR4 (N222, N214, N99, N109, N194);
nor NOR2 (N223, N221, N141);
and AND3 (N224, N223, N124, N78);
not NOT1 (N225, N210);
xor XOR2 (N226, N217, N62);
nor NOR3 (N227, N218, N58, N225);
nand NAND3 (N228, N74, N199, N46);
nor NOR4 (N229, N203, N67, N1, N194);
nand NAND2 (N230, N222, N99);
nor NOR2 (N231, N228, N113);
nand NAND4 (N232, N231, N84, N219, N118);
xor XOR2 (N233, N224, N207);
xor XOR2 (N234, N229, N230);
nor NOR3 (N235, N76, N49, N107);
buf BUF1 (N236, N232);
buf BUF1 (N237, N213);
buf BUF1 (N238, N227);
buf BUF1 (N239, N220);
not NOT1 (N240, N239);
nor NOR2 (N241, N240, N93);
buf BUF1 (N242, N236);
nand NAND4 (N243, N234, N16, N149, N117);
and AND3 (N244, N242, N108, N47);
and AND3 (N245, N226, N7, N51);
and AND4 (N246, N237, N131, N129, N96);
buf BUF1 (N247, N244);
not NOT1 (N248, N247);
xor XOR2 (N249, N215, N164);
buf BUF1 (N250, N249);
nor NOR2 (N251, N246, N6);
xor XOR2 (N252, N233, N144);
and AND3 (N253, N235, N184, N2);
and AND3 (N254, N250, N71, N214);
xor XOR2 (N255, N238, N158);
or OR4 (N256, N245, N122, N159, N120);
or OR4 (N257, N254, N254, N46, N44);
nand NAND3 (N258, N176, N224, N143);
buf BUF1 (N259, N241);
nand NAND2 (N260, N253, N157);
nor NOR3 (N261, N257, N220, N102);
not NOT1 (N262, N260);
and AND3 (N263, N248, N72, N115);
or OR2 (N264, N243, N147);
buf BUF1 (N265, N261);
nor NOR2 (N266, N258, N23);
or OR3 (N267, N262, N74, N61);
or OR4 (N268, N252, N208, N179, N243);
nand NAND2 (N269, N256, N161);
and AND3 (N270, N255, N66, N188);
nor NOR4 (N271, N263, N14, N125, N24);
not NOT1 (N272, N259);
and AND4 (N273, N266, N147, N193, N170);
nand NAND4 (N274, N273, N32, N178, N203);
xor XOR2 (N275, N270, N212);
not NOT1 (N276, N272);
or OR3 (N277, N271, N97, N106);
nand NAND3 (N278, N268, N39, N265);
xor XOR2 (N279, N260, N242);
or OR2 (N280, N264, N228);
buf BUF1 (N281, N269);
nand NAND3 (N282, N279, N80, N118);
xor XOR2 (N283, N280, N196);
or OR4 (N284, N281, N189, N53, N197);
nand NAND2 (N285, N277, N45);
nor NOR4 (N286, N267, N140, N193, N178);
nor NOR3 (N287, N275, N161, N184);
buf BUF1 (N288, N274);
buf BUF1 (N289, N282);
and AND2 (N290, N289, N67);
not NOT1 (N291, N284);
xor XOR2 (N292, N286, N57);
nor NOR3 (N293, N292, N104, N94);
xor XOR2 (N294, N290, N189);
buf BUF1 (N295, N288);
and AND2 (N296, N251, N59);
nor NOR4 (N297, N283, N260, N173, N7);
not NOT1 (N298, N276);
or OR4 (N299, N285, N49, N10, N139);
xor XOR2 (N300, N297, N59);
or OR4 (N301, N295, N183, N174, N163);
not NOT1 (N302, N291);
nand NAND4 (N303, N278, N165, N208, N259);
not NOT1 (N304, N300);
not NOT1 (N305, N302);
xor XOR2 (N306, N299, N17);
nand NAND3 (N307, N304, N104, N6);
or OR2 (N308, N307, N261);
not NOT1 (N309, N305);
not NOT1 (N310, N301);
and AND4 (N311, N293, N98, N6, N102);
not NOT1 (N312, N309);
xor XOR2 (N313, N308, N297);
buf BUF1 (N314, N310);
or OR2 (N315, N306, N27);
nand NAND4 (N316, N312, N36, N124, N14);
nand NAND2 (N317, N315, N223);
buf BUF1 (N318, N316);
and AND2 (N319, N303, N115);
not NOT1 (N320, N294);
nand NAND3 (N321, N298, N65, N251);
nand NAND2 (N322, N320, N80);
nand NAND2 (N323, N319, N131);
not NOT1 (N324, N321);
xor XOR2 (N325, N322, N314);
buf BUF1 (N326, N150);
and AND4 (N327, N318, N95, N134, N210);
and AND3 (N328, N325, N314, N66);
and AND4 (N329, N311, N275, N239, N318);
or OR2 (N330, N324, N210);
not NOT1 (N331, N317);
buf BUF1 (N332, N326);
and AND4 (N333, N296, N203, N303, N130);
and AND3 (N334, N329, N173, N91);
xor XOR2 (N335, N327, N122);
and AND4 (N336, N334, N325, N40, N89);
not NOT1 (N337, N328);
nand NAND2 (N338, N330, N2);
nor NOR4 (N339, N335, N14, N42, N147);
not NOT1 (N340, N323);
not NOT1 (N341, N337);
or OR4 (N342, N341, N323, N220, N47);
nor NOR2 (N343, N332, N155);
or OR4 (N344, N340, N74, N111, N158);
xor XOR2 (N345, N344, N176);
nor NOR4 (N346, N339, N51, N167, N210);
not NOT1 (N347, N313);
or OR2 (N348, N342, N81);
and AND2 (N349, N343, N244);
nor NOR3 (N350, N346, N268, N80);
buf BUF1 (N351, N331);
not NOT1 (N352, N351);
xor XOR2 (N353, N352, N269);
xor XOR2 (N354, N347, N145);
or OR3 (N355, N348, N352, N112);
xor XOR2 (N356, N355, N45);
xor XOR2 (N357, N354, N8);
and AND2 (N358, N336, N143);
and AND3 (N359, N338, N315, N126);
and AND4 (N360, N287, N92, N182, N65);
xor XOR2 (N361, N350, N286);
nand NAND3 (N362, N349, N340, N88);
nand NAND4 (N363, N345, N17, N216, N329);
and AND2 (N364, N359, N67);
xor XOR2 (N365, N356, N215);
not NOT1 (N366, N360);
not NOT1 (N367, N366);
or OR2 (N368, N357, N59);
buf BUF1 (N369, N333);
and AND3 (N370, N362, N188, N369);
not NOT1 (N371, N265);
and AND4 (N372, N367, N184, N7, N309);
not NOT1 (N373, N370);
xor XOR2 (N374, N372, N273);
xor XOR2 (N375, N358, N66);
xor XOR2 (N376, N365, N60);
or OR3 (N377, N375, N131, N351);
nand NAND4 (N378, N373, N29, N163, N223);
nand NAND4 (N379, N377, N363, N160, N201);
or OR3 (N380, N364, N261, N100);
xor XOR2 (N381, N33, N315);
xor XOR2 (N382, N353, N362);
or OR3 (N383, N378, N17, N203);
nand NAND4 (N384, N382, N347, N220, N98);
or OR4 (N385, N379, N28, N138, N301);
and AND2 (N386, N383, N146);
not NOT1 (N387, N381);
or OR2 (N388, N368, N114);
and AND2 (N389, N387, N302);
buf BUF1 (N390, N388);
or OR4 (N391, N385, N111, N269, N329);
nor NOR2 (N392, N374, N44);
xor XOR2 (N393, N390, N299);
or OR4 (N394, N392, N343, N62, N383);
and AND2 (N395, N391, N94);
xor XOR2 (N396, N380, N10);
not NOT1 (N397, N361);
nor NOR3 (N398, N386, N373, N34);
buf BUF1 (N399, N393);
nor NOR2 (N400, N396, N179);
not NOT1 (N401, N371);
nand NAND2 (N402, N397, N157);
or OR3 (N403, N398, N300, N127);
not NOT1 (N404, N400);
or OR2 (N405, N376, N156);
buf BUF1 (N406, N384);
or OR2 (N407, N394, N175);
xor XOR2 (N408, N401, N233);
and AND2 (N409, N399, N15);
nor NOR2 (N410, N409, N230);
or OR3 (N411, N405, N112, N134);
and AND2 (N412, N402, N130);
buf BUF1 (N413, N407);
or OR4 (N414, N389, N115, N250, N314);
xor XOR2 (N415, N413, N104);
nand NAND2 (N416, N404, N403);
and AND4 (N417, N222, N222, N50, N6);
and AND2 (N418, N415, N264);
xor XOR2 (N419, N395, N205);
nand NAND3 (N420, N408, N6, N374);
and AND4 (N421, N412, N318, N137, N58);
not NOT1 (N422, N416);
nor NOR3 (N423, N414, N363, N22);
nand NAND2 (N424, N421, N111);
nand NAND2 (N425, N423, N63);
buf BUF1 (N426, N420);
or OR3 (N427, N417, N343, N337);
nand NAND2 (N428, N419, N25);
not NOT1 (N429, N424);
nand NAND4 (N430, N425, N379, N109, N20);
nor NOR4 (N431, N429, N289, N123, N195);
xor XOR2 (N432, N430, N253);
buf BUF1 (N433, N427);
buf BUF1 (N434, N418);
and AND4 (N435, N428, N17, N73, N279);
not NOT1 (N436, N431);
not NOT1 (N437, N422);
nor NOR2 (N438, N432, N32);
nand NAND2 (N439, N406, N20);
and AND3 (N440, N433, N195, N280);
not NOT1 (N441, N440);
or OR4 (N442, N441, N14, N337, N188);
xor XOR2 (N443, N439, N436);
not NOT1 (N444, N12);
buf BUF1 (N445, N434);
or OR2 (N446, N443, N262);
nor NOR4 (N447, N438, N315, N337, N301);
and AND3 (N448, N442, N362, N151);
and AND2 (N449, N411, N243);
or OR3 (N450, N410, N263, N174);
and AND4 (N451, N447, N276, N344, N50);
and AND2 (N452, N448, N157);
or OR3 (N453, N444, N391, N204);
or OR4 (N454, N435, N234, N270, N374);
or OR4 (N455, N450, N90, N305, N396);
nand NAND3 (N456, N455, N98, N198);
xor XOR2 (N457, N426, N246);
not NOT1 (N458, N453);
not NOT1 (N459, N446);
buf BUF1 (N460, N451);
buf BUF1 (N461, N452);
buf BUF1 (N462, N454);
nand NAND2 (N463, N457, N184);
not NOT1 (N464, N456);
nand NAND4 (N465, N460, N58, N252, N175);
not NOT1 (N466, N465);
nand NAND2 (N467, N458, N413);
buf BUF1 (N468, N467);
nand NAND3 (N469, N449, N254, N7);
nor NOR3 (N470, N459, N337, N72);
nand NAND2 (N471, N437, N440);
or OR4 (N472, N470, N86, N159, N140);
not NOT1 (N473, N468);
nand NAND4 (N474, N471, N449, N208, N469);
or OR2 (N475, N35, N75);
or OR2 (N476, N466, N295);
not NOT1 (N477, N476);
or OR2 (N478, N473, N130);
and AND3 (N479, N445, N278, N147);
nand NAND3 (N480, N474, N75, N478);
and AND3 (N481, N318, N388, N259);
nand NAND3 (N482, N481, N308, N194);
and AND3 (N483, N472, N86, N204);
buf BUF1 (N484, N461);
or OR4 (N485, N480, N478, N321, N5);
and AND2 (N486, N462, N332);
nor NOR4 (N487, N483, N46, N115, N424);
xor XOR2 (N488, N477, N374);
or OR4 (N489, N463, N316, N75, N79);
nor NOR2 (N490, N489, N16);
nor NOR2 (N491, N482, N197);
not NOT1 (N492, N490);
buf BUF1 (N493, N487);
buf BUF1 (N494, N491);
nor NOR4 (N495, N475, N152, N402, N222);
nor NOR4 (N496, N492, N476, N366, N64);
or OR4 (N497, N493, N428, N224, N466);
xor XOR2 (N498, N464, N164);
not NOT1 (N499, N498);
and AND3 (N500, N479, N71, N279);
nor NOR4 (N501, N486, N104, N224, N431);
buf BUF1 (N502, N497);
nor NOR3 (N503, N501, N223, N490);
xor XOR2 (N504, N502, N191);
or OR3 (N505, N494, N368, N189);
buf BUF1 (N506, N505);
buf BUF1 (N507, N500);
nand NAND4 (N508, N506, N446, N147, N229);
buf BUF1 (N509, N504);
nand NAND2 (N510, N495, N487);
or OR4 (N511, N484, N142, N226, N247);
xor XOR2 (N512, N509, N328);
not NOT1 (N513, N511);
xor XOR2 (N514, N510, N157);
or OR2 (N515, N514, N317);
xor XOR2 (N516, N485, N109);
not NOT1 (N517, N503);
and AND2 (N518, N516, N432);
or OR4 (N519, N517, N398, N448, N17);
buf BUF1 (N520, N508);
not NOT1 (N521, N520);
not NOT1 (N522, N515);
or OR4 (N523, N512, N496, N30, N30);
buf BUF1 (N524, N380);
xor XOR2 (N525, N518, N417);
or OR2 (N526, N523, N138);
and AND3 (N527, N522, N209, N184);
buf BUF1 (N528, N527);
buf BUF1 (N529, N513);
or OR3 (N530, N488, N201, N475);
or OR4 (N531, N499, N6, N177, N432);
buf BUF1 (N532, N528);
or OR2 (N533, N529, N462);
or OR3 (N534, N519, N270, N217);
nand NAND2 (N535, N507, N486);
nor NOR4 (N536, N525, N109, N201, N133);
or OR2 (N537, N534, N220);
and AND4 (N538, N533, N490, N354, N312);
and AND2 (N539, N524, N290);
nor NOR2 (N540, N526, N173);
nor NOR4 (N541, N536, N270, N109, N435);
not NOT1 (N542, N538);
and AND2 (N543, N535, N72);
xor XOR2 (N544, N521, N11);
or OR3 (N545, N537, N239, N427);
buf BUF1 (N546, N531);
buf BUF1 (N547, N546);
and AND4 (N548, N532, N102, N179, N193);
nor NOR2 (N549, N540, N5);
xor XOR2 (N550, N542, N277);
nand NAND2 (N551, N544, N54);
buf BUF1 (N552, N543);
and AND3 (N553, N549, N70, N30);
not NOT1 (N554, N547);
nand NAND4 (N555, N552, N230, N18, N508);
nor NOR2 (N556, N539, N322);
and AND3 (N557, N541, N271, N155);
nor NOR2 (N558, N548, N289);
nor NOR2 (N559, N545, N6);
and AND3 (N560, N530, N107, N331);
xor XOR2 (N561, N554, N448);
nand NAND4 (N562, N555, N23, N26, N304);
nor NOR3 (N563, N561, N269, N173);
xor XOR2 (N564, N558, N312);
and AND3 (N565, N563, N77, N211);
and AND2 (N566, N550, N483);
nor NOR3 (N567, N551, N105, N217);
nor NOR2 (N568, N553, N107);
nor NOR3 (N569, N557, N211, N316);
or OR3 (N570, N559, N334, N122);
nor NOR4 (N571, N569, N269, N68, N246);
buf BUF1 (N572, N564);
xor XOR2 (N573, N568, N114);
and AND2 (N574, N567, N488);
buf BUF1 (N575, N560);
buf BUF1 (N576, N556);
xor XOR2 (N577, N573, N92);
or OR3 (N578, N570, N147, N139);
not NOT1 (N579, N576);
and AND2 (N580, N575, N524);
or OR3 (N581, N572, N358, N46);
nand NAND4 (N582, N571, N146, N540, N214);
and AND3 (N583, N582, N146, N321);
and AND4 (N584, N579, N395, N86, N439);
nand NAND2 (N585, N584, N365);
and AND4 (N586, N585, N251, N454, N55);
xor XOR2 (N587, N566, N260);
xor XOR2 (N588, N580, N271);
buf BUF1 (N589, N581);
and AND3 (N590, N587, N142, N194);
buf BUF1 (N591, N562);
xor XOR2 (N592, N586, N438);
xor XOR2 (N593, N578, N410);
and AND3 (N594, N583, N20, N504);
nand NAND3 (N595, N593, N472, N102);
not NOT1 (N596, N589);
and AND4 (N597, N595, N79, N117, N17);
nand NAND4 (N598, N594, N547, N227, N340);
xor XOR2 (N599, N590, N92);
buf BUF1 (N600, N574);
or OR2 (N601, N598, N525);
nor NOR3 (N602, N599, N202, N526);
not NOT1 (N603, N588);
nand NAND2 (N604, N592, N125);
and AND3 (N605, N577, N69, N570);
not NOT1 (N606, N601);
buf BUF1 (N607, N606);
nor NOR2 (N608, N607, N477);
not NOT1 (N609, N603);
and AND3 (N610, N596, N180, N209);
nand NAND3 (N611, N591, N448, N54);
or OR4 (N612, N608, N596, N386, N179);
xor XOR2 (N613, N610, N434);
or OR4 (N614, N605, N91, N602, N151);
buf BUF1 (N615, N18);
nor NOR3 (N616, N612, N434, N163);
and AND3 (N617, N614, N89, N352);
not NOT1 (N618, N617);
nor NOR4 (N619, N615, N491, N350, N439);
not NOT1 (N620, N565);
or OR3 (N621, N619, N296, N441);
or OR3 (N622, N616, N367, N92);
or OR2 (N623, N618, N420);
not NOT1 (N624, N600);
or OR2 (N625, N613, N299);
buf BUF1 (N626, N622);
nand NAND4 (N627, N621, N181, N300, N76);
buf BUF1 (N628, N626);
nor NOR3 (N629, N623, N278, N563);
or OR2 (N630, N627, N445);
and AND3 (N631, N620, N256, N110);
xor XOR2 (N632, N597, N340);
xor XOR2 (N633, N631, N118);
xor XOR2 (N634, N625, N358);
nand NAND4 (N635, N624, N364, N259, N472);
nand NAND4 (N636, N609, N459, N13, N127);
xor XOR2 (N637, N634, N427);
buf BUF1 (N638, N611);
not NOT1 (N639, N629);
or OR4 (N640, N638, N171, N526, N203);
or OR4 (N641, N630, N530, N576, N205);
nor NOR2 (N642, N636, N363);
or OR3 (N643, N635, N27, N124);
and AND3 (N644, N643, N297, N53);
or OR4 (N645, N640, N288, N266, N250);
nor NOR2 (N646, N628, N432);
not NOT1 (N647, N645);
or OR4 (N648, N633, N61, N506, N561);
and AND2 (N649, N639, N132);
buf BUF1 (N650, N641);
not NOT1 (N651, N647);
or OR4 (N652, N649, N49, N243, N166);
nor NOR3 (N653, N642, N440, N82);
or OR2 (N654, N646, N111);
xor XOR2 (N655, N653, N598);
nor NOR2 (N656, N604, N98);
xor XOR2 (N657, N654, N137);
and AND2 (N658, N637, N100);
buf BUF1 (N659, N652);
nand NAND4 (N660, N659, N252, N438, N72);
nand NAND2 (N661, N660, N180);
not NOT1 (N662, N651);
nand NAND3 (N663, N632, N604, N434);
and AND3 (N664, N663, N216, N357);
nand NAND2 (N665, N664, N498);
buf BUF1 (N666, N650);
and AND2 (N667, N658, N449);
not NOT1 (N668, N661);
and AND4 (N669, N648, N394, N269, N536);
buf BUF1 (N670, N655);
nor NOR3 (N671, N666, N608, N142);
nand NAND4 (N672, N667, N474, N509, N136);
or OR3 (N673, N668, N588, N485);
and AND2 (N674, N656, N189);
buf BUF1 (N675, N644);
nand NAND2 (N676, N669, N400);
nor NOR2 (N677, N676, N330);
nor NOR3 (N678, N665, N586, N175);
not NOT1 (N679, N662);
nand NAND3 (N680, N679, N553, N202);
or OR3 (N681, N677, N496, N671);
nand NAND2 (N682, N331, N234);
and AND4 (N683, N680, N186, N390, N651);
not NOT1 (N684, N683);
nor NOR3 (N685, N681, N671, N276);
or OR3 (N686, N673, N449, N369);
or OR2 (N687, N684, N402);
or OR2 (N688, N672, N684);
and AND3 (N689, N674, N300, N32);
nor NOR4 (N690, N687, N599, N267, N590);
not NOT1 (N691, N685);
or OR2 (N692, N678, N271);
or OR4 (N693, N689, N302, N460, N206);
nor NOR2 (N694, N657, N173);
nand NAND3 (N695, N694, N370, N243);
nor NOR4 (N696, N675, N386, N108, N402);
and AND3 (N697, N690, N577, N617);
and AND4 (N698, N697, N98, N629, N460);
and AND2 (N699, N688, N14);
nand NAND3 (N700, N682, N651, N164);
nor NOR4 (N701, N686, N577, N126, N24);
and AND4 (N702, N699, N216, N422, N541);
and AND3 (N703, N698, N185, N44);
nor NOR3 (N704, N670, N71, N472);
nor NOR2 (N705, N700, N571);
and AND2 (N706, N701, N132);
and AND2 (N707, N705, N246);
buf BUF1 (N708, N707);
nor NOR2 (N709, N706, N196);
buf BUF1 (N710, N709);
or OR4 (N711, N703, N82, N537, N209);
and AND4 (N712, N711, N514, N58, N52);
or OR4 (N713, N704, N266, N248, N691);
nor NOR3 (N714, N600, N27, N654);
not NOT1 (N715, N712);
buf BUF1 (N716, N695);
buf BUF1 (N717, N716);
nor NOR4 (N718, N693, N423, N671, N312);
and AND3 (N719, N714, N269, N201);
buf BUF1 (N720, N719);
nand NAND4 (N721, N713, N524, N552, N379);
nand NAND3 (N722, N702, N709, N137);
or OR2 (N723, N720, N462);
buf BUF1 (N724, N721);
nor NOR3 (N725, N722, N170, N507);
nand NAND3 (N726, N692, N240, N646);
nor NOR2 (N727, N715, N271);
not NOT1 (N728, N725);
and AND2 (N729, N723, N603);
or OR3 (N730, N718, N242, N384);
and AND4 (N731, N728, N630, N209, N532);
and AND2 (N732, N696, N73);
not NOT1 (N733, N727);
and AND2 (N734, N729, N63);
not NOT1 (N735, N724);
nor NOR4 (N736, N730, N384, N564, N208);
not NOT1 (N737, N731);
nor NOR3 (N738, N732, N185, N682);
buf BUF1 (N739, N737);
and AND3 (N740, N736, N89, N547);
nand NAND3 (N741, N726, N64, N555);
nor NOR2 (N742, N740, N668);
and AND4 (N743, N742, N320, N437, N98);
xor XOR2 (N744, N733, N39);
and AND2 (N745, N735, N510);
not NOT1 (N746, N738);
nand NAND4 (N747, N746, N712, N182, N666);
xor XOR2 (N748, N734, N661);
buf BUF1 (N749, N744);
nor NOR4 (N750, N717, N559, N379, N73);
not NOT1 (N751, N743);
and AND2 (N752, N710, N488);
buf BUF1 (N753, N708);
nand NAND2 (N754, N753, N157);
or OR2 (N755, N750, N412);
and AND3 (N756, N747, N477, N556);
xor XOR2 (N757, N739, N79);
nor NOR4 (N758, N749, N259, N86, N257);
and AND3 (N759, N752, N643, N546);
nand NAND3 (N760, N754, N542, N124);
nor NOR3 (N761, N745, N283, N567);
buf BUF1 (N762, N756);
and AND4 (N763, N757, N482, N204, N673);
nor NOR2 (N764, N758, N549);
nand NAND2 (N765, N741, N91);
xor XOR2 (N766, N762, N644);
nand NAND2 (N767, N760, N561);
not NOT1 (N768, N761);
buf BUF1 (N769, N765);
and AND3 (N770, N768, N514, N763);
buf BUF1 (N771, N70);
and AND4 (N772, N771, N613, N663, N187);
buf BUF1 (N773, N759);
nand NAND4 (N774, N770, N688, N2, N373);
not NOT1 (N775, N773);
nor NOR4 (N776, N772, N53, N413, N620);
xor XOR2 (N777, N769, N327);
buf BUF1 (N778, N776);
nand NAND3 (N779, N774, N611, N539);
nand NAND2 (N780, N779, N487);
not NOT1 (N781, N764);
and AND2 (N782, N780, N619);
or OR2 (N783, N778, N522);
and AND4 (N784, N755, N106, N61, N735);
nor NOR3 (N785, N751, N308, N404);
or OR4 (N786, N782, N333, N374, N389);
xor XOR2 (N787, N785, N78);
xor XOR2 (N788, N783, N25);
nand NAND3 (N789, N766, N677, N128);
or OR4 (N790, N777, N532, N179, N775);
or OR3 (N791, N494, N597, N210);
or OR3 (N792, N787, N783, N638);
nand NAND3 (N793, N788, N439, N619);
buf BUF1 (N794, N790);
nor NOR4 (N795, N791, N423, N432, N447);
nor NOR3 (N796, N748, N792, N771);
or OR2 (N797, N520, N227);
buf BUF1 (N798, N794);
nand NAND2 (N799, N784, N305);
not NOT1 (N800, N793);
buf BUF1 (N801, N786);
buf BUF1 (N802, N797);
nor NOR4 (N803, N789, N91, N211, N407);
buf BUF1 (N804, N799);
and AND2 (N805, N803, N140);
not NOT1 (N806, N796);
and AND2 (N807, N805, N259);
and AND2 (N808, N807, N55);
buf BUF1 (N809, N781);
and AND3 (N810, N795, N60, N213);
not NOT1 (N811, N809);
or OR2 (N812, N801, N624);
buf BUF1 (N813, N767);
and AND2 (N814, N808, N768);
and AND4 (N815, N813, N289, N585, N513);
nand NAND3 (N816, N806, N117, N451);
or OR2 (N817, N804, N510);
endmodule