// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21;

output N1519,N1514,N1516,N1518,N1520,N1504,N1508,N1505,N1512,N1521;

nand NAND2 (N22, N6, N21);
and AND2 (N23, N21, N4);
nor NOR2 (N24, N14, N11);
xor XOR2 (N25, N12, N22);
and AND4 (N26, N10, N1, N5, N13);
and AND2 (N27, N25, N8);
not NOT1 (N28, N19);
nand NAND4 (N29, N26, N15, N21, N6);
or OR4 (N30, N15, N19, N17, N25);
xor XOR2 (N31, N28, N28);
nand NAND3 (N32, N1, N7, N22);
or OR4 (N33, N27, N19, N29, N22);
nand NAND4 (N34, N13, N12, N10, N8);
nand NAND2 (N35, N30, N5);
xor XOR2 (N36, N12, N3);
xor XOR2 (N37, N8, N9);
not NOT1 (N38, N34);
nand NAND2 (N39, N17, N10);
buf BUF1 (N40, N38);
nand NAND3 (N41, N40, N35, N30);
and AND3 (N42, N25, N23, N40);
xor XOR2 (N43, N35, N26);
nand NAND2 (N44, N31, N37);
buf BUF1 (N45, N7);
nor NOR2 (N46, N36, N25);
and AND2 (N47, N43, N9);
not NOT1 (N48, N41);
and AND4 (N49, N44, N44, N11, N39);
and AND4 (N50, N29, N27, N16, N12);
xor XOR2 (N51, N24, N46);
or OR2 (N52, N43, N14);
nor NOR4 (N53, N47, N31, N43, N42);
buf BUF1 (N54, N5);
nor NOR3 (N55, N50, N27, N5);
xor XOR2 (N56, N53, N14);
or OR2 (N57, N32, N31);
xor XOR2 (N58, N54, N56);
buf BUF1 (N59, N14);
nand NAND2 (N60, N51, N56);
xor XOR2 (N61, N48, N44);
not NOT1 (N62, N45);
xor XOR2 (N63, N55, N59);
or OR2 (N64, N52, N29);
or OR2 (N65, N47, N42);
buf BUF1 (N66, N64);
buf BUF1 (N67, N33);
nand NAND4 (N68, N66, N3, N38, N40);
and AND3 (N69, N58, N54, N33);
and AND2 (N70, N57, N8);
not NOT1 (N71, N60);
nor NOR3 (N72, N63, N42, N55);
nand NAND4 (N73, N70, N27, N14, N63);
not NOT1 (N74, N71);
or OR4 (N75, N73, N61, N1, N73);
nand NAND2 (N76, N64, N64);
and AND4 (N77, N72, N2, N29, N57);
nand NAND4 (N78, N75, N65, N43, N8);
nor NOR2 (N79, N70, N8);
and AND3 (N80, N69, N48, N13);
not NOT1 (N81, N68);
or OR4 (N82, N80, N77, N61, N9);
nor NOR2 (N83, N8, N81);
buf BUF1 (N84, N68);
or OR3 (N85, N76, N23, N47);
not NOT1 (N86, N62);
xor XOR2 (N87, N85, N60);
xor XOR2 (N88, N78, N21);
buf BUF1 (N89, N67);
or OR4 (N90, N84, N15, N50, N63);
or OR2 (N91, N89, N32);
xor XOR2 (N92, N74, N69);
nand NAND4 (N93, N83, N39, N47, N39);
xor XOR2 (N94, N88, N62);
or OR3 (N95, N82, N52, N21);
and AND2 (N96, N95, N19);
and AND4 (N97, N94, N26, N53, N31);
nor NOR2 (N98, N87, N79);
and AND4 (N99, N98, N8, N96, N38);
and AND3 (N100, N56, N64, N11);
not NOT1 (N101, N89);
nand NAND3 (N102, N93, N51, N72);
and AND2 (N103, N91, N2);
nor NOR3 (N104, N97, N40, N75);
and AND3 (N105, N101, N90, N87);
xor XOR2 (N106, N54, N41);
not NOT1 (N107, N100);
or OR2 (N108, N99, N59);
nor NOR2 (N109, N108, N75);
nor NOR3 (N110, N107, N71, N31);
and AND2 (N111, N104, N39);
buf BUF1 (N112, N111);
nand NAND3 (N113, N92, N51, N26);
buf BUF1 (N114, N86);
nor NOR4 (N115, N112, N106, N50, N107);
not NOT1 (N116, N5);
and AND4 (N117, N102, N38, N19, N66);
nand NAND3 (N118, N114, N9, N64);
and AND4 (N119, N103, N58, N66, N9);
nor NOR2 (N120, N105, N78);
xor XOR2 (N121, N119, N89);
nor NOR4 (N122, N118, N117, N26, N1);
nand NAND4 (N123, N76, N25, N22, N37);
nor NOR2 (N124, N110, N67);
or OR2 (N125, N116, N105);
or OR3 (N126, N115, N93, N92);
buf BUF1 (N127, N124);
nand NAND2 (N128, N49, N95);
nor NOR3 (N129, N125, N92, N55);
nand NAND3 (N130, N121, N45, N96);
and AND2 (N131, N130, N102);
nand NAND3 (N132, N122, N109, N83);
and AND4 (N133, N106, N35, N37, N30);
xor XOR2 (N134, N131, N59);
and AND4 (N135, N113, N17, N76, N20);
nor NOR3 (N136, N120, N92, N87);
xor XOR2 (N137, N136, N60);
xor XOR2 (N138, N129, N97);
buf BUF1 (N139, N134);
not NOT1 (N140, N133);
buf BUF1 (N141, N126);
nand NAND3 (N142, N140, N136, N1);
or OR4 (N143, N127, N48, N97, N7);
not NOT1 (N144, N128);
nand NAND2 (N145, N137, N54);
not NOT1 (N146, N132);
xor XOR2 (N147, N123, N106);
not NOT1 (N148, N145);
and AND4 (N149, N146, N50, N113, N37);
nand NAND2 (N150, N143, N63);
xor XOR2 (N151, N147, N49);
not NOT1 (N152, N135);
nand NAND3 (N153, N150, N29, N35);
buf BUF1 (N154, N141);
xor XOR2 (N155, N144, N4);
and AND2 (N156, N155, N33);
and AND3 (N157, N139, N85, N113);
nor NOR3 (N158, N149, N76, N37);
not NOT1 (N159, N157);
or OR4 (N160, N153, N11, N122, N25);
and AND2 (N161, N156, N26);
or OR2 (N162, N158, N89);
nand NAND4 (N163, N142, N48, N13, N149);
not NOT1 (N164, N148);
not NOT1 (N165, N164);
not NOT1 (N166, N165);
nand NAND2 (N167, N152, N135);
not NOT1 (N168, N167);
and AND3 (N169, N151, N18, N29);
and AND2 (N170, N154, N51);
or OR2 (N171, N168, N167);
or OR2 (N172, N170, N144);
nor NOR3 (N173, N166, N33, N49);
not NOT1 (N174, N162);
xor XOR2 (N175, N161, N167);
or OR4 (N176, N160, N76, N144, N145);
not NOT1 (N177, N173);
nor NOR3 (N178, N174, N115, N157);
xor XOR2 (N179, N159, N83);
buf BUF1 (N180, N178);
or OR4 (N181, N138, N83, N140, N72);
xor XOR2 (N182, N171, N66);
buf BUF1 (N183, N176);
or OR4 (N184, N181, N98, N80, N12);
and AND3 (N185, N172, N90, N11);
xor XOR2 (N186, N180, N62);
xor XOR2 (N187, N183, N88);
and AND3 (N188, N177, N150, N166);
nor NOR4 (N189, N188, N106, N160, N182);
buf BUF1 (N190, N83);
nor NOR3 (N191, N186, N148, N29);
nand NAND4 (N192, N187, N190, N57, N139);
nor NOR3 (N193, N119, N120, N8);
buf BUF1 (N194, N185);
and AND2 (N195, N191, N135);
xor XOR2 (N196, N175, N16);
or OR2 (N197, N184, N33);
and AND3 (N198, N179, N46, N137);
and AND4 (N199, N193, N159, N150, N196);
buf BUF1 (N200, N10);
nand NAND2 (N201, N189, N59);
nor NOR2 (N202, N194, N101);
nand NAND3 (N203, N202, N90, N129);
or OR2 (N204, N195, N64);
xor XOR2 (N205, N201, N118);
nand NAND4 (N206, N163, N157, N67, N158);
not NOT1 (N207, N192);
buf BUF1 (N208, N204);
or OR4 (N209, N206, N10, N148, N18);
xor XOR2 (N210, N207, N54);
buf BUF1 (N211, N169);
or OR2 (N212, N209, N113);
not NOT1 (N213, N208);
or OR4 (N214, N213, N120, N47, N117);
buf BUF1 (N215, N197);
xor XOR2 (N216, N203, N164);
nand NAND3 (N217, N205, N146, N106);
not NOT1 (N218, N200);
nand NAND3 (N219, N199, N66, N62);
and AND4 (N220, N198, N41, N186, N107);
not NOT1 (N221, N217);
or OR2 (N222, N212, N138);
and AND4 (N223, N211, N3, N29, N180);
xor XOR2 (N224, N216, N132);
nor NOR4 (N225, N210, N8, N187, N179);
or OR3 (N226, N218, N37, N29);
xor XOR2 (N227, N220, N38);
nand NAND2 (N228, N221, N114);
xor XOR2 (N229, N215, N100);
or OR3 (N230, N228, N163, N180);
not NOT1 (N231, N229);
and AND2 (N232, N223, N91);
nand NAND4 (N233, N230, N170, N211, N138);
not NOT1 (N234, N231);
xor XOR2 (N235, N234, N45);
not NOT1 (N236, N226);
and AND3 (N237, N224, N80, N89);
buf BUF1 (N238, N214);
nor NOR4 (N239, N227, N63, N164, N133);
buf BUF1 (N240, N238);
and AND3 (N241, N240, N38, N31);
nor NOR3 (N242, N235, N86, N225);
nand NAND2 (N243, N238, N119);
xor XOR2 (N244, N233, N159);
not NOT1 (N245, N237);
xor XOR2 (N246, N232, N219);
nor NOR4 (N247, N60, N216, N189, N135);
xor XOR2 (N248, N242, N109);
not NOT1 (N249, N222);
xor XOR2 (N250, N249, N142);
nor NOR3 (N251, N243, N26, N59);
not NOT1 (N252, N247);
nor NOR4 (N253, N239, N41, N231, N189);
and AND2 (N254, N236, N74);
not NOT1 (N255, N254);
nand NAND2 (N256, N251, N203);
or OR2 (N257, N252, N214);
or OR4 (N258, N248, N245, N94, N74);
not NOT1 (N259, N137);
not NOT1 (N260, N246);
not NOT1 (N261, N241);
xor XOR2 (N262, N258, N229);
nand NAND4 (N263, N262, N129, N201, N184);
xor XOR2 (N264, N255, N26);
buf BUF1 (N265, N264);
not NOT1 (N266, N261);
or OR3 (N267, N260, N174, N110);
or OR3 (N268, N263, N51, N192);
buf BUF1 (N269, N265);
not NOT1 (N270, N256);
and AND4 (N271, N270, N69, N63, N86);
xor XOR2 (N272, N257, N89);
and AND2 (N273, N272, N160);
and AND4 (N274, N266, N144, N68, N206);
nor NOR2 (N275, N253, N245);
not NOT1 (N276, N273);
xor XOR2 (N277, N250, N68);
not NOT1 (N278, N275);
not NOT1 (N279, N278);
buf BUF1 (N280, N276);
nand NAND3 (N281, N277, N66, N274);
not NOT1 (N282, N150);
xor XOR2 (N283, N268, N223);
nor NOR4 (N284, N282, N30, N102, N193);
nor NOR3 (N285, N269, N82, N24);
xor XOR2 (N286, N271, N32);
xor XOR2 (N287, N285, N191);
buf BUF1 (N288, N287);
buf BUF1 (N289, N284);
buf BUF1 (N290, N286);
nor NOR2 (N291, N281, N280);
not NOT1 (N292, N9);
nor NOR4 (N293, N292, N108, N173, N267);
and AND4 (N294, N61, N215, N230, N200);
and AND4 (N295, N290, N128, N145, N75);
buf BUF1 (N296, N279);
and AND3 (N297, N283, N222, N53);
nand NAND2 (N298, N289, N20);
nand NAND4 (N299, N259, N7, N170, N43);
nand NAND2 (N300, N297, N38);
xor XOR2 (N301, N299, N165);
nand NAND4 (N302, N288, N174, N161, N199);
and AND4 (N303, N244, N35, N34, N291);
or OR2 (N304, N246, N201);
not NOT1 (N305, N302);
nand NAND2 (N306, N294, N71);
nor NOR4 (N307, N306, N296, N28, N4);
or OR3 (N308, N260, N58, N150);
or OR2 (N309, N295, N215);
xor XOR2 (N310, N309, N56);
buf BUF1 (N311, N308);
nand NAND3 (N312, N307, N166, N8);
and AND3 (N313, N303, N51, N115);
and AND4 (N314, N311, N62, N270, N18);
nor NOR4 (N315, N304, N263, N126, N231);
nand NAND2 (N316, N312, N310);
nor NOR4 (N317, N128, N78, N77, N55);
or OR2 (N318, N293, N49);
nand NAND4 (N319, N316, N165, N192, N7);
nor NOR4 (N320, N318, N142, N274, N118);
and AND2 (N321, N315, N150);
buf BUF1 (N322, N314);
or OR2 (N323, N320, N60);
or OR3 (N324, N305, N319, N16);
xor XOR2 (N325, N274, N151);
nor NOR2 (N326, N321, N225);
xor XOR2 (N327, N313, N233);
nor NOR4 (N328, N322, N96, N194, N258);
nor NOR2 (N329, N298, N225);
not NOT1 (N330, N328);
xor XOR2 (N331, N326, N182);
nor NOR4 (N332, N300, N255, N233, N163);
nor NOR3 (N333, N331, N276, N75);
and AND2 (N334, N332, N117);
or OR2 (N335, N329, N204);
nor NOR4 (N336, N324, N48, N275, N38);
not NOT1 (N337, N301);
buf BUF1 (N338, N330);
nor NOR3 (N339, N337, N180, N163);
buf BUF1 (N340, N335);
not NOT1 (N341, N340);
xor XOR2 (N342, N336, N174);
nand NAND4 (N343, N327, N282, N264, N287);
not NOT1 (N344, N317);
nor NOR2 (N345, N339, N73);
nand NAND4 (N346, N334, N325, N234, N185);
or OR3 (N347, N76, N78, N53);
buf BUF1 (N348, N341);
or OR2 (N349, N323, N100);
xor XOR2 (N350, N344, N119);
buf BUF1 (N351, N350);
nor NOR2 (N352, N347, N40);
nand NAND2 (N353, N343, N243);
buf BUF1 (N354, N338);
or OR2 (N355, N353, N16);
or OR4 (N356, N333, N281, N71, N98);
buf BUF1 (N357, N342);
or OR3 (N358, N348, N237, N254);
xor XOR2 (N359, N351, N301);
nand NAND2 (N360, N359, N6);
nand NAND4 (N361, N360, N115, N314, N356);
nor NOR4 (N362, N11, N240, N68, N243);
and AND2 (N363, N345, N59);
not NOT1 (N364, N352);
buf BUF1 (N365, N354);
xor XOR2 (N366, N349, N202);
not NOT1 (N367, N366);
not NOT1 (N368, N361);
and AND2 (N369, N365, N320);
or OR4 (N370, N357, N205, N212, N265);
not NOT1 (N371, N370);
or OR4 (N372, N367, N205, N242, N255);
xor XOR2 (N373, N358, N247);
nand NAND3 (N374, N372, N62, N238);
buf BUF1 (N375, N369);
and AND4 (N376, N363, N246, N51, N200);
buf BUF1 (N377, N374);
xor XOR2 (N378, N362, N219);
nand NAND3 (N379, N378, N130, N205);
xor XOR2 (N380, N375, N260);
xor XOR2 (N381, N364, N119);
and AND3 (N382, N381, N158, N329);
nor NOR2 (N383, N346, N357);
and AND2 (N384, N382, N67);
nand NAND2 (N385, N379, N144);
not NOT1 (N386, N377);
buf BUF1 (N387, N383);
nor NOR2 (N388, N373, N369);
or OR2 (N389, N387, N19);
and AND3 (N390, N386, N257, N135);
and AND4 (N391, N371, N292, N265, N35);
nand NAND2 (N392, N388, N4);
nand NAND2 (N393, N390, N32);
nand NAND4 (N394, N391, N67, N4, N224);
and AND3 (N395, N393, N304, N252);
and AND4 (N396, N384, N378, N170, N14);
nor NOR4 (N397, N396, N282, N93, N234);
nand NAND2 (N398, N392, N214);
or OR2 (N399, N395, N237);
or OR4 (N400, N397, N296, N347, N265);
and AND4 (N401, N389, N128, N325, N199);
not NOT1 (N402, N380);
nor NOR3 (N403, N400, N294, N356);
buf BUF1 (N404, N398);
buf BUF1 (N405, N403);
buf BUF1 (N406, N394);
or OR2 (N407, N404, N268);
not NOT1 (N408, N406);
and AND3 (N409, N399, N250, N141);
not NOT1 (N410, N405);
nor NOR2 (N411, N410, N102);
nor NOR2 (N412, N408, N62);
buf BUF1 (N413, N355);
and AND3 (N414, N413, N223, N177);
and AND3 (N415, N412, N49, N201);
or OR2 (N416, N411, N363);
not NOT1 (N417, N402);
not NOT1 (N418, N417);
not NOT1 (N419, N401);
xor XOR2 (N420, N419, N224);
or OR3 (N421, N409, N34, N180);
or OR3 (N422, N407, N275, N228);
xor XOR2 (N423, N368, N372);
and AND4 (N424, N416, N267, N52, N375);
and AND3 (N425, N376, N373, N183);
or OR2 (N426, N415, N19);
xor XOR2 (N427, N414, N174);
nand NAND4 (N428, N421, N293, N208, N117);
or OR4 (N429, N428, N197, N27, N130);
and AND3 (N430, N424, N88, N100);
buf BUF1 (N431, N425);
xor XOR2 (N432, N418, N347);
buf BUF1 (N433, N423);
and AND4 (N434, N429, N62, N290, N125);
or OR2 (N435, N422, N290);
xor XOR2 (N436, N435, N429);
xor XOR2 (N437, N427, N82);
and AND4 (N438, N433, N324, N187, N135);
or OR4 (N439, N434, N267, N27, N33);
and AND3 (N440, N432, N253, N5);
not NOT1 (N441, N439);
nor NOR2 (N442, N437, N350);
or OR2 (N443, N440, N395);
not NOT1 (N444, N420);
xor XOR2 (N445, N436, N269);
or OR3 (N446, N385, N344, N327);
buf BUF1 (N447, N445);
nor NOR4 (N448, N426, N398, N291, N352);
nor NOR2 (N449, N438, N261);
or OR3 (N450, N443, N1, N58);
xor XOR2 (N451, N448, N429);
xor XOR2 (N452, N431, N211);
or OR4 (N453, N441, N156, N317, N238);
not NOT1 (N454, N452);
nand NAND2 (N455, N453, N318);
and AND3 (N456, N444, N384, N116);
or OR3 (N457, N454, N116, N217);
buf BUF1 (N458, N450);
and AND2 (N459, N447, N183);
not NOT1 (N460, N459);
xor XOR2 (N461, N456, N304);
not NOT1 (N462, N457);
nor NOR3 (N463, N462, N35, N172);
nand NAND4 (N464, N461, N167, N463, N206);
buf BUF1 (N465, N446);
nor NOR2 (N466, N149, N25);
nor NOR3 (N467, N442, N160, N365);
xor XOR2 (N468, N430, N18);
xor XOR2 (N469, N455, N10);
xor XOR2 (N470, N466, N240);
xor XOR2 (N471, N458, N45);
and AND4 (N472, N468, N370, N470, N241);
and AND2 (N473, N98, N420);
nand NAND2 (N474, N469, N425);
xor XOR2 (N475, N451, N346);
xor XOR2 (N476, N472, N415);
not NOT1 (N477, N475);
or OR2 (N478, N476, N436);
and AND3 (N479, N474, N310, N418);
buf BUF1 (N480, N465);
not NOT1 (N481, N477);
xor XOR2 (N482, N479, N381);
nor NOR4 (N483, N481, N357, N253, N150);
nand NAND2 (N484, N480, N147);
and AND3 (N485, N478, N116, N428);
buf BUF1 (N486, N449);
and AND3 (N487, N486, N393, N17);
buf BUF1 (N488, N483);
or OR4 (N489, N460, N465, N208, N436);
not NOT1 (N490, N482);
or OR4 (N491, N484, N55, N472, N276);
nor NOR3 (N492, N464, N148, N321);
and AND4 (N493, N488, N427, N478, N358);
xor XOR2 (N494, N489, N72);
nand NAND2 (N495, N490, N433);
nand NAND4 (N496, N471, N432, N410, N321);
and AND2 (N497, N496, N23);
not NOT1 (N498, N467);
and AND3 (N499, N485, N331, N338);
or OR3 (N500, N498, N281, N405);
and AND4 (N501, N497, N137, N33, N428);
and AND3 (N502, N487, N99, N464);
xor XOR2 (N503, N494, N422);
and AND4 (N504, N493, N298, N385, N258);
xor XOR2 (N505, N491, N90);
nand NAND2 (N506, N492, N495);
and AND3 (N507, N158, N350, N385);
nand NAND4 (N508, N500, N107, N300, N438);
nor NOR4 (N509, N501, N400, N304, N94);
or OR3 (N510, N504, N181, N353);
nand NAND2 (N511, N508, N329);
nand NAND2 (N512, N503, N176);
nand NAND2 (N513, N506, N51);
nor NOR2 (N514, N512, N365);
not NOT1 (N515, N473);
buf BUF1 (N516, N502);
and AND2 (N517, N510, N497);
nor NOR4 (N518, N511, N253, N93, N342);
xor XOR2 (N519, N517, N17);
or OR3 (N520, N516, N67, N438);
buf BUF1 (N521, N520);
buf BUF1 (N522, N509);
not NOT1 (N523, N522);
nor NOR4 (N524, N521, N482, N47, N507);
not NOT1 (N525, N69);
xor XOR2 (N526, N514, N404);
xor XOR2 (N527, N524, N94);
nor NOR4 (N528, N525, N161, N426, N284);
buf BUF1 (N529, N519);
nand NAND3 (N530, N523, N475, N268);
nor NOR2 (N531, N499, N108);
nor NOR3 (N532, N527, N350, N364);
and AND4 (N533, N518, N235, N200, N364);
or OR2 (N534, N513, N157);
nor NOR3 (N535, N515, N18, N386);
buf BUF1 (N536, N531);
not NOT1 (N537, N505);
xor XOR2 (N538, N532, N54);
and AND4 (N539, N528, N431, N276, N372);
nand NAND3 (N540, N535, N119, N6);
and AND4 (N541, N540, N286, N526, N146);
not NOT1 (N542, N474);
nor NOR3 (N543, N539, N159, N486);
and AND3 (N544, N530, N527, N124);
or OR3 (N545, N544, N366, N289);
and AND3 (N546, N542, N524, N56);
xor XOR2 (N547, N546, N66);
nand NAND3 (N548, N536, N15, N344);
or OR4 (N549, N534, N163, N316, N138);
or OR4 (N550, N549, N412, N205, N13);
nor NOR3 (N551, N538, N368, N428);
or OR4 (N552, N550, N9, N474, N525);
not NOT1 (N553, N552);
nor NOR2 (N554, N545, N433);
not NOT1 (N555, N547);
xor XOR2 (N556, N543, N314);
and AND3 (N557, N548, N420, N74);
and AND4 (N558, N533, N450, N536, N386);
buf BUF1 (N559, N541);
or OR3 (N560, N529, N95, N10);
nor NOR3 (N561, N551, N428, N15);
xor XOR2 (N562, N555, N378);
not NOT1 (N563, N560);
and AND2 (N564, N554, N534);
buf BUF1 (N565, N562);
nor NOR4 (N566, N537, N276, N3, N400);
nand NAND4 (N567, N556, N355, N514, N396);
xor XOR2 (N568, N557, N16);
not NOT1 (N569, N566);
nand NAND2 (N570, N565, N544);
not NOT1 (N571, N567);
nand NAND3 (N572, N561, N369, N160);
not NOT1 (N573, N563);
nand NAND4 (N574, N559, N104, N123, N378);
and AND4 (N575, N553, N486, N524, N336);
xor XOR2 (N576, N558, N356);
not NOT1 (N577, N574);
nand NAND3 (N578, N570, N91, N128);
nor NOR3 (N579, N576, N142, N193);
xor XOR2 (N580, N571, N74);
buf BUF1 (N581, N577);
buf BUF1 (N582, N569);
xor XOR2 (N583, N572, N417);
nor NOR3 (N584, N568, N240, N73);
nor NOR4 (N585, N580, N341, N382, N45);
buf BUF1 (N586, N581);
nor NOR2 (N587, N585, N302);
or OR4 (N588, N586, N31, N442, N544);
nand NAND4 (N589, N583, N140, N43, N442);
nand NAND2 (N590, N573, N441);
not NOT1 (N591, N582);
xor XOR2 (N592, N578, N69);
buf BUF1 (N593, N588);
and AND3 (N594, N591, N8, N207);
not NOT1 (N595, N590);
nor NOR4 (N596, N595, N62, N441, N503);
nand NAND2 (N597, N593, N558);
not NOT1 (N598, N596);
buf BUF1 (N599, N592);
not NOT1 (N600, N575);
not NOT1 (N601, N589);
or OR3 (N602, N594, N317, N153);
buf BUF1 (N603, N587);
buf BUF1 (N604, N600);
nand NAND3 (N605, N597, N430, N496);
xor XOR2 (N606, N599, N179);
and AND2 (N607, N584, N85);
or OR4 (N608, N606, N238, N100, N450);
buf BUF1 (N609, N579);
not NOT1 (N610, N601);
not NOT1 (N611, N607);
xor XOR2 (N612, N603, N549);
xor XOR2 (N613, N605, N597);
buf BUF1 (N614, N613);
nand NAND4 (N615, N610, N258, N240, N74);
nor NOR2 (N616, N609, N516);
or OR2 (N617, N616, N447);
not NOT1 (N618, N598);
nand NAND2 (N619, N615, N389);
or OR4 (N620, N619, N26, N503, N505);
not NOT1 (N621, N614);
or OR4 (N622, N602, N389, N459, N461);
and AND2 (N623, N621, N27);
not NOT1 (N624, N608);
not NOT1 (N625, N612);
and AND4 (N626, N620, N285, N563, N439);
xor XOR2 (N627, N622, N76);
nand NAND4 (N628, N617, N625, N498, N46);
buf BUF1 (N629, N419);
not NOT1 (N630, N629);
nand NAND2 (N631, N630, N361);
or OR3 (N632, N627, N409, N476);
nand NAND4 (N633, N626, N335, N185, N447);
nor NOR4 (N634, N611, N161, N379, N260);
buf BUF1 (N635, N631);
buf BUF1 (N636, N624);
buf BUF1 (N637, N633);
and AND2 (N638, N635, N521);
and AND3 (N639, N638, N612, N290);
nor NOR4 (N640, N632, N283, N632, N261);
nor NOR3 (N641, N564, N501, N224);
nand NAND3 (N642, N618, N625, N437);
nor NOR4 (N643, N641, N310, N604, N16);
buf BUF1 (N644, N44);
buf BUF1 (N645, N623);
nor NOR2 (N646, N640, N380);
or OR3 (N647, N646, N599, N512);
or OR4 (N648, N636, N295, N147, N641);
buf BUF1 (N649, N647);
nor NOR3 (N650, N642, N520, N69);
and AND2 (N651, N650, N213);
and AND2 (N652, N649, N263);
not NOT1 (N653, N644);
or OR2 (N654, N648, N85);
nand NAND3 (N655, N637, N202, N492);
not NOT1 (N656, N653);
not NOT1 (N657, N651);
xor XOR2 (N658, N645, N67);
and AND2 (N659, N658, N25);
or OR3 (N660, N652, N33, N460);
nor NOR2 (N661, N655, N557);
xor XOR2 (N662, N639, N652);
buf BUF1 (N663, N656);
not NOT1 (N664, N663);
buf BUF1 (N665, N664);
nand NAND3 (N666, N660, N170, N547);
not NOT1 (N667, N662);
nor NOR3 (N668, N657, N439, N602);
or OR3 (N669, N659, N524, N240);
buf BUF1 (N670, N668);
buf BUF1 (N671, N654);
nor NOR2 (N672, N643, N636);
nand NAND4 (N673, N665, N315, N424, N250);
not NOT1 (N674, N667);
xor XOR2 (N675, N661, N365);
not NOT1 (N676, N628);
xor XOR2 (N677, N673, N391);
nand NAND3 (N678, N666, N564, N559);
nor NOR2 (N679, N634, N660);
nor NOR3 (N680, N678, N114, N97);
nor NOR3 (N681, N679, N232, N277);
xor XOR2 (N682, N670, N597);
not NOT1 (N683, N674);
or OR4 (N684, N682, N545, N609, N397);
or OR2 (N685, N680, N208);
nor NOR2 (N686, N675, N658);
xor XOR2 (N687, N683, N670);
nand NAND3 (N688, N671, N175, N543);
not NOT1 (N689, N681);
buf BUF1 (N690, N686);
nor NOR3 (N691, N676, N684, N122);
buf BUF1 (N692, N486);
or OR3 (N693, N677, N274, N489);
or OR3 (N694, N691, N635, N419);
or OR2 (N695, N694, N246);
buf BUF1 (N696, N685);
xor XOR2 (N697, N695, N8);
buf BUF1 (N698, N672);
nand NAND4 (N699, N696, N24, N565, N229);
nand NAND2 (N700, N688, N620);
xor XOR2 (N701, N698, N688);
or OR4 (N702, N689, N181, N190, N496);
nand NAND3 (N703, N687, N325, N519);
xor XOR2 (N704, N701, N555);
xor XOR2 (N705, N699, N37);
or OR4 (N706, N702, N589, N577, N704);
and AND2 (N707, N158, N580);
and AND4 (N708, N692, N615, N509, N445);
or OR4 (N709, N708, N682, N9, N80);
buf BUF1 (N710, N706);
buf BUF1 (N711, N669);
xor XOR2 (N712, N697, N191);
or OR3 (N713, N709, N460, N182);
not NOT1 (N714, N707);
nand NAND2 (N715, N690, N140);
xor XOR2 (N716, N712, N380);
or OR2 (N717, N711, N44);
not NOT1 (N718, N703);
or OR4 (N719, N717, N124, N686, N561);
nand NAND3 (N720, N719, N403, N137);
not NOT1 (N721, N720);
nand NAND2 (N722, N718, N470);
and AND2 (N723, N721, N426);
and AND2 (N724, N723, N27);
xor XOR2 (N725, N693, N486);
or OR4 (N726, N724, N502, N50, N354);
or OR3 (N727, N726, N391, N246);
not NOT1 (N728, N716);
nor NOR3 (N729, N715, N517, N205);
or OR4 (N730, N727, N282, N66, N484);
and AND4 (N731, N722, N349, N289, N226);
not NOT1 (N732, N729);
or OR2 (N733, N714, N162);
nor NOR2 (N734, N731, N643);
xor XOR2 (N735, N700, N423);
not NOT1 (N736, N713);
xor XOR2 (N737, N725, N639);
and AND4 (N738, N733, N261, N383, N79);
or OR3 (N739, N732, N253, N404);
nor NOR3 (N740, N730, N310, N472);
buf BUF1 (N741, N736);
not NOT1 (N742, N728);
not NOT1 (N743, N740);
not NOT1 (N744, N705);
not NOT1 (N745, N734);
buf BUF1 (N746, N710);
or OR3 (N747, N746, N587, N717);
and AND2 (N748, N738, N308);
or OR3 (N749, N748, N712, N620);
xor XOR2 (N750, N745, N13);
and AND4 (N751, N749, N299, N273, N378);
or OR3 (N752, N743, N323, N395);
and AND3 (N753, N737, N76, N339);
nand NAND2 (N754, N735, N515);
xor XOR2 (N755, N739, N695);
or OR2 (N756, N755, N63);
nand NAND2 (N757, N741, N43);
nor NOR4 (N758, N753, N36, N479, N495);
nor NOR2 (N759, N757, N401);
nor NOR4 (N760, N742, N260, N357, N742);
buf BUF1 (N761, N754);
xor XOR2 (N762, N752, N63);
nand NAND4 (N763, N756, N588, N275, N547);
nand NAND2 (N764, N750, N461);
or OR2 (N765, N744, N386);
nor NOR4 (N766, N763, N534, N717, N431);
or OR2 (N767, N751, N151);
or OR2 (N768, N761, N533);
nand NAND3 (N769, N765, N246, N706);
or OR2 (N770, N758, N545);
xor XOR2 (N771, N766, N549);
or OR4 (N772, N768, N284, N302, N368);
nor NOR2 (N773, N770, N671);
or OR2 (N774, N769, N219);
not NOT1 (N775, N774);
buf BUF1 (N776, N775);
buf BUF1 (N777, N760);
nor NOR4 (N778, N771, N754, N709, N595);
buf BUF1 (N779, N762);
nand NAND3 (N780, N767, N700, N517);
not NOT1 (N781, N779);
nand NAND2 (N782, N772, N311);
not NOT1 (N783, N773);
nand NAND4 (N784, N781, N492, N658, N674);
buf BUF1 (N785, N783);
buf BUF1 (N786, N747);
and AND3 (N787, N785, N245, N568);
nand NAND2 (N788, N784, N62);
buf BUF1 (N789, N777);
and AND3 (N790, N778, N190, N329);
nand NAND2 (N791, N787, N173);
not NOT1 (N792, N764);
not NOT1 (N793, N790);
nand NAND4 (N794, N788, N54, N699, N780);
xor XOR2 (N795, N751, N338);
not NOT1 (N796, N794);
or OR4 (N797, N795, N546, N187, N413);
xor XOR2 (N798, N792, N315);
not NOT1 (N799, N789);
xor XOR2 (N800, N797, N159);
buf BUF1 (N801, N791);
buf BUF1 (N802, N759);
nor NOR4 (N803, N782, N410, N690, N688);
not NOT1 (N804, N786);
not NOT1 (N805, N776);
nor NOR3 (N806, N800, N795, N148);
not NOT1 (N807, N803);
nor NOR4 (N808, N807, N681, N622, N1);
and AND4 (N809, N805, N756, N30, N499);
buf BUF1 (N810, N808);
and AND2 (N811, N796, N470);
nand NAND2 (N812, N811, N593);
nand NAND3 (N813, N809, N112, N219);
buf BUF1 (N814, N812);
and AND4 (N815, N799, N512, N253, N481);
and AND4 (N816, N801, N414, N348, N308);
not NOT1 (N817, N814);
nor NOR2 (N818, N804, N217);
and AND2 (N819, N815, N648);
nor NOR4 (N820, N810, N488, N216, N780);
and AND3 (N821, N818, N594, N45);
not NOT1 (N822, N802);
or OR2 (N823, N820, N66);
not NOT1 (N824, N793);
nand NAND4 (N825, N817, N159, N671, N708);
and AND4 (N826, N798, N588, N302, N88);
and AND4 (N827, N819, N572, N294, N410);
or OR3 (N828, N827, N300, N410);
or OR4 (N829, N828, N125, N262, N207);
buf BUF1 (N830, N825);
or OR2 (N831, N822, N542);
not NOT1 (N832, N806);
nand NAND2 (N833, N832, N624);
and AND3 (N834, N823, N492, N776);
not NOT1 (N835, N824);
nor NOR2 (N836, N830, N153);
nand NAND3 (N837, N816, N674, N628);
buf BUF1 (N838, N834);
nor NOR2 (N839, N836, N101);
not NOT1 (N840, N826);
nor NOR3 (N841, N839, N213, N312);
nand NAND4 (N842, N838, N623, N791, N125);
nor NOR2 (N843, N842, N410);
nand NAND3 (N844, N841, N586, N605);
or OR2 (N845, N831, N438);
nand NAND4 (N846, N844, N234, N193, N499);
and AND3 (N847, N843, N223, N529);
or OR4 (N848, N840, N591, N155, N547);
nand NAND3 (N849, N835, N218, N728);
and AND2 (N850, N833, N656);
buf BUF1 (N851, N821);
nand NAND3 (N852, N850, N235, N668);
buf BUF1 (N853, N851);
nor NOR2 (N854, N847, N280);
xor XOR2 (N855, N829, N589);
or OR2 (N856, N849, N428);
xor XOR2 (N857, N856, N239);
xor XOR2 (N858, N852, N487);
and AND2 (N859, N854, N502);
buf BUF1 (N860, N845);
nand NAND2 (N861, N858, N735);
buf BUF1 (N862, N861);
xor XOR2 (N863, N857, N10);
nand NAND4 (N864, N853, N228, N643, N762);
not NOT1 (N865, N862);
nand NAND2 (N866, N863, N627);
or OR2 (N867, N848, N503);
nor NOR3 (N868, N864, N505, N677);
nor NOR4 (N869, N860, N112, N793, N89);
nor NOR4 (N870, N813, N856, N355, N516);
and AND4 (N871, N865, N833, N384, N484);
xor XOR2 (N872, N846, N507);
or OR2 (N873, N837, N607);
and AND2 (N874, N855, N786);
xor XOR2 (N875, N867, N871);
not NOT1 (N876, N739);
xor XOR2 (N877, N876, N336);
or OR2 (N878, N875, N152);
or OR3 (N879, N874, N455, N88);
and AND3 (N880, N866, N874, N401);
and AND2 (N881, N869, N342);
xor XOR2 (N882, N873, N541);
xor XOR2 (N883, N872, N439);
buf BUF1 (N884, N870);
nor NOR3 (N885, N859, N214, N409);
nand NAND3 (N886, N878, N822, N879);
xor XOR2 (N887, N74, N314);
not NOT1 (N888, N884);
nor NOR4 (N889, N880, N173, N411, N90);
not NOT1 (N890, N885);
nand NAND3 (N891, N881, N718, N866);
and AND2 (N892, N891, N231);
and AND3 (N893, N868, N824, N337);
xor XOR2 (N894, N893, N761);
xor XOR2 (N895, N882, N855);
and AND4 (N896, N888, N691, N223, N767);
or OR4 (N897, N877, N299, N129, N537);
or OR2 (N898, N883, N601);
xor XOR2 (N899, N887, N448);
or OR2 (N900, N889, N199);
or OR3 (N901, N900, N796, N288);
and AND3 (N902, N896, N267, N775);
nor NOR3 (N903, N901, N877, N225);
or OR3 (N904, N898, N245, N155);
nor NOR2 (N905, N903, N802);
buf BUF1 (N906, N892);
or OR3 (N907, N897, N598, N495);
nand NAND4 (N908, N894, N595, N254, N633);
or OR2 (N909, N899, N844);
xor XOR2 (N910, N890, N183);
and AND3 (N911, N910, N745, N573);
nor NOR2 (N912, N909, N398);
nor NOR3 (N913, N895, N730, N628);
xor XOR2 (N914, N907, N567);
or OR4 (N915, N914, N745, N261, N36);
buf BUF1 (N916, N912);
and AND2 (N917, N902, N454);
buf BUF1 (N918, N886);
buf BUF1 (N919, N918);
xor XOR2 (N920, N905, N851);
not NOT1 (N921, N906);
xor XOR2 (N922, N913, N596);
or OR3 (N923, N919, N630, N909);
xor XOR2 (N924, N904, N891);
nor NOR2 (N925, N911, N786);
nand NAND2 (N926, N922, N228);
nor NOR2 (N927, N917, N830);
and AND2 (N928, N927, N126);
and AND2 (N929, N915, N790);
nand NAND2 (N930, N923, N116);
nand NAND3 (N931, N928, N483, N599);
buf BUF1 (N932, N921);
buf BUF1 (N933, N930);
nand NAND4 (N934, N933, N348, N505, N446);
not NOT1 (N935, N934);
xor XOR2 (N936, N920, N859);
nor NOR2 (N937, N908, N619);
nand NAND2 (N938, N926, N477);
nand NAND3 (N939, N925, N799, N267);
xor XOR2 (N940, N929, N811);
or OR3 (N941, N940, N233, N841);
xor XOR2 (N942, N932, N140);
nand NAND4 (N943, N924, N634, N240, N208);
nand NAND3 (N944, N931, N670, N695);
nand NAND4 (N945, N941, N83, N761, N225);
buf BUF1 (N946, N945);
nand NAND4 (N947, N942, N653, N782, N500);
buf BUF1 (N948, N935);
xor XOR2 (N949, N948, N214);
nand NAND3 (N950, N916, N73, N122);
not NOT1 (N951, N939);
xor XOR2 (N952, N946, N681);
and AND3 (N953, N949, N437, N158);
or OR4 (N954, N938, N689, N531, N186);
nand NAND3 (N955, N953, N837, N679);
nand NAND3 (N956, N943, N764, N32);
nor NOR2 (N957, N936, N539);
buf BUF1 (N958, N950);
nor NOR3 (N959, N957, N700, N508);
xor XOR2 (N960, N947, N329);
xor XOR2 (N961, N937, N947);
nor NOR3 (N962, N961, N302, N72);
buf BUF1 (N963, N960);
nor NOR2 (N964, N952, N729);
nor NOR4 (N965, N944, N867, N741, N431);
buf BUF1 (N966, N954);
not NOT1 (N967, N964);
nor NOR2 (N968, N958, N242);
or OR3 (N969, N968, N923, N390);
nand NAND4 (N970, N963, N838, N48, N524);
xor XOR2 (N971, N967, N670);
nor NOR2 (N972, N965, N836);
xor XOR2 (N973, N955, N870);
nor NOR3 (N974, N959, N530, N49);
nand NAND2 (N975, N974, N473);
and AND2 (N976, N969, N210);
buf BUF1 (N977, N970);
buf BUF1 (N978, N951);
nor NOR2 (N979, N972, N330);
and AND4 (N980, N978, N745, N200, N498);
nand NAND3 (N981, N971, N403, N5);
or OR3 (N982, N975, N959, N234);
or OR3 (N983, N962, N263, N490);
nor NOR2 (N984, N979, N847);
nor NOR2 (N985, N977, N841);
nor NOR4 (N986, N980, N124, N619, N853);
or OR3 (N987, N966, N439, N469);
or OR4 (N988, N987, N461, N396, N434);
nor NOR3 (N989, N976, N339, N950);
or OR3 (N990, N956, N93, N102);
nand NAND2 (N991, N985, N755);
nand NAND2 (N992, N991, N697);
or OR4 (N993, N992, N939, N971, N46);
not NOT1 (N994, N986);
nand NAND2 (N995, N984, N950);
nor NOR3 (N996, N983, N753, N639);
nor NOR4 (N997, N993, N303, N683, N246);
or OR3 (N998, N995, N742, N5);
xor XOR2 (N999, N990, N21);
and AND2 (N1000, N973, N150);
nand NAND3 (N1001, N998, N726, N77);
and AND3 (N1002, N996, N191, N684);
and AND2 (N1003, N994, N359);
xor XOR2 (N1004, N988, N986);
or OR4 (N1005, N981, N355, N420, N313);
buf BUF1 (N1006, N1005);
buf BUF1 (N1007, N1001);
xor XOR2 (N1008, N1002, N663);
nand NAND4 (N1009, N1000, N502, N526, N44);
xor XOR2 (N1010, N1003, N851);
and AND4 (N1011, N1009, N1007, N237, N923);
nand NAND4 (N1012, N902, N727, N353, N939);
and AND2 (N1013, N1006, N186);
not NOT1 (N1014, N1011);
not NOT1 (N1015, N1014);
and AND2 (N1016, N997, N688);
xor XOR2 (N1017, N1013, N560);
not NOT1 (N1018, N982);
not NOT1 (N1019, N1010);
and AND4 (N1020, N1018, N195, N285, N762);
or OR3 (N1021, N1004, N384, N982);
and AND3 (N1022, N989, N145, N603);
xor XOR2 (N1023, N1008, N927);
not NOT1 (N1024, N1012);
or OR3 (N1025, N1016, N52, N324);
nor NOR3 (N1026, N1017, N717, N318);
buf BUF1 (N1027, N1023);
or OR3 (N1028, N1022, N64, N624);
nand NAND4 (N1029, N1026, N372, N256, N923);
and AND2 (N1030, N1020, N447);
nand NAND3 (N1031, N1027, N908, N233);
not NOT1 (N1032, N1029);
buf BUF1 (N1033, N1019);
or OR3 (N1034, N1033, N346, N467);
xor XOR2 (N1035, N1030, N202);
buf BUF1 (N1036, N1035);
or OR2 (N1037, N1028, N988);
buf BUF1 (N1038, N999);
or OR3 (N1039, N1036, N277, N13);
xor XOR2 (N1040, N1037, N373);
buf BUF1 (N1041, N1040);
or OR3 (N1042, N1039, N964, N244);
and AND4 (N1043, N1038, N861, N301, N904);
nand NAND2 (N1044, N1032, N229);
and AND4 (N1045, N1044, N762, N801, N646);
and AND4 (N1046, N1031, N285, N104, N711);
buf BUF1 (N1047, N1024);
xor XOR2 (N1048, N1043, N579);
not NOT1 (N1049, N1046);
buf BUF1 (N1050, N1021);
nor NOR2 (N1051, N1041, N410);
not NOT1 (N1052, N1047);
or OR2 (N1053, N1050, N308);
not NOT1 (N1054, N1049);
not NOT1 (N1055, N1015);
nand NAND3 (N1056, N1055, N273, N324);
and AND3 (N1057, N1056, N270, N24);
or OR2 (N1058, N1045, N895);
buf BUF1 (N1059, N1052);
buf BUF1 (N1060, N1048);
xor XOR2 (N1061, N1058, N803);
xor XOR2 (N1062, N1059, N435);
or OR4 (N1063, N1051, N105, N1009, N776);
and AND2 (N1064, N1061, N960);
or OR2 (N1065, N1063, N810);
or OR2 (N1066, N1057, N452);
xor XOR2 (N1067, N1053, N808);
xor XOR2 (N1068, N1065, N185);
or OR2 (N1069, N1067, N340);
xor XOR2 (N1070, N1066, N180);
xor XOR2 (N1071, N1042, N372);
not NOT1 (N1072, N1062);
and AND2 (N1073, N1068, N314);
xor XOR2 (N1074, N1071, N998);
not NOT1 (N1075, N1072);
nand NAND4 (N1076, N1034, N716, N640, N297);
and AND3 (N1077, N1069, N643, N426);
not NOT1 (N1078, N1073);
not NOT1 (N1079, N1076);
buf BUF1 (N1080, N1070);
buf BUF1 (N1081, N1079);
not NOT1 (N1082, N1054);
nand NAND4 (N1083, N1080, N410, N176, N650);
nor NOR4 (N1084, N1025, N254, N380, N802);
xor XOR2 (N1085, N1082, N495);
nand NAND4 (N1086, N1083, N445, N316, N349);
nand NAND4 (N1087, N1077, N194, N297, N458);
not NOT1 (N1088, N1064);
xor XOR2 (N1089, N1087, N792);
buf BUF1 (N1090, N1074);
buf BUF1 (N1091, N1060);
buf BUF1 (N1092, N1088);
nand NAND4 (N1093, N1091, N650, N357, N1077);
buf BUF1 (N1094, N1081);
xor XOR2 (N1095, N1078, N13);
nor NOR4 (N1096, N1090, N166, N944, N171);
or OR3 (N1097, N1075, N113, N980);
nor NOR3 (N1098, N1086, N1049, N1043);
buf BUF1 (N1099, N1097);
nand NAND2 (N1100, N1096, N731);
nor NOR4 (N1101, N1092, N502, N851, N366);
nor NOR4 (N1102, N1099, N57, N255, N759);
not NOT1 (N1103, N1093);
nand NAND4 (N1104, N1102, N175, N837, N703);
nor NOR3 (N1105, N1094, N683, N1038);
and AND4 (N1106, N1098, N242, N157, N740);
not NOT1 (N1107, N1085);
buf BUF1 (N1108, N1103);
nor NOR3 (N1109, N1105, N54, N28);
buf BUF1 (N1110, N1084);
xor XOR2 (N1111, N1095, N224);
not NOT1 (N1112, N1107);
nor NOR4 (N1113, N1112, N1092, N738, N825);
xor XOR2 (N1114, N1101, N125);
xor XOR2 (N1115, N1109, N969);
or OR3 (N1116, N1108, N267, N797);
nor NOR4 (N1117, N1115, N780, N467, N983);
nor NOR2 (N1118, N1110, N479);
and AND3 (N1119, N1106, N555, N941);
not NOT1 (N1120, N1118);
nand NAND3 (N1121, N1111, N1005, N386);
not NOT1 (N1122, N1117);
or OR4 (N1123, N1121, N654, N969, N160);
buf BUF1 (N1124, N1123);
buf BUF1 (N1125, N1122);
nor NOR2 (N1126, N1113, N921);
or OR2 (N1127, N1120, N656);
and AND2 (N1128, N1126, N355);
not NOT1 (N1129, N1124);
or OR2 (N1130, N1104, N604);
nor NOR3 (N1131, N1089, N817, N515);
not NOT1 (N1132, N1116);
xor XOR2 (N1133, N1125, N727);
xor XOR2 (N1134, N1119, N543);
xor XOR2 (N1135, N1100, N122);
xor XOR2 (N1136, N1134, N71);
nand NAND4 (N1137, N1127, N618, N334, N798);
nor NOR2 (N1138, N1129, N272);
xor XOR2 (N1139, N1135, N66);
buf BUF1 (N1140, N1114);
buf BUF1 (N1141, N1137);
nor NOR4 (N1142, N1132, N638, N882, N1074);
or OR2 (N1143, N1142, N862);
or OR3 (N1144, N1128, N609, N351);
xor XOR2 (N1145, N1144, N619);
or OR3 (N1146, N1145, N726, N359);
xor XOR2 (N1147, N1131, N587);
nor NOR2 (N1148, N1130, N769);
buf BUF1 (N1149, N1133);
not NOT1 (N1150, N1146);
nand NAND3 (N1151, N1138, N1059, N271);
not NOT1 (N1152, N1150);
nand NAND4 (N1153, N1139, N531, N478, N570);
nor NOR3 (N1154, N1143, N573, N44);
or OR4 (N1155, N1154, N447, N767, N350);
buf BUF1 (N1156, N1140);
not NOT1 (N1157, N1148);
not NOT1 (N1158, N1152);
nand NAND2 (N1159, N1155, N880);
or OR2 (N1160, N1153, N462);
xor XOR2 (N1161, N1158, N935);
and AND3 (N1162, N1136, N968, N1150);
or OR2 (N1163, N1157, N724);
buf BUF1 (N1164, N1149);
nor NOR3 (N1165, N1161, N1064, N538);
buf BUF1 (N1166, N1156);
nand NAND4 (N1167, N1166, N62, N740, N344);
nand NAND2 (N1168, N1151, N589);
and AND2 (N1169, N1168, N617);
xor XOR2 (N1170, N1160, N59);
or OR3 (N1171, N1141, N1108, N18);
or OR2 (N1172, N1147, N265);
nor NOR3 (N1173, N1162, N399, N580);
and AND2 (N1174, N1172, N833);
not NOT1 (N1175, N1169);
or OR2 (N1176, N1159, N501);
or OR4 (N1177, N1164, N1059, N933, N741);
or OR2 (N1178, N1174, N1061);
nor NOR3 (N1179, N1176, N916, N580);
nand NAND2 (N1180, N1175, N880);
buf BUF1 (N1181, N1173);
and AND4 (N1182, N1178, N874, N599, N190);
xor XOR2 (N1183, N1180, N816);
buf BUF1 (N1184, N1165);
xor XOR2 (N1185, N1171, N130);
buf BUF1 (N1186, N1167);
not NOT1 (N1187, N1177);
or OR3 (N1188, N1183, N101, N840);
xor XOR2 (N1189, N1170, N688);
xor XOR2 (N1190, N1185, N734);
nor NOR2 (N1191, N1186, N310);
not NOT1 (N1192, N1179);
or OR3 (N1193, N1188, N993, N257);
nor NOR2 (N1194, N1191, N566);
buf BUF1 (N1195, N1184);
not NOT1 (N1196, N1194);
buf BUF1 (N1197, N1187);
buf BUF1 (N1198, N1163);
or OR2 (N1199, N1182, N1052);
xor XOR2 (N1200, N1189, N534);
buf BUF1 (N1201, N1193);
and AND3 (N1202, N1200, N627, N254);
nand NAND2 (N1203, N1202, N906);
nor NOR2 (N1204, N1203, N1159);
buf BUF1 (N1205, N1195);
nand NAND3 (N1206, N1199, N169, N1169);
and AND2 (N1207, N1197, N414);
buf BUF1 (N1208, N1198);
buf BUF1 (N1209, N1192);
nor NOR3 (N1210, N1207, N686, N110);
buf BUF1 (N1211, N1210);
or OR4 (N1212, N1205, N673, N28, N702);
and AND2 (N1213, N1181, N1120);
xor XOR2 (N1214, N1196, N916);
nand NAND4 (N1215, N1212, N142, N699, N88);
and AND2 (N1216, N1204, N715);
not NOT1 (N1217, N1190);
nand NAND2 (N1218, N1217, N818);
or OR4 (N1219, N1208, N982, N595, N686);
nand NAND2 (N1220, N1211, N658);
not NOT1 (N1221, N1209);
nor NOR2 (N1222, N1220, N691);
xor XOR2 (N1223, N1206, N96);
or OR3 (N1224, N1221, N1179, N382);
nor NOR3 (N1225, N1213, N946, N1099);
xor XOR2 (N1226, N1223, N542);
and AND4 (N1227, N1218, N455, N446, N1014);
buf BUF1 (N1228, N1214);
and AND2 (N1229, N1216, N297);
xor XOR2 (N1230, N1219, N141);
not NOT1 (N1231, N1201);
not NOT1 (N1232, N1228);
not NOT1 (N1233, N1224);
not NOT1 (N1234, N1230);
nand NAND2 (N1235, N1233, N888);
and AND2 (N1236, N1229, N298);
and AND4 (N1237, N1226, N1140, N1199, N266);
nor NOR4 (N1238, N1231, N1133, N1137, N368);
and AND4 (N1239, N1238, N824, N220, N1115);
xor XOR2 (N1240, N1232, N705);
nor NOR2 (N1241, N1225, N840);
not NOT1 (N1242, N1241);
nor NOR2 (N1243, N1240, N186);
xor XOR2 (N1244, N1222, N520);
not NOT1 (N1245, N1243);
and AND4 (N1246, N1244, N205, N799, N273);
nand NAND3 (N1247, N1237, N497, N610);
not NOT1 (N1248, N1245);
nor NOR3 (N1249, N1247, N629, N227);
nand NAND2 (N1250, N1234, N588);
buf BUF1 (N1251, N1246);
nand NAND4 (N1252, N1236, N520, N441, N1127);
and AND2 (N1253, N1251, N862);
buf BUF1 (N1254, N1242);
or OR4 (N1255, N1239, N553, N731, N1039);
xor XOR2 (N1256, N1250, N1035);
xor XOR2 (N1257, N1253, N122);
and AND4 (N1258, N1249, N537, N525, N700);
and AND3 (N1259, N1227, N900, N1109);
and AND2 (N1260, N1259, N338);
and AND3 (N1261, N1255, N957, N668);
not NOT1 (N1262, N1235);
or OR4 (N1263, N1260, N670, N1074, N1256);
nor NOR4 (N1264, N19, N769, N1244, N983);
buf BUF1 (N1265, N1248);
xor XOR2 (N1266, N1215, N336);
nand NAND2 (N1267, N1264, N908);
or OR3 (N1268, N1257, N1023, N202);
buf BUF1 (N1269, N1261);
xor XOR2 (N1270, N1266, N807);
xor XOR2 (N1271, N1268, N530);
or OR3 (N1272, N1269, N720, N1253);
or OR2 (N1273, N1254, N896);
not NOT1 (N1274, N1271);
nand NAND4 (N1275, N1262, N867, N914, N953);
and AND3 (N1276, N1275, N1133, N1131);
buf BUF1 (N1277, N1276);
not NOT1 (N1278, N1263);
and AND3 (N1279, N1258, N145, N960);
or OR4 (N1280, N1277, N612, N1051, N1056);
nand NAND3 (N1281, N1274, N1017, N311);
and AND4 (N1282, N1272, N507, N426, N165);
not NOT1 (N1283, N1281);
nor NOR3 (N1284, N1265, N1094, N14);
nor NOR4 (N1285, N1273, N1058, N829, N8);
buf BUF1 (N1286, N1282);
and AND2 (N1287, N1278, N647);
xor XOR2 (N1288, N1279, N306);
and AND3 (N1289, N1267, N704, N1162);
nor NOR3 (N1290, N1287, N1212, N821);
buf BUF1 (N1291, N1280);
nand NAND3 (N1292, N1285, N562, N333);
and AND4 (N1293, N1288, N1207, N792, N67);
xor XOR2 (N1294, N1283, N919);
nor NOR2 (N1295, N1252, N587);
not NOT1 (N1296, N1284);
nor NOR2 (N1297, N1292, N867);
xor XOR2 (N1298, N1270, N1166);
xor XOR2 (N1299, N1293, N669);
nand NAND3 (N1300, N1299, N225, N997);
or OR3 (N1301, N1290, N1232, N1084);
xor XOR2 (N1302, N1295, N439);
nand NAND3 (N1303, N1300, N129, N1087);
or OR3 (N1304, N1301, N1272, N82);
xor XOR2 (N1305, N1294, N650);
or OR4 (N1306, N1296, N1064, N1296, N75);
and AND4 (N1307, N1291, N582, N685, N485);
nor NOR4 (N1308, N1289, N313, N425, N1279);
buf BUF1 (N1309, N1307);
nor NOR2 (N1310, N1297, N85);
nand NAND4 (N1311, N1304, N841, N509, N984);
buf BUF1 (N1312, N1302);
not NOT1 (N1313, N1310);
buf BUF1 (N1314, N1308);
not NOT1 (N1315, N1303);
xor XOR2 (N1316, N1312, N870);
or OR2 (N1317, N1286, N253);
xor XOR2 (N1318, N1315, N256);
and AND4 (N1319, N1306, N341, N1096, N79);
nand NAND2 (N1320, N1318, N685);
xor XOR2 (N1321, N1317, N926);
nand NAND4 (N1322, N1321, N874, N281, N346);
and AND3 (N1323, N1316, N1192, N295);
xor XOR2 (N1324, N1322, N653);
or OR2 (N1325, N1324, N1186);
or OR2 (N1326, N1325, N402);
or OR4 (N1327, N1305, N252, N846, N148);
not NOT1 (N1328, N1323);
buf BUF1 (N1329, N1314);
not NOT1 (N1330, N1298);
not NOT1 (N1331, N1326);
or OR2 (N1332, N1309, N76);
buf BUF1 (N1333, N1328);
xor XOR2 (N1334, N1313, N1004);
and AND4 (N1335, N1333, N1232, N531, N1220);
or OR2 (N1336, N1335, N362);
or OR4 (N1337, N1320, N1234, N1075, N938);
xor XOR2 (N1338, N1337, N1083);
nor NOR4 (N1339, N1319, N1062, N166, N149);
and AND2 (N1340, N1338, N149);
not NOT1 (N1341, N1340);
nor NOR4 (N1342, N1336, N571, N1251, N1196);
not NOT1 (N1343, N1332);
nand NAND4 (N1344, N1343, N731, N778, N235);
or OR4 (N1345, N1327, N103, N992, N11);
buf BUF1 (N1346, N1345);
nor NOR2 (N1347, N1342, N352);
or OR4 (N1348, N1329, N40, N862, N835);
nor NOR3 (N1349, N1339, N398, N716);
nor NOR4 (N1350, N1348, N300, N1057, N318);
nor NOR4 (N1351, N1341, N509, N111, N9);
nand NAND3 (N1352, N1347, N1087, N443);
nand NAND4 (N1353, N1311, N1257, N487, N738);
nor NOR3 (N1354, N1352, N1124, N298);
not NOT1 (N1355, N1349);
or OR4 (N1356, N1334, N890, N410, N1166);
nand NAND3 (N1357, N1351, N1219, N298);
and AND2 (N1358, N1350, N349);
xor XOR2 (N1359, N1353, N879);
and AND2 (N1360, N1344, N169);
nand NAND3 (N1361, N1346, N924, N369);
not NOT1 (N1362, N1359);
nor NOR2 (N1363, N1358, N725);
or OR4 (N1364, N1361, N157, N934, N1156);
nand NAND3 (N1365, N1356, N578, N643);
or OR2 (N1366, N1355, N69);
buf BUF1 (N1367, N1362);
or OR3 (N1368, N1357, N601, N1025);
not NOT1 (N1369, N1354);
and AND2 (N1370, N1364, N842);
not NOT1 (N1371, N1363);
not NOT1 (N1372, N1371);
xor XOR2 (N1373, N1372, N858);
nor NOR2 (N1374, N1369, N335);
nor NOR4 (N1375, N1366, N368, N1170, N621);
or OR4 (N1376, N1331, N1032, N1105, N1214);
buf BUF1 (N1377, N1367);
or OR3 (N1378, N1376, N1069, N691);
buf BUF1 (N1379, N1368);
nor NOR2 (N1380, N1360, N170);
buf BUF1 (N1381, N1377);
nor NOR3 (N1382, N1365, N321, N1250);
nor NOR4 (N1383, N1382, N1238, N433, N1061);
or OR2 (N1384, N1330, N485);
buf BUF1 (N1385, N1373);
and AND4 (N1386, N1385, N365, N1104, N95);
xor XOR2 (N1387, N1370, N763);
buf BUF1 (N1388, N1383);
xor XOR2 (N1389, N1381, N637);
buf BUF1 (N1390, N1386);
buf BUF1 (N1391, N1388);
nand NAND3 (N1392, N1389, N968, N390);
not NOT1 (N1393, N1378);
nand NAND2 (N1394, N1390, N64);
or OR2 (N1395, N1380, N520);
nand NAND3 (N1396, N1391, N264, N380);
xor XOR2 (N1397, N1374, N1376);
and AND2 (N1398, N1397, N797);
and AND4 (N1399, N1392, N1071, N1347, N837);
or OR2 (N1400, N1395, N1057);
and AND3 (N1401, N1398, N966, N648);
and AND4 (N1402, N1399, N1361, N891, N1117);
not NOT1 (N1403, N1375);
nand NAND2 (N1404, N1401, N870);
nand NAND4 (N1405, N1402, N568, N962, N574);
nand NAND2 (N1406, N1379, N574);
not NOT1 (N1407, N1394);
and AND3 (N1408, N1387, N168, N166);
or OR4 (N1409, N1404, N246, N632, N469);
or OR3 (N1410, N1396, N814, N522);
not NOT1 (N1411, N1408);
not NOT1 (N1412, N1411);
nand NAND3 (N1413, N1403, N14, N1051);
nand NAND2 (N1414, N1407, N596);
not NOT1 (N1415, N1400);
buf BUF1 (N1416, N1384);
or OR3 (N1417, N1412, N10, N542);
not NOT1 (N1418, N1414);
nand NAND4 (N1419, N1415, N1141, N1133, N89);
xor XOR2 (N1420, N1417, N1389);
xor XOR2 (N1421, N1418, N36);
not NOT1 (N1422, N1419);
buf BUF1 (N1423, N1405);
not NOT1 (N1424, N1421);
nand NAND4 (N1425, N1422, N600, N15, N678);
xor XOR2 (N1426, N1393, N1312);
nor NOR3 (N1427, N1426, N994, N1060);
or OR4 (N1428, N1420, N1281, N897, N263);
and AND4 (N1429, N1425, N459, N605, N828);
or OR4 (N1430, N1416, N740, N1139, N565);
nand NAND4 (N1431, N1406, N822, N672, N921);
and AND2 (N1432, N1413, N1403);
nand NAND3 (N1433, N1431, N718, N57);
and AND3 (N1434, N1430, N134, N495);
xor XOR2 (N1435, N1428, N1073);
or OR3 (N1436, N1434, N78, N54);
nand NAND2 (N1437, N1432, N103);
and AND2 (N1438, N1423, N285);
not NOT1 (N1439, N1437);
xor XOR2 (N1440, N1427, N472);
or OR2 (N1441, N1440, N1054);
xor XOR2 (N1442, N1435, N1089);
nand NAND3 (N1443, N1409, N182, N1096);
not NOT1 (N1444, N1433);
and AND4 (N1445, N1444, N469, N863, N561);
and AND4 (N1446, N1445, N1099, N481, N604);
or OR4 (N1447, N1436, N1164, N176, N1367);
xor XOR2 (N1448, N1439, N1440);
xor XOR2 (N1449, N1442, N442);
and AND3 (N1450, N1446, N745, N1284);
buf BUF1 (N1451, N1448);
not NOT1 (N1452, N1447);
nand NAND2 (N1453, N1451, N647);
and AND4 (N1454, N1443, N763, N512, N491);
nor NOR4 (N1455, N1410, N577, N211, N536);
xor XOR2 (N1456, N1454, N1036);
and AND2 (N1457, N1456, N626);
and AND2 (N1458, N1455, N138);
nand NAND4 (N1459, N1438, N249, N1152, N705);
xor XOR2 (N1460, N1424, N1244);
xor XOR2 (N1461, N1453, N1333);
not NOT1 (N1462, N1457);
xor XOR2 (N1463, N1462, N345);
nor NOR4 (N1464, N1463, N332, N301, N1034);
or OR3 (N1465, N1441, N778, N949);
nor NOR3 (N1466, N1464, N1367, N240);
buf BUF1 (N1467, N1449);
or OR4 (N1468, N1465, N86, N1032, N329);
and AND3 (N1469, N1467, N73, N628);
nand NAND2 (N1470, N1429, N270);
nor NOR2 (N1471, N1461, N1155);
buf BUF1 (N1472, N1470);
nor NOR4 (N1473, N1468, N85, N928, N397);
xor XOR2 (N1474, N1473, N18);
xor XOR2 (N1475, N1459, N966);
nor NOR4 (N1476, N1471, N518, N500, N84);
nand NAND2 (N1477, N1450, N1052);
xor XOR2 (N1478, N1466, N1209);
buf BUF1 (N1479, N1474);
nand NAND4 (N1480, N1475, N552, N124, N1155);
not NOT1 (N1481, N1472);
buf BUF1 (N1482, N1479);
nand NAND2 (N1483, N1482, N1467);
buf BUF1 (N1484, N1483);
not NOT1 (N1485, N1478);
and AND3 (N1486, N1485, N1018, N1037);
or OR3 (N1487, N1460, N693, N325);
buf BUF1 (N1488, N1469);
nand NAND2 (N1489, N1476, N1111);
nor NOR2 (N1490, N1481, N1104);
nor NOR3 (N1491, N1487, N1176, N504);
and AND3 (N1492, N1489, N560, N101);
buf BUF1 (N1493, N1458);
buf BUF1 (N1494, N1480);
buf BUF1 (N1495, N1452);
nand NAND3 (N1496, N1492, N315, N407);
buf BUF1 (N1497, N1477);
not NOT1 (N1498, N1493);
or OR2 (N1499, N1494, N900);
nand NAND4 (N1500, N1484, N357, N17, N656);
nor NOR3 (N1501, N1491, N226, N439);
nand NAND4 (N1502, N1500, N890, N506, N969);
or OR2 (N1503, N1502, N734);
buf BUF1 (N1504, N1490);
not NOT1 (N1505, N1488);
not NOT1 (N1506, N1486);
and AND3 (N1507, N1499, N96, N1219);
not NOT1 (N1508, N1496);
and AND3 (N1509, N1506, N226, N785);
or OR2 (N1510, N1495, N1011);
nand NAND3 (N1511, N1497, N449, N137);
and AND3 (N1512, N1509, N566, N1057);
buf BUF1 (N1513, N1503);
and AND3 (N1514, N1511, N960, N403);
nor NOR4 (N1515, N1513, N357, N295, N175);
or OR3 (N1516, N1510, N284, N550);
and AND3 (N1517, N1501, N368, N905);
buf BUF1 (N1518, N1507);
nand NAND3 (N1519, N1517, N1241, N63);
not NOT1 (N1520, N1515);
buf BUF1 (N1521, N1498);
endmodule