// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13;

output N3503,N3504,N3506,N3508,N3511,N3512,N3500,N3507,N3485,N3513;

or OR3 (N14, N9, N7, N3);
buf BUF1 (N15, N1);
and AND3 (N16, N15, N12, N2);
nor NOR2 (N17, N15, N8);
or OR3 (N18, N11, N10, N17);
xor XOR2 (N19, N17, N13);
and AND4 (N20, N11, N8, N12, N11);
or OR2 (N21, N20, N17);
nor NOR4 (N22, N8, N10, N2, N7);
not NOT1 (N23, N1);
not NOT1 (N24, N3);
and AND2 (N25, N10, N9);
buf BUF1 (N26, N2);
nor NOR2 (N27, N14, N5);
nand NAND3 (N28, N27, N20, N20);
nor NOR4 (N29, N18, N15, N28, N21);
buf BUF1 (N30, N8);
not NOT1 (N31, N27);
xor XOR2 (N32, N23, N2);
or OR3 (N33, N26, N23, N32);
not NOT1 (N34, N18);
not NOT1 (N35, N24);
and AND3 (N36, N22, N19, N24);
xor XOR2 (N37, N21, N2);
nand NAND3 (N38, N29, N16, N33);
and AND2 (N39, N1, N22);
not NOT1 (N40, N25);
nor NOR3 (N41, N38, N32, N15);
nand NAND4 (N42, N13, N26, N18, N9);
nor NOR2 (N43, N40, N11);
buf BUF1 (N44, N41);
xor XOR2 (N45, N30, N27);
buf BUF1 (N46, N39);
nor NOR2 (N47, N31, N40);
not NOT1 (N48, N44);
not NOT1 (N49, N48);
buf BUF1 (N50, N46);
nor NOR4 (N51, N43, N22, N7, N39);
nor NOR2 (N52, N42, N20);
xor XOR2 (N53, N49, N12);
xor XOR2 (N54, N45, N31);
and AND4 (N55, N34, N41, N51, N43);
nor NOR2 (N56, N38, N33);
xor XOR2 (N57, N55, N19);
or OR3 (N58, N52, N5, N40);
and AND4 (N59, N50, N26, N22, N43);
nand NAND4 (N60, N36, N36, N53, N18);
xor XOR2 (N61, N42, N56);
xor XOR2 (N62, N57, N10);
buf BUF1 (N63, N27);
or OR2 (N64, N60, N36);
xor XOR2 (N65, N64, N56);
buf BUF1 (N66, N35);
nand NAND2 (N67, N59, N57);
nand NAND3 (N68, N54, N52, N64);
buf BUF1 (N69, N62);
or OR3 (N70, N68, N62, N67);
and AND2 (N71, N41, N13);
nor NOR3 (N72, N66, N68, N11);
nand NAND4 (N73, N61, N26, N35, N35);
xor XOR2 (N74, N73, N10);
and AND4 (N75, N72, N67, N51, N8);
and AND2 (N76, N37, N18);
xor XOR2 (N77, N63, N70);
or OR4 (N78, N38, N1, N30, N60);
nor NOR4 (N79, N76, N6, N30, N21);
xor XOR2 (N80, N74, N79);
nor NOR2 (N81, N76, N14);
xor XOR2 (N82, N80, N57);
or OR4 (N83, N47, N34, N47, N50);
buf BUF1 (N84, N58);
or OR3 (N85, N84, N31, N14);
not NOT1 (N86, N69);
nor NOR3 (N87, N78, N86, N17);
or OR3 (N88, N73, N30, N74);
xor XOR2 (N89, N77, N14);
nand NAND4 (N90, N83, N70, N68, N75);
not NOT1 (N91, N75);
and AND4 (N92, N90, N73, N46, N12);
and AND3 (N93, N89, N11, N28);
and AND2 (N94, N85, N62);
or OR2 (N95, N82, N39);
or OR3 (N96, N94, N72, N11);
not NOT1 (N97, N87);
xor XOR2 (N98, N81, N83);
nor NOR4 (N99, N96, N27, N30, N54);
or OR4 (N100, N88, N38, N29, N5);
nor NOR4 (N101, N99, N68, N70, N57);
and AND2 (N102, N100, N7);
nand NAND4 (N103, N71, N17, N92, N71);
nor NOR2 (N104, N94, N37);
or OR2 (N105, N65, N92);
nor NOR2 (N106, N103, N99);
buf BUF1 (N107, N101);
buf BUF1 (N108, N98);
not NOT1 (N109, N91);
nand NAND4 (N110, N107, N84, N99, N13);
not NOT1 (N111, N97);
nor NOR4 (N112, N109, N100, N72, N66);
nand NAND3 (N113, N108, N57, N95);
nor NOR4 (N114, N104, N62, N112, N25);
and AND4 (N115, N52, N87, N40, N96);
xor XOR2 (N116, N74, N41);
nand NAND2 (N117, N105, N96);
or OR4 (N118, N116, N88, N57, N25);
not NOT1 (N119, N102);
buf BUF1 (N120, N93);
and AND2 (N121, N115, N100);
and AND2 (N122, N119, N102);
not NOT1 (N123, N118);
or OR4 (N124, N113, N3, N82, N65);
xor XOR2 (N125, N124, N92);
nor NOR4 (N126, N110, N43, N89, N107);
buf BUF1 (N127, N123);
nand NAND4 (N128, N125, N13, N70, N1);
nand NAND2 (N129, N120, N52);
buf BUF1 (N130, N111);
nor NOR3 (N131, N122, N39, N83);
and AND2 (N132, N117, N44);
or OR3 (N133, N129, N122, N19);
or OR3 (N134, N114, N69, N58);
nand NAND3 (N135, N106, N30, N1);
and AND2 (N136, N135, N40);
buf BUF1 (N137, N121);
xor XOR2 (N138, N134, N7);
and AND4 (N139, N128, N63, N134, N127);
not NOT1 (N140, N134);
and AND3 (N141, N136, N119, N38);
buf BUF1 (N142, N138);
or OR4 (N143, N131, N8, N12, N91);
buf BUF1 (N144, N143);
not NOT1 (N145, N133);
not NOT1 (N146, N139);
or OR2 (N147, N137, N14);
xor XOR2 (N148, N141, N48);
and AND2 (N149, N145, N146);
or OR3 (N150, N22, N144, N136);
not NOT1 (N151, N148);
and AND3 (N152, N35, N122, N98);
nor NOR3 (N153, N140, N43, N18);
or OR4 (N154, N132, N30, N150, N82);
nand NAND3 (N155, N118, N44, N50);
or OR3 (N156, N151, N131, N132);
nand NAND2 (N157, N155, N156);
not NOT1 (N158, N123);
nand NAND2 (N159, N130, N38);
nor NOR2 (N160, N158, N19);
nand NAND3 (N161, N157, N33, N63);
nand NAND4 (N162, N153, N126, N83, N71);
xor XOR2 (N163, N20, N30);
and AND3 (N164, N154, N155, N16);
nand NAND4 (N165, N152, N122, N130, N5);
or OR2 (N166, N149, N60);
or OR3 (N167, N159, N152, N166);
nand NAND4 (N168, N6, N74, N130, N138);
buf BUF1 (N169, N142);
not NOT1 (N170, N165);
xor XOR2 (N171, N168, N147);
nand NAND2 (N172, N96, N99);
and AND3 (N173, N163, N59, N40);
xor XOR2 (N174, N162, N87);
or OR2 (N175, N169, N50);
or OR4 (N176, N173, N71, N139, N84);
xor XOR2 (N177, N172, N6);
buf BUF1 (N178, N170);
or OR3 (N179, N167, N112, N84);
buf BUF1 (N180, N164);
nand NAND4 (N181, N179, N78, N53, N94);
and AND2 (N182, N174, N39);
nand NAND4 (N183, N180, N106, N44, N143);
not NOT1 (N184, N160);
buf BUF1 (N185, N181);
nor NOR3 (N186, N171, N140, N29);
nor NOR3 (N187, N177, N78, N90);
and AND2 (N188, N186, N35);
xor XOR2 (N189, N183, N64);
buf BUF1 (N190, N176);
xor XOR2 (N191, N178, N178);
nor NOR4 (N192, N175, N172, N66, N12);
not NOT1 (N193, N189);
not NOT1 (N194, N187);
buf BUF1 (N195, N188);
nand NAND4 (N196, N161, N19, N109, N146);
nand NAND3 (N197, N191, N73, N92);
nor NOR4 (N198, N193, N11, N165, N45);
and AND3 (N199, N198, N133, N190);
or OR3 (N200, N128, N7, N174);
nor NOR4 (N201, N185, N67, N63, N149);
nor NOR2 (N202, N182, N64);
or OR4 (N203, N195, N18, N90, N133);
nor NOR3 (N204, N184, N18, N58);
and AND4 (N205, N199, N105, N39, N49);
nand NAND4 (N206, N192, N186, N6, N149);
buf BUF1 (N207, N204);
or OR2 (N208, N201, N82);
and AND4 (N209, N202, N66, N194, N143);
xor XOR2 (N210, N189, N151);
buf BUF1 (N211, N205);
xor XOR2 (N212, N207, N188);
nor NOR2 (N213, N206, N56);
nor NOR2 (N214, N211, N180);
buf BUF1 (N215, N213);
buf BUF1 (N216, N196);
not NOT1 (N217, N209);
buf BUF1 (N218, N200);
or OR3 (N219, N214, N207, N45);
and AND4 (N220, N210, N53, N2, N127);
and AND2 (N221, N216, N186);
buf BUF1 (N222, N219);
not NOT1 (N223, N218);
nor NOR2 (N224, N203, N50);
nand NAND4 (N225, N208, N180, N15, N46);
nand NAND4 (N226, N224, N157, N42, N112);
nor NOR3 (N227, N222, N6, N103);
buf BUF1 (N228, N227);
buf BUF1 (N229, N221);
nor NOR4 (N230, N223, N1, N8, N176);
xor XOR2 (N231, N220, N5);
buf BUF1 (N232, N230);
and AND2 (N233, N225, N106);
nor NOR3 (N234, N231, N187, N137);
or OR2 (N235, N228, N153);
xor XOR2 (N236, N215, N225);
xor XOR2 (N237, N234, N96);
not NOT1 (N238, N197);
nor NOR2 (N239, N232, N220);
nor NOR4 (N240, N217, N41, N172, N108);
nand NAND4 (N241, N229, N219, N73, N84);
and AND4 (N242, N212, N237, N86, N44);
nand NAND3 (N243, N108, N69, N60);
and AND2 (N244, N226, N33);
not NOT1 (N245, N236);
not NOT1 (N246, N240);
not NOT1 (N247, N239);
nand NAND2 (N248, N241, N150);
and AND2 (N249, N246, N115);
or OR3 (N250, N248, N89, N144);
nand NAND3 (N251, N238, N242, N170);
buf BUF1 (N252, N242);
xor XOR2 (N253, N251, N127);
not NOT1 (N254, N235);
nand NAND2 (N255, N244, N230);
not NOT1 (N256, N233);
and AND3 (N257, N249, N249, N85);
nand NAND3 (N258, N245, N182, N105);
and AND3 (N259, N243, N246, N186);
buf BUF1 (N260, N252);
or OR2 (N261, N247, N182);
nand NAND2 (N262, N255, N193);
not NOT1 (N263, N258);
xor XOR2 (N264, N253, N248);
or OR4 (N265, N263, N181, N67, N16);
or OR4 (N266, N259, N187, N241, N205);
not NOT1 (N267, N262);
nor NOR3 (N268, N267, N105, N159);
xor XOR2 (N269, N256, N80);
not NOT1 (N270, N257);
nand NAND4 (N271, N261, N54, N259, N159);
not NOT1 (N272, N268);
or OR4 (N273, N254, N227, N221, N171);
or OR4 (N274, N273, N91, N62, N81);
buf BUF1 (N275, N266);
nor NOR3 (N276, N272, N76, N152);
nor NOR2 (N277, N270, N202);
nor NOR2 (N278, N277, N243);
and AND2 (N279, N271, N77);
nor NOR3 (N280, N274, N28, N32);
or OR3 (N281, N279, N3, N79);
not NOT1 (N282, N269);
or OR2 (N283, N265, N111);
not NOT1 (N284, N280);
xor XOR2 (N285, N250, N230);
not NOT1 (N286, N260);
and AND4 (N287, N264, N139, N177, N256);
not NOT1 (N288, N281);
not NOT1 (N289, N278);
xor XOR2 (N290, N282, N170);
or OR4 (N291, N276, N134, N237, N234);
or OR2 (N292, N287, N8);
and AND2 (N293, N284, N57);
or OR2 (N294, N290, N134);
nand NAND2 (N295, N294, N273);
not NOT1 (N296, N293);
buf BUF1 (N297, N292);
nor NOR3 (N298, N288, N202, N175);
buf BUF1 (N299, N297);
nor NOR4 (N300, N298, N216, N124, N272);
or OR3 (N301, N283, N254, N205);
xor XOR2 (N302, N301, N104);
not NOT1 (N303, N289);
buf BUF1 (N304, N286);
nand NAND4 (N305, N275, N17, N301, N108);
not NOT1 (N306, N302);
nand NAND4 (N307, N300, N34, N55, N297);
nor NOR3 (N308, N304, N57, N36);
and AND4 (N309, N307, N26, N209, N77);
not NOT1 (N310, N291);
not NOT1 (N311, N308);
xor XOR2 (N312, N299, N3);
xor XOR2 (N313, N296, N310);
nor NOR2 (N314, N222, N190);
and AND4 (N315, N313, N176, N178, N72);
not NOT1 (N316, N309);
or OR2 (N317, N315, N18);
and AND3 (N318, N285, N220, N184);
or OR4 (N319, N305, N145, N72, N298);
nor NOR2 (N320, N306, N38);
buf BUF1 (N321, N319);
xor XOR2 (N322, N312, N187);
buf BUF1 (N323, N295);
or OR3 (N324, N323, N188, N110);
not NOT1 (N325, N317);
nand NAND2 (N326, N303, N104);
buf BUF1 (N327, N325);
or OR2 (N328, N321, N51);
nor NOR4 (N329, N326, N205, N116, N35);
xor XOR2 (N330, N328, N16);
nand NAND3 (N331, N329, N66, N308);
xor XOR2 (N332, N331, N104);
and AND4 (N333, N322, N298, N95, N290);
buf BUF1 (N334, N316);
buf BUF1 (N335, N330);
nor NOR2 (N336, N335, N319);
not NOT1 (N337, N318);
not NOT1 (N338, N337);
or OR2 (N339, N338, N298);
nand NAND2 (N340, N311, N80);
or OR2 (N341, N334, N17);
nand NAND2 (N342, N324, N232);
xor XOR2 (N343, N336, N9);
nor NOR2 (N344, N314, N151);
nor NOR4 (N345, N332, N91, N195, N7);
nor NOR4 (N346, N339, N121, N13, N87);
and AND2 (N347, N342, N243);
and AND2 (N348, N327, N14);
nand NAND3 (N349, N340, N187, N201);
nand NAND3 (N350, N341, N207, N330);
buf BUF1 (N351, N350);
or OR2 (N352, N349, N224);
or OR4 (N353, N345, N89, N241, N114);
and AND4 (N354, N320, N248, N296, N16);
not NOT1 (N355, N346);
nand NAND4 (N356, N352, N347, N264, N74);
buf BUF1 (N357, N20);
and AND3 (N358, N356, N143, N8);
nand NAND4 (N359, N358, N166, N153, N258);
nand NAND3 (N360, N354, N120, N173);
nand NAND2 (N361, N353, N198);
nand NAND3 (N362, N348, N126, N101);
not NOT1 (N363, N351);
buf BUF1 (N364, N343);
xor XOR2 (N365, N357, N232);
or OR4 (N366, N364, N78, N333, N112);
not NOT1 (N367, N220);
not NOT1 (N368, N365);
and AND4 (N369, N367, N49, N210, N307);
nand NAND2 (N370, N355, N52);
or OR4 (N371, N360, N270, N194, N216);
xor XOR2 (N372, N366, N300);
xor XOR2 (N373, N369, N28);
not NOT1 (N374, N344);
buf BUF1 (N375, N373);
not NOT1 (N376, N362);
nand NAND2 (N377, N374, N150);
not NOT1 (N378, N372);
and AND3 (N379, N377, N101, N213);
xor XOR2 (N380, N368, N111);
not NOT1 (N381, N371);
nand NAND2 (N382, N380, N67);
nand NAND3 (N383, N376, N94, N282);
buf BUF1 (N384, N359);
and AND4 (N385, N379, N29, N200, N84);
nand NAND2 (N386, N363, N85);
nor NOR2 (N387, N361, N220);
or OR2 (N388, N384, N161);
buf BUF1 (N389, N388);
not NOT1 (N390, N381);
or OR3 (N391, N378, N153, N26);
and AND2 (N392, N391, N301);
nor NOR3 (N393, N385, N19, N178);
nand NAND3 (N394, N390, N268, N229);
xor XOR2 (N395, N392, N121);
or OR4 (N396, N383, N219, N335, N210);
not NOT1 (N397, N370);
not NOT1 (N398, N396);
nand NAND2 (N399, N389, N175);
or OR2 (N400, N387, N202);
or OR2 (N401, N395, N215);
xor XOR2 (N402, N386, N354);
and AND4 (N403, N402, N72, N398, N142);
and AND4 (N404, N104, N318, N328, N26);
xor XOR2 (N405, N399, N256);
nand NAND3 (N406, N375, N298, N302);
nor NOR3 (N407, N382, N137, N260);
not NOT1 (N408, N403);
or OR2 (N409, N408, N19);
xor XOR2 (N410, N394, N340);
or OR3 (N411, N407, N364, N149);
and AND3 (N412, N401, N94, N267);
xor XOR2 (N413, N406, N123);
not NOT1 (N414, N405);
or OR2 (N415, N413, N262);
nand NAND4 (N416, N411, N400, N300, N22);
buf BUF1 (N417, N247);
nand NAND4 (N418, N404, N210, N125, N89);
buf BUF1 (N419, N418);
xor XOR2 (N420, N414, N75);
nor NOR2 (N421, N415, N63);
or OR4 (N422, N416, N355, N232, N416);
or OR3 (N423, N412, N131, N215);
nor NOR4 (N424, N420, N122, N106, N372);
and AND2 (N425, N423, N170);
or OR3 (N426, N417, N4, N34);
not NOT1 (N427, N393);
nor NOR2 (N428, N425, N124);
nand NAND3 (N429, N421, N323, N332);
not NOT1 (N430, N397);
and AND4 (N431, N422, N5, N5, N294);
or OR4 (N432, N429, N263, N306, N165);
buf BUF1 (N433, N410);
not NOT1 (N434, N427);
nand NAND2 (N435, N430, N419);
buf BUF1 (N436, N178);
or OR3 (N437, N432, N330, N161);
xor XOR2 (N438, N431, N52);
nor NOR2 (N439, N409, N115);
not NOT1 (N440, N439);
not NOT1 (N441, N438);
xor XOR2 (N442, N435, N375);
nand NAND4 (N443, N424, N188, N100, N209);
nor NOR3 (N444, N437, N428, N359);
or OR2 (N445, N44, N438);
xor XOR2 (N446, N445, N64);
and AND3 (N447, N433, N393, N353);
nor NOR3 (N448, N426, N186, N211);
not NOT1 (N449, N440);
xor XOR2 (N450, N444, N64);
or OR3 (N451, N450, N426, N259);
or OR3 (N452, N449, N210, N156);
or OR4 (N453, N443, N76, N370, N39);
nor NOR2 (N454, N441, N121);
nand NAND4 (N455, N454, N122, N71, N408);
nor NOR3 (N456, N455, N275, N126);
nor NOR3 (N457, N452, N411, N304);
and AND3 (N458, N446, N368, N358);
nand NAND2 (N459, N448, N432);
buf BUF1 (N460, N459);
and AND4 (N461, N456, N84, N51, N210);
xor XOR2 (N462, N451, N251);
nand NAND3 (N463, N460, N43, N362);
xor XOR2 (N464, N463, N128);
nand NAND2 (N465, N434, N249);
xor XOR2 (N466, N442, N345);
or OR4 (N467, N458, N123, N397, N171);
and AND2 (N468, N464, N195);
not NOT1 (N469, N467);
nor NOR3 (N470, N466, N369, N381);
buf BUF1 (N471, N453);
buf BUF1 (N472, N465);
nor NOR2 (N473, N436, N106);
buf BUF1 (N474, N461);
nor NOR4 (N475, N470, N338, N361, N56);
not NOT1 (N476, N474);
buf BUF1 (N477, N475);
not NOT1 (N478, N477);
xor XOR2 (N479, N478, N293);
nor NOR4 (N480, N447, N461, N33, N403);
not NOT1 (N481, N473);
nor NOR3 (N482, N476, N154, N353);
or OR4 (N483, N457, N56, N27, N205);
or OR3 (N484, N471, N254, N221);
nor NOR3 (N485, N468, N100, N59);
xor XOR2 (N486, N482, N326);
buf BUF1 (N487, N485);
xor XOR2 (N488, N481, N351);
and AND3 (N489, N462, N387, N176);
and AND3 (N490, N486, N133, N38);
xor XOR2 (N491, N488, N239);
xor XOR2 (N492, N483, N323);
nand NAND4 (N493, N484, N75, N118, N253);
and AND2 (N494, N472, N278);
nor NOR2 (N495, N487, N61);
nand NAND4 (N496, N492, N336, N90, N214);
or OR4 (N497, N495, N464, N139, N155);
and AND3 (N498, N493, N350, N381);
not NOT1 (N499, N491);
not NOT1 (N500, N499);
or OR4 (N501, N469, N478, N314, N418);
not NOT1 (N502, N489);
not NOT1 (N503, N479);
and AND3 (N504, N497, N109, N227);
nor NOR2 (N505, N500, N241);
or OR3 (N506, N494, N14, N502);
xor XOR2 (N507, N465, N145);
not NOT1 (N508, N506);
not NOT1 (N509, N496);
nand NAND4 (N510, N503, N76, N281, N347);
and AND4 (N511, N480, N108, N227, N5);
buf BUF1 (N512, N511);
nor NOR4 (N513, N507, N201, N295, N121);
not NOT1 (N514, N508);
nor NOR2 (N515, N505, N414);
and AND3 (N516, N504, N25, N246);
not NOT1 (N517, N490);
not NOT1 (N518, N515);
nand NAND3 (N519, N517, N206, N285);
buf BUF1 (N520, N509);
not NOT1 (N521, N516);
buf BUF1 (N522, N520);
not NOT1 (N523, N513);
or OR4 (N524, N519, N229, N42, N211);
nor NOR3 (N525, N512, N188, N290);
not NOT1 (N526, N523);
not NOT1 (N527, N525);
nor NOR2 (N528, N518, N92);
buf BUF1 (N529, N527);
or OR4 (N530, N498, N190, N238, N139);
not NOT1 (N531, N514);
not NOT1 (N532, N522);
or OR4 (N533, N501, N451, N60, N413);
buf BUF1 (N534, N533);
xor XOR2 (N535, N526, N5);
buf BUF1 (N536, N534);
and AND4 (N537, N529, N186, N82, N301);
xor XOR2 (N538, N537, N378);
buf BUF1 (N539, N521);
not NOT1 (N540, N535);
nor NOR4 (N541, N524, N202, N191, N462);
buf BUF1 (N542, N536);
buf BUF1 (N543, N531);
xor XOR2 (N544, N541, N336);
and AND2 (N545, N528, N466);
xor XOR2 (N546, N544, N395);
and AND4 (N547, N546, N51, N378, N301);
nand NAND2 (N548, N547, N141);
and AND3 (N549, N538, N144, N115);
xor XOR2 (N550, N548, N361);
buf BUF1 (N551, N530);
not NOT1 (N552, N545);
xor XOR2 (N553, N543, N244);
buf BUF1 (N554, N551);
nand NAND2 (N555, N510, N319);
nor NOR3 (N556, N540, N166, N539);
nand NAND2 (N557, N546, N266);
and AND2 (N558, N552, N355);
buf BUF1 (N559, N532);
buf BUF1 (N560, N554);
xor XOR2 (N561, N553, N289);
not NOT1 (N562, N549);
nor NOR2 (N563, N557, N507);
buf BUF1 (N564, N542);
buf BUF1 (N565, N560);
or OR4 (N566, N565, N494, N166, N243);
nor NOR3 (N567, N555, N433, N230);
or OR4 (N568, N556, N111, N59, N532);
nor NOR2 (N569, N563, N515);
or OR4 (N570, N569, N509, N32, N520);
nor NOR2 (N571, N562, N455);
buf BUF1 (N572, N570);
xor XOR2 (N573, N572, N419);
xor XOR2 (N574, N559, N358);
xor XOR2 (N575, N566, N541);
not NOT1 (N576, N574);
or OR3 (N577, N564, N167, N18);
and AND4 (N578, N550, N540, N191, N40);
nor NOR3 (N579, N576, N316, N104);
not NOT1 (N580, N558);
nor NOR3 (N581, N580, N59, N48);
xor XOR2 (N582, N571, N180);
buf BUF1 (N583, N575);
or OR4 (N584, N568, N407, N484, N224);
or OR4 (N585, N582, N537, N148, N77);
buf BUF1 (N586, N579);
buf BUF1 (N587, N577);
or OR3 (N588, N586, N542, N374);
nor NOR3 (N589, N581, N159, N24);
xor XOR2 (N590, N587, N488);
nand NAND2 (N591, N561, N303);
or OR3 (N592, N584, N485, N293);
and AND4 (N593, N591, N5, N123, N454);
nor NOR2 (N594, N578, N307);
nand NAND2 (N595, N590, N310);
nand NAND3 (N596, N592, N143, N276);
not NOT1 (N597, N589);
xor XOR2 (N598, N593, N151);
buf BUF1 (N599, N595);
xor XOR2 (N600, N588, N16);
not NOT1 (N601, N585);
buf BUF1 (N602, N573);
and AND4 (N603, N602, N146, N294, N442);
xor XOR2 (N604, N603, N14);
not NOT1 (N605, N594);
and AND3 (N606, N601, N117, N182);
xor XOR2 (N607, N600, N548);
or OR3 (N608, N606, N503, N407);
xor XOR2 (N609, N604, N136);
not NOT1 (N610, N596);
or OR4 (N611, N567, N465, N145, N332);
xor XOR2 (N612, N598, N247);
nand NAND2 (N613, N609, N100);
nand NAND2 (N614, N605, N148);
nand NAND2 (N615, N612, N608);
buf BUF1 (N616, N517);
or OR3 (N617, N611, N401, N82);
nor NOR2 (N618, N613, N25);
and AND2 (N619, N614, N605);
buf BUF1 (N620, N610);
xor XOR2 (N621, N607, N187);
or OR3 (N622, N620, N160, N568);
nand NAND4 (N623, N615, N577, N144, N434);
and AND4 (N624, N618, N142, N408, N74);
xor XOR2 (N625, N623, N439);
not NOT1 (N626, N624);
not NOT1 (N627, N622);
nor NOR4 (N628, N621, N292, N90, N68);
not NOT1 (N629, N583);
buf BUF1 (N630, N627);
not NOT1 (N631, N626);
or OR4 (N632, N597, N622, N524, N234);
or OR4 (N633, N632, N542, N161, N3);
buf BUF1 (N634, N616);
nand NAND2 (N635, N634, N581);
buf BUF1 (N636, N633);
nand NAND2 (N637, N630, N77);
and AND2 (N638, N619, N561);
xor XOR2 (N639, N637, N189);
nand NAND4 (N640, N636, N390, N62, N205);
and AND3 (N641, N640, N264, N171);
and AND2 (N642, N641, N298);
nor NOR2 (N643, N635, N290);
nor NOR2 (N644, N631, N444);
or OR4 (N645, N643, N78, N604, N353);
xor XOR2 (N646, N644, N37);
xor XOR2 (N647, N639, N562);
and AND2 (N648, N646, N565);
xor XOR2 (N649, N625, N540);
not NOT1 (N650, N628);
not NOT1 (N651, N650);
nor NOR2 (N652, N651, N49);
nor NOR3 (N653, N638, N62, N117);
buf BUF1 (N654, N647);
not NOT1 (N655, N652);
buf BUF1 (N656, N629);
buf BUF1 (N657, N642);
buf BUF1 (N658, N599);
or OR3 (N659, N656, N631, N221);
or OR4 (N660, N659, N417, N297, N486);
xor XOR2 (N661, N660, N349);
xor XOR2 (N662, N648, N455);
buf BUF1 (N663, N662);
xor XOR2 (N664, N657, N586);
nor NOR2 (N665, N617, N180);
xor XOR2 (N666, N645, N167);
not NOT1 (N667, N655);
and AND4 (N668, N661, N443, N39, N262);
or OR4 (N669, N666, N597, N107, N484);
nand NAND4 (N670, N663, N464, N405, N77);
buf BUF1 (N671, N670);
nor NOR2 (N672, N665, N104);
buf BUF1 (N673, N669);
xor XOR2 (N674, N658, N70);
not NOT1 (N675, N654);
nand NAND3 (N676, N671, N370, N382);
nand NAND2 (N677, N667, N515);
nor NOR4 (N678, N664, N114, N650, N568);
xor XOR2 (N679, N677, N237);
nor NOR2 (N680, N679, N476);
not NOT1 (N681, N668);
not NOT1 (N682, N653);
buf BUF1 (N683, N678);
and AND3 (N684, N675, N119, N539);
nor NOR3 (N685, N683, N635, N604);
nand NAND3 (N686, N685, N624, N29);
or OR3 (N687, N676, N42, N616);
buf BUF1 (N688, N686);
xor XOR2 (N689, N688, N106);
nor NOR2 (N690, N687, N243);
and AND3 (N691, N680, N471, N116);
or OR4 (N692, N689, N127, N611, N585);
and AND2 (N693, N649, N181);
and AND3 (N694, N684, N319, N282);
nand NAND4 (N695, N690, N429, N689, N349);
and AND3 (N696, N694, N340, N360);
buf BUF1 (N697, N672);
and AND4 (N698, N692, N67, N251, N116);
xor XOR2 (N699, N674, N83);
xor XOR2 (N700, N697, N666);
not NOT1 (N701, N673);
xor XOR2 (N702, N693, N286);
not NOT1 (N703, N702);
xor XOR2 (N704, N703, N154);
not NOT1 (N705, N695);
nor NOR2 (N706, N698, N386);
and AND4 (N707, N691, N11, N135, N165);
nor NOR2 (N708, N682, N136);
buf BUF1 (N709, N708);
or OR3 (N710, N706, N291, N394);
nand NAND3 (N711, N707, N434, N32);
and AND2 (N712, N699, N502);
or OR3 (N713, N709, N550, N708);
or OR4 (N714, N710, N583, N70, N440);
and AND4 (N715, N701, N609, N403, N383);
nor NOR4 (N716, N696, N488, N547, N238);
and AND4 (N717, N714, N181, N193, N53);
and AND2 (N718, N716, N405);
xor XOR2 (N719, N715, N226);
or OR3 (N720, N711, N154, N608);
nand NAND4 (N721, N713, N581, N210, N29);
buf BUF1 (N722, N718);
xor XOR2 (N723, N721, N263);
buf BUF1 (N724, N720);
not NOT1 (N725, N719);
and AND3 (N726, N700, N446, N132);
not NOT1 (N727, N723);
nor NOR2 (N728, N727, N240);
buf BUF1 (N729, N717);
xor XOR2 (N730, N681, N434);
not NOT1 (N731, N726);
nand NAND2 (N732, N728, N356);
buf BUF1 (N733, N732);
and AND2 (N734, N729, N461);
nor NOR3 (N735, N704, N297, N96);
xor XOR2 (N736, N722, N243);
nor NOR4 (N737, N731, N333, N508, N70);
or OR3 (N738, N730, N247, N683);
or OR3 (N739, N734, N682, N618);
nor NOR4 (N740, N736, N564, N333, N326);
nand NAND3 (N741, N725, N216, N504);
not NOT1 (N742, N712);
xor XOR2 (N743, N741, N740);
not NOT1 (N744, N74);
buf BUF1 (N745, N735);
nor NOR4 (N746, N733, N77, N642, N4);
or OR3 (N747, N743, N144, N212);
and AND3 (N748, N744, N669, N559);
nor NOR3 (N749, N739, N447, N86);
and AND4 (N750, N705, N742, N330, N549);
xor XOR2 (N751, N710, N499);
buf BUF1 (N752, N749);
nand NAND2 (N753, N745, N738);
and AND3 (N754, N180, N541, N89);
nor NOR3 (N755, N747, N698, N325);
nand NAND2 (N756, N746, N87);
xor XOR2 (N757, N737, N165);
nand NAND4 (N758, N750, N338, N546, N184);
nand NAND3 (N759, N753, N274, N716);
and AND4 (N760, N752, N694, N231, N342);
not NOT1 (N761, N756);
nor NOR3 (N762, N724, N633, N88);
xor XOR2 (N763, N754, N390);
nand NAND4 (N764, N759, N696, N380, N556);
not NOT1 (N765, N748);
nand NAND3 (N766, N757, N131, N756);
buf BUF1 (N767, N755);
nor NOR3 (N768, N751, N537, N17);
buf BUF1 (N769, N758);
nor NOR3 (N770, N764, N628, N169);
xor XOR2 (N771, N770, N737);
and AND2 (N772, N765, N534);
nor NOR4 (N773, N769, N81, N506, N161);
not NOT1 (N774, N772);
or OR2 (N775, N766, N366);
or OR2 (N776, N774, N278);
nand NAND3 (N777, N768, N419, N104);
nor NOR2 (N778, N762, N375);
not NOT1 (N779, N778);
nor NOR4 (N780, N771, N381, N673, N413);
buf BUF1 (N781, N780);
nor NOR3 (N782, N760, N154, N115);
nor NOR3 (N783, N779, N565, N619);
nor NOR4 (N784, N783, N82, N185, N289);
or OR2 (N785, N767, N554);
and AND4 (N786, N785, N504, N250, N406);
nand NAND4 (N787, N773, N624, N328, N8);
or OR3 (N788, N777, N494, N83);
and AND4 (N789, N775, N465, N25, N546);
or OR3 (N790, N781, N457, N217);
buf BUF1 (N791, N788);
xor XOR2 (N792, N786, N324);
nor NOR3 (N793, N784, N485, N367);
nor NOR4 (N794, N782, N257, N675, N9);
or OR2 (N795, N794, N243);
nand NAND3 (N796, N793, N521, N413);
buf BUF1 (N797, N787);
not NOT1 (N798, N789);
buf BUF1 (N799, N795);
nor NOR4 (N800, N798, N200, N704, N682);
and AND2 (N801, N761, N603);
or OR3 (N802, N799, N467, N109);
nand NAND4 (N803, N792, N123, N497, N211);
nor NOR2 (N804, N763, N124);
and AND2 (N805, N797, N150);
nand NAND2 (N806, N802, N60);
nand NAND4 (N807, N790, N576, N681, N714);
or OR2 (N808, N807, N150);
and AND2 (N809, N808, N489);
or OR2 (N810, N800, N12);
buf BUF1 (N811, N801);
nor NOR4 (N812, N811, N612, N360, N540);
xor XOR2 (N813, N809, N727);
nand NAND2 (N814, N813, N789);
not NOT1 (N815, N803);
buf BUF1 (N816, N814);
not NOT1 (N817, N805);
not NOT1 (N818, N812);
buf BUF1 (N819, N796);
or OR2 (N820, N816, N359);
and AND3 (N821, N820, N522, N278);
or OR2 (N822, N818, N547);
xor XOR2 (N823, N817, N622);
nor NOR4 (N824, N791, N802, N490, N529);
xor XOR2 (N825, N815, N256);
nand NAND4 (N826, N810, N93, N820, N547);
nand NAND2 (N827, N776, N514);
buf BUF1 (N828, N804);
nor NOR3 (N829, N806, N233, N266);
nand NAND4 (N830, N823, N276, N554, N568);
xor XOR2 (N831, N824, N554);
and AND3 (N832, N826, N87, N643);
buf BUF1 (N833, N832);
nor NOR4 (N834, N827, N476, N793, N785);
or OR2 (N835, N829, N765);
not NOT1 (N836, N833);
nor NOR4 (N837, N830, N358, N39, N69);
buf BUF1 (N838, N836);
buf BUF1 (N839, N834);
nor NOR4 (N840, N819, N423, N73, N701);
not NOT1 (N841, N840);
xor XOR2 (N842, N831, N275);
nand NAND2 (N843, N839, N823);
nand NAND4 (N844, N838, N154, N279, N650);
nand NAND2 (N845, N821, N767);
nand NAND2 (N846, N835, N518);
nor NOR3 (N847, N828, N335, N611);
nand NAND4 (N848, N825, N833, N29, N66);
not NOT1 (N849, N847);
and AND3 (N850, N845, N425, N846);
not NOT1 (N851, N247);
or OR3 (N852, N837, N660, N163);
xor XOR2 (N853, N850, N197);
or OR3 (N854, N843, N303, N793);
nor NOR4 (N855, N848, N444, N109, N431);
or OR3 (N856, N853, N209, N604);
or OR3 (N857, N841, N416, N682);
xor XOR2 (N858, N856, N276);
not NOT1 (N859, N857);
and AND3 (N860, N849, N299, N637);
or OR3 (N861, N844, N127, N294);
and AND3 (N862, N860, N592, N32);
nand NAND3 (N863, N861, N620, N419);
xor XOR2 (N864, N855, N144);
nor NOR3 (N865, N864, N569, N525);
nand NAND2 (N866, N863, N30);
xor XOR2 (N867, N866, N277);
xor XOR2 (N868, N867, N596);
not NOT1 (N869, N865);
xor XOR2 (N870, N842, N404);
and AND3 (N871, N869, N16, N123);
nor NOR3 (N872, N871, N415, N92);
and AND3 (N873, N854, N611, N606);
buf BUF1 (N874, N851);
nand NAND3 (N875, N858, N553, N179);
and AND2 (N876, N868, N224);
buf BUF1 (N877, N872);
and AND2 (N878, N852, N838);
not NOT1 (N879, N870);
buf BUF1 (N880, N874);
buf BUF1 (N881, N873);
xor XOR2 (N882, N877, N654);
nand NAND3 (N883, N880, N543, N66);
or OR2 (N884, N859, N743);
nor NOR3 (N885, N882, N162, N873);
and AND2 (N886, N822, N426);
and AND3 (N887, N885, N788, N329);
nand NAND3 (N888, N878, N451, N859);
nor NOR3 (N889, N887, N572, N688);
nand NAND2 (N890, N886, N477);
or OR2 (N891, N883, N645);
nor NOR2 (N892, N888, N505);
not NOT1 (N893, N889);
xor XOR2 (N894, N884, N783);
buf BUF1 (N895, N875);
not NOT1 (N896, N881);
not NOT1 (N897, N890);
xor XOR2 (N898, N893, N745);
nor NOR2 (N899, N892, N413);
xor XOR2 (N900, N896, N355);
xor XOR2 (N901, N899, N336);
nand NAND2 (N902, N891, N752);
xor XOR2 (N903, N879, N712);
and AND3 (N904, N902, N357, N193);
or OR3 (N905, N894, N629, N575);
nor NOR4 (N906, N876, N798, N732, N232);
not NOT1 (N907, N901);
or OR2 (N908, N907, N97);
nand NAND4 (N909, N905, N748, N413, N503);
nand NAND2 (N910, N900, N388);
nor NOR4 (N911, N895, N647, N267, N668);
and AND4 (N912, N908, N524, N43, N5);
xor XOR2 (N913, N906, N478);
or OR4 (N914, N903, N801, N417, N368);
and AND3 (N915, N904, N579, N755);
and AND4 (N916, N910, N577, N291, N772);
not NOT1 (N917, N862);
and AND3 (N918, N915, N681, N63);
and AND4 (N919, N916, N457, N648, N636);
and AND2 (N920, N913, N92);
xor XOR2 (N921, N919, N559);
not NOT1 (N922, N917);
or OR2 (N923, N922, N403);
nor NOR4 (N924, N897, N81, N549, N708);
nor NOR4 (N925, N924, N484, N195, N575);
not NOT1 (N926, N920);
not NOT1 (N927, N918);
and AND3 (N928, N912, N347, N461);
and AND3 (N929, N911, N775, N536);
nand NAND4 (N930, N928, N733, N392, N429);
nand NAND2 (N931, N927, N779);
not NOT1 (N932, N931);
not NOT1 (N933, N930);
not NOT1 (N934, N926);
or OR4 (N935, N921, N715, N550, N480);
buf BUF1 (N936, N934);
nor NOR2 (N937, N933, N329);
xor XOR2 (N938, N932, N933);
not NOT1 (N939, N935);
not NOT1 (N940, N923);
buf BUF1 (N941, N914);
or OR3 (N942, N936, N510, N607);
nand NAND2 (N943, N937, N505);
nor NOR2 (N944, N929, N156);
not NOT1 (N945, N898);
nand NAND2 (N946, N945, N438);
xor XOR2 (N947, N940, N428);
or OR4 (N948, N938, N612, N703, N917);
or OR3 (N949, N943, N817, N612);
nand NAND2 (N950, N944, N235);
nor NOR4 (N951, N947, N663, N945, N307);
buf BUF1 (N952, N942);
nor NOR3 (N953, N948, N853, N269);
xor XOR2 (N954, N941, N273);
nor NOR3 (N955, N951, N199, N555);
nor NOR3 (N956, N954, N469, N205);
buf BUF1 (N957, N956);
and AND2 (N958, N946, N276);
and AND2 (N959, N957, N12);
nand NAND2 (N960, N950, N299);
not NOT1 (N961, N925);
buf BUF1 (N962, N959);
and AND2 (N963, N953, N353);
not NOT1 (N964, N955);
buf BUF1 (N965, N909);
buf BUF1 (N966, N961);
or OR4 (N967, N962, N301, N875, N408);
not NOT1 (N968, N960);
buf BUF1 (N969, N967);
nor NOR2 (N970, N968, N291);
xor XOR2 (N971, N952, N111);
nor NOR3 (N972, N958, N676, N339);
or OR2 (N973, N972, N457);
nor NOR4 (N974, N973, N926, N330, N80);
or OR3 (N975, N965, N194, N111);
xor XOR2 (N976, N974, N12);
nand NAND3 (N977, N969, N850, N663);
xor XOR2 (N978, N939, N958);
buf BUF1 (N979, N949);
and AND2 (N980, N975, N776);
and AND2 (N981, N966, N266);
or OR2 (N982, N980, N361);
not NOT1 (N983, N982);
xor XOR2 (N984, N963, N260);
buf BUF1 (N985, N981);
xor XOR2 (N986, N979, N601);
and AND2 (N987, N984, N413);
buf BUF1 (N988, N987);
nor NOR2 (N989, N983, N227);
and AND4 (N990, N985, N339, N29, N980);
or OR4 (N991, N970, N691, N231, N100);
nand NAND4 (N992, N986, N846, N45, N687);
nand NAND3 (N993, N989, N228, N84);
or OR2 (N994, N988, N576);
nor NOR2 (N995, N994, N976);
buf BUF1 (N996, N630);
not NOT1 (N997, N993);
buf BUF1 (N998, N995);
not NOT1 (N999, N996);
buf BUF1 (N1000, N999);
nand NAND2 (N1001, N971, N535);
or OR2 (N1002, N997, N740);
nor NOR3 (N1003, N1001, N238, N295);
not NOT1 (N1004, N991);
xor XOR2 (N1005, N977, N577);
nor NOR3 (N1006, N992, N151, N608);
and AND4 (N1007, N1004, N174, N382, N359);
not NOT1 (N1008, N964);
and AND4 (N1009, N1003, N296, N633, N638);
or OR3 (N1010, N1005, N57, N914);
not NOT1 (N1011, N1006);
and AND2 (N1012, N1011, N124);
and AND4 (N1013, N990, N874, N618, N855);
nor NOR2 (N1014, N1013, N200);
nor NOR4 (N1015, N1002, N338, N225, N926);
nor NOR3 (N1016, N998, N154, N297);
or OR4 (N1017, N1015, N471, N449, N367);
nor NOR4 (N1018, N1008, N313, N314, N106);
xor XOR2 (N1019, N1018, N648);
nand NAND4 (N1020, N978, N173, N578, N818);
nor NOR3 (N1021, N1012, N192, N1009);
xor XOR2 (N1022, N303, N987);
nand NAND3 (N1023, N1017, N812, N207);
buf BUF1 (N1024, N1022);
not NOT1 (N1025, N1000);
nand NAND4 (N1026, N1016, N93, N512, N285);
buf BUF1 (N1027, N1023);
nand NAND3 (N1028, N1021, N72, N169);
buf BUF1 (N1029, N1028);
or OR4 (N1030, N1024, N964, N412, N149);
and AND3 (N1031, N1014, N616, N257);
nor NOR4 (N1032, N1031, N216, N641, N505);
and AND4 (N1033, N1027, N555, N517, N795);
xor XOR2 (N1034, N1029, N459);
nand NAND2 (N1035, N1026, N477);
nor NOR2 (N1036, N1032, N946);
and AND2 (N1037, N1036, N477);
and AND3 (N1038, N1035, N967, N491);
nor NOR3 (N1039, N1010, N87, N4);
nand NAND4 (N1040, N1007, N378, N938, N688);
and AND3 (N1041, N1019, N293, N980);
or OR4 (N1042, N1025, N452, N659, N867);
not NOT1 (N1043, N1040);
not NOT1 (N1044, N1041);
not NOT1 (N1045, N1034);
buf BUF1 (N1046, N1033);
or OR4 (N1047, N1045, N892, N314, N166);
xor XOR2 (N1048, N1039, N996);
nand NAND3 (N1049, N1044, N126, N696);
nand NAND4 (N1050, N1037, N31, N403, N545);
nand NAND3 (N1051, N1050, N769, N751);
nand NAND4 (N1052, N1038, N1007, N968, N796);
nand NAND3 (N1053, N1048, N192, N944);
not NOT1 (N1054, N1053);
buf BUF1 (N1055, N1049);
xor XOR2 (N1056, N1052, N383);
nand NAND3 (N1057, N1046, N879, N784);
nand NAND4 (N1058, N1043, N67, N747, N661);
xor XOR2 (N1059, N1030, N26);
not NOT1 (N1060, N1051);
xor XOR2 (N1061, N1054, N898);
and AND4 (N1062, N1060, N243, N468, N879);
buf BUF1 (N1063, N1056);
and AND4 (N1064, N1055, N303, N249, N54);
or OR2 (N1065, N1061, N590);
buf BUF1 (N1066, N1065);
nand NAND2 (N1067, N1066, N541);
not NOT1 (N1068, N1058);
nor NOR3 (N1069, N1020, N457, N819);
nand NAND4 (N1070, N1059, N20, N723, N234);
nor NOR2 (N1071, N1057, N851);
xor XOR2 (N1072, N1070, N489);
and AND2 (N1073, N1072, N730);
buf BUF1 (N1074, N1068);
and AND2 (N1075, N1047, N1063);
nand NAND4 (N1076, N71, N540, N1027, N706);
xor XOR2 (N1077, N1075, N720);
not NOT1 (N1078, N1076);
or OR2 (N1079, N1064, N1033);
xor XOR2 (N1080, N1077, N81);
and AND2 (N1081, N1042, N570);
and AND2 (N1082, N1074, N257);
or OR3 (N1083, N1082, N27, N278);
xor XOR2 (N1084, N1081, N619);
nor NOR4 (N1085, N1078, N1022, N872, N498);
buf BUF1 (N1086, N1083);
nand NAND3 (N1087, N1085, N649, N219);
or OR4 (N1088, N1079, N620, N767, N340);
not NOT1 (N1089, N1080);
and AND3 (N1090, N1088, N489, N750);
or OR2 (N1091, N1071, N692);
buf BUF1 (N1092, N1086);
buf BUF1 (N1093, N1067);
or OR4 (N1094, N1069, N384, N535, N268);
not NOT1 (N1095, N1062);
nand NAND3 (N1096, N1092, N794, N665);
and AND2 (N1097, N1095, N884);
not NOT1 (N1098, N1084);
nor NOR4 (N1099, N1094, N353, N553, N857);
nor NOR2 (N1100, N1091, N773);
nand NAND3 (N1101, N1099, N927, N637);
buf BUF1 (N1102, N1097);
not NOT1 (N1103, N1087);
nand NAND2 (N1104, N1098, N715);
nor NOR4 (N1105, N1096, N155, N706, N72);
xor XOR2 (N1106, N1093, N33);
and AND4 (N1107, N1102, N396, N142, N718);
and AND4 (N1108, N1105, N396, N892, N339);
nor NOR2 (N1109, N1104, N895);
nor NOR3 (N1110, N1106, N641, N555);
not NOT1 (N1111, N1103);
or OR3 (N1112, N1101, N617, N829);
or OR3 (N1113, N1111, N869, N126);
nand NAND3 (N1114, N1107, N217, N321);
not NOT1 (N1115, N1073);
and AND2 (N1116, N1100, N852);
nand NAND4 (N1117, N1089, N944, N906, N237);
xor XOR2 (N1118, N1116, N27);
or OR4 (N1119, N1117, N738, N341, N197);
or OR3 (N1120, N1115, N802, N641);
buf BUF1 (N1121, N1118);
xor XOR2 (N1122, N1114, N570);
and AND2 (N1123, N1119, N982);
nand NAND2 (N1124, N1090, N817);
nor NOR3 (N1125, N1121, N315, N39);
nor NOR4 (N1126, N1110, N612, N136, N730);
not NOT1 (N1127, N1126);
or OR3 (N1128, N1123, N151, N934);
or OR3 (N1129, N1113, N781, N252);
xor XOR2 (N1130, N1120, N349);
buf BUF1 (N1131, N1109);
xor XOR2 (N1132, N1124, N892);
or OR2 (N1133, N1131, N128);
nor NOR2 (N1134, N1133, N808);
nand NAND3 (N1135, N1125, N608, N579);
not NOT1 (N1136, N1130);
buf BUF1 (N1137, N1132);
or OR3 (N1138, N1122, N876, N489);
nand NAND2 (N1139, N1108, N967);
or OR2 (N1140, N1136, N648);
or OR4 (N1141, N1134, N344, N16, N523);
nand NAND2 (N1142, N1128, N938);
xor XOR2 (N1143, N1112, N865);
or OR2 (N1144, N1139, N768);
nand NAND2 (N1145, N1135, N496);
and AND2 (N1146, N1143, N708);
xor XOR2 (N1147, N1140, N416);
nand NAND2 (N1148, N1141, N430);
nand NAND4 (N1149, N1144, N187, N906, N257);
buf BUF1 (N1150, N1142);
or OR4 (N1151, N1149, N535, N196, N890);
nor NOR3 (N1152, N1146, N873, N1052);
not NOT1 (N1153, N1145);
xor XOR2 (N1154, N1148, N784);
nor NOR3 (N1155, N1147, N762, N108);
not NOT1 (N1156, N1151);
or OR3 (N1157, N1129, N822, N260);
not NOT1 (N1158, N1155);
xor XOR2 (N1159, N1150, N1057);
nor NOR2 (N1160, N1158, N287);
nor NOR4 (N1161, N1138, N177, N61, N1002);
xor XOR2 (N1162, N1152, N49);
or OR3 (N1163, N1160, N665, N914);
nor NOR2 (N1164, N1127, N109);
and AND2 (N1165, N1164, N191);
or OR3 (N1166, N1163, N779, N1137);
buf BUF1 (N1167, N567);
nand NAND3 (N1168, N1154, N993, N460);
nand NAND4 (N1169, N1153, N122, N728, N713);
nor NOR2 (N1170, N1165, N190);
buf BUF1 (N1171, N1157);
buf BUF1 (N1172, N1156);
and AND4 (N1173, N1171, N2, N7, N752);
not NOT1 (N1174, N1172);
buf BUF1 (N1175, N1159);
buf BUF1 (N1176, N1169);
nor NOR3 (N1177, N1162, N1070, N147);
xor XOR2 (N1178, N1174, N983);
nor NOR4 (N1179, N1166, N1064, N798, N1132);
nand NAND3 (N1180, N1179, N600, N163);
and AND3 (N1181, N1161, N732, N975);
and AND2 (N1182, N1168, N715);
not NOT1 (N1183, N1170);
buf BUF1 (N1184, N1180);
nor NOR2 (N1185, N1183, N922);
xor XOR2 (N1186, N1178, N1095);
buf BUF1 (N1187, N1185);
xor XOR2 (N1188, N1173, N122);
xor XOR2 (N1189, N1182, N899);
buf BUF1 (N1190, N1181);
nor NOR2 (N1191, N1188, N921);
not NOT1 (N1192, N1189);
or OR2 (N1193, N1192, N557);
buf BUF1 (N1194, N1177);
nand NAND2 (N1195, N1176, N422);
nor NOR2 (N1196, N1194, N958);
not NOT1 (N1197, N1193);
not NOT1 (N1198, N1190);
not NOT1 (N1199, N1196);
or OR3 (N1200, N1199, N1112, N754);
not NOT1 (N1201, N1200);
not NOT1 (N1202, N1187);
buf BUF1 (N1203, N1198);
buf BUF1 (N1204, N1191);
nand NAND4 (N1205, N1186, N359, N699, N343);
nand NAND3 (N1206, N1175, N778, N617);
buf BUF1 (N1207, N1202);
nor NOR4 (N1208, N1201, N128, N564, N56);
xor XOR2 (N1209, N1208, N21);
and AND3 (N1210, N1204, N603, N285);
not NOT1 (N1211, N1184);
and AND3 (N1212, N1205, N895, N187);
and AND3 (N1213, N1211, N307, N306);
nand NAND2 (N1214, N1207, N180);
not NOT1 (N1215, N1209);
and AND4 (N1216, N1167, N39, N527, N27);
or OR2 (N1217, N1213, N946);
buf BUF1 (N1218, N1210);
not NOT1 (N1219, N1216);
nand NAND4 (N1220, N1203, N139, N1161, N181);
nand NAND4 (N1221, N1214, N729, N356, N637);
and AND4 (N1222, N1219, N281, N487, N579);
or OR3 (N1223, N1221, N447, N727);
and AND2 (N1224, N1220, N600);
nor NOR4 (N1225, N1195, N1088, N1145, N1011);
nand NAND2 (N1226, N1222, N586);
or OR2 (N1227, N1225, N164);
nor NOR2 (N1228, N1223, N1044);
nand NAND3 (N1229, N1226, N1227, N769);
nor NOR2 (N1230, N194, N648);
xor XOR2 (N1231, N1224, N1101);
or OR3 (N1232, N1212, N1094, N798);
nor NOR2 (N1233, N1197, N289);
and AND2 (N1234, N1217, N710);
or OR2 (N1235, N1234, N796);
not NOT1 (N1236, N1233);
or OR4 (N1237, N1230, N111, N710, N77);
and AND4 (N1238, N1229, N694, N635, N405);
or OR2 (N1239, N1228, N181);
nor NOR3 (N1240, N1235, N712, N671);
and AND4 (N1241, N1215, N260, N67, N185);
buf BUF1 (N1242, N1218);
nand NAND2 (N1243, N1236, N408);
nor NOR4 (N1244, N1237, N474, N728, N542);
not NOT1 (N1245, N1239);
or OR4 (N1246, N1231, N1128, N663, N785);
and AND2 (N1247, N1241, N689);
xor XOR2 (N1248, N1243, N15);
not NOT1 (N1249, N1206);
nand NAND4 (N1250, N1249, N28, N1154, N423);
or OR2 (N1251, N1242, N949);
or OR4 (N1252, N1240, N389, N196, N1);
nor NOR2 (N1253, N1247, N43);
nor NOR2 (N1254, N1232, N641);
or OR4 (N1255, N1238, N953, N195, N1123);
or OR2 (N1256, N1246, N353);
buf BUF1 (N1257, N1256);
or OR2 (N1258, N1251, N544);
xor XOR2 (N1259, N1257, N281);
not NOT1 (N1260, N1259);
buf BUF1 (N1261, N1244);
and AND3 (N1262, N1254, N84, N951);
not NOT1 (N1263, N1255);
not NOT1 (N1264, N1245);
buf BUF1 (N1265, N1262);
or OR2 (N1266, N1253, N382);
nand NAND4 (N1267, N1252, N245, N876, N461);
not NOT1 (N1268, N1263);
nor NOR3 (N1269, N1267, N438, N419);
nor NOR3 (N1270, N1266, N641, N103);
or OR3 (N1271, N1258, N828, N1083);
nor NOR4 (N1272, N1268, N739, N583, N164);
and AND4 (N1273, N1265, N988, N436, N1057);
buf BUF1 (N1274, N1273);
buf BUF1 (N1275, N1264);
not NOT1 (N1276, N1261);
nor NOR2 (N1277, N1276, N475);
and AND2 (N1278, N1248, N983);
and AND3 (N1279, N1269, N94, N641);
xor XOR2 (N1280, N1260, N267);
nand NAND2 (N1281, N1278, N902);
buf BUF1 (N1282, N1280);
or OR4 (N1283, N1281, N887, N806, N176);
or OR4 (N1284, N1277, N470, N698, N531);
nor NOR3 (N1285, N1283, N1172, N494);
not NOT1 (N1286, N1272);
not NOT1 (N1287, N1285);
or OR4 (N1288, N1275, N189, N1005, N1273);
or OR2 (N1289, N1274, N662);
nand NAND4 (N1290, N1286, N1032, N485, N364);
nor NOR4 (N1291, N1288, N572, N544, N814);
nand NAND4 (N1292, N1282, N416, N963, N913);
not NOT1 (N1293, N1271);
and AND4 (N1294, N1293, N960, N232, N1006);
nor NOR2 (N1295, N1294, N409);
and AND2 (N1296, N1250, N1217);
nand NAND2 (N1297, N1289, N7);
or OR3 (N1298, N1270, N1181, N1076);
nand NAND4 (N1299, N1296, N586, N1012, N122);
nand NAND2 (N1300, N1298, N315);
buf BUF1 (N1301, N1297);
and AND4 (N1302, N1287, N948, N880, N854);
not NOT1 (N1303, N1301);
buf BUF1 (N1304, N1299);
or OR4 (N1305, N1290, N779, N72, N716);
buf BUF1 (N1306, N1304);
buf BUF1 (N1307, N1284);
buf BUF1 (N1308, N1307);
buf BUF1 (N1309, N1302);
buf BUF1 (N1310, N1309);
or OR3 (N1311, N1295, N1166, N791);
and AND2 (N1312, N1291, N627);
not NOT1 (N1313, N1303);
xor XOR2 (N1314, N1305, N345);
or OR2 (N1315, N1313, N1124);
and AND4 (N1316, N1306, N549, N291, N1119);
buf BUF1 (N1317, N1315);
nor NOR4 (N1318, N1314, N595, N312, N1129);
buf BUF1 (N1319, N1300);
not NOT1 (N1320, N1318);
nor NOR2 (N1321, N1320, N357);
not NOT1 (N1322, N1308);
nor NOR4 (N1323, N1292, N713, N961, N123);
and AND3 (N1324, N1311, N1094, N521);
or OR2 (N1325, N1319, N555);
nand NAND2 (N1326, N1325, N766);
nand NAND3 (N1327, N1312, N222, N903);
xor XOR2 (N1328, N1327, N969);
or OR2 (N1329, N1310, N467);
xor XOR2 (N1330, N1324, N1065);
buf BUF1 (N1331, N1317);
and AND4 (N1332, N1321, N446, N590, N685);
not NOT1 (N1333, N1328);
or OR3 (N1334, N1323, N907, N1249);
nor NOR2 (N1335, N1279, N678);
xor XOR2 (N1336, N1334, N1081);
or OR2 (N1337, N1330, N3);
nor NOR4 (N1338, N1329, N172, N77, N101);
buf BUF1 (N1339, N1331);
nand NAND4 (N1340, N1316, N1119, N957, N200);
not NOT1 (N1341, N1322);
nand NAND4 (N1342, N1341, N396, N976, N703);
or OR2 (N1343, N1333, N1281);
not NOT1 (N1344, N1332);
xor XOR2 (N1345, N1338, N2);
xor XOR2 (N1346, N1326, N842);
not NOT1 (N1347, N1342);
xor XOR2 (N1348, N1339, N663);
buf BUF1 (N1349, N1340);
nor NOR4 (N1350, N1345, N53, N509, N523);
nor NOR2 (N1351, N1343, N834);
buf BUF1 (N1352, N1344);
xor XOR2 (N1353, N1335, N1004);
xor XOR2 (N1354, N1336, N1243);
buf BUF1 (N1355, N1350);
buf BUF1 (N1356, N1354);
buf BUF1 (N1357, N1352);
buf BUF1 (N1358, N1337);
and AND2 (N1359, N1348, N452);
not NOT1 (N1360, N1347);
xor XOR2 (N1361, N1359, N631);
nand NAND2 (N1362, N1351, N74);
nor NOR4 (N1363, N1360, N1314, N1297, N109);
nand NAND4 (N1364, N1353, N159, N848, N595);
or OR4 (N1365, N1364, N1188, N65, N976);
nand NAND2 (N1366, N1361, N905);
buf BUF1 (N1367, N1358);
nor NOR4 (N1368, N1346, N638, N1249, N945);
and AND3 (N1369, N1362, N727, N22);
and AND3 (N1370, N1367, N811, N335);
buf BUF1 (N1371, N1365);
xor XOR2 (N1372, N1357, N542);
not NOT1 (N1373, N1371);
nand NAND4 (N1374, N1349, N1026, N1134, N1079);
and AND2 (N1375, N1363, N614);
and AND3 (N1376, N1356, N289, N588);
buf BUF1 (N1377, N1373);
xor XOR2 (N1378, N1366, N1070);
xor XOR2 (N1379, N1376, N267);
nor NOR4 (N1380, N1369, N1160, N1188, N435);
and AND4 (N1381, N1380, N138, N605, N58);
or OR4 (N1382, N1370, N439, N262, N767);
nor NOR3 (N1383, N1372, N1120, N818);
or OR3 (N1384, N1379, N973, N240);
and AND4 (N1385, N1355, N401, N493, N495);
or OR3 (N1386, N1382, N319, N48);
nor NOR2 (N1387, N1377, N572);
and AND4 (N1388, N1387, N625, N1215, N1332);
xor XOR2 (N1389, N1368, N1129);
or OR4 (N1390, N1389, N1007, N439, N1277);
buf BUF1 (N1391, N1378);
xor XOR2 (N1392, N1384, N1328);
xor XOR2 (N1393, N1388, N83);
xor XOR2 (N1394, N1375, N746);
or OR3 (N1395, N1381, N195, N622);
or OR3 (N1396, N1395, N1045, N255);
or OR2 (N1397, N1393, N680);
nor NOR4 (N1398, N1383, N1133, N900, N311);
and AND4 (N1399, N1386, N364, N1062, N180);
buf BUF1 (N1400, N1374);
not NOT1 (N1401, N1385);
or OR2 (N1402, N1394, N1098);
nand NAND2 (N1403, N1392, N116);
not NOT1 (N1404, N1398);
or OR4 (N1405, N1397, N79, N75, N702);
not NOT1 (N1406, N1404);
not NOT1 (N1407, N1403);
xor XOR2 (N1408, N1390, N175);
or OR3 (N1409, N1400, N1142, N144);
or OR3 (N1410, N1407, N41, N32);
nor NOR4 (N1411, N1410, N972, N698, N28);
xor XOR2 (N1412, N1409, N841);
xor XOR2 (N1413, N1402, N1251);
nor NOR3 (N1414, N1391, N1014, N1112);
xor XOR2 (N1415, N1405, N1414);
nand NAND3 (N1416, N391, N1406, N1399);
not NOT1 (N1417, N199);
buf BUF1 (N1418, N587);
buf BUF1 (N1419, N1401);
buf BUF1 (N1420, N1411);
nor NOR3 (N1421, N1415, N70, N670);
and AND4 (N1422, N1413, N767, N761, N1286);
nand NAND4 (N1423, N1420, N600, N902, N1159);
nand NAND3 (N1424, N1416, N585, N264);
or OR3 (N1425, N1422, N872, N294);
buf BUF1 (N1426, N1418);
nor NOR2 (N1427, N1421, N1065);
not NOT1 (N1428, N1408);
and AND4 (N1429, N1425, N471, N1282, N797);
xor XOR2 (N1430, N1396, N923);
or OR3 (N1431, N1424, N1416, N1104);
xor XOR2 (N1432, N1431, N1216);
and AND2 (N1433, N1419, N110);
or OR3 (N1434, N1428, N956, N536);
nor NOR3 (N1435, N1432, N240, N267);
or OR3 (N1436, N1417, N40, N1252);
buf BUF1 (N1437, N1430);
or OR2 (N1438, N1435, N148);
not NOT1 (N1439, N1437);
buf BUF1 (N1440, N1412);
buf BUF1 (N1441, N1434);
nor NOR2 (N1442, N1429, N753);
xor XOR2 (N1443, N1439, N921);
nor NOR3 (N1444, N1441, N835, N426);
not NOT1 (N1445, N1433);
xor XOR2 (N1446, N1442, N1390);
nand NAND4 (N1447, N1426, N1302, N617, N74);
nand NAND4 (N1448, N1440, N1260, N394, N669);
not NOT1 (N1449, N1444);
or OR4 (N1450, N1438, N280, N905, N958);
not NOT1 (N1451, N1445);
xor XOR2 (N1452, N1436, N509);
or OR4 (N1453, N1452, N396, N1444, N361);
nor NOR2 (N1454, N1448, N1418);
nand NAND4 (N1455, N1446, N593, N313, N988);
and AND2 (N1456, N1450, N409);
and AND3 (N1457, N1427, N655, N937);
nand NAND4 (N1458, N1449, N1308, N1417, N235);
buf BUF1 (N1459, N1453);
or OR2 (N1460, N1447, N607);
buf BUF1 (N1461, N1455);
buf BUF1 (N1462, N1457);
and AND2 (N1463, N1462, N495);
or OR4 (N1464, N1454, N620, N455, N1343);
and AND3 (N1465, N1451, N1207, N875);
or OR3 (N1466, N1459, N1165, N1098);
and AND3 (N1467, N1443, N1185, N139);
nor NOR3 (N1468, N1460, N220, N740);
or OR3 (N1469, N1466, N157, N354);
buf BUF1 (N1470, N1468);
not NOT1 (N1471, N1458);
or OR2 (N1472, N1467, N372);
nor NOR4 (N1473, N1469, N542, N693, N1147);
and AND4 (N1474, N1464, N404, N496, N351);
not NOT1 (N1475, N1461);
xor XOR2 (N1476, N1470, N734);
nor NOR4 (N1477, N1463, N1284, N1458, N668);
xor XOR2 (N1478, N1474, N422);
nand NAND4 (N1479, N1478, N244, N202, N774);
xor XOR2 (N1480, N1465, N126);
and AND3 (N1481, N1477, N56, N550);
nor NOR2 (N1482, N1475, N1428);
nand NAND3 (N1483, N1482, N967, N1333);
xor XOR2 (N1484, N1483, N1284);
and AND3 (N1485, N1481, N648, N498);
or OR4 (N1486, N1473, N50, N830, N195);
nor NOR4 (N1487, N1480, N148, N672, N1179);
and AND4 (N1488, N1484, N1046, N1158, N807);
or OR3 (N1489, N1486, N1413, N991);
nand NAND3 (N1490, N1471, N1172, N974);
or OR3 (N1491, N1472, N174, N354);
or OR2 (N1492, N1476, N243);
buf BUF1 (N1493, N1492);
nor NOR4 (N1494, N1488, N1223, N133, N935);
or OR4 (N1495, N1487, N422, N430, N1028);
xor XOR2 (N1496, N1485, N617);
xor XOR2 (N1497, N1491, N1304);
nor NOR2 (N1498, N1456, N842);
or OR4 (N1499, N1495, N1490, N1125, N1306);
buf BUF1 (N1500, N355);
or OR4 (N1501, N1500, N624, N231, N926);
not NOT1 (N1502, N1499);
not NOT1 (N1503, N1502);
not NOT1 (N1504, N1503);
buf BUF1 (N1505, N1423);
and AND2 (N1506, N1489, N945);
and AND2 (N1507, N1496, N1430);
buf BUF1 (N1508, N1493);
nand NAND2 (N1509, N1506, N1390);
nand NAND4 (N1510, N1508, N1389, N1385, N312);
or OR3 (N1511, N1507, N1163, N567);
and AND3 (N1512, N1498, N392, N779);
not NOT1 (N1513, N1497);
nor NOR3 (N1514, N1494, N49, N47);
buf BUF1 (N1515, N1501);
nor NOR2 (N1516, N1479, N1381);
buf BUF1 (N1517, N1515);
buf BUF1 (N1518, N1505);
xor XOR2 (N1519, N1510, N829);
buf BUF1 (N1520, N1513);
nor NOR4 (N1521, N1511, N862, N954, N273);
buf BUF1 (N1522, N1521);
xor XOR2 (N1523, N1512, N1074);
and AND2 (N1524, N1517, N1395);
or OR4 (N1525, N1519, N979, N168, N80);
nor NOR3 (N1526, N1522, N526, N720);
and AND4 (N1527, N1504, N630, N213, N806);
not NOT1 (N1528, N1516);
xor XOR2 (N1529, N1520, N645);
nand NAND3 (N1530, N1514, N1306, N1444);
nand NAND2 (N1531, N1530, N1480);
nand NAND3 (N1532, N1524, N1048, N986);
not NOT1 (N1533, N1532);
nor NOR4 (N1534, N1509, N290, N1372, N1026);
buf BUF1 (N1535, N1525);
not NOT1 (N1536, N1518);
and AND3 (N1537, N1533, N737, N1268);
buf BUF1 (N1538, N1527);
nand NAND2 (N1539, N1538, N1434);
not NOT1 (N1540, N1539);
nand NAND4 (N1541, N1529, N848, N594, N121);
xor XOR2 (N1542, N1540, N1007);
xor XOR2 (N1543, N1537, N519);
not NOT1 (N1544, N1542);
not NOT1 (N1545, N1523);
xor XOR2 (N1546, N1528, N712);
not NOT1 (N1547, N1536);
xor XOR2 (N1548, N1547, N834);
and AND3 (N1549, N1535, N500, N1484);
nand NAND3 (N1550, N1531, N967, N865);
and AND4 (N1551, N1546, N33, N711, N54);
not NOT1 (N1552, N1549);
nand NAND2 (N1553, N1544, N318);
not NOT1 (N1554, N1541);
not NOT1 (N1555, N1554);
nand NAND2 (N1556, N1555, N1050);
buf BUF1 (N1557, N1553);
xor XOR2 (N1558, N1534, N426);
or OR3 (N1559, N1548, N258, N809);
and AND4 (N1560, N1550, N831, N30, N995);
nand NAND4 (N1561, N1545, N1029, N93, N1088);
nand NAND4 (N1562, N1560, N317, N619, N982);
and AND3 (N1563, N1556, N1281, N752);
not NOT1 (N1564, N1552);
nor NOR4 (N1565, N1543, N837, N1135, N1);
or OR2 (N1566, N1564, N1281);
buf BUF1 (N1567, N1557);
nand NAND4 (N1568, N1558, N2, N1240, N1114);
and AND3 (N1569, N1566, N515, N1436);
xor XOR2 (N1570, N1559, N877);
nor NOR2 (N1571, N1562, N1412);
nand NAND2 (N1572, N1570, N956);
not NOT1 (N1573, N1569);
nand NAND2 (N1574, N1565, N946);
xor XOR2 (N1575, N1574, N831);
and AND2 (N1576, N1571, N929);
nor NOR4 (N1577, N1561, N1103, N1030, N1344);
xor XOR2 (N1578, N1572, N1371);
or OR3 (N1579, N1575, N213, N1150);
nor NOR2 (N1580, N1573, N1509);
nand NAND2 (N1581, N1568, N1028);
not NOT1 (N1582, N1578);
nor NOR2 (N1583, N1580, N640);
buf BUF1 (N1584, N1526);
xor XOR2 (N1585, N1576, N1388);
buf BUF1 (N1586, N1579);
nor NOR3 (N1587, N1581, N1451, N821);
nor NOR3 (N1588, N1582, N1180, N647);
and AND4 (N1589, N1567, N359, N454, N217);
xor XOR2 (N1590, N1588, N488);
and AND2 (N1591, N1590, N1114);
nor NOR2 (N1592, N1551, N735);
buf BUF1 (N1593, N1587);
nand NAND2 (N1594, N1585, N295);
xor XOR2 (N1595, N1594, N854);
nand NAND4 (N1596, N1595, N697, N1443, N254);
not NOT1 (N1597, N1584);
nor NOR4 (N1598, N1563, N1563, N1160, N745);
and AND4 (N1599, N1591, N4, N334, N122);
buf BUF1 (N1600, N1599);
nand NAND3 (N1601, N1593, N548, N877);
nand NAND2 (N1602, N1596, N574);
not NOT1 (N1603, N1589);
nand NAND4 (N1604, N1601, N252, N1533, N1004);
or OR2 (N1605, N1603, N359);
or OR4 (N1606, N1583, N126, N345, N1019);
xor XOR2 (N1607, N1606, N1350);
nand NAND4 (N1608, N1592, N697, N439, N632);
and AND4 (N1609, N1577, N843, N773, N104);
not NOT1 (N1610, N1607);
and AND3 (N1611, N1609, N671, N658);
nand NAND3 (N1612, N1586, N725, N1191);
buf BUF1 (N1613, N1610);
xor XOR2 (N1614, N1608, N619);
nor NOR4 (N1615, N1614, N516, N1012, N813);
or OR4 (N1616, N1600, N1192, N591, N177);
nand NAND3 (N1617, N1598, N649, N1331);
and AND3 (N1618, N1605, N36, N268);
nand NAND2 (N1619, N1615, N1316);
or OR2 (N1620, N1597, N1540);
nand NAND3 (N1621, N1618, N1215, N1340);
nor NOR3 (N1622, N1620, N1360, N366);
nor NOR3 (N1623, N1617, N377, N1305);
nor NOR4 (N1624, N1613, N550, N756, N934);
xor XOR2 (N1625, N1611, N19);
not NOT1 (N1626, N1616);
not NOT1 (N1627, N1602);
buf BUF1 (N1628, N1604);
nand NAND4 (N1629, N1619, N1062, N141, N349);
buf BUF1 (N1630, N1624);
nand NAND3 (N1631, N1621, N1061, N1278);
xor XOR2 (N1632, N1631, N1011);
or OR3 (N1633, N1630, N77, N1152);
nand NAND2 (N1634, N1626, N616);
and AND2 (N1635, N1622, N240);
or OR4 (N1636, N1627, N1231, N1034, N1366);
buf BUF1 (N1637, N1636);
or OR2 (N1638, N1623, N1534);
nor NOR4 (N1639, N1629, N784, N1457, N202);
nor NOR4 (N1640, N1638, N1486, N689, N781);
not NOT1 (N1641, N1634);
buf BUF1 (N1642, N1641);
and AND4 (N1643, N1637, N606, N619, N558);
not NOT1 (N1644, N1612);
not NOT1 (N1645, N1639);
or OR3 (N1646, N1635, N318, N1096);
nand NAND3 (N1647, N1625, N1609, N1398);
or OR3 (N1648, N1643, N1082, N1414);
xor XOR2 (N1649, N1646, N1250);
nand NAND2 (N1650, N1645, N459);
xor XOR2 (N1651, N1644, N151);
nand NAND4 (N1652, N1642, N1324, N1098, N556);
buf BUF1 (N1653, N1648);
nor NOR3 (N1654, N1647, N971, N1267);
nand NAND2 (N1655, N1632, N1022);
and AND4 (N1656, N1653, N1505, N1398, N105);
nor NOR4 (N1657, N1628, N95, N218, N397);
or OR2 (N1658, N1649, N723);
nand NAND2 (N1659, N1658, N621);
nor NOR3 (N1660, N1656, N569, N393);
and AND2 (N1661, N1660, N27);
and AND4 (N1662, N1651, N652, N1075, N668);
xor XOR2 (N1663, N1659, N329);
nand NAND4 (N1664, N1663, N1541, N986, N628);
or OR2 (N1665, N1640, N599);
buf BUF1 (N1666, N1650);
or OR3 (N1667, N1652, N1662, N186);
nand NAND3 (N1668, N471, N1645, N553);
nand NAND4 (N1669, N1661, N733, N50, N996);
nor NOR4 (N1670, N1633, N1336, N1566, N228);
or OR3 (N1671, N1664, N986, N1030);
xor XOR2 (N1672, N1654, N550);
xor XOR2 (N1673, N1667, N1460);
xor XOR2 (N1674, N1657, N1529);
nand NAND3 (N1675, N1665, N891, N987);
nor NOR3 (N1676, N1666, N572, N1359);
and AND3 (N1677, N1668, N327, N238);
nand NAND3 (N1678, N1676, N191, N135);
nor NOR2 (N1679, N1677, N1631);
nor NOR2 (N1680, N1679, N1284);
or OR4 (N1681, N1669, N443, N1427, N172);
and AND2 (N1682, N1681, N401);
nand NAND4 (N1683, N1682, N1216, N911, N1306);
not NOT1 (N1684, N1672);
not NOT1 (N1685, N1670);
nor NOR4 (N1686, N1678, N203, N1535, N1280);
and AND4 (N1687, N1686, N1091, N1136, N356);
xor XOR2 (N1688, N1674, N1096);
xor XOR2 (N1689, N1680, N96);
and AND2 (N1690, N1688, N1517);
nor NOR4 (N1691, N1675, N982, N470, N1469);
xor XOR2 (N1692, N1689, N412);
nand NAND2 (N1693, N1692, N1190);
and AND4 (N1694, N1690, N1446, N311, N501);
and AND4 (N1695, N1684, N1561, N1210, N666);
nor NOR4 (N1696, N1685, N965, N588, N151);
nor NOR2 (N1697, N1695, N676);
xor XOR2 (N1698, N1671, N1258);
buf BUF1 (N1699, N1691);
xor XOR2 (N1700, N1683, N239);
nor NOR3 (N1701, N1655, N1298, N463);
nor NOR3 (N1702, N1697, N1505, N449);
nand NAND2 (N1703, N1702, N272);
xor XOR2 (N1704, N1687, N757);
xor XOR2 (N1705, N1696, N1452);
xor XOR2 (N1706, N1705, N148);
nor NOR2 (N1707, N1701, N625);
and AND3 (N1708, N1704, N1178, N1617);
or OR2 (N1709, N1700, N1639);
nor NOR2 (N1710, N1693, N316);
not NOT1 (N1711, N1699);
not NOT1 (N1712, N1710);
xor XOR2 (N1713, N1707, N1662);
not NOT1 (N1714, N1694);
or OR3 (N1715, N1714, N1018, N713);
or OR4 (N1716, N1708, N450, N1314, N1656);
and AND3 (N1717, N1709, N1198, N65);
or OR3 (N1718, N1703, N598, N291);
and AND3 (N1719, N1673, N69, N945);
or OR3 (N1720, N1698, N1708, N90);
xor XOR2 (N1721, N1718, N509);
buf BUF1 (N1722, N1717);
not NOT1 (N1723, N1716);
and AND4 (N1724, N1720, N1137, N1614, N708);
xor XOR2 (N1725, N1712, N737);
or OR2 (N1726, N1722, N1547);
not NOT1 (N1727, N1715);
and AND2 (N1728, N1721, N1314);
not NOT1 (N1729, N1727);
buf BUF1 (N1730, N1706);
or OR2 (N1731, N1725, N1428);
not NOT1 (N1732, N1719);
not NOT1 (N1733, N1723);
xor XOR2 (N1734, N1713, N1554);
not NOT1 (N1735, N1726);
or OR2 (N1736, N1732, N376);
not NOT1 (N1737, N1728);
buf BUF1 (N1738, N1711);
nand NAND4 (N1739, N1733, N1420, N512, N543);
nand NAND2 (N1740, N1736, N657);
not NOT1 (N1741, N1737);
buf BUF1 (N1742, N1739);
buf BUF1 (N1743, N1741);
not NOT1 (N1744, N1730);
nand NAND4 (N1745, N1729, N1365, N1719, N154);
nor NOR4 (N1746, N1744, N1184, N29, N445);
nand NAND3 (N1747, N1734, N1027, N1275);
nor NOR4 (N1748, N1742, N153, N1298, N1314);
xor XOR2 (N1749, N1738, N202);
xor XOR2 (N1750, N1735, N893);
or OR2 (N1751, N1748, N301);
buf BUF1 (N1752, N1745);
not NOT1 (N1753, N1731);
xor XOR2 (N1754, N1740, N257);
not NOT1 (N1755, N1749);
not NOT1 (N1756, N1755);
and AND4 (N1757, N1753, N1068, N1132, N792);
or OR3 (N1758, N1751, N1481, N612);
or OR2 (N1759, N1758, N585);
and AND4 (N1760, N1743, N1202, N810, N112);
xor XOR2 (N1761, N1724, N731);
nand NAND3 (N1762, N1756, N123, N372);
buf BUF1 (N1763, N1757);
and AND4 (N1764, N1762, N1107, N476, N1420);
or OR3 (N1765, N1761, N947, N1276);
xor XOR2 (N1766, N1754, N1208);
nor NOR4 (N1767, N1763, N1271, N1741, N778);
nand NAND4 (N1768, N1764, N894, N1353, N524);
nor NOR3 (N1769, N1768, N1423, N1763);
not NOT1 (N1770, N1750);
and AND4 (N1771, N1767, N228, N1576, N1424);
not NOT1 (N1772, N1766);
xor XOR2 (N1773, N1771, N985);
or OR4 (N1774, N1772, N868, N280, N1312);
xor XOR2 (N1775, N1770, N491);
not NOT1 (N1776, N1774);
or OR3 (N1777, N1759, N676, N1259);
or OR3 (N1778, N1769, N980, N1251);
buf BUF1 (N1779, N1773);
nor NOR4 (N1780, N1765, N1473, N389, N865);
xor XOR2 (N1781, N1775, N1024);
and AND2 (N1782, N1752, N1060);
xor XOR2 (N1783, N1779, N553);
not NOT1 (N1784, N1780);
or OR3 (N1785, N1760, N1338, N1272);
not NOT1 (N1786, N1782);
buf BUF1 (N1787, N1785);
and AND3 (N1788, N1777, N1646, N1459);
nor NOR2 (N1789, N1786, N71);
xor XOR2 (N1790, N1784, N1595);
not NOT1 (N1791, N1781);
or OR4 (N1792, N1783, N504, N669, N1278);
or OR4 (N1793, N1778, N1124, N320, N1651);
xor XOR2 (N1794, N1746, N160);
nand NAND4 (N1795, N1793, N715, N51, N1545);
xor XOR2 (N1796, N1787, N366);
xor XOR2 (N1797, N1792, N273);
and AND4 (N1798, N1790, N592, N1439, N543);
xor XOR2 (N1799, N1798, N1593);
buf BUF1 (N1800, N1799);
nor NOR3 (N1801, N1789, N553, N577);
and AND4 (N1802, N1795, N739, N753, N1344);
and AND2 (N1803, N1794, N1127);
xor XOR2 (N1804, N1802, N951);
not NOT1 (N1805, N1747);
nand NAND3 (N1806, N1801, N434, N115);
not NOT1 (N1807, N1776);
or OR3 (N1808, N1803, N1319, N1530);
and AND4 (N1809, N1791, N1322, N49, N1555);
not NOT1 (N1810, N1807);
buf BUF1 (N1811, N1797);
or OR4 (N1812, N1809, N382, N969, N928);
nand NAND3 (N1813, N1804, N1431, N662);
nor NOR3 (N1814, N1810, N1172, N798);
not NOT1 (N1815, N1812);
nor NOR3 (N1816, N1815, N964, N1641);
and AND4 (N1817, N1788, N1690, N1197, N1535);
nand NAND3 (N1818, N1817, N1178, N1464);
nor NOR4 (N1819, N1818, N237, N975, N1298);
nand NAND4 (N1820, N1819, N524, N975, N271);
xor XOR2 (N1821, N1800, N841);
or OR4 (N1822, N1821, N1227, N323, N1366);
and AND4 (N1823, N1822, N1568, N760, N730);
not NOT1 (N1824, N1808);
nand NAND2 (N1825, N1820, N1303);
and AND4 (N1826, N1824, N1358, N257, N221);
and AND2 (N1827, N1823, N114);
buf BUF1 (N1828, N1806);
nand NAND2 (N1829, N1796, N1522);
and AND3 (N1830, N1813, N177, N665);
xor XOR2 (N1831, N1828, N1533);
not NOT1 (N1832, N1825);
buf BUF1 (N1833, N1816);
not NOT1 (N1834, N1811);
or OR4 (N1835, N1826, N317, N1379, N1651);
nand NAND4 (N1836, N1829, N209, N634, N1598);
nor NOR3 (N1837, N1832, N878, N505);
xor XOR2 (N1838, N1836, N136);
nor NOR4 (N1839, N1827, N1389, N947, N1411);
not NOT1 (N1840, N1835);
not NOT1 (N1841, N1839);
nor NOR2 (N1842, N1805, N355);
or OR3 (N1843, N1830, N524, N1058);
nand NAND4 (N1844, N1834, N537, N260, N1705);
and AND2 (N1845, N1833, N638);
and AND4 (N1846, N1845, N227, N240, N503);
and AND3 (N1847, N1843, N118, N868);
or OR4 (N1848, N1837, N1304, N327, N1414);
buf BUF1 (N1849, N1841);
nor NOR3 (N1850, N1814, N1225, N423);
nand NAND3 (N1851, N1848, N524, N1639);
buf BUF1 (N1852, N1838);
nand NAND2 (N1853, N1840, N472);
and AND4 (N1854, N1844, N1128, N333, N425);
nor NOR4 (N1855, N1850, N31, N414, N1343);
buf BUF1 (N1856, N1842);
nand NAND4 (N1857, N1831, N1573, N377, N182);
or OR4 (N1858, N1851, N813, N564, N129);
xor XOR2 (N1859, N1856, N135);
xor XOR2 (N1860, N1857, N522);
xor XOR2 (N1861, N1853, N1344);
not NOT1 (N1862, N1847);
nand NAND3 (N1863, N1855, N1849, N667);
nand NAND2 (N1864, N1592, N992);
or OR3 (N1865, N1846, N1103, N624);
and AND4 (N1866, N1865, N1616, N321, N131);
and AND2 (N1867, N1864, N920);
and AND2 (N1868, N1858, N882);
nor NOR4 (N1869, N1863, N735, N24, N1118);
and AND2 (N1870, N1861, N352);
or OR2 (N1871, N1852, N1178);
nor NOR4 (N1872, N1868, N195, N835, N1789);
nor NOR4 (N1873, N1859, N1419, N298, N1293);
not NOT1 (N1874, N1871);
buf BUF1 (N1875, N1854);
buf BUF1 (N1876, N1860);
nor NOR4 (N1877, N1872, N1154, N1431, N323);
buf BUF1 (N1878, N1866);
xor XOR2 (N1879, N1862, N1194);
nor NOR4 (N1880, N1874, N1634, N1425, N879);
nor NOR4 (N1881, N1879, N304, N884, N84);
or OR3 (N1882, N1869, N733, N1727);
xor XOR2 (N1883, N1875, N365);
nand NAND3 (N1884, N1867, N670, N1721);
or OR4 (N1885, N1876, N495, N713, N115);
nand NAND4 (N1886, N1882, N766, N740, N1611);
not NOT1 (N1887, N1883);
nand NAND4 (N1888, N1877, N294, N863, N1334);
and AND4 (N1889, N1888, N1846, N1499, N1413);
nand NAND3 (N1890, N1884, N1188, N1837);
nor NOR2 (N1891, N1885, N1233);
and AND2 (N1892, N1887, N1061);
buf BUF1 (N1893, N1878);
or OR4 (N1894, N1892, N516, N1186, N180);
not NOT1 (N1895, N1880);
or OR2 (N1896, N1873, N1128);
or OR3 (N1897, N1881, N1420, N1546);
buf BUF1 (N1898, N1890);
nor NOR4 (N1899, N1897, N1165, N1868, N1017);
buf BUF1 (N1900, N1895);
xor XOR2 (N1901, N1896, N1582);
xor XOR2 (N1902, N1898, N899);
xor XOR2 (N1903, N1900, N217);
not NOT1 (N1904, N1891);
nor NOR4 (N1905, N1894, N516, N1885, N1598);
nand NAND2 (N1906, N1904, N1280);
nor NOR4 (N1907, N1902, N52, N743, N1278);
xor XOR2 (N1908, N1907, N483);
not NOT1 (N1909, N1886);
and AND2 (N1910, N1889, N185);
xor XOR2 (N1911, N1906, N960);
nor NOR4 (N1912, N1901, N1613, N1000, N1621);
nor NOR3 (N1913, N1870, N1215, N649);
not NOT1 (N1914, N1893);
and AND3 (N1915, N1914, N1384, N1458);
nand NAND3 (N1916, N1915, N1747, N1540);
nand NAND4 (N1917, N1913, N786, N1829, N1495);
xor XOR2 (N1918, N1903, N419);
nor NOR4 (N1919, N1908, N837, N887, N291);
and AND4 (N1920, N1918, N1688, N1128, N430);
xor XOR2 (N1921, N1919, N1412);
or OR4 (N1922, N1912, N401, N1540, N1716);
xor XOR2 (N1923, N1911, N1766);
nor NOR4 (N1924, N1905, N747, N912, N1073);
xor XOR2 (N1925, N1921, N144);
buf BUF1 (N1926, N1924);
not NOT1 (N1927, N1909);
and AND2 (N1928, N1916, N67);
xor XOR2 (N1929, N1927, N744);
not NOT1 (N1930, N1899);
nand NAND4 (N1931, N1929, N1868, N1799, N86);
nand NAND4 (N1932, N1910, N1881, N890, N185);
xor XOR2 (N1933, N1923, N257);
or OR2 (N1934, N1931, N720);
nand NAND3 (N1935, N1922, N1080, N1714);
not NOT1 (N1936, N1925);
or OR2 (N1937, N1933, N110);
not NOT1 (N1938, N1937);
or OR4 (N1939, N1936, N560, N1764, N1718);
nand NAND3 (N1940, N1928, N1168, N108);
not NOT1 (N1941, N1939);
nand NAND3 (N1942, N1934, N386, N1702);
nand NAND4 (N1943, N1917, N1451, N1405, N1766);
buf BUF1 (N1944, N1941);
buf BUF1 (N1945, N1932);
or OR4 (N1946, N1944, N1099, N346, N1590);
not NOT1 (N1947, N1946);
nor NOR2 (N1948, N1938, N1569);
nand NAND4 (N1949, N1948, N1203, N889, N1591);
not NOT1 (N1950, N1945);
buf BUF1 (N1951, N1943);
nor NOR3 (N1952, N1935, N1255, N1269);
and AND3 (N1953, N1920, N1807, N1720);
buf BUF1 (N1954, N1947);
xor XOR2 (N1955, N1952, N742);
and AND4 (N1956, N1954, N1362, N37, N1143);
xor XOR2 (N1957, N1949, N1088);
and AND2 (N1958, N1953, N242);
nor NOR2 (N1959, N1955, N348);
xor XOR2 (N1960, N1940, N1484);
nand NAND2 (N1961, N1926, N847);
and AND3 (N1962, N1956, N1692, N363);
buf BUF1 (N1963, N1962);
nor NOR2 (N1964, N1963, N1826);
not NOT1 (N1965, N1942);
and AND3 (N1966, N1964, N825, N143);
nand NAND4 (N1967, N1930, N1198, N1223, N865);
nand NAND3 (N1968, N1950, N569, N1667);
and AND2 (N1969, N1958, N373);
not NOT1 (N1970, N1968);
nand NAND3 (N1971, N1961, N1157, N1452);
not NOT1 (N1972, N1965);
buf BUF1 (N1973, N1971);
nand NAND4 (N1974, N1966, N320, N398, N1514);
or OR4 (N1975, N1967, N1650, N913, N1481);
not NOT1 (N1976, N1957);
nor NOR3 (N1977, N1970, N1066, N793);
nand NAND4 (N1978, N1959, N1490, N1910, N695);
xor XOR2 (N1979, N1978, N1644);
xor XOR2 (N1980, N1972, N1254);
xor XOR2 (N1981, N1977, N1655);
not NOT1 (N1982, N1980);
nand NAND3 (N1983, N1982, N795, N1026);
xor XOR2 (N1984, N1975, N714);
or OR2 (N1985, N1984, N1392);
or OR4 (N1986, N1979, N1409, N852, N908);
xor XOR2 (N1987, N1986, N1073);
nor NOR4 (N1988, N1973, N1511, N1457, N922);
or OR2 (N1989, N1974, N456);
or OR3 (N1990, N1976, N215, N1301);
not NOT1 (N1991, N1983);
not NOT1 (N1992, N1951);
nor NOR3 (N1993, N1992, N1655, N206);
xor XOR2 (N1994, N1987, N1903);
xor XOR2 (N1995, N1990, N1767);
buf BUF1 (N1996, N1995);
nor NOR3 (N1997, N1969, N900, N1648);
nand NAND2 (N1998, N1993, N933);
and AND2 (N1999, N1991, N1387);
and AND2 (N2000, N1999, N46);
buf BUF1 (N2001, N1989);
buf BUF1 (N2002, N1981);
xor XOR2 (N2003, N1994, N1641);
buf BUF1 (N2004, N1997);
nand NAND3 (N2005, N2004, N1467, N1033);
nand NAND2 (N2006, N1988, N856);
nand NAND4 (N2007, N1998, N1861, N1225, N573);
buf BUF1 (N2008, N1960);
not NOT1 (N2009, N2008);
buf BUF1 (N2010, N1985);
nor NOR4 (N2011, N2002, N719, N18, N275);
and AND3 (N2012, N2010, N906, N191);
xor XOR2 (N2013, N2000, N1287);
buf BUF1 (N2014, N2011);
or OR2 (N2015, N2013, N1138);
or OR3 (N2016, N2003, N729, N411);
nor NOR4 (N2017, N2007, N365, N1228, N637);
or OR2 (N2018, N2016, N40);
nand NAND3 (N2019, N2005, N888, N118);
not NOT1 (N2020, N2015);
buf BUF1 (N2021, N2018);
nand NAND2 (N2022, N2009, N1111);
or OR3 (N2023, N2014, N886, N1463);
nand NAND2 (N2024, N2020, N1408);
buf BUF1 (N2025, N2017);
xor XOR2 (N2026, N2022, N884);
and AND2 (N2027, N2019, N263);
or OR2 (N2028, N2012, N933);
and AND4 (N2029, N2006, N820, N910, N1616);
buf BUF1 (N2030, N2023);
not NOT1 (N2031, N2030);
nand NAND4 (N2032, N2001, N1064, N1503, N469);
not NOT1 (N2033, N2024);
buf BUF1 (N2034, N2025);
xor XOR2 (N2035, N2021, N1438);
xor XOR2 (N2036, N2031, N933);
nand NAND3 (N2037, N2032, N1327, N905);
and AND2 (N2038, N2036, N923);
nor NOR2 (N2039, N2035, N477);
nand NAND2 (N2040, N2034, N1527);
and AND2 (N2041, N2027, N1592);
or OR3 (N2042, N2029, N337, N1671);
nor NOR4 (N2043, N2041, N608, N477, N1766);
nand NAND4 (N2044, N2037, N1685, N1146, N1870);
xor XOR2 (N2045, N2026, N419);
nand NAND3 (N2046, N2045, N63, N1588);
nor NOR2 (N2047, N2046, N507);
nor NOR3 (N2048, N2033, N385, N192);
buf BUF1 (N2049, N2048);
xor XOR2 (N2050, N2028, N604);
xor XOR2 (N2051, N1996, N1341);
or OR4 (N2052, N2039, N318, N1566, N1652);
not NOT1 (N2053, N2038);
nand NAND2 (N2054, N2043, N811);
and AND4 (N2055, N2050, N1213, N1572, N1346);
not NOT1 (N2056, N2047);
buf BUF1 (N2057, N2044);
nand NAND4 (N2058, N2042, N162, N707, N791);
not NOT1 (N2059, N2055);
buf BUF1 (N2060, N2059);
not NOT1 (N2061, N2051);
nand NAND4 (N2062, N2049, N723, N612, N725);
or OR2 (N2063, N2058, N2022);
nor NOR4 (N2064, N2057, N1811, N782, N1711);
not NOT1 (N2065, N2060);
or OR2 (N2066, N2053, N1669);
nand NAND2 (N2067, N2064, N1943);
nand NAND4 (N2068, N2040, N503, N1356, N1094);
or OR2 (N2069, N2068, N1824);
not NOT1 (N2070, N2062);
not NOT1 (N2071, N2070);
nand NAND3 (N2072, N2069, N1421, N1163);
not NOT1 (N2073, N2067);
nand NAND2 (N2074, N2061, N1075);
nand NAND2 (N2075, N2066, N2044);
nor NOR3 (N2076, N2071, N2065, N64);
nand NAND3 (N2077, N1228, N2016, N167);
and AND3 (N2078, N2063, N850, N1499);
nor NOR3 (N2079, N2052, N370, N1909);
xor XOR2 (N2080, N2054, N2035);
and AND4 (N2081, N2076, N1218, N1334, N230);
xor XOR2 (N2082, N2080, N622);
and AND4 (N2083, N2073, N2040, N717, N2056);
not NOT1 (N2084, N380);
buf BUF1 (N2085, N2082);
nor NOR2 (N2086, N2078, N1474);
buf BUF1 (N2087, N2072);
not NOT1 (N2088, N2084);
nand NAND3 (N2089, N2081, N57, N1744);
nand NAND4 (N2090, N2083, N1310, N820, N1527);
xor XOR2 (N2091, N2079, N783);
nand NAND4 (N2092, N2087, N621, N1294, N1830);
buf BUF1 (N2093, N2092);
not NOT1 (N2094, N2085);
not NOT1 (N2095, N2075);
nor NOR3 (N2096, N2094, N1876, N656);
nor NOR4 (N2097, N2093, N1397, N1479, N42);
or OR3 (N2098, N2091, N1356, N1481);
nand NAND4 (N2099, N2090, N345, N81, N1356);
and AND4 (N2100, N2099, N2, N1378, N2022);
buf BUF1 (N2101, N2096);
and AND3 (N2102, N2098, N963, N1424);
nand NAND2 (N2103, N2100, N527);
xor XOR2 (N2104, N2086, N1287);
nor NOR3 (N2105, N2095, N2002, N865);
buf BUF1 (N2106, N2074);
or OR2 (N2107, N2104, N703);
nor NOR4 (N2108, N2089, N1194, N1476, N1574);
or OR3 (N2109, N2106, N1229, N1461);
xor XOR2 (N2110, N2077, N1446);
xor XOR2 (N2111, N2103, N1671);
nand NAND2 (N2112, N2101, N402);
xor XOR2 (N2113, N2110, N1227);
xor XOR2 (N2114, N2112, N1583);
nand NAND3 (N2115, N2105, N822, N600);
nor NOR3 (N2116, N2102, N1205, N657);
and AND4 (N2117, N2097, N832, N1818, N1739);
xor XOR2 (N2118, N2111, N239);
buf BUF1 (N2119, N2113);
nand NAND4 (N2120, N2108, N623, N2040, N1882);
xor XOR2 (N2121, N2114, N200);
buf BUF1 (N2122, N2120);
nor NOR3 (N2123, N2119, N1302, N1545);
and AND4 (N2124, N2115, N1511, N525, N117);
nand NAND2 (N2125, N2116, N736);
nand NAND3 (N2126, N2125, N1922, N486);
nand NAND4 (N2127, N2088, N789, N401, N1787);
nand NAND3 (N2128, N2123, N2046, N295);
xor XOR2 (N2129, N2122, N1627);
nor NOR4 (N2130, N2126, N1041, N1521, N1127);
and AND2 (N2131, N2129, N1161);
not NOT1 (N2132, N2130);
xor XOR2 (N2133, N2127, N598);
xor XOR2 (N2134, N2121, N114);
nand NAND4 (N2135, N2117, N788, N1186, N642);
or OR4 (N2136, N2131, N1317, N1257, N898);
or OR3 (N2137, N2135, N359, N66);
not NOT1 (N2138, N2132);
not NOT1 (N2139, N2107);
buf BUF1 (N2140, N2124);
and AND3 (N2141, N2138, N1680, N1908);
nand NAND4 (N2142, N2134, N2083, N128, N745);
xor XOR2 (N2143, N2142, N614);
nor NOR2 (N2144, N2133, N382);
xor XOR2 (N2145, N2140, N1012);
and AND4 (N2146, N2109, N1163, N2100, N1948);
nor NOR2 (N2147, N2118, N54);
xor XOR2 (N2148, N2141, N1648);
xor XOR2 (N2149, N2145, N1642);
and AND3 (N2150, N2144, N1360, N874);
nor NOR4 (N2151, N2149, N1854, N821, N556);
nor NOR3 (N2152, N2128, N1372, N1557);
or OR3 (N2153, N2147, N1177, N1415);
xor XOR2 (N2154, N2146, N1471);
xor XOR2 (N2155, N2153, N199);
and AND2 (N2156, N2151, N855);
not NOT1 (N2157, N2148);
buf BUF1 (N2158, N2152);
nor NOR2 (N2159, N2156, N696);
and AND3 (N2160, N2139, N622, N1551);
not NOT1 (N2161, N2136);
xor XOR2 (N2162, N2143, N10);
nor NOR2 (N2163, N2159, N850);
buf BUF1 (N2164, N2155);
nor NOR2 (N2165, N2158, N294);
xor XOR2 (N2166, N2150, N1579);
not NOT1 (N2167, N2160);
xor XOR2 (N2168, N2164, N685);
or OR3 (N2169, N2168, N1455, N701);
and AND2 (N2170, N2161, N519);
buf BUF1 (N2171, N2163);
nor NOR2 (N2172, N2137, N2118);
buf BUF1 (N2173, N2169);
buf BUF1 (N2174, N2154);
or OR4 (N2175, N2170, N951, N1662, N2157);
and AND3 (N2176, N221, N549, N1731);
nor NOR2 (N2177, N2173, N816);
or OR4 (N2178, N2171, N1024, N488, N180);
xor XOR2 (N2179, N2175, N641);
or OR2 (N2180, N2177, N1320);
buf BUF1 (N2181, N2180);
or OR3 (N2182, N2178, N861, N2076);
buf BUF1 (N2183, N2165);
xor XOR2 (N2184, N2162, N1918);
not NOT1 (N2185, N2167);
xor XOR2 (N2186, N2182, N14);
and AND4 (N2187, N2172, N406, N847, N720);
nand NAND4 (N2188, N2184, N1094, N1105, N1457);
nand NAND2 (N2189, N2166, N2127);
and AND3 (N2190, N2183, N2153, N201);
xor XOR2 (N2191, N2174, N481);
nand NAND3 (N2192, N2190, N879, N1420);
xor XOR2 (N2193, N2187, N831);
or OR2 (N2194, N2179, N1149);
nor NOR3 (N2195, N2194, N242, N66);
and AND2 (N2196, N2188, N1813);
nand NAND3 (N2197, N2193, N1278, N470);
buf BUF1 (N2198, N2191);
and AND2 (N2199, N2198, N651);
and AND3 (N2200, N2181, N1078, N246);
nand NAND2 (N2201, N2195, N1515);
or OR2 (N2202, N2201, N1694);
and AND2 (N2203, N2202, N2086);
not NOT1 (N2204, N2189);
xor XOR2 (N2205, N2176, N112);
nor NOR3 (N2206, N2185, N1979, N145);
buf BUF1 (N2207, N2199);
xor XOR2 (N2208, N2205, N444);
not NOT1 (N2209, N2207);
nand NAND3 (N2210, N2196, N881, N1893);
xor XOR2 (N2211, N2197, N1287);
xor XOR2 (N2212, N2210, N2002);
nor NOR3 (N2213, N2212, N811, N859);
buf BUF1 (N2214, N2200);
not NOT1 (N2215, N2206);
not NOT1 (N2216, N2204);
or OR3 (N2217, N2213, N891, N870);
buf BUF1 (N2218, N2186);
not NOT1 (N2219, N2214);
nor NOR3 (N2220, N2203, N1222, N512);
not NOT1 (N2221, N2217);
nor NOR2 (N2222, N2216, N1552);
not NOT1 (N2223, N2219);
buf BUF1 (N2224, N2209);
xor XOR2 (N2225, N2218, N502);
and AND2 (N2226, N2224, N1405);
or OR3 (N2227, N2220, N1599, N2099);
not NOT1 (N2228, N2222);
nor NOR3 (N2229, N2225, N608, N2024);
xor XOR2 (N2230, N2227, N2127);
not NOT1 (N2231, N2228);
not NOT1 (N2232, N2215);
not NOT1 (N2233, N2232);
buf BUF1 (N2234, N2211);
not NOT1 (N2235, N2229);
not NOT1 (N2236, N2231);
xor XOR2 (N2237, N2236, N819);
or OR4 (N2238, N2223, N797, N1375, N1386);
xor XOR2 (N2239, N2235, N1075);
not NOT1 (N2240, N2234);
not NOT1 (N2241, N2230);
buf BUF1 (N2242, N2221);
buf BUF1 (N2243, N2239);
and AND2 (N2244, N2233, N1067);
and AND2 (N2245, N2241, N874);
xor XOR2 (N2246, N2208, N489);
xor XOR2 (N2247, N2243, N1414);
xor XOR2 (N2248, N2226, N374);
xor XOR2 (N2249, N2240, N1561);
or OR4 (N2250, N2237, N1735, N543, N621);
nand NAND3 (N2251, N2250, N544, N919);
or OR4 (N2252, N2247, N1303, N510, N487);
or OR3 (N2253, N2244, N2095, N925);
nand NAND4 (N2254, N2238, N1709, N1780, N1804);
or OR3 (N2255, N2248, N1930, N4);
or OR2 (N2256, N2253, N341);
buf BUF1 (N2257, N2252);
or OR4 (N2258, N2249, N1842, N867, N388);
nor NOR3 (N2259, N2257, N1268, N2163);
xor XOR2 (N2260, N2256, N981);
nand NAND3 (N2261, N2251, N2083, N21);
and AND3 (N2262, N2254, N1043, N2236);
xor XOR2 (N2263, N2261, N234);
buf BUF1 (N2264, N2262);
or OR4 (N2265, N2245, N1013, N2236, N2212);
nand NAND2 (N2266, N2246, N1162);
buf BUF1 (N2267, N2263);
nor NOR2 (N2268, N2192, N1254);
nand NAND4 (N2269, N2266, N978, N191, N1273);
not NOT1 (N2270, N2268);
or OR4 (N2271, N2260, N1577, N2139, N813);
nand NAND2 (N2272, N2255, N198);
nand NAND4 (N2273, N2272, N408, N1742, N1897);
or OR3 (N2274, N2267, N1694, N1109);
xor XOR2 (N2275, N2258, N1824);
buf BUF1 (N2276, N2275);
buf BUF1 (N2277, N2265);
xor XOR2 (N2278, N2277, N231);
not NOT1 (N2279, N2270);
buf BUF1 (N2280, N2279);
xor XOR2 (N2281, N2242, N1665);
or OR3 (N2282, N2280, N1038, N2080);
not NOT1 (N2283, N2274);
and AND2 (N2284, N2281, N574);
nor NOR2 (N2285, N2271, N733);
and AND3 (N2286, N2276, N520, N1746);
and AND3 (N2287, N2259, N1936, N505);
or OR3 (N2288, N2283, N1981, N153);
nor NOR3 (N2289, N2278, N2024, N2066);
and AND3 (N2290, N2282, N1645, N960);
xor XOR2 (N2291, N2284, N1975);
and AND4 (N2292, N2269, N311, N1160, N1390);
and AND4 (N2293, N2287, N239, N1331, N973);
nor NOR4 (N2294, N2290, N1978, N1263, N1886);
xor XOR2 (N2295, N2289, N421);
or OR2 (N2296, N2291, N1311);
nor NOR2 (N2297, N2293, N1076);
xor XOR2 (N2298, N2292, N1009);
nand NAND2 (N2299, N2286, N1995);
nand NAND4 (N2300, N2298, N1796, N1940, N102);
or OR2 (N2301, N2299, N460);
nor NOR4 (N2302, N2300, N2038, N448, N1304);
or OR4 (N2303, N2296, N1689, N1374, N115);
nor NOR3 (N2304, N2303, N194, N686);
or OR3 (N2305, N2288, N70, N237);
nor NOR2 (N2306, N2273, N1851);
or OR3 (N2307, N2294, N420, N1279);
nand NAND3 (N2308, N2285, N206, N1463);
and AND3 (N2309, N2302, N236, N1122);
buf BUF1 (N2310, N2305);
xor XOR2 (N2311, N2301, N1885);
xor XOR2 (N2312, N2264, N77);
not NOT1 (N2313, N2304);
and AND4 (N2314, N2308, N416, N2103, N773);
or OR3 (N2315, N2297, N28, N2038);
xor XOR2 (N2316, N2306, N363);
and AND4 (N2317, N2295, N471, N1325, N1490);
xor XOR2 (N2318, N2317, N270);
buf BUF1 (N2319, N2314);
and AND4 (N2320, N2311, N772, N1272, N2131);
nand NAND4 (N2321, N2320, N743, N489, N385);
nand NAND3 (N2322, N2319, N1351, N1598);
buf BUF1 (N2323, N2309);
xor XOR2 (N2324, N2318, N1812);
or OR3 (N2325, N2316, N1885, N240);
or OR4 (N2326, N2315, N658, N1998, N500);
buf BUF1 (N2327, N2321);
and AND2 (N2328, N2323, N972);
or OR4 (N2329, N2324, N1401, N84, N1367);
nand NAND2 (N2330, N2325, N1279);
or OR4 (N2331, N2312, N433, N1300, N16);
not NOT1 (N2332, N2326);
or OR2 (N2333, N2330, N1332);
or OR3 (N2334, N2310, N1698, N2046);
nor NOR4 (N2335, N2322, N350, N1956, N389);
nor NOR4 (N2336, N2329, N93, N1921, N587);
buf BUF1 (N2337, N2331);
buf BUF1 (N2338, N2335);
or OR3 (N2339, N2334, N971, N1417);
not NOT1 (N2340, N2339);
and AND4 (N2341, N2327, N1713, N1137, N319);
not NOT1 (N2342, N2338);
not NOT1 (N2343, N2328);
or OR2 (N2344, N2340, N938);
xor XOR2 (N2345, N2336, N981);
xor XOR2 (N2346, N2333, N2120);
nand NAND4 (N2347, N2307, N1664, N771, N2338);
buf BUF1 (N2348, N2332);
buf BUF1 (N2349, N2313);
nand NAND3 (N2350, N2337, N1927, N1492);
buf BUF1 (N2351, N2344);
nand NAND3 (N2352, N2343, N2235, N1143);
not NOT1 (N2353, N2350);
nand NAND4 (N2354, N2341, N2115, N1863, N756);
or OR4 (N2355, N2346, N378, N1633, N2229);
and AND4 (N2356, N2348, N2233, N1616, N1485);
and AND3 (N2357, N2354, N1422, N1362);
not NOT1 (N2358, N2355);
nand NAND4 (N2359, N2347, N1125, N763, N1971);
xor XOR2 (N2360, N2359, N1143);
nor NOR2 (N2361, N2342, N863);
nor NOR2 (N2362, N2352, N1783);
nor NOR3 (N2363, N2358, N838, N549);
nand NAND4 (N2364, N2363, N879, N1330, N1140);
buf BUF1 (N2365, N2345);
nor NOR4 (N2366, N2357, N1336, N1249, N1309);
nand NAND2 (N2367, N2366, N1884);
buf BUF1 (N2368, N2367);
or OR2 (N2369, N2362, N408);
or OR4 (N2370, N2364, N506, N1645, N2335);
nand NAND2 (N2371, N2365, N351);
nand NAND4 (N2372, N2369, N510, N1419, N1956);
and AND3 (N2373, N2353, N589, N1014);
not NOT1 (N2374, N2360);
and AND4 (N2375, N2356, N745, N200, N922);
or OR3 (N2376, N2351, N2340, N243);
nor NOR3 (N2377, N2349, N1801, N424);
and AND4 (N2378, N2374, N429, N100, N2167);
or OR4 (N2379, N2361, N26, N831, N1718);
nor NOR4 (N2380, N2377, N1626, N322, N303);
and AND2 (N2381, N2372, N1520);
not NOT1 (N2382, N2370);
xor XOR2 (N2383, N2368, N356);
or OR2 (N2384, N2380, N723);
nand NAND2 (N2385, N2376, N1165);
nor NOR4 (N2386, N2381, N1938, N1807, N2312);
xor XOR2 (N2387, N2379, N1978);
nand NAND3 (N2388, N2371, N914, N1748);
buf BUF1 (N2389, N2386);
not NOT1 (N2390, N2383);
and AND3 (N2391, N2378, N1377, N1067);
nor NOR2 (N2392, N2390, N418);
nor NOR4 (N2393, N2375, N263, N2179, N2337);
or OR2 (N2394, N2393, N525);
not NOT1 (N2395, N2382);
nor NOR3 (N2396, N2373, N355, N1291);
nor NOR3 (N2397, N2387, N199, N2388);
nand NAND3 (N2398, N1469, N241, N1002);
xor XOR2 (N2399, N2397, N1066);
or OR2 (N2400, N2395, N635);
nor NOR3 (N2401, N2384, N2346, N1212);
and AND4 (N2402, N2394, N354, N1826, N222);
not NOT1 (N2403, N2398);
nor NOR2 (N2404, N2402, N1590);
or OR2 (N2405, N2392, N391);
xor XOR2 (N2406, N2404, N1013);
nand NAND2 (N2407, N2391, N878);
and AND4 (N2408, N2407, N2092, N1404, N1558);
nor NOR3 (N2409, N2406, N1892, N2106);
buf BUF1 (N2410, N2396);
nand NAND4 (N2411, N2399, N739, N793, N591);
xor XOR2 (N2412, N2408, N1307);
buf BUF1 (N2413, N2412);
buf BUF1 (N2414, N2400);
xor XOR2 (N2415, N2413, N2239);
nor NOR2 (N2416, N2385, N2342);
not NOT1 (N2417, N2415);
not NOT1 (N2418, N2409);
nand NAND3 (N2419, N2401, N157, N2224);
nor NOR3 (N2420, N2403, N375, N2175);
nor NOR4 (N2421, N2414, N1042, N1107, N974);
nand NAND2 (N2422, N2416, N1989);
and AND2 (N2423, N2410, N1929);
and AND2 (N2424, N2411, N1171);
nand NAND4 (N2425, N2421, N1857, N85, N158);
or OR4 (N2426, N2425, N90, N716, N56);
or OR3 (N2427, N2419, N2024, N687);
or OR4 (N2428, N2389, N384, N1478, N532);
and AND4 (N2429, N2426, N581, N1823, N424);
not NOT1 (N2430, N2423);
not NOT1 (N2431, N2405);
or OR2 (N2432, N2417, N1850);
nand NAND4 (N2433, N2428, N856, N1690, N2006);
nand NAND3 (N2434, N2422, N1331, N921);
xor XOR2 (N2435, N2424, N2251);
and AND3 (N2436, N2430, N1917, N375);
or OR3 (N2437, N2433, N672, N1063);
nand NAND2 (N2438, N2435, N1671);
buf BUF1 (N2439, N2418);
nand NAND3 (N2440, N2431, N2249, N1895);
nor NOR4 (N2441, N2420, N1593, N2009, N1400);
nand NAND2 (N2442, N2439, N1052);
or OR4 (N2443, N2442, N1609, N2046, N2324);
or OR2 (N2444, N2440, N849);
or OR4 (N2445, N2438, N2051, N1470, N445);
or OR4 (N2446, N2441, N526, N980, N794);
buf BUF1 (N2447, N2444);
nor NOR3 (N2448, N2432, N2372, N1896);
not NOT1 (N2449, N2436);
nor NOR3 (N2450, N2448, N432, N677);
not NOT1 (N2451, N2437);
buf BUF1 (N2452, N2445);
not NOT1 (N2453, N2449);
xor XOR2 (N2454, N2446, N1689);
nor NOR3 (N2455, N2443, N1796, N97);
xor XOR2 (N2456, N2429, N916);
not NOT1 (N2457, N2434);
not NOT1 (N2458, N2457);
xor XOR2 (N2459, N2456, N103);
and AND2 (N2460, N2458, N97);
or OR3 (N2461, N2450, N76, N808);
not NOT1 (N2462, N2453);
and AND3 (N2463, N2461, N1453, N1261);
not NOT1 (N2464, N2463);
or OR2 (N2465, N2459, N208);
nor NOR2 (N2466, N2452, N56);
or OR2 (N2467, N2464, N1348);
or OR4 (N2468, N2467, N2354, N387, N2150);
not NOT1 (N2469, N2468);
nand NAND3 (N2470, N2447, N1433, N1319);
and AND2 (N2471, N2454, N936);
and AND2 (N2472, N2469, N225);
xor XOR2 (N2473, N2470, N1910);
and AND4 (N2474, N2460, N1449, N180, N2134);
nand NAND2 (N2475, N2462, N2242);
or OR3 (N2476, N2474, N438, N732);
xor XOR2 (N2477, N2451, N2332);
not NOT1 (N2478, N2427);
nand NAND3 (N2479, N2465, N1008, N894);
nand NAND3 (N2480, N2477, N1141, N1800);
nand NAND4 (N2481, N2473, N1746, N766, N2104);
nand NAND3 (N2482, N2455, N1969, N882);
nor NOR4 (N2483, N2481, N2479, N1854, N1718);
and AND3 (N2484, N1140, N949, N1908);
and AND2 (N2485, N2475, N1010);
xor XOR2 (N2486, N2466, N1411);
not NOT1 (N2487, N2471);
and AND2 (N2488, N2478, N2411);
buf BUF1 (N2489, N2484);
nor NOR4 (N2490, N2488, N1258, N1702, N2221);
and AND4 (N2491, N2476, N2163, N2176, N1697);
and AND2 (N2492, N2491, N2402);
xor XOR2 (N2493, N2480, N723);
not NOT1 (N2494, N2489);
or OR2 (N2495, N2482, N1269);
nand NAND3 (N2496, N2490, N1164, N2315);
nand NAND3 (N2497, N2496, N11, N451);
and AND2 (N2498, N2483, N2378);
xor XOR2 (N2499, N2497, N2436);
nor NOR4 (N2500, N2487, N1296, N847, N1604);
xor XOR2 (N2501, N2495, N1937);
nor NOR3 (N2502, N2486, N213, N228);
nand NAND2 (N2503, N2502, N593);
nor NOR3 (N2504, N2499, N1206, N374);
or OR3 (N2505, N2501, N2495, N2149);
or OR2 (N2506, N2494, N207);
not NOT1 (N2507, N2498);
buf BUF1 (N2508, N2485);
not NOT1 (N2509, N2492);
buf BUF1 (N2510, N2500);
nand NAND3 (N2511, N2506, N217, N2426);
not NOT1 (N2512, N2472);
or OR3 (N2513, N2511, N2224, N2284);
not NOT1 (N2514, N2510);
and AND2 (N2515, N2513, N2408);
nor NOR3 (N2516, N2503, N1509, N757);
and AND2 (N2517, N2507, N2107);
and AND4 (N2518, N2508, N702, N830, N2126);
nor NOR3 (N2519, N2516, N1417, N2235);
nor NOR2 (N2520, N2493, N1895);
not NOT1 (N2521, N2519);
not NOT1 (N2522, N2515);
nor NOR4 (N2523, N2514, N76, N1905, N454);
and AND4 (N2524, N2505, N2354, N1036, N94);
not NOT1 (N2525, N2518);
not NOT1 (N2526, N2525);
xor XOR2 (N2527, N2522, N522);
not NOT1 (N2528, N2521);
nor NOR3 (N2529, N2526, N1805, N1945);
buf BUF1 (N2530, N2524);
nand NAND3 (N2531, N2528, N1113, N957);
xor XOR2 (N2532, N2504, N2356);
nor NOR2 (N2533, N2517, N1232);
nor NOR4 (N2534, N2529, N1741, N1749, N1465);
nor NOR4 (N2535, N2531, N1999, N416, N2115);
not NOT1 (N2536, N2534);
nor NOR2 (N2537, N2520, N547);
nand NAND3 (N2538, N2533, N2408, N2125);
and AND2 (N2539, N2537, N2485);
buf BUF1 (N2540, N2539);
xor XOR2 (N2541, N2538, N2469);
nand NAND4 (N2542, N2527, N282, N2441, N1675);
and AND3 (N2543, N2523, N1519, N2231);
buf BUF1 (N2544, N2509);
buf BUF1 (N2545, N2544);
and AND2 (N2546, N2543, N382);
xor XOR2 (N2547, N2541, N544);
and AND2 (N2548, N2542, N1343);
not NOT1 (N2549, N2536);
or OR4 (N2550, N2540, N2336, N474, N1442);
not NOT1 (N2551, N2548);
not NOT1 (N2552, N2550);
not NOT1 (N2553, N2552);
or OR2 (N2554, N2547, N2391);
or OR3 (N2555, N2535, N1160, N420);
buf BUF1 (N2556, N2546);
nor NOR2 (N2557, N2530, N275);
buf BUF1 (N2558, N2512);
not NOT1 (N2559, N2549);
buf BUF1 (N2560, N2551);
buf BUF1 (N2561, N2558);
buf BUF1 (N2562, N2555);
not NOT1 (N2563, N2554);
nand NAND3 (N2564, N2562, N937, N1115);
nor NOR4 (N2565, N2532, N2331, N1187, N1318);
nor NOR4 (N2566, N2553, N1852, N1719, N1856);
nand NAND3 (N2567, N2564, N922, N1036);
or OR2 (N2568, N2560, N1070);
or OR3 (N2569, N2565, N1144, N1765);
and AND4 (N2570, N2561, N32, N130, N2307);
nor NOR3 (N2571, N2556, N345, N456);
xor XOR2 (N2572, N2563, N2294);
nor NOR2 (N2573, N2572, N894);
xor XOR2 (N2574, N2571, N1814);
not NOT1 (N2575, N2570);
buf BUF1 (N2576, N2574);
nand NAND2 (N2577, N2566, N1431);
nand NAND2 (N2578, N2575, N516);
xor XOR2 (N2579, N2559, N939);
xor XOR2 (N2580, N2569, N701);
or OR4 (N2581, N2567, N941, N686, N643);
and AND2 (N2582, N2573, N912);
xor XOR2 (N2583, N2568, N1362);
and AND4 (N2584, N2583, N2355, N1275, N45);
not NOT1 (N2585, N2545);
xor XOR2 (N2586, N2576, N1653);
nor NOR3 (N2587, N2557, N1164, N51);
xor XOR2 (N2588, N2580, N229);
and AND2 (N2589, N2577, N1714);
and AND4 (N2590, N2585, N563, N1898, N2392);
nand NAND2 (N2591, N2589, N2506);
not NOT1 (N2592, N2587);
or OR3 (N2593, N2586, N2166, N822);
or OR4 (N2594, N2591, N2229, N1544, N1012);
xor XOR2 (N2595, N2584, N1638);
nor NOR3 (N2596, N2590, N922, N2519);
xor XOR2 (N2597, N2596, N648);
and AND2 (N2598, N2593, N2245);
and AND4 (N2599, N2594, N2047, N1455, N1728);
not NOT1 (N2600, N2581);
buf BUF1 (N2601, N2578);
not NOT1 (N2602, N2597);
nor NOR3 (N2603, N2588, N1742, N1816);
and AND4 (N2604, N2579, N1151, N828, N2500);
not NOT1 (N2605, N2604);
or OR2 (N2606, N2595, N2016);
or OR2 (N2607, N2600, N1376);
buf BUF1 (N2608, N2602);
buf BUF1 (N2609, N2605);
xor XOR2 (N2610, N2607, N213);
nand NAND3 (N2611, N2598, N47, N703);
nor NOR4 (N2612, N2582, N146, N221, N359);
xor XOR2 (N2613, N2603, N331);
xor XOR2 (N2614, N2610, N2376);
or OR2 (N2615, N2613, N718);
or OR3 (N2616, N2608, N49, N803);
nor NOR2 (N2617, N2601, N1570);
nand NAND4 (N2618, N2617, N574, N2549, N697);
buf BUF1 (N2619, N2592);
not NOT1 (N2620, N2606);
and AND2 (N2621, N2609, N1422);
nand NAND3 (N2622, N2599, N658, N2499);
nand NAND4 (N2623, N2611, N2157, N1095, N602);
buf BUF1 (N2624, N2615);
nor NOR4 (N2625, N2619, N712, N1539, N916);
xor XOR2 (N2626, N2612, N1018);
and AND4 (N2627, N2614, N1702, N1633, N879);
xor XOR2 (N2628, N2626, N1828);
not NOT1 (N2629, N2627);
or OR2 (N2630, N2629, N2199);
and AND4 (N2631, N2628, N2230, N2187, N54);
buf BUF1 (N2632, N2630);
nor NOR2 (N2633, N2622, N1376);
and AND3 (N2634, N2618, N170, N706);
xor XOR2 (N2635, N2625, N484);
buf BUF1 (N2636, N2620);
xor XOR2 (N2637, N2636, N2531);
buf BUF1 (N2638, N2634);
and AND2 (N2639, N2616, N1959);
or OR3 (N2640, N2624, N804, N1651);
nor NOR2 (N2641, N2632, N1391);
not NOT1 (N2642, N2635);
buf BUF1 (N2643, N2638);
or OR3 (N2644, N2631, N1134, N1341);
or OR2 (N2645, N2641, N1215);
nor NOR3 (N2646, N2621, N1109, N964);
not NOT1 (N2647, N2637);
nand NAND4 (N2648, N2640, N2441, N1327, N205);
nor NOR2 (N2649, N2623, N1913);
nand NAND2 (N2650, N2642, N1562);
nand NAND3 (N2651, N2648, N2378, N112);
buf BUF1 (N2652, N2633);
nand NAND4 (N2653, N2650, N1414, N1831, N349);
or OR2 (N2654, N2649, N1061);
buf BUF1 (N2655, N2652);
or OR2 (N2656, N2644, N249);
or OR3 (N2657, N2654, N784, N1441);
xor XOR2 (N2658, N2656, N1574);
and AND4 (N2659, N2651, N1089, N456, N2242);
nand NAND3 (N2660, N2646, N300, N1281);
and AND3 (N2661, N2660, N675, N2124);
not NOT1 (N2662, N2661);
or OR3 (N2663, N2653, N2551, N763);
or OR3 (N2664, N2639, N2283, N1130);
nor NOR4 (N2665, N2658, N2167, N946, N409);
nand NAND2 (N2666, N2655, N2557);
nand NAND3 (N2667, N2663, N2006, N2183);
nor NOR4 (N2668, N2647, N1561, N1749, N592);
not NOT1 (N2669, N2643);
nor NOR2 (N2670, N2659, N1298);
xor XOR2 (N2671, N2669, N2574);
not NOT1 (N2672, N2668);
nand NAND3 (N2673, N2666, N687, N1312);
buf BUF1 (N2674, N2657);
not NOT1 (N2675, N2662);
xor XOR2 (N2676, N2664, N1598);
nor NOR4 (N2677, N2673, N1983, N1213, N1697);
or OR3 (N2678, N2675, N2342, N1782);
buf BUF1 (N2679, N2667);
nand NAND4 (N2680, N2678, N1201, N1723, N759);
buf BUF1 (N2681, N2676);
or OR4 (N2682, N2680, N1921, N1968, N738);
nor NOR4 (N2683, N2672, N2119, N2397, N509);
xor XOR2 (N2684, N2645, N1349);
and AND2 (N2685, N2670, N145);
and AND3 (N2686, N2671, N2401, N1788);
or OR4 (N2687, N2679, N2542, N1256, N2670);
nor NOR3 (N2688, N2683, N1308, N1892);
buf BUF1 (N2689, N2686);
nand NAND4 (N2690, N2685, N2470, N1358, N918);
buf BUF1 (N2691, N2689);
and AND4 (N2692, N2691, N2132, N1916, N129);
not NOT1 (N2693, N2665);
not NOT1 (N2694, N2677);
or OR4 (N2695, N2688, N2271, N1651, N249);
buf BUF1 (N2696, N2694);
or OR4 (N2697, N2693, N2313, N2022, N2123);
nor NOR2 (N2698, N2692, N1350);
and AND2 (N2699, N2697, N2463);
buf BUF1 (N2700, N2674);
nor NOR4 (N2701, N2690, N1096, N347, N869);
nor NOR3 (N2702, N2701, N374, N1447);
not NOT1 (N2703, N2695);
and AND3 (N2704, N2700, N416, N2098);
not NOT1 (N2705, N2687);
nor NOR3 (N2706, N2703, N1411, N2403);
nor NOR4 (N2707, N2704, N1840, N2247, N1011);
xor XOR2 (N2708, N2705, N2215);
not NOT1 (N2709, N2682);
not NOT1 (N2710, N2709);
or OR4 (N2711, N2708, N481, N833, N2535);
or OR3 (N2712, N2699, N2110, N509);
nand NAND3 (N2713, N2707, N1007, N2464);
not NOT1 (N2714, N2706);
not NOT1 (N2715, N2713);
not NOT1 (N2716, N2712);
nor NOR4 (N2717, N2698, N1342, N698, N654);
xor XOR2 (N2718, N2714, N1125);
nor NOR3 (N2719, N2684, N2656, N1156);
not NOT1 (N2720, N2681);
not NOT1 (N2721, N2711);
nor NOR3 (N2722, N2715, N786, N1597);
nand NAND2 (N2723, N2702, N759);
xor XOR2 (N2724, N2718, N2537);
and AND3 (N2725, N2716, N465, N1038);
and AND3 (N2726, N2725, N1649, N1881);
nor NOR3 (N2727, N2722, N1519, N1989);
nand NAND2 (N2728, N2696, N1728);
xor XOR2 (N2729, N2719, N1879);
or OR3 (N2730, N2723, N1354, N995);
or OR4 (N2731, N2728, N1229, N1302, N1837);
buf BUF1 (N2732, N2729);
nand NAND4 (N2733, N2727, N52, N1769, N1003);
and AND3 (N2734, N2732, N1381, N2683);
nand NAND2 (N2735, N2724, N1662);
nor NOR2 (N2736, N2721, N2278);
or OR4 (N2737, N2720, N640, N2712, N1861);
nand NAND4 (N2738, N2735, N2007, N2535, N2507);
xor XOR2 (N2739, N2734, N1203);
nand NAND4 (N2740, N2733, N565, N1801, N277);
not NOT1 (N2741, N2717);
nor NOR3 (N2742, N2736, N1374, N1202);
xor XOR2 (N2743, N2737, N942);
nor NOR3 (N2744, N2742, N521, N2203);
buf BUF1 (N2745, N2731);
nand NAND4 (N2746, N2741, N728, N1800, N1235);
nor NOR4 (N2747, N2710, N397, N2452, N2069);
xor XOR2 (N2748, N2747, N397);
xor XOR2 (N2749, N2743, N229);
and AND2 (N2750, N2746, N2233);
nor NOR4 (N2751, N2745, N2196, N710, N101);
or OR4 (N2752, N2739, N2225, N1088, N1313);
xor XOR2 (N2753, N2730, N2365);
not NOT1 (N2754, N2738);
nand NAND2 (N2755, N2753, N2245);
buf BUF1 (N2756, N2744);
buf BUF1 (N2757, N2754);
and AND4 (N2758, N2740, N2433, N1619, N90);
not NOT1 (N2759, N2758);
xor XOR2 (N2760, N2756, N689);
or OR3 (N2761, N2760, N409, N2013);
xor XOR2 (N2762, N2751, N1321);
buf BUF1 (N2763, N2748);
or OR3 (N2764, N2750, N841, N1660);
buf BUF1 (N2765, N2726);
buf BUF1 (N2766, N2755);
not NOT1 (N2767, N2752);
or OR4 (N2768, N2757, N1175, N2749, N2335);
buf BUF1 (N2769, N1362);
or OR3 (N2770, N2769, N596, N2292);
buf BUF1 (N2771, N2759);
xor XOR2 (N2772, N2765, N1929);
or OR4 (N2773, N2766, N1598, N269, N386);
buf BUF1 (N2774, N2772);
nand NAND2 (N2775, N2764, N1459);
nor NOR2 (N2776, N2761, N2725);
buf BUF1 (N2777, N2763);
nor NOR3 (N2778, N2775, N331, N1062);
buf BUF1 (N2779, N2773);
and AND4 (N2780, N2774, N1901, N1053, N999);
and AND3 (N2781, N2780, N1509, N329);
nand NAND2 (N2782, N2777, N2275);
and AND2 (N2783, N2770, N493);
nand NAND2 (N2784, N2783, N1293);
not NOT1 (N2785, N2762);
and AND4 (N2786, N2781, N2526, N1802, N44);
and AND4 (N2787, N2784, N1632, N474, N130);
or OR4 (N2788, N2771, N1675, N1717, N191);
nand NAND3 (N2789, N2787, N2178, N949);
nor NOR3 (N2790, N2768, N2169, N941);
buf BUF1 (N2791, N2779);
not NOT1 (N2792, N2788);
not NOT1 (N2793, N2778);
nand NAND2 (N2794, N2789, N1736);
not NOT1 (N2795, N2767);
xor XOR2 (N2796, N2794, N638);
nor NOR3 (N2797, N2776, N2590, N1335);
buf BUF1 (N2798, N2782);
and AND3 (N2799, N2785, N1125, N2743);
nand NAND4 (N2800, N2791, N502, N2214, N1006);
xor XOR2 (N2801, N2793, N755);
or OR2 (N2802, N2792, N123);
and AND3 (N2803, N2801, N1507, N2353);
xor XOR2 (N2804, N2798, N1409);
or OR4 (N2805, N2786, N1182, N659, N87);
nor NOR3 (N2806, N2800, N62, N2078);
nor NOR4 (N2807, N2806, N1905, N1001, N1773);
and AND2 (N2808, N2805, N316);
buf BUF1 (N2809, N2799);
xor XOR2 (N2810, N2795, N763);
nor NOR4 (N2811, N2810, N1608, N2732, N722);
buf BUF1 (N2812, N2807);
nand NAND3 (N2813, N2797, N1862, N610);
not NOT1 (N2814, N2808);
and AND2 (N2815, N2814, N1370);
not NOT1 (N2816, N2811);
xor XOR2 (N2817, N2802, N267);
xor XOR2 (N2818, N2804, N2590);
xor XOR2 (N2819, N2796, N487);
xor XOR2 (N2820, N2809, N2288);
nand NAND2 (N2821, N2812, N2158);
xor XOR2 (N2822, N2820, N1116);
and AND2 (N2823, N2790, N2234);
buf BUF1 (N2824, N2803);
nand NAND4 (N2825, N2823, N2505, N2074, N1303);
buf BUF1 (N2826, N2824);
or OR4 (N2827, N2817, N474, N462, N2774);
not NOT1 (N2828, N2816);
buf BUF1 (N2829, N2827);
and AND4 (N2830, N2813, N937, N40, N1303);
and AND4 (N2831, N2826, N615, N734, N1161);
or OR3 (N2832, N2822, N2168, N1179);
nor NOR2 (N2833, N2830, N2366);
nand NAND3 (N2834, N2821, N2493, N264);
nor NOR2 (N2835, N2825, N2173);
not NOT1 (N2836, N2831);
or OR2 (N2837, N2819, N1808);
or OR4 (N2838, N2836, N1926, N1622, N1657);
nand NAND3 (N2839, N2829, N1660, N885);
nor NOR2 (N2840, N2833, N1108);
and AND3 (N2841, N2815, N970, N1466);
nor NOR2 (N2842, N2837, N763);
and AND4 (N2843, N2835, N2087, N779, N2625);
or OR3 (N2844, N2834, N1817, N2522);
xor XOR2 (N2845, N2840, N1025);
nor NOR2 (N2846, N2838, N2449);
nand NAND2 (N2847, N2842, N2050);
and AND3 (N2848, N2843, N2554, N1766);
nand NAND3 (N2849, N2818, N2661, N2848);
nor NOR2 (N2850, N2384, N2422);
not NOT1 (N2851, N2844);
nand NAND2 (N2852, N2839, N2660);
nor NOR2 (N2853, N2850, N1382);
xor XOR2 (N2854, N2841, N2222);
nor NOR4 (N2855, N2847, N789, N969, N2460);
nor NOR2 (N2856, N2846, N2325);
not NOT1 (N2857, N2845);
nor NOR2 (N2858, N2828, N122);
nor NOR2 (N2859, N2849, N468);
not NOT1 (N2860, N2852);
buf BUF1 (N2861, N2860);
and AND3 (N2862, N2832, N148, N358);
buf BUF1 (N2863, N2857);
or OR3 (N2864, N2859, N1523, N1187);
buf BUF1 (N2865, N2853);
and AND3 (N2866, N2862, N1599, N1634);
not NOT1 (N2867, N2863);
nand NAND2 (N2868, N2861, N187);
buf BUF1 (N2869, N2864);
buf BUF1 (N2870, N2869);
or OR4 (N2871, N2866, N661, N823, N501);
and AND4 (N2872, N2858, N2854, N2825, N2274);
nor NOR4 (N2873, N1851, N408, N1590, N2755);
nor NOR2 (N2874, N2851, N1132);
nand NAND3 (N2875, N2871, N2419, N1737);
or OR2 (N2876, N2855, N2086);
buf BUF1 (N2877, N2872);
not NOT1 (N2878, N2856);
and AND4 (N2879, N2875, N182, N1843, N2328);
or OR2 (N2880, N2870, N154);
or OR2 (N2881, N2880, N1151);
buf BUF1 (N2882, N2874);
buf BUF1 (N2883, N2879);
nor NOR4 (N2884, N2868, N1787, N1344, N58);
not NOT1 (N2885, N2865);
or OR4 (N2886, N2882, N2422, N1957, N580);
nor NOR4 (N2887, N2883, N2629, N793, N161);
not NOT1 (N2888, N2884);
or OR3 (N2889, N2877, N708, N2375);
nand NAND4 (N2890, N2886, N515, N597, N1110);
xor XOR2 (N2891, N2881, N2180);
or OR3 (N2892, N2873, N2555, N1448);
nand NAND2 (N2893, N2888, N2117);
and AND2 (N2894, N2878, N131);
or OR2 (N2895, N2892, N1866);
nor NOR4 (N2896, N2895, N2616, N2007, N1850);
and AND3 (N2897, N2885, N1577, N779);
or OR2 (N2898, N2896, N634);
or OR2 (N2899, N2891, N2640);
nand NAND3 (N2900, N2887, N334, N1497);
not NOT1 (N2901, N2899);
xor XOR2 (N2902, N2893, N383);
xor XOR2 (N2903, N2894, N317);
not NOT1 (N2904, N2902);
nand NAND2 (N2905, N2889, N2450);
nand NAND3 (N2906, N2867, N529, N1493);
or OR4 (N2907, N2905, N631, N1676, N1000);
not NOT1 (N2908, N2898);
buf BUF1 (N2909, N2900);
buf BUF1 (N2910, N2906);
nor NOR4 (N2911, N2901, N1260, N2065, N756);
nand NAND3 (N2912, N2897, N1731, N402);
buf BUF1 (N2913, N2908);
or OR4 (N2914, N2903, N114, N2457, N2108);
or OR2 (N2915, N2907, N2768);
or OR2 (N2916, N2876, N1626);
buf BUF1 (N2917, N2913);
nand NAND3 (N2918, N2915, N2716, N2171);
nor NOR4 (N2919, N2910, N2881, N2329, N763);
not NOT1 (N2920, N2890);
xor XOR2 (N2921, N2912, N2652);
nand NAND3 (N2922, N2920, N59, N989);
not NOT1 (N2923, N2911);
buf BUF1 (N2924, N2917);
and AND4 (N2925, N2909, N958, N2356, N2494);
or OR2 (N2926, N2919, N2243);
and AND4 (N2927, N2918, N1683, N2449, N2724);
buf BUF1 (N2928, N2921);
or OR2 (N2929, N2922, N2355);
not NOT1 (N2930, N2928);
nand NAND2 (N2931, N2914, N196);
nand NAND2 (N2932, N2930, N1097);
or OR4 (N2933, N2916, N447, N1035, N1233);
nand NAND3 (N2934, N2924, N790, N916);
xor XOR2 (N2935, N2904, N2109);
not NOT1 (N2936, N2932);
buf BUF1 (N2937, N2925);
buf BUF1 (N2938, N2923);
nor NOR3 (N2939, N2938, N134, N2611);
nand NAND2 (N2940, N2939, N1911);
or OR4 (N2941, N2936, N815, N2588, N794);
and AND4 (N2942, N2935, N1767, N516, N718);
xor XOR2 (N2943, N2942, N180);
xor XOR2 (N2944, N2937, N2289);
not NOT1 (N2945, N2943);
or OR3 (N2946, N2940, N2747, N1608);
and AND3 (N2947, N2944, N2346, N2057);
or OR3 (N2948, N2947, N747, N1285);
buf BUF1 (N2949, N2946);
not NOT1 (N2950, N2948);
or OR3 (N2951, N2950, N758, N2668);
buf BUF1 (N2952, N2933);
buf BUF1 (N2953, N2927);
xor XOR2 (N2954, N2929, N629);
and AND4 (N2955, N2926, N1389, N1699, N370);
nand NAND2 (N2956, N2934, N2729);
buf BUF1 (N2957, N2945);
xor XOR2 (N2958, N2957, N2645);
not NOT1 (N2959, N2953);
xor XOR2 (N2960, N2931, N2137);
xor XOR2 (N2961, N2955, N1135);
not NOT1 (N2962, N2952);
and AND3 (N2963, N2954, N419, N684);
or OR2 (N2964, N2949, N1837);
buf BUF1 (N2965, N2951);
xor XOR2 (N2966, N2958, N2241);
nand NAND3 (N2967, N2962, N2507, N177);
not NOT1 (N2968, N2965);
or OR4 (N2969, N2963, N2596, N2625, N2437);
and AND3 (N2970, N2956, N2110, N547);
and AND2 (N2971, N2968, N498);
nand NAND2 (N2972, N2967, N423);
buf BUF1 (N2973, N2969);
xor XOR2 (N2974, N2941, N1160);
nand NAND3 (N2975, N2972, N2350, N757);
buf BUF1 (N2976, N2964);
xor XOR2 (N2977, N2975, N2870);
nand NAND4 (N2978, N2977, N1670, N1673, N677);
buf BUF1 (N2979, N2960);
nor NOR4 (N2980, N2979, N1216, N1562, N539);
not NOT1 (N2981, N2966);
buf BUF1 (N2982, N2959);
nor NOR4 (N2983, N2961, N918, N2516, N1878);
nand NAND3 (N2984, N2974, N2457, N1895);
nand NAND4 (N2985, N2973, N2557, N1726, N2555);
and AND3 (N2986, N2978, N2097, N1563);
xor XOR2 (N2987, N2985, N2522);
buf BUF1 (N2988, N2984);
or OR2 (N2989, N2970, N603);
buf BUF1 (N2990, N2988);
or OR2 (N2991, N2980, N2976);
or OR4 (N2992, N874, N194, N1793, N2234);
or OR4 (N2993, N2989, N2302, N37, N1647);
or OR3 (N2994, N2982, N1357, N1902);
nand NAND2 (N2995, N2993, N1772);
nand NAND4 (N2996, N2983, N2516, N2881, N67);
nor NOR4 (N2997, N2992, N1895, N2344, N457);
nor NOR2 (N2998, N2991, N942);
xor XOR2 (N2999, N2986, N1674);
or OR4 (N3000, N2998, N1887, N2974, N1387);
xor XOR2 (N3001, N2990, N1290);
not NOT1 (N3002, N2994);
or OR4 (N3003, N2971, N201, N1184, N2492);
nand NAND4 (N3004, N3003, N1469, N2541, N1340);
nand NAND4 (N3005, N3000, N1660, N2236, N2470);
not NOT1 (N3006, N2981);
nor NOR4 (N3007, N2996, N1950, N345, N263);
not NOT1 (N3008, N3002);
or OR2 (N3009, N3001, N1666);
nand NAND2 (N3010, N3008, N547);
or OR3 (N3011, N3009, N2116, N2681);
buf BUF1 (N3012, N2999);
not NOT1 (N3013, N2997);
buf BUF1 (N3014, N3011);
nor NOR2 (N3015, N3006, N741);
and AND3 (N3016, N2987, N2714, N1998);
nand NAND3 (N3017, N3015, N2821, N575);
and AND2 (N3018, N3005, N456);
and AND3 (N3019, N3010, N1159, N2562);
buf BUF1 (N3020, N3014);
buf BUF1 (N3021, N2995);
not NOT1 (N3022, N3021);
not NOT1 (N3023, N3018);
nand NAND3 (N3024, N3016, N1115, N2118);
not NOT1 (N3025, N3017);
not NOT1 (N3026, N3022);
nor NOR4 (N3027, N3019, N2445, N2723, N678);
nand NAND2 (N3028, N3023, N836);
buf BUF1 (N3029, N3013);
and AND4 (N3030, N3027, N112, N1615, N777);
nor NOR3 (N3031, N3029, N2375, N1066);
not NOT1 (N3032, N3012);
or OR4 (N3033, N3026, N1958, N660, N1458);
not NOT1 (N3034, N3030);
and AND4 (N3035, N3007, N2139, N709, N2051);
or OR2 (N3036, N3025, N1874);
or OR3 (N3037, N3036, N2060, N390);
nand NAND2 (N3038, N3024, N1644);
xor XOR2 (N3039, N3031, N1526);
and AND2 (N3040, N3039, N1481);
not NOT1 (N3041, N3004);
or OR3 (N3042, N3037, N2393, N952);
nor NOR3 (N3043, N3042, N2907, N112);
and AND3 (N3044, N3035, N558, N1791);
not NOT1 (N3045, N3038);
buf BUF1 (N3046, N3044);
buf BUF1 (N3047, N3046);
nand NAND3 (N3048, N3043, N2364, N1141);
nor NOR2 (N3049, N3047, N1265);
buf BUF1 (N3050, N3045);
or OR4 (N3051, N3041, N1900, N381, N2153);
not NOT1 (N3052, N3049);
buf BUF1 (N3053, N3050);
nor NOR3 (N3054, N3040, N1980, N2368);
xor XOR2 (N3055, N3032, N2513);
buf BUF1 (N3056, N3053);
nor NOR2 (N3057, N3028, N341);
and AND3 (N3058, N3048, N2445, N492);
xor XOR2 (N3059, N3033, N2379);
nor NOR2 (N3060, N3055, N1665);
not NOT1 (N3061, N3034);
not NOT1 (N3062, N3051);
nor NOR4 (N3063, N3059, N1679, N1879, N1562);
or OR3 (N3064, N3054, N1066, N1448);
nand NAND3 (N3065, N3060, N854, N174);
not NOT1 (N3066, N3062);
buf BUF1 (N3067, N3057);
nor NOR3 (N3068, N3058, N1667, N1943);
and AND2 (N3069, N3065, N748);
buf BUF1 (N3070, N3063);
buf BUF1 (N3071, N3020);
nor NOR4 (N3072, N3064, N1798, N4, N1832);
xor XOR2 (N3073, N3061, N962);
xor XOR2 (N3074, N3052, N1600);
buf BUF1 (N3075, N3069);
or OR2 (N3076, N3071, N195);
not NOT1 (N3077, N3074);
nor NOR3 (N3078, N3076, N1212, N2388);
xor XOR2 (N3079, N3066, N1085);
not NOT1 (N3080, N3078);
xor XOR2 (N3081, N3068, N1414);
nand NAND3 (N3082, N3079, N1336, N790);
nor NOR3 (N3083, N3073, N2121, N2614);
or OR4 (N3084, N3080, N2472, N593, N2494);
not NOT1 (N3085, N3081);
not NOT1 (N3086, N3085);
buf BUF1 (N3087, N3067);
or OR2 (N3088, N3084, N334);
buf BUF1 (N3089, N3083);
and AND4 (N3090, N3082, N2834, N1082, N2483);
not NOT1 (N3091, N3089);
not NOT1 (N3092, N3075);
not NOT1 (N3093, N3091);
nor NOR2 (N3094, N3072, N2682);
and AND4 (N3095, N3093, N2944, N792, N487);
nand NAND2 (N3096, N3094, N3002);
or OR4 (N3097, N3086, N2014, N3091, N1367);
nor NOR2 (N3098, N3092, N2593);
and AND4 (N3099, N3056, N2455, N1012, N1893);
nor NOR4 (N3100, N3097, N2189, N782, N1198);
xor XOR2 (N3101, N3099, N2041);
xor XOR2 (N3102, N3088, N2692);
nor NOR3 (N3103, N3098, N432, N814);
xor XOR2 (N3104, N3090, N1905);
nor NOR3 (N3105, N3087, N2094, N1376);
not NOT1 (N3106, N3101);
xor XOR2 (N3107, N3105, N357);
buf BUF1 (N3108, N3107);
and AND2 (N3109, N3106, N803);
and AND2 (N3110, N3070, N1393);
or OR2 (N3111, N3102, N226);
xor XOR2 (N3112, N3077, N2644);
nand NAND4 (N3113, N3096, N2842, N1688, N387);
xor XOR2 (N3114, N3113, N2049);
not NOT1 (N3115, N3114);
xor XOR2 (N3116, N3100, N2940);
or OR3 (N3117, N3116, N2420, N1546);
not NOT1 (N3118, N3112);
nor NOR3 (N3119, N3095, N1977, N477);
nand NAND3 (N3120, N3103, N2985, N1835);
buf BUF1 (N3121, N3111);
or OR4 (N3122, N3104, N732, N2622, N568);
nand NAND3 (N3123, N3108, N846, N2813);
and AND2 (N3124, N3115, N406);
xor XOR2 (N3125, N3118, N669);
not NOT1 (N3126, N3122);
buf BUF1 (N3127, N3110);
nor NOR2 (N3128, N3123, N169);
not NOT1 (N3129, N3128);
xor XOR2 (N3130, N3129, N1658);
not NOT1 (N3131, N3119);
nand NAND4 (N3132, N3109, N997, N1379, N1271);
and AND3 (N3133, N3131, N1939, N1060);
or OR2 (N3134, N3127, N538);
nor NOR2 (N3135, N3124, N1276);
nand NAND4 (N3136, N3121, N974, N2586, N2492);
nor NOR4 (N3137, N3117, N1872, N336, N2229);
not NOT1 (N3138, N3130);
and AND2 (N3139, N3135, N2176);
not NOT1 (N3140, N3126);
not NOT1 (N3141, N3139);
or OR2 (N3142, N3120, N1075);
xor XOR2 (N3143, N3142, N35);
nand NAND3 (N3144, N3136, N1979, N832);
buf BUF1 (N3145, N3132);
nor NOR3 (N3146, N3137, N191, N2375);
or OR2 (N3147, N3133, N2074);
nor NOR2 (N3148, N3140, N1061);
xor XOR2 (N3149, N3134, N1698);
not NOT1 (N3150, N3148);
xor XOR2 (N3151, N3150, N2202);
nor NOR2 (N3152, N3144, N670);
xor XOR2 (N3153, N3152, N2330);
nand NAND2 (N3154, N3149, N1666);
and AND2 (N3155, N3151, N467);
not NOT1 (N3156, N3154);
or OR2 (N3157, N3138, N1907);
nor NOR2 (N3158, N3125, N2280);
or OR2 (N3159, N3158, N2347);
and AND4 (N3160, N3145, N2847, N2616, N1579);
nor NOR4 (N3161, N3160, N485, N860, N2011);
nand NAND2 (N3162, N3141, N1568);
nand NAND4 (N3163, N3161, N2457, N368, N1732);
and AND3 (N3164, N3159, N30, N2030);
or OR4 (N3165, N3162, N1443, N336, N2785);
nor NOR3 (N3166, N3147, N1518, N2744);
xor XOR2 (N3167, N3153, N1037);
xor XOR2 (N3168, N3165, N2840);
xor XOR2 (N3169, N3164, N2517);
xor XOR2 (N3170, N3169, N408);
nor NOR4 (N3171, N3168, N2716, N2940, N2016);
and AND4 (N3172, N3157, N683, N2668, N868);
and AND3 (N3173, N3155, N1956, N557);
buf BUF1 (N3174, N3163);
nor NOR2 (N3175, N3170, N483);
xor XOR2 (N3176, N3174, N1474);
xor XOR2 (N3177, N3143, N1025);
or OR4 (N3178, N3175, N1433, N1342, N1658);
nor NOR3 (N3179, N3177, N1442, N2445);
not NOT1 (N3180, N3179);
nor NOR3 (N3181, N3172, N208, N2107);
nand NAND2 (N3182, N3146, N404);
nand NAND2 (N3183, N3166, N2367);
not NOT1 (N3184, N3183);
or OR4 (N3185, N3182, N2282, N3147, N753);
xor XOR2 (N3186, N3180, N736);
and AND3 (N3187, N3176, N2373, N2704);
and AND3 (N3188, N3186, N2839, N322);
buf BUF1 (N3189, N3171);
or OR3 (N3190, N3178, N2483, N2339);
not NOT1 (N3191, N3184);
and AND3 (N3192, N3185, N1854, N2490);
nand NAND2 (N3193, N3192, N1884);
and AND4 (N3194, N3181, N2744, N767, N2245);
not NOT1 (N3195, N3189);
or OR2 (N3196, N3188, N155);
xor XOR2 (N3197, N3195, N2952);
not NOT1 (N3198, N3156);
and AND2 (N3199, N3190, N1836);
nand NAND3 (N3200, N3193, N1524, N1469);
xor XOR2 (N3201, N3167, N14);
and AND4 (N3202, N3198, N1011, N3110, N1566);
not NOT1 (N3203, N3191);
and AND2 (N3204, N3202, N1985);
nor NOR4 (N3205, N3173, N2292, N500, N521);
and AND4 (N3206, N3194, N2051, N2569, N8);
nor NOR2 (N3207, N3206, N1414);
and AND3 (N3208, N3207, N3203, N1731);
not NOT1 (N3209, N1267);
or OR3 (N3210, N3200, N1628, N1214);
buf BUF1 (N3211, N3204);
nand NAND4 (N3212, N3209, N389, N1918, N1899);
and AND4 (N3213, N3208, N2004, N123, N637);
xor XOR2 (N3214, N3213, N2290);
and AND3 (N3215, N3212, N665, N2614);
nor NOR4 (N3216, N3197, N281, N2528, N2711);
nor NOR4 (N3217, N3201, N1383, N207, N2475);
nor NOR4 (N3218, N3215, N280, N2148, N1270);
nor NOR2 (N3219, N3210, N879);
buf BUF1 (N3220, N3214);
or OR3 (N3221, N3220, N1318, N362);
xor XOR2 (N3222, N3205, N2814);
or OR4 (N3223, N3219, N201, N1372, N2242);
nand NAND2 (N3224, N3223, N1908);
buf BUF1 (N3225, N3199);
xor XOR2 (N3226, N3187, N956);
nor NOR3 (N3227, N3221, N2750, N1167);
nand NAND3 (N3228, N3217, N312, N1254);
xor XOR2 (N3229, N3228, N1293);
xor XOR2 (N3230, N3229, N3203);
xor XOR2 (N3231, N3230, N1106);
not NOT1 (N3232, N3211);
not NOT1 (N3233, N3231);
and AND4 (N3234, N3226, N893, N209, N2288);
or OR4 (N3235, N3216, N2446, N1800, N1772);
buf BUF1 (N3236, N3196);
and AND3 (N3237, N3222, N1058, N876);
buf BUF1 (N3238, N3235);
or OR2 (N3239, N3218, N2977);
and AND3 (N3240, N3238, N899, N1889);
nor NOR4 (N3241, N3234, N739, N2228, N1358);
and AND3 (N3242, N3240, N478, N1236);
xor XOR2 (N3243, N3227, N1621);
and AND3 (N3244, N3239, N2573, N2393);
nand NAND2 (N3245, N3232, N1504);
or OR4 (N3246, N3224, N1229, N708, N2289);
buf BUF1 (N3247, N3244);
nand NAND4 (N3248, N3243, N2030, N1988, N1393);
buf BUF1 (N3249, N3247);
nor NOR2 (N3250, N3245, N806);
and AND2 (N3251, N3237, N2370);
xor XOR2 (N3252, N3248, N522);
buf BUF1 (N3253, N3233);
or OR2 (N3254, N3249, N2163);
nor NOR2 (N3255, N3254, N1035);
nor NOR3 (N3256, N3241, N537, N2270);
or OR4 (N3257, N3251, N2912, N2183, N314);
buf BUF1 (N3258, N3246);
nand NAND2 (N3259, N3225, N1081);
or OR3 (N3260, N3259, N3224, N431);
nand NAND4 (N3261, N3255, N2700, N544, N2528);
or OR2 (N3262, N3250, N63);
and AND2 (N3263, N3256, N2520);
not NOT1 (N3264, N3258);
xor XOR2 (N3265, N3262, N762);
not NOT1 (N3266, N3261);
nand NAND4 (N3267, N3266, N1712, N2772, N174);
nand NAND3 (N3268, N3252, N2268, N2913);
and AND2 (N3269, N3268, N122);
nor NOR4 (N3270, N3253, N1619, N879, N3089);
or OR2 (N3271, N3264, N2574);
nand NAND3 (N3272, N3236, N2813, N744);
nand NAND3 (N3273, N3267, N283, N427);
or OR3 (N3274, N3271, N1601, N945);
xor XOR2 (N3275, N3260, N219);
nand NAND3 (N3276, N3273, N1721, N2849);
or OR4 (N3277, N3263, N2987, N1351, N2713);
or OR3 (N3278, N3272, N1642, N2797);
nor NOR2 (N3279, N3277, N2857);
buf BUF1 (N3280, N3269);
xor XOR2 (N3281, N3275, N3209);
nand NAND2 (N3282, N3281, N3257);
buf BUF1 (N3283, N743);
or OR3 (N3284, N3283, N260, N122);
or OR4 (N3285, N3270, N1763, N1195, N488);
not NOT1 (N3286, N3265);
buf BUF1 (N3287, N3285);
or OR3 (N3288, N3284, N2474, N2080);
not NOT1 (N3289, N3287);
or OR3 (N3290, N3278, N799, N2763);
nand NAND4 (N3291, N3274, N20, N1002, N2821);
and AND3 (N3292, N3289, N1328, N1354);
nand NAND3 (N3293, N3280, N3245, N2644);
or OR3 (N3294, N3293, N2381, N2289);
and AND4 (N3295, N3286, N524, N665, N1300);
nor NOR3 (N3296, N3292, N45, N627);
buf BUF1 (N3297, N3279);
buf BUF1 (N3298, N3282);
nand NAND2 (N3299, N3288, N1491);
xor XOR2 (N3300, N3297, N2618);
nor NOR2 (N3301, N3298, N782);
or OR2 (N3302, N3301, N603);
xor XOR2 (N3303, N3302, N3115);
or OR3 (N3304, N3290, N2544, N1328);
and AND4 (N3305, N3242, N2408, N2134, N1778);
nand NAND2 (N3306, N3296, N2187);
or OR2 (N3307, N3305, N2165);
xor XOR2 (N3308, N3304, N1726);
or OR2 (N3309, N3291, N3091);
xor XOR2 (N3310, N3299, N1957);
nand NAND3 (N3311, N3276, N2195, N987);
xor XOR2 (N3312, N3308, N1893);
xor XOR2 (N3313, N3312, N2047);
buf BUF1 (N3314, N3309);
buf BUF1 (N3315, N3313);
buf BUF1 (N3316, N3307);
not NOT1 (N3317, N3316);
nor NOR3 (N3318, N3294, N1948, N2212);
nor NOR2 (N3319, N3310, N1735);
nand NAND3 (N3320, N3295, N1608, N1388);
and AND2 (N3321, N3303, N2121);
xor XOR2 (N3322, N3320, N28);
and AND2 (N3323, N3315, N2736);
nor NOR3 (N3324, N3311, N1028, N2118);
not NOT1 (N3325, N3300);
nand NAND2 (N3326, N3319, N3217);
and AND2 (N3327, N3318, N1626);
not NOT1 (N3328, N3317);
nor NOR4 (N3329, N3321, N452, N1889, N3138);
or OR4 (N3330, N3306, N3122, N2984, N975);
nor NOR3 (N3331, N3324, N2148, N2190);
not NOT1 (N3332, N3314);
nor NOR3 (N3333, N3331, N2306, N2854);
and AND4 (N3334, N3327, N1327, N985, N226);
not NOT1 (N3335, N3329);
nor NOR3 (N3336, N3326, N499, N1920);
nor NOR2 (N3337, N3325, N2398);
nor NOR2 (N3338, N3323, N2487);
xor XOR2 (N3339, N3336, N645);
buf BUF1 (N3340, N3334);
or OR3 (N3341, N3332, N922, N155);
nor NOR2 (N3342, N3335, N359);
nor NOR2 (N3343, N3328, N433);
nand NAND4 (N3344, N3338, N1575, N157, N3144);
buf BUF1 (N3345, N3340);
buf BUF1 (N3346, N3339);
nand NAND4 (N3347, N3346, N2097, N1349, N366);
nand NAND3 (N3348, N3341, N23, N957);
nor NOR2 (N3349, N3345, N2706);
nand NAND4 (N3350, N3343, N1113, N3349, N1665);
or OR4 (N3351, N1328, N32, N2655, N1294);
or OR2 (N3352, N3333, N1718);
nand NAND3 (N3353, N3322, N543, N201);
buf BUF1 (N3354, N3351);
xor XOR2 (N3355, N3348, N879);
xor XOR2 (N3356, N3353, N3029);
nor NOR2 (N3357, N3342, N1961);
nand NAND3 (N3358, N3347, N2876, N3149);
nand NAND3 (N3359, N3352, N3076, N3215);
xor XOR2 (N3360, N3330, N874);
or OR4 (N3361, N3355, N2301, N168, N2271);
nand NAND4 (N3362, N3350, N1972, N3126, N2101);
nand NAND3 (N3363, N3358, N554, N226);
nor NOR3 (N3364, N3337, N2587, N730);
and AND3 (N3365, N3361, N1232, N2394);
or OR3 (N3366, N3364, N2118, N2686);
buf BUF1 (N3367, N3362);
nand NAND4 (N3368, N3366, N2593, N1690, N1467);
or OR3 (N3369, N3360, N2996, N939);
and AND3 (N3370, N3344, N1619, N576);
not NOT1 (N3371, N3368);
not NOT1 (N3372, N3371);
xor XOR2 (N3373, N3357, N2309);
buf BUF1 (N3374, N3369);
buf BUF1 (N3375, N3373);
and AND3 (N3376, N3375, N452, N1461);
or OR3 (N3377, N3365, N1615, N937);
nor NOR3 (N3378, N3372, N2868, N581);
buf BUF1 (N3379, N3377);
or OR3 (N3380, N3359, N576, N913);
nand NAND4 (N3381, N3376, N265, N1760, N421);
and AND4 (N3382, N3374, N3116, N652, N2697);
xor XOR2 (N3383, N3367, N964);
nor NOR2 (N3384, N3382, N2270);
not NOT1 (N3385, N3354);
and AND4 (N3386, N3383, N2290, N2345, N1894);
nand NAND3 (N3387, N3381, N682, N816);
nand NAND3 (N3388, N3356, N64, N1746);
buf BUF1 (N3389, N3386);
nand NAND4 (N3390, N3389, N569, N2551, N3210);
nand NAND3 (N3391, N3380, N577, N3003);
nor NOR4 (N3392, N3379, N1068, N27, N3200);
not NOT1 (N3393, N3392);
xor XOR2 (N3394, N3385, N2857);
or OR4 (N3395, N3394, N2512, N3058, N1915);
nand NAND4 (N3396, N3384, N709, N2399, N1648);
not NOT1 (N3397, N3391);
nand NAND2 (N3398, N3370, N3285);
xor XOR2 (N3399, N3387, N396);
nor NOR2 (N3400, N3378, N3037);
not NOT1 (N3401, N3388);
buf BUF1 (N3402, N3390);
and AND3 (N3403, N3399, N1920, N375);
nand NAND3 (N3404, N3393, N2594, N1395);
nor NOR2 (N3405, N3400, N1132);
not NOT1 (N3406, N3402);
not NOT1 (N3407, N3403);
and AND4 (N3408, N3395, N502, N1778, N1415);
not NOT1 (N3409, N3406);
nand NAND4 (N3410, N3408, N2215, N421, N1971);
buf BUF1 (N3411, N3401);
and AND4 (N3412, N3411, N1606, N24, N1516);
xor XOR2 (N3413, N3363, N2003);
or OR4 (N3414, N3409, N3295, N679, N2762);
and AND3 (N3415, N3407, N2627, N97);
nand NAND2 (N3416, N3405, N3279);
or OR3 (N3417, N3415, N1443, N349);
buf BUF1 (N3418, N3414);
nor NOR2 (N3419, N3397, N247);
buf BUF1 (N3420, N3417);
xor XOR2 (N3421, N3419, N2042);
nor NOR2 (N3422, N3410, N1055);
buf BUF1 (N3423, N3421);
buf BUF1 (N3424, N3422);
xor XOR2 (N3425, N3418, N3409);
buf BUF1 (N3426, N3398);
and AND2 (N3427, N3412, N1574);
xor XOR2 (N3428, N3396, N257);
nor NOR3 (N3429, N3426, N117, N2298);
and AND2 (N3430, N3423, N277);
not NOT1 (N3431, N3427);
nand NAND3 (N3432, N3413, N2131, N1147);
buf BUF1 (N3433, N3432);
nand NAND3 (N3434, N3425, N430, N1666);
or OR2 (N3435, N3424, N1191);
buf BUF1 (N3436, N3429);
nand NAND2 (N3437, N3431, N1734);
nor NOR2 (N3438, N3435, N74);
nand NAND2 (N3439, N3416, N508);
buf BUF1 (N3440, N3438);
not NOT1 (N3441, N3437);
nand NAND3 (N3442, N3436, N1775, N3009);
not NOT1 (N3443, N3434);
not NOT1 (N3444, N3443);
not NOT1 (N3445, N3442);
not NOT1 (N3446, N3404);
xor XOR2 (N3447, N3446, N874);
nand NAND4 (N3448, N3444, N2957, N507, N2295);
and AND4 (N3449, N3439, N3090, N1563, N314);
buf BUF1 (N3450, N3428);
xor XOR2 (N3451, N3433, N2990);
not NOT1 (N3452, N3420);
buf BUF1 (N3453, N3445);
nor NOR2 (N3454, N3447, N736);
nand NAND2 (N3455, N3448, N1424);
or OR3 (N3456, N3453, N838, N2982);
buf BUF1 (N3457, N3456);
xor XOR2 (N3458, N3450, N515);
buf BUF1 (N3459, N3457);
xor XOR2 (N3460, N3440, N3341);
and AND2 (N3461, N3454, N2880);
nand NAND3 (N3462, N3458, N3211, N1086);
nand NAND4 (N3463, N3452, N2408, N674, N3310);
buf BUF1 (N3464, N3461);
nand NAND3 (N3465, N3430, N622, N1504);
nand NAND3 (N3466, N3460, N1673, N2698);
and AND2 (N3467, N3441, N2350);
nand NAND4 (N3468, N3463, N2068, N2082, N1466);
nand NAND3 (N3469, N3467, N826, N1058);
buf BUF1 (N3470, N3469);
nand NAND3 (N3471, N3464, N54, N454);
not NOT1 (N3472, N3471);
or OR4 (N3473, N3472, N35, N3232, N1222);
xor XOR2 (N3474, N3462, N194);
or OR4 (N3475, N3455, N575, N1456, N2552);
nor NOR4 (N3476, N3473, N339, N1667, N1110);
nor NOR3 (N3477, N3468, N2601, N2010);
or OR2 (N3478, N3474, N448);
and AND3 (N3479, N3449, N3371, N455);
nor NOR2 (N3480, N3477, N572);
and AND3 (N3481, N3480, N2199, N3321);
buf BUF1 (N3482, N3479);
and AND4 (N3483, N3475, N159, N2916, N2469);
and AND3 (N3484, N3483, N700, N2459);
and AND4 (N3485, N3470, N1176, N2512, N2681);
not NOT1 (N3486, N3482);
nor NOR4 (N3487, N3451, N1315, N201, N3440);
nor NOR4 (N3488, N3486, N339, N2045, N1405);
nand NAND2 (N3489, N3466, N287);
nand NAND2 (N3490, N3487, N787);
nand NAND4 (N3491, N3489, N3226, N309, N3445);
buf BUF1 (N3492, N3459);
buf BUF1 (N3493, N3491);
nor NOR2 (N3494, N3493, N211);
nand NAND2 (N3495, N3492, N96);
and AND2 (N3496, N3488, N1288);
or OR4 (N3497, N3496, N458, N1148, N1434);
not NOT1 (N3498, N3484);
nand NAND3 (N3499, N3494, N127, N3274);
nand NAND4 (N3500, N3476, N2605, N748, N3192);
not NOT1 (N3501, N3490);
nor NOR2 (N3502, N3499, N1806);
or OR3 (N3503, N3495, N2515, N2691);
nor NOR4 (N3504, N3498, N2286, N9, N457);
nor NOR3 (N3505, N3478, N3473, N3464);
or OR3 (N3506, N3501, N2545, N2876);
nor NOR3 (N3507, N3502, N1854, N393);
and AND3 (N3508, N3481, N1176, N2387);
not NOT1 (N3509, N3497);
nor NOR2 (N3510, N3465, N1901);
nor NOR4 (N3511, N3510, N506, N1198, N1938);
xor XOR2 (N3512, N3509, N764);
buf BUF1 (N3513, N3505);
endmodule