// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24;

output N6415,N6413,N6423,N6392,N6419,N6410,N6420,N6407,N6422,N6424;

or OR2 (N25, N13, N21);
not NOT1 (N26, N22);
or OR3 (N27, N22, N12, N12);
buf BUF1 (N28, N10);
not NOT1 (N29, N3);
nor NOR4 (N30, N11, N10, N17, N12);
nand NAND4 (N31, N13, N7, N3, N27);
not NOT1 (N32, N2);
not NOT1 (N33, N27);
buf BUF1 (N34, N24);
nand NAND2 (N35, N25, N31);
nand NAND2 (N36, N5, N17);
buf BUF1 (N37, N5);
or OR3 (N38, N28, N27, N24);
xor XOR2 (N39, N37, N36);
nand NAND4 (N40, N24, N8, N25, N27);
nand NAND2 (N41, N29, N3);
nor NOR3 (N42, N41, N31, N26);
not NOT1 (N43, N29);
or OR4 (N44, N39, N33, N25, N36);
buf BUF1 (N45, N22);
buf BUF1 (N46, N32);
and AND4 (N47, N34, N28, N2, N33);
not NOT1 (N48, N40);
or OR4 (N49, N46, N15, N5, N35);
or OR2 (N50, N32, N16);
and AND2 (N51, N38, N39);
nand NAND2 (N52, N43, N35);
xor XOR2 (N53, N49, N50);
buf BUF1 (N54, N18);
nand NAND2 (N55, N48, N47);
nor NOR2 (N56, N49, N24);
and AND4 (N57, N52, N28, N6, N56);
or OR3 (N58, N26, N16, N10);
not NOT1 (N59, N57);
and AND4 (N60, N45, N46, N1, N50);
and AND3 (N61, N54, N24, N12);
nand NAND3 (N62, N44, N51, N20);
xor XOR2 (N63, N46, N23);
nand NAND2 (N64, N58, N60);
nor NOR3 (N65, N42, N51, N34);
nand NAND4 (N66, N27, N23, N40, N4);
or OR4 (N67, N53, N22, N19, N11);
nand NAND3 (N68, N66, N58, N7);
nand NAND2 (N69, N61, N34);
and AND2 (N70, N67, N5);
nor NOR2 (N71, N70, N66);
or OR4 (N72, N62, N9, N68, N38);
xor XOR2 (N73, N34, N35);
and AND3 (N74, N55, N65, N63);
nor NOR2 (N75, N16, N26);
xor XOR2 (N76, N68, N72);
xor XOR2 (N77, N49, N26);
not NOT1 (N78, N77);
nor NOR2 (N79, N30, N42);
buf BUF1 (N80, N73);
xor XOR2 (N81, N69, N74);
nor NOR4 (N82, N63, N55, N11, N16);
or OR3 (N83, N71, N6, N33);
or OR2 (N84, N80, N19);
or OR3 (N85, N79, N58, N25);
nand NAND2 (N86, N64, N17);
nand NAND4 (N87, N75, N6, N57, N45);
not NOT1 (N88, N86);
xor XOR2 (N89, N78, N9);
and AND3 (N90, N87, N11, N47);
nor NOR3 (N91, N89, N5, N16);
nor NOR3 (N92, N76, N4, N5);
or OR4 (N93, N92, N47, N31, N67);
nand NAND2 (N94, N59, N7);
and AND4 (N95, N90, N46, N45, N16);
xor XOR2 (N96, N83, N74);
and AND3 (N97, N84, N7, N40);
buf BUF1 (N98, N97);
nand NAND3 (N99, N85, N45, N34);
nand NAND2 (N100, N93, N37);
and AND3 (N101, N81, N23, N34);
xor XOR2 (N102, N100, N32);
and AND3 (N103, N102, N23, N71);
and AND2 (N104, N82, N39);
xor XOR2 (N105, N98, N51);
and AND3 (N106, N94, N65, N46);
buf BUF1 (N107, N95);
or OR4 (N108, N101, N27, N96, N100);
and AND3 (N109, N5, N91, N94);
not NOT1 (N110, N89);
or OR4 (N111, N108, N85, N46, N97);
not NOT1 (N112, N99);
not NOT1 (N113, N111);
buf BUF1 (N114, N112);
buf BUF1 (N115, N104);
nor NOR4 (N116, N106, N63, N16, N24);
not NOT1 (N117, N116);
and AND2 (N118, N105, N73);
and AND3 (N119, N114, N92, N15);
xor XOR2 (N120, N118, N90);
or OR4 (N121, N120, N97, N25, N29);
nand NAND3 (N122, N110, N30, N94);
and AND3 (N123, N103, N100, N120);
buf BUF1 (N124, N115);
not NOT1 (N125, N117);
xor XOR2 (N126, N88, N18);
or OR3 (N127, N113, N91, N65);
and AND4 (N128, N126, N50, N39, N67);
buf BUF1 (N129, N128);
buf BUF1 (N130, N125);
xor XOR2 (N131, N123, N1);
xor XOR2 (N132, N109, N29);
xor XOR2 (N133, N119, N111);
buf BUF1 (N134, N131);
or OR4 (N135, N127, N102, N23, N36);
nor NOR4 (N136, N132, N122, N39, N9);
xor XOR2 (N137, N76, N116);
or OR4 (N138, N130, N55, N101, N5);
nand NAND3 (N139, N121, N59, N123);
nand NAND3 (N140, N124, N97, N55);
nand NAND3 (N141, N134, N53, N44);
or OR2 (N142, N141, N134);
nor NOR3 (N143, N139, N80, N126);
or OR4 (N144, N107, N45, N36, N52);
buf BUF1 (N145, N138);
nor NOR4 (N146, N135, N143, N99, N92);
or OR3 (N147, N95, N24, N11);
not NOT1 (N148, N140);
and AND4 (N149, N147, N117, N19, N68);
or OR2 (N150, N146, N53);
nor NOR4 (N151, N148, N10, N38, N93);
xor XOR2 (N152, N133, N9);
nor NOR4 (N153, N136, N27, N69, N34);
xor XOR2 (N154, N129, N125);
nor NOR4 (N155, N149, N3, N33, N108);
not NOT1 (N156, N150);
buf BUF1 (N157, N144);
or OR4 (N158, N153, N1, N111, N74);
not NOT1 (N159, N152);
nor NOR3 (N160, N157, N119, N76);
xor XOR2 (N161, N154, N26);
or OR2 (N162, N145, N104);
nand NAND2 (N163, N151, N7);
xor XOR2 (N164, N158, N8);
buf BUF1 (N165, N162);
or OR3 (N166, N160, N100, N147);
nand NAND2 (N167, N137, N103);
nand NAND2 (N168, N163, N96);
buf BUF1 (N169, N166);
xor XOR2 (N170, N167, N119);
nand NAND4 (N171, N168, N113, N169, N144);
xor XOR2 (N172, N95, N36);
xor XOR2 (N173, N172, N122);
and AND3 (N174, N170, N20, N63);
not NOT1 (N175, N174);
nand NAND4 (N176, N164, N14, N77, N21);
nor NOR4 (N177, N161, N136, N171, N148);
not NOT1 (N178, N64);
nand NAND3 (N179, N142, N81, N101);
buf BUF1 (N180, N177);
or OR4 (N181, N156, N157, N85, N135);
nor NOR3 (N182, N159, N8, N147);
nor NOR4 (N183, N182, N154, N114, N14);
nor NOR4 (N184, N183, N171, N109, N131);
nand NAND2 (N185, N179, N131);
nor NOR2 (N186, N185, N88);
buf BUF1 (N187, N176);
xor XOR2 (N188, N178, N118);
xor XOR2 (N189, N173, N129);
nor NOR2 (N190, N181, N172);
and AND4 (N191, N186, N130, N90, N39);
buf BUF1 (N192, N184);
xor XOR2 (N193, N188, N17);
nand NAND2 (N194, N193, N176);
buf BUF1 (N195, N187);
not NOT1 (N196, N190);
not NOT1 (N197, N192);
not NOT1 (N198, N191);
or OR4 (N199, N165, N120, N9, N43);
nor NOR2 (N200, N180, N97);
or OR2 (N201, N194, N47);
buf BUF1 (N202, N196);
xor XOR2 (N203, N200, N59);
not NOT1 (N204, N175);
and AND2 (N205, N189, N111);
nand NAND3 (N206, N195, N54, N124);
or OR3 (N207, N199, N112, N127);
nor NOR3 (N208, N206, N169, N45);
not NOT1 (N209, N202);
nor NOR2 (N210, N207, N208);
or OR3 (N211, N177, N20, N33);
or OR2 (N212, N155, N68);
nor NOR2 (N213, N209, N178);
and AND4 (N214, N201, N183, N82, N81);
xor XOR2 (N215, N203, N212);
buf BUF1 (N216, N28);
xor XOR2 (N217, N198, N115);
buf BUF1 (N218, N216);
and AND3 (N219, N204, N180, N158);
or OR4 (N220, N215, N55, N125, N125);
not NOT1 (N221, N219);
nand NAND4 (N222, N220, N149, N209, N14);
nor NOR4 (N223, N218, N122, N192, N147);
nor NOR4 (N224, N223, N150, N93, N161);
nor NOR4 (N225, N222, N160, N178, N41);
not NOT1 (N226, N213);
or OR2 (N227, N205, N15);
not NOT1 (N228, N211);
not NOT1 (N229, N217);
and AND3 (N230, N225, N135, N216);
xor XOR2 (N231, N214, N148);
nand NAND4 (N232, N221, N77, N112, N56);
and AND2 (N233, N224, N100);
buf BUF1 (N234, N197);
and AND2 (N235, N210, N52);
xor XOR2 (N236, N234, N94);
or OR2 (N237, N226, N84);
buf BUF1 (N238, N228);
xor XOR2 (N239, N237, N65);
not NOT1 (N240, N235);
xor XOR2 (N241, N236, N103);
xor XOR2 (N242, N232, N161);
nand NAND3 (N243, N227, N172, N221);
and AND4 (N244, N229, N104, N219, N6);
buf BUF1 (N245, N231);
buf BUF1 (N246, N244);
buf BUF1 (N247, N241);
or OR2 (N248, N247, N161);
and AND3 (N249, N248, N101, N160);
nor NOR2 (N250, N245, N138);
not NOT1 (N251, N238);
and AND3 (N252, N242, N5, N19);
or OR2 (N253, N233, N118);
nand NAND4 (N254, N251, N186, N238, N106);
not NOT1 (N255, N250);
xor XOR2 (N256, N254, N151);
nor NOR3 (N257, N230, N208, N2);
or OR4 (N258, N253, N79, N253, N53);
nand NAND2 (N259, N239, N187);
not NOT1 (N260, N246);
nor NOR4 (N261, N260, N213, N224, N74);
buf BUF1 (N262, N257);
and AND2 (N263, N249, N232);
buf BUF1 (N264, N258);
or OR3 (N265, N243, N7, N184);
or OR4 (N266, N263, N241, N128, N202);
buf BUF1 (N267, N252);
and AND2 (N268, N265, N198);
not NOT1 (N269, N266);
not NOT1 (N270, N268);
xor XOR2 (N271, N255, N141);
not NOT1 (N272, N269);
buf BUF1 (N273, N262);
nor NOR2 (N274, N240, N160);
or OR4 (N275, N267, N266, N214, N160);
nand NAND3 (N276, N273, N65, N209);
not NOT1 (N277, N261);
and AND2 (N278, N264, N8);
xor XOR2 (N279, N274, N5);
buf BUF1 (N280, N279);
and AND3 (N281, N276, N188, N134);
nand NAND2 (N282, N259, N50);
nor NOR4 (N283, N282, N270, N203, N168);
nor NOR4 (N284, N29, N106, N143, N263);
not NOT1 (N285, N275);
xor XOR2 (N286, N280, N275);
nand NAND4 (N287, N285, N116, N34, N286);
and AND2 (N288, N23, N265);
buf BUF1 (N289, N288);
nor NOR3 (N290, N278, N133, N108);
xor XOR2 (N291, N281, N28);
not NOT1 (N292, N284);
nor NOR4 (N293, N291, N77, N234, N36);
nand NAND2 (N294, N283, N167);
xor XOR2 (N295, N256, N164);
or OR4 (N296, N294, N220, N41, N37);
buf BUF1 (N297, N295);
nand NAND3 (N298, N296, N271, N297);
not NOT1 (N299, N113);
buf BUF1 (N300, N270);
nor NOR2 (N301, N299, N10);
buf BUF1 (N302, N287);
xor XOR2 (N303, N301, N238);
not NOT1 (N304, N290);
not NOT1 (N305, N289);
nand NAND2 (N306, N302, N76);
or OR2 (N307, N306, N32);
buf BUF1 (N308, N304);
or OR2 (N309, N292, N71);
or OR3 (N310, N277, N18, N262);
and AND3 (N311, N310, N63, N155);
not NOT1 (N312, N311);
not NOT1 (N313, N305);
not NOT1 (N314, N309);
xor XOR2 (N315, N307, N28);
nand NAND2 (N316, N272, N122);
buf BUF1 (N317, N314);
nor NOR3 (N318, N317, N58, N34);
not NOT1 (N319, N316);
or OR4 (N320, N308, N266, N37, N267);
buf BUF1 (N321, N303);
nor NOR3 (N322, N300, N187, N170);
buf BUF1 (N323, N321);
or OR4 (N324, N318, N189, N169, N256);
nand NAND4 (N325, N324, N79, N173, N23);
nand NAND2 (N326, N323, N191);
nand NAND3 (N327, N293, N277, N113);
nor NOR4 (N328, N322, N33, N124, N161);
buf BUF1 (N329, N298);
buf BUF1 (N330, N328);
or OR4 (N331, N326, N109, N38, N225);
xor XOR2 (N332, N315, N211);
or OR3 (N333, N325, N85, N300);
xor XOR2 (N334, N331, N333);
not NOT1 (N335, N70);
and AND4 (N336, N313, N323, N75, N194);
and AND3 (N337, N327, N27, N94);
not NOT1 (N338, N329);
nand NAND3 (N339, N334, N306, N58);
nor NOR3 (N340, N339, N105, N295);
or OR2 (N341, N319, N104);
buf BUF1 (N342, N312);
not NOT1 (N343, N338);
or OR3 (N344, N342, N144, N30);
not NOT1 (N345, N332);
and AND2 (N346, N341, N114);
or OR4 (N347, N340, N209, N117, N63);
buf BUF1 (N348, N336);
and AND4 (N349, N344, N213, N53, N345);
nand NAND4 (N350, N60, N13, N327, N36);
nor NOR2 (N351, N349, N146);
nand NAND3 (N352, N351, N117, N312);
or OR4 (N353, N347, N292, N134, N60);
not NOT1 (N354, N330);
nand NAND2 (N355, N350, N266);
buf BUF1 (N356, N354);
nor NOR4 (N357, N320, N67, N315, N293);
not NOT1 (N358, N346);
nor NOR4 (N359, N358, N216, N348, N121);
or OR2 (N360, N173, N209);
buf BUF1 (N361, N335);
xor XOR2 (N362, N353, N220);
xor XOR2 (N363, N362, N22);
or OR2 (N364, N360, N124);
nor NOR4 (N365, N356, N40, N201, N162);
not NOT1 (N366, N359);
nand NAND4 (N367, N361, N329, N140, N221);
xor XOR2 (N368, N352, N265);
and AND4 (N369, N364, N24, N49, N228);
buf BUF1 (N370, N365);
nor NOR4 (N371, N369, N151, N334, N125);
or OR4 (N372, N357, N97, N342, N17);
or OR4 (N373, N355, N357, N17, N296);
xor XOR2 (N374, N367, N329);
buf BUF1 (N375, N371);
nand NAND2 (N376, N363, N254);
nor NOR4 (N377, N343, N5, N168, N369);
not NOT1 (N378, N374);
not NOT1 (N379, N375);
not NOT1 (N380, N372);
and AND4 (N381, N373, N172, N315, N32);
nand NAND3 (N382, N378, N48, N22);
or OR4 (N383, N370, N314, N191, N295);
buf BUF1 (N384, N382);
or OR3 (N385, N337, N208, N24);
xor XOR2 (N386, N368, N125);
buf BUF1 (N387, N380);
or OR3 (N388, N387, N53, N341);
nor NOR4 (N389, N366, N123, N3, N67);
not NOT1 (N390, N376);
buf BUF1 (N391, N384);
nand NAND2 (N392, N385, N34);
not NOT1 (N393, N377);
and AND2 (N394, N383, N139);
buf BUF1 (N395, N386);
or OR3 (N396, N379, N296, N35);
nor NOR2 (N397, N388, N241);
or OR2 (N398, N390, N46);
not NOT1 (N399, N391);
or OR3 (N400, N392, N327, N163);
not NOT1 (N401, N399);
buf BUF1 (N402, N398);
nor NOR2 (N403, N401, N361);
buf BUF1 (N404, N403);
xor XOR2 (N405, N397, N265);
nand NAND4 (N406, N394, N2, N329, N107);
and AND3 (N407, N402, N82, N210);
buf BUF1 (N408, N381);
nand NAND4 (N409, N405, N254, N293, N58);
buf BUF1 (N410, N393);
xor XOR2 (N411, N406, N303);
nor NOR2 (N412, N404, N133);
and AND4 (N413, N407, N225, N12, N198);
not NOT1 (N414, N413);
or OR2 (N415, N408, N112);
nor NOR2 (N416, N410, N264);
nand NAND3 (N417, N412, N301, N337);
and AND3 (N418, N409, N375, N295);
nor NOR3 (N419, N418, N148, N7);
or OR2 (N420, N415, N88);
xor XOR2 (N421, N419, N183);
or OR3 (N422, N411, N90, N4);
xor XOR2 (N423, N396, N1);
not NOT1 (N424, N421);
nor NOR2 (N425, N423, N411);
or OR4 (N426, N425, N241, N147, N236);
buf BUF1 (N427, N389);
nor NOR3 (N428, N427, N383, N110);
xor XOR2 (N429, N395, N295);
buf BUF1 (N430, N417);
xor XOR2 (N431, N426, N288);
not NOT1 (N432, N428);
and AND2 (N433, N400, N11);
nor NOR4 (N434, N420, N207, N402, N375);
or OR4 (N435, N422, N113, N54, N134);
xor XOR2 (N436, N432, N264);
buf BUF1 (N437, N431);
xor XOR2 (N438, N416, N366);
nor NOR3 (N439, N435, N426, N327);
buf BUF1 (N440, N430);
nor NOR2 (N441, N436, N193);
and AND3 (N442, N414, N183, N272);
not NOT1 (N443, N442);
nor NOR4 (N444, N441, N433, N360, N400);
not NOT1 (N445, N198);
and AND2 (N446, N438, N407);
buf BUF1 (N447, N446);
nor NOR4 (N448, N443, N2, N355, N113);
nor NOR4 (N449, N448, N395, N23, N150);
and AND3 (N450, N447, N404, N227);
nand NAND2 (N451, N445, N57);
buf BUF1 (N452, N444);
buf BUF1 (N453, N450);
not NOT1 (N454, N439);
not NOT1 (N455, N449);
nor NOR4 (N456, N437, N416, N235, N250);
xor XOR2 (N457, N451, N307);
and AND3 (N458, N455, N268, N299);
nor NOR4 (N459, N424, N126, N285, N358);
nand NAND2 (N460, N458, N98);
nor NOR4 (N461, N459, N199, N61, N422);
or OR2 (N462, N457, N372);
xor XOR2 (N463, N454, N325);
nand NAND4 (N464, N462, N115, N413, N384);
buf BUF1 (N465, N440);
buf BUF1 (N466, N429);
buf BUF1 (N467, N461);
xor XOR2 (N468, N466, N326);
or OR3 (N469, N468, N220, N126);
nor NOR2 (N470, N464, N388);
nor NOR4 (N471, N463, N117, N196, N350);
buf BUF1 (N472, N460);
or OR4 (N473, N452, N21, N238, N2);
nor NOR3 (N474, N456, N248, N169);
nand NAND4 (N475, N471, N65, N107, N188);
and AND4 (N476, N434, N187, N43, N206);
nor NOR2 (N477, N470, N356);
nor NOR2 (N478, N465, N428);
buf BUF1 (N479, N478);
xor XOR2 (N480, N476, N446);
or OR2 (N481, N477, N273);
not NOT1 (N482, N473);
not NOT1 (N483, N475);
or OR2 (N484, N482, N471);
buf BUF1 (N485, N481);
or OR2 (N486, N474, N283);
nand NAND2 (N487, N486, N71);
nor NOR3 (N488, N453, N448, N66);
nand NAND2 (N489, N488, N322);
not NOT1 (N490, N479);
xor XOR2 (N491, N480, N88);
not NOT1 (N492, N469);
nand NAND3 (N493, N489, N162, N46);
nor NOR2 (N494, N492, N38);
and AND2 (N495, N472, N130);
or OR3 (N496, N490, N305, N247);
or OR3 (N497, N493, N473, N436);
nand NAND4 (N498, N495, N158, N360, N77);
nor NOR2 (N499, N491, N404);
xor XOR2 (N500, N487, N277);
nand NAND4 (N501, N484, N24, N149, N298);
or OR3 (N502, N483, N81, N218);
buf BUF1 (N503, N501);
xor XOR2 (N504, N494, N39);
nand NAND2 (N505, N498, N10);
not NOT1 (N506, N505);
buf BUF1 (N507, N497);
or OR2 (N508, N507, N441);
buf BUF1 (N509, N508);
nand NAND4 (N510, N509, N303, N448, N361);
nor NOR2 (N511, N502, N48);
not NOT1 (N512, N506);
or OR4 (N513, N503, N108, N473, N402);
and AND3 (N514, N511, N401, N236);
not NOT1 (N515, N512);
or OR4 (N516, N510, N373, N404, N193);
nor NOR2 (N517, N499, N398);
buf BUF1 (N518, N504);
or OR3 (N519, N485, N128, N10);
nand NAND3 (N520, N467, N191, N470);
xor XOR2 (N521, N520, N357);
not NOT1 (N522, N517);
not NOT1 (N523, N496);
nor NOR3 (N524, N516, N22, N399);
buf BUF1 (N525, N515);
nand NAND4 (N526, N525, N91, N15, N437);
nor NOR2 (N527, N500, N388);
nand NAND3 (N528, N521, N189, N452);
nand NAND3 (N529, N523, N33, N21);
or OR3 (N530, N529, N162, N2);
and AND3 (N531, N513, N154, N144);
not NOT1 (N532, N530);
nand NAND3 (N533, N524, N215, N51);
not NOT1 (N534, N533);
xor XOR2 (N535, N522, N429);
and AND2 (N536, N532, N166);
nor NOR4 (N537, N534, N534, N424, N305);
nand NAND2 (N538, N531, N423);
not NOT1 (N539, N526);
nor NOR3 (N540, N528, N55, N306);
nor NOR2 (N541, N536, N486);
nand NAND4 (N542, N539, N354, N334, N231);
or OR4 (N543, N527, N84, N75, N70);
or OR4 (N544, N542, N128, N359, N438);
xor XOR2 (N545, N544, N142);
not NOT1 (N546, N519);
and AND4 (N547, N541, N490, N192, N545);
nand NAND2 (N548, N392, N348);
nor NOR2 (N549, N538, N155);
or OR4 (N550, N543, N294, N528, N315);
or OR2 (N551, N535, N54);
nor NOR2 (N552, N518, N454);
or OR4 (N553, N547, N208, N86, N526);
nand NAND3 (N554, N550, N494, N445);
not NOT1 (N555, N549);
buf BUF1 (N556, N546);
nand NAND2 (N557, N553, N518);
and AND3 (N558, N537, N55, N109);
nand NAND2 (N559, N558, N488);
buf BUF1 (N560, N555);
or OR4 (N561, N559, N341, N241, N332);
xor XOR2 (N562, N561, N145);
nand NAND2 (N563, N560, N48);
not NOT1 (N564, N556);
or OR4 (N565, N563, N129, N206, N227);
nor NOR4 (N566, N562, N489, N387, N137);
nand NAND4 (N567, N540, N166, N454, N300);
and AND2 (N568, N566, N271);
buf BUF1 (N569, N514);
or OR3 (N570, N567, N82, N113);
not NOT1 (N571, N568);
not NOT1 (N572, N557);
nand NAND2 (N573, N569, N239);
nand NAND3 (N574, N552, N142, N332);
and AND3 (N575, N574, N569, N95);
nor NOR4 (N576, N548, N81, N351, N157);
nand NAND2 (N577, N570, N160);
and AND3 (N578, N573, N373, N31);
nor NOR3 (N579, N554, N103, N196);
or OR4 (N580, N551, N554, N108, N477);
and AND3 (N581, N575, N421, N449);
or OR2 (N582, N579, N394);
and AND2 (N583, N576, N471);
xor XOR2 (N584, N571, N261);
not NOT1 (N585, N578);
xor XOR2 (N586, N565, N261);
or OR4 (N587, N586, N317, N225, N73);
and AND4 (N588, N564, N220, N431, N257);
nand NAND4 (N589, N583, N62, N101, N356);
nand NAND3 (N590, N589, N352, N240);
buf BUF1 (N591, N585);
buf BUF1 (N592, N580);
or OR3 (N593, N581, N450, N310);
buf BUF1 (N594, N577);
xor XOR2 (N595, N590, N553);
nand NAND2 (N596, N587, N265);
and AND2 (N597, N593, N165);
not NOT1 (N598, N591);
and AND3 (N599, N588, N507, N40);
and AND3 (N600, N599, N144, N476);
not NOT1 (N601, N596);
xor XOR2 (N602, N600, N146);
or OR4 (N603, N584, N267, N578, N30);
nor NOR4 (N604, N595, N218, N358, N19);
or OR2 (N605, N594, N282);
buf BUF1 (N606, N604);
xor XOR2 (N607, N572, N561);
or OR2 (N608, N607, N161);
buf BUF1 (N609, N592);
nand NAND3 (N610, N597, N225, N213);
buf BUF1 (N611, N603);
nand NAND3 (N612, N602, N32, N510);
not NOT1 (N613, N612);
not NOT1 (N614, N601);
or OR3 (N615, N609, N123, N324);
not NOT1 (N616, N582);
nand NAND2 (N617, N605, N291);
not NOT1 (N618, N617);
buf BUF1 (N619, N608);
not NOT1 (N620, N610);
and AND2 (N621, N619, N409);
nand NAND4 (N622, N618, N67, N153, N574);
or OR3 (N623, N613, N121, N281);
xor XOR2 (N624, N616, N94);
nand NAND2 (N625, N614, N248);
or OR4 (N626, N611, N159, N282, N425);
nor NOR3 (N627, N620, N379, N573);
not NOT1 (N628, N598);
nand NAND3 (N629, N615, N327, N628);
nor NOR3 (N630, N360, N53, N143);
xor XOR2 (N631, N623, N184);
nand NAND2 (N632, N627, N148);
nand NAND3 (N633, N630, N336, N50);
not NOT1 (N634, N624);
or OR3 (N635, N606, N293, N581);
not NOT1 (N636, N622);
nand NAND3 (N637, N635, N111, N348);
xor XOR2 (N638, N626, N465);
buf BUF1 (N639, N621);
nor NOR3 (N640, N631, N122, N532);
and AND3 (N641, N638, N159, N595);
buf BUF1 (N642, N636);
and AND3 (N643, N640, N577, N369);
and AND4 (N644, N642, N510, N100, N51);
buf BUF1 (N645, N632);
buf BUF1 (N646, N645);
and AND4 (N647, N643, N538, N317, N98);
xor XOR2 (N648, N646, N613);
buf BUF1 (N649, N625);
xor XOR2 (N650, N649, N538);
nand NAND4 (N651, N647, N225, N147, N596);
and AND2 (N652, N637, N551);
buf BUF1 (N653, N629);
not NOT1 (N654, N650);
and AND2 (N655, N651, N641);
or OR4 (N656, N25, N64, N365, N112);
not NOT1 (N657, N654);
nand NAND2 (N658, N644, N359);
or OR3 (N659, N639, N3, N364);
and AND4 (N660, N634, N398, N603, N538);
or OR4 (N661, N659, N182, N16, N500);
buf BUF1 (N662, N648);
or OR3 (N663, N652, N409, N178);
or OR3 (N664, N663, N663, N408);
and AND3 (N665, N657, N408, N97);
not NOT1 (N666, N653);
xor XOR2 (N667, N661, N500);
or OR2 (N668, N665, N6);
nor NOR4 (N669, N667, N134, N324, N438);
not NOT1 (N670, N664);
and AND2 (N671, N633, N99);
and AND2 (N672, N666, N206);
nand NAND3 (N673, N658, N654, N550);
buf BUF1 (N674, N672);
xor XOR2 (N675, N655, N173);
buf BUF1 (N676, N669);
or OR3 (N677, N675, N321, N372);
buf BUF1 (N678, N660);
buf BUF1 (N679, N668);
or OR2 (N680, N676, N488);
not NOT1 (N681, N662);
or OR2 (N682, N674, N600);
and AND3 (N683, N681, N682, N365);
not NOT1 (N684, N595);
nand NAND3 (N685, N679, N627, N138);
xor XOR2 (N686, N683, N217);
xor XOR2 (N687, N677, N153);
nor NOR4 (N688, N687, N276, N585, N508);
nor NOR4 (N689, N670, N284, N197, N309);
or OR3 (N690, N656, N213, N675);
nand NAND2 (N691, N688, N244);
xor XOR2 (N692, N680, N571);
xor XOR2 (N693, N692, N237);
xor XOR2 (N694, N690, N147);
buf BUF1 (N695, N691);
not NOT1 (N696, N694);
or OR2 (N697, N678, N525);
nor NOR3 (N698, N684, N63, N251);
or OR4 (N699, N673, N242, N241, N507);
nand NAND2 (N700, N693, N193);
and AND2 (N701, N689, N527);
buf BUF1 (N702, N699);
xor XOR2 (N703, N671, N433);
and AND4 (N704, N686, N692, N143, N553);
nand NAND2 (N705, N704, N431);
nor NOR4 (N706, N702, N622, N529, N153);
and AND3 (N707, N698, N572, N236);
and AND4 (N708, N685, N558, N117, N414);
xor XOR2 (N709, N705, N539);
not NOT1 (N710, N706);
and AND4 (N711, N696, N84, N222, N364);
not NOT1 (N712, N700);
nand NAND4 (N713, N707, N542, N667, N110);
xor XOR2 (N714, N695, N254);
nand NAND3 (N715, N710, N676, N362);
and AND2 (N716, N703, N207);
buf BUF1 (N717, N711);
xor XOR2 (N718, N712, N315);
not NOT1 (N719, N709);
and AND2 (N720, N697, N445);
nor NOR4 (N721, N716, N301, N84, N124);
and AND4 (N722, N721, N200, N665, N38);
and AND4 (N723, N708, N197, N267, N24);
xor XOR2 (N724, N720, N213);
not NOT1 (N725, N714);
buf BUF1 (N726, N723);
not NOT1 (N727, N719);
or OR3 (N728, N722, N681, N309);
nor NOR3 (N729, N726, N630, N667);
not NOT1 (N730, N715);
and AND4 (N731, N724, N319, N121, N648);
and AND4 (N732, N729, N373, N686, N655);
xor XOR2 (N733, N731, N607);
nand NAND2 (N734, N733, N518);
buf BUF1 (N735, N728);
or OR2 (N736, N734, N372);
nor NOR2 (N737, N730, N632);
buf BUF1 (N738, N732);
buf BUF1 (N739, N713);
or OR2 (N740, N727, N470);
nand NAND2 (N741, N718, N561);
not NOT1 (N742, N737);
nand NAND3 (N743, N701, N477, N204);
and AND3 (N744, N735, N74, N219);
or OR3 (N745, N742, N323, N655);
buf BUF1 (N746, N738);
nor NOR4 (N747, N717, N63, N236, N167);
buf BUF1 (N748, N747);
or OR2 (N749, N746, N718);
not NOT1 (N750, N749);
nand NAND2 (N751, N740, N195);
buf BUF1 (N752, N748);
nand NAND4 (N753, N745, N735, N179, N232);
buf BUF1 (N754, N751);
xor XOR2 (N755, N736, N753);
nor NOR3 (N756, N498, N173, N709);
xor XOR2 (N757, N750, N201);
or OR4 (N758, N755, N131, N19, N98);
and AND4 (N759, N758, N641, N575, N313);
and AND4 (N760, N754, N274, N286, N600);
xor XOR2 (N761, N744, N165);
xor XOR2 (N762, N756, N76);
nand NAND3 (N763, N759, N661, N409);
buf BUF1 (N764, N757);
and AND4 (N765, N761, N387, N305, N343);
nand NAND2 (N766, N760, N406);
and AND4 (N767, N741, N489, N533, N553);
xor XOR2 (N768, N762, N220);
nor NOR2 (N769, N765, N582);
nand NAND2 (N770, N766, N394);
xor XOR2 (N771, N752, N298);
and AND4 (N772, N770, N44, N155, N671);
nor NOR2 (N773, N772, N186);
or OR2 (N774, N773, N751);
not NOT1 (N775, N774);
not NOT1 (N776, N743);
and AND2 (N777, N769, N719);
nand NAND2 (N778, N763, N86);
nand NAND4 (N779, N767, N397, N80, N131);
and AND4 (N780, N775, N12, N591, N700);
buf BUF1 (N781, N779);
or OR4 (N782, N776, N685, N44, N525);
nor NOR2 (N783, N778, N529);
and AND4 (N784, N764, N564, N661, N271);
not NOT1 (N785, N739);
or OR2 (N786, N777, N634);
buf BUF1 (N787, N781);
nand NAND2 (N788, N771, N724);
and AND4 (N789, N786, N371, N148, N745);
nor NOR2 (N790, N782, N336);
or OR4 (N791, N784, N221, N790, N601);
buf BUF1 (N792, N201);
buf BUF1 (N793, N783);
xor XOR2 (N794, N725, N668);
buf BUF1 (N795, N780);
not NOT1 (N796, N794);
nand NAND3 (N797, N787, N640, N686);
nand NAND4 (N798, N792, N324, N154, N609);
buf BUF1 (N799, N768);
not NOT1 (N800, N785);
nor NOR2 (N801, N791, N252);
and AND2 (N802, N799, N296);
nand NAND2 (N803, N788, N772);
and AND3 (N804, N797, N112, N37);
not NOT1 (N805, N789);
and AND4 (N806, N803, N151, N62, N317);
not NOT1 (N807, N795);
nor NOR3 (N808, N801, N192, N535);
nor NOR4 (N809, N808, N543, N805, N721);
buf BUF1 (N810, N486);
and AND3 (N811, N800, N371, N353);
nand NAND4 (N812, N793, N600, N197, N611);
nand NAND2 (N813, N809, N218);
buf BUF1 (N814, N811);
nor NOR4 (N815, N796, N208, N73, N591);
nand NAND3 (N816, N798, N282, N503);
nand NAND2 (N817, N804, N475);
not NOT1 (N818, N812);
nand NAND4 (N819, N814, N797, N310, N55);
buf BUF1 (N820, N819);
xor XOR2 (N821, N807, N511);
or OR3 (N822, N820, N374, N116);
buf BUF1 (N823, N822);
or OR3 (N824, N821, N560, N576);
nand NAND2 (N825, N824, N31);
nor NOR2 (N826, N802, N700);
or OR2 (N827, N817, N57);
buf BUF1 (N828, N816);
or OR4 (N829, N828, N504, N291, N676);
xor XOR2 (N830, N810, N39);
xor XOR2 (N831, N826, N321);
buf BUF1 (N832, N815);
nor NOR2 (N833, N829, N483);
and AND4 (N834, N806, N520, N639, N690);
nand NAND4 (N835, N832, N140, N270, N206);
buf BUF1 (N836, N835);
nand NAND2 (N837, N827, N469);
or OR3 (N838, N825, N524, N171);
nand NAND4 (N839, N834, N550, N816, N293);
buf BUF1 (N840, N836);
nor NOR4 (N841, N839, N746, N717, N183);
xor XOR2 (N842, N838, N674);
nand NAND4 (N843, N813, N472, N601, N374);
nand NAND2 (N844, N843, N146);
or OR3 (N845, N833, N438, N107);
nand NAND4 (N846, N831, N361, N553, N651);
xor XOR2 (N847, N840, N729);
nor NOR2 (N848, N837, N540);
nor NOR2 (N849, N847, N458);
xor XOR2 (N850, N849, N119);
or OR3 (N851, N844, N425, N537);
or OR2 (N852, N818, N674);
nand NAND3 (N853, N851, N147, N205);
or OR4 (N854, N823, N16, N849, N62);
nor NOR2 (N855, N853, N164);
xor XOR2 (N856, N854, N745);
nor NOR4 (N857, N845, N412, N113, N626);
buf BUF1 (N858, N842);
and AND2 (N859, N848, N589);
xor XOR2 (N860, N850, N399);
nor NOR3 (N861, N856, N33, N292);
or OR3 (N862, N855, N325, N681);
xor XOR2 (N863, N857, N107);
nor NOR2 (N864, N830, N495);
or OR2 (N865, N841, N837);
buf BUF1 (N866, N865);
and AND4 (N867, N846, N833, N266, N251);
xor XOR2 (N868, N852, N843);
buf BUF1 (N869, N858);
xor XOR2 (N870, N866, N508);
nor NOR3 (N871, N863, N659, N564);
nor NOR2 (N872, N871, N765);
and AND2 (N873, N867, N802);
and AND3 (N874, N859, N334, N677);
or OR4 (N875, N864, N611, N595, N690);
buf BUF1 (N876, N874);
nor NOR4 (N877, N870, N5, N323, N836);
not NOT1 (N878, N869);
nor NOR3 (N879, N875, N427, N281);
and AND3 (N880, N879, N403, N363);
not NOT1 (N881, N877);
or OR4 (N882, N868, N115, N297, N813);
buf BUF1 (N883, N878);
or OR3 (N884, N883, N645, N835);
and AND2 (N885, N880, N244);
nor NOR2 (N886, N873, N301);
xor XOR2 (N887, N872, N870);
not NOT1 (N888, N860);
nor NOR3 (N889, N881, N331, N479);
nand NAND3 (N890, N876, N519, N296);
nand NAND2 (N891, N861, N458);
nand NAND4 (N892, N889, N629, N670, N209);
nand NAND2 (N893, N890, N733);
xor XOR2 (N894, N887, N378);
nand NAND2 (N895, N885, N326);
nor NOR2 (N896, N892, N828);
not NOT1 (N897, N891);
and AND3 (N898, N862, N392, N599);
buf BUF1 (N899, N894);
and AND4 (N900, N888, N665, N337, N312);
xor XOR2 (N901, N900, N533);
nor NOR2 (N902, N886, N693);
nor NOR2 (N903, N893, N189);
and AND3 (N904, N884, N558, N790);
and AND3 (N905, N899, N390, N530);
nor NOR2 (N906, N903, N416);
xor XOR2 (N907, N905, N221);
nand NAND3 (N908, N882, N830, N533);
nor NOR3 (N909, N901, N636, N189);
nand NAND2 (N910, N895, N594);
nand NAND4 (N911, N904, N881, N651, N249);
nor NOR2 (N912, N897, N390);
buf BUF1 (N913, N896);
or OR4 (N914, N910, N111, N200, N651);
not NOT1 (N915, N906);
nor NOR4 (N916, N907, N562, N539, N366);
or OR2 (N917, N913, N142);
nor NOR3 (N918, N911, N475, N895);
and AND2 (N919, N917, N447);
nor NOR3 (N920, N914, N594, N905);
buf BUF1 (N921, N919);
xor XOR2 (N922, N918, N471);
buf BUF1 (N923, N909);
and AND4 (N924, N902, N509, N682, N247);
not NOT1 (N925, N920);
and AND2 (N926, N915, N576);
buf BUF1 (N927, N924);
not NOT1 (N928, N912);
nor NOR2 (N929, N925, N502);
xor XOR2 (N930, N916, N648);
nand NAND3 (N931, N908, N434, N360);
xor XOR2 (N932, N922, N243);
buf BUF1 (N933, N929);
nand NAND4 (N934, N928, N794, N66, N301);
not NOT1 (N935, N931);
or OR4 (N936, N898, N331, N381, N587);
nand NAND3 (N937, N935, N563, N237);
nor NOR2 (N938, N937, N188);
or OR2 (N939, N926, N558);
and AND4 (N940, N930, N64, N826, N444);
nand NAND4 (N941, N921, N920, N516, N358);
nor NOR3 (N942, N939, N400, N546);
xor XOR2 (N943, N941, N932);
and AND2 (N944, N783, N860);
nand NAND4 (N945, N938, N245, N414, N164);
and AND3 (N946, N923, N61, N599);
nor NOR2 (N947, N933, N108);
xor XOR2 (N948, N942, N331);
nor NOR2 (N949, N934, N26);
buf BUF1 (N950, N936);
xor XOR2 (N951, N943, N260);
buf BUF1 (N952, N948);
nand NAND4 (N953, N947, N746, N11, N547);
xor XOR2 (N954, N951, N801);
buf BUF1 (N955, N952);
buf BUF1 (N956, N954);
and AND2 (N957, N950, N691);
nand NAND3 (N958, N927, N850, N501);
or OR4 (N959, N946, N203, N362, N544);
buf BUF1 (N960, N949);
nand NAND3 (N961, N957, N750, N671);
not NOT1 (N962, N956);
buf BUF1 (N963, N955);
buf BUF1 (N964, N962);
buf BUF1 (N965, N960);
buf BUF1 (N966, N953);
buf BUF1 (N967, N940);
nor NOR2 (N968, N964, N887);
xor XOR2 (N969, N966, N709);
nand NAND2 (N970, N945, N656);
or OR3 (N971, N965, N455, N497);
not NOT1 (N972, N970);
nand NAND4 (N973, N963, N691, N514, N897);
nand NAND4 (N974, N961, N701, N461, N816);
not NOT1 (N975, N973);
nand NAND4 (N976, N974, N208, N679, N302);
or OR3 (N977, N976, N653, N339);
or OR2 (N978, N977, N34);
nor NOR3 (N979, N978, N99, N364);
xor XOR2 (N980, N979, N812);
or OR4 (N981, N971, N876, N30, N732);
xor XOR2 (N982, N968, N192);
not NOT1 (N983, N958);
nand NAND2 (N984, N982, N977);
or OR2 (N985, N980, N761);
xor XOR2 (N986, N969, N91);
nand NAND2 (N987, N975, N406);
nand NAND3 (N988, N967, N892, N274);
or OR4 (N989, N944, N955, N182, N185);
and AND4 (N990, N981, N854, N321, N530);
nor NOR3 (N991, N988, N100, N918);
nand NAND2 (N992, N986, N978);
nand NAND2 (N993, N972, N584);
xor XOR2 (N994, N983, N31);
not NOT1 (N995, N959);
buf BUF1 (N996, N995);
and AND2 (N997, N989, N646);
and AND4 (N998, N992, N376, N320, N261);
nor NOR2 (N999, N990, N538);
nor NOR2 (N1000, N994, N936);
nor NOR2 (N1001, N996, N460);
nand NAND4 (N1002, N1000, N585, N390, N590);
nor NOR2 (N1003, N998, N327);
or OR4 (N1004, N1001, N516, N195, N674);
nor NOR2 (N1005, N1003, N914);
not NOT1 (N1006, N985);
and AND4 (N1007, N1004, N981, N460, N210);
and AND4 (N1008, N993, N634, N66, N59);
buf BUF1 (N1009, N1005);
and AND3 (N1010, N1002, N594, N619);
xor XOR2 (N1011, N999, N518);
nand NAND4 (N1012, N1006, N759, N412, N556);
xor XOR2 (N1013, N987, N121);
xor XOR2 (N1014, N991, N12);
buf BUF1 (N1015, N1009);
or OR4 (N1016, N1015, N155, N612, N325);
xor XOR2 (N1017, N984, N216);
buf BUF1 (N1018, N997);
xor XOR2 (N1019, N1014, N1007);
xor XOR2 (N1020, N78, N731);
nor NOR3 (N1021, N1017, N326, N215);
nand NAND2 (N1022, N1021, N980);
xor XOR2 (N1023, N1012, N89);
or OR2 (N1024, N1019, N146);
buf BUF1 (N1025, N1008);
or OR4 (N1026, N1016, N347, N162, N401);
and AND2 (N1027, N1025, N679);
buf BUF1 (N1028, N1011);
not NOT1 (N1029, N1020);
and AND4 (N1030, N1024, N387, N149, N511);
and AND2 (N1031, N1018, N343);
or OR2 (N1032, N1028, N1027);
not NOT1 (N1033, N283);
xor XOR2 (N1034, N1022, N909);
xor XOR2 (N1035, N1034, N165);
nand NAND4 (N1036, N1035, N152, N724, N391);
and AND4 (N1037, N1029, N323, N424, N704);
nand NAND2 (N1038, N1031, N630);
and AND3 (N1039, N1013, N79, N12);
or OR2 (N1040, N1037, N679);
nand NAND2 (N1041, N1010, N605);
xor XOR2 (N1042, N1040, N932);
or OR2 (N1043, N1039, N470);
xor XOR2 (N1044, N1038, N518);
xor XOR2 (N1045, N1043, N305);
nand NAND3 (N1046, N1044, N126, N9);
buf BUF1 (N1047, N1030);
buf BUF1 (N1048, N1033);
or OR2 (N1049, N1045, N463);
nor NOR2 (N1050, N1047, N569);
buf BUF1 (N1051, N1046);
buf BUF1 (N1052, N1051);
nor NOR3 (N1053, N1036, N169, N252);
or OR2 (N1054, N1023, N351);
and AND4 (N1055, N1049, N116, N618, N501);
and AND4 (N1056, N1050, N113, N277, N459);
or OR2 (N1057, N1026, N99);
buf BUF1 (N1058, N1053);
xor XOR2 (N1059, N1052, N427);
nor NOR2 (N1060, N1058, N999);
buf BUF1 (N1061, N1056);
not NOT1 (N1062, N1060);
and AND3 (N1063, N1054, N968, N159);
not NOT1 (N1064, N1041);
not NOT1 (N1065, N1061);
nor NOR2 (N1066, N1057, N848);
xor XOR2 (N1067, N1063, N310);
nand NAND4 (N1068, N1065, N162, N1044, N259);
and AND3 (N1069, N1066, N663, N691);
buf BUF1 (N1070, N1059);
and AND3 (N1071, N1068, N774, N268);
nor NOR3 (N1072, N1070, N282, N429);
xor XOR2 (N1073, N1062, N924);
buf BUF1 (N1074, N1073);
not NOT1 (N1075, N1071);
nand NAND4 (N1076, N1069, N112, N505, N651);
nor NOR3 (N1077, N1067, N433, N666);
nor NOR4 (N1078, N1048, N429, N882, N516);
nand NAND3 (N1079, N1078, N264, N931);
xor XOR2 (N1080, N1042, N67);
not NOT1 (N1081, N1079);
not NOT1 (N1082, N1055);
not NOT1 (N1083, N1076);
xor XOR2 (N1084, N1082, N222);
nor NOR4 (N1085, N1032, N371, N1, N420);
and AND4 (N1086, N1083, N93, N468, N867);
nor NOR2 (N1087, N1077, N399);
nor NOR4 (N1088, N1064, N291, N910, N966);
nand NAND4 (N1089, N1084, N896, N306, N125);
or OR3 (N1090, N1086, N596, N453);
and AND3 (N1091, N1072, N980, N324);
or OR3 (N1092, N1089, N639, N353);
not NOT1 (N1093, N1074);
nand NAND2 (N1094, N1092, N30);
or OR4 (N1095, N1075, N764, N87, N503);
buf BUF1 (N1096, N1090);
nor NOR4 (N1097, N1087, N299, N488, N727);
xor XOR2 (N1098, N1088, N754);
buf BUF1 (N1099, N1095);
nor NOR2 (N1100, N1085, N265);
buf BUF1 (N1101, N1097);
xor XOR2 (N1102, N1101, N222);
xor XOR2 (N1103, N1096, N598);
nor NOR3 (N1104, N1093, N1049, N180);
buf BUF1 (N1105, N1091);
buf BUF1 (N1106, N1080);
not NOT1 (N1107, N1094);
not NOT1 (N1108, N1104);
not NOT1 (N1109, N1108);
and AND2 (N1110, N1105, N119);
and AND3 (N1111, N1102, N371, N435);
not NOT1 (N1112, N1109);
or OR4 (N1113, N1112, N174, N401, N491);
buf BUF1 (N1114, N1107);
and AND3 (N1115, N1113, N23, N454);
or OR2 (N1116, N1114, N811);
xor XOR2 (N1117, N1098, N473);
or OR4 (N1118, N1100, N840, N499, N418);
nand NAND3 (N1119, N1118, N786, N2);
nor NOR3 (N1120, N1110, N586, N125);
or OR2 (N1121, N1117, N467);
nand NAND4 (N1122, N1081, N276, N121, N571);
nand NAND3 (N1123, N1121, N666, N186);
nand NAND2 (N1124, N1116, N776);
not NOT1 (N1125, N1115);
and AND4 (N1126, N1122, N483, N588, N336);
not NOT1 (N1127, N1124);
nor NOR2 (N1128, N1127, N171);
xor XOR2 (N1129, N1123, N921);
buf BUF1 (N1130, N1099);
buf BUF1 (N1131, N1119);
or OR4 (N1132, N1130, N630, N198, N144);
or OR3 (N1133, N1126, N756, N904);
xor XOR2 (N1134, N1106, N232);
and AND2 (N1135, N1131, N743);
or OR4 (N1136, N1120, N770, N807, N701);
nand NAND3 (N1137, N1136, N450, N793);
buf BUF1 (N1138, N1137);
nor NOR2 (N1139, N1111, N350);
nand NAND3 (N1140, N1134, N473, N280);
buf BUF1 (N1141, N1135);
or OR3 (N1142, N1103, N496, N405);
xor XOR2 (N1143, N1140, N549);
xor XOR2 (N1144, N1139, N341);
or OR4 (N1145, N1142, N429, N476, N1016);
nand NAND2 (N1146, N1132, N850);
and AND4 (N1147, N1125, N393, N676, N577);
and AND3 (N1148, N1141, N437, N694);
xor XOR2 (N1149, N1145, N741);
and AND2 (N1150, N1149, N386);
buf BUF1 (N1151, N1144);
nand NAND2 (N1152, N1150, N790);
or OR4 (N1153, N1128, N969, N197, N841);
nor NOR2 (N1154, N1143, N375);
nor NOR3 (N1155, N1153, N203, N44);
buf BUF1 (N1156, N1148);
and AND3 (N1157, N1156, N787, N609);
and AND4 (N1158, N1146, N238, N648, N356);
buf BUF1 (N1159, N1133);
xor XOR2 (N1160, N1152, N778);
or OR2 (N1161, N1147, N605);
buf BUF1 (N1162, N1159);
nand NAND3 (N1163, N1154, N849, N839);
buf BUF1 (N1164, N1158);
nand NAND3 (N1165, N1161, N293, N283);
buf BUF1 (N1166, N1151);
xor XOR2 (N1167, N1129, N873);
xor XOR2 (N1168, N1162, N1087);
or OR2 (N1169, N1167, N766);
buf BUF1 (N1170, N1166);
xor XOR2 (N1171, N1164, N781);
xor XOR2 (N1172, N1138, N1027);
or OR2 (N1173, N1163, N526);
and AND2 (N1174, N1165, N875);
buf BUF1 (N1175, N1155);
nor NOR3 (N1176, N1170, N918, N703);
not NOT1 (N1177, N1175);
or OR3 (N1178, N1174, N324, N832);
not NOT1 (N1179, N1176);
or OR3 (N1180, N1160, N151, N878);
nor NOR3 (N1181, N1168, N169, N453);
nand NAND2 (N1182, N1169, N985);
or OR4 (N1183, N1157, N311, N965, N505);
not NOT1 (N1184, N1179);
xor XOR2 (N1185, N1172, N868);
or OR4 (N1186, N1180, N790, N97, N490);
and AND3 (N1187, N1186, N370, N622);
not NOT1 (N1188, N1183);
not NOT1 (N1189, N1188);
not NOT1 (N1190, N1178);
and AND2 (N1191, N1189, N407);
and AND3 (N1192, N1173, N477, N1106);
not NOT1 (N1193, N1184);
xor XOR2 (N1194, N1193, N85);
nor NOR2 (N1195, N1181, N484);
buf BUF1 (N1196, N1182);
buf BUF1 (N1197, N1185);
buf BUF1 (N1198, N1196);
xor XOR2 (N1199, N1198, N332);
nor NOR3 (N1200, N1191, N1087, N769);
or OR4 (N1201, N1200, N621, N632, N1139);
nand NAND2 (N1202, N1195, N158);
and AND4 (N1203, N1171, N367, N1061, N763);
nor NOR4 (N1204, N1190, N339, N716, N7);
not NOT1 (N1205, N1177);
nand NAND2 (N1206, N1194, N94);
nor NOR2 (N1207, N1187, N865);
buf BUF1 (N1208, N1207);
nor NOR3 (N1209, N1208, N756, N930);
xor XOR2 (N1210, N1201, N70);
buf BUF1 (N1211, N1209);
and AND4 (N1212, N1206, N298, N641, N570);
nand NAND2 (N1213, N1202, N910);
or OR4 (N1214, N1199, N408, N36, N699);
nor NOR2 (N1215, N1212, N797);
buf BUF1 (N1216, N1205);
xor XOR2 (N1217, N1192, N790);
not NOT1 (N1218, N1217);
and AND2 (N1219, N1210, N617);
or OR2 (N1220, N1211, N30);
or OR2 (N1221, N1215, N442);
xor XOR2 (N1222, N1203, N849);
and AND4 (N1223, N1216, N355, N235, N738);
xor XOR2 (N1224, N1219, N897);
nor NOR3 (N1225, N1224, N976, N377);
and AND3 (N1226, N1218, N534, N1057);
nor NOR4 (N1227, N1222, N723, N99, N649);
or OR2 (N1228, N1221, N850);
not NOT1 (N1229, N1197);
nor NOR2 (N1230, N1220, N1212);
nor NOR3 (N1231, N1225, N988, N829);
nand NAND4 (N1232, N1204, N102, N915, N240);
buf BUF1 (N1233, N1214);
nor NOR2 (N1234, N1231, N512);
and AND4 (N1235, N1232, N502, N860, N9);
nor NOR3 (N1236, N1227, N788, N1185);
not NOT1 (N1237, N1228);
xor XOR2 (N1238, N1229, N620);
buf BUF1 (N1239, N1213);
nor NOR2 (N1240, N1223, N306);
and AND4 (N1241, N1239, N48, N1034, N315);
xor XOR2 (N1242, N1236, N1122);
xor XOR2 (N1243, N1237, N1103);
and AND4 (N1244, N1240, N630, N645, N113);
nand NAND4 (N1245, N1241, N520, N1183, N56);
not NOT1 (N1246, N1235);
xor XOR2 (N1247, N1238, N608);
buf BUF1 (N1248, N1246);
and AND4 (N1249, N1248, N1042, N60, N913);
and AND3 (N1250, N1249, N394, N533);
or OR3 (N1251, N1233, N669, N885);
nor NOR3 (N1252, N1244, N829, N364);
or OR4 (N1253, N1251, N1099, N2, N129);
or OR4 (N1254, N1253, N487, N602, N329);
nor NOR4 (N1255, N1242, N1054, N13, N1180);
not NOT1 (N1256, N1243);
and AND3 (N1257, N1226, N1003, N891);
or OR2 (N1258, N1257, N973);
nor NOR4 (N1259, N1234, N309, N407, N304);
nand NAND4 (N1260, N1252, N269, N1137, N212);
not NOT1 (N1261, N1230);
not NOT1 (N1262, N1245);
not NOT1 (N1263, N1255);
and AND3 (N1264, N1260, N340, N935);
and AND4 (N1265, N1262, N788, N961, N892);
nor NOR4 (N1266, N1259, N383, N414, N873);
nand NAND2 (N1267, N1264, N298);
not NOT1 (N1268, N1258);
buf BUF1 (N1269, N1263);
or OR4 (N1270, N1268, N534, N825, N979);
nor NOR4 (N1271, N1270, N615, N119, N962);
nor NOR4 (N1272, N1271, N938, N748, N327);
or OR4 (N1273, N1254, N1258, N392, N317);
not NOT1 (N1274, N1265);
xor XOR2 (N1275, N1274, N646);
buf BUF1 (N1276, N1250);
nor NOR4 (N1277, N1276, N658, N239, N581);
nor NOR2 (N1278, N1275, N1243);
buf BUF1 (N1279, N1273);
nor NOR2 (N1280, N1278, N734);
nand NAND2 (N1281, N1279, N1189);
and AND4 (N1282, N1272, N434, N666, N757);
not NOT1 (N1283, N1256);
or OR2 (N1284, N1269, N359);
not NOT1 (N1285, N1281);
not NOT1 (N1286, N1261);
xor XOR2 (N1287, N1286, N722);
buf BUF1 (N1288, N1266);
nor NOR2 (N1289, N1247, N844);
xor XOR2 (N1290, N1287, N373);
nand NAND3 (N1291, N1283, N990, N145);
nor NOR4 (N1292, N1291, N114, N917, N1122);
or OR2 (N1293, N1284, N1045);
not NOT1 (N1294, N1288);
and AND2 (N1295, N1289, N706);
buf BUF1 (N1296, N1295);
and AND3 (N1297, N1285, N740, N795);
xor XOR2 (N1298, N1296, N137);
buf BUF1 (N1299, N1267);
or OR3 (N1300, N1277, N888, N275);
nand NAND4 (N1301, N1299, N416, N471, N1203);
nor NOR2 (N1302, N1297, N593);
nor NOR4 (N1303, N1302, N1067, N932, N939);
buf BUF1 (N1304, N1292);
xor XOR2 (N1305, N1303, N1042);
xor XOR2 (N1306, N1305, N1039);
not NOT1 (N1307, N1293);
xor XOR2 (N1308, N1282, N436);
xor XOR2 (N1309, N1307, N1230);
or OR4 (N1310, N1309, N1014, N61, N815);
and AND2 (N1311, N1308, N477);
and AND4 (N1312, N1310, N496, N1092, N410);
not NOT1 (N1313, N1301);
and AND4 (N1314, N1306, N75, N1127, N678);
and AND3 (N1315, N1311, N304, N110);
not NOT1 (N1316, N1304);
xor XOR2 (N1317, N1280, N1284);
not NOT1 (N1318, N1315);
or OR4 (N1319, N1316, N280, N969, N1098);
and AND3 (N1320, N1298, N771, N1029);
nand NAND3 (N1321, N1314, N571, N1021);
buf BUF1 (N1322, N1313);
nor NOR2 (N1323, N1319, N111);
not NOT1 (N1324, N1290);
not NOT1 (N1325, N1321);
nand NAND3 (N1326, N1318, N456, N1280);
not NOT1 (N1327, N1294);
xor XOR2 (N1328, N1325, N922);
buf BUF1 (N1329, N1327);
buf BUF1 (N1330, N1328);
buf BUF1 (N1331, N1323);
not NOT1 (N1332, N1326);
nand NAND4 (N1333, N1332, N353, N394, N125);
and AND3 (N1334, N1333, N937, N521);
and AND4 (N1335, N1300, N1036, N980, N533);
or OR2 (N1336, N1335, N322);
buf BUF1 (N1337, N1312);
xor XOR2 (N1338, N1322, N985);
nor NOR3 (N1339, N1329, N444, N590);
not NOT1 (N1340, N1320);
or OR4 (N1341, N1330, N420, N1298, N214);
nor NOR2 (N1342, N1339, N105);
and AND2 (N1343, N1337, N560);
and AND4 (N1344, N1340, N921, N401, N70);
not NOT1 (N1345, N1344);
nor NOR4 (N1346, N1324, N1263, N1190, N596);
buf BUF1 (N1347, N1334);
or OR2 (N1348, N1341, N641);
nor NOR2 (N1349, N1331, N902);
buf BUF1 (N1350, N1349);
not NOT1 (N1351, N1348);
not NOT1 (N1352, N1346);
or OR4 (N1353, N1350, N1178, N1084, N685);
buf BUF1 (N1354, N1352);
and AND2 (N1355, N1343, N27);
not NOT1 (N1356, N1353);
nand NAND2 (N1357, N1347, N872);
or OR4 (N1358, N1355, N238, N433, N398);
buf BUF1 (N1359, N1317);
xor XOR2 (N1360, N1345, N973);
or OR2 (N1361, N1357, N870);
xor XOR2 (N1362, N1354, N1187);
nor NOR3 (N1363, N1338, N47, N1229);
or OR4 (N1364, N1363, N969, N804, N1257);
and AND2 (N1365, N1336, N303);
xor XOR2 (N1366, N1342, N389);
nor NOR3 (N1367, N1360, N697, N954);
nor NOR3 (N1368, N1365, N167, N1192);
and AND3 (N1369, N1364, N1119, N1155);
or OR2 (N1370, N1366, N1294);
and AND3 (N1371, N1369, N255, N990);
nand NAND2 (N1372, N1371, N235);
and AND3 (N1373, N1361, N1341, N193);
xor XOR2 (N1374, N1356, N632);
nor NOR2 (N1375, N1359, N1243);
nor NOR4 (N1376, N1372, N884, N276, N742);
and AND2 (N1377, N1358, N365);
nor NOR2 (N1378, N1376, N642);
buf BUF1 (N1379, N1375);
and AND4 (N1380, N1367, N1231, N985, N92);
buf BUF1 (N1381, N1373);
not NOT1 (N1382, N1362);
nand NAND3 (N1383, N1377, N1260, N218);
or OR3 (N1384, N1380, N66, N1372);
not NOT1 (N1385, N1368);
and AND4 (N1386, N1351, N662, N450, N43);
or OR2 (N1387, N1379, N1171);
xor XOR2 (N1388, N1386, N845);
buf BUF1 (N1389, N1370);
not NOT1 (N1390, N1389);
buf BUF1 (N1391, N1381);
nor NOR4 (N1392, N1378, N50, N517, N222);
buf BUF1 (N1393, N1390);
xor XOR2 (N1394, N1383, N153);
nand NAND4 (N1395, N1391, N523, N319, N486);
or OR3 (N1396, N1388, N610, N491);
nor NOR3 (N1397, N1374, N925, N1283);
or OR4 (N1398, N1384, N1332, N245, N745);
nand NAND3 (N1399, N1394, N116, N1133);
or OR2 (N1400, N1395, N175);
nand NAND2 (N1401, N1385, N471);
buf BUF1 (N1402, N1387);
and AND3 (N1403, N1398, N633, N3);
not NOT1 (N1404, N1392);
nor NOR4 (N1405, N1403, N1132, N1245, N1187);
or OR2 (N1406, N1393, N793);
not NOT1 (N1407, N1399);
or OR3 (N1408, N1396, N893, N1058);
xor XOR2 (N1409, N1402, N89);
buf BUF1 (N1410, N1400);
nor NOR3 (N1411, N1407, N866, N1362);
xor XOR2 (N1412, N1406, N114);
nor NOR2 (N1413, N1405, N1248);
not NOT1 (N1414, N1397);
and AND2 (N1415, N1410, N338);
nand NAND3 (N1416, N1404, N665, N601);
xor XOR2 (N1417, N1409, N606);
and AND2 (N1418, N1382, N140);
xor XOR2 (N1419, N1417, N1144);
and AND3 (N1420, N1412, N891, N998);
nor NOR4 (N1421, N1420, N1213, N980, N1000);
or OR2 (N1422, N1421, N1279);
and AND4 (N1423, N1411, N76, N963, N951);
nor NOR3 (N1424, N1413, N1140, N209);
buf BUF1 (N1425, N1418);
xor XOR2 (N1426, N1408, N218);
and AND4 (N1427, N1415, N455, N1339, N865);
xor XOR2 (N1428, N1427, N611);
nand NAND4 (N1429, N1423, N97, N590, N1199);
nand NAND2 (N1430, N1426, N557);
or OR3 (N1431, N1414, N418, N1173);
not NOT1 (N1432, N1428);
not NOT1 (N1433, N1429);
and AND3 (N1434, N1419, N13, N728);
and AND4 (N1435, N1431, N1371, N627, N1100);
nor NOR3 (N1436, N1432, N519, N291);
and AND3 (N1437, N1436, N897, N1022);
and AND3 (N1438, N1437, N580, N82);
buf BUF1 (N1439, N1425);
nand NAND2 (N1440, N1439, N111);
nor NOR3 (N1441, N1430, N182, N172);
xor XOR2 (N1442, N1434, N716);
nand NAND3 (N1443, N1433, N1112, N593);
or OR3 (N1444, N1401, N1062, N381);
buf BUF1 (N1445, N1438);
nand NAND2 (N1446, N1424, N836);
nor NOR4 (N1447, N1446, N866, N1348, N1222);
or OR2 (N1448, N1441, N1238);
and AND3 (N1449, N1445, N652, N945);
not NOT1 (N1450, N1435);
not NOT1 (N1451, N1442);
xor XOR2 (N1452, N1448, N960);
nor NOR3 (N1453, N1449, N336, N1335);
xor XOR2 (N1454, N1444, N1028);
not NOT1 (N1455, N1453);
nor NOR4 (N1456, N1416, N74, N769, N751);
not NOT1 (N1457, N1454);
and AND2 (N1458, N1452, N244);
and AND2 (N1459, N1443, N1193);
or OR2 (N1460, N1440, N911);
nand NAND3 (N1461, N1456, N412, N107);
buf BUF1 (N1462, N1461);
xor XOR2 (N1463, N1459, N820);
or OR3 (N1464, N1422, N1229, N157);
nor NOR3 (N1465, N1457, N1221, N24);
xor XOR2 (N1466, N1460, N184);
xor XOR2 (N1467, N1466, N746);
nand NAND3 (N1468, N1455, N1079, N42);
or OR4 (N1469, N1450, N170, N687, N1267);
and AND3 (N1470, N1469, N416, N1281);
or OR3 (N1471, N1458, N21, N456);
not NOT1 (N1472, N1462);
not NOT1 (N1473, N1465);
buf BUF1 (N1474, N1473);
nand NAND3 (N1475, N1447, N660, N214);
or OR4 (N1476, N1474, N736, N1175, N610);
nand NAND3 (N1477, N1476, N418, N480);
and AND4 (N1478, N1463, N1352, N501, N579);
or OR4 (N1479, N1478, N1468, N964, N989);
or OR4 (N1480, N356, N745, N801, N479);
not NOT1 (N1481, N1470);
or OR4 (N1482, N1479, N991, N1442, N720);
or OR4 (N1483, N1471, N877, N1381, N334);
not NOT1 (N1484, N1451);
or OR2 (N1485, N1482, N832);
nand NAND2 (N1486, N1484, N262);
nor NOR3 (N1487, N1481, N215, N1418);
nor NOR3 (N1488, N1480, N1036, N1282);
nor NOR2 (N1489, N1483, N696);
nand NAND3 (N1490, N1486, N428, N184);
or OR4 (N1491, N1467, N84, N771, N1139);
or OR4 (N1492, N1490, N908, N900, N240);
or OR4 (N1493, N1492, N772, N496, N1023);
buf BUF1 (N1494, N1488);
and AND2 (N1495, N1475, N732);
and AND4 (N1496, N1472, N1204, N268, N1154);
xor XOR2 (N1497, N1489, N690);
nand NAND3 (N1498, N1477, N1447, N4);
and AND4 (N1499, N1493, N565, N105, N343);
buf BUF1 (N1500, N1487);
and AND4 (N1501, N1498, N275, N197, N1358);
nor NOR4 (N1502, N1495, N55, N1256, N945);
and AND3 (N1503, N1496, N1063, N1258);
or OR4 (N1504, N1464, N1015, N1280, N300);
not NOT1 (N1505, N1494);
nand NAND3 (N1506, N1503, N621, N1058);
buf BUF1 (N1507, N1491);
not NOT1 (N1508, N1500);
and AND2 (N1509, N1505, N839);
and AND4 (N1510, N1502, N1057, N1290, N769);
nor NOR2 (N1511, N1501, N502);
not NOT1 (N1512, N1510);
nand NAND4 (N1513, N1507, N869, N967, N779);
xor XOR2 (N1514, N1485, N1474);
or OR3 (N1515, N1508, N878, N1112);
and AND3 (N1516, N1504, N1030, N1205);
not NOT1 (N1517, N1512);
nor NOR2 (N1518, N1497, N806);
nand NAND3 (N1519, N1518, N82, N955);
or OR4 (N1520, N1509, N569, N163, N923);
and AND3 (N1521, N1514, N702, N1462);
nor NOR2 (N1522, N1516, N344);
or OR4 (N1523, N1519, N42, N254, N657);
not NOT1 (N1524, N1499);
buf BUF1 (N1525, N1523);
nand NAND3 (N1526, N1517, N107, N443);
nand NAND3 (N1527, N1506, N93, N401);
not NOT1 (N1528, N1522);
nor NOR2 (N1529, N1513, N524);
and AND4 (N1530, N1529, N577, N1144, N817);
and AND4 (N1531, N1524, N198, N349, N880);
buf BUF1 (N1532, N1528);
not NOT1 (N1533, N1526);
or OR4 (N1534, N1515, N1201, N1399, N276);
or OR4 (N1535, N1511, N793, N742, N1303);
xor XOR2 (N1536, N1521, N1256);
xor XOR2 (N1537, N1520, N519);
buf BUF1 (N1538, N1530);
nor NOR4 (N1539, N1533, N292, N316, N1287);
buf BUF1 (N1540, N1525);
nor NOR4 (N1541, N1540, N1404, N1274, N1247);
not NOT1 (N1542, N1534);
not NOT1 (N1543, N1538);
buf BUF1 (N1544, N1532);
xor XOR2 (N1545, N1543, N1063);
and AND2 (N1546, N1531, N738);
or OR4 (N1547, N1542, N1150, N595, N129);
nand NAND4 (N1548, N1539, N1320, N305, N595);
not NOT1 (N1549, N1548);
or OR2 (N1550, N1527, N211);
nor NOR2 (N1551, N1541, N702);
nor NOR2 (N1552, N1536, N644);
or OR4 (N1553, N1549, N365, N1132, N916);
nor NOR2 (N1554, N1546, N846);
and AND4 (N1555, N1537, N603, N660, N388);
not NOT1 (N1556, N1553);
not NOT1 (N1557, N1547);
xor XOR2 (N1558, N1552, N644);
not NOT1 (N1559, N1556);
buf BUF1 (N1560, N1557);
or OR2 (N1561, N1544, N1494);
nand NAND3 (N1562, N1550, N1428, N965);
and AND3 (N1563, N1535, N807, N203);
nor NOR4 (N1564, N1559, N1468, N587, N1533);
xor XOR2 (N1565, N1561, N1283);
buf BUF1 (N1566, N1562);
nor NOR3 (N1567, N1560, N404, N1474);
or OR3 (N1568, N1558, N628, N534);
buf BUF1 (N1569, N1545);
buf BUF1 (N1570, N1554);
buf BUF1 (N1571, N1551);
or OR3 (N1572, N1555, N1097, N886);
buf BUF1 (N1573, N1566);
nand NAND3 (N1574, N1570, N1177, N106);
nand NAND4 (N1575, N1565, N1235, N669, N825);
buf BUF1 (N1576, N1571);
not NOT1 (N1577, N1569);
nand NAND4 (N1578, N1572, N1549, N1533, N1345);
not NOT1 (N1579, N1575);
buf BUF1 (N1580, N1568);
not NOT1 (N1581, N1578);
nand NAND2 (N1582, N1573, N947);
or OR2 (N1583, N1567, N646);
nand NAND2 (N1584, N1580, N388);
xor XOR2 (N1585, N1583, N18);
and AND3 (N1586, N1581, N477, N539);
xor XOR2 (N1587, N1563, N585);
and AND3 (N1588, N1577, N156, N491);
and AND3 (N1589, N1584, N125, N629);
and AND3 (N1590, N1585, N1197, N415);
nand NAND4 (N1591, N1589, N180, N137, N208);
and AND3 (N1592, N1576, N737, N645);
and AND2 (N1593, N1586, N52);
xor XOR2 (N1594, N1564, N1276);
nor NOR2 (N1595, N1590, N90);
not NOT1 (N1596, N1593);
xor XOR2 (N1597, N1596, N216);
not NOT1 (N1598, N1582);
buf BUF1 (N1599, N1574);
xor XOR2 (N1600, N1594, N1330);
or OR4 (N1601, N1597, N978, N1518, N699);
nor NOR4 (N1602, N1600, N1098, N1361, N1217);
not NOT1 (N1603, N1595);
and AND3 (N1604, N1588, N1482, N911);
nand NAND3 (N1605, N1587, N768, N623);
and AND2 (N1606, N1602, N441);
nand NAND2 (N1607, N1591, N584);
nor NOR4 (N1608, N1604, N647, N748, N686);
and AND3 (N1609, N1601, N1320, N1483);
and AND3 (N1610, N1592, N202, N548);
not NOT1 (N1611, N1598);
or OR2 (N1612, N1603, N633);
or OR4 (N1613, N1612, N241, N1247, N758);
nor NOR3 (N1614, N1613, N1440, N1332);
xor XOR2 (N1615, N1605, N967);
buf BUF1 (N1616, N1579);
or OR2 (N1617, N1610, N99);
nor NOR4 (N1618, N1614, N284, N1611, N663);
or OR3 (N1619, N115, N1098, N125);
xor XOR2 (N1620, N1609, N533);
nand NAND2 (N1621, N1608, N531);
and AND2 (N1622, N1606, N1299);
nand NAND4 (N1623, N1617, N1418, N1465, N990);
xor XOR2 (N1624, N1616, N726);
xor XOR2 (N1625, N1615, N963);
or OR2 (N1626, N1599, N205);
or OR2 (N1627, N1626, N1062);
or OR4 (N1628, N1618, N421, N1287, N847);
xor XOR2 (N1629, N1624, N1147);
nor NOR3 (N1630, N1629, N1574, N1460);
nand NAND2 (N1631, N1607, N1066);
buf BUF1 (N1632, N1621);
nand NAND2 (N1633, N1628, N575);
nand NAND3 (N1634, N1631, N210, N610);
nand NAND4 (N1635, N1625, N455, N1335, N1326);
nand NAND4 (N1636, N1622, N1406, N375, N942);
xor XOR2 (N1637, N1619, N1000);
nand NAND3 (N1638, N1637, N918, N1536);
xor XOR2 (N1639, N1632, N425);
nor NOR2 (N1640, N1634, N368);
xor XOR2 (N1641, N1636, N1257);
not NOT1 (N1642, N1620);
xor XOR2 (N1643, N1635, N152);
nand NAND3 (N1644, N1630, N580, N613);
buf BUF1 (N1645, N1639);
and AND2 (N1646, N1643, N1243);
nand NAND2 (N1647, N1644, N113);
and AND4 (N1648, N1640, N615, N920, N280);
nand NAND2 (N1649, N1642, N1029);
and AND2 (N1650, N1638, N986);
buf BUF1 (N1651, N1623);
nand NAND2 (N1652, N1633, N1550);
nor NOR4 (N1653, N1648, N991, N1195, N815);
or OR2 (N1654, N1653, N1063);
xor XOR2 (N1655, N1646, N1235);
or OR3 (N1656, N1641, N1336, N151);
or OR2 (N1657, N1647, N749);
not NOT1 (N1658, N1649);
nor NOR2 (N1659, N1656, N1327);
or OR4 (N1660, N1658, N884, N1589, N1168);
or OR4 (N1661, N1645, N736, N848, N350);
xor XOR2 (N1662, N1655, N196);
or OR3 (N1663, N1627, N150, N155);
xor XOR2 (N1664, N1661, N1414);
and AND4 (N1665, N1660, N1207, N1051, N409);
buf BUF1 (N1666, N1659);
xor XOR2 (N1667, N1657, N349);
buf BUF1 (N1668, N1665);
buf BUF1 (N1669, N1668);
nor NOR4 (N1670, N1650, N870, N40, N259);
not NOT1 (N1671, N1666);
xor XOR2 (N1672, N1671, N1019);
nand NAND4 (N1673, N1669, N1400, N22, N1613);
xor XOR2 (N1674, N1673, N1218);
and AND2 (N1675, N1651, N591);
or OR3 (N1676, N1672, N1482, N1019);
not NOT1 (N1677, N1662);
buf BUF1 (N1678, N1676);
nor NOR2 (N1679, N1663, N834);
not NOT1 (N1680, N1675);
and AND4 (N1681, N1667, N1206, N1459, N1584);
and AND2 (N1682, N1654, N1508);
not NOT1 (N1683, N1674);
not NOT1 (N1684, N1679);
xor XOR2 (N1685, N1652, N1098);
xor XOR2 (N1686, N1677, N744);
xor XOR2 (N1687, N1686, N638);
xor XOR2 (N1688, N1664, N12);
or OR2 (N1689, N1682, N355);
and AND4 (N1690, N1688, N1670, N1637, N757);
nor NOR2 (N1691, N846, N1158);
or OR2 (N1692, N1681, N1294);
xor XOR2 (N1693, N1691, N610);
nor NOR3 (N1694, N1687, N539, N1119);
not NOT1 (N1695, N1678);
xor XOR2 (N1696, N1693, N1439);
and AND4 (N1697, N1696, N49, N721, N1094);
nor NOR3 (N1698, N1697, N1649, N1639);
xor XOR2 (N1699, N1680, N353);
nand NAND3 (N1700, N1695, N1076, N949);
buf BUF1 (N1701, N1699);
not NOT1 (N1702, N1689);
buf BUF1 (N1703, N1702);
and AND2 (N1704, N1698, N201);
nand NAND2 (N1705, N1683, N310);
nor NOR2 (N1706, N1692, N89);
buf BUF1 (N1707, N1704);
xor XOR2 (N1708, N1700, N884);
nand NAND4 (N1709, N1684, N1247, N1495, N528);
nand NAND2 (N1710, N1705, N692);
or OR4 (N1711, N1694, N269, N823, N1347);
nand NAND2 (N1712, N1706, N193);
or OR4 (N1713, N1703, N1075, N379, N1403);
xor XOR2 (N1714, N1713, N963);
xor XOR2 (N1715, N1701, N735);
and AND2 (N1716, N1715, N439);
buf BUF1 (N1717, N1714);
buf BUF1 (N1718, N1716);
not NOT1 (N1719, N1718);
buf BUF1 (N1720, N1708);
or OR3 (N1721, N1685, N19, N1549);
nand NAND4 (N1722, N1721, N202, N68, N705);
and AND4 (N1723, N1719, N59, N942, N691);
nor NOR4 (N1724, N1711, N373, N1317, N996);
xor XOR2 (N1725, N1724, N537);
nor NOR2 (N1726, N1707, N43);
nand NAND4 (N1727, N1710, N817, N1713, N268);
xor XOR2 (N1728, N1720, N1725);
or OR4 (N1729, N1328, N107, N544, N1673);
nand NAND3 (N1730, N1729, N639, N530);
xor XOR2 (N1731, N1709, N1015);
not NOT1 (N1732, N1726);
buf BUF1 (N1733, N1732);
and AND2 (N1734, N1723, N1013);
and AND2 (N1735, N1730, N1712);
buf BUF1 (N1736, N240);
nand NAND3 (N1737, N1722, N940, N539);
xor XOR2 (N1738, N1731, N141);
nand NAND2 (N1739, N1737, N206);
or OR4 (N1740, N1690, N1593, N1467, N1449);
not NOT1 (N1741, N1728);
xor XOR2 (N1742, N1738, N133);
nand NAND2 (N1743, N1734, N1684);
nand NAND4 (N1744, N1717, N757, N1581, N995);
or OR2 (N1745, N1744, N489);
nor NOR2 (N1746, N1735, N382);
nand NAND2 (N1747, N1743, N167);
buf BUF1 (N1748, N1742);
buf BUF1 (N1749, N1740);
nand NAND2 (N1750, N1736, N133);
nor NOR3 (N1751, N1745, N1589, N417);
nor NOR3 (N1752, N1746, N873, N187);
xor XOR2 (N1753, N1727, N889);
nand NAND2 (N1754, N1733, N321);
and AND3 (N1755, N1741, N395, N1684);
or OR2 (N1756, N1749, N78);
nor NOR3 (N1757, N1747, N1559, N1358);
nor NOR3 (N1758, N1739, N14, N343);
and AND2 (N1759, N1755, N194);
xor XOR2 (N1760, N1757, N1272);
nor NOR2 (N1761, N1756, N163);
xor XOR2 (N1762, N1760, N53);
nand NAND4 (N1763, N1762, N1583, N1021, N876);
buf BUF1 (N1764, N1750);
nand NAND4 (N1765, N1748, N1285, N1232, N2);
not NOT1 (N1766, N1764);
and AND3 (N1767, N1753, N1383, N439);
nand NAND3 (N1768, N1752, N323, N1662);
and AND4 (N1769, N1766, N269, N125, N1577);
nand NAND2 (N1770, N1759, N907);
xor XOR2 (N1771, N1769, N1353);
nor NOR2 (N1772, N1765, N57);
nand NAND2 (N1773, N1768, N1310);
buf BUF1 (N1774, N1758);
xor XOR2 (N1775, N1767, N1202);
or OR2 (N1776, N1751, N1375);
not NOT1 (N1777, N1770);
and AND4 (N1778, N1777, N1221, N1713, N161);
not NOT1 (N1779, N1763);
not NOT1 (N1780, N1774);
nor NOR2 (N1781, N1779, N569);
xor XOR2 (N1782, N1761, N1157);
and AND3 (N1783, N1773, N540, N1459);
and AND3 (N1784, N1772, N240, N403);
and AND3 (N1785, N1778, N1285, N1378);
buf BUF1 (N1786, N1775);
nor NOR4 (N1787, N1780, N768, N1121, N1608);
or OR4 (N1788, N1781, N946, N776, N735);
nor NOR4 (N1789, N1788, N25, N425, N809);
nor NOR2 (N1790, N1782, N893);
xor XOR2 (N1791, N1789, N1392);
and AND2 (N1792, N1784, N1557);
nor NOR2 (N1793, N1787, N1378);
nor NOR2 (N1794, N1793, N1789);
nand NAND2 (N1795, N1794, N577);
and AND3 (N1796, N1785, N835, N357);
not NOT1 (N1797, N1786);
xor XOR2 (N1798, N1797, N827);
buf BUF1 (N1799, N1754);
not NOT1 (N1800, N1783);
nand NAND2 (N1801, N1792, N1677);
buf BUF1 (N1802, N1796);
nand NAND4 (N1803, N1798, N319, N987, N1778);
nand NAND4 (N1804, N1776, N423, N140, N1226);
nor NOR4 (N1805, N1791, N984, N487, N778);
or OR3 (N1806, N1800, N1462, N517);
buf BUF1 (N1807, N1804);
or OR4 (N1808, N1803, N622, N994, N1210);
buf BUF1 (N1809, N1790);
not NOT1 (N1810, N1801);
not NOT1 (N1811, N1802);
and AND2 (N1812, N1771, N1581);
and AND2 (N1813, N1811, N1682);
or OR4 (N1814, N1812, N1755, N35, N641);
or OR2 (N1815, N1805, N1512);
nor NOR3 (N1816, N1806, N1029, N1536);
and AND3 (N1817, N1813, N1732, N647);
or OR2 (N1818, N1809, N1141);
not NOT1 (N1819, N1799);
xor XOR2 (N1820, N1808, N941);
not NOT1 (N1821, N1820);
or OR2 (N1822, N1818, N1200);
not NOT1 (N1823, N1814);
not NOT1 (N1824, N1815);
not NOT1 (N1825, N1821);
not NOT1 (N1826, N1816);
and AND3 (N1827, N1817, N313, N1785);
not NOT1 (N1828, N1819);
and AND3 (N1829, N1795, N538, N1550);
buf BUF1 (N1830, N1829);
not NOT1 (N1831, N1807);
not NOT1 (N1832, N1822);
xor XOR2 (N1833, N1823, N1292);
nor NOR3 (N1834, N1831, N787, N1560);
or OR3 (N1835, N1827, N1626, N532);
xor XOR2 (N1836, N1826, N1184);
not NOT1 (N1837, N1810);
buf BUF1 (N1838, N1828);
not NOT1 (N1839, N1824);
not NOT1 (N1840, N1834);
xor XOR2 (N1841, N1833, N1207);
and AND3 (N1842, N1830, N797, N1010);
and AND4 (N1843, N1836, N930, N972, N690);
nand NAND2 (N1844, N1840, N133);
not NOT1 (N1845, N1837);
not NOT1 (N1846, N1832);
nand NAND4 (N1847, N1838, N1402, N826, N10);
and AND3 (N1848, N1835, N168, N246);
nand NAND3 (N1849, N1844, N1435, N1311);
nand NAND4 (N1850, N1845, N1170, N653, N1094);
or OR4 (N1851, N1847, N71, N1081, N618);
xor XOR2 (N1852, N1841, N1500);
and AND3 (N1853, N1842, N1418, N1019);
nor NOR4 (N1854, N1851, N459, N671, N1274);
and AND3 (N1855, N1843, N1065, N1764);
xor XOR2 (N1856, N1853, N1170);
xor XOR2 (N1857, N1850, N462);
xor XOR2 (N1858, N1857, N1495);
xor XOR2 (N1859, N1854, N522);
nor NOR3 (N1860, N1855, N1793, N1505);
nand NAND3 (N1861, N1860, N1253, N1512);
nor NOR3 (N1862, N1848, N1634, N1825);
nand NAND4 (N1863, N363, N1702, N400, N1176);
nor NOR3 (N1864, N1858, N676, N696);
not NOT1 (N1865, N1846);
or OR3 (N1866, N1862, N1818, N702);
nor NOR3 (N1867, N1859, N734, N1008);
buf BUF1 (N1868, N1866);
nor NOR2 (N1869, N1849, N901);
or OR4 (N1870, N1868, N1763, N560, N839);
nor NOR4 (N1871, N1864, N1802, N755, N207);
and AND2 (N1872, N1852, N1777);
xor XOR2 (N1873, N1869, N215);
or OR4 (N1874, N1870, N923, N1102, N1398);
and AND2 (N1875, N1863, N245);
buf BUF1 (N1876, N1872);
not NOT1 (N1877, N1876);
xor XOR2 (N1878, N1861, N445);
xor XOR2 (N1879, N1878, N495);
nand NAND4 (N1880, N1875, N104, N1162, N1699);
nand NAND3 (N1881, N1865, N771, N798);
buf BUF1 (N1882, N1839);
nor NOR4 (N1883, N1856, N1365, N612, N1514);
nor NOR4 (N1884, N1874, N561, N18, N421);
nor NOR4 (N1885, N1882, N967, N1852, N937);
buf BUF1 (N1886, N1871);
nand NAND2 (N1887, N1884, N784);
buf BUF1 (N1888, N1867);
or OR2 (N1889, N1880, N1780);
nor NOR3 (N1890, N1889, N1069, N199);
buf BUF1 (N1891, N1877);
nor NOR2 (N1892, N1891, N204);
nor NOR3 (N1893, N1879, N502, N1425);
nand NAND2 (N1894, N1892, N1635);
and AND4 (N1895, N1885, N204, N1687, N174);
not NOT1 (N1896, N1883);
nand NAND2 (N1897, N1894, N1147);
and AND3 (N1898, N1888, N433, N1717);
nor NOR2 (N1899, N1896, N412);
nor NOR4 (N1900, N1897, N1399, N463, N173);
xor XOR2 (N1901, N1890, N984);
nand NAND2 (N1902, N1898, N553);
or OR3 (N1903, N1901, N27, N202);
or OR2 (N1904, N1886, N1499);
or OR3 (N1905, N1893, N957, N1518);
or OR2 (N1906, N1895, N97);
not NOT1 (N1907, N1905);
or OR3 (N1908, N1907, N336, N1507);
or OR2 (N1909, N1904, N1697);
xor XOR2 (N1910, N1902, N480);
buf BUF1 (N1911, N1906);
or OR4 (N1912, N1908, N1766, N1142, N1805);
and AND3 (N1913, N1887, N862, N31);
not NOT1 (N1914, N1900);
not NOT1 (N1915, N1899);
nand NAND2 (N1916, N1873, N1032);
nor NOR3 (N1917, N1881, N276, N64);
xor XOR2 (N1918, N1914, N234);
or OR4 (N1919, N1909, N427, N1431, N1694);
or OR4 (N1920, N1915, N1404, N540, N746);
not NOT1 (N1921, N1910);
nor NOR3 (N1922, N1920, N900, N165);
or OR2 (N1923, N1917, N895);
not NOT1 (N1924, N1918);
nand NAND4 (N1925, N1903, N703, N1545, N918);
xor XOR2 (N1926, N1922, N814);
nor NOR2 (N1927, N1926, N974);
and AND4 (N1928, N1911, N1830, N1026, N86);
not NOT1 (N1929, N1916);
not NOT1 (N1930, N1928);
buf BUF1 (N1931, N1924);
and AND4 (N1932, N1931, N815, N1561, N1196);
xor XOR2 (N1933, N1929, N331);
nor NOR4 (N1934, N1933, N1617, N1153, N764);
and AND4 (N1935, N1925, N1592, N655, N198);
nor NOR3 (N1936, N1930, N928, N1183);
not NOT1 (N1937, N1912);
and AND4 (N1938, N1932, N187, N1750, N341);
or OR4 (N1939, N1921, N133, N1720, N1384);
and AND2 (N1940, N1913, N681);
nor NOR3 (N1941, N1923, N1204, N1750);
xor XOR2 (N1942, N1940, N303);
xor XOR2 (N1943, N1938, N730);
not NOT1 (N1944, N1919);
nor NOR4 (N1945, N1937, N1777, N728, N910);
or OR4 (N1946, N1942, N386, N1607, N1794);
nand NAND4 (N1947, N1936, N914, N1213, N917);
buf BUF1 (N1948, N1935);
xor XOR2 (N1949, N1946, N719);
not NOT1 (N1950, N1934);
and AND4 (N1951, N1944, N102, N1382, N1835);
nand NAND3 (N1952, N1948, N1892, N188);
buf BUF1 (N1953, N1945);
nand NAND4 (N1954, N1941, N358, N1199, N20);
and AND4 (N1955, N1950, N1071, N1014, N195);
buf BUF1 (N1956, N1954);
buf BUF1 (N1957, N1939);
or OR4 (N1958, N1949, N1322, N1720, N1806);
nand NAND2 (N1959, N1953, N622);
buf BUF1 (N1960, N1956);
xor XOR2 (N1961, N1958, N338);
not NOT1 (N1962, N1961);
buf BUF1 (N1963, N1952);
buf BUF1 (N1964, N1951);
not NOT1 (N1965, N1962);
xor XOR2 (N1966, N1959, N951);
nand NAND3 (N1967, N1957, N54, N1009);
nand NAND2 (N1968, N1927, N454);
or OR4 (N1969, N1960, N983, N1345, N1686);
and AND3 (N1970, N1966, N509, N151);
buf BUF1 (N1971, N1968);
nand NAND3 (N1972, N1955, N1024, N376);
nor NOR3 (N1973, N1964, N499, N1072);
nor NOR2 (N1974, N1970, N1138);
xor XOR2 (N1975, N1947, N32);
and AND2 (N1976, N1969, N1612);
nand NAND3 (N1977, N1973, N1335, N867);
not NOT1 (N1978, N1974);
xor XOR2 (N1979, N1965, N892);
buf BUF1 (N1980, N1979);
buf BUF1 (N1981, N1967);
or OR4 (N1982, N1971, N924, N1018, N95);
nor NOR2 (N1983, N1972, N23);
nor NOR2 (N1984, N1980, N1112);
and AND2 (N1985, N1983, N800);
buf BUF1 (N1986, N1975);
buf BUF1 (N1987, N1977);
xor XOR2 (N1988, N1963, N1548);
buf BUF1 (N1989, N1943);
nand NAND3 (N1990, N1988, N1894, N1928);
nor NOR2 (N1991, N1984, N1742);
buf BUF1 (N1992, N1990);
and AND3 (N1993, N1976, N885, N1968);
buf BUF1 (N1994, N1992);
buf BUF1 (N1995, N1982);
xor XOR2 (N1996, N1986, N841);
nand NAND2 (N1997, N1987, N10);
or OR2 (N1998, N1996, N858);
buf BUF1 (N1999, N1994);
and AND3 (N2000, N1978, N1838, N1871);
xor XOR2 (N2001, N1995, N1266);
buf BUF1 (N2002, N1993);
buf BUF1 (N2003, N2002);
nand NAND2 (N2004, N1991, N939);
buf BUF1 (N2005, N2003);
xor XOR2 (N2006, N1985, N417);
xor XOR2 (N2007, N2006, N1468);
buf BUF1 (N2008, N1989);
nor NOR3 (N2009, N2007, N995, N617);
nor NOR4 (N2010, N1998, N1676, N763, N41);
xor XOR2 (N2011, N1999, N963);
xor XOR2 (N2012, N2004, N1984);
not NOT1 (N2013, N2010);
nand NAND2 (N2014, N2009, N1513);
nand NAND2 (N2015, N2014, N370);
buf BUF1 (N2016, N2005);
buf BUF1 (N2017, N2008);
buf BUF1 (N2018, N2013);
buf BUF1 (N2019, N1981);
nand NAND4 (N2020, N1997, N936, N1942, N326);
or OR3 (N2021, N2020, N337, N432);
xor XOR2 (N2022, N2001, N503);
not NOT1 (N2023, N2022);
not NOT1 (N2024, N2023);
and AND4 (N2025, N2018, N1942, N1860, N867);
buf BUF1 (N2026, N2017);
or OR4 (N2027, N2012, N798, N924, N1322);
xor XOR2 (N2028, N2026, N1091);
and AND4 (N2029, N2028, N1393, N848, N289);
or OR3 (N2030, N2029, N521, N1252);
not NOT1 (N2031, N2019);
and AND4 (N2032, N2000, N1895, N602, N1923);
nor NOR4 (N2033, N2016, N1688, N1128, N589);
not NOT1 (N2034, N2024);
not NOT1 (N2035, N2032);
xor XOR2 (N2036, N2030, N15);
buf BUF1 (N2037, N2035);
nand NAND2 (N2038, N2011, N1394);
xor XOR2 (N2039, N2015, N1919);
and AND3 (N2040, N2031, N380, N1620);
and AND2 (N2041, N2027, N1822);
and AND2 (N2042, N2040, N639);
or OR3 (N2043, N2034, N651, N1412);
and AND2 (N2044, N2041, N284);
buf BUF1 (N2045, N2043);
buf BUF1 (N2046, N2037);
or OR4 (N2047, N2036, N68, N679, N868);
not NOT1 (N2048, N2039);
not NOT1 (N2049, N2045);
or OR4 (N2050, N2038, N485, N1164, N1228);
not NOT1 (N2051, N2042);
buf BUF1 (N2052, N2025);
not NOT1 (N2053, N2021);
or OR2 (N2054, N2053, N901);
buf BUF1 (N2055, N2054);
or OR4 (N2056, N2049, N240, N823, N537);
nor NOR3 (N2057, N2051, N1208, N699);
not NOT1 (N2058, N2033);
nand NAND4 (N2059, N2057, N412, N1603, N1216);
xor XOR2 (N2060, N2056, N822);
buf BUF1 (N2061, N2052);
nor NOR4 (N2062, N2058, N1559, N1401, N317);
and AND2 (N2063, N2059, N532);
and AND3 (N2064, N2063, N1639, N291);
xor XOR2 (N2065, N2061, N106);
or OR4 (N2066, N2062, N528, N202, N11);
buf BUF1 (N2067, N2065);
xor XOR2 (N2068, N2055, N1337);
nor NOR4 (N2069, N2044, N1881, N1040, N679);
or OR3 (N2070, N2060, N1761, N1487);
nor NOR4 (N2071, N2067, N669, N784, N758);
nand NAND4 (N2072, N2048, N779, N1386, N1065);
or OR2 (N2073, N2066, N1854);
not NOT1 (N2074, N2073);
buf BUF1 (N2075, N2064);
xor XOR2 (N2076, N2072, N1675);
or OR2 (N2077, N2069, N1955);
nor NOR2 (N2078, N2077, N1380);
buf BUF1 (N2079, N2071);
xor XOR2 (N2080, N2075, N2038);
nand NAND4 (N2081, N2078, N1406, N829, N1859);
buf BUF1 (N2082, N2079);
buf BUF1 (N2083, N2076);
buf BUF1 (N2084, N2080);
nor NOR3 (N2085, N2050, N1170, N216);
and AND3 (N2086, N2068, N693, N659);
and AND3 (N2087, N2084, N698, N1210);
nor NOR4 (N2088, N2083, N70, N1529, N1038);
and AND4 (N2089, N2082, N115, N1764, N1658);
or OR2 (N2090, N2086, N1664);
buf BUF1 (N2091, N2046);
and AND3 (N2092, N2087, N696, N1999);
not NOT1 (N2093, N2091);
not NOT1 (N2094, N2085);
and AND2 (N2095, N2089, N1188);
or OR4 (N2096, N2088, N141, N1885, N1827);
nor NOR4 (N2097, N2090, N1625, N584, N464);
not NOT1 (N2098, N2093);
or OR2 (N2099, N2096, N456);
buf BUF1 (N2100, N2095);
or OR3 (N2101, N2047, N1393, N1673);
nand NAND4 (N2102, N2081, N1714, N1424, N1114);
buf BUF1 (N2103, N2101);
or OR2 (N2104, N2100, N1432);
nor NOR2 (N2105, N2097, N1640);
nand NAND4 (N2106, N2105, N1116, N677, N108);
buf BUF1 (N2107, N2094);
or OR2 (N2108, N2074, N1039);
buf BUF1 (N2109, N2107);
nand NAND3 (N2110, N2106, N1749, N249);
buf BUF1 (N2111, N2104);
nand NAND3 (N2112, N2102, N571, N1365);
not NOT1 (N2113, N2110);
or OR4 (N2114, N2111, N364, N1138, N1884);
nand NAND2 (N2115, N2112, N13);
not NOT1 (N2116, N2070);
nor NOR3 (N2117, N2115, N1846, N1043);
nor NOR3 (N2118, N2092, N1996, N945);
buf BUF1 (N2119, N2117);
xor XOR2 (N2120, N2119, N1031);
nand NAND4 (N2121, N2113, N1262, N888, N794);
not NOT1 (N2122, N2121);
buf BUF1 (N2123, N2114);
and AND4 (N2124, N2116, N1377, N995, N401);
not NOT1 (N2125, N2098);
nor NOR4 (N2126, N2120, N1592, N1527, N1632);
or OR2 (N2127, N2122, N114);
not NOT1 (N2128, N2127);
xor XOR2 (N2129, N2123, N1025);
nand NAND2 (N2130, N2108, N728);
buf BUF1 (N2131, N2109);
nand NAND3 (N2132, N2130, N1786, N1803);
or OR3 (N2133, N2099, N154, N1197);
xor XOR2 (N2134, N2132, N482);
nand NAND2 (N2135, N2128, N1549);
not NOT1 (N2136, N2131);
and AND2 (N2137, N2126, N1089);
nand NAND2 (N2138, N2137, N1147);
nand NAND4 (N2139, N2136, N1686, N392, N940);
and AND4 (N2140, N2129, N505, N2069, N875);
nor NOR4 (N2141, N2139, N427, N709, N724);
or OR3 (N2142, N2135, N2089, N1325);
and AND2 (N2143, N2118, N1725);
buf BUF1 (N2144, N2124);
not NOT1 (N2145, N2140);
and AND4 (N2146, N2145, N774, N1470, N893);
nand NAND4 (N2147, N2134, N1249, N1091, N131);
not NOT1 (N2148, N2146);
nor NOR3 (N2149, N2144, N735, N2051);
and AND3 (N2150, N2138, N1283, N664);
and AND2 (N2151, N2148, N29);
nand NAND3 (N2152, N2151, N807, N859);
nor NOR3 (N2153, N2142, N1390, N1594);
xor XOR2 (N2154, N2133, N1088);
xor XOR2 (N2155, N2143, N1877);
or OR3 (N2156, N2125, N1128, N1006);
xor XOR2 (N2157, N2155, N1493);
nor NOR2 (N2158, N2147, N1294);
nand NAND3 (N2159, N2141, N1505, N758);
not NOT1 (N2160, N2157);
not NOT1 (N2161, N2160);
buf BUF1 (N2162, N2149);
not NOT1 (N2163, N2158);
xor XOR2 (N2164, N2156, N458);
nand NAND4 (N2165, N2161, N1677, N449, N1562);
or OR4 (N2166, N2165, N2158, N1751, N302);
nand NAND2 (N2167, N2166, N1584);
not NOT1 (N2168, N2103);
and AND2 (N2169, N2154, N1749);
nand NAND4 (N2170, N2168, N1643, N952, N1628);
buf BUF1 (N2171, N2159);
nor NOR3 (N2172, N2162, N2110, N1677);
xor XOR2 (N2173, N2150, N2053);
nand NAND4 (N2174, N2164, N1689, N61, N1501);
nand NAND4 (N2175, N2169, N1960, N1054, N674);
or OR2 (N2176, N2153, N85);
nor NOR3 (N2177, N2167, N690, N994);
or OR2 (N2178, N2170, N611);
buf BUF1 (N2179, N2152);
buf BUF1 (N2180, N2171);
nor NOR2 (N2181, N2172, N237);
and AND4 (N2182, N2163, N503, N1122, N1618);
buf BUF1 (N2183, N2177);
nor NOR2 (N2184, N2176, N2134);
nand NAND3 (N2185, N2183, N212, N850);
and AND4 (N2186, N2174, N325, N1316, N983);
xor XOR2 (N2187, N2179, N646);
or OR4 (N2188, N2173, N1473, N257, N2153);
nor NOR2 (N2189, N2186, N1579);
and AND3 (N2190, N2188, N1890, N1399);
and AND4 (N2191, N2182, N658, N1872, N1281);
xor XOR2 (N2192, N2189, N1858);
or OR3 (N2193, N2192, N476, N1479);
xor XOR2 (N2194, N2178, N1354);
or OR3 (N2195, N2180, N1420, N1389);
buf BUF1 (N2196, N2181);
xor XOR2 (N2197, N2190, N1730);
not NOT1 (N2198, N2196);
buf BUF1 (N2199, N2175);
not NOT1 (N2200, N2187);
xor XOR2 (N2201, N2185, N816);
buf BUF1 (N2202, N2200);
nor NOR2 (N2203, N2193, N1926);
and AND3 (N2204, N2195, N1596, N1533);
not NOT1 (N2205, N2198);
xor XOR2 (N2206, N2201, N1827);
or OR2 (N2207, N2206, N1398);
nor NOR2 (N2208, N2203, N373);
nor NOR2 (N2209, N2194, N1834);
buf BUF1 (N2210, N2205);
not NOT1 (N2211, N2210);
nor NOR4 (N2212, N2207, N432, N1955, N20);
nand NAND3 (N2213, N2191, N340, N300);
nand NAND2 (N2214, N2204, N2050);
nand NAND3 (N2215, N2209, N2021, N828);
xor XOR2 (N2216, N2208, N1062);
nand NAND4 (N2217, N2213, N953, N1740, N914);
buf BUF1 (N2218, N2199);
xor XOR2 (N2219, N2215, N814);
buf BUF1 (N2220, N2197);
nand NAND3 (N2221, N2220, N552, N176);
nor NOR3 (N2222, N2212, N675, N866);
not NOT1 (N2223, N2222);
nor NOR3 (N2224, N2219, N1819, N1983);
not NOT1 (N2225, N2218);
xor XOR2 (N2226, N2225, N1586);
xor XOR2 (N2227, N2221, N769);
or OR4 (N2228, N2223, N1113, N1712, N1398);
not NOT1 (N2229, N2184);
xor XOR2 (N2230, N2217, N1221);
nor NOR4 (N2231, N2229, N1663, N1096, N1390);
nand NAND3 (N2232, N2216, N145, N2148);
or OR3 (N2233, N2228, N48, N973);
buf BUF1 (N2234, N2227);
or OR4 (N2235, N2233, N910, N1456, N835);
and AND3 (N2236, N2231, N968, N1870);
or OR2 (N2237, N2232, N182);
nor NOR3 (N2238, N2234, N334, N1373);
xor XOR2 (N2239, N2238, N744);
or OR4 (N2240, N2235, N86, N148, N1149);
xor XOR2 (N2241, N2239, N187);
or OR4 (N2242, N2236, N2115, N1483, N1369);
nor NOR4 (N2243, N2214, N1486, N474, N812);
or OR4 (N2244, N2241, N27, N1736, N83);
nor NOR2 (N2245, N2244, N1876);
not NOT1 (N2246, N2242);
xor XOR2 (N2247, N2211, N1950);
xor XOR2 (N2248, N2245, N839);
nor NOR2 (N2249, N2247, N1592);
nor NOR2 (N2250, N2202, N1695);
buf BUF1 (N2251, N2226);
or OR3 (N2252, N2224, N714, N909);
nand NAND4 (N2253, N2240, N2154, N664, N2033);
not NOT1 (N2254, N2250);
buf BUF1 (N2255, N2246);
not NOT1 (N2256, N2252);
nor NOR4 (N2257, N2230, N1884, N1925, N400);
and AND2 (N2258, N2237, N1055);
nand NAND3 (N2259, N2257, N1740, N2051);
buf BUF1 (N2260, N2258);
xor XOR2 (N2261, N2251, N279);
xor XOR2 (N2262, N2261, N531);
nor NOR2 (N2263, N2253, N1813);
nor NOR3 (N2264, N2255, N1196, N338);
nor NOR2 (N2265, N2249, N1787);
nand NAND2 (N2266, N2243, N185);
and AND3 (N2267, N2262, N1008, N317);
not NOT1 (N2268, N2248);
not NOT1 (N2269, N2266);
or OR3 (N2270, N2267, N538, N173);
nand NAND4 (N2271, N2268, N229, N203, N1121);
or OR3 (N2272, N2256, N1904, N1581);
and AND2 (N2273, N2265, N2178);
buf BUF1 (N2274, N2263);
xor XOR2 (N2275, N2259, N1631);
nand NAND3 (N2276, N2273, N52, N2190);
nand NAND2 (N2277, N2274, N1153);
nand NAND4 (N2278, N2272, N1669, N1477, N591);
nand NAND4 (N2279, N2276, N1899, N1844, N673);
and AND4 (N2280, N2260, N385, N1189, N1984);
buf BUF1 (N2281, N2270);
not NOT1 (N2282, N2269);
buf BUF1 (N2283, N2282);
nand NAND4 (N2284, N2283, N1362, N1893, N482);
and AND4 (N2285, N2280, N726, N1218, N23);
nor NOR2 (N2286, N2278, N1536);
not NOT1 (N2287, N2275);
or OR2 (N2288, N2264, N731);
xor XOR2 (N2289, N2281, N213);
nand NAND4 (N2290, N2287, N723, N753, N1317);
not NOT1 (N2291, N2277);
nor NOR4 (N2292, N2284, N968, N1067, N883);
not NOT1 (N2293, N2290);
nor NOR2 (N2294, N2292, N1772);
xor XOR2 (N2295, N2285, N791);
xor XOR2 (N2296, N2271, N387);
nand NAND4 (N2297, N2289, N319, N444, N894);
buf BUF1 (N2298, N2293);
nor NOR2 (N2299, N2291, N1377);
and AND2 (N2300, N2298, N935);
or OR2 (N2301, N2286, N1107);
not NOT1 (N2302, N2279);
buf BUF1 (N2303, N2288);
xor XOR2 (N2304, N2295, N146);
buf BUF1 (N2305, N2299);
and AND3 (N2306, N2302, N1761, N1167);
buf BUF1 (N2307, N2306);
xor XOR2 (N2308, N2294, N2032);
nor NOR3 (N2309, N2296, N878, N445);
buf BUF1 (N2310, N2300);
xor XOR2 (N2311, N2305, N1649);
buf BUF1 (N2312, N2311);
and AND3 (N2313, N2304, N1231, N973);
not NOT1 (N2314, N2308);
xor XOR2 (N2315, N2310, N1139);
or OR2 (N2316, N2297, N1234);
buf BUF1 (N2317, N2312);
xor XOR2 (N2318, N2307, N2023);
not NOT1 (N2319, N2303);
and AND4 (N2320, N2317, N753, N1214, N1050);
buf BUF1 (N2321, N2254);
nand NAND4 (N2322, N2320, N175, N1077, N1165);
buf BUF1 (N2323, N2318);
nand NAND3 (N2324, N2309, N26, N1914);
nand NAND4 (N2325, N2316, N397, N489, N1054);
and AND4 (N2326, N2325, N733, N1282, N1735);
nand NAND2 (N2327, N2322, N1910);
not NOT1 (N2328, N2313);
xor XOR2 (N2329, N2328, N1362);
buf BUF1 (N2330, N2319);
xor XOR2 (N2331, N2326, N233);
not NOT1 (N2332, N2323);
nor NOR4 (N2333, N2301, N1160, N2073, N365);
xor XOR2 (N2334, N2327, N1407);
buf BUF1 (N2335, N2331);
not NOT1 (N2336, N2321);
nor NOR3 (N2337, N2314, N401, N90);
buf BUF1 (N2338, N2324);
and AND3 (N2339, N2333, N150, N1572);
nor NOR4 (N2340, N2334, N312, N1462, N80);
buf BUF1 (N2341, N2332);
nand NAND4 (N2342, N2338, N940, N2220, N1814);
nor NOR3 (N2343, N2315, N888, N1733);
not NOT1 (N2344, N2341);
nor NOR4 (N2345, N2337, N1442, N1789, N549);
nor NOR2 (N2346, N2336, N1608);
nand NAND3 (N2347, N2330, N2064, N31);
buf BUF1 (N2348, N2340);
and AND4 (N2349, N2348, N421, N1902, N672);
xor XOR2 (N2350, N2346, N1628);
and AND3 (N2351, N2350, N214, N484);
not NOT1 (N2352, N2351);
or OR4 (N2353, N2347, N1037, N1545, N1762);
and AND4 (N2354, N2329, N1662, N1768, N2107);
nand NAND3 (N2355, N2339, N1912, N1302);
not NOT1 (N2356, N2345);
and AND4 (N2357, N2342, N2114, N371, N126);
xor XOR2 (N2358, N2349, N11);
xor XOR2 (N2359, N2352, N845);
or OR2 (N2360, N2355, N922);
nor NOR2 (N2361, N2360, N1707);
xor XOR2 (N2362, N2354, N1504);
xor XOR2 (N2363, N2357, N2046);
and AND3 (N2364, N2353, N2143, N1237);
buf BUF1 (N2365, N2356);
and AND2 (N2366, N2362, N17);
nand NAND3 (N2367, N2343, N1973, N1937);
nor NOR2 (N2368, N2335, N2231);
and AND4 (N2369, N2367, N154, N1792, N2338);
buf BUF1 (N2370, N2365);
or OR4 (N2371, N2363, N382, N1385, N166);
buf BUF1 (N2372, N2370);
nand NAND2 (N2373, N2358, N1030);
not NOT1 (N2374, N2369);
buf BUF1 (N2375, N2359);
and AND4 (N2376, N2373, N1515, N611, N1904);
nor NOR2 (N2377, N2375, N148);
not NOT1 (N2378, N2344);
nor NOR4 (N2379, N2374, N1762, N1280, N1706);
or OR2 (N2380, N2377, N1709);
and AND2 (N2381, N2372, N1894);
or OR2 (N2382, N2379, N1542);
and AND2 (N2383, N2371, N2330);
or OR2 (N2384, N2381, N258);
or OR2 (N2385, N2366, N1682);
or OR3 (N2386, N2376, N1819, N2075);
or OR4 (N2387, N2383, N58, N20, N555);
and AND3 (N2388, N2378, N693, N2252);
not NOT1 (N2389, N2380);
and AND4 (N2390, N2387, N1347, N285, N2278);
nor NOR2 (N2391, N2389, N1449);
xor XOR2 (N2392, N2391, N534);
nor NOR3 (N2393, N2385, N1130, N929);
not NOT1 (N2394, N2368);
not NOT1 (N2395, N2390);
nor NOR3 (N2396, N2395, N786, N1255);
and AND4 (N2397, N2382, N893, N1327, N2178);
buf BUF1 (N2398, N2388);
and AND4 (N2399, N2364, N570, N505, N909);
or OR3 (N2400, N2399, N1660, N319);
nor NOR2 (N2401, N2392, N2037);
and AND3 (N2402, N2397, N1809, N441);
nor NOR3 (N2403, N2396, N462, N2241);
nor NOR4 (N2404, N2361, N344, N174, N305);
and AND3 (N2405, N2398, N1179, N2348);
xor XOR2 (N2406, N2403, N56);
buf BUF1 (N2407, N2405);
nor NOR4 (N2408, N2407, N1084, N2043, N668);
buf BUF1 (N2409, N2384);
nand NAND4 (N2410, N2393, N555, N1435, N1491);
buf BUF1 (N2411, N2394);
xor XOR2 (N2412, N2386, N711);
xor XOR2 (N2413, N2406, N2156);
and AND3 (N2414, N2413, N2343, N2375);
nor NOR2 (N2415, N2412, N2394);
and AND2 (N2416, N2404, N1504);
not NOT1 (N2417, N2408);
buf BUF1 (N2418, N2411);
not NOT1 (N2419, N2409);
xor XOR2 (N2420, N2417, N2322);
buf BUF1 (N2421, N2400);
nor NOR4 (N2422, N2419, N2014, N1429, N2288);
not NOT1 (N2423, N2418);
and AND2 (N2424, N2416, N1718);
buf BUF1 (N2425, N2415);
or OR3 (N2426, N2423, N2014, N758);
or OR4 (N2427, N2420, N651, N2172, N332);
or OR2 (N2428, N2421, N741);
buf BUF1 (N2429, N2410);
xor XOR2 (N2430, N2427, N975);
or OR3 (N2431, N2428, N1233, N1153);
or OR4 (N2432, N2422, N579, N42, N1933);
not NOT1 (N2433, N2431);
buf BUF1 (N2434, N2433);
and AND2 (N2435, N2432, N10);
buf BUF1 (N2436, N2429);
nor NOR4 (N2437, N2426, N1931, N2362, N2015);
not NOT1 (N2438, N2401);
not NOT1 (N2439, N2430);
nor NOR2 (N2440, N2439, N1567);
nor NOR3 (N2441, N2440, N1771, N1320);
and AND3 (N2442, N2441, N2426, N612);
buf BUF1 (N2443, N2435);
nand NAND3 (N2444, N2424, N2243, N1729);
not NOT1 (N2445, N2442);
not NOT1 (N2446, N2443);
and AND2 (N2447, N2437, N1784);
xor XOR2 (N2448, N2414, N311);
nand NAND4 (N2449, N2445, N1605, N1374, N488);
buf BUF1 (N2450, N2449);
not NOT1 (N2451, N2436);
and AND4 (N2452, N2434, N988, N334, N527);
and AND2 (N2453, N2450, N636);
buf BUF1 (N2454, N2444);
buf BUF1 (N2455, N2425);
xor XOR2 (N2456, N2452, N749);
not NOT1 (N2457, N2456);
not NOT1 (N2458, N2447);
nor NOR4 (N2459, N2448, N1247, N146, N774);
buf BUF1 (N2460, N2438);
or OR4 (N2461, N2460, N920, N400, N1451);
and AND2 (N2462, N2458, N211);
nor NOR3 (N2463, N2457, N990, N2143);
nand NAND4 (N2464, N2446, N871, N883, N2260);
nand NAND4 (N2465, N2454, N702, N2243, N2423);
nand NAND3 (N2466, N2462, N648, N1398);
or OR2 (N2467, N2461, N1960);
buf BUF1 (N2468, N2455);
or OR3 (N2469, N2466, N1143, N1719);
nor NOR4 (N2470, N2467, N1241, N57, N36);
buf BUF1 (N2471, N2464);
nor NOR2 (N2472, N2402, N256);
buf BUF1 (N2473, N2472);
or OR4 (N2474, N2469, N983, N901, N2133);
xor XOR2 (N2475, N2474, N246);
or OR3 (N2476, N2453, N1430, N850);
buf BUF1 (N2477, N2459);
nand NAND2 (N2478, N2475, N1186);
xor XOR2 (N2479, N2477, N1992);
and AND3 (N2480, N2473, N2462, N976);
xor XOR2 (N2481, N2465, N1182);
and AND4 (N2482, N2471, N764, N1080, N1270);
and AND2 (N2483, N2470, N2436);
xor XOR2 (N2484, N2480, N1370);
nand NAND2 (N2485, N2479, N1665);
nor NOR4 (N2486, N2463, N1702, N1309, N579);
not NOT1 (N2487, N2486);
xor XOR2 (N2488, N2482, N1920);
and AND4 (N2489, N2484, N1026, N311, N399);
not NOT1 (N2490, N2487);
buf BUF1 (N2491, N2481);
not NOT1 (N2492, N2489);
not NOT1 (N2493, N2468);
not NOT1 (N2494, N2490);
not NOT1 (N2495, N2476);
not NOT1 (N2496, N2491);
nor NOR2 (N2497, N2494, N1464);
nor NOR4 (N2498, N2488, N1581, N248, N824);
not NOT1 (N2499, N2478);
nand NAND3 (N2500, N2499, N770, N2060);
buf BUF1 (N2501, N2500);
xor XOR2 (N2502, N2493, N841);
not NOT1 (N2503, N2496);
buf BUF1 (N2504, N2503);
nand NAND2 (N2505, N2497, N1490);
or OR4 (N2506, N2498, N1594, N1452, N712);
or OR2 (N2507, N2485, N1897);
buf BUF1 (N2508, N2507);
nor NOR3 (N2509, N2502, N1758, N1209);
or OR2 (N2510, N2509, N1253);
and AND2 (N2511, N2508, N1865);
buf BUF1 (N2512, N2483);
or OR3 (N2513, N2510, N547, N1181);
not NOT1 (N2514, N2451);
nor NOR4 (N2515, N2514, N601, N618, N558);
buf BUF1 (N2516, N2515);
and AND3 (N2517, N2506, N600, N752);
not NOT1 (N2518, N2513);
nor NOR4 (N2519, N2504, N1719, N618, N596);
xor XOR2 (N2520, N2519, N2346);
not NOT1 (N2521, N2516);
nor NOR4 (N2522, N2520, N1988, N1983, N2392);
and AND4 (N2523, N2511, N19, N2050, N526);
xor XOR2 (N2524, N2521, N677);
not NOT1 (N2525, N2495);
or OR4 (N2526, N2522, N1527, N958, N369);
or OR4 (N2527, N2501, N1851, N1506, N515);
xor XOR2 (N2528, N2517, N1746);
or OR2 (N2529, N2523, N1930);
not NOT1 (N2530, N2528);
or OR3 (N2531, N2530, N1085, N292);
xor XOR2 (N2532, N2525, N2264);
nand NAND3 (N2533, N2532, N923, N2417);
nor NOR4 (N2534, N2524, N1291, N741, N533);
not NOT1 (N2535, N2505);
and AND2 (N2536, N2518, N53);
nor NOR4 (N2537, N2531, N2132, N99, N97);
and AND4 (N2538, N2535, N1008, N756, N1508);
and AND3 (N2539, N2529, N2, N471);
or OR3 (N2540, N2492, N873, N1379);
or OR2 (N2541, N2538, N2176);
nand NAND3 (N2542, N2534, N988, N2054);
nor NOR4 (N2543, N2540, N704, N656, N647);
and AND4 (N2544, N2542, N201, N2392, N130);
nor NOR2 (N2545, N2537, N2235);
or OR3 (N2546, N2544, N2069, N2270);
buf BUF1 (N2547, N2539);
nand NAND3 (N2548, N2546, N1926, N133);
xor XOR2 (N2549, N2536, N2141);
not NOT1 (N2550, N2512);
buf BUF1 (N2551, N2547);
nor NOR3 (N2552, N2533, N2351, N1583);
not NOT1 (N2553, N2541);
and AND2 (N2554, N2551, N1948);
xor XOR2 (N2555, N2549, N887);
nand NAND4 (N2556, N2555, N779, N1353, N489);
buf BUF1 (N2557, N2545);
or OR4 (N2558, N2548, N651, N1836, N602);
not NOT1 (N2559, N2553);
or OR2 (N2560, N2526, N1505);
buf BUF1 (N2561, N2527);
buf BUF1 (N2562, N2550);
buf BUF1 (N2563, N2552);
not NOT1 (N2564, N2562);
and AND4 (N2565, N2543, N1497, N1563, N2480);
xor XOR2 (N2566, N2557, N1906);
buf BUF1 (N2567, N2560);
nor NOR4 (N2568, N2567, N428, N1827, N1589);
or OR2 (N2569, N2568, N1146);
nor NOR4 (N2570, N2563, N748, N2294, N939);
buf BUF1 (N2571, N2569);
and AND3 (N2572, N2565, N350, N288);
xor XOR2 (N2573, N2571, N1576);
and AND2 (N2574, N2564, N1457);
xor XOR2 (N2575, N2574, N675);
not NOT1 (N2576, N2573);
not NOT1 (N2577, N2559);
buf BUF1 (N2578, N2558);
nand NAND3 (N2579, N2556, N2334, N2504);
xor XOR2 (N2580, N2570, N1871);
nand NAND4 (N2581, N2554, N2541, N2360, N1575);
and AND3 (N2582, N2577, N2075, N1237);
buf BUF1 (N2583, N2576);
nor NOR2 (N2584, N2582, N230);
nand NAND2 (N2585, N2578, N2352);
nor NOR2 (N2586, N2581, N2255);
nand NAND4 (N2587, N2584, N700, N2314, N1785);
nand NAND3 (N2588, N2579, N1316, N671);
nor NOR4 (N2589, N2588, N1956, N1574, N1703);
or OR3 (N2590, N2589, N1355, N2034);
xor XOR2 (N2591, N2585, N2590);
xor XOR2 (N2592, N358, N591);
or OR4 (N2593, N2580, N2022, N593, N427);
nor NOR4 (N2594, N2575, N202, N1933, N265);
nand NAND3 (N2595, N2591, N2523, N1734);
nand NAND4 (N2596, N2572, N48, N1030, N1030);
buf BUF1 (N2597, N2561);
or OR3 (N2598, N2583, N1872, N104);
buf BUF1 (N2599, N2594);
xor XOR2 (N2600, N2592, N1898);
not NOT1 (N2601, N2596);
or OR2 (N2602, N2598, N1111);
xor XOR2 (N2603, N2602, N1091);
or OR4 (N2604, N2599, N861, N523, N813);
not NOT1 (N2605, N2587);
nand NAND3 (N2606, N2601, N959, N1345);
nor NOR2 (N2607, N2606, N314);
nand NAND2 (N2608, N2593, N1858);
or OR3 (N2609, N2595, N1091, N259);
not NOT1 (N2610, N2603);
and AND4 (N2611, N2610, N1405, N2143, N2200);
and AND2 (N2612, N2600, N2379);
nand NAND4 (N2613, N2609, N2177, N1359, N2573);
or OR2 (N2614, N2613, N2602);
or OR3 (N2615, N2566, N214, N2386);
buf BUF1 (N2616, N2607);
xor XOR2 (N2617, N2605, N1728);
buf BUF1 (N2618, N2586);
buf BUF1 (N2619, N2597);
and AND3 (N2620, N2614, N2210, N1792);
and AND3 (N2621, N2619, N927, N562);
or OR4 (N2622, N2608, N1038, N2272, N1566);
xor XOR2 (N2623, N2621, N1068);
xor XOR2 (N2624, N2618, N281);
and AND2 (N2625, N2623, N878);
nand NAND4 (N2626, N2604, N2602, N110, N1226);
and AND4 (N2627, N2616, N1455, N1841, N1010);
not NOT1 (N2628, N2624);
not NOT1 (N2629, N2620);
buf BUF1 (N2630, N2617);
and AND3 (N2631, N2630, N2059, N2583);
or OR3 (N2632, N2622, N358, N346);
nand NAND2 (N2633, N2629, N227);
nor NOR4 (N2634, N2628, N1361, N1091, N771);
and AND4 (N2635, N2612, N758, N2091, N197);
or OR3 (N2636, N2633, N2339, N1759);
buf BUF1 (N2637, N2611);
and AND2 (N2638, N2615, N1166);
and AND4 (N2639, N2631, N1806, N413, N1157);
nand NAND4 (N2640, N2634, N2539, N2329, N1782);
not NOT1 (N2641, N2627);
not NOT1 (N2642, N2625);
and AND2 (N2643, N2637, N1);
nand NAND4 (N2644, N2632, N1305, N1528, N527);
xor XOR2 (N2645, N2640, N1250);
not NOT1 (N2646, N2645);
or OR4 (N2647, N2636, N2635, N33, N2170);
nand NAND2 (N2648, N1301, N2005);
xor XOR2 (N2649, N2638, N2069);
xor XOR2 (N2650, N2641, N1687);
nor NOR3 (N2651, N2646, N2074, N2290);
buf BUF1 (N2652, N2642);
not NOT1 (N2653, N2647);
or OR2 (N2654, N2651, N302);
nand NAND2 (N2655, N2652, N91);
buf BUF1 (N2656, N2653);
and AND2 (N2657, N2626, N1234);
and AND4 (N2658, N2650, N65, N2595, N1761);
buf BUF1 (N2659, N2657);
buf BUF1 (N2660, N2655);
nand NAND4 (N2661, N2660, N1677, N1919, N231);
nor NOR4 (N2662, N2644, N1121, N2041, N2661);
nand NAND3 (N2663, N2625, N2246, N1774);
nand NAND2 (N2664, N2662, N1219);
and AND2 (N2665, N2663, N2660);
or OR2 (N2666, N2659, N2594);
nor NOR3 (N2667, N2656, N1706, N1409);
not NOT1 (N2668, N2667);
xor XOR2 (N2669, N2639, N1321);
xor XOR2 (N2670, N2649, N293);
nor NOR3 (N2671, N2669, N684, N270);
not NOT1 (N2672, N2666);
not NOT1 (N2673, N2665);
buf BUF1 (N2674, N2673);
nand NAND3 (N2675, N2671, N2240, N2592);
nand NAND3 (N2676, N2643, N144, N1266);
buf BUF1 (N2677, N2658);
or OR2 (N2678, N2664, N1010);
and AND2 (N2679, N2676, N2533);
or OR4 (N2680, N2677, N2366, N2285, N2179);
xor XOR2 (N2681, N2675, N872);
xor XOR2 (N2682, N2668, N186);
xor XOR2 (N2683, N2648, N2525);
nand NAND3 (N2684, N2672, N998, N2552);
nand NAND2 (N2685, N2654, N574);
buf BUF1 (N2686, N2682);
not NOT1 (N2687, N2681);
buf BUF1 (N2688, N2674);
or OR2 (N2689, N2680, N1937);
or OR4 (N2690, N2679, N219, N2539, N411);
or OR4 (N2691, N2670, N1825, N669, N1734);
or OR4 (N2692, N2683, N189, N2474, N1461);
xor XOR2 (N2693, N2686, N2371);
nand NAND2 (N2694, N2688, N2011);
buf BUF1 (N2695, N2691);
nand NAND2 (N2696, N2692, N1145);
nor NOR2 (N2697, N2690, N832);
nand NAND4 (N2698, N2695, N2343, N441, N666);
or OR4 (N2699, N2684, N2072, N444, N2549);
buf BUF1 (N2700, N2685);
and AND3 (N2701, N2694, N857, N2149);
xor XOR2 (N2702, N2700, N728);
xor XOR2 (N2703, N2701, N1701);
nor NOR2 (N2704, N2699, N1678);
nand NAND4 (N2705, N2698, N1509, N2050, N744);
not NOT1 (N2706, N2693);
or OR4 (N2707, N2705, N1755, N557, N1645);
not NOT1 (N2708, N2706);
nor NOR4 (N2709, N2703, N1983, N40, N1);
xor XOR2 (N2710, N2704, N2039);
nand NAND2 (N2711, N2708, N510);
nand NAND3 (N2712, N2710, N94, N997);
nand NAND3 (N2713, N2697, N332, N1076);
buf BUF1 (N2714, N2707);
or OR3 (N2715, N2702, N880, N2590);
or OR3 (N2716, N2678, N534, N2188);
or OR2 (N2717, N2711, N2302);
and AND3 (N2718, N2717, N2337, N1079);
and AND3 (N2719, N2715, N1358, N1996);
or OR3 (N2720, N2689, N1396, N2700);
and AND4 (N2721, N2719, N272, N466, N1496);
or OR3 (N2722, N2687, N1163, N1361);
nor NOR2 (N2723, N2696, N1286);
nor NOR2 (N2724, N2709, N711);
nand NAND4 (N2725, N2712, N1672, N469, N2399);
nor NOR3 (N2726, N2713, N1275, N2098);
or OR4 (N2727, N2725, N1152, N1386, N1670);
not NOT1 (N2728, N2721);
not NOT1 (N2729, N2718);
not NOT1 (N2730, N2716);
buf BUF1 (N2731, N2726);
nor NOR2 (N2732, N2722, N136);
buf BUF1 (N2733, N2731);
xor XOR2 (N2734, N2714, N2497);
not NOT1 (N2735, N2734);
or OR2 (N2736, N2728, N2052);
nor NOR3 (N2737, N2720, N1464, N766);
not NOT1 (N2738, N2730);
not NOT1 (N2739, N2733);
or OR2 (N2740, N2736, N1749);
and AND2 (N2741, N2738, N2462);
nor NOR4 (N2742, N2737, N1482, N307, N1818);
buf BUF1 (N2743, N2735);
xor XOR2 (N2744, N2732, N2733);
buf BUF1 (N2745, N2744);
buf BUF1 (N2746, N2723);
not NOT1 (N2747, N2740);
nor NOR4 (N2748, N2729, N1367, N958, N2206);
and AND4 (N2749, N2741, N1983, N2219, N850);
and AND4 (N2750, N2739, N1650, N1537, N772);
not NOT1 (N2751, N2748);
nand NAND3 (N2752, N2747, N1175, N2720);
or OR2 (N2753, N2742, N2698);
buf BUF1 (N2754, N2752);
buf BUF1 (N2755, N2751);
nor NOR2 (N2756, N2745, N282);
nand NAND3 (N2757, N2755, N2510, N1374);
not NOT1 (N2758, N2753);
nor NOR4 (N2759, N2727, N856, N1960, N2433);
buf BUF1 (N2760, N2749);
buf BUF1 (N2761, N2760);
nand NAND4 (N2762, N2743, N524, N2115, N2061);
or OR2 (N2763, N2750, N670);
xor XOR2 (N2764, N2757, N1053);
nand NAND2 (N2765, N2746, N1592);
xor XOR2 (N2766, N2758, N2472);
nor NOR4 (N2767, N2761, N1155, N601, N15);
not NOT1 (N2768, N2762);
nand NAND3 (N2769, N2724, N443, N2091);
nor NOR3 (N2770, N2766, N1175, N581);
xor XOR2 (N2771, N2756, N2284);
and AND4 (N2772, N2754, N2119, N141, N2650);
nor NOR3 (N2773, N2764, N887, N2263);
or OR2 (N2774, N2772, N2491);
nor NOR4 (N2775, N2763, N1380, N288, N1087);
not NOT1 (N2776, N2767);
and AND3 (N2777, N2770, N486, N2564);
and AND3 (N2778, N2771, N1248, N1136);
nor NOR4 (N2779, N2765, N2618, N2048, N1550);
not NOT1 (N2780, N2777);
nand NAND2 (N2781, N2779, N114);
buf BUF1 (N2782, N2778);
or OR4 (N2783, N2773, N1033, N463, N1569);
nand NAND4 (N2784, N2768, N202, N2673, N1254);
not NOT1 (N2785, N2776);
nor NOR4 (N2786, N2780, N2005, N2343, N264);
buf BUF1 (N2787, N2774);
and AND3 (N2788, N2782, N1497, N1979);
nor NOR3 (N2789, N2785, N1523, N2674);
or OR4 (N2790, N2783, N2034, N2620, N1341);
or OR3 (N2791, N2775, N1360, N1121);
not NOT1 (N2792, N2786);
and AND2 (N2793, N2790, N1091);
not NOT1 (N2794, N2788);
not NOT1 (N2795, N2784);
and AND2 (N2796, N2794, N749);
buf BUF1 (N2797, N2796);
not NOT1 (N2798, N2791);
and AND4 (N2799, N2798, N210, N361, N1623);
nand NAND2 (N2800, N2787, N2409);
nor NOR3 (N2801, N2800, N838, N1380);
xor XOR2 (N2802, N2759, N1557);
buf BUF1 (N2803, N2789);
buf BUF1 (N2804, N2781);
buf BUF1 (N2805, N2795);
nand NAND3 (N2806, N2802, N305, N2793);
nor NOR3 (N2807, N676, N822, N2168);
buf BUF1 (N2808, N2803);
and AND3 (N2809, N2804, N1909, N324);
or OR3 (N2810, N2806, N244, N504);
buf BUF1 (N2811, N2799);
not NOT1 (N2812, N2807);
xor XOR2 (N2813, N2811, N2139);
buf BUF1 (N2814, N2813);
not NOT1 (N2815, N2769);
xor XOR2 (N2816, N2797, N2302);
xor XOR2 (N2817, N2808, N287);
nand NAND4 (N2818, N2801, N2357, N991, N96);
and AND3 (N2819, N2816, N1098, N1401);
nand NAND2 (N2820, N2809, N616);
nand NAND3 (N2821, N2817, N1395, N509);
buf BUF1 (N2822, N2792);
xor XOR2 (N2823, N2805, N1575);
nor NOR2 (N2824, N2823, N382);
nor NOR4 (N2825, N2824, N1267, N680, N302);
not NOT1 (N2826, N2818);
nor NOR2 (N2827, N2820, N1651);
not NOT1 (N2828, N2814);
nor NOR4 (N2829, N2815, N2007, N919, N1219);
not NOT1 (N2830, N2825);
buf BUF1 (N2831, N2827);
nand NAND4 (N2832, N2831, N1585, N239, N2757);
nor NOR4 (N2833, N2812, N1347, N1618, N377);
and AND4 (N2834, N2821, N463, N1494, N310);
or OR4 (N2835, N2810, N4, N2690, N1743);
nor NOR2 (N2836, N2829, N17);
buf BUF1 (N2837, N2833);
not NOT1 (N2838, N2837);
buf BUF1 (N2839, N2832);
buf BUF1 (N2840, N2838);
or OR4 (N2841, N2835, N587, N1655, N2427);
nor NOR3 (N2842, N2834, N95, N2405);
nand NAND4 (N2843, N2822, N2737, N2769, N2050);
or OR4 (N2844, N2826, N556, N696, N890);
or OR2 (N2845, N2819, N2524);
nand NAND3 (N2846, N2844, N1174, N1511);
xor XOR2 (N2847, N2830, N1198);
not NOT1 (N2848, N2840);
nand NAND4 (N2849, N2848, N1057, N213, N1054);
xor XOR2 (N2850, N2843, N1140);
nor NOR2 (N2851, N2847, N2130);
nor NOR2 (N2852, N2850, N2280);
nor NOR3 (N2853, N2841, N518, N2276);
nand NAND3 (N2854, N2846, N794, N109);
and AND3 (N2855, N2851, N361, N1608);
xor XOR2 (N2856, N2854, N2479);
nor NOR4 (N2857, N2839, N2722, N2679, N1903);
and AND3 (N2858, N2852, N2046, N1135);
not NOT1 (N2859, N2856);
xor XOR2 (N2860, N2855, N161);
not NOT1 (N2861, N2853);
nand NAND4 (N2862, N2857, N1208, N1551, N791);
xor XOR2 (N2863, N2842, N613);
nor NOR2 (N2864, N2849, N715);
xor XOR2 (N2865, N2836, N146);
not NOT1 (N2866, N2863);
not NOT1 (N2867, N2862);
nand NAND4 (N2868, N2860, N1171, N1651, N102);
or OR4 (N2869, N2859, N403, N978, N2223);
or OR4 (N2870, N2867, N374, N433, N608);
xor XOR2 (N2871, N2864, N2513);
buf BUF1 (N2872, N2866);
nand NAND2 (N2873, N2861, N980);
nor NOR3 (N2874, N2828, N2757, N126);
nand NAND3 (N2875, N2865, N1349, N997);
not NOT1 (N2876, N2868);
buf BUF1 (N2877, N2845);
nor NOR3 (N2878, N2876, N2289, N1905);
or OR2 (N2879, N2878, N2842);
not NOT1 (N2880, N2873);
not NOT1 (N2881, N2870);
buf BUF1 (N2882, N2877);
nand NAND3 (N2883, N2874, N1887, N1042);
and AND2 (N2884, N2882, N1087);
buf BUF1 (N2885, N2872);
nand NAND4 (N2886, N2875, N1864, N2585, N2703);
nor NOR4 (N2887, N2884, N157, N2378, N1525);
nor NOR2 (N2888, N2883, N449);
buf BUF1 (N2889, N2858);
not NOT1 (N2890, N2885);
or OR4 (N2891, N2890, N1016, N1838, N2112);
xor XOR2 (N2892, N2871, N2535);
not NOT1 (N2893, N2886);
and AND2 (N2894, N2892, N148);
and AND2 (N2895, N2880, N2056);
and AND3 (N2896, N2894, N209, N541);
buf BUF1 (N2897, N2895);
not NOT1 (N2898, N2893);
and AND4 (N2899, N2881, N1387, N260, N635);
buf BUF1 (N2900, N2896);
and AND4 (N2901, N2889, N399, N1226, N1147);
buf BUF1 (N2902, N2900);
or OR3 (N2903, N2887, N72, N463);
xor XOR2 (N2904, N2898, N1851);
nor NOR4 (N2905, N2904, N724, N1284, N2577);
buf BUF1 (N2906, N2888);
not NOT1 (N2907, N2879);
or OR2 (N2908, N2907, N2824);
nor NOR2 (N2909, N2901, N1241);
and AND4 (N2910, N2905, N1098, N1203, N2541);
nand NAND2 (N2911, N2903, N774);
buf BUF1 (N2912, N2911);
buf BUF1 (N2913, N2902);
or OR3 (N2914, N2899, N232, N690);
buf BUF1 (N2915, N2913);
or OR3 (N2916, N2914, N2563, N2275);
buf BUF1 (N2917, N2912);
nand NAND3 (N2918, N2897, N204, N2452);
and AND2 (N2919, N2906, N1719);
xor XOR2 (N2920, N2919, N792);
nand NAND3 (N2921, N2917, N2245, N1418);
not NOT1 (N2922, N2891);
nand NAND4 (N2923, N2916, N2875, N1718, N80);
nor NOR3 (N2924, N2909, N2503, N2342);
or OR4 (N2925, N2924, N1674, N1013, N1783);
xor XOR2 (N2926, N2920, N357);
xor XOR2 (N2927, N2921, N231);
nor NOR3 (N2928, N2869, N1532, N358);
and AND2 (N2929, N2915, N2665);
buf BUF1 (N2930, N2918);
or OR2 (N2931, N2923, N1624);
or OR3 (N2932, N2910, N2218, N1718);
not NOT1 (N2933, N2928);
not NOT1 (N2934, N2927);
buf BUF1 (N2935, N2931);
nand NAND2 (N2936, N2930, N1682);
xor XOR2 (N2937, N2925, N2785);
xor XOR2 (N2938, N2932, N2055);
or OR4 (N2939, N2933, N2691, N1761, N1950);
and AND3 (N2940, N2929, N632, N1937);
nor NOR4 (N2941, N2940, N2313, N2664, N1019);
nor NOR2 (N2942, N2936, N71);
buf BUF1 (N2943, N2937);
and AND4 (N2944, N2941, N2448, N29, N1202);
nand NAND3 (N2945, N2934, N106, N891);
not NOT1 (N2946, N2945);
nor NOR4 (N2947, N2926, N1952, N390, N1044);
nand NAND4 (N2948, N2943, N136, N1595, N571);
nor NOR3 (N2949, N2922, N739, N2786);
nand NAND4 (N2950, N2949, N689, N534, N420);
nor NOR4 (N2951, N2944, N1853, N515, N1368);
nand NAND4 (N2952, N2951, N2309, N2576, N1202);
and AND3 (N2953, N2938, N2821, N296);
or OR3 (N2954, N2935, N91, N241);
not NOT1 (N2955, N2953);
xor XOR2 (N2956, N2950, N1050);
buf BUF1 (N2957, N2946);
or OR3 (N2958, N2939, N2730, N703);
nor NOR2 (N2959, N2952, N2187);
xor XOR2 (N2960, N2954, N2246);
buf BUF1 (N2961, N2960);
and AND2 (N2962, N2961, N894);
xor XOR2 (N2963, N2956, N2571);
buf BUF1 (N2964, N2908);
not NOT1 (N2965, N2959);
xor XOR2 (N2966, N2957, N2644);
not NOT1 (N2967, N2955);
nor NOR2 (N2968, N2942, N281);
buf BUF1 (N2969, N2963);
xor XOR2 (N2970, N2966, N2495);
and AND3 (N2971, N2958, N2121, N2539);
and AND2 (N2972, N2967, N1334);
nor NOR2 (N2973, N2962, N1280);
or OR4 (N2974, N2947, N601, N2286, N1146);
and AND4 (N2975, N2973, N1167, N2437, N345);
not NOT1 (N2976, N2971);
and AND2 (N2977, N2976, N1045);
and AND2 (N2978, N2965, N917);
not NOT1 (N2979, N2977);
not NOT1 (N2980, N2968);
not NOT1 (N2981, N2980);
buf BUF1 (N2982, N2948);
or OR4 (N2983, N2964, N1243, N2828, N659);
buf BUF1 (N2984, N2972);
and AND4 (N2985, N2978, N63, N200, N2671);
and AND2 (N2986, N2984, N1441);
and AND4 (N2987, N2985, N2813, N920, N1003);
or OR2 (N2988, N2970, N2754);
or OR3 (N2989, N2982, N2490, N2488);
nand NAND4 (N2990, N2979, N510, N2743, N193);
nor NOR2 (N2991, N2969, N196);
xor XOR2 (N2992, N2991, N1341);
buf BUF1 (N2993, N2990);
xor XOR2 (N2994, N2993, N1776);
or OR2 (N2995, N2983, N1513);
not NOT1 (N2996, N2974);
nor NOR4 (N2997, N2992, N1835, N1295, N16);
not NOT1 (N2998, N2988);
nor NOR4 (N2999, N2989, N2647, N1856, N68);
buf BUF1 (N3000, N2981);
nor NOR3 (N3001, N2975, N943, N1845);
and AND3 (N3002, N2995, N1590, N1266);
buf BUF1 (N3003, N2998);
nor NOR2 (N3004, N3000, N2105);
not NOT1 (N3005, N2997);
xor XOR2 (N3006, N2999, N2500);
xor XOR2 (N3007, N2996, N1185);
buf BUF1 (N3008, N3006);
and AND4 (N3009, N3008, N2144, N1502, N2902);
or OR2 (N3010, N3007, N2639);
buf BUF1 (N3011, N2994);
nand NAND4 (N3012, N3010, N489, N1814, N1033);
buf BUF1 (N3013, N3012);
or OR2 (N3014, N3005, N2792);
xor XOR2 (N3015, N3004, N2529);
nand NAND2 (N3016, N3013, N378);
buf BUF1 (N3017, N3016);
and AND2 (N3018, N3015, N1097);
xor XOR2 (N3019, N3003, N2087);
or OR4 (N3020, N3002, N2400, N335, N2861);
xor XOR2 (N3021, N3009, N221);
nand NAND4 (N3022, N3020, N976, N2742, N988);
or OR4 (N3023, N3017, N2637, N1359, N2286);
not NOT1 (N3024, N3022);
nand NAND3 (N3025, N2986, N670, N696);
nand NAND3 (N3026, N3011, N2352, N1269);
xor XOR2 (N3027, N3001, N2073);
xor XOR2 (N3028, N2987, N2586);
nand NAND3 (N3029, N3019, N2968, N708);
buf BUF1 (N3030, N3018);
nand NAND4 (N3031, N3030, N1622, N2238, N1974);
or OR3 (N3032, N3029, N1206, N1058);
buf BUF1 (N3033, N3031);
or OR2 (N3034, N3033, N1347);
and AND2 (N3035, N3028, N235);
xor XOR2 (N3036, N3021, N143);
not NOT1 (N3037, N3024);
nor NOR2 (N3038, N3026, N1612);
not NOT1 (N3039, N3025);
nor NOR4 (N3040, N3032, N364, N112, N1088);
not NOT1 (N3041, N3023);
nand NAND2 (N3042, N3038, N2787);
nor NOR3 (N3043, N3037, N2838, N809);
not NOT1 (N3044, N3036);
nor NOR3 (N3045, N3041, N258, N1835);
or OR2 (N3046, N3034, N1667);
buf BUF1 (N3047, N3046);
and AND4 (N3048, N3047, N2982, N1948, N47);
not NOT1 (N3049, N3042);
or OR2 (N3050, N3014, N2021);
and AND4 (N3051, N3049, N531, N230, N186);
or OR3 (N3052, N3040, N394, N831);
nand NAND4 (N3053, N3052, N198, N1788, N1081);
nor NOR4 (N3054, N3035, N2802, N68, N1129);
nand NAND2 (N3055, N3048, N1138);
not NOT1 (N3056, N3044);
or OR4 (N3057, N3043, N3030, N1294, N2118);
xor XOR2 (N3058, N3051, N2971);
and AND3 (N3059, N3055, N2875, N377);
nand NAND2 (N3060, N3054, N433);
and AND4 (N3061, N3060, N1646, N2303, N657);
xor XOR2 (N3062, N3057, N389);
and AND3 (N3063, N3056, N853, N650);
or OR2 (N3064, N3062, N583);
and AND4 (N3065, N3058, N848, N1253, N3004);
and AND2 (N3066, N3061, N1739);
xor XOR2 (N3067, N3053, N95);
nor NOR4 (N3068, N3045, N1300, N1581, N1847);
xor XOR2 (N3069, N3065, N1489);
buf BUF1 (N3070, N3067);
nor NOR3 (N3071, N3027, N621, N499);
nor NOR3 (N3072, N3064, N2914, N1809);
nand NAND3 (N3073, N3071, N1337, N2175);
not NOT1 (N3074, N3072);
or OR2 (N3075, N3070, N571);
not NOT1 (N3076, N3069);
and AND2 (N3077, N3059, N1917);
not NOT1 (N3078, N3050);
and AND3 (N3079, N3068, N136, N548);
not NOT1 (N3080, N3066);
nor NOR2 (N3081, N3063, N2387);
and AND4 (N3082, N3073, N212, N553, N540);
nand NAND2 (N3083, N3039, N746);
nand NAND2 (N3084, N3078, N3065);
nor NOR2 (N3085, N3076, N642);
or OR4 (N3086, N3085, N543, N1204, N2402);
and AND4 (N3087, N3084, N1536, N13, N177);
nand NAND2 (N3088, N3080, N2106);
not NOT1 (N3089, N3088);
nor NOR4 (N3090, N3077, N1156, N2137, N620);
xor XOR2 (N3091, N3089, N1381);
not NOT1 (N3092, N3074);
not NOT1 (N3093, N3086);
not NOT1 (N3094, N3087);
not NOT1 (N3095, N3090);
buf BUF1 (N3096, N3094);
nand NAND2 (N3097, N3075, N2596);
not NOT1 (N3098, N3091);
not NOT1 (N3099, N3096);
nor NOR4 (N3100, N3092, N782, N1578, N2218);
nand NAND3 (N3101, N3079, N2288, N1254);
and AND2 (N3102, N3095, N1788);
not NOT1 (N3103, N3101);
buf BUF1 (N3104, N3082);
buf BUF1 (N3105, N3093);
not NOT1 (N3106, N3083);
and AND2 (N3107, N3100, N498);
not NOT1 (N3108, N3103);
nand NAND4 (N3109, N3105, N388, N1564, N2972);
not NOT1 (N3110, N3097);
or OR3 (N3111, N3110, N1397, N2711);
not NOT1 (N3112, N3099);
buf BUF1 (N3113, N3098);
and AND3 (N3114, N3102, N1648, N2860);
nand NAND2 (N3115, N3108, N320);
buf BUF1 (N3116, N3114);
xor XOR2 (N3117, N3081, N1584);
nand NAND3 (N3118, N3113, N1066, N1005);
buf BUF1 (N3119, N3112);
or OR2 (N3120, N3106, N681);
nor NOR4 (N3121, N3104, N392, N928, N730);
not NOT1 (N3122, N3107);
nand NAND2 (N3123, N3111, N2333);
not NOT1 (N3124, N3117);
or OR4 (N3125, N3115, N154, N895, N2212);
or OR3 (N3126, N3119, N684, N2304);
and AND2 (N3127, N3123, N125);
xor XOR2 (N3128, N3127, N2617);
nand NAND4 (N3129, N3124, N1802, N2327, N144);
or OR3 (N3130, N3120, N2294, N1058);
nand NAND4 (N3131, N3121, N2738, N1800, N1410);
and AND3 (N3132, N3122, N1506, N1314);
nand NAND4 (N3133, N3118, N1475, N1944, N1926);
buf BUF1 (N3134, N3131);
nor NOR2 (N3135, N3125, N1076);
nor NOR3 (N3136, N3130, N3004, N1682);
nand NAND3 (N3137, N3135, N1705, N735);
nor NOR4 (N3138, N3116, N1416, N1099, N3049);
or OR4 (N3139, N3128, N2974, N439, N424);
nand NAND4 (N3140, N3132, N1042, N2544, N1960);
not NOT1 (N3141, N3137);
or OR4 (N3142, N3136, N2344, N2370, N2110);
and AND3 (N3143, N3141, N4, N174);
not NOT1 (N3144, N3126);
not NOT1 (N3145, N3144);
nand NAND3 (N3146, N3143, N175, N306);
and AND2 (N3147, N3139, N2390);
nor NOR3 (N3148, N3146, N1757, N2129);
nor NOR4 (N3149, N3129, N2905, N2071, N2433);
or OR4 (N3150, N3133, N2385, N163, N408);
or OR3 (N3151, N3142, N1929, N937);
nand NAND4 (N3152, N3145, N1574, N1066, N418);
or OR3 (N3153, N3109, N744, N1883);
nand NAND2 (N3154, N3149, N3003);
and AND2 (N3155, N3138, N1277);
or OR3 (N3156, N3134, N348, N76);
buf BUF1 (N3157, N3150);
nor NOR4 (N3158, N3154, N615, N1455, N788);
buf BUF1 (N3159, N3157);
or OR2 (N3160, N3156, N1469);
nand NAND3 (N3161, N3160, N1155, N1392);
nor NOR2 (N3162, N3152, N2869);
and AND3 (N3163, N3140, N2529, N661);
buf BUF1 (N3164, N3159);
nand NAND4 (N3165, N3163, N648, N792, N808);
or OR4 (N3166, N3165, N1896, N1925, N927);
buf BUF1 (N3167, N3158);
nor NOR3 (N3168, N3162, N2841, N55);
xor XOR2 (N3169, N3153, N2937);
xor XOR2 (N3170, N3167, N810);
not NOT1 (N3171, N3147);
or OR4 (N3172, N3161, N194, N533, N1719);
buf BUF1 (N3173, N3151);
nand NAND4 (N3174, N3171, N1321, N2807, N2086);
xor XOR2 (N3175, N3169, N2428);
buf BUF1 (N3176, N3166);
xor XOR2 (N3177, N3170, N2449);
and AND2 (N3178, N3175, N1604);
buf BUF1 (N3179, N3164);
not NOT1 (N3180, N3178);
buf BUF1 (N3181, N3176);
nor NOR2 (N3182, N3168, N461);
xor XOR2 (N3183, N3182, N1865);
and AND4 (N3184, N3183, N2782, N3045, N1465);
or OR3 (N3185, N3180, N2781, N1898);
or OR2 (N3186, N3155, N1736);
nand NAND4 (N3187, N3148, N753, N676, N3155);
and AND3 (N3188, N3187, N2868, N2662);
nand NAND4 (N3189, N3181, N843, N3036, N1857);
xor XOR2 (N3190, N3173, N1908);
and AND4 (N3191, N3184, N1963, N2154, N884);
nand NAND3 (N3192, N3188, N1440, N3079);
not NOT1 (N3193, N3179);
or OR4 (N3194, N3186, N458, N2703, N1544);
nand NAND2 (N3195, N3189, N953);
or OR4 (N3196, N3185, N438, N22, N1155);
nor NOR2 (N3197, N3193, N232);
xor XOR2 (N3198, N3172, N1005);
nand NAND2 (N3199, N3196, N2618);
buf BUF1 (N3200, N3198);
nand NAND2 (N3201, N3199, N1421);
nor NOR2 (N3202, N3192, N1781);
and AND3 (N3203, N3201, N2388, N752);
buf BUF1 (N3204, N3197);
and AND4 (N3205, N3200, N1347, N1359, N1548);
nand NAND3 (N3206, N3194, N3157, N1971);
nor NOR4 (N3207, N3202, N946, N2714, N564);
nand NAND2 (N3208, N3204, N858);
buf BUF1 (N3209, N3208);
nand NAND2 (N3210, N3177, N1743);
and AND2 (N3211, N3210, N3133);
or OR2 (N3212, N3203, N2762);
nand NAND2 (N3213, N3206, N1339);
nor NOR3 (N3214, N3191, N1183, N1822);
not NOT1 (N3215, N3213);
buf BUF1 (N3216, N3205);
nand NAND2 (N3217, N3190, N1537);
nor NOR3 (N3218, N3216, N2922, N1136);
nor NOR4 (N3219, N3174, N1851, N2098, N2563);
nor NOR4 (N3220, N3218, N1516, N2860, N998);
or OR4 (N3221, N3214, N1005, N147, N1111);
buf BUF1 (N3222, N3209);
or OR4 (N3223, N3212, N2093, N1453, N1217);
nand NAND3 (N3224, N3221, N2808, N119);
nor NOR3 (N3225, N3207, N1225, N2349);
nor NOR2 (N3226, N3211, N354);
xor XOR2 (N3227, N3220, N2069);
and AND2 (N3228, N3223, N1190);
xor XOR2 (N3229, N3227, N1346);
not NOT1 (N3230, N3226);
and AND3 (N3231, N3195, N54, N2152);
xor XOR2 (N3232, N3215, N38);
xor XOR2 (N3233, N3232, N115);
buf BUF1 (N3234, N3231);
buf BUF1 (N3235, N3217);
nand NAND3 (N3236, N3230, N1214, N1648);
buf BUF1 (N3237, N3224);
and AND4 (N3238, N3236, N993, N869, N1352);
nor NOR4 (N3239, N3228, N3139, N2988, N485);
or OR4 (N3240, N3238, N1478, N2172, N574);
buf BUF1 (N3241, N3222);
buf BUF1 (N3242, N3225);
xor XOR2 (N3243, N3229, N2902);
not NOT1 (N3244, N3233);
not NOT1 (N3245, N3237);
xor XOR2 (N3246, N3243, N2742);
and AND4 (N3247, N3240, N895, N472, N253);
buf BUF1 (N3248, N3235);
not NOT1 (N3249, N3234);
buf BUF1 (N3250, N3242);
buf BUF1 (N3251, N3241);
nand NAND2 (N3252, N3249, N306);
or OR3 (N3253, N3247, N1701, N2743);
nor NOR4 (N3254, N3245, N2758, N11, N473);
or OR2 (N3255, N3253, N1863);
not NOT1 (N3256, N3244);
or OR2 (N3257, N3251, N1564);
nor NOR2 (N3258, N3255, N28);
buf BUF1 (N3259, N3257);
xor XOR2 (N3260, N3250, N186);
buf BUF1 (N3261, N3246);
nand NAND3 (N3262, N3252, N2691, N2884);
buf BUF1 (N3263, N3219);
xor XOR2 (N3264, N3256, N780);
xor XOR2 (N3265, N3264, N717);
buf BUF1 (N3266, N3260);
buf BUF1 (N3267, N3259);
xor XOR2 (N3268, N3266, N1380);
buf BUF1 (N3269, N3239);
or OR4 (N3270, N3267, N2044, N971, N2760);
and AND2 (N3271, N3270, N1576);
and AND2 (N3272, N3268, N2294);
not NOT1 (N3273, N3261);
not NOT1 (N3274, N3271);
not NOT1 (N3275, N3265);
nand NAND3 (N3276, N3254, N1880, N2471);
not NOT1 (N3277, N3262);
nor NOR4 (N3278, N3276, N2475, N487, N2605);
and AND4 (N3279, N3277, N1766, N3041, N2280);
and AND3 (N3280, N3269, N2779, N2731);
or OR3 (N3281, N3248, N1961, N1134);
not NOT1 (N3282, N3281);
buf BUF1 (N3283, N3263);
xor XOR2 (N3284, N3279, N57);
buf BUF1 (N3285, N3282);
nor NOR4 (N3286, N3272, N2443, N1011, N1028);
or OR2 (N3287, N3286, N1514);
nor NOR3 (N3288, N3285, N3064, N1431);
nand NAND3 (N3289, N3284, N2255, N1475);
buf BUF1 (N3290, N3275);
buf BUF1 (N3291, N3290);
or OR3 (N3292, N3283, N1885, N235);
nor NOR2 (N3293, N3291, N3236);
xor XOR2 (N3294, N3287, N3126);
not NOT1 (N3295, N3273);
nor NOR3 (N3296, N3280, N283, N15);
buf BUF1 (N3297, N3274);
and AND4 (N3298, N3296, N2008, N430, N1355);
nor NOR2 (N3299, N3292, N1877);
or OR4 (N3300, N3294, N3148, N2927, N2021);
and AND2 (N3301, N3295, N2893);
and AND2 (N3302, N3297, N735);
nand NAND4 (N3303, N3301, N2761, N2487, N3105);
and AND2 (N3304, N3302, N2663);
or OR2 (N3305, N3298, N2581);
and AND3 (N3306, N3258, N1294, N1291);
nand NAND4 (N3307, N3300, N1594, N1630, N1293);
xor XOR2 (N3308, N3278, N547);
nor NOR4 (N3309, N3308, N777, N1099, N2523);
or OR2 (N3310, N3309, N920);
nor NOR2 (N3311, N3310, N197);
and AND3 (N3312, N3307, N128, N968);
nand NAND2 (N3313, N3288, N2718);
xor XOR2 (N3314, N3304, N13);
buf BUF1 (N3315, N3303);
buf BUF1 (N3316, N3314);
xor XOR2 (N3317, N3306, N2963);
buf BUF1 (N3318, N3317);
and AND2 (N3319, N3318, N2316);
or OR3 (N3320, N3289, N2978, N1537);
xor XOR2 (N3321, N3305, N2716);
not NOT1 (N3322, N3321);
buf BUF1 (N3323, N3322);
and AND2 (N3324, N3312, N183);
buf BUF1 (N3325, N3299);
xor XOR2 (N3326, N3311, N2241);
xor XOR2 (N3327, N3313, N373);
nor NOR2 (N3328, N3324, N1208);
buf BUF1 (N3329, N3323);
nor NOR2 (N3330, N3320, N147);
or OR4 (N3331, N3327, N447, N1550, N1510);
nor NOR3 (N3332, N3319, N346, N1572);
nor NOR3 (N3333, N3293, N1089, N1612);
and AND2 (N3334, N3315, N2578);
nor NOR3 (N3335, N3330, N905, N1193);
nor NOR3 (N3336, N3325, N3179, N2631);
buf BUF1 (N3337, N3336);
buf BUF1 (N3338, N3333);
or OR2 (N3339, N3331, N3174);
nor NOR2 (N3340, N3329, N1751);
xor XOR2 (N3341, N3332, N1398);
not NOT1 (N3342, N3335);
nand NAND2 (N3343, N3340, N631);
and AND4 (N3344, N3343, N3335, N246, N3256);
xor XOR2 (N3345, N3337, N1662);
nor NOR2 (N3346, N3316, N1498);
or OR3 (N3347, N3339, N788, N1804);
or OR4 (N3348, N3344, N1575, N1268, N1191);
not NOT1 (N3349, N3345);
or OR2 (N3350, N3348, N2532);
not NOT1 (N3351, N3346);
xor XOR2 (N3352, N3351, N1962);
nand NAND4 (N3353, N3342, N3341, N948, N2470);
xor XOR2 (N3354, N1078, N1107);
and AND2 (N3355, N3349, N3305);
and AND4 (N3356, N3334, N3203, N3287, N143);
not NOT1 (N3357, N3338);
and AND3 (N3358, N3350, N2684, N1796);
not NOT1 (N3359, N3328);
or OR4 (N3360, N3356, N1613, N2770, N2888);
not NOT1 (N3361, N3352);
and AND4 (N3362, N3357, N2858, N1020, N2303);
buf BUF1 (N3363, N3347);
nor NOR2 (N3364, N3355, N894);
or OR2 (N3365, N3359, N2560);
nor NOR3 (N3366, N3326, N696, N2424);
xor XOR2 (N3367, N3364, N884);
or OR4 (N3368, N3354, N3357, N1428, N2623);
nand NAND3 (N3369, N3368, N3180, N376);
not NOT1 (N3370, N3360);
buf BUF1 (N3371, N3363);
xor XOR2 (N3372, N3358, N3295);
and AND4 (N3373, N3365, N787, N1602, N964);
buf BUF1 (N3374, N3367);
and AND4 (N3375, N3371, N1272, N392, N1887);
nor NOR4 (N3376, N3373, N1515, N884, N305);
and AND3 (N3377, N3370, N388, N199);
or OR4 (N3378, N3361, N1712, N852, N1038);
nand NAND4 (N3379, N3375, N3241, N2489, N2531);
nand NAND2 (N3380, N3372, N342);
not NOT1 (N3381, N3374);
not NOT1 (N3382, N3376);
buf BUF1 (N3383, N3366);
or OR2 (N3384, N3362, N1250);
and AND4 (N3385, N3383, N2725, N1891, N905);
xor XOR2 (N3386, N3379, N2032);
nand NAND3 (N3387, N3384, N2438, N1479);
nand NAND4 (N3388, N3385, N1558, N2217, N2116);
not NOT1 (N3389, N3380);
or OR2 (N3390, N3381, N1687);
and AND3 (N3391, N3386, N3389, N238);
or OR2 (N3392, N1421, N3081);
xor XOR2 (N3393, N3390, N1311);
and AND4 (N3394, N3369, N1398, N593, N815);
not NOT1 (N3395, N3353);
buf BUF1 (N3396, N3388);
nand NAND2 (N3397, N3391, N2803);
nor NOR4 (N3398, N3382, N1096, N133, N2925);
xor XOR2 (N3399, N3387, N58);
nor NOR4 (N3400, N3377, N1267, N2507, N159);
or OR4 (N3401, N3398, N1290, N1459, N2762);
not NOT1 (N3402, N3378);
buf BUF1 (N3403, N3401);
nand NAND2 (N3404, N3402, N3272);
not NOT1 (N3405, N3393);
or OR2 (N3406, N3405, N800);
not NOT1 (N3407, N3403);
xor XOR2 (N3408, N3397, N301);
and AND4 (N3409, N3394, N304, N837, N2835);
and AND2 (N3410, N3399, N1352);
not NOT1 (N3411, N3400);
xor XOR2 (N3412, N3406, N433);
not NOT1 (N3413, N3392);
or OR4 (N3414, N3395, N556, N499, N2424);
not NOT1 (N3415, N3411);
buf BUF1 (N3416, N3412);
xor XOR2 (N3417, N3396, N1510);
buf BUF1 (N3418, N3413);
or OR4 (N3419, N3404, N365, N24, N1621);
nand NAND3 (N3420, N3408, N2038, N303);
and AND2 (N3421, N3407, N2271);
xor XOR2 (N3422, N3410, N1286);
nand NAND4 (N3423, N3422, N1593, N1052, N386);
xor XOR2 (N3424, N3414, N110);
buf BUF1 (N3425, N3420);
and AND4 (N3426, N3415, N3306, N973, N1818);
nand NAND2 (N3427, N3423, N1262);
nand NAND3 (N3428, N3425, N1212, N2700);
or OR3 (N3429, N3419, N113, N1883);
or OR4 (N3430, N3421, N2224, N2793, N2848);
nor NOR4 (N3431, N3427, N3233, N3037, N2781);
and AND2 (N3432, N3431, N3186);
xor XOR2 (N3433, N3426, N1296);
and AND4 (N3434, N3409, N2119, N3237, N810);
not NOT1 (N3435, N3418);
buf BUF1 (N3436, N3424);
not NOT1 (N3437, N3430);
nor NOR4 (N3438, N3432, N1253, N3149, N292);
nor NOR2 (N3439, N3436, N2476);
and AND4 (N3440, N3439, N3385, N3014, N606);
nor NOR4 (N3441, N3435, N2814, N2511, N1768);
xor XOR2 (N3442, N3428, N2162);
nor NOR3 (N3443, N3417, N3357, N2660);
buf BUF1 (N3444, N3416);
buf BUF1 (N3445, N3443);
nor NOR4 (N3446, N3438, N1502, N3441, N1885);
not NOT1 (N3447, N2997);
buf BUF1 (N3448, N3442);
xor XOR2 (N3449, N3433, N3347);
and AND4 (N3450, N3444, N449, N903, N983);
buf BUF1 (N3451, N3440);
and AND4 (N3452, N3450, N1810, N3115, N1706);
and AND3 (N3453, N3447, N3313, N2971);
and AND4 (N3454, N3434, N1663, N799, N3373);
buf BUF1 (N3455, N3446);
nand NAND3 (N3456, N3455, N535, N2675);
and AND3 (N3457, N3454, N1889, N3167);
and AND4 (N3458, N3449, N1739, N1616, N2264);
xor XOR2 (N3459, N3452, N1825);
buf BUF1 (N3460, N3445);
and AND4 (N3461, N3451, N1605, N835, N3271);
not NOT1 (N3462, N3448);
nor NOR4 (N3463, N3462, N1805, N2427, N3176);
and AND4 (N3464, N3460, N199, N2518, N650);
not NOT1 (N3465, N3461);
nand NAND4 (N3466, N3437, N2409, N450, N2218);
nor NOR3 (N3467, N3465, N837, N1215);
or OR2 (N3468, N3463, N2465);
nor NOR3 (N3469, N3464, N2403, N3435);
nand NAND2 (N3470, N3467, N1737);
and AND3 (N3471, N3458, N140, N3186);
nor NOR3 (N3472, N3471, N2098, N1494);
or OR3 (N3473, N3469, N2509, N86);
buf BUF1 (N3474, N3456);
xor XOR2 (N3475, N3457, N2920);
or OR4 (N3476, N3474, N2853, N3062, N1173);
xor XOR2 (N3477, N3472, N2427);
xor XOR2 (N3478, N3429, N2396);
or OR2 (N3479, N3475, N368);
not NOT1 (N3480, N3473);
nand NAND2 (N3481, N3453, N2438);
or OR3 (N3482, N3476, N1007, N936);
and AND2 (N3483, N3459, N1180);
or OR3 (N3484, N3477, N2781, N2823);
and AND4 (N3485, N3484, N2260, N1354, N1118);
or OR4 (N3486, N3470, N2152, N1155, N2715);
xor XOR2 (N3487, N3483, N216);
nor NOR3 (N3488, N3480, N675, N2389);
buf BUF1 (N3489, N3487);
nor NOR3 (N3490, N3468, N153, N2417);
or OR2 (N3491, N3466, N582);
nand NAND3 (N3492, N3481, N3459, N720);
or OR4 (N3493, N3478, N2226, N3174, N130);
and AND2 (N3494, N3482, N1425);
nor NOR4 (N3495, N3479, N549, N2936, N2838);
nor NOR4 (N3496, N3490, N1383, N2362, N2381);
buf BUF1 (N3497, N3486);
not NOT1 (N3498, N3488);
or OR3 (N3499, N3493, N126, N1561);
or OR4 (N3500, N3485, N2226, N1213, N3037);
and AND3 (N3501, N3489, N2936, N673);
nand NAND3 (N3502, N3492, N1338, N2457);
buf BUF1 (N3503, N3491);
and AND2 (N3504, N3502, N3102);
and AND3 (N3505, N3501, N2053, N3296);
not NOT1 (N3506, N3503);
and AND4 (N3507, N3496, N2831, N1834, N288);
xor XOR2 (N3508, N3495, N3086);
buf BUF1 (N3509, N3500);
not NOT1 (N3510, N3497);
buf BUF1 (N3511, N3504);
not NOT1 (N3512, N3498);
buf BUF1 (N3513, N3506);
buf BUF1 (N3514, N3509);
not NOT1 (N3515, N3494);
nor NOR3 (N3516, N3510, N1241, N2410);
and AND4 (N3517, N3499, N247, N2209, N2875);
xor XOR2 (N3518, N3508, N3388);
and AND3 (N3519, N3514, N2708, N1796);
nor NOR4 (N3520, N3515, N1107, N1783, N48);
nand NAND2 (N3521, N3505, N2228);
nand NAND3 (N3522, N3518, N462, N58);
buf BUF1 (N3523, N3512);
nor NOR2 (N3524, N3523, N1432);
xor XOR2 (N3525, N3521, N2384);
nor NOR4 (N3526, N3516, N3498, N2449, N1955);
not NOT1 (N3527, N3526);
nor NOR4 (N3528, N3513, N3175, N751, N2777);
buf BUF1 (N3529, N3524);
not NOT1 (N3530, N3520);
nand NAND3 (N3531, N3507, N1700, N3039);
or OR2 (N3532, N3525, N1246);
xor XOR2 (N3533, N3528, N1015);
and AND4 (N3534, N3529, N2771, N308, N1580);
xor XOR2 (N3535, N3522, N2219);
and AND4 (N3536, N3532, N2172, N234, N1632);
xor XOR2 (N3537, N3535, N148);
xor XOR2 (N3538, N3537, N2562);
xor XOR2 (N3539, N3527, N3421);
nand NAND4 (N3540, N3534, N3084, N1116, N971);
xor XOR2 (N3541, N3519, N3302);
buf BUF1 (N3542, N3517);
or OR2 (N3543, N3538, N3107);
nand NAND4 (N3544, N3542, N1431, N2334, N774);
not NOT1 (N3545, N3533);
and AND2 (N3546, N3545, N493);
xor XOR2 (N3547, N3546, N305);
or OR3 (N3548, N3541, N1681, N1820);
and AND3 (N3549, N3531, N2791, N2258);
or OR3 (N3550, N3539, N1977, N863);
not NOT1 (N3551, N3511);
not NOT1 (N3552, N3530);
nor NOR4 (N3553, N3552, N2060, N3552, N2861);
not NOT1 (N3554, N3536);
xor XOR2 (N3555, N3553, N2147);
xor XOR2 (N3556, N3548, N2553);
xor XOR2 (N3557, N3550, N2690);
not NOT1 (N3558, N3557);
xor XOR2 (N3559, N3556, N3480);
or OR2 (N3560, N3555, N891);
and AND3 (N3561, N3547, N636, N3064);
buf BUF1 (N3562, N3551);
xor XOR2 (N3563, N3554, N799);
xor XOR2 (N3564, N3561, N2826);
nand NAND3 (N3565, N3564, N1913, N533);
not NOT1 (N3566, N3563);
or OR3 (N3567, N3544, N1886, N890);
xor XOR2 (N3568, N3543, N970);
buf BUF1 (N3569, N3562);
nor NOR2 (N3570, N3558, N1430);
or OR4 (N3571, N3560, N356, N2267, N1577);
or OR2 (N3572, N3565, N3321);
xor XOR2 (N3573, N3566, N3306);
or OR4 (N3574, N3573, N227, N3304, N3147);
buf BUF1 (N3575, N3559);
nand NAND2 (N3576, N3571, N12);
buf BUF1 (N3577, N3569);
buf BUF1 (N3578, N3567);
and AND2 (N3579, N3575, N1985);
xor XOR2 (N3580, N3572, N2230);
or OR3 (N3581, N3576, N2547, N2635);
nor NOR3 (N3582, N3540, N2495, N346);
not NOT1 (N3583, N3581);
not NOT1 (N3584, N3574);
nand NAND4 (N3585, N3583, N49, N667, N2379);
nor NOR4 (N3586, N3549, N672, N797, N3521);
buf BUF1 (N3587, N3570);
nor NOR3 (N3588, N3586, N3252, N2647);
and AND2 (N3589, N3577, N1818);
nor NOR3 (N3590, N3584, N400, N2114);
and AND3 (N3591, N3589, N685, N419);
xor XOR2 (N3592, N3590, N3054);
or OR2 (N3593, N3585, N544);
and AND4 (N3594, N3578, N2315, N1371, N41);
buf BUF1 (N3595, N3580);
or OR2 (N3596, N3591, N3333);
or OR3 (N3597, N3588, N1673, N42);
and AND2 (N3598, N3593, N731);
nor NOR4 (N3599, N3587, N733, N2524, N2446);
buf BUF1 (N3600, N3597);
nand NAND2 (N3601, N3599, N2858);
not NOT1 (N3602, N3582);
nand NAND3 (N3603, N3594, N3065, N540);
nand NAND4 (N3604, N3568, N1316, N3406, N1099);
not NOT1 (N3605, N3598);
buf BUF1 (N3606, N3596);
and AND3 (N3607, N3595, N533, N1426);
not NOT1 (N3608, N3600);
xor XOR2 (N3609, N3606, N3009);
nand NAND3 (N3610, N3609, N1337, N3163);
not NOT1 (N3611, N3607);
and AND3 (N3612, N3603, N2916, N3445);
not NOT1 (N3613, N3602);
nand NAND2 (N3614, N3608, N81);
nor NOR4 (N3615, N3579, N1493, N1657, N201);
buf BUF1 (N3616, N3615);
not NOT1 (N3617, N3613);
nor NOR2 (N3618, N3610, N821);
not NOT1 (N3619, N3611);
nand NAND3 (N3620, N3592, N1506, N2582);
xor XOR2 (N3621, N3605, N1172);
xor XOR2 (N3622, N3618, N3174);
buf BUF1 (N3623, N3621);
not NOT1 (N3624, N3619);
buf BUF1 (N3625, N3623);
buf BUF1 (N3626, N3620);
and AND2 (N3627, N3622, N2010);
not NOT1 (N3628, N3616);
or OR2 (N3629, N3604, N738);
and AND2 (N3630, N3601, N2022);
buf BUF1 (N3631, N3624);
and AND2 (N3632, N3627, N477);
nor NOR2 (N3633, N3628, N1723);
not NOT1 (N3634, N3631);
or OR3 (N3635, N3614, N2621, N1717);
xor XOR2 (N3636, N3612, N3609);
nand NAND3 (N3637, N3635, N2249, N3440);
nor NOR3 (N3638, N3633, N697, N2708);
nor NOR3 (N3639, N3637, N2040, N1498);
and AND4 (N3640, N3636, N393, N1278, N632);
and AND3 (N3641, N3629, N172, N79);
or OR2 (N3642, N3634, N155);
nand NAND2 (N3643, N3638, N567);
or OR2 (N3644, N3625, N3416);
or OR4 (N3645, N3644, N3410, N713, N1267);
nand NAND4 (N3646, N3617, N2738, N701, N3641);
and AND2 (N3647, N2523, N229);
nand NAND3 (N3648, N3647, N2073, N700);
and AND4 (N3649, N3642, N2800, N104, N3190);
xor XOR2 (N3650, N3639, N2290);
nand NAND4 (N3651, N3626, N2378, N978, N1019);
not NOT1 (N3652, N3645);
or OR4 (N3653, N3646, N2180, N3187, N229);
not NOT1 (N3654, N3640);
not NOT1 (N3655, N3643);
and AND3 (N3656, N3652, N24, N1559);
not NOT1 (N3657, N3630);
nor NOR2 (N3658, N3653, N3572);
and AND2 (N3659, N3655, N3394);
buf BUF1 (N3660, N3654);
nor NOR2 (N3661, N3648, N566);
buf BUF1 (N3662, N3656);
buf BUF1 (N3663, N3657);
not NOT1 (N3664, N3659);
not NOT1 (N3665, N3663);
not NOT1 (N3666, N3662);
xor XOR2 (N3667, N3658, N937);
and AND2 (N3668, N3651, N1437);
nor NOR4 (N3669, N3665, N2417, N2908, N1434);
buf BUF1 (N3670, N3667);
nor NOR4 (N3671, N3632, N1114, N2535, N36);
nand NAND3 (N3672, N3671, N1646, N3197);
and AND2 (N3673, N3670, N1479);
nand NAND4 (N3674, N3649, N1283, N2803, N3476);
nor NOR2 (N3675, N3660, N1648);
xor XOR2 (N3676, N3675, N1491);
buf BUF1 (N3677, N3668);
nor NOR4 (N3678, N3666, N1455, N991, N2638);
or OR2 (N3679, N3664, N751);
or OR3 (N3680, N3650, N273, N2486);
buf BUF1 (N3681, N3673);
or OR3 (N3682, N3677, N3243, N2539);
nor NOR2 (N3683, N3680, N237);
and AND3 (N3684, N3674, N2059, N107);
and AND2 (N3685, N3672, N580);
not NOT1 (N3686, N3681);
buf BUF1 (N3687, N3676);
buf BUF1 (N3688, N3661);
xor XOR2 (N3689, N3688, N1542);
buf BUF1 (N3690, N3686);
nand NAND2 (N3691, N3679, N805);
buf BUF1 (N3692, N3691);
and AND4 (N3693, N3690, N965, N1503, N2267);
buf BUF1 (N3694, N3685);
nor NOR4 (N3695, N3684, N3451, N3684, N3608);
not NOT1 (N3696, N3695);
not NOT1 (N3697, N3693);
xor XOR2 (N3698, N3696, N762);
and AND4 (N3699, N3692, N1886, N1889, N605);
nor NOR4 (N3700, N3697, N1803, N3450, N2368);
and AND2 (N3701, N3689, N1159);
or OR2 (N3702, N3699, N2762);
xor XOR2 (N3703, N3683, N258);
nand NAND3 (N3704, N3682, N1540, N3114);
xor XOR2 (N3705, N3702, N2555);
nand NAND2 (N3706, N3705, N2525);
nor NOR4 (N3707, N3706, N608, N112, N13);
xor XOR2 (N3708, N3669, N2308);
nand NAND3 (N3709, N3678, N2161, N703);
xor XOR2 (N3710, N3707, N3231);
not NOT1 (N3711, N3687);
buf BUF1 (N3712, N3710);
and AND4 (N3713, N3712, N2100, N2277, N2004);
xor XOR2 (N3714, N3713, N75);
nor NOR4 (N3715, N3700, N2941, N3545, N1134);
xor XOR2 (N3716, N3704, N1115);
xor XOR2 (N3717, N3714, N2033);
nor NOR3 (N3718, N3709, N2152, N2894);
or OR3 (N3719, N3703, N2579, N1645);
nor NOR4 (N3720, N3719, N1599, N2117, N3015);
and AND3 (N3721, N3708, N3283, N2954);
not NOT1 (N3722, N3720);
nand NAND4 (N3723, N3717, N1047, N3434, N1377);
nor NOR3 (N3724, N3723, N311, N2752);
buf BUF1 (N3725, N3715);
not NOT1 (N3726, N3721);
buf BUF1 (N3727, N3698);
and AND3 (N3728, N3701, N2886, N1450);
nor NOR4 (N3729, N3725, N1165, N1345, N1428);
and AND2 (N3730, N3718, N2642);
xor XOR2 (N3731, N3694, N2415);
not NOT1 (N3732, N3716);
buf BUF1 (N3733, N3726);
and AND3 (N3734, N3733, N2920, N2301);
nor NOR4 (N3735, N3724, N2294, N788, N739);
and AND4 (N3736, N3731, N3321, N3117, N83);
and AND4 (N3737, N3727, N1455, N2017, N1744);
not NOT1 (N3738, N3722);
nand NAND4 (N3739, N3732, N1355, N1571, N2044);
not NOT1 (N3740, N3729);
nand NAND4 (N3741, N3728, N3629, N291, N891);
nor NOR3 (N3742, N3739, N59, N390);
or OR2 (N3743, N3734, N3704);
and AND3 (N3744, N3742, N1810, N1540);
nor NOR4 (N3745, N3741, N1705, N1386, N2035);
not NOT1 (N3746, N3711);
xor XOR2 (N3747, N3735, N1729);
and AND4 (N3748, N3747, N2986, N3676, N1943);
xor XOR2 (N3749, N3730, N3362);
nor NOR2 (N3750, N3748, N2336);
xor XOR2 (N3751, N3746, N3164);
not NOT1 (N3752, N3738);
and AND3 (N3753, N3745, N1354, N2261);
xor XOR2 (N3754, N3744, N3143);
xor XOR2 (N3755, N3753, N810);
xor XOR2 (N3756, N3754, N2058);
buf BUF1 (N3757, N3752);
or OR3 (N3758, N3743, N1043, N301);
nor NOR2 (N3759, N3737, N1599);
not NOT1 (N3760, N3736);
nor NOR4 (N3761, N3758, N2660, N2000, N1288);
and AND3 (N3762, N3750, N2258, N2090);
nand NAND3 (N3763, N3762, N3165, N260);
nand NAND2 (N3764, N3763, N3138);
nor NOR4 (N3765, N3760, N2726, N3462, N3206);
xor XOR2 (N3766, N3751, N457);
buf BUF1 (N3767, N3757);
xor XOR2 (N3768, N3759, N1777);
nand NAND3 (N3769, N3749, N990, N1536);
not NOT1 (N3770, N3769);
and AND3 (N3771, N3770, N1891, N2200);
and AND3 (N3772, N3761, N1614, N94);
xor XOR2 (N3773, N3756, N3277);
xor XOR2 (N3774, N3767, N2590);
or OR2 (N3775, N3764, N2827);
buf BUF1 (N3776, N3771);
buf BUF1 (N3777, N3765);
nand NAND2 (N3778, N3740, N1549);
buf BUF1 (N3779, N3775);
nor NOR2 (N3780, N3755, N2651);
xor XOR2 (N3781, N3780, N2095);
or OR3 (N3782, N3773, N441, N536);
not NOT1 (N3783, N3768);
nand NAND2 (N3784, N3783, N3129);
nand NAND4 (N3785, N3782, N312, N1367, N3368);
or OR3 (N3786, N3781, N2002, N2390);
or OR2 (N3787, N3772, N2337);
and AND3 (N3788, N3776, N1274, N435);
and AND2 (N3789, N3784, N1268);
nor NOR4 (N3790, N3785, N3299, N937, N3248);
not NOT1 (N3791, N3790);
buf BUF1 (N3792, N3787);
nor NOR4 (N3793, N3792, N3533, N346, N5);
not NOT1 (N3794, N3777);
nand NAND4 (N3795, N3791, N3392, N1543, N2653);
and AND3 (N3796, N3793, N1475, N1857);
nor NOR4 (N3797, N3795, N105, N2797, N2569);
and AND3 (N3798, N3786, N274, N729);
nand NAND3 (N3799, N3789, N3269, N3787);
not NOT1 (N3800, N3797);
xor XOR2 (N3801, N3774, N83);
buf BUF1 (N3802, N3801);
buf BUF1 (N3803, N3778);
nor NOR3 (N3804, N3794, N3662, N3);
or OR4 (N3805, N3779, N1519, N3394, N3328);
and AND4 (N3806, N3799, N3234, N2967, N3780);
xor XOR2 (N3807, N3766, N3660);
nand NAND2 (N3808, N3806, N68);
or OR4 (N3809, N3798, N3733, N2536, N47);
not NOT1 (N3810, N3807);
nor NOR3 (N3811, N3805, N73, N3233);
or OR3 (N3812, N3809, N3784, N2504);
nor NOR4 (N3813, N3800, N3414, N3020, N3221);
not NOT1 (N3814, N3804);
xor XOR2 (N3815, N3808, N2908);
and AND3 (N3816, N3810, N3012, N1390);
not NOT1 (N3817, N3788);
and AND2 (N3818, N3815, N2100);
not NOT1 (N3819, N3818);
nor NOR2 (N3820, N3816, N2159);
nand NAND4 (N3821, N3813, N2463, N2302, N1628);
or OR3 (N3822, N3819, N64, N3527);
not NOT1 (N3823, N3814);
or OR4 (N3824, N3817, N440, N1993, N83);
buf BUF1 (N3825, N3821);
or OR4 (N3826, N3823, N1797, N1277, N1289);
buf BUF1 (N3827, N3824);
xor XOR2 (N3828, N3820, N370);
not NOT1 (N3829, N3803);
nand NAND3 (N3830, N3828, N3609, N851);
or OR4 (N3831, N3796, N1674, N543, N2665);
nand NAND3 (N3832, N3827, N3604, N2454);
buf BUF1 (N3833, N3812);
and AND3 (N3834, N3831, N1548, N1557);
nor NOR4 (N3835, N3802, N1387, N3105, N1004);
buf BUF1 (N3836, N3826);
or OR3 (N3837, N3825, N1940, N2702);
nor NOR2 (N3838, N3835, N404);
and AND4 (N3839, N3832, N208, N2872, N1956);
buf BUF1 (N3840, N3838);
not NOT1 (N3841, N3822);
nor NOR3 (N3842, N3836, N3032, N3743);
and AND3 (N3843, N3839, N2698, N1614);
buf BUF1 (N3844, N3811);
nor NOR4 (N3845, N3844, N1270, N579, N2140);
buf BUF1 (N3846, N3833);
and AND4 (N3847, N3834, N736, N515, N1903);
not NOT1 (N3848, N3845);
buf BUF1 (N3849, N3830);
or OR4 (N3850, N3842, N2499, N2191, N3667);
and AND2 (N3851, N3847, N1249);
not NOT1 (N3852, N3840);
or OR3 (N3853, N3841, N3424, N1236);
nor NOR3 (N3854, N3849, N3196, N2046);
and AND4 (N3855, N3850, N2579, N1978, N3091);
or OR2 (N3856, N3848, N3262);
and AND2 (N3857, N3851, N2262);
buf BUF1 (N3858, N3846);
not NOT1 (N3859, N3853);
or OR4 (N3860, N3829, N1457, N1198, N297);
buf BUF1 (N3861, N3858);
xor XOR2 (N3862, N3859, N1093);
buf BUF1 (N3863, N3856);
nand NAND4 (N3864, N3855, N2579, N3675, N88);
nor NOR2 (N3865, N3862, N134);
and AND4 (N3866, N3865, N1116, N2377, N1589);
nor NOR2 (N3867, N3864, N426);
buf BUF1 (N3868, N3861);
nor NOR2 (N3869, N3837, N1902);
buf BUF1 (N3870, N3868);
and AND3 (N3871, N3869, N1472, N1404);
not NOT1 (N3872, N3860);
nand NAND3 (N3873, N3857, N775, N1196);
buf BUF1 (N3874, N3873);
not NOT1 (N3875, N3874);
buf BUF1 (N3876, N3854);
buf BUF1 (N3877, N3863);
buf BUF1 (N3878, N3867);
or OR3 (N3879, N3872, N1694, N2078);
not NOT1 (N3880, N3876);
buf BUF1 (N3881, N3871);
buf BUF1 (N3882, N3875);
not NOT1 (N3883, N3843);
and AND4 (N3884, N3882, N2263, N951, N2838);
not NOT1 (N3885, N3852);
buf BUF1 (N3886, N3881);
or OR2 (N3887, N3878, N2307);
and AND3 (N3888, N3879, N1288, N3196);
and AND2 (N3889, N3880, N2332);
xor XOR2 (N3890, N3888, N2805);
nor NOR2 (N3891, N3889, N667);
buf BUF1 (N3892, N3891);
and AND2 (N3893, N3890, N1699);
and AND3 (N3894, N3866, N1344, N193);
nor NOR4 (N3895, N3892, N300, N1766, N1016);
or OR3 (N3896, N3870, N2849, N871);
or OR2 (N3897, N3895, N2213);
or OR2 (N3898, N3884, N2677);
nand NAND2 (N3899, N3898, N2267);
and AND2 (N3900, N3877, N3564);
buf BUF1 (N3901, N3883);
not NOT1 (N3902, N3886);
not NOT1 (N3903, N3897);
nor NOR4 (N3904, N3901, N178, N637, N959);
or OR4 (N3905, N3893, N2898, N1665, N2613);
and AND4 (N3906, N3900, N230, N1153, N1265);
not NOT1 (N3907, N3894);
xor XOR2 (N3908, N3906, N2779);
nand NAND4 (N3909, N3896, N40, N1557, N1878);
and AND4 (N3910, N3905, N3152, N95, N2318);
buf BUF1 (N3911, N3908);
not NOT1 (N3912, N3902);
and AND2 (N3913, N3909, N1213);
nor NOR4 (N3914, N3899, N3056, N2539, N3098);
or OR4 (N3915, N3903, N328, N144, N421);
buf BUF1 (N3916, N3915);
buf BUF1 (N3917, N3887);
or OR2 (N3918, N3916, N717);
and AND4 (N3919, N3911, N65, N220, N3542);
or OR4 (N3920, N3914, N55, N2577, N1926);
buf BUF1 (N3921, N3910);
and AND3 (N3922, N3913, N3862, N3100);
xor XOR2 (N3923, N3919, N502);
not NOT1 (N3924, N3912);
and AND2 (N3925, N3907, N302);
buf BUF1 (N3926, N3925);
buf BUF1 (N3927, N3920);
nor NOR4 (N3928, N3885, N2498, N1864, N3827);
not NOT1 (N3929, N3926);
or OR4 (N3930, N3927, N1351, N3429, N3048);
nand NAND2 (N3931, N3928, N2934);
and AND4 (N3932, N3930, N880, N2346, N3698);
and AND3 (N3933, N3921, N1347, N917);
xor XOR2 (N3934, N3917, N1954);
not NOT1 (N3935, N3933);
and AND2 (N3936, N3935, N2265);
buf BUF1 (N3937, N3923);
nor NOR3 (N3938, N3918, N2436, N2468);
nand NAND4 (N3939, N3922, N2438, N2157, N2202);
and AND4 (N3940, N3931, N1969, N2847, N2817);
buf BUF1 (N3941, N3929);
or OR3 (N3942, N3938, N3206, N3689);
buf BUF1 (N3943, N3904);
xor XOR2 (N3944, N3942, N2099);
and AND2 (N3945, N3937, N220);
or OR2 (N3946, N3932, N389);
or OR4 (N3947, N3946, N1603, N1214, N3600);
xor XOR2 (N3948, N3944, N732);
or OR2 (N3949, N3943, N349);
not NOT1 (N3950, N3945);
not NOT1 (N3951, N3941);
nand NAND3 (N3952, N3951, N1927, N3657);
buf BUF1 (N3953, N3949);
nor NOR4 (N3954, N3940, N238, N3377, N3064);
xor XOR2 (N3955, N3948, N3804);
and AND4 (N3956, N3934, N1351, N2341, N2342);
buf BUF1 (N3957, N3936);
nor NOR3 (N3958, N3955, N276, N3083);
not NOT1 (N3959, N3954);
not NOT1 (N3960, N3959);
nor NOR2 (N3961, N3956, N235);
and AND2 (N3962, N3961, N650);
not NOT1 (N3963, N3939);
xor XOR2 (N3964, N3962, N461);
not NOT1 (N3965, N3952);
buf BUF1 (N3966, N3960);
and AND3 (N3967, N3947, N3262, N134);
nand NAND4 (N3968, N3958, N2723, N2839, N3915);
nor NOR3 (N3969, N3950, N2577, N2660);
nor NOR4 (N3970, N3966, N1622, N2579, N1745);
not NOT1 (N3971, N3965);
or OR3 (N3972, N3953, N573, N1831);
nor NOR4 (N3973, N3924, N624, N697, N1969);
nand NAND3 (N3974, N3967, N2665, N982);
nor NOR3 (N3975, N3964, N82, N400);
or OR2 (N3976, N3968, N1101);
not NOT1 (N3977, N3974);
or OR2 (N3978, N3975, N2779);
nand NAND3 (N3979, N3976, N595, N1895);
nand NAND4 (N3980, N3979, N1855, N1909, N3226);
buf BUF1 (N3981, N3980);
not NOT1 (N3982, N3978);
and AND2 (N3983, N3971, N3658);
or OR3 (N3984, N3970, N2449, N3138);
and AND3 (N3985, N3969, N806, N2928);
not NOT1 (N3986, N3983);
buf BUF1 (N3987, N3972);
nand NAND3 (N3988, N3982, N1181, N1669);
nand NAND3 (N3989, N3957, N1272, N50);
nand NAND4 (N3990, N3973, N2440, N867, N2073);
buf BUF1 (N3991, N3981);
not NOT1 (N3992, N3989);
nor NOR4 (N3993, N3977, N2392, N2996, N566);
nor NOR3 (N3994, N3985, N3914, N3208);
buf BUF1 (N3995, N3992);
not NOT1 (N3996, N3994);
xor XOR2 (N3997, N3984, N1076);
buf BUF1 (N3998, N3988);
and AND2 (N3999, N3987, N271);
nor NOR4 (N4000, N3990, N2537, N2854, N201);
nor NOR4 (N4001, N3999, N853, N3219, N492);
nand NAND3 (N4002, N3998, N1042, N178);
buf BUF1 (N4003, N3996);
nor NOR2 (N4004, N3986, N2448);
nand NAND4 (N4005, N3997, N3269, N347, N885);
xor XOR2 (N4006, N3995, N2358);
buf BUF1 (N4007, N4005);
nand NAND3 (N4008, N4006, N2634, N2024);
not NOT1 (N4009, N4004);
or OR4 (N4010, N3991, N2297, N208, N1284);
nand NAND3 (N4011, N4001, N2410, N783);
and AND3 (N4012, N4008, N617, N2671);
nor NOR2 (N4013, N4000, N1494);
not NOT1 (N4014, N4010);
or OR4 (N4015, N4003, N2735, N3656, N3624);
and AND3 (N4016, N4012, N2907, N808);
nor NOR2 (N4017, N4007, N377);
not NOT1 (N4018, N4011);
nand NAND3 (N4019, N3993, N3322, N3702);
nor NOR4 (N4020, N4018, N2472, N1499, N1424);
nor NOR2 (N4021, N4013, N1325);
nand NAND3 (N4022, N4014, N1185, N2459);
nor NOR2 (N4023, N4020, N319);
xor XOR2 (N4024, N3963, N1974);
or OR3 (N4025, N4021, N704, N2790);
nand NAND4 (N4026, N4015, N86, N3720, N595);
not NOT1 (N4027, N4016);
not NOT1 (N4028, N4002);
nand NAND3 (N4029, N4026, N2647, N2848);
or OR4 (N4030, N4023, N1967, N2788, N2451);
and AND2 (N4031, N4017, N3492);
and AND3 (N4032, N4024, N109, N1303);
nand NAND2 (N4033, N4030, N3739);
xor XOR2 (N4034, N4025, N2767);
xor XOR2 (N4035, N4033, N1925);
nor NOR3 (N4036, N4022, N3313, N3110);
nor NOR3 (N4037, N4034, N709, N1634);
xor XOR2 (N4038, N4036, N1949);
and AND2 (N4039, N4019, N192);
nand NAND2 (N4040, N4039, N3050);
not NOT1 (N4041, N4031);
and AND3 (N4042, N4029, N692, N2017);
and AND4 (N4043, N4035, N3686, N464, N1475);
buf BUF1 (N4044, N4038);
not NOT1 (N4045, N4041);
and AND4 (N4046, N4028, N3807, N123, N2647);
xor XOR2 (N4047, N4032, N1875);
not NOT1 (N4048, N4009);
or OR2 (N4049, N4043, N1601);
or OR4 (N4050, N4027, N592, N936, N2018);
and AND3 (N4051, N4045, N2880, N2017);
not NOT1 (N4052, N4048);
or OR2 (N4053, N4051, N1483);
nand NAND3 (N4054, N4052, N2237, N2870);
and AND2 (N4055, N4040, N2977);
nand NAND4 (N4056, N4047, N1680, N219, N741);
buf BUF1 (N4057, N4037);
xor XOR2 (N4058, N4042, N375);
and AND3 (N4059, N4055, N3916, N2516);
or OR4 (N4060, N4049, N1728, N3794, N2672);
and AND4 (N4061, N4059, N1386, N1641, N179);
nand NAND3 (N4062, N4053, N1369, N1617);
nor NOR2 (N4063, N4058, N3947);
nand NAND2 (N4064, N4057, N422);
buf BUF1 (N4065, N4064);
not NOT1 (N4066, N4062);
xor XOR2 (N4067, N4056, N2271);
nand NAND3 (N4068, N4067, N3922, N2465);
xor XOR2 (N4069, N4063, N2455);
nand NAND3 (N4070, N4066, N1174, N1493);
buf BUF1 (N4071, N4054);
buf BUF1 (N4072, N4070);
nand NAND2 (N4073, N4072, N3240);
and AND4 (N4074, N4050, N1936, N1951, N1641);
nor NOR4 (N4075, N4068, N2310, N1376, N1626);
nand NAND2 (N4076, N4075, N3124);
not NOT1 (N4077, N4073);
nor NOR3 (N4078, N4046, N1751, N3427);
and AND3 (N4079, N4061, N339, N2315);
xor XOR2 (N4080, N4077, N3837);
and AND2 (N4081, N4076, N3577);
or OR3 (N4082, N4044, N2246, N2217);
not NOT1 (N4083, N4080);
not NOT1 (N4084, N4069);
not NOT1 (N4085, N4065);
xor XOR2 (N4086, N4085, N1558);
xor XOR2 (N4087, N4086, N694);
nand NAND2 (N4088, N4060, N2203);
nor NOR4 (N4089, N4084, N2494, N2044, N2873);
nor NOR4 (N4090, N4082, N3975, N744, N3334);
xor XOR2 (N4091, N4079, N3121);
nor NOR2 (N4092, N4087, N3847);
or OR4 (N4093, N4092, N3520, N1539, N2806);
nand NAND4 (N4094, N4088, N1804, N1918, N2969);
and AND2 (N4095, N4071, N3487);
not NOT1 (N4096, N4089);
not NOT1 (N4097, N4074);
nor NOR3 (N4098, N4096, N1001, N3248);
nand NAND2 (N4099, N4090, N1047);
and AND3 (N4100, N4093, N2106, N2394);
or OR3 (N4101, N4094, N3607, N3523);
buf BUF1 (N4102, N4091);
nand NAND3 (N4103, N4100, N771, N4019);
xor XOR2 (N4104, N4081, N1239);
xor XOR2 (N4105, N4102, N2150);
xor XOR2 (N4106, N4098, N85);
or OR2 (N4107, N4099, N3636);
nand NAND3 (N4108, N4095, N2596, N2026);
nor NOR4 (N4109, N4101, N3367, N3248, N1237);
buf BUF1 (N4110, N4107);
nor NOR3 (N4111, N4108, N1442, N148);
buf BUF1 (N4112, N4110);
and AND2 (N4113, N4109, N3721);
buf BUF1 (N4114, N4106);
nor NOR4 (N4115, N4083, N2453, N199, N3981);
xor XOR2 (N4116, N4115, N489);
nand NAND3 (N4117, N4104, N1369, N2118);
nand NAND4 (N4118, N4113, N1899, N1017, N1847);
buf BUF1 (N4119, N4103);
buf BUF1 (N4120, N4119);
or OR2 (N4121, N4105, N2181);
nand NAND3 (N4122, N4111, N1887, N2877);
nand NAND3 (N4123, N4118, N2863, N1784);
nand NAND2 (N4124, N4097, N3751);
xor XOR2 (N4125, N4123, N3699);
nand NAND2 (N4126, N4078, N2495);
xor XOR2 (N4127, N4117, N2042);
nor NOR3 (N4128, N4112, N188, N3639);
and AND2 (N4129, N4124, N1319);
buf BUF1 (N4130, N4114);
nand NAND4 (N4131, N4128, N533, N324, N343);
and AND2 (N4132, N4121, N2526);
nor NOR2 (N4133, N4129, N228);
xor XOR2 (N4134, N4132, N2995);
not NOT1 (N4135, N4126);
xor XOR2 (N4136, N4130, N3683);
not NOT1 (N4137, N4125);
not NOT1 (N4138, N4136);
not NOT1 (N4139, N4120);
nand NAND2 (N4140, N4131, N610);
and AND4 (N4141, N4138, N1537, N2784, N2800);
nor NOR3 (N4142, N4134, N3838, N3338);
buf BUF1 (N4143, N4133);
and AND3 (N4144, N4141, N708, N169);
or OR4 (N4145, N4142, N1064, N3109, N2348);
and AND3 (N4146, N4135, N1391, N3866);
nand NAND2 (N4147, N4139, N804);
buf BUF1 (N4148, N4122);
buf BUF1 (N4149, N4137);
and AND2 (N4150, N4116, N131);
and AND4 (N4151, N4127, N2396, N3748, N3820);
or OR2 (N4152, N4146, N1385);
and AND2 (N4153, N4145, N745);
and AND2 (N4154, N4149, N238);
xor XOR2 (N4155, N4148, N1945);
or OR4 (N4156, N4147, N1925, N3847, N1653);
or OR3 (N4157, N4156, N1909, N734);
nand NAND4 (N4158, N4150, N2357, N520, N1113);
nor NOR4 (N4159, N4158, N2819, N1881, N3079);
nand NAND3 (N4160, N4153, N3379, N3319);
and AND4 (N4161, N4152, N1676, N970, N3125);
nor NOR3 (N4162, N4140, N161, N665);
buf BUF1 (N4163, N4160);
buf BUF1 (N4164, N4154);
buf BUF1 (N4165, N4155);
nand NAND3 (N4166, N4163, N808, N1336);
nand NAND3 (N4167, N4164, N1397, N465);
and AND2 (N4168, N4159, N1632);
nor NOR3 (N4169, N4166, N1202, N2687);
or OR4 (N4170, N4143, N1782, N3389, N437);
or OR2 (N4171, N4144, N17);
or OR4 (N4172, N4151, N3591, N3663, N1943);
xor XOR2 (N4173, N4157, N3579);
buf BUF1 (N4174, N4162);
not NOT1 (N4175, N4170);
not NOT1 (N4176, N4168);
nand NAND4 (N4177, N4167, N1433, N691, N434);
or OR2 (N4178, N4171, N644);
not NOT1 (N4179, N4161);
buf BUF1 (N4180, N4177);
or OR3 (N4181, N4176, N2524, N4110);
not NOT1 (N4182, N4175);
and AND4 (N4183, N4174, N2991, N3982, N2927);
nor NOR4 (N4184, N4181, N3438, N77, N3349);
nor NOR2 (N4185, N4182, N3688);
nor NOR2 (N4186, N4172, N1321);
nor NOR4 (N4187, N4178, N118, N2379, N2525);
or OR3 (N4188, N4185, N2682, N292);
xor XOR2 (N4189, N4183, N2242);
buf BUF1 (N4190, N4187);
or OR3 (N4191, N4190, N379, N3664);
nor NOR4 (N4192, N4188, N986, N1279, N2291);
nor NOR3 (N4193, N4169, N745, N1348);
buf BUF1 (N4194, N4173);
and AND4 (N4195, N4191, N1740, N660, N3659);
xor XOR2 (N4196, N4179, N3722);
xor XOR2 (N4197, N4186, N1141);
buf BUF1 (N4198, N4180);
xor XOR2 (N4199, N4184, N1272);
and AND4 (N4200, N4193, N278, N1937, N3351);
nand NAND4 (N4201, N4196, N2097, N4147, N89);
not NOT1 (N4202, N4192);
nor NOR4 (N4203, N4165, N2697, N1880, N4035);
nor NOR2 (N4204, N4195, N1639);
nor NOR2 (N4205, N4202, N869);
nor NOR2 (N4206, N4197, N3937);
buf BUF1 (N4207, N4205);
or OR2 (N4208, N4203, N3872);
not NOT1 (N4209, N4208);
buf BUF1 (N4210, N4209);
buf BUF1 (N4211, N4194);
buf BUF1 (N4212, N4204);
buf BUF1 (N4213, N4198);
or OR3 (N4214, N4189, N3197, N843);
nor NOR2 (N4215, N4206, N1064);
or OR2 (N4216, N4210, N2691);
and AND3 (N4217, N4207, N455, N639);
or OR3 (N4218, N4214, N717, N294);
or OR2 (N4219, N4199, N781);
not NOT1 (N4220, N4217);
xor XOR2 (N4221, N4213, N259);
nand NAND4 (N4222, N4215, N1726, N1519, N1640);
xor XOR2 (N4223, N4201, N1520);
buf BUF1 (N4224, N4221);
and AND2 (N4225, N4212, N710);
and AND3 (N4226, N4223, N1640, N1157);
nand NAND3 (N4227, N4224, N633, N3251);
or OR2 (N4228, N4211, N3133);
and AND3 (N4229, N4218, N2141, N211);
buf BUF1 (N4230, N4226);
not NOT1 (N4231, N4225);
buf BUF1 (N4232, N4216);
xor XOR2 (N4233, N4230, N1509);
and AND2 (N4234, N4219, N1866);
or OR2 (N4235, N4229, N550);
xor XOR2 (N4236, N4232, N1837);
buf BUF1 (N4237, N4233);
or OR3 (N4238, N4220, N1623, N1805);
not NOT1 (N4239, N4231);
or OR3 (N4240, N4227, N32, N3820);
buf BUF1 (N4241, N4239);
buf BUF1 (N4242, N4240);
not NOT1 (N4243, N4235);
nand NAND4 (N4244, N4238, N2881, N2045, N1930);
not NOT1 (N4245, N4228);
nor NOR2 (N4246, N4245, N390);
buf BUF1 (N4247, N4241);
not NOT1 (N4248, N4236);
and AND2 (N4249, N4242, N1178);
and AND2 (N4250, N4247, N2309);
nand NAND3 (N4251, N4234, N109, N2224);
or OR2 (N4252, N4222, N3754);
not NOT1 (N4253, N4237);
or OR4 (N4254, N4248, N327, N1441, N4052);
buf BUF1 (N4255, N4251);
nand NAND2 (N4256, N4255, N4250);
xor XOR2 (N4257, N229, N828);
and AND4 (N4258, N4246, N2943, N1999, N3224);
or OR4 (N4259, N4254, N1590, N1993, N1367);
nor NOR2 (N4260, N4257, N3291);
xor XOR2 (N4261, N4259, N3395);
or OR3 (N4262, N4258, N1198, N3091);
and AND2 (N4263, N4262, N2178);
buf BUF1 (N4264, N4261);
buf BUF1 (N4265, N4200);
nor NOR4 (N4266, N4260, N2662, N4090, N3300);
buf BUF1 (N4267, N4265);
buf BUF1 (N4268, N4249);
xor XOR2 (N4269, N4264, N1624);
xor XOR2 (N4270, N4267, N169);
nor NOR3 (N4271, N4269, N2595, N2529);
not NOT1 (N4272, N4243);
and AND2 (N4273, N4272, N3996);
nand NAND2 (N4274, N4244, N612);
nor NOR2 (N4275, N4263, N1685);
xor XOR2 (N4276, N4253, N4049);
or OR3 (N4277, N4256, N1013, N3100);
xor XOR2 (N4278, N4268, N3);
nand NAND4 (N4279, N4274, N880, N1243, N2269);
nor NOR4 (N4280, N4278, N2957, N1292, N3917);
buf BUF1 (N4281, N4266);
nand NAND4 (N4282, N4276, N2276, N3327, N4217);
nand NAND4 (N4283, N4270, N2141, N56, N3358);
nor NOR2 (N4284, N4279, N2037);
not NOT1 (N4285, N4281);
buf BUF1 (N4286, N4285);
not NOT1 (N4287, N4252);
or OR3 (N4288, N4287, N3489, N1754);
nand NAND3 (N4289, N4284, N2888, N2781);
and AND4 (N4290, N4282, N2861, N2332, N3127);
buf BUF1 (N4291, N4273);
nand NAND4 (N4292, N4275, N2651, N3746, N58);
or OR4 (N4293, N4277, N186, N1820, N2086);
xor XOR2 (N4294, N4291, N579);
not NOT1 (N4295, N4280);
xor XOR2 (N4296, N4271, N4184);
not NOT1 (N4297, N4292);
nand NAND2 (N4298, N4294, N2645);
or OR4 (N4299, N4295, N3232, N4055, N1041);
buf BUF1 (N4300, N4286);
xor XOR2 (N4301, N4298, N590);
buf BUF1 (N4302, N4293);
buf BUF1 (N4303, N4300);
and AND2 (N4304, N4289, N340);
xor XOR2 (N4305, N4301, N3826);
or OR4 (N4306, N4305, N784, N3658, N490);
nor NOR3 (N4307, N4306, N3443, N1443);
nand NAND2 (N4308, N4302, N1624);
and AND4 (N4309, N4299, N745, N694, N3155);
or OR2 (N4310, N4307, N2048);
buf BUF1 (N4311, N4309);
xor XOR2 (N4312, N4304, N3417);
or OR3 (N4313, N4312, N8, N3345);
and AND2 (N4314, N4311, N3012);
nor NOR2 (N4315, N4310, N2172);
and AND4 (N4316, N4314, N2393, N2856, N2436);
xor XOR2 (N4317, N4290, N1515);
buf BUF1 (N4318, N4317);
buf BUF1 (N4319, N4303);
or OR2 (N4320, N4288, N3485);
xor XOR2 (N4321, N4297, N113);
nor NOR3 (N4322, N4296, N3825, N3708);
not NOT1 (N4323, N4315);
nand NAND4 (N4324, N4318, N2894, N4121, N760);
nand NAND3 (N4325, N4323, N2314, N2085);
buf BUF1 (N4326, N4283);
and AND4 (N4327, N4308, N1016, N134, N2159);
xor XOR2 (N4328, N4320, N3190);
and AND4 (N4329, N4325, N506, N3532, N4267);
nand NAND2 (N4330, N4326, N3028);
and AND2 (N4331, N4327, N1056);
nor NOR2 (N4332, N4313, N3870);
xor XOR2 (N4333, N4316, N2376);
and AND3 (N4334, N4333, N769, N3239);
nand NAND3 (N4335, N4328, N4303, N3538);
or OR3 (N4336, N4330, N4219, N925);
buf BUF1 (N4337, N4332);
nor NOR3 (N4338, N4337, N3070, N2344);
not NOT1 (N4339, N4329);
nand NAND2 (N4340, N4321, N3855);
or OR3 (N4341, N4335, N4212, N1942);
xor XOR2 (N4342, N4322, N1190);
not NOT1 (N4343, N4331);
not NOT1 (N4344, N4339);
or OR3 (N4345, N4340, N2622, N10);
nand NAND2 (N4346, N4344, N1379);
and AND4 (N4347, N4324, N3342, N1144, N3134);
xor XOR2 (N4348, N4342, N2680);
nand NAND3 (N4349, N4348, N1109, N893);
xor XOR2 (N4350, N4349, N3725);
and AND2 (N4351, N4334, N1976);
nand NAND3 (N4352, N4319, N999, N2359);
nor NOR2 (N4353, N4338, N4011);
xor XOR2 (N4354, N4336, N3159);
nor NOR3 (N4355, N4352, N434, N1262);
nor NOR2 (N4356, N4351, N2734);
nor NOR4 (N4357, N4347, N2799, N3341, N266);
and AND3 (N4358, N4341, N116, N3182);
nand NAND3 (N4359, N4346, N1826, N3958);
not NOT1 (N4360, N4357);
and AND2 (N4361, N4359, N2642);
not NOT1 (N4362, N4350);
xor XOR2 (N4363, N4355, N373);
nor NOR3 (N4364, N4356, N3578, N628);
not NOT1 (N4365, N4358);
nor NOR2 (N4366, N4354, N53);
or OR2 (N4367, N4364, N1372);
buf BUF1 (N4368, N4367);
and AND4 (N4369, N4362, N3212, N2969, N1463);
and AND4 (N4370, N4363, N2094, N3223, N3615);
xor XOR2 (N4371, N4353, N1585);
buf BUF1 (N4372, N4360);
nand NAND4 (N4373, N4343, N2339, N412, N3932);
nor NOR4 (N4374, N4372, N2175, N1969, N1427);
nand NAND4 (N4375, N4366, N4226, N421, N3194);
buf BUF1 (N4376, N4373);
buf BUF1 (N4377, N4370);
xor XOR2 (N4378, N4377, N3041);
nor NOR3 (N4379, N4374, N2682, N2321);
not NOT1 (N4380, N4376);
or OR3 (N4381, N4378, N3228, N3436);
nand NAND3 (N4382, N4371, N3830, N1252);
xor XOR2 (N4383, N4345, N3220);
nor NOR2 (N4384, N4382, N217);
xor XOR2 (N4385, N4381, N1689);
xor XOR2 (N4386, N4369, N1525);
xor XOR2 (N4387, N4386, N2388);
nand NAND3 (N4388, N4384, N2245, N2957);
nor NOR3 (N4389, N4361, N724, N4121);
buf BUF1 (N4390, N4388);
xor XOR2 (N4391, N4380, N1863);
xor XOR2 (N4392, N4389, N4028);
not NOT1 (N4393, N4368);
xor XOR2 (N4394, N4393, N2535);
or OR4 (N4395, N4379, N1253, N4178, N4387);
xor XOR2 (N4396, N3496, N3813);
buf BUF1 (N4397, N4375);
buf BUF1 (N4398, N4397);
nand NAND4 (N4399, N4395, N1881, N3886, N2416);
or OR2 (N4400, N4365, N3189);
or OR4 (N4401, N4385, N1068, N1521, N2289);
and AND4 (N4402, N4398, N3981, N3008, N221);
not NOT1 (N4403, N4400);
and AND3 (N4404, N4396, N1247, N253);
not NOT1 (N4405, N4404);
not NOT1 (N4406, N4401);
not NOT1 (N4407, N4402);
or OR4 (N4408, N4390, N4067, N4062, N1076);
or OR4 (N4409, N4407, N3942, N3921, N395);
and AND4 (N4410, N4408, N4073, N1746, N1540);
nor NOR3 (N4411, N4399, N3220, N2809);
buf BUF1 (N4412, N4405);
and AND2 (N4413, N4411, N2459);
nor NOR3 (N4414, N4392, N427, N2803);
and AND2 (N4415, N4406, N3966);
not NOT1 (N4416, N4403);
or OR4 (N4417, N4394, N420, N1696, N2702);
not NOT1 (N4418, N4391);
xor XOR2 (N4419, N4383, N2920);
not NOT1 (N4420, N4419);
or OR4 (N4421, N4413, N4056, N1793, N1330);
or OR4 (N4422, N4410, N1566, N1209, N3470);
buf BUF1 (N4423, N4414);
or OR3 (N4424, N4409, N2033, N4128);
nor NOR2 (N4425, N4416, N2409);
or OR3 (N4426, N4423, N1802, N1873);
nand NAND4 (N4427, N4424, N1440, N450, N2062);
xor XOR2 (N4428, N4425, N3813);
and AND4 (N4429, N4427, N4045, N1982, N2376);
xor XOR2 (N4430, N4429, N1782);
and AND3 (N4431, N4417, N4414, N2210);
nor NOR2 (N4432, N4431, N1326);
nor NOR4 (N4433, N4426, N3587, N804, N1706);
not NOT1 (N4434, N4433);
buf BUF1 (N4435, N4420);
buf BUF1 (N4436, N4432);
nor NOR4 (N4437, N4418, N4206, N2256, N2010);
or OR3 (N4438, N4422, N4245, N74);
nand NAND2 (N4439, N4428, N3212);
nor NOR4 (N4440, N4430, N931, N2381, N1770);
not NOT1 (N4441, N4421);
buf BUF1 (N4442, N4434);
not NOT1 (N4443, N4436);
buf BUF1 (N4444, N4437);
and AND3 (N4445, N4444, N3534, N2104);
nand NAND2 (N4446, N4435, N4022);
not NOT1 (N4447, N4446);
or OR2 (N4448, N4445, N4273);
nand NAND4 (N4449, N4415, N2440, N3089, N1755);
nor NOR2 (N4450, N4448, N4358);
xor XOR2 (N4451, N4441, N437);
not NOT1 (N4452, N4443);
xor XOR2 (N4453, N4450, N939);
xor XOR2 (N4454, N4449, N3491);
xor XOR2 (N4455, N4442, N1552);
nor NOR3 (N4456, N4455, N3887, N1731);
nand NAND4 (N4457, N4412, N2089, N3175, N2532);
or OR2 (N4458, N4439, N3405);
nand NAND3 (N4459, N4438, N4456, N2754);
and AND3 (N4460, N2504, N2046, N2117);
nor NOR2 (N4461, N4453, N187);
nand NAND2 (N4462, N4457, N371);
buf BUF1 (N4463, N4462);
nor NOR3 (N4464, N4440, N3263, N928);
nor NOR4 (N4465, N4458, N2868, N98, N1965);
nor NOR4 (N4466, N4463, N1542, N3265, N787);
xor XOR2 (N4467, N4452, N552);
xor XOR2 (N4468, N4459, N3251);
nand NAND4 (N4469, N4467, N1500, N4157, N1521);
nor NOR3 (N4470, N4461, N791, N2260);
and AND3 (N4471, N4460, N2027, N1460);
or OR4 (N4472, N4471, N695, N2317, N3894);
and AND3 (N4473, N4466, N3412, N1626);
not NOT1 (N4474, N4465);
xor XOR2 (N4475, N4474, N2001);
or OR2 (N4476, N4475, N3919);
nor NOR2 (N4477, N4470, N3598);
xor XOR2 (N4478, N4472, N2742);
or OR4 (N4479, N4478, N1131, N4352, N1804);
nor NOR4 (N4480, N4451, N513, N348, N4128);
buf BUF1 (N4481, N4476);
nand NAND3 (N4482, N4477, N3513, N3828);
nor NOR2 (N4483, N4468, N1786);
nor NOR4 (N4484, N4482, N2718, N1244, N2969);
nand NAND3 (N4485, N4481, N451, N788);
not NOT1 (N4486, N4483);
not NOT1 (N4487, N4484);
xor XOR2 (N4488, N4485, N2190);
buf BUF1 (N4489, N4447);
nand NAND2 (N4490, N4486, N1178);
nand NAND2 (N4491, N4464, N3713);
xor XOR2 (N4492, N4488, N4098);
not NOT1 (N4493, N4492);
nand NAND3 (N4494, N4487, N3771, N2866);
and AND3 (N4495, N4469, N1466, N644);
nand NAND2 (N4496, N4494, N4156);
xor XOR2 (N4497, N4480, N2548);
buf BUF1 (N4498, N4479);
nand NAND3 (N4499, N4493, N892, N2413);
xor XOR2 (N4500, N4473, N1276);
not NOT1 (N4501, N4454);
nand NAND2 (N4502, N4501, N1007);
or OR3 (N4503, N4495, N1481, N2275);
or OR3 (N4504, N4500, N4478, N464);
nand NAND2 (N4505, N4504, N1394);
or OR2 (N4506, N4497, N3611);
xor XOR2 (N4507, N4498, N3852);
or OR3 (N4508, N4506, N2562, N2393);
nor NOR2 (N4509, N4489, N2724);
nand NAND3 (N4510, N4499, N3562, N3759);
nand NAND3 (N4511, N4490, N875, N3547);
nand NAND2 (N4512, N4496, N4437);
or OR3 (N4513, N4512, N855, N243);
not NOT1 (N4514, N4502);
not NOT1 (N4515, N4503);
buf BUF1 (N4516, N4491);
buf BUF1 (N4517, N4514);
buf BUF1 (N4518, N4515);
not NOT1 (N4519, N4505);
xor XOR2 (N4520, N4513, N2072);
and AND3 (N4521, N4520, N2875, N1431);
or OR3 (N4522, N4519, N2019, N1095);
buf BUF1 (N4523, N4511);
nor NOR3 (N4524, N4510, N2907, N3487);
buf BUF1 (N4525, N4517);
or OR3 (N4526, N4523, N2429, N2200);
nor NOR2 (N4527, N4518, N4299);
not NOT1 (N4528, N4525);
xor XOR2 (N4529, N4508, N38);
or OR4 (N4530, N4507, N4157, N3115, N617);
or OR2 (N4531, N4527, N813);
or OR2 (N4532, N4529, N307);
nor NOR3 (N4533, N4530, N291, N3584);
nor NOR4 (N4534, N4532, N2196, N2204, N1762);
nand NAND2 (N4535, N4516, N5);
not NOT1 (N4536, N4521);
not NOT1 (N4537, N4531);
nor NOR2 (N4538, N4535, N4125);
nand NAND3 (N4539, N4534, N3457, N939);
nand NAND3 (N4540, N4539, N3019, N3780);
nor NOR3 (N4541, N4524, N4131, N2740);
xor XOR2 (N4542, N4538, N1696);
or OR2 (N4543, N4542, N1424);
xor XOR2 (N4544, N4541, N300);
buf BUF1 (N4545, N4543);
buf BUF1 (N4546, N4537);
nand NAND4 (N4547, N4536, N2608, N558, N3925);
or OR3 (N4548, N4509, N1477, N3727);
xor XOR2 (N4549, N4526, N3921);
not NOT1 (N4550, N4546);
buf BUF1 (N4551, N4533);
or OR3 (N4552, N4549, N3898, N3490);
or OR2 (N4553, N4552, N1793);
nand NAND2 (N4554, N4553, N141);
and AND3 (N4555, N4547, N3579, N2622);
xor XOR2 (N4556, N4544, N3011);
and AND3 (N4557, N4550, N681, N2354);
nor NOR3 (N4558, N4557, N1308, N3986);
buf BUF1 (N4559, N4551);
and AND3 (N4560, N4528, N4517, N4502);
or OR3 (N4561, N4554, N3922, N868);
xor XOR2 (N4562, N4522, N776);
or OR4 (N4563, N4558, N2137, N1687, N3761);
and AND2 (N4564, N4540, N2048);
nor NOR4 (N4565, N4560, N520, N2847, N1248);
nand NAND2 (N4566, N4564, N2456);
and AND3 (N4567, N4561, N680, N275);
nand NAND4 (N4568, N4566, N95, N1432, N831);
buf BUF1 (N4569, N4545);
xor XOR2 (N4570, N4555, N2537);
not NOT1 (N4571, N4556);
buf BUF1 (N4572, N4563);
not NOT1 (N4573, N4571);
nand NAND3 (N4574, N4568, N21, N1378);
or OR3 (N4575, N4548, N1024, N2099);
not NOT1 (N4576, N4562);
nor NOR3 (N4577, N4572, N2574, N1678);
or OR4 (N4578, N4574, N3519, N12, N1888);
nor NOR2 (N4579, N4575, N4173);
xor XOR2 (N4580, N4579, N3254);
not NOT1 (N4581, N4576);
nor NOR3 (N4582, N4578, N2046, N2998);
or OR2 (N4583, N4582, N1351);
nand NAND3 (N4584, N4569, N823, N802);
not NOT1 (N4585, N4559);
nor NOR4 (N4586, N4580, N4406, N4014, N782);
or OR2 (N4587, N4570, N1790);
and AND2 (N4588, N4565, N2864);
or OR4 (N4589, N4567, N4409, N275, N926);
or OR3 (N4590, N4583, N452, N1169);
not NOT1 (N4591, N4587);
xor XOR2 (N4592, N4586, N1950);
and AND2 (N4593, N4588, N3688);
and AND3 (N4594, N4577, N1989, N1953);
xor XOR2 (N4595, N4590, N736);
not NOT1 (N4596, N4593);
xor XOR2 (N4597, N4581, N470);
and AND4 (N4598, N4584, N2521, N598, N2908);
or OR2 (N4599, N4598, N1274);
xor XOR2 (N4600, N4597, N3719);
nand NAND2 (N4601, N4585, N4270);
and AND4 (N4602, N4592, N2424, N3233, N1197);
or OR4 (N4603, N4602, N2662, N1207, N1481);
not NOT1 (N4604, N4596);
nor NOR2 (N4605, N4603, N4022);
and AND3 (N4606, N4601, N4273, N2510);
and AND2 (N4607, N4605, N3894);
and AND3 (N4608, N4594, N1742, N2203);
not NOT1 (N4609, N4573);
nand NAND3 (N4610, N4606, N1265, N3167);
xor XOR2 (N4611, N4609, N1739);
or OR2 (N4612, N4604, N4281);
nor NOR2 (N4613, N4608, N2186);
buf BUF1 (N4614, N4591);
and AND3 (N4615, N4589, N4300, N704);
xor XOR2 (N4616, N4615, N867);
nor NOR3 (N4617, N4599, N420, N682);
buf BUF1 (N4618, N4610);
buf BUF1 (N4619, N4617);
buf BUF1 (N4620, N4612);
not NOT1 (N4621, N4618);
and AND3 (N4622, N4620, N3730, N1045);
xor XOR2 (N4623, N4611, N2790);
buf BUF1 (N4624, N4614);
nand NAND3 (N4625, N4619, N912, N1690);
nor NOR3 (N4626, N4613, N754, N795);
not NOT1 (N4627, N4622);
and AND2 (N4628, N4627, N2382);
buf BUF1 (N4629, N4628);
nand NAND4 (N4630, N4600, N3787, N2163, N3334);
and AND3 (N4631, N4616, N1463, N681);
xor XOR2 (N4632, N4625, N3092);
or OR3 (N4633, N4621, N3535, N1481);
not NOT1 (N4634, N4607);
buf BUF1 (N4635, N4632);
nor NOR3 (N4636, N4624, N307, N553);
or OR3 (N4637, N4629, N4303, N1515);
nor NOR3 (N4638, N4595, N3780, N4625);
or OR4 (N4639, N4633, N1558, N2683, N3877);
not NOT1 (N4640, N4631);
nand NAND3 (N4641, N4640, N3164, N3768);
buf BUF1 (N4642, N4639);
and AND4 (N4643, N4636, N3132, N2248, N2267);
and AND4 (N4644, N4637, N3746, N2318, N227);
buf BUF1 (N4645, N4635);
and AND2 (N4646, N4623, N1425);
nand NAND3 (N4647, N4643, N2817, N4053);
or OR3 (N4648, N4634, N1517, N3475);
buf BUF1 (N4649, N4642);
or OR3 (N4650, N4630, N1089, N2114);
and AND4 (N4651, N4638, N219, N2669, N1662);
buf BUF1 (N4652, N4650);
nor NOR3 (N4653, N4645, N1650, N1094);
xor XOR2 (N4654, N4649, N4077);
not NOT1 (N4655, N4626);
or OR4 (N4656, N4653, N4170, N3023, N2606);
buf BUF1 (N4657, N4641);
not NOT1 (N4658, N4651);
nor NOR4 (N4659, N4655, N4304, N3863, N923);
not NOT1 (N4660, N4644);
xor XOR2 (N4661, N4657, N4224);
nand NAND3 (N4662, N4660, N4540, N3285);
buf BUF1 (N4663, N4658);
and AND2 (N4664, N4663, N4376);
nand NAND2 (N4665, N4646, N1684);
nand NAND3 (N4666, N4656, N697, N3227);
nor NOR2 (N4667, N4654, N3207);
not NOT1 (N4668, N4664);
and AND3 (N4669, N4647, N1471, N80);
nand NAND3 (N4670, N4662, N3409, N1634);
nor NOR2 (N4671, N4667, N2540);
nand NAND2 (N4672, N4669, N1053);
buf BUF1 (N4673, N4665);
not NOT1 (N4674, N4659);
or OR4 (N4675, N4661, N1640, N2191, N1180);
xor XOR2 (N4676, N4672, N4649);
not NOT1 (N4677, N4670);
nor NOR2 (N4678, N4676, N4388);
and AND4 (N4679, N4648, N1541, N2843, N3607);
xor XOR2 (N4680, N4677, N4329);
nor NOR3 (N4681, N4673, N572, N153);
or OR2 (N4682, N4666, N3561);
buf BUF1 (N4683, N4682);
nor NOR3 (N4684, N4683, N512, N2038);
nand NAND4 (N4685, N4668, N1884, N4316, N493);
nand NAND2 (N4686, N4685, N378);
not NOT1 (N4687, N4675);
nor NOR3 (N4688, N4671, N4347, N346);
nor NOR3 (N4689, N4678, N3843, N2787);
and AND3 (N4690, N4652, N139, N4277);
buf BUF1 (N4691, N4690);
not NOT1 (N4692, N4691);
and AND4 (N4693, N4681, N4001, N2578, N1683);
buf BUF1 (N4694, N4674);
nor NOR4 (N4695, N4679, N3987, N2563, N4654);
not NOT1 (N4696, N4687);
buf BUF1 (N4697, N4692);
buf BUF1 (N4698, N4689);
or OR2 (N4699, N4693, N2961);
xor XOR2 (N4700, N4688, N3084);
or OR3 (N4701, N4684, N804, N665);
nand NAND2 (N4702, N4694, N4677);
xor XOR2 (N4703, N4700, N2646);
nor NOR2 (N4704, N4703, N511);
or OR4 (N4705, N4696, N3829, N1479, N729);
or OR3 (N4706, N4704, N632, N912);
and AND4 (N4707, N4699, N918, N3929, N520);
buf BUF1 (N4708, N4706);
buf BUF1 (N4709, N4707);
or OR2 (N4710, N4698, N1732);
nor NOR3 (N4711, N4686, N526, N1703);
xor XOR2 (N4712, N4711, N1229);
not NOT1 (N4713, N4697);
nor NOR2 (N4714, N4708, N2838);
not NOT1 (N4715, N4702);
buf BUF1 (N4716, N4714);
and AND3 (N4717, N4680, N916, N394);
xor XOR2 (N4718, N4716, N2119);
and AND3 (N4719, N4710, N1972, N3319);
buf BUF1 (N4720, N4715);
nor NOR4 (N4721, N4720, N3265, N2617, N521);
buf BUF1 (N4722, N4709);
or OR3 (N4723, N4701, N2548, N447);
nand NAND4 (N4724, N4723, N3756, N468, N3763);
not NOT1 (N4725, N4705);
nor NOR2 (N4726, N4722, N1410);
not NOT1 (N4727, N4718);
not NOT1 (N4728, N4695);
or OR3 (N4729, N4719, N3908, N2309);
nand NAND3 (N4730, N4729, N2870, N3278);
and AND4 (N4731, N4730, N3446, N3119, N3631);
buf BUF1 (N4732, N4727);
not NOT1 (N4733, N4728);
buf BUF1 (N4734, N4721);
xor XOR2 (N4735, N4732, N827);
nand NAND3 (N4736, N4734, N1266, N811);
xor XOR2 (N4737, N4736, N1156);
xor XOR2 (N4738, N4733, N305);
buf BUF1 (N4739, N4725);
nor NOR2 (N4740, N4731, N19);
not NOT1 (N4741, N4726);
buf BUF1 (N4742, N4739);
nor NOR3 (N4743, N4735, N2538, N4439);
nor NOR2 (N4744, N4741, N609);
xor XOR2 (N4745, N4712, N3767);
buf BUF1 (N4746, N4745);
nor NOR4 (N4747, N4744, N1943, N3998, N1005);
not NOT1 (N4748, N4747);
not NOT1 (N4749, N4748);
not NOT1 (N4750, N4746);
not NOT1 (N4751, N4724);
nor NOR3 (N4752, N4742, N389, N4519);
nand NAND2 (N4753, N4737, N3488);
or OR3 (N4754, N4749, N3948, N3254);
nand NAND2 (N4755, N4750, N3118);
and AND2 (N4756, N4754, N1941);
xor XOR2 (N4757, N4755, N2274);
and AND3 (N4758, N4756, N1773, N2472);
nor NOR3 (N4759, N4752, N797, N2324);
buf BUF1 (N4760, N4740);
nand NAND3 (N4761, N4751, N35, N2866);
nor NOR3 (N4762, N4758, N2652, N3612);
xor XOR2 (N4763, N4743, N4467);
nand NAND2 (N4764, N4762, N4153);
xor XOR2 (N4765, N4759, N1044);
not NOT1 (N4766, N4757);
or OR4 (N4767, N4713, N1595, N416, N1777);
buf BUF1 (N4768, N4738);
buf BUF1 (N4769, N4717);
or OR2 (N4770, N4753, N4341);
or OR3 (N4771, N4769, N3992, N836);
and AND2 (N4772, N4763, N3305);
nor NOR3 (N4773, N4766, N35, N4698);
and AND2 (N4774, N4765, N1679);
and AND2 (N4775, N4773, N3304);
buf BUF1 (N4776, N4774);
not NOT1 (N4777, N4771);
and AND4 (N4778, N4760, N4593, N3768, N82);
or OR4 (N4779, N4767, N1209, N4269, N1135);
nor NOR4 (N4780, N4776, N2470, N4603, N2840);
and AND3 (N4781, N4779, N4602, N2748);
xor XOR2 (N4782, N4777, N1969);
nand NAND2 (N4783, N4781, N1812);
not NOT1 (N4784, N4780);
not NOT1 (N4785, N4783);
nor NOR2 (N4786, N4770, N722);
xor XOR2 (N4787, N4786, N3844);
xor XOR2 (N4788, N4782, N3956);
nor NOR4 (N4789, N4761, N1558, N1892, N2169);
nand NAND4 (N4790, N4785, N1078, N3885, N2271);
nand NAND4 (N4791, N4772, N4298, N2445, N4785);
nor NOR3 (N4792, N4775, N2645, N3437);
not NOT1 (N4793, N4778);
or OR4 (N4794, N4791, N4665, N1488, N2089);
and AND2 (N4795, N4787, N2474);
not NOT1 (N4796, N4764);
and AND2 (N4797, N4796, N1949);
not NOT1 (N4798, N4794);
not NOT1 (N4799, N4789);
nor NOR4 (N4800, N4784, N990, N2583, N1727);
nor NOR4 (N4801, N4800, N788, N158, N214);
nand NAND2 (N4802, N4790, N3250);
nand NAND3 (N4803, N4799, N3022, N2616);
and AND4 (N4804, N4802, N114, N630, N361);
not NOT1 (N4805, N4768);
and AND2 (N4806, N4793, N2907);
buf BUF1 (N4807, N4798);
nor NOR3 (N4808, N4804, N3945, N818);
or OR3 (N4809, N4801, N4682, N379);
buf BUF1 (N4810, N4805);
xor XOR2 (N4811, N4795, N3519);
nor NOR2 (N4812, N4797, N104);
buf BUF1 (N4813, N4812);
xor XOR2 (N4814, N4806, N2358);
nand NAND4 (N4815, N4808, N4316, N3417, N369);
nor NOR3 (N4816, N4813, N2922, N3050);
xor XOR2 (N4817, N4807, N3871);
xor XOR2 (N4818, N4817, N1595);
nand NAND2 (N4819, N4810, N83);
nor NOR4 (N4820, N4803, N31, N914, N2844);
buf BUF1 (N4821, N4815);
nand NAND3 (N4822, N4821, N589, N400);
nor NOR3 (N4823, N4820, N1823, N792);
buf BUF1 (N4824, N4788);
or OR3 (N4825, N4824, N3799, N3902);
nand NAND4 (N4826, N4823, N1394, N2474, N3261);
not NOT1 (N4827, N4809);
xor XOR2 (N4828, N4816, N3470);
or OR3 (N4829, N4827, N2285, N2981);
and AND2 (N4830, N4829, N2696);
or OR4 (N4831, N4792, N1166, N2790, N290);
nor NOR2 (N4832, N4818, N4039);
nor NOR4 (N4833, N4822, N1013, N1893, N2961);
and AND3 (N4834, N4814, N3577, N3556);
nor NOR4 (N4835, N4833, N884, N2540, N3424);
or OR2 (N4836, N4828, N1243);
and AND3 (N4837, N4825, N3266, N410);
buf BUF1 (N4838, N4819);
or OR4 (N4839, N4811, N2082, N755, N3552);
and AND3 (N4840, N4838, N1995, N1272);
or OR3 (N4841, N4836, N1483, N819);
buf BUF1 (N4842, N4831);
and AND3 (N4843, N4826, N1343, N396);
and AND2 (N4844, N4835, N1075);
buf BUF1 (N4845, N4832);
buf BUF1 (N4846, N4837);
buf BUF1 (N4847, N4830);
buf BUF1 (N4848, N4845);
xor XOR2 (N4849, N4834, N4587);
or OR4 (N4850, N4848, N618, N1046, N1548);
and AND2 (N4851, N4843, N2587);
buf BUF1 (N4852, N4851);
not NOT1 (N4853, N4839);
nor NOR2 (N4854, N4852, N4096);
buf BUF1 (N4855, N4844);
xor XOR2 (N4856, N4847, N2980);
buf BUF1 (N4857, N4850);
not NOT1 (N4858, N4849);
not NOT1 (N4859, N4842);
not NOT1 (N4860, N4841);
and AND2 (N4861, N4857, N1162);
or OR4 (N4862, N4854, N639, N4103, N4432);
buf BUF1 (N4863, N4860);
or OR4 (N4864, N4855, N2801, N1762, N1316);
nor NOR3 (N4865, N4862, N4197, N316);
xor XOR2 (N4866, N4865, N4361);
not NOT1 (N4867, N4866);
buf BUF1 (N4868, N4867);
and AND2 (N4869, N4840, N4675);
or OR3 (N4870, N4864, N3019, N4023);
nand NAND4 (N4871, N4853, N1282, N1556, N4621);
nand NAND3 (N4872, N4871, N3032, N4771);
nor NOR2 (N4873, N4858, N3249);
not NOT1 (N4874, N4846);
nand NAND3 (N4875, N4863, N2914, N2115);
not NOT1 (N4876, N4868);
xor XOR2 (N4877, N4859, N1472);
and AND2 (N4878, N4861, N2306);
and AND4 (N4879, N4873, N3718, N36, N1136);
xor XOR2 (N4880, N4874, N580);
nand NAND2 (N4881, N4880, N1267);
nand NAND4 (N4882, N4878, N517, N1613, N187);
nand NAND4 (N4883, N4879, N3853, N59, N3688);
nand NAND2 (N4884, N4883, N2534);
buf BUF1 (N4885, N4884);
xor XOR2 (N4886, N4877, N815);
nor NOR4 (N4887, N4856, N1785, N1624, N3081);
and AND2 (N4888, N4876, N642);
buf BUF1 (N4889, N4869);
xor XOR2 (N4890, N4885, N2759);
and AND3 (N4891, N4872, N3854, N3005);
xor XOR2 (N4892, N4888, N3545);
not NOT1 (N4893, N4881);
not NOT1 (N4894, N4882);
not NOT1 (N4895, N4891);
or OR2 (N4896, N4875, N4070);
nor NOR2 (N4897, N4895, N97);
nand NAND3 (N4898, N4870, N1270, N3353);
buf BUF1 (N4899, N4890);
and AND4 (N4900, N4896, N3659, N1211, N818);
xor XOR2 (N4901, N4900, N3207);
or OR2 (N4902, N4901, N2694);
and AND4 (N4903, N4898, N631, N2205, N159);
buf BUF1 (N4904, N4886);
buf BUF1 (N4905, N4903);
nor NOR3 (N4906, N4899, N1932, N3617);
nor NOR3 (N4907, N4905, N3136, N2855);
not NOT1 (N4908, N4906);
or OR3 (N4909, N4887, N3007, N2407);
xor XOR2 (N4910, N4908, N2252);
and AND2 (N4911, N4909, N871);
and AND2 (N4912, N4907, N3451);
nand NAND3 (N4913, N4912, N360, N3311);
xor XOR2 (N4914, N4910, N3298);
xor XOR2 (N4915, N4892, N2273);
nor NOR2 (N4916, N4914, N4422);
and AND2 (N4917, N4894, N3435);
or OR3 (N4918, N4915, N1167, N3883);
buf BUF1 (N4919, N4904);
nor NOR2 (N4920, N4889, N2489);
nand NAND3 (N4921, N4893, N4486, N1303);
and AND3 (N4922, N4917, N1268, N873);
xor XOR2 (N4923, N4921, N4378);
nor NOR2 (N4924, N4897, N545);
or OR3 (N4925, N4911, N2199, N598);
nor NOR3 (N4926, N4924, N1982, N3650);
nor NOR2 (N4927, N4919, N2544);
nor NOR4 (N4928, N4922, N1712, N3467, N3354);
and AND4 (N4929, N4916, N1068, N3215, N921);
buf BUF1 (N4930, N4926);
buf BUF1 (N4931, N4918);
nand NAND2 (N4932, N4920, N2915);
and AND2 (N4933, N4928, N3999);
nand NAND2 (N4934, N4902, N80);
nand NAND3 (N4935, N4933, N2488, N1228);
xor XOR2 (N4936, N4929, N789);
and AND3 (N4937, N4923, N3076, N749);
nand NAND3 (N4938, N4932, N1021, N4845);
not NOT1 (N4939, N4938);
nand NAND2 (N4940, N4930, N3604);
or OR4 (N4941, N4939, N4376, N3094, N1744);
buf BUF1 (N4942, N4937);
not NOT1 (N4943, N4935);
buf BUF1 (N4944, N4925);
buf BUF1 (N4945, N4913);
nor NOR2 (N4946, N4942, N4115);
nor NOR3 (N4947, N4934, N295, N2533);
xor XOR2 (N4948, N4940, N4425);
and AND4 (N4949, N4927, N4749, N2760, N763);
xor XOR2 (N4950, N4931, N4643);
nor NOR2 (N4951, N4941, N2043);
and AND4 (N4952, N4943, N353, N3407, N1970);
not NOT1 (N4953, N4944);
buf BUF1 (N4954, N4951);
xor XOR2 (N4955, N4945, N2238);
nand NAND2 (N4956, N4949, N3236);
nor NOR3 (N4957, N4953, N242, N3410);
not NOT1 (N4958, N4956);
nand NAND4 (N4959, N4947, N1481, N2532, N4626);
buf BUF1 (N4960, N4959);
nor NOR4 (N4961, N4958, N993, N610, N4631);
xor XOR2 (N4962, N4955, N720);
not NOT1 (N4963, N4936);
nand NAND4 (N4964, N4954, N4622, N3251, N3237);
buf BUF1 (N4965, N4962);
not NOT1 (N4966, N4948);
nor NOR2 (N4967, N4963, N1486);
nor NOR2 (N4968, N4960, N2658);
nand NAND2 (N4969, N4965, N4902);
nand NAND2 (N4970, N4950, N1408);
or OR3 (N4971, N4964, N1892, N2721);
not NOT1 (N4972, N4952);
and AND4 (N4973, N4957, N3937, N773, N4431);
and AND2 (N4974, N4972, N3477);
buf BUF1 (N4975, N4973);
or OR3 (N4976, N4967, N1814, N3369);
nand NAND4 (N4977, N4975, N4630, N2670, N2169);
not NOT1 (N4978, N4968);
nand NAND4 (N4979, N4969, N1255, N1884, N1007);
or OR3 (N4980, N4961, N626, N2531);
and AND3 (N4981, N4970, N1395, N4306);
buf BUF1 (N4982, N4976);
nand NAND3 (N4983, N4977, N784, N2560);
not NOT1 (N4984, N4974);
and AND4 (N4985, N4966, N3349, N1955, N3906);
not NOT1 (N4986, N4946);
or OR4 (N4987, N4985, N3995, N1754, N573);
buf BUF1 (N4988, N4971);
nand NAND2 (N4989, N4986, N1643);
nand NAND3 (N4990, N4978, N4248, N1031);
nand NAND4 (N4991, N4979, N4113, N228, N4026);
and AND3 (N4992, N4982, N625, N969);
not NOT1 (N4993, N4987);
or OR4 (N4994, N4984, N590, N3700, N2940);
or OR2 (N4995, N4993, N1347);
buf BUF1 (N4996, N4988);
buf BUF1 (N4997, N4983);
and AND4 (N4998, N4997, N1533, N4967, N4431);
or OR2 (N4999, N4989, N748);
nand NAND2 (N5000, N4996, N4472);
not NOT1 (N5001, N4999);
not NOT1 (N5002, N4980);
xor XOR2 (N5003, N4995, N2244);
xor XOR2 (N5004, N4981, N882);
nand NAND2 (N5005, N5004, N2688);
not NOT1 (N5006, N5001);
or OR2 (N5007, N5005, N1368);
nand NAND3 (N5008, N4991, N4137, N3194);
or OR2 (N5009, N4994, N2065);
or OR4 (N5010, N5000, N1901, N1065, N16);
not NOT1 (N5011, N5003);
buf BUF1 (N5012, N5002);
nand NAND2 (N5013, N5011, N3525);
buf BUF1 (N5014, N5012);
nand NAND2 (N5015, N5014, N92);
or OR2 (N5016, N5006, N1518);
or OR2 (N5017, N5016, N2152);
not NOT1 (N5018, N5013);
not NOT1 (N5019, N5015);
nand NAND4 (N5020, N5007, N188, N1876, N778);
xor XOR2 (N5021, N5010, N4737);
buf BUF1 (N5022, N4990);
xor XOR2 (N5023, N5018, N4745);
or OR3 (N5024, N5017, N4971, N3553);
or OR3 (N5025, N4992, N1048, N3496);
and AND3 (N5026, N5023, N1175, N4013);
not NOT1 (N5027, N5026);
nand NAND2 (N5028, N5009, N375);
nor NOR3 (N5029, N5020, N1087, N2787);
or OR2 (N5030, N5025, N622);
not NOT1 (N5031, N5019);
nor NOR4 (N5032, N5024, N4723, N3913, N4741);
and AND4 (N5033, N5022, N3013, N2959, N1446);
xor XOR2 (N5034, N5021, N1750);
or OR3 (N5035, N5008, N489, N148);
or OR3 (N5036, N5033, N3788, N1067);
xor XOR2 (N5037, N5030, N1119);
and AND2 (N5038, N5031, N2722);
xor XOR2 (N5039, N5032, N2821);
nor NOR2 (N5040, N5034, N390);
xor XOR2 (N5041, N5039, N1164);
nand NAND4 (N5042, N5028, N3003, N2661, N139);
buf BUF1 (N5043, N5041);
buf BUF1 (N5044, N4998);
buf BUF1 (N5045, N5036);
and AND2 (N5046, N5027, N4457);
or OR4 (N5047, N5035, N2649, N263, N4847);
nor NOR3 (N5048, N5045, N3760, N2927);
and AND3 (N5049, N5042, N637, N3779);
or OR4 (N5050, N5038, N1325, N508, N2819);
not NOT1 (N5051, N5047);
nand NAND4 (N5052, N5040, N4272, N2040, N1159);
or OR4 (N5053, N5037, N492, N459, N4817);
buf BUF1 (N5054, N5049);
xor XOR2 (N5055, N5053, N753);
or OR4 (N5056, N5054, N388, N1957, N2219);
or OR2 (N5057, N5050, N3514);
or OR2 (N5058, N5048, N3188);
xor XOR2 (N5059, N5029, N2989);
nand NAND2 (N5060, N5059, N1608);
nand NAND3 (N5061, N5055, N349, N997);
nor NOR3 (N5062, N5046, N2977, N3629);
nand NAND2 (N5063, N5060, N4263);
buf BUF1 (N5064, N5063);
buf BUF1 (N5065, N5061);
buf BUF1 (N5066, N5056);
buf BUF1 (N5067, N5065);
nand NAND2 (N5068, N5051, N1790);
nand NAND2 (N5069, N5066, N2286);
not NOT1 (N5070, N5052);
nor NOR2 (N5071, N5067, N356);
buf BUF1 (N5072, N5070);
not NOT1 (N5073, N5058);
and AND3 (N5074, N5062, N3431, N879);
or OR4 (N5075, N5072, N4237, N3480, N1054);
not NOT1 (N5076, N5064);
and AND2 (N5077, N5075, N1849);
not NOT1 (N5078, N5074);
nor NOR4 (N5079, N5077, N1661, N809, N1952);
buf BUF1 (N5080, N5073);
not NOT1 (N5081, N5044);
not NOT1 (N5082, N5081);
not NOT1 (N5083, N5082);
buf BUF1 (N5084, N5079);
nor NOR3 (N5085, N5076, N1040, N3468);
xor XOR2 (N5086, N5084, N1205);
and AND2 (N5087, N5071, N238);
and AND4 (N5088, N5085, N2366, N3190, N603);
buf BUF1 (N5089, N5083);
not NOT1 (N5090, N5068);
buf BUF1 (N5091, N5087);
or OR2 (N5092, N5043, N4961);
nor NOR3 (N5093, N5057, N2317, N4442);
buf BUF1 (N5094, N5091);
nand NAND4 (N5095, N5080, N995, N1303, N808);
nor NOR4 (N5096, N5069, N993, N2151, N3171);
nor NOR3 (N5097, N5094, N4374, N16);
nor NOR4 (N5098, N5093, N4904, N2764, N1212);
and AND2 (N5099, N5089, N532);
nor NOR3 (N5100, N5097, N2842, N920);
nand NAND3 (N5101, N5078, N1248, N2721);
and AND2 (N5102, N5090, N1358);
nor NOR2 (N5103, N5095, N4356);
nor NOR3 (N5104, N5098, N2923, N2163);
and AND4 (N5105, N5101, N4267, N2154, N3324);
or OR3 (N5106, N5092, N3775, N2157);
nand NAND2 (N5107, N5106, N2910);
xor XOR2 (N5108, N5105, N240);
xor XOR2 (N5109, N5100, N2829);
xor XOR2 (N5110, N5102, N805);
nor NOR3 (N5111, N5110, N1837, N2621);
not NOT1 (N5112, N5088);
and AND3 (N5113, N5109, N3120, N3241);
and AND3 (N5114, N5104, N384, N1610);
xor XOR2 (N5115, N5112, N2675);
and AND4 (N5116, N5086, N678, N317, N4103);
or OR4 (N5117, N5113, N3266, N2493, N2256);
buf BUF1 (N5118, N5108);
and AND3 (N5119, N5107, N2742, N741);
nand NAND2 (N5120, N5115, N4531);
nand NAND2 (N5121, N5111, N2919);
nand NAND4 (N5122, N5120, N4565, N3860, N2559);
and AND4 (N5123, N5117, N4159, N4147, N1611);
buf BUF1 (N5124, N5096);
and AND2 (N5125, N5118, N2622);
or OR2 (N5126, N5121, N4095);
or OR3 (N5127, N5125, N1572, N3662);
nand NAND4 (N5128, N5123, N1309, N3408, N4192);
nand NAND2 (N5129, N5103, N2293);
nand NAND3 (N5130, N5126, N1225, N2451);
xor XOR2 (N5131, N5127, N1662);
xor XOR2 (N5132, N5124, N4543);
xor XOR2 (N5133, N5122, N184);
nand NAND4 (N5134, N5130, N5030, N4050, N690);
xor XOR2 (N5135, N5133, N5062);
nand NAND2 (N5136, N5132, N5115);
or OR3 (N5137, N5099, N4015, N4150);
buf BUF1 (N5138, N5114);
and AND3 (N5139, N5116, N4151, N4837);
not NOT1 (N5140, N5135);
buf BUF1 (N5141, N5139);
xor XOR2 (N5142, N5136, N4589);
and AND3 (N5143, N5142, N2205, N406);
xor XOR2 (N5144, N5143, N3407);
or OR2 (N5145, N5141, N782);
not NOT1 (N5146, N5119);
nand NAND3 (N5147, N5145, N1465, N2635);
xor XOR2 (N5148, N5134, N544);
and AND4 (N5149, N5138, N4347, N1412, N1426);
and AND2 (N5150, N5148, N234);
nand NAND3 (N5151, N5150, N4518, N9);
buf BUF1 (N5152, N5144);
not NOT1 (N5153, N5151);
xor XOR2 (N5154, N5137, N217);
and AND2 (N5155, N5149, N4872);
not NOT1 (N5156, N5152);
not NOT1 (N5157, N5129);
xor XOR2 (N5158, N5153, N3773);
and AND2 (N5159, N5157, N1575);
not NOT1 (N5160, N5158);
buf BUF1 (N5161, N5155);
not NOT1 (N5162, N5128);
and AND4 (N5163, N5156, N1774, N1612, N3003);
nor NOR2 (N5164, N5154, N3925);
nor NOR4 (N5165, N5159, N2465, N2651, N4418);
and AND4 (N5166, N5146, N216, N3944, N1875);
nor NOR3 (N5167, N5161, N471, N5023);
buf BUF1 (N5168, N5166);
nor NOR4 (N5169, N5131, N4878, N3711, N1263);
and AND4 (N5170, N5163, N3387, N214, N2816);
not NOT1 (N5171, N5167);
buf BUF1 (N5172, N5147);
xor XOR2 (N5173, N5164, N816);
not NOT1 (N5174, N5168);
nor NOR2 (N5175, N5165, N3425);
xor XOR2 (N5176, N5170, N250);
and AND3 (N5177, N5160, N3928, N3181);
not NOT1 (N5178, N5162);
buf BUF1 (N5179, N5175);
xor XOR2 (N5180, N5173, N3211);
xor XOR2 (N5181, N5177, N962);
and AND3 (N5182, N5181, N927, N3735);
xor XOR2 (N5183, N5174, N2518);
buf BUF1 (N5184, N5176);
or OR4 (N5185, N5171, N188, N2510, N2769);
xor XOR2 (N5186, N5178, N2377);
or OR4 (N5187, N5183, N4079, N1945, N1770);
xor XOR2 (N5188, N5182, N3896);
nor NOR4 (N5189, N5184, N3807, N3514, N3797);
and AND4 (N5190, N5140, N5151, N1837, N1166);
xor XOR2 (N5191, N5187, N2123);
not NOT1 (N5192, N5172);
and AND2 (N5193, N5186, N4974);
nand NAND2 (N5194, N5169, N4754);
nand NAND2 (N5195, N5193, N3419);
or OR3 (N5196, N5192, N4099, N1162);
nand NAND2 (N5197, N5196, N4680);
and AND4 (N5198, N5197, N1622, N760, N327);
xor XOR2 (N5199, N5194, N2107);
nand NAND3 (N5200, N5185, N1966, N1366);
or OR4 (N5201, N5180, N1852, N2417, N2691);
nand NAND4 (N5202, N5190, N3321, N862, N3347);
buf BUF1 (N5203, N5191);
buf BUF1 (N5204, N5200);
nand NAND3 (N5205, N5204, N441, N4224);
xor XOR2 (N5206, N5179, N415);
and AND3 (N5207, N5202, N3900, N3591);
nand NAND2 (N5208, N5207, N2674);
or OR2 (N5209, N5195, N1410);
or OR4 (N5210, N5203, N3608, N1227, N4888);
buf BUF1 (N5211, N5201);
not NOT1 (N5212, N5210);
buf BUF1 (N5213, N5189);
or OR4 (N5214, N5213, N180, N4732, N1802);
or OR3 (N5215, N5198, N2350, N4415);
xor XOR2 (N5216, N5212, N2121);
nand NAND3 (N5217, N5209, N950, N4297);
nor NOR4 (N5218, N5205, N4935, N1390, N1979);
not NOT1 (N5219, N5216);
not NOT1 (N5220, N5215);
and AND4 (N5221, N5188, N16, N1405, N3821);
buf BUF1 (N5222, N5199);
and AND4 (N5223, N5220, N2088, N1608, N339);
and AND4 (N5224, N5222, N2313, N1525, N428);
and AND4 (N5225, N5208, N2691, N4514, N4609);
buf BUF1 (N5226, N5224);
xor XOR2 (N5227, N5214, N3972);
nor NOR4 (N5228, N5225, N3796, N4266, N126);
or OR3 (N5229, N5219, N552, N702);
and AND4 (N5230, N5218, N2892, N4699, N1839);
and AND4 (N5231, N5221, N2417, N3222, N401);
or OR4 (N5232, N5228, N913, N1306, N1672);
or OR3 (N5233, N5230, N3547, N2720);
buf BUF1 (N5234, N5223);
buf BUF1 (N5235, N5217);
buf BUF1 (N5236, N5226);
not NOT1 (N5237, N5206);
or OR4 (N5238, N5235, N3723, N5118, N3);
buf BUF1 (N5239, N5238);
xor XOR2 (N5240, N5229, N3893);
buf BUF1 (N5241, N5236);
buf BUF1 (N5242, N5227);
buf BUF1 (N5243, N5233);
and AND4 (N5244, N5242, N3748, N68, N1019);
or OR4 (N5245, N5234, N2194, N2056, N4499);
or OR3 (N5246, N5244, N4247, N2437);
xor XOR2 (N5247, N5240, N1409);
or OR4 (N5248, N5239, N2053, N4568, N1016);
or OR2 (N5249, N5248, N1499);
or OR3 (N5250, N5247, N286, N3325);
buf BUF1 (N5251, N5232);
nand NAND2 (N5252, N5245, N260);
xor XOR2 (N5253, N5250, N4090);
and AND3 (N5254, N5243, N4952, N510);
buf BUF1 (N5255, N5254);
buf BUF1 (N5256, N5231);
xor XOR2 (N5257, N5251, N2223);
and AND4 (N5258, N5246, N805, N3789, N1153);
and AND4 (N5259, N5249, N4600, N347, N2056);
xor XOR2 (N5260, N5259, N1943);
or OR4 (N5261, N5211, N406, N4549, N1149);
not NOT1 (N5262, N5260);
xor XOR2 (N5263, N5241, N994);
or OR3 (N5264, N5255, N2758, N4648);
or OR4 (N5265, N5256, N1247, N4304, N3690);
or OR2 (N5266, N5262, N116);
xor XOR2 (N5267, N5261, N717);
or OR2 (N5268, N5265, N253);
and AND3 (N5269, N5257, N974, N3544);
and AND3 (N5270, N5253, N3576, N3449);
nor NOR2 (N5271, N5237, N1630);
xor XOR2 (N5272, N5271, N4638);
nand NAND3 (N5273, N5272, N3583, N649);
or OR4 (N5274, N5269, N917, N3362, N4782);
xor XOR2 (N5275, N5264, N4058);
and AND4 (N5276, N5263, N1841, N3502, N5060);
buf BUF1 (N5277, N5275);
nand NAND2 (N5278, N5274, N3381);
nand NAND4 (N5279, N5267, N432, N4553, N1664);
and AND3 (N5280, N5276, N48, N741);
or OR4 (N5281, N5268, N746, N1733, N4954);
buf BUF1 (N5282, N5252);
buf BUF1 (N5283, N5278);
nand NAND4 (N5284, N5258, N1058, N4050, N700);
nor NOR3 (N5285, N5279, N351, N2872);
xor XOR2 (N5286, N5284, N1208);
buf BUF1 (N5287, N5285);
buf BUF1 (N5288, N5281);
xor XOR2 (N5289, N5283, N1428);
nor NOR4 (N5290, N5286, N4766, N2420, N176);
xor XOR2 (N5291, N5282, N294);
or OR2 (N5292, N5291, N20);
and AND3 (N5293, N5280, N2668, N4847);
or OR4 (N5294, N5266, N2094, N1298, N1110);
and AND3 (N5295, N5287, N2621, N2942);
nand NAND2 (N5296, N5290, N1408);
and AND4 (N5297, N5296, N2615, N1572, N829);
or OR2 (N5298, N5270, N2181);
nand NAND4 (N5299, N5294, N4519, N3284, N1361);
nand NAND4 (N5300, N5298, N1164, N1085, N5299);
buf BUF1 (N5301, N2958);
nand NAND4 (N5302, N5273, N908, N4784, N1565);
nor NOR3 (N5303, N5289, N1724, N817);
xor XOR2 (N5304, N5303, N2076);
and AND3 (N5305, N5302, N3492, N2949);
xor XOR2 (N5306, N5300, N221);
buf BUF1 (N5307, N5277);
not NOT1 (N5308, N5295);
buf BUF1 (N5309, N5293);
and AND2 (N5310, N5308, N2608);
nor NOR4 (N5311, N5310, N3021, N4868, N1148);
nor NOR4 (N5312, N5301, N3349, N1669, N5174);
and AND4 (N5313, N5305, N3659, N2331, N3479);
or OR2 (N5314, N5288, N1819);
not NOT1 (N5315, N5311);
nor NOR2 (N5316, N5297, N1483);
xor XOR2 (N5317, N5292, N1435);
nor NOR3 (N5318, N5316, N1804, N3105);
buf BUF1 (N5319, N5313);
buf BUF1 (N5320, N5304);
xor XOR2 (N5321, N5307, N3159);
and AND3 (N5322, N5315, N4229, N880);
nor NOR4 (N5323, N5312, N4133, N4796, N2369);
or OR3 (N5324, N5318, N2549, N2043);
nor NOR2 (N5325, N5319, N2289);
or OR4 (N5326, N5320, N3748, N727, N4691);
buf BUF1 (N5327, N5314);
or OR2 (N5328, N5323, N3540);
and AND2 (N5329, N5309, N4077);
and AND4 (N5330, N5322, N3989, N352, N4770);
or OR2 (N5331, N5321, N201);
not NOT1 (N5332, N5328);
buf BUF1 (N5333, N5327);
xor XOR2 (N5334, N5326, N3172);
or OR2 (N5335, N5333, N2255);
xor XOR2 (N5336, N5331, N170);
or OR2 (N5337, N5332, N1039);
buf BUF1 (N5338, N5330);
xor XOR2 (N5339, N5325, N1896);
nand NAND3 (N5340, N5338, N2663, N2558);
xor XOR2 (N5341, N5324, N4802);
nor NOR2 (N5342, N5306, N3086);
or OR4 (N5343, N5340, N2408, N1774, N1391);
and AND4 (N5344, N5334, N2265, N3410, N910);
and AND2 (N5345, N5341, N4210);
or OR3 (N5346, N5342, N4547, N1922);
nor NOR3 (N5347, N5336, N3831, N5079);
nand NAND4 (N5348, N5346, N3869, N1632, N1726);
or OR2 (N5349, N5343, N4357);
not NOT1 (N5350, N5339);
not NOT1 (N5351, N5347);
xor XOR2 (N5352, N5348, N2787);
xor XOR2 (N5353, N5350, N3682);
xor XOR2 (N5354, N5317, N854);
nand NAND3 (N5355, N5344, N3686, N5133);
not NOT1 (N5356, N5351);
not NOT1 (N5357, N5355);
or OR3 (N5358, N5329, N1128, N5129);
buf BUF1 (N5359, N5356);
nor NOR2 (N5360, N5345, N2611);
nor NOR3 (N5361, N5358, N3187, N4156);
buf BUF1 (N5362, N5353);
nor NOR4 (N5363, N5349, N2718, N5320, N932);
not NOT1 (N5364, N5362);
not NOT1 (N5365, N5361);
or OR4 (N5366, N5335, N585, N3144, N4290);
nor NOR4 (N5367, N5352, N4090, N522, N4395);
nand NAND2 (N5368, N5359, N3639);
nand NAND2 (N5369, N5365, N2462);
and AND4 (N5370, N5368, N4844, N1579, N1094);
xor XOR2 (N5371, N5370, N389);
or OR2 (N5372, N5360, N1642);
not NOT1 (N5373, N5372);
nand NAND4 (N5374, N5363, N1134, N2531, N748);
nor NOR3 (N5375, N5374, N4711, N1446);
and AND4 (N5376, N5371, N1199, N4146, N4706);
and AND4 (N5377, N5337, N2330, N1089, N2816);
or OR4 (N5378, N5377, N3877, N2950, N1671);
or OR2 (N5379, N5354, N2125);
xor XOR2 (N5380, N5364, N1747);
nand NAND4 (N5381, N5379, N4730, N2003, N3526);
nand NAND3 (N5382, N5373, N1799, N538);
buf BUF1 (N5383, N5357);
nand NAND3 (N5384, N5380, N2602, N2380);
buf BUF1 (N5385, N5376);
or OR2 (N5386, N5382, N3198);
or OR2 (N5387, N5385, N3603);
not NOT1 (N5388, N5369);
nor NOR2 (N5389, N5383, N5263);
nor NOR2 (N5390, N5389, N2159);
nand NAND4 (N5391, N5366, N4123, N493, N2962);
or OR4 (N5392, N5367, N2288, N4498, N2321);
nand NAND4 (N5393, N5392, N4445, N2133, N2007);
nor NOR2 (N5394, N5393, N1759);
xor XOR2 (N5395, N5394, N3514);
nand NAND2 (N5396, N5386, N2056);
xor XOR2 (N5397, N5378, N2588);
buf BUF1 (N5398, N5391);
and AND3 (N5399, N5398, N4385, N4454);
xor XOR2 (N5400, N5390, N247);
nor NOR4 (N5401, N5399, N1608, N2374, N3310);
buf BUF1 (N5402, N5381);
or OR4 (N5403, N5396, N3693, N403, N1557);
and AND3 (N5404, N5387, N2080, N1328);
nand NAND4 (N5405, N5375, N3635, N2739, N2602);
nand NAND2 (N5406, N5402, N3698);
or OR3 (N5407, N5395, N940, N1875);
buf BUF1 (N5408, N5407);
nor NOR2 (N5409, N5401, N3198);
xor XOR2 (N5410, N5408, N3879);
buf BUF1 (N5411, N5405);
or OR4 (N5412, N5409, N3761, N4417, N1338);
xor XOR2 (N5413, N5384, N5115);
not NOT1 (N5414, N5400);
and AND2 (N5415, N5410, N3444);
nand NAND2 (N5416, N5414, N3973);
nand NAND4 (N5417, N5406, N5162, N66, N1064);
buf BUF1 (N5418, N5417);
nand NAND2 (N5419, N5416, N2774);
and AND3 (N5420, N5404, N3600, N1594);
not NOT1 (N5421, N5415);
not NOT1 (N5422, N5403);
nand NAND4 (N5423, N5412, N3812, N2490, N3317);
and AND4 (N5424, N5411, N1147, N2084, N1511);
and AND3 (N5425, N5419, N1239, N622);
nand NAND2 (N5426, N5425, N2104);
xor XOR2 (N5427, N5420, N823);
not NOT1 (N5428, N5421);
not NOT1 (N5429, N5422);
nor NOR2 (N5430, N5388, N2501);
nor NOR3 (N5431, N5423, N4129, N2054);
or OR2 (N5432, N5431, N1490);
and AND4 (N5433, N5428, N2564, N709, N4781);
and AND2 (N5434, N5432, N2023);
xor XOR2 (N5435, N5427, N4762);
or OR2 (N5436, N5426, N2635);
and AND2 (N5437, N5413, N2792);
buf BUF1 (N5438, N5429);
buf BUF1 (N5439, N5430);
not NOT1 (N5440, N5437);
nor NOR3 (N5441, N5435, N4571, N4274);
nand NAND2 (N5442, N5397, N2741);
xor XOR2 (N5443, N5441, N2510);
or OR2 (N5444, N5439, N183);
buf BUF1 (N5445, N5442);
nor NOR4 (N5446, N5434, N1817, N3849, N27);
xor XOR2 (N5447, N5436, N3396);
buf BUF1 (N5448, N5424);
buf BUF1 (N5449, N5418);
and AND4 (N5450, N5447, N632, N3798, N1923);
nand NAND3 (N5451, N5446, N5168, N3993);
xor XOR2 (N5452, N5448, N2036);
buf BUF1 (N5453, N5438);
buf BUF1 (N5454, N5443);
nand NAND2 (N5455, N5440, N2819);
buf BUF1 (N5456, N5433);
buf BUF1 (N5457, N5449);
and AND2 (N5458, N5444, N206);
or OR3 (N5459, N5450, N3524, N3860);
or OR3 (N5460, N5451, N66, N4746);
not NOT1 (N5461, N5455);
nand NAND3 (N5462, N5459, N2194, N460);
nor NOR4 (N5463, N5458, N3145, N2339, N5155);
or OR4 (N5464, N5461, N2405, N1205, N781);
and AND3 (N5465, N5462, N416, N1519);
not NOT1 (N5466, N5454);
not NOT1 (N5467, N5464);
buf BUF1 (N5468, N5456);
and AND2 (N5469, N5452, N3574);
nand NAND2 (N5470, N5463, N192);
nand NAND4 (N5471, N5457, N5368, N4327, N3949);
xor XOR2 (N5472, N5466, N5266);
nand NAND4 (N5473, N5468, N4343, N721, N1666);
nand NAND2 (N5474, N5460, N5074);
nor NOR3 (N5475, N5465, N2060, N3541);
nor NOR3 (N5476, N5473, N4593, N3233);
and AND4 (N5477, N5453, N367, N2122, N489);
nand NAND3 (N5478, N5477, N906, N4732);
xor XOR2 (N5479, N5476, N1797);
nor NOR3 (N5480, N5474, N2785, N1518);
or OR3 (N5481, N5467, N464, N1131);
not NOT1 (N5482, N5471);
nand NAND3 (N5483, N5481, N1800, N4117);
or OR2 (N5484, N5470, N2162);
buf BUF1 (N5485, N5469);
or OR3 (N5486, N5475, N720, N1823);
and AND2 (N5487, N5479, N4100);
or OR4 (N5488, N5485, N300, N4383, N5355);
and AND4 (N5489, N5484, N5424, N5339, N2514);
and AND2 (N5490, N5488, N5169);
buf BUF1 (N5491, N5489);
or OR4 (N5492, N5483, N2871, N728, N4372);
nor NOR3 (N5493, N5482, N5481, N135);
not NOT1 (N5494, N5490);
nand NAND2 (N5495, N5486, N2319);
buf BUF1 (N5496, N5480);
buf BUF1 (N5497, N5487);
nand NAND4 (N5498, N5472, N3295, N666, N2106);
and AND3 (N5499, N5493, N1058, N4833);
buf BUF1 (N5500, N5495);
buf BUF1 (N5501, N5496);
buf BUF1 (N5502, N5445);
or OR3 (N5503, N5499, N4753, N4224);
nor NOR2 (N5504, N5501, N3268);
xor XOR2 (N5505, N5491, N3916);
nor NOR2 (N5506, N5502, N959);
buf BUF1 (N5507, N5504);
nand NAND3 (N5508, N5507, N4279, N4579);
nor NOR4 (N5509, N5505, N4414, N1491, N5235);
nand NAND4 (N5510, N5508, N366, N2011, N4099);
or OR4 (N5511, N5503, N4846, N2412, N2982);
not NOT1 (N5512, N5506);
nand NAND3 (N5513, N5509, N2699, N4809);
buf BUF1 (N5514, N5497);
not NOT1 (N5515, N5500);
xor XOR2 (N5516, N5511, N3518);
nand NAND2 (N5517, N5512, N1965);
nor NOR4 (N5518, N5510, N3191, N3642, N3582);
buf BUF1 (N5519, N5514);
buf BUF1 (N5520, N5513);
xor XOR2 (N5521, N5516, N3510);
xor XOR2 (N5522, N5494, N132);
nand NAND2 (N5523, N5519, N2398);
or OR4 (N5524, N5520, N4534, N3210, N1640);
not NOT1 (N5525, N5517);
and AND2 (N5526, N5524, N542);
and AND3 (N5527, N5523, N1414, N3380);
nor NOR3 (N5528, N5518, N4923, N603);
nor NOR4 (N5529, N5522, N1547, N4351, N4050);
and AND4 (N5530, N5492, N4749, N1412, N685);
nor NOR2 (N5531, N5515, N1550);
buf BUF1 (N5532, N5525);
not NOT1 (N5533, N5527);
not NOT1 (N5534, N5521);
not NOT1 (N5535, N5478);
xor XOR2 (N5536, N5498, N3948);
or OR4 (N5537, N5533, N902, N5000, N4457);
xor XOR2 (N5538, N5534, N673);
buf BUF1 (N5539, N5531);
xor XOR2 (N5540, N5530, N2396);
not NOT1 (N5541, N5537);
nand NAND2 (N5542, N5535, N375);
nor NOR2 (N5543, N5540, N3378);
or OR3 (N5544, N5539, N4590, N4157);
not NOT1 (N5545, N5536);
or OR4 (N5546, N5532, N4053, N2445, N3899);
nand NAND2 (N5547, N5543, N426);
nand NAND3 (N5548, N5542, N2942, N4844);
nand NAND3 (N5549, N5544, N2711, N1190);
and AND3 (N5550, N5545, N3919, N3788);
xor XOR2 (N5551, N5528, N1703);
not NOT1 (N5552, N5541);
not NOT1 (N5553, N5546);
nand NAND4 (N5554, N5547, N1448, N1177, N105);
not NOT1 (N5555, N5553);
or OR3 (N5556, N5550, N5441, N2302);
buf BUF1 (N5557, N5548);
nand NAND4 (N5558, N5557, N1114, N4427, N2127);
buf BUF1 (N5559, N5551);
buf BUF1 (N5560, N5555);
or OR4 (N5561, N5526, N5043, N1809, N5235);
xor XOR2 (N5562, N5559, N1520);
not NOT1 (N5563, N5529);
buf BUF1 (N5564, N5552);
and AND3 (N5565, N5554, N3518, N3418);
nand NAND2 (N5566, N5538, N2071);
not NOT1 (N5567, N5561);
nor NOR4 (N5568, N5567, N1927, N4081, N4369);
xor XOR2 (N5569, N5563, N2166);
nand NAND4 (N5570, N5562, N5459, N2266, N1762);
nor NOR3 (N5571, N5568, N4539, N4552);
nand NAND4 (N5572, N5570, N286, N2327, N3366);
nor NOR3 (N5573, N5566, N410, N4680);
buf BUF1 (N5574, N5564);
nand NAND4 (N5575, N5572, N4956, N2856, N1695);
or OR2 (N5576, N5549, N3086);
and AND3 (N5577, N5576, N4491, N1885);
nor NOR2 (N5578, N5577, N4735);
nand NAND2 (N5579, N5571, N1084);
or OR3 (N5580, N5574, N1636, N5356);
not NOT1 (N5581, N5573);
xor XOR2 (N5582, N5558, N5361);
xor XOR2 (N5583, N5575, N5524);
xor XOR2 (N5584, N5580, N490);
and AND3 (N5585, N5569, N4105, N5292);
or OR3 (N5586, N5579, N3473, N640);
or OR3 (N5587, N5578, N1412, N2969);
nor NOR2 (N5588, N5587, N306);
buf BUF1 (N5589, N5584);
nor NOR4 (N5590, N5583, N4567, N703, N5145);
not NOT1 (N5591, N5565);
not NOT1 (N5592, N5586);
xor XOR2 (N5593, N5581, N3297);
buf BUF1 (N5594, N5560);
and AND2 (N5595, N5592, N1338);
and AND4 (N5596, N5593, N3960, N2774, N883);
buf BUF1 (N5597, N5582);
nor NOR2 (N5598, N5594, N667);
and AND3 (N5599, N5590, N1575, N1880);
xor XOR2 (N5600, N5596, N2098);
buf BUF1 (N5601, N5597);
not NOT1 (N5602, N5595);
buf BUF1 (N5603, N5556);
nand NAND3 (N5604, N5589, N1358, N3780);
nor NOR2 (N5605, N5600, N510);
and AND3 (N5606, N5601, N4395, N1347);
not NOT1 (N5607, N5604);
or OR4 (N5608, N5598, N2599, N2063, N1391);
xor XOR2 (N5609, N5585, N4737);
and AND2 (N5610, N5602, N972);
and AND2 (N5611, N5605, N1301);
buf BUF1 (N5612, N5611);
nor NOR3 (N5613, N5610, N3559, N2282);
buf BUF1 (N5614, N5612);
nor NOR2 (N5615, N5606, N3723);
buf BUF1 (N5616, N5591);
and AND3 (N5617, N5613, N228, N4515);
xor XOR2 (N5618, N5588, N23);
or OR2 (N5619, N5608, N120);
xor XOR2 (N5620, N5616, N3693);
xor XOR2 (N5621, N5614, N2032);
xor XOR2 (N5622, N5617, N2731);
nor NOR2 (N5623, N5607, N3208);
and AND4 (N5624, N5615, N4120, N5173, N938);
or OR2 (N5625, N5622, N1909);
or OR3 (N5626, N5621, N176, N2280);
not NOT1 (N5627, N5619);
xor XOR2 (N5628, N5618, N5454);
nand NAND2 (N5629, N5627, N706);
not NOT1 (N5630, N5599);
buf BUF1 (N5631, N5603);
not NOT1 (N5632, N5623);
or OR4 (N5633, N5620, N3573, N5034, N4131);
not NOT1 (N5634, N5609);
nor NOR4 (N5635, N5630, N4793, N2989, N5332);
xor XOR2 (N5636, N5629, N1858);
nand NAND3 (N5637, N5633, N1601, N4209);
or OR2 (N5638, N5626, N1835);
buf BUF1 (N5639, N5631);
xor XOR2 (N5640, N5637, N436);
or OR2 (N5641, N5635, N2789);
buf BUF1 (N5642, N5624);
nand NAND3 (N5643, N5636, N5484, N5165);
nand NAND4 (N5644, N5639, N3617, N3575, N2285);
buf BUF1 (N5645, N5632);
and AND3 (N5646, N5638, N1337, N4817);
xor XOR2 (N5647, N5628, N496);
xor XOR2 (N5648, N5640, N3350);
not NOT1 (N5649, N5648);
xor XOR2 (N5650, N5641, N1895);
xor XOR2 (N5651, N5649, N2843);
nor NOR3 (N5652, N5634, N3779, N2882);
not NOT1 (N5653, N5645);
xor XOR2 (N5654, N5644, N3167);
buf BUF1 (N5655, N5653);
and AND4 (N5656, N5654, N851, N2595, N766);
not NOT1 (N5657, N5651);
nand NAND4 (N5658, N5656, N2820, N3494, N4728);
and AND3 (N5659, N5643, N139, N3363);
and AND4 (N5660, N5658, N5348, N1100, N839);
and AND2 (N5661, N5655, N2430);
or OR2 (N5662, N5650, N3446);
buf BUF1 (N5663, N5652);
xor XOR2 (N5664, N5642, N5546);
and AND4 (N5665, N5646, N3201, N1754, N5664);
nand NAND2 (N5666, N82, N240);
not NOT1 (N5667, N5663);
nand NAND4 (N5668, N5657, N3458, N1345, N4965);
not NOT1 (N5669, N5667);
or OR3 (N5670, N5669, N2013, N3071);
or OR3 (N5671, N5659, N1534, N4652);
xor XOR2 (N5672, N5662, N136);
not NOT1 (N5673, N5665);
not NOT1 (N5674, N5666);
nor NOR4 (N5675, N5625, N4606, N845, N4348);
buf BUF1 (N5676, N5675);
or OR2 (N5677, N5668, N3316);
xor XOR2 (N5678, N5673, N3423);
xor XOR2 (N5679, N5660, N1646);
and AND4 (N5680, N5674, N5176, N5280, N2446);
xor XOR2 (N5681, N5677, N4257);
buf BUF1 (N5682, N5678);
or OR3 (N5683, N5647, N3330, N440);
not NOT1 (N5684, N5681);
and AND2 (N5685, N5661, N4984);
or OR2 (N5686, N5685, N3344);
nor NOR3 (N5687, N5680, N2360, N1145);
nand NAND2 (N5688, N5671, N4177);
and AND4 (N5689, N5672, N5430, N898, N5461);
buf BUF1 (N5690, N5684);
not NOT1 (N5691, N5690);
or OR4 (N5692, N5689, N1384, N2013, N1218);
or OR3 (N5693, N5691, N5635, N1642);
nor NOR2 (N5694, N5693, N2831);
and AND3 (N5695, N5682, N3343, N5675);
buf BUF1 (N5696, N5692);
and AND2 (N5697, N5695, N3543);
nor NOR3 (N5698, N5683, N5231, N2462);
not NOT1 (N5699, N5670);
xor XOR2 (N5700, N5676, N3649);
and AND4 (N5701, N5686, N4321, N4494, N2823);
not NOT1 (N5702, N5687);
buf BUF1 (N5703, N5696);
or OR2 (N5704, N5679, N738);
not NOT1 (N5705, N5701);
not NOT1 (N5706, N5688);
or OR2 (N5707, N5703, N4374);
nand NAND2 (N5708, N5700, N5069);
xor XOR2 (N5709, N5705, N2377);
xor XOR2 (N5710, N5694, N4017);
not NOT1 (N5711, N5704);
buf BUF1 (N5712, N5698);
and AND3 (N5713, N5699, N2460, N4395);
nand NAND4 (N5714, N5697, N4166, N5592, N5372);
nand NAND3 (N5715, N5710, N2761, N5439);
buf BUF1 (N5716, N5712);
and AND4 (N5717, N5713, N1994, N3362, N906);
nor NOR3 (N5718, N5716, N499, N3230);
or OR4 (N5719, N5702, N4611, N4379, N4814);
and AND4 (N5720, N5718, N1602, N294, N4171);
or OR4 (N5721, N5719, N2559, N1, N3732);
nor NOR3 (N5722, N5711, N4900, N5597);
and AND4 (N5723, N5707, N2798, N1346, N1100);
or OR2 (N5724, N5717, N4372);
or OR4 (N5725, N5714, N1711, N5260, N4033);
not NOT1 (N5726, N5721);
nand NAND3 (N5727, N5720, N1881, N824);
xor XOR2 (N5728, N5726, N2232);
not NOT1 (N5729, N5728);
nand NAND3 (N5730, N5727, N2064, N4639);
nand NAND2 (N5731, N5729, N1184);
or OR3 (N5732, N5715, N4562, N1900);
buf BUF1 (N5733, N5722);
xor XOR2 (N5734, N5732, N2780);
or OR3 (N5735, N5708, N4540, N5194);
nor NOR3 (N5736, N5730, N1534, N4741);
not NOT1 (N5737, N5735);
nor NOR3 (N5738, N5724, N4376, N595);
and AND3 (N5739, N5738, N1843, N1932);
not NOT1 (N5740, N5723);
buf BUF1 (N5741, N5709);
or OR3 (N5742, N5739, N4234, N3674);
nand NAND4 (N5743, N5733, N2242, N1208, N3348);
and AND4 (N5744, N5743, N39, N3997, N2594);
buf BUF1 (N5745, N5737);
and AND3 (N5746, N5744, N989, N184);
and AND4 (N5747, N5741, N1186, N2179, N4065);
nand NAND2 (N5748, N5745, N4783);
not NOT1 (N5749, N5725);
or OR2 (N5750, N5706, N1413);
nor NOR4 (N5751, N5750, N4692, N302, N4355);
nor NOR3 (N5752, N5734, N1917, N2015);
xor XOR2 (N5753, N5736, N1795);
xor XOR2 (N5754, N5740, N1760);
and AND3 (N5755, N5742, N4821, N3185);
or OR2 (N5756, N5751, N2928);
not NOT1 (N5757, N5753);
buf BUF1 (N5758, N5752);
xor XOR2 (N5759, N5755, N1521);
buf BUF1 (N5760, N5731);
not NOT1 (N5761, N5760);
not NOT1 (N5762, N5759);
not NOT1 (N5763, N5762);
or OR4 (N5764, N5758, N3809, N4675, N2134);
not NOT1 (N5765, N5746);
and AND3 (N5766, N5748, N1793, N198);
and AND2 (N5767, N5764, N3485);
and AND3 (N5768, N5754, N1666, N3516);
not NOT1 (N5769, N5766);
not NOT1 (N5770, N5769);
xor XOR2 (N5771, N5747, N3170);
nand NAND3 (N5772, N5756, N2376, N5754);
buf BUF1 (N5773, N5770);
xor XOR2 (N5774, N5771, N1120);
buf BUF1 (N5775, N5761);
not NOT1 (N5776, N5765);
not NOT1 (N5777, N5763);
buf BUF1 (N5778, N5767);
or OR2 (N5779, N5773, N4090);
and AND2 (N5780, N5776, N4540);
nand NAND4 (N5781, N5757, N1095, N4426, N70);
nand NAND2 (N5782, N5777, N2604);
buf BUF1 (N5783, N5779);
buf BUF1 (N5784, N5749);
nand NAND4 (N5785, N5782, N2006, N3403, N13);
buf BUF1 (N5786, N5775);
nor NOR2 (N5787, N5784, N1575);
and AND3 (N5788, N5774, N677, N1849);
xor XOR2 (N5789, N5781, N1809);
nor NOR4 (N5790, N5772, N4143, N411, N655);
nand NAND4 (N5791, N5768, N3146, N141, N3935);
nor NOR3 (N5792, N5786, N5220, N5115);
nand NAND4 (N5793, N5791, N1935, N1968, N572);
buf BUF1 (N5794, N5790);
nor NOR4 (N5795, N5792, N526, N41, N1323);
or OR3 (N5796, N5778, N4389, N974);
buf BUF1 (N5797, N5789);
and AND2 (N5798, N5787, N5466);
xor XOR2 (N5799, N5783, N4731);
or OR3 (N5800, N5780, N5567, N3778);
nand NAND4 (N5801, N5797, N5509, N4308, N5109);
buf BUF1 (N5802, N5800);
and AND4 (N5803, N5793, N2279, N457, N199);
xor XOR2 (N5804, N5802, N1523);
and AND4 (N5805, N5804, N4735, N3424, N5279);
not NOT1 (N5806, N5801);
xor XOR2 (N5807, N5806, N707);
and AND3 (N5808, N5807, N374, N2112);
not NOT1 (N5809, N5794);
xor XOR2 (N5810, N5785, N1219);
xor XOR2 (N5811, N5803, N627);
and AND3 (N5812, N5805, N168, N3244);
or OR2 (N5813, N5799, N3690);
and AND2 (N5814, N5798, N5423);
buf BUF1 (N5815, N5810);
xor XOR2 (N5816, N5796, N1531);
nand NAND2 (N5817, N5808, N4204);
xor XOR2 (N5818, N5795, N183);
or OR2 (N5819, N5812, N2555);
not NOT1 (N5820, N5811);
buf BUF1 (N5821, N5819);
and AND4 (N5822, N5813, N4896, N2856, N4776);
not NOT1 (N5823, N5816);
not NOT1 (N5824, N5822);
buf BUF1 (N5825, N5824);
and AND2 (N5826, N5820, N4524);
or OR4 (N5827, N5825, N4945, N5305, N4431);
nor NOR4 (N5828, N5814, N1935, N1479, N4199);
xor XOR2 (N5829, N5809, N3892);
not NOT1 (N5830, N5788);
xor XOR2 (N5831, N5828, N143);
nor NOR2 (N5832, N5830, N1307);
xor XOR2 (N5833, N5831, N754);
xor XOR2 (N5834, N5829, N159);
nand NAND2 (N5835, N5834, N5286);
or OR3 (N5836, N5826, N4137, N2913);
xor XOR2 (N5837, N5832, N4769);
nand NAND4 (N5838, N5837, N887, N4810, N4951);
buf BUF1 (N5839, N5818);
xor XOR2 (N5840, N5835, N3542);
nand NAND3 (N5841, N5827, N5764, N1250);
or OR3 (N5842, N5838, N2825, N3783);
buf BUF1 (N5843, N5817);
nor NOR3 (N5844, N5815, N4756, N4986);
xor XOR2 (N5845, N5821, N507);
and AND3 (N5846, N5836, N5118, N2212);
buf BUF1 (N5847, N5845);
nand NAND4 (N5848, N5840, N1511, N977, N2684);
not NOT1 (N5849, N5848);
not NOT1 (N5850, N5846);
not NOT1 (N5851, N5847);
buf BUF1 (N5852, N5841);
or OR2 (N5853, N5823, N4388);
buf BUF1 (N5854, N5844);
and AND3 (N5855, N5839, N650, N5056);
or OR2 (N5856, N5842, N4123);
or OR4 (N5857, N5852, N5046, N4051, N3497);
and AND3 (N5858, N5850, N3377, N1153);
and AND4 (N5859, N5843, N5753, N2009, N787);
buf BUF1 (N5860, N5833);
xor XOR2 (N5861, N5860, N1940);
nor NOR3 (N5862, N5859, N654, N5482);
nand NAND4 (N5863, N5858, N407, N5722, N1537);
not NOT1 (N5864, N5861);
or OR2 (N5865, N5863, N749);
xor XOR2 (N5866, N5865, N3721);
and AND4 (N5867, N5854, N2973, N1475, N3143);
buf BUF1 (N5868, N5862);
or OR3 (N5869, N5868, N3536, N1978);
or OR4 (N5870, N5864, N4706, N4537, N4498);
nor NOR3 (N5871, N5851, N2889, N3865);
nand NAND4 (N5872, N5870, N834, N2710, N518);
not NOT1 (N5873, N5871);
nand NAND3 (N5874, N5857, N1741, N480);
nand NAND3 (N5875, N5867, N5335, N5414);
or OR3 (N5876, N5856, N5076, N1680);
not NOT1 (N5877, N5849);
or OR4 (N5878, N5866, N4678, N3058, N2191);
or OR2 (N5879, N5869, N402);
not NOT1 (N5880, N5875);
buf BUF1 (N5881, N5853);
or OR4 (N5882, N5876, N3600, N352, N2280);
buf BUF1 (N5883, N5877);
nor NOR2 (N5884, N5879, N4860);
and AND4 (N5885, N5878, N2555, N4558, N4070);
or OR4 (N5886, N5874, N4007, N4396, N5721);
buf BUF1 (N5887, N5886);
xor XOR2 (N5888, N5872, N654);
and AND3 (N5889, N5882, N3911, N4276);
nand NAND4 (N5890, N5883, N1923, N979, N2399);
nor NOR3 (N5891, N5890, N566, N116);
or OR2 (N5892, N5873, N4300);
and AND2 (N5893, N5892, N4114);
nand NAND4 (N5894, N5855, N4639, N1575, N5115);
nor NOR4 (N5895, N5894, N1418, N4567, N439);
xor XOR2 (N5896, N5881, N2737);
nor NOR3 (N5897, N5889, N5514, N603);
nand NAND4 (N5898, N5880, N5129, N5017, N5823);
and AND3 (N5899, N5898, N588, N3530);
buf BUF1 (N5900, N5884);
buf BUF1 (N5901, N5897);
not NOT1 (N5902, N5901);
xor XOR2 (N5903, N5885, N5885);
or OR2 (N5904, N5891, N2028);
nand NAND2 (N5905, N5887, N4590);
and AND3 (N5906, N5888, N1236, N326);
not NOT1 (N5907, N5895);
buf BUF1 (N5908, N5903);
or OR3 (N5909, N5902, N627, N1585);
nor NOR4 (N5910, N5906, N875, N5708, N3520);
and AND2 (N5911, N5905, N3599);
or OR2 (N5912, N5893, N4898);
nor NOR2 (N5913, N5904, N243);
buf BUF1 (N5914, N5911);
not NOT1 (N5915, N5900);
and AND4 (N5916, N5913, N5424, N4736, N4014);
not NOT1 (N5917, N5896);
xor XOR2 (N5918, N5914, N4222);
nor NOR2 (N5919, N5907, N602);
nand NAND3 (N5920, N5916, N5026, N3564);
or OR2 (N5921, N5909, N4104);
buf BUF1 (N5922, N5899);
and AND4 (N5923, N5921, N5191, N76, N541);
and AND2 (N5924, N5910, N2502);
not NOT1 (N5925, N5919);
nor NOR3 (N5926, N5912, N2714, N579);
not NOT1 (N5927, N5925);
nor NOR3 (N5928, N5922, N2401, N2846);
buf BUF1 (N5929, N5924);
nor NOR2 (N5930, N5915, N93);
and AND2 (N5931, N5928, N3983);
buf BUF1 (N5932, N5918);
not NOT1 (N5933, N5931);
nor NOR4 (N5934, N5908, N4242, N53, N2756);
nor NOR2 (N5935, N5933, N1707);
buf BUF1 (N5936, N5927);
nand NAND3 (N5937, N5926, N3436, N2798);
and AND3 (N5938, N5917, N691, N255);
or OR4 (N5939, N5932, N2642, N4477, N2809);
or OR3 (N5940, N5934, N5739, N5045);
buf BUF1 (N5941, N5935);
nand NAND3 (N5942, N5938, N1062, N618);
xor XOR2 (N5943, N5920, N2063);
and AND3 (N5944, N5942, N4003, N1142);
and AND2 (N5945, N5941, N2376);
and AND3 (N5946, N5923, N4186, N1196);
not NOT1 (N5947, N5944);
or OR2 (N5948, N5940, N5359);
nor NOR4 (N5949, N5943, N3335, N1299, N4384);
nor NOR3 (N5950, N5945, N5016, N494);
and AND3 (N5951, N5930, N4896, N4988);
xor XOR2 (N5952, N5948, N5806);
not NOT1 (N5953, N5946);
buf BUF1 (N5954, N5953);
xor XOR2 (N5955, N5950, N1625);
nand NAND3 (N5956, N5929, N3899, N3124);
not NOT1 (N5957, N5949);
not NOT1 (N5958, N5954);
buf BUF1 (N5959, N5957);
nand NAND2 (N5960, N5959, N3756);
nor NOR3 (N5961, N5955, N995, N420);
nor NOR4 (N5962, N5960, N482, N5786, N1330);
or OR2 (N5963, N5951, N2256);
and AND4 (N5964, N5937, N952, N3153, N468);
and AND4 (N5965, N5962, N1900, N700, N1221);
not NOT1 (N5966, N5964);
buf BUF1 (N5967, N5966);
nand NAND4 (N5968, N5967, N4999, N2671, N4407);
nand NAND2 (N5969, N5939, N4440);
and AND3 (N5970, N5968, N651, N2505);
nor NOR3 (N5971, N5952, N2359, N5128);
or OR2 (N5972, N5963, N958);
not NOT1 (N5973, N5956);
xor XOR2 (N5974, N5970, N3718);
or OR4 (N5975, N5971, N4757, N1911, N133);
xor XOR2 (N5976, N5972, N4620);
or OR3 (N5977, N5969, N2911, N5660);
xor XOR2 (N5978, N5965, N2491);
nand NAND3 (N5979, N5974, N3025, N5227);
xor XOR2 (N5980, N5961, N2173);
nand NAND4 (N5981, N5975, N4442, N3843, N3980);
nand NAND2 (N5982, N5936, N3325);
buf BUF1 (N5983, N5982);
or OR3 (N5984, N5978, N4259, N383);
nand NAND2 (N5985, N5984, N110);
or OR3 (N5986, N5977, N5765, N2233);
nand NAND4 (N5987, N5958, N3185, N4413, N4446);
and AND3 (N5988, N5985, N1359, N2786);
nor NOR4 (N5989, N5988, N4035, N4871, N4377);
and AND4 (N5990, N5947, N1777, N5492, N2939);
and AND3 (N5991, N5980, N1225, N419);
buf BUF1 (N5992, N5983);
not NOT1 (N5993, N5992);
and AND3 (N5994, N5989, N4229, N4808);
and AND4 (N5995, N5993, N4491, N45, N4500);
nand NAND2 (N5996, N5973, N658);
xor XOR2 (N5997, N5995, N4397);
nand NAND2 (N5998, N5996, N3204);
not NOT1 (N5999, N5981);
buf BUF1 (N6000, N5986);
xor XOR2 (N6001, N5997, N4913);
xor XOR2 (N6002, N6001, N1804);
nand NAND4 (N6003, N5976, N3808, N1049, N3885);
and AND3 (N6004, N6000, N5480, N513);
and AND3 (N6005, N5979, N31, N2858);
nand NAND4 (N6006, N5990, N3361, N5328, N928);
nor NOR3 (N6007, N5998, N1777, N2997);
nand NAND2 (N6008, N6007, N3025);
and AND4 (N6009, N6006, N2963, N3793, N3954);
or OR4 (N6010, N5991, N776, N4867, N1842);
buf BUF1 (N6011, N5987);
nand NAND3 (N6012, N6009, N5646, N5784);
and AND2 (N6013, N6002, N3810);
not NOT1 (N6014, N6010);
buf BUF1 (N6015, N6013);
or OR2 (N6016, N6015, N40);
buf BUF1 (N6017, N6008);
nand NAND4 (N6018, N6004, N763, N5715, N803);
buf BUF1 (N6019, N6017);
not NOT1 (N6020, N6019);
or OR4 (N6021, N5999, N192, N391, N2319);
and AND4 (N6022, N6012, N3418, N2896, N520);
and AND2 (N6023, N6021, N2520);
buf BUF1 (N6024, N6014);
buf BUF1 (N6025, N6003);
xor XOR2 (N6026, N6005, N4964);
buf BUF1 (N6027, N5994);
buf BUF1 (N6028, N6018);
nor NOR3 (N6029, N6016, N1170, N2097);
or OR2 (N6030, N6028, N613);
xor XOR2 (N6031, N6025, N2442);
nor NOR3 (N6032, N6026, N1983, N2083);
and AND4 (N6033, N6032, N4878, N5123, N806);
and AND2 (N6034, N6033, N3840);
xor XOR2 (N6035, N6024, N3978);
nor NOR3 (N6036, N6031, N1085, N3247);
and AND4 (N6037, N6023, N773, N3538, N2693);
and AND3 (N6038, N6020, N2045, N3771);
xor XOR2 (N6039, N6027, N4401);
not NOT1 (N6040, N6036);
not NOT1 (N6041, N6029);
or OR4 (N6042, N6038, N5954, N112, N1707);
or OR4 (N6043, N6022, N719, N1844, N102);
or OR3 (N6044, N6043, N3955, N2461);
nand NAND2 (N6045, N6042, N4241);
nand NAND4 (N6046, N6035, N4046, N515, N4909);
buf BUF1 (N6047, N6037);
nor NOR2 (N6048, N6034, N5880);
or OR4 (N6049, N6039, N2284, N200, N4964);
nand NAND2 (N6050, N6011, N1442);
not NOT1 (N6051, N6044);
not NOT1 (N6052, N6045);
or OR4 (N6053, N6049, N141, N2944, N3400);
nor NOR2 (N6054, N6050, N2121);
buf BUF1 (N6055, N6041);
xor XOR2 (N6056, N6048, N2349);
buf BUF1 (N6057, N6052);
or OR3 (N6058, N6056, N109, N4575);
xor XOR2 (N6059, N6053, N3571);
or OR4 (N6060, N6040, N3278, N1579, N5864);
nand NAND4 (N6061, N6054, N3727, N4775, N5298);
nor NOR2 (N6062, N6060, N4422);
xor XOR2 (N6063, N6062, N4201);
and AND4 (N6064, N6051, N743, N4384, N3126);
xor XOR2 (N6065, N6046, N476);
nand NAND3 (N6066, N6057, N790, N1980);
nor NOR3 (N6067, N6055, N238, N4750);
or OR4 (N6068, N6058, N3887, N1352, N68);
buf BUF1 (N6069, N6067);
nor NOR2 (N6070, N6047, N4821);
and AND3 (N6071, N6065, N5750, N1302);
or OR4 (N6072, N6069, N2478, N205, N510);
not NOT1 (N6073, N6063);
xor XOR2 (N6074, N6064, N5210);
not NOT1 (N6075, N6061);
nor NOR2 (N6076, N6073, N5094);
xor XOR2 (N6077, N6070, N3922);
not NOT1 (N6078, N6071);
and AND3 (N6079, N6075, N2292, N5187);
nand NAND2 (N6080, N6077, N4290);
xor XOR2 (N6081, N6080, N4563);
nor NOR3 (N6082, N6068, N857, N174);
or OR3 (N6083, N6078, N4222, N6041);
nand NAND3 (N6084, N6059, N4011, N700);
nor NOR3 (N6085, N6076, N3756, N4635);
and AND3 (N6086, N6085, N3367, N4007);
nand NAND2 (N6087, N6083, N1569);
nor NOR4 (N6088, N6030, N4156, N4058, N5894);
and AND3 (N6089, N6084, N3809, N2543);
buf BUF1 (N6090, N6087);
nor NOR3 (N6091, N6072, N5476, N3388);
nand NAND3 (N6092, N6082, N3223, N5862);
nand NAND4 (N6093, N6089, N2778, N2881, N4702);
or OR2 (N6094, N6081, N3599);
not NOT1 (N6095, N6091);
not NOT1 (N6096, N6088);
buf BUF1 (N6097, N6079);
not NOT1 (N6098, N6090);
or OR3 (N6099, N6097, N4300, N462);
not NOT1 (N6100, N6066);
and AND3 (N6101, N6093, N290, N1523);
and AND3 (N6102, N6074, N1897, N2802);
or OR4 (N6103, N6095, N258, N5180, N1201);
and AND3 (N6104, N6094, N930, N4816);
not NOT1 (N6105, N6098);
nor NOR2 (N6106, N6092, N5713);
or OR4 (N6107, N6103, N4001, N4555, N4889);
buf BUF1 (N6108, N6100);
nor NOR2 (N6109, N6104, N4416);
nand NAND4 (N6110, N6099, N637, N4017, N5464);
or OR2 (N6111, N6086, N4652);
or OR3 (N6112, N6108, N3487, N2732);
nand NAND4 (N6113, N6105, N4738, N3734, N3308);
and AND2 (N6114, N6111, N3168);
buf BUF1 (N6115, N6106);
buf BUF1 (N6116, N6096);
nor NOR3 (N6117, N6101, N4793, N221);
not NOT1 (N6118, N6117);
xor XOR2 (N6119, N6114, N2565);
not NOT1 (N6120, N6118);
and AND3 (N6121, N6120, N3959, N3295);
buf BUF1 (N6122, N6113);
or OR3 (N6123, N6102, N36, N137);
nand NAND4 (N6124, N6115, N406, N1372, N4223);
nand NAND4 (N6125, N6119, N4888, N863, N1563);
buf BUF1 (N6126, N6122);
nand NAND2 (N6127, N6123, N1924);
not NOT1 (N6128, N6107);
or OR2 (N6129, N6124, N1981);
and AND2 (N6130, N6125, N1267);
xor XOR2 (N6131, N6116, N524);
or OR2 (N6132, N6109, N1635);
and AND4 (N6133, N6110, N5287, N1192, N1069);
or OR4 (N6134, N6121, N2899, N385, N5993);
buf BUF1 (N6135, N6134);
buf BUF1 (N6136, N6130);
nand NAND2 (N6137, N6131, N2817);
not NOT1 (N6138, N6127);
or OR3 (N6139, N6136, N2664, N3919);
nor NOR2 (N6140, N6139, N2950);
xor XOR2 (N6141, N6133, N639);
or OR2 (N6142, N6128, N3683);
buf BUF1 (N6143, N6142);
buf BUF1 (N6144, N6126);
nand NAND4 (N6145, N6138, N3911, N3747, N2274);
not NOT1 (N6146, N6143);
nor NOR3 (N6147, N6137, N4495, N1720);
nor NOR3 (N6148, N6144, N2117, N643);
xor XOR2 (N6149, N6135, N5495);
buf BUF1 (N6150, N6147);
not NOT1 (N6151, N6148);
nand NAND4 (N6152, N6140, N4355, N5097, N4979);
not NOT1 (N6153, N6150);
or OR2 (N6154, N6129, N32);
or OR2 (N6155, N6152, N1686);
not NOT1 (N6156, N6154);
nor NOR2 (N6157, N6156, N3436);
xor XOR2 (N6158, N6151, N4716);
buf BUF1 (N6159, N6157);
not NOT1 (N6160, N6145);
or OR3 (N6161, N6158, N2105, N5954);
nor NOR4 (N6162, N6160, N4993, N945, N4895);
not NOT1 (N6163, N6149);
not NOT1 (N6164, N6155);
or OR4 (N6165, N6161, N2550, N4999, N4758);
xor XOR2 (N6166, N6153, N1698);
nor NOR3 (N6167, N6141, N5931, N2063);
or OR2 (N6168, N6167, N1339);
buf BUF1 (N6169, N6168);
buf BUF1 (N6170, N6166);
not NOT1 (N6171, N6159);
or OR2 (N6172, N6171, N4730);
not NOT1 (N6173, N6172);
nand NAND3 (N6174, N6165, N5446, N4504);
buf BUF1 (N6175, N6170);
buf BUF1 (N6176, N6162);
nand NAND2 (N6177, N6174, N4369);
xor XOR2 (N6178, N6112, N5714);
not NOT1 (N6179, N6169);
nor NOR3 (N6180, N6173, N760, N5263);
nand NAND2 (N6181, N6164, N2071);
nand NAND4 (N6182, N6132, N403, N4388, N3661);
nand NAND2 (N6183, N6146, N5192);
nand NAND2 (N6184, N6181, N4130);
nor NOR2 (N6185, N6176, N2713);
and AND3 (N6186, N6177, N1839, N3660);
buf BUF1 (N6187, N6179);
xor XOR2 (N6188, N6163, N3235);
and AND2 (N6189, N6182, N2608);
nand NAND3 (N6190, N6189, N1573, N4476);
buf BUF1 (N6191, N6190);
nand NAND2 (N6192, N6180, N4164);
nor NOR3 (N6193, N6188, N173, N26);
or OR3 (N6194, N6175, N4932, N1126);
xor XOR2 (N6195, N6192, N528);
xor XOR2 (N6196, N6185, N1916);
not NOT1 (N6197, N6186);
and AND3 (N6198, N6195, N3119, N4100);
or OR2 (N6199, N6194, N5610);
or OR2 (N6200, N6199, N2129);
and AND4 (N6201, N6196, N4203, N2443, N337);
nor NOR2 (N6202, N6198, N4559);
xor XOR2 (N6203, N6191, N1594);
nand NAND4 (N6204, N6183, N1249, N6162, N2754);
not NOT1 (N6205, N6187);
xor XOR2 (N6206, N6201, N2966);
xor XOR2 (N6207, N6197, N3203);
or OR4 (N6208, N6184, N641, N1411, N5551);
not NOT1 (N6209, N6205);
or OR3 (N6210, N6206, N5287, N619);
buf BUF1 (N6211, N6207);
nor NOR2 (N6212, N6178, N3265);
not NOT1 (N6213, N6193);
nor NOR4 (N6214, N6213, N3273, N4260, N1262);
xor XOR2 (N6215, N6212, N3585);
xor XOR2 (N6216, N6204, N4157);
not NOT1 (N6217, N6200);
nand NAND4 (N6218, N6209, N5723, N5326, N418);
or OR3 (N6219, N6211, N5646, N5773);
not NOT1 (N6220, N6216);
nor NOR2 (N6221, N6208, N320);
and AND4 (N6222, N6203, N4028, N2984, N1421);
buf BUF1 (N6223, N6210);
not NOT1 (N6224, N6220);
nor NOR2 (N6225, N6222, N1688);
buf BUF1 (N6226, N6224);
xor XOR2 (N6227, N6225, N4003);
not NOT1 (N6228, N6218);
nor NOR2 (N6229, N6215, N2839);
and AND4 (N6230, N6217, N4615, N3540, N3303);
xor XOR2 (N6231, N6227, N5996);
or OR3 (N6232, N6231, N1694, N5376);
nor NOR2 (N6233, N6232, N4201);
nor NOR4 (N6234, N6202, N5786, N6090, N6005);
or OR3 (N6235, N6221, N4760, N1594);
and AND2 (N6236, N6223, N2590);
buf BUF1 (N6237, N6234);
xor XOR2 (N6238, N6229, N2412);
buf BUF1 (N6239, N6230);
or OR2 (N6240, N6235, N1154);
nor NOR2 (N6241, N6214, N3568);
or OR4 (N6242, N6240, N1415, N1676, N5029);
or OR3 (N6243, N6226, N4196, N5115);
buf BUF1 (N6244, N6228);
buf BUF1 (N6245, N6239);
xor XOR2 (N6246, N6236, N3457);
buf BUF1 (N6247, N6243);
or OR2 (N6248, N6219, N545);
xor XOR2 (N6249, N6245, N3824);
and AND2 (N6250, N6246, N1922);
not NOT1 (N6251, N6242);
nor NOR3 (N6252, N6237, N3104, N2616);
xor XOR2 (N6253, N6249, N2100);
not NOT1 (N6254, N6247);
or OR3 (N6255, N6248, N4021, N4002);
or OR3 (N6256, N6244, N5793, N3834);
not NOT1 (N6257, N6253);
nor NOR4 (N6258, N6257, N4473, N624, N4066);
nor NOR2 (N6259, N6255, N2854);
buf BUF1 (N6260, N6251);
nor NOR2 (N6261, N6252, N4419);
nor NOR4 (N6262, N6238, N2192, N242, N536);
nand NAND3 (N6263, N6250, N2070, N2916);
not NOT1 (N6264, N6259);
nand NAND2 (N6265, N6262, N2757);
buf BUF1 (N6266, N6264);
or OR4 (N6267, N6241, N2399, N5703, N5501);
nor NOR4 (N6268, N6265, N5006, N5786, N800);
and AND4 (N6269, N6254, N409, N483, N4402);
not NOT1 (N6270, N6267);
buf BUF1 (N6271, N6261);
nor NOR3 (N6272, N6269, N1205, N3574);
and AND4 (N6273, N6260, N5804, N3617, N5676);
not NOT1 (N6274, N6273);
and AND4 (N6275, N6272, N5410, N3549, N525);
xor XOR2 (N6276, N6258, N5024);
not NOT1 (N6277, N6266);
not NOT1 (N6278, N6233);
nand NAND3 (N6279, N6274, N192, N6276);
xor XOR2 (N6280, N1225, N3017);
xor XOR2 (N6281, N6278, N1484);
xor XOR2 (N6282, N6275, N974);
not NOT1 (N6283, N6268);
buf BUF1 (N6284, N6282);
or OR4 (N6285, N6256, N5489, N4940, N5403);
buf BUF1 (N6286, N6263);
xor XOR2 (N6287, N6281, N5713);
or OR4 (N6288, N6287, N5871, N2095, N87);
nand NAND3 (N6289, N6280, N2709, N2779);
nor NOR2 (N6290, N6277, N207);
or OR3 (N6291, N6286, N2645, N5479);
and AND4 (N6292, N6283, N2172, N1604, N6016);
or OR3 (N6293, N6271, N2128, N2704);
nor NOR3 (N6294, N6289, N1649, N3745);
buf BUF1 (N6295, N6279);
or OR3 (N6296, N6284, N393, N2624);
xor XOR2 (N6297, N6293, N4993);
xor XOR2 (N6298, N6285, N5255);
buf BUF1 (N6299, N6290);
nand NAND4 (N6300, N6270, N872, N5307, N5514);
or OR4 (N6301, N6300, N3583, N3750, N6296);
nor NOR4 (N6302, N5402, N4018, N3114, N2554);
or OR2 (N6303, N6288, N889);
xor XOR2 (N6304, N6298, N4367);
nor NOR4 (N6305, N6297, N5384, N4166, N5307);
or OR3 (N6306, N6304, N1703, N2679);
nand NAND3 (N6307, N6302, N568, N2507);
not NOT1 (N6308, N6307);
nor NOR4 (N6309, N6299, N3416, N4761, N1497);
not NOT1 (N6310, N6303);
or OR2 (N6311, N6292, N4371);
or OR4 (N6312, N6311, N3280, N4953, N1482);
or OR3 (N6313, N6294, N1310, N4638);
nand NAND2 (N6314, N6306, N2746);
and AND4 (N6315, N6313, N212, N5846, N6098);
nand NAND2 (N6316, N6305, N3447);
nor NOR2 (N6317, N6291, N689);
nor NOR3 (N6318, N6312, N817, N1758);
not NOT1 (N6319, N6318);
nand NAND3 (N6320, N6315, N3347, N1069);
nand NAND4 (N6321, N6317, N5833, N4258, N1840);
xor XOR2 (N6322, N6321, N1179);
and AND2 (N6323, N6322, N398);
nand NAND2 (N6324, N6295, N3602);
or OR3 (N6325, N6323, N6015, N2251);
or OR2 (N6326, N6316, N828);
or OR3 (N6327, N6309, N918, N2853);
nor NOR3 (N6328, N6320, N1438, N4216);
or OR3 (N6329, N6308, N3205, N3285);
nand NAND4 (N6330, N6329, N93, N2605, N3653);
or OR3 (N6331, N6314, N4156, N516);
nor NOR2 (N6332, N6301, N4364);
nor NOR3 (N6333, N6324, N4221, N4197);
buf BUF1 (N6334, N6330);
nor NOR4 (N6335, N6333, N5844, N4244, N5247);
xor XOR2 (N6336, N6310, N2962);
xor XOR2 (N6337, N6319, N5964);
or OR4 (N6338, N6327, N2131, N4396, N4442);
or OR3 (N6339, N6337, N3707, N1642);
buf BUF1 (N6340, N6336);
xor XOR2 (N6341, N6335, N1318);
or OR4 (N6342, N6340, N4765, N1857, N1945);
not NOT1 (N6343, N6328);
not NOT1 (N6344, N6343);
buf BUF1 (N6345, N6332);
buf BUF1 (N6346, N6338);
not NOT1 (N6347, N6346);
not NOT1 (N6348, N6326);
xor XOR2 (N6349, N6344, N5216);
or OR4 (N6350, N6349, N6236, N2412, N6288);
buf BUF1 (N6351, N6345);
nand NAND4 (N6352, N6347, N5544, N2606, N4331);
buf BUF1 (N6353, N6325);
nand NAND4 (N6354, N6342, N5357, N2915, N2363);
buf BUF1 (N6355, N6351);
or OR3 (N6356, N6339, N1536, N3456);
xor XOR2 (N6357, N6355, N2002);
nand NAND2 (N6358, N6348, N1351);
buf BUF1 (N6359, N6354);
nor NOR2 (N6360, N6352, N485);
and AND4 (N6361, N6341, N5815, N1388, N2601);
buf BUF1 (N6362, N6353);
buf BUF1 (N6363, N6359);
buf BUF1 (N6364, N6363);
or OR4 (N6365, N6360, N1501, N3633, N468);
or OR4 (N6366, N6361, N1941, N1678, N4433);
xor XOR2 (N6367, N6350, N5289);
nor NOR2 (N6368, N6367, N1190);
nor NOR3 (N6369, N6365, N443, N293);
nand NAND3 (N6370, N6356, N186, N3343);
nor NOR2 (N6371, N6370, N663);
buf BUF1 (N6372, N6369);
not NOT1 (N6373, N6334);
and AND4 (N6374, N6331, N5154, N4327, N6229);
or OR4 (N6375, N6358, N3108, N1338, N2467);
or OR3 (N6376, N6368, N4432, N1014);
nor NOR2 (N6377, N6357, N4437);
or OR2 (N6378, N6366, N1745);
not NOT1 (N6379, N6375);
not NOT1 (N6380, N6372);
buf BUF1 (N6381, N6376);
nand NAND2 (N6382, N6364, N5903);
and AND4 (N6383, N6362, N2057, N3761, N1640);
xor XOR2 (N6384, N6381, N1055);
not NOT1 (N6385, N6382);
xor XOR2 (N6386, N6383, N440);
not NOT1 (N6387, N6380);
nor NOR2 (N6388, N6371, N5885);
not NOT1 (N6389, N6388);
buf BUF1 (N6390, N6377);
buf BUF1 (N6391, N6378);
not NOT1 (N6392, N6390);
and AND3 (N6393, N6384, N3744, N5347);
or OR4 (N6394, N6391, N2613, N4798, N2396);
and AND4 (N6395, N6373, N3076, N1719, N5527);
buf BUF1 (N6396, N6387);
or OR4 (N6397, N6385, N2015, N3754, N2709);
or OR2 (N6398, N6389, N4194);
buf BUF1 (N6399, N6374);
nor NOR2 (N6400, N6397, N4949);
not NOT1 (N6401, N6399);
and AND2 (N6402, N6400, N2518);
or OR3 (N6403, N6379, N407, N3397);
nand NAND3 (N6404, N6386, N895, N3800);
nor NOR4 (N6405, N6404, N6156, N5236, N5698);
buf BUF1 (N6406, N6398);
not NOT1 (N6407, N6403);
nor NOR2 (N6408, N6395, N5075);
or OR4 (N6409, N6405, N1679, N5644, N1885);
not NOT1 (N6410, N6401);
xor XOR2 (N6411, N6406, N3745);
xor XOR2 (N6412, N6411, N4610);
nand NAND2 (N6413, N6408, N4372);
nand NAND3 (N6414, N6412, N710, N4777);
or OR4 (N6415, N6409, N4682, N2632, N5167);
xor XOR2 (N6416, N6414, N5611);
nor NOR4 (N6417, N6394, N5966, N1665, N1179);
xor XOR2 (N6418, N6402, N4690);
and AND4 (N6419, N6417, N6196, N5945, N2675);
nand NAND3 (N6420, N6393, N5632, N3173);
not NOT1 (N6421, N6396);
nand NAND3 (N6422, N6418, N3824, N2934);
xor XOR2 (N6423, N6421, N6214);
nand NAND2 (N6424, N6416, N4438);
endmodule