// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11;

output N3009,N2969,N2954,N3003,N3001,N3002,N2985,N2999,N3006,N3011;

not NOT1 (N12, N5);
and AND3 (N13, N6, N5, N5);
nor NOR3 (N14, N9, N13, N6);
not NOT1 (N15, N2);
and AND2 (N16, N4, N11);
or OR3 (N17, N12, N4, N15);
nand NAND2 (N18, N13, N13);
buf BUF1 (N19, N6);
buf BUF1 (N20, N17);
or OR3 (N21, N18, N20, N4);
buf BUF1 (N22, N21);
buf BUF1 (N23, N7);
not NOT1 (N24, N4);
buf BUF1 (N25, N24);
and AND4 (N26, N13, N5, N19, N19);
or OR4 (N27, N24, N3, N2, N14);
nor NOR3 (N28, N13, N24, N27);
or OR2 (N29, N7, N25);
nand NAND3 (N30, N17, N15, N28);
xor XOR2 (N31, N28, N30);
not NOT1 (N32, N24);
or OR4 (N33, N8, N5, N29, N29);
nor NOR3 (N34, N17, N15, N5);
not NOT1 (N35, N5);
nand NAND2 (N36, N20, N16);
buf BUF1 (N37, N13);
not NOT1 (N38, N32);
nor NOR4 (N39, N23, N7, N22, N13);
and AND2 (N40, N37, N5);
buf BUF1 (N41, N36);
xor XOR2 (N42, N28, N19);
nand NAND2 (N43, N40, N42);
and AND2 (N44, N11, N20);
xor XOR2 (N45, N39, N6);
and AND2 (N46, N34, N25);
buf BUF1 (N47, N33);
or OR2 (N48, N44, N34);
or OR4 (N49, N26, N23, N33, N12);
buf BUF1 (N50, N47);
nand NAND4 (N51, N50, N20, N45, N11);
xor XOR2 (N52, N41, N30);
nor NOR4 (N53, N48, N22, N31, N40);
or OR4 (N54, N34, N13, N45, N49);
not NOT1 (N55, N43);
nor NOR3 (N56, N3, N24, N10);
nand NAND2 (N57, N15, N12);
buf BUF1 (N58, N56);
nor NOR3 (N59, N53, N14, N47);
xor XOR2 (N60, N58, N12);
xor XOR2 (N61, N57, N17);
or OR3 (N62, N55, N4, N29);
nor NOR2 (N63, N60, N2);
xor XOR2 (N64, N63, N30);
not NOT1 (N65, N59);
nand NAND2 (N66, N38, N32);
or OR4 (N67, N62, N17, N45, N52);
xor XOR2 (N68, N8, N27);
xor XOR2 (N69, N46, N20);
not NOT1 (N70, N67);
or OR4 (N71, N64, N2, N55, N23);
not NOT1 (N72, N35);
or OR2 (N73, N72, N25);
xor XOR2 (N74, N54, N46);
or OR4 (N75, N71, N29, N15, N38);
not NOT1 (N76, N69);
not NOT1 (N77, N51);
xor XOR2 (N78, N65, N46);
xor XOR2 (N79, N77, N2);
nand NAND4 (N80, N78, N12, N12, N12);
nor NOR3 (N81, N75, N77, N78);
not NOT1 (N82, N61);
nor NOR4 (N83, N79, N16, N27, N22);
and AND4 (N84, N82, N32, N22, N32);
nor NOR2 (N85, N74, N40);
xor XOR2 (N86, N81, N63);
and AND3 (N87, N76, N11, N50);
not NOT1 (N88, N85);
buf BUF1 (N89, N70);
buf BUF1 (N90, N66);
or OR4 (N91, N88, N6, N17, N52);
buf BUF1 (N92, N87);
xor XOR2 (N93, N68, N6);
not NOT1 (N94, N84);
nand NAND3 (N95, N89, N35, N82);
and AND4 (N96, N91, N3, N20, N83);
nand NAND2 (N97, N13, N57);
and AND2 (N98, N97, N50);
and AND2 (N99, N98, N48);
buf BUF1 (N100, N93);
and AND2 (N101, N92, N30);
nand NAND3 (N102, N101, N7, N77);
nor NOR3 (N103, N73, N98, N87);
or OR3 (N104, N102, N32, N79);
and AND3 (N105, N99, N32, N104);
nor NOR3 (N106, N43, N16, N54);
nor NOR2 (N107, N90, N36);
nand NAND2 (N108, N103, N23);
not NOT1 (N109, N105);
xor XOR2 (N110, N94, N99);
nor NOR2 (N111, N107, N96);
buf BUF1 (N112, N86);
nor NOR3 (N113, N61, N79, N70);
buf BUF1 (N114, N113);
xor XOR2 (N115, N95, N50);
and AND3 (N116, N108, N60, N12);
xor XOR2 (N117, N114, N34);
buf BUF1 (N118, N115);
or OR3 (N119, N117, N32, N96);
or OR4 (N120, N100, N16, N7, N62);
nor NOR4 (N121, N118, N17, N77, N27);
and AND4 (N122, N119, N81, N36, N83);
xor XOR2 (N123, N106, N58);
nand NAND2 (N124, N111, N49);
nand NAND4 (N125, N116, N79, N27, N103);
nor NOR3 (N126, N110, N37, N14);
buf BUF1 (N127, N120);
and AND2 (N128, N123, N37);
not NOT1 (N129, N112);
buf BUF1 (N130, N125);
buf BUF1 (N131, N130);
buf BUF1 (N132, N80);
xor XOR2 (N133, N131, N54);
buf BUF1 (N134, N121);
nor NOR2 (N135, N126, N72);
or OR3 (N136, N128, N73, N87);
xor XOR2 (N137, N127, N59);
buf BUF1 (N138, N135);
buf BUF1 (N139, N109);
or OR2 (N140, N129, N95);
and AND3 (N141, N140, N63, N136);
or OR2 (N142, N137, N76);
xor XOR2 (N143, N76, N79);
not NOT1 (N144, N141);
not NOT1 (N145, N124);
nor NOR3 (N146, N132, N55, N31);
buf BUF1 (N147, N144);
not NOT1 (N148, N139);
nand NAND2 (N149, N147, N128);
nor NOR2 (N150, N149, N133);
nand NAND3 (N151, N126, N61, N73);
xor XOR2 (N152, N138, N102);
and AND3 (N153, N143, N91, N6);
buf BUF1 (N154, N152);
not NOT1 (N155, N142);
buf BUF1 (N156, N146);
buf BUF1 (N157, N148);
or OR3 (N158, N151, N98, N113);
nand NAND2 (N159, N153, N48);
and AND4 (N160, N134, N87, N9, N33);
nand NAND4 (N161, N158, N4, N101, N141);
buf BUF1 (N162, N156);
nand NAND4 (N163, N154, N110, N58, N44);
buf BUF1 (N164, N122);
or OR2 (N165, N162, N134);
nand NAND3 (N166, N165, N165, N37);
buf BUF1 (N167, N150);
nand NAND2 (N168, N164, N83);
buf BUF1 (N169, N167);
or OR3 (N170, N166, N160, N139);
nor NOR3 (N171, N164, N36, N103);
buf BUF1 (N172, N169);
or OR3 (N173, N157, N32, N82);
nor NOR4 (N174, N155, N19, N90, N110);
nand NAND2 (N175, N159, N81);
nor NOR2 (N176, N171, N55);
and AND2 (N177, N170, N97);
nand NAND2 (N178, N177, N132);
nor NOR3 (N179, N172, N8, N8);
nand NAND3 (N180, N163, N164, N174);
nor NOR3 (N181, N172, N28, N13);
nand NAND3 (N182, N178, N113, N56);
not NOT1 (N183, N181);
and AND3 (N184, N180, N68, N35);
nand NAND2 (N185, N175, N113);
xor XOR2 (N186, N173, N176);
not NOT1 (N187, N182);
and AND4 (N188, N121, N28, N103, N89);
or OR2 (N189, N185, N185);
not NOT1 (N190, N161);
buf BUF1 (N191, N190);
or OR3 (N192, N145, N110, N142);
and AND2 (N193, N184, N11);
and AND4 (N194, N187, N118, N84, N28);
nand NAND3 (N195, N193, N165, N112);
and AND2 (N196, N194, N32);
or OR3 (N197, N196, N12, N42);
and AND3 (N198, N191, N155, N117);
buf BUF1 (N199, N189);
not NOT1 (N200, N195);
or OR2 (N201, N183, N77);
nor NOR4 (N202, N188, N38, N123, N87);
nor NOR2 (N203, N199, N45);
nor NOR4 (N204, N200, N166, N78, N83);
buf BUF1 (N205, N186);
and AND2 (N206, N202, N74);
nand NAND2 (N207, N192, N62);
nor NOR2 (N208, N207, N159);
buf BUF1 (N209, N179);
and AND2 (N210, N201, N28);
xor XOR2 (N211, N197, N180);
nor NOR4 (N212, N208, N54, N56, N15);
xor XOR2 (N213, N209, N104);
not NOT1 (N214, N203);
or OR3 (N215, N168, N60, N204);
buf BUF1 (N216, N44);
not NOT1 (N217, N198);
buf BUF1 (N218, N212);
and AND4 (N219, N214, N33, N158, N78);
buf BUF1 (N220, N211);
nor NOR3 (N221, N220, N193, N187);
and AND2 (N222, N219, N68);
xor XOR2 (N223, N210, N200);
nor NOR4 (N224, N213, N153, N46, N157);
or OR2 (N225, N221, N214);
not NOT1 (N226, N216);
xor XOR2 (N227, N217, N118);
and AND2 (N228, N223, N196);
or OR4 (N229, N206, N26, N47, N38);
or OR2 (N230, N226, N106);
buf BUF1 (N231, N229);
and AND3 (N232, N228, N14, N120);
or OR4 (N233, N232, N72, N95, N44);
or OR4 (N234, N222, N202, N15, N178);
buf BUF1 (N235, N234);
xor XOR2 (N236, N218, N121);
not NOT1 (N237, N225);
nand NAND4 (N238, N224, N207, N183, N11);
and AND2 (N239, N233, N226);
nand NAND4 (N240, N235, N122, N172, N91);
nand NAND2 (N241, N237, N158);
nand NAND3 (N242, N238, N84, N60);
or OR3 (N243, N215, N135, N163);
buf BUF1 (N244, N239);
buf BUF1 (N245, N243);
xor XOR2 (N246, N245, N38);
buf BUF1 (N247, N241);
not NOT1 (N248, N246);
nand NAND4 (N249, N227, N131, N157, N184);
buf BUF1 (N250, N244);
or OR4 (N251, N247, N178, N248, N178);
buf BUF1 (N252, N56);
not NOT1 (N253, N251);
not NOT1 (N254, N242);
nand NAND3 (N255, N236, N247, N1);
and AND4 (N256, N240, N181, N45, N210);
and AND4 (N257, N230, N130, N119, N233);
nand NAND3 (N258, N250, N224, N81);
xor XOR2 (N259, N205, N90);
not NOT1 (N260, N253);
xor XOR2 (N261, N257, N127);
nand NAND4 (N262, N258, N115, N79, N25);
or OR3 (N263, N261, N63, N155);
not NOT1 (N264, N262);
and AND3 (N265, N260, N179, N41);
and AND2 (N266, N255, N254);
nand NAND4 (N267, N134, N217, N149, N100);
nand NAND4 (N268, N256, N147, N241, N55);
not NOT1 (N269, N263);
nor NOR2 (N270, N269, N68);
nand NAND2 (N271, N267, N110);
buf BUF1 (N272, N271);
or OR2 (N273, N266, N89);
not NOT1 (N274, N264);
xor XOR2 (N275, N270, N84);
and AND4 (N276, N259, N124, N190, N87);
nand NAND2 (N277, N273, N138);
buf BUF1 (N278, N275);
not NOT1 (N279, N277);
and AND3 (N280, N268, N208, N178);
buf BUF1 (N281, N272);
nand NAND4 (N282, N278, N121, N35, N61);
not NOT1 (N283, N276);
nor NOR3 (N284, N280, N200, N267);
not NOT1 (N285, N274);
nor NOR2 (N286, N281, N41);
nand NAND2 (N287, N279, N19);
or OR3 (N288, N287, N188, N161);
not NOT1 (N289, N249);
and AND3 (N290, N252, N3, N187);
xor XOR2 (N291, N284, N242);
xor XOR2 (N292, N282, N34);
nand NAND3 (N293, N285, N146, N64);
nor NOR2 (N294, N288, N228);
buf BUF1 (N295, N283);
not NOT1 (N296, N292);
nor NOR4 (N297, N296, N180, N52, N240);
nand NAND2 (N298, N294, N112);
nand NAND3 (N299, N297, N62, N242);
nor NOR2 (N300, N295, N105);
or OR4 (N301, N291, N130, N125, N281);
nor NOR3 (N302, N290, N54, N44);
nand NAND3 (N303, N301, N19, N263);
nand NAND4 (N304, N303, N281, N32, N207);
xor XOR2 (N305, N265, N159);
nor NOR3 (N306, N300, N265, N116);
nor NOR4 (N307, N302, N165, N19, N108);
or OR4 (N308, N298, N191, N39, N198);
or OR4 (N309, N299, N244, N179, N12);
nand NAND3 (N310, N308, N150, N49);
not NOT1 (N311, N307);
nand NAND2 (N312, N289, N263);
buf BUF1 (N313, N309);
buf BUF1 (N314, N304);
or OR3 (N315, N286, N63, N107);
and AND4 (N316, N314, N117, N198, N222);
nor NOR3 (N317, N293, N305, N70);
and AND4 (N318, N182, N274, N312, N257);
nand NAND2 (N319, N58, N160);
or OR2 (N320, N306, N55);
nand NAND4 (N321, N320, N162, N172, N234);
nand NAND3 (N322, N319, N131, N121);
nor NOR4 (N323, N322, N311, N201, N251);
nand NAND3 (N324, N124, N253, N118);
nand NAND4 (N325, N318, N30, N290, N60);
nand NAND2 (N326, N323, N51);
nand NAND3 (N327, N310, N243, N116);
xor XOR2 (N328, N327, N230);
not NOT1 (N329, N315);
xor XOR2 (N330, N317, N49);
buf BUF1 (N331, N329);
nor NOR4 (N332, N328, N192, N282, N284);
buf BUF1 (N333, N331);
or OR2 (N334, N231, N125);
and AND2 (N335, N321, N19);
and AND2 (N336, N330, N37);
buf BUF1 (N337, N313);
nand NAND3 (N338, N334, N57, N14);
or OR3 (N339, N338, N244, N161);
and AND3 (N340, N333, N45, N78);
or OR3 (N341, N335, N332, N51);
nor NOR4 (N342, N226, N261, N102, N77);
or OR3 (N343, N337, N113, N129);
not NOT1 (N344, N340);
not NOT1 (N345, N325);
buf BUF1 (N346, N336);
or OR2 (N347, N344, N78);
and AND4 (N348, N345, N304, N81, N4);
nor NOR3 (N349, N324, N334, N312);
nor NOR2 (N350, N339, N309);
nand NAND2 (N351, N350, N81);
not NOT1 (N352, N316);
xor XOR2 (N353, N351, N213);
not NOT1 (N354, N342);
nor NOR3 (N355, N348, N145, N47);
not NOT1 (N356, N355);
not NOT1 (N357, N353);
and AND2 (N358, N357, N213);
nand NAND2 (N359, N343, N190);
or OR3 (N360, N359, N30, N168);
nor NOR2 (N361, N341, N312);
xor XOR2 (N362, N346, N356);
buf BUF1 (N363, N290);
or OR2 (N364, N347, N290);
or OR4 (N365, N358, N71, N227, N212);
and AND2 (N366, N349, N181);
or OR2 (N367, N365, N203);
xor XOR2 (N368, N352, N261);
nand NAND4 (N369, N354, N305, N79, N239);
nand NAND2 (N370, N364, N264);
xor XOR2 (N371, N366, N282);
and AND2 (N372, N360, N127);
or OR4 (N373, N363, N69, N300, N116);
buf BUF1 (N374, N369);
and AND2 (N375, N368, N361);
not NOT1 (N376, N225);
not NOT1 (N377, N375);
and AND4 (N378, N374, N48, N307, N314);
buf BUF1 (N379, N326);
not NOT1 (N380, N371);
xor XOR2 (N381, N376, N103);
and AND4 (N382, N378, N150, N207, N311);
or OR2 (N383, N372, N128);
or OR4 (N384, N377, N260, N103, N281);
nor NOR3 (N385, N382, N219, N104);
not NOT1 (N386, N362);
xor XOR2 (N387, N370, N262);
nand NAND2 (N388, N379, N163);
xor XOR2 (N389, N385, N148);
nor NOR3 (N390, N386, N260, N37);
xor XOR2 (N391, N388, N218);
not NOT1 (N392, N389);
nand NAND4 (N393, N381, N295, N388, N271);
buf BUF1 (N394, N387);
buf BUF1 (N395, N394);
buf BUF1 (N396, N391);
and AND4 (N397, N380, N70, N56, N115);
nand NAND3 (N398, N367, N246, N186);
nor NOR4 (N399, N383, N204, N66, N102);
nand NAND4 (N400, N384, N348, N88, N210);
xor XOR2 (N401, N400, N373);
and AND4 (N402, N6, N324, N261, N83);
xor XOR2 (N403, N399, N340);
or OR2 (N404, N402, N360);
not NOT1 (N405, N395);
buf BUF1 (N406, N392);
nor NOR4 (N407, N406, N131, N240, N79);
xor XOR2 (N408, N405, N17);
or OR4 (N409, N393, N280, N108, N288);
nand NAND4 (N410, N403, N223, N264, N122);
nor NOR3 (N411, N410, N311, N301);
nand NAND4 (N412, N401, N211, N91, N294);
and AND4 (N413, N407, N138, N409, N380);
not NOT1 (N414, N191);
nor NOR4 (N415, N404, N271, N84, N39);
nand NAND2 (N416, N411, N323);
nand NAND2 (N417, N415, N162);
or OR3 (N418, N390, N395, N174);
buf BUF1 (N419, N416);
nand NAND4 (N420, N414, N14, N264, N251);
not NOT1 (N421, N408);
xor XOR2 (N422, N412, N244);
nor NOR3 (N423, N413, N74, N320);
nand NAND3 (N424, N396, N162, N323);
xor XOR2 (N425, N398, N215);
buf BUF1 (N426, N419);
nor NOR3 (N427, N397, N417, N298);
nand NAND2 (N428, N280, N324);
xor XOR2 (N429, N418, N96);
or OR3 (N430, N425, N153, N67);
not NOT1 (N431, N422);
nor NOR4 (N432, N424, N331, N61, N271);
and AND4 (N433, N427, N72, N404, N398);
buf BUF1 (N434, N433);
or OR2 (N435, N432, N414);
and AND3 (N436, N428, N166, N267);
or OR3 (N437, N434, N235, N396);
nand NAND2 (N438, N431, N13);
or OR4 (N439, N421, N2, N211, N185);
and AND2 (N440, N423, N202);
nand NAND4 (N441, N438, N221, N283, N127);
or OR2 (N442, N436, N20);
xor XOR2 (N443, N442, N422);
nand NAND4 (N444, N430, N223, N69, N115);
buf BUF1 (N445, N444);
not NOT1 (N446, N429);
nor NOR3 (N447, N443, N130, N282);
nor NOR4 (N448, N440, N386, N92, N250);
xor XOR2 (N449, N435, N230);
nand NAND3 (N450, N448, N277, N90);
buf BUF1 (N451, N420);
xor XOR2 (N452, N426, N12);
nand NAND2 (N453, N450, N348);
nor NOR4 (N454, N437, N235, N376, N403);
and AND2 (N455, N449, N159);
and AND4 (N456, N453, N373, N454, N335);
and AND4 (N457, N174, N410, N340, N363);
nand NAND3 (N458, N445, N399, N148);
buf BUF1 (N459, N457);
xor XOR2 (N460, N452, N192);
nor NOR3 (N461, N456, N58, N459);
and AND3 (N462, N79, N209, N220);
and AND3 (N463, N455, N24, N345);
not NOT1 (N464, N463);
xor XOR2 (N465, N439, N156);
not NOT1 (N466, N462);
not NOT1 (N467, N441);
and AND4 (N468, N466, N384, N386, N144);
or OR3 (N469, N458, N451, N30);
xor XOR2 (N470, N365, N239);
or OR2 (N471, N465, N239);
xor XOR2 (N472, N447, N330);
not NOT1 (N473, N461);
not NOT1 (N474, N472);
or OR2 (N475, N474, N400);
xor XOR2 (N476, N464, N177);
or OR2 (N477, N470, N373);
not NOT1 (N478, N460);
and AND2 (N479, N469, N241);
buf BUF1 (N480, N476);
or OR4 (N481, N467, N369, N33, N410);
nand NAND3 (N482, N468, N280, N357);
not NOT1 (N483, N481);
buf BUF1 (N484, N482);
buf BUF1 (N485, N475);
nor NOR2 (N486, N471, N200);
nor NOR3 (N487, N483, N375, N425);
not NOT1 (N488, N484);
and AND2 (N489, N487, N481);
xor XOR2 (N490, N489, N114);
xor XOR2 (N491, N446, N277);
buf BUF1 (N492, N479);
or OR2 (N493, N486, N110);
or OR3 (N494, N480, N380, N97);
xor XOR2 (N495, N492, N410);
nor NOR3 (N496, N491, N425, N200);
nand NAND4 (N497, N485, N178, N103, N293);
xor XOR2 (N498, N473, N106);
and AND3 (N499, N495, N409, N168);
or OR2 (N500, N494, N231);
not NOT1 (N501, N488);
and AND2 (N502, N493, N42);
xor XOR2 (N503, N502, N502);
not NOT1 (N504, N498);
not NOT1 (N505, N478);
xor XOR2 (N506, N505, N499);
nand NAND4 (N507, N114, N282, N303, N72);
buf BUF1 (N508, N507);
or OR3 (N509, N504, N367, N427);
nor NOR3 (N510, N503, N290, N392);
nand NAND2 (N511, N496, N88);
xor XOR2 (N512, N497, N368);
buf BUF1 (N513, N506);
and AND4 (N514, N477, N279, N415, N246);
nor NOR2 (N515, N490, N440);
not NOT1 (N516, N512);
and AND2 (N517, N500, N397);
buf BUF1 (N518, N510);
not NOT1 (N519, N509);
nand NAND3 (N520, N515, N97, N425);
nand NAND2 (N521, N519, N275);
buf BUF1 (N522, N516);
and AND3 (N523, N522, N398, N502);
and AND4 (N524, N523, N231, N75, N161);
not NOT1 (N525, N513);
nor NOR2 (N526, N517, N350);
nand NAND2 (N527, N511, N232);
nor NOR3 (N528, N508, N178, N152);
xor XOR2 (N529, N526, N351);
and AND3 (N530, N529, N362, N207);
nor NOR4 (N531, N514, N35, N82, N30);
or OR2 (N532, N520, N513);
and AND3 (N533, N528, N155, N87);
nand NAND2 (N534, N532, N243);
or OR3 (N535, N533, N9, N351);
xor XOR2 (N536, N521, N197);
not NOT1 (N537, N531);
and AND2 (N538, N535, N113);
not NOT1 (N539, N530);
not NOT1 (N540, N524);
nand NAND2 (N541, N538, N291);
or OR2 (N542, N534, N228);
buf BUF1 (N543, N537);
xor XOR2 (N544, N542, N284);
xor XOR2 (N545, N541, N414);
nand NAND3 (N546, N525, N219, N168);
xor XOR2 (N547, N539, N273);
and AND2 (N548, N527, N184);
nor NOR2 (N549, N548, N179);
not NOT1 (N550, N543);
nor NOR4 (N551, N536, N240, N200, N481);
nor NOR4 (N552, N550, N181, N419, N374);
xor XOR2 (N553, N544, N190);
or OR3 (N554, N545, N269, N255);
buf BUF1 (N555, N553);
buf BUF1 (N556, N546);
buf BUF1 (N557, N556);
or OR4 (N558, N551, N361, N181, N532);
buf BUF1 (N559, N554);
or OR4 (N560, N558, N459, N279, N435);
xor XOR2 (N561, N518, N522);
xor XOR2 (N562, N552, N122);
and AND4 (N563, N501, N157, N344, N283);
or OR2 (N564, N561, N60);
nor NOR4 (N565, N562, N384, N373, N59);
not NOT1 (N566, N563);
nor NOR2 (N567, N559, N221);
not NOT1 (N568, N557);
nand NAND2 (N569, N560, N393);
or OR3 (N570, N567, N19, N484);
or OR4 (N571, N555, N73, N271, N443);
xor XOR2 (N572, N547, N494);
nand NAND2 (N573, N572, N199);
and AND3 (N574, N566, N350, N91);
not NOT1 (N575, N574);
not NOT1 (N576, N575);
xor XOR2 (N577, N571, N147);
or OR3 (N578, N568, N269, N79);
and AND3 (N579, N573, N282, N235);
xor XOR2 (N580, N577, N197);
nand NAND4 (N581, N570, N199, N51, N262);
buf BUF1 (N582, N580);
xor XOR2 (N583, N579, N163);
and AND4 (N584, N576, N361, N400, N98);
and AND3 (N585, N564, N251, N224);
not NOT1 (N586, N585);
and AND4 (N587, N565, N535, N464, N191);
or OR2 (N588, N582, N19);
buf BUF1 (N589, N588);
or OR3 (N590, N578, N102, N240);
nand NAND3 (N591, N581, N291, N311);
buf BUF1 (N592, N587);
xor XOR2 (N593, N591, N191);
nand NAND3 (N594, N593, N97, N108);
or OR3 (N595, N583, N513, N3);
and AND4 (N596, N592, N511, N557, N25);
and AND4 (N597, N549, N247, N551, N261);
and AND4 (N598, N540, N253, N552, N45);
not NOT1 (N599, N590);
and AND3 (N600, N586, N222, N435);
buf BUF1 (N601, N569);
nand NAND2 (N602, N596, N75);
nor NOR2 (N603, N601, N452);
xor XOR2 (N604, N603, N603);
or OR2 (N605, N604, N294);
buf BUF1 (N606, N595);
xor XOR2 (N607, N602, N307);
nor NOR3 (N608, N589, N133, N39);
and AND3 (N609, N599, N173, N543);
or OR3 (N610, N598, N266, N472);
xor XOR2 (N611, N600, N36);
nand NAND2 (N612, N584, N53);
nor NOR4 (N613, N612, N491, N191, N367);
nand NAND4 (N614, N608, N532, N55, N486);
buf BUF1 (N615, N611);
or OR2 (N616, N609, N119);
nor NOR2 (N617, N606, N364);
nand NAND4 (N618, N610, N375, N48, N273);
or OR3 (N619, N618, N127, N32);
nand NAND4 (N620, N619, N290, N262, N146);
nor NOR2 (N621, N617, N263);
xor XOR2 (N622, N605, N191);
or OR4 (N623, N607, N104, N113, N166);
xor XOR2 (N624, N613, N314);
nand NAND2 (N625, N616, N515);
xor XOR2 (N626, N625, N103);
or OR2 (N627, N597, N528);
or OR3 (N628, N627, N406, N497);
xor XOR2 (N629, N614, N295);
buf BUF1 (N630, N621);
not NOT1 (N631, N594);
nor NOR2 (N632, N626, N374);
nand NAND4 (N633, N622, N490, N494, N222);
buf BUF1 (N634, N630);
and AND2 (N635, N615, N511);
not NOT1 (N636, N632);
and AND3 (N637, N635, N234, N351);
not NOT1 (N638, N620);
buf BUF1 (N639, N623);
or OR4 (N640, N628, N1, N53, N368);
nor NOR4 (N641, N638, N172, N485, N536);
buf BUF1 (N642, N634);
xor XOR2 (N643, N637, N627);
not NOT1 (N644, N636);
or OR2 (N645, N633, N410);
not NOT1 (N646, N629);
or OR2 (N647, N631, N362);
nor NOR4 (N648, N646, N105, N83, N491);
buf BUF1 (N649, N642);
nor NOR4 (N650, N641, N299, N462, N303);
nand NAND2 (N651, N643, N316);
buf BUF1 (N652, N649);
xor XOR2 (N653, N650, N313);
nor NOR2 (N654, N651, N545);
nand NAND3 (N655, N654, N261, N487);
or OR4 (N656, N640, N125, N638, N320);
nand NAND4 (N657, N655, N253, N533, N618);
nor NOR2 (N658, N652, N377);
buf BUF1 (N659, N653);
nand NAND4 (N660, N648, N358, N119, N537);
nor NOR3 (N661, N656, N14, N101);
and AND2 (N662, N658, N17);
not NOT1 (N663, N661);
nor NOR2 (N664, N662, N206);
and AND3 (N665, N660, N568, N33);
and AND4 (N666, N663, N228, N562, N449);
nand NAND2 (N667, N647, N429);
or OR2 (N668, N664, N312);
nand NAND3 (N669, N639, N455, N170);
not NOT1 (N670, N666);
buf BUF1 (N671, N667);
not NOT1 (N672, N665);
or OR2 (N673, N657, N303);
buf BUF1 (N674, N645);
nand NAND2 (N675, N674, N89);
xor XOR2 (N676, N672, N130);
or OR3 (N677, N624, N217, N182);
nor NOR2 (N678, N675, N653);
not NOT1 (N679, N671);
xor XOR2 (N680, N669, N504);
nor NOR3 (N681, N677, N514, N646);
xor XOR2 (N682, N681, N470);
nand NAND3 (N683, N644, N260, N609);
buf BUF1 (N684, N683);
and AND4 (N685, N679, N118, N209, N189);
buf BUF1 (N686, N668);
or OR2 (N687, N685, N504);
nor NOR2 (N688, N686, N324);
not NOT1 (N689, N678);
xor XOR2 (N690, N689, N41);
or OR4 (N691, N680, N502, N606, N249);
buf BUF1 (N692, N684);
nor NOR4 (N693, N676, N474, N275, N281);
xor XOR2 (N694, N691, N419);
xor XOR2 (N695, N673, N236);
and AND3 (N696, N695, N198, N166);
nor NOR3 (N697, N659, N472, N412);
xor XOR2 (N698, N694, N258);
nor NOR2 (N699, N698, N75);
not NOT1 (N700, N688);
not NOT1 (N701, N682);
or OR4 (N702, N693, N272, N653, N586);
not NOT1 (N703, N696);
buf BUF1 (N704, N670);
nand NAND3 (N705, N690, N695, N122);
nand NAND4 (N706, N699, N571, N424, N323);
xor XOR2 (N707, N692, N25);
nand NAND4 (N708, N697, N34, N585, N695);
and AND3 (N709, N700, N455, N115);
or OR3 (N710, N706, N81, N369);
nand NAND2 (N711, N704, N321);
nor NOR2 (N712, N702, N118);
xor XOR2 (N713, N703, N415);
nand NAND3 (N714, N707, N646, N99);
xor XOR2 (N715, N705, N289);
not NOT1 (N716, N711);
or OR4 (N717, N710, N95, N329, N233);
xor XOR2 (N718, N713, N383);
and AND4 (N719, N717, N476, N656, N100);
or OR4 (N720, N701, N293, N644, N170);
buf BUF1 (N721, N708);
not NOT1 (N722, N714);
nor NOR4 (N723, N720, N14, N553, N576);
and AND4 (N724, N709, N332, N664, N269);
nor NOR4 (N725, N721, N44, N666, N307);
not NOT1 (N726, N712);
or OR4 (N727, N725, N200, N148, N54);
xor XOR2 (N728, N687, N718);
nand NAND3 (N729, N543, N251, N248);
or OR4 (N730, N724, N26, N274, N312);
or OR3 (N731, N722, N589, N352);
nand NAND4 (N732, N716, N526, N622, N560);
not NOT1 (N733, N732);
and AND3 (N734, N719, N397, N660);
nor NOR2 (N735, N733, N696);
buf BUF1 (N736, N730);
not NOT1 (N737, N728);
and AND4 (N738, N731, N650, N688, N512);
and AND4 (N739, N737, N486, N589, N440);
or OR2 (N740, N726, N142);
and AND3 (N741, N735, N391, N572);
and AND3 (N742, N736, N139, N411);
nor NOR4 (N743, N739, N110, N645, N506);
or OR3 (N744, N743, N4, N212);
buf BUF1 (N745, N742);
nand NAND2 (N746, N738, N86);
not NOT1 (N747, N741);
nand NAND3 (N748, N729, N424, N291);
buf BUF1 (N749, N715);
buf BUF1 (N750, N745);
xor XOR2 (N751, N748, N187);
nand NAND4 (N752, N727, N272, N358, N569);
nand NAND2 (N753, N723, N532);
xor XOR2 (N754, N740, N366);
and AND2 (N755, N753, N153);
nand NAND2 (N756, N747, N720);
xor XOR2 (N757, N756, N239);
buf BUF1 (N758, N734);
nand NAND4 (N759, N744, N107, N346, N731);
nor NOR3 (N760, N750, N423, N549);
not NOT1 (N761, N746);
nand NAND3 (N762, N759, N252, N393);
nor NOR4 (N763, N757, N604, N717, N627);
nor NOR3 (N764, N763, N756, N749);
or OR3 (N765, N543, N147, N324);
nand NAND2 (N766, N752, N626);
or OR4 (N767, N766, N1, N90, N514);
or OR4 (N768, N754, N615, N251, N25);
nand NAND3 (N769, N755, N41, N592);
and AND3 (N770, N762, N266, N375);
nor NOR3 (N771, N758, N300, N288);
or OR4 (N772, N760, N533, N79, N111);
not NOT1 (N773, N767);
or OR2 (N774, N771, N286);
xor XOR2 (N775, N769, N400);
buf BUF1 (N776, N764);
nor NOR4 (N777, N772, N531, N449, N606);
or OR3 (N778, N773, N197, N209);
buf BUF1 (N779, N778);
and AND4 (N780, N770, N358, N118, N272);
not NOT1 (N781, N768);
or OR3 (N782, N765, N349, N467);
and AND4 (N783, N781, N220, N120, N141);
xor XOR2 (N784, N779, N254);
nand NAND3 (N785, N776, N572, N319);
nor NOR3 (N786, N751, N763, N402);
not NOT1 (N787, N784);
and AND2 (N788, N786, N212);
nand NAND2 (N789, N775, N620);
not NOT1 (N790, N787);
not NOT1 (N791, N782);
nand NAND4 (N792, N761, N116, N14, N523);
buf BUF1 (N793, N777);
xor XOR2 (N794, N788, N693);
nand NAND3 (N795, N774, N705, N369);
nand NAND2 (N796, N794, N511);
and AND2 (N797, N785, N185);
buf BUF1 (N798, N793);
xor XOR2 (N799, N796, N126);
nand NAND4 (N800, N783, N598, N309, N580);
or OR3 (N801, N799, N83, N359);
not NOT1 (N802, N780);
xor XOR2 (N803, N798, N60);
buf BUF1 (N804, N789);
not NOT1 (N805, N800);
buf BUF1 (N806, N797);
not NOT1 (N807, N792);
not NOT1 (N808, N795);
and AND4 (N809, N808, N247, N707, N677);
nor NOR3 (N810, N802, N529, N240);
nand NAND2 (N811, N790, N122);
buf BUF1 (N812, N809);
xor XOR2 (N813, N801, N566);
nand NAND2 (N814, N806, N215);
nor NOR3 (N815, N804, N196, N596);
not NOT1 (N816, N812);
or OR3 (N817, N813, N481, N518);
or OR4 (N818, N807, N482, N577, N98);
or OR3 (N819, N805, N687, N526);
nand NAND2 (N820, N811, N233);
not NOT1 (N821, N814);
or OR3 (N822, N817, N120, N579);
not NOT1 (N823, N816);
or OR3 (N824, N819, N114, N695);
and AND3 (N825, N815, N89, N186);
nor NOR3 (N826, N810, N691, N439);
and AND4 (N827, N824, N577, N380, N591);
nand NAND2 (N828, N822, N763);
not NOT1 (N829, N791);
nand NAND3 (N830, N828, N280, N401);
not NOT1 (N831, N818);
nand NAND4 (N832, N825, N570, N731, N337);
and AND2 (N833, N831, N427);
and AND2 (N834, N823, N152);
or OR4 (N835, N803, N144, N350, N651);
xor XOR2 (N836, N835, N46);
and AND4 (N837, N826, N762, N10, N90);
and AND3 (N838, N827, N528, N290);
nand NAND3 (N839, N833, N184, N84);
nand NAND2 (N840, N820, N499);
buf BUF1 (N841, N840);
buf BUF1 (N842, N838);
nor NOR4 (N843, N832, N751, N820, N803);
buf BUF1 (N844, N837);
nor NOR3 (N845, N830, N672, N230);
nand NAND2 (N846, N839, N685);
nor NOR3 (N847, N841, N836, N275);
xor XOR2 (N848, N363, N559);
and AND4 (N849, N829, N601, N561, N369);
and AND2 (N850, N849, N55);
buf BUF1 (N851, N843);
nand NAND2 (N852, N844, N330);
nand NAND3 (N853, N842, N552, N792);
buf BUF1 (N854, N845);
buf BUF1 (N855, N848);
not NOT1 (N856, N850);
nand NAND4 (N857, N821, N282, N852, N670);
nor NOR4 (N858, N229, N659, N403, N532);
or OR4 (N859, N846, N699, N510, N90);
nor NOR2 (N860, N856, N562);
or OR3 (N861, N834, N850, N220);
nor NOR4 (N862, N857, N473, N748, N68);
and AND2 (N863, N861, N631);
xor XOR2 (N864, N853, N596);
buf BUF1 (N865, N855);
xor XOR2 (N866, N854, N790);
or OR3 (N867, N847, N776, N431);
nor NOR4 (N868, N866, N154, N799, N832);
not NOT1 (N869, N851);
buf BUF1 (N870, N869);
xor XOR2 (N871, N862, N361);
nand NAND2 (N872, N867, N460);
nand NAND2 (N873, N865, N309);
and AND2 (N874, N873, N263);
not NOT1 (N875, N871);
and AND4 (N876, N864, N222, N495, N176);
not NOT1 (N877, N872);
nor NOR4 (N878, N868, N50, N459, N292);
or OR4 (N879, N863, N407, N458, N165);
and AND2 (N880, N870, N163);
xor XOR2 (N881, N874, N138);
not NOT1 (N882, N876);
buf BUF1 (N883, N879);
and AND4 (N884, N882, N640, N649, N520);
nor NOR3 (N885, N877, N309, N443);
xor XOR2 (N886, N878, N584);
not NOT1 (N887, N880);
nor NOR3 (N888, N881, N856, N361);
nor NOR2 (N889, N859, N752);
and AND2 (N890, N888, N351);
xor XOR2 (N891, N886, N730);
not NOT1 (N892, N884);
buf BUF1 (N893, N885);
not NOT1 (N894, N891);
or OR4 (N895, N887, N178, N817, N512);
xor XOR2 (N896, N895, N518);
xor XOR2 (N897, N883, N694);
nand NAND2 (N898, N897, N728);
xor XOR2 (N899, N875, N877);
not NOT1 (N900, N894);
xor XOR2 (N901, N893, N482);
xor XOR2 (N902, N898, N348);
and AND2 (N903, N892, N353);
xor XOR2 (N904, N900, N674);
nor NOR2 (N905, N860, N694);
nor NOR2 (N906, N905, N100);
nand NAND2 (N907, N899, N132);
and AND2 (N908, N903, N178);
not NOT1 (N909, N907);
and AND3 (N910, N890, N573, N76);
and AND3 (N911, N909, N470, N868);
xor XOR2 (N912, N910, N257);
buf BUF1 (N913, N911);
nor NOR4 (N914, N912, N732, N171, N322);
and AND4 (N915, N904, N80, N711, N612);
or OR4 (N916, N914, N834, N638, N771);
xor XOR2 (N917, N908, N342);
xor XOR2 (N918, N858, N764);
xor XOR2 (N919, N902, N333);
buf BUF1 (N920, N918);
xor XOR2 (N921, N915, N147);
xor XOR2 (N922, N889, N593);
nand NAND3 (N923, N919, N201, N27);
xor XOR2 (N924, N916, N334);
nor NOR4 (N925, N906, N104, N96, N374);
and AND3 (N926, N896, N378, N630);
nand NAND4 (N927, N922, N365, N891, N258);
or OR4 (N928, N901, N342, N182, N710);
xor XOR2 (N929, N921, N198);
and AND2 (N930, N920, N427);
not NOT1 (N931, N930);
not NOT1 (N932, N925);
nor NOR3 (N933, N923, N216, N531);
nand NAND4 (N934, N928, N89, N770, N664);
nor NOR2 (N935, N932, N869);
nand NAND4 (N936, N931, N496, N55, N527);
nand NAND4 (N937, N926, N118, N641, N205);
xor XOR2 (N938, N927, N618);
xor XOR2 (N939, N935, N404);
not NOT1 (N940, N917);
not NOT1 (N941, N924);
buf BUF1 (N942, N934);
buf BUF1 (N943, N933);
nor NOR3 (N944, N940, N68, N406);
nor NOR2 (N945, N939, N828);
buf BUF1 (N946, N943);
or OR3 (N947, N945, N773, N639);
nor NOR3 (N948, N941, N915, N212);
and AND3 (N949, N946, N505, N697);
and AND3 (N950, N938, N849, N32);
or OR2 (N951, N942, N249);
nor NOR4 (N952, N949, N535, N397, N670);
nor NOR3 (N953, N948, N453, N546);
or OR4 (N954, N947, N541, N142, N907);
nor NOR3 (N955, N936, N870, N812);
xor XOR2 (N956, N952, N338);
or OR3 (N957, N954, N301, N937);
and AND2 (N958, N795, N908);
nand NAND4 (N959, N929, N46, N535, N449);
not NOT1 (N960, N958);
nand NAND4 (N961, N944, N56, N692, N384);
and AND4 (N962, N955, N251, N680, N224);
and AND4 (N963, N961, N622, N396, N105);
and AND2 (N964, N960, N523);
or OR3 (N965, N913, N893, N271);
xor XOR2 (N966, N964, N634);
buf BUF1 (N967, N965);
or OR4 (N968, N956, N759, N549, N206);
or OR3 (N969, N967, N160, N35);
not NOT1 (N970, N968);
or OR2 (N971, N957, N869);
and AND2 (N972, N966, N91);
or OR3 (N973, N950, N722, N726);
nor NOR2 (N974, N972, N331);
xor XOR2 (N975, N973, N291);
nor NOR3 (N976, N969, N952, N939);
nor NOR2 (N977, N976, N757);
buf BUF1 (N978, N951);
or OR3 (N979, N959, N364, N296);
not NOT1 (N980, N963);
nand NAND4 (N981, N978, N109, N778, N278);
nand NAND4 (N982, N979, N321, N905, N547);
buf BUF1 (N983, N971);
buf BUF1 (N984, N982);
nand NAND3 (N985, N977, N139, N395);
and AND2 (N986, N953, N303);
buf BUF1 (N987, N975);
not NOT1 (N988, N983);
buf BUF1 (N989, N986);
nand NAND2 (N990, N985, N924);
or OR3 (N991, N987, N484, N676);
nand NAND4 (N992, N984, N206, N53, N392);
and AND2 (N993, N980, N266);
nand NAND3 (N994, N990, N121, N226);
nor NOR4 (N995, N992, N709, N208, N6);
not NOT1 (N996, N988);
not NOT1 (N997, N974);
or OR3 (N998, N991, N915, N681);
and AND3 (N999, N995, N283, N237);
or OR4 (N1000, N996, N249, N414, N301);
and AND3 (N1001, N994, N792, N783);
xor XOR2 (N1002, N1001, N145);
not NOT1 (N1003, N981);
buf BUF1 (N1004, N997);
not NOT1 (N1005, N993);
or OR3 (N1006, N998, N522, N77);
nand NAND3 (N1007, N970, N454, N284);
buf BUF1 (N1008, N1005);
xor XOR2 (N1009, N989, N1);
not NOT1 (N1010, N1007);
not NOT1 (N1011, N999);
buf BUF1 (N1012, N1000);
buf BUF1 (N1013, N1011);
nor NOR4 (N1014, N1006, N619, N954, N779);
or OR4 (N1015, N1004, N737, N877, N940);
not NOT1 (N1016, N1013);
or OR4 (N1017, N1002, N129, N890, N62);
nand NAND3 (N1018, N1003, N1006, N777);
or OR3 (N1019, N1008, N250, N722);
or OR3 (N1020, N1018, N621, N161);
buf BUF1 (N1021, N1020);
xor XOR2 (N1022, N1021, N753);
xor XOR2 (N1023, N1014, N607);
nand NAND3 (N1024, N1009, N609, N58);
nor NOR2 (N1025, N1015, N784);
and AND3 (N1026, N1010, N921, N427);
buf BUF1 (N1027, N1017);
or OR2 (N1028, N962, N555);
and AND4 (N1029, N1022, N664, N418, N42);
nor NOR3 (N1030, N1025, N541, N807);
buf BUF1 (N1031, N1016);
or OR4 (N1032, N1029, N882, N111, N590);
and AND4 (N1033, N1023, N268, N95, N891);
nor NOR4 (N1034, N1019, N292, N79, N189);
xor XOR2 (N1035, N1026, N978);
buf BUF1 (N1036, N1024);
nand NAND3 (N1037, N1028, N849, N669);
buf BUF1 (N1038, N1037);
nor NOR3 (N1039, N1034, N22, N253);
nand NAND4 (N1040, N1036, N623, N563, N532);
nor NOR3 (N1041, N1031, N84, N237);
not NOT1 (N1042, N1041);
or OR2 (N1043, N1038, N568);
nand NAND4 (N1044, N1027, N973, N230, N519);
and AND3 (N1045, N1033, N264, N85);
and AND2 (N1046, N1035, N445);
not NOT1 (N1047, N1046);
nand NAND3 (N1048, N1039, N388, N1006);
xor XOR2 (N1049, N1048, N785);
not NOT1 (N1050, N1042);
and AND3 (N1051, N1040, N413, N542);
not NOT1 (N1052, N1045);
nand NAND4 (N1053, N1049, N333, N29, N11);
nand NAND4 (N1054, N1043, N1003, N903, N882);
and AND3 (N1055, N1050, N188, N351);
not NOT1 (N1056, N1044);
xor XOR2 (N1057, N1056, N904);
and AND3 (N1058, N1032, N210, N103);
not NOT1 (N1059, N1053);
or OR2 (N1060, N1012, N687);
not NOT1 (N1061, N1052);
not NOT1 (N1062, N1057);
nor NOR2 (N1063, N1054, N440);
and AND3 (N1064, N1063, N1051, N718);
xor XOR2 (N1065, N2, N380);
xor XOR2 (N1066, N1064, N22);
xor XOR2 (N1067, N1062, N297);
nor NOR3 (N1068, N1058, N685, N571);
nor NOR3 (N1069, N1066, N634, N514);
or OR2 (N1070, N1068, N1026);
nor NOR2 (N1071, N1055, N821);
nand NAND3 (N1072, N1059, N878, N286);
and AND2 (N1073, N1061, N802);
not NOT1 (N1074, N1065);
and AND3 (N1075, N1072, N745, N936);
or OR2 (N1076, N1060, N462);
buf BUF1 (N1077, N1074);
buf BUF1 (N1078, N1067);
xor XOR2 (N1079, N1071, N548);
nor NOR2 (N1080, N1078, N392);
nor NOR3 (N1081, N1073, N59, N98);
nor NOR4 (N1082, N1075, N667, N590, N584);
or OR2 (N1083, N1082, N368);
or OR4 (N1084, N1047, N665, N416, N702);
nand NAND2 (N1085, N1083, N195);
and AND4 (N1086, N1030, N925, N470, N424);
xor XOR2 (N1087, N1081, N189);
or OR2 (N1088, N1086, N619);
nand NAND3 (N1089, N1080, N1032, N342);
and AND2 (N1090, N1088, N792);
nor NOR2 (N1091, N1084, N612);
xor XOR2 (N1092, N1091, N131);
nand NAND4 (N1093, N1076, N782, N490, N437);
buf BUF1 (N1094, N1077);
and AND4 (N1095, N1093, N668, N519, N78);
and AND3 (N1096, N1089, N21, N327);
nand NAND4 (N1097, N1070, N945, N245, N505);
or OR2 (N1098, N1087, N538);
or OR3 (N1099, N1090, N142, N897);
nand NAND4 (N1100, N1092, N943, N842, N326);
and AND3 (N1101, N1097, N603, N770);
not NOT1 (N1102, N1069);
and AND4 (N1103, N1094, N599, N174, N485);
not NOT1 (N1104, N1095);
nand NAND4 (N1105, N1103, N1099, N860, N802);
nor NOR2 (N1106, N950, N887);
xor XOR2 (N1107, N1079, N29);
nand NAND3 (N1108, N1098, N121, N11);
xor XOR2 (N1109, N1101, N1103);
buf BUF1 (N1110, N1085);
not NOT1 (N1111, N1108);
buf BUF1 (N1112, N1105);
buf BUF1 (N1113, N1096);
buf BUF1 (N1114, N1109);
and AND4 (N1115, N1106, N766, N44, N678);
nor NOR3 (N1116, N1111, N146, N1084);
nand NAND2 (N1117, N1104, N38);
and AND3 (N1118, N1110, N989, N74);
and AND4 (N1119, N1114, N1019, N146, N278);
nor NOR4 (N1120, N1118, N473, N785, N1072);
nand NAND2 (N1121, N1115, N508);
nand NAND3 (N1122, N1116, N877, N764);
nand NAND3 (N1123, N1100, N33, N848);
or OR4 (N1124, N1113, N684, N859, N932);
or OR2 (N1125, N1120, N214);
xor XOR2 (N1126, N1117, N969);
and AND3 (N1127, N1107, N111, N245);
xor XOR2 (N1128, N1122, N939);
not NOT1 (N1129, N1128);
or OR3 (N1130, N1129, N154, N905);
nand NAND4 (N1131, N1125, N380, N930, N369);
xor XOR2 (N1132, N1127, N992);
nand NAND3 (N1133, N1131, N404, N991);
or OR2 (N1134, N1102, N447);
not NOT1 (N1135, N1119);
xor XOR2 (N1136, N1135, N984);
xor XOR2 (N1137, N1124, N1076);
or OR2 (N1138, N1137, N551);
and AND3 (N1139, N1126, N611, N570);
nand NAND4 (N1140, N1136, N259, N823, N977);
or OR2 (N1141, N1138, N888);
xor XOR2 (N1142, N1139, N888);
buf BUF1 (N1143, N1123);
buf BUF1 (N1144, N1142);
xor XOR2 (N1145, N1141, N901);
xor XOR2 (N1146, N1143, N469);
xor XOR2 (N1147, N1132, N206);
not NOT1 (N1148, N1121);
buf BUF1 (N1149, N1133);
and AND4 (N1150, N1112, N777, N3, N669);
xor XOR2 (N1151, N1150, N579);
buf BUF1 (N1152, N1140);
or OR3 (N1153, N1130, N329, N932);
or OR3 (N1154, N1144, N718, N772);
and AND2 (N1155, N1145, N1077);
nand NAND3 (N1156, N1154, N427, N752);
nand NAND4 (N1157, N1147, N451, N325, N1028);
and AND3 (N1158, N1153, N942, N394);
and AND3 (N1159, N1146, N1154, N542);
or OR3 (N1160, N1134, N694, N160);
xor XOR2 (N1161, N1158, N408);
nand NAND4 (N1162, N1152, N850, N285, N108);
or OR2 (N1163, N1148, N778);
or OR2 (N1164, N1157, N464);
or OR2 (N1165, N1155, N434);
not NOT1 (N1166, N1149);
nand NAND4 (N1167, N1156, N408, N121, N745);
or OR2 (N1168, N1164, N12);
buf BUF1 (N1169, N1168);
xor XOR2 (N1170, N1162, N56);
or OR4 (N1171, N1161, N508, N679, N995);
or OR3 (N1172, N1170, N241, N649);
nand NAND4 (N1173, N1159, N254, N953, N457);
and AND4 (N1174, N1166, N290, N175, N1002);
and AND2 (N1175, N1151, N32);
xor XOR2 (N1176, N1169, N743);
buf BUF1 (N1177, N1167);
nor NOR3 (N1178, N1173, N859, N504);
nand NAND4 (N1179, N1177, N982, N1137, N476);
and AND4 (N1180, N1179, N181, N876, N969);
buf BUF1 (N1181, N1175);
and AND3 (N1182, N1181, N1120, N805);
xor XOR2 (N1183, N1160, N3);
and AND4 (N1184, N1172, N749, N983, N28);
or OR2 (N1185, N1184, N1043);
nor NOR4 (N1186, N1174, N740, N736, N963);
not NOT1 (N1187, N1182);
and AND2 (N1188, N1176, N186);
nor NOR3 (N1189, N1180, N54, N817);
nor NOR2 (N1190, N1171, N833);
not NOT1 (N1191, N1183);
nor NOR3 (N1192, N1165, N596, N303);
nand NAND2 (N1193, N1191, N723);
not NOT1 (N1194, N1187);
not NOT1 (N1195, N1185);
nor NOR4 (N1196, N1189, N576, N1183, N131);
nor NOR4 (N1197, N1195, N1062, N245, N739);
or OR4 (N1198, N1193, N1102, N1018, N978);
and AND2 (N1199, N1192, N437);
nor NOR3 (N1200, N1196, N583, N840);
and AND2 (N1201, N1190, N944);
buf BUF1 (N1202, N1194);
nor NOR3 (N1203, N1199, N247, N368);
xor XOR2 (N1204, N1203, N466);
and AND2 (N1205, N1201, N331);
nor NOR3 (N1206, N1178, N1094, N327);
not NOT1 (N1207, N1188);
and AND3 (N1208, N1198, N1095, N777);
nor NOR4 (N1209, N1208, N991, N857, N612);
buf BUF1 (N1210, N1186);
buf BUF1 (N1211, N1200);
xor XOR2 (N1212, N1205, N195);
and AND4 (N1213, N1212, N822, N48, N830);
or OR4 (N1214, N1206, N547, N89, N357);
or OR4 (N1215, N1210, N23, N535, N258);
nor NOR4 (N1216, N1204, N140, N999, N531);
xor XOR2 (N1217, N1211, N110);
nor NOR2 (N1218, N1215, N156);
or OR2 (N1219, N1216, N520);
nor NOR2 (N1220, N1219, N478);
nor NOR4 (N1221, N1197, N1013, N167, N650);
not NOT1 (N1222, N1202);
nand NAND4 (N1223, N1217, N293, N869, N1097);
xor XOR2 (N1224, N1222, N1168);
nor NOR3 (N1225, N1214, N657, N1109);
and AND3 (N1226, N1209, N353, N913);
not NOT1 (N1227, N1220);
or OR4 (N1228, N1221, N455, N7, N701);
nand NAND4 (N1229, N1163, N572, N310, N209);
buf BUF1 (N1230, N1229);
buf BUF1 (N1231, N1227);
and AND3 (N1232, N1218, N144, N1197);
or OR2 (N1233, N1230, N1223);
and AND2 (N1234, N490, N482);
nor NOR3 (N1235, N1207, N576, N1050);
or OR4 (N1236, N1232, N1030, N480, N867);
buf BUF1 (N1237, N1231);
nor NOR4 (N1238, N1236, N747, N362, N1014);
and AND3 (N1239, N1234, N681, N648);
nor NOR2 (N1240, N1225, N294);
or OR3 (N1241, N1228, N266, N411);
nor NOR4 (N1242, N1213, N542, N432, N1142);
buf BUF1 (N1243, N1233);
xor XOR2 (N1244, N1241, N636);
or OR3 (N1245, N1226, N601, N321);
buf BUF1 (N1246, N1224);
not NOT1 (N1247, N1235);
nor NOR4 (N1248, N1238, N234, N465, N1077);
or OR2 (N1249, N1242, N385);
xor XOR2 (N1250, N1240, N523);
or OR2 (N1251, N1237, N535);
buf BUF1 (N1252, N1239);
nor NOR2 (N1253, N1244, N256);
nand NAND3 (N1254, N1251, N938, N375);
buf BUF1 (N1255, N1250);
buf BUF1 (N1256, N1254);
or OR4 (N1257, N1252, N1152, N828, N243);
not NOT1 (N1258, N1243);
and AND4 (N1259, N1255, N226, N402, N938);
buf BUF1 (N1260, N1249);
not NOT1 (N1261, N1258);
xor XOR2 (N1262, N1246, N1008);
nor NOR4 (N1263, N1259, N177, N848, N538);
nor NOR4 (N1264, N1245, N558, N248, N54);
or OR2 (N1265, N1248, N868);
and AND3 (N1266, N1262, N592, N289);
nor NOR2 (N1267, N1264, N322);
nand NAND4 (N1268, N1267, N876, N696, N328);
nand NAND4 (N1269, N1268, N716, N183, N453);
not NOT1 (N1270, N1247);
buf BUF1 (N1271, N1261);
nand NAND2 (N1272, N1266, N168);
or OR2 (N1273, N1272, N265);
nor NOR4 (N1274, N1260, N201, N1099, N58);
not NOT1 (N1275, N1274);
and AND2 (N1276, N1270, N660);
xor XOR2 (N1277, N1265, N964);
or OR2 (N1278, N1275, N334);
nand NAND2 (N1279, N1276, N917);
nor NOR3 (N1280, N1273, N484, N456);
nand NAND2 (N1281, N1280, N493);
and AND3 (N1282, N1253, N695, N209);
not NOT1 (N1283, N1281);
buf BUF1 (N1284, N1256);
not NOT1 (N1285, N1284);
nand NAND4 (N1286, N1282, N669, N493, N448);
or OR3 (N1287, N1278, N660, N364);
and AND2 (N1288, N1285, N1136);
nor NOR2 (N1289, N1279, N179);
or OR3 (N1290, N1289, N857, N110);
nor NOR3 (N1291, N1277, N561, N1040);
and AND3 (N1292, N1291, N805, N26);
nor NOR2 (N1293, N1292, N732);
and AND4 (N1294, N1293, N1002, N866, N1136);
nor NOR3 (N1295, N1288, N1285, N695);
or OR2 (N1296, N1271, N74);
nand NAND4 (N1297, N1295, N127, N1187, N637);
buf BUF1 (N1298, N1283);
nand NAND4 (N1299, N1269, N845, N892, N205);
not NOT1 (N1300, N1290);
and AND3 (N1301, N1257, N977, N445);
nand NAND2 (N1302, N1287, N977);
and AND3 (N1303, N1298, N693, N369);
or OR3 (N1304, N1303, N1047, N33);
buf BUF1 (N1305, N1294);
buf BUF1 (N1306, N1297);
or OR2 (N1307, N1286, N1017);
nor NOR2 (N1308, N1300, N496);
buf BUF1 (N1309, N1306);
and AND4 (N1310, N1296, N484, N1232, N1112);
or OR4 (N1311, N1310, N1194, N1117, N1223);
nand NAND2 (N1312, N1299, N998);
nand NAND4 (N1313, N1263, N1225, N731, N1000);
nor NOR4 (N1314, N1311, N920, N84, N1242);
or OR4 (N1315, N1308, N409, N440, N971);
nand NAND3 (N1316, N1313, N917, N1113);
and AND4 (N1317, N1316, N920, N1010, N383);
or OR3 (N1318, N1304, N95, N878);
nand NAND2 (N1319, N1314, N1309);
buf BUF1 (N1320, N829);
and AND2 (N1321, N1319, N597);
and AND2 (N1322, N1318, N757);
and AND2 (N1323, N1321, N410);
or OR2 (N1324, N1305, N748);
not NOT1 (N1325, N1320);
not NOT1 (N1326, N1323);
buf BUF1 (N1327, N1326);
or OR3 (N1328, N1315, N851, N713);
buf BUF1 (N1329, N1328);
and AND4 (N1330, N1324, N79, N980, N505);
not NOT1 (N1331, N1302);
or OR2 (N1332, N1301, N392);
xor XOR2 (N1333, N1307, N581);
or OR3 (N1334, N1333, N1332, N613);
nor NOR3 (N1335, N61, N730, N593);
nand NAND4 (N1336, N1329, N920, N1076, N692);
nand NAND3 (N1337, N1336, N1041, N754);
not NOT1 (N1338, N1317);
nand NAND2 (N1339, N1312, N994);
not NOT1 (N1340, N1337);
or OR4 (N1341, N1327, N214, N745, N1310);
nand NAND2 (N1342, N1335, N911);
or OR3 (N1343, N1330, N544, N1227);
and AND4 (N1344, N1339, N1120, N707, N392);
nand NAND3 (N1345, N1343, N935, N605);
xor XOR2 (N1346, N1341, N747);
or OR3 (N1347, N1322, N1137, N246);
and AND3 (N1348, N1347, N1037, N683);
xor XOR2 (N1349, N1348, N1329);
nor NOR3 (N1350, N1344, N40, N694);
xor XOR2 (N1351, N1331, N725);
nand NAND4 (N1352, N1350, N114, N471, N525);
nor NOR4 (N1353, N1351, N947, N763, N364);
buf BUF1 (N1354, N1334);
nor NOR2 (N1355, N1342, N820);
nand NAND4 (N1356, N1352, N500, N86, N1224);
not NOT1 (N1357, N1338);
not NOT1 (N1358, N1346);
nor NOR3 (N1359, N1353, N512, N81);
or OR4 (N1360, N1359, N644, N689, N29);
nand NAND2 (N1361, N1360, N1253);
and AND2 (N1362, N1325, N640);
buf BUF1 (N1363, N1345);
nor NOR3 (N1364, N1363, N585, N273);
nor NOR4 (N1365, N1349, N761, N649, N975);
and AND2 (N1366, N1356, N13);
nand NAND3 (N1367, N1365, N1038, N527);
xor XOR2 (N1368, N1367, N380);
buf BUF1 (N1369, N1358);
or OR2 (N1370, N1368, N686);
nand NAND2 (N1371, N1355, N772);
xor XOR2 (N1372, N1361, N1196);
and AND2 (N1373, N1362, N1062);
nor NOR4 (N1374, N1354, N660, N226, N1120);
xor XOR2 (N1375, N1372, N1335);
nor NOR2 (N1376, N1340, N121);
or OR4 (N1377, N1369, N459, N52, N210);
nor NOR2 (N1378, N1377, N462);
xor XOR2 (N1379, N1375, N43);
not NOT1 (N1380, N1374);
nand NAND2 (N1381, N1376, N177);
xor XOR2 (N1382, N1381, N908);
nand NAND2 (N1383, N1373, N56);
not NOT1 (N1384, N1366);
not NOT1 (N1385, N1379);
or OR4 (N1386, N1357, N597, N343, N122);
nor NOR2 (N1387, N1380, N376);
xor XOR2 (N1388, N1370, N882);
not NOT1 (N1389, N1364);
nand NAND3 (N1390, N1386, N737, N1104);
buf BUF1 (N1391, N1384);
nor NOR2 (N1392, N1391, N776);
and AND2 (N1393, N1390, N4);
nor NOR2 (N1394, N1393, N431);
not NOT1 (N1395, N1394);
nor NOR3 (N1396, N1389, N337, N1041);
buf BUF1 (N1397, N1383);
nand NAND4 (N1398, N1382, N782, N507, N243);
or OR2 (N1399, N1392, N1353);
nand NAND3 (N1400, N1385, N1200, N657);
buf BUF1 (N1401, N1400);
and AND2 (N1402, N1397, N1172);
xor XOR2 (N1403, N1402, N1229);
and AND4 (N1404, N1399, N398, N416, N1323);
nand NAND4 (N1405, N1401, N1236, N324, N130);
nor NOR2 (N1406, N1404, N1203);
and AND3 (N1407, N1396, N198, N632);
and AND4 (N1408, N1395, N652, N632, N443);
buf BUF1 (N1409, N1398);
nand NAND2 (N1410, N1407, N495);
not NOT1 (N1411, N1408);
nor NOR3 (N1412, N1409, N913, N241);
nand NAND4 (N1413, N1378, N161, N482, N719);
buf BUF1 (N1414, N1371);
buf BUF1 (N1415, N1403);
and AND4 (N1416, N1414, N259, N260, N56);
nor NOR4 (N1417, N1410, N1313, N1188, N302);
nand NAND2 (N1418, N1415, N499);
not NOT1 (N1419, N1417);
and AND2 (N1420, N1419, N1356);
not NOT1 (N1421, N1406);
not NOT1 (N1422, N1405);
not NOT1 (N1423, N1416);
nand NAND3 (N1424, N1422, N82, N371);
or OR4 (N1425, N1411, N950, N1081, N290);
not NOT1 (N1426, N1418);
or OR2 (N1427, N1421, N559);
or OR2 (N1428, N1387, N738);
nor NOR4 (N1429, N1428, N818, N118, N763);
xor XOR2 (N1430, N1423, N57);
nand NAND2 (N1431, N1425, N1398);
buf BUF1 (N1432, N1431);
or OR4 (N1433, N1413, N439, N682, N1404);
buf BUF1 (N1434, N1432);
nor NOR4 (N1435, N1427, N996, N1065, N521);
or OR3 (N1436, N1388, N132, N225);
and AND4 (N1437, N1436, N279, N1058, N1363);
or OR4 (N1438, N1433, N577, N1283, N116);
xor XOR2 (N1439, N1434, N270);
not NOT1 (N1440, N1435);
or OR2 (N1441, N1420, N290);
and AND4 (N1442, N1439, N453, N1356, N425);
not NOT1 (N1443, N1412);
or OR3 (N1444, N1430, N1164, N1187);
xor XOR2 (N1445, N1442, N1041);
nand NAND2 (N1446, N1443, N627);
buf BUF1 (N1447, N1429);
not NOT1 (N1448, N1437);
buf BUF1 (N1449, N1438);
buf BUF1 (N1450, N1440);
nand NAND2 (N1451, N1441, N361);
nor NOR4 (N1452, N1450, N349, N178, N202);
buf BUF1 (N1453, N1448);
nand NAND2 (N1454, N1426, N370);
xor XOR2 (N1455, N1451, N730);
nor NOR3 (N1456, N1445, N233, N343);
or OR2 (N1457, N1447, N1445);
xor XOR2 (N1458, N1457, N1116);
and AND4 (N1459, N1449, N659, N443, N607);
nor NOR2 (N1460, N1454, N200);
nor NOR3 (N1461, N1452, N266, N379);
buf BUF1 (N1462, N1459);
and AND3 (N1463, N1424, N737, N116);
buf BUF1 (N1464, N1444);
nor NOR3 (N1465, N1456, N259, N603);
not NOT1 (N1466, N1455);
nand NAND2 (N1467, N1453, N763);
xor XOR2 (N1468, N1458, N987);
not NOT1 (N1469, N1468);
nor NOR2 (N1470, N1467, N119);
nand NAND4 (N1471, N1463, N1081, N141, N1434);
and AND2 (N1472, N1465, N1209);
nor NOR2 (N1473, N1472, N1003);
nor NOR4 (N1474, N1466, N862, N444, N784);
or OR2 (N1475, N1461, N46);
buf BUF1 (N1476, N1470);
nor NOR3 (N1477, N1475, N24, N1224);
or OR3 (N1478, N1464, N1113, N62);
buf BUF1 (N1479, N1471);
not NOT1 (N1480, N1477);
nand NAND4 (N1481, N1473, N1118, N765, N200);
and AND2 (N1482, N1481, N1356);
or OR3 (N1483, N1479, N1016, N1171);
nand NAND2 (N1484, N1478, N282);
buf BUF1 (N1485, N1480);
nor NOR4 (N1486, N1462, N562, N88, N1244);
xor XOR2 (N1487, N1484, N1326);
nor NOR3 (N1488, N1474, N400, N730);
nand NAND3 (N1489, N1482, N635, N1448);
nand NAND3 (N1490, N1446, N427, N529);
xor XOR2 (N1491, N1485, N903);
and AND4 (N1492, N1491, N1110, N330, N1321);
and AND3 (N1493, N1488, N740, N119);
nand NAND3 (N1494, N1476, N1003, N1252);
nand NAND3 (N1495, N1469, N17, N233);
not NOT1 (N1496, N1492);
not NOT1 (N1497, N1495);
nand NAND4 (N1498, N1486, N261, N39, N391);
not NOT1 (N1499, N1460);
xor XOR2 (N1500, N1497, N1107);
nand NAND2 (N1501, N1489, N539);
nor NOR2 (N1502, N1496, N893);
xor XOR2 (N1503, N1501, N1177);
and AND4 (N1504, N1493, N463, N604, N243);
not NOT1 (N1505, N1487);
xor XOR2 (N1506, N1494, N942);
or OR2 (N1507, N1502, N871);
not NOT1 (N1508, N1498);
and AND4 (N1509, N1500, N67, N1346, N230);
nand NAND2 (N1510, N1507, N267);
xor XOR2 (N1511, N1509, N591);
xor XOR2 (N1512, N1508, N611);
nand NAND2 (N1513, N1512, N234);
nor NOR2 (N1514, N1499, N940);
not NOT1 (N1515, N1503);
and AND2 (N1516, N1513, N1029);
or OR2 (N1517, N1511, N1059);
not NOT1 (N1518, N1506);
buf BUF1 (N1519, N1516);
and AND3 (N1520, N1514, N682, N1444);
nand NAND4 (N1521, N1483, N1219, N563, N185);
nor NOR2 (N1522, N1521, N1267);
or OR3 (N1523, N1490, N116, N1089);
xor XOR2 (N1524, N1523, N113);
and AND4 (N1525, N1504, N1195, N773, N181);
nand NAND4 (N1526, N1525, N1089, N736, N642);
and AND3 (N1527, N1505, N122, N650);
xor XOR2 (N1528, N1527, N1048);
or OR2 (N1529, N1522, N652);
nand NAND4 (N1530, N1526, N227, N128, N1063);
not NOT1 (N1531, N1510);
xor XOR2 (N1532, N1515, N1009);
buf BUF1 (N1533, N1518);
or OR2 (N1534, N1519, N1223);
nor NOR4 (N1535, N1531, N1120, N982, N493);
and AND3 (N1536, N1533, N636, N1187);
buf BUF1 (N1537, N1536);
nor NOR4 (N1538, N1517, N1162, N253, N735);
and AND4 (N1539, N1538, N1116, N483, N1207);
buf BUF1 (N1540, N1535);
and AND2 (N1541, N1534, N1004);
nor NOR2 (N1542, N1520, N292);
xor XOR2 (N1543, N1542, N594);
xor XOR2 (N1544, N1530, N551);
not NOT1 (N1545, N1537);
nand NAND3 (N1546, N1528, N779, N1522);
buf BUF1 (N1547, N1529);
xor XOR2 (N1548, N1543, N1159);
or OR4 (N1549, N1544, N59, N939, N729);
and AND3 (N1550, N1548, N1482, N536);
or OR4 (N1551, N1546, N589, N605, N483);
buf BUF1 (N1552, N1550);
or OR3 (N1553, N1545, N1317, N213);
xor XOR2 (N1554, N1553, N742);
nand NAND3 (N1555, N1524, N350, N313);
xor XOR2 (N1556, N1547, N430);
nor NOR4 (N1557, N1556, N30, N716, N1137);
xor XOR2 (N1558, N1532, N819);
or OR2 (N1559, N1541, N332);
buf BUF1 (N1560, N1558);
and AND2 (N1561, N1555, N173);
not NOT1 (N1562, N1552);
not NOT1 (N1563, N1559);
xor XOR2 (N1564, N1554, N1038);
buf BUF1 (N1565, N1563);
buf BUF1 (N1566, N1557);
buf BUF1 (N1567, N1560);
buf BUF1 (N1568, N1565);
and AND3 (N1569, N1540, N413, N808);
not NOT1 (N1570, N1561);
buf BUF1 (N1571, N1568);
nor NOR4 (N1572, N1570, N295, N1428, N981);
xor XOR2 (N1573, N1569, N630);
buf BUF1 (N1574, N1564);
nand NAND2 (N1575, N1567, N89);
and AND3 (N1576, N1571, N752, N405);
or OR4 (N1577, N1576, N256, N208, N1466);
nor NOR2 (N1578, N1549, N533);
nand NAND3 (N1579, N1566, N1230, N1555);
buf BUF1 (N1580, N1562);
xor XOR2 (N1581, N1579, N755);
and AND3 (N1582, N1572, N1027, N225);
buf BUF1 (N1583, N1582);
buf BUF1 (N1584, N1575);
nor NOR2 (N1585, N1551, N501);
and AND2 (N1586, N1573, N161);
not NOT1 (N1587, N1580);
buf BUF1 (N1588, N1578);
xor XOR2 (N1589, N1584, N1568);
and AND3 (N1590, N1539, N868, N1168);
or OR2 (N1591, N1590, N133);
or OR3 (N1592, N1591, N1449, N1002);
and AND2 (N1593, N1588, N691);
not NOT1 (N1594, N1583);
and AND3 (N1595, N1589, N35, N1082);
not NOT1 (N1596, N1593);
or OR3 (N1597, N1581, N233, N871);
and AND4 (N1598, N1585, N401, N524, N239);
or OR4 (N1599, N1592, N239, N1345, N1315);
buf BUF1 (N1600, N1599);
xor XOR2 (N1601, N1598, N973);
not NOT1 (N1602, N1595);
and AND2 (N1603, N1586, N781);
or OR2 (N1604, N1596, N608);
buf BUF1 (N1605, N1603);
buf BUF1 (N1606, N1604);
and AND3 (N1607, N1597, N802, N632);
and AND2 (N1608, N1574, N1008);
not NOT1 (N1609, N1606);
and AND4 (N1610, N1605, N1125, N124, N1453);
not NOT1 (N1611, N1607);
buf BUF1 (N1612, N1601);
nand NAND4 (N1613, N1612, N1130, N337, N1611);
nor NOR2 (N1614, N844, N1348);
not NOT1 (N1615, N1609);
and AND4 (N1616, N1602, N550, N577, N444);
and AND3 (N1617, N1610, N1196, N1372);
xor XOR2 (N1618, N1594, N449);
and AND3 (N1619, N1618, N453, N464);
and AND3 (N1620, N1608, N1156, N505);
and AND2 (N1621, N1617, N1008);
nand NAND3 (N1622, N1587, N874, N502);
xor XOR2 (N1623, N1600, N387);
nand NAND3 (N1624, N1614, N1099, N1023);
not NOT1 (N1625, N1613);
not NOT1 (N1626, N1624);
nor NOR2 (N1627, N1625, N72);
or OR2 (N1628, N1626, N784);
nor NOR4 (N1629, N1621, N311, N1114, N52);
nand NAND4 (N1630, N1628, N621, N46, N154);
and AND4 (N1631, N1629, N1115, N313, N1140);
buf BUF1 (N1632, N1619);
not NOT1 (N1633, N1620);
nand NAND3 (N1634, N1615, N955, N1483);
buf BUF1 (N1635, N1632);
nand NAND3 (N1636, N1622, N506, N1369);
buf BUF1 (N1637, N1633);
nor NOR2 (N1638, N1631, N68);
xor XOR2 (N1639, N1635, N978);
nand NAND4 (N1640, N1634, N1009, N242, N387);
or OR4 (N1641, N1577, N352, N1088, N1399);
nor NOR2 (N1642, N1641, N1519);
xor XOR2 (N1643, N1623, N102);
nand NAND4 (N1644, N1627, N597, N284, N5);
or OR4 (N1645, N1640, N504, N253, N746);
nor NOR2 (N1646, N1643, N320);
and AND3 (N1647, N1642, N1580, N499);
nand NAND4 (N1648, N1646, N1299, N1173, N17);
xor XOR2 (N1649, N1647, N1448);
nor NOR2 (N1650, N1639, N1270);
or OR4 (N1651, N1649, N1072, N1252, N1165);
xor XOR2 (N1652, N1636, N535);
buf BUF1 (N1653, N1644);
nand NAND2 (N1654, N1651, N852);
not NOT1 (N1655, N1637);
buf BUF1 (N1656, N1630);
not NOT1 (N1657, N1652);
nand NAND4 (N1658, N1656, N92, N1489, N1451);
xor XOR2 (N1659, N1616, N823);
nand NAND4 (N1660, N1653, N1435, N717, N47);
xor XOR2 (N1661, N1645, N870);
and AND3 (N1662, N1638, N496, N926);
or OR2 (N1663, N1658, N217);
or OR2 (N1664, N1662, N1000);
buf BUF1 (N1665, N1650);
buf BUF1 (N1666, N1665);
and AND3 (N1667, N1666, N387, N361);
nor NOR2 (N1668, N1655, N1606);
not NOT1 (N1669, N1654);
nor NOR2 (N1670, N1657, N1336);
and AND2 (N1671, N1669, N385);
not NOT1 (N1672, N1664);
not NOT1 (N1673, N1661);
buf BUF1 (N1674, N1660);
xor XOR2 (N1675, N1671, N1429);
buf BUF1 (N1676, N1675);
and AND3 (N1677, N1648, N1094, N1289);
xor XOR2 (N1678, N1668, N882);
not NOT1 (N1679, N1659);
or OR2 (N1680, N1678, N620);
nand NAND3 (N1681, N1673, N1043, N918);
not NOT1 (N1682, N1677);
nor NOR3 (N1683, N1682, N696, N961);
not NOT1 (N1684, N1670);
nand NAND3 (N1685, N1667, N124, N1136);
and AND3 (N1686, N1684, N337, N398);
nor NOR3 (N1687, N1683, N1524, N184);
or OR2 (N1688, N1672, N4);
nand NAND3 (N1689, N1687, N1653, N290);
nand NAND4 (N1690, N1674, N486, N154, N486);
and AND3 (N1691, N1680, N544, N1212);
nand NAND2 (N1692, N1685, N1011);
not NOT1 (N1693, N1663);
buf BUF1 (N1694, N1689);
and AND2 (N1695, N1691, N461);
and AND3 (N1696, N1679, N644, N961);
buf BUF1 (N1697, N1695);
or OR4 (N1698, N1690, N1409, N898, N237);
not NOT1 (N1699, N1676);
nor NOR4 (N1700, N1696, N1248, N1545, N1314);
and AND4 (N1701, N1688, N883, N701, N27);
not NOT1 (N1702, N1699);
nand NAND4 (N1703, N1692, N118, N14, N1253);
nor NOR3 (N1704, N1693, N942, N499);
not NOT1 (N1705, N1698);
or OR3 (N1706, N1700, N713, N915);
nor NOR3 (N1707, N1702, N707, N63);
nand NAND2 (N1708, N1703, N1162);
nor NOR2 (N1709, N1705, N1448);
or OR2 (N1710, N1694, N844);
nor NOR4 (N1711, N1697, N703, N267, N1272);
xor XOR2 (N1712, N1706, N387);
not NOT1 (N1713, N1712);
not NOT1 (N1714, N1711);
nand NAND4 (N1715, N1709, N291, N1428, N209);
or OR3 (N1716, N1715, N108, N595);
nor NOR3 (N1717, N1710, N1620, N1396);
nor NOR4 (N1718, N1714, N10, N1342, N121);
not NOT1 (N1719, N1707);
xor XOR2 (N1720, N1704, N118);
buf BUF1 (N1721, N1681);
not NOT1 (N1722, N1719);
xor XOR2 (N1723, N1686, N1062);
or OR4 (N1724, N1701, N916, N1232, N1712);
nand NAND4 (N1725, N1708, N886, N1079, N435);
nor NOR3 (N1726, N1725, N320, N729);
or OR3 (N1727, N1724, N688, N466);
not NOT1 (N1728, N1718);
nand NAND3 (N1729, N1720, N1621, N1586);
nand NAND4 (N1730, N1726, N1506, N91, N1652);
or OR4 (N1731, N1716, N1001, N814, N243);
and AND2 (N1732, N1723, N457);
and AND3 (N1733, N1730, N367, N1020);
and AND4 (N1734, N1732, N1020, N1078, N1620);
nand NAND2 (N1735, N1721, N1662);
nand NAND2 (N1736, N1729, N1684);
nand NAND3 (N1737, N1713, N1235, N739);
xor XOR2 (N1738, N1737, N1);
xor XOR2 (N1739, N1717, N122);
xor XOR2 (N1740, N1738, N20);
xor XOR2 (N1741, N1728, N488);
nor NOR2 (N1742, N1736, N607);
and AND4 (N1743, N1734, N1213, N1105, N961);
nand NAND4 (N1744, N1731, N1144, N945, N1666);
nor NOR2 (N1745, N1733, N1461);
nor NOR3 (N1746, N1735, N1120, N1021);
nand NAND4 (N1747, N1742, N1277, N873, N1087);
nor NOR4 (N1748, N1741, N479, N389, N849);
not NOT1 (N1749, N1739);
nor NOR4 (N1750, N1749, N1694, N1521, N1730);
and AND2 (N1751, N1727, N1167);
xor XOR2 (N1752, N1747, N1139);
nor NOR3 (N1753, N1746, N229, N923);
xor XOR2 (N1754, N1744, N539);
nand NAND4 (N1755, N1752, N1481, N1407, N379);
or OR3 (N1756, N1755, N1506, N149);
nand NAND3 (N1757, N1722, N209, N593);
and AND4 (N1758, N1754, N13, N718, N900);
xor XOR2 (N1759, N1751, N1678);
not NOT1 (N1760, N1758);
or OR3 (N1761, N1750, N700, N885);
buf BUF1 (N1762, N1743);
nand NAND2 (N1763, N1740, N15);
nand NAND2 (N1764, N1753, N797);
or OR3 (N1765, N1762, N808, N1015);
buf BUF1 (N1766, N1760);
buf BUF1 (N1767, N1757);
nor NOR3 (N1768, N1767, N1270, N1480);
or OR2 (N1769, N1764, N937);
buf BUF1 (N1770, N1763);
nor NOR3 (N1771, N1765, N1507, N972);
and AND3 (N1772, N1745, N257, N922);
or OR2 (N1773, N1768, N39);
nand NAND4 (N1774, N1769, N1236, N385, N804);
or OR4 (N1775, N1756, N928, N132, N1702);
nand NAND3 (N1776, N1761, N295, N1532);
nand NAND2 (N1777, N1772, N272);
and AND3 (N1778, N1775, N577, N1592);
nor NOR2 (N1779, N1766, N1615);
nand NAND4 (N1780, N1774, N289, N837, N95);
and AND2 (N1781, N1778, N1579);
or OR4 (N1782, N1776, N1269, N1729, N94);
and AND2 (N1783, N1759, N1180);
or OR3 (N1784, N1780, N120, N92);
or OR4 (N1785, N1779, N1550, N890, N1547);
buf BUF1 (N1786, N1782);
nor NOR3 (N1787, N1777, N889, N1364);
not NOT1 (N1788, N1785);
xor XOR2 (N1789, N1773, N915);
not NOT1 (N1790, N1787);
not NOT1 (N1791, N1783);
xor XOR2 (N1792, N1784, N79);
and AND2 (N1793, N1788, N60);
not NOT1 (N1794, N1791);
xor XOR2 (N1795, N1786, N191);
and AND2 (N1796, N1794, N223);
xor XOR2 (N1797, N1795, N1470);
not NOT1 (N1798, N1796);
nand NAND3 (N1799, N1770, N1682, N647);
and AND3 (N1800, N1790, N906, N261);
nor NOR4 (N1801, N1748, N209, N191, N1133);
or OR3 (N1802, N1798, N808, N1072);
xor XOR2 (N1803, N1799, N1102);
and AND2 (N1804, N1792, N1660);
nand NAND4 (N1805, N1802, N267, N1662, N510);
not NOT1 (N1806, N1789);
not NOT1 (N1807, N1806);
and AND3 (N1808, N1801, N208, N372);
or OR4 (N1809, N1803, N522, N1409, N549);
and AND3 (N1810, N1771, N170, N1010);
and AND2 (N1811, N1800, N1396);
nor NOR3 (N1812, N1809, N227, N1428);
buf BUF1 (N1813, N1807);
xor XOR2 (N1814, N1810, N1406);
xor XOR2 (N1815, N1797, N990);
buf BUF1 (N1816, N1804);
or OR3 (N1817, N1812, N743, N107);
not NOT1 (N1818, N1815);
and AND3 (N1819, N1793, N1712, N1390);
nand NAND4 (N1820, N1781, N649, N1735, N1557);
and AND2 (N1821, N1818, N600);
xor XOR2 (N1822, N1813, N1105);
or OR2 (N1823, N1819, N886);
not NOT1 (N1824, N1823);
nand NAND3 (N1825, N1814, N1536, N1237);
buf BUF1 (N1826, N1808);
and AND4 (N1827, N1820, N1546, N990, N140);
not NOT1 (N1828, N1821);
or OR4 (N1829, N1826, N1231, N908, N1194);
nand NAND3 (N1830, N1817, N935, N668);
nor NOR3 (N1831, N1811, N747, N1653);
buf BUF1 (N1832, N1825);
nand NAND2 (N1833, N1827, N461);
xor XOR2 (N1834, N1816, N1548);
or OR4 (N1835, N1832, N457, N128, N1115);
nor NOR2 (N1836, N1833, N602);
and AND4 (N1837, N1831, N130, N1247, N1444);
xor XOR2 (N1838, N1829, N668);
nor NOR4 (N1839, N1830, N1709, N516, N206);
buf BUF1 (N1840, N1835);
not NOT1 (N1841, N1839);
xor XOR2 (N1842, N1805, N1548);
not NOT1 (N1843, N1836);
nor NOR3 (N1844, N1828, N1187, N643);
nand NAND2 (N1845, N1843, N1806);
buf BUF1 (N1846, N1837);
not NOT1 (N1847, N1846);
or OR3 (N1848, N1824, N72, N1658);
nor NOR4 (N1849, N1841, N1830, N55, N369);
or OR3 (N1850, N1849, N1382, N419);
and AND4 (N1851, N1822, N1186, N920, N580);
and AND3 (N1852, N1844, N1128, N1127);
not NOT1 (N1853, N1850);
buf BUF1 (N1854, N1842);
xor XOR2 (N1855, N1847, N1604);
not NOT1 (N1856, N1834);
not NOT1 (N1857, N1845);
xor XOR2 (N1858, N1853, N951);
or OR2 (N1859, N1858, N635);
buf BUF1 (N1860, N1838);
and AND4 (N1861, N1851, N804, N561, N253);
nand NAND4 (N1862, N1855, N1359, N108, N598);
not NOT1 (N1863, N1860);
nor NOR2 (N1864, N1862, N326);
nor NOR4 (N1865, N1863, N1554, N1108, N635);
not NOT1 (N1866, N1856);
nand NAND3 (N1867, N1840, N1165, N505);
nor NOR3 (N1868, N1854, N1617, N1398);
nand NAND2 (N1869, N1867, N1133);
buf BUF1 (N1870, N1865);
and AND4 (N1871, N1859, N1022, N943, N1278);
xor XOR2 (N1872, N1869, N452);
xor XOR2 (N1873, N1864, N533);
xor XOR2 (N1874, N1848, N1277);
buf BUF1 (N1875, N1857);
nand NAND3 (N1876, N1872, N106, N958);
nor NOR2 (N1877, N1870, N1692);
buf BUF1 (N1878, N1866);
buf BUF1 (N1879, N1878);
buf BUF1 (N1880, N1868);
or OR4 (N1881, N1876, N1805, N388, N318);
or OR4 (N1882, N1881, N1846, N568, N1560);
nor NOR3 (N1883, N1877, N1773, N1071);
nor NOR2 (N1884, N1861, N1756);
or OR2 (N1885, N1884, N157);
and AND4 (N1886, N1885, N1435, N1047, N1376);
nand NAND3 (N1887, N1880, N1664, N1463);
or OR2 (N1888, N1879, N867);
xor XOR2 (N1889, N1874, N1369);
and AND3 (N1890, N1888, N1484, N173);
nor NOR3 (N1891, N1887, N1002, N460);
not NOT1 (N1892, N1882);
buf BUF1 (N1893, N1892);
nand NAND4 (N1894, N1893, N154, N1544, N696);
or OR3 (N1895, N1889, N1790, N1814);
buf BUF1 (N1896, N1871);
nand NAND2 (N1897, N1890, N732);
nand NAND4 (N1898, N1894, N1371, N278, N271);
xor XOR2 (N1899, N1898, N1692);
nor NOR2 (N1900, N1895, N1063);
xor XOR2 (N1901, N1883, N799);
and AND3 (N1902, N1875, N35, N113);
nor NOR4 (N1903, N1896, N292, N1373, N86);
xor XOR2 (N1904, N1886, N85);
or OR4 (N1905, N1897, N605, N1724, N1873);
buf BUF1 (N1906, N1712);
xor XOR2 (N1907, N1852, N924);
nand NAND2 (N1908, N1900, N1558);
nor NOR2 (N1909, N1903, N1667);
nor NOR4 (N1910, N1907, N285, N94, N1900);
nor NOR4 (N1911, N1909, N784, N348, N1105);
not NOT1 (N1912, N1904);
and AND2 (N1913, N1899, N1357);
buf BUF1 (N1914, N1913);
xor XOR2 (N1915, N1912, N1821);
and AND3 (N1916, N1915, N1400, N1897);
or OR4 (N1917, N1891, N124, N882, N1369);
nand NAND4 (N1918, N1916, N1639, N1080, N886);
nand NAND4 (N1919, N1905, N1905, N787, N1421);
and AND4 (N1920, N1918, N888, N877, N557);
and AND2 (N1921, N1920, N1771);
buf BUF1 (N1922, N1910);
not NOT1 (N1923, N1906);
nor NOR3 (N1924, N1902, N634, N1217);
nand NAND4 (N1925, N1919, N1647, N705, N161);
xor XOR2 (N1926, N1921, N1206);
not NOT1 (N1927, N1924);
xor XOR2 (N1928, N1908, N635);
buf BUF1 (N1929, N1925);
or OR2 (N1930, N1926, N577);
buf BUF1 (N1931, N1929);
or OR2 (N1932, N1911, N1104);
and AND4 (N1933, N1931, N1839, N406, N926);
and AND4 (N1934, N1932, N597, N1526, N643);
xor XOR2 (N1935, N1923, N1321);
nor NOR4 (N1936, N1914, N113, N409, N1804);
buf BUF1 (N1937, N1934);
or OR3 (N1938, N1922, N557, N250);
nand NAND4 (N1939, N1901, N471, N952, N297);
nor NOR3 (N1940, N1927, N1751, N1773);
or OR4 (N1941, N1917, N756, N73, N1513);
buf BUF1 (N1942, N1941);
nand NAND4 (N1943, N1928, N346, N270, N1534);
nor NOR3 (N1944, N1935, N1613, N584);
xor XOR2 (N1945, N1930, N721);
nand NAND4 (N1946, N1937, N1513, N330, N1636);
not NOT1 (N1947, N1938);
nor NOR2 (N1948, N1942, N379);
buf BUF1 (N1949, N1944);
not NOT1 (N1950, N1948);
nand NAND2 (N1951, N1949, N1401);
not NOT1 (N1952, N1936);
nand NAND4 (N1953, N1946, N356, N213, N1634);
and AND3 (N1954, N1952, N760, N14);
buf BUF1 (N1955, N1951);
nand NAND3 (N1956, N1943, N469, N1595);
xor XOR2 (N1957, N1950, N821);
and AND3 (N1958, N1939, N452, N1386);
not NOT1 (N1959, N1945);
or OR2 (N1960, N1957, N1087);
or OR4 (N1961, N1954, N1639, N252, N1637);
buf BUF1 (N1962, N1955);
nor NOR2 (N1963, N1961, N193);
xor XOR2 (N1964, N1940, N1021);
not NOT1 (N1965, N1960);
buf BUF1 (N1966, N1953);
and AND3 (N1967, N1966, N1195, N775);
and AND4 (N1968, N1967, N1154, N1916, N82);
xor XOR2 (N1969, N1968, N663);
or OR2 (N1970, N1964, N1609);
not NOT1 (N1971, N1965);
and AND4 (N1972, N1956, N1127, N1228, N250);
or OR2 (N1973, N1933, N1322);
not NOT1 (N1974, N1958);
nor NOR3 (N1975, N1970, N1205, N1167);
nor NOR3 (N1976, N1972, N628, N192);
and AND4 (N1977, N1969, N199, N623, N1676);
and AND3 (N1978, N1977, N707, N151);
xor XOR2 (N1979, N1976, N493);
not NOT1 (N1980, N1973);
nor NOR3 (N1981, N1971, N401, N1350);
buf BUF1 (N1982, N1962);
not NOT1 (N1983, N1974);
xor XOR2 (N1984, N1979, N466);
nand NAND2 (N1985, N1982, N1764);
or OR3 (N1986, N1985, N1161, N1196);
xor XOR2 (N1987, N1947, N524);
or OR4 (N1988, N1984, N1874, N1243, N1265);
buf BUF1 (N1989, N1983);
xor XOR2 (N1990, N1988, N1238);
nor NOR3 (N1991, N1990, N114, N1884);
xor XOR2 (N1992, N1986, N577);
xor XOR2 (N1993, N1989, N1516);
nand NAND3 (N1994, N1978, N1121, N1499);
nor NOR4 (N1995, N1991, N628, N998, N1725);
not NOT1 (N1996, N1992);
buf BUF1 (N1997, N1963);
not NOT1 (N1998, N1997);
or OR2 (N1999, N1987, N1731);
not NOT1 (N2000, N1975);
xor XOR2 (N2001, N1995, N79);
and AND3 (N2002, N1959, N31, N866);
not NOT1 (N2003, N1981);
not NOT1 (N2004, N2000);
and AND3 (N2005, N2002, N1092, N56);
and AND2 (N2006, N2005, N1812);
xor XOR2 (N2007, N1996, N401);
nand NAND2 (N2008, N2004, N1648);
xor XOR2 (N2009, N1999, N254);
and AND3 (N2010, N1998, N456, N847);
buf BUF1 (N2011, N2010);
and AND2 (N2012, N2008, N294);
nand NAND2 (N2013, N2011, N875);
not NOT1 (N2014, N1993);
nor NOR2 (N2015, N2007, N514);
not NOT1 (N2016, N2006);
nand NAND2 (N2017, N2009, N1692);
xor XOR2 (N2018, N2016, N12);
or OR4 (N2019, N2001, N1236, N829, N276);
not NOT1 (N2020, N2019);
or OR3 (N2021, N2013, N93, N355);
nand NAND3 (N2022, N2018, N1105, N1724);
nand NAND2 (N2023, N1994, N104);
or OR2 (N2024, N2023, N1632);
or OR3 (N2025, N2017, N719, N38);
or OR2 (N2026, N2003, N2001);
nand NAND3 (N2027, N2025, N1063, N181);
nand NAND3 (N2028, N2015, N574, N208);
and AND2 (N2029, N2028, N1439);
buf BUF1 (N2030, N2012);
not NOT1 (N2031, N2027);
and AND4 (N2032, N2022, N714, N1176, N688);
buf BUF1 (N2033, N2014);
nand NAND2 (N2034, N2024, N845);
or OR4 (N2035, N2031, N880, N1261, N88);
xor XOR2 (N2036, N2026, N1306);
nor NOR2 (N2037, N2033, N84);
xor XOR2 (N2038, N2030, N1367);
nor NOR2 (N2039, N1980, N1795);
or OR4 (N2040, N2036, N1770, N1254, N710);
or OR3 (N2041, N2038, N478, N713);
buf BUF1 (N2042, N2032);
nand NAND4 (N2043, N2034, N526, N479, N934);
xor XOR2 (N2044, N2040, N1294);
and AND4 (N2045, N2037, N1474, N1859, N87);
not NOT1 (N2046, N2035);
or OR4 (N2047, N2029, N1037, N1267, N421);
nor NOR4 (N2048, N2043, N1315, N735, N1900);
nand NAND3 (N2049, N2044, N24, N836);
or OR3 (N2050, N2021, N132, N1005);
xor XOR2 (N2051, N2039, N2014);
nor NOR2 (N2052, N2048, N1529);
nor NOR3 (N2053, N2046, N395, N1044);
buf BUF1 (N2054, N2053);
not NOT1 (N2055, N2042);
and AND4 (N2056, N2055, N1194, N344, N881);
buf BUF1 (N2057, N2041);
not NOT1 (N2058, N2020);
nand NAND4 (N2059, N2057, N14, N1197, N909);
and AND4 (N2060, N2052, N1299, N458, N174);
or OR4 (N2061, N2051, N1486, N1196, N786);
or OR4 (N2062, N2059, N297, N970, N562);
and AND2 (N2063, N2050, N1563);
nand NAND3 (N2064, N2054, N1445, N1861);
not NOT1 (N2065, N2061);
nor NOR2 (N2066, N2047, N768);
xor XOR2 (N2067, N2064, N600);
xor XOR2 (N2068, N2049, N1995);
or OR4 (N2069, N2068, N293, N317, N1447);
nor NOR4 (N2070, N2069, N723, N1066, N139);
nor NOR4 (N2071, N2067, N821, N911, N943);
and AND4 (N2072, N2065, N559, N76, N1697);
xor XOR2 (N2073, N2066, N752);
and AND2 (N2074, N2045, N1216);
or OR2 (N2075, N2060, N1206);
buf BUF1 (N2076, N2072);
nor NOR4 (N2077, N2056, N1968, N207, N1221);
nand NAND3 (N2078, N2063, N285, N1663);
not NOT1 (N2079, N2076);
or OR3 (N2080, N2058, N1115, N650);
or OR4 (N2081, N2077, N2072, N1006, N833);
xor XOR2 (N2082, N2071, N1830);
nor NOR4 (N2083, N2075, N1869, N1968, N311);
buf BUF1 (N2084, N2073);
buf BUF1 (N2085, N2078);
not NOT1 (N2086, N2079);
buf BUF1 (N2087, N2082);
buf BUF1 (N2088, N2087);
nand NAND2 (N2089, N2083, N246);
nor NOR4 (N2090, N2070, N518, N713, N1362);
nor NOR4 (N2091, N2081, N2082, N612, N1255);
xor XOR2 (N2092, N2088, N102);
or OR3 (N2093, N2085, N888, N108);
nor NOR3 (N2094, N2084, N1925, N739);
xor XOR2 (N2095, N2074, N757);
nand NAND3 (N2096, N2092, N1732, N482);
nand NAND4 (N2097, N2090, N77, N1629, N1768);
nor NOR3 (N2098, N2062, N1039, N1183);
nor NOR3 (N2099, N2089, N659, N89);
and AND2 (N2100, N2098, N44);
not NOT1 (N2101, N2093);
xor XOR2 (N2102, N2095, N530);
or OR2 (N2103, N2094, N954);
xor XOR2 (N2104, N2080, N655);
xor XOR2 (N2105, N2086, N615);
nand NAND3 (N2106, N2091, N438, N558);
nand NAND2 (N2107, N2104, N1711);
nand NAND4 (N2108, N2106, N201, N1535, N945);
and AND3 (N2109, N2102, N1795, N1630);
and AND2 (N2110, N2096, N1961);
nor NOR4 (N2111, N2110, N1618, N911, N1976);
or OR4 (N2112, N2101, N505, N781, N952);
or OR3 (N2113, N2100, N13, N870);
buf BUF1 (N2114, N2113);
not NOT1 (N2115, N2111);
or OR3 (N2116, N2097, N447, N1079);
and AND2 (N2117, N2108, N546);
not NOT1 (N2118, N2109);
not NOT1 (N2119, N2112);
nand NAND3 (N2120, N2119, N375, N1774);
and AND3 (N2121, N2120, N1148, N1074);
not NOT1 (N2122, N2116);
buf BUF1 (N2123, N2118);
and AND2 (N2124, N2121, N2067);
xor XOR2 (N2125, N2122, N2010);
or OR2 (N2126, N2115, N2105);
nor NOR3 (N2127, N1149, N538, N425);
buf BUF1 (N2128, N2124);
and AND4 (N2129, N2125, N1541, N1913, N1461);
or OR4 (N2130, N2123, N838, N1898, N1117);
or OR3 (N2131, N2103, N1971, N684);
buf BUF1 (N2132, N2127);
and AND3 (N2133, N2129, N591, N985);
xor XOR2 (N2134, N2128, N1322);
or OR4 (N2135, N2126, N942, N934, N1300);
not NOT1 (N2136, N2134);
nand NAND2 (N2137, N2099, N1026);
or OR4 (N2138, N2131, N1494, N199, N467);
nand NAND3 (N2139, N2132, N641, N1387);
xor XOR2 (N2140, N2135, N1144);
or OR4 (N2141, N2117, N444, N1897, N934);
not NOT1 (N2142, N2136);
and AND2 (N2143, N2142, N1066);
or OR2 (N2144, N2133, N1072);
not NOT1 (N2145, N2130);
or OR3 (N2146, N2144, N1345, N1722);
buf BUF1 (N2147, N2114);
nand NAND3 (N2148, N2137, N1758, N2115);
or OR3 (N2149, N2139, N702, N449);
and AND3 (N2150, N2138, N674, N593);
buf BUF1 (N2151, N2148);
nand NAND2 (N2152, N2145, N683);
nand NAND3 (N2153, N2107, N857, N1152);
or OR3 (N2154, N2152, N833, N162);
or OR3 (N2155, N2149, N1316, N241);
xor XOR2 (N2156, N2146, N1185);
xor XOR2 (N2157, N2150, N127);
not NOT1 (N2158, N2143);
or OR2 (N2159, N2147, N1977);
nand NAND3 (N2160, N2153, N1726, N2121);
or OR2 (N2161, N2141, N1512);
or OR2 (N2162, N2154, N972);
not NOT1 (N2163, N2155);
nand NAND3 (N2164, N2163, N370, N1010);
nor NOR3 (N2165, N2159, N803, N1107);
not NOT1 (N2166, N2156);
buf BUF1 (N2167, N2164);
or OR3 (N2168, N2157, N1662, N194);
buf BUF1 (N2169, N2162);
nand NAND2 (N2170, N2160, N662);
not NOT1 (N2171, N2161);
nor NOR3 (N2172, N2158, N1717, N346);
or OR3 (N2173, N2170, N1601, N1979);
and AND2 (N2174, N2151, N1897);
not NOT1 (N2175, N2174);
xor XOR2 (N2176, N2172, N1750);
buf BUF1 (N2177, N2168);
or OR3 (N2178, N2169, N210, N460);
not NOT1 (N2179, N2178);
or OR3 (N2180, N2165, N1049, N341);
not NOT1 (N2181, N2166);
or OR3 (N2182, N2177, N1501, N924);
xor XOR2 (N2183, N2175, N1978);
nand NAND3 (N2184, N2183, N1795, N848);
nand NAND2 (N2185, N2173, N1337);
and AND4 (N2186, N2171, N1972, N230, N2184);
buf BUF1 (N2187, N507);
nand NAND4 (N2188, N2187, N1710, N1176, N1849);
nor NOR3 (N2189, N2180, N1675, N942);
xor XOR2 (N2190, N2188, N303);
nor NOR3 (N2191, N2190, N650, N2015);
and AND3 (N2192, N2191, N977, N334);
xor XOR2 (N2193, N2167, N2067);
nor NOR4 (N2194, N2179, N1079, N48, N1550);
nand NAND3 (N2195, N2176, N1675, N417);
xor XOR2 (N2196, N2192, N201);
not NOT1 (N2197, N2189);
nand NAND3 (N2198, N2140, N1692, N1283);
nor NOR2 (N2199, N2197, N1001);
xor XOR2 (N2200, N2193, N1381);
or OR2 (N2201, N2200, N471);
nand NAND4 (N2202, N2201, N286, N47, N1592);
buf BUF1 (N2203, N2195);
nand NAND2 (N2204, N2202, N544);
and AND2 (N2205, N2194, N755);
not NOT1 (N2206, N2205);
and AND3 (N2207, N2203, N790, N980);
nand NAND4 (N2208, N2182, N218, N1695, N439);
nor NOR3 (N2209, N2207, N832, N258);
or OR2 (N2210, N2198, N134);
or OR3 (N2211, N2208, N1600, N1102);
and AND4 (N2212, N2196, N1873, N257, N261);
nand NAND3 (N2213, N2212, N2005, N2058);
nand NAND2 (N2214, N2181, N1400);
xor XOR2 (N2215, N2206, N1382);
nor NOR2 (N2216, N2199, N1398);
and AND2 (N2217, N2215, N2164);
not NOT1 (N2218, N2186);
nor NOR2 (N2219, N2213, N813);
nor NOR2 (N2220, N2210, N2177);
xor XOR2 (N2221, N2216, N1821);
or OR3 (N2222, N2185, N557, N968);
not NOT1 (N2223, N2221);
buf BUF1 (N2224, N2222);
not NOT1 (N2225, N2214);
nand NAND4 (N2226, N2204, N2023, N474, N72);
not NOT1 (N2227, N2209);
not NOT1 (N2228, N2223);
xor XOR2 (N2229, N2228, N808);
and AND2 (N2230, N2219, N588);
and AND2 (N2231, N2218, N1834);
nand NAND4 (N2232, N2226, N988, N437, N765);
and AND2 (N2233, N2225, N1154);
nor NOR4 (N2234, N2227, N2182, N1952, N913);
not NOT1 (N2235, N2217);
and AND4 (N2236, N2233, N2219, N542, N421);
nand NAND2 (N2237, N2234, N821);
nor NOR4 (N2238, N2237, N1998, N1794, N2149);
xor XOR2 (N2239, N2211, N1909);
nor NOR4 (N2240, N2231, N451, N2116, N1522);
xor XOR2 (N2241, N2235, N131);
or OR3 (N2242, N2241, N2155, N1677);
xor XOR2 (N2243, N2224, N2164);
and AND3 (N2244, N2236, N1784, N1670);
or OR2 (N2245, N2230, N1297);
xor XOR2 (N2246, N2242, N223);
or OR2 (N2247, N2243, N1460);
buf BUF1 (N2248, N2238);
not NOT1 (N2249, N2240);
xor XOR2 (N2250, N2220, N836);
xor XOR2 (N2251, N2248, N1091);
and AND2 (N2252, N2247, N474);
buf BUF1 (N2253, N2246);
and AND3 (N2254, N2250, N590, N1527);
and AND2 (N2255, N2253, N460);
not NOT1 (N2256, N2255);
xor XOR2 (N2257, N2244, N1655);
buf BUF1 (N2258, N2254);
xor XOR2 (N2259, N2251, N2217);
not NOT1 (N2260, N2258);
and AND4 (N2261, N2260, N1623, N1089, N848);
not NOT1 (N2262, N2257);
nand NAND3 (N2263, N2256, N1204, N804);
xor XOR2 (N2264, N2261, N593);
buf BUF1 (N2265, N2239);
nor NOR2 (N2266, N2263, N253);
or OR4 (N2267, N2266, N330, N672, N1344);
and AND4 (N2268, N2249, N1310, N945, N276);
nor NOR2 (N2269, N2265, N354);
not NOT1 (N2270, N2267);
buf BUF1 (N2271, N2269);
nand NAND2 (N2272, N2270, N625);
xor XOR2 (N2273, N2259, N1576);
nor NOR4 (N2274, N2245, N1879, N1285, N1883);
xor XOR2 (N2275, N2229, N270);
xor XOR2 (N2276, N2272, N83);
not NOT1 (N2277, N2252);
buf BUF1 (N2278, N2262);
xor XOR2 (N2279, N2274, N255);
or OR4 (N2280, N2268, N1104, N220, N1450);
nor NOR4 (N2281, N2278, N1060, N859, N382);
and AND2 (N2282, N2279, N269);
nand NAND2 (N2283, N2275, N1337);
and AND4 (N2284, N2283, N1367, N1668, N1802);
nand NAND3 (N2285, N2282, N1524, N741);
and AND4 (N2286, N2284, N1477, N244, N1839);
not NOT1 (N2287, N2277);
nor NOR4 (N2288, N2285, N703, N60, N134);
nor NOR4 (N2289, N2271, N780, N774, N267);
xor XOR2 (N2290, N2281, N1630);
nand NAND2 (N2291, N2264, N664);
nor NOR4 (N2292, N2232, N2286, N2112, N970);
nand NAND3 (N2293, N907, N378, N2265);
and AND2 (N2294, N2289, N2192);
nor NOR4 (N2295, N2273, N1877, N479, N48);
nor NOR3 (N2296, N2292, N772, N1238);
nand NAND3 (N2297, N2280, N1393, N2255);
and AND4 (N2298, N2291, N2061, N105, N1408);
nand NAND4 (N2299, N2287, N2113, N1685, N958);
nand NAND2 (N2300, N2295, N2136);
or OR2 (N2301, N2294, N255);
nand NAND4 (N2302, N2276, N1196, N163, N1741);
or OR3 (N2303, N2302, N1517, N2106);
and AND4 (N2304, N2298, N2027, N858, N701);
and AND4 (N2305, N2300, N1802, N1155, N2087);
buf BUF1 (N2306, N2296);
buf BUF1 (N2307, N2290);
buf BUF1 (N2308, N2299);
nand NAND2 (N2309, N2303, N2208);
or OR3 (N2310, N2308, N1686, N2083);
or OR3 (N2311, N2309, N209, N884);
nor NOR4 (N2312, N2297, N595, N1445, N2190);
or OR2 (N2313, N2311, N1907);
or OR4 (N2314, N2310, N1663, N617, N1041);
buf BUF1 (N2315, N2312);
xor XOR2 (N2316, N2313, N578);
not NOT1 (N2317, N2315);
nor NOR3 (N2318, N2317, N388, N121);
not NOT1 (N2319, N2301);
xor XOR2 (N2320, N2318, N714);
buf BUF1 (N2321, N2304);
nand NAND4 (N2322, N2293, N1269, N761, N1786);
or OR4 (N2323, N2314, N1929, N1360, N1158);
nor NOR2 (N2324, N2323, N75);
not NOT1 (N2325, N2288);
or OR4 (N2326, N2322, N1188, N326, N1248);
buf BUF1 (N2327, N2325);
nor NOR4 (N2328, N2306, N1733, N1514, N1835);
buf BUF1 (N2329, N2320);
buf BUF1 (N2330, N2326);
or OR3 (N2331, N2327, N364, N1057);
xor XOR2 (N2332, N2328, N120);
or OR2 (N2333, N2319, N125);
nand NAND4 (N2334, N2330, N1722, N2086, N1053);
not NOT1 (N2335, N2331);
nor NOR2 (N2336, N2324, N1639);
or OR3 (N2337, N2329, N54, N907);
not NOT1 (N2338, N2305);
not NOT1 (N2339, N2335);
xor XOR2 (N2340, N2338, N701);
buf BUF1 (N2341, N2316);
nand NAND4 (N2342, N2334, N1577, N1821, N1247);
not NOT1 (N2343, N2342);
and AND3 (N2344, N2307, N2341, N154);
buf BUF1 (N2345, N689);
buf BUF1 (N2346, N2332);
and AND2 (N2347, N2337, N439);
not NOT1 (N2348, N2336);
or OR2 (N2349, N2344, N1936);
buf BUF1 (N2350, N2345);
nor NOR4 (N2351, N2346, N204, N2054, N1051);
xor XOR2 (N2352, N2349, N456);
or OR2 (N2353, N2321, N1592);
buf BUF1 (N2354, N2347);
not NOT1 (N2355, N2339);
not NOT1 (N2356, N2351);
buf BUF1 (N2357, N2340);
nand NAND4 (N2358, N2348, N1110, N1511, N2115);
nand NAND2 (N2359, N2356, N385);
nand NAND4 (N2360, N2359, N1716, N900, N458);
buf BUF1 (N2361, N2350);
not NOT1 (N2362, N2355);
or OR2 (N2363, N2353, N1222);
nor NOR2 (N2364, N2360, N2001);
not NOT1 (N2365, N2354);
or OR2 (N2366, N2365, N638);
nor NOR3 (N2367, N2357, N26, N1540);
not NOT1 (N2368, N2361);
and AND2 (N2369, N2364, N349);
and AND3 (N2370, N2352, N110, N749);
and AND4 (N2371, N2368, N813, N2157, N415);
or OR4 (N2372, N2358, N1250, N1182, N850);
and AND3 (N2373, N2362, N1648, N2333);
nand NAND2 (N2374, N604, N896);
xor XOR2 (N2375, N2373, N412);
xor XOR2 (N2376, N2367, N137);
nor NOR3 (N2377, N2366, N952, N638);
and AND2 (N2378, N2370, N182);
buf BUF1 (N2379, N2372);
nor NOR4 (N2380, N2376, N1295, N2136, N148);
nand NAND4 (N2381, N2371, N1845, N275, N1323);
buf BUF1 (N2382, N2375);
xor XOR2 (N2383, N2380, N877);
buf BUF1 (N2384, N2383);
and AND2 (N2385, N2369, N625);
xor XOR2 (N2386, N2343, N2336);
nor NOR2 (N2387, N2384, N81);
xor XOR2 (N2388, N2377, N2253);
or OR3 (N2389, N2387, N925, N2197);
buf BUF1 (N2390, N2382);
and AND2 (N2391, N2388, N2309);
or OR4 (N2392, N2390, N1447, N846, N56);
buf BUF1 (N2393, N2379);
xor XOR2 (N2394, N2363, N629);
nor NOR3 (N2395, N2392, N1604, N444);
xor XOR2 (N2396, N2395, N608);
xor XOR2 (N2397, N2391, N968);
not NOT1 (N2398, N2389);
or OR3 (N2399, N2393, N1654, N1675);
nor NOR4 (N2400, N2378, N2086, N127, N1278);
and AND3 (N2401, N2386, N594, N1967);
buf BUF1 (N2402, N2381);
not NOT1 (N2403, N2396);
and AND2 (N2404, N2397, N1081);
or OR3 (N2405, N2399, N680, N112);
and AND3 (N2406, N2404, N883, N1360);
and AND4 (N2407, N2398, N2353, N870, N1238);
buf BUF1 (N2408, N2394);
and AND3 (N2409, N2374, N1207, N1579);
nor NOR4 (N2410, N2406, N325, N670, N956);
and AND4 (N2411, N2405, N712, N46, N71);
nand NAND2 (N2412, N2411, N1700);
nand NAND3 (N2413, N2385, N22, N166);
not NOT1 (N2414, N2412);
not NOT1 (N2415, N2402);
xor XOR2 (N2416, N2408, N1219);
and AND3 (N2417, N2400, N1793, N2171);
or OR4 (N2418, N2407, N1055, N2279, N2113);
not NOT1 (N2419, N2415);
nor NOR3 (N2420, N2413, N1237, N2383);
nor NOR3 (N2421, N2417, N657, N1450);
nand NAND4 (N2422, N2409, N538, N2332, N1933);
nand NAND2 (N2423, N2414, N57);
xor XOR2 (N2424, N2401, N1381);
and AND2 (N2425, N2419, N450);
buf BUF1 (N2426, N2423);
xor XOR2 (N2427, N2403, N1371);
or OR4 (N2428, N2424, N821, N1407, N1886);
or OR2 (N2429, N2421, N40);
or OR2 (N2430, N2425, N1032);
nand NAND3 (N2431, N2416, N1594, N2182);
or OR2 (N2432, N2428, N2219);
nor NOR2 (N2433, N2427, N2314);
buf BUF1 (N2434, N2422);
xor XOR2 (N2435, N2434, N1607);
nand NAND2 (N2436, N2435, N2087);
or OR2 (N2437, N2410, N1869);
and AND2 (N2438, N2433, N2356);
and AND2 (N2439, N2426, N359);
not NOT1 (N2440, N2420);
and AND4 (N2441, N2431, N1078, N929, N1436);
and AND2 (N2442, N2439, N1915);
not NOT1 (N2443, N2429);
buf BUF1 (N2444, N2418);
and AND2 (N2445, N2444, N1702);
or OR4 (N2446, N2445, N1849, N387, N601);
nor NOR3 (N2447, N2437, N1958, N1828);
buf BUF1 (N2448, N2438);
buf BUF1 (N2449, N2442);
and AND2 (N2450, N2443, N625);
or OR4 (N2451, N2441, N1162, N2438, N979);
buf BUF1 (N2452, N2432);
buf BUF1 (N2453, N2451);
nand NAND3 (N2454, N2453, N583, N1988);
and AND4 (N2455, N2448, N962, N1927, N1606);
nor NOR3 (N2456, N2447, N1654, N1487);
nand NAND2 (N2457, N2456, N2034);
not NOT1 (N2458, N2440);
and AND4 (N2459, N2454, N1198, N378, N1703);
or OR3 (N2460, N2457, N1768, N773);
nor NOR4 (N2461, N2458, N2064, N2130, N69);
nor NOR4 (N2462, N2446, N1583, N1370, N64);
not NOT1 (N2463, N2462);
not NOT1 (N2464, N2461);
buf BUF1 (N2465, N2449);
and AND3 (N2466, N2436, N961, N1882);
not NOT1 (N2467, N2459);
or OR4 (N2468, N2430, N1710, N1678, N394);
and AND3 (N2469, N2452, N343, N292);
not NOT1 (N2470, N2467);
buf BUF1 (N2471, N2460);
or OR2 (N2472, N2470, N1058);
xor XOR2 (N2473, N2465, N1203);
or OR4 (N2474, N2469, N1516, N1578, N620);
xor XOR2 (N2475, N2471, N2180);
and AND2 (N2476, N2463, N2026);
or OR3 (N2477, N2475, N2022, N1838);
xor XOR2 (N2478, N2464, N1055);
not NOT1 (N2479, N2472);
not NOT1 (N2480, N2468);
or OR4 (N2481, N2476, N2107, N321, N2170);
buf BUF1 (N2482, N2481);
nor NOR3 (N2483, N2473, N1335, N1682);
and AND3 (N2484, N2478, N1893, N1746);
or OR2 (N2485, N2474, N2373);
nor NOR3 (N2486, N2484, N73, N1253);
not NOT1 (N2487, N2483);
xor XOR2 (N2488, N2486, N673);
xor XOR2 (N2489, N2466, N1893);
or OR3 (N2490, N2479, N1344, N665);
nand NAND2 (N2491, N2450, N1408);
xor XOR2 (N2492, N2480, N1875);
or OR4 (N2493, N2489, N353, N814, N1539);
nand NAND4 (N2494, N2492, N111, N986, N751);
buf BUF1 (N2495, N2493);
nor NOR2 (N2496, N2477, N1780);
and AND3 (N2497, N2491, N86, N1794);
buf BUF1 (N2498, N2494);
buf BUF1 (N2499, N2497);
and AND2 (N2500, N2488, N656);
nor NOR2 (N2501, N2500, N2384);
not NOT1 (N2502, N2501);
nor NOR2 (N2503, N2496, N12);
nor NOR3 (N2504, N2503, N1570, N1250);
not NOT1 (N2505, N2499);
not NOT1 (N2506, N2455);
xor XOR2 (N2507, N2502, N2130);
buf BUF1 (N2508, N2490);
or OR3 (N2509, N2485, N1549, N530);
xor XOR2 (N2510, N2495, N2003);
nand NAND4 (N2511, N2507, N471, N694, N449);
nor NOR2 (N2512, N2506, N1131);
nand NAND2 (N2513, N2498, N2167);
not NOT1 (N2514, N2509);
and AND2 (N2515, N2487, N1043);
xor XOR2 (N2516, N2515, N1695);
or OR4 (N2517, N2510, N1559, N1523, N1077);
xor XOR2 (N2518, N2513, N1194);
buf BUF1 (N2519, N2504);
nor NOR3 (N2520, N2518, N476, N1619);
and AND4 (N2521, N2512, N724, N2401, N259);
nor NOR3 (N2522, N2520, N1372, N101);
or OR3 (N2523, N2482, N635, N341);
not NOT1 (N2524, N2516);
xor XOR2 (N2525, N2524, N1443);
buf BUF1 (N2526, N2523);
or OR2 (N2527, N2526, N1448);
xor XOR2 (N2528, N2521, N1731);
buf BUF1 (N2529, N2519);
and AND3 (N2530, N2505, N1631, N1186);
nand NAND3 (N2531, N2514, N477, N1100);
buf BUF1 (N2532, N2531);
nor NOR2 (N2533, N2532, N1939);
not NOT1 (N2534, N2529);
and AND3 (N2535, N2517, N67, N945);
not NOT1 (N2536, N2522);
nor NOR3 (N2537, N2525, N583, N563);
buf BUF1 (N2538, N2530);
not NOT1 (N2539, N2535);
and AND4 (N2540, N2533, N790, N23, N1319);
not NOT1 (N2541, N2508);
nand NAND4 (N2542, N2538, N1732, N1927, N1728);
nor NOR3 (N2543, N2527, N829, N2522);
xor XOR2 (N2544, N2542, N893);
xor XOR2 (N2545, N2534, N1319);
xor XOR2 (N2546, N2511, N1733);
buf BUF1 (N2547, N2536);
buf BUF1 (N2548, N2546);
nand NAND4 (N2549, N2541, N1330, N1206, N2076);
or OR4 (N2550, N2549, N418, N1527, N212);
nand NAND2 (N2551, N2550, N991);
or OR4 (N2552, N2545, N2308, N691, N1771);
xor XOR2 (N2553, N2544, N73);
nor NOR3 (N2554, N2537, N295, N1121);
xor XOR2 (N2555, N2543, N1070);
nand NAND2 (N2556, N2547, N2386);
or OR2 (N2557, N2555, N1266);
and AND3 (N2558, N2552, N395, N2255);
not NOT1 (N2559, N2548);
nor NOR3 (N2560, N2559, N892, N1552);
or OR4 (N2561, N2558, N432, N1115, N2328);
xor XOR2 (N2562, N2551, N24);
and AND4 (N2563, N2560, N2403, N1633, N253);
nand NAND3 (N2564, N2528, N343, N382);
nor NOR2 (N2565, N2562, N350);
or OR4 (N2566, N2557, N1302, N1360, N35);
xor XOR2 (N2567, N2540, N2388);
and AND3 (N2568, N2567, N1776, N1057);
and AND3 (N2569, N2563, N906, N345);
xor XOR2 (N2570, N2566, N56);
nand NAND2 (N2571, N2564, N1759);
and AND3 (N2572, N2554, N1764, N1155);
nor NOR3 (N2573, N2572, N1651, N999);
xor XOR2 (N2574, N2570, N1035);
nor NOR3 (N2575, N2556, N1650, N35);
and AND4 (N2576, N2573, N650, N2104, N462);
or OR3 (N2577, N2574, N415, N2431);
buf BUF1 (N2578, N2575);
nor NOR3 (N2579, N2568, N1069, N469);
not NOT1 (N2580, N2565);
not NOT1 (N2581, N2580);
and AND2 (N2582, N2571, N280);
nor NOR4 (N2583, N2561, N199, N356, N350);
nand NAND2 (N2584, N2581, N421);
or OR2 (N2585, N2569, N692);
xor XOR2 (N2586, N2578, N1740);
xor XOR2 (N2587, N2583, N1271);
nor NOR2 (N2588, N2553, N1463);
nor NOR2 (N2589, N2539, N556);
not NOT1 (N2590, N2579);
and AND4 (N2591, N2582, N304, N1251, N193);
nor NOR3 (N2592, N2590, N1919, N2477);
xor XOR2 (N2593, N2586, N2315);
and AND4 (N2594, N2577, N594, N1146, N26);
xor XOR2 (N2595, N2576, N2371);
and AND3 (N2596, N2584, N1278, N1345);
nor NOR2 (N2597, N2593, N1557);
xor XOR2 (N2598, N2597, N2042);
nand NAND4 (N2599, N2592, N577, N2348, N1652);
xor XOR2 (N2600, N2599, N199);
and AND4 (N2601, N2585, N1022, N641, N1877);
nand NAND3 (N2602, N2600, N752, N778);
or OR3 (N2603, N2601, N1175, N1210);
and AND3 (N2604, N2591, N220, N1849);
nand NAND4 (N2605, N2598, N2101, N2458, N1957);
nor NOR2 (N2606, N2594, N2497);
not NOT1 (N2607, N2605);
xor XOR2 (N2608, N2602, N1189);
nand NAND3 (N2609, N2607, N1650, N125);
nand NAND4 (N2610, N2608, N1432, N800, N1311);
or OR2 (N2611, N2589, N2013);
not NOT1 (N2612, N2611);
nand NAND3 (N2613, N2587, N2056, N576);
nand NAND2 (N2614, N2613, N321);
buf BUF1 (N2615, N2588);
buf BUF1 (N2616, N2603);
buf BUF1 (N2617, N2609);
or OR2 (N2618, N2612, N2563);
and AND4 (N2619, N2615, N390, N1757, N1519);
buf BUF1 (N2620, N2595);
xor XOR2 (N2621, N2617, N667);
nor NOR4 (N2622, N2618, N1085, N1495, N535);
not NOT1 (N2623, N2622);
not NOT1 (N2624, N2620);
xor XOR2 (N2625, N2606, N416);
buf BUF1 (N2626, N2621);
nor NOR3 (N2627, N2619, N2247, N159);
nor NOR4 (N2628, N2626, N1718, N2241, N172);
not NOT1 (N2629, N2614);
not NOT1 (N2630, N2610);
nor NOR2 (N2631, N2604, N726);
and AND4 (N2632, N2630, N118, N1129, N458);
and AND2 (N2633, N2629, N1772);
buf BUF1 (N2634, N2625);
nand NAND2 (N2635, N2634, N1603);
xor XOR2 (N2636, N2628, N1185);
or OR2 (N2637, N2633, N1926);
nand NAND4 (N2638, N2596, N1010, N3, N2492);
not NOT1 (N2639, N2638);
nor NOR3 (N2640, N2637, N1195, N2338);
not NOT1 (N2641, N2636);
and AND3 (N2642, N2640, N2534, N55);
and AND3 (N2643, N2642, N2407, N1858);
nand NAND4 (N2644, N2643, N1367, N2289, N256);
nand NAND3 (N2645, N2623, N2224, N1350);
or OR4 (N2646, N2631, N1357, N803, N383);
or OR2 (N2647, N2646, N258);
buf BUF1 (N2648, N2632);
nand NAND3 (N2649, N2647, N660, N2644);
xor XOR2 (N2650, N2233, N20);
or OR3 (N2651, N2639, N2432, N1235);
buf BUF1 (N2652, N2645);
buf BUF1 (N2653, N2635);
nor NOR4 (N2654, N2641, N223, N2409, N1465);
not NOT1 (N2655, N2652);
nand NAND4 (N2656, N2649, N1149, N289, N808);
nand NAND2 (N2657, N2654, N2069);
nor NOR4 (N2658, N2624, N2024, N495, N2101);
xor XOR2 (N2659, N2650, N1920);
not NOT1 (N2660, N2656);
nor NOR2 (N2661, N2658, N2514);
or OR2 (N2662, N2616, N2161);
and AND4 (N2663, N2657, N2352, N137, N750);
xor XOR2 (N2664, N2627, N1459);
nand NAND3 (N2665, N2662, N1925, N1164);
nand NAND4 (N2666, N2660, N2147, N2135, N1634);
buf BUF1 (N2667, N2651);
xor XOR2 (N2668, N2667, N199);
and AND4 (N2669, N2664, N750, N1924, N621);
or OR3 (N2670, N2665, N394, N608);
buf BUF1 (N2671, N2666);
nor NOR4 (N2672, N2669, N2219, N620, N902);
and AND2 (N2673, N2668, N684);
buf BUF1 (N2674, N2653);
and AND4 (N2675, N2674, N1146, N1719, N1662);
not NOT1 (N2676, N2663);
and AND3 (N2677, N2659, N1869, N127);
and AND3 (N2678, N2670, N392, N66);
or OR4 (N2679, N2671, N1426, N438, N2021);
nand NAND3 (N2680, N2679, N88, N1498);
and AND3 (N2681, N2655, N2482, N412);
or OR2 (N2682, N2677, N1050);
and AND3 (N2683, N2678, N999, N2674);
and AND4 (N2684, N2675, N1806, N2042, N200);
or OR2 (N2685, N2648, N1501);
not NOT1 (N2686, N2684);
xor XOR2 (N2687, N2686, N1289);
xor XOR2 (N2688, N2673, N2040);
not NOT1 (N2689, N2685);
nor NOR2 (N2690, N2687, N1147);
xor XOR2 (N2691, N2661, N913);
or OR2 (N2692, N2681, N681);
and AND4 (N2693, N2688, N1584, N1272, N2588);
nor NOR4 (N2694, N2691, N1673, N673, N8);
nor NOR2 (N2695, N2692, N2174);
or OR2 (N2696, N2689, N293);
buf BUF1 (N2697, N2694);
buf BUF1 (N2698, N2683);
nor NOR3 (N2699, N2693, N1039, N2314);
not NOT1 (N2700, N2676);
or OR4 (N2701, N2698, N2215, N355, N503);
nand NAND3 (N2702, N2696, N394, N1861);
nor NOR2 (N2703, N2680, N930);
and AND2 (N2704, N2702, N879);
nand NAND3 (N2705, N2672, N520, N2188);
nor NOR3 (N2706, N2695, N125, N1317);
not NOT1 (N2707, N2704);
nand NAND4 (N2708, N2699, N1609, N2660, N1280);
buf BUF1 (N2709, N2701);
or OR2 (N2710, N2705, N377);
not NOT1 (N2711, N2690);
or OR2 (N2712, N2711, N376);
buf BUF1 (N2713, N2709);
nand NAND4 (N2714, N2710, N1400, N927, N1018);
nor NOR4 (N2715, N2703, N462, N893, N1402);
nor NOR4 (N2716, N2697, N485, N648, N1386);
and AND2 (N2717, N2700, N12);
or OR3 (N2718, N2717, N1668, N1940);
nor NOR2 (N2719, N2712, N1921);
buf BUF1 (N2720, N2706);
and AND2 (N2721, N2707, N905);
and AND3 (N2722, N2682, N1547, N2638);
xor XOR2 (N2723, N2718, N2007);
not NOT1 (N2724, N2708);
or OR3 (N2725, N2719, N1095, N1391);
buf BUF1 (N2726, N2723);
nand NAND4 (N2727, N2722, N1635, N1941, N1071);
nand NAND3 (N2728, N2725, N2191, N2573);
nor NOR2 (N2729, N2715, N1014);
or OR4 (N2730, N2716, N462, N906, N441);
not NOT1 (N2731, N2721);
or OR2 (N2732, N2730, N13);
nor NOR3 (N2733, N2728, N2193, N837);
nor NOR3 (N2734, N2733, N1464, N1433);
buf BUF1 (N2735, N2734);
not NOT1 (N2736, N2726);
not NOT1 (N2737, N2720);
nand NAND3 (N2738, N2727, N1124, N350);
nand NAND2 (N2739, N2732, N2134);
and AND4 (N2740, N2729, N1825, N920, N734);
or OR2 (N2741, N2713, N1470);
and AND4 (N2742, N2731, N239, N1541, N1039);
or OR4 (N2743, N2738, N507, N213, N2514);
not NOT1 (N2744, N2743);
and AND4 (N2745, N2744, N459, N1366, N1591);
not NOT1 (N2746, N2745);
not NOT1 (N2747, N2746);
buf BUF1 (N2748, N2740);
nor NOR4 (N2749, N2735, N1510, N692, N2272);
or OR4 (N2750, N2747, N966, N1819, N457);
and AND2 (N2751, N2749, N1260);
and AND2 (N2752, N2736, N461);
xor XOR2 (N2753, N2741, N2488);
and AND4 (N2754, N2751, N2029, N1378, N705);
buf BUF1 (N2755, N2748);
buf BUF1 (N2756, N2714);
buf BUF1 (N2757, N2750);
and AND3 (N2758, N2753, N1555, N29);
nand NAND4 (N2759, N2752, N1257, N2259, N1183);
buf BUF1 (N2760, N2758);
nor NOR2 (N2761, N2755, N2110);
or OR4 (N2762, N2757, N2368, N2295, N691);
xor XOR2 (N2763, N2754, N2632);
nor NOR2 (N2764, N2760, N286);
and AND4 (N2765, N2763, N1080, N1616, N1905);
nor NOR2 (N2766, N2737, N602);
nand NAND3 (N2767, N2764, N1460, N1917);
not NOT1 (N2768, N2739);
nor NOR2 (N2769, N2765, N868);
nand NAND3 (N2770, N2761, N2544, N719);
or OR4 (N2771, N2724, N1531, N444, N1677);
or OR3 (N2772, N2770, N454, N1715);
or OR4 (N2773, N2769, N2020, N890, N415);
not NOT1 (N2774, N2773);
or OR3 (N2775, N2772, N1524, N431);
or OR4 (N2776, N2762, N1048, N2074, N1241);
buf BUF1 (N2777, N2742);
or OR3 (N2778, N2775, N2069, N2255);
xor XOR2 (N2779, N2778, N590);
not NOT1 (N2780, N2771);
not NOT1 (N2781, N2768);
xor XOR2 (N2782, N2780, N1706);
nand NAND4 (N2783, N2779, N1372, N1066, N284);
nor NOR3 (N2784, N2766, N2588, N1659);
nor NOR3 (N2785, N2759, N2159, N1556);
and AND4 (N2786, N2774, N1345, N1174, N1568);
not NOT1 (N2787, N2782);
not NOT1 (N2788, N2777);
not NOT1 (N2789, N2767);
not NOT1 (N2790, N2756);
or OR4 (N2791, N2788, N2483, N304, N2702);
or OR3 (N2792, N2784, N524, N2535);
xor XOR2 (N2793, N2787, N1014);
xor XOR2 (N2794, N2789, N2170);
xor XOR2 (N2795, N2786, N1136);
and AND2 (N2796, N2794, N2595);
nand NAND2 (N2797, N2796, N2183);
nand NAND3 (N2798, N2792, N1647, N2496);
nand NAND4 (N2799, N2785, N1042, N553, N1610);
and AND2 (N2800, N2798, N1873);
xor XOR2 (N2801, N2791, N2671);
or OR2 (N2802, N2776, N660);
nand NAND3 (N2803, N2799, N2734, N2479);
xor XOR2 (N2804, N2795, N2515);
and AND3 (N2805, N2802, N904, N1435);
or OR3 (N2806, N2803, N2550, N1973);
or OR2 (N2807, N2781, N2306);
xor XOR2 (N2808, N2801, N1171);
not NOT1 (N2809, N2808);
nand NAND4 (N2810, N2783, N1866, N1233, N1526);
nand NAND3 (N2811, N2806, N431, N1038);
not NOT1 (N2812, N2811);
xor XOR2 (N2813, N2809, N2684);
xor XOR2 (N2814, N2812, N1091);
buf BUF1 (N2815, N2797);
xor XOR2 (N2816, N2804, N2594);
nand NAND2 (N2817, N2807, N1204);
nand NAND4 (N2818, N2813, N2588, N2631, N2195);
and AND2 (N2819, N2805, N2786);
or OR4 (N2820, N2819, N668, N742, N2365);
not NOT1 (N2821, N2790);
not NOT1 (N2822, N2810);
or OR2 (N2823, N2793, N382);
buf BUF1 (N2824, N2815);
xor XOR2 (N2825, N2814, N2549);
and AND4 (N2826, N2817, N89, N470, N1040);
nor NOR2 (N2827, N2825, N1916);
not NOT1 (N2828, N2826);
and AND3 (N2829, N2816, N2006, N2044);
or OR2 (N2830, N2827, N2757);
not NOT1 (N2831, N2820);
xor XOR2 (N2832, N2818, N1163);
nor NOR3 (N2833, N2831, N133, N2647);
xor XOR2 (N2834, N2824, N2498);
xor XOR2 (N2835, N2823, N950);
buf BUF1 (N2836, N2833);
nor NOR4 (N2837, N2832, N1500, N1537, N1649);
or OR3 (N2838, N2835, N641, N362);
buf BUF1 (N2839, N2822);
buf BUF1 (N2840, N2830);
nor NOR3 (N2841, N2800, N1968, N400);
nand NAND3 (N2842, N2834, N735, N1379);
not NOT1 (N2843, N2838);
nor NOR4 (N2844, N2840, N259, N122, N1635);
nand NAND4 (N2845, N2837, N1838, N1356, N1240);
or OR2 (N2846, N2842, N256);
buf BUF1 (N2847, N2845);
buf BUF1 (N2848, N2846);
not NOT1 (N2849, N2841);
nand NAND4 (N2850, N2828, N8, N481, N2089);
not NOT1 (N2851, N2843);
and AND4 (N2852, N2829, N889, N1056, N384);
or OR2 (N2853, N2848, N672);
or OR2 (N2854, N2844, N1520);
nand NAND2 (N2855, N2849, N1877);
or OR3 (N2856, N2821, N1289, N272);
and AND4 (N2857, N2839, N620, N2244, N1717);
xor XOR2 (N2858, N2856, N2157);
xor XOR2 (N2859, N2850, N875);
buf BUF1 (N2860, N2847);
xor XOR2 (N2861, N2853, N1088);
nor NOR3 (N2862, N2859, N2058, N1863);
or OR3 (N2863, N2860, N98, N2702);
nor NOR3 (N2864, N2858, N1460, N1228);
or OR3 (N2865, N2864, N1451, N2222);
not NOT1 (N2866, N2863);
not NOT1 (N2867, N2861);
nor NOR4 (N2868, N2867, N2093, N1942, N1531);
not NOT1 (N2869, N2855);
or OR2 (N2870, N2869, N1932);
or OR2 (N2871, N2868, N308);
xor XOR2 (N2872, N2851, N1761);
or OR4 (N2873, N2870, N945, N1887, N597);
nor NOR4 (N2874, N2854, N1316, N1244, N1428);
xor XOR2 (N2875, N2836, N1711);
buf BUF1 (N2876, N2865);
or OR3 (N2877, N2875, N795, N2610);
and AND2 (N2878, N2852, N1306);
not NOT1 (N2879, N2876);
xor XOR2 (N2880, N2877, N2069);
or OR4 (N2881, N2872, N54, N2582, N1763);
or OR4 (N2882, N2878, N2767, N2871, N1125);
and AND3 (N2883, N607, N1914, N1656);
buf BUF1 (N2884, N2862);
xor XOR2 (N2885, N2874, N1800);
or OR3 (N2886, N2881, N669, N123);
and AND2 (N2887, N2873, N985);
xor XOR2 (N2888, N2883, N2703);
or OR3 (N2889, N2887, N1035, N2785);
buf BUF1 (N2890, N2885);
nor NOR2 (N2891, N2880, N2494);
nand NAND2 (N2892, N2889, N66);
nand NAND2 (N2893, N2884, N633);
or OR3 (N2894, N2893, N642, N2496);
or OR2 (N2895, N2882, N1593);
or OR3 (N2896, N2891, N1620, N2289);
xor XOR2 (N2897, N2896, N1045);
and AND4 (N2898, N2886, N928, N1070, N2773);
buf BUF1 (N2899, N2892);
nand NAND4 (N2900, N2898, N2381, N674, N1812);
buf BUF1 (N2901, N2890);
not NOT1 (N2902, N2901);
not NOT1 (N2903, N2888);
nand NAND4 (N2904, N2902, N1409, N2692, N1454);
or OR3 (N2905, N2897, N1262, N2619);
nand NAND2 (N2906, N2903, N2340);
buf BUF1 (N2907, N2879);
nand NAND2 (N2908, N2900, N2315);
nor NOR3 (N2909, N2866, N47, N605);
xor XOR2 (N2910, N2895, N2411);
or OR2 (N2911, N2908, N1184);
xor XOR2 (N2912, N2911, N232);
and AND3 (N2913, N2857, N1470, N2664);
nand NAND2 (N2914, N2909, N2202);
xor XOR2 (N2915, N2907, N929);
xor XOR2 (N2916, N2906, N1606);
nor NOR4 (N2917, N2914, N2225, N2567, N2791);
xor XOR2 (N2918, N2917, N2353);
and AND3 (N2919, N2894, N2389, N821);
nand NAND3 (N2920, N2918, N1591, N736);
not NOT1 (N2921, N2913);
nand NAND2 (N2922, N2910, N452);
xor XOR2 (N2923, N2919, N1318);
xor XOR2 (N2924, N2921, N2545);
not NOT1 (N2925, N2904);
or OR2 (N2926, N2912, N2289);
not NOT1 (N2927, N2916);
xor XOR2 (N2928, N2899, N2029);
buf BUF1 (N2929, N2922);
xor XOR2 (N2930, N2926, N365);
nand NAND2 (N2931, N2915, N703);
buf BUF1 (N2932, N2905);
nand NAND4 (N2933, N2932, N1995, N2311, N1111);
not NOT1 (N2934, N2930);
xor XOR2 (N2935, N2931, N1624);
xor XOR2 (N2936, N2934, N344);
not NOT1 (N2937, N2936);
not NOT1 (N2938, N2935);
not NOT1 (N2939, N2924);
or OR3 (N2940, N2933, N1645, N223);
buf BUF1 (N2941, N2928);
not NOT1 (N2942, N2941);
and AND4 (N2943, N2939, N900, N765, N2822);
and AND3 (N2944, N2940, N2196, N2280);
or OR3 (N2945, N2937, N2130, N850);
nor NOR4 (N2946, N2943, N637, N1247, N2500);
buf BUF1 (N2947, N2927);
or OR4 (N2948, N2938, N756, N1771, N1279);
and AND2 (N2949, N2947, N78);
and AND2 (N2950, N2923, N2478);
or OR3 (N2951, N2944, N931, N1615);
xor XOR2 (N2952, N2949, N1933);
xor XOR2 (N2953, N2952, N85);
nand NAND4 (N2954, N2925, N2107, N811, N1353);
xor XOR2 (N2955, N2946, N1654);
nand NAND2 (N2956, N2951, N1128);
or OR3 (N2957, N2950, N2217, N2338);
and AND4 (N2958, N2942, N70, N2202, N691);
xor XOR2 (N2959, N2948, N2198);
and AND2 (N2960, N2956, N627);
buf BUF1 (N2961, N2957);
not NOT1 (N2962, N2945);
and AND4 (N2963, N2920, N2490, N1453, N2863);
not NOT1 (N2964, N2955);
and AND4 (N2965, N2958, N1544, N2925, N2957);
or OR3 (N2966, N2965, N2750, N1796);
or OR3 (N2967, N2953, N2281, N2598);
xor XOR2 (N2968, N2963, N1058);
not NOT1 (N2969, N2929);
nor NOR4 (N2970, N2959, N474, N1727, N485);
xor XOR2 (N2971, N2962, N222);
and AND2 (N2972, N2960, N263);
and AND3 (N2973, N2968, N1472, N1132);
not NOT1 (N2974, N2966);
nor NOR3 (N2975, N2967, N2476, N1164);
and AND4 (N2976, N2975, N1888, N2391, N1261);
xor XOR2 (N2977, N2973, N2596);
not NOT1 (N2978, N2976);
buf BUF1 (N2979, N2961);
and AND2 (N2980, N2978, N1098);
nand NAND4 (N2981, N2977, N21, N1531, N1329);
not NOT1 (N2982, N2979);
and AND2 (N2983, N2970, N2176);
buf BUF1 (N2984, N2971);
or OR3 (N2985, N2972, N1138, N662);
buf BUF1 (N2986, N2964);
nand NAND2 (N2987, N2986, N692);
nand NAND3 (N2988, N2980, N2482, N2543);
nor NOR2 (N2989, N2981, N1728);
or OR3 (N2990, N2984, N167, N162);
nand NAND2 (N2991, N2988, N1883);
nor NOR3 (N2992, N2983, N2737, N1120);
buf BUF1 (N2993, N2974);
xor XOR2 (N2994, N2990, N1123);
or OR4 (N2995, N2987, N2175, N2081, N923);
or OR4 (N2996, N2989, N813, N1520, N67);
or OR4 (N2997, N2993, N208, N1454, N1515);
and AND4 (N2998, N2992, N1331, N2166, N644);
xor XOR2 (N2999, N2998, N329);
nand NAND3 (N3000, N2991, N2107, N550);
or OR4 (N3001, N2996, N917, N2855, N1409);
or OR2 (N3002, N2994, N1712);
nor NOR4 (N3003, N3000, N1284, N2422, N2569);
xor XOR2 (N3004, N2982, N539);
nand NAND4 (N3005, N2995, N1211, N1142, N3000);
and AND3 (N3006, N3005, N118, N2852);
not NOT1 (N3007, N2997);
xor XOR2 (N3008, N3007, N2402);
buf BUF1 (N3009, N3008);
nand NAND2 (N3010, N3004, N1796);
and AND2 (N3011, N3010, N1748);
endmodule