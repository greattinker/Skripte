// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18;

output N416,N404,N417,N415,N411,N406,N414,N380,N412,N418;

nand NAND2 (N19, N18, N15);
and AND4 (N20, N3, N18, N16, N11);
xor XOR2 (N21, N9, N20);
xor XOR2 (N22, N4, N6);
nor NOR4 (N23, N22, N12, N21, N18);
not NOT1 (N24, N23);
buf BUF1 (N25, N17);
and AND3 (N26, N23, N1, N4);
and AND4 (N27, N8, N11, N19, N20);
nor NOR2 (N28, N25, N10);
buf BUF1 (N29, N11);
nand NAND2 (N30, N3, N24);
or OR3 (N31, N24, N3, N28);
and AND3 (N32, N26, N10, N25);
or OR2 (N33, N23, N18);
buf BUF1 (N34, N4);
not NOT1 (N35, N12);
nand NAND4 (N36, N4, N11, N14, N35);
nand NAND4 (N37, N2, N26, N31, N3);
nand NAND2 (N38, N17, N4);
or OR3 (N39, N2, N9, N35);
buf BUF1 (N40, N38);
not NOT1 (N41, N30);
nor NOR2 (N42, N34, N21);
and AND3 (N43, N29, N31, N20);
or OR3 (N44, N40, N41, N36);
buf BUF1 (N45, N28);
xor XOR2 (N46, N34, N26);
nand NAND2 (N47, N46, N44);
nand NAND4 (N48, N8, N23, N24, N33);
nor NOR4 (N49, N46, N15, N36, N18);
nor NOR2 (N50, N49, N15);
nand NAND4 (N51, N42, N46, N8, N6);
xor XOR2 (N52, N43, N43);
nor NOR4 (N53, N51, N12, N4, N2);
nor NOR3 (N54, N52, N46, N15);
not NOT1 (N55, N47);
not NOT1 (N56, N50);
buf BUF1 (N57, N27);
nand NAND3 (N58, N48, N31, N17);
xor XOR2 (N59, N39, N49);
xor XOR2 (N60, N37, N39);
nand NAND4 (N61, N53, N28, N46, N1);
buf BUF1 (N62, N59);
xor XOR2 (N63, N54, N2);
or OR2 (N64, N57, N59);
buf BUF1 (N65, N61);
nand NAND2 (N66, N55, N16);
or OR4 (N67, N58, N28, N44, N10);
or OR4 (N68, N62, N18, N13, N39);
xor XOR2 (N69, N68, N28);
buf BUF1 (N70, N65);
nor NOR3 (N71, N66, N52, N31);
nor NOR4 (N72, N45, N53, N3, N21);
buf BUF1 (N73, N60);
nor NOR4 (N74, N72, N26, N67, N28);
nand NAND4 (N75, N3, N14, N72, N51);
nor NOR4 (N76, N56, N6, N5, N33);
and AND2 (N77, N70, N22);
xor XOR2 (N78, N63, N40);
and AND3 (N79, N78, N39, N9);
or OR3 (N80, N64, N32, N42);
not NOT1 (N81, N43);
nor NOR3 (N82, N69, N56, N20);
nor NOR3 (N83, N76, N71, N56);
xor XOR2 (N84, N66, N33);
and AND2 (N85, N75, N12);
nand NAND2 (N86, N83, N24);
nor NOR4 (N87, N73, N12, N50, N64);
xor XOR2 (N88, N81, N67);
nand NAND2 (N89, N80, N54);
nor NOR3 (N90, N79, N63, N42);
and AND3 (N91, N90, N82, N75);
buf BUF1 (N92, N58);
xor XOR2 (N93, N87, N55);
and AND4 (N94, N89, N68, N52, N56);
xor XOR2 (N95, N94, N36);
nor NOR4 (N96, N85, N90, N48, N72);
xor XOR2 (N97, N77, N14);
and AND2 (N98, N74, N43);
nand NAND2 (N99, N91, N52);
nor NOR4 (N100, N86, N18, N64, N61);
or OR2 (N101, N95, N92);
and AND4 (N102, N72, N1, N8, N47);
nor NOR3 (N103, N98, N54, N12);
nor NOR2 (N104, N101, N82);
nor NOR4 (N105, N93, N28, N43, N48);
and AND2 (N106, N96, N48);
and AND4 (N107, N99, N85, N30, N30);
and AND3 (N108, N102, N40, N76);
nor NOR3 (N109, N97, N44, N53);
nor NOR2 (N110, N84, N48);
xor XOR2 (N111, N104, N43);
or OR2 (N112, N106, N8);
xor XOR2 (N113, N103, N21);
nor NOR2 (N114, N108, N20);
nand NAND4 (N115, N114, N50, N26, N22);
or OR4 (N116, N109, N32, N43, N99);
nor NOR4 (N117, N111, N70, N50, N47);
buf BUF1 (N118, N100);
xor XOR2 (N119, N112, N60);
buf BUF1 (N120, N115);
and AND3 (N121, N88, N18, N118);
not NOT1 (N122, N67);
or OR3 (N123, N110, N47, N93);
not NOT1 (N124, N119);
and AND4 (N125, N122, N84, N119, N69);
or OR2 (N126, N105, N38);
nor NOR4 (N127, N124, N56, N39, N98);
nor NOR3 (N128, N123, N112, N11);
nor NOR2 (N129, N121, N12);
not NOT1 (N130, N128);
buf BUF1 (N131, N125);
and AND2 (N132, N120, N7);
buf BUF1 (N133, N131);
nand NAND3 (N134, N132, N86, N30);
nor NOR3 (N135, N113, N29, N75);
not NOT1 (N136, N107);
nand NAND4 (N137, N134, N124, N2, N59);
nand NAND4 (N138, N129, N124, N86, N110);
nand NAND4 (N139, N116, N9, N122, N96);
nor NOR3 (N140, N136, N14, N66);
buf BUF1 (N141, N133);
nand NAND2 (N142, N130, N26);
buf BUF1 (N143, N126);
nand NAND3 (N144, N138, N54, N87);
or OR2 (N145, N127, N121);
and AND3 (N146, N137, N1, N118);
and AND2 (N147, N143, N146);
buf BUF1 (N148, N75);
not NOT1 (N149, N117);
xor XOR2 (N150, N142, N119);
and AND4 (N151, N149, N114, N64, N39);
and AND2 (N152, N140, N34);
not NOT1 (N153, N144);
or OR2 (N154, N141, N58);
not NOT1 (N155, N150);
or OR4 (N156, N152, N59, N2, N94);
and AND2 (N157, N156, N58);
nand NAND2 (N158, N153, N140);
xor XOR2 (N159, N151, N49);
nor NOR4 (N160, N155, N109, N57, N153);
not NOT1 (N161, N145);
nand NAND3 (N162, N139, N5, N156);
nand NAND3 (N163, N159, N123, N89);
nand NAND2 (N164, N162, N78);
xor XOR2 (N165, N148, N36);
xor XOR2 (N166, N154, N17);
not NOT1 (N167, N147);
buf BUF1 (N168, N158);
buf BUF1 (N169, N135);
nor NOR4 (N170, N157, N12, N31, N86);
xor XOR2 (N171, N160, N83);
and AND3 (N172, N163, N36, N49);
and AND4 (N173, N161, N111, N164, N54);
and AND2 (N174, N56, N11);
or OR4 (N175, N167, N121, N69, N105);
buf BUF1 (N176, N174);
nand NAND2 (N177, N171, N105);
and AND2 (N178, N177, N125);
not NOT1 (N179, N169);
nor NOR3 (N180, N165, N39, N97);
nor NOR2 (N181, N175, N171);
nand NAND4 (N182, N168, N33, N151, N37);
nand NAND2 (N183, N182, N29);
and AND3 (N184, N179, N139, N161);
or OR2 (N185, N178, N133);
and AND4 (N186, N184, N158, N153, N56);
and AND4 (N187, N181, N3, N22, N92);
nor NOR3 (N188, N173, N74, N36);
nand NAND3 (N189, N180, N179, N184);
and AND3 (N190, N170, N154, N172);
nor NOR3 (N191, N138, N132, N92);
and AND4 (N192, N176, N118, N117, N72);
xor XOR2 (N193, N166, N75);
buf BUF1 (N194, N185);
not NOT1 (N195, N194);
and AND4 (N196, N186, N81, N75, N10);
buf BUF1 (N197, N191);
and AND4 (N198, N183, N119, N174, N66);
xor XOR2 (N199, N198, N178);
nor NOR2 (N200, N190, N103);
not NOT1 (N201, N187);
or OR4 (N202, N188, N152, N199, N106);
not NOT1 (N203, N103);
xor XOR2 (N204, N200, N79);
xor XOR2 (N205, N189, N6);
nand NAND3 (N206, N196, N204, N80);
nand NAND2 (N207, N39, N160);
not NOT1 (N208, N202);
and AND3 (N209, N205, N156, N134);
or OR2 (N210, N192, N100);
or OR4 (N211, N209, N129, N175, N145);
not NOT1 (N212, N201);
nor NOR4 (N213, N211, N205, N12, N141);
buf BUF1 (N214, N213);
or OR3 (N215, N206, N13, N147);
nand NAND2 (N216, N210, N58);
buf BUF1 (N217, N212);
nor NOR4 (N218, N207, N175, N2, N189);
and AND3 (N219, N193, N23, N163);
not NOT1 (N220, N214);
buf BUF1 (N221, N215);
nand NAND3 (N222, N195, N127, N160);
and AND3 (N223, N217, N18, N178);
xor XOR2 (N224, N218, N153);
xor XOR2 (N225, N216, N133);
buf BUF1 (N226, N221);
nor NOR3 (N227, N197, N54, N81);
and AND3 (N228, N220, N38, N9);
buf BUF1 (N229, N219);
nor NOR4 (N230, N208, N20, N74, N20);
nor NOR3 (N231, N224, N59, N69);
or OR2 (N232, N230, N65);
nand NAND2 (N233, N229, N129);
xor XOR2 (N234, N203, N3);
xor XOR2 (N235, N225, N45);
or OR3 (N236, N234, N47, N181);
nor NOR2 (N237, N222, N61);
nor NOR4 (N238, N232, N111, N169, N150);
nand NAND4 (N239, N238, N181, N39, N139);
not NOT1 (N240, N228);
and AND2 (N241, N240, N197);
nand NAND3 (N242, N236, N158, N82);
or OR3 (N243, N242, N121, N158);
nor NOR2 (N244, N233, N30);
and AND2 (N245, N244, N77);
buf BUF1 (N246, N237);
buf BUF1 (N247, N239);
xor XOR2 (N248, N246, N231);
buf BUF1 (N249, N199);
or OR3 (N250, N248, N213, N191);
nand NAND2 (N251, N235, N205);
not NOT1 (N252, N247);
not NOT1 (N253, N251);
not NOT1 (N254, N250);
buf BUF1 (N255, N241);
and AND2 (N256, N226, N117);
nand NAND3 (N257, N223, N157, N63);
buf BUF1 (N258, N253);
buf BUF1 (N259, N245);
nor NOR4 (N260, N256, N53, N226, N169);
buf BUF1 (N261, N252);
xor XOR2 (N262, N259, N169);
not NOT1 (N263, N260);
buf BUF1 (N264, N262);
not NOT1 (N265, N249);
not NOT1 (N266, N263);
buf BUF1 (N267, N264);
nand NAND2 (N268, N265, N173);
or OR4 (N269, N254, N21, N250, N163);
buf BUF1 (N270, N227);
nor NOR4 (N271, N258, N133, N7, N182);
buf BUF1 (N272, N271);
not NOT1 (N273, N268);
not NOT1 (N274, N261);
and AND4 (N275, N273, N79, N264, N36);
buf BUF1 (N276, N255);
not NOT1 (N277, N257);
or OR3 (N278, N270, N214, N41);
not NOT1 (N279, N275);
nor NOR3 (N280, N266, N159, N166);
nand NAND2 (N281, N267, N78);
not NOT1 (N282, N280);
nor NOR4 (N283, N278, N212, N78, N134);
nor NOR3 (N284, N276, N213, N230);
not NOT1 (N285, N282);
nand NAND4 (N286, N283, N226, N86, N220);
nand NAND2 (N287, N281, N112);
buf BUF1 (N288, N272);
buf BUF1 (N289, N277);
or OR2 (N290, N243, N224);
xor XOR2 (N291, N288, N131);
and AND4 (N292, N291, N157, N8, N188);
or OR3 (N293, N286, N14, N221);
not NOT1 (N294, N285);
nor NOR4 (N295, N274, N67, N187, N156);
nand NAND3 (N296, N290, N292, N21);
nand NAND4 (N297, N194, N25, N253, N274);
buf BUF1 (N298, N279);
xor XOR2 (N299, N294, N167);
buf BUF1 (N300, N284);
nor NOR3 (N301, N295, N208, N49);
or OR2 (N302, N300, N114);
xor XOR2 (N303, N287, N133);
buf BUF1 (N304, N269);
xor XOR2 (N305, N293, N174);
not NOT1 (N306, N297);
and AND3 (N307, N305, N199, N18);
nand NAND3 (N308, N299, N253, N307);
buf BUF1 (N309, N275);
buf BUF1 (N310, N309);
not NOT1 (N311, N298);
buf BUF1 (N312, N302);
buf BUF1 (N313, N311);
not NOT1 (N314, N303);
buf BUF1 (N315, N306);
nor NOR2 (N316, N304, N140);
or OR2 (N317, N296, N134);
buf BUF1 (N318, N310);
buf BUF1 (N319, N315);
nor NOR3 (N320, N316, N282, N127);
not NOT1 (N321, N289);
buf BUF1 (N322, N313);
nand NAND2 (N323, N301, N71);
not NOT1 (N324, N314);
nor NOR3 (N325, N324, N153, N160);
xor XOR2 (N326, N323, N16);
nand NAND2 (N327, N320, N235);
nor NOR4 (N328, N326, N62, N17, N324);
buf BUF1 (N329, N318);
xor XOR2 (N330, N308, N15);
buf BUF1 (N331, N312);
or OR4 (N332, N328, N61, N121, N94);
buf BUF1 (N333, N329);
or OR3 (N334, N333, N78, N156);
buf BUF1 (N335, N331);
nand NAND2 (N336, N325, N72);
xor XOR2 (N337, N322, N234);
buf BUF1 (N338, N319);
not NOT1 (N339, N317);
nand NAND3 (N340, N336, N22, N45);
nand NAND2 (N341, N337, N64);
and AND4 (N342, N340, N93, N152, N332);
xor XOR2 (N343, N132, N188);
and AND3 (N344, N335, N105, N64);
and AND4 (N345, N330, N328, N293, N230);
and AND3 (N346, N342, N118, N185);
and AND3 (N347, N344, N136, N236);
and AND3 (N348, N338, N95, N40);
xor XOR2 (N349, N346, N313);
buf BUF1 (N350, N341);
or OR4 (N351, N349, N53, N313, N303);
nand NAND3 (N352, N321, N139, N211);
nand NAND2 (N353, N352, N123);
xor XOR2 (N354, N345, N204);
or OR4 (N355, N351, N219, N172, N270);
and AND2 (N356, N353, N131);
not NOT1 (N357, N339);
buf BUF1 (N358, N356);
nor NOR4 (N359, N347, N268, N136, N87);
not NOT1 (N360, N327);
buf BUF1 (N361, N350);
xor XOR2 (N362, N348, N92);
buf BUF1 (N363, N357);
or OR2 (N364, N343, N128);
or OR3 (N365, N361, N113, N284);
and AND4 (N366, N334, N128, N114, N142);
nor NOR2 (N367, N364, N49);
buf BUF1 (N368, N355);
buf BUF1 (N369, N365);
or OR2 (N370, N369, N94);
not NOT1 (N371, N370);
not NOT1 (N372, N367);
xor XOR2 (N373, N368, N325);
nand NAND2 (N374, N372, N156);
or OR2 (N375, N371, N240);
or OR4 (N376, N358, N217, N198, N197);
and AND3 (N377, N360, N290, N178);
buf BUF1 (N378, N359);
and AND2 (N379, N377, N124);
not NOT1 (N380, N362);
not NOT1 (N381, N378);
nor NOR4 (N382, N366, N229, N64, N225);
or OR2 (N383, N374, N278);
or OR3 (N384, N381, N92, N160);
xor XOR2 (N385, N373, N158);
buf BUF1 (N386, N382);
nand NAND3 (N387, N384, N178, N148);
buf BUF1 (N388, N354);
xor XOR2 (N389, N379, N149);
xor XOR2 (N390, N388, N37);
and AND3 (N391, N390, N113, N39);
or OR4 (N392, N389, N143, N329, N99);
or OR3 (N393, N375, N386, N337);
nand NAND2 (N394, N236, N353);
not NOT1 (N395, N394);
nand NAND3 (N396, N391, N174, N210);
nor NOR2 (N397, N396, N72);
or OR3 (N398, N395, N195, N263);
nor NOR3 (N399, N376, N6, N198);
nor NOR2 (N400, N383, N244);
xor XOR2 (N401, N363, N105);
not NOT1 (N402, N385);
and AND4 (N403, N400, N383, N371, N266);
not NOT1 (N404, N403);
nor NOR2 (N405, N392, N155);
not NOT1 (N406, N398);
xor XOR2 (N407, N405, N157);
or OR2 (N408, N387, N15);
nor NOR2 (N409, N393, N133);
nand NAND2 (N410, N397, N385);
xor XOR2 (N411, N409, N119);
not NOT1 (N412, N408);
not NOT1 (N413, N410);
nor NOR2 (N414, N407, N293);
nand NAND3 (N415, N401, N158, N301);
not NOT1 (N416, N399);
nand NAND3 (N417, N402, N128, N81);
and AND3 (N418, N413, N186, N84);
endmodule