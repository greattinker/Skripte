// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16;

output N1493,N1515,N1503,N1468,N1504,N1508,N1507,N1509,N1492,N1516;

xor XOR2 (N17, N4, N11);
or OR3 (N18, N16, N2, N7);
xor XOR2 (N19, N6, N6);
and AND3 (N20, N15, N16, N19);
and AND4 (N21, N5, N9, N13, N5);
buf BUF1 (N22, N12);
xor XOR2 (N23, N4, N1);
nand NAND3 (N24, N11, N12, N20);
xor XOR2 (N25, N4, N17);
xor XOR2 (N26, N16, N11);
buf BUF1 (N27, N2);
or OR4 (N28, N3, N16, N23, N3);
buf BUF1 (N29, N22);
buf BUF1 (N30, N1);
not NOT1 (N31, N2);
nand NAND3 (N32, N21, N14, N11);
nor NOR4 (N33, N26, N32, N25, N5);
xor XOR2 (N34, N8, N12);
nor NOR4 (N35, N20, N9, N7, N5);
nand NAND4 (N36, N33, N19, N8, N21);
and AND4 (N37, N27, N10, N1, N9);
and AND2 (N38, N37, N4);
or OR2 (N39, N28, N6);
nand NAND2 (N40, N39, N1);
nor NOR4 (N41, N18, N3, N12, N33);
buf BUF1 (N42, N36);
nand NAND4 (N43, N38, N19, N42, N39);
nand NAND4 (N44, N36, N3, N20, N43);
nand NAND2 (N45, N6, N35);
nand NAND4 (N46, N33, N14, N38, N14);
or OR4 (N47, N34, N44, N42, N21);
nor NOR2 (N48, N29, N6);
or OR4 (N49, N45, N42, N23, N46);
and AND4 (N50, N40, N36, N8, N3);
not NOT1 (N51, N6);
xor XOR2 (N52, N13, N38);
not NOT1 (N53, N41);
or OR2 (N54, N47, N19);
and AND3 (N55, N31, N41, N28);
nor NOR4 (N56, N49, N48, N54, N31);
not NOT1 (N57, N14);
buf BUF1 (N58, N28);
nand NAND3 (N59, N52, N22, N6);
not NOT1 (N60, N24);
or OR4 (N61, N56, N7, N28, N18);
and AND2 (N62, N50, N55);
not NOT1 (N63, N21);
nor NOR4 (N64, N30, N19, N19, N60);
not NOT1 (N65, N44);
xor XOR2 (N66, N61, N31);
nand NAND3 (N67, N65, N8, N37);
xor XOR2 (N68, N66, N34);
nand NAND2 (N69, N53, N13);
buf BUF1 (N70, N64);
or OR4 (N71, N51, N42, N58, N58);
or OR2 (N72, N54, N70);
not NOT1 (N73, N38);
nand NAND4 (N74, N68, N13, N21, N66);
and AND2 (N75, N59, N61);
nand NAND2 (N76, N57, N62);
xor XOR2 (N77, N74, N62);
xor XOR2 (N78, N57, N55);
and AND2 (N79, N76, N62);
buf BUF1 (N80, N79);
buf BUF1 (N81, N63);
and AND3 (N82, N78, N14, N78);
nor NOR4 (N83, N77, N62, N23, N33);
and AND3 (N84, N83, N10, N59);
and AND3 (N85, N69, N48, N22);
and AND2 (N86, N84, N75);
nand NAND4 (N87, N79, N83, N53, N67);
xor XOR2 (N88, N26, N6);
not NOT1 (N89, N72);
buf BUF1 (N90, N87);
or OR3 (N91, N90, N44, N45);
and AND4 (N92, N71, N2, N17, N83);
buf BUF1 (N93, N89);
not NOT1 (N94, N93);
or OR2 (N95, N80, N25);
xor XOR2 (N96, N86, N58);
not NOT1 (N97, N73);
buf BUF1 (N98, N82);
nand NAND2 (N99, N92, N34);
xor XOR2 (N100, N96, N94);
nand NAND2 (N101, N88, N30);
nor NOR2 (N102, N4, N17);
or OR2 (N103, N95, N39);
and AND3 (N104, N102, N80, N11);
or OR3 (N105, N85, N29, N70);
nor NOR4 (N106, N97, N49, N82, N39);
buf BUF1 (N107, N104);
xor XOR2 (N108, N107, N72);
not NOT1 (N109, N108);
and AND4 (N110, N81, N40, N48, N50);
or OR4 (N111, N100, N62, N37, N87);
nor NOR3 (N112, N99, N89, N99);
xor XOR2 (N113, N103, N79);
nor NOR3 (N114, N98, N45, N13);
buf BUF1 (N115, N113);
nand NAND3 (N116, N109, N89, N36);
nand NAND4 (N117, N111, N86, N81, N57);
and AND3 (N118, N112, N55, N115);
buf BUF1 (N119, N74);
xor XOR2 (N120, N116, N70);
nor NOR3 (N121, N91, N68, N57);
nor NOR2 (N122, N121, N54);
xor XOR2 (N123, N117, N48);
or OR3 (N124, N106, N25, N57);
not NOT1 (N125, N119);
not NOT1 (N126, N120);
not NOT1 (N127, N105);
or OR4 (N128, N110, N25, N51, N6);
not NOT1 (N129, N124);
nor NOR2 (N130, N118, N118);
nor NOR2 (N131, N101, N99);
or OR4 (N132, N129, N98, N72, N74);
not NOT1 (N133, N132);
nor NOR2 (N134, N122, N111);
or OR2 (N135, N131, N42);
nand NAND2 (N136, N130, N43);
xor XOR2 (N137, N125, N51);
nand NAND2 (N138, N126, N137);
and AND3 (N139, N117, N63, N17);
or OR3 (N140, N127, N75, N101);
nor NOR4 (N141, N138, N120, N5, N136);
xor XOR2 (N142, N13, N11);
and AND2 (N143, N114, N1);
and AND3 (N144, N128, N131, N86);
nor NOR2 (N145, N123, N65);
not NOT1 (N146, N144);
and AND3 (N147, N135, N101, N87);
nand NAND4 (N148, N145, N31, N138, N80);
or OR3 (N149, N141, N8, N68);
or OR3 (N150, N133, N111, N74);
not NOT1 (N151, N134);
not NOT1 (N152, N150);
and AND4 (N153, N147, N150, N94, N64);
nor NOR2 (N154, N142, N119);
xor XOR2 (N155, N149, N141);
and AND2 (N156, N146, N42);
buf BUF1 (N157, N139);
xor XOR2 (N158, N152, N69);
nand NAND2 (N159, N158, N112);
and AND2 (N160, N159, N69);
xor XOR2 (N161, N151, N147);
buf BUF1 (N162, N154);
or OR2 (N163, N155, N100);
xor XOR2 (N164, N160, N62);
buf BUF1 (N165, N143);
or OR2 (N166, N140, N145);
not NOT1 (N167, N165);
nand NAND2 (N168, N156, N143);
xor XOR2 (N169, N164, N11);
buf BUF1 (N170, N168);
or OR3 (N171, N170, N128, N153);
and AND3 (N172, N82, N21, N157);
nand NAND3 (N173, N154, N96, N13);
xor XOR2 (N174, N161, N92);
or OR4 (N175, N162, N171, N110, N113);
and AND2 (N176, N95, N86);
xor XOR2 (N177, N173, N58);
buf BUF1 (N178, N172);
not NOT1 (N179, N148);
xor XOR2 (N180, N166, N47);
xor XOR2 (N181, N175, N6);
not NOT1 (N182, N181);
xor XOR2 (N183, N178, N45);
or OR4 (N184, N182, N158, N122, N56);
not NOT1 (N185, N180);
buf BUF1 (N186, N179);
xor XOR2 (N187, N169, N120);
not NOT1 (N188, N183);
nand NAND2 (N189, N174, N27);
and AND2 (N190, N186, N113);
nor NOR2 (N191, N189, N66);
nand NAND4 (N192, N188, N61, N113, N150);
and AND3 (N193, N191, N136, N23);
or OR2 (N194, N192, N158);
buf BUF1 (N195, N177);
xor XOR2 (N196, N190, N19);
not NOT1 (N197, N195);
xor XOR2 (N198, N193, N172);
nand NAND3 (N199, N196, N109, N165);
or OR4 (N200, N199, N54, N108, N26);
and AND4 (N201, N167, N106, N114, N15);
not NOT1 (N202, N185);
nand NAND4 (N203, N187, N80, N147, N70);
nor NOR2 (N204, N194, N118);
not NOT1 (N205, N176);
nand NAND4 (N206, N197, N151, N44, N12);
nor NOR4 (N207, N203, N79, N171, N83);
and AND2 (N208, N200, N83);
or OR3 (N209, N206, N130, N153);
buf BUF1 (N210, N204);
xor XOR2 (N211, N202, N72);
not NOT1 (N212, N209);
buf BUF1 (N213, N163);
nand NAND2 (N214, N213, N116);
nor NOR3 (N215, N201, N100, N60);
and AND4 (N216, N212, N78, N33, N46);
or OR3 (N217, N216, N136, N28);
or OR2 (N218, N210, N20);
xor XOR2 (N219, N205, N148);
nand NAND4 (N220, N211, N47, N32, N134);
nand NAND3 (N221, N214, N4, N161);
or OR4 (N222, N207, N213, N32, N202);
or OR2 (N223, N222, N23);
not NOT1 (N224, N223);
buf BUF1 (N225, N208);
and AND4 (N226, N184, N49, N161, N132);
not NOT1 (N227, N219);
buf BUF1 (N228, N221);
xor XOR2 (N229, N215, N11);
not NOT1 (N230, N198);
buf BUF1 (N231, N227);
nand NAND3 (N232, N228, N129, N11);
and AND4 (N233, N229, N135, N12, N46);
or OR3 (N234, N217, N56, N206);
and AND2 (N235, N232, N202);
nand NAND4 (N236, N226, N184, N161, N21);
or OR4 (N237, N231, N62, N28, N170);
not NOT1 (N238, N218);
buf BUF1 (N239, N225);
or OR2 (N240, N234, N85);
buf BUF1 (N241, N224);
or OR3 (N242, N237, N136, N88);
nand NAND3 (N243, N220, N30, N236);
or OR4 (N244, N232, N59, N214, N8);
nand NAND3 (N245, N241, N79, N164);
or OR3 (N246, N242, N188, N51);
and AND4 (N247, N240, N176, N121, N38);
and AND3 (N248, N243, N160, N97);
and AND2 (N249, N245, N6);
not NOT1 (N250, N248);
buf BUF1 (N251, N250);
and AND3 (N252, N233, N67, N78);
nand NAND4 (N253, N246, N20, N166, N238);
and AND3 (N254, N252, N141, N69);
nand NAND4 (N255, N251, N196, N200, N219);
xor XOR2 (N256, N63, N15);
buf BUF1 (N257, N249);
or OR2 (N258, N256, N193);
buf BUF1 (N259, N230);
nand NAND2 (N260, N257, N188);
nand NAND4 (N261, N258, N144, N148, N117);
not NOT1 (N262, N259);
buf BUF1 (N263, N260);
and AND2 (N264, N247, N219);
and AND2 (N265, N255, N93);
or OR2 (N266, N263, N117);
buf BUF1 (N267, N262);
buf BUF1 (N268, N266);
nand NAND3 (N269, N265, N58, N59);
and AND3 (N270, N235, N36, N182);
and AND2 (N271, N254, N240);
xor XOR2 (N272, N244, N251);
or OR4 (N273, N239, N6, N93, N10);
buf BUF1 (N274, N270);
not NOT1 (N275, N261);
nand NAND3 (N276, N264, N49, N142);
not NOT1 (N277, N271);
nand NAND2 (N278, N272, N153);
or OR3 (N279, N268, N83, N16);
and AND4 (N280, N276, N83, N117, N21);
and AND4 (N281, N280, N163, N252, N250);
and AND3 (N282, N278, N278, N173);
xor XOR2 (N283, N253, N278);
and AND2 (N284, N275, N8);
and AND2 (N285, N267, N162);
nand NAND4 (N286, N273, N269, N209, N25);
or OR4 (N287, N168, N243, N146, N95);
not NOT1 (N288, N282);
not NOT1 (N289, N283);
and AND2 (N290, N279, N100);
nor NOR4 (N291, N274, N10, N33, N34);
or OR4 (N292, N284, N120, N218, N253);
not NOT1 (N293, N290);
xor XOR2 (N294, N291, N235);
nand NAND2 (N295, N277, N173);
nand NAND2 (N296, N292, N125);
or OR4 (N297, N294, N173, N211, N243);
not NOT1 (N298, N281);
or OR4 (N299, N286, N137, N209, N257);
nor NOR4 (N300, N295, N206, N39, N155);
xor XOR2 (N301, N296, N240);
and AND2 (N302, N300, N257);
and AND4 (N303, N302, N136, N51, N39);
or OR4 (N304, N285, N283, N40, N117);
not NOT1 (N305, N299);
or OR4 (N306, N293, N286, N94, N252);
or OR2 (N307, N305, N255);
nor NOR2 (N308, N288, N14);
not NOT1 (N309, N304);
or OR4 (N310, N289, N87, N60, N119);
nand NAND3 (N311, N298, N22, N57);
and AND2 (N312, N303, N73);
nand NAND3 (N313, N297, N287, N268);
buf BUF1 (N314, N95);
nand NAND3 (N315, N310, N80, N74);
not NOT1 (N316, N309);
not NOT1 (N317, N313);
nand NAND3 (N318, N306, N317, N105);
and AND2 (N319, N64, N156);
not NOT1 (N320, N312);
buf BUF1 (N321, N318);
nand NAND2 (N322, N301, N23);
nor NOR4 (N323, N320, N222, N140, N32);
buf BUF1 (N324, N308);
or OR4 (N325, N319, N50, N210, N324);
buf BUF1 (N326, N186);
xor XOR2 (N327, N326, N283);
and AND3 (N328, N307, N97, N240);
buf BUF1 (N329, N323);
and AND4 (N330, N315, N166, N104, N32);
nor NOR2 (N331, N314, N288);
nor NOR4 (N332, N328, N303, N36, N104);
not NOT1 (N333, N321);
nor NOR2 (N334, N331, N44);
buf BUF1 (N335, N334);
nand NAND3 (N336, N332, N121, N68);
buf BUF1 (N337, N336);
not NOT1 (N338, N322);
and AND3 (N339, N325, N319, N63);
not NOT1 (N340, N338);
nand NAND4 (N341, N316, N40, N254, N223);
nand NAND4 (N342, N341, N308, N144, N115);
and AND4 (N343, N340, N99, N280, N178);
xor XOR2 (N344, N339, N35);
and AND3 (N345, N337, N145, N117);
xor XOR2 (N346, N343, N74);
nor NOR4 (N347, N345, N227, N103, N36);
nand NAND4 (N348, N335, N148, N106, N185);
buf BUF1 (N349, N347);
and AND4 (N350, N346, N64, N294, N177);
xor XOR2 (N351, N344, N292);
buf BUF1 (N352, N327);
nor NOR2 (N353, N330, N59);
buf BUF1 (N354, N351);
not NOT1 (N355, N354);
nor NOR2 (N356, N311, N56);
or OR2 (N357, N329, N70);
not NOT1 (N358, N356);
xor XOR2 (N359, N353, N313);
nor NOR3 (N360, N355, N209, N248);
not NOT1 (N361, N352);
buf BUF1 (N362, N357);
and AND3 (N363, N342, N83, N271);
or OR4 (N364, N350, N66, N269, N286);
or OR3 (N365, N360, N192, N162);
buf BUF1 (N366, N359);
nor NOR2 (N367, N348, N322);
or OR3 (N368, N367, N98, N113);
buf BUF1 (N369, N362);
not NOT1 (N370, N366);
buf BUF1 (N371, N370);
and AND2 (N372, N333, N225);
buf BUF1 (N373, N371);
buf BUF1 (N374, N349);
nor NOR4 (N375, N373, N26, N116, N167);
buf BUF1 (N376, N363);
nor NOR2 (N377, N364, N214);
nor NOR3 (N378, N377, N203, N333);
xor XOR2 (N379, N368, N339);
xor XOR2 (N380, N375, N313);
buf BUF1 (N381, N361);
buf BUF1 (N382, N365);
not NOT1 (N383, N369);
and AND3 (N384, N372, N8, N27);
xor XOR2 (N385, N384, N349);
or OR4 (N386, N380, N230, N187, N5);
not NOT1 (N387, N383);
xor XOR2 (N388, N379, N123);
and AND2 (N389, N374, N3);
buf BUF1 (N390, N381);
or OR4 (N391, N385, N216, N125, N195);
nor NOR4 (N392, N386, N297, N262, N142);
xor XOR2 (N393, N382, N3);
nand NAND3 (N394, N387, N99, N350);
buf BUF1 (N395, N393);
nand NAND3 (N396, N388, N99, N263);
buf BUF1 (N397, N391);
buf BUF1 (N398, N358);
nor NOR3 (N399, N378, N111, N90);
nand NAND2 (N400, N394, N128);
and AND4 (N401, N400, N238, N95, N262);
xor XOR2 (N402, N392, N150);
not NOT1 (N403, N376);
not NOT1 (N404, N389);
and AND4 (N405, N401, N142, N384, N291);
buf BUF1 (N406, N395);
nand NAND4 (N407, N403, N348, N252, N170);
not NOT1 (N408, N406);
buf BUF1 (N409, N405);
nand NAND4 (N410, N397, N57, N286, N234);
not NOT1 (N411, N407);
or OR2 (N412, N396, N288);
or OR4 (N413, N398, N302, N136, N52);
buf BUF1 (N414, N402);
or OR3 (N415, N409, N254, N274);
and AND2 (N416, N408, N186);
or OR3 (N417, N399, N280, N94);
nand NAND3 (N418, N416, N326, N291);
nor NOR2 (N419, N417, N288);
and AND3 (N420, N390, N237, N387);
not NOT1 (N421, N418);
xor XOR2 (N422, N404, N58);
xor XOR2 (N423, N419, N63);
buf BUF1 (N424, N413);
or OR2 (N425, N411, N42);
xor XOR2 (N426, N423, N60);
not NOT1 (N427, N420);
xor XOR2 (N428, N412, N156);
nor NOR3 (N429, N421, N296, N315);
nor NOR2 (N430, N425, N370);
and AND4 (N431, N427, N363, N396, N160);
not NOT1 (N432, N430);
buf BUF1 (N433, N424);
and AND4 (N434, N433, N63, N255, N153);
or OR2 (N435, N432, N273);
xor XOR2 (N436, N434, N357);
or OR2 (N437, N410, N255);
and AND3 (N438, N422, N67, N293);
not NOT1 (N439, N431);
nand NAND3 (N440, N426, N305, N178);
nor NOR4 (N441, N414, N117, N298, N283);
and AND2 (N442, N441, N336);
not NOT1 (N443, N439);
not NOT1 (N444, N438);
nor NOR2 (N445, N429, N310);
and AND2 (N446, N440, N434);
nand NAND2 (N447, N446, N120);
nor NOR2 (N448, N436, N244);
nand NAND2 (N449, N448, N259);
or OR4 (N450, N437, N60, N321, N413);
or OR3 (N451, N442, N105, N378);
and AND3 (N452, N450, N353, N281);
and AND2 (N453, N449, N83);
nor NOR4 (N454, N447, N149, N241, N60);
not NOT1 (N455, N445);
not NOT1 (N456, N454);
buf BUF1 (N457, N455);
not NOT1 (N458, N415);
not NOT1 (N459, N443);
or OR2 (N460, N457, N243);
buf BUF1 (N461, N451);
nand NAND4 (N462, N461, N407, N33, N274);
not NOT1 (N463, N462);
xor XOR2 (N464, N459, N348);
xor XOR2 (N465, N428, N357);
nor NOR3 (N466, N453, N38, N101);
or OR2 (N467, N435, N136);
and AND3 (N468, N467, N166, N392);
buf BUF1 (N469, N468);
xor XOR2 (N470, N466, N205);
and AND2 (N471, N470, N75);
nor NOR2 (N472, N460, N62);
nand NAND3 (N473, N469, N433, N428);
nor NOR2 (N474, N471, N225);
or OR2 (N475, N464, N190);
buf BUF1 (N476, N472);
xor XOR2 (N477, N465, N61);
nor NOR3 (N478, N463, N393, N466);
and AND4 (N479, N476, N214, N105, N99);
not NOT1 (N480, N474);
xor XOR2 (N481, N452, N121);
not NOT1 (N482, N444);
nand NAND2 (N483, N473, N191);
nor NOR3 (N484, N478, N390, N46);
nand NAND3 (N485, N484, N372, N42);
nor NOR2 (N486, N482, N79);
xor XOR2 (N487, N479, N251);
not NOT1 (N488, N458);
xor XOR2 (N489, N477, N246);
or OR4 (N490, N488, N272, N400, N401);
or OR2 (N491, N490, N436);
nand NAND2 (N492, N483, N158);
not NOT1 (N493, N481);
nor NOR3 (N494, N493, N75, N247);
or OR3 (N495, N486, N94, N95);
nor NOR2 (N496, N494, N442);
and AND2 (N497, N489, N253);
nor NOR2 (N498, N491, N427);
xor XOR2 (N499, N456, N149);
and AND4 (N500, N499, N428, N392, N415);
buf BUF1 (N501, N497);
not NOT1 (N502, N485);
not NOT1 (N503, N475);
xor XOR2 (N504, N480, N97);
buf BUF1 (N505, N487);
nand NAND4 (N506, N505, N383, N273, N128);
xor XOR2 (N507, N495, N402);
nand NAND3 (N508, N492, N417, N491);
and AND4 (N509, N504, N422, N25, N69);
buf BUF1 (N510, N496);
and AND2 (N511, N501, N322);
buf BUF1 (N512, N498);
and AND3 (N513, N508, N308, N280);
nand NAND4 (N514, N512, N380, N7, N338);
nor NOR2 (N515, N511, N316);
and AND3 (N516, N507, N58, N13);
and AND4 (N517, N502, N348, N398, N490);
buf BUF1 (N518, N517);
not NOT1 (N519, N509);
buf BUF1 (N520, N518);
not NOT1 (N521, N520);
nor NOR3 (N522, N514, N182, N236);
nand NAND3 (N523, N519, N348, N84);
buf BUF1 (N524, N516);
and AND3 (N525, N515, N235, N123);
nor NOR4 (N526, N523, N414, N32, N368);
and AND3 (N527, N510, N239, N276);
and AND4 (N528, N527, N287, N292, N241);
buf BUF1 (N529, N521);
or OR4 (N530, N506, N435, N226, N343);
and AND3 (N531, N522, N266, N173);
not NOT1 (N532, N530);
xor XOR2 (N533, N525, N143);
not NOT1 (N534, N533);
or OR3 (N535, N500, N101, N148);
nor NOR4 (N536, N532, N308, N223, N348);
nor NOR3 (N537, N534, N131, N497);
nor NOR3 (N538, N524, N389, N136);
buf BUF1 (N539, N538);
not NOT1 (N540, N529);
nand NAND3 (N541, N539, N290, N303);
nand NAND3 (N542, N540, N529, N174);
not NOT1 (N543, N531);
buf BUF1 (N544, N513);
not NOT1 (N545, N541);
nand NAND3 (N546, N503, N533, N321);
xor XOR2 (N547, N545, N546);
nor NOR3 (N548, N454, N452, N272);
nor NOR2 (N549, N544, N532);
xor XOR2 (N550, N542, N544);
not NOT1 (N551, N535);
xor XOR2 (N552, N536, N150);
or OR4 (N553, N543, N77, N524, N238);
not NOT1 (N554, N549);
nor NOR2 (N555, N528, N426);
and AND2 (N556, N555, N158);
xor XOR2 (N557, N550, N45);
buf BUF1 (N558, N554);
or OR3 (N559, N537, N339, N337);
or OR2 (N560, N553, N224);
nor NOR3 (N561, N526, N185, N87);
and AND2 (N562, N561, N414);
not NOT1 (N563, N556);
xor XOR2 (N564, N562, N36);
and AND3 (N565, N563, N405, N468);
not NOT1 (N566, N559);
buf BUF1 (N567, N547);
xor XOR2 (N568, N567, N552);
and AND2 (N569, N310, N543);
or OR2 (N570, N564, N244);
nand NAND4 (N571, N560, N401, N250, N503);
xor XOR2 (N572, N557, N277);
not NOT1 (N573, N548);
not NOT1 (N574, N571);
not NOT1 (N575, N570);
buf BUF1 (N576, N568);
nor NOR3 (N577, N572, N455, N387);
or OR3 (N578, N576, N434, N444);
nand NAND4 (N579, N575, N536, N577, N368);
nand NAND2 (N580, N263, N386);
xor XOR2 (N581, N579, N269);
nand NAND4 (N582, N565, N204, N171, N36);
not NOT1 (N583, N566);
nor NOR3 (N584, N573, N73, N32);
or OR4 (N585, N581, N514, N547, N144);
buf BUF1 (N586, N578);
not NOT1 (N587, N558);
buf BUF1 (N588, N587);
not NOT1 (N589, N583);
and AND3 (N590, N580, N42, N4);
buf BUF1 (N591, N584);
nor NOR4 (N592, N569, N510, N64, N424);
buf BUF1 (N593, N551);
buf BUF1 (N594, N586);
and AND2 (N595, N593, N93);
xor XOR2 (N596, N595, N349);
xor XOR2 (N597, N592, N516);
xor XOR2 (N598, N594, N431);
buf BUF1 (N599, N597);
and AND2 (N600, N585, N283);
nor NOR4 (N601, N590, N598, N198, N19);
nand NAND2 (N602, N300, N429);
buf BUF1 (N603, N591);
not NOT1 (N604, N582);
xor XOR2 (N605, N596, N437);
or OR4 (N606, N599, N254, N155, N60);
or OR3 (N607, N574, N601, N489);
or OR2 (N608, N14, N380);
xor XOR2 (N609, N604, N127);
buf BUF1 (N610, N588);
nand NAND2 (N611, N605, N335);
not NOT1 (N612, N608);
nand NAND3 (N613, N612, N367, N76);
nand NAND4 (N614, N602, N171, N166, N313);
nand NAND2 (N615, N606, N22);
and AND2 (N616, N603, N326);
and AND2 (N617, N614, N336);
or OR3 (N618, N617, N397, N264);
nand NAND3 (N619, N600, N82, N343);
buf BUF1 (N620, N615);
not NOT1 (N621, N613);
nor NOR3 (N622, N620, N271, N306);
buf BUF1 (N623, N621);
nand NAND2 (N624, N622, N24);
not NOT1 (N625, N611);
xor XOR2 (N626, N619, N34);
buf BUF1 (N627, N610);
buf BUF1 (N628, N625);
xor XOR2 (N629, N624, N333);
buf BUF1 (N630, N626);
xor XOR2 (N631, N628, N38);
not NOT1 (N632, N623);
nor NOR3 (N633, N631, N454, N394);
nand NAND2 (N634, N589, N51);
and AND4 (N635, N609, N271, N103, N300);
not NOT1 (N636, N627);
and AND2 (N637, N618, N291);
not NOT1 (N638, N637);
xor XOR2 (N639, N607, N576);
or OR2 (N640, N634, N569);
nor NOR4 (N641, N638, N605, N425, N50);
nand NAND3 (N642, N633, N251, N49);
or OR2 (N643, N641, N63);
and AND4 (N644, N616, N293, N111, N523);
xor XOR2 (N645, N644, N369);
nor NOR3 (N646, N642, N316, N206);
xor XOR2 (N647, N629, N269);
not NOT1 (N648, N647);
and AND2 (N649, N639, N254);
nand NAND4 (N650, N643, N221, N546, N181);
and AND2 (N651, N650, N504);
nor NOR2 (N652, N636, N434);
nand NAND2 (N653, N645, N367);
buf BUF1 (N654, N640);
xor XOR2 (N655, N651, N84);
and AND2 (N656, N652, N461);
xor XOR2 (N657, N655, N359);
not NOT1 (N658, N656);
nor NOR4 (N659, N646, N593, N63, N502);
not NOT1 (N660, N657);
buf BUF1 (N661, N635);
nand NAND2 (N662, N630, N190);
xor XOR2 (N663, N662, N579);
xor XOR2 (N664, N659, N87);
xor XOR2 (N665, N654, N184);
nor NOR4 (N666, N663, N375, N328, N289);
nor NOR3 (N667, N665, N618, N225);
buf BUF1 (N668, N648);
or OR4 (N669, N666, N142, N28, N81);
buf BUF1 (N670, N669);
buf BUF1 (N671, N632);
nand NAND3 (N672, N661, N624, N113);
not NOT1 (N673, N653);
nand NAND3 (N674, N672, N530, N188);
nand NAND2 (N675, N668, N399);
nor NOR2 (N676, N667, N195);
nand NAND3 (N677, N664, N240, N634);
and AND3 (N678, N671, N667, N182);
or OR2 (N679, N660, N497);
not NOT1 (N680, N677);
not NOT1 (N681, N676);
buf BUF1 (N682, N678);
nand NAND3 (N683, N680, N491, N203);
or OR2 (N684, N673, N650);
not NOT1 (N685, N675);
and AND4 (N686, N658, N297, N470, N373);
and AND2 (N687, N682, N62);
and AND3 (N688, N679, N30, N180);
nand NAND4 (N689, N684, N141, N536, N575);
and AND4 (N690, N683, N37, N292, N295);
nor NOR4 (N691, N687, N680, N169, N108);
nor NOR4 (N692, N670, N348, N573, N557);
not NOT1 (N693, N688);
or OR3 (N694, N693, N272, N383);
buf BUF1 (N695, N689);
or OR4 (N696, N674, N518, N449, N540);
xor XOR2 (N697, N694, N680);
nor NOR3 (N698, N681, N244, N132);
xor XOR2 (N699, N685, N667);
nand NAND4 (N700, N686, N231, N603, N130);
buf BUF1 (N701, N698);
or OR3 (N702, N691, N162, N231);
or OR4 (N703, N701, N217, N336, N657);
or OR4 (N704, N690, N428, N36, N169);
not NOT1 (N705, N702);
nand NAND3 (N706, N695, N385, N635);
or OR2 (N707, N649, N20);
nand NAND4 (N708, N703, N506, N183, N157);
or OR4 (N709, N708, N218, N499, N187);
nor NOR3 (N710, N692, N644, N121);
and AND2 (N711, N707, N404);
nor NOR3 (N712, N699, N239, N101);
nor NOR2 (N713, N712, N58);
not NOT1 (N714, N696);
and AND3 (N715, N700, N61, N111);
nor NOR4 (N716, N709, N581, N192, N676);
buf BUF1 (N717, N716);
or OR4 (N718, N711, N636, N642, N594);
and AND4 (N719, N704, N45, N451, N530);
xor XOR2 (N720, N705, N47);
and AND2 (N721, N720, N305);
nor NOR4 (N722, N697, N557, N626, N653);
buf BUF1 (N723, N717);
buf BUF1 (N724, N723);
xor XOR2 (N725, N724, N394);
nor NOR4 (N726, N715, N89, N209, N512);
nor NOR3 (N727, N719, N715, N16);
xor XOR2 (N728, N726, N680);
or OR4 (N729, N706, N269, N582, N638);
nor NOR4 (N730, N714, N295, N230, N353);
xor XOR2 (N731, N729, N430);
xor XOR2 (N732, N722, N701);
or OR2 (N733, N731, N584);
buf BUF1 (N734, N732);
buf BUF1 (N735, N733);
buf BUF1 (N736, N718);
nor NOR2 (N737, N736, N305);
buf BUF1 (N738, N730);
or OR3 (N739, N713, N486, N645);
xor XOR2 (N740, N727, N450);
nor NOR2 (N741, N721, N571);
buf BUF1 (N742, N728);
or OR3 (N743, N710, N668, N724);
buf BUF1 (N744, N741);
xor XOR2 (N745, N725, N397);
nand NAND3 (N746, N743, N417, N506);
and AND4 (N747, N734, N714, N524, N440);
and AND3 (N748, N744, N622, N289);
not NOT1 (N749, N745);
or OR4 (N750, N739, N83, N384, N324);
nor NOR2 (N751, N738, N42);
buf BUF1 (N752, N740);
not NOT1 (N753, N749);
nor NOR4 (N754, N737, N747, N691, N700);
or OR3 (N755, N642, N503, N693);
nand NAND2 (N756, N746, N302);
nand NAND3 (N757, N754, N536, N111);
nor NOR3 (N758, N735, N445, N299);
nand NAND4 (N759, N753, N441, N668, N712);
and AND4 (N760, N758, N225, N470, N636);
nand NAND3 (N761, N757, N112, N664);
nand NAND2 (N762, N756, N7);
not NOT1 (N763, N760);
or OR4 (N764, N742, N308, N414, N728);
nor NOR4 (N765, N750, N521, N484, N37);
buf BUF1 (N766, N755);
nor NOR2 (N767, N761, N306);
and AND4 (N768, N767, N737, N135, N423);
buf BUF1 (N769, N764);
xor XOR2 (N770, N762, N596);
xor XOR2 (N771, N752, N364);
or OR3 (N772, N751, N435, N487);
buf BUF1 (N773, N772);
xor XOR2 (N774, N768, N600);
buf BUF1 (N775, N748);
not NOT1 (N776, N773);
buf BUF1 (N777, N765);
not NOT1 (N778, N776);
nand NAND3 (N779, N769, N323, N644);
nand NAND3 (N780, N774, N395, N734);
not NOT1 (N781, N778);
nand NAND4 (N782, N759, N682, N127, N446);
or OR3 (N783, N781, N601, N271);
not NOT1 (N784, N779);
not NOT1 (N785, N784);
xor XOR2 (N786, N783, N593);
or OR4 (N787, N785, N758, N752, N138);
and AND2 (N788, N770, N301);
xor XOR2 (N789, N775, N409);
nor NOR3 (N790, N763, N633, N688);
or OR3 (N791, N790, N180, N731);
and AND2 (N792, N777, N733);
buf BUF1 (N793, N780);
or OR4 (N794, N793, N10, N102, N749);
buf BUF1 (N795, N786);
or OR4 (N796, N787, N475, N420, N146);
or OR3 (N797, N791, N682, N394);
nand NAND3 (N798, N789, N128, N338);
buf BUF1 (N799, N792);
nand NAND4 (N800, N799, N703, N405, N423);
buf BUF1 (N801, N800);
not NOT1 (N802, N796);
xor XOR2 (N803, N788, N443);
or OR2 (N804, N801, N431);
nand NAND4 (N805, N782, N548, N343, N171);
and AND4 (N806, N794, N236, N224, N76);
not NOT1 (N807, N802);
buf BUF1 (N808, N766);
nor NOR2 (N809, N803, N91);
not NOT1 (N810, N805);
buf BUF1 (N811, N795);
nor NOR2 (N812, N798, N176);
or OR3 (N813, N809, N806, N131);
nor NOR3 (N814, N387, N227, N801);
and AND3 (N815, N808, N85, N399);
and AND4 (N816, N813, N164, N772, N39);
xor XOR2 (N817, N804, N255);
buf BUF1 (N818, N771);
or OR2 (N819, N817, N603);
nand NAND4 (N820, N812, N439, N436, N390);
nand NAND2 (N821, N807, N419);
nor NOR2 (N822, N816, N44);
buf BUF1 (N823, N821);
buf BUF1 (N824, N822);
or OR2 (N825, N824, N513);
and AND2 (N826, N823, N628);
nor NOR2 (N827, N811, N320);
buf BUF1 (N828, N815);
or OR4 (N829, N825, N791, N15, N671);
nor NOR3 (N830, N827, N391, N569);
xor XOR2 (N831, N814, N739);
nand NAND3 (N832, N797, N97, N713);
not NOT1 (N833, N830);
buf BUF1 (N834, N826);
or OR4 (N835, N828, N385, N762, N515);
nor NOR3 (N836, N833, N745, N326);
buf BUF1 (N837, N829);
xor XOR2 (N838, N832, N15);
or OR3 (N839, N831, N118, N736);
not NOT1 (N840, N837);
not NOT1 (N841, N810);
xor XOR2 (N842, N820, N534);
xor XOR2 (N843, N839, N293);
nor NOR2 (N844, N842, N659);
nor NOR4 (N845, N843, N548, N556, N254);
or OR2 (N846, N818, N581);
not NOT1 (N847, N819);
nor NOR4 (N848, N845, N379, N76, N13);
or OR3 (N849, N847, N165, N273);
and AND4 (N850, N838, N348, N755, N223);
nor NOR2 (N851, N846, N498);
not NOT1 (N852, N840);
and AND4 (N853, N848, N5, N618, N103);
not NOT1 (N854, N853);
nor NOR4 (N855, N836, N376, N5, N304);
nor NOR4 (N856, N849, N26, N312, N482);
or OR4 (N857, N844, N3, N311, N235);
or OR4 (N858, N855, N390, N668, N189);
not NOT1 (N859, N850);
nor NOR2 (N860, N835, N770);
and AND4 (N861, N854, N387, N797, N341);
not NOT1 (N862, N841);
and AND4 (N863, N860, N267, N210, N6);
not NOT1 (N864, N863);
nand NAND3 (N865, N862, N125, N652);
nor NOR3 (N866, N856, N274, N19);
xor XOR2 (N867, N858, N191);
nand NAND4 (N868, N852, N617, N558, N274);
not NOT1 (N869, N867);
not NOT1 (N870, N865);
xor XOR2 (N871, N834, N863);
and AND3 (N872, N864, N473, N788);
nand NAND2 (N873, N859, N795);
xor XOR2 (N874, N870, N693);
or OR4 (N875, N869, N439, N395, N296);
or OR3 (N876, N875, N545, N639);
not NOT1 (N877, N851);
or OR3 (N878, N872, N145, N758);
buf BUF1 (N879, N873);
and AND3 (N880, N857, N876, N748);
nand NAND2 (N881, N281, N598);
nor NOR4 (N882, N879, N190, N589, N695);
and AND2 (N883, N871, N641);
nand NAND4 (N884, N882, N852, N689, N26);
or OR3 (N885, N881, N827, N456);
and AND3 (N886, N861, N659, N89);
xor XOR2 (N887, N868, N866);
nand NAND4 (N888, N772, N111, N112, N95);
nor NOR3 (N889, N888, N235, N588);
not NOT1 (N890, N884);
xor XOR2 (N891, N887, N619);
not NOT1 (N892, N878);
xor XOR2 (N893, N889, N127);
or OR2 (N894, N890, N440);
buf BUF1 (N895, N885);
or OR4 (N896, N886, N431, N322, N472);
not NOT1 (N897, N894);
nor NOR4 (N898, N877, N291, N166, N555);
nor NOR2 (N899, N895, N894);
nand NAND4 (N900, N893, N698, N265, N827);
nor NOR4 (N901, N891, N416, N116, N360);
and AND4 (N902, N892, N506, N293, N825);
nand NAND4 (N903, N883, N5, N321, N802);
and AND3 (N904, N897, N301, N555);
nand NAND4 (N905, N904, N765, N494, N522);
not NOT1 (N906, N898);
nand NAND4 (N907, N905, N753, N156, N618);
nor NOR4 (N908, N907, N741, N521, N574);
and AND4 (N909, N908, N460, N327, N543);
nor NOR4 (N910, N874, N323, N290, N804);
xor XOR2 (N911, N900, N694);
not NOT1 (N912, N910);
buf BUF1 (N913, N906);
xor XOR2 (N914, N911, N628);
not NOT1 (N915, N909);
nand NAND2 (N916, N902, N721);
or OR3 (N917, N914, N908, N51);
or OR2 (N918, N896, N66);
and AND3 (N919, N915, N698, N575);
nor NOR2 (N920, N917, N77);
buf BUF1 (N921, N899);
nand NAND4 (N922, N901, N560, N123, N442);
nand NAND2 (N923, N913, N523);
or OR3 (N924, N923, N210, N302);
nand NAND2 (N925, N920, N283);
xor XOR2 (N926, N921, N16);
and AND2 (N927, N925, N745);
and AND4 (N928, N880, N280, N711, N347);
or OR3 (N929, N903, N12, N473);
nand NAND2 (N930, N912, N612);
nand NAND4 (N931, N929, N689, N451, N443);
not NOT1 (N932, N930);
xor XOR2 (N933, N922, N330);
or OR4 (N934, N924, N378, N539, N262);
nor NOR3 (N935, N931, N526, N908);
and AND4 (N936, N927, N323, N449, N353);
nor NOR2 (N937, N916, N903);
and AND4 (N938, N933, N383, N293, N237);
or OR2 (N939, N918, N850);
xor XOR2 (N940, N939, N120);
nor NOR3 (N941, N938, N777, N176);
nor NOR4 (N942, N935, N930, N691, N547);
not NOT1 (N943, N919);
xor XOR2 (N944, N943, N46);
buf BUF1 (N945, N934);
nor NOR3 (N946, N941, N436, N36);
xor XOR2 (N947, N945, N13);
nor NOR4 (N948, N947, N921, N92, N931);
or OR3 (N949, N946, N624, N106);
nand NAND4 (N950, N942, N887, N81, N198);
and AND2 (N951, N940, N751);
or OR2 (N952, N937, N326);
xor XOR2 (N953, N928, N811);
or OR4 (N954, N951, N531, N35, N867);
and AND4 (N955, N952, N668, N810, N891);
or OR2 (N956, N944, N637);
xor XOR2 (N957, N949, N470);
and AND3 (N958, N948, N798, N664);
xor XOR2 (N959, N936, N545);
not NOT1 (N960, N932);
nand NAND4 (N961, N926, N426, N268, N601);
and AND3 (N962, N950, N260, N369);
nor NOR2 (N963, N953, N625);
buf BUF1 (N964, N962);
and AND2 (N965, N954, N790);
or OR4 (N966, N955, N741, N861, N40);
xor XOR2 (N967, N956, N730);
xor XOR2 (N968, N965, N887);
and AND3 (N969, N968, N385, N944);
buf BUF1 (N970, N963);
buf BUF1 (N971, N970);
buf BUF1 (N972, N969);
nand NAND3 (N973, N971, N768, N143);
or OR4 (N974, N957, N184, N932, N181);
or OR4 (N975, N973, N14, N358, N440);
buf BUF1 (N976, N964);
and AND2 (N977, N972, N82);
xor XOR2 (N978, N960, N887);
xor XOR2 (N979, N958, N666);
nand NAND2 (N980, N979, N386);
buf BUF1 (N981, N975);
and AND3 (N982, N966, N216, N371);
not NOT1 (N983, N974);
xor XOR2 (N984, N982, N664);
not NOT1 (N985, N981);
not NOT1 (N986, N985);
buf BUF1 (N987, N978);
and AND2 (N988, N984, N398);
nand NAND3 (N989, N977, N959, N23);
buf BUF1 (N990, N517);
not NOT1 (N991, N986);
nor NOR2 (N992, N983, N801);
or OR2 (N993, N990, N124);
buf BUF1 (N994, N992);
nor NOR2 (N995, N993, N294);
nand NAND2 (N996, N976, N461);
nand NAND4 (N997, N996, N352, N764, N153);
or OR3 (N998, N987, N86, N174);
nand NAND4 (N999, N961, N884, N28, N639);
and AND4 (N1000, N999, N208, N438, N496);
xor XOR2 (N1001, N1000, N920);
not NOT1 (N1002, N997);
buf BUF1 (N1003, N1001);
nor NOR3 (N1004, N967, N615, N600);
xor XOR2 (N1005, N989, N744);
or OR3 (N1006, N988, N319, N964);
nor NOR2 (N1007, N1004, N752);
or OR2 (N1008, N1003, N234);
not NOT1 (N1009, N1007);
not NOT1 (N1010, N994);
nor NOR2 (N1011, N991, N440);
xor XOR2 (N1012, N1005, N381);
and AND3 (N1013, N1002, N660, N856);
nand NAND2 (N1014, N1008, N523);
nand NAND2 (N1015, N998, N850);
and AND2 (N1016, N1009, N739);
or OR2 (N1017, N1013, N433);
nor NOR4 (N1018, N1006, N373, N1017, N254);
xor XOR2 (N1019, N891, N451);
or OR3 (N1020, N1011, N425, N747);
not NOT1 (N1021, N980);
and AND2 (N1022, N1014, N486);
nor NOR2 (N1023, N995, N764);
xor XOR2 (N1024, N1010, N564);
xor XOR2 (N1025, N1023, N188);
nand NAND3 (N1026, N1022, N584, N583);
and AND2 (N1027, N1026, N274);
and AND3 (N1028, N1019, N105, N287);
nor NOR3 (N1029, N1027, N909, N10);
buf BUF1 (N1030, N1024);
and AND3 (N1031, N1030, N168, N419);
xor XOR2 (N1032, N1015, N147);
not NOT1 (N1033, N1016);
not NOT1 (N1034, N1021);
and AND3 (N1035, N1031, N126, N758);
not NOT1 (N1036, N1033);
not NOT1 (N1037, N1034);
xor XOR2 (N1038, N1025, N487);
xor XOR2 (N1039, N1012, N683);
nand NAND3 (N1040, N1029, N748, N419);
and AND4 (N1041, N1040, N1022, N360, N226);
xor XOR2 (N1042, N1032, N604);
nor NOR4 (N1043, N1041, N432, N732, N1018);
nand NAND3 (N1044, N21, N792, N1031);
or OR3 (N1045, N1039, N128, N383);
buf BUF1 (N1046, N1028);
not NOT1 (N1047, N1020);
not NOT1 (N1048, N1037);
buf BUF1 (N1049, N1043);
xor XOR2 (N1050, N1048, N532);
xor XOR2 (N1051, N1050, N629);
xor XOR2 (N1052, N1036, N170);
buf BUF1 (N1053, N1042);
or OR3 (N1054, N1051, N487, N676);
nor NOR2 (N1055, N1035, N148);
xor XOR2 (N1056, N1047, N181);
buf BUF1 (N1057, N1055);
xor XOR2 (N1058, N1038, N701);
buf BUF1 (N1059, N1053);
and AND4 (N1060, N1058, N568, N1036, N899);
nand NAND3 (N1061, N1054, N588, N466);
xor XOR2 (N1062, N1057, N532);
buf BUF1 (N1063, N1056);
and AND2 (N1064, N1059, N968);
or OR4 (N1065, N1052, N103, N137, N67);
not NOT1 (N1066, N1065);
nor NOR2 (N1067, N1060, N209);
nand NAND3 (N1068, N1064, N200, N456);
not NOT1 (N1069, N1045);
nand NAND3 (N1070, N1063, N388, N993);
not NOT1 (N1071, N1046);
nor NOR3 (N1072, N1049, N825, N628);
or OR2 (N1073, N1071, N458);
buf BUF1 (N1074, N1067);
nor NOR4 (N1075, N1068, N456, N555, N527);
nor NOR2 (N1076, N1075, N408);
nand NAND2 (N1077, N1061, N184);
or OR2 (N1078, N1044, N435);
not NOT1 (N1079, N1070);
nand NAND2 (N1080, N1079, N71);
or OR2 (N1081, N1080, N969);
not NOT1 (N1082, N1077);
nor NOR3 (N1083, N1076, N976, N765);
nand NAND4 (N1084, N1081, N975, N29, N305);
nor NOR2 (N1085, N1078, N317);
and AND4 (N1086, N1083, N895, N440, N352);
or OR4 (N1087, N1072, N685, N1053, N273);
xor XOR2 (N1088, N1066, N615);
and AND2 (N1089, N1082, N15);
nor NOR2 (N1090, N1062, N167);
and AND3 (N1091, N1088, N829, N1006);
buf BUF1 (N1092, N1085);
not NOT1 (N1093, N1091);
nand NAND2 (N1094, N1087, N508);
xor XOR2 (N1095, N1086, N472);
nand NAND2 (N1096, N1069, N805);
and AND2 (N1097, N1092, N705);
nand NAND3 (N1098, N1096, N92, N749);
buf BUF1 (N1099, N1094);
nand NAND4 (N1100, N1084, N438, N22, N868);
nor NOR2 (N1101, N1097, N887);
xor XOR2 (N1102, N1089, N146);
nor NOR3 (N1103, N1090, N735, N601);
nand NAND2 (N1104, N1093, N707);
and AND2 (N1105, N1103, N770);
nand NAND3 (N1106, N1074, N540, N329);
buf BUF1 (N1107, N1098);
not NOT1 (N1108, N1106);
or OR2 (N1109, N1100, N231);
nand NAND2 (N1110, N1109, N901);
and AND2 (N1111, N1102, N644);
or OR4 (N1112, N1104, N99, N521, N528);
and AND4 (N1113, N1101, N542, N720, N216);
xor XOR2 (N1114, N1112, N101);
nor NOR3 (N1115, N1095, N1111, N1026);
and AND3 (N1116, N1068, N499, N351);
not NOT1 (N1117, N1114);
or OR3 (N1118, N1110, N924, N594);
buf BUF1 (N1119, N1107);
xor XOR2 (N1120, N1105, N115);
buf BUF1 (N1121, N1119);
not NOT1 (N1122, N1115);
nor NOR2 (N1123, N1099, N986);
nand NAND4 (N1124, N1113, N696, N888, N284);
xor XOR2 (N1125, N1123, N46);
xor XOR2 (N1126, N1124, N926);
and AND3 (N1127, N1073, N1015, N1008);
or OR2 (N1128, N1116, N482);
or OR4 (N1129, N1128, N665, N540, N229);
nand NAND3 (N1130, N1117, N1028, N92);
xor XOR2 (N1131, N1120, N61);
not NOT1 (N1132, N1131);
and AND2 (N1133, N1127, N178);
nand NAND4 (N1134, N1133, N644, N141, N834);
not NOT1 (N1135, N1126);
or OR2 (N1136, N1122, N1082);
not NOT1 (N1137, N1134);
nand NAND4 (N1138, N1121, N58, N238, N611);
and AND3 (N1139, N1138, N130, N1101);
and AND3 (N1140, N1132, N346, N51);
nand NAND2 (N1141, N1137, N821);
not NOT1 (N1142, N1139);
not NOT1 (N1143, N1118);
or OR4 (N1144, N1142, N270, N585, N27);
not NOT1 (N1145, N1135);
not NOT1 (N1146, N1108);
not NOT1 (N1147, N1125);
buf BUF1 (N1148, N1136);
not NOT1 (N1149, N1148);
and AND3 (N1150, N1149, N498, N143);
xor XOR2 (N1151, N1140, N842);
buf BUF1 (N1152, N1146);
nand NAND4 (N1153, N1147, N110, N834, N1145);
buf BUF1 (N1154, N942);
nand NAND2 (N1155, N1154, N523);
nor NOR4 (N1156, N1130, N665, N692, N263);
nand NAND4 (N1157, N1152, N1155, N1112, N1024);
nor NOR2 (N1158, N66, N978);
or OR4 (N1159, N1144, N413, N847, N1028);
nor NOR3 (N1160, N1153, N102, N865);
and AND3 (N1161, N1159, N542, N361);
nor NOR2 (N1162, N1156, N41);
not NOT1 (N1163, N1129);
buf BUF1 (N1164, N1162);
or OR4 (N1165, N1163, N576, N739, N918);
or OR2 (N1166, N1164, N1138);
buf BUF1 (N1167, N1165);
buf BUF1 (N1168, N1150);
xor XOR2 (N1169, N1143, N44);
nor NOR2 (N1170, N1151, N172);
and AND3 (N1171, N1157, N467, N177);
or OR2 (N1172, N1169, N576);
and AND3 (N1173, N1161, N667, N441);
not NOT1 (N1174, N1173);
or OR4 (N1175, N1172, N954, N217, N406);
nand NAND3 (N1176, N1167, N635, N829);
nor NOR2 (N1177, N1160, N1075);
nand NAND2 (N1178, N1171, N730);
and AND2 (N1179, N1177, N231);
nand NAND2 (N1180, N1175, N770);
nand NAND2 (N1181, N1178, N518);
nor NOR3 (N1182, N1168, N461, N207);
nand NAND3 (N1183, N1174, N842, N831);
xor XOR2 (N1184, N1180, N813);
and AND4 (N1185, N1158, N1150, N969, N539);
not NOT1 (N1186, N1184);
buf BUF1 (N1187, N1181);
nand NAND4 (N1188, N1183, N484, N1075, N1031);
not NOT1 (N1189, N1179);
and AND4 (N1190, N1176, N863, N787, N835);
nand NAND4 (N1191, N1189, N428, N386, N1145);
xor XOR2 (N1192, N1166, N722);
nor NOR2 (N1193, N1170, N317);
xor XOR2 (N1194, N1182, N611);
nor NOR2 (N1195, N1186, N281);
and AND3 (N1196, N1187, N977, N477);
nand NAND3 (N1197, N1141, N963, N853);
buf BUF1 (N1198, N1194);
nor NOR4 (N1199, N1198, N160, N281, N113);
nand NAND3 (N1200, N1191, N927, N704);
buf BUF1 (N1201, N1192);
nor NOR2 (N1202, N1196, N1043);
or OR2 (N1203, N1190, N659);
buf BUF1 (N1204, N1185);
buf BUF1 (N1205, N1193);
nor NOR4 (N1206, N1200, N704, N248, N812);
xor XOR2 (N1207, N1203, N898);
nand NAND3 (N1208, N1202, N271, N675);
buf BUF1 (N1209, N1207);
buf BUF1 (N1210, N1204);
nand NAND4 (N1211, N1188, N866, N1154, N1196);
nand NAND4 (N1212, N1209, N536, N1135, N1171);
nor NOR3 (N1213, N1208, N1029, N903);
nor NOR4 (N1214, N1206, N860, N837, N1011);
nor NOR2 (N1215, N1213, N274);
and AND2 (N1216, N1199, N686);
and AND3 (N1217, N1197, N1173, N250);
xor XOR2 (N1218, N1212, N609);
buf BUF1 (N1219, N1215);
buf BUF1 (N1220, N1195);
not NOT1 (N1221, N1217);
nor NOR3 (N1222, N1221, N1055, N1029);
nor NOR3 (N1223, N1216, N999, N235);
nor NOR3 (N1224, N1214, N1055, N745);
nand NAND4 (N1225, N1224, N945, N155, N865);
and AND4 (N1226, N1210, N1087, N1107, N923);
nor NOR3 (N1227, N1226, N915, N962);
xor XOR2 (N1228, N1218, N1118);
nor NOR2 (N1229, N1227, N1142);
xor XOR2 (N1230, N1225, N392);
buf BUF1 (N1231, N1230);
nor NOR2 (N1232, N1205, N866);
nor NOR3 (N1233, N1220, N174, N744);
not NOT1 (N1234, N1233);
nor NOR3 (N1235, N1222, N39, N697);
and AND2 (N1236, N1211, N680);
xor XOR2 (N1237, N1201, N197);
buf BUF1 (N1238, N1231);
or OR2 (N1239, N1219, N418);
nand NAND2 (N1240, N1229, N731);
nand NAND2 (N1241, N1237, N1152);
or OR3 (N1242, N1239, N948, N1158);
nor NOR2 (N1243, N1241, N432);
nand NAND3 (N1244, N1236, N788, N932);
nand NAND3 (N1245, N1223, N711, N960);
xor XOR2 (N1246, N1238, N968);
nand NAND2 (N1247, N1246, N48);
not NOT1 (N1248, N1234);
buf BUF1 (N1249, N1242);
not NOT1 (N1250, N1247);
buf BUF1 (N1251, N1250);
and AND4 (N1252, N1240, N902, N1223, N398);
xor XOR2 (N1253, N1248, N613);
not NOT1 (N1254, N1235);
and AND3 (N1255, N1252, N657, N1002);
nor NOR3 (N1256, N1251, N298, N422);
buf BUF1 (N1257, N1256);
xor XOR2 (N1258, N1244, N301);
nand NAND4 (N1259, N1257, N668, N839, N658);
and AND3 (N1260, N1228, N572, N1179);
nand NAND4 (N1261, N1258, N337, N415, N422);
and AND4 (N1262, N1259, N1213, N668, N991);
xor XOR2 (N1263, N1255, N443);
and AND4 (N1264, N1262, N481, N1020, N581);
xor XOR2 (N1265, N1243, N1200);
nor NOR2 (N1266, N1264, N42);
xor XOR2 (N1267, N1266, N469);
nand NAND3 (N1268, N1249, N1125, N514);
buf BUF1 (N1269, N1267);
and AND4 (N1270, N1232, N1251, N325, N829);
and AND3 (N1271, N1245, N1034, N552);
or OR4 (N1272, N1261, N651, N252, N74);
nor NOR2 (N1273, N1253, N50);
buf BUF1 (N1274, N1260);
or OR4 (N1275, N1269, N505, N1033, N421);
and AND2 (N1276, N1271, N1191);
xor XOR2 (N1277, N1270, N816);
not NOT1 (N1278, N1265);
and AND2 (N1279, N1273, N250);
buf BUF1 (N1280, N1254);
and AND4 (N1281, N1263, N951, N135, N228);
buf BUF1 (N1282, N1278);
or OR2 (N1283, N1277, N464);
xor XOR2 (N1284, N1281, N353);
and AND2 (N1285, N1275, N288);
or OR2 (N1286, N1279, N802);
buf BUF1 (N1287, N1274);
or OR2 (N1288, N1272, N683);
buf BUF1 (N1289, N1286);
buf BUF1 (N1290, N1284);
buf BUF1 (N1291, N1290);
xor XOR2 (N1292, N1282, N437);
buf BUF1 (N1293, N1276);
xor XOR2 (N1294, N1285, N512);
or OR3 (N1295, N1287, N919, N680);
or OR4 (N1296, N1293, N158, N151, N402);
or OR4 (N1297, N1268, N1265, N483, N963);
or OR2 (N1298, N1291, N1170);
nand NAND2 (N1299, N1295, N533);
not NOT1 (N1300, N1289);
or OR4 (N1301, N1299, N305, N33, N431);
xor XOR2 (N1302, N1280, N581);
and AND3 (N1303, N1288, N1246, N201);
or OR4 (N1304, N1298, N1133, N1184, N896);
nor NOR2 (N1305, N1283, N559);
xor XOR2 (N1306, N1300, N435);
or OR2 (N1307, N1294, N1038);
buf BUF1 (N1308, N1302);
and AND2 (N1309, N1303, N1286);
buf BUF1 (N1310, N1305);
xor XOR2 (N1311, N1309, N162);
xor XOR2 (N1312, N1308, N924);
not NOT1 (N1313, N1301);
not NOT1 (N1314, N1292);
buf BUF1 (N1315, N1313);
buf BUF1 (N1316, N1296);
nand NAND4 (N1317, N1311, N1071, N81, N500);
nand NAND2 (N1318, N1304, N1312);
xor XOR2 (N1319, N599, N371);
xor XOR2 (N1320, N1319, N388);
xor XOR2 (N1321, N1314, N33);
buf BUF1 (N1322, N1307);
xor XOR2 (N1323, N1310, N1229);
buf BUF1 (N1324, N1322);
or OR3 (N1325, N1317, N659, N1157);
nor NOR3 (N1326, N1316, N30, N747);
xor XOR2 (N1327, N1306, N970);
xor XOR2 (N1328, N1327, N1297);
buf BUF1 (N1329, N813);
not NOT1 (N1330, N1329);
nand NAND2 (N1331, N1320, N983);
or OR2 (N1332, N1315, N651);
nor NOR2 (N1333, N1318, N778);
or OR2 (N1334, N1328, N482);
and AND2 (N1335, N1331, N1209);
buf BUF1 (N1336, N1324);
not NOT1 (N1337, N1333);
and AND3 (N1338, N1330, N233, N374);
or OR4 (N1339, N1326, N669, N425, N1265);
or OR3 (N1340, N1338, N851, N587);
and AND4 (N1341, N1340, N311, N996, N419);
or OR4 (N1342, N1336, N1098, N625, N238);
not NOT1 (N1343, N1325);
and AND4 (N1344, N1342, N986, N1285, N384);
or OR4 (N1345, N1343, N551, N947, N325);
nand NAND3 (N1346, N1345, N611, N626);
xor XOR2 (N1347, N1335, N295);
buf BUF1 (N1348, N1334);
or OR2 (N1349, N1341, N1114);
and AND4 (N1350, N1339, N613, N250, N747);
buf BUF1 (N1351, N1321);
buf BUF1 (N1352, N1344);
xor XOR2 (N1353, N1323, N827);
xor XOR2 (N1354, N1353, N712);
and AND2 (N1355, N1349, N240);
nand NAND2 (N1356, N1332, N1348);
and AND4 (N1357, N314, N328, N24, N438);
buf BUF1 (N1358, N1347);
nand NAND3 (N1359, N1350, N70, N745);
or OR2 (N1360, N1352, N595);
nor NOR3 (N1361, N1356, N682, N1253);
not NOT1 (N1362, N1337);
or OR4 (N1363, N1346, N53, N809, N607);
nor NOR4 (N1364, N1357, N99, N1044, N1229);
buf BUF1 (N1365, N1362);
buf BUF1 (N1366, N1359);
nand NAND3 (N1367, N1366, N1353, N1254);
nand NAND2 (N1368, N1354, N206);
or OR4 (N1369, N1363, N1161, N1077, N658);
xor XOR2 (N1370, N1351, N1112);
xor XOR2 (N1371, N1358, N1298);
and AND3 (N1372, N1361, N623, N208);
nor NOR2 (N1373, N1369, N827);
nand NAND2 (N1374, N1365, N602);
xor XOR2 (N1375, N1372, N569);
nand NAND3 (N1376, N1364, N1365, N892);
nand NAND3 (N1377, N1367, N547, N723);
buf BUF1 (N1378, N1355);
nor NOR3 (N1379, N1370, N288, N140);
and AND4 (N1380, N1375, N453, N1265, N572);
and AND4 (N1381, N1371, N798, N1218, N536);
and AND3 (N1382, N1378, N745, N917);
buf BUF1 (N1383, N1373);
nand NAND3 (N1384, N1381, N165, N272);
nor NOR4 (N1385, N1382, N1368, N278, N979);
and AND4 (N1386, N945, N578, N1207, N100);
or OR2 (N1387, N1377, N116);
and AND3 (N1388, N1374, N1315, N25);
not NOT1 (N1389, N1379);
or OR4 (N1390, N1380, N792, N1188, N55);
xor XOR2 (N1391, N1376, N1093);
nor NOR4 (N1392, N1383, N1149, N194, N690);
nor NOR3 (N1393, N1390, N484, N137);
nand NAND3 (N1394, N1385, N882, N96);
nor NOR3 (N1395, N1386, N805, N660);
buf BUF1 (N1396, N1389);
nand NAND2 (N1397, N1395, N1017);
not NOT1 (N1398, N1387);
or OR2 (N1399, N1397, N1004);
nand NAND3 (N1400, N1392, N799, N1194);
buf BUF1 (N1401, N1360);
buf BUF1 (N1402, N1401);
buf BUF1 (N1403, N1398);
and AND4 (N1404, N1399, N1132, N1156, N574);
not NOT1 (N1405, N1388);
not NOT1 (N1406, N1402);
not NOT1 (N1407, N1384);
nand NAND3 (N1408, N1404, N671, N973);
not NOT1 (N1409, N1405);
buf BUF1 (N1410, N1403);
buf BUF1 (N1411, N1394);
buf BUF1 (N1412, N1406);
nor NOR2 (N1413, N1396, N1250);
buf BUF1 (N1414, N1410);
and AND4 (N1415, N1393, N1354, N604, N1374);
not NOT1 (N1416, N1391);
buf BUF1 (N1417, N1413);
or OR3 (N1418, N1417, N60, N1383);
not NOT1 (N1419, N1411);
xor XOR2 (N1420, N1418, N469);
nand NAND4 (N1421, N1400, N640, N152, N116);
buf BUF1 (N1422, N1416);
nor NOR2 (N1423, N1412, N563);
nand NAND3 (N1424, N1421, N1400, N915);
or OR2 (N1425, N1407, N649);
xor XOR2 (N1426, N1420, N534);
xor XOR2 (N1427, N1426, N25);
nand NAND4 (N1428, N1422, N1108, N330, N338);
xor XOR2 (N1429, N1419, N731);
or OR2 (N1430, N1415, N562);
buf BUF1 (N1431, N1428);
not NOT1 (N1432, N1424);
nand NAND3 (N1433, N1429, N1087, N657);
not NOT1 (N1434, N1427);
nand NAND4 (N1435, N1430, N914, N1372, N1382);
or OR3 (N1436, N1423, N841, N327);
xor XOR2 (N1437, N1434, N110);
nor NOR3 (N1438, N1425, N469, N235);
or OR2 (N1439, N1436, N260);
nand NAND4 (N1440, N1435, N184, N132, N1131);
nor NOR3 (N1441, N1437, N1061, N336);
not NOT1 (N1442, N1433);
nand NAND4 (N1443, N1441, N281, N1238, N437);
not NOT1 (N1444, N1409);
xor XOR2 (N1445, N1442, N419);
or OR2 (N1446, N1445, N46);
nand NAND3 (N1447, N1438, N687, N1129);
buf BUF1 (N1448, N1431);
nand NAND3 (N1449, N1448, N728, N998);
not NOT1 (N1450, N1440);
and AND2 (N1451, N1450, N881);
and AND4 (N1452, N1446, N1376, N706, N1345);
buf BUF1 (N1453, N1414);
buf BUF1 (N1454, N1408);
nor NOR3 (N1455, N1451, N542, N205);
not NOT1 (N1456, N1447);
not NOT1 (N1457, N1455);
nand NAND3 (N1458, N1454, N1236, N1003);
or OR2 (N1459, N1439, N727);
nor NOR3 (N1460, N1453, N609, N871);
buf BUF1 (N1461, N1460);
buf BUF1 (N1462, N1458);
or OR3 (N1463, N1461, N1153, N78);
or OR2 (N1464, N1457, N660);
or OR3 (N1465, N1432, N606, N501);
nor NOR2 (N1466, N1449, N592);
and AND3 (N1467, N1456, N903, N859);
xor XOR2 (N1468, N1467, N761);
and AND4 (N1469, N1444, N983, N490, N336);
nor NOR2 (N1470, N1443, N1295);
not NOT1 (N1471, N1464);
or OR4 (N1472, N1462, N1080, N706, N369);
not NOT1 (N1473, N1452);
and AND3 (N1474, N1463, N1197, N343);
buf BUF1 (N1475, N1471);
not NOT1 (N1476, N1459);
or OR3 (N1477, N1469, N1382, N275);
and AND3 (N1478, N1470, N554, N597);
or OR3 (N1479, N1476, N1005, N1136);
not NOT1 (N1480, N1477);
buf BUF1 (N1481, N1480);
nor NOR3 (N1482, N1472, N1462, N426);
not NOT1 (N1483, N1466);
nand NAND4 (N1484, N1474, N1206, N1384, N1097);
and AND4 (N1485, N1483, N400, N824, N1379);
nand NAND4 (N1486, N1484, N864, N760, N704);
xor XOR2 (N1487, N1465, N1133);
not NOT1 (N1488, N1482);
or OR3 (N1489, N1479, N896, N1217);
buf BUF1 (N1490, N1486);
buf BUF1 (N1491, N1475);
buf BUF1 (N1492, N1485);
and AND2 (N1493, N1473, N225);
not NOT1 (N1494, N1491);
buf BUF1 (N1495, N1488);
nor NOR4 (N1496, N1489, N833, N72, N1038);
nor NOR3 (N1497, N1478, N746, N1077);
nand NAND4 (N1498, N1487, N337, N947, N289);
nand NAND3 (N1499, N1495, N609, N1046);
not NOT1 (N1500, N1494);
not NOT1 (N1501, N1496);
and AND3 (N1502, N1490, N1232, N394);
and AND4 (N1503, N1481, N40, N824, N1337);
xor XOR2 (N1504, N1497, N1408);
buf BUF1 (N1505, N1499);
buf BUF1 (N1506, N1505);
nor NOR3 (N1507, N1506, N808, N464);
or OR3 (N1508, N1501, N1033, N816);
buf BUF1 (N1509, N1498);
nor NOR3 (N1510, N1500, N1500, N1045);
and AND4 (N1511, N1502, N1138, N768, N252);
buf BUF1 (N1512, N1511);
xor XOR2 (N1513, N1512, N1);
and AND2 (N1514, N1510, N604);
or OR4 (N1515, N1513, N119, N189, N462);
xor XOR2 (N1516, N1514, N1335);
endmodule