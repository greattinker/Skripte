// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21;

output N12805,N12819,N12815,N12809,N12810,N12820,N12814,N12816,N12811,N12821;

or OR2 (N22, N18, N15);
and AND4 (N23, N18, N16, N2, N7);
xor XOR2 (N24, N9, N14);
nand NAND4 (N25, N9, N21, N24, N17);
buf BUF1 (N26, N17);
buf BUF1 (N27, N18);
buf BUF1 (N28, N5);
or OR2 (N29, N19, N18);
and AND3 (N30, N11, N1, N29);
buf BUF1 (N31, N24);
nor NOR2 (N32, N22, N25);
xor XOR2 (N33, N9, N19);
xor XOR2 (N34, N18, N9);
and AND2 (N35, N15, N4);
xor XOR2 (N36, N26, N24);
not NOT1 (N37, N23);
not NOT1 (N38, N34);
nor NOR4 (N39, N33, N26, N8, N19);
or OR2 (N40, N28, N37);
nand NAND3 (N41, N25, N21, N40);
or OR3 (N42, N34, N38, N17);
or OR3 (N43, N7, N2, N11);
and AND4 (N44, N27, N41, N38, N39);
buf BUF1 (N45, N30);
buf BUF1 (N46, N3);
nand NAND3 (N47, N10, N3, N19);
nor NOR2 (N48, N32, N25);
xor XOR2 (N49, N43, N45);
buf BUF1 (N50, N5);
nand NAND3 (N51, N49, N45, N50);
xor XOR2 (N52, N10, N25);
and AND4 (N53, N47, N44, N20, N47);
nand NAND2 (N54, N36, N53);
buf BUF1 (N55, N6);
nor NOR4 (N56, N52, N22, N32, N16);
nor NOR2 (N57, N12, N14);
or OR4 (N58, N55, N41, N29, N25);
and AND4 (N59, N31, N4, N10, N44);
not NOT1 (N60, N56);
buf BUF1 (N61, N57);
not NOT1 (N62, N48);
or OR2 (N63, N58, N18);
not NOT1 (N64, N61);
buf BUF1 (N65, N35);
not NOT1 (N66, N42);
and AND4 (N67, N65, N37, N64, N53);
not NOT1 (N68, N4);
nor NOR2 (N69, N68, N3);
nand NAND2 (N70, N60, N67);
buf BUF1 (N71, N60);
xor XOR2 (N72, N46, N53);
buf BUF1 (N73, N63);
not NOT1 (N74, N62);
nor NOR2 (N75, N73, N52);
xor XOR2 (N76, N74, N21);
or OR2 (N77, N54, N12);
not NOT1 (N78, N51);
and AND2 (N79, N71, N71);
not NOT1 (N80, N78);
buf BUF1 (N81, N80);
nor NOR2 (N82, N66, N62);
nand NAND4 (N83, N77, N30, N27, N82);
or OR2 (N84, N63, N82);
or OR3 (N85, N79, N2, N11);
xor XOR2 (N86, N76, N53);
buf BUF1 (N87, N70);
or OR4 (N88, N84, N13, N20, N37);
or OR2 (N89, N81, N82);
not NOT1 (N90, N59);
xor XOR2 (N91, N72, N85);
xor XOR2 (N92, N30, N64);
not NOT1 (N93, N69);
nand NAND2 (N94, N89, N20);
nand NAND3 (N95, N93, N9, N50);
nor NOR2 (N96, N94, N21);
or OR3 (N97, N86, N3, N70);
not NOT1 (N98, N92);
xor XOR2 (N99, N88, N46);
xor XOR2 (N100, N91, N80);
not NOT1 (N101, N90);
not NOT1 (N102, N101);
nor NOR2 (N103, N75, N65);
buf BUF1 (N104, N83);
xor XOR2 (N105, N96, N79);
xor XOR2 (N106, N98, N101);
or OR3 (N107, N105, N92, N23);
not NOT1 (N108, N107);
buf BUF1 (N109, N99);
xor XOR2 (N110, N104, N52);
nor NOR2 (N111, N108, N79);
not NOT1 (N112, N97);
xor XOR2 (N113, N112, N83);
nor NOR4 (N114, N100, N11, N90, N110);
nand NAND3 (N115, N109, N81, N14);
xor XOR2 (N116, N61, N94);
buf BUF1 (N117, N114);
not NOT1 (N118, N106);
not NOT1 (N119, N87);
nor NOR4 (N120, N116, N43, N97, N42);
or OR4 (N121, N111, N55, N111, N20);
or OR4 (N122, N95, N89, N83, N40);
nand NAND2 (N123, N102, N69);
xor XOR2 (N124, N113, N116);
not NOT1 (N125, N117);
and AND2 (N126, N115, N29);
and AND4 (N127, N119, N18, N23, N74);
or OR2 (N128, N123, N35);
xor XOR2 (N129, N120, N9);
nand NAND2 (N130, N124, N49);
nand NAND4 (N131, N125, N23, N56, N108);
nor NOR4 (N132, N126, N12, N6, N86);
nand NAND4 (N133, N132, N104, N92, N61);
and AND3 (N134, N121, N38, N64);
xor XOR2 (N135, N131, N81);
nand NAND4 (N136, N134, N79, N5, N18);
xor XOR2 (N137, N133, N113);
not NOT1 (N138, N135);
or OR4 (N139, N136, N123, N81, N77);
not NOT1 (N140, N122);
nand NAND3 (N141, N139, N117, N20);
not NOT1 (N142, N127);
nand NAND4 (N143, N141, N19, N111, N126);
nand NAND2 (N144, N103, N53);
and AND4 (N145, N144, N117, N101, N54);
xor XOR2 (N146, N130, N53);
not NOT1 (N147, N129);
nand NAND4 (N148, N140, N18, N71, N129);
not NOT1 (N149, N137);
buf BUF1 (N150, N146);
buf BUF1 (N151, N143);
not NOT1 (N152, N151);
nor NOR3 (N153, N118, N106, N114);
xor XOR2 (N154, N148, N109);
and AND2 (N155, N138, N36);
not NOT1 (N156, N150);
buf BUF1 (N157, N154);
and AND4 (N158, N128, N132, N50, N107);
and AND3 (N159, N149, N125, N22);
xor XOR2 (N160, N142, N56);
or OR4 (N161, N157, N77, N79, N29);
buf BUF1 (N162, N153);
buf BUF1 (N163, N161);
and AND4 (N164, N160, N16, N37, N4);
or OR4 (N165, N156, N44, N157, N13);
not NOT1 (N166, N145);
not NOT1 (N167, N159);
nand NAND3 (N168, N158, N102, N54);
nand NAND2 (N169, N152, N108);
nor NOR2 (N170, N162, N136);
xor XOR2 (N171, N165, N28);
xor XOR2 (N172, N168, N6);
nor NOR2 (N173, N172, N132);
nor NOR4 (N174, N167, N128, N33, N97);
or OR3 (N175, N171, N51, N80);
and AND3 (N176, N164, N159, N81);
nor NOR2 (N177, N173, N14);
and AND4 (N178, N174, N172, N22, N66);
not NOT1 (N179, N155);
nor NOR4 (N180, N178, N7, N29, N136);
xor XOR2 (N181, N166, N45);
nand NAND4 (N182, N147, N177, N55, N181);
nand NAND2 (N183, N154, N136);
and AND3 (N184, N138, N105, N146);
nor NOR4 (N185, N175, N108, N78, N177);
or OR4 (N186, N185, N97, N25, N33);
xor XOR2 (N187, N169, N37);
buf BUF1 (N188, N170);
not NOT1 (N189, N179);
or OR4 (N190, N188, N74, N119, N68);
xor XOR2 (N191, N182, N186);
xor XOR2 (N192, N27, N104);
xor XOR2 (N193, N189, N143);
and AND3 (N194, N193, N174, N174);
buf BUF1 (N195, N194);
not NOT1 (N196, N184);
xor XOR2 (N197, N196, N77);
buf BUF1 (N198, N163);
nor NOR4 (N199, N197, N109, N194, N93);
buf BUF1 (N200, N195);
not NOT1 (N201, N191);
nand NAND4 (N202, N183, N185, N118, N27);
xor XOR2 (N203, N187, N166);
and AND3 (N204, N198, N79, N22);
nand NAND3 (N205, N201, N185, N148);
not NOT1 (N206, N199);
xor XOR2 (N207, N205, N49);
nor NOR3 (N208, N206, N198, N201);
buf BUF1 (N209, N207);
not NOT1 (N210, N208);
buf BUF1 (N211, N180);
not NOT1 (N212, N190);
buf BUF1 (N213, N209);
nand NAND3 (N214, N200, N24, N99);
xor XOR2 (N215, N212, N29);
or OR4 (N216, N203, N50, N61, N59);
or OR2 (N217, N215, N11);
and AND4 (N218, N192, N170, N135, N155);
and AND4 (N219, N216, N28, N122, N126);
and AND4 (N220, N218, N44, N138, N182);
nand NAND2 (N221, N211, N63);
or OR3 (N222, N176, N14, N164);
and AND3 (N223, N210, N20, N71);
or OR2 (N224, N202, N128);
not NOT1 (N225, N213);
or OR4 (N226, N219, N7, N71, N206);
buf BUF1 (N227, N222);
nor NOR4 (N228, N224, N9, N177, N219);
nor NOR4 (N229, N214, N209, N92, N208);
nor NOR3 (N230, N227, N158, N182);
buf BUF1 (N231, N223);
nor NOR2 (N232, N230, N223);
not NOT1 (N233, N204);
buf BUF1 (N234, N233);
xor XOR2 (N235, N234, N45);
or OR3 (N236, N232, N180, N137);
nand NAND3 (N237, N221, N70, N23);
buf BUF1 (N238, N236);
and AND2 (N239, N238, N10);
buf BUF1 (N240, N235);
buf BUF1 (N241, N228);
xor XOR2 (N242, N231, N136);
or OR4 (N243, N217, N48, N210, N212);
or OR2 (N244, N225, N92);
nor NOR2 (N245, N241, N196);
and AND3 (N246, N243, N53, N70);
buf BUF1 (N247, N220);
and AND4 (N248, N247, N203, N203, N160);
nor NOR3 (N249, N242, N184, N216);
or OR3 (N250, N249, N217, N101);
buf BUF1 (N251, N240);
nand NAND4 (N252, N226, N78, N40, N196);
nor NOR3 (N253, N237, N211, N228);
buf BUF1 (N254, N253);
xor XOR2 (N255, N248, N249);
and AND4 (N256, N252, N209, N117, N239);
and AND3 (N257, N119, N20, N127);
nand NAND2 (N258, N254, N113);
buf BUF1 (N259, N246);
xor XOR2 (N260, N251, N50);
and AND3 (N261, N245, N50, N139);
buf BUF1 (N262, N244);
not NOT1 (N263, N262);
buf BUF1 (N264, N258);
nor NOR4 (N265, N257, N72, N71, N174);
not NOT1 (N266, N256);
buf BUF1 (N267, N266);
not NOT1 (N268, N267);
or OR4 (N269, N229, N193, N1, N154);
not NOT1 (N270, N260);
not NOT1 (N271, N270);
xor XOR2 (N272, N263, N191);
not NOT1 (N273, N261);
buf BUF1 (N274, N268);
or OR3 (N275, N250, N20, N47);
and AND3 (N276, N264, N86, N22);
nand NAND2 (N277, N275, N94);
and AND3 (N278, N273, N148, N231);
nand NAND3 (N279, N271, N195, N216);
or OR2 (N280, N278, N131);
nand NAND2 (N281, N259, N18);
and AND4 (N282, N276, N177, N248, N267);
nand NAND4 (N283, N255, N19, N154, N124);
nand NAND4 (N284, N279, N253, N4, N203);
not NOT1 (N285, N272);
nand NAND3 (N286, N280, N275, N249);
nor NOR4 (N287, N274, N14, N31, N204);
nor NOR3 (N288, N265, N242, N206);
not NOT1 (N289, N269);
or OR2 (N290, N281, N140);
and AND2 (N291, N283, N152);
or OR3 (N292, N288, N274, N270);
not NOT1 (N293, N289);
nor NOR4 (N294, N287, N250, N219, N170);
not NOT1 (N295, N292);
and AND4 (N296, N284, N60, N287, N49);
not NOT1 (N297, N285);
or OR3 (N298, N290, N201, N230);
or OR4 (N299, N294, N175, N56, N104);
xor XOR2 (N300, N286, N152);
or OR2 (N301, N295, N138);
nor NOR3 (N302, N299, N169, N197);
buf BUF1 (N303, N297);
and AND2 (N304, N302, N52);
not NOT1 (N305, N301);
nand NAND4 (N306, N298, N229, N165, N290);
buf BUF1 (N307, N296);
nand NAND3 (N308, N305, N226, N130);
or OR3 (N309, N293, N117, N124);
nand NAND4 (N310, N277, N66, N80, N117);
buf BUF1 (N311, N308);
not NOT1 (N312, N307);
and AND3 (N313, N309, N229, N16);
not NOT1 (N314, N311);
not NOT1 (N315, N312);
and AND4 (N316, N313, N291, N261, N180);
and AND4 (N317, N70, N279, N304, N164);
xor XOR2 (N318, N23, N12);
not NOT1 (N319, N318);
nor NOR4 (N320, N303, N136, N162, N33);
nand NAND2 (N321, N314, N223);
nor NOR3 (N322, N315, N14, N277);
nor NOR4 (N323, N322, N177, N100, N69);
not NOT1 (N324, N319);
not NOT1 (N325, N306);
and AND4 (N326, N321, N32, N199, N161);
xor XOR2 (N327, N317, N174);
not NOT1 (N328, N325);
not NOT1 (N329, N328);
and AND2 (N330, N310, N124);
buf BUF1 (N331, N300);
and AND2 (N332, N323, N192);
and AND4 (N333, N326, N232, N146, N246);
buf BUF1 (N334, N320);
not NOT1 (N335, N334);
or OR4 (N336, N316, N208, N326, N120);
not NOT1 (N337, N335);
xor XOR2 (N338, N324, N135);
xor XOR2 (N339, N338, N228);
and AND3 (N340, N337, N284, N43);
nor NOR2 (N341, N329, N77);
nor NOR3 (N342, N331, N108, N179);
or OR2 (N343, N342, N51);
buf BUF1 (N344, N343);
nand NAND3 (N345, N282, N196, N237);
or OR3 (N346, N333, N135, N126);
or OR3 (N347, N341, N75, N12);
xor XOR2 (N348, N327, N255);
and AND4 (N349, N340, N169, N136, N148);
not NOT1 (N350, N349);
nor NOR2 (N351, N350, N113);
or OR3 (N352, N339, N90, N305);
and AND2 (N353, N348, N180);
nor NOR3 (N354, N336, N306, N149);
not NOT1 (N355, N354);
or OR4 (N356, N330, N307, N7, N32);
buf BUF1 (N357, N355);
xor XOR2 (N358, N356, N90);
not NOT1 (N359, N346);
nor NOR3 (N360, N353, N106, N329);
nor NOR4 (N361, N357, N115, N322, N143);
buf BUF1 (N362, N345);
nor NOR2 (N363, N361, N212);
buf BUF1 (N364, N358);
not NOT1 (N365, N360);
nor NOR4 (N366, N352, N336, N187, N164);
xor XOR2 (N367, N332, N153);
or OR2 (N368, N365, N262);
and AND4 (N369, N363, N78, N58, N350);
or OR3 (N370, N366, N320, N163);
xor XOR2 (N371, N368, N226);
and AND3 (N372, N351, N225, N193);
not NOT1 (N373, N359);
or OR2 (N374, N373, N154);
nor NOR4 (N375, N367, N305, N167, N297);
or OR4 (N376, N370, N282, N292, N216);
not NOT1 (N377, N375);
xor XOR2 (N378, N347, N314);
or OR4 (N379, N371, N165, N352, N120);
nand NAND4 (N380, N369, N254, N132, N67);
xor XOR2 (N381, N378, N162);
not NOT1 (N382, N379);
xor XOR2 (N383, N380, N72);
and AND4 (N384, N377, N234, N365, N177);
xor XOR2 (N385, N383, N29);
xor XOR2 (N386, N382, N360);
buf BUF1 (N387, N344);
xor XOR2 (N388, N384, N62);
and AND4 (N389, N374, N153, N344, N141);
and AND2 (N390, N385, N85);
nand NAND2 (N391, N386, N146);
not NOT1 (N392, N387);
xor XOR2 (N393, N388, N251);
nand NAND4 (N394, N364, N239, N85, N242);
nor NOR2 (N395, N376, N301);
or OR4 (N396, N391, N297, N39, N293);
and AND3 (N397, N362, N248, N328);
nor NOR2 (N398, N397, N289);
nor NOR3 (N399, N390, N209, N296);
xor XOR2 (N400, N398, N210);
nor NOR2 (N401, N392, N16);
and AND4 (N402, N394, N291, N138, N84);
nor NOR3 (N403, N401, N346, N127);
and AND2 (N404, N372, N344);
nand NAND2 (N405, N402, N61);
buf BUF1 (N406, N404);
and AND4 (N407, N406, N284, N86, N327);
xor XOR2 (N408, N400, N285);
nand NAND2 (N409, N389, N108);
and AND2 (N410, N399, N323);
not NOT1 (N411, N408);
or OR3 (N412, N409, N326, N301);
nand NAND3 (N413, N412, N22, N295);
or OR2 (N414, N393, N26);
buf BUF1 (N415, N396);
buf BUF1 (N416, N381);
nand NAND3 (N417, N414, N31, N38);
buf BUF1 (N418, N405);
buf BUF1 (N419, N415);
nor NOR3 (N420, N419, N362, N56);
xor XOR2 (N421, N407, N361);
not NOT1 (N422, N410);
nand NAND3 (N423, N411, N408, N410);
nand NAND4 (N424, N416, N124, N362, N393);
xor XOR2 (N425, N403, N403);
xor XOR2 (N426, N395, N246);
not NOT1 (N427, N423);
buf BUF1 (N428, N422);
nor NOR2 (N429, N428, N311);
nand NAND4 (N430, N413, N85, N48, N428);
nor NOR3 (N431, N418, N334, N422);
buf BUF1 (N432, N426);
and AND3 (N433, N424, N326, N296);
xor XOR2 (N434, N431, N319);
and AND2 (N435, N429, N430);
and AND3 (N436, N192, N88, N19);
nand NAND2 (N437, N420, N218);
or OR2 (N438, N435, N107);
nor NOR3 (N439, N436, N116, N356);
xor XOR2 (N440, N432, N243);
xor XOR2 (N441, N433, N99);
buf BUF1 (N442, N439);
and AND3 (N443, N421, N347, N361);
not NOT1 (N444, N442);
xor XOR2 (N445, N443, N45);
and AND2 (N446, N440, N77);
and AND4 (N447, N446, N42, N139, N374);
nand NAND4 (N448, N444, N162, N162, N302);
buf BUF1 (N449, N417);
nor NOR4 (N450, N437, N313, N4, N136);
buf BUF1 (N451, N445);
or OR3 (N452, N448, N271, N209);
nand NAND4 (N453, N449, N398, N86, N419);
or OR2 (N454, N450, N88);
nor NOR4 (N455, N425, N147, N121, N73);
nand NAND3 (N456, N452, N450, N302);
nand NAND2 (N457, N427, N41);
or OR3 (N458, N434, N173, N69);
not NOT1 (N459, N454);
nand NAND4 (N460, N457, N152, N175, N205);
nor NOR3 (N461, N453, N394, N93);
buf BUF1 (N462, N441);
and AND3 (N463, N458, N89, N398);
buf BUF1 (N464, N455);
not NOT1 (N465, N463);
nand NAND3 (N466, N447, N72, N78);
and AND4 (N467, N462, N187, N385, N233);
buf BUF1 (N468, N456);
or OR3 (N469, N466, N394, N41);
or OR3 (N470, N451, N372, N171);
nand NAND4 (N471, N464, N252, N48, N344);
nand NAND3 (N472, N465, N441, N10);
not NOT1 (N473, N461);
not NOT1 (N474, N470);
xor XOR2 (N475, N471, N446);
buf BUF1 (N476, N474);
buf BUF1 (N477, N438);
xor XOR2 (N478, N469, N23);
xor XOR2 (N479, N472, N459);
xor XOR2 (N480, N281, N275);
buf BUF1 (N481, N476);
buf BUF1 (N482, N467);
nor NOR2 (N483, N482, N210);
or OR4 (N484, N479, N427, N181, N328);
not NOT1 (N485, N483);
nand NAND2 (N486, N484, N449);
buf BUF1 (N487, N477);
or OR3 (N488, N475, N246, N326);
and AND2 (N489, N485, N158);
xor XOR2 (N490, N473, N68);
or OR2 (N491, N488, N460);
xor XOR2 (N492, N181, N148);
not NOT1 (N493, N490);
not NOT1 (N494, N492);
nor NOR4 (N495, N494, N17, N447, N51);
nor NOR3 (N496, N491, N384, N401);
nand NAND3 (N497, N480, N121, N71);
not NOT1 (N498, N495);
or OR2 (N499, N481, N428);
not NOT1 (N500, N497);
or OR3 (N501, N493, N22, N81);
not NOT1 (N502, N486);
not NOT1 (N503, N502);
buf BUF1 (N504, N498);
nand NAND3 (N505, N489, N222, N207);
nor NOR2 (N506, N468, N448);
or OR3 (N507, N503, N234, N337);
nor NOR4 (N508, N507, N178, N74, N440);
not NOT1 (N509, N487);
or OR4 (N510, N508, N443, N274, N306);
not NOT1 (N511, N478);
buf BUF1 (N512, N505);
not NOT1 (N513, N500);
nand NAND4 (N514, N499, N203, N240, N60);
and AND3 (N515, N511, N357, N315);
nor NOR3 (N516, N504, N149, N125);
not NOT1 (N517, N516);
nand NAND3 (N518, N512, N481, N172);
buf BUF1 (N519, N518);
nor NOR2 (N520, N515, N161);
not NOT1 (N521, N517);
or OR2 (N522, N521, N348);
or OR2 (N523, N519, N208);
buf BUF1 (N524, N509);
and AND2 (N525, N510, N40);
nand NAND2 (N526, N501, N227);
nor NOR3 (N527, N514, N56, N246);
xor XOR2 (N528, N496, N191);
and AND3 (N529, N506, N61, N244);
nor NOR3 (N530, N513, N207, N123);
xor XOR2 (N531, N520, N410);
and AND2 (N532, N523, N53);
or OR3 (N533, N532, N344, N227);
nor NOR3 (N534, N531, N58, N40);
and AND2 (N535, N528, N301);
nand NAND3 (N536, N527, N329, N430);
buf BUF1 (N537, N524);
nand NAND2 (N538, N526, N191);
xor XOR2 (N539, N533, N282);
xor XOR2 (N540, N529, N93);
not NOT1 (N541, N525);
buf BUF1 (N542, N534);
not NOT1 (N543, N538);
and AND4 (N544, N535, N64, N280, N253);
nand NAND3 (N545, N542, N460, N245);
or OR4 (N546, N545, N108, N247, N241);
nand NAND2 (N547, N543, N227);
nor NOR4 (N548, N539, N354, N409, N56);
or OR4 (N549, N547, N156, N120, N85);
not NOT1 (N550, N544);
nor NOR4 (N551, N530, N308, N40, N26);
nand NAND2 (N552, N549, N320);
xor XOR2 (N553, N540, N411);
xor XOR2 (N554, N537, N434);
xor XOR2 (N555, N553, N163);
buf BUF1 (N556, N546);
nand NAND4 (N557, N548, N185, N391, N149);
xor XOR2 (N558, N554, N446);
and AND2 (N559, N551, N157);
or OR3 (N560, N558, N534, N113);
xor XOR2 (N561, N550, N128);
xor XOR2 (N562, N552, N261);
xor XOR2 (N563, N559, N539);
not NOT1 (N564, N555);
and AND4 (N565, N563, N313, N70, N356);
xor XOR2 (N566, N560, N420);
nand NAND3 (N567, N541, N381, N169);
xor XOR2 (N568, N557, N529);
buf BUF1 (N569, N556);
buf BUF1 (N570, N561);
not NOT1 (N571, N568);
xor XOR2 (N572, N566, N504);
and AND2 (N573, N571, N140);
xor XOR2 (N574, N573, N7);
or OR4 (N575, N574, N356, N509, N186);
or OR3 (N576, N565, N561, N385);
and AND3 (N577, N564, N507, N420);
or OR2 (N578, N575, N536);
and AND4 (N579, N210, N7, N498, N244);
buf BUF1 (N580, N578);
nand NAND2 (N581, N576, N362);
xor XOR2 (N582, N577, N339);
buf BUF1 (N583, N569);
not NOT1 (N584, N522);
xor XOR2 (N585, N583, N536);
buf BUF1 (N586, N580);
nor NOR3 (N587, N562, N131, N473);
and AND3 (N588, N572, N293, N383);
buf BUF1 (N589, N581);
nand NAND2 (N590, N582, N463);
buf BUF1 (N591, N584);
xor XOR2 (N592, N587, N162);
buf BUF1 (N593, N586);
buf BUF1 (N594, N589);
xor XOR2 (N595, N591, N462);
nor NOR2 (N596, N595, N570);
and AND2 (N597, N316, N340);
nand NAND4 (N598, N567, N31, N494, N500);
not NOT1 (N599, N579);
not NOT1 (N600, N599);
not NOT1 (N601, N592);
nor NOR4 (N602, N598, N387, N160, N106);
xor XOR2 (N603, N593, N3);
and AND4 (N604, N600, N181, N527, N211);
nand NAND4 (N605, N588, N196, N78, N223);
and AND2 (N606, N604, N521);
or OR3 (N607, N602, N521, N210);
nor NOR4 (N608, N594, N499, N280, N109);
nor NOR3 (N609, N590, N4, N190);
and AND2 (N610, N601, N602);
or OR3 (N611, N585, N368, N545);
not NOT1 (N612, N605);
nor NOR2 (N613, N608, N71);
nor NOR3 (N614, N606, N185, N251);
nor NOR3 (N615, N612, N512, N314);
nor NOR4 (N616, N614, N555, N117, N473);
nand NAND4 (N617, N610, N465, N359, N180);
and AND3 (N618, N616, N538, N374);
or OR3 (N619, N596, N440, N310);
nand NAND3 (N620, N597, N449, N486);
and AND3 (N621, N613, N122, N208);
or OR2 (N622, N603, N319);
not NOT1 (N623, N619);
buf BUF1 (N624, N609);
not NOT1 (N625, N617);
not NOT1 (N626, N618);
and AND4 (N627, N626, N252, N147, N113);
xor XOR2 (N628, N623, N79);
nor NOR2 (N629, N622, N139);
or OR4 (N630, N615, N562, N312, N413);
nor NOR2 (N631, N607, N525);
nand NAND3 (N632, N621, N59, N379);
and AND2 (N633, N625, N262);
or OR3 (N634, N630, N414, N419);
or OR2 (N635, N628, N35);
xor XOR2 (N636, N635, N323);
xor XOR2 (N637, N629, N342);
and AND3 (N638, N637, N336, N303);
or OR3 (N639, N636, N1, N231);
nor NOR4 (N640, N632, N199, N5, N258);
not NOT1 (N641, N638);
buf BUF1 (N642, N620);
or OR4 (N643, N639, N272, N534, N1);
buf BUF1 (N644, N641);
xor XOR2 (N645, N633, N546);
buf BUF1 (N646, N611);
or OR3 (N647, N644, N344, N172);
nor NOR2 (N648, N646, N531);
not NOT1 (N649, N640);
nand NAND3 (N650, N627, N440, N291);
buf BUF1 (N651, N645);
and AND4 (N652, N642, N260, N373, N106);
nand NAND2 (N653, N648, N443);
not NOT1 (N654, N624);
or OR2 (N655, N634, N488);
nand NAND2 (N656, N653, N188);
not NOT1 (N657, N654);
or OR2 (N658, N650, N530);
and AND4 (N659, N652, N562, N186, N200);
nor NOR2 (N660, N631, N624);
or OR4 (N661, N655, N140, N329, N294);
and AND2 (N662, N658, N591);
nand NAND2 (N663, N643, N294);
and AND4 (N664, N659, N364, N576, N125);
buf BUF1 (N665, N657);
not NOT1 (N666, N661);
nor NOR4 (N667, N663, N502, N216, N221);
and AND2 (N668, N649, N278);
xor XOR2 (N669, N656, N129);
not NOT1 (N670, N660);
not NOT1 (N671, N670);
not NOT1 (N672, N668);
and AND3 (N673, N651, N257, N187);
and AND4 (N674, N672, N452, N608, N150);
buf BUF1 (N675, N665);
nor NOR4 (N676, N675, N6, N107, N504);
and AND3 (N677, N669, N286, N387);
nand NAND4 (N678, N666, N621, N475, N422);
or OR2 (N679, N664, N447);
not NOT1 (N680, N678);
not NOT1 (N681, N647);
buf BUF1 (N682, N676);
nor NOR3 (N683, N673, N374, N617);
not NOT1 (N684, N680);
xor XOR2 (N685, N683, N569);
nand NAND3 (N686, N679, N320, N598);
not NOT1 (N687, N686);
nor NOR2 (N688, N667, N15);
not NOT1 (N689, N684);
nand NAND2 (N690, N689, N460);
nand NAND2 (N691, N688, N305);
or OR3 (N692, N687, N401, N528);
nor NOR3 (N693, N662, N411, N213);
or OR4 (N694, N693, N611, N315, N262);
not NOT1 (N695, N694);
not NOT1 (N696, N671);
nand NAND3 (N697, N681, N172, N235);
nand NAND3 (N698, N677, N647, N238);
nor NOR4 (N699, N695, N267, N271, N423);
nor NOR3 (N700, N685, N653, N206);
nor NOR2 (N701, N690, N329);
and AND2 (N702, N692, N523);
and AND2 (N703, N699, N143);
nor NOR3 (N704, N702, N7, N255);
or OR4 (N705, N703, N545, N271, N104);
nor NOR4 (N706, N698, N624, N638, N524);
nand NAND3 (N707, N704, N533, N212);
buf BUF1 (N708, N682);
nand NAND3 (N709, N705, N237, N351);
and AND3 (N710, N697, N441, N312);
nand NAND4 (N711, N701, N381, N537, N277);
buf BUF1 (N712, N674);
not NOT1 (N713, N700);
and AND4 (N714, N696, N200, N3, N620);
not NOT1 (N715, N710);
and AND2 (N716, N715, N148);
and AND4 (N717, N713, N5, N54, N349);
not NOT1 (N718, N691);
nand NAND4 (N719, N718, N716, N635, N162);
buf BUF1 (N720, N104);
nand NAND3 (N721, N709, N629, N499);
xor XOR2 (N722, N720, N287);
xor XOR2 (N723, N722, N668);
nor NOR4 (N724, N706, N410, N22, N409);
nor NOR3 (N725, N717, N664, N622);
nor NOR3 (N726, N721, N627, N236);
nor NOR2 (N727, N723, N25);
nor NOR3 (N728, N711, N171, N408);
buf BUF1 (N729, N726);
nand NAND2 (N730, N712, N648);
buf BUF1 (N731, N719);
and AND3 (N732, N730, N457, N100);
and AND3 (N733, N724, N149, N74);
buf BUF1 (N734, N727);
not NOT1 (N735, N707);
and AND4 (N736, N714, N732, N495, N591);
nor NOR3 (N737, N131, N104, N549);
nand NAND4 (N738, N731, N639, N584, N419);
xor XOR2 (N739, N725, N190);
buf BUF1 (N740, N728);
nand NAND3 (N741, N737, N722, N640);
xor XOR2 (N742, N735, N312);
not NOT1 (N743, N739);
nor NOR4 (N744, N729, N13, N222, N161);
nor NOR2 (N745, N733, N548);
buf BUF1 (N746, N738);
nor NOR3 (N747, N742, N335, N262);
buf BUF1 (N748, N744);
and AND4 (N749, N745, N592, N20, N379);
buf BUF1 (N750, N734);
nor NOR3 (N751, N747, N176, N448);
buf BUF1 (N752, N741);
not NOT1 (N753, N743);
nand NAND4 (N754, N740, N684, N166, N243);
or OR4 (N755, N708, N474, N581, N699);
nand NAND2 (N756, N755, N491);
nor NOR2 (N757, N756, N357);
nor NOR2 (N758, N754, N507);
nor NOR3 (N759, N757, N590, N623);
xor XOR2 (N760, N752, N750);
and AND3 (N761, N91, N57, N257);
buf BUF1 (N762, N759);
buf BUF1 (N763, N753);
buf BUF1 (N764, N758);
not NOT1 (N765, N762);
xor XOR2 (N766, N749, N459);
nand NAND2 (N767, N766, N688);
not NOT1 (N768, N761);
xor XOR2 (N769, N760, N230);
xor XOR2 (N770, N763, N67);
not NOT1 (N771, N767);
buf BUF1 (N772, N770);
and AND2 (N773, N764, N711);
nor NOR2 (N774, N751, N511);
not NOT1 (N775, N773);
or OR4 (N776, N774, N33, N717, N549);
buf BUF1 (N777, N771);
xor XOR2 (N778, N748, N377);
buf BUF1 (N779, N772);
nor NOR2 (N780, N776, N741);
not NOT1 (N781, N780);
xor XOR2 (N782, N775, N279);
xor XOR2 (N783, N765, N375);
nor NOR3 (N784, N777, N38, N699);
not NOT1 (N785, N769);
nor NOR2 (N786, N768, N322);
or OR4 (N787, N778, N566, N301, N135);
buf BUF1 (N788, N746);
buf BUF1 (N789, N786);
nand NAND2 (N790, N788, N210);
nor NOR2 (N791, N736, N737);
nor NOR4 (N792, N790, N468, N623, N19);
nor NOR4 (N793, N781, N743, N742, N59);
not NOT1 (N794, N779);
or OR3 (N795, N784, N349, N718);
or OR2 (N796, N791, N794);
and AND3 (N797, N616, N404, N198);
nand NAND2 (N798, N787, N644);
not NOT1 (N799, N795);
nand NAND3 (N800, N782, N62, N775);
nand NAND2 (N801, N797, N537);
xor XOR2 (N802, N792, N588);
buf BUF1 (N803, N796);
and AND2 (N804, N789, N36);
buf BUF1 (N805, N799);
xor XOR2 (N806, N798, N490);
nor NOR3 (N807, N801, N265, N408);
and AND3 (N808, N785, N464, N516);
xor XOR2 (N809, N808, N371);
buf BUF1 (N810, N793);
xor XOR2 (N811, N803, N782);
nor NOR4 (N812, N800, N362, N793, N108);
and AND4 (N813, N809, N444, N737, N186);
buf BUF1 (N814, N805);
or OR3 (N815, N810, N673, N105);
nand NAND4 (N816, N802, N753, N75, N589);
xor XOR2 (N817, N813, N638);
nand NAND4 (N818, N807, N523, N337, N65);
and AND4 (N819, N783, N317, N510, N139);
not NOT1 (N820, N811);
nor NOR2 (N821, N818, N718);
nor NOR2 (N822, N815, N418);
or OR3 (N823, N817, N803, N447);
not NOT1 (N824, N816);
nand NAND4 (N825, N820, N355, N126, N659);
and AND2 (N826, N824, N481);
buf BUF1 (N827, N804);
nor NOR2 (N828, N826, N490);
and AND3 (N829, N825, N258, N293);
buf BUF1 (N830, N822);
buf BUF1 (N831, N821);
and AND2 (N832, N819, N568);
or OR2 (N833, N828, N510);
and AND4 (N834, N814, N650, N625, N53);
not NOT1 (N835, N830);
or OR3 (N836, N812, N75, N51);
and AND3 (N837, N829, N502, N202);
not NOT1 (N838, N823);
or OR4 (N839, N838, N709, N419, N541);
and AND2 (N840, N831, N319);
xor XOR2 (N841, N806, N283);
not NOT1 (N842, N833);
not NOT1 (N843, N835);
or OR3 (N844, N834, N134, N264);
and AND3 (N845, N843, N484, N362);
nor NOR2 (N846, N827, N697);
or OR4 (N847, N837, N139, N74, N781);
buf BUF1 (N848, N846);
buf BUF1 (N849, N840);
xor XOR2 (N850, N847, N116);
nor NOR4 (N851, N850, N109, N811, N758);
nor NOR3 (N852, N844, N798, N119);
and AND4 (N853, N832, N210, N531, N395);
and AND4 (N854, N842, N279, N127, N510);
and AND2 (N855, N854, N165);
and AND3 (N856, N836, N231, N48);
not NOT1 (N857, N849);
buf BUF1 (N858, N857);
nor NOR4 (N859, N839, N835, N703, N34);
and AND3 (N860, N855, N365, N31);
nand NAND3 (N861, N859, N577, N812);
buf BUF1 (N862, N848);
and AND2 (N863, N856, N52);
nor NOR2 (N864, N852, N235);
not NOT1 (N865, N845);
and AND4 (N866, N865, N220, N433, N14);
not NOT1 (N867, N864);
buf BUF1 (N868, N867);
not NOT1 (N869, N851);
xor XOR2 (N870, N860, N468);
nand NAND2 (N871, N869, N111);
or OR4 (N872, N841, N729, N356, N239);
nand NAND3 (N873, N863, N680, N57);
and AND2 (N874, N868, N624);
nand NAND3 (N875, N861, N70, N436);
nand NAND4 (N876, N872, N43, N647, N766);
nor NOR2 (N877, N874, N785);
nand NAND4 (N878, N877, N699, N305, N806);
nand NAND2 (N879, N870, N741);
nor NOR2 (N880, N866, N438);
or OR3 (N881, N873, N185, N779);
nand NAND3 (N882, N875, N29, N540);
and AND2 (N883, N862, N32);
buf BUF1 (N884, N881);
nor NOR2 (N885, N876, N445);
nand NAND3 (N886, N882, N804, N107);
xor XOR2 (N887, N853, N319);
not NOT1 (N888, N886);
or OR2 (N889, N884, N451);
xor XOR2 (N890, N885, N114);
buf BUF1 (N891, N883);
or OR2 (N892, N880, N431);
and AND4 (N893, N879, N287, N276, N563);
and AND4 (N894, N887, N256, N38, N396);
and AND4 (N895, N888, N295, N875, N97);
nand NAND2 (N896, N889, N528);
xor XOR2 (N897, N896, N196);
not NOT1 (N898, N871);
buf BUF1 (N899, N890);
and AND4 (N900, N895, N622, N738, N40);
nand NAND4 (N901, N900, N152, N113, N232);
xor XOR2 (N902, N891, N721);
not NOT1 (N903, N893);
xor XOR2 (N904, N898, N563);
nor NOR3 (N905, N904, N86, N533);
nor NOR2 (N906, N878, N272);
buf BUF1 (N907, N899);
nor NOR4 (N908, N892, N283, N268, N651);
buf BUF1 (N909, N901);
nor NOR4 (N910, N858, N681, N404, N102);
or OR2 (N911, N897, N460);
not NOT1 (N912, N910);
not NOT1 (N913, N912);
and AND2 (N914, N911, N478);
and AND3 (N915, N906, N914, N314);
nand NAND3 (N916, N651, N34, N664);
nor NOR2 (N917, N902, N363);
not NOT1 (N918, N908);
nor NOR4 (N919, N913, N181, N844, N260);
and AND4 (N920, N903, N763, N769, N696);
or OR3 (N921, N918, N404, N895);
or OR4 (N922, N905, N90, N742, N531);
xor XOR2 (N923, N915, N103);
not NOT1 (N924, N919);
xor XOR2 (N925, N924, N19);
not NOT1 (N926, N907);
not NOT1 (N927, N920);
xor XOR2 (N928, N927, N426);
not NOT1 (N929, N928);
not NOT1 (N930, N923);
buf BUF1 (N931, N917);
not NOT1 (N932, N922);
and AND2 (N933, N931, N257);
not NOT1 (N934, N932);
not NOT1 (N935, N926);
not NOT1 (N936, N925);
or OR4 (N937, N921, N33, N751, N668);
xor XOR2 (N938, N937, N237);
nand NAND2 (N939, N936, N320);
nor NOR4 (N940, N916, N670, N211, N859);
buf BUF1 (N941, N935);
xor XOR2 (N942, N929, N800);
and AND4 (N943, N941, N48, N14, N59);
not NOT1 (N944, N909);
nand NAND2 (N945, N942, N325);
and AND4 (N946, N894, N503, N98, N826);
xor XOR2 (N947, N943, N317);
buf BUF1 (N948, N934);
and AND2 (N949, N940, N581);
nor NOR2 (N950, N933, N816);
nor NOR2 (N951, N938, N937);
and AND3 (N952, N947, N754, N306);
not NOT1 (N953, N939);
and AND3 (N954, N930, N205, N27);
nand NAND4 (N955, N945, N921, N478, N940);
or OR4 (N956, N949, N17, N384, N445);
nor NOR3 (N957, N944, N512, N432);
or OR3 (N958, N946, N921, N319);
nor NOR3 (N959, N954, N793, N818);
nor NOR3 (N960, N956, N384, N138);
nand NAND4 (N961, N950, N663, N894, N841);
nand NAND2 (N962, N953, N508);
nand NAND4 (N963, N955, N816, N701, N865);
xor XOR2 (N964, N959, N109);
buf BUF1 (N965, N948);
buf BUF1 (N966, N963);
or OR2 (N967, N958, N15);
buf BUF1 (N968, N951);
and AND4 (N969, N966, N482, N129, N573);
and AND3 (N970, N965, N291, N181);
buf BUF1 (N971, N957);
and AND2 (N972, N969, N507);
nor NOR2 (N973, N972, N812);
xor XOR2 (N974, N967, N434);
not NOT1 (N975, N968);
or OR3 (N976, N973, N431, N313);
or OR4 (N977, N970, N825, N144, N510);
nor NOR4 (N978, N961, N848, N435, N804);
xor XOR2 (N979, N978, N398);
and AND2 (N980, N975, N800);
and AND2 (N981, N976, N420);
xor XOR2 (N982, N974, N190);
and AND4 (N983, N971, N863, N804, N67);
and AND4 (N984, N952, N419, N380, N826);
buf BUF1 (N985, N984);
xor XOR2 (N986, N981, N401);
or OR3 (N987, N982, N163, N631);
xor XOR2 (N988, N985, N262);
nor NOR4 (N989, N987, N136, N405, N925);
xor XOR2 (N990, N960, N375);
not NOT1 (N991, N989);
and AND2 (N992, N983, N740);
nor NOR3 (N993, N991, N410, N167);
or OR2 (N994, N962, N499);
or OR3 (N995, N993, N474, N142);
nor NOR4 (N996, N988, N19, N771, N420);
and AND3 (N997, N994, N274, N326);
xor XOR2 (N998, N995, N496);
nor NOR2 (N999, N992, N1);
or OR2 (N1000, N997, N263);
and AND3 (N1001, N979, N59, N209);
buf BUF1 (N1002, N1001);
xor XOR2 (N1003, N964, N712);
nor NOR2 (N1004, N990, N127);
and AND3 (N1005, N986, N132, N949);
and AND4 (N1006, N1000, N679, N888, N202);
not NOT1 (N1007, N1003);
xor XOR2 (N1008, N1004, N44);
and AND4 (N1009, N1002, N657, N384, N400);
not NOT1 (N1010, N977);
nor NOR3 (N1011, N1007, N148, N241);
not NOT1 (N1012, N1010);
or OR4 (N1013, N1009, N523, N49, N536);
nand NAND4 (N1014, N998, N668, N2, N214);
nand NAND4 (N1015, N999, N352, N977, N107);
or OR2 (N1016, N1006, N311);
not NOT1 (N1017, N1015);
or OR2 (N1018, N1017, N124);
or OR3 (N1019, N1012, N486, N1001);
nor NOR3 (N1020, N1005, N102, N178);
and AND3 (N1021, N1020, N168, N688);
or OR2 (N1022, N1021, N645);
buf BUF1 (N1023, N1013);
buf BUF1 (N1024, N980);
buf BUF1 (N1025, N1024);
nor NOR3 (N1026, N1011, N730, N980);
buf BUF1 (N1027, N1019);
and AND2 (N1028, N1023, N313);
nand NAND3 (N1029, N1028, N40, N248);
nand NAND4 (N1030, N1026, N945, N168, N385);
and AND3 (N1031, N1016, N201, N552);
or OR3 (N1032, N1029, N900, N393);
and AND3 (N1033, N1025, N314, N145);
or OR4 (N1034, N996, N1007, N233, N631);
or OR4 (N1035, N1008, N42, N358, N217);
buf BUF1 (N1036, N1033);
xor XOR2 (N1037, N1031, N431);
buf BUF1 (N1038, N1022);
and AND4 (N1039, N1032, N522, N608, N187);
nor NOR2 (N1040, N1027, N347);
xor XOR2 (N1041, N1037, N401);
nor NOR3 (N1042, N1040, N38, N276);
or OR4 (N1043, N1018, N569, N311, N522);
buf BUF1 (N1044, N1034);
nor NOR4 (N1045, N1044, N753, N676, N71);
not NOT1 (N1046, N1038);
not NOT1 (N1047, N1043);
nand NAND3 (N1048, N1047, N303, N41);
nor NOR3 (N1049, N1041, N176, N638);
or OR4 (N1050, N1048, N597, N1030, N752);
not NOT1 (N1051, N631);
nor NOR4 (N1052, N1049, N230, N505, N542);
not NOT1 (N1053, N1052);
and AND3 (N1054, N1036, N909, N482);
nor NOR4 (N1055, N1014, N295, N384, N682);
or OR2 (N1056, N1039, N743);
or OR2 (N1057, N1053, N586);
and AND2 (N1058, N1035, N172);
nand NAND4 (N1059, N1046, N901, N621, N22);
not NOT1 (N1060, N1054);
nand NAND3 (N1061, N1058, N81, N210);
nand NAND2 (N1062, N1042, N953);
not NOT1 (N1063, N1059);
xor XOR2 (N1064, N1062, N432);
nor NOR3 (N1065, N1051, N572, N832);
nand NAND4 (N1066, N1057, N373, N707, N118);
or OR3 (N1067, N1066, N31, N247);
xor XOR2 (N1068, N1056, N542);
buf BUF1 (N1069, N1060);
not NOT1 (N1070, N1068);
nor NOR2 (N1071, N1065, N1026);
nand NAND4 (N1072, N1069, N1013, N275, N402);
buf BUF1 (N1073, N1055);
nand NAND3 (N1074, N1063, N757, N359);
xor XOR2 (N1075, N1064, N433);
buf BUF1 (N1076, N1067);
xor XOR2 (N1077, N1076, N365);
xor XOR2 (N1078, N1071, N186);
or OR2 (N1079, N1073, N945);
buf BUF1 (N1080, N1072);
or OR3 (N1081, N1079, N724, N877);
nor NOR4 (N1082, N1077, N180, N333, N863);
nand NAND2 (N1083, N1081, N641);
or OR3 (N1084, N1080, N133, N382);
or OR3 (N1085, N1070, N915, N565);
nand NAND4 (N1086, N1082, N415, N191, N88);
not NOT1 (N1087, N1078);
nor NOR4 (N1088, N1085, N821, N995, N16);
nand NAND2 (N1089, N1045, N53);
and AND2 (N1090, N1086, N189);
buf BUF1 (N1091, N1088);
xor XOR2 (N1092, N1090, N464);
or OR3 (N1093, N1061, N293, N242);
not NOT1 (N1094, N1092);
not NOT1 (N1095, N1083);
or OR3 (N1096, N1089, N242, N727);
xor XOR2 (N1097, N1050, N705);
and AND3 (N1098, N1074, N135, N1016);
and AND2 (N1099, N1097, N242);
nor NOR2 (N1100, N1091, N483);
or OR4 (N1101, N1099, N31, N644, N1038);
xor XOR2 (N1102, N1096, N219);
nor NOR2 (N1103, N1084, N268);
xor XOR2 (N1104, N1101, N711);
and AND4 (N1105, N1102, N12, N763, N443);
or OR3 (N1106, N1104, N299, N744);
xor XOR2 (N1107, N1087, N713);
and AND3 (N1108, N1098, N460, N1009);
and AND3 (N1109, N1103, N427, N1050);
or OR2 (N1110, N1106, N115);
and AND4 (N1111, N1108, N355, N619, N403);
nand NAND4 (N1112, N1094, N1064, N60, N631);
buf BUF1 (N1113, N1100);
and AND4 (N1114, N1109, N794, N514, N1063);
xor XOR2 (N1115, N1093, N75);
nor NOR4 (N1116, N1111, N545, N1043, N901);
xor XOR2 (N1117, N1115, N611);
and AND2 (N1118, N1116, N236);
or OR4 (N1119, N1107, N867, N553, N573);
and AND2 (N1120, N1112, N710);
nor NOR4 (N1121, N1118, N509, N67, N1094);
nor NOR2 (N1122, N1075, N18);
not NOT1 (N1123, N1110);
nand NAND2 (N1124, N1105, N1059);
and AND2 (N1125, N1120, N996);
nand NAND2 (N1126, N1125, N214);
nor NOR3 (N1127, N1113, N121, N291);
buf BUF1 (N1128, N1127);
xor XOR2 (N1129, N1126, N203);
nor NOR2 (N1130, N1117, N438);
xor XOR2 (N1131, N1119, N713);
not NOT1 (N1132, N1130);
or OR4 (N1133, N1131, N1099, N143, N320);
xor XOR2 (N1134, N1095, N599);
and AND3 (N1135, N1122, N358, N551);
nor NOR4 (N1136, N1133, N899, N928, N611);
not NOT1 (N1137, N1135);
nand NAND4 (N1138, N1124, N76, N909, N275);
not NOT1 (N1139, N1129);
buf BUF1 (N1140, N1132);
or OR2 (N1141, N1134, N77);
and AND3 (N1142, N1140, N660, N999);
or OR3 (N1143, N1141, N774, N938);
nand NAND4 (N1144, N1138, N916, N125, N293);
buf BUF1 (N1145, N1142);
not NOT1 (N1146, N1144);
nand NAND4 (N1147, N1128, N113, N317, N1079);
nor NOR3 (N1148, N1114, N70, N1043);
xor XOR2 (N1149, N1123, N612);
or OR2 (N1150, N1147, N658);
and AND2 (N1151, N1150, N227);
buf BUF1 (N1152, N1145);
nor NOR4 (N1153, N1152, N177, N1011, N223);
and AND2 (N1154, N1136, N134);
nand NAND4 (N1155, N1146, N171, N211, N543);
or OR3 (N1156, N1153, N897, N531);
or OR2 (N1157, N1137, N407);
or OR2 (N1158, N1156, N862);
nor NOR3 (N1159, N1151, N1138, N844);
buf BUF1 (N1160, N1159);
buf BUF1 (N1161, N1139);
xor XOR2 (N1162, N1148, N512);
xor XOR2 (N1163, N1162, N612);
or OR4 (N1164, N1121, N1095, N749, N840);
not NOT1 (N1165, N1157);
xor XOR2 (N1166, N1154, N681);
xor XOR2 (N1167, N1158, N746);
or OR3 (N1168, N1149, N983, N162);
nand NAND2 (N1169, N1143, N913);
not NOT1 (N1170, N1163);
and AND2 (N1171, N1167, N1093);
nand NAND3 (N1172, N1169, N425, N1115);
nand NAND3 (N1173, N1172, N704, N186);
not NOT1 (N1174, N1171);
nor NOR3 (N1175, N1164, N357, N86);
buf BUF1 (N1176, N1170);
and AND2 (N1177, N1165, N603);
not NOT1 (N1178, N1174);
nor NOR2 (N1179, N1168, N1061);
and AND3 (N1180, N1161, N1036, N1056);
xor XOR2 (N1181, N1155, N432);
or OR2 (N1182, N1180, N203);
or OR2 (N1183, N1179, N469);
and AND4 (N1184, N1173, N65, N76, N1);
nand NAND4 (N1185, N1178, N997, N465, N431);
not NOT1 (N1186, N1177);
not NOT1 (N1187, N1183);
nand NAND4 (N1188, N1160, N681, N1141, N854);
or OR2 (N1189, N1186, N245);
xor XOR2 (N1190, N1182, N82);
and AND4 (N1191, N1187, N845, N915, N705);
buf BUF1 (N1192, N1176);
and AND3 (N1193, N1184, N90, N593);
buf BUF1 (N1194, N1181);
not NOT1 (N1195, N1166);
nand NAND2 (N1196, N1175, N975);
nor NOR4 (N1197, N1188, N309, N1010, N1115);
and AND3 (N1198, N1190, N241, N1062);
or OR4 (N1199, N1195, N879, N82, N710);
and AND4 (N1200, N1196, N210, N701, N591);
not NOT1 (N1201, N1200);
xor XOR2 (N1202, N1185, N672);
nand NAND3 (N1203, N1202, N881, N1151);
buf BUF1 (N1204, N1197);
nand NAND3 (N1205, N1194, N522, N933);
and AND4 (N1206, N1193, N207, N282, N69);
or OR3 (N1207, N1191, N421, N767);
nand NAND3 (N1208, N1201, N556, N618);
xor XOR2 (N1209, N1206, N456);
or OR4 (N1210, N1189, N131, N873, N13);
buf BUF1 (N1211, N1198);
buf BUF1 (N1212, N1192);
or OR4 (N1213, N1208, N957, N687, N895);
and AND3 (N1214, N1207, N821, N642);
or OR2 (N1215, N1209, N40);
not NOT1 (N1216, N1210);
or OR4 (N1217, N1205, N741, N169, N905);
xor XOR2 (N1218, N1214, N766);
not NOT1 (N1219, N1211);
buf BUF1 (N1220, N1204);
buf BUF1 (N1221, N1220);
buf BUF1 (N1222, N1213);
or OR3 (N1223, N1216, N1187, N1191);
buf BUF1 (N1224, N1215);
nand NAND2 (N1225, N1203, N53);
buf BUF1 (N1226, N1223);
nor NOR2 (N1227, N1224, N804);
not NOT1 (N1228, N1217);
xor XOR2 (N1229, N1222, N90);
nor NOR4 (N1230, N1228, N1150, N478, N60);
or OR3 (N1231, N1230, N520, N808);
not NOT1 (N1232, N1199);
nand NAND4 (N1233, N1231, N168, N49, N629);
xor XOR2 (N1234, N1219, N25);
xor XOR2 (N1235, N1233, N725);
not NOT1 (N1236, N1225);
nor NOR4 (N1237, N1226, N472, N948, N1154);
not NOT1 (N1238, N1237);
nand NAND2 (N1239, N1232, N585);
not NOT1 (N1240, N1234);
and AND4 (N1241, N1240, N1052, N379, N1203);
or OR2 (N1242, N1212, N224);
nor NOR2 (N1243, N1218, N727);
xor XOR2 (N1244, N1221, N118);
buf BUF1 (N1245, N1227);
buf BUF1 (N1246, N1229);
nand NAND3 (N1247, N1241, N208, N577);
not NOT1 (N1248, N1245);
not NOT1 (N1249, N1239);
and AND2 (N1250, N1243, N717);
nand NAND2 (N1251, N1247, N1184);
or OR2 (N1252, N1242, N1232);
nand NAND4 (N1253, N1249, N143, N394, N689);
buf BUF1 (N1254, N1253);
buf BUF1 (N1255, N1250);
xor XOR2 (N1256, N1235, N25);
buf BUF1 (N1257, N1246);
xor XOR2 (N1258, N1238, N1005);
nor NOR3 (N1259, N1255, N842, N691);
nor NOR2 (N1260, N1258, N837);
and AND4 (N1261, N1260, N135, N594, N564);
or OR2 (N1262, N1251, N888);
not NOT1 (N1263, N1256);
xor XOR2 (N1264, N1254, N477);
and AND2 (N1265, N1236, N901);
and AND2 (N1266, N1248, N727);
nor NOR4 (N1267, N1262, N1202, N7, N1266);
or OR2 (N1268, N121, N274);
nor NOR4 (N1269, N1252, N511, N448, N667);
nand NAND3 (N1270, N1244, N511, N377);
nand NAND3 (N1271, N1261, N1094, N834);
and AND4 (N1272, N1268, N92, N956, N1238);
xor XOR2 (N1273, N1269, N291);
or OR4 (N1274, N1271, N1009, N908, N1035);
or OR3 (N1275, N1257, N551, N332);
or OR2 (N1276, N1263, N837);
nor NOR2 (N1277, N1270, N421);
nor NOR4 (N1278, N1264, N507, N482, N848);
xor XOR2 (N1279, N1278, N395);
and AND4 (N1280, N1279, N1001, N636, N456);
and AND4 (N1281, N1259, N1179, N630, N1048);
nor NOR3 (N1282, N1275, N259, N679);
nor NOR4 (N1283, N1281, N421, N979, N817);
or OR4 (N1284, N1276, N93, N100, N356);
and AND2 (N1285, N1284, N251);
or OR4 (N1286, N1283, N871, N655, N294);
nor NOR3 (N1287, N1272, N231, N392);
nor NOR3 (N1288, N1274, N1, N1054);
or OR3 (N1289, N1280, N142, N568);
and AND4 (N1290, N1265, N144, N607, N672);
not NOT1 (N1291, N1273);
or OR3 (N1292, N1289, N1217, N724);
not NOT1 (N1293, N1287);
nand NAND2 (N1294, N1282, N592);
buf BUF1 (N1295, N1294);
not NOT1 (N1296, N1291);
and AND2 (N1297, N1293, N1111);
not NOT1 (N1298, N1295);
not NOT1 (N1299, N1267);
or OR2 (N1300, N1292, N1287);
and AND4 (N1301, N1298, N311, N40, N747);
xor XOR2 (N1302, N1277, N421);
and AND3 (N1303, N1285, N996, N509);
nand NAND4 (N1304, N1300, N18, N1187, N1199);
not NOT1 (N1305, N1301);
nor NOR3 (N1306, N1288, N574, N730);
nor NOR2 (N1307, N1297, N851);
or OR2 (N1308, N1305, N1051);
xor XOR2 (N1309, N1290, N1176);
and AND4 (N1310, N1309, N1284, N279, N1254);
nand NAND2 (N1311, N1296, N1261);
buf BUF1 (N1312, N1311);
nand NAND4 (N1313, N1306, N904, N1021, N1152);
nand NAND4 (N1314, N1313, N274, N456, N1197);
nor NOR2 (N1315, N1307, N1077);
or OR3 (N1316, N1299, N1213, N824);
xor XOR2 (N1317, N1302, N736);
or OR3 (N1318, N1317, N941, N91);
or OR2 (N1319, N1303, N789);
xor XOR2 (N1320, N1316, N1289);
or OR3 (N1321, N1320, N237, N344);
and AND4 (N1322, N1304, N1040, N1120, N803);
xor XOR2 (N1323, N1319, N692);
nand NAND3 (N1324, N1286, N1280, N356);
nor NOR4 (N1325, N1324, N149, N578, N587);
nor NOR2 (N1326, N1310, N1266);
not NOT1 (N1327, N1312);
not NOT1 (N1328, N1314);
not NOT1 (N1329, N1328);
buf BUF1 (N1330, N1329);
buf BUF1 (N1331, N1315);
xor XOR2 (N1332, N1321, N880);
buf BUF1 (N1333, N1325);
not NOT1 (N1334, N1308);
and AND2 (N1335, N1327, N827);
buf BUF1 (N1336, N1334);
nor NOR3 (N1337, N1326, N375, N494);
or OR3 (N1338, N1337, N640, N1131);
nor NOR4 (N1339, N1330, N917, N651, N862);
or OR2 (N1340, N1339, N49);
nor NOR4 (N1341, N1332, N797, N1163, N745);
and AND4 (N1342, N1340, N1305, N364, N1012);
nor NOR3 (N1343, N1323, N466, N933);
or OR3 (N1344, N1341, N993, N170);
and AND2 (N1345, N1335, N234);
xor XOR2 (N1346, N1333, N414);
nand NAND4 (N1347, N1343, N469, N1247, N498);
nor NOR3 (N1348, N1342, N588, N1114);
xor XOR2 (N1349, N1347, N505);
or OR2 (N1350, N1348, N1281);
or OR2 (N1351, N1322, N979);
nand NAND4 (N1352, N1346, N389, N641, N1150);
nor NOR3 (N1353, N1349, N1153, N415);
not NOT1 (N1354, N1336);
not NOT1 (N1355, N1318);
and AND4 (N1356, N1345, N570, N299, N591);
nand NAND3 (N1357, N1338, N1087, N603);
buf BUF1 (N1358, N1357);
nor NOR3 (N1359, N1356, N460, N1351);
and AND4 (N1360, N752, N231, N1117, N715);
nor NOR3 (N1361, N1360, N843, N1097);
nand NAND2 (N1362, N1350, N426);
nand NAND4 (N1363, N1352, N360, N240, N1321);
nor NOR4 (N1364, N1353, N267, N397, N377);
nor NOR2 (N1365, N1331, N1080);
buf BUF1 (N1366, N1364);
buf BUF1 (N1367, N1366);
buf BUF1 (N1368, N1354);
or OR2 (N1369, N1355, N135);
xor XOR2 (N1370, N1358, N2);
buf BUF1 (N1371, N1359);
buf BUF1 (N1372, N1370);
xor XOR2 (N1373, N1371, N917);
nand NAND2 (N1374, N1344, N1140);
and AND3 (N1375, N1372, N426, N161);
or OR3 (N1376, N1367, N660, N972);
nand NAND4 (N1377, N1368, N1236, N1335, N710);
and AND3 (N1378, N1374, N1110, N435);
nand NAND4 (N1379, N1362, N819, N812, N227);
buf BUF1 (N1380, N1377);
not NOT1 (N1381, N1363);
nand NAND3 (N1382, N1378, N405, N963);
and AND3 (N1383, N1361, N980, N498);
nor NOR2 (N1384, N1382, N685);
buf BUF1 (N1385, N1376);
not NOT1 (N1386, N1373);
or OR3 (N1387, N1381, N368, N103);
nand NAND4 (N1388, N1387, N754, N1048, N383);
xor XOR2 (N1389, N1383, N516);
xor XOR2 (N1390, N1380, N158);
not NOT1 (N1391, N1379);
xor XOR2 (N1392, N1388, N1085);
buf BUF1 (N1393, N1391);
not NOT1 (N1394, N1365);
xor XOR2 (N1395, N1389, N62);
nand NAND4 (N1396, N1386, N1393, N396, N203);
buf BUF1 (N1397, N77);
nand NAND3 (N1398, N1390, N583, N936);
or OR2 (N1399, N1394, N382);
nor NOR2 (N1400, N1384, N205);
nor NOR2 (N1401, N1395, N416);
nand NAND3 (N1402, N1375, N364, N532);
buf BUF1 (N1403, N1385);
buf BUF1 (N1404, N1402);
nand NAND4 (N1405, N1404, N1046, N72, N1160);
not NOT1 (N1406, N1403);
and AND4 (N1407, N1392, N467, N960, N1404);
buf BUF1 (N1408, N1406);
and AND2 (N1409, N1400, N1396);
xor XOR2 (N1410, N374, N1043);
buf BUF1 (N1411, N1399);
or OR4 (N1412, N1408, N87, N334, N1111);
and AND4 (N1413, N1405, N720, N1027, N509);
buf BUF1 (N1414, N1410);
or OR2 (N1415, N1411, N372);
xor XOR2 (N1416, N1413, N1102);
xor XOR2 (N1417, N1414, N976);
not NOT1 (N1418, N1412);
buf BUF1 (N1419, N1416);
nand NAND2 (N1420, N1415, N1358);
and AND4 (N1421, N1417, N1205, N1018, N705);
buf BUF1 (N1422, N1420);
nand NAND2 (N1423, N1421, N747);
xor XOR2 (N1424, N1409, N237);
buf BUF1 (N1425, N1407);
nand NAND4 (N1426, N1422, N683, N1416, N564);
xor XOR2 (N1427, N1424, N486);
nor NOR4 (N1428, N1426, N899, N70, N300);
buf BUF1 (N1429, N1398);
nor NOR4 (N1430, N1397, N1030, N667, N246);
nand NAND4 (N1431, N1419, N1127, N1223, N1178);
buf BUF1 (N1432, N1401);
and AND4 (N1433, N1431, N675, N875, N86);
nor NOR4 (N1434, N1430, N958, N1135, N89);
xor XOR2 (N1435, N1425, N70);
and AND4 (N1436, N1433, N992, N749, N880);
not NOT1 (N1437, N1423);
or OR4 (N1438, N1418, N675, N1247, N971);
nor NOR4 (N1439, N1435, N752, N863, N1236);
nand NAND3 (N1440, N1437, N571, N883);
xor XOR2 (N1441, N1436, N878);
nor NOR4 (N1442, N1434, N1032, N282, N130);
or OR2 (N1443, N1432, N269);
nor NOR2 (N1444, N1429, N176);
or OR3 (N1445, N1444, N1166, N880);
nor NOR4 (N1446, N1441, N1352, N1262, N576);
xor XOR2 (N1447, N1442, N826);
buf BUF1 (N1448, N1427);
nor NOR4 (N1449, N1445, N971, N782, N108);
xor XOR2 (N1450, N1443, N353);
and AND4 (N1451, N1369, N608, N1099, N1289);
not NOT1 (N1452, N1439);
not NOT1 (N1453, N1440);
xor XOR2 (N1454, N1448, N663);
nand NAND4 (N1455, N1438, N270, N1288, N1148);
or OR2 (N1456, N1446, N1384);
and AND4 (N1457, N1451, N1345, N75, N280);
and AND4 (N1458, N1453, N1305, N329, N976);
or OR3 (N1459, N1447, N632, N712);
nand NAND3 (N1460, N1449, N485, N560);
and AND2 (N1461, N1457, N268);
buf BUF1 (N1462, N1459);
or OR3 (N1463, N1428, N1358, N1341);
buf BUF1 (N1464, N1455);
and AND2 (N1465, N1458, N379);
nand NAND2 (N1466, N1456, N1144);
or OR2 (N1467, N1466, N733);
nor NOR2 (N1468, N1460, N1197);
or OR3 (N1469, N1462, N920, N618);
nor NOR4 (N1470, N1469, N1387, N962, N932);
nand NAND4 (N1471, N1461, N1424, N455, N165);
nor NOR2 (N1472, N1470, N415);
buf BUF1 (N1473, N1472);
buf BUF1 (N1474, N1464);
nor NOR2 (N1475, N1450, N1119);
buf BUF1 (N1476, N1475);
nor NOR3 (N1477, N1473, N164, N215);
or OR2 (N1478, N1471, N34);
nor NOR4 (N1479, N1465, N1192, N823, N834);
nand NAND4 (N1480, N1454, N194, N1137, N508);
nand NAND2 (N1481, N1476, N891);
nor NOR3 (N1482, N1474, N109, N1133);
and AND3 (N1483, N1479, N433, N714);
xor XOR2 (N1484, N1468, N668);
xor XOR2 (N1485, N1481, N354);
buf BUF1 (N1486, N1480);
or OR4 (N1487, N1463, N447, N1153, N298);
or OR3 (N1488, N1477, N224, N749);
not NOT1 (N1489, N1478);
xor XOR2 (N1490, N1467, N981);
and AND4 (N1491, N1486, N895, N695, N511);
nor NOR3 (N1492, N1484, N1038, N745);
and AND4 (N1493, N1492, N365, N924, N1316);
or OR2 (N1494, N1482, N84);
nor NOR2 (N1495, N1489, N1419);
nor NOR3 (N1496, N1491, N989, N644);
xor XOR2 (N1497, N1495, N627);
nor NOR4 (N1498, N1452, N967, N1156, N340);
xor XOR2 (N1499, N1485, N1155);
xor XOR2 (N1500, N1488, N483);
xor XOR2 (N1501, N1498, N1470);
or OR3 (N1502, N1496, N516, N382);
xor XOR2 (N1503, N1483, N567);
nand NAND3 (N1504, N1503, N1089, N6);
and AND3 (N1505, N1499, N545, N473);
nor NOR4 (N1506, N1490, N982, N352, N1409);
nand NAND2 (N1507, N1504, N895);
and AND2 (N1508, N1497, N1126);
or OR3 (N1509, N1507, N1502, N961);
not NOT1 (N1510, N1005);
buf BUF1 (N1511, N1494);
and AND2 (N1512, N1501, N81);
or OR4 (N1513, N1493, N439, N531, N566);
nor NOR3 (N1514, N1510, N1170, N995);
or OR4 (N1515, N1509, N527, N36, N741);
nand NAND2 (N1516, N1512, N1491);
or OR4 (N1517, N1500, N936, N747, N1242);
xor XOR2 (N1518, N1515, N613);
not NOT1 (N1519, N1487);
nand NAND4 (N1520, N1517, N123, N1366, N625);
xor XOR2 (N1521, N1513, N1359);
buf BUF1 (N1522, N1506);
and AND3 (N1523, N1505, N20, N1140);
or OR3 (N1524, N1516, N110, N1009);
and AND3 (N1525, N1511, N565, N1003);
and AND4 (N1526, N1525, N1416, N575, N1056);
or OR4 (N1527, N1514, N1199, N1487, N1065);
not NOT1 (N1528, N1521);
not NOT1 (N1529, N1520);
and AND2 (N1530, N1526, N394);
nor NOR2 (N1531, N1522, N244);
and AND2 (N1532, N1524, N1065);
and AND3 (N1533, N1527, N499, N1242);
not NOT1 (N1534, N1531);
buf BUF1 (N1535, N1508);
not NOT1 (N1536, N1530);
xor XOR2 (N1537, N1532, N446);
not NOT1 (N1538, N1523);
buf BUF1 (N1539, N1533);
nor NOR3 (N1540, N1518, N1262, N1163);
nor NOR4 (N1541, N1529, N848, N227, N417);
buf BUF1 (N1542, N1540);
nor NOR3 (N1543, N1539, N171, N1459);
not NOT1 (N1544, N1535);
and AND4 (N1545, N1542, N22, N696, N572);
xor XOR2 (N1546, N1541, N784);
or OR3 (N1547, N1519, N211, N874);
or OR4 (N1548, N1543, N625, N1127, N252);
xor XOR2 (N1549, N1544, N931);
xor XOR2 (N1550, N1534, N540);
or OR3 (N1551, N1546, N1193, N1499);
nor NOR3 (N1552, N1547, N135, N90);
nand NAND2 (N1553, N1550, N739);
nand NAND2 (N1554, N1549, N347);
xor XOR2 (N1555, N1553, N1545);
nand NAND4 (N1556, N282, N623, N1553, N560);
buf BUF1 (N1557, N1555);
and AND3 (N1558, N1548, N409, N45);
nor NOR3 (N1559, N1557, N1503, N210);
nor NOR2 (N1560, N1537, N860);
not NOT1 (N1561, N1554);
nor NOR4 (N1562, N1559, N1340, N900, N704);
not NOT1 (N1563, N1536);
not NOT1 (N1564, N1552);
and AND3 (N1565, N1551, N363, N1227);
nand NAND3 (N1566, N1528, N1400, N435);
xor XOR2 (N1567, N1561, N309);
nor NOR4 (N1568, N1556, N1121, N683, N138);
and AND3 (N1569, N1538, N1119, N629);
and AND2 (N1570, N1567, N1080);
and AND2 (N1571, N1565, N1289);
and AND2 (N1572, N1558, N100);
or OR3 (N1573, N1564, N1358, N164);
or OR3 (N1574, N1560, N1411, N1493);
and AND2 (N1575, N1563, N531);
xor XOR2 (N1576, N1572, N1444);
nand NAND3 (N1577, N1566, N502, N245);
xor XOR2 (N1578, N1574, N824);
xor XOR2 (N1579, N1569, N779);
nor NOR3 (N1580, N1579, N1026, N850);
or OR4 (N1581, N1577, N999, N1216, N55);
or OR3 (N1582, N1571, N1428, N435);
and AND2 (N1583, N1576, N830);
nor NOR2 (N1584, N1570, N125);
not NOT1 (N1585, N1583);
not NOT1 (N1586, N1584);
nor NOR3 (N1587, N1578, N354, N802);
nor NOR4 (N1588, N1585, N259, N309, N701);
buf BUF1 (N1589, N1587);
nor NOR2 (N1590, N1588, N1033);
or OR2 (N1591, N1581, N1579);
xor XOR2 (N1592, N1575, N1004);
nand NAND4 (N1593, N1580, N560, N1523, N349);
xor XOR2 (N1594, N1592, N792);
and AND4 (N1595, N1589, N1512, N1479, N1308);
nor NOR2 (N1596, N1568, N573);
nand NAND3 (N1597, N1593, N1083, N818);
xor XOR2 (N1598, N1597, N22);
or OR3 (N1599, N1562, N406, N967);
xor XOR2 (N1600, N1582, N948);
nor NOR3 (N1601, N1600, N1340, N1311);
xor XOR2 (N1602, N1599, N69);
or OR3 (N1603, N1586, N1267, N1154);
not NOT1 (N1604, N1596);
buf BUF1 (N1605, N1601);
not NOT1 (N1606, N1602);
not NOT1 (N1607, N1573);
not NOT1 (N1608, N1606);
not NOT1 (N1609, N1605);
not NOT1 (N1610, N1598);
buf BUF1 (N1611, N1603);
nand NAND4 (N1612, N1595, N461, N368, N738);
nand NAND4 (N1613, N1608, N1563, N923, N1490);
buf BUF1 (N1614, N1604);
not NOT1 (N1615, N1614);
buf BUF1 (N1616, N1615);
nand NAND3 (N1617, N1607, N1208, N876);
and AND4 (N1618, N1591, N1332, N1120, N1133);
nor NOR4 (N1619, N1611, N1426, N1389, N356);
buf BUF1 (N1620, N1618);
nand NAND2 (N1621, N1620, N234);
or OR3 (N1622, N1590, N97, N212);
buf BUF1 (N1623, N1621);
not NOT1 (N1624, N1622);
buf BUF1 (N1625, N1609);
buf BUF1 (N1626, N1594);
or OR2 (N1627, N1626, N801);
xor XOR2 (N1628, N1612, N1604);
nand NAND3 (N1629, N1619, N1529, N823);
or OR4 (N1630, N1623, N871, N48, N297);
not NOT1 (N1631, N1630);
buf BUF1 (N1632, N1631);
or OR3 (N1633, N1629, N803, N1251);
buf BUF1 (N1634, N1628);
or OR2 (N1635, N1633, N757);
and AND3 (N1636, N1634, N181, N496);
not NOT1 (N1637, N1632);
and AND2 (N1638, N1616, N669);
not NOT1 (N1639, N1636);
and AND2 (N1640, N1624, N1560);
and AND4 (N1641, N1637, N1052, N1002, N51);
xor XOR2 (N1642, N1625, N1533);
and AND3 (N1643, N1641, N1487, N792);
or OR2 (N1644, N1617, N1512);
buf BUF1 (N1645, N1642);
nand NAND3 (N1646, N1635, N1390, N48);
nor NOR2 (N1647, N1643, N1405);
buf BUF1 (N1648, N1640);
not NOT1 (N1649, N1645);
xor XOR2 (N1650, N1649, N1116);
and AND3 (N1651, N1627, N1638, N513);
nor NOR3 (N1652, N1387, N764, N1123);
or OR3 (N1653, N1644, N814, N1000);
buf BUF1 (N1654, N1653);
nor NOR2 (N1655, N1651, N815);
buf BUF1 (N1656, N1646);
nor NOR2 (N1657, N1652, N945);
nand NAND3 (N1658, N1639, N1285, N1006);
or OR3 (N1659, N1647, N902, N72);
nor NOR4 (N1660, N1648, N888, N1562, N29);
and AND2 (N1661, N1610, N633);
and AND3 (N1662, N1650, N1084, N1171);
nor NOR3 (N1663, N1655, N670, N47);
or OR3 (N1664, N1662, N1430, N34);
nor NOR2 (N1665, N1613, N270);
not NOT1 (N1666, N1659);
and AND2 (N1667, N1657, N1000);
and AND3 (N1668, N1666, N1131, N1166);
nor NOR3 (N1669, N1658, N568, N1194);
not NOT1 (N1670, N1663);
or OR3 (N1671, N1669, N304, N875);
nand NAND2 (N1672, N1660, N1134);
nor NOR2 (N1673, N1668, N1210);
not NOT1 (N1674, N1673);
or OR3 (N1675, N1670, N1064, N410);
xor XOR2 (N1676, N1675, N66);
not NOT1 (N1677, N1672);
nand NAND2 (N1678, N1654, N429);
xor XOR2 (N1679, N1678, N1446);
not NOT1 (N1680, N1679);
nor NOR3 (N1681, N1680, N821, N1086);
or OR4 (N1682, N1656, N766, N982, N202);
or OR4 (N1683, N1676, N498, N1458, N287);
nand NAND2 (N1684, N1682, N1353);
and AND3 (N1685, N1665, N1512, N1404);
xor XOR2 (N1686, N1667, N373);
buf BUF1 (N1687, N1681);
buf BUF1 (N1688, N1687);
or OR3 (N1689, N1661, N832, N1614);
xor XOR2 (N1690, N1688, N1514);
nand NAND4 (N1691, N1664, N1646, N470, N1121);
nand NAND4 (N1692, N1686, N970, N845, N204);
and AND3 (N1693, N1684, N431, N1459);
nor NOR3 (N1694, N1674, N902, N771);
not NOT1 (N1695, N1694);
buf BUF1 (N1696, N1671);
xor XOR2 (N1697, N1683, N1225);
xor XOR2 (N1698, N1685, N226);
buf BUF1 (N1699, N1695);
buf BUF1 (N1700, N1697);
not NOT1 (N1701, N1689);
nand NAND3 (N1702, N1693, N783, N559);
buf BUF1 (N1703, N1698);
or OR2 (N1704, N1702, N1117);
not NOT1 (N1705, N1703);
or OR2 (N1706, N1691, N757);
xor XOR2 (N1707, N1699, N692);
and AND3 (N1708, N1696, N740, N1430);
and AND2 (N1709, N1708, N1499);
xor XOR2 (N1710, N1690, N1125);
buf BUF1 (N1711, N1701);
and AND4 (N1712, N1677, N1574, N532, N693);
buf BUF1 (N1713, N1707);
nand NAND4 (N1714, N1706, N919, N537, N781);
not NOT1 (N1715, N1709);
nor NOR3 (N1716, N1715, N530, N1285);
not NOT1 (N1717, N1692);
nand NAND2 (N1718, N1700, N1008);
nand NAND4 (N1719, N1705, N659, N1714, N1496);
xor XOR2 (N1720, N214, N1134);
nor NOR3 (N1721, N1719, N765, N493);
xor XOR2 (N1722, N1710, N1553);
not NOT1 (N1723, N1713);
nand NAND3 (N1724, N1721, N1099, N1436);
nand NAND4 (N1725, N1716, N867, N390, N508);
nor NOR2 (N1726, N1717, N930);
buf BUF1 (N1727, N1726);
nand NAND3 (N1728, N1704, N276, N1632);
not NOT1 (N1729, N1711);
xor XOR2 (N1730, N1720, N1413);
nor NOR2 (N1731, N1729, N462);
xor XOR2 (N1732, N1725, N302);
and AND3 (N1733, N1718, N1576, N1280);
and AND3 (N1734, N1733, N1272, N812);
nand NAND3 (N1735, N1727, N264, N1371);
buf BUF1 (N1736, N1712);
or OR4 (N1737, N1736, N571, N1130, N1232);
not NOT1 (N1738, N1735);
nand NAND4 (N1739, N1738, N6, N469, N586);
buf BUF1 (N1740, N1731);
nand NAND4 (N1741, N1723, N1442, N1460, N345);
buf BUF1 (N1742, N1741);
nor NOR4 (N1743, N1737, N151, N550, N1072);
nand NAND3 (N1744, N1732, N1665, N309);
nand NAND4 (N1745, N1742, N1227, N1427, N1438);
nor NOR4 (N1746, N1745, N1063, N910, N300);
not NOT1 (N1747, N1722);
not NOT1 (N1748, N1744);
nor NOR2 (N1749, N1724, N394);
or OR4 (N1750, N1728, N896, N805, N474);
or OR4 (N1751, N1747, N1595, N1524, N1298);
xor XOR2 (N1752, N1743, N935);
nand NAND3 (N1753, N1740, N250, N1606);
not NOT1 (N1754, N1739);
nand NAND3 (N1755, N1750, N202, N366);
and AND2 (N1756, N1752, N1185);
and AND4 (N1757, N1734, N1729, N252, N621);
buf BUF1 (N1758, N1746);
and AND4 (N1759, N1758, N982, N1454, N1527);
not NOT1 (N1760, N1754);
nor NOR2 (N1761, N1759, N563);
buf BUF1 (N1762, N1748);
nor NOR3 (N1763, N1753, N976, N1466);
or OR3 (N1764, N1730, N79, N1549);
or OR3 (N1765, N1761, N10, N886);
and AND3 (N1766, N1755, N1710, N485);
not NOT1 (N1767, N1765);
or OR2 (N1768, N1760, N431);
or OR2 (N1769, N1764, N1217);
xor XOR2 (N1770, N1756, N304);
xor XOR2 (N1771, N1763, N1600);
nand NAND3 (N1772, N1749, N1330, N715);
and AND4 (N1773, N1772, N1128, N633, N845);
not NOT1 (N1774, N1757);
xor XOR2 (N1775, N1769, N1461);
buf BUF1 (N1776, N1762);
not NOT1 (N1777, N1768);
xor XOR2 (N1778, N1776, N89);
xor XOR2 (N1779, N1774, N956);
buf BUF1 (N1780, N1773);
nand NAND4 (N1781, N1777, N1380, N114, N1709);
xor XOR2 (N1782, N1778, N114);
and AND3 (N1783, N1780, N201, N1464);
or OR4 (N1784, N1771, N1180, N701, N1269);
not NOT1 (N1785, N1767);
buf BUF1 (N1786, N1782);
nor NOR4 (N1787, N1779, N855, N1497, N603);
nor NOR4 (N1788, N1785, N1295, N612, N633);
not NOT1 (N1789, N1784);
buf BUF1 (N1790, N1787);
and AND4 (N1791, N1786, N1082, N1222, N1261);
xor XOR2 (N1792, N1781, N1513);
and AND4 (N1793, N1766, N1328, N33, N1368);
nand NAND4 (N1794, N1770, N930, N767, N1213);
buf BUF1 (N1795, N1751);
nand NAND3 (N1796, N1789, N1764, N187);
buf BUF1 (N1797, N1793);
xor XOR2 (N1798, N1795, N371);
nand NAND3 (N1799, N1792, N1564, N250);
not NOT1 (N1800, N1790);
buf BUF1 (N1801, N1798);
xor XOR2 (N1802, N1791, N509);
nor NOR3 (N1803, N1796, N204, N480);
nor NOR3 (N1804, N1797, N488, N1433);
nand NAND3 (N1805, N1775, N1486, N153);
buf BUF1 (N1806, N1803);
and AND2 (N1807, N1783, N872);
not NOT1 (N1808, N1801);
not NOT1 (N1809, N1804);
buf BUF1 (N1810, N1794);
buf BUF1 (N1811, N1800);
buf BUF1 (N1812, N1807);
buf BUF1 (N1813, N1812);
nor NOR2 (N1814, N1808, N925);
xor XOR2 (N1815, N1806, N1121);
and AND2 (N1816, N1788, N960);
buf BUF1 (N1817, N1814);
nand NAND2 (N1818, N1809, N1747);
buf BUF1 (N1819, N1810);
buf BUF1 (N1820, N1817);
xor XOR2 (N1821, N1799, N526);
not NOT1 (N1822, N1818);
nor NOR4 (N1823, N1813, N200, N1414, N27);
xor XOR2 (N1824, N1823, N1386);
buf BUF1 (N1825, N1819);
nand NAND3 (N1826, N1805, N405, N1818);
xor XOR2 (N1827, N1822, N1607);
buf BUF1 (N1828, N1802);
nor NOR4 (N1829, N1825, N686, N1035, N241);
xor XOR2 (N1830, N1811, N237);
nand NAND3 (N1831, N1821, N758, N537);
not NOT1 (N1832, N1820);
nor NOR2 (N1833, N1828, N1336);
nor NOR4 (N1834, N1831, N1669, N1261, N476);
or OR4 (N1835, N1824, N808, N204, N257);
nand NAND4 (N1836, N1829, N1274, N951, N1160);
nand NAND4 (N1837, N1826, N1244, N1216, N1713);
not NOT1 (N1838, N1815);
not NOT1 (N1839, N1834);
or OR2 (N1840, N1838, N1500);
or OR3 (N1841, N1840, N890, N436);
not NOT1 (N1842, N1827);
nand NAND2 (N1843, N1839, N616);
nor NOR4 (N1844, N1841, N736, N1547, N1531);
xor XOR2 (N1845, N1842, N179);
or OR4 (N1846, N1844, N1267, N176, N570);
nor NOR3 (N1847, N1835, N377, N1461);
or OR2 (N1848, N1847, N457);
nand NAND4 (N1849, N1845, N490, N354, N1093);
and AND4 (N1850, N1816, N254, N600, N1600);
buf BUF1 (N1851, N1849);
nand NAND2 (N1852, N1850, N126);
nor NOR4 (N1853, N1836, N985, N366, N1362);
xor XOR2 (N1854, N1851, N331);
and AND2 (N1855, N1846, N559);
and AND4 (N1856, N1855, N1269, N258, N643);
nor NOR2 (N1857, N1848, N1503);
not NOT1 (N1858, N1857);
nor NOR3 (N1859, N1853, N1472, N772);
xor XOR2 (N1860, N1858, N1459);
or OR4 (N1861, N1852, N24, N1434, N1365);
or OR2 (N1862, N1833, N443);
and AND2 (N1863, N1837, N293);
and AND2 (N1864, N1843, N109);
and AND4 (N1865, N1860, N804, N1259, N1505);
not NOT1 (N1866, N1856);
buf BUF1 (N1867, N1864);
nand NAND2 (N1868, N1830, N1814);
not NOT1 (N1869, N1861);
xor XOR2 (N1870, N1859, N373);
and AND4 (N1871, N1862, N948, N276, N1750);
nor NOR2 (N1872, N1869, N35);
xor XOR2 (N1873, N1867, N54);
and AND2 (N1874, N1870, N332);
or OR2 (N1875, N1872, N378);
or OR4 (N1876, N1874, N1861, N734, N1385);
or OR3 (N1877, N1871, N549, N1004);
xor XOR2 (N1878, N1873, N1540);
nand NAND4 (N1879, N1878, N1065, N561, N1104);
not NOT1 (N1880, N1854);
buf BUF1 (N1881, N1863);
buf BUF1 (N1882, N1875);
nor NOR2 (N1883, N1865, N625);
buf BUF1 (N1884, N1876);
and AND4 (N1885, N1883, N1696, N350, N1473);
nor NOR3 (N1886, N1877, N1111, N1723);
and AND3 (N1887, N1881, N77, N1719);
or OR2 (N1888, N1880, N1107);
or OR3 (N1889, N1887, N1519, N1795);
or OR3 (N1890, N1879, N644, N516);
xor XOR2 (N1891, N1888, N1253);
nor NOR4 (N1892, N1890, N491, N845, N336);
nor NOR3 (N1893, N1868, N692, N997);
nor NOR3 (N1894, N1891, N1747, N1280);
nand NAND4 (N1895, N1892, N1204, N601, N504);
nor NOR2 (N1896, N1832, N9);
and AND3 (N1897, N1889, N229, N1684);
buf BUF1 (N1898, N1895);
not NOT1 (N1899, N1866);
nand NAND2 (N1900, N1894, N203);
buf BUF1 (N1901, N1882);
and AND2 (N1902, N1898, N1503);
buf BUF1 (N1903, N1886);
nor NOR4 (N1904, N1903, N1797, N1697, N119);
and AND4 (N1905, N1900, N1505, N1642, N1780);
nor NOR3 (N1906, N1901, N1710, N1881);
nand NAND2 (N1907, N1896, N920);
nor NOR3 (N1908, N1893, N178, N1510);
xor XOR2 (N1909, N1907, N463);
not NOT1 (N1910, N1885);
nand NAND3 (N1911, N1902, N934, N1879);
or OR3 (N1912, N1905, N1709, N1699);
nor NOR4 (N1913, N1897, N182, N220, N423);
and AND4 (N1914, N1884, N221, N1144, N1804);
nand NAND3 (N1915, N1911, N1450, N868);
buf BUF1 (N1916, N1899);
buf BUF1 (N1917, N1914);
buf BUF1 (N1918, N1915);
not NOT1 (N1919, N1913);
and AND2 (N1920, N1917, N1859);
or OR2 (N1921, N1906, N1213);
or OR4 (N1922, N1910, N860, N1546, N889);
xor XOR2 (N1923, N1909, N153);
not NOT1 (N1924, N1904);
nand NAND3 (N1925, N1919, N187, N1621);
xor XOR2 (N1926, N1922, N1164);
buf BUF1 (N1927, N1920);
not NOT1 (N1928, N1912);
and AND4 (N1929, N1926, N721, N652, N1748);
nand NAND2 (N1930, N1927, N187);
not NOT1 (N1931, N1908);
not NOT1 (N1932, N1929);
nand NAND2 (N1933, N1928, N1592);
and AND2 (N1934, N1924, N1445);
nand NAND3 (N1935, N1934, N869, N164);
nand NAND3 (N1936, N1918, N1437, N635);
nor NOR4 (N1937, N1933, N713, N1809, N1441);
or OR4 (N1938, N1936, N1008, N1422, N194);
nor NOR4 (N1939, N1930, N623, N230, N902);
not NOT1 (N1940, N1938);
nor NOR2 (N1941, N1916, N1476);
not NOT1 (N1942, N1931);
nand NAND2 (N1943, N1941, N1477);
nand NAND4 (N1944, N1932, N1784, N886, N1326);
xor XOR2 (N1945, N1923, N104);
buf BUF1 (N1946, N1944);
xor XOR2 (N1947, N1925, N635);
xor XOR2 (N1948, N1942, N394);
xor XOR2 (N1949, N1935, N440);
not NOT1 (N1950, N1940);
buf BUF1 (N1951, N1945);
and AND4 (N1952, N1937, N424, N1360, N1531);
not NOT1 (N1953, N1943);
nand NAND3 (N1954, N1951, N303, N1628);
xor XOR2 (N1955, N1954, N644);
xor XOR2 (N1956, N1953, N962);
buf BUF1 (N1957, N1949);
not NOT1 (N1958, N1956);
not NOT1 (N1959, N1921);
nand NAND4 (N1960, N1957, N781, N1212, N297);
or OR4 (N1961, N1939, N125, N161, N1159);
and AND3 (N1962, N1960, N570, N1421);
nor NOR4 (N1963, N1952, N1673, N1598, N436);
and AND3 (N1964, N1961, N226, N1133);
buf BUF1 (N1965, N1963);
buf BUF1 (N1966, N1948);
nand NAND4 (N1967, N1959, N1097, N750, N1386);
nand NAND3 (N1968, N1965, N473, N1479);
nand NAND4 (N1969, N1967, N1967, N1019, N1340);
nand NAND2 (N1970, N1955, N1277);
or OR4 (N1971, N1962, N1323, N1803, N470);
or OR4 (N1972, N1950, N562, N565, N1435);
or OR4 (N1973, N1966, N1417, N1798, N1771);
xor XOR2 (N1974, N1964, N80);
xor XOR2 (N1975, N1968, N158);
nand NAND3 (N1976, N1970, N1172, N281);
not NOT1 (N1977, N1958);
buf BUF1 (N1978, N1971);
nor NOR4 (N1979, N1947, N1216, N881, N1021);
or OR2 (N1980, N1977, N809);
buf BUF1 (N1981, N1980);
buf BUF1 (N1982, N1981);
xor XOR2 (N1983, N1982, N674);
not NOT1 (N1984, N1979);
or OR2 (N1985, N1974, N220);
not NOT1 (N1986, N1976);
nand NAND4 (N1987, N1975, N1929, N461, N403);
or OR2 (N1988, N1973, N620);
or OR2 (N1989, N1985, N1988);
nor NOR3 (N1990, N1372, N292, N1402);
or OR2 (N1991, N1984, N269);
nand NAND3 (N1992, N1969, N1751, N1681);
and AND2 (N1993, N1990, N1642);
buf BUF1 (N1994, N1993);
xor XOR2 (N1995, N1983, N1744);
and AND4 (N1996, N1992, N1652, N1650, N1003);
not NOT1 (N1997, N1994);
buf BUF1 (N1998, N1997);
not NOT1 (N1999, N1986);
buf BUF1 (N2000, N1972);
xor XOR2 (N2001, N1995, N1220);
xor XOR2 (N2002, N1989, N25);
buf BUF1 (N2003, N2002);
and AND3 (N2004, N2003, N1228, N1787);
or OR3 (N2005, N2004, N1316, N897);
not NOT1 (N2006, N1978);
buf BUF1 (N2007, N1946);
or OR3 (N2008, N2001, N406, N1020);
nand NAND2 (N2009, N1987, N299);
nor NOR4 (N2010, N1998, N1136, N1561, N1671);
and AND3 (N2011, N2008, N354, N502);
not NOT1 (N2012, N2010);
buf BUF1 (N2013, N2000);
nor NOR2 (N2014, N2012, N933);
xor XOR2 (N2015, N2014, N66);
or OR2 (N2016, N1996, N1425);
not NOT1 (N2017, N2005);
and AND3 (N2018, N2017, N751, N543);
or OR4 (N2019, N2011, N792, N1178, N432);
buf BUF1 (N2020, N1991);
buf BUF1 (N2021, N2013);
xor XOR2 (N2022, N2016, N637);
buf BUF1 (N2023, N2006);
nand NAND3 (N2024, N2023, N1754, N892);
nor NOR4 (N2025, N2022, N244, N1461, N1940);
nor NOR2 (N2026, N2021, N1356);
not NOT1 (N2027, N2009);
or OR3 (N2028, N2018, N1527, N1994);
buf BUF1 (N2029, N2020);
and AND2 (N2030, N2028, N1451);
xor XOR2 (N2031, N2027, N1328);
nand NAND2 (N2032, N2019, N1900);
buf BUF1 (N2033, N2030);
not NOT1 (N2034, N2024);
and AND2 (N2035, N2031, N1964);
not NOT1 (N2036, N2029);
and AND2 (N2037, N1999, N1700);
nor NOR3 (N2038, N2015, N145, N1429);
nand NAND4 (N2039, N2037, N1832, N342, N1511);
not NOT1 (N2040, N2033);
or OR3 (N2041, N2036, N1763, N436);
or OR4 (N2042, N2038, N1151, N612, N395);
nand NAND4 (N2043, N2035, N1156, N141, N1354);
buf BUF1 (N2044, N2025);
and AND4 (N2045, N2041, N1713, N379, N268);
not NOT1 (N2046, N2040);
xor XOR2 (N2047, N2007, N1125);
nor NOR3 (N2048, N2043, N372, N1277);
xor XOR2 (N2049, N2032, N1876);
and AND3 (N2050, N2047, N123, N890);
buf BUF1 (N2051, N2042);
buf BUF1 (N2052, N2049);
xor XOR2 (N2053, N2045, N1268);
nor NOR4 (N2054, N2048, N1469, N948, N1968);
nor NOR3 (N2055, N2054, N1604, N1729);
nand NAND4 (N2056, N2052, N721, N950, N1197);
buf BUF1 (N2057, N2050);
xor XOR2 (N2058, N2055, N1800);
nand NAND4 (N2059, N2051, N1181, N341, N84);
nor NOR4 (N2060, N2059, N686, N291, N1217);
not NOT1 (N2061, N2060);
nor NOR4 (N2062, N2057, N139, N2001, N604);
nor NOR3 (N2063, N2056, N335, N971);
buf BUF1 (N2064, N2026);
nand NAND3 (N2065, N2063, N1481, N280);
nand NAND4 (N2066, N2044, N1974, N1123, N811);
xor XOR2 (N2067, N2058, N1666);
not NOT1 (N2068, N2067);
nor NOR2 (N2069, N2066, N1087);
nand NAND2 (N2070, N2069, N422);
not NOT1 (N2071, N2065);
nor NOR4 (N2072, N2061, N438, N1185, N1841);
buf BUF1 (N2073, N2046);
nand NAND3 (N2074, N2068, N1736, N577);
not NOT1 (N2075, N2034);
and AND2 (N2076, N2064, N662);
or OR4 (N2077, N2039, N1802, N1583, N952);
not NOT1 (N2078, N2076);
nand NAND3 (N2079, N2074, N1512, N1740);
and AND4 (N2080, N2073, N1375, N1305, N1963);
not NOT1 (N2081, N2053);
nor NOR3 (N2082, N2081, N1431, N292);
and AND3 (N2083, N2080, N207, N377);
buf BUF1 (N2084, N2078);
not NOT1 (N2085, N2071);
not NOT1 (N2086, N2079);
nor NOR2 (N2087, N2070, N338);
or OR3 (N2088, N2062, N424, N1265);
not NOT1 (N2089, N2085);
not NOT1 (N2090, N2083);
nor NOR3 (N2091, N2072, N734, N512);
nand NAND2 (N2092, N2089, N2041);
nand NAND3 (N2093, N2086, N623, N234);
nand NAND4 (N2094, N2092, N1249, N6, N436);
xor XOR2 (N2095, N2091, N1032);
buf BUF1 (N2096, N2093);
nand NAND4 (N2097, N2077, N391, N1783, N1955);
or OR3 (N2098, N2090, N1018, N109);
nand NAND4 (N2099, N2087, N1072, N334, N1090);
not NOT1 (N2100, N2082);
or OR3 (N2101, N2100, N386, N160);
not NOT1 (N2102, N2084);
buf BUF1 (N2103, N2102);
nor NOR4 (N2104, N2075, N360, N17, N1571);
nand NAND4 (N2105, N2097, N631, N782, N1319);
nand NAND2 (N2106, N2104, N636);
not NOT1 (N2107, N2105);
nor NOR2 (N2108, N2088, N1260);
buf BUF1 (N2109, N2103);
xor XOR2 (N2110, N2095, N1231);
nand NAND4 (N2111, N2108, N832, N1345, N801);
not NOT1 (N2112, N2110);
xor XOR2 (N2113, N2098, N1682);
and AND4 (N2114, N2109, N627, N706, N747);
not NOT1 (N2115, N2113);
buf BUF1 (N2116, N2096);
and AND2 (N2117, N2112, N1079);
nand NAND2 (N2118, N2094, N17);
xor XOR2 (N2119, N2118, N1751);
or OR3 (N2120, N2107, N1864, N195);
nand NAND3 (N2121, N2106, N1646, N1516);
buf BUF1 (N2122, N2099);
or OR4 (N2123, N2120, N978, N1300, N1967);
and AND2 (N2124, N2101, N786);
and AND2 (N2125, N2111, N1147);
nor NOR3 (N2126, N2124, N1580, N835);
nand NAND4 (N2127, N2116, N1101, N2122, N1778);
xor XOR2 (N2128, N434, N1117);
or OR2 (N2129, N2127, N1099);
not NOT1 (N2130, N2129);
nand NAND4 (N2131, N2130, N1927, N2099, N1442);
or OR4 (N2132, N2123, N1475, N843, N974);
nand NAND2 (N2133, N2128, N1930);
nand NAND3 (N2134, N2132, N85, N62);
or OR2 (N2135, N2125, N1543);
nand NAND3 (N2136, N2131, N1114, N719);
xor XOR2 (N2137, N2126, N1940);
nor NOR4 (N2138, N2115, N63, N898, N1716);
not NOT1 (N2139, N2121);
not NOT1 (N2140, N2136);
or OR2 (N2141, N2138, N1614);
nand NAND4 (N2142, N2137, N639, N36, N747);
buf BUF1 (N2143, N2119);
or OR3 (N2144, N2133, N1629, N1954);
and AND2 (N2145, N2140, N1035);
xor XOR2 (N2146, N2143, N614);
buf BUF1 (N2147, N2134);
nor NOR4 (N2148, N2114, N1260, N1519, N493);
and AND2 (N2149, N2135, N641);
nor NOR4 (N2150, N2148, N1183, N1740, N924);
nor NOR3 (N2151, N2141, N1167, N1386);
or OR4 (N2152, N2139, N1925, N1062, N1318);
and AND2 (N2153, N2144, N919);
nor NOR2 (N2154, N2142, N1339);
xor XOR2 (N2155, N2154, N80);
buf BUF1 (N2156, N2151);
nand NAND4 (N2157, N2150, N2099, N1327, N1973);
and AND4 (N2158, N2156, N559, N1931, N778);
xor XOR2 (N2159, N2147, N1804);
not NOT1 (N2160, N2159);
xor XOR2 (N2161, N2146, N1838);
nand NAND2 (N2162, N2152, N1358);
or OR2 (N2163, N2162, N965);
nand NAND4 (N2164, N2163, N1130, N1071, N2072);
nand NAND4 (N2165, N2117, N2100, N542, N1499);
and AND4 (N2166, N2149, N715, N1617, N304);
xor XOR2 (N2167, N2164, N892);
and AND3 (N2168, N2166, N312, N1636);
buf BUF1 (N2169, N2145);
nand NAND2 (N2170, N2157, N939);
buf BUF1 (N2171, N2168);
buf BUF1 (N2172, N2158);
nand NAND2 (N2173, N2165, N1715);
nand NAND3 (N2174, N2172, N2167, N1528);
or OR2 (N2175, N1756, N1700);
nor NOR3 (N2176, N2161, N1154, N1394);
buf BUF1 (N2177, N2153);
or OR4 (N2178, N2155, N124, N355, N1467);
nand NAND4 (N2179, N2169, N802, N962, N1924);
or OR3 (N2180, N2160, N718, N900);
or OR4 (N2181, N2173, N2157, N440, N355);
and AND3 (N2182, N2181, N2033, N10);
not NOT1 (N2183, N2179);
nand NAND4 (N2184, N2176, N1154, N94, N1550);
and AND2 (N2185, N2171, N429);
or OR2 (N2186, N2183, N23);
nand NAND3 (N2187, N2182, N1390, N848);
nand NAND2 (N2188, N2187, N979);
or OR4 (N2189, N2174, N657, N1330, N1766);
nor NOR3 (N2190, N2186, N27, N787);
not NOT1 (N2191, N2177);
nor NOR4 (N2192, N2189, N2073, N406, N1521);
nand NAND4 (N2193, N2180, N541, N1950, N2136);
buf BUF1 (N2194, N2185);
buf BUF1 (N2195, N2194);
nor NOR2 (N2196, N2170, N1738);
and AND4 (N2197, N2196, N2139, N468, N238);
nor NOR3 (N2198, N2197, N2183, N583);
and AND2 (N2199, N2191, N362);
buf BUF1 (N2200, N2198);
xor XOR2 (N2201, N2184, N798);
nor NOR3 (N2202, N2201, N440, N214);
nand NAND3 (N2203, N2188, N2116, N696);
nand NAND3 (N2204, N2192, N1825, N2107);
and AND4 (N2205, N2178, N1381, N1032, N929);
nand NAND2 (N2206, N2202, N831);
and AND4 (N2207, N2199, N54, N850, N69);
or OR4 (N2208, N2204, N1125, N1337, N665);
not NOT1 (N2209, N2206);
xor XOR2 (N2210, N2207, N1401);
nor NOR4 (N2211, N2203, N2018, N2065, N829);
nand NAND2 (N2212, N2209, N754);
xor XOR2 (N2213, N2211, N920);
nand NAND3 (N2214, N2210, N221, N2112);
buf BUF1 (N2215, N2205);
xor XOR2 (N2216, N2195, N1550);
xor XOR2 (N2217, N2215, N784);
nor NOR3 (N2218, N2175, N1006, N2078);
or OR4 (N2219, N2190, N754, N42, N1957);
or OR4 (N2220, N2213, N936, N844, N611);
and AND2 (N2221, N2212, N1214);
buf BUF1 (N2222, N2193);
xor XOR2 (N2223, N2208, N1511);
nand NAND2 (N2224, N2217, N408);
nand NAND4 (N2225, N2224, N2188, N1484, N372);
nor NOR4 (N2226, N2222, N2138, N380, N1874);
nand NAND2 (N2227, N2214, N598);
nor NOR3 (N2228, N2225, N1996, N2097);
or OR4 (N2229, N2220, N1403, N1382, N699);
nand NAND2 (N2230, N2216, N1862);
buf BUF1 (N2231, N2223);
xor XOR2 (N2232, N2218, N1546);
nand NAND3 (N2233, N2221, N1189, N1384);
xor XOR2 (N2234, N2219, N1166);
nor NOR4 (N2235, N2227, N1886, N1171, N441);
not NOT1 (N2236, N2231);
and AND2 (N2237, N2233, N2121);
nand NAND3 (N2238, N2237, N357, N2181);
not NOT1 (N2239, N2238);
buf BUF1 (N2240, N2200);
buf BUF1 (N2241, N2226);
nand NAND4 (N2242, N2236, N1814, N642, N97);
and AND3 (N2243, N2242, N2062, N2183);
nor NOR4 (N2244, N2235, N1458, N1463, N1203);
nor NOR4 (N2245, N2234, N749, N166, N811);
nor NOR3 (N2246, N2232, N1246, N1091);
buf BUF1 (N2247, N2228);
or OR2 (N2248, N2239, N792);
and AND4 (N2249, N2246, N335, N34, N1756);
nor NOR2 (N2250, N2245, N1631);
nand NAND3 (N2251, N2250, N965, N500);
nand NAND3 (N2252, N2229, N761, N2040);
or OR2 (N2253, N2240, N2091);
nand NAND3 (N2254, N2249, N114, N1161);
nor NOR2 (N2255, N2243, N1760);
or OR4 (N2256, N2230, N766, N357, N1231);
or OR2 (N2257, N2254, N1921);
nand NAND4 (N2258, N2247, N2257, N1863, N1321);
or OR3 (N2259, N1745, N470, N87);
nand NAND4 (N2260, N2253, N1121, N1492, N1422);
buf BUF1 (N2261, N2244);
xor XOR2 (N2262, N2252, N895);
buf BUF1 (N2263, N2255);
buf BUF1 (N2264, N2261);
nand NAND3 (N2265, N2251, N1388, N252);
nand NAND4 (N2266, N2260, N1601, N968, N1423);
and AND2 (N2267, N2248, N1090);
nand NAND3 (N2268, N2265, N557, N1016);
buf BUF1 (N2269, N2263);
not NOT1 (N2270, N2268);
nor NOR3 (N2271, N2270, N380, N2173);
not NOT1 (N2272, N2269);
buf BUF1 (N2273, N2259);
buf BUF1 (N2274, N2272);
nor NOR4 (N2275, N2241, N481, N1621, N502);
xor XOR2 (N2276, N2273, N2151);
nor NOR2 (N2277, N2275, N2076);
nor NOR3 (N2278, N2256, N277, N1729);
nand NAND4 (N2279, N2274, N90, N2241, N1086);
and AND4 (N2280, N2271, N1272, N1951, N181);
nor NOR2 (N2281, N2278, N159);
not NOT1 (N2282, N2276);
buf BUF1 (N2283, N2281);
or OR2 (N2284, N2264, N480);
or OR4 (N2285, N2283, N1699, N2057, N1618);
nor NOR2 (N2286, N2267, N239);
and AND2 (N2287, N2286, N261);
nand NAND4 (N2288, N2285, N614, N1990, N1202);
not NOT1 (N2289, N2284);
not NOT1 (N2290, N2279);
nand NAND4 (N2291, N2277, N625, N1382, N1103);
and AND2 (N2292, N2258, N1038);
xor XOR2 (N2293, N2280, N887);
nor NOR2 (N2294, N2289, N39);
and AND3 (N2295, N2262, N1840, N1412);
xor XOR2 (N2296, N2282, N961);
xor XOR2 (N2297, N2290, N1855);
and AND3 (N2298, N2288, N2149, N628);
not NOT1 (N2299, N2297);
xor XOR2 (N2300, N2292, N1854);
xor XOR2 (N2301, N2291, N1491);
xor XOR2 (N2302, N2298, N608);
xor XOR2 (N2303, N2294, N560);
buf BUF1 (N2304, N2266);
xor XOR2 (N2305, N2304, N626);
not NOT1 (N2306, N2300);
nor NOR2 (N2307, N2305, N1739);
or OR3 (N2308, N2287, N45, N2271);
buf BUF1 (N2309, N2307);
nand NAND4 (N2310, N2296, N389, N1234, N1869);
xor XOR2 (N2311, N2306, N774);
nor NOR3 (N2312, N2302, N1025, N945);
nor NOR4 (N2313, N2301, N1003, N1121, N1205);
xor XOR2 (N2314, N2293, N1766);
not NOT1 (N2315, N2303);
xor XOR2 (N2316, N2309, N2184);
nand NAND4 (N2317, N2311, N2177, N2072, N2249);
or OR3 (N2318, N2308, N1224, N2127);
nand NAND4 (N2319, N2313, N1932, N134, N1034);
and AND4 (N2320, N2299, N256, N629, N1072);
buf BUF1 (N2321, N2318);
and AND2 (N2322, N2295, N2220);
not NOT1 (N2323, N2312);
nand NAND2 (N2324, N2321, N689);
and AND3 (N2325, N2315, N1830, N254);
and AND2 (N2326, N2314, N1088);
and AND4 (N2327, N2319, N1278, N432, N1829);
not NOT1 (N2328, N2323);
and AND3 (N2329, N2326, N1673, N686);
not NOT1 (N2330, N2317);
nor NOR4 (N2331, N2330, N436, N2330, N1182);
and AND3 (N2332, N2324, N422, N1584);
nand NAND3 (N2333, N2310, N1047, N2131);
buf BUF1 (N2334, N2325);
buf BUF1 (N2335, N2329);
and AND3 (N2336, N2331, N337, N1118);
nand NAND2 (N2337, N2316, N1975);
nor NOR2 (N2338, N2322, N1574);
not NOT1 (N2339, N2327);
and AND3 (N2340, N2328, N2259, N1767);
nand NAND3 (N2341, N2320, N713, N1224);
xor XOR2 (N2342, N2334, N2117);
nand NAND3 (N2343, N2333, N952, N839);
and AND3 (N2344, N2342, N1053, N694);
and AND4 (N2345, N2343, N1486, N982, N476);
buf BUF1 (N2346, N2338);
not NOT1 (N2347, N2335);
and AND4 (N2348, N2332, N312, N1939, N1126);
xor XOR2 (N2349, N2340, N598);
nor NOR2 (N2350, N2337, N2112);
xor XOR2 (N2351, N2336, N292);
not NOT1 (N2352, N2345);
nor NOR2 (N2353, N2341, N2175);
buf BUF1 (N2354, N2350);
buf BUF1 (N2355, N2351);
buf BUF1 (N2356, N2347);
nor NOR3 (N2357, N2353, N1616, N2066);
buf BUF1 (N2358, N2357);
and AND3 (N2359, N2339, N2347, N1747);
nor NOR3 (N2360, N2355, N1358, N522);
xor XOR2 (N2361, N2359, N1379);
not NOT1 (N2362, N2344);
nor NOR2 (N2363, N2354, N230);
nor NOR3 (N2364, N2349, N907, N1812);
nand NAND2 (N2365, N2358, N746);
and AND4 (N2366, N2363, N283, N480, N1213);
buf BUF1 (N2367, N2362);
or OR4 (N2368, N2346, N2220, N393, N755);
or OR2 (N2369, N2348, N995);
buf BUF1 (N2370, N2364);
buf BUF1 (N2371, N2356);
and AND3 (N2372, N2361, N1568, N1570);
not NOT1 (N2373, N2371);
nor NOR4 (N2374, N2360, N40, N724, N656);
and AND2 (N2375, N2367, N1873);
and AND4 (N2376, N2366, N1518, N864, N818);
not NOT1 (N2377, N2374);
or OR2 (N2378, N2375, N1987);
and AND3 (N2379, N2368, N2015, N422);
xor XOR2 (N2380, N2372, N852);
and AND4 (N2381, N2376, N808, N1060, N1575);
or OR4 (N2382, N2377, N541, N1436, N99);
or OR4 (N2383, N2381, N107, N824, N2321);
and AND4 (N2384, N2370, N802, N1468, N268);
and AND2 (N2385, N2380, N1067);
or OR2 (N2386, N2383, N606);
and AND3 (N2387, N2378, N1847, N285);
xor XOR2 (N2388, N2386, N1381);
or OR2 (N2389, N2387, N1189);
and AND2 (N2390, N2352, N1455);
nand NAND4 (N2391, N2384, N1843, N1640, N1604);
or OR2 (N2392, N2369, N1038);
and AND3 (N2393, N2388, N1268, N465);
or OR3 (N2394, N2379, N802, N2274);
xor XOR2 (N2395, N2373, N817);
and AND3 (N2396, N2393, N239, N1284);
buf BUF1 (N2397, N2365);
not NOT1 (N2398, N2391);
buf BUF1 (N2399, N2395);
nand NAND4 (N2400, N2399, N926, N1132, N507);
not NOT1 (N2401, N2397);
xor XOR2 (N2402, N2401, N1817);
not NOT1 (N2403, N2389);
xor XOR2 (N2404, N2392, N2272);
xor XOR2 (N2405, N2403, N449);
buf BUF1 (N2406, N2396);
not NOT1 (N2407, N2405);
and AND4 (N2408, N2394, N339, N1534, N1560);
nor NOR2 (N2409, N2400, N934);
not NOT1 (N2410, N2382);
not NOT1 (N2411, N2398);
nor NOR2 (N2412, N2411, N2073);
and AND2 (N2413, N2390, N541);
nand NAND3 (N2414, N2385, N218, N1827);
not NOT1 (N2415, N2407);
nor NOR4 (N2416, N2415, N162, N1845, N2164);
buf BUF1 (N2417, N2404);
not NOT1 (N2418, N2409);
and AND3 (N2419, N2414, N711, N1688);
not NOT1 (N2420, N2418);
buf BUF1 (N2421, N2408);
or OR3 (N2422, N2421, N1969, N2127);
buf BUF1 (N2423, N2406);
or OR2 (N2424, N2416, N1011);
xor XOR2 (N2425, N2412, N1489);
nor NOR3 (N2426, N2424, N718, N2026);
nor NOR2 (N2427, N2402, N788);
xor XOR2 (N2428, N2419, N1969);
and AND3 (N2429, N2427, N1872, N140);
buf BUF1 (N2430, N2426);
xor XOR2 (N2431, N2422, N2352);
buf BUF1 (N2432, N2430);
nand NAND2 (N2433, N2420, N227);
and AND2 (N2434, N2433, N432);
or OR2 (N2435, N2432, N1107);
and AND3 (N2436, N2435, N1999, N833);
buf BUF1 (N2437, N2410);
and AND2 (N2438, N2431, N1339);
not NOT1 (N2439, N2428);
not NOT1 (N2440, N2438);
nor NOR3 (N2441, N2425, N1228, N930);
nand NAND3 (N2442, N2434, N1493, N839);
or OR4 (N2443, N2439, N148, N1746, N952);
not NOT1 (N2444, N2436);
or OR3 (N2445, N2413, N1101, N261);
nor NOR3 (N2446, N2445, N532, N475);
or OR4 (N2447, N2437, N1906, N2268, N295);
xor XOR2 (N2448, N2447, N555);
and AND3 (N2449, N2441, N2072, N297);
nor NOR3 (N2450, N2442, N2025, N1872);
buf BUF1 (N2451, N2423);
xor XOR2 (N2452, N2417, N1688);
nor NOR2 (N2453, N2452, N294);
buf BUF1 (N2454, N2449);
and AND2 (N2455, N2444, N173);
buf BUF1 (N2456, N2453);
and AND2 (N2457, N2456, N1416);
or OR2 (N2458, N2455, N240);
not NOT1 (N2459, N2457);
xor XOR2 (N2460, N2451, N950);
not NOT1 (N2461, N2443);
not NOT1 (N2462, N2454);
nand NAND4 (N2463, N2450, N1938, N1959, N373);
not NOT1 (N2464, N2448);
and AND2 (N2465, N2463, N449);
and AND3 (N2466, N2446, N606, N1031);
nand NAND3 (N2467, N2464, N1615, N2156);
buf BUF1 (N2468, N2458);
xor XOR2 (N2469, N2465, N472);
buf BUF1 (N2470, N2461);
nor NOR3 (N2471, N2467, N1442, N1726);
nor NOR3 (N2472, N2470, N1316, N194);
or OR2 (N2473, N2429, N1075);
buf BUF1 (N2474, N2468);
not NOT1 (N2475, N2472);
not NOT1 (N2476, N2471);
not NOT1 (N2477, N2474);
and AND2 (N2478, N2476, N1671);
or OR2 (N2479, N2478, N1959);
not NOT1 (N2480, N2469);
and AND2 (N2481, N2466, N883);
not NOT1 (N2482, N2440);
and AND2 (N2483, N2459, N827);
nor NOR4 (N2484, N2482, N2202, N575, N21);
nand NAND2 (N2485, N2460, N1394);
nand NAND3 (N2486, N2477, N2419, N2105);
and AND3 (N2487, N2475, N775, N1394);
xor XOR2 (N2488, N2483, N954);
or OR4 (N2489, N2473, N2000, N2268, N646);
nand NAND2 (N2490, N2487, N405);
xor XOR2 (N2491, N2490, N906);
nand NAND2 (N2492, N2481, N824);
nand NAND2 (N2493, N2485, N1256);
or OR3 (N2494, N2489, N342, N476);
buf BUF1 (N2495, N2491);
or OR3 (N2496, N2479, N2266, N1417);
not NOT1 (N2497, N2488);
and AND2 (N2498, N2492, N31);
nor NOR3 (N2499, N2496, N1224, N1092);
nand NAND3 (N2500, N2499, N832, N427);
and AND2 (N2501, N2480, N2133);
nor NOR3 (N2502, N2495, N896, N223);
and AND2 (N2503, N2502, N818);
and AND3 (N2504, N2493, N222, N1828);
or OR3 (N2505, N2500, N1550, N2191);
or OR4 (N2506, N2503, N729, N702, N2296);
buf BUF1 (N2507, N2486);
xor XOR2 (N2508, N2497, N1892);
or OR3 (N2509, N2484, N575, N1560);
nand NAND4 (N2510, N2498, N1932, N740, N1188);
not NOT1 (N2511, N2507);
or OR2 (N2512, N2508, N1804);
xor XOR2 (N2513, N2506, N1522);
not NOT1 (N2514, N2504);
nor NOR3 (N2515, N2514, N769, N2312);
not NOT1 (N2516, N2512);
and AND3 (N2517, N2462, N1201, N2331);
nor NOR4 (N2518, N2516, N639, N684, N1509);
and AND3 (N2519, N2494, N669, N1701);
nand NAND4 (N2520, N2519, N317, N1434, N2273);
nor NOR4 (N2521, N2515, N918, N1205, N1480);
buf BUF1 (N2522, N2520);
xor XOR2 (N2523, N2521, N1168);
nor NOR3 (N2524, N2522, N2305, N1632);
not NOT1 (N2525, N2518);
xor XOR2 (N2526, N2525, N552);
xor XOR2 (N2527, N2501, N1106);
nor NOR3 (N2528, N2511, N1248, N1271);
nand NAND3 (N2529, N2523, N2187, N1824);
or OR2 (N2530, N2528, N1457);
and AND3 (N2531, N2529, N681, N2353);
buf BUF1 (N2532, N2524);
and AND2 (N2533, N2517, N467);
buf BUF1 (N2534, N2530);
xor XOR2 (N2535, N2531, N1677);
nand NAND4 (N2536, N2505, N870, N649, N1912);
nor NOR3 (N2537, N2534, N715, N1941);
and AND3 (N2538, N2513, N1124, N1203);
not NOT1 (N2539, N2526);
not NOT1 (N2540, N2509);
and AND4 (N2541, N2535, N1673, N1493, N831);
buf BUF1 (N2542, N2533);
buf BUF1 (N2543, N2536);
nand NAND4 (N2544, N2527, N1539, N2460, N1429);
nor NOR2 (N2545, N2540, N2284);
buf BUF1 (N2546, N2543);
xor XOR2 (N2547, N2510, N1117);
nor NOR2 (N2548, N2537, N490);
nor NOR4 (N2549, N2541, N1908, N2386, N1812);
or OR4 (N2550, N2548, N989, N1031, N2345);
or OR4 (N2551, N2549, N195, N1789, N2503);
and AND3 (N2552, N2542, N182, N797);
nor NOR4 (N2553, N2546, N1911, N784, N1387);
nand NAND4 (N2554, N2539, N1947, N1343, N2335);
xor XOR2 (N2555, N2532, N967);
buf BUF1 (N2556, N2538);
not NOT1 (N2557, N2552);
xor XOR2 (N2558, N2555, N2263);
xor XOR2 (N2559, N2547, N2256);
nand NAND4 (N2560, N2553, N2390, N619, N2238);
nor NOR2 (N2561, N2554, N86);
nor NOR3 (N2562, N2544, N899, N1075);
nand NAND2 (N2563, N2562, N1263);
or OR2 (N2564, N2561, N118);
xor XOR2 (N2565, N2557, N998);
nand NAND3 (N2566, N2558, N1831, N925);
nand NAND2 (N2567, N2559, N2420);
and AND3 (N2568, N2560, N1460, N358);
not NOT1 (N2569, N2563);
nand NAND4 (N2570, N2565, N959, N1343, N1870);
nor NOR3 (N2571, N2545, N1490, N5);
nor NOR4 (N2572, N2570, N1249, N645, N749);
not NOT1 (N2573, N2568);
nor NOR2 (N2574, N2573, N2336);
xor XOR2 (N2575, N2569, N1901);
and AND3 (N2576, N2551, N617, N2280);
buf BUF1 (N2577, N2566);
xor XOR2 (N2578, N2574, N1164);
not NOT1 (N2579, N2571);
not NOT1 (N2580, N2564);
or OR2 (N2581, N2572, N1701);
buf BUF1 (N2582, N2576);
and AND3 (N2583, N2579, N654, N295);
buf BUF1 (N2584, N2577);
or OR2 (N2585, N2583, N2563);
buf BUF1 (N2586, N2556);
xor XOR2 (N2587, N2581, N1249);
not NOT1 (N2588, N2584);
or OR2 (N2589, N2580, N2140);
nor NOR4 (N2590, N2585, N2381, N2355, N2001);
nor NOR3 (N2591, N2586, N506, N1403);
buf BUF1 (N2592, N2578);
nand NAND4 (N2593, N2587, N1812, N267, N765);
nand NAND2 (N2594, N2575, N1371);
xor XOR2 (N2595, N2591, N2102);
or OR3 (N2596, N2550, N1993, N1702);
not NOT1 (N2597, N2582);
nor NOR3 (N2598, N2595, N1236, N1038);
buf BUF1 (N2599, N2594);
buf BUF1 (N2600, N2592);
nor NOR3 (N2601, N2590, N1378, N1696);
and AND3 (N2602, N2593, N368, N2435);
or OR4 (N2603, N2589, N1750, N1708, N379);
not NOT1 (N2604, N2598);
nor NOR3 (N2605, N2596, N1343, N1248);
nor NOR4 (N2606, N2600, N744, N1720, N1037);
nand NAND3 (N2607, N2597, N481, N1490);
nand NAND3 (N2608, N2605, N2316, N984);
nor NOR4 (N2609, N2602, N2107, N332, N1600);
nand NAND4 (N2610, N2609, N2189, N773, N156);
not NOT1 (N2611, N2608);
nor NOR4 (N2612, N2567, N2088, N2597, N663);
and AND4 (N2613, N2610, N2480, N1525, N1105);
nor NOR4 (N2614, N2604, N950, N924, N1430);
buf BUF1 (N2615, N2613);
and AND4 (N2616, N2599, N1884, N1210, N224);
nand NAND2 (N2617, N2614, N189);
buf BUF1 (N2618, N2601);
nor NOR3 (N2619, N2615, N2554, N2116);
nand NAND3 (N2620, N2606, N2036, N145);
nand NAND3 (N2621, N2616, N1285, N1275);
not NOT1 (N2622, N2618);
not NOT1 (N2623, N2588);
buf BUF1 (N2624, N2622);
xor XOR2 (N2625, N2620, N1349);
and AND4 (N2626, N2603, N1176, N1752, N2584);
not NOT1 (N2627, N2624);
not NOT1 (N2628, N2627);
not NOT1 (N2629, N2623);
buf BUF1 (N2630, N2617);
buf BUF1 (N2631, N2611);
nand NAND4 (N2632, N2630, N1396, N844, N2542);
and AND3 (N2633, N2621, N1574, N1451);
nand NAND2 (N2634, N2632, N1775);
not NOT1 (N2635, N2628);
xor XOR2 (N2636, N2634, N2072);
or OR4 (N2637, N2631, N149, N2359, N2140);
or OR3 (N2638, N2629, N772, N297);
xor XOR2 (N2639, N2635, N1436);
nand NAND4 (N2640, N2637, N2168, N1153, N1760);
not NOT1 (N2641, N2633);
not NOT1 (N2642, N2638);
buf BUF1 (N2643, N2642);
or OR3 (N2644, N2607, N19, N819);
nor NOR2 (N2645, N2644, N2422);
xor XOR2 (N2646, N2645, N1743);
xor XOR2 (N2647, N2626, N1646);
nand NAND4 (N2648, N2640, N309, N804, N2602);
nor NOR4 (N2649, N2625, N1779, N66, N211);
and AND4 (N2650, N2649, N1533, N2371, N2106);
nor NOR2 (N2651, N2643, N646);
not NOT1 (N2652, N2639);
and AND4 (N2653, N2646, N2055, N1719, N699);
and AND2 (N2654, N2612, N786);
xor XOR2 (N2655, N2650, N1982);
nand NAND2 (N2656, N2651, N1587);
buf BUF1 (N2657, N2619);
nor NOR3 (N2658, N2654, N2618, N620);
nor NOR3 (N2659, N2653, N2381, N2376);
and AND2 (N2660, N2636, N947);
nand NAND2 (N2661, N2648, N1305);
buf BUF1 (N2662, N2655);
and AND4 (N2663, N2656, N2464, N414, N2449);
or OR4 (N2664, N2657, N2286, N1936, N1023);
xor XOR2 (N2665, N2641, N529);
or OR4 (N2666, N2665, N2105, N2029, N113);
buf BUF1 (N2667, N2661);
nand NAND2 (N2668, N2667, N974);
and AND3 (N2669, N2647, N1981, N956);
buf BUF1 (N2670, N2660);
not NOT1 (N2671, N2666);
nor NOR4 (N2672, N2670, N552, N729, N1788);
or OR2 (N2673, N2663, N1455);
or OR3 (N2674, N2662, N2558, N1467);
nand NAND2 (N2675, N2671, N38);
nor NOR3 (N2676, N2674, N2427, N1272);
nor NOR3 (N2677, N2676, N744, N141);
buf BUF1 (N2678, N2672);
buf BUF1 (N2679, N2673);
nand NAND4 (N2680, N2652, N984, N85, N497);
xor XOR2 (N2681, N2669, N1492);
nor NOR4 (N2682, N2675, N302, N1243, N2018);
not NOT1 (N2683, N2668);
or OR4 (N2684, N2664, N1119, N1785, N2376);
not NOT1 (N2685, N2684);
buf BUF1 (N2686, N2682);
nand NAND4 (N2687, N2681, N1639, N2172, N2268);
or OR3 (N2688, N2659, N583, N2086);
xor XOR2 (N2689, N2677, N1845);
buf BUF1 (N2690, N2683);
xor XOR2 (N2691, N2658, N681);
nand NAND4 (N2692, N2679, N1349, N918, N4);
buf BUF1 (N2693, N2678);
nor NOR4 (N2694, N2680, N1126, N492, N526);
and AND3 (N2695, N2688, N1383, N1597);
buf BUF1 (N2696, N2689);
nor NOR2 (N2697, N2691, N1387);
or OR4 (N2698, N2694, N341, N738, N1646);
nand NAND2 (N2699, N2686, N2450);
nand NAND4 (N2700, N2698, N1687, N2489, N2255);
nor NOR3 (N2701, N2693, N2039, N2398);
xor XOR2 (N2702, N2701, N2200);
or OR2 (N2703, N2696, N1162);
buf BUF1 (N2704, N2697);
and AND2 (N2705, N2695, N230);
xor XOR2 (N2706, N2685, N1803);
or OR2 (N2707, N2706, N544);
and AND2 (N2708, N2705, N1011);
not NOT1 (N2709, N2687);
xor XOR2 (N2710, N2707, N2497);
and AND2 (N2711, N2710, N2382);
or OR2 (N2712, N2690, N493);
buf BUF1 (N2713, N2700);
and AND2 (N2714, N2703, N2390);
nor NOR4 (N2715, N2704, N1526, N199, N866);
not NOT1 (N2716, N2714);
or OR3 (N2717, N2716, N336, N1120);
buf BUF1 (N2718, N2717);
buf BUF1 (N2719, N2692);
nor NOR2 (N2720, N2702, N511);
nor NOR2 (N2721, N2708, N795);
buf BUF1 (N2722, N2718);
buf BUF1 (N2723, N2712);
xor XOR2 (N2724, N2713, N1694);
or OR3 (N2725, N2723, N2252, N1198);
not NOT1 (N2726, N2715);
xor XOR2 (N2727, N2699, N2498);
nor NOR3 (N2728, N2722, N1629, N2615);
buf BUF1 (N2729, N2727);
not NOT1 (N2730, N2728);
nand NAND4 (N2731, N2724, N746, N2040, N620);
buf BUF1 (N2732, N2731);
or OR3 (N2733, N2720, N1719, N2551);
nor NOR2 (N2734, N2719, N582);
nor NOR3 (N2735, N2733, N2391, N1038);
nand NAND3 (N2736, N2711, N1843, N857);
not NOT1 (N2737, N2734);
or OR2 (N2738, N2729, N2156);
or OR2 (N2739, N2709, N1154);
nand NAND2 (N2740, N2738, N1462);
nand NAND3 (N2741, N2730, N640, N2069);
xor XOR2 (N2742, N2726, N1440);
or OR4 (N2743, N2725, N1853, N130, N2647);
buf BUF1 (N2744, N2740);
nand NAND3 (N2745, N2736, N2234, N441);
and AND2 (N2746, N2745, N2437);
not NOT1 (N2747, N2721);
nor NOR2 (N2748, N2743, N369);
nor NOR4 (N2749, N2735, N2240, N1449, N1384);
not NOT1 (N2750, N2749);
nor NOR2 (N2751, N2744, N2026);
and AND4 (N2752, N2739, N1672, N2102, N2641);
and AND2 (N2753, N2752, N560);
not NOT1 (N2754, N2747);
buf BUF1 (N2755, N2754);
or OR2 (N2756, N2746, N26);
nand NAND2 (N2757, N2737, N136);
and AND3 (N2758, N2756, N421, N329);
not NOT1 (N2759, N2753);
not NOT1 (N2760, N2742);
nor NOR2 (N2761, N2748, N2101);
nand NAND3 (N2762, N2741, N2008, N1071);
nor NOR2 (N2763, N2762, N2538);
or OR2 (N2764, N2751, N2551);
not NOT1 (N2765, N2758);
or OR3 (N2766, N2759, N1831, N2503);
nor NOR2 (N2767, N2764, N1506);
or OR4 (N2768, N2750, N2523, N2232, N2526);
or OR2 (N2769, N2761, N1134);
nor NOR2 (N2770, N2760, N459);
nand NAND3 (N2771, N2769, N2029, N2454);
buf BUF1 (N2772, N2768);
nand NAND3 (N2773, N2770, N2747, N1295);
not NOT1 (N2774, N2757);
and AND4 (N2775, N2765, N138, N1309, N2629);
or OR3 (N2776, N2732, N1974, N732);
or OR3 (N2777, N2774, N692, N2258);
or OR2 (N2778, N2755, N847);
nand NAND3 (N2779, N2777, N1426, N714);
and AND2 (N2780, N2771, N1275);
buf BUF1 (N2781, N2780);
nor NOR3 (N2782, N2779, N2173, N1609);
nor NOR2 (N2783, N2763, N2241);
buf BUF1 (N2784, N2773);
buf BUF1 (N2785, N2776);
and AND3 (N2786, N2785, N1134, N1551);
nor NOR2 (N2787, N2778, N1092);
and AND2 (N2788, N2781, N2082);
not NOT1 (N2789, N2787);
buf BUF1 (N2790, N2767);
xor XOR2 (N2791, N2789, N2642);
not NOT1 (N2792, N2775);
not NOT1 (N2793, N2783);
buf BUF1 (N2794, N2786);
nand NAND3 (N2795, N2790, N596, N1316);
buf BUF1 (N2796, N2788);
xor XOR2 (N2797, N2791, N417);
xor XOR2 (N2798, N2792, N1525);
xor XOR2 (N2799, N2794, N587);
nand NAND2 (N2800, N2798, N1342);
and AND3 (N2801, N2799, N487, N1276);
nor NOR2 (N2802, N2784, N2367);
nand NAND4 (N2803, N2800, N2100, N2140, N600);
buf BUF1 (N2804, N2802);
nor NOR2 (N2805, N2796, N970);
and AND2 (N2806, N2793, N817);
buf BUF1 (N2807, N2772);
buf BUF1 (N2808, N2801);
not NOT1 (N2809, N2803);
buf BUF1 (N2810, N2804);
or OR4 (N2811, N2766, N1662, N1082, N2360);
or OR3 (N2812, N2795, N2618, N564);
not NOT1 (N2813, N2807);
buf BUF1 (N2814, N2806);
not NOT1 (N2815, N2813);
xor XOR2 (N2816, N2808, N2261);
not NOT1 (N2817, N2809);
buf BUF1 (N2818, N2817);
buf BUF1 (N2819, N2810);
nor NOR4 (N2820, N2805, N2428, N1250, N1546);
and AND2 (N2821, N2815, N116);
xor XOR2 (N2822, N2820, N371);
buf BUF1 (N2823, N2822);
nand NAND4 (N2824, N2816, N1493, N2147, N2525);
buf BUF1 (N2825, N2823);
nor NOR2 (N2826, N2818, N1215);
nor NOR2 (N2827, N2826, N411);
or OR2 (N2828, N2825, N987);
nor NOR4 (N2829, N2819, N2214, N1591, N2145);
nand NAND3 (N2830, N2782, N1221, N973);
nor NOR2 (N2831, N2829, N1823);
nor NOR4 (N2832, N2812, N77, N941, N804);
or OR4 (N2833, N2814, N2178, N1814, N3);
nand NAND4 (N2834, N2828, N2661, N66, N2798);
buf BUF1 (N2835, N2831);
nor NOR4 (N2836, N2821, N158, N909, N1746);
or OR2 (N2837, N2836, N544);
buf BUF1 (N2838, N2832);
nor NOR2 (N2839, N2811, N652);
nor NOR2 (N2840, N2839, N153);
or OR4 (N2841, N2827, N1531, N1387, N1080);
nor NOR4 (N2842, N2797, N1624, N1107, N2417);
or OR3 (N2843, N2837, N2091, N1061);
nor NOR4 (N2844, N2824, N1720, N1730, N1614);
xor XOR2 (N2845, N2841, N2560);
nand NAND4 (N2846, N2835, N1580, N189, N2600);
nand NAND2 (N2847, N2830, N272);
or OR4 (N2848, N2845, N59, N2530, N5);
nand NAND4 (N2849, N2848, N319, N1269, N813);
xor XOR2 (N2850, N2838, N598);
nor NOR2 (N2851, N2847, N2345);
nor NOR4 (N2852, N2833, N1667, N2029, N2766);
or OR3 (N2853, N2849, N530, N1487);
not NOT1 (N2854, N2853);
or OR4 (N2855, N2843, N1056, N1822, N1492);
not NOT1 (N2856, N2846);
nand NAND2 (N2857, N2844, N880);
nor NOR2 (N2858, N2851, N2214);
and AND2 (N2859, N2854, N1492);
or OR3 (N2860, N2855, N1225, N2357);
buf BUF1 (N2861, N2857);
and AND2 (N2862, N2856, N1825);
nand NAND2 (N2863, N2859, N1483);
xor XOR2 (N2864, N2860, N1240);
not NOT1 (N2865, N2852);
buf BUF1 (N2866, N2834);
or OR4 (N2867, N2858, N999, N875, N2388);
not NOT1 (N2868, N2842);
buf BUF1 (N2869, N2850);
or OR4 (N2870, N2862, N2109, N1814, N269);
nand NAND2 (N2871, N2867, N573);
not NOT1 (N2872, N2868);
nor NOR4 (N2873, N2840, N858, N2480, N1879);
xor XOR2 (N2874, N2864, N2418);
or OR2 (N2875, N2871, N345);
not NOT1 (N2876, N2874);
and AND2 (N2877, N2863, N2388);
and AND4 (N2878, N2872, N1001, N312, N1789);
not NOT1 (N2879, N2866);
and AND4 (N2880, N2879, N1805, N1151, N850);
xor XOR2 (N2881, N2873, N2228);
not NOT1 (N2882, N2876);
or OR3 (N2883, N2882, N78, N2602);
xor XOR2 (N2884, N2883, N1990);
not NOT1 (N2885, N2870);
not NOT1 (N2886, N2885);
and AND4 (N2887, N2869, N1073, N1, N921);
nand NAND4 (N2888, N2886, N2864, N801, N1283);
nor NOR4 (N2889, N2888, N435, N1012, N2047);
or OR4 (N2890, N2865, N1403, N2611, N957);
or OR4 (N2891, N2875, N1285, N859, N2071);
buf BUF1 (N2892, N2887);
xor XOR2 (N2893, N2892, N697);
and AND4 (N2894, N2861, N479, N2234, N46);
and AND4 (N2895, N2881, N452, N1031, N1321);
or OR4 (N2896, N2880, N1903, N1559, N1287);
buf BUF1 (N2897, N2884);
xor XOR2 (N2898, N2897, N8);
and AND2 (N2899, N2890, N497);
nand NAND2 (N2900, N2877, N2123);
buf BUF1 (N2901, N2889);
or OR4 (N2902, N2893, N792, N2342, N2104);
and AND3 (N2903, N2896, N1966, N1038);
or OR2 (N2904, N2901, N2165);
and AND2 (N2905, N2904, N348);
nor NOR2 (N2906, N2905, N1063);
nand NAND3 (N2907, N2891, N240, N2182);
not NOT1 (N2908, N2900);
nand NAND2 (N2909, N2903, N2660);
nor NOR4 (N2910, N2909, N900, N844, N2313);
not NOT1 (N2911, N2878);
and AND3 (N2912, N2894, N533, N2252);
or OR4 (N2913, N2898, N674, N114, N1852);
not NOT1 (N2914, N2899);
xor XOR2 (N2915, N2912, N923);
not NOT1 (N2916, N2907);
nor NOR2 (N2917, N2911, N27);
xor XOR2 (N2918, N2917, N1085);
buf BUF1 (N2919, N2908);
xor XOR2 (N2920, N2915, N1506);
nor NOR4 (N2921, N2906, N1858, N1104, N599);
nand NAND4 (N2922, N2921, N1483, N1391, N1776);
and AND2 (N2923, N2913, N2224);
not NOT1 (N2924, N2910);
not NOT1 (N2925, N2924);
buf BUF1 (N2926, N2914);
not NOT1 (N2927, N2916);
nand NAND2 (N2928, N2895, N2673);
buf BUF1 (N2929, N2923);
buf BUF1 (N2930, N2927);
nor NOR3 (N2931, N2930, N2436, N115);
nor NOR4 (N2932, N2918, N175, N1625, N962);
or OR4 (N2933, N2902, N1422, N2015, N2698);
buf BUF1 (N2934, N2919);
nor NOR3 (N2935, N2928, N1569, N2546);
buf BUF1 (N2936, N2932);
and AND3 (N2937, N2936, N2810, N78);
not NOT1 (N2938, N2929);
buf BUF1 (N2939, N2935);
buf BUF1 (N2940, N2937);
not NOT1 (N2941, N2934);
nand NAND3 (N2942, N2926, N1768, N415);
xor XOR2 (N2943, N2942, N1092);
and AND2 (N2944, N2925, N2514);
and AND4 (N2945, N2939, N2764, N1117, N1307);
or OR3 (N2946, N2945, N2799, N1496);
and AND2 (N2947, N2938, N435);
and AND4 (N2948, N2947, N1814, N1642, N1303);
nor NOR4 (N2949, N2922, N2235, N1945, N2072);
not NOT1 (N2950, N2946);
or OR3 (N2951, N2941, N1128, N363);
nor NOR3 (N2952, N2951, N1290, N2708);
or OR3 (N2953, N2920, N2626, N2054);
nor NOR4 (N2954, N2943, N1301, N549, N2284);
buf BUF1 (N2955, N2952);
buf BUF1 (N2956, N2950);
not NOT1 (N2957, N2933);
nand NAND2 (N2958, N2953, N844);
xor XOR2 (N2959, N2931, N879);
xor XOR2 (N2960, N2954, N795);
or OR4 (N2961, N2955, N190, N1700, N824);
not NOT1 (N2962, N2944);
nand NAND4 (N2963, N2961, N1144, N87, N2010);
and AND4 (N2964, N2960, N372, N681, N1027);
xor XOR2 (N2965, N2959, N2840);
xor XOR2 (N2966, N2940, N488);
xor XOR2 (N2967, N2962, N459);
and AND2 (N2968, N2967, N1791);
and AND4 (N2969, N2948, N2637, N2116, N322);
nor NOR2 (N2970, N2958, N1324);
xor XOR2 (N2971, N2966, N1352);
or OR3 (N2972, N2971, N833, N1648);
xor XOR2 (N2973, N2956, N570);
not NOT1 (N2974, N2965);
buf BUF1 (N2975, N2949);
nand NAND2 (N2976, N2968, N2146);
or OR3 (N2977, N2974, N2204, N2803);
buf BUF1 (N2978, N2970);
xor XOR2 (N2979, N2969, N1153);
and AND3 (N2980, N2973, N1643, N2730);
or OR4 (N2981, N2972, N1749, N2418, N1866);
not NOT1 (N2982, N2980);
and AND4 (N2983, N2975, N1186, N1992, N1878);
not NOT1 (N2984, N2978);
not NOT1 (N2985, N2976);
buf BUF1 (N2986, N2983);
nor NOR4 (N2987, N2986, N102, N392, N1871);
xor XOR2 (N2988, N2963, N2585);
nor NOR3 (N2989, N2987, N1101, N1896);
xor XOR2 (N2990, N2981, N2396);
buf BUF1 (N2991, N2957);
and AND2 (N2992, N2988, N2525);
nand NAND3 (N2993, N2984, N2494, N688);
xor XOR2 (N2994, N2964, N276);
xor XOR2 (N2995, N2982, N2296);
xor XOR2 (N2996, N2985, N859);
nor NOR3 (N2997, N2993, N1237, N1975);
buf BUF1 (N2998, N2992);
not NOT1 (N2999, N2990);
buf BUF1 (N3000, N2989);
xor XOR2 (N3001, N2996, N1122);
buf BUF1 (N3002, N2999);
not NOT1 (N3003, N3001);
nor NOR3 (N3004, N2991, N2463, N2390);
not NOT1 (N3005, N3003);
or OR4 (N3006, N2979, N722, N552, N793);
not NOT1 (N3007, N3002);
and AND4 (N3008, N3005, N1905, N1492, N1021);
or OR2 (N3009, N2977, N2778);
and AND4 (N3010, N2994, N855, N364, N1652);
or OR2 (N3011, N2998, N188);
not NOT1 (N3012, N2995);
xor XOR2 (N3013, N3012, N138);
and AND3 (N3014, N3010, N1724, N444);
nor NOR3 (N3015, N3013, N2770, N2956);
xor XOR2 (N3016, N3004, N1217);
or OR2 (N3017, N3009, N1806);
xor XOR2 (N3018, N3017, N1109);
not NOT1 (N3019, N2997);
and AND4 (N3020, N3016, N2487, N2977, N465);
buf BUF1 (N3021, N3006);
nand NAND4 (N3022, N3014, N2977, N2045, N1233);
buf BUF1 (N3023, N3021);
or OR4 (N3024, N3011, N756, N1338, N1280);
and AND3 (N3025, N3015, N2169, N2407);
and AND2 (N3026, N3018, N2270);
buf BUF1 (N3027, N3000);
and AND4 (N3028, N3023, N1729, N1159, N1883);
not NOT1 (N3029, N3007);
nor NOR2 (N3030, N3020, N55);
not NOT1 (N3031, N3028);
buf BUF1 (N3032, N3030);
or OR2 (N3033, N3027, N1252);
nand NAND3 (N3034, N3026, N1023, N506);
nand NAND4 (N3035, N3019, N338, N1379, N977);
nand NAND4 (N3036, N3031, N2064, N2582, N305);
buf BUF1 (N3037, N3036);
buf BUF1 (N3038, N3024);
nor NOR2 (N3039, N3037, N720);
or OR2 (N3040, N3035, N557);
buf BUF1 (N3041, N3029);
nor NOR2 (N3042, N3039, N1234);
or OR2 (N3043, N3008, N1059);
nor NOR4 (N3044, N3034, N467, N2121, N1357);
and AND3 (N3045, N3025, N754, N2392);
and AND4 (N3046, N3022, N1204, N2673, N2316);
nor NOR2 (N3047, N3044, N2237);
and AND4 (N3048, N3041, N108, N331, N466);
not NOT1 (N3049, N3033);
buf BUF1 (N3050, N3047);
not NOT1 (N3051, N3042);
or OR2 (N3052, N3038, N921);
or OR4 (N3053, N3032, N2631, N2116, N2332);
and AND3 (N3054, N3052, N2946, N516);
xor XOR2 (N3055, N3040, N1784);
and AND2 (N3056, N3050, N1620);
not NOT1 (N3057, N3043);
xor XOR2 (N3058, N3057, N1414);
nor NOR3 (N3059, N3049, N2932, N575);
and AND4 (N3060, N3055, N1839, N938, N249);
or OR2 (N3061, N3045, N874);
buf BUF1 (N3062, N3058);
not NOT1 (N3063, N3062);
nor NOR3 (N3064, N3051, N948, N328);
nor NOR2 (N3065, N3061, N974);
nor NOR3 (N3066, N3060, N1362, N2172);
not NOT1 (N3067, N3059);
not NOT1 (N3068, N3053);
and AND2 (N3069, N3063, N2735);
nand NAND3 (N3070, N3068, N1907, N2432);
or OR4 (N3071, N3056, N2177, N801, N2717);
not NOT1 (N3072, N3070);
buf BUF1 (N3073, N3069);
or OR3 (N3074, N3046, N3006, N453);
nand NAND2 (N3075, N3066, N1637);
nor NOR2 (N3076, N3075, N1791);
xor XOR2 (N3077, N3065, N1337);
xor XOR2 (N3078, N3074, N1071);
buf BUF1 (N3079, N3076);
buf BUF1 (N3080, N3064);
and AND4 (N3081, N3078, N897, N1475, N1358);
buf BUF1 (N3082, N3081);
and AND4 (N3083, N3080, N2798, N2889, N950);
not NOT1 (N3084, N3072);
not NOT1 (N3085, N3071);
and AND2 (N3086, N3073, N367);
xor XOR2 (N3087, N3082, N1700);
nor NOR3 (N3088, N3084, N1128, N2238);
nand NAND4 (N3089, N3054, N2749, N1794, N265);
and AND3 (N3090, N3079, N603, N2689);
buf BUF1 (N3091, N3048);
not NOT1 (N3092, N3089);
or OR3 (N3093, N3067, N941, N2496);
nor NOR2 (N3094, N3090, N537);
buf BUF1 (N3095, N3093);
and AND3 (N3096, N3094, N2445, N2963);
and AND4 (N3097, N3083, N1566, N1431, N2497);
xor XOR2 (N3098, N3091, N1297);
and AND2 (N3099, N3077, N2205);
not NOT1 (N3100, N3087);
or OR4 (N3101, N3097, N1477, N2527, N1158);
nor NOR3 (N3102, N3092, N1688, N1032);
xor XOR2 (N3103, N3096, N1995);
xor XOR2 (N3104, N3102, N2524);
or OR2 (N3105, N3098, N1108);
and AND3 (N3106, N3095, N2041, N2525);
nor NOR2 (N3107, N3085, N1226);
nand NAND4 (N3108, N3100, N1701, N247, N599);
and AND2 (N3109, N3088, N2604);
xor XOR2 (N3110, N3101, N599);
xor XOR2 (N3111, N3108, N1314);
and AND2 (N3112, N3099, N2353);
buf BUF1 (N3113, N3107);
nand NAND2 (N3114, N3112, N992);
xor XOR2 (N3115, N3086, N2752);
nor NOR3 (N3116, N3106, N1697, N680);
buf BUF1 (N3117, N3109);
nand NAND2 (N3118, N3111, N268);
buf BUF1 (N3119, N3118);
not NOT1 (N3120, N3113);
or OR3 (N3121, N3114, N2730, N1804);
nor NOR3 (N3122, N3117, N1970, N408);
xor XOR2 (N3123, N3104, N826);
and AND2 (N3124, N3115, N762);
not NOT1 (N3125, N3121);
not NOT1 (N3126, N3124);
and AND4 (N3127, N3105, N2021, N491, N2718);
and AND3 (N3128, N3125, N2288, N2758);
xor XOR2 (N3129, N3126, N3009);
nor NOR4 (N3130, N3123, N2896, N2082, N1866);
nor NOR4 (N3131, N3110, N2417, N83, N1896);
and AND2 (N3132, N3127, N268);
and AND4 (N3133, N3129, N2294, N2259, N1720);
and AND4 (N3134, N3120, N1052, N650, N1979);
nand NAND3 (N3135, N3130, N1918, N871);
not NOT1 (N3136, N3116);
not NOT1 (N3137, N3119);
nand NAND3 (N3138, N3137, N2124, N2310);
and AND3 (N3139, N3128, N3039, N1758);
nor NOR4 (N3140, N3131, N1872, N2231, N710);
not NOT1 (N3141, N3132);
not NOT1 (N3142, N3103);
buf BUF1 (N3143, N3140);
not NOT1 (N3144, N3135);
nand NAND2 (N3145, N3142, N1236);
and AND2 (N3146, N3136, N72);
nand NAND4 (N3147, N3133, N453, N1050, N1212);
not NOT1 (N3148, N3146);
and AND4 (N3149, N3134, N2947, N1819, N1169);
buf BUF1 (N3150, N3149);
or OR2 (N3151, N3139, N1045);
xor XOR2 (N3152, N3141, N1991);
and AND3 (N3153, N3150, N2199, N1394);
buf BUF1 (N3154, N3145);
nand NAND4 (N3155, N3151, N2582, N1735, N1394);
not NOT1 (N3156, N3143);
nor NOR3 (N3157, N3148, N1406, N1165);
and AND3 (N3158, N3157, N1389, N136);
or OR4 (N3159, N3144, N156, N2575, N2835);
buf BUF1 (N3160, N3147);
buf BUF1 (N3161, N3155);
xor XOR2 (N3162, N3152, N2762);
or OR2 (N3163, N3153, N466);
buf BUF1 (N3164, N3138);
and AND2 (N3165, N3122, N37);
or OR3 (N3166, N3160, N1786, N1864);
or OR4 (N3167, N3159, N2017, N2678, N2574);
or OR3 (N3168, N3164, N1408, N518);
nand NAND4 (N3169, N3163, N2510, N2267, N1641);
or OR3 (N3170, N3166, N1667, N1225);
nor NOR4 (N3171, N3168, N1357, N1098, N156);
nor NOR4 (N3172, N3162, N1124, N2572, N2998);
nor NOR3 (N3173, N3167, N207, N1982);
or OR2 (N3174, N3172, N664);
nand NAND2 (N3175, N3158, N2969);
not NOT1 (N3176, N3156);
or OR2 (N3177, N3171, N2075);
and AND4 (N3178, N3154, N1989, N479, N681);
xor XOR2 (N3179, N3169, N2073);
nor NOR2 (N3180, N3173, N2966);
and AND2 (N3181, N3179, N1754);
buf BUF1 (N3182, N3180);
buf BUF1 (N3183, N3177);
or OR4 (N3184, N3165, N2280, N2721, N303);
and AND3 (N3185, N3176, N480, N275);
or OR4 (N3186, N3175, N2388, N67, N2901);
not NOT1 (N3187, N3174);
nor NOR4 (N3188, N3185, N1117, N1603, N434);
nand NAND2 (N3189, N3182, N2959);
not NOT1 (N3190, N3184);
buf BUF1 (N3191, N3190);
not NOT1 (N3192, N3188);
not NOT1 (N3193, N3161);
buf BUF1 (N3194, N3181);
buf BUF1 (N3195, N3170);
or OR4 (N3196, N3178, N483, N16, N2986);
xor XOR2 (N3197, N3193, N1648);
not NOT1 (N3198, N3183);
and AND4 (N3199, N3197, N32, N1301, N2368);
and AND2 (N3200, N3189, N1066);
not NOT1 (N3201, N3187);
and AND2 (N3202, N3198, N2493);
xor XOR2 (N3203, N3202, N2932);
nor NOR2 (N3204, N3192, N2604);
and AND4 (N3205, N3195, N1490, N2649, N1560);
xor XOR2 (N3206, N3204, N2144);
nor NOR3 (N3207, N3205, N2652, N1849);
and AND4 (N3208, N3201, N3029, N2137, N593);
and AND3 (N3209, N3186, N3174, N3033);
xor XOR2 (N3210, N3207, N952);
buf BUF1 (N3211, N3194);
nor NOR3 (N3212, N3211, N1297, N1035);
nand NAND4 (N3213, N3210, N2121, N128, N489);
and AND4 (N3214, N3203, N2085, N2657, N1528);
or OR4 (N3215, N3196, N946, N2423, N1533);
xor XOR2 (N3216, N3191, N1356);
nor NOR4 (N3217, N3206, N2958, N104, N1994);
and AND2 (N3218, N3209, N225);
nor NOR4 (N3219, N3215, N322, N1528, N2849);
or OR4 (N3220, N3214, N2737, N3107, N1977);
not NOT1 (N3221, N3212);
nor NOR4 (N3222, N3217, N966, N280, N1720);
xor XOR2 (N3223, N3222, N138);
nor NOR3 (N3224, N3219, N2318, N2429);
nand NAND4 (N3225, N3223, N1650, N152, N45);
xor XOR2 (N3226, N3199, N869);
or OR4 (N3227, N3213, N1789, N168, N1703);
buf BUF1 (N3228, N3200);
not NOT1 (N3229, N3226);
buf BUF1 (N3230, N3216);
nand NAND2 (N3231, N3229, N496);
or OR2 (N3232, N3227, N40);
not NOT1 (N3233, N3230);
nor NOR2 (N3234, N3228, N1654);
nor NOR4 (N3235, N3234, N2659, N71, N12);
or OR2 (N3236, N3225, N1826);
buf BUF1 (N3237, N3231);
and AND2 (N3238, N3233, N1055);
nand NAND3 (N3239, N3220, N2162, N1269);
nand NAND2 (N3240, N3238, N1649);
nor NOR4 (N3241, N3239, N1502, N1221, N117);
xor XOR2 (N3242, N3235, N1704);
xor XOR2 (N3243, N3242, N394);
and AND3 (N3244, N3237, N31, N2199);
nor NOR2 (N3245, N3232, N2477);
xor XOR2 (N3246, N3241, N1332);
buf BUF1 (N3247, N3243);
buf BUF1 (N3248, N3246);
buf BUF1 (N3249, N3236);
xor XOR2 (N3250, N3224, N1743);
buf BUF1 (N3251, N3244);
buf BUF1 (N3252, N3248);
buf BUF1 (N3253, N3221);
or OR3 (N3254, N3252, N603, N2821);
xor XOR2 (N3255, N3250, N2292);
not NOT1 (N3256, N3255);
and AND3 (N3257, N3247, N1044, N901);
and AND4 (N3258, N3251, N665, N1907, N1575);
not NOT1 (N3259, N3218);
nand NAND3 (N3260, N3259, N753, N103);
not NOT1 (N3261, N3258);
nand NAND3 (N3262, N3249, N2522, N3221);
not NOT1 (N3263, N3208);
nand NAND4 (N3264, N3261, N1203, N2723, N293);
and AND4 (N3265, N3253, N1312, N853, N723);
nand NAND4 (N3266, N3254, N1686, N1674, N2051);
or OR4 (N3267, N3265, N314, N2878, N871);
or OR4 (N3268, N3266, N2375, N838, N2336);
xor XOR2 (N3269, N3257, N1261);
nand NAND4 (N3270, N3256, N1230, N3106, N1025);
and AND2 (N3271, N3268, N663);
nor NOR3 (N3272, N3270, N2032, N2014);
nor NOR4 (N3273, N3267, N1612, N2175, N1032);
and AND2 (N3274, N3264, N249);
nand NAND3 (N3275, N3263, N333, N2304);
or OR2 (N3276, N3272, N1401);
or OR3 (N3277, N3260, N1607, N1711);
and AND3 (N3278, N3271, N1454, N495);
nand NAND4 (N3279, N3274, N259, N1616, N245);
or OR3 (N3280, N3245, N1157, N2070);
nand NAND2 (N3281, N3279, N2431);
nand NAND2 (N3282, N3240, N810);
nand NAND3 (N3283, N3262, N2971, N987);
nand NAND3 (N3284, N3283, N1998, N206);
buf BUF1 (N3285, N3277);
xor XOR2 (N3286, N3284, N2983);
buf BUF1 (N3287, N3275);
buf BUF1 (N3288, N3286);
and AND4 (N3289, N3287, N2134, N612, N537);
nor NOR4 (N3290, N3288, N1038, N650, N1406);
nor NOR3 (N3291, N3282, N1276, N1468);
nor NOR3 (N3292, N3285, N1318, N775);
or OR3 (N3293, N3290, N2363, N2798);
xor XOR2 (N3294, N3278, N3123);
nand NAND4 (N3295, N3281, N1033, N3248, N1324);
and AND4 (N3296, N3294, N2179, N1940, N806);
nor NOR4 (N3297, N3293, N2308, N1798, N2312);
not NOT1 (N3298, N3297);
buf BUF1 (N3299, N3291);
nor NOR4 (N3300, N3298, N946, N30, N695);
nor NOR3 (N3301, N3289, N1179, N1667);
buf BUF1 (N3302, N3295);
or OR4 (N3303, N3299, N3006, N658, N2299);
or OR4 (N3304, N3301, N1695, N2478, N1752);
nor NOR2 (N3305, N3292, N1397);
and AND4 (N3306, N3303, N2380, N1713, N698);
nand NAND3 (N3307, N3304, N124, N1540);
nor NOR4 (N3308, N3276, N68, N1647, N2895);
nand NAND3 (N3309, N3269, N3076, N1508);
nor NOR3 (N3310, N3280, N2957, N1713);
nand NAND3 (N3311, N3307, N364, N1408);
and AND4 (N3312, N3296, N2661, N2338, N3212);
or OR3 (N3313, N3310, N1318, N2617);
xor XOR2 (N3314, N3312, N2091);
or OR2 (N3315, N3309, N497);
xor XOR2 (N3316, N3305, N647);
nand NAND4 (N3317, N3273, N364, N3003, N260);
not NOT1 (N3318, N3311);
nor NOR3 (N3319, N3306, N902, N232);
xor XOR2 (N3320, N3313, N2553);
nand NAND2 (N3321, N3315, N472);
buf BUF1 (N3322, N3320);
or OR3 (N3323, N3314, N3196, N2799);
or OR3 (N3324, N3302, N2733, N71);
buf BUF1 (N3325, N3316);
not NOT1 (N3326, N3323);
nor NOR3 (N3327, N3321, N192, N2816);
not NOT1 (N3328, N3318);
and AND4 (N3329, N3300, N2161, N1015, N2634);
xor XOR2 (N3330, N3325, N3150);
not NOT1 (N3331, N3327);
nor NOR2 (N3332, N3328, N2343);
buf BUF1 (N3333, N3329);
nor NOR4 (N3334, N3326, N1090, N1561, N2279);
nor NOR4 (N3335, N3332, N3310, N2603, N1939);
buf BUF1 (N3336, N3317);
nor NOR3 (N3337, N3308, N817, N1517);
xor XOR2 (N3338, N3336, N1261);
and AND4 (N3339, N3333, N3207, N1782, N268);
nand NAND3 (N3340, N3334, N2672, N1791);
and AND3 (N3341, N3339, N1319, N1274);
not NOT1 (N3342, N3337);
or OR3 (N3343, N3342, N1308, N2408);
nor NOR3 (N3344, N3340, N2784, N1513);
not NOT1 (N3345, N3343);
xor XOR2 (N3346, N3345, N1027);
nor NOR4 (N3347, N3322, N454, N468, N661);
and AND3 (N3348, N3331, N2598, N1654);
nand NAND2 (N3349, N3324, N1437);
not NOT1 (N3350, N3338);
buf BUF1 (N3351, N3344);
not NOT1 (N3352, N3350);
or OR2 (N3353, N3349, N309);
xor XOR2 (N3354, N3335, N2649);
or OR4 (N3355, N3353, N2892, N2616, N3237);
buf BUF1 (N3356, N3319);
nand NAND4 (N3357, N3348, N1348, N2936, N2475);
and AND3 (N3358, N3346, N756, N2700);
nand NAND2 (N3359, N3356, N584);
nor NOR3 (N3360, N3347, N2725, N2307);
buf BUF1 (N3361, N3352);
nand NAND4 (N3362, N3355, N219, N3273, N2796);
and AND4 (N3363, N3360, N3107, N2530, N3123);
or OR4 (N3364, N3330, N3276, N3141, N1388);
not NOT1 (N3365, N3354);
xor XOR2 (N3366, N3351, N2481);
nand NAND4 (N3367, N3358, N2947, N2543, N3291);
not NOT1 (N3368, N3359);
not NOT1 (N3369, N3364);
buf BUF1 (N3370, N3357);
nand NAND4 (N3371, N3363, N2288, N2196, N3269);
not NOT1 (N3372, N3361);
nor NOR2 (N3373, N3365, N222);
nor NOR4 (N3374, N3341, N1015, N1778, N1052);
or OR3 (N3375, N3374, N2067, N3157);
buf BUF1 (N3376, N3372);
buf BUF1 (N3377, N3376);
not NOT1 (N3378, N3368);
nor NOR3 (N3379, N3366, N1410, N1123);
nor NOR4 (N3380, N3370, N1587, N2851, N1802);
and AND3 (N3381, N3375, N1085, N244);
buf BUF1 (N3382, N3381);
nor NOR2 (N3383, N3373, N2053);
not NOT1 (N3384, N3380);
nand NAND2 (N3385, N3379, N472);
nor NOR2 (N3386, N3367, N1459);
or OR2 (N3387, N3362, N3253);
or OR2 (N3388, N3382, N2995);
nand NAND3 (N3389, N3371, N2320, N2224);
or OR2 (N3390, N3369, N2050);
nor NOR2 (N3391, N3389, N1149);
and AND3 (N3392, N3378, N974, N2724);
buf BUF1 (N3393, N3386);
buf BUF1 (N3394, N3387);
nand NAND4 (N3395, N3394, N2875, N1619, N3284);
nor NOR3 (N3396, N3385, N3345, N968);
and AND4 (N3397, N3392, N1293, N2567, N1285);
xor XOR2 (N3398, N3377, N286);
not NOT1 (N3399, N3398);
buf BUF1 (N3400, N3384);
nor NOR2 (N3401, N3383, N1047);
nor NOR2 (N3402, N3399, N165);
buf BUF1 (N3403, N3395);
not NOT1 (N3404, N3397);
and AND4 (N3405, N3390, N2398, N3014, N712);
buf BUF1 (N3406, N3401);
nor NOR4 (N3407, N3400, N948, N1296, N3145);
buf BUF1 (N3408, N3407);
nor NOR4 (N3409, N3402, N355, N819, N956);
nand NAND2 (N3410, N3406, N1204);
buf BUF1 (N3411, N3410);
nor NOR3 (N3412, N3409, N2839, N2808);
nor NOR3 (N3413, N3391, N1480, N1000);
not NOT1 (N3414, N3396);
nor NOR2 (N3415, N3413, N2751);
nor NOR4 (N3416, N3405, N2974, N2755, N2348);
nor NOR3 (N3417, N3412, N2391, N834);
or OR4 (N3418, N3416, N1527, N2826, N387);
not NOT1 (N3419, N3411);
xor XOR2 (N3420, N3418, N2693);
or OR3 (N3421, N3417, N3188, N278);
not NOT1 (N3422, N3393);
and AND4 (N3423, N3421, N2450, N1065, N1602);
or OR3 (N3424, N3420, N1799, N3154);
and AND3 (N3425, N3423, N1648, N3400);
not NOT1 (N3426, N3404);
nor NOR2 (N3427, N3426, N2657);
and AND3 (N3428, N3427, N2956, N722);
not NOT1 (N3429, N3388);
buf BUF1 (N3430, N3429);
and AND2 (N3431, N3408, N1094);
buf BUF1 (N3432, N3403);
nand NAND3 (N3433, N3432, N1403, N729);
nand NAND4 (N3434, N3431, N2566, N4, N1913);
buf BUF1 (N3435, N3433);
buf BUF1 (N3436, N3414);
buf BUF1 (N3437, N3419);
xor XOR2 (N3438, N3415, N1593);
xor XOR2 (N3439, N3438, N940);
xor XOR2 (N3440, N3428, N2957);
or OR4 (N3441, N3439, N744, N1679, N1678);
nor NOR4 (N3442, N3422, N848, N1088, N203);
not NOT1 (N3443, N3442);
xor XOR2 (N3444, N3424, N1806);
nand NAND4 (N3445, N3436, N168, N2221, N1421);
not NOT1 (N3446, N3435);
or OR4 (N3447, N3441, N608, N3058, N439);
and AND2 (N3448, N3437, N2932);
buf BUF1 (N3449, N3447);
not NOT1 (N3450, N3443);
xor XOR2 (N3451, N3440, N832);
and AND4 (N3452, N3451, N2730, N2069, N3232);
and AND4 (N3453, N3450, N1399, N1897, N3234);
nand NAND4 (N3454, N3446, N1000, N970, N2330);
or OR4 (N3455, N3444, N2052, N3270, N2408);
not NOT1 (N3456, N3449);
and AND4 (N3457, N3452, N885, N1675, N3226);
and AND4 (N3458, N3448, N2536, N2821, N2787);
nor NOR4 (N3459, N3434, N233, N500, N1474);
buf BUF1 (N3460, N3459);
xor XOR2 (N3461, N3460, N3315);
or OR4 (N3462, N3454, N2672, N3056, N3164);
xor XOR2 (N3463, N3458, N1572);
nor NOR3 (N3464, N3425, N2869, N1708);
nand NAND2 (N3465, N3453, N2217);
buf BUF1 (N3466, N3455);
nor NOR2 (N3467, N3462, N1449);
buf BUF1 (N3468, N3430);
xor XOR2 (N3469, N3463, N1384);
not NOT1 (N3470, N3467);
nand NAND2 (N3471, N3456, N1532);
or OR4 (N3472, N3461, N1606, N2598, N3400);
xor XOR2 (N3473, N3469, N1482);
not NOT1 (N3474, N3472);
nand NAND4 (N3475, N3445, N1214, N1709, N2657);
or OR3 (N3476, N3475, N104, N2816);
nor NOR2 (N3477, N3457, N687);
not NOT1 (N3478, N3470);
or OR4 (N3479, N3465, N351, N1845, N774);
buf BUF1 (N3480, N3478);
buf BUF1 (N3481, N3477);
xor XOR2 (N3482, N3473, N1784);
nand NAND2 (N3483, N3474, N3478);
buf BUF1 (N3484, N3482);
and AND4 (N3485, N3484, N2601, N1706, N2220);
buf BUF1 (N3486, N3471);
buf BUF1 (N3487, N3480);
buf BUF1 (N3488, N3466);
not NOT1 (N3489, N3476);
buf BUF1 (N3490, N3483);
nor NOR4 (N3491, N3485, N2470, N1907, N2389);
xor XOR2 (N3492, N3488, N1667);
nor NOR3 (N3493, N3481, N302, N320);
and AND2 (N3494, N3479, N3130);
and AND4 (N3495, N3468, N2642, N2153, N927);
and AND2 (N3496, N3495, N2632);
buf BUF1 (N3497, N3493);
xor XOR2 (N3498, N3494, N2353);
nor NOR2 (N3499, N3490, N2916);
xor XOR2 (N3500, N3497, N2665);
nor NOR3 (N3501, N3498, N1307, N3008);
not NOT1 (N3502, N3496);
nand NAND3 (N3503, N3492, N779, N1739);
not NOT1 (N3504, N3464);
buf BUF1 (N3505, N3501);
or OR3 (N3506, N3487, N2745, N3396);
xor XOR2 (N3507, N3489, N3125);
and AND3 (N3508, N3491, N2057, N536);
nor NOR4 (N3509, N3503, N444, N2090, N1956);
xor XOR2 (N3510, N3509, N905);
nand NAND4 (N3511, N3502, N2339, N980, N1960);
xor XOR2 (N3512, N3508, N542);
not NOT1 (N3513, N3504);
buf BUF1 (N3514, N3510);
and AND3 (N3515, N3506, N2195, N143);
nand NAND3 (N3516, N3514, N984, N1066);
nand NAND3 (N3517, N3500, N2686, N2072);
nand NAND2 (N3518, N3512, N2932);
nor NOR4 (N3519, N3513, N2290, N2783, N2278);
not NOT1 (N3520, N3518);
and AND4 (N3521, N3507, N2849, N507, N2735);
buf BUF1 (N3522, N3505);
xor XOR2 (N3523, N3499, N2328);
and AND3 (N3524, N3486, N1933, N2928);
nor NOR2 (N3525, N3523, N767);
nor NOR2 (N3526, N3517, N1195);
xor XOR2 (N3527, N3526, N2979);
and AND3 (N3528, N3520, N2061, N2760);
buf BUF1 (N3529, N3519);
or OR2 (N3530, N3524, N372);
nor NOR2 (N3531, N3516, N43);
or OR3 (N3532, N3522, N3211, N707);
or OR2 (N3533, N3528, N971);
not NOT1 (N3534, N3511);
nand NAND2 (N3535, N3533, N1279);
nor NOR2 (N3536, N3530, N121);
buf BUF1 (N3537, N3525);
buf BUF1 (N3538, N3535);
nand NAND2 (N3539, N3531, N1472);
and AND2 (N3540, N3529, N333);
or OR2 (N3541, N3521, N389);
buf BUF1 (N3542, N3532);
xor XOR2 (N3543, N3534, N2154);
and AND4 (N3544, N3538, N944, N915, N1936);
not NOT1 (N3545, N3527);
not NOT1 (N3546, N3543);
and AND4 (N3547, N3515, N1023, N2600, N1049);
or OR4 (N3548, N3536, N2460, N1452, N530);
xor XOR2 (N3549, N3541, N854);
not NOT1 (N3550, N3548);
nand NAND3 (N3551, N3537, N3458, N866);
xor XOR2 (N3552, N3549, N3075);
not NOT1 (N3553, N3552);
nand NAND2 (N3554, N3550, N784);
xor XOR2 (N3555, N3553, N310);
or OR3 (N3556, N3540, N615, N2140);
not NOT1 (N3557, N3551);
or OR2 (N3558, N3554, N1718);
nor NOR4 (N3559, N3539, N3075, N92, N3210);
nand NAND2 (N3560, N3544, N1322);
nand NAND4 (N3561, N3557, N467, N2462, N1874);
nor NOR3 (N3562, N3555, N3514, N1918);
nand NAND2 (N3563, N3562, N2707);
nand NAND3 (N3564, N3559, N1952, N1281);
or OR4 (N3565, N3546, N1114, N3358, N1749);
and AND3 (N3566, N3564, N1979, N2399);
xor XOR2 (N3567, N3563, N2981);
not NOT1 (N3568, N3556);
nand NAND3 (N3569, N3567, N712, N830);
nor NOR3 (N3570, N3561, N1468, N3188);
buf BUF1 (N3571, N3547);
or OR4 (N3572, N3545, N3025, N2169, N2475);
nor NOR2 (N3573, N3568, N1655);
not NOT1 (N3574, N3569);
nor NOR3 (N3575, N3574, N2747, N1224);
buf BUF1 (N3576, N3571);
buf BUF1 (N3577, N3573);
or OR2 (N3578, N3560, N2674);
nor NOR2 (N3579, N3572, N1981);
nor NOR2 (N3580, N3577, N2247);
xor XOR2 (N3581, N3570, N1050);
and AND2 (N3582, N3565, N320);
nand NAND3 (N3583, N3542, N2551, N1415);
or OR2 (N3584, N3578, N2509);
nand NAND2 (N3585, N3579, N1688);
nand NAND3 (N3586, N3576, N1723, N3467);
buf BUF1 (N3587, N3558);
or OR2 (N3588, N3584, N3042);
nand NAND3 (N3589, N3582, N1746, N1784);
or OR4 (N3590, N3588, N15, N2305, N2746);
xor XOR2 (N3591, N3566, N148);
nand NAND3 (N3592, N3580, N503, N849);
xor XOR2 (N3593, N3591, N3381);
xor XOR2 (N3594, N3585, N3210);
nand NAND4 (N3595, N3586, N603, N1432, N3178);
nor NOR2 (N3596, N3575, N2944);
xor XOR2 (N3597, N3593, N3226);
xor XOR2 (N3598, N3590, N2618);
or OR4 (N3599, N3589, N738, N1746, N1332);
buf BUF1 (N3600, N3597);
buf BUF1 (N3601, N3581);
xor XOR2 (N3602, N3592, N1197);
xor XOR2 (N3603, N3587, N703);
buf BUF1 (N3604, N3601);
buf BUF1 (N3605, N3583);
xor XOR2 (N3606, N3600, N173);
or OR3 (N3607, N3603, N404, N2046);
or OR3 (N3608, N3604, N2877, N3155);
buf BUF1 (N3609, N3606);
not NOT1 (N3610, N3595);
or OR4 (N3611, N3609, N958, N2579, N1390);
not NOT1 (N3612, N3605);
buf BUF1 (N3613, N3598);
nand NAND3 (N3614, N3599, N2453, N818);
not NOT1 (N3615, N3594);
not NOT1 (N3616, N3607);
and AND4 (N3617, N3614, N3504, N934, N2551);
nand NAND4 (N3618, N3611, N3439, N1155, N482);
xor XOR2 (N3619, N3596, N2827);
or OR3 (N3620, N3608, N2534, N1622);
nand NAND3 (N3621, N3616, N599, N2105);
nor NOR2 (N3622, N3617, N1837);
nand NAND3 (N3623, N3615, N127, N978);
not NOT1 (N3624, N3619);
or OR3 (N3625, N3613, N2743, N1914);
and AND3 (N3626, N3623, N1422, N2811);
xor XOR2 (N3627, N3622, N10);
nor NOR4 (N3628, N3626, N857, N1489, N186);
or OR3 (N3629, N3612, N1870, N3588);
xor XOR2 (N3630, N3624, N1316);
or OR3 (N3631, N3628, N3101, N2680);
not NOT1 (N3632, N3629);
xor XOR2 (N3633, N3630, N909);
nor NOR2 (N3634, N3602, N3578);
nor NOR2 (N3635, N3621, N1142);
not NOT1 (N3636, N3633);
and AND2 (N3637, N3618, N2443);
or OR4 (N3638, N3620, N3287, N3420, N1135);
not NOT1 (N3639, N3636);
nand NAND4 (N3640, N3627, N2448, N556, N340);
nor NOR2 (N3641, N3637, N3160);
buf BUF1 (N3642, N3634);
nor NOR2 (N3643, N3610, N2450);
buf BUF1 (N3644, N3641);
or OR3 (N3645, N3640, N2004, N2598);
buf BUF1 (N3646, N3635);
nor NOR2 (N3647, N3625, N628);
nor NOR4 (N3648, N3646, N3376, N959, N3205);
nor NOR2 (N3649, N3632, N1992);
and AND3 (N3650, N3645, N2723, N3003);
buf BUF1 (N3651, N3649);
or OR3 (N3652, N3651, N3186, N2200);
not NOT1 (N3653, N3639);
and AND3 (N3654, N3643, N2300, N892);
buf BUF1 (N3655, N3631);
xor XOR2 (N3656, N3647, N2948);
not NOT1 (N3657, N3654);
and AND4 (N3658, N3644, N3151, N1480, N1998);
buf BUF1 (N3659, N3653);
nand NAND3 (N3660, N3656, N1694, N3272);
buf BUF1 (N3661, N3658);
xor XOR2 (N3662, N3660, N1529);
or OR2 (N3663, N3662, N2512);
and AND3 (N3664, N3648, N2457, N3017);
or OR2 (N3665, N3663, N777);
buf BUF1 (N3666, N3661);
and AND3 (N3667, N3657, N2129, N126);
nand NAND3 (N3668, N3650, N2864, N2538);
xor XOR2 (N3669, N3668, N1687);
xor XOR2 (N3670, N3638, N2764);
or OR3 (N3671, N3642, N2240, N1156);
nand NAND2 (N3672, N3664, N3051);
xor XOR2 (N3673, N3659, N262);
nand NAND3 (N3674, N3652, N1161, N556);
or OR4 (N3675, N3670, N2158, N214, N1828);
xor XOR2 (N3676, N3673, N3305);
buf BUF1 (N3677, N3667);
not NOT1 (N3678, N3674);
not NOT1 (N3679, N3677);
xor XOR2 (N3680, N3671, N890);
and AND4 (N3681, N3666, N98, N2246, N3548);
nand NAND3 (N3682, N3679, N1873, N1275);
and AND3 (N3683, N3655, N2806, N1320);
xor XOR2 (N3684, N3665, N2178);
nor NOR3 (N3685, N3676, N1986, N5);
nand NAND4 (N3686, N3672, N2045, N34, N751);
nor NOR2 (N3687, N3678, N1608);
xor XOR2 (N3688, N3683, N476);
and AND3 (N3689, N3681, N189, N2693);
buf BUF1 (N3690, N3686);
buf BUF1 (N3691, N3669);
not NOT1 (N3692, N3690);
xor XOR2 (N3693, N3685, N919);
nand NAND4 (N3694, N3692, N3022, N3631, N3520);
nor NOR3 (N3695, N3675, N1117, N567);
xor XOR2 (N3696, N3687, N1095);
buf BUF1 (N3697, N3696);
and AND2 (N3698, N3697, N481);
nor NOR4 (N3699, N3680, N3360, N2439, N1053);
and AND2 (N3700, N3699, N2122);
not NOT1 (N3701, N3695);
not NOT1 (N3702, N3701);
buf BUF1 (N3703, N3688);
and AND3 (N3704, N3698, N1661, N399);
or OR3 (N3705, N3689, N148, N186);
not NOT1 (N3706, N3693);
and AND2 (N3707, N3705, N1562);
or OR4 (N3708, N3682, N545, N1644, N2903);
or OR2 (N3709, N3684, N2810);
nand NAND2 (N3710, N3704, N752);
xor XOR2 (N3711, N3700, N1635);
nand NAND4 (N3712, N3706, N1090, N1653, N867);
nand NAND3 (N3713, N3702, N184, N2287);
buf BUF1 (N3714, N3703);
or OR4 (N3715, N3714, N490, N3658, N1537);
and AND4 (N3716, N3711, N2214, N3436, N272);
or OR4 (N3717, N3709, N2883, N480, N1543);
buf BUF1 (N3718, N3715);
nor NOR2 (N3719, N3694, N1858);
buf BUF1 (N3720, N3713);
buf BUF1 (N3721, N3708);
xor XOR2 (N3722, N3721, N1169);
or OR3 (N3723, N3719, N792, N2588);
buf BUF1 (N3724, N3722);
nand NAND4 (N3725, N3716, N1450, N1245, N3352);
buf BUF1 (N3726, N3723);
nor NOR4 (N3727, N3725, N364, N1194, N3304);
not NOT1 (N3728, N3724);
or OR4 (N3729, N3726, N393, N2574, N1691);
xor XOR2 (N3730, N3718, N1089);
or OR2 (N3731, N3717, N986);
not NOT1 (N3732, N3729);
or OR3 (N3733, N3727, N2796, N951);
buf BUF1 (N3734, N3728);
buf BUF1 (N3735, N3731);
xor XOR2 (N3736, N3712, N3655);
xor XOR2 (N3737, N3735, N2919);
buf BUF1 (N3738, N3736);
or OR3 (N3739, N3707, N1745, N3342);
or OR4 (N3740, N3710, N1593, N1554, N160);
not NOT1 (N3741, N3720);
buf BUF1 (N3742, N3734);
nor NOR3 (N3743, N3732, N3575, N3661);
nand NAND2 (N3744, N3738, N1901);
nor NOR3 (N3745, N3740, N1845, N469);
or OR4 (N3746, N3741, N2220, N931, N1247);
or OR2 (N3747, N3744, N580);
not NOT1 (N3748, N3747);
and AND2 (N3749, N3691, N3658);
nor NOR4 (N3750, N3737, N2277, N1835, N2757);
nand NAND3 (N3751, N3748, N369, N611);
buf BUF1 (N3752, N3733);
buf BUF1 (N3753, N3750);
or OR3 (N3754, N3730, N1698, N2475);
nor NOR4 (N3755, N3751, N3191, N1515, N781);
nor NOR2 (N3756, N3742, N452);
xor XOR2 (N3757, N3755, N825);
not NOT1 (N3758, N3739);
and AND3 (N3759, N3754, N899, N2897);
nand NAND2 (N3760, N3756, N979);
and AND4 (N3761, N3758, N1539, N1522, N1309);
nor NOR4 (N3762, N3761, N2838, N269, N2037);
or OR3 (N3763, N3743, N696, N452);
buf BUF1 (N3764, N3753);
not NOT1 (N3765, N3764);
xor XOR2 (N3766, N3745, N3223);
not NOT1 (N3767, N3746);
and AND2 (N3768, N3757, N3220);
buf BUF1 (N3769, N3749);
or OR3 (N3770, N3767, N3192, N1871);
nand NAND4 (N3771, N3759, N3241, N86, N2466);
buf BUF1 (N3772, N3760);
and AND3 (N3773, N3772, N2896, N3359);
or OR4 (N3774, N3769, N1535, N846, N1025);
and AND2 (N3775, N3765, N1306);
and AND3 (N3776, N3768, N1774, N3048);
nor NOR4 (N3777, N3771, N3299, N84, N3303);
not NOT1 (N3778, N3776);
not NOT1 (N3779, N3775);
or OR2 (N3780, N3763, N353);
not NOT1 (N3781, N3777);
xor XOR2 (N3782, N3752, N2081);
xor XOR2 (N3783, N3773, N3428);
or OR2 (N3784, N3781, N2866);
and AND2 (N3785, N3783, N3474);
not NOT1 (N3786, N3766);
and AND3 (N3787, N3780, N3086, N667);
buf BUF1 (N3788, N3784);
buf BUF1 (N3789, N3770);
not NOT1 (N3790, N3774);
and AND3 (N3791, N3786, N2076, N178);
nand NAND2 (N3792, N3778, N729);
or OR4 (N3793, N3787, N2261, N3194, N2819);
not NOT1 (N3794, N3789);
nor NOR2 (N3795, N3793, N2520);
not NOT1 (N3796, N3782);
and AND4 (N3797, N3794, N1571, N893, N419);
not NOT1 (N3798, N3788);
nor NOR4 (N3799, N3785, N1435, N3560, N2299);
nand NAND4 (N3800, N3796, N2970, N811, N2537);
xor XOR2 (N3801, N3790, N1792);
and AND3 (N3802, N3791, N3777, N1998);
nor NOR2 (N3803, N3799, N666);
and AND2 (N3804, N3797, N873);
xor XOR2 (N3805, N3792, N3081);
nor NOR3 (N3806, N3798, N1346, N2198);
or OR2 (N3807, N3779, N2797);
xor XOR2 (N3808, N3800, N3314);
not NOT1 (N3809, N3795);
xor XOR2 (N3810, N3805, N3301);
or OR2 (N3811, N3801, N3294);
buf BUF1 (N3812, N3811);
nor NOR3 (N3813, N3802, N372, N1413);
nand NAND4 (N3814, N3809, N2131, N1048, N102);
nor NOR3 (N3815, N3814, N762, N671);
buf BUF1 (N3816, N3813);
xor XOR2 (N3817, N3803, N3388);
nand NAND4 (N3818, N3808, N1411, N2463, N3779);
nand NAND4 (N3819, N3817, N685, N3541, N3652);
nand NAND3 (N3820, N3804, N1273, N2083);
or OR3 (N3821, N3815, N3293, N3225);
buf BUF1 (N3822, N3806);
nand NAND4 (N3823, N3821, N1837, N1180, N2719);
nor NOR3 (N3824, N3816, N3622, N2117);
and AND3 (N3825, N3824, N2821, N1331);
nor NOR3 (N3826, N3822, N2257, N91);
nand NAND2 (N3827, N3807, N3611);
not NOT1 (N3828, N3819);
not NOT1 (N3829, N3820);
not NOT1 (N3830, N3825);
nand NAND2 (N3831, N3829, N2077);
buf BUF1 (N3832, N3826);
buf BUF1 (N3833, N3812);
or OR3 (N3834, N3810, N1057, N100);
xor XOR2 (N3835, N3833, N1075);
buf BUF1 (N3836, N3762);
nand NAND3 (N3837, N3834, N1875, N1639);
xor XOR2 (N3838, N3828, N3753);
buf BUF1 (N3839, N3837);
xor XOR2 (N3840, N3836, N2121);
nand NAND2 (N3841, N3830, N3021);
buf BUF1 (N3842, N3839);
buf BUF1 (N3843, N3841);
buf BUF1 (N3844, N3818);
and AND4 (N3845, N3832, N1194, N3458, N3507);
xor XOR2 (N3846, N3840, N2002);
or OR4 (N3847, N3844, N2833, N1210, N852);
nand NAND2 (N3848, N3845, N3611);
or OR2 (N3849, N3827, N3432);
nor NOR4 (N3850, N3846, N794, N2204, N3154);
buf BUF1 (N3851, N3847);
nor NOR4 (N3852, N3848, N3197, N2271, N540);
or OR4 (N3853, N3831, N3537, N3110, N106);
buf BUF1 (N3854, N3849);
and AND2 (N3855, N3851, N1476);
not NOT1 (N3856, N3855);
not NOT1 (N3857, N3838);
buf BUF1 (N3858, N3854);
nor NOR2 (N3859, N3853, N1033);
or OR3 (N3860, N3859, N987, N2701);
nor NOR2 (N3861, N3860, N2618);
not NOT1 (N3862, N3856);
xor XOR2 (N3863, N3858, N2216);
nand NAND3 (N3864, N3835, N1387, N1353);
nand NAND2 (N3865, N3852, N1627);
nor NOR3 (N3866, N3864, N414, N2330);
nor NOR2 (N3867, N3857, N1302);
not NOT1 (N3868, N3865);
xor XOR2 (N3869, N3862, N1672);
buf BUF1 (N3870, N3823);
xor XOR2 (N3871, N3842, N1268);
nor NOR4 (N3872, N3869, N1688, N377, N2196);
and AND4 (N3873, N3861, N3376, N3750, N1423);
nand NAND3 (N3874, N3850, N3047, N2506);
nor NOR3 (N3875, N3866, N1845, N710);
nand NAND2 (N3876, N3875, N1052);
nor NOR4 (N3877, N3876, N3394, N2785, N3488);
nand NAND3 (N3878, N3872, N2999, N2373);
xor XOR2 (N3879, N3871, N2370);
nor NOR3 (N3880, N3843, N3731, N1617);
not NOT1 (N3881, N3877);
buf BUF1 (N3882, N3867);
nor NOR4 (N3883, N3873, N3080, N1357, N1188);
not NOT1 (N3884, N3863);
nand NAND2 (N3885, N3879, N2376);
nor NOR3 (N3886, N3882, N519, N2807);
and AND3 (N3887, N3881, N1578, N384);
xor XOR2 (N3888, N3870, N3134);
buf BUF1 (N3889, N3874);
or OR2 (N3890, N3889, N111);
nand NAND4 (N3891, N3883, N1109, N2995, N128);
nor NOR4 (N3892, N3887, N887, N507, N3554);
and AND3 (N3893, N3884, N103, N155);
and AND2 (N3894, N3892, N3869);
nor NOR4 (N3895, N3890, N671, N2897, N238);
or OR2 (N3896, N3880, N813);
nand NAND3 (N3897, N3868, N319, N981);
nand NAND3 (N3898, N3895, N1972, N1229);
nand NAND2 (N3899, N3886, N2638);
and AND3 (N3900, N3899, N81, N759);
buf BUF1 (N3901, N3894);
nand NAND2 (N3902, N3901, N3480);
xor XOR2 (N3903, N3893, N3730);
nor NOR3 (N3904, N3891, N2874, N2282);
nor NOR3 (N3905, N3898, N2333, N373);
xor XOR2 (N3906, N3902, N2854);
or OR2 (N3907, N3906, N3181);
buf BUF1 (N3908, N3878);
buf BUF1 (N3909, N3888);
nand NAND3 (N3910, N3896, N2966, N974);
xor XOR2 (N3911, N3909, N3346);
buf BUF1 (N3912, N3905);
or OR4 (N3913, N3897, N3849, N179, N561);
not NOT1 (N3914, N3900);
and AND2 (N3915, N3911, N2513);
xor XOR2 (N3916, N3915, N2134);
not NOT1 (N3917, N3910);
xor XOR2 (N3918, N3914, N549);
nand NAND2 (N3919, N3904, N3187);
or OR2 (N3920, N3916, N1434);
xor XOR2 (N3921, N3908, N213);
not NOT1 (N3922, N3917);
buf BUF1 (N3923, N3913);
or OR3 (N3924, N3921, N1183, N2424);
xor XOR2 (N3925, N3907, N1909);
and AND2 (N3926, N3903, N44);
xor XOR2 (N3927, N3924, N2417);
nor NOR2 (N3928, N3922, N2322);
nor NOR2 (N3929, N3923, N3619);
and AND4 (N3930, N3925, N3255, N3078, N1812);
xor XOR2 (N3931, N3929, N1396);
buf BUF1 (N3932, N3918);
xor XOR2 (N3933, N3927, N879);
xor XOR2 (N3934, N3928, N3004);
nand NAND2 (N3935, N3919, N2918);
buf BUF1 (N3936, N3912);
xor XOR2 (N3937, N3885, N1509);
not NOT1 (N3938, N3934);
not NOT1 (N3939, N3933);
or OR2 (N3940, N3930, N588);
buf BUF1 (N3941, N3932);
buf BUF1 (N3942, N3940);
nor NOR3 (N3943, N3935, N1269, N199);
nor NOR4 (N3944, N3943, N254, N336, N2352);
buf BUF1 (N3945, N3931);
and AND3 (N3946, N3938, N3388, N2259);
nand NAND4 (N3947, N3939, N179, N1008, N1007);
nor NOR4 (N3948, N3946, N358, N668, N3378);
or OR3 (N3949, N3947, N711, N3419);
and AND2 (N3950, N3948, N1013);
buf BUF1 (N3951, N3945);
xor XOR2 (N3952, N3949, N1423);
or OR4 (N3953, N3941, N1087, N2150, N1690);
not NOT1 (N3954, N3920);
or OR3 (N3955, N3926, N417, N498);
or OR3 (N3956, N3944, N3364, N94);
buf BUF1 (N3957, N3952);
nor NOR3 (N3958, N3951, N1137, N2407);
buf BUF1 (N3959, N3958);
nor NOR3 (N3960, N3953, N813, N2342);
nor NOR4 (N3961, N3959, N3376, N1971, N2557);
not NOT1 (N3962, N3956);
xor XOR2 (N3963, N3957, N3018);
nor NOR4 (N3964, N3955, N1240, N3660, N1541);
nor NOR3 (N3965, N3937, N1125, N1083);
or OR3 (N3966, N3950, N3631, N1227);
not NOT1 (N3967, N3961);
and AND2 (N3968, N3964, N1230);
and AND3 (N3969, N3963, N190, N1640);
or OR2 (N3970, N3967, N1133);
or OR2 (N3971, N3936, N3742);
xor XOR2 (N3972, N3965, N1390);
nor NOR3 (N3973, N3968, N2071, N791);
buf BUF1 (N3974, N3973);
nand NAND2 (N3975, N3970, N3724);
not NOT1 (N3976, N3974);
or OR2 (N3977, N3942, N635);
or OR3 (N3978, N3977, N495, N2819);
and AND2 (N3979, N3966, N683);
and AND2 (N3980, N3969, N1745);
not NOT1 (N3981, N3960);
nor NOR2 (N3982, N3978, N2540);
nor NOR2 (N3983, N3971, N2543);
and AND2 (N3984, N3983, N2674);
buf BUF1 (N3985, N3984);
xor XOR2 (N3986, N3982, N2125);
nor NOR4 (N3987, N3972, N1097, N1156, N785);
or OR3 (N3988, N3985, N1726, N3381);
xor XOR2 (N3989, N3988, N3311);
buf BUF1 (N3990, N3980);
or OR3 (N3991, N3981, N3201, N2401);
not NOT1 (N3992, N3986);
or OR2 (N3993, N3990, N1174);
buf BUF1 (N3994, N3954);
buf BUF1 (N3995, N3975);
and AND4 (N3996, N3994, N3709, N2587, N454);
buf BUF1 (N3997, N3996);
or OR4 (N3998, N3993, N1801, N2543, N1044);
nor NOR4 (N3999, N3992, N3729, N48, N1092);
buf BUF1 (N4000, N3999);
xor XOR2 (N4001, N3995, N1457);
not NOT1 (N4002, N3989);
nor NOR3 (N4003, N3987, N1059, N3758);
or OR2 (N4004, N4000, N3137);
and AND3 (N4005, N3979, N3139, N2145);
nand NAND4 (N4006, N4001, N3226, N89, N1645);
or OR3 (N4007, N3976, N2259, N3532);
and AND2 (N4008, N4002, N1910);
buf BUF1 (N4009, N3991);
nor NOR3 (N4010, N3962, N1751, N3141);
xor XOR2 (N4011, N4004, N832);
buf BUF1 (N4012, N4011);
buf BUF1 (N4013, N4005);
or OR4 (N4014, N4003, N1253, N1320, N1600);
buf BUF1 (N4015, N4006);
or OR3 (N4016, N4010, N1601, N3559);
nor NOR3 (N4017, N4008, N205, N3913);
xor XOR2 (N4018, N4016, N3166);
nand NAND4 (N4019, N4013, N2552, N2665, N3448);
and AND2 (N4020, N3998, N965);
and AND3 (N4021, N3997, N1198, N1284);
and AND2 (N4022, N4020, N2884);
xor XOR2 (N4023, N4019, N1512);
buf BUF1 (N4024, N4023);
and AND4 (N4025, N4018, N3622, N77, N2376);
nand NAND3 (N4026, N4024, N3811, N232);
xor XOR2 (N4027, N4025, N1564);
xor XOR2 (N4028, N4017, N1784);
nor NOR3 (N4029, N4012, N1349, N1973);
and AND3 (N4030, N4015, N2864, N289);
or OR4 (N4031, N4030, N1868, N2122, N3816);
nand NAND2 (N4032, N4009, N1950);
and AND2 (N4033, N4031, N3559);
nand NAND4 (N4034, N4021, N2283, N2584, N1942);
or OR4 (N4035, N4033, N2324, N3999, N693);
and AND4 (N4036, N4034, N2610, N3996, N2602);
nor NOR3 (N4037, N4035, N3485, N34);
not NOT1 (N4038, N4022);
buf BUF1 (N4039, N4014);
or OR3 (N4040, N4038, N2062, N9);
nand NAND3 (N4041, N4028, N2803, N2450);
xor XOR2 (N4042, N4039, N172);
buf BUF1 (N4043, N4027);
not NOT1 (N4044, N4032);
buf BUF1 (N4045, N4041);
xor XOR2 (N4046, N4029, N2282);
nor NOR3 (N4047, N4044, N2608, N2041);
nor NOR3 (N4048, N4026, N2521, N3420);
nor NOR4 (N4049, N4048, N107, N3005, N845);
buf BUF1 (N4050, N4045);
nor NOR3 (N4051, N4043, N98, N3605);
nor NOR3 (N4052, N4046, N1637, N663);
buf BUF1 (N4053, N4049);
and AND2 (N4054, N4042, N2596);
nor NOR4 (N4055, N4050, N3932, N3759, N1299);
xor XOR2 (N4056, N4053, N2256);
buf BUF1 (N4057, N4051);
or OR4 (N4058, N4047, N2626, N188, N3195);
nand NAND4 (N4059, N4036, N480, N1010, N3619);
not NOT1 (N4060, N4059);
nor NOR2 (N4061, N4007, N2480);
buf BUF1 (N4062, N4060);
or OR2 (N4063, N4057, N2449);
or OR4 (N4064, N4055, N2969, N2969, N3394);
buf BUF1 (N4065, N4052);
not NOT1 (N4066, N4056);
and AND3 (N4067, N4062, N1164, N2949);
xor XOR2 (N4068, N4066, N8);
not NOT1 (N4069, N4040);
and AND3 (N4070, N4054, N2149, N2746);
not NOT1 (N4071, N4065);
xor XOR2 (N4072, N4063, N2445);
xor XOR2 (N4073, N4061, N1078);
nor NOR2 (N4074, N4069, N226);
xor XOR2 (N4075, N4067, N2651);
and AND2 (N4076, N4058, N804);
nand NAND3 (N4077, N4070, N2563, N2400);
xor XOR2 (N4078, N4074, N2878);
or OR3 (N4079, N4064, N1477, N2360);
xor XOR2 (N4080, N4072, N3704);
nand NAND2 (N4081, N4079, N1037);
nor NOR2 (N4082, N4081, N1942);
xor XOR2 (N4083, N4080, N1719);
buf BUF1 (N4084, N4075);
and AND4 (N4085, N4076, N1240, N1206, N3704);
nor NOR4 (N4086, N4083, N475, N2686, N1720);
and AND3 (N4087, N4073, N1686, N2612);
not NOT1 (N4088, N4037);
xor XOR2 (N4089, N4078, N3316);
nor NOR2 (N4090, N4085, N1234);
and AND4 (N4091, N4071, N1382, N3661, N1018);
nand NAND3 (N4092, N4082, N2343, N1243);
and AND4 (N4093, N4090, N2690, N1067, N1373);
xor XOR2 (N4094, N4092, N2890);
not NOT1 (N4095, N4088);
nand NAND3 (N4096, N4084, N320, N1055);
buf BUF1 (N4097, N4086);
xor XOR2 (N4098, N4087, N2946);
and AND3 (N4099, N4093, N3275, N902);
nor NOR3 (N4100, N4099, N3047, N547);
and AND4 (N4101, N4068, N759, N836, N516);
not NOT1 (N4102, N4097);
and AND2 (N4103, N4096, N431);
not NOT1 (N4104, N4100);
not NOT1 (N4105, N4103);
nor NOR2 (N4106, N4091, N2591);
or OR4 (N4107, N4106, N1587, N1294, N282);
nand NAND3 (N4108, N4101, N518, N233);
and AND4 (N4109, N4107, N2439, N2622, N584);
not NOT1 (N4110, N4094);
nand NAND4 (N4111, N4089, N3001, N128, N642);
not NOT1 (N4112, N4108);
buf BUF1 (N4113, N4110);
buf BUF1 (N4114, N4112);
nor NOR3 (N4115, N4104, N651, N1855);
and AND2 (N4116, N4077, N609);
nor NOR4 (N4117, N4095, N2180, N425, N1339);
and AND4 (N4118, N4111, N1502, N3444, N2692);
and AND3 (N4119, N4109, N776, N512);
nand NAND3 (N4120, N4105, N3247, N2252);
buf BUF1 (N4121, N4114);
and AND3 (N4122, N4119, N3736, N1942);
and AND4 (N4123, N4116, N1842, N433, N2460);
or OR3 (N4124, N4117, N1841, N2429);
nor NOR2 (N4125, N4102, N449);
or OR4 (N4126, N4115, N4041, N3631, N2464);
or OR4 (N4127, N4122, N877, N2209, N3915);
and AND4 (N4128, N4123, N3324, N1954, N1126);
not NOT1 (N4129, N4126);
buf BUF1 (N4130, N4113);
or OR4 (N4131, N4125, N1694, N3146, N293);
or OR4 (N4132, N4129, N3705, N1368, N2002);
nand NAND2 (N4133, N4098, N2142);
or OR4 (N4134, N4118, N1333, N3203, N2982);
nor NOR3 (N4135, N4132, N2821, N146);
and AND3 (N4136, N4135, N4040, N1730);
nor NOR4 (N4137, N4121, N3547, N3457, N2446);
nor NOR2 (N4138, N4120, N5);
and AND2 (N4139, N4137, N1100);
or OR4 (N4140, N4124, N2127, N276, N3645);
not NOT1 (N4141, N4140);
nand NAND4 (N4142, N4139, N3720, N80, N522);
nand NAND2 (N4143, N4138, N3119);
buf BUF1 (N4144, N4143);
not NOT1 (N4145, N4142);
not NOT1 (N4146, N4131);
or OR3 (N4147, N4134, N2883, N2889);
buf BUF1 (N4148, N4127);
nor NOR2 (N4149, N4133, N1037);
nor NOR4 (N4150, N4145, N3764, N2217, N2778);
not NOT1 (N4151, N4149);
not NOT1 (N4152, N4141);
xor XOR2 (N4153, N4128, N1881);
not NOT1 (N4154, N4151);
xor XOR2 (N4155, N4146, N4128);
buf BUF1 (N4156, N4144);
not NOT1 (N4157, N4156);
xor XOR2 (N4158, N4154, N298);
nand NAND3 (N4159, N4147, N2993, N1825);
buf BUF1 (N4160, N4150);
and AND2 (N4161, N4152, N542);
or OR2 (N4162, N4161, N732);
buf BUF1 (N4163, N4153);
xor XOR2 (N4164, N4155, N3428);
nand NAND3 (N4165, N4148, N2035, N3741);
nor NOR4 (N4166, N4136, N2588, N1601, N2074);
nor NOR3 (N4167, N4130, N2079, N1539);
buf BUF1 (N4168, N4157);
buf BUF1 (N4169, N4163);
nand NAND4 (N4170, N4166, N4006, N585, N1162);
or OR2 (N4171, N4167, N26);
nand NAND2 (N4172, N4162, N1398);
xor XOR2 (N4173, N4168, N2992);
not NOT1 (N4174, N4170);
and AND4 (N4175, N4172, N1218, N3769, N3838);
xor XOR2 (N4176, N4173, N3661);
xor XOR2 (N4177, N4171, N2564);
nand NAND4 (N4178, N4159, N3539, N1921, N2954);
buf BUF1 (N4179, N4169);
xor XOR2 (N4180, N4179, N199);
nor NOR3 (N4181, N4175, N49, N2610);
nand NAND4 (N4182, N4165, N2527, N3725, N1923);
and AND4 (N4183, N4176, N1, N1431, N2531);
and AND4 (N4184, N4182, N21, N2468, N2988);
not NOT1 (N4185, N4177);
nor NOR3 (N4186, N4184, N1837, N291);
nand NAND2 (N4187, N4174, N888);
nand NAND3 (N4188, N4186, N1799, N3634);
not NOT1 (N4189, N4160);
xor XOR2 (N4190, N4187, N113);
and AND3 (N4191, N4188, N1275, N1665);
or OR2 (N4192, N4185, N2124);
and AND4 (N4193, N4164, N1826, N1325, N3452);
and AND4 (N4194, N4193, N775, N1559, N3365);
or OR2 (N4195, N4180, N1831);
xor XOR2 (N4196, N4158, N3588);
and AND2 (N4197, N4183, N273);
xor XOR2 (N4198, N4181, N883);
or OR2 (N4199, N4195, N4103);
nand NAND4 (N4200, N4194, N948, N1524, N1687);
nand NAND3 (N4201, N4189, N1192, N253);
not NOT1 (N4202, N4196);
nand NAND3 (N4203, N4178, N3127, N3321);
not NOT1 (N4204, N4190);
or OR4 (N4205, N4191, N2512, N3360, N63);
buf BUF1 (N4206, N4198);
or OR3 (N4207, N4202, N1456, N3881);
not NOT1 (N4208, N4205);
or OR3 (N4209, N4199, N498, N1125);
xor XOR2 (N4210, N4208, N2114);
and AND2 (N4211, N4206, N1504);
and AND3 (N4212, N4210, N3790, N1639);
not NOT1 (N4213, N4212);
and AND3 (N4214, N4204, N932, N1337);
not NOT1 (N4215, N4214);
nor NOR4 (N4216, N4207, N2916, N603, N195);
nor NOR3 (N4217, N4200, N3851, N700);
and AND4 (N4218, N4209, N3520, N431, N926);
buf BUF1 (N4219, N4218);
not NOT1 (N4220, N4203);
xor XOR2 (N4221, N4213, N2605);
not NOT1 (N4222, N4219);
or OR4 (N4223, N4215, N2871, N3880, N3426);
buf BUF1 (N4224, N4221);
nor NOR3 (N4225, N4216, N2315, N2533);
or OR2 (N4226, N4211, N1135);
not NOT1 (N4227, N4223);
not NOT1 (N4228, N4227);
not NOT1 (N4229, N4217);
or OR3 (N4230, N4225, N3473, N320);
buf BUF1 (N4231, N4192);
not NOT1 (N4232, N4220);
not NOT1 (N4233, N4201);
not NOT1 (N4234, N4229);
or OR2 (N4235, N4230, N1534);
not NOT1 (N4236, N4231);
buf BUF1 (N4237, N4228);
or OR3 (N4238, N4232, N3211, N3534);
nor NOR4 (N4239, N4234, N1011, N3928, N3695);
buf BUF1 (N4240, N4237);
buf BUF1 (N4241, N4238);
nor NOR2 (N4242, N4241, N1392);
not NOT1 (N4243, N4242);
buf BUF1 (N4244, N4236);
and AND2 (N4245, N4235, N2540);
and AND3 (N4246, N4244, N1385, N2685);
buf BUF1 (N4247, N4243);
xor XOR2 (N4248, N4222, N759);
not NOT1 (N4249, N4247);
and AND2 (N4250, N4245, N2405);
buf BUF1 (N4251, N4226);
or OR4 (N4252, N4224, N1049, N1339, N2789);
not NOT1 (N4253, N4249);
xor XOR2 (N4254, N4251, N797);
buf BUF1 (N4255, N4254);
xor XOR2 (N4256, N4239, N4232);
nor NOR3 (N4257, N4255, N886, N1314);
and AND3 (N4258, N4246, N1594, N344);
nand NAND2 (N4259, N4248, N2095);
xor XOR2 (N4260, N4259, N2344);
or OR3 (N4261, N4258, N1786, N3150);
xor XOR2 (N4262, N4252, N3085);
nand NAND2 (N4263, N4257, N3922);
nand NAND2 (N4264, N4240, N1628);
nor NOR2 (N4265, N4260, N3077);
nand NAND2 (N4266, N4233, N3703);
xor XOR2 (N4267, N4266, N3822);
nand NAND4 (N4268, N4265, N3322, N31, N3225);
and AND4 (N4269, N4268, N1544, N201, N2927);
nor NOR2 (N4270, N4197, N198);
nor NOR2 (N4271, N4269, N3828);
or OR2 (N4272, N4270, N3288);
nor NOR2 (N4273, N4263, N1763);
and AND4 (N4274, N4261, N3852, N1292, N2271);
nor NOR2 (N4275, N4267, N3320);
or OR4 (N4276, N4262, N1229, N1847, N3217);
xor XOR2 (N4277, N4256, N4077);
not NOT1 (N4278, N4264);
buf BUF1 (N4279, N4253);
and AND2 (N4280, N4278, N1929);
xor XOR2 (N4281, N4250, N2711);
or OR4 (N4282, N4271, N3811, N2010, N3480);
and AND4 (N4283, N4280, N1208, N370, N1311);
not NOT1 (N4284, N4275);
buf BUF1 (N4285, N4277);
buf BUF1 (N4286, N4272);
nor NOR2 (N4287, N4276, N2546);
buf BUF1 (N4288, N4284);
xor XOR2 (N4289, N4287, N3745);
or OR2 (N4290, N4286, N1427);
and AND2 (N4291, N4281, N3580);
not NOT1 (N4292, N4288);
buf BUF1 (N4293, N4279);
or OR3 (N4294, N4293, N899, N3522);
buf BUF1 (N4295, N4289);
nor NOR2 (N4296, N4274, N832);
buf BUF1 (N4297, N4292);
xor XOR2 (N4298, N4291, N1040);
nor NOR4 (N4299, N4273, N1739, N3810, N1279);
nor NOR2 (N4300, N4296, N3526);
xor XOR2 (N4301, N4297, N90);
nand NAND4 (N4302, N4299, N3707, N397, N3451);
buf BUF1 (N4303, N4282);
xor XOR2 (N4304, N4283, N938);
not NOT1 (N4305, N4303);
or OR3 (N4306, N4290, N1841, N3809);
and AND4 (N4307, N4302, N1498, N3265, N2611);
xor XOR2 (N4308, N4300, N3880);
nand NAND4 (N4309, N4305, N3682, N3321, N3069);
nor NOR3 (N4310, N4301, N1371, N3500);
nand NAND2 (N4311, N4294, N3816);
nand NAND3 (N4312, N4310, N3264, N705);
buf BUF1 (N4313, N4285);
and AND4 (N4314, N4304, N839, N3050, N3235);
not NOT1 (N4315, N4312);
buf BUF1 (N4316, N4307);
xor XOR2 (N4317, N4295, N2808);
buf BUF1 (N4318, N4311);
not NOT1 (N4319, N4306);
buf BUF1 (N4320, N4308);
xor XOR2 (N4321, N4320, N2163);
or OR2 (N4322, N4315, N1834);
nor NOR2 (N4323, N4313, N662);
and AND3 (N4324, N4317, N1660, N2248);
nor NOR4 (N4325, N4309, N413, N2363, N438);
and AND4 (N4326, N4321, N145, N1541, N1355);
and AND4 (N4327, N4326, N1711, N1945, N2159);
xor XOR2 (N4328, N4325, N2144);
or OR3 (N4329, N4319, N1260, N922);
nor NOR4 (N4330, N4314, N524, N3156, N1435);
buf BUF1 (N4331, N4324);
nand NAND3 (N4332, N4329, N1815, N923);
xor XOR2 (N4333, N4330, N241);
not NOT1 (N4334, N4298);
nand NAND3 (N4335, N4332, N3722, N3346);
or OR2 (N4336, N4318, N227);
nand NAND4 (N4337, N4336, N1854, N4027, N430);
buf BUF1 (N4338, N4323);
not NOT1 (N4339, N4331);
or OR2 (N4340, N4339, N3008);
buf BUF1 (N4341, N4337);
buf BUF1 (N4342, N4335);
xor XOR2 (N4343, N4340, N642);
nand NAND4 (N4344, N4334, N307, N2617, N4160);
buf BUF1 (N4345, N4333);
nor NOR2 (N4346, N4338, N476);
and AND4 (N4347, N4316, N2176, N1217, N539);
and AND2 (N4348, N4347, N535);
nor NOR2 (N4349, N4348, N729);
not NOT1 (N4350, N4342);
buf BUF1 (N4351, N4343);
nor NOR3 (N4352, N4322, N2796, N1511);
and AND3 (N4353, N4328, N3581, N1141);
and AND2 (N4354, N4345, N3643);
buf BUF1 (N4355, N4353);
or OR2 (N4356, N4351, N1419);
or OR3 (N4357, N4349, N1250, N2181);
buf BUF1 (N4358, N4327);
xor XOR2 (N4359, N4358, N2143);
nor NOR3 (N4360, N4341, N4270, N1791);
not NOT1 (N4361, N4350);
nor NOR2 (N4362, N4346, N1687);
buf BUF1 (N4363, N4357);
buf BUF1 (N4364, N4359);
xor XOR2 (N4365, N4344, N107);
nand NAND4 (N4366, N4354, N2547, N25, N4217);
not NOT1 (N4367, N4355);
nand NAND3 (N4368, N4367, N985, N2146);
and AND2 (N4369, N4362, N1598);
xor XOR2 (N4370, N4352, N335);
or OR3 (N4371, N4364, N4260, N1691);
nand NAND2 (N4372, N4363, N306);
buf BUF1 (N4373, N4368);
nor NOR2 (N4374, N4356, N3468);
buf BUF1 (N4375, N4374);
nor NOR3 (N4376, N4375, N3456, N1259);
or OR3 (N4377, N4376, N2639, N2680);
or OR2 (N4378, N4365, N2016);
nand NAND2 (N4379, N4366, N1611);
nand NAND3 (N4380, N4373, N1310, N2024);
nor NOR3 (N4381, N4380, N2281, N2084);
nor NOR2 (N4382, N4377, N3258);
or OR2 (N4383, N4360, N3698);
nor NOR3 (N4384, N4369, N1033, N3190);
or OR3 (N4385, N4370, N700, N2664);
or OR3 (N4386, N4381, N757, N3277);
not NOT1 (N4387, N4385);
nor NOR2 (N4388, N4372, N2309);
and AND3 (N4389, N4386, N258, N4323);
not NOT1 (N4390, N4383);
nand NAND3 (N4391, N4389, N2402, N4214);
not NOT1 (N4392, N4378);
nor NOR3 (N4393, N4387, N638, N3348);
xor XOR2 (N4394, N4391, N120);
or OR4 (N4395, N4388, N2922, N2451, N3127);
not NOT1 (N4396, N4382);
not NOT1 (N4397, N4392);
and AND3 (N4398, N4396, N2656, N1845);
xor XOR2 (N4399, N4371, N1126);
or OR2 (N4400, N4397, N4262);
buf BUF1 (N4401, N4400);
and AND2 (N4402, N4390, N299);
not NOT1 (N4403, N4394);
nand NAND3 (N4404, N4403, N3151, N215);
buf BUF1 (N4405, N4395);
nand NAND2 (N4406, N4404, N3247);
and AND4 (N4407, N4384, N1142, N55, N620);
xor XOR2 (N4408, N4406, N3939);
not NOT1 (N4409, N4408);
not NOT1 (N4410, N4361);
xor XOR2 (N4411, N4407, N1510);
buf BUF1 (N4412, N4411);
and AND2 (N4413, N4379, N1717);
buf BUF1 (N4414, N4398);
or OR3 (N4415, N4401, N2999, N2324);
xor XOR2 (N4416, N4413, N3021);
or OR2 (N4417, N4393, N1770);
xor XOR2 (N4418, N4409, N2718);
xor XOR2 (N4419, N4399, N2122);
xor XOR2 (N4420, N4419, N3235);
and AND3 (N4421, N4418, N998, N1935);
nor NOR4 (N4422, N4421, N2273, N1835, N4162);
or OR3 (N4423, N4405, N2884, N1139);
not NOT1 (N4424, N4417);
nor NOR3 (N4425, N4423, N1718, N613);
nor NOR3 (N4426, N4414, N404, N1079);
buf BUF1 (N4427, N4415);
xor XOR2 (N4428, N4420, N1774);
buf BUF1 (N4429, N4422);
not NOT1 (N4430, N4426);
and AND4 (N4431, N4410, N262, N480, N1841);
not NOT1 (N4432, N4425);
nor NOR2 (N4433, N4416, N2860);
buf BUF1 (N4434, N4433);
nor NOR4 (N4435, N4429, N1806, N606, N478);
and AND3 (N4436, N4434, N1478, N2637);
nand NAND2 (N4437, N4427, N3157);
xor XOR2 (N4438, N4424, N3307);
nand NAND2 (N4439, N4428, N450);
nand NAND2 (N4440, N4432, N3395);
and AND4 (N4441, N4438, N1429, N395, N16);
or OR4 (N4442, N4441, N1002, N3374, N1344);
nor NOR2 (N4443, N4431, N1745);
xor XOR2 (N4444, N4435, N2924);
buf BUF1 (N4445, N4436);
buf BUF1 (N4446, N4402);
xor XOR2 (N4447, N4443, N4308);
xor XOR2 (N4448, N4446, N2502);
xor XOR2 (N4449, N4430, N950);
not NOT1 (N4450, N4440);
xor XOR2 (N4451, N4439, N2456);
nor NOR3 (N4452, N4451, N4241, N1133);
not NOT1 (N4453, N4447);
nor NOR3 (N4454, N4450, N3559, N195);
buf BUF1 (N4455, N4412);
buf BUF1 (N4456, N4448);
nand NAND2 (N4457, N4449, N4452);
or OR4 (N4458, N4209, N1641, N2306, N2913);
buf BUF1 (N4459, N4444);
nand NAND4 (N4460, N4442, N3140, N137, N2931);
and AND3 (N4461, N4459, N1, N4368);
buf BUF1 (N4462, N4456);
and AND3 (N4463, N4454, N1294, N4317);
xor XOR2 (N4464, N4437, N2777);
not NOT1 (N4465, N4461);
or OR3 (N4466, N4460, N2045, N1435);
not NOT1 (N4467, N4466);
xor XOR2 (N4468, N4464, N1951);
or OR2 (N4469, N4445, N145);
and AND3 (N4470, N4469, N3196, N1964);
nor NOR2 (N4471, N4455, N1281);
nor NOR2 (N4472, N4467, N456);
buf BUF1 (N4473, N4453);
buf BUF1 (N4474, N4473);
or OR3 (N4475, N4465, N4474, N474);
xor XOR2 (N4476, N2889, N1630);
nor NOR2 (N4477, N4471, N1501);
buf BUF1 (N4478, N4476);
nor NOR3 (N4479, N4472, N1003, N1735);
nand NAND2 (N4480, N4475, N2304);
and AND3 (N4481, N4479, N430, N4473);
xor XOR2 (N4482, N4481, N2696);
xor XOR2 (N4483, N4482, N4374);
buf BUF1 (N4484, N4457);
or OR4 (N4485, N4483, N400, N3311, N208);
not NOT1 (N4486, N4478);
nor NOR3 (N4487, N4486, N3615, N1642);
nand NAND2 (N4488, N4468, N1272);
not NOT1 (N4489, N4463);
nand NAND3 (N4490, N4485, N2662, N3057);
or OR3 (N4491, N4480, N3657, N719);
or OR3 (N4492, N4488, N532, N2755);
nand NAND3 (N4493, N4490, N1096, N2064);
buf BUF1 (N4494, N4462);
or OR2 (N4495, N4458, N3367);
and AND3 (N4496, N4477, N2592, N525);
not NOT1 (N4497, N4489);
nor NOR4 (N4498, N4495, N1823, N940, N2019);
buf BUF1 (N4499, N4492);
and AND3 (N4500, N4499, N93, N1689);
not NOT1 (N4501, N4496);
or OR4 (N4502, N4501, N101, N666, N3670);
xor XOR2 (N4503, N4497, N1297);
or OR3 (N4504, N4500, N3560, N1352);
not NOT1 (N4505, N4504);
nor NOR2 (N4506, N4503, N3020);
and AND3 (N4507, N4487, N988, N2629);
and AND3 (N4508, N4491, N1565, N994);
or OR4 (N4509, N4507, N2225, N2920, N2557);
nand NAND4 (N4510, N4470, N1847, N4073, N4323);
nand NAND2 (N4511, N4494, N3302);
not NOT1 (N4512, N4505);
xor XOR2 (N4513, N4512, N4420);
nand NAND2 (N4514, N4484, N4329);
or OR2 (N4515, N4511, N3503);
nand NAND2 (N4516, N4508, N2088);
xor XOR2 (N4517, N4509, N1983);
nor NOR3 (N4518, N4510, N1519, N3434);
nand NAND4 (N4519, N4493, N3557, N2819, N1596);
and AND2 (N4520, N4518, N4129);
buf BUF1 (N4521, N4520);
nor NOR2 (N4522, N4521, N558);
not NOT1 (N4523, N4515);
nor NOR4 (N4524, N4513, N1484, N1731, N4210);
or OR4 (N4525, N4517, N987, N1369, N3336);
and AND2 (N4526, N4522, N1866);
and AND3 (N4527, N4524, N2652, N1859);
buf BUF1 (N4528, N4525);
not NOT1 (N4529, N4506);
not NOT1 (N4530, N4502);
xor XOR2 (N4531, N4529, N336);
nor NOR2 (N4532, N4514, N1820);
or OR2 (N4533, N4523, N1130);
buf BUF1 (N4534, N4533);
not NOT1 (N4535, N4530);
xor XOR2 (N4536, N4516, N14);
nor NOR2 (N4537, N4531, N4471);
not NOT1 (N4538, N4534);
or OR4 (N4539, N4498, N2754, N2901, N424);
and AND2 (N4540, N4539, N2228);
or OR4 (N4541, N4535, N2752, N11, N2356);
buf BUF1 (N4542, N4532);
xor XOR2 (N4543, N4542, N3706);
xor XOR2 (N4544, N4541, N4025);
and AND2 (N4545, N4519, N2622);
xor XOR2 (N4546, N4540, N2210);
not NOT1 (N4547, N4537);
nand NAND3 (N4548, N4527, N20, N3569);
or OR4 (N4549, N4547, N2253, N1174, N2340);
nor NOR4 (N4550, N4538, N555, N3948, N824);
and AND4 (N4551, N4545, N547, N2829, N2592);
buf BUF1 (N4552, N4543);
or OR2 (N4553, N4544, N2293);
buf BUF1 (N4554, N4536);
nor NOR2 (N4555, N4548, N3952);
nor NOR4 (N4556, N4553, N1425, N2611, N565);
or OR3 (N4557, N4552, N1208, N2909);
not NOT1 (N4558, N4550);
not NOT1 (N4559, N4551);
or OR3 (N4560, N4528, N461, N2424);
nand NAND3 (N4561, N4549, N2829, N1547);
nand NAND4 (N4562, N4554, N3181, N3406, N1350);
or OR2 (N4563, N4555, N3962);
not NOT1 (N4564, N4562);
not NOT1 (N4565, N4560);
and AND3 (N4566, N4559, N4302, N1904);
buf BUF1 (N4567, N4546);
not NOT1 (N4568, N4561);
not NOT1 (N4569, N4565);
not NOT1 (N4570, N4526);
not NOT1 (N4571, N4564);
nor NOR4 (N4572, N4567, N2979, N3770, N3887);
buf BUF1 (N4573, N4572);
not NOT1 (N4574, N4557);
not NOT1 (N4575, N4563);
and AND2 (N4576, N4566, N3600);
buf BUF1 (N4577, N4570);
and AND2 (N4578, N4558, N3059);
not NOT1 (N4579, N4571);
nand NAND2 (N4580, N4577, N3528);
and AND4 (N4581, N4573, N3391, N3315, N939);
or OR2 (N4582, N4574, N1573);
xor XOR2 (N4583, N4576, N534);
or OR2 (N4584, N4569, N1188);
xor XOR2 (N4585, N4583, N1339);
not NOT1 (N4586, N4580);
nand NAND4 (N4587, N4582, N2484, N2015, N2200);
or OR2 (N4588, N4586, N1852);
not NOT1 (N4589, N4584);
or OR4 (N4590, N4568, N1175, N2269, N816);
or OR3 (N4591, N4590, N3518, N3468);
not NOT1 (N4592, N4581);
xor XOR2 (N4593, N4575, N4061);
nor NOR4 (N4594, N4585, N3734, N1310, N2726);
and AND4 (N4595, N4588, N580, N764, N2489);
or OR2 (N4596, N4587, N3059);
not NOT1 (N4597, N4596);
nand NAND3 (N4598, N4556, N3332, N1629);
buf BUF1 (N4599, N4594);
nor NOR4 (N4600, N4598, N2595, N223, N4060);
and AND4 (N4601, N4589, N364, N2673, N2406);
xor XOR2 (N4602, N4599, N15);
and AND4 (N4603, N4602, N2892, N11, N4482);
or OR3 (N4604, N4579, N1119, N623);
xor XOR2 (N4605, N4595, N265);
nand NAND4 (N4606, N4591, N1781, N2768, N4248);
not NOT1 (N4607, N4597);
nand NAND4 (N4608, N4603, N2815, N3480, N191);
or OR3 (N4609, N4578, N3859, N1858);
or OR3 (N4610, N4600, N254, N1997);
or OR4 (N4611, N4605, N621, N1116, N33);
or OR2 (N4612, N4610, N752);
not NOT1 (N4613, N4606);
nand NAND2 (N4614, N4604, N3770);
xor XOR2 (N4615, N4613, N3450);
or OR4 (N4616, N4614, N203, N4223, N2660);
xor XOR2 (N4617, N4612, N3296);
and AND2 (N4618, N4617, N2571);
buf BUF1 (N4619, N4601);
and AND2 (N4620, N4619, N1618);
not NOT1 (N4621, N4618);
and AND3 (N4622, N4608, N1806, N3495);
not NOT1 (N4623, N4620);
buf BUF1 (N4624, N4607);
and AND2 (N4625, N4615, N119);
nand NAND2 (N4626, N4623, N2951);
not NOT1 (N4627, N4621);
buf BUF1 (N4628, N4611);
and AND2 (N4629, N4624, N1423);
and AND4 (N4630, N4616, N631, N309, N503);
xor XOR2 (N4631, N4629, N427);
or OR3 (N4632, N4626, N3415, N1335);
and AND4 (N4633, N4627, N1062, N1308, N3708);
buf BUF1 (N4634, N4631);
or OR2 (N4635, N4593, N1665);
xor XOR2 (N4636, N4625, N3023);
xor XOR2 (N4637, N4609, N1019);
buf BUF1 (N4638, N4622);
and AND2 (N4639, N4638, N2667);
buf BUF1 (N4640, N4634);
nand NAND3 (N4641, N4592, N2793, N329);
or OR2 (N4642, N4641, N2640);
nand NAND4 (N4643, N4637, N1409, N2867, N181);
nand NAND2 (N4644, N4635, N3428);
xor XOR2 (N4645, N4632, N464);
or OR3 (N4646, N4639, N1432, N2022);
and AND4 (N4647, N4644, N3509, N886, N706);
nand NAND2 (N4648, N4645, N431);
and AND2 (N4649, N4630, N1864);
nand NAND2 (N4650, N4642, N2593);
and AND2 (N4651, N4650, N3126);
or OR4 (N4652, N4647, N66, N1179, N3616);
xor XOR2 (N4653, N4648, N2988);
xor XOR2 (N4654, N4628, N4598);
not NOT1 (N4655, N4654);
nand NAND3 (N4656, N4649, N3850, N1672);
not NOT1 (N4657, N4653);
nand NAND3 (N4658, N4656, N3254, N1370);
nand NAND2 (N4659, N4633, N542);
nor NOR3 (N4660, N4646, N3660, N3556);
and AND2 (N4661, N4659, N2024);
not NOT1 (N4662, N4660);
xor XOR2 (N4663, N4643, N391);
buf BUF1 (N4664, N4661);
xor XOR2 (N4665, N4664, N4442);
xor XOR2 (N4666, N4665, N400);
buf BUF1 (N4667, N4658);
xor XOR2 (N4668, N4663, N4094);
nor NOR3 (N4669, N4662, N83, N3097);
buf BUF1 (N4670, N4651);
nand NAND2 (N4671, N4636, N2290);
or OR4 (N4672, N4669, N2212, N562, N1272);
nand NAND4 (N4673, N4652, N4546, N398, N932);
and AND3 (N4674, N4668, N4657, N3942);
nor NOR2 (N4675, N1710, N3846);
xor XOR2 (N4676, N4671, N2421);
xor XOR2 (N4677, N4655, N2628);
or OR2 (N4678, N4676, N1429);
buf BUF1 (N4679, N4670);
nand NAND2 (N4680, N4678, N2537);
not NOT1 (N4681, N4672);
buf BUF1 (N4682, N4675);
buf BUF1 (N4683, N4667);
buf BUF1 (N4684, N4680);
buf BUF1 (N4685, N4684);
or OR3 (N4686, N4674, N2765, N3334);
nor NOR2 (N4687, N4681, N4341);
nor NOR3 (N4688, N4685, N4125, N3851);
nand NAND4 (N4689, N4687, N1620, N3075, N3055);
and AND3 (N4690, N4673, N3338, N2950);
or OR3 (N4691, N4686, N2103, N597);
not NOT1 (N4692, N4677);
xor XOR2 (N4693, N4691, N1915);
buf BUF1 (N4694, N4688);
buf BUF1 (N4695, N4693);
or OR3 (N4696, N4692, N4425, N4344);
not NOT1 (N4697, N4696);
or OR3 (N4698, N4640, N1786, N1072);
or OR3 (N4699, N4689, N4000, N2786);
buf BUF1 (N4700, N4666);
nand NAND4 (N4701, N4698, N1178, N4187, N2094);
buf BUF1 (N4702, N4690);
buf BUF1 (N4703, N4702);
or OR4 (N4704, N4700, N2731, N2700, N362);
nand NAND3 (N4705, N4701, N272, N705);
nor NOR2 (N4706, N4682, N3364);
nand NAND2 (N4707, N4695, N2064);
or OR4 (N4708, N4699, N2204, N1655, N1509);
and AND3 (N4709, N4683, N291, N3148);
or OR3 (N4710, N4697, N3709, N2078);
or OR3 (N4711, N4703, N3353, N1759);
not NOT1 (N4712, N4707);
not NOT1 (N4713, N4679);
xor XOR2 (N4714, N4713, N3502);
not NOT1 (N4715, N4710);
or OR4 (N4716, N4704, N766, N1339, N3400);
nor NOR2 (N4717, N4711, N2387);
or OR2 (N4718, N4705, N772);
xor XOR2 (N4719, N4716, N4389);
not NOT1 (N4720, N4706);
not NOT1 (N4721, N4718);
nor NOR4 (N4722, N4694, N2996, N3943, N1961);
nand NAND2 (N4723, N4717, N2684);
and AND3 (N4724, N4722, N590, N882);
not NOT1 (N4725, N4724);
buf BUF1 (N4726, N4709);
or OR4 (N4727, N4708, N453, N3186, N4346);
and AND4 (N4728, N4721, N2609, N1543, N765);
nand NAND2 (N4729, N4715, N4434);
nand NAND3 (N4730, N4714, N2053, N4645);
or OR4 (N4731, N4726, N489, N3039, N3450);
nor NOR2 (N4732, N4725, N215);
buf BUF1 (N4733, N4728);
or OR2 (N4734, N4730, N2279);
or OR4 (N4735, N4732, N2589, N1540, N2994);
nor NOR3 (N4736, N4727, N3815, N3611);
xor XOR2 (N4737, N4720, N4631);
nor NOR3 (N4738, N4734, N3506, N1900);
buf BUF1 (N4739, N4731);
xor XOR2 (N4740, N4736, N3907);
buf BUF1 (N4741, N4733);
xor XOR2 (N4742, N4712, N4713);
not NOT1 (N4743, N4741);
nand NAND3 (N4744, N4737, N799, N826);
buf BUF1 (N4745, N4743);
nor NOR3 (N4746, N4729, N2678, N1496);
not NOT1 (N4747, N4745);
buf BUF1 (N4748, N4742);
buf BUF1 (N4749, N4744);
or OR4 (N4750, N4735, N908, N4239, N3301);
not NOT1 (N4751, N4749);
nand NAND2 (N4752, N4719, N1995);
buf BUF1 (N4753, N4751);
xor XOR2 (N4754, N4750, N4557);
xor XOR2 (N4755, N4747, N3258);
xor XOR2 (N4756, N4753, N3763);
xor XOR2 (N4757, N4738, N1332);
buf BUF1 (N4758, N4757);
buf BUF1 (N4759, N4723);
buf BUF1 (N4760, N4759);
not NOT1 (N4761, N4755);
buf BUF1 (N4762, N4754);
and AND4 (N4763, N4762, N130, N2855, N3482);
or OR3 (N4764, N4748, N3000, N2245);
buf BUF1 (N4765, N4756);
buf BUF1 (N4766, N4746);
or OR3 (N4767, N4739, N2109, N2024);
buf BUF1 (N4768, N4764);
xor XOR2 (N4769, N4761, N3236);
nand NAND2 (N4770, N4767, N656);
nand NAND3 (N4771, N4752, N2961, N1509);
buf BUF1 (N4772, N4763);
buf BUF1 (N4773, N4772);
and AND4 (N4774, N4758, N2039, N3408, N2886);
buf BUF1 (N4775, N4770);
buf BUF1 (N4776, N4774);
nor NOR3 (N4777, N4766, N2698, N3489);
xor XOR2 (N4778, N4740, N2159);
or OR3 (N4779, N4768, N684, N4686);
nor NOR2 (N4780, N4760, N3082);
not NOT1 (N4781, N4771);
xor XOR2 (N4782, N4779, N1143);
nor NOR2 (N4783, N4778, N534);
not NOT1 (N4784, N4782);
and AND4 (N4785, N4781, N147, N2073, N1160);
xor XOR2 (N4786, N4765, N362);
nand NAND4 (N4787, N4777, N3978, N3939, N568);
not NOT1 (N4788, N4776);
xor XOR2 (N4789, N4787, N312);
buf BUF1 (N4790, N4775);
nand NAND3 (N4791, N4790, N3680, N3163);
xor XOR2 (N4792, N4791, N3654);
not NOT1 (N4793, N4769);
and AND3 (N4794, N4783, N4469, N3756);
and AND2 (N4795, N4788, N1047);
not NOT1 (N4796, N4792);
not NOT1 (N4797, N4785);
nor NOR4 (N4798, N4773, N1005, N4520, N974);
and AND2 (N4799, N4784, N2703);
buf BUF1 (N4800, N4793);
or OR4 (N4801, N4799, N631, N331, N1296);
or OR3 (N4802, N4798, N4072, N2916);
buf BUF1 (N4803, N4802);
nor NOR3 (N4804, N4803, N2545, N2727);
or OR2 (N4805, N4801, N3259);
and AND4 (N4806, N4789, N1951, N1216, N72);
nand NAND2 (N4807, N4806, N3995);
nor NOR4 (N4808, N4794, N881, N1700, N4254);
or OR2 (N4809, N4800, N4394);
nor NOR3 (N4810, N4796, N325, N3302);
nor NOR3 (N4811, N4797, N3664, N1459);
nand NAND2 (N4812, N4811, N3059);
buf BUF1 (N4813, N4809);
not NOT1 (N4814, N4795);
or OR4 (N4815, N4814, N2620, N3437, N2603);
xor XOR2 (N4816, N4812, N3889);
nand NAND4 (N4817, N4780, N267, N3920, N598);
nand NAND2 (N4818, N4813, N1874);
nor NOR3 (N4819, N4808, N3138, N1325);
and AND3 (N4820, N4805, N1746, N2945);
or OR4 (N4821, N4804, N3691, N215, N3145);
nor NOR2 (N4822, N4818, N144);
buf BUF1 (N4823, N4815);
nand NAND3 (N4824, N4821, N778, N2099);
or OR4 (N4825, N4819, N1656, N2584, N148);
buf BUF1 (N4826, N4824);
and AND2 (N4827, N4816, N428);
xor XOR2 (N4828, N4786, N2130);
xor XOR2 (N4829, N4828, N3162);
and AND2 (N4830, N4829, N1065);
buf BUF1 (N4831, N4826);
buf BUF1 (N4832, N4817);
and AND3 (N4833, N4825, N1448, N3431);
buf BUF1 (N4834, N4827);
nor NOR2 (N4835, N4831, N3832);
or OR2 (N4836, N4835, N1201);
or OR3 (N4837, N4832, N4226, N1326);
nand NAND2 (N4838, N4834, N1124);
nor NOR2 (N4839, N4836, N1716);
and AND2 (N4840, N4830, N2690);
nor NOR3 (N4841, N4838, N3424, N8);
nor NOR2 (N4842, N4833, N1964);
or OR3 (N4843, N4822, N4, N2375);
not NOT1 (N4844, N4843);
buf BUF1 (N4845, N4840);
not NOT1 (N4846, N4839);
nand NAND3 (N4847, N4823, N3978, N64);
and AND4 (N4848, N4820, N24, N1844, N4453);
nor NOR3 (N4849, N4844, N4825, N1825);
not NOT1 (N4850, N4807);
or OR2 (N4851, N4842, N2000);
not NOT1 (N4852, N4837);
nand NAND2 (N4853, N4847, N1988);
nor NOR3 (N4854, N4841, N1398, N973);
nor NOR2 (N4855, N4854, N819);
xor XOR2 (N4856, N4851, N2538);
xor XOR2 (N4857, N4855, N956);
buf BUF1 (N4858, N4857);
or OR3 (N4859, N4856, N2036, N2331);
not NOT1 (N4860, N4853);
nand NAND3 (N4861, N4860, N226, N566);
buf BUF1 (N4862, N4810);
xor XOR2 (N4863, N4848, N1678);
and AND2 (N4864, N4852, N4001);
nor NOR2 (N4865, N4845, N1567);
nor NOR4 (N4866, N4849, N3150, N3873, N624);
xor XOR2 (N4867, N4863, N2685);
buf BUF1 (N4868, N4850);
or OR2 (N4869, N4862, N1143);
buf BUF1 (N4870, N4866);
nand NAND2 (N4871, N4870, N985);
nand NAND2 (N4872, N4865, N3522);
buf BUF1 (N4873, N4868);
not NOT1 (N4874, N4867);
and AND2 (N4875, N4858, N1678);
nor NOR3 (N4876, N4869, N3157, N3224);
nand NAND4 (N4877, N4859, N3823, N1790, N1903);
xor XOR2 (N4878, N4876, N3678);
and AND4 (N4879, N4872, N148, N4486, N1912);
and AND4 (N4880, N4879, N151, N2786, N1643);
nand NAND2 (N4881, N4874, N2955);
and AND2 (N4882, N4873, N4627);
nand NAND3 (N4883, N4881, N1081, N4834);
xor XOR2 (N4884, N4878, N4086);
and AND3 (N4885, N4882, N1522, N136);
xor XOR2 (N4886, N4885, N2823);
not NOT1 (N4887, N4846);
and AND2 (N4888, N4877, N3525);
xor XOR2 (N4889, N4887, N472);
xor XOR2 (N4890, N4888, N3619);
or OR3 (N4891, N4861, N3151, N3881);
xor XOR2 (N4892, N4884, N1645);
or OR3 (N4893, N4875, N1586, N3954);
or OR3 (N4894, N4892, N2946, N4172);
buf BUF1 (N4895, N4889);
buf BUF1 (N4896, N4890);
nand NAND2 (N4897, N4891, N3015);
nor NOR2 (N4898, N4897, N2989);
and AND2 (N4899, N4893, N41);
not NOT1 (N4900, N4864);
nor NOR4 (N4901, N4899, N4518, N412, N4844);
not NOT1 (N4902, N4900);
not NOT1 (N4903, N4895);
buf BUF1 (N4904, N4886);
not NOT1 (N4905, N4883);
and AND2 (N4906, N4901, N3160);
or OR4 (N4907, N4896, N939, N4207, N2427);
not NOT1 (N4908, N4906);
and AND2 (N4909, N4905, N945);
or OR4 (N4910, N4880, N1061, N3891, N4156);
xor XOR2 (N4911, N4908, N696);
not NOT1 (N4912, N4871);
nor NOR4 (N4913, N4894, N3345, N3768, N4316);
nand NAND2 (N4914, N4903, N3161);
and AND3 (N4915, N4898, N3477, N126);
xor XOR2 (N4916, N4913, N817);
buf BUF1 (N4917, N4916);
buf BUF1 (N4918, N4902);
nand NAND3 (N4919, N4910, N4727, N3123);
buf BUF1 (N4920, N4904);
nand NAND2 (N4921, N4917, N3856);
or OR3 (N4922, N4915, N4047, N104);
or OR3 (N4923, N4919, N2306, N2705);
and AND2 (N4924, N4912, N1863);
buf BUF1 (N4925, N4920);
xor XOR2 (N4926, N4907, N4490);
nor NOR2 (N4927, N4925, N4682);
or OR2 (N4928, N4918, N4792);
buf BUF1 (N4929, N4923);
buf BUF1 (N4930, N4928);
or OR4 (N4931, N4927, N2867, N239, N281);
xor XOR2 (N4932, N4931, N1169);
nor NOR4 (N4933, N4922, N3990, N2627, N2583);
and AND3 (N4934, N4933, N4269, N787);
buf BUF1 (N4935, N4932);
nor NOR4 (N4936, N4930, N1752, N1053, N2955);
nor NOR3 (N4937, N4935, N2382, N255);
buf BUF1 (N4938, N4936);
not NOT1 (N4939, N4924);
xor XOR2 (N4940, N4929, N2207);
buf BUF1 (N4941, N4909);
and AND2 (N4942, N4937, N3147);
nor NOR2 (N4943, N4941, N849);
not NOT1 (N4944, N4934);
nor NOR4 (N4945, N4939, N3483, N2333, N1193);
xor XOR2 (N4946, N4943, N110);
buf BUF1 (N4947, N4942);
xor XOR2 (N4948, N4946, N4501);
nor NOR2 (N4949, N4945, N3746);
buf BUF1 (N4950, N4938);
buf BUF1 (N4951, N4914);
not NOT1 (N4952, N4940);
not NOT1 (N4953, N4926);
nor NOR3 (N4954, N4944, N2944, N2919);
and AND2 (N4955, N4951, N4536);
and AND3 (N4956, N4950, N1991, N396);
or OR4 (N4957, N4956, N1280, N2228, N2267);
not NOT1 (N4958, N4921);
nand NAND3 (N4959, N4948, N4404, N3025);
nand NAND4 (N4960, N4957, N4592, N3641, N3376);
nand NAND2 (N4961, N4954, N1640);
and AND2 (N4962, N4952, N904);
buf BUF1 (N4963, N4958);
and AND3 (N4964, N4953, N408, N76);
not NOT1 (N4965, N4949);
nand NAND2 (N4966, N4911, N1404);
and AND2 (N4967, N4960, N4185);
not NOT1 (N4968, N4947);
nor NOR3 (N4969, N4966, N3223, N4258);
and AND2 (N4970, N4955, N1017);
not NOT1 (N4971, N4968);
or OR2 (N4972, N4969, N3012);
buf BUF1 (N4973, N4972);
or OR2 (N4974, N4967, N842);
nand NAND2 (N4975, N4974, N3722);
buf BUF1 (N4976, N4975);
and AND3 (N4977, N4961, N3421, N3386);
or OR4 (N4978, N4976, N1613, N4118, N2448);
not NOT1 (N4979, N4962);
nor NOR2 (N4980, N4977, N229);
not NOT1 (N4981, N4963);
nor NOR3 (N4982, N4971, N31, N4471);
xor XOR2 (N4983, N4979, N3838);
xor XOR2 (N4984, N4959, N1090);
or OR4 (N4985, N4981, N918, N204, N3698);
and AND2 (N4986, N4980, N2787);
nand NAND3 (N4987, N4982, N738, N4645);
buf BUF1 (N4988, N4970);
or OR3 (N4989, N4983, N2377, N3328);
buf BUF1 (N4990, N4964);
nand NAND4 (N4991, N4985, N3620, N2247, N4910);
and AND2 (N4992, N4989, N2067);
not NOT1 (N4993, N4992);
xor XOR2 (N4994, N4978, N2847);
nand NAND2 (N4995, N4965, N2492);
not NOT1 (N4996, N4993);
not NOT1 (N4997, N4995);
or OR4 (N4998, N4988, N2028, N4351, N3068);
nand NAND2 (N4999, N4984, N1551);
buf BUF1 (N5000, N4991);
nor NOR4 (N5001, N4999, N4692, N1474, N2498);
buf BUF1 (N5002, N4997);
not NOT1 (N5003, N4998);
nor NOR4 (N5004, N4996, N4547, N3421, N3805);
not NOT1 (N5005, N4987);
nor NOR2 (N5006, N4994, N3969);
nand NAND4 (N5007, N5000, N1208, N4345, N4819);
nor NOR4 (N5008, N5006, N2464, N2571, N1267);
xor XOR2 (N5009, N5004, N3007);
nand NAND4 (N5010, N5007, N1399, N2015, N3456);
buf BUF1 (N5011, N5001);
buf BUF1 (N5012, N5010);
nor NOR2 (N5013, N5011, N1072);
xor XOR2 (N5014, N5012, N3322);
not NOT1 (N5015, N4986);
xor XOR2 (N5016, N5014, N4221);
nor NOR3 (N5017, N5003, N1697, N4322);
nor NOR3 (N5018, N5013, N2287, N4155);
and AND2 (N5019, N4973, N3503);
buf BUF1 (N5020, N5019);
buf BUF1 (N5021, N5009);
buf BUF1 (N5022, N5016);
and AND2 (N5023, N5015, N4645);
nor NOR3 (N5024, N5005, N4403, N822);
not NOT1 (N5025, N5020);
nand NAND4 (N5026, N5018, N4775, N414, N2835);
buf BUF1 (N5027, N5021);
not NOT1 (N5028, N5027);
buf BUF1 (N5029, N5024);
not NOT1 (N5030, N5017);
not NOT1 (N5031, N5023);
and AND3 (N5032, N5025, N2277, N4033);
xor XOR2 (N5033, N5022, N2968);
and AND3 (N5034, N5032, N3639, N3328);
xor XOR2 (N5035, N5030, N4211);
and AND4 (N5036, N5029, N2383, N1802, N169);
xor XOR2 (N5037, N5002, N4412);
nand NAND3 (N5038, N5034, N445, N904);
xor XOR2 (N5039, N4990, N845);
nand NAND4 (N5040, N5026, N1602, N3376, N3407);
or OR2 (N5041, N5039, N3524);
or OR4 (N5042, N5033, N650, N4372, N2281);
buf BUF1 (N5043, N5036);
and AND2 (N5044, N5038, N1347);
nor NOR4 (N5045, N5042, N124, N417, N4399);
xor XOR2 (N5046, N5031, N1311);
buf BUF1 (N5047, N5008);
buf BUF1 (N5048, N5047);
buf BUF1 (N5049, N5037);
and AND3 (N5050, N5044, N3725, N3077);
nand NAND2 (N5051, N5050, N4731);
nand NAND4 (N5052, N5041, N2481, N3291, N4647);
not NOT1 (N5053, N5043);
buf BUF1 (N5054, N5035);
and AND2 (N5055, N5040, N1055);
buf BUF1 (N5056, N5054);
buf BUF1 (N5057, N5045);
not NOT1 (N5058, N5053);
or OR2 (N5059, N5049, N106);
nor NOR3 (N5060, N5058, N31, N811);
buf BUF1 (N5061, N5046);
not NOT1 (N5062, N5056);
or OR4 (N5063, N5048, N4320, N516, N1020);
xor XOR2 (N5064, N5057, N1511);
xor XOR2 (N5065, N5062, N4595);
xor XOR2 (N5066, N5051, N4383);
nand NAND4 (N5067, N5065, N4514, N3434, N5066);
and AND3 (N5068, N4067, N3188, N4998);
or OR2 (N5069, N5067, N4001);
xor XOR2 (N5070, N5059, N195);
and AND4 (N5071, N5068, N1911, N2334, N1474);
xor XOR2 (N5072, N5061, N3172);
and AND4 (N5073, N5072, N4544, N1685, N4772);
not NOT1 (N5074, N5060);
or OR4 (N5075, N5070, N1168, N3739, N3470);
xor XOR2 (N5076, N5052, N3305);
not NOT1 (N5077, N5055);
and AND2 (N5078, N5028, N1624);
nand NAND3 (N5079, N5078, N148, N2614);
or OR3 (N5080, N5076, N3939, N877);
nor NOR2 (N5081, N5074, N3281);
buf BUF1 (N5082, N5079);
buf BUF1 (N5083, N5081);
nor NOR3 (N5084, N5077, N3346, N1389);
buf BUF1 (N5085, N5082);
not NOT1 (N5086, N5071);
or OR4 (N5087, N5063, N2493, N870, N3178);
or OR2 (N5088, N5064, N3092);
buf BUF1 (N5089, N5087);
not NOT1 (N5090, N5085);
or OR4 (N5091, N5069, N2616, N4227, N2513);
or OR4 (N5092, N5090, N1962, N2243, N2236);
nand NAND2 (N5093, N5073, N4139);
buf BUF1 (N5094, N5091);
or OR3 (N5095, N5089, N3885, N1229);
and AND3 (N5096, N5080, N3645, N122);
nand NAND4 (N5097, N5094, N1356, N4839, N2564);
buf BUF1 (N5098, N5075);
and AND2 (N5099, N5088, N458);
and AND2 (N5100, N5093, N2387);
nor NOR3 (N5101, N5092, N4945, N1094);
not NOT1 (N5102, N5099);
or OR2 (N5103, N5101, N1828);
nand NAND2 (N5104, N5084, N2819);
xor XOR2 (N5105, N5102, N2560);
or OR3 (N5106, N5100, N1112, N2866);
and AND4 (N5107, N5104, N1374, N1758, N599);
or OR4 (N5108, N5103, N76, N1260, N4871);
not NOT1 (N5109, N5086);
xor XOR2 (N5110, N5105, N2701);
nor NOR3 (N5111, N5096, N2650, N3617);
xor XOR2 (N5112, N5098, N2133);
buf BUF1 (N5113, N5083);
or OR4 (N5114, N5110, N2304, N3313, N4556);
xor XOR2 (N5115, N5107, N4719);
not NOT1 (N5116, N5112);
buf BUF1 (N5117, N5114);
buf BUF1 (N5118, N5097);
xor XOR2 (N5119, N5109, N3625);
xor XOR2 (N5120, N5111, N4918);
xor XOR2 (N5121, N5118, N3902);
or OR3 (N5122, N5106, N784, N617);
not NOT1 (N5123, N5095);
nand NAND2 (N5124, N5123, N408);
and AND4 (N5125, N5122, N5055, N1171, N1456);
or OR4 (N5126, N5120, N1769, N4919, N673);
nor NOR3 (N5127, N5121, N478, N1497);
and AND3 (N5128, N5108, N1266, N3267);
nor NOR3 (N5129, N5127, N2304, N2755);
nor NOR2 (N5130, N5125, N1433);
nor NOR4 (N5131, N5130, N825, N942, N2263);
xor XOR2 (N5132, N5116, N793);
or OR2 (N5133, N5117, N4252);
nor NOR3 (N5134, N5131, N4343, N3636);
and AND4 (N5135, N5124, N5032, N1050, N1762);
buf BUF1 (N5136, N5119);
or OR3 (N5137, N5133, N815, N83);
and AND4 (N5138, N5115, N4842, N2632, N639);
xor XOR2 (N5139, N5129, N2809);
xor XOR2 (N5140, N5137, N4341);
not NOT1 (N5141, N5138);
or OR4 (N5142, N5126, N4888, N2250, N2062);
and AND2 (N5143, N5136, N159);
not NOT1 (N5144, N5139);
xor XOR2 (N5145, N5144, N3236);
nand NAND4 (N5146, N5135, N3004, N2729, N2714);
nand NAND4 (N5147, N5128, N3977, N1256, N3912);
and AND4 (N5148, N5142, N4064, N336, N4712);
nand NAND3 (N5149, N5145, N4237, N5073);
nor NOR3 (N5150, N5148, N2793, N1515);
nor NOR2 (N5151, N5132, N3410);
or OR2 (N5152, N5150, N1995);
buf BUF1 (N5153, N5151);
xor XOR2 (N5154, N5152, N4454);
nor NOR4 (N5155, N5143, N245, N2274, N1507);
buf BUF1 (N5156, N5155);
buf BUF1 (N5157, N5156);
nand NAND3 (N5158, N5146, N1825, N3749);
nor NOR4 (N5159, N5141, N1171, N3261, N4983);
and AND2 (N5160, N5154, N1185);
and AND3 (N5161, N5140, N971, N247);
xor XOR2 (N5162, N5160, N1941);
nor NOR2 (N5163, N5113, N1847);
not NOT1 (N5164, N5162);
not NOT1 (N5165, N5159);
buf BUF1 (N5166, N5134);
buf BUF1 (N5167, N5163);
xor XOR2 (N5168, N5166, N641);
nand NAND2 (N5169, N5167, N1752);
and AND2 (N5170, N5153, N2695);
not NOT1 (N5171, N5161);
nand NAND4 (N5172, N5171, N1162, N1466, N1164);
not NOT1 (N5173, N5165);
buf BUF1 (N5174, N5164);
buf BUF1 (N5175, N5149);
nor NOR3 (N5176, N5175, N4148, N226);
not NOT1 (N5177, N5158);
and AND4 (N5178, N5174, N553, N3538, N2965);
nand NAND2 (N5179, N5157, N37);
xor XOR2 (N5180, N5170, N1152);
nand NAND3 (N5181, N5176, N2815, N5169);
not NOT1 (N5182, N1798);
or OR2 (N5183, N5182, N46);
or OR4 (N5184, N5178, N4673, N2537, N3731);
nand NAND3 (N5185, N5181, N4934, N331);
or OR2 (N5186, N5173, N2096);
xor XOR2 (N5187, N5168, N920);
xor XOR2 (N5188, N5180, N200);
not NOT1 (N5189, N5184);
buf BUF1 (N5190, N5186);
not NOT1 (N5191, N5147);
buf BUF1 (N5192, N5189);
nor NOR3 (N5193, N5179, N2190, N4170);
nor NOR2 (N5194, N5185, N4587);
buf BUF1 (N5195, N5194);
buf BUF1 (N5196, N5172);
or OR3 (N5197, N5195, N4618, N2529);
not NOT1 (N5198, N5190);
or OR2 (N5199, N5198, N229);
buf BUF1 (N5200, N5183);
or OR4 (N5201, N5177, N2009, N2650, N1432);
xor XOR2 (N5202, N5191, N3545);
and AND3 (N5203, N5202, N1545, N3701);
or OR2 (N5204, N5196, N1643);
not NOT1 (N5205, N5187);
and AND4 (N5206, N5203, N3213, N2916, N2277);
nor NOR3 (N5207, N5206, N2188, N4382);
and AND2 (N5208, N5193, N1022);
not NOT1 (N5209, N5192);
buf BUF1 (N5210, N5204);
xor XOR2 (N5211, N5201, N1099);
nand NAND3 (N5212, N5207, N4762, N3022);
and AND3 (N5213, N5188, N4477, N407);
buf BUF1 (N5214, N5212);
or OR4 (N5215, N5210, N4520, N302, N2088);
and AND3 (N5216, N5215, N1622, N2019);
xor XOR2 (N5217, N5211, N1066);
and AND2 (N5218, N5209, N331);
xor XOR2 (N5219, N5217, N1999);
xor XOR2 (N5220, N5208, N3156);
and AND4 (N5221, N5197, N3458, N5182, N869);
or OR2 (N5222, N5221, N4715);
or OR2 (N5223, N5213, N4972);
not NOT1 (N5224, N5199);
xor XOR2 (N5225, N5219, N3915);
nor NOR4 (N5226, N5224, N888, N818, N2777);
xor XOR2 (N5227, N5218, N3809);
buf BUF1 (N5228, N5226);
or OR4 (N5229, N5214, N2930, N124, N3788);
not NOT1 (N5230, N5228);
and AND4 (N5231, N5220, N996, N2126, N2737);
nand NAND4 (N5232, N5231, N4445, N2884, N3909);
nand NAND3 (N5233, N5229, N2475, N1665);
not NOT1 (N5234, N5233);
nand NAND4 (N5235, N5216, N3359, N2009, N5117);
and AND2 (N5236, N5205, N4723);
nand NAND4 (N5237, N5200, N1961, N2322, N1596);
nand NAND4 (N5238, N5235, N4904, N2981, N848);
or OR3 (N5239, N5237, N1826, N5088);
buf BUF1 (N5240, N5236);
nor NOR2 (N5241, N5230, N137);
nor NOR3 (N5242, N5222, N2028, N2610);
buf BUF1 (N5243, N5238);
nand NAND4 (N5244, N5239, N2688, N3148, N1767);
nand NAND4 (N5245, N5232, N4602, N247, N107);
buf BUF1 (N5246, N5241);
buf BUF1 (N5247, N5223);
buf BUF1 (N5248, N5240);
and AND3 (N5249, N5248, N1388, N3609);
not NOT1 (N5250, N5245);
or OR3 (N5251, N5234, N1569, N189);
and AND2 (N5252, N5242, N739);
nand NAND3 (N5253, N5252, N4730, N2745);
not NOT1 (N5254, N5251);
buf BUF1 (N5255, N5243);
nor NOR2 (N5256, N5227, N487);
or OR2 (N5257, N5253, N3046);
not NOT1 (N5258, N5244);
buf BUF1 (N5259, N5258);
and AND2 (N5260, N5256, N576);
xor XOR2 (N5261, N5254, N4345);
or OR3 (N5262, N5261, N4532, N3701);
xor XOR2 (N5263, N5259, N3839);
and AND3 (N5264, N5255, N2680, N1396);
and AND3 (N5265, N5262, N1586, N4986);
not NOT1 (N5266, N5250);
and AND4 (N5267, N5264, N4793, N223, N2344);
buf BUF1 (N5268, N5263);
not NOT1 (N5269, N5267);
and AND2 (N5270, N5269, N813);
nor NOR4 (N5271, N5249, N1821, N2897, N2500);
not NOT1 (N5272, N5270);
nand NAND4 (N5273, N5225, N3767, N3394, N4666);
xor XOR2 (N5274, N5273, N3388);
buf BUF1 (N5275, N5274);
nor NOR2 (N5276, N5275, N650);
xor XOR2 (N5277, N5265, N3913);
not NOT1 (N5278, N5272);
not NOT1 (N5279, N5266);
not NOT1 (N5280, N5277);
and AND4 (N5281, N5271, N726, N4418, N4635);
nand NAND4 (N5282, N5260, N3029, N4934, N2042);
not NOT1 (N5283, N5276);
or OR4 (N5284, N5278, N2021, N152, N192);
nor NOR3 (N5285, N5282, N1698, N4734);
not NOT1 (N5286, N5280);
nand NAND2 (N5287, N5247, N2178);
or OR2 (N5288, N5286, N4296);
nor NOR4 (N5289, N5288, N792, N5243, N5270);
nand NAND2 (N5290, N5268, N2019);
nand NAND4 (N5291, N5283, N3773, N3779, N2205);
buf BUF1 (N5292, N5281);
not NOT1 (N5293, N5246);
not NOT1 (N5294, N5289);
buf BUF1 (N5295, N5287);
buf BUF1 (N5296, N5293);
or OR4 (N5297, N5291, N1261, N4076, N1781);
or OR2 (N5298, N5284, N867);
or OR4 (N5299, N5257, N4246, N2556, N4839);
xor XOR2 (N5300, N5290, N547);
nor NOR2 (N5301, N5296, N4298);
nand NAND4 (N5302, N5295, N1441, N4869, N2976);
buf BUF1 (N5303, N5299);
nor NOR2 (N5304, N5301, N3860);
or OR2 (N5305, N5292, N4091);
xor XOR2 (N5306, N5304, N1753);
buf BUF1 (N5307, N5297);
xor XOR2 (N5308, N5300, N552);
xor XOR2 (N5309, N5298, N727);
xor XOR2 (N5310, N5307, N3484);
and AND2 (N5311, N5294, N1882);
or OR2 (N5312, N5308, N3862);
nor NOR4 (N5313, N5303, N1586, N1672, N739);
xor XOR2 (N5314, N5313, N2833);
buf BUF1 (N5315, N5302);
and AND4 (N5316, N5310, N3188, N555, N5103);
and AND4 (N5317, N5315, N3884, N5155, N4045);
nor NOR4 (N5318, N5316, N1022, N3482, N4498);
and AND2 (N5319, N5279, N2047);
nand NAND3 (N5320, N5318, N1109, N4697);
not NOT1 (N5321, N5314);
or OR3 (N5322, N5285, N521, N5066);
nor NOR4 (N5323, N5311, N3533, N3352, N4777);
or OR2 (N5324, N5323, N3356);
not NOT1 (N5325, N5319);
nand NAND2 (N5326, N5325, N4383);
buf BUF1 (N5327, N5321);
nand NAND2 (N5328, N5324, N4493);
nor NOR3 (N5329, N5312, N3644, N3478);
nor NOR3 (N5330, N5309, N451, N496);
or OR4 (N5331, N5327, N5186, N3668, N995);
not NOT1 (N5332, N5326);
or OR2 (N5333, N5305, N4044);
nand NAND3 (N5334, N5317, N83, N331);
nor NOR3 (N5335, N5332, N444, N3353);
xor XOR2 (N5336, N5328, N3165);
and AND4 (N5337, N5336, N555, N2977, N1898);
or OR4 (N5338, N5335, N4433, N4758, N3205);
nor NOR2 (N5339, N5333, N2172);
or OR4 (N5340, N5338, N829, N2730, N1485);
nor NOR4 (N5341, N5337, N4187, N4432, N3812);
and AND2 (N5342, N5306, N138);
or OR2 (N5343, N5340, N4619);
and AND4 (N5344, N5341, N1020, N3848, N1114);
and AND3 (N5345, N5344, N4459, N3362);
and AND3 (N5346, N5334, N604, N4157);
not NOT1 (N5347, N5345);
nor NOR2 (N5348, N5342, N3683);
nand NAND3 (N5349, N5346, N4507, N1035);
xor XOR2 (N5350, N5329, N177);
not NOT1 (N5351, N5320);
buf BUF1 (N5352, N5339);
or OR3 (N5353, N5331, N3320, N5066);
and AND2 (N5354, N5348, N1141);
and AND4 (N5355, N5322, N4528, N4275, N640);
nand NAND3 (N5356, N5330, N2714, N3768);
xor XOR2 (N5357, N5349, N1236);
and AND3 (N5358, N5351, N1670, N2534);
not NOT1 (N5359, N5357);
or OR3 (N5360, N5355, N2045, N4312);
and AND3 (N5361, N5352, N402, N5006);
and AND2 (N5362, N5343, N4258);
xor XOR2 (N5363, N5362, N2022);
xor XOR2 (N5364, N5359, N3676);
and AND2 (N5365, N5363, N997);
nand NAND2 (N5366, N5354, N2753);
and AND3 (N5367, N5350, N1024, N2865);
nor NOR3 (N5368, N5360, N3310, N1428);
nor NOR4 (N5369, N5364, N975, N2147, N660);
or OR2 (N5370, N5369, N1424);
not NOT1 (N5371, N5365);
xor XOR2 (N5372, N5361, N2077);
nand NAND2 (N5373, N5347, N4509);
not NOT1 (N5374, N5356);
buf BUF1 (N5375, N5371);
not NOT1 (N5376, N5353);
and AND2 (N5377, N5366, N794);
xor XOR2 (N5378, N5367, N1289);
and AND4 (N5379, N5372, N3838, N2758, N4228);
not NOT1 (N5380, N5377);
nand NAND2 (N5381, N5379, N375);
nand NAND3 (N5382, N5370, N2196, N3780);
and AND2 (N5383, N5382, N1104);
or OR2 (N5384, N5378, N11);
buf BUF1 (N5385, N5383);
nor NOR3 (N5386, N5373, N2970, N306);
and AND3 (N5387, N5374, N4364, N89);
buf BUF1 (N5388, N5368);
not NOT1 (N5389, N5375);
nor NOR2 (N5390, N5385, N1538);
xor XOR2 (N5391, N5358, N1928);
nor NOR2 (N5392, N5381, N916);
nor NOR4 (N5393, N5391, N1847, N1515, N787);
nor NOR3 (N5394, N5388, N4671, N43);
xor XOR2 (N5395, N5384, N1509);
not NOT1 (N5396, N5380);
buf BUF1 (N5397, N5395);
buf BUF1 (N5398, N5376);
xor XOR2 (N5399, N5398, N5210);
not NOT1 (N5400, N5392);
buf BUF1 (N5401, N5393);
xor XOR2 (N5402, N5394, N4568);
xor XOR2 (N5403, N5401, N995);
xor XOR2 (N5404, N5397, N3313);
nand NAND3 (N5405, N5402, N1110, N1078);
xor XOR2 (N5406, N5390, N4660);
buf BUF1 (N5407, N5387);
or OR3 (N5408, N5400, N1441, N5303);
or OR4 (N5409, N5407, N3642, N414, N4274);
buf BUF1 (N5410, N5403);
and AND3 (N5411, N5396, N1315, N4291);
xor XOR2 (N5412, N5406, N2455);
buf BUF1 (N5413, N5408);
not NOT1 (N5414, N5411);
xor XOR2 (N5415, N5413, N5003);
nand NAND2 (N5416, N5399, N195);
xor XOR2 (N5417, N5412, N521);
nand NAND4 (N5418, N5404, N1999, N647, N1456);
or OR3 (N5419, N5418, N3927, N4684);
and AND2 (N5420, N5410, N2073);
nand NAND4 (N5421, N5417, N5306, N1192, N1632);
not NOT1 (N5422, N5405);
nor NOR4 (N5423, N5419, N1705, N2792, N3102);
not NOT1 (N5424, N5416);
not NOT1 (N5425, N5409);
xor XOR2 (N5426, N5414, N4690);
xor XOR2 (N5427, N5421, N3905);
nand NAND2 (N5428, N5420, N999);
or OR3 (N5429, N5428, N1315, N4867);
nand NAND2 (N5430, N5427, N1960);
nand NAND4 (N5431, N5423, N2407, N1251, N3823);
and AND3 (N5432, N5386, N234, N1527);
nor NOR4 (N5433, N5430, N4485, N937, N687);
and AND2 (N5434, N5415, N5240);
xor XOR2 (N5435, N5389, N2649);
xor XOR2 (N5436, N5433, N3657);
and AND2 (N5437, N5435, N4926);
nor NOR4 (N5438, N5434, N3391, N903, N1104);
xor XOR2 (N5439, N5437, N2052);
xor XOR2 (N5440, N5432, N3951);
and AND4 (N5441, N5436, N3408, N1861, N1818);
nand NAND4 (N5442, N5424, N4702, N2974, N1417);
nand NAND2 (N5443, N5426, N2904);
and AND3 (N5444, N5442, N818, N3836);
nor NOR3 (N5445, N5444, N2937, N2038);
nor NOR4 (N5446, N5438, N4449, N3762, N2256);
or OR4 (N5447, N5422, N5105, N4228, N4623);
buf BUF1 (N5448, N5446);
buf BUF1 (N5449, N5440);
nor NOR4 (N5450, N5449, N2406, N1436, N2963);
nor NOR2 (N5451, N5441, N737);
xor XOR2 (N5452, N5443, N2957);
and AND2 (N5453, N5445, N2451);
and AND2 (N5454, N5450, N5042);
nor NOR2 (N5455, N5451, N3534);
xor XOR2 (N5456, N5447, N2331);
buf BUF1 (N5457, N5425);
nand NAND2 (N5458, N5431, N4537);
not NOT1 (N5459, N5454);
nand NAND3 (N5460, N5429, N278, N475);
nor NOR4 (N5461, N5456, N5190, N3980, N2205);
not NOT1 (N5462, N5461);
not NOT1 (N5463, N5462);
or OR2 (N5464, N5458, N3052);
buf BUF1 (N5465, N5464);
nor NOR2 (N5466, N5457, N3118);
xor XOR2 (N5467, N5452, N4836);
not NOT1 (N5468, N5466);
not NOT1 (N5469, N5459);
nand NAND4 (N5470, N5439, N1259, N4969, N1003);
buf BUF1 (N5471, N5470);
buf BUF1 (N5472, N5471);
xor XOR2 (N5473, N5453, N2271);
nand NAND2 (N5474, N5468, N4880);
nor NOR3 (N5475, N5469, N1747, N3746);
nor NOR2 (N5476, N5475, N4662);
buf BUF1 (N5477, N5460);
nor NOR3 (N5478, N5474, N2236, N2975);
not NOT1 (N5479, N5465);
nor NOR2 (N5480, N5467, N4721);
nor NOR4 (N5481, N5463, N2814, N2640, N4433);
or OR3 (N5482, N5480, N1818, N3512);
or OR4 (N5483, N5481, N5170, N1328, N846);
buf BUF1 (N5484, N5473);
nor NOR3 (N5485, N5455, N2109, N3847);
buf BUF1 (N5486, N5448);
or OR2 (N5487, N5482, N1550);
not NOT1 (N5488, N5476);
nor NOR3 (N5489, N5488, N4656, N1116);
nor NOR3 (N5490, N5489, N3019, N2691);
nand NAND4 (N5491, N5478, N2851, N3426, N3);
and AND2 (N5492, N5490, N2022);
xor XOR2 (N5493, N5483, N4243);
nor NOR2 (N5494, N5492, N1601);
and AND4 (N5495, N5491, N3537, N5000, N4630);
not NOT1 (N5496, N5486);
and AND3 (N5497, N5496, N4410, N1136);
nor NOR4 (N5498, N5484, N2989, N1824, N612);
nor NOR3 (N5499, N5487, N1429, N2702);
not NOT1 (N5500, N5479);
or OR3 (N5501, N5499, N1731, N3607);
buf BUF1 (N5502, N5498);
nor NOR4 (N5503, N5502, N470, N2558, N1036);
nor NOR3 (N5504, N5472, N1818, N1848);
buf BUF1 (N5505, N5500);
not NOT1 (N5506, N5505);
or OR2 (N5507, N5495, N3631);
or OR2 (N5508, N5497, N4735);
xor XOR2 (N5509, N5494, N25);
and AND2 (N5510, N5504, N715);
nor NOR3 (N5511, N5506, N5192, N2550);
and AND3 (N5512, N5508, N3721, N396);
or OR3 (N5513, N5509, N3916, N751);
buf BUF1 (N5514, N5512);
xor XOR2 (N5515, N5513, N5043);
xor XOR2 (N5516, N5507, N3725);
nand NAND3 (N5517, N5511, N2914, N2822);
not NOT1 (N5518, N5516);
nor NOR3 (N5519, N5477, N4085, N4380);
not NOT1 (N5520, N5485);
xor XOR2 (N5521, N5519, N3327);
not NOT1 (N5522, N5514);
or OR2 (N5523, N5493, N921);
xor XOR2 (N5524, N5517, N3931);
nand NAND3 (N5525, N5523, N5192, N2165);
and AND2 (N5526, N5510, N1425);
nor NOR4 (N5527, N5515, N3956, N3042, N399);
nand NAND3 (N5528, N5522, N4800, N2958);
or OR4 (N5529, N5518, N2502, N1730, N3666);
not NOT1 (N5530, N5520);
or OR3 (N5531, N5525, N3637, N2265);
and AND3 (N5532, N5528, N4534, N959);
or OR3 (N5533, N5531, N5469, N172);
or OR2 (N5534, N5533, N3282);
not NOT1 (N5535, N5532);
xor XOR2 (N5536, N5530, N2796);
xor XOR2 (N5537, N5501, N4032);
nor NOR4 (N5538, N5535, N3234, N193, N5513);
xor XOR2 (N5539, N5537, N802);
buf BUF1 (N5540, N5529);
and AND2 (N5541, N5539, N518);
nand NAND4 (N5542, N5536, N2714, N5483, N627);
not NOT1 (N5543, N5542);
nand NAND4 (N5544, N5526, N3636, N518, N3331);
nor NOR2 (N5545, N5534, N3597);
nor NOR2 (N5546, N5503, N1348);
and AND2 (N5547, N5524, N4408);
nor NOR2 (N5548, N5544, N5017);
nor NOR3 (N5549, N5545, N4433, N2966);
buf BUF1 (N5550, N5538);
or OR2 (N5551, N5543, N3472);
not NOT1 (N5552, N5551);
and AND2 (N5553, N5550, N2913);
xor XOR2 (N5554, N5521, N3609);
buf BUF1 (N5555, N5547);
not NOT1 (N5556, N5555);
nor NOR4 (N5557, N5556, N2261, N4621, N5457);
nand NAND2 (N5558, N5546, N4895);
nor NOR3 (N5559, N5548, N1354, N598);
not NOT1 (N5560, N5559);
buf BUF1 (N5561, N5553);
xor XOR2 (N5562, N5557, N1705);
buf BUF1 (N5563, N5554);
xor XOR2 (N5564, N5540, N2398);
and AND2 (N5565, N5549, N642);
or OR3 (N5566, N5558, N1925, N4450);
and AND4 (N5567, N5566, N5301, N558, N4853);
not NOT1 (N5568, N5527);
nor NOR2 (N5569, N5541, N3487);
or OR4 (N5570, N5565, N1364, N354, N3543);
xor XOR2 (N5571, N5567, N1495);
and AND3 (N5572, N5571, N840, N88);
xor XOR2 (N5573, N5572, N4760);
buf BUF1 (N5574, N5568);
nor NOR4 (N5575, N5562, N4604, N953, N1061);
nand NAND2 (N5576, N5560, N2739);
nor NOR3 (N5577, N5563, N1274, N1693);
nor NOR2 (N5578, N5570, N2136);
nor NOR3 (N5579, N5573, N1376, N5001);
or OR2 (N5580, N5569, N944);
buf BUF1 (N5581, N5564);
nand NAND3 (N5582, N5579, N1392, N2113);
buf BUF1 (N5583, N5561);
nor NOR3 (N5584, N5581, N4050, N2059);
or OR2 (N5585, N5578, N110);
xor XOR2 (N5586, N5575, N902);
and AND3 (N5587, N5552, N5089, N4728);
xor XOR2 (N5588, N5582, N2635);
xor XOR2 (N5589, N5577, N1083);
or OR2 (N5590, N5583, N31);
xor XOR2 (N5591, N5587, N1872);
nor NOR2 (N5592, N5580, N459);
buf BUF1 (N5593, N5591);
or OR2 (N5594, N5576, N5508);
buf BUF1 (N5595, N5574);
buf BUF1 (N5596, N5593);
and AND4 (N5597, N5588, N2816, N1956, N668);
nand NAND3 (N5598, N5584, N3525, N3266);
buf BUF1 (N5599, N5594);
nand NAND4 (N5600, N5585, N4598, N829, N5025);
nand NAND4 (N5601, N5589, N2578, N3522, N703);
not NOT1 (N5602, N5586);
not NOT1 (N5603, N5598);
not NOT1 (N5604, N5590);
nor NOR4 (N5605, N5595, N5143, N5546, N2552);
not NOT1 (N5606, N5602);
nand NAND4 (N5607, N5601, N1304, N2939, N1789);
not NOT1 (N5608, N5606);
nand NAND3 (N5609, N5605, N2149, N2955);
not NOT1 (N5610, N5609);
nor NOR2 (N5611, N5603, N1224);
and AND4 (N5612, N5604, N604, N3761, N1948);
or OR4 (N5613, N5608, N1663, N2432, N4707);
xor XOR2 (N5614, N5596, N855);
or OR3 (N5615, N5592, N465, N564);
nor NOR4 (N5616, N5610, N5555, N5028, N3579);
nand NAND3 (N5617, N5611, N584, N4199);
buf BUF1 (N5618, N5600);
or OR3 (N5619, N5597, N3516, N3330);
nor NOR2 (N5620, N5618, N5596);
xor XOR2 (N5621, N5617, N2043);
xor XOR2 (N5622, N5599, N5221);
nand NAND2 (N5623, N5607, N1700);
buf BUF1 (N5624, N5615);
not NOT1 (N5625, N5614);
and AND2 (N5626, N5625, N3390);
nand NAND4 (N5627, N5623, N4948, N3577, N1656);
not NOT1 (N5628, N5627);
nand NAND3 (N5629, N5624, N3274, N5151);
or OR4 (N5630, N5619, N2439, N3528, N3689);
xor XOR2 (N5631, N5630, N4);
buf BUF1 (N5632, N5616);
xor XOR2 (N5633, N5612, N4985);
not NOT1 (N5634, N5632);
and AND2 (N5635, N5634, N4445);
buf BUF1 (N5636, N5629);
nor NOR3 (N5637, N5628, N5507, N20);
buf BUF1 (N5638, N5635);
and AND3 (N5639, N5620, N980, N574);
or OR4 (N5640, N5621, N1550, N914, N4094);
xor XOR2 (N5641, N5636, N2235);
buf BUF1 (N5642, N5641);
not NOT1 (N5643, N5637);
not NOT1 (N5644, N5643);
nor NOR3 (N5645, N5644, N4211, N913);
and AND2 (N5646, N5642, N4254);
buf BUF1 (N5647, N5646);
not NOT1 (N5648, N5639);
nor NOR4 (N5649, N5645, N5608, N5593, N1955);
buf BUF1 (N5650, N5622);
and AND4 (N5651, N5633, N5129, N201, N1093);
nand NAND2 (N5652, N5651, N4111);
buf BUF1 (N5653, N5613);
nand NAND2 (N5654, N5652, N2858);
nor NOR4 (N5655, N5653, N2682, N1483, N3359);
nand NAND4 (N5656, N5640, N137, N3777, N1427);
or OR2 (N5657, N5648, N813);
xor XOR2 (N5658, N5656, N2640);
or OR3 (N5659, N5655, N4399, N5025);
buf BUF1 (N5660, N5626);
xor XOR2 (N5661, N5650, N5273);
nor NOR2 (N5662, N5654, N2580);
or OR4 (N5663, N5649, N2537, N2208, N4675);
not NOT1 (N5664, N5647);
and AND2 (N5665, N5638, N5289);
and AND4 (N5666, N5664, N4507, N4433, N4379);
buf BUF1 (N5667, N5631);
not NOT1 (N5668, N5661);
or OR4 (N5669, N5659, N1612, N3950, N1270);
not NOT1 (N5670, N5663);
or OR2 (N5671, N5662, N5614);
nand NAND3 (N5672, N5657, N3840, N5310);
nor NOR2 (N5673, N5667, N896);
and AND4 (N5674, N5671, N616, N3801, N5118);
not NOT1 (N5675, N5660);
buf BUF1 (N5676, N5658);
buf BUF1 (N5677, N5674);
xor XOR2 (N5678, N5666, N1819);
nor NOR4 (N5679, N5668, N3153, N1634, N3488);
nand NAND4 (N5680, N5676, N5225, N768, N2438);
or OR3 (N5681, N5665, N4073, N2547);
not NOT1 (N5682, N5677);
buf BUF1 (N5683, N5680);
not NOT1 (N5684, N5679);
not NOT1 (N5685, N5675);
buf BUF1 (N5686, N5670);
buf BUF1 (N5687, N5669);
not NOT1 (N5688, N5685);
nand NAND2 (N5689, N5682, N4875);
xor XOR2 (N5690, N5689, N4837);
nor NOR3 (N5691, N5678, N2914, N3483);
xor XOR2 (N5692, N5683, N3478);
nor NOR2 (N5693, N5686, N4469);
nand NAND4 (N5694, N5684, N319, N4468, N231);
buf BUF1 (N5695, N5692);
xor XOR2 (N5696, N5695, N4858);
nor NOR3 (N5697, N5690, N461, N3792);
not NOT1 (N5698, N5688);
not NOT1 (N5699, N5681);
nand NAND3 (N5700, N5673, N1388, N3402);
nor NOR3 (N5701, N5697, N5304, N2386);
not NOT1 (N5702, N5700);
nand NAND4 (N5703, N5694, N1385, N2575, N3010);
xor XOR2 (N5704, N5701, N374);
not NOT1 (N5705, N5702);
xor XOR2 (N5706, N5693, N4049);
and AND3 (N5707, N5706, N5610, N3478);
buf BUF1 (N5708, N5672);
or OR3 (N5709, N5696, N1523, N190);
and AND3 (N5710, N5704, N675, N5486);
buf BUF1 (N5711, N5691);
buf BUF1 (N5712, N5698);
buf BUF1 (N5713, N5699);
and AND2 (N5714, N5687, N1665);
nand NAND3 (N5715, N5713, N100, N2856);
nand NAND4 (N5716, N5715, N4983, N2541, N1156);
and AND3 (N5717, N5714, N404, N1422);
not NOT1 (N5718, N5717);
nor NOR2 (N5719, N5712, N230);
nor NOR3 (N5720, N5709, N1049, N41);
and AND3 (N5721, N5718, N2162, N2232);
nand NAND3 (N5722, N5707, N3701, N5717);
not NOT1 (N5723, N5722);
buf BUF1 (N5724, N5711);
nand NAND3 (N5725, N5705, N119, N5258);
or OR4 (N5726, N5710, N5031, N1588, N206);
nand NAND2 (N5727, N5721, N1980);
buf BUF1 (N5728, N5724);
xor XOR2 (N5729, N5727, N942);
and AND2 (N5730, N5725, N4768);
buf BUF1 (N5731, N5730);
and AND2 (N5732, N5703, N1467);
buf BUF1 (N5733, N5728);
xor XOR2 (N5734, N5732, N2254);
nor NOR2 (N5735, N5726, N4902);
xor XOR2 (N5736, N5723, N3476);
or OR2 (N5737, N5729, N2039);
not NOT1 (N5738, N5719);
and AND3 (N5739, N5733, N1979, N244);
xor XOR2 (N5740, N5708, N5036);
buf BUF1 (N5741, N5738);
or OR3 (N5742, N5740, N4141, N238);
not NOT1 (N5743, N5720);
xor XOR2 (N5744, N5741, N4618);
and AND3 (N5745, N5734, N1317, N2062);
or OR4 (N5746, N5716, N2985, N709, N1625);
and AND2 (N5747, N5735, N4998);
not NOT1 (N5748, N5736);
or OR4 (N5749, N5746, N4168, N3981, N2418);
buf BUF1 (N5750, N5731);
and AND4 (N5751, N5748, N2445, N2794, N4931);
or OR3 (N5752, N5743, N3878, N2650);
nand NAND4 (N5753, N5747, N4441, N1037, N1026);
xor XOR2 (N5754, N5737, N23);
and AND2 (N5755, N5742, N3334);
nand NAND4 (N5756, N5754, N1752, N2260, N1754);
buf BUF1 (N5757, N5739);
buf BUF1 (N5758, N5755);
nand NAND2 (N5759, N5753, N4484);
not NOT1 (N5760, N5750);
nand NAND2 (N5761, N5745, N718);
or OR3 (N5762, N5756, N2372, N214);
or OR2 (N5763, N5752, N2908);
and AND4 (N5764, N5760, N1992, N1418, N2192);
and AND4 (N5765, N5764, N1833, N387, N222);
xor XOR2 (N5766, N5763, N5180);
or OR4 (N5767, N5757, N3580, N3969, N4695);
or OR3 (N5768, N5765, N2799, N1958);
buf BUF1 (N5769, N5767);
buf BUF1 (N5770, N5744);
nand NAND4 (N5771, N5766, N3186, N5621, N3601);
nand NAND3 (N5772, N5769, N4367, N1486);
buf BUF1 (N5773, N5761);
nor NOR4 (N5774, N5772, N4423, N2412, N4223);
nand NAND4 (N5775, N5771, N5216, N2533, N383);
or OR2 (N5776, N5759, N175);
and AND3 (N5777, N5770, N3796, N5201);
xor XOR2 (N5778, N5777, N1523);
buf BUF1 (N5779, N5758);
nor NOR4 (N5780, N5762, N1364, N3667, N1569);
xor XOR2 (N5781, N5749, N132);
or OR4 (N5782, N5778, N3292, N5207, N463);
nor NOR3 (N5783, N5773, N64, N4522);
xor XOR2 (N5784, N5776, N1614);
nor NOR2 (N5785, N5768, N4073);
nand NAND3 (N5786, N5779, N3439, N673);
buf BUF1 (N5787, N5780);
not NOT1 (N5788, N5781);
xor XOR2 (N5789, N5775, N2784);
xor XOR2 (N5790, N5751, N1724);
buf BUF1 (N5791, N5785);
or OR3 (N5792, N5783, N4814, N3360);
xor XOR2 (N5793, N5774, N1035);
or OR2 (N5794, N5792, N5501);
nand NAND4 (N5795, N5784, N368, N275, N1566);
xor XOR2 (N5796, N5794, N5748);
or OR4 (N5797, N5790, N757, N5242, N1232);
xor XOR2 (N5798, N5788, N1402);
buf BUF1 (N5799, N5786);
nand NAND4 (N5800, N5787, N286, N5197, N2611);
nand NAND4 (N5801, N5798, N1155, N3806, N1099);
nor NOR2 (N5802, N5800, N2383);
xor XOR2 (N5803, N5793, N282);
xor XOR2 (N5804, N5791, N4641);
not NOT1 (N5805, N5804);
not NOT1 (N5806, N5797);
or OR2 (N5807, N5801, N2979);
nor NOR3 (N5808, N5806, N2414, N1544);
or OR2 (N5809, N5796, N2936);
and AND2 (N5810, N5808, N3295);
nand NAND2 (N5811, N5799, N5658);
buf BUF1 (N5812, N5807);
nor NOR4 (N5813, N5805, N1552, N3495, N1473);
not NOT1 (N5814, N5795);
and AND4 (N5815, N5782, N5573, N5077, N2903);
or OR2 (N5816, N5815, N2000);
buf BUF1 (N5817, N5803);
nor NOR2 (N5818, N5816, N2766);
not NOT1 (N5819, N5802);
xor XOR2 (N5820, N5814, N4770);
or OR2 (N5821, N5819, N557);
or OR2 (N5822, N5821, N3045);
buf BUF1 (N5823, N5811);
buf BUF1 (N5824, N5813);
buf BUF1 (N5825, N5824);
nand NAND4 (N5826, N5817, N4574, N2470, N875);
xor XOR2 (N5827, N5789, N2133);
and AND2 (N5828, N5822, N950);
nor NOR2 (N5829, N5828, N399);
nand NAND3 (N5830, N5812, N2878, N735);
or OR3 (N5831, N5810, N3438, N3445);
xor XOR2 (N5832, N5809, N2359);
not NOT1 (N5833, N5830);
nor NOR4 (N5834, N5826, N2195, N2184, N732);
and AND4 (N5835, N5823, N1178, N5620, N2830);
buf BUF1 (N5836, N5827);
or OR4 (N5837, N5834, N2434, N1747, N3064);
or OR4 (N5838, N5833, N2226, N4761, N3041);
nor NOR4 (N5839, N5836, N5135, N3950, N2622);
not NOT1 (N5840, N5820);
or OR4 (N5841, N5835, N1169, N4257, N957);
or OR4 (N5842, N5818, N3428, N4600, N4009);
not NOT1 (N5843, N5839);
and AND3 (N5844, N5825, N4656, N646);
nand NAND4 (N5845, N5838, N3423, N1943, N5698);
and AND2 (N5846, N5831, N426);
and AND2 (N5847, N5842, N601);
nor NOR3 (N5848, N5837, N683, N1127);
not NOT1 (N5849, N5845);
or OR3 (N5850, N5840, N889, N31);
not NOT1 (N5851, N5832);
not NOT1 (N5852, N5829);
nand NAND2 (N5853, N5852, N5518);
nand NAND4 (N5854, N5841, N5074, N2751, N2935);
nand NAND4 (N5855, N5843, N354, N3001, N5763);
not NOT1 (N5856, N5848);
nand NAND4 (N5857, N5847, N2141, N5804, N1599);
nor NOR4 (N5858, N5846, N5114, N232, N347);
and AND2 (N5859, N5850, N2266);
nor NOR3 (N5860, N5851, N94, N288);
not NOT1 (N5861, N5844);
or OR2 (N5862, N5855, N2245);
or OR2 (N5863, N5857, N1478);
xor XOR2 (N5864, N5860, N2521);
nor NOR4 (N5865, N5863, N4309, N3353, N2153);
nand NAND2 (N5866, N5858, N2706);
xor XOR2 (N5867, N5854, N5749);
or OR2 (N5868, N5859, N1457);
nor NOR2 (N5869, N5862, N1786);
nand NAND3 (N5870, N5869, N2447, N508);
not NOT1 (N5871, N5861);
nor NOR4 (N5872, N5864, N2124, N5778, N2512);
nor NOR2 (N5873, N5872, N452);
nand NAND2 (N5874, N5856, N306);
nor NOR3 (N5875, N5873, N3055, N5596);
and AND2 (N5876, N5865, N4633);
buf BUF1 (N5877, N5876);
buf BUF1 (N5878, N5871);
buf BUF1 (N5879, N5874);
buf BUF1 (N5880, N5866);
not NOT1 (N5881, N5853);
xor XOR2 (N5882, N5867, N3870);
or OR3 (N5883, N5870, N5370, N3934);
buf BUF1 (N5884, N5880);
not NOT1 (N5885, N5881);
and AND3 (N5886, N5877, N5115, N5367);
or OR3 (N5887, N5849, N5145, N3558);
buf BUF1 (N5888, N5878);
not NOT1 (N5889, N5888);
nor NOR3 (N5890, N5887, N4335, N3313);
nor NOR4 (N5891, N5875, N2361, N3361, N1970);
and AND4 (N5892, N5883, N1801, N3958, N3449);
or OR3 (N5893, N5892, N2058, N3752);
and AND3 (N5894, N5886, N1114, N3992);
nor NOR2 (N5895, N5868, N2150);
buf BUF1 (N5896, N5884);
nor NOR2 (N5897, N5879, N153);
xor XOR2 (N5898, N5895, N5565);
and AND3 (N5899, N5898, N2444, N3934);
nand NAND3 (N5900, N5897, N902, N142);
buf BUF1 (N5901, N5900);
nand NAND4 (N5902, N5890, N1570, N1950, N4864);
nor NOR3 (N5903, N5896, N5360, N4757);
not NOT1 (N5904, N5891);
or OR4 (N5905, N5901, N714, N2056, N5353);
xor XOR2 (N5906, N5885, N3534);
xor XOR2 (N5907, N5882, N1824);
nor NOR2 (N5908, N5889, N3814);
buf BUF1 (N5909, N5904);
and AND4 (N5910, N5905, N2319, N4985, N1218);
not NOT1 (N5911, N5909);
xor XOR2 (N5912, N5910, N5157);
buf BUF1 (N5913, N5893);
xor XOR2 (N5914, N5902, N1606);
nand NAND2 (N5915, N5894, N4794);
nand NAND3 (N5916, N5908, N775, N5863);
nor NOR4 (N5917, N5906, N2100, N2559, N2653);
nor NOR3 (N5918, N5911, N2417, N2041);
or OR2 (N5919, N5916, N288);
or OR2 (N5920, N5899, N4795);
nor NOR2 (N5921, N5914, N1900);
and AND3 (N5922, N5920, N42, N2214);
and AND3 (N5923, N5907, N480, N875);
nand NAND3 (N5924, N5913, N3703, N5034);
or OR2 (N5925, N5919, N5745);
not NOT1 (N5926, N5917);
nor NOR2 (N5927, N5924, N5600);
nor NOR3 (N5928, N5926, N3278, N4270);
and AND4 (N5929, N5928, N5038, N5343, N2576);
not NOT1 (N5930, N5922);
or OR4 (N5931, N5923, N1342, N1650, N2565);
xor XOR2 (N5932, N5927, N2379);
nand NAND4 (N5933, N5931, N3239, N128, N5774);
not NOT1 (N5934, N5912);
or OR2 (N5935, N5921, N4923);
not NOT1 (N5936, N5934);
or OR2 (N5937, N5915, N4299);
nand NAND3 (N5938, N5925, N5383, N2268);
and AND2 (N5939, N5918, N1471);
buf BUF1 (N5940, N5936);
or OR3 (N5941, N5903, N1326, N4193);
buf BUF1 (N5942, N5938);
nor NOR4 (N5943, N5933, N2964, N3609, N1825);
nor NOR4 (N5944, N5930, N4100, N3263, N5487);
nor NOR3 (N5945, N5932, N5710, N2758);
or OR2 (N5946, N5942, N2824);
and AND2 (N5947, N5943, N2789);
nor NOR3 (N5948, N5945, N2760, N3770);
or OR3 (N5949, N5946, N1661, N3797);
xor XOR2 (N5950, N5947, N2583);
xor XOR2 (N5951, N5939, N4688);
xor XOR2 (N5952, N5935, N2325);
xor XOR2 (N5953, N5940, N3909);
xor XOR2 (N5954, N5953, N4698);
xor XOR2 (N5955, N5937, N997);
xor XOR2 (N5956, N5929, N4693);
and AND2 (N5957, N5950, N3093);
or OR4 (N5958, N5954, N2713, N701, N4188);
buf BUF1 (N5959, N5952);
nor NOR2 (N5960, N5944, N1374);
and AND4 (N5961, N5955, N3117, N2931, N4861);
nand NAND4 (N5962, N5948, N3904, N3053, N5447);
buf BUF1 (N5963, N5951);
not NOT1 (N5964, N5949);
or OR4 (N5965, N5957, N182, N3642, N1616);
nand NAND4 (N5966, N5964, N2916, N2145, N2698);
nor NOR3 (N5967, N5956, N4668, N2796);
not NOT1 (N5968, N5941);
not NOT1 (N5969, N5958);
xor XOR2 (N5970, N5960, N2631);
or OR2 (N5971, N5959, N3288);
nor NOR4 (N5972, N5962, N2776, N5177, N4860);
xor XOR2 (N5973, N5970, N3134);
or OR2 (N5974, N5968, N1237);
nand NAND4 (N5975, N5963, N4635, N1814, N3517);
buf BUF1 (N5976, N5974);
nor NOR2 (N5977, N5973, N2820);
xor XOR2 (N5978, N5965, N4951);
not NOT1 (N5979, N5966);
and AND2 (N5980, N5976, N5543);
nor NOR4 (N5981, N5978, N5361, N5476, N4880);
not NOT1 (N5982, N5972);
or OR3 (N5983, N5969, N4228, N59);
nand NAND4 (N5984, N5975, N3064, N734, N1556);
or OR2 (N5985, N5981, N5443);
buf BUF1 (N5986, N5983);
buf BUF1 (N5987, N5979);
xor XOR2 (N5988, N5980, N3380);
nor NOR3 (N5989, N5982, N1453, N1258);
xor XOR2 (N5990, N5987, N4228);
not NOT1 (N5991, N5961);
not NOT1 (N5992, N5985);
buf BUF1 (N5993, N5971);
xor XOR2 (N5994, N5988, N5953);
xor XOR2 (N5995, N5977, N907);
buf BUF1 (N5996, N5967);
nor NOR4 (N5997, N5993, N4777, N5349, N4803);
xor XOR2 (N5998, N5996, N245);
buf BUF1 (N5999, N5991);
nand NAND2 (N6000, N5997, N911);
or OR3 (N6001, N5994, N3004, N214);
nor NOR2 (N6002, N5999, N5037);
xor XOR2 (N6003, N6001, N5286);
nand NAND2 (N6004, N5992, N2333);
and AND3 (N6005, N5986, N1490, N591);
nor NOR2 (N6006, N6004, N2573);
not NOT1 (N6007, N5998);
nor NOR4 (N6008, N5989, N1627, N3181, N2179);
nand NAND4 (N6009, N5990, N5352, N1871, N2421);
and AND4 (N6010, N6002, N469, N704, N3844);
nor NOR3 (N6011, N5984, N3883, N5278);
nand NAND2 (N6012, N6006, N3271);
xor XOR2 (N6013, N6012, N3304);
or OR3 (N6014, N6011, N900, N5546);
nor NOR2 (N6015, N6009, N1417);
or OR3 (N6016, N6014, N2144, N3776);
nor NOR3 (N6017, N6013, N221, N4387);
buf BUF1 (N6018, N6000);
nand NAND3 (N6019, N5995, N5973, N351);
not NOT1 (N6020, N6007);
xor XOR2 (N6021, N6017, N729);
nor NOR4 (N6022, N6021, N4703, N3024, N2299);
buf BUF1 (N6023, N6008);
nand NAND3 (N6024, N6020, N660, N1679);
xor XOR2 (N6025, N6015, N1466);
nand NAND4 (N6026, N6016, N3141, N826, N4427);
nand NAND3 (N6027, N6010, N4005, N253);
and AND4 (N6028, N6003, N2090, N5092, N2033);
xor XOR2 (N6029, N6019, N1899);
not NOT1 (N6030, N6022);
not NOT1 (N6031, N6018);
not NOT1 (N6032, N6024);
nand NAND3 (N6033, N6028, N4873, N75);
xor XOR2 (N6034, N6005, N3870);
or OR2 (N6035, N6027, N2622);
or OR4 (N6036, N6026, N5809, N3675, N5776);
and AND3 (N6037, N6030, N4812, N5503);
xor XOR2 (N6038, N6025, N5901);
nor NOR4 (N6039, N6029, N3876, N2029, N3164);
not NOT1 (N6040, N6031);
nand NAND4 (N6041, N6039, N3139, N4841, N5698);
or OR2 (N6042, N6023, N4152);
buf BUF1 (N6043, N6041);
buf BUF1 (N6044, N6042);
buf BUF1 (N6045, N6038);
nor NOR4 (N6046, N6043, N5643, N3635, N1764);
and AND2 (N6047, N6032, N4571);
not NOT1 (N6048, N6047);
nand NAND4 (N6049, N6045, N2007, N1181, N5032);
or OR4 (N6050, N6048, N4205, N1340, N5736);
nor NOR3 (N6051, N6046, N4210, N4400);
not NOT1 (N6052, N6034);
nor NOR4 (N6053, N6036, N1109, N3081, N3765);
nor NOR2 (N6054, N6052, N3363);
xor XOR2 (N6055, N6033, N4351);
nor NOR3 (N6056, N6053, N2286, N5949);
buf BUF1 (N6057, N6055);
nand NAND3 (N6058, N6049, N5204, N943);
nand NAND2 (N6059, N6037, N719);
and AND2 (N6060, N6051, N1051);
and AND4 (N6061, N6057, N3005, N816, N5900);
or OR3 (N6062, N6056, N4991, N883);
buf BUF1 (N6063, N6044);
buf BUF1 (N6064, N6054);
buf BUF1 (N6065, N6062);
buf BUF1 (N6066, N6040);
buf BUF1 (N6067, N6059);
xor XOR2 (N6068, N6035, N3770);
nor NOR3 (N6069, N6050, N4830, N920);
and AND3 (N6070, N6058, N1622, N3464);
xor XOR2 (N6071, N6063, N5744);
nand NAND4 (N6072, N6070, N2018, N1913, N1990);
and AND2 (N6073, N6067, N4605);
nand NAND3 (N6074, N6072, N5345, N3512);
nor NOR2 (N6075, N6073, N2390);
nand NAND4 (N6076, N6068, N1276, N4497, N381);
nor NOR2 (N6077, N6061, N1540);
nand NAND2 (N6078, N6069, N4);
nand NAND2 (N6079, N6075, N4649);
xor XOR2 (N6080, N6078, N1732);
nor NOR3 (N6081, N6064, N3792, N4421);
or OR3 (N6082, N6071, N2068, N5230);
buf BUF1 (N6083, N6076);
and AND4 (N6084, N6074, N3204, N486, N4865);
nand NAND4 (N6085, N6084, N365, N877, N670);
not NOT1 (N6086, N6077);
buf BUF1 (N6087, N6085);
nand NAND3 (N6088, N6083, N4531, N1654);
and AND4 (N6089, N6087, N4857, N5691, N1896);
xor XOR2 (N6090, N6079, N2454);
nor NOR3 (N6091, N6089, N2136, N4129);
not NOT1 (N6092, N6080);
or OR4 (N6093, N6092, N4774, N3774, N702);
not NOT1 (N6094, N6066);
xor XOR2 (N6095, N6060, N4527);
or OR3 (N6096, N6088, N595, N3132);
nor NOR3 (N6097, N6086, N2417, N4194);
not NOT1 (N6098, N6081);
nor NOR2 (N6099, N6096, N5938);
and AND2 (N6100, N6095, N3179);
or OR2 (N6101, N6082, N92);
and AND2 (N6102, N6097, N3171);
nand NAND3 (N6103, N6094, N305, N4501);
and AND3 (N6104, N6099, N1230, N5504);
nor NOR2 (N6105, N6100, N5595);
nand NAND2 (N6106, N6098, N4196);
nand NAND4 (N6107, N6091, N22, N3125, N34);
nand NAND2 (N6108, N6103, N5849);
buf BUF1 (N6109, N6105);
buf BUF1 (N6110, N6109);
and AND4 (N6111, N6101, N1241, N5821, N2557);
buf BUF1 (N6112, N6107);
xor XOR2 (N6113, N6106, N5648);
buf BUF1 (N6114, N6093);
buf BUF1 (N6115, N6112);
xor XOR2 (N6116, N6113, N1794);
nor NOR4 (N6117, N6065, N848, N2126, N4694);
nor NOR4 (N6118, N6110, N2051, N4936, N3811);
nor NOR2 (N6119, N6102, N947);
nor NOR3 (N6120, N6111, N3565, N6006);
not NOT1 (N6121, N6090);
or OR3 (N6122, N6114, N4868, N3989);
or OR3 (N6123, N6122, N1280, N153);
or OR2 (N6124, N6119, N4713);
buf BUF1 (N6125, N6115);
nor NOR4 (N6126, N6108, N5416, N3475, N1224);
nand NAND3 (N6127, N6104, N4807, N174);
xor XOR2 (N6128, N6116, N3265);
or OR3 (N6129, N6128, N441, N1795);
buf BUF1 (N6130, N6123);
nand NAND4 (N6131, N6126, N5187, N2858, N396);
not NOT1 (N6132, N6117);
nor NOR2 (N6133, N6118, N5816);
xor XOR2 (N6134, N6131, N341);
nand NAND3 (N6135, N6125, N1414, N1949);
and AND4 (N6136, N6127, N3266, N3768, N5759);
not NOT1 (N6137, N6132);
nand NAND2 (N6138, N6120, N5591);
xor XOR2 (N6139, N6133, N3692);
and AND4 (N6140, N6136, N1872, N1425, N1096);
not NOT1 (N6141, N6138);
nor NOR2 (N6142, N6141, N5214);
nand NAND4 (N6143, N6137, N3026, N2448, N3644);
buf BUF1 (N6144, N6134);
nor NOR2 (N6145, N6140, N2276);
nor NOR2 (N6146, N6129, N6053);
nor NOR4 (N6147, N6145, N3093, N5816, N4792);
not NOT1 (N6148, N6124);
xor XOR2 (N6149, N6121, N1812);
not NOT1 (N6150, N6148);
nand NAND4 (N6151, N6144, N2801, N256, N1718);
xor XOR2 (N6152, N6135, N769);
and AND3 (N6153, N6142, N3447, N5543);
buf BUF1 (N6154, N6150);
or OR2 (N6155, N6146, N6026);
not NOT1 (N6156, N6143);
xor XOR2 (N6157, N6147, N4325);
or OR4 (N6158, N6154, N5578, N1531, N8);
and AND3 (N6159, N6149, N4928, N611);
not NOT1 (N6160, N6155);
nand NAND4 (N6161, N6130, N3173, N1835, N2239);
buf BUF1 (N6162, N6161);
xor XOR2 (N6163, N6152, N2828);
buf BUF1 (N6164, N6159);
nor NOR4 (N6165, N6158, N2636, N3918, N1074);
nor NOR3 (N6166, N6153, N2440, N722);
or OR4 (N6167, N6162, N5582, N263, N2679);
nor NOR2 (N6168, N6164, N6037);
nand NAND3 (N6169, N6156, N714, N2071);
buf BUF1 (N6170, N6151);
buf BUF1 (N6171, N6168);
buf BUF1 (N6172, N6165);
or OR4 (N6173, N6170, N3971, N3169, N2858);
not NOT1 (N6174, N6169);
or OR4 (N6175, N6160, N1977, N5455, N1867);
nor NOR3 (N6176, N6139, N4636, N420);
and AND3 (N6177, N6176, N4237, N2088);
nor NOR2 (N6178, N6167, N1654);
nor NOR3 (N6179, N6157, N4744, N3057);
and AND3 (N6180, N6175, N4850, N5425);
buf BUF1 (N6181, N6177);
xor XOR2 (N6182, N6173, N5273);
and AND3 (N6183, N6178, N1441, N3790);
xor XOR2 (N6184, N6166, N2969);
nand NAND4 (N6185, N6182, N2734, N5574, N4231);
not NOT1 (N6186, N6183);
nand NAND4 (N6187, N6185, N1645, N1304, N1063);
nor NOR2 (N6188, N6174, N5206);
or OR3 (N6189, N6180, N4762, N1622);
and AND2 (N6190, N6181, N2144);
nand NAND3 (N6191, N6186, N4290, N332);
or OR4 (N6192, N6171, N4503, N3331, N2522);
nand NAND3 (N6193, N6163, N4670, N3258);
and AND2 (N6194, N6188, N2316);
and AND4 (N6195, N6193, N4007, N1403, N201);
nand NAND2 (N6196, N6184, N2345);
nand NAND3 (N6197, N6194, N3503, N3156);
xor XOR2 (N6198, N6197, N2399);
and AND2 (N6199, N6189, N5003);
or OR3 (N6200, N6190, N2653, N4852);
and AND2 (N6201, N6200, N5328);
buf BUF1 (N6202, N6187);
xor XOR2 (N6203, N6191, N2372);
nand NAND2 (N6204, N6201, N6168);
or OR3 (N6205, N6199, N4365, N4016);
not NOT1 (N6206, N6192);
or OR2 (N6207, N6203, N2443);
not NOT1 (N6208, N6172);
nor NOR3 (N6209, N6202, N3158, N5471);
and AND4 (N6210, N6209, N3186, N137, N5225);
buf BUF1 (N6211, N6195);
and AND4 (N6212, N6204, N3047, N4491, N5210);
buf BUF1 (N6213, N6179);
not NOT1 (N6214, N6213);
nor NOR3 (N6215, N6196, N3694, N3933);
or OR3 (N6216, N6210, N5783, N4112);
not NOT1 (N6217, N6215);
or OR2 (N6218, N6211, N2568);
and AND2 (N6219, N6205, N3889);
xor XOR2 (N6220, N6217, N4562);
buf BUF1 (N6221, N6206);
and AND2 (N6222, N6216, N3997);
nor NOR3 (N6223, N6221, N688, N231);
or OR4 (N6224, N6212, N447, N4073, N323);
not NOT1 (N6225, N6208);
not NOT1 (N6226, N6224);
and AND3 (N6227, N6218, N3568, N490);
not NOT1 (N6228, N6222);
or OR4 (N6229, N6227, N2646, N224, N3450);
or OR2 (N6230, N6226, N5480);
nand NAND2 (N6231, N6214, N1042);
not NOT1 (N6232, N6231);
buf BUF1 (N6233, N6230);
nand NAND3 (N6234, N6233, N4815, N4154);
nor NOR2 (N6235, N6219, N3808);
and AND2 (N6236, N6232, N3679);
or OR4 (N6237, N6234, N4751, N1408, N4389);
and AND2 (N6238, N6225, N5826);
nor NOR4 (N6239, N6237, N5111, N1210, N5146);
and AND3 (N6240, N6239, N6158, N2013);
or OR3 (N6241, N6198, N1570, N3755);
buf BUF1 (N6242, N6207);
nor NOR3 (N6243, N6241, N3641, N4455);
xor XOR2 (N6244, N6223, N3102);
or OR2 (N6245, N6243, N4864);
not NOT1 (N6246, N6220);
and AND4 (N6247, N6229, N4812, N1554, N1545);
and AND4 (N6248, N6242, N4849, N535, N4125);
buf BUF1 (N6249, N6247);
xor XOR2 (N6250, N6249, N5608);
buf BUF1 (N6251, N6236);
not NOT1 (N6252, N6250);
not NOT1 (N6253, N6248);
nand NAND4 (N6254, N6228, N410, N235, N2222);
xor XOR2 (N6255, N6251, N3637);
nand NAND2 (N6256, N6238, N4824);
nand NAND4 (N6257, N6244, N4961, N523, N4167);
xor XOR2 (N6258, N6245, N5399);
not NOT1 (N6259, N6252);
or OR3 (N6260, N6257, N4668, N4320);
xor XOR2 (N6261, N6254, N4586);
or OR3 (N6262, N6258, N2650, N655);
nor NOR2 (N6263, N6259, N2648);
nand NAND4 (N6264, N6246, N4197, N2728, N2546);
and AND2 (N6265, N6263, N3221);
and AND3 (N6266, N6260, N2789, N2661);
not NOT1 (N6267, N6255);
or OR3 (N6268, N6262, N2022, N877);
or OR4 (N6269, N6268, N3863, N317, N5164);
nand NAND2 (N6270, N6235, N4045);
nor NOR2 (N6271, N6253, N296);
not NOT1 (N6272, N6270);
and AND2 (N6273, N6264, N3626);
not NOT1 (N6274, N6256);
or OR3 (N6275, N6266, N1731, N5685);
not NOT1 (N6276, N6272);
nand NAND2 (N6277, N6274, N4978);
xor XOR2 (N6278, N6277, N1935);
buf BUF1 (N6279, N6240);
or OR2 (N6280, N6276, N3695);
not NOT1 (N6281, N6273);
buf BUF1 (N6282, N6265);
and AND3 (N6283, N6267, N1446, N5130);
buf BUF1 (N6284, N6269);
buf BUF1 (N6285, N6283);
nand NAND3 (N6286, N6261, N5021, N2722);
xor XOR2 (N6287, N6278, N1116);
buf BUF1 (N6288, N6282);
and AND3 (N6289, N6271, N4361, N1132);
xor XOR2 (N6290, N6275, N1947);
buf BUF1 (N6291, N6284);
xor XOR2 (N6292, N6286, N666);
xor XOR2 (N6293, N6279, N737);
not NOT1 (N6294, N6287);
or OR4 (N6295, N6292, N390, N2723, N877);
or OR4 (N6296, N6285, N2905, N4882, N328);
nand NAND3 (N6297, N6281, N5595, N5285);
xor XOR2 (N6298, N6294, N4882);
or OR2 (N6299, N6280, N5862);
or OR4 (N6300, N6289, N4968, N4029, N3478);
not NOT1 (N6301, N6295);
nor NOR4 (N6302, N6290, N5706, N1842, N4341);
buf BUF1 (N6303, N6297);
and AND2 (N6304, N6303, N3127);
and AND3 (N6305, N6293, N1416, N4624);
xor XOR2 (N6306, N6304, N2451);
or OR2 (N6307, N6291, N113);
and AND2 (N6308, N6302, N407);
buf BUF1 (N6309, N6298);
not NOT1 (N6310, N6301);
and AND4 (N6311, N6309, N1404, N3018, N1207);
not NOT1 (N6312, N6300);
nand NAND3 (N6313, N6310, N4028, N2510);
buf BUF1 (N6314, N6312);
buf BUF1 (N6315, N6313);
buf BUF1 (N6316, N6296);
xor XOR2 (N6317, N6288, N5867);
xor XOR2 (N6318, N6308, N4612);
xor XOR2 (N6319, N6305, N3139);
and AND4 (N6320, N6315, N3006, N2772, N6207);
and AND2 (N6321, N6319, N4489);
nor NOR2 (N6322, N6307, N332);
not NOT1 (N6323, N6306);
nand NAND2 (N6324, N6321, N3624);
nor NOR3 (N6325, N6324, N5085, N4902);
nand NAND3 (N6326, N6325, N6056, N2350);
xor XOR2 (N6327, N6323, N2295);
buf BUF1 (N6328, N6327);
nor NOR2 (N6329, N6326, N1742);
and AND4 (N6330, N6299, N4385, N1116, N2889);
nand NAND4 (N6331, N6318, N4249, N4941, N3392);
or OR2 (N6332, N6311, N291);
not NOT1 (N6333, N6314);
nand NAND2 (N6334, N6328, N5160);
nor NOR3 (N6335, N6331, N5035, N1994);
buf BUF1 (N6336, N6320);
nand NAND3 (N6337, N6330, N560, N1265);
buf BUF1 (N6338, N6316);
nand NAND2 (N6339, N6336, N5717);
buf BUF1 (N6340, N6334);
and AND2 (N6341, N6322, N5527);
xor XOR2 (N6342, N6333, N1084);
or OR2 (N6343, N6335, N5795);
buf BUF1 (N6344, N6338);
and AND3 (N6345, N6342, N2168, N4937);
and AND4 (N6346, N6344, N5868, N4519, N941);
xor XOR2 (N6347, N6343, N5022);
nor NOR4 (N6348, N6337, N2421, N5217, N2003);
and AND3 (N6349, N6329, N839, N3884);
nor NOR4 (N6350, N6341, N1399, N4217, N945);
buf BUF1 (N6351, N6349);
and AND2 (N6352, N6339, N1484);
or OR3 (N6353, N6348, N832, N5155);
nand NAND2 (N6354, N6352, N5540);
or OR2 (N6355, N6345, N4319);
and AND2 (N6356, N6317, N3899);
buf BUF1 (N6357, N6340);
not NOT1 (N6358, N6350);
and AND2 (N6359, N6351, N487);
nand NAND3 (N6360, N6356, N4778, N194);
xor XOR2 (N6361, N6357, N1246);
nor NOR3 (N6362, N6361, N584, N2567);
nand NAND4 (N6363, N6360, N1519, N4221, N2396);
and AND2 (N6364, N6362, N3489);
not NOT1 (N6365, N6347);
nor NOR2 (N6366, N6365, N2751);
xor XOR2 (N6367, N6359, N2842);
and AND3 (N6368, N6355, N4499, N5479);
not NOT1 (N6369, N6364);
nor NOR4 (N6370, N6368, N4909, N4517, N2182);
buf BUF1 (N6371, N6346);
nor NOR2 (N6372, N6367, N2679);
not NOT1 (N6373, N6370);
and AND4 (N6374, N6372, N5705, N4849, N6008);
and AND2 (N6375, N6369, N5301);
nand NAND2 (N6376, N6371, N5503);
nor NOR4 (N6377, N6363, N5669, N5154, N3701);
not NOT1 (N6378, N6376);
nor NOR3 (N6379, N6354, N1982, N459);
not NOT1 (N6380, N6374);
buf BUF1 (N6381, N6375);
nor NOR2 (N6382, N6379, N3658);
or OR4 (N6383, N6377, N2080, N2334, N5228);
buf BUF1 (N6384, N6381);
nand NAND2 (N6385, N6382, N10);
nand NAND3 (N6386, N6353, N845, N2469);
and AND4 (N6387, N6386, N3277, N6055, N5183);
buf BUF1 (N6388, N6358);
xor XOR2 (N6389, N6366, N1723);
nor NOR2 (N6390, N6380, N678);
buf BUF1 (N6391, N6383);
not NOT1 (N6392, N6332);
not NOT1 (N6393, N6392);
nand NAND2 (N6394, N6385, N5080);
or OR3 (N6395, N6373, N3661, N4926);
buf BUF1 (N6396, N6395);
and AND3 (N6397, N6393, N3097, N1667);
xor XOR2 (N6398, N6389, N4036);
or OR2 (N6399, N6387, N1457);
nand NAND2 (N6400, N6398, N5728);
nand NAND3 (N6401, N6399, N1034, N5291);
not NOT1 (N6402, N6401);
not NOT1 (N6403, N6391);
nor NOR2 (N6404, N6402, N283);
buf BUF1 (N6405, N6397);
xor XOR2 (N6406, N6404, N514);
xor XOR2 (N6407, N6388, N535);
buf BUF1 (N6408, N6400);
not NOT1 (N6409, N6407);
nor NOR4 (N6410, N6408, N549, N1203, N3561);
and AND3 (N6411, N6410, N2324, N6061);
or OR3 (N6412, N6378, N517, N2138);
xor XOR2 (N6413, N6405, N5662);
xor XOR2 (N6414, N6412, N2392);
nor NOR3 (N6415, N6403, N5342, N1871);
nor NOR4 (N6416, N6411, N4483, N4094, N2649);
not NOT1 (N6417, N6394);
or OR4 (N6418, N6414, N1316, N5463, N4212);
nor NOR2 (N6419, N6390, N458);
nor NOR2 (N6420, N6396, N436);
not NOT1 (N6421, N6420);
buf BUF1 (N6422, N6409);
xor XOR2 (N6423, N6415, N2705);
or OR4 (N6424, N6418, N5691, N556, N3420);
or OR4 (N6425, N6416, N4304, N2054, N559);
nor NOR4 (N6426, N6423, N908, N5757, N1242);
nand NAND2 (N6427, N6424, N6304);
and AND2 (N6428, N6419, N4133);
xor XOR2 (N6429, N6428, N3388);
or OR4 (N6430, N6413, N726, N714, N4054);
xor XOR2 (N6431, N6384, N1666);
nor NOR2 (N6432, N6430, N5662);
nor NOR3 (N6433, N6425, N426, N3292);
buf BUF1 (N6434, N6417);
buf BUF1 (N6435, N6422);
not NOT1 (N6436, N6406);
nand NAND2 (N6437, N6421, N2683);
or OR4 (N6438, N6436, N71, N4375, N5077);
and AND4 (N6439, N6426, N4018, N2707, N2967);
or OR4 (N6440, N6429, N3884, N5918, N249);
xor XOR2 (N6441, N6432, N2356);
or OR4 (N6442, N6427, N4319, N2795, N1688);
xor XOR2 (N6443, N6441, N3096);
nor NOR4 (N6444, N6443, N754, N2099, N3874);
xor XOR2 (N6445, N6434, N3464);
or OR2 (N6446, N6444, N4624);
buf BUF1 (N6447, N6442);
nand NAND4 (N6448, N6437, N4293, N1968, N821);
and AND3 (N6449, N6440, N1439, N205);
xor XOR2 (N6450, N6435, N2340);
not NOT1 (N6451, N6446);
nor NOR3 (N6452, N6445, N1262, N4717);
and AND4 (N6453, N6448, N3025, N5642, N5676);
or OR2 (N6454, N6451, N719);
or OR4 (N6455, N6447, N5401, N3460, N6328);
or OR3 (N6456, N6438, N502, N2803);
xor XOR2 (N6457, N6453, N2332);
or OR3 (N6458, N6456, N5588, N5663);
and AND3 (N6459, N6433, N105, N5262);
xor XOR2 (N6460, N6459, N2952);
and AND2 (N6461, N6450, N4678);
buf BUF1 (N6462, N6431);
not NOT1 (N6463, N6452);
and AND3 (N6464, N6463, N955, N2958);
xor XOR2 (N6465, N6449, N2057);
buf BUF1 (N6466, N6464);
nand NAND4 (N6467, N6457, N6167, N120, N5870);
buf BUF1 (N6468, N6467);
or OR3 (N6469, N6458, N3929, N3963);
nand NAND2 (N6470, N6439, N2601);
nand NAND4 (N6471, N6460, N690, N2325, N6380);
and AND2 (N6472, N6455, N2489);
not NOT1 (N6473, N6471);
not NOT1 (N6474, N6465);
nor NOR2 (N6475, N6469, N914);
nand NAND2 (N6476, N6474, N16);
not NOT1 (N6477, N6461);
not NOT1 (N6478, N6462);
buf BUF1 (N6479, N6454);
and AND4 (N6480, N6479, N3043, N1202, N4231);
not NOT1 (N6481, N6470);
nand NAND2 (N6482, N6466, N2155);
nor NOR3 (N6483, N6473, N1065, N3811);
buf BUF1 (N6484, N6483);
nor NOR3 (N6485, N6468, N4544, N2366);
xor XOR2 (N6486, N6478, N5846);
or OR2 (N6487, N6486, N3189);
and AND4 (N6488, N6480, N4113, N2817, N5219);
not NOT1 (N6489, N6484);
xor XOR2 (N6490, N6488, N2058);
xor XOR2 (N6491, N6485, N6112);
nand NAND4 (N6492, N6481, N1198, N4591, N2199);
or OR3 (N6493, N6477, N699, N3199);
nor NOR4 (N6494, N6476, N3697, N1574, N1266);
nand NAND2 (N6495, N6487, N2012);
nor NOR4 (N6496, N6495, N6430, N4006, N1481);
or OR3 (N6497, N6494, N1070, N3755);
xor XOR2 (N6498, N6491, N588);
buf BUF1 (N6499, N6498);
buf BUF1 (N6500, N6492);
not NOT1 (N6501, N6496);
nand NAND4 (N6502, N6499, N3234, N1301, N3966);
or OR2 (N6503, N6502, N4422);
and AND3 (N6504, N6475, N4424, N4587);
nand NAND3 (N6505, N6489, N651, N2428);
nor NOR4 (N6506, N6493, N4210, N5720, N2995);
nor NOR3 (N6507, N6504, N6048, N5812);
buf BUF1 (N6508, N6507);
and AND3 (N6509, N6503, N293, N3429);
xor XOR2 (N6510, N6490, N3909);
and AND2 (N6511, N6500, N687);
not NOT1 (N6512, N6506);
or OR2 (N6513, N6510, N5131);
buf BUF1 (N6514, N6472);
nor NOR2 (N6515, N6514, N1155);
nand NAND3 (N6516, N6508, N6248, N5854);
not NOT1 (N6517, N6497);
and AND2 (N6518, N6501, N2998);
or OR2 (N6519, N6509, N10);
nand NAND2 (N6520, N6512, N1737);
and AND2 (N6521, N6516, N1164);
or OR3 (N6522, N6505, N4723, N993);
or OR3 (N6523, N6517, N613, N3125);
nand NAND4 (N6524, N6520, N2111, N3829, N6029);
nor NOR2 (N6525, N6522, N3532);
or OR2 (N6526, N6513, N4818);
nand NAND4 (N6527, N6511, N269, N6109, N3687);
buf BUF1 (N6528, N6527);
xor XOR2 (N6529, N6525, N5347);
nor NOR3 (N6530, N6482, N3146, N5502);
xor XOR2 (N6531, N6529, N4830);
not NOT1 (N6532, N6521);
nand NAND2 (N6533, N6526, N2131);
xor XOR2 (N6534, N6531, N4818);
nand NAND3 (N6535, N6515, N2079, N4170);
nand NAND2 (N6536, N6530, N2850);
nand NAND4 (N6537, N6518, N113, N2060, N12);
and AND2 (N6538, N6535, N5290);
and AND3 (N6539, N6538, N1244, N1323);
and AND3 (N6540, N6534, N254, N465);
nand NAND2 (N6541, N6519, N5969);
buf BUF1 (N6542, N6539);
xor XOR2 (N6543, N6523, N6075);
xor XOR2 (N6544, N6540, N3633);
nand NAND2 (N6545, N6537, N1776);
or OR3 (N6546, N6543, N6417, N5338);
nor NOR2 (N6547, N6541, N477);
buf BUF1 (N6548, N6545);
not NOT1 (N6549, N6536);
nor NOR4 (N6550, N6542, N3276, N6364, N5531);
xor XOR2 (N6551, N6532, N1132);
xor XOR2 (N6552, N6551, N3342);
and AND2 (N6553, N6549, N3166);
buf BUF1 (N6554, N6547);
and AND4 (N6555, N6528, N1155, N3537, N5654);
nand NAND2 (N6556, N6533, N4633);
buf BUF1 (N6557, N6552);
or OR3 (N6558, N6524, N3738, N705);
and AND4 (N6559, N6548, N2360, N3316, N2640);
and AND3 (N6560, N6544, N667, N3252);
and AND3 (N6561, N6556, N2099, N4330);
nor NOR4 (N6562, N6561, N4369, N2562, N3042);
nor NOR4 (N6563, N6560, N4029, N4796, N957);
buf BUF1 (N6564, N6554);
nor NOR3 (N6565, N6557, N3997, N3007);
and AND2 (N6566, N6565, N3325);
not NOT1 (N6567, N6558);
or OR2 (N6568, N6566, N5603);
xor XOR2 (N6569, N6546, N179);
xor XOR2 (N6570, N6567, N4240);
buf BUF1 (N6571, N6563);
not NOT1 (N6572, N6568);
or OR3 (N6573, N6569, N3930, N4996);
not NOT1 (N6574, N6559);
nand NAND2 (N6575, N6564, N3928);
nand NAND4 (N6576, N6570, N3565, N1610, N2905);
nand NAND2 (N6577, N6573, N1269);
and AND4 (N6578, N6550, N2586, N4514, N2164);
nand NAND4 (N6579, N6562, N2522, N1787, N4869);
or OR2 (N6580, N6577, N4954);
nand NAND2 (N6581, N6574, N147);
nand NAND4 (N6582, N6575, N4597, N4339, N1124);
or OR4 (N6583, N6555, N604, N2517, N5390);
not NOT1 (N6584, N6553);
and AND2 (N6585, N6571, N4363);
buf BUF1 (N6586, N6581);
and AND4 (N6587, N6579, N2720, N2352, N3760);
and AND4 (N6588, N6572, N2780, N1546, N5591);
and AND4 (N6589, N6582, N4377, N3380, N6437);
or OR3 (N6590, N6588, N6232, N4464);
xor XOR2 (N6591, N6587, N1053);
xor XOR2 (N6592, N6576, N6245);
xor XOR2 (N6593, N6584, N1124);
xor XOR2 (N6594, N6591, N771);
buf BUF1 (N6595, N6593);
nor NOR3 (N6596, N6583, N1353, N4221);
or OR2 (N6597, N6586, N1716);
and AND4 (N6598, N6597, N1064, N2108, N922);
and AND3 (N6599, N6592, N5726, N1820);
nand NAND4 (N6600, N6590, N3385, N4296, N5851);
xor XOR2 (N6601, N6578, N6456);
buf BUF1 (N6602, N6595);
buf BUF1 (N6603, N6602);
buf BUF1 (N6604, N6603);
buf BUF1 (N6605, N6580);
nor NOR4 (N6606, N6585, N5710, N2219, N5718);
nand NAND3 (N6607, N6600, N764, N1060);
or OR3 (N6608, N6598, N5439, N4327);
xor XOR2 (N6609, N6599, N258);
nand NAND2 (N6610, N6608, N1686);
buf BUF1 (N6611, N6610);
or OR4 (N6612, N6589, N2251, N3228, N4766);
nor NOR4 (N6613, N6607, N4040, N1477, N597);
or OR4 (N6614, N6612, N6341, N1034, N6128);
nor NOR3 (N6615, N6601, N2949, N1233);
xor XOR2 (N6616, N6611, N5457);
xor XOR2 (N6617, N6605, N482);
buf BUF1 (N6618, N6613);
and AND3 (N6619, N6594, N5892, N3532);
buf BUF1 (N6620, N6606);
or OR3 (N6621, N6619, N3750, N2329);
and AND2 (N6622, N6621, N5674);
xor XOR2 (N6623, N6618, N3512);
nor NOR2 (N6624, N6604, N4429);
and AND3 (N6625, N6622, N6361, N2996);
not NOT1 (N6626, N6609);
xor XOR2 (N6627, N6616, N3907);
nor NOR3 (N6628, N6623, N5940, N835);
buf BUF1 (N6629, N6626);
buf BUF1 (N6630, N6617);
or OR4 (N6631, N6630, N1991, N5662, N4001);
nor NOR4 (N6632, N6629, N5098, N6572, N6467);
buf BUF1 (N6633, N6632);
or OR3 (N6634, N6615, N861, N302);
buf BUF1 (N6635, N6596);
or OR2 (N6636, N6631, N5207);
or OR2 (N6637, N6620, N1746);
and AND3 (N6638, N6636, N4942, N3477);
buf BUF1 (N6639, N6638);
not NOT1 (N6640, N6614);
xor XOR2 (N6641, N6633, N4845);
and AND3 (N6642, N6641, N5213, N5086);
or OR4 (N6643, N6642, N2670, N3606, N3726);
xor XOR2 (N6644, N6640, N710);
buf BUF1 (N6645, N6643);
nand NAND4 (N6646, N6634, N6538, N6468, N2284);
nand NAND2 (N6647, N6644, N5696);
nand NAND4 (N6648, N6645, N4766, N895, N312);
xor XOR2 (N6649, N6625, N523);
not NOT1 (N6650, N6648);
and AND3 (N6651, N6649, N5836, N2654);
and AND3 (N6652, N6635, N4335, N2262);
and AND2 (N6653, N6637, N1243);
nand NAND4 (N6654, N6639, N238, N408, N4997);
nand NAND4 (N6655, N6647, N954, N2487, N3619);
not NOT1 (N6656, N6654);
xor XOR2 (N6657, N6655, N4266);
nand NAND4 (N6658, N6652, N2556, N5596, N3116);
nor NOR3 (N6659, N6657, N6447, N3028);
nand NAND3 (N6660, N6646, N3887, N6633);
and AND3 (N6661, N6650, N3641, N2055);
nor NOR2 (N6662, N6659, N1271);
not NOT1 (N6663, N6661);
buf BUF1 (N6664, N6662);
xor XOR2 (N6665, N6624, N4373);
not NOT1 (N6666, N6628);
nor NOR2 (N6667, N6653, N5979);
nor NOR4 (N6668, N6651, N1940, N3495, N5167);
buf BUF1 (N6669, N6663);
xor XOR2 (N6670, N6668, N5467);
not NOT1 (N6671, N6669);
not NOT1 (N6672, N6656);
xor XOR2 (N6673, N6672, N6601);
nor NOR3 (N6674, N6664, N3395, N5921);
nor NOR4 (N6675, N6671, N3184, N1021, N434);
buf BUF1 (N6676, N6674);
and AND2 (N6677, N6627, N5828);
nand NAND4 (N6678, N6670, N2749, N334, N3496);
or OR4 (N6679, N6667, N4578, N4800, N4963);
xor XOR2 (N6680, N6678, N1316);
not NOT1 (N6681, N6673);
nor NOR4 (N6682, N6677, N2019, N4423, N4163);
and AND3 (N6683, N6682, N6635, N3881);
or OR2 (N6684, N6681, N2528);
or OR3 (N6685, N6680, N6503, N1573);
and AND3 (N6686, N6676, N3542, N1334);
or OR4 (N6687, N6665, N5659, N4499, N1043);
or OR3 (N6688, N6666, N6504, N2085);
xor XOR2 (N6689, N6686, N4244);
and AND3 (N6690, N6685, N5640, N1005);
not NOT1 (N6691, N6660);
nor NOR2 (N6692, N6691, N2467);
nor NOR3 (N6693, N6690, N1350, N711);
or OR4 (N6694, N6675, N5387, N5985, N2187);
not NOT1 (N6695, N6684);
nor NOR3 (N6696, N6679, N3095, N5620);
not NOT1 (N6697, N6688);
buf BUF1 (N6698, N6693);
not NOT1 (N6699, N6697);
nand NAND3 (N6700, N6694, N2706, N2699);
and AND3 (N6701, N6695, N2569, N6213);
nor NOR4 (N6702, N6689, N1584, N2919, N4834);
nor NOR2 (N6703, N6683, N6603);
nor NOR2 (N6704, N6699, N4807);
nor NOR2 (N6705, N6700, N4179);
xor XOR2 (N6706, N6658, N5948);
xor XOR2 (N6707, N6696, N1454);
buf BUF1 (N6708, N6687);
not NOT1 (N6709, N6701);
buf BUF1 (N6710, N6703);
and AND3 (N6711, N6702, N1958, N580);
nand NAND4 (N6712, N6706, N379, N4105, N2691);
nor NOR3 (N6713, N6711, N3473, N795);
nand NAND3 (N6714, N6698, N4456, N3858);
nand NAND3 (N6715, N6692, N4279, N4227);
and AND3 (N6716, N6714, N3870, N2778);
and AND3 (N6717, N6704, N1579, N4357);
not NOT1 (N6718, N6716);
not NOT1 (N6719, N6715);
nor NOR4 (N6720, N6713, N3489, N5095, N5887);
xor XOR2 (N6721, N6709, N1829);
xor XOR2 (N6722, N6719, N278);
not NOT1 (N6723, N6720);
nor NOR4 (N6724, N6717, N3339, N4234, N3215);
nand NAND4 (N6725, N6712, N4244, N6293, N5596);
xor XOR2 (N6726, N6707, N5499);
or OR2 (N6727, N6722, N527);
xor XOR2 (N6728, N6723, N2054);
or OR2 (N6729, N6726, N119);
nand NAND2 (N6730, N6728, N1551);
nor NOR3 (N6731, N6708, N4027, N1502);
nand NAND3 (N6732, N6705, N5222, N3362);
not NOT1 (N6733, N6710);
or OR3 (N6734, N6721, N2527, N4766);
buf BUF1 (N6735, N6732);
buf BUF1 (N6736, N6727);
xor XOR2 (N6737, N6729, N4941);
not NOT1 (N6738, N6735);
and AND3 (N6739, N6734, N2860, N975);
not NOT1 (N6740, N6725);
and AND4 (N6741, N6733, N1914, N2426, N5846);
nor NOR2 (N6742, N6730, N1050);
nand NAND4 (N6743, N6739, N3817, N6512, N1489);
buf BUF1 (N6744, N6718);
or OR3 (N6745, N6741, N5453, N344);
or OR2 (N6746, N6731, N3312);
xor XOR2 (N6747, N6736, N5661);
and AND2 (N6748, N6747, N1013);
buf BUF1 (N6749, N6744);
xor XOR2 (N6750, N6746, N1791);
or OR2 (N6751, N6749, N4388);
and AND2 (N6752, N6745, N6296);
xor XOR2 (N6753, N6748, N5483);
xor XOR2 (N6754, N6737, N5637);
not NOT1 (N6755, N6740);
nand NAND2 (N6756, N6755, N751);
xor XOR2 (N6757, N6750, N6209);
buf BUF1 (N6758, N6724);
nand NAND2 (N6759, N6738, N2942);
nand NAND4 (N6760, N6742, N134, N4584, N1654);
not NOT1 (N6761, N6751);
nand NAND2 (N6762, N6760, N4136);
buf BUF1 (N6763, N6743);
xor XOR2 (N6764, N6756, N95);
nor NOR3 (N6765, N6757, N438, N1220);
xor XOR2 (N6766, N6759, N2696);
buf BUF1 (N6767, N6754);
xor XOR2 (N6768, N6764, N4576);
not NOT1 (N6769, N6753);
not NOT1 (N6770, N6758);
not NOT1 (N6771, N6752);
nand NAND4 (N6772, N6763, N4589, N5081, N5718);
nor NOR3 (N6773, N6772, N2068, N5551);
or OR3 (N6774, N6765, N5218, N5906);
not NOT1 (N6775, N6773);
nand NAND3 (N6776, N6766, N5062, N4496);
nand NAND4 (N6777, N6769, N93, N1129, N2697);
or OR3 (N6778, N6776, N2148, N5830);
buf BUF1 (N6779, N6775);
buf BUF1 (N6780, N6778);
not NOT1 (N6781, N6768);
and AND3 (N6782, N6770, N5293, N790);
xor XOR2 (N6783, N6779, N1838);
xor XOR2 (N6784, N6774, N1094);
nand NAND4 (N6785, N6767, N2441, N4432, N6559);
or OR3 (N6786, N6761, N5030, N5245);
or OR3 (N6787, N6783, N6232, N4957);
buf BUF1 (N6788, N6780);
xor XOR2 (N6789, N6762, N3509);
nor NOR4 (N6790, N6786, N4705, N1582, N336);
and AND2 (N6791, N6777, N367);
not NOT1 (N6792, N6787);
not NOT1 (N6793, N6789);
or OR4 (N6794, N6784, N2372, N1028, N921);
buf BUF1 (N6795, N6791);
not NOT1 (N6796, N6771);
nand NAND2 (N6797, N6795, N6456);
and AND2 (N6798, N6790, N5675);
not NOT1 (N6799, N6792);
nand NAND2 (N6800, N6782, N734);
xor XOR2 (N6801, N6799, N4433);
buf BUF1 (N6802, N6798);
nor NOR2 (N6803, N6788, N1931);
and AND4 (N6804, N6801, N2565, N839, N6799);
nor NOR4 (N6805, N6802, N1592, N4738, N3738);
nor NOR4 (N6806, N6794, N6800, N811, N5577);
not NOT1 (N6807, N1579);
not NOT1 (N6808, N6793);
buf BUF1 (N6809, N6803);
not NOT1 (N6810, N6807);
not NOT1 (N6811, N6805);
or OR3 (N6812, N6811, N3408, N4622);
or OR4 (N6813, N6810, N993, N6497, N1052);
buf BUF1 (N6814, N6813);
not NOT1 (N6815, N6808);
nand NAND3 (N6816, N6781, N6417, N5720);
or OR2 (N6817, N6809, N6010);
and AND3 (N6818, N6806, N4744, N87);
buf BUF1 (N6819, N6816);
nand NAND4 (N6820, N6815, N6228, N3819, N5354);
nand NAND4 (N6821, N6812, N722, N5711, N644);
nor NOR2 (N6822, N6821, N6084);
not NOT1 (N6823, N6804);
and AND2 (N6824, N6817, N4287);
buf BUF1 (N6825, N6819);
nand NAND3 (N6826, N6824, N2893, N582);
not NOT1 (N6827, N6823);
xor XOR2 (N6828, N6796, N320);
nand NAND2 (N6829, N6820, N3102);
nand NAND4 (N6830, N6822, N5075, N2980, N143);
not NOT1 (N6831, N6827);
buf BUF1 (N6832, N6826);
buf BUF1 (N6833, N6829);
nand NAND4 (N6834, N6831, N3840, N560, N2285);
nand NAND3 (N6835, N6814, N1102, N5867);
nand NAND4 (N6836, N6834, N6744, N4952, N5349);
or OR3 (N6837, N6830, N4470, N4502);
or OR2 (N6838, N6832, N6106);
buf BUF1 (N6839, N6785);
buf BUF1 (N6840, N6833);
xor XOR2 (N6841, N6840, N1701);
or OR2 (N6842, N6841, N5883);
or OR2 (N6843, N6825, N4385);
xor XOR2 (N6844, N6797, N2297);
xor XOR2 (N6845, N6838, N4977);
nand NAND4 (N6846, N6837, N1454, N4518, N5590);
nand NAND2 (N6847, N6836, N2518);
nand NAND4 (N6848, N6842, N2218, N664, N4722);
buf BUF1 (N6849, N6835);
and AND2 (N6850, N6847, N331);
nand NAND2 (N6851, N6846, N6071);
not NOT1 (N6852, N6839);
xor XOR2 (N6853, N6851, N2545);
not NOT1 (N6854, N6843);
or OR2 (N6855, N6848, N744);
xor XOR2 (N6856, N6855, N255);
and AND3 (N6857, N6845, N383, N4200);
nor NOR3 (N6858, N6857, N278, N2991);
not NOT1 (N6859, N6818);
nand NAND2 (N6860, N6828, N1732);
or OR3 (N6861, N6856, N87, N2006);
nor NOR3 (N6862, N6849, N2769, N4758);
nor NOR3 (N6863, N6859, N6856, N112);
nand NAND3 (N6864, N6863, N1941, N1286);
or OR3 (N6865, N6852, N782, N6633);
and AND3 (N6866, N6864, N4361, N2887);
and AND3 (N6867, N6854, N638, N4167);
buf BUF1 (N6868, N6862);
and AND3 (N6869, N6868, N4107, N1143);
nand NAND3 (N6870, N6850, N287, N1649);
buf BUF1 (N6871, N6867);
xor XOR2 (N6872, N6869, N888);
xor XOR2 (N6873, N6866, N1277);
xor XOR2 (N6874, N6873, N4844);
and AND4 (N6875, N6844, N4260, N1091, N1867);
buf BUF1 (N6876, N6875);
or OR3 (N6877, N6871, N6115, N5312);
nand NAND4 (N6878, N6858, N4937, N438, N870);
xor XOR2 (N6879, N6865, N1570);
nor NOR2 (N6880, N6876, N2178);
buf BUF1 (N6881, N6877);
and AND4 (N6882, N6872, N6749, N4893, N3541);
not NOT1 (N6883, N6880);
xor XOR2 (N6884, N6860, N142);
or OR3 (N6885, N6882, N6109, N833);
not NOT1 (N6886, N6881);
and AND3 (N6887, N6861, N4319, N3926);
nand NAND2 (N6888, N6878, N582);
and AND3 (N6889, N6887, N2486, N5371);
or OR4 (N6890, N6885, N2742, N449, N6270);
nand NAND3 (N6891, N6879, N2817, N3076);
nand NAND3 (N6892, N6889, N5613, N6272);
not NOT1 (N6893, N6886);
xor XOR2 (N6894, N6888, N5143);
and AND4 (N6895, N6893, N3508, N5990, N384);
buf BUF1 (N6896, N6890);
not NOT1 (N6897, N6853);
nor NOR3 (N6898, N6896, N2558, N3);
buf BUF1 (N6899, N6891);
xor XOR2 (N6900, N6884, N3080);
xor XOR2 (N6901, N6895, N754);
xor XOR2 (N6902, N6898, N2797);
nor NOR3 (N6903, N6894, N6640, N5158);
or OR3 (N6904, N6897, N5767, N779);
or OR3 (N6905, N6883, N4173, N3345);
nor NOR3 (N6906, N6903, N2995, N6601);
and AND4 (N6907, N6902, N2253, N835, N3003);
buf BUF1 (N6908, N6906);
buf BUF1 (N6909, N6900);
or OR2 (N6910, N6870, N2709);
buf BUF1 (N6911, N6910);
or OR3 (N6912, N6911, N2363, N502);
or OR2 (N6913, N6892, N132);
buf BUF1 (N6914, N6912);
xor XOR2 (N6915, N6904, N1296);
and AND3 (N6916, N6915, N3191, N3169);
not NOT1 (N6917, N6908);
nor NOR4 (N6918, N6917, N944, N3761, N4707);
xor XOR2 (N6919, N6874, N6178);
not NOT1 (N6920, N6899);
not NOT1 (N6921, N6919);
or OR4 (N6922, N6901, N5185, N4726, N6323);
xor XOR2 (N6923, N6913, N3361);
buf BUF1 (N6924, N6916);
not NOT1 (N6925, N6920);
buf BUF1 (N6926, N6907);
buf BUF1 (N6927, N6905);
buf BUF1 (N6928, N6926);
nor NOR4 (N6929, N6925, N1814, N2665, N259);
buf BUF1 (N6930, N6921);
xor XOR2 (N6931, N6923, N1865);
or OR4 (N6932, N6914, N6154, N1143, N6144);
or OR2 (N6933, N6930, N4902);
xor XOR2 (N6934, N6929, N5476);
or OR3 (N6935, N6909, N5667, N5317);
not NOT1 (N6936, N6931);
and AND3 (N6937, N6935, N5950, N1113);
nor NOR4 (N6938, N6928, N6350, N3588, N6395);
nor NOR4 (N6939, N6932, N5204, N3100, N1519);
buf BUF1 (N6940, N6937);
not NOT1 (N6941, N6933);
nand NAND4 (N6942, N6934, N2308, N5992, N1312);
or OR2 (N6943, N6922, N1480);
not NOT1 (N6944, N6938);
and AND4 (N6945, N6924, N61, N6367, N5638);
buf BUF1 (N6946, N6936);
buf BUF1 (N6947, N6944);
xor XOR2 (N6948, N6941, N5584);
not NOT1 (N6949, N6918);
or OR2 (N6950, N6942, N2442);
nor NOR4 (N6951, N6947, N1735, N2954, N651);
not NOT1 (N6952, N6939);
xor XOR2 (N6953, N6951, N6639);
or OR3 (N6954, N6940, N1612, N1929);
xor XOR2 (N6955, N6945, N6589);
xor XOR2 (N6956, N6953, N1688);
buf BUF1 (N6957, N6952);
or OR3 (N6958, N6956, N1068, N1505);
not NOT1 (N6959, N6943);
and AND3 (N6960, N6957, N2246, N4476);
nor NOR3 (N6961, N6955, N3348, N6617);
nand NAND2 (N6962, N6954, N729);
xor XOR2 (N6963, N6949, N2271);
xor XOR2 (N6964, N6962, N1744);
and AND4 (N6965, N6958, N1543, N3794, N1093);
xor XOR2 (N6966, N6950, N6914);
and AND4 (N6967, N6927, N1373, N4360, N5148);
xor XOR2 (N6968, N6959, N6276);
and AND2 (N6969, N6963, N252);
not NOT1 (N6970, N6961);
not NOT1 (N6971, N6965);
or OR2 (N6972, N6966, N2161);
nor NOR2 (N6973, N6970, N732);
nand NAND3 (N6974, N6964, N3396, N6400);
xor XOR2 (N6975, N6967, N2580);
nor NOR4 (N6976, N6972, N5714, N1206, N4857);
and AND2 (N6977, N6976, N5906);
and AND3 (N6978, N6973, N6174, N3919);
nor NOR3 (N6979, N6978, N263, N2423);
not NOT1 (N6980, N6946);
xor XOR2 (N6981, N6977, N831);
or OR4 (N6982, N6975, N2883, N5442, N2451);
xor XOR2 (N6983, N6979, N6117);
xor XOR2 (N6984, N6971, N10);
not NOT1 (N6985, N6983);
or OR4 (N6986, N6981, N727, N2954, N3103);
xor XOR2 (N6987, N6960, N6251);
xor XOR2 (N6988, N6982, N5622);
not NOT1 (N6989, N6985);
buf BUF1 (N6990, N6986);
buf BUF1 (N6991, N6987);
xor XOR2 (N6992, N6988, N3165);
buf BUF1 (N6993, N6991);
not NOT1 (N6994, N6948);
nor NOR4 (N6995, N6969, N5230, N3209, N5703);
not NOT1 (N6996, N6984);
or OR2 (N6997, N6995, N2183);
buf BUF1 (N6998, N6997);
xor XOR2 (N6999, N6990, N3042);
nor NOR3 (N7000, N6989, N6911, N1114);
nand NAND3 (N7001, N6999, N5745, N6356);
buf BUF1 (N7002, N6992);
xor XOR2 (N7003, N7001, N4557);
or OR4 (N7004, N7003, N6326, N1284, N6957);
or OR2 (N7005, N7000, N6976);
and AND4 (N7006, N6993, N3969, N4835, N1298);
not NOT1 (N7007, N6968);
not NOT1 (N7008, N6996);
buf BUF1 (N7009, N7006);
and AND4 (N7010, N7005, N2189, N2841, N5332);
nand NAND2 (N7011, N7010, N3304);
nand NAND4 (N7012, N7002, N2297, N4757, N5873);
and AND3 (N7013, N7009, N167, N6109);
nor NOR2 (N7014, N6994, N5260);
xor XOR2 (N7015, N6974, N3111);
buf BUF1 (N7016, N7013);
buf BUF1 (N7017, N7008);
and AND3 (N7018, N6980, N2015, N6618);
not NOT1 (N7019, N7016);
buf BUF1 (N7020, N7004);
buf BUF1 (N7021, N7015);
nor NOR4 (N7022, N7014, N6373, N3011, N5701);
xor XOR2 (N7023, N7018, N4694);
not NOT1 (N7024, N7022);
and AND4 (N7025, N7024, N299, N6467, N5147);
and AND2 (N7026, N6998, N5579);
buf BUF1 (N7027, N7019);
not NOT1 (N7028, N7027);
not NOT1 (N7029, N7025);
nor NOR4 (N7030, N7012, N6708, N3678, N4992);
nand NAND4 (N7031, N7030, N1973, N1171, N5654);
buf BUF1 (N7032, N7017);
not NOT1 (N7033, N7023);
nand NAND4 (N7034, N7011, N6867, N1020, N631);
xor XOR2 (N7035, N7032, N256);
nand NAND4 (N7036, N7031, N4528, N6390, N853);
buf BUF1 (N7037, N7029);
nand NAND3 (N7038, N7021, N119, N4313);
buf BUF1 (N7039, N7020);
nor NOR3 (N7040, N7036, N832, N6986);
not NOT1 (N7041, N7038);
or OR4 (N7042, N7028, N1367, N3352, N30);
xor XOR2 (N7043, N7007, N963);
nor NOR4 (N7044, N7042, N4719, N3762, N6031);
and AND4 (N7045, N7043, N6949, N6984, N2080);
not NOT1 (N7046, N7037);
nor NOR2 (N7047, N7026, N4504);
or OR2 (N7048, N7046, N5604);
buf BUF1 (N7049, N7041);
nand NAND4 (N7050, N7033, N116, N2369, N4730);
nand NAND4 (N7051, N7049, N5026, N6110, N3087);
or OR4 (N7052, N7047, N981, N5734, N4923);
nand NAND3 (N7053, N7040, N1179, N3307);
not NOT1 (N7054, N7053);
buf BUF1 (N7055, N7045);
nor NOR2 (N7056, N7044, N6727);
xor XOR2 (N7057, N7039, N3536);
nor NOR4 (N7058, N7056, N6880, N612, N479);
not NOT1 (N7059, N7054);
and AND2 (N7060, N7057, N2295);
xor XOR2 (N7061, N7051, N2825);
nand NAND3 (N7062, N7058, N4692, N358);
buf BUF1 (N7063, N7048);
buf BUF1 (N7064, N7060);
not NOT1 (N7065, N7035);
or OR3 (N7066, N7034, N5373, N5343);
xor XOR2 (N7067, N7050, N1027);
or OR4 (N7068, N7052, N261, N21, N845);
and AND3 (N7069, N7061, N2974, N240);
nor NOR2 (N7070, N7069, N93);
and AND4 (N7071, N7070, N137, N6261, N2624);
not NOT1 (N7072, N7063);
not NOT1 (N7073, N7071);
buf BUF1 (N7074, N7072);
not NOT1 (N7075, N7064);
not NOT1 (N7076, N7065);
not NOT1 (N7077, N7055);
not NOT1 (N7078, N7074);
and AND3 (N7079, N7059, N2059, N2636);
not NOT1 (N7080, N7076);
buf BUF1 (N7081, N7062);
or OR4 (N7082, N7067, N3655, N7040, N493);
nand NAND4 (N7083, N7080, N2489, N2704, N37);
not NOT1 (N7084, N7077);
nor NOR4 (N7085, N7066, N810, N2559, N824);
xor XOR2 (N7086, N7075, N176);
and AND4 (N7087, N7083, N3190, N665, N7081);
not NOT1 (N7088, N1007);
nor NOR3 (N7089, N7087, N3002, N6298);
or OR4 (N7090, N7068, N1270, N1315, N6447);
or OR3 (N7091, N7085, N6816, N4704);
not NOT1 (N7092, N7073);
nand NAND4 (N7093, N7090, N3150, N6965, N2285);
not NOT1 (N7094, N7093);
or OR4 (N7095, N7091, N739, N6343, N549);
and AND4 (N7096, N7095, N5927, N2893, N1494);
and AND4 (N7097, N7086, N363, N3992, N4265);
and AND2 (N7098, N7084, N4089);
buf BUF1 (N7099, N7079);
xor XOR2 (N7100, N7088, N533);
or OR4 (N7101, N7100, N5809, N4149, N446);
or OR4 (N7102, N7101, N6874, N2655, N6460);
and AND3 (N7103, N7094, N1624, N6187);
nor NOR3 (N7104, N7103, N4513, N7001);
and AND2 (N7105, N7102, N3656);
not NOT1 (N7106, N7098);
nand NAND2 (N7107, N7082, N5006);
not NOT1 (N7108, N7078);
or OR2 (N7109, N7108, N7012);
nand NAND3 (N7110, N7107, N1051, N4180);
buf BUF1 (N7111, N7110);
not NOT1 (N7112, N7105);
nand NAND2 (N7113, N7089, N4112);
xor XOR2 (N7114, N7109, N2846);
and AND4 (N7115, N7096, N6335, N4649, N6818);
or OR2 (N7116, N7097, N4849);
nor NOR2 (N7117, N7115, N2747);
nor NOR4 (N7118, N7104, N361, N5574, N929);
nor NOR3 (N7119, N7111, N1096, N5850);
xor XOR2 (N7120, N7092, N320);
buf BUF1 (N7121, N7116);
or OR4 (N7122, N7117, N5157, N6099, N6032);
not NOT1 (N7123, N7106);
xor XOR2 (N7124, N7114, N4911);
or OR2 (N7125, N7119, N5241);
buf BUF1 (N7126, N7099);
or OR3 (N7127, N7118, N1032, N4840);
or OR4 (N7128, N7127, N6577, N2319, N6350);
nor NOR4 (N7129, N7121, N1450, N2418, N7031);
xor XOR2 (N7130, N7123, N3990);
buf BUF1 (N7131, N7122);
nand NAND3 (N7132, N7129, N2641, N864);
not NOT1 (N7133, N7131);
xor XOR2 (N7134, N7128, N5875);
nand NAND4 (N7135, N7132, N3183, N877, N6766);
not NOT1 (N7136, N7113);
nand NAND2 (N7137, N7133, N5532);
buf BUF1 (N7138, N7135);
or OR3 (N7139, N7130, N5557, N3192);
nand NAND3 (N7140, N7137, N4873, N3805);
nor NOR4 (N7141, N7112, N5560, N6263, N6403);
and AND3 (N7142, N7140, N741, N4943);
not NOT1 (N7143, N7139);
and AND2 (N7144, N7143, N1397);
nand NAND3 (N7145, N7136, N6529, N6214);
and AND3 (N7146, N7124, N5363, N2016);
nand NAND4 (N7147, N7146, N424, N3034, N2539);
xor XOR2 (N7148, N7147, N511);
buf BUF1 (N7149, N7138);
xor XOR2 (N7150, N7134, N1461);
xor XOR2 (N7151, N7142, N6605);
or OR3 (N7152, N7148, N3927, N5677);
not NOT1 (N7153, N7120);
and AND3 (N7154, N7153, N50, N1448);
nand NAND3 (N7155, N7126, N3405, N1529);
xor XOR2 (N7156, N7151, N5382);
not NOT1 (N7157, N7141);
nand NAND4 (N7158, N7156, N6489, N3462, N188);
buf BUF1 (N7159, N7154);
nand NAND4 (N7160, N7150, N2039, N280, N3420);
buf BUF1 (N7161, N7157);
nor NOR2 (N7162, N7125, N1303);
nand NAND4 (N7163, N7159, N3011, N822, N3591);
or OR3 (N7164, N7161, N4086, N5809);
buf BUF1 (N7165, N7164);
buf BUF1 (N7166, N7149);
or OR4 (N7167, N7152, N1184, N7163, N5334);
and AND2 (N7168, N1103, N6502);
xor XOR2 (N7169, N7168, N2152);
or OR3 (N7170, N7169, N3100, N4969);
or OR4 (N7171, N7155, N7158, N6704, N1754);
buf BUF1 (N7172, N6781);
buf BUF1 (N7173, N7165);
nand NAND4 (N7174, N7171, N6452, N1144, N6881);
and AND2 (N7175, N7162, N5136);
buf BUF1 (N7176, N7174);
and AND3 (N7177, N7172, N1958, N1821);
xor XOR2 (N7178, N7176, N1035);
buf BUF1 (N7179, N7175);
buf BUF1 (N7180, N7170);
nor NOR2 (N7181, N7180, N1330);
nor NOR4 (N7182, N7177, N273, N4960, N4170);
xor XOR2 (N7183, N7145, N3371);
buf BUF1 (N7184, N7160);
nor NOR3 (N7185, N7179, N2450, N40);
or OR4 (N7186, N7182, N6337, N5245, N1460);
and AND3 (N7187, N7178, N6449, N953);
xor XOR2 (N7188, N7185, N32);
or OR4 (N7189, N7187, N4738, N167, N2335);
nor NOR4 (N7190, N7144, N4481, N271, N682);
xor XOR2 (N7191, N7190, N1827);
and AND4 (N7192, N7183, N5634, N93, N1318);
or OR3 (N7193, N7166, N3064, N5501);
and AND3 (N7194, N7181, N1755, N5426);
nor NOR3 (N7195, N7191, N4496, N4217);
nand NAND3 (N7196, N7167, N6826, N4458);
buf BUF1 (N7197, N7173);
or OR2 (N7198, N7192, N1287);
nor NOR4 (N7199, N7186, N2055, N818, N4452);
or OR3 (N7200, N7193, N7022, N228);
nor NOR2 (N7201, N7196, N573);
nand NAND4 (N7202, N7184, N3756, N4308, N3049);
buf BUF1 (N7203, N7188);
not NOT1 (N7204, N7197);
xor XOR2 (N7205, N7202, N844);
and AND3 (N7206, N7200, N2595, N3923);
and AND3 (N7207, N7199, N3444, N3079);
not NOT1 (N7208, N7189);
nor NOR3 (N7209, N7206, N4618, N4080);
buf BUF1 (N7210, N7204);
or OR2 (N7211, N7209, N6782);
and AND4 (N7212, N7194, N588, N3341, N4437);
nor NOR3 (N7213, N7212, N5110, N5180);
or OR3 (N7214, N7213, N1963, N5433);
nor NOR4 (N7215, N7210, N3196, N7063, N240);
and AND3 (N7216, N7195, N4519, N2889);
nand NAND3 (N7217, N7201, N5103, N1121);
not NOT1 (N7218, N7217);
and AND3 (N7219, N7215, N2228, N1903);
buf BUF1 (N7220, N7214);
not NOT1 (N7221, N7218);
and AND4 (N7222, N7203, N1812, N6558, N5743);
nand NAND4 (N7223, N7222, N259, N702, N1453);
not NOT1 (N7224, N7205);
buf BUF1 (N7225, N7219);
or OR4 (N7226, N7224, N2343, N4870, N5447);
or OR4 (N7227, N7221, N6620, N4360, N633);
not NOT1 (N7228, N7208);
nand NAND2 (N7229, N7226, N4898);
buf BUF1 (N7230, N7229);
or OR3 (N7231, N7223, N5435, N1549);
nand NAND3 (N7232, N7225, N2969, N765);
buf BUF1 (N7233, N7228);
buf BUF1 (N7234, N7230);
buf BUF1 (N7235, N7207);
buf BUF1 (N7236, N7235);
nand NAND2 (N7237, N7211, N4344);
nand NAND2 (N7238, N7220, N6012);
xor XOR2 (N7239, N7231, N7072);
or OR2 (N7240, N7198, N6604);
or OR4 (N7241, N7234, N7193, N3890, N28);
xor XOR2 (N7242, N7238, N764);
not NOT1 (N7243, N7236);
buf BUF1 (N7244, N7240);
xor XOR2 (N7245, N7244, N6010);
nand NAND4 (N7246, N7241, N2911, N7189, N4632);
and AND2 (N7247, N7232, N3798);
buf BUF1 (N7248, N7246);
nand NAND3 (N7249, N7227, N4242, N5831);
nor NOR2 (N7250, N7239, N6327);
xor XOR2 (N7251, N7243, N2398);
nor NOR3 (N7252, N7248, N1048, N5137);
and AND2 (N7253, N7250, N6644);
xor XOR2 (N7254, N7242, N4933);
nor NOR4 (N7255, N7252, N7060, N1289, N2062);
nand NAND3 (N7256, N7237, N6758, N418);
buf BUF1 (N7257, N7247);
nor NOR4 (N7258, N7249, N1651, N3401, N373);
and AND2 (N7259, N7257, N5115);
not NOT1 (N7260, N7258);
or OR2 (N7261, N7251, N6237);
buf BUF1 (N7262, N7245);
not NOT1 (N7263, N7254);
and AND3 (N7264, N7263, N3676, N5843);
or OR2 (N7265, N7260, N6795);
and AND3 (N7266, N7262, N3272, N6464);
nor NOR4 (N7267, N7253, N1718, N6017, N2419);
nor NOR2 (N7268, N7216, N5130);
xor XOR2 (N7269, N7261, N4261);
nand NAND2 (N7270, N7256, N1041);
or OR4 (N7271, N7255, N1152, N1201, N3399);
nor NOR4 (N7272, N7269, N3750, N6378, N2806);
buf BUF1 (N7273, N7267);
nor NOR3 (N7274, N7271, N1708, N6482);
xor XOR2 (N7275, N7265, N1304);
xor XOR2 (N7276, N7270, N4461);
xor XOR2 (N7277, N7276, N7230);
and AND3 (N7278, N7272, N3319, N6104);
xor XOR2 (N7279, N7278, N1082);
buf BUF1 (N7280, N7274);
xor XOR2 (N7281, N7277, N6356);
buf BUF1 (N7282, N7233);
buf BUF1 (N7283, N7266);
buf BUF1 (N7284, N7275);
nand NAND4 (N7285, N7264, N1936, N1628, N2967);
nor NOR3 (N7286, N7285, N1233, N1119);
and AND2 (N7287, N7280, N3970);
xor XOR2 (N7288, N7273, N7000);
or OR3 (N7289, N7282, N6207, N503);
or OR4 (N7290, N7289, N4200, N2950, N4007);
or OR4 (N7291, N7288, N4637, N3726, N1272);
buf BUF1 (N7292, N7291);
buf BUF1 (N7293, N7279);
xor XOR2 (N7294, N7286, N5693);
xor XOR2 (N7295, N7281, N6538);
and AND2 (N7296, N7283, N2117);
nand NAND3 (N7297, N7296, N171, N7214);
nor NOR4 (N7298, N7287, N1623, N1695, N7204);
xor XOR2 (N7299, N7297, N6347);
nor NOR2 (N7300, N7294, N4982);
not NOT1 (N7301, N7298);
xor XOR2 (N7302, N7301, N6318);
or OR2 (N7303, N7284, N4519);
xor XOR2 (N7304, N7293, N6517);
and AND2 (N7305, N7303, N7216);
nor NOR2 (N7306, N7259, N6268);
and AND2 (N7307, N7306, N1211);
nor NOR3 (N7308, N7302, N1799, N1203);
nor NOR3 (N7309, N7307, N7219, N5603);
and AND4 (N7310, N7304, N3553, N1695, N5489);
buf BUF1 (N7311, N7300);
nor NOR3 (N7312, N7310, N3886, N707);
nand NAND3 (N7313, N7312, N6590, N6825);
and AND3 (N7314, N7268, N369, N525);
and AND3 (N7315, N7295, N4047, N3702);
and AND2 (N7316, N7313, N4905);
buf BUF1 (N7317, N7290);
buf BUF1 (N7318, N7316);
buf BUF1 (N7319, N7292);
or OR3 (N7320, N7309, N1796, N584);
and AND4 (N7321, N7319, N3594, N1830, N5919);
not NOT1 (N7322, N7317);
and AND2 (N7323, N7305, N4730);
buf BUF1 (N7324, N7321);
xor XOR2 (N7325, N7308, N1204);
xor XOR2 (N7326, N7320, N1910);
xor XOR2 (N7327, N7299, N6847);
and AND2 (N7328, N7315, N2547);
nand NAND3 (N7329, N7323, N735, N793);
xor XOR2 (N7330, N7314, N3184);
or OR4 (N7331, N7328, N639, N6899, N2089);
xor XOR2 (N7332, N7327, N2378);
or OR4 (N7333, N7324, N5262, N1577, N6251);
nor NOR3 (N7334, N7331, N7207, N7024);
nand NAND3 (N7335, N7330, N7004, N332);
xor XOR2 (N7336, N7325, N5795);
nand NAND3 (N7337, N7318, N7236, N3865);
xor XOR2 (N7338, N7332, N783);
xor XOR2 (N7339, N7326, N1676);
and AND4 (N7340, N7339, N5237, N1396, N567);
or OR3 (N7341, N7329, N6056, N7282);
and AND3 (N7342, N7333, N3495, N2417);
xor XOR2 (N7343, N7341, N6839);
or OR3 (N7344, N7337, N407, N6448);
and AND4 (N7345, N7334, N5530, N906, N5733);
not NOT1 (N7346, N7342);
nand NAND3 (N7347, N7338, N6926, N4718);
buf BUF1 (N7348, N7336);
nand NAND4 (N7349, N7343, N5845, N3126, N4885);
and AND4 (N7350, N7345, N2367, N543, N6415);
nor NOR4 (N7351, N7335, N1663, N5647, N6651);
not NOT1 (N7352, N7348);
and AND4 (N7353, N7349, N2576, N47, N750);
nand NAND2 (N7354, N7346, N6312);
and AND3 (N7355, N7354, N3095, N7094);
xor XOR2 (N7356, N7344, N661);
buf BUF1 (N7357, N7353);
nor NOR3 (N7358, N7322, N5404, N7248);
and AND4 (N7359, N7355, N5082, N4067, N1431);
nor NOR2 (N7360, N7350, N7317);
or OR2 (N7361, N7340, N5384);
xor XOR2 (N7362, N7351, N1642);
nor NOR2 (N7363, N7356, N2206);
and AND2 (N7364, N7311, N5604);
not NOT1 (N7365, N7359);
and AND2 (N7366, N7364, N1693);
nor NOR4 (N7367, N7360, N2681, N1368, N1231);
nor NOR4 (N7368, N7366, N3279, N432, N5017);
or OR4 (N7369, N7365, N6853, N531, N4100);
buf BUF1 (N7370, N7363);
xor XOR2 (N7371, N7367, N4100);
buf BUF1 (N7372, N7371);
not NOT1 (N7373, N7357);
nand NAND3 (N7374, N7361, N2904, N2500);
xor XOR2 (N7375, N7374, N1987);
or OR3 (N7376, N7369, N4912, N2207);
buf BUF1 (N7377, N7376);
nor NOR3 (N7378, N7362, N2146, N1884);
nand NAND3 (N7379, N7370, N6773, N3211);
nor NOR3 (N7380, N7378, N2404, N4793);
buf BUF1 (N7381, N7380);
not NOT1 (N7382, N7373);
not NOT1 (N7383, N7368);
buf BUF1 (N7384, N7383);
buf BUF1 (N7385, N7347);
nor NOR3 (N7386, N7372, N4893, N6643);
buf BUF1 (N7387, N7379);
xor XOR2 (N7388, N7386, N1256);
nand NAND2 (N7389, N7385, N3809);
or OR2 (N7390, N7352, N1586);
buf BUF1 (N7391, N7387);
nand NAND2 (N7392, N7390, N3851);
buf BUF1 (N7393, N7375);
nor NOR3 (N7394, N7358, N1702, N1966);
buf BUF1 (N7395, N7394);
xor XOR2 (N7396, N7382, N4626);
buf BUF1 (N7397, N7393);
and AND3 (N7398, N7381, N2027, N2764);
or OR3 (N7399, N7389, N4384, N6480);
buf BUF1 (N7400, N7388);
buf BUF1 (N7401, N7398);
xor XOR2 (N7402, N7396, N4298);
buf BUF1 (N7403, N7391);
xor XOR2 (N7404, N7400, N4873);
buf BUF1 (N7405, N7377);
and AND2 (N7406, N7401, N307);
nor NOR2 (N7407, N7392, N1780);
nor NOR3 (N7408, N7407, N3715, N4357);
buf BUF1 (N7409, N7397);
buf BUF1 (N7410, N7409);
and AND3 (N7411, N7395, N264, N46);
not NOT1 (N7412, N7384);
buf BUF1 (N7413, N7412);
buf BUF1 (N7414, N7406);
buf BUF1 (N7415, N7405);
and AND4 (N7416, N7403, N4287, N1591, N4837);
or OR2 (N7417, N7411, N4426);
and AND4 (N7418, N7414, N5255, N4888, N5864);
nand NAND3 (N7419, N7404, N7127, N6027);
and AND2 (N7420, N7417, N4857);
not NOT1 (N7421, N7410);
not NOT1 (N7422, N7402);
nor NOR3 (N7423, N7413, N3970, N6812);
nand NAND3 (N7424, N7419, N3557, N6093);
buf BUF1 (N7425, N7415);
buf BUF1 (N7426, N7418);
buf BUF1 (N7427, N7422);
buf BUF1 (N7428, N7423);
xor XOR2 (N7429, N7427, N432);
nor NOR2 (N7430, N7428, N4498);
nand NAND4 (N7431, N7424, N199, N1860, N2891);
not NOT1 (N7432, N7426);
or OR4 (N7433, N7416, N7184, N3655, N4708);
xor XOR2 (N7434, N7421, N3765);
and AND4 (N7435, N7432, N233, N4964, N6389);
xor XOR2 (N7436, N7433, N3653);
xor XOR2 (N7437, N7435, N1064);
and AND4 (N7438, N7408, N162, N1292, N281);
not NOT1 (N7439, N7429);
xor XOR2 (N7440, N7399, N4216);
nand NAND3 (N7441, N7420, N1854, N5341);
xor XOR2 (N7442, N7438, N4670);
nand NAND2 (N7443, N7439, N1692);
and AND2 (N7444, N7440, N4886);
xor XOR2 (N7445, N7431, N1198);
nand NAND4 (N7446, N7445, N1108, N4164, N766);
or OR3 (N7447, N7430, N6042, N2617);
not NOT1 (N7448, N7444);
nand NAND3 (N7449, N7434, N5028, N4387);
not NOT1 (N7450, N7425);
and AND4 (N7451, N7448, N1542, N1653, N2314);
nor NOR4 (N7452, N7449, N4508, N1564, N5371);
buf BUF1 (N7453, N7441);
nand NAND3 (N7454, N7437, N2186, N1859);
xor XOR2 (N7455, N7436, N1656);
nand NAND2 (N7456, N7453, N7159);
not NOT1 (N7457, N7452);
or OR2 (N7458, N7442, N4254);
and AND4 (N7459, N7457, N2138, N733, N6544);
nor NOR4 (N7460, N7458, N6036, N805, N2166);
buf BUF1 (N7461, N7456);
buf BUF1 (N7462, N7459);
nor NOR2 (N7463, N7443, N4339);
nand NAND2 (N7464, N7447, N4121);
or OR4 (N7465, N7454, N6147, N4374, N3392);
nand NAND4 (N7466, N7463, N3207, N3450, N1604);
nor NOR3 (N7467, N7464, N185, N7066);
buf BUF1 (N7468, N7451);
and AND2 (N7469, N7460, N2265);
xor XOR2 (N7470, N7455, N345);
or OR4 (N7471, N7450, N668, N1674, N1213);
nor NOR4 (N7472, N7462, N1518, N6684, N3185);
and AND4 (N7473, N7468, N7045, N6926, N5618);
or OR4 (N7474, N7471, N6284, N5355, N5016);
nand NAND4 (N7475, N7473, N4516, N1737, N6496);
nand NAND3 (N7476, N7465, N7091, N1412);
nor NOR3 (N7477, N7470, N3865, N1292);
buf BUF1 (N7478, N7469);
nor NOR4 (N7479, N7467, N952, N1880, N5093);
and AND3 (N7480, N7475, N6045, N436);
and AND2 (N7481, N7478, N4852);
or OR3 (N7482, N7480, N2746, N6621);
and AND2 (N7483, N7477, N7422);
xor XOR2 (N7484, N7466, N3200);
not NOT1 (N7485, N7472);
not NOT1 (N7486, N7476);
or OR4 (N7487, N7485, N2624, N6693, N748);
nand NAND3 (N7488, N7487, N446, N4100);
buf BUF1 (N7489, N7446);
and AND2 (N7490, N7489, N4385);
buf BUF1 (N7491, N7486);
and AND3 (N7492, N7484, N629, N2989);
or OR3 (N7493, N7492, N2047, N1016);
and AND3 (N7494, N7493, N7373, N5103);
or OR4 (N7495, N7479, N5139, N1102, N4944);
buf BUF1 (N7496, N7494);
nand NAND2 (N7497, N7481, N4503);
and AND4 (N7498, N7497, N1398, N3475, N4101);
nand NAND3 (N7499, N7491, N2650, N1047);
or OR3 (N7500, N7498, N4275, N4077);
xor XOR2 (N7501, N7499, N2016);
buf BUF1 (N7502, N7495);
buf BUF1 (N7503, N7500);
or OR4 (N7504, N7503, N1310, N1797, N5256);
or OR3 (N7505, N7502, N1586, N3782);
buf BUF1 (N7506, N7461);
not NOT1 (N7507, N7490);
xor XOR2 (N7508, N7506, N7063);
nor NOR4 (N7509, N7501, N6664, N6340, N6858);
buf BUF1 (N7510, N7483);
not NOT1 (N7511, N7504);
nand NAND3 (N7512, N7507, N3074, N5009);
not NOT1 (N7513, N7509);
nand NAND4 (N7514, N7511, N4309, N3754, N6071);
or OR3 (N7515, N7496, N3908, N5848);
nor NOR3 (N7516, N7474, N5195, N4308);
xor XOR2 (N7517, N7514, N5803);
or OR4 (N7518, N7482, N7443, N3080, N2895);
or OR2 (N7519, N7513, N7446);
or OR3 (N7520, N7512, N1492, N389);
nand NAND4 (N7521, N7488, N1250, N4706, N2048);
or OR4 (N7522, N7519, N7271, N3704, N6752);
not NOT1 (N7523, N7505);
xor XOR2 (N7524, N7520, N2303);
xor XOR2 (N7525, N7524, N3998);
nor NOR2 (N7526, N7510, N630);
and AND2 (N7527, N7518, N5720);
or OR4 (N7528, N7525, N1765, N4808, N2885);
buf BUF1 (N7529, N7523);
and AND3 (N7530, N7527, N4571, N16);
buf BUF1 (N7531, N7516);
buf BUF1 (N7532, N7529);
nor NOR2 (N7533, N7530, N3929);
or OR2 (N7534, N7521, N22);
not NOT1 (N7535, N7528);
not NOT1 (N7536, N7531);
nor NOR3 (N7537, N7517, N3092, N1745);
buf BUF1 (N7538, N7526);
buf BUF1 (N7539, N7522);
not NOT1 (N7540, N7515);
or OR2 (N7541, N7533, N3832);
nor NOR4 (N7542, N7538, N4285, N2739, N2618);
xor XOR2 (N7543, N7537, N2869);
nor NOR3 (N7544, N7543, N6608, N2387);
or OR4 (N7545, N7536, N457, N1608, N5690);
buf BUF1 (N7546, N7540);
not NOT1 (N7547, N7546);
nor NOR3 (N7548, N7542, N3612, N1843);
not NOT1 (N7549, N7508);
not NOT1 (N7550, N7547);
or OR4 (N7551, N7534, N2338, N4319, N662);
nor NOR3 (N7552, N7535, N7223, N4099);
xor XOR2 (N7553, N7552, N643);
or OR3 (N7554, N7541, N6720, N2766);
nor NOR2 (N7555, N7539, N42);
or OR4 (N7556, N7532, N3080, N1025, N4844);
not NOT1 (N7557, N7554);
xor XOR2 (N7558, N7550, N3717);
nand NAND2 (N7559, N7545, N6821);
nor NOR4 (N7560, N7553, N994, N3280, N4917);
buf BUF1 (N7561, N7559);
not NOT1 (N7562, N7549);
or OR2 (N7563, N7555, N6619);
not NOT1 (N7564, N7556);
or OR3 (N7565, N7564, N3196, N7515);
xor XOR2 (N7566, N7557, N6506);
buf BUF1 (N7567, N7548);
buf BUF1 (N7568, N7562);
nand NAND2 (N7569, N7565, N6605);
not NOT1 (N7570, N7561);
buf BUF1 (N7571, N7570);
nor NOR2 (N7572, N7569, N4051);
nand NAND3 (N7573, N7567, N1501, N4258);
and AND2 (N7574, N7563, N5521);
nor NOR4 (N7575, N7544, N725, N537, N269);
nand NAND4 (N7576, N7573, N866, N3633, N4557);
or OR2 (N7577, N7558, N3143);
nand NAND3 (N7578, N7551, N6370, N6708);
and AND3 (N7579, N7571, N4293, N1092);
buf BUF1 (N7580, N7572);
xor XOR2 (N7581, N7566, N4918);
xor XOR2 (N7582, N7575, N57);
not NOT1 (N7583, N7560);
buf BUF1 (N7584, N7583);
nor NOR2 (N7585, N7568, N6632);
nor NOR4 (N7586, N7584, N5613, N1120, N2023);
nor NOR2 (N7587, N7576, N2870);
xor XOR2 (N7588, N7585, N7497);
nand NAND4 (N7589, N7580, N2468, N4104, N4504);
nor NOR4 (N7590, N7586, N4600, N3056, N3512);
or OR2 (N7591, N7574, N126);
xor XOR2 (N7592, N7591, N858);
buf BUF1 (N7593, N7589);
xor XOR2 (N7594, N7579, N562);
xor XOR2 (N7595, N7578, N818);
nand NAND4 (N7596, N7593, N3519, N3448, N1682);
xor XOR2 (N7597, N7581, N7475);
xor XOR2 (N7598, N7577, N6350);
nand NAND3 (N7599, N7582, N5536, N2732);
buf BUF1 (N7600, N7592);
and AND4 (N7601, N7597, N1949, N5370, N1476);
nand NAND3 (N7602, N7600, N1772, N7109);
or OR4 (N7603, N7588, N5900, N3808, N301);
nor NOR2 (N7604, N7595, N4388);
not NOT1 (N7605, N7598);
or OR2 (N7606, N7596, N4546);
nor NOR3 (N7607, N7587, N1263, N2129);
not NOT1 (N7608, N7599);
nand NAND3 (N7609, N7602, N4689, N2139);
not NOT1 (N7610, N7606);
xor XOR2 (N7611, N7609, N88);
nand NAND2 (N7612, N7601, N6538);
or OR2 (N7613, N7607, N6661);
nor NOR2 (N7614, N7613, N7294);
xor XOR2 (N7615, N7610, N4074);
and AND4 (N7616, N7614, N4329, N454, N3154);
nor NOR2 (N7617, N7616, N2988);
and AND2 (N7618, N7608, N570);
not NOT1 (N7619, N7594);
buf BUF1 (N7620, N7590);
xor XOR2 (N7621, N7617, N1743);
xor XOR2 (N7622, N7603, N4647);
or OR2 (N7623, N7622, N2019);
nor NOR2 (N7624, N7623, N1915);
and AND4 (N7625, N7604, N7373, N3585, N2839);
nand NAND2 (N7626, N7605, N2043);
buf BUF1 (N7627, N7620);
and AND2 (N7628, N7618, N7302);
nor NOR2 (N7629, N7628, N2737);
buf BUF1 (N7630, N7619);
and AND3 (N7631, N7612, N5839, N3461);
xor XOR2 (N7632, N7627, N3135);
xor XOR2 (N7633, N7621, N3061);
or OR4 (N7634, N7611, N1939, N1564, N2589);
not NOT1 (N7635, N7625);
and AND4 (N7636, N7629, N2632, N946, N5789);
or OR2 (N7637, N7626, N4702);
buf BUF1 (N7638, N7633);
not NOT1 (N7639, N7615);
nand NAND2 (N7640, N7637, N540);
nor NOR2 (N7641, N7635, N190);
or OR4 (N7642, N7631, N655, N2438, N3495);
or OR2 (N7643, N7624, N6255);
nand NAND3 (N7644, N7640, N7056, N7011);
nor NOR4 (N7645, N7636, N6219, N1750, N4635);
or OR4 (N7646, N7642, N553, N1303, N4560);
or OR3 (N7647, N7641, N4634, N2931);
and AND4 (N7648, N7632, N6924, N5057, N5561);
not NOT1 (N7649, N7634);
nand NAND4 (N7650, N7639, N4689, N6284, N475);
xor XOR2 (N7651, N7645, N415);
buf BUF1 (N7652, N7646);
buf BUF1 (N7653, N7650);
nor NOR2 (N7654, N7648, N192);
and AND3 (N7655, N7647, N1539, N2943);
not NOT1 (N7656, N7630);
nor NOR3 (N7657, N7649, N3927, N6663);
and AND4 (N7658, N7656, N6194, N781, N5210);
xor XOR2 (N7659, N7653, N2313);
not NOT1 (N7660, N7654);
nand NAND2 (N7661, N7657, N6508);
nand NAND3 (N7662, N7644, N2722, N4176);
and AND3 (N7663, N7643, N4114, N1357);
nor NOR3 (N7664, N7638, N4086, N1644);
nor NOR4 (N7665, N7651, N4531, N5445, N74);
xor XOR2 (N7666, N7664, N4636);
or OR4 (N7667, N7662, N4886, N2035, N7302);
and AND2 (N7668, N7667, N6279);
or OR2 (N7669, N7655, N1193);
nand NAND3 (N7670, N7668, N2859, N2521);
or OR2 (N7671, N7659, N4419);
xor XOR2 (N7672, N7663, N843);
and AND2 (N7673, N7660, N6765);
xor XOR2 (N7674, N7670, N2202);
nor NOR4 (N7675, N7674, N2254, N3000, N5147);
not NOT1 (N7676, N7666);
or OR2 (N7677, N7652, N2420);
nand NAND2 (N7678, N7669, N2307);
buf BUF1 (N7679, N7676);
xor XOR2 (N7680, N7661, N4928);
nor NOR2 (N7681, N7672, N6154);
and AND4 (N7682, N7678, N2904, N5024, N4759);
buf BUF1 (N7683, N7658);
not NOT1 (N7684, N7679);
xor XOR2 (N7685, N7677, N4523);
nand NAND2 (N7686, N7682, N1436);
and AND2 (N7687, N7671, N2129);
buf BUF1 (N7688, N7675);
not NOT1 (N7689, N7673);
not NOT1 (N7690, N7683);
and AND2 (N7691, N7688, N7284);
not NOT1 (N7692, N7685);
buf BUF1 (N7693, N7665);
or OR2 (N7694, N7686, N4276);
nand NAND3 (N7695, N7692, N5379, N679);
nor NOR4 (N7696, N7693, N6266, N5439, N1149);
or OR4 (N7697, N7694, N1170, N5664, N4802);
nor NOR3 (N7698, N7681, N1264, N4958);
nor NOR4 (N7699, N7698, N1935, N309, N2748);
xor XOR2 (N7700, N7684, N2785);
not NOT1 (N7701, N7696);
xor XOR2 (N7702, N7697, N6969);
not NOT1 (N7703, N7687);
buf BUF1 (N7704, N7701);
and AND2 (N7705, N7704, N3438);
and AND2 (N7706, N7700, N1120);
or OR2 (N7707, N7680, N4425);
xor XOR2 (N7708, N7695, N3121);
nand NAND4 (N7709, N7690, N3669, N7515, N172);
or OR3 (N7710, N7691, N6987, N2155);
nand NAND3 (N7711, N7706, N276, N2300);
and AND3 (N7712, N7689, N7271, N2317);
nor NOR3 (N7713, N7699, N1215, N3705);
and AND2 (N7714, N7705, N7603);
or OR2 (N7715, N7710, N6836);
nor NOR3 (N7716, N7708, N3133, N4516);
not NOT1 (N7717, N7713);
or OR2 (N7718, N7709, N1470);
nor NOR4 (N7719, N7714, N7604, N243, N3131);
not NOT1 (N7720, N7719);
and AND3 (N7721, N7715, N5396, N5794);
nand NAND4 (N7722, N7716, N3991, N909, N59);
nor NOR2 (N7723, N7712, N5669);
xor XOR2 (N7724, N7707, N2299);
nand NAND2 (N7725, N7724, N6165);
not NOT1 (N7726, N7718);
xor XOR2 (N7727, N7711, N2369);
xor XOR2 (N7728, N7727, N6337);
or OR4 (N7729, N7720, N2308, N1991, N7562);
or OR3 (N7730, N7703, N7265, N3874);
xor XOR2 (N7731, N7728, N5793);
xor XOR2 (N7732, N7721, N5479);
buf BUF1 (N7733, N7726);
nor NOR2 (N7734, N7717, N1879);
nand NAND2 (N7735, N7734, N398);
not NOT1 (N7736, N7733);
buf BUF1 (N7737, N7702);
nand NAND2 (N7738, N7735, N7044);
xor XOR2 (N7739, N7738, N46);
and AND4 (N7740, N7730, N3151, N6796, N5935);
buf BUF1 (N7741, N7732);
and AND3 (N7742, N7725, N1598, N2238);
buf BUF1 (N7743, N7740);
not NOT1 (N7744, N7736);
nor NOR3 (N7745, N7722, N1101, N2545);
or OR4 (N7746, N7745, N1534, N2797, N5812);
and AND3 (N7747, N7731, N3860, N5427);
not NOT1 (N7748, N7747);
nand NAND4 (N7749, N7737, N6568, N4003, N7143);
nor NOR2 (N7750, N7744, N4483);
buf BUF1 (N7751, N7729);
nor NOR2 (N7752, N7742, N6088);
buf BUF1 (N7753, N7739);
buf BUF1 (N7754, N7749);
or OR3 (N7755, N7741, N3351, N3205);
not NOT1 (N7756, N7754);
and AND2 (N7757, N7746, N2687);
not NOT1 (N7758, N7751);
buf BUF1 (N7759, N7748);
nand NAND2 (N7760, N7753, N5595);
buf BUF1 (N7761, N7757);
or OR2 (N7762, N7723, N1787);
buf BUF1 (N7763, N7750);
xor XOR2 (N7764, N7763, N1882);
nor NOR2 (N7765, N7758, N4211);
and AND3 (N7766, N7743, N1379, N7214);
buf BUF1 (N7767, N7764);
and AND4 (N7768, N7762, N3902, N6497, N1812);
or OR4 (N7769, N7760, N7597, N411, N3379);
nor NOR2 (N7770, N7755, N2412);
or OR4 (N7771, N7752, N3391, N291, N5851);
nor NOR3 (N7772, N7759, N134, N1101);
nand NAND2 (N7773, N7770, N2030);
buf BUF1 (N7774, N7773);
and AND4 (N7775, N7766, N5406, N5603, N6853);
and AND4 (N7776, N7765, N2915, N5622, N5866);
nand NAND2 (N7777, N7768, N1175);
nand NAND2 (N7778, N7777, N3855);
buf BUF1 (N7779, N7771);
or OR3 (N7780, N7776, N6644, N7652);
nand NAND4 (N7781, N7769, N706, N6297, N905);
or OR3 (N7782, N7779, N4201, N821);
nor NOR2 (N7783, N7780, N6288);
nor NOR2 (N7784, N7782, N1223);
nand NAND4 (N7785, N7772, N6222, N2503, N341);
xor XOR2 (N7786, N7767, N7653);
or OR3 (N7787, N7786, N7283, N2020);
xor XOR2 (N7788, N7785, N6122);
and AND2 (N7789, N7787, N7594);
or OR2 (N7790, N7784, N7503);
not NOT1 (N7791, N7790);
and AND4 (N7792, N7778, N5642, N7779, N2193);
nor NOR2 (N7793, N7774, N2874);
or OR4 (N7794, N7761, N6791, N502, N3684);
nor NOR3 (N7795, N7789, N6038, N6988);
nand NAND2 (N7796, N7783, N2842);
or OR4 (N7797, N7792, N6996, N2539, N2158);
or OR4 (N7798, N7797, N3974, N7593, N3716);
buf BUF1 (N7799, N7796);
or OR4 (N7800, N7788, N3293, N4214, N6183);
xor XOR2 (N7801, N7799, N3907);
not NOT1 (N7802, N7781);
nand NAND2 (N7803, N7794, N1978);
or OR2 (N7804, N7756, N5020);
nand NAND4 (N7805, N7791, N7380, N5576, N4568);
nor NOR4 (N7806, N7775, N432, N651, N2854);
xor XOR2 (N7807, N7802, N6574);
nor NOR4 (N7808, N7804, N7254, N6102, N4446);
buf BUF1 (N7809, N7800);
and AND2 (N7810, N7807, N1293);
and AND4 (N7811, N7809, N2287, N2960, N3593);
not NOT1 (N7812, N7801);
not NOT1 (N7813, N7798);
xor XOR2 (N7814, N7793, N1753);
nor NOR2 (N7815, N7806, N2487);
or OR2 (N7816, N7812, N3594);
xor XOR2 (N7817, N7811, N7070);
buf BUF1 (N7818, N7815);
or OR3 (N7819, N7817, N930, N1472);
buf BUF1 (N7820, N7810);
nor NOR3 (N7821, N7820, N1911, N2266);
not NOT1 (N7822, N7808);
not NOT1 (N7823, N7822);
and AND3 (N7824, N7795, N809, N5990);
or OR2 (N7825, N7814, N6976);
xor XOR2 (N7826, N7816, N6246);
nor NOR2 (N7827, N7826, N4502);
nor NOR2 (N7828, N7824, N3687);
or OR3 (N7829, N7805, N5106, N7597);
xor XOR2 (N7830, N7827, N3054);
nand NAND4 (N7831, N7830, N2959, N1230, N6828);
not NOT1 (N7832, N7818);
xor XOR2 (N7833, N7825, N4817);
nor NOR3 (N7834, N7831, N5967, N3898);
buf BUF1 (N7835, N7833);
or OR3 (N7836, N7821, N6748, N6023);
or OR3 (N7837, N7813, N7021, N5279);
or OR3 (N7838, N7832, N5374, N5087);
xor XOR2 (N7839, N7828, N2231);
buf BUF1 (N7840, N7829);
nor NOR3 (N7841, N7803, N2641, N1740);
and AND3 (N7842, N7837, N4684, N2765);
nand NAND4 (N7843, N7841, N5283, N329, N4163);
xor XOR2 (N7844, N7843, N29);
nor NOR4 (N7845, N7835, N1376, N1646, N1955);
nand NAND3 (N7846, N7823, N3212, N2870);
xor XOR2 (N7847, N7845, N2424);
nor NOR4 (N7848, N7838, N4567, N4390, N4996);
xor XOR2 (N7849, N7839, N2868);
and AND3 (N7850, N7836, N127, N4275);
xor XOR2 (N7851, N7842, N704);
nor NOR3 (N7852, N7851, N1836, N4465);
or OR2 (N7853, N7849, N4196);
buf BUF1 (N7854, N7853);
nand NAND3 (N7855, N7819, N724, N7389);
nand NAND2 (N7856, N7848, N1271);
buf BUF1 (N7857, N7854);
buf BUF1 (N7858, N7855);
nor NOR4 (N7859, N7857, N2553, N3294, N3558);
and AND4 (N7860, N7844, N3958, N396, N7619);
and AND2 (N7861, N7858, N4678);
and AND4 (N7862, N7852, N2341, N7335, N4761);
buf BUF1 (N7863, N7861);
not NOT1 (N7864, N7850);
nand NAND2 (N7865, N7834, N2297);
nor NOR2 (N7866, N7860, N1139);
buf BUF1 (N7867, N7862);
not NOT1 (N7868, N7840);
not NOT1 (N7869, N7847);
and AND4 (N7870, N7866, N7834, N5466, N5997);
not NOT1 (N7871, N7846);
xor XOR2 (N7872, N7863, N4686);
buf BUF1 (N7873, N7864);
or OR4 (N7874, N7868, N5982, N1472, N6924);
and AND2 (N7875, N7859, N2820);
buf BUF1 (N7876, N7871);
nor NOR4 (N7877, N7876, N5751, N6856, N5596);
and AND2 (N7878, N7877, N7254);
nand NAND3 (N7879, N7873, N3061, N717);
nand NAND2 (N7880, N7865, N7625);
or OR4 (N7881, N7872, N6986, N1554, N2141);
and AND3 (N7882, N7878, N6952, N7392);
nor NOR4 (N7883, N7870, N4073, N2022, N6105);
nand NAND3 (N7884, N7875, N618, N3757);
xor XOR2 (N7885, N7874, N6857);
or OR4 (N7886, N7856, N6633, N4285, N3077);
nand NAND3 (N7887, N7884, N4505, N1073);
nand NAND3 (N7888, N7882, N1261, N6006);
not NOT1 (N7889, N7888);
xor XOR2 (N7890, N7879, N3185);
or OR4 (N7891, N7887, N1692, N1839, N3896);
nand NAND4 (N7892, N7889, N836, N4672, N1705);
and AND3 (N7893, N7869, N7271, N7834);
buf BUF1 (N7894, N7891);
buf BUF1 (N7895, N7885);
not NOT1 (N7896, N7894);
xor XOR2 (N7897, N7886, N228);
and AND4 (N7898, N7881, N4108, N6932, N354);
nand NAND3 (N7899, N7883, N2937, N1653);
and AND4 (N7900, N7890, N7722, N664, N2987);
nor NOR4 (N7901, N7898, N5508, N7398, N5907);
buf BUF1 (N7902, N7880);
not NOT1 (N7903, N7893);
and AND4 (N7904, N7903, N5849, N5403, N3357);
buf BUF1 (N7905, N7892);
or OR2 (N7906, N7904, N1712);
xor XOR2 (N7907, N7905, N1401);
nor NOR2 (N7908, N7901, N404);
not NOT1 (N7909, N7867);
and AND3 (N7910, N7906, N368, N5733);
and AND3 (N7911, N7909, N2005, N7257);
or OR4 (N7912, N7908, N5262, N7582, N1725);
buf BUF1 (N7913, N7897);
and AND2 (N7914, N7907, N6586);
buf BUF1 (N7915, N7900);
buf BUF1 (N7916, N7895);
and AND3 (N7917, N7911, N2206, N7548);
xor XOR2 (N7918, N7916, N2107);
buf BUF1 (N7919, N7910);
or OR4 (N7920, N7912, N6736, N7792, N4176);
buf BUF1 (N7921, N7914);
nand NAND4 (N7922, N7919, N6224, N4556, N4642);
buf BUF1 (N7923, N7918);
nand NAND4 (N7924, N7920, N2815, N146, N7118);
buf BUF1 (N7925, N7899);
or OR4 (N7926, N7915, N7410, N2731, N5937);
buf BUF1 (N7927, N7917);
nand NAND3 (N7928, N7927, N7389, N1539);
nand NAND4 (N7929, N7925, N1713, N1417, N5855);
xor XOR2 (N7930, N7923, N3138);
or OR2 (N7931, N7922, N2053);
or OR4 (N7932, N7896, N429, N1058, N7287);
nand NAND3 (N7933, N7924, N3041, N4624);
and AND2 (N7934, N7932, N5370);
xor XOR2 (N7935, N7926, N872);
not NOT1 (N7936, N7935);
nor NOR2 (N7937, N7930, N3247);
not NOT1 (N7938, N7928);
or OR4 (N7939, N7902, N3218, N2711, N1440);
nand NAND4 (N7940, N7929, N2698, N1166, N4865);
not NOT1 (N7941, N7934);
not NOT1 (N7942, N7933);
and AND2 (N7943, N7941, N4022);
nor NOR2 (N7944, N7939, N4079);
xor XOR2 (N7945, N7944, N6122);
nor NOR3 (N7946, N7913, N2602, N923);
nand NAND4 (N7947, N7940, N926, N4572, N5143);
or OR2 (N7948, N7945, N3938);
or OR3 (N7949, N7948, N5331, N5956);
buf BUF1 (N7950, N7949);
nand NAND3 (N7951, N7946, N4768, N456);
not NOT1 (N7952, N7936);
nand NAND2 (N7953, N7942, N6545);
xor XOR2 (N7954, N7950, N3035);
nand NAND3 (N7955, N7951, N2692, N6008);
buf BUF1 (N7956, N7937);
buf BUF1 (N7957, N7954);
nand NAND2 (N7958, N7931, N6839);
nand NAND2 (N7959, N7958, N2762);
and AND2 (N7960, N7943, N5709);
and AND2 (N7961, N7938, N2875);
or OR2 (N7962, N7955, N2659);
nor NOR3 (N7963, N7953, N2988, N5491);
buf BUF1 (N7964, N7963);
nor NOR4 (N7965, N7960, N4402, N6166, N6175);
not NOT1 (N7966, N7964);
and AND3 (N7967, N7921, N3015, N1368);
nand NAND2 (N7968, N7961, N461);
or OR3 (N7969, N7952, N4931, N5037);
and AND2 (N7970, N7962, N731);
not NOT1 (N7971, N7959);
or OR3 (N7972, N7956, N2387, N1474);
nand NAND4 (N7973, N7966, N3064, N3803, N5312);
and AND2 (N7974, N7947, N2986);
and AND2 (N7975, N7970, N3238);
nor NOR4 (N7976, N7967, N2958, N926, N5631);
not NOT1 (N7977, N7974);
xor XOR2 (N7978, N7968, N6435);
or OR2 (N7979, N7975, N7688);
nor NOR3 (N7980, N7965, N912, N404);
not NOT1 (N7981, N7977);
xor XOR2 (N7982, N7978, N1625);
or OR2 (N7983, N7981, N4697);
not NOT1 (N7984, N7983);
nand NAND2 (N7985, N7979, N3398);
buf BUF1 (N7986, N7976);
or OR2 (N7987, N7985, N1376);
nand NAND3 (N7988, N7987, N1651, N1507);
xor XOR2 (N7989, N7982, N6362);
xor XOR2 (N7990, N7972, N7840);
nor NOR2 (N7991, N7990, N6940);
nor NOR2 (N7992, N7957, N3521);
and AND4 (N7993, N7971, N3841, N6124, N3348);
nand NAND4 (N7994, N7980, N981, N1821, N2572);
not NOT1 (N7995, N7994);
not NOT1 (N7996, N7988);
nand NAND4 (N7997, N7996, N7473, N246, N2990);
not NOT1 (N7998, N7984);
nand NAND4 (N7999, N7969, N3496, N6700, N4376);
xor XOR2 (N8000, N7993, N7645);
not NOT1 (N8001, N8000);
and AND4 (N8002, N8001, N7044, N273, N2634);
and AND4 (N8003, N7998, N7881, N971, N4338);
nand NAND2 (N8004, N7991, N7989);
nor NOR4 (N8005, N4670, N690, N3539, N1045);
buf BUF1 (N8006, N8004);
xor XOR2 (N8007, N7995, N4212);
nand NAND2 (N8008, N7992, N839);
buf BUF1 (N8009, N7997);
not NOT1 (N8010, N8006);
nand NAND4 (N8011, N8010, N6008, N4589, N149);
nor NOR3 (N8012, N8005, N5315, N5835);
or OR3 (N8013, N7986, N4352, N4313);
xor XOR2 (N8014, N8012, N3678);
or OR4 (N8015, N8003, N5319, N4556, N4296);
and AND4 (N8016, N8009, N1547, N3506, N176);
nor NOR3 (N8017, N8011, N1211, N1162);
xor XOR2 (N8018, N7973, N7703);
nor NOR3 (N8019, N8002, N3599, N6234);
or OR2 (N8020, N8019, N4781);
xor XOR2 (N8021, N8017, N8020);
xor XOR2 (N8022, N3385, N3297);
not NOT1 (N8023, N8016);
or OR3 (N8024, N8023, N3792, N7646);
or OR2 (N8025, N8024, N3308);
nand NAND3 (N8026, N7999, N2873, N2104);
buf BUF1 (N8027, N8007);
xor XOR2 (N8028, N8025, N5396);
and AND2 (N8029, N8015, N5696);
nand NAND3 (N8030, N8029, N7624, N5278);
or OR4 (N8031, N8028, N7707, N243, N5651);
or OR2 (N8032, N8026, N3732);
buf BUF1 (N8033, N8008);
nand NAND2 (N8034, N8018, N6570);
and AND3 (N8035, N8033, N4458, N914);
or OR3 (N8036, N8021, N6523, N7595);
or OR4 (N8037, N8034, N1227, N1052, N5152);
xor XOR2 (N8038, N8030, N2377);
or OR3 (N8039, N8022, N5292, N3447);
nand NAND3 (N8040, N8035, N6729, N4135);
nor NOR2 (N8041, N8032, N6469);
not NOT1 (N8042, N8038);
buf BUF1 (N8043, N8042);
buf BUF1 (N8044, N8027);
nand NAND2 (N8045, N8014, N2315);
nand NAND3 (N8046, N8031, N816, N4984);
nand NAND3 (N8047, N8044, N3289, N6363);
or OR3 (N8048, N8036, N848, N6755);
or OR4 (N8049, N8048, N6564, N4966, N185);
nor NOR2 (N8050, N8049, N3421);
not NOT1 (N8051, N8045);
and AND4 (N8052, N8013, N6195, N5219, N3275);
or OR4 (N8053, N8039, N7466, N4527, N4737);
and AND3 (N8054, N8043, N850, N1629);
xor XOR2 (N8055, N8041, N5898);
nand NAND3 (N8056, N8047, N5920, N1785);
nor NOR4 (N8057, N8052, N5210, N4401, N2025);
and AND3 (N8058, N8040, N4969, N2614);
and AND4 (N8059, N8055, N7803, N3131, N1583);
nand NAND2 (N8060, N8037, N1806);
buf BUF1 (N8061, N8050);
and AND2 (N8062, N8056, N6563);
and AND2 (N8063, N8061, N1975);
xor XOR2 (N8064, N8054, N4172);
nand NAND2 (N8065, N8059, N6214);
nand NAND3 (N8066, N8046, N6055, N6696);
buf BUF1 (N8067, N8065);
not NOT1 (N8068, N8064);
nand NAND3 (N8069, N8057, N809, N6115);
nor NOR2 (N8070, N8069, N1727);
nor NOR3 (N8071, N8062, N3658, N5267);
and AND3 (N8072, N8067, N5403, N3926);
nor NOR2 (N8073, N8068, N4469);
or OR2 (N8074, N8072, N1504);
or OR3 (N8075, N8074, N4163, N6698);
buf BUF1 (N8076, N8073);
nor NOR3 (N8077, N8075, N5215, N3492);
nor NOR3 (N8078, N8053, N3663, N920);
nand NAND2 (N8079, N8071, N7200);
nor NOR2 (N8080, N8066, N1833);
buf BUF1 (N8081, N8051);
xor XOR2 (N8082, N8078, N1431);
or OR2 (N8083, N8058, N3664);
or OR4 (N8084, N8063, N7377, N6448, N5486);
nor NOR2 (N8085, N8079, N6593);
nand NAND4 (N8086, N8082, N5833, N5212, N3911);
and AND3 (N8087, N8083, N3132, N6738);
buf BUF1 (N8088, N8076);
nand NAND3 (N8089, N8085, N3304, N4005);
buf BUF1 (N8090, N8060);
xor XOR2 (N8091, N8089, N4176);
not NOT1 (N8092, N8087);
xor XOR2 (N8093, N8081, N2539);
not NOT1 (N8094, N8077);
or OR2 (N8095, N8088, N3021);
xor XOR2 (N8096, N8090, N105);
xor XOR2 (N8097, N8080, N5109);
not NOT1 (N8098, N8070);
and AND2 (N8099, N8094, N8014);
nand NAND4 (N8100, N8084, N6186, N3787, N3389);
nor NOR4 (N8101, N8086, N731, N7732, N66);
and AND2 (N8102, N8098, N340);
not NOT1 (N8103, N8091);
or OR3 (N8104, N8092, N4125, N4928);
xor XOR2 (N8105, N8102, N2606);
buf BUF1 (N8106, N8104);
and AND3 (N8107, N8096, N4645, N1686);
and AND4 (N8108, N8107, N3367, N6112, N5622);
xor XOR2 (N8109, N8093, N868);
nor NOR2 (N8110, N8097, N1855);
buf BUF1 (N8111, N8108);
nor NOR3 (N8112, N8099, N532, N142);
xor XOR2 (N8113, N8110, N5416);
and AND4 (N8114, N8111, N8097, N4204, N325);
and AND3 (N8115, N8101, N7259, N854);
not NOT1 (N8116, N8113);
xor XOR2 (N8117, N8095, N3294);
buf BUF1 (N8118, N8116);
xor XOR2 (N8119, N8114, N7927);
buf BUF1 (N8120, N8115);
not NOT1 (N8121, N8117);
nand NAND4 (N8122, N8118, N6739, N1346, N6676);
buf BUF1 (N8123, N8105);
not NOT1 (N8124, N8119);
not NOT1 (N8125, N8103);
or OR2 (N8126, N8121, N941);
nand NAND3 (N8127, N8109, N3904, N812);
and AND2 (N8128, N8100, N5640);
nand NAND4 (N8129, N8127, N654, N4001, N7809);
or OR4 (N8130, N8123, N555, N1427, N1792);
nor NOR4 (N8131, N8122, N8043, N3567, N4030);
nor NOR3 (N8132, N8130, N609, N2565);
and AND3 (N8133, N8106, N8015, N7949);
buf BUF1 (N8134, N8112);
xor XOR2 (N8135, N8125, N6713);
and AND4 (N8136, N8135, N3017, N3263, N7398);
not NOT1 (N8137, N8126);
not NOT1 (N8138, N8129);
not NOT1 (N8139, N8132);
not NOT1 (N8140, N8124);
not NOT1 (N8141, N8140);
xor XOR2 (N8142, N8133, N4992);
and AND3 (N8143, N8138, N4538, N2300);
buf BUF1 (N8144, N8143);
nor NOR2 (N8145, N8120, N2641);
xor XOR2 (N8146, N8142, N278);
and AND2 (N8147, N8128, N3634);
and AND3 (N8148, N8136, N6262, N4649);
nor NOR4 (N8149, N8137, N7249, N4865, N7448);
and AND2 (N8150, N8149, N2360);
buf BUF1 (N8151, N8144);
and AND4 (N8152, N8147, N4014, N6078, N2156);
xor XOR2 (N8153, N8141, N2515);
or OR4 (N8154, N8145, N4698, N1749, N5293);
nand NAND4 (N8155, N8134, N6584, N1712, N7613);
not NOT1 (N8156, N8150);
nor NOR3 (N8157, N8148, N1727, N3810);
buf BUF1 (N8158, N8146);
not NOT1 (N8159, N8155);
xor XOR2 (N8160, N8139, N8065);
and AND2 (N8161, N8160, N4825);
and AND3 (N8162, N8157, N2404, N3573);
nand NAND2 (N8163, N8152, N7454);
xor XOR2 (N8164, N8151, N2534);
nor NOR4 (N8165, N8164, N4815, N4677, N6206);
or OR3 (N8166, N8156, N5502, N696);
buf BUF1 (N8167, N8159);
buf BUF1 (N8168, N8158);
nor NOR4 (N8169, N8161, N2237, N412, N6110);
or OR4 (N8170, N8169, N7915, N7158, N1551);
and AND3 (N8171, N8153, N6819, N3198);
or OR2 (N8172, N8163, N1076);
and AND4 (N8173, N8162, N4210, N137, N3589);
nor NOR4 (N8174, N8154, N3752, N4619, N5904);
not NOT1 (N8175, N8173);
and AND4 (N8176, N8168, N2154, N3140, N3240);
and AND3 (N8177, N8175, N3658, N7353);
buf BUF1 (N8178, N8131);
not NOT1 (N8179, N8165);
and AND3 (N8180, N8177, N3282, N6402);
and AND2 (N8181, N8179, N7793);
buf BUF1 (N8182, N8178);
xor XOR2 (N8183, N8174, N7513);
not NOT1 (N8184, N8180);
nor NOR3 (N8185, N8181, N5661, N360);
or OR3 (N8186, N8170, N6011, N1650);
not NOT1 (N8187, N8176);
and AND4 (N8188, N8184, N2926, N3306, N6691);
nand NAND2 (N8189, N8187, N4325);
nand NAND2 (N8190, N8166, N214);
not NOT1 (N8191, N8185);
xor XOR2 (N8192, N8182, N8030);
nand NAND3 (N8193, N8192, N2151, N3109);
and AND4 (N8194, N8190, N1298, N1765, N6139);
nand NAND2 (N8195, N8172, N4369);
nor NOR3 (N8196, N8189, N5996, N2277);
nor NOR3 (N8197, N8186, N5779, N6679);
or OR2 (N8198, N8188, N7484);
or OR3 (N8199, N8197, N5827, N205);
nand NAND2 (N8200, N8191, N5103);
or OR2 (N8201, N8167, N592);
nand NAND4 (N8202, N8183, N1142, N6834, N5279);
xor XOR2 (N8203, N8201, N7934);
nor NOR2 (N8204, N8193, N5531);
nand NAND3 (N8205, N8196, N7077, N6792);
xor XOR2 (N8206, N8205, N1802);
nand NAND3 (N8207, N8200, N5094, N1964);
not NOT1 (N8208, N8207);
or OR3 (N8209, N8202, N1512, N3122);
and AND3 (N8210, N8203, N1261, N5974);
nor NOR2 (N8211, N8194, N6226);
nor NOR2 (N8212, N8199, N6196);
nor NOR4 (N8213, N8206, N2235, N2033, N6113);
nand NAND3 (N8214, N8210, N4255, N6802);
nand NAND2 (N8215, N8213, N3604);
not NOT1 (N8216, N8195);
nand NAND3 (N8217, N8216, N5847, N1719);
and AND4 (N8218, N8211, N4851, N6471, N7682);
nand NAND3 (N8219, N8171, N4302, N7569);
xor XOR2 (N8220, N8219, N330);
nor NOR2 (N8221, N8204, N299);
nor NOR3 (N8222, N8214, N1112, N2352);
nor NOR2 (N8223, N8208, N7203);
nand NAND2 (N8224, N8215, N118);
and AND2 (N8225, N8198, N5083);
xor XOR2 (N8226, N8222, N1098);
buf BUF1 (N8227, N8209);
buf BUF1 (N8228, N8227);
buf BUF1 (N8229, N8212);
nand NAND4 (N8230, N8228, N8111, N4174, N4847);
or OR4 (N8231, N8224, N1702, N1989, N4455);
or OR4 (N8232, N8231, N5177, N6569, N7781);
buf BUF1 (N8233, N8225);
xor XOR2 (N8234, N8226, N3931);
xor XOR2 (N8235, N8223, N7871);
and AND2 (N8236, N8232, N6155);
and AND2 (N8237, N8236, N8122);
nor NOR3 (N8238, N8221, N6276, N1072);
nor NOR3 (N8239, N8218, N1448, N5474);
not NOT1 (N8240, N8237);
nand NAND4 (N8241, N8239, N7775, N2400, N5473);
nand NAND3 (N8242, N8241, N5194, N1520);
buf BUF1 (N8243, N8242);
nor NOR3 (N8244, N8217, N2898, N1661);
nand NAND2 (N8245, N8238, N101);
and AND3 (N8246, N8220, N3872, N5179);
nor NOR3 (N8247, N8235, N3052, N6144);
and AND2 (N8248, N8233, N4132);
nand NAND2 (N8249, N8240, N715);
nand NAND2 (N8250, N8245, N4596);
xor XOR2 (N8251, N8246, N2183);
and AND3 (N8252, N8230, N5940, N3754);
or OR3 (N8253, N8252, N7959, N713);
not NOT1 (N8254, N8253);
nor NOR2 (N8255, N8248, N3952);
and AND2 (N8256, N8244, N5912);
buf BUF1 (N8257, N8254);
or OR3 (N8258, N8251, N5974, N6572);
and AND4 (N8259, N8234, N8216, N6429, N961);
nor NOR2 (N8260, N8229, N4356);
not NOT1 (N8261, N8257);
nand NAND2 (N8262, N8250, N3461);
and AND4 (N8263, N8249, N4030, N1568, N6935);
or OR2 (N8264, N8256, N1617);
xor XOR2 (N8265, N8247, N1469);
nor NOR4 (N8266, N8258, N7573, N7630, N5299);
not NOT1 (N8267, N8265);
nand NAND3 (N8268, N8264, N4111, N162);
not NOT1 (N8269, N8263);
and AND2 (N8270, N8268, N6514);
nor NOR2 (N8271, N8269, N7651);
or OR3 (N8272, N8255, N4612, N4997);
or OR2 (N8273, N8260, N4833);
not NOT1 (N8274, N8270);
nor NOR4 (N8275, N8273, N7188, N3892, N4583);
buf BUF1 (N8276, N8275);
buf BUF1 (N8277, N8243);
and AND4 (N8278, N8266, N1432, N5972, N7441);
nor NOR4 (N8279, N8261, N3195, N736, N1761);
not NOT1 (N8280, N8274);
nor NOR2 (N8281, N8267, N6834);
and AND3 (N8282, N8272, N8260, N724);
and AND3 (N8283, N8262, N3009, N5176);
buf BUF1 (N8284, N8280);
buf BUF1 (N8285, N8278);
nand NAND4 (N8286, N8284, N7575, N5883, N3207);
and AND2 (N8287, N8277, N5089);
or OR4 (N8288, N8287, N6516, N4861, N5076);
buf BUF1 (N8289, N8271);
nand NAND4 (N8290, N8289, N7771, N40, N5836);
xor XOR2 (N8291, N8282, N538);
buf BUF1 (N8292, N8276);
nand NAND3 (N8293, N8279, N4397, N2236);
buf BUF1 (N8294, N8285);
nand NAND2 (N8295, N8283, N3102);
not NOT1 (N8296, N8288);
and AND2 (N8297, N8295, N6883);
nor NOR4 (N8298, N8293, N3198, N7344, N1355);
nor NOR4 (N8299, N8298, N292, N6956, N239);
xor XOR2 (N8300, N8290, N6417);
not NOT1 (N8301, N8300);
buf BUF1 (N8302, N8281);
nand NAND4 (N8303, N8294, N3354, N2595, N2075);
nor NOR4 (N8304, N8296, N6542, N3778, N834);
and AND4 (N8305, N8297, N3086, N5206, N5456);
nor NOR3 (N8306, N8301, N3209, N3464);
buf BUF1 (N8307, N8305);
and AND2 (N8308, N8307, N1093);
nand NAND2 (N8309, N8306, N5362);
not NOT1 (N8310, N8308);
buf BUF1 (N8311, N8302);
nor NOR3 (N8312, N8310, N5050, N6917);
nor NOR3 (N8313, N8259, N1237, N7475);
nor NOR4 (N8314, N8286, N5117, N4313, N2690);
and AND3 (N8315, N8291, N3047, N6316);
nand NAND2 (N8316, N8311, N2046);
buf BUF1 (N8317, N8315);
buf BUF1 (N8318, N8314);
not NOT1 (N8319, N8304);
nor NOR2 (N8320, N8303, N248);
nor NOR2 (N8321, N8318, N4139);
nand NAND2 (N8322, N8317, N1534);
or OR4 (N8323, N8312, N218, N5127, N2621);
and AND3 (N8324, N8321, N6696, N4703);
nand NAND4 (N8325, N8319, N5260, N5000, N2417);
and AND3 (N8326, N8316, N4761, N2402);
nand NAND4 (N8327, N8313, N7932, N3212, N5084);
or OR2 (N8328, N8320, N2738);
buf BUF1 (N8329, N8324);
nor NOR2 (N8330, N8299, N3758);
nand NAND4 (N8331, N8322, N3422, N4239, N5917);
buf BUF1 (N8332, N8309);
not NOT1 (N8333, N8331);
nor NOR4 (N8334, N8333, N2037, N4822, N3287);
and AND4 (N8335, N8332, N2170, N887, N5184);
and AND2 (N8336, N8292, N2383);
buf BUF1 (N8337, N8327);
nand NAND3 (N8338, N8336, N1261, N2697);
nor NOR4 (N8339, N8326, N403, N440, N5246);
xor XOR2 (N8340, N8328, N1573);
not NOT1 (N8341, N8330);
buf BUF1 (N8342, N8339);
and AND2 (N8343, N8337, N5966);
not NOT1 (N8344, N8335);
nor NOR4 (N8345, N8342, N8273, N8154, N1427);
and AND2 (N8346, N8334, N543);
nand NAND3 (N8347, N8344, N4353, N5854);
or OR3 (N8348, N8341, N3293, N3616);
nor NOR4 (N8349, N8340, N5880, N684, N3612);
buf BUF1 (N8350, N8343);
and AND3 (N8351, N8345, N6602, N5898);
not NOT1 (N8352, N8348);
nor NOR2 (N8353, N8346, N583);
nand NAND2 (N8354, N8347, N3882);
nor NOR2 (N8355, N8351, N5708);
xor XOR2 (N8356, N8355, N4383);
xor XOR2 (N8357, N8352, N4149);
or OR2 (N8358, N8329, N1168);
or OR4 (N8359, N8349, N2683, N7558, N7576);
not NOT1 (N8360, N8354);
nand NAND4 (N8361, N8338, N666, N273, N464);
and AND4 (N8362, N8360, N3824, N7712, N2465);
or OR2 (N8363, N8358, N1104);
or OR3 (N8364, N8359, N5984, N2437);
and AND4 (N8365, N8364, N2887, N4465, N7860);
buf BUF1 (N8366, N8356);
xor XOR2 (N8367, N8357, N5629);
and AND2 (N8368, N8361, N1663);
and AND4 (N8369, N8323, N3437, N779, N4814);
buf BUF1 (N8370, N8369);
or OR4 (N8371, N8362, N2194, N9, N4323);
nor NOR2 (N8372, N8371, N4266);
and AND3 (N8373, N8363, N3629, N3637);
nor NOR4 (N8374, N8325, N1822, N3940, N7401);
or OR2 (N8375, N8368, N2299);
xor XOR2 (N8376, N8373, N7404);
or OR2 (N8377, N8350, N7790);
or OR4 (N8378, N8365, N2924, N2460, N5457);
nor NOR3 (N8379, N8367, N5365, N6517);
xor XOR2 (N8380, N8378, N3420);
nand NAND4 (N8381, N8375, N3804, N5713, N7794);
and AND2 (N8382, N8366, N1509);
nor NOR4 (N8383, N8353, N2033, N7820, N6288);
not NOT1 (N8384, N8381);
nor NOR4 (N8385, N8382, N661, N1982, N2339);
or OR2 (N8386, N8383, N2144);
and AND4 (N8387, N8374, N5712, N5577, N2391);
or OR4 (N8388, N8372, N6324, N1971, N3178);
buf BUF1 (N8389, N8387);
not NOT1 (N8390, N8370);
nor NOR3 (N8391, N8388, N5336, N8010);
buf BUF1 (N8392, N8379);
nor NOR2 (N8393, N8392, N1754);
and AND2 (N8394, N8384, N70);
and AND3 (N8395, N8376, N1212, N7895);
buf BUF1 (N8396, N8395);
not NOT1 (N8397, N8396);
not NOT1 (N8398, N8393);
or OR3 (N8399, N8386, N6554, N6780);
nor NOR3 (N8400, N8399, N5891, N7524);
or OR2 (N8401, N8380, N8248);
not NOT1 (N8402, N8390);
nand NAND4 (N8403, N8398, N7685, N2865, N5683);
xor XOR2 (N8404, N8389, N1315);
nor NOR3 (N8405, N8394, N6627, N1603);
nor NOR4 (N8406, N8401, N5629, N1483, N3130);
buf BUF1 (N8407, N8377);
or OR2 (N8408, N8404, N569);
xor XOR2 (N8409, N8405, N5782);
nand NAND4 (N8410, N8407, N7481, N8063, N5918);
nor NOR3 (N8411, N8403, N6874, N3458);
or OR4 (N8412, N8400, N186, N5487, N6960);
nand NAND3 (N8413, N8402, N3095, N7980);
or OR3 (N8414, N8411, N3088, N3150);
and AND4 (N8415, N8414, N8099, N6227, N888);
nor NOR2 (N8416, N8397, N8382);
nor NOR4 (N8417, N8413, N2237, N5194, N2289);
nand NAND2 (N8418, N8385, N3954);
nand NAND3 (N8419, N8418, N4027, N8018);
nor NOR4 (N8420, N8415, N5602, N5887, N6664);
and AND3 (N8421, N8408, N5201, N6717);
buf BUF1 (N8422, N8410);
nand NAND3 (N8423, N8409, N4859, N1474);
nor NOR4 (N8424, N8423, N4220, N181, N4980);
nor NOR3 (N8425, N8417, N2657, N4176);
nand NAND3 (N8426, N8420, N1939, N2543);
or OR2 (N8427, N8419, N3864);
xor XOR2 (N8428, N8391, N4552);
not NOT1 (N8429, N8406);
nand NAND3 (N8430, N8421, N1187, N6312);
and AND4 (N8431, N8430, N7812, N8051, N7997);
nand NAND3 (N8432, N8424, N1109, N4877);
and AND2 (N8433, N8431, N136);
xor XOR2 (N8434, N8432, N5728);
nand NAND2 (N8435, N8425, N7135);
and AND2 (N8436, N8426, N3888);
nor NOR3 (N8437, N8416, N1601, N1889);
not NOT1 (N8438, N8422);
nor NOR3 (N8439, N8436, N1320, N8026);
and AND4 (N8440, N8437, N3673, N3683, N4989);
buf BUF1 (N8441, N8433);
or OR3 (N8442, N8429, N1129, N4648);
nor NOR4 (N8443, N8428, N6913, N1516, N8362);
nor NOR2 (N8444, N8427, N4641);
not NOT1 (N8445, N8440);
xor XOR2 (N8446, N8439, N3032);
and AND3 (N8447, N8434, N2478, N4314);
and AND4 (N8448, N8412, N560, N4838, N1269);
buf BUF1 (N8449, N8438);
xor XOR2 (N8450, N8444, N2049);
not NOT1 (N8451, N8449);
nand NAND4 (N8452, N8447, N8298, N5679, N7669);
buf BUF1 (N8453, N8442);
xor XOR2 (N8454, N8450, N8283);
buf BUF1 (N8455, N8453);
nor NOR2 (N8456, N8452, N8176);
or OR4 (N8457, N8445, N56, N3979, N485);
buf BUF1 (N8458, N8448);
and AND3 (N8459, N8456, N4563, N3091);
nor NOR3 (N8460, N8454, N747, N1732);
nand NAND4 (N8461, N8460, N3831, N5869, N6979);
not NOT1 (N8462, N8441);
not NOT1 (N8463, N8461);
or OR2 (N8464, N8435, N7139);
not NOT1 (N8465, N8457);
nand NAND2 (N8466, N8463, N964);
xor XOR2 (N8467, N8462, N6935);
and AND3 (N8468, N8464, N1424, N5070);
xor XOR2 (N8469, N8451, N4159);
nand NAND2 (N8470, N8469, N575);
nor NOR3 (N8471, N8455, N7338, N926);
nand NAND4 (N8472, N8458, N60, N4170, N5640);
nand NAND4 (N8473, N8466, N5460, N7134, N7551);
nand NAND4 (N8474, N8473, N3559, N5007, N971);
not NOT1 (N8475, N8467);
and AND2 (N8476, N8446, N1775);
buf BUF1 (N8477, N8476);
nor NOR3 (N8478, N8470, N3042, N2848);
or OR2 (N8479, N8474, N3439);
nand NAND2 (N8480, N8443, N7859);
nand NAND4 (N8481, N8478, N1066, N4754, N3175);
or OR2 (N8482, N8468, N1009);
or OR2 (N8483, N8459, N1947);
and AND4 (N8484, N8482, N158, N4909, N1501);
and AND2 (N8485, N8471, N4523);
or OR2 (N8486, N8475, N3642);
nand NAND2 (N8487, N8486, N3635);
or OR2 (N8488, N8480, N78);
nand NAND3 (N8489, N8465, N103, N3518);
xor XOR2 (N8490, N8489, N4885);
buf BUF1 (N8491, N8483);
and AND2 (N8492, N8481, N6893);
not NOT1 (N8493, N8485);
xor XOR2 (N8494, N8487, N8253);
buf BUF1 (N8495, N8472);
not NOT1 (N8496, N8490);
and AND2 (N8497, N8496, N5851);
nand NAND2 (N8498, N8491, N44);
nor NOR2 (N8499, N8488, N4710);
not NOT1 (N8500, N8484);
and AND4 (N8501, N8500, N6546, N7098, N2919);
xor XOR2 (N8502, N8494, N4103);
or OR3 (N8503, N8492, N3465, N5916);
not NOT1 (N8504, N8493);
xor XOR2 (N8505, N8497, N2009);
nor NOR2 (N8506, N8479, N1246);
nand NAND4 (N8507, N8502, N7108, N929, N5544);
nand NAND4 (N8508, N8503, N5620, N6409, N5767);
nor NOR3 (N8509, N8507, N1218, N7992);
nand NAND2 (N8510, N8505, N8416);
buf BUF1 (N8511, N8506);
xor XOR2 (N8512, N8509, N2484);
not NOT1 (N8513, N8498);
and AND3 (N8514, N8513, N3141, N298);
and AND4 (N8515, N8477, N5380, N7215, N991);
nor NOR3 (N8516, N8512, N54, N1939);
not NOT1 (N8517, N8495);
and AND2 (N8518, N8515, N7176);
buf BUF1 (N8519, N8510);
nand NAND2 (N8520, N8504, N897);
xor XOR2 (N8521, N8508, N888);
not NOT1 (N8522, N8501);
xor XOR2 (N8523, N8521, N7749);
buf BUF1 (N8524, N8514);
buf BUF1 (N8525, N8499);
and AND4 (N8526, N8525, N6368, N7178, N7361);
nand NAND2 (N8527, N8517, N6486);
or OR2 (N8528, N8526, N3139);
and AND3 (N8529, N8528, N2992, N2238);
xor XOR2 (N8530, N8523, N2295);
or OR2 (N8531, N8524, N5100);
buf BUF1 (N8532, N8511);
xor XOR2 (N8533, N8530, N5022);
nor NOR2 (N8534, N8516, N5945);
nor NOR2 (N8535, N8527, N4729);
and AND4 (N8536, N8534, N4259, N1366, N8376);
nand NAND4 (N8537, N8520, N31, N2433, N579);
or OR4 (N8538, N8531, N6846, N6622, N2140);
xor XOR2 (N8539, N8537, N645);
nand NAND4 (N8540, N8522, N193, N2370, N2606);
and AND4 (N8541, N8529, N5970, N5805, N7922);
not NOT1 (N8542, N8518);
not NOT1 (N8543, N8538);
or OR2 (N8544, N8539, N5929);
buf BUF1 (N8545, N8533);
nor NOR4 (N8546, N8540, N6784, N3404, N4220);
and AND4 (N8547, N8541, N7759, N4899, N5637);
or OR2 (N8548, N8543, N162);
or OR4 (N8549, N8536, N786, N4330, N1034);
buf BUF1 (N8550, N8547);
nor NOR4 (N8551, N8549, N7374, N1682, N1772);
nor NOR3 (N8552, N8550, N7063, N6167);
xor XOR2 (N8553, N8544, N141);
nor NOR4 (N8554, N8546, N4749, N4336, N864);
xor XOR2 (N8555, N8532, N4324);
nor NOR3 (N8556, N8519, N519, N5597);
or OR2 (N8557, N8545, N7105);
nor NOR3 (N8558, N8554, N3656, N5068);
buf BUF1 (N8559, N8553);
nor NOR4 (N8560, N8548, N5117, N7143, N915);
nor NOR4 (N8561, N8552, N8252, N3161, N7534);
not NOT1 (N8562, N8535);
and AND4 (N8563, N8558, N4209, N4054, N2933);
xor XOR2 (N8564, N8556, N1866);
not NOT1 (N8565, N8563);
or OR2 (N8566, N8562, N3435);
xor XOR2 (N8567, N8564, N6587);
nand NAND4 (N8568, N8542, N4352, N5308, N2784);
not NOT1 (N8569, N8560);
xor XOR2 (N8570, N8565, N2848);
xor XOR2 (N8571, N8555, N58);
not NOT1 (N8572, N8570);
buf BUF1 (N8573, N8567);
nor NOR3 (N8574, N8571, N793, N1446);
and AND2 (N8575, N8561, N2599);
and AND2 (N8576, N8569, N2817);
nor NOR3 (N8577, N8568, N2904, N4056);
nor NOR2 (N8578, N8557, N4852);
buf BUF1 (N8579, N8574);
nor NOR3 (N8580, N8551, N1699, N7099);
and AND2 (N8581, N8577, N7507);
xor XOR2 (N8582, N8572, N5023);
buf BUF1 (N8583, N8580);
nand NAND2 (N8584, N8573, N5538);
nor NOR2 (N8585, N8583, N1129);
xor XOR2 (N8586, N8576, N710);
and AND3 (N8587, N8566, N6145, N4465);
nor NOR4 (N8588, N8587, N380, N1447, N5994);
nand NAND3 (N8589, N8588, N4707, N6671);
xor XOR2 (N8590, N8585, N1152);
not NOT1 (N8591, N8559);
and AND4 (N8592, N8581, N6218, N5217, N3459);
buf BUF1 (N8593, N8582);
not NOT1 (N8594, N8575);
nand NAND2 (N8595, N8593, N6610);
xor XOR2 (N8596, N8578, N143);
or OR2 (N8597, N8579, N8062);
not NOT1 (N8598, N8596);
not NOT1 (N8599, N8594);
nand NAND4 (N8600, N8590, N1008, N4043, N6441);
buf BUF1 (N8601, N8595);
and AND3 (N8602, N8600, N3357, N1455);
nor NOR2 (N8603, N8601, N1439);
buf BUF1 (N8604, N8586);
buf BUF1 (N8605, N8597);
not NOT1 (N8606, N8592);
and AND3 (N8607, N8584, N5811, N663);
buf BUF1 (N8608, N8599);
not NOT1 (N8609, N8605);
or OR2 (N8610, N8604, N3259);
or OR3 (N8611, N8598, N639, N6282);
xor XOR2 (N8612, N8591, N6955);
nand NAND2 (N8613, N8608, N6624);
xor XOR2 (N8614, N8589, N7832);
and AND2 (N8615, N8603, N7817);
nor NOR3 (N8616, N8613, N4640, N2699);
xor XOR2 (N8617, N8610, N2288);
buf BUF1 (N8618, N8602);
xor XOR2 (N8619, N8617, N1769);
and AND4 (N8620, N8609, N136, N8472, N4895);
nand NAND3 (N8621, N8616, N7477, N8470);
buf BUF1 (N8622, N8611);
nor NOR3 (N8623, N8606, N3358, N2706);
not NOT1 (N8624, N8621);
nand NAND4 (N8625, N8607, N5615, N1386, N7506);
xor XOR2 (N8626, N8615, N6941);
buf BUF1 (N8627, N8620);
buf BUF1 (N8628, N8626);
nand NAND4 (N8629, N8618, N4963, N3021, N4713);
or OR3 (N8630, N8612, N1230, N6960);
and AND2 (N8631, N8614, N965);
nand NAND3 (N8632, N8627, N4910, N1131);
or OR3 (N8633, N8619, N6177, N8218);
nand NAND2 (N8634, N8630, N1795);
or OR2 (N8635, N8623, N7047);
not NOT1 (N8636, N8625);
buf BUF1 (N8637, N8632);
buf BUF1 (N8638, N8624);
nor NOR4 (N8639, N8633, N4903, N2395, N7814);
xor XOR2 (N8640, N8635, N5348);
nor NOR2 (N8641, N8628, N5327);
buf BUF1 (N8642, N8641);
nor NOR4 (N8643, N8636, N803, N386, N6990);
not NOT1 (N8644, N8622);
and AND3 (N8645, N8631, N1286, N720);
buf BUF1 (N8646, N8640);
and AND3 (N8647, N8629, N7110, N3194);
not NOT1 (N8648, N8644);
and AND3 (N8649, N8648, N1730, N7770);
nor NOR3 (N8650, N8634, N2237, N1389);
and AND2 (N8651, N8649, N5295);
buf BUF1 (N8652, N8646);
nand NAND4 (N8653, N8639, N3924, N6298, N1118);
and AND3 (N8654, N8651, N2740, N6829);
or OR2 (N8655, N8654, N454);
or OR3 (N8656, N8643, N3191, N772);
and AND3 (N8657, N8650, N8313, N3832);
buf BUF1 (N8658, N8647);
or OR4 (N8659, N8645, N4200, N5533, N8457);
buf BUF1 (N8660, N8657);
nand NAND2 (N8661, N8660, N3845);
nor NOR2 (N8662, N8638, N1105);
and AND3 (N8663, N8637, N6489, N6972);
and AND2 (N8664, N8659, N4777);
buf BUF1 (N8665, N8642);
xor XOR2 (N8666, N8662, N3352);
buf BUF1 (N8667, N8665);
and AND2 (N8668, N8653, N4691);
nor NOR4 (N8669, N8664, N6122, N1761, N68);
not NOT1 (N8670, N8661);
nand NAND3 (N8671, N8669, N7083, N8448);
buf BUF1 (N8672, N8666);
nand NAND4 (N8673, N8656, N5978, N7175, N2761);
or OR3 (N8674, N8663, N7267, N3907);
not NOT1 (N8675, N8671);
and AND3 (N8676, N8675, N3788, N844);
or OR2 (N8677, N8658, N3557);
nand NAND4 (N8678, N8670, N2376, N3211, N3313);
buf BUF1 (N8679, N8678);
and AND2 (N8680, N8679, N1393);
nor NOR3 (N8681, N8676, N7383, N1934);
nor NOR2 (N8682, N8674, N2327);
not NOT1 (N8683, N8672);
nand NAND2 (N8684, N8667, N3703);
not NOT1 (N8685, N8652);
nor NOR3 (N8686, N8680, N175, N7083);
buf BUF1 (N8687, N8668);
and AND4 (N8688, N8682, N4093, N2048, N7520);
nand NAND4 (N8689, N8655, N3352, N284, N3904);
or OR3 (N8690, N8686, N8433, N4833);
not NOT1 (N8691, N8685);
or OR4 (N8692, N8683, N2838, N818, N210);
or OR2 (N8693, N8673, N7782);
or OR3 (N8694, N8692, N5836, N5181);
nor NOR4 (N8695, N8690, N7842, N7340, N1863);
nor NOR2 (N8696, N8693, N5574);
buf BUF1 (N8697, N8696);
xor XOR2 (N8698, N8677, N2905);
buf BUF1 (N8699, N8694);
nand NAND2 (N8700, N8688, N1629);
and AND3 (N8701, N8697, N3717, N5222);
and AND2 (N8702, N8695, N2631);
buf BUF1 (N8703, N8681);
nand NAND2 (N8704, N8699, N7229);
buf BUF1 (N8705, N8691);
or OR3 (N8706, N8698, N1403, N3815);
xor XOR2 (N8707, N8701, N4413);
and AND4 (N8708, N8700, N5921, N2038, N7825);
or OR4 (N8709, N8689, N7795, N1238, N465);
and AND2 (N8710, N8707, N8028);
not NOT1 (N8711, N8708);
and AND2 (N8712, N8710, N3398);
and AND2 (N8713, N8703, N1873);
nor NOR2 (N8714, N8705, N4598);
and AND3 (N8715, N8712, N349, N464);
not NOT1 (N8716, N8706);
nand NAND2 (N8717, N8711, N538);
or OR3 (N8718, N8709, N1015, N2317);
xor XOR2 (N8719, N8684, N2052);
buf BUF1 (N8720, N8687);
not NOT1 (N8721, N8717);
and AND3 (N8722, N8702, N3248, N415);
nand NAND4 (N8723, N8713, N7616, N4238, N8059);
or OR3 (N8724, N8721, N8434, N5910);
and AND4 (N8725, N8724, N5344, N5376, N7519);
nand NAND2 (N8726, N8718, N7168);
and AND3 (N8727, N8704, N3379, N3616);
and AND3 (N8728, N8720, N6468, N4271);
xor XOR2 (N8729, N8715, N5926);
nor NOR3 (N8730, N8714, N8268, N99);
and AND2 (N8731, N8716, N3862);
not NOT1 (N8732, N8719);
xor XOR2 (N8733, N8732, N5007);
xor XOR2 (N8734, N8733, N6920);
buf BUF1 (N8735, N8729);
xor XOR2 (N8736, N8734, N496);
not NOT1 (N8737, N8727);
nor NOR3 (N8738, N8730, N7109, N7640);
xor XOR2 (N8739, N8725, N1766);
xor XOR2 (N8740, N8722, N350);
not NOT1 (N8741, N8739);
or OR3 (N8742, N8738, N8209, N6554);
nor NOR3 (N8743, N8731, N4343, N7562);
and AND3 (N8744, N8726, N830, N8641);
and AND3 (N8745, N8743, N92, N2539);
buf BUF1 (N8746, N8728);
nand NAND4 (N8747, N8735, N7854, N4555, N2811);
nand NAND3 (N8748, N8747, N5033, N772);
nand NAND4 (N8749, N8745, N2498, N5272, N6661);
not NOT1 (N8750, N8723);
buf BUF1 (N8751, N8748);
or OR4 (N8752, N8751, N5934, N2394, N5375);
nor NOR3 (N8753, N8744, N5759, N7300);
not NOT1 (N8754, N8742);
buf BUF1 (N8755, N8741);
xor XOR2 (N8756, N8736, N7870);
xor XOR2 (N8757, N8752, N6344);
xor XOR2 (N8758, N8753, N1121);
xor XOR2 (N8759, N8750, N6045);
nor NOR2 (N8760, N8758, N4108);
xor XOR2 (N8761, N8737, N5385);
or OR4 (N8762, N8754, N626, N7936, N5146);
xor XOR2 (N8763, N8749, N3931);
or OR2 (N8764, N8757, N2382);
not NOT1 (N8765, N8764);
not NOT1 (N8766, N8746);
nor NOR4 (N8767, N8763, N7498, N6251, N3353);
xor XOR2 (N8768, N8759, N8091);
or OR3 (N8769, N8761, N1258, N3109);
and AND2 (N8770, N8760, N7170);
nand NAND4 (N8771, N8769, N1928, N3641, N6667);
not NOT1 (N8772, N8756);
not NOT1 (N8773, N8770);
buf BUF1 (N8774, N8767);
nor NOR3 (N8775, N8773, N6351, N7099);
or OR2 (N8776, N8755, N2327);
not NOT1 (N8777, N8766);
buf BUF1 (N8778, N8765);
nor NOR2 (N8779, N8774, N3515);
buf BUF1 (N8780, N8768);
nor NOR4 (N8781, N8771, N2904, N229, N2716);
buf BUF1 (N8782, N8780);
nor NOR2 (N8783, N8777, N3711);
nor NOR4 (N8784, N8782, N843, N3995, N4985);
not NOT1 (N8785, N8784);
or OR4 (N8786, N8779, N6546, N3375, N557);
and AND4 (N8787, N8778, N6867, N591, N4994);
buf BUF1 (N8788, N8762);
buf BUF1 (N8789, N8740);
and AND2 (N8790, N8772, N692);
or OR4 (N8791, N8776, N388, N8248, N2966);
or OR2 (N8792, N8781, N5996);
not NOT1 (N8793, N8788);
nor NOR2 (N8794, N8785, N2313);
and AND3 (N8795, N8790, N3719, N8272);
nor NOR2 (N8796, N8789, N6770);
nor NOR2 (N8797, N8791, N4970);
not NOT1 (N8798, N8786);
not NOT1 (N8799, N8798);
xor XOR2 (N8800, N8787, N4571);
xor XOR2 (N8801, N8793, N8705);
and AND4 (N8802, N8795, N7854, N6252, N8195);
xor XOR2 (N8803, N8794, N6117);
xor XOR2 (N8804, N8797, N11);
xor XOR2 (N8805, N8796, N7021);
nor NOR4 (N8806, N8792, N7487, N5691, N7276);
and AND4 (N8807, N8783, N4269, N8470, N6532);
not NOT1 (N8808, N8775);
and AND2 (N8809, N8802, N1073);
xor XOR2 (N8810, N8806, N7993);
and AND4 (N8811, N8810, N6803, N920, N4162);
and AND2 (N8812, N8805, N3061);
nor NOR3 (N8813, N8807, N1237, N2121);
not NOT1 (N8814, N8804);
and AND3 (N8815, N8813, N4131, N171);
not NOT1 (N8816, N8800);
xor XOR2 (N8817, N8801, N5157);
xor XOR2 (N8818, N8812, N3862);
buf BUF1 (N8819, N8817);
xor XOR2 (N8820, N8809, N8631);
buf BUF1 (N8821, N8811);
xor XOR2 (N8822, N8814, N950);
or OR3 (N8823, N8799, N70, N3368);
nor NOR2 (N8824, N8820, N2951);
or OR2 (N8825, N8815, N3273);
buf BUF1 (N8826, N8823);
and AND3 (N8827, N8821, N3812, N1791);
not NOT1 (N8828, N8827);
or OR4 (N8829, N8828, N4039, N8111, N4318);
nand NAND4 (N8830, N8824, N3204, N2319, N8827);
buf BUF1 (N8831, N8803);
nor NOR2 (N8832, N8829, N6361);
xor XOR2 (N8833, N8831, N7849);
and AND4 (N8834, N8808, N339, N8256, N4618);
not NOT1 (N8835, N8816);
and AND4 (N8836, N8834, N1982, N7116, N3401);
buf BUF1 (N8837, N8822);
or OR3 (N8838, N8836, N3024, N7916);
or OR2 (N8839, N8833, N7803);
nand NAND2 (N8840, N8818, N1573);
buf BUF1 (N8841, N8838);
nand NAND3 (N8842, N8839, N2391, N2193);
not NOT1 (N8843, N8840);
and AND2 (N8844, N8843, N3480);
not NOT1 (N8845, N8842);
or OR4 (N8846, N8832, N731, N7525, N4294);
and AND4 (N8847, N8837, N5676, N1685, N1769);
not NOT1 (N8848, N8841);
buf BUF1 (N8849, N8845);
buf BUF1 (N8850, N8844);
or OR3 (N8851, N8846, N2663, N2134);
not NOT1 (N8852, N8825);
buf BUF1 (N8853, N8826);
nor NOR4 (N8854, N8819, N8845, N7934, N4819);
buf BUF1 (N8855, N8850);
nor NOR4 (N8856, N8855, N3042, N2316, N1889);
and AND2 (N8857, N8856, N3526);
not NOT1 (N8858, N8854);
nand NAND4 (N8859, N8857, N2895, N3965, N8713);
not NOT1 (N8860, N8830);
and AND3 (N8861, N8852, N4591, N5092);
not NOT1 (N8862, N8860);
or OR3 (N8863, N8858, N3479, N73);
or OR2 (N8864, N8847, N5977);
nand NAND3 (N8865, N8863, N5101, N3353);
nor NOR2 (N8866, N8848, N2826);
nand NAND2 (N8867, N8862, N3837);
or OR3 (N8868, N8866, N4775, N7515);
xor XOR2 (N8869, N8861, N7097);
buf BUF1 (N8870, N8853);
and AND4 (N8871, N8859, N1351, N1357, N2658);
buf BUF1 (N8872, N8865);
not NOT1 (N8873, N8849);
and AND2 (N8874, N8870, N6013);
buf BUF1 (N8875, N8869);
nor NOR4 (N8876, N8874, N5063, N6485, N4003);
nor NOR2 (N8877, N8864, N5984);
nor NOR2 (N8878, N8876, N3154);
and AND2 (N8879, N8835, N5984);
not NOT1 (N8880, N8877);
and AND3 (N8881, N8851, N4171, N85);
xor XOR2 (N8882, N8878, N2064);
buf BUF1 (N8883, N8881);
nor NOR3 (N8884, N8882, N5571, N2450);
not NOT1 (N8885, N8867);
nand NAND4 (N8886, N8884, N6540, N7430, N4895);
xor XOR2 (N8887, N8879, N4472);
xor XOR2 (N8888, N8885, N7153);
nand NAND2 (N8889, N8888, N8706);
xor XOR2 (N8890, N8868, N4498);
and AND2 (N8891, N8889, N6525);
not NOT1 (N8892, N8875);
not NOT1 (N8893, N8891);
or OR2 (N8894, N8892, N5835);
nand NAND3 (N8895, N8872, N2796, N7286);
not NOT1 (N8896, N8890);
nor NOR3 (N8897, N8871, N2083, N3670);
nand NAND2 (N8898, N8895, N3363);
buf BUF1 (N8899, N8886);
not NOT1 (N8900, N8873);
and AND4 (N8901, N8887, N4548, N1762, N4960);
nand NAND4 (N8902, N8899, N3280, N3107, N5652);
and AND4 (N8903, N8896, N1023, N6319, N1701);
buf BUF1 (N8904, N8901);
not NOT1 (N8905, N8894);
nor NOR2 (N8906, N8880, N7632);
or OR4 (N8907, N8904, N4127, N8055, N2079);
or OR4 (N8908, N8907, N2586, N5530, N8789);
nand NAND2 (N8909, N8900, N3379);
xor XOR2 (N8910, N8898, N6113);
xor XOR2 (N8911, N8905, N7846);
xor XOR2 (N8912, N8883, N1222);
or OR3 (N8913, N8908, N7184, N5287);
not NOT1 (N8914, N8909);
nand NAND4 (N8915, N8910, N6570, N3189, N7644);
buf BUF1 (N8916, N8911);
or OR4 (N8917, N8893, N7134, N4401, N5609);
and AND3 (N8918, N8906, N5757, N8811);
buf BUF1 (N8919, N8914);
buf BUF1 (N8920, N8903);
and AND4 (N8921, N8913, N6435, N472, N1054);
not NOT1 (N8922, N8917);
nor NOR2 (N8923, N8918, N8759);
nand NAND4 (N8924, N8912, N1901, N5412, N4438);
buf BUF1 (N8925, N8922);
nand NAND3 (N8926, N8923, N7645, N5812);
xor XOR2 (N8927, N8902, N4995);
and AND3 (N8928, N8919, N5048, N2459);
and AND3 (N8929, N8927, N8092, N4402);
and AND2 (N8930, N8921, N6469);
not NOT1 (N8931, N8930);
buf BUF1 (N8932, N8916);
buf BUF1 (N8933, N8932);
nor NOR3 (N8934, N8915, N8133, N6988);
nor NOR3 (N8935, N8934, N5457, N1734);
not NOT1 (N8936, N8925);
not NOT1 (N8937, N8920);
not NOT1 (N8938, N8931);
nand NAND4 (N8939, N8924, N4644, N7871, N2170);
or OR2 (N8940, N8926, N6888);
buf BUF1 (N8941, N8939);
or OR4 (N8942, N8936, N1911, N8521, N4191);
or OR3 (N8943, N8897, N2190, N8850);
nor NOR2 (N8944, N8941, N1667);
and AND2 (N8945, N8937, N1716);
or OR3 (N8946, N8943, N4723, N3332);
or OR4 (N8947, N8945, N7518, N7125, N5761);
nand NAND2 (N8948, N8946, N3403);
buf BUF1 (N8949, N8938);
or OR2 (N8950, N8933, N4150);
and AND4 (N8951, N8947, N8026, N4408, N8442);
buf BUF1 (N8952, N8942);
buf BUF1 (N8953, N8940);
nand NAND4 (N8954, N8935, N2438, N5131, N5916);
and AND2 (N8955, N8928, N2474);
or OR3 (N8956, N8951, N1585, N1593);
or OR4 (N8957, N8949, N2493, N7021, N6680);
nand NAND3 (N8958, N8954, N3937, N5511);
xor XOR2 (N8959, N8948, N933);
nor NOR4 (N8960, N8956, N4719, N6781, N5587);
nor NOR4 (N8961, N8959, N8422, N8812, N359);
or OR3 (N8962, N8953, N8237, N2507);
buf BUF1 (N8963, N8960);
and AND3 (N8964, N8962, N7959, N8507);
buf BUF1 (N8965, N8961);
or OR2 (N8966, N8952, N4416);
nor NOR3 (N8967, N8964, N8246, N8137);
nor NOR2 (N8968, N8966, N5914);
and AND2 (N8969, N8967, N8186);
nor NOR4 (N8970, N8929, N6028, N7152, N6261);
nand NAND3 (N8971, N8970, N5154, N1363);
or OR2 (N8972, N8969, N4912);
or OR4 (N8973, N8971, N1136, N1252, N4187);
and AND2 (N8974, N8955, N8640);
nand NAND3 (N8975, N8973, N8411, N5036);
buf BUF1 (N8976, N8958);
and AND3 (N8977, N8963, N8633, N6701);
not NOT1 (N8978, N8972);
buf BUF1 (N8979, N8950);
nand NAND2 (N8980, N8979, N27);
nand NAND4 (N8981, N8974, N1047, N3274, N2933);
or OR4 (N8982, N8976, N8127, N2984, N7987);
xor XOR2 (N8983, N8944, N5361);
or OR2 (N8984, N8975, N3244);
buf BUF1 (N8985, N8982);
buf BUF1 (N8986, N8985);
buf BUF1 (N8987, N8984);
nor NOR4 (N8988, N8965, N6675, N6768, N7605);
nand NAND2 (N8989, N8968, N3059);
not NOT1 (N8990, N8988);
nor NOR2 (N8991, N8990, N249);
nand NAND3 (N8992, N8981, N4376, N4477);
nand NAND3 (N8993, N8957, N1485, N1440);
buf BUF1 (N8994, N8986);
xor XOR2 (N8995, N8980, N4155);
nand NAND2 (N8996, N8989, N3366);
nand NAND4 (N8997, N8995, N930, N4114, N6303);
and AND2 (N8998, N8993, N1514);
buf BUF1 (N8999, N8991);
and AND3 (N9000, N8999, N5677, N414);
xor XOR2 (N9001, N8992, N2049);
xor XOR2 (N9002, N8978, N3224);
buf BUF1 (N9003, N8987);
xor XOR2 (N9004, N9003, N2698);
or OR2 (N9005, N8996, N5982);
and AND2 (N9006, N8983, N4039);
nand NAND3 (N9007, N8998, N6071, N7590);
and AND3 (N9008, N9000, N6678, N789);
nor NOR3 (N9009, N9008, N8644, N1123);
not NOT1 (N9010, N9001);
nand NAND3 (N9011, N8997, N7151, N4315);
nand NAND2 (N9012, N8994, N6404);
xor XOR2 (N9013, N9009, N5694);
nor NOR4 (N9014, N9010, N1801, N1719, N2089);
xor XOR2 (N9015, N9007, N1818);
not NOT1 (N9016, N8977);
xor XOR2 (N9017, N9006, N3146);
and AND3 (N9018, N9016, N660, N4128);
nor NOR3 (N9019, N9013, N8194, N3380);
not NOT1 (N9020, N9002);
xor XOR2 (N9021, N9019, N5523);
nand NAND2 (N9022, N9005, N241);
nand NAND2 (N9023, N9017, N7562);
and AND4 (N9024, N9022, N7115, N3192, N8773);
or OR4 (N9025, N9023, N5721, N8561, N1270);
not NOT1 (N9026, N9012);
or OR3 (N9027, N9020, N3952, N5434);
buf BUF1 (N9028, N9021);
not NOT1 (N9029, N9018);
or OR4 (N9030, N9027, N5686, N5944, N1391);
or OR3 (N9031, N9004, N4256, N6440);
nor NOR3 (N9032, N9014, N4985, N3710);
buf BUF1 (N9033, N9031);
not NOT1 (N9034, N9028);
nor NOR2 (N9035, N9015, N5844);
nor NOR4 (N9036, N9024, N2238, N5691, N8977);
buf BUF1 (N9037, N9030);
xor XOR2 (N9038, N9011, N1676);
not NOT1 (N9039, N9032);
or OR3 (N9040, N9029, N2639, N889);
xor XOR2 (N9041, N9038, N7410);
nand NAND2 (N9042, N9026, N5504);
not NOT1 (N9043, N9041);
buf BUF1 (N9044, N9034);
nor NOR2 (N9045, N9025, N2617);
and AND4 (N9046, N9040, N3356, N1526, N5932);
or OR2 (N9047, N9044, N6271);
nor NOR4 (N9048, N9037, N541, N6157, N3505);
buf BUF1 (N9049, N9048);
nor NOR3 (N9050, N9033, N5028, N5868);
buf BUF1 (N9051, N9035);
or OR4 (N9052, N9045, N8122, N1052, N1137);
and AND4 (N9053, N9049, N2543, N7873, N6359);
or OR3 (N9054, N9053, N6046, N7647);
not NOT1 (N9055, N9047);
and AND4 (N9056, N9039, N7327, N8461, N859);
nand NAND3 (N9057, N9054, N6060, N6967);
nand NAND2 (N9058, N9043, N3511);
buf BUF1 (N9059, N9055);
or OR2 (N9060, N9050, N3624);
nand NAND3 (N9061, N9058, N6148, N8986);
nor NOR4 (N9062, N9057, N4334, N6286, N7104);
buf BUF1 (N9063, N9042);
buf BUF1 (N9064, N9046);
not NOT1 (N9065, N9063);
and AND3 (N9066, N9065, N6054, N7003);
nand NAND2 (N9067, N9061, N5933);
buf BUF1 (N9068, N9064);
nor NOR2 (N9069, N9060, N2368);
or OR3 (N9070, N9051, N1779, N4441);
xor XOR2 (N9071, N9069, N5042);
or OR3 (N9072, N9059, N2746, N5168);
or OR4 (N9073, N9066, N2212, N2931, N287);
nand NAND2 (N9074, N9062, N4865);
and AND4 (N9075, N9068, N8939, N672, N4479);
buf BUF1 (N9076, N9070);
or OR2 (N9077, N9052, N1175);
xor XOR2 (N9078, N9072, N5175);
or OR4 (N9079, N9036, N603, N5694, N7929);
and AND4 (N9080, N9071, N4249, N6444, N3352);
nor NOR2 (N9081, N9080, N4064);
not NOT1 (N9082, N9081);
not NOT1 (N9083, N9056);
nand NAND4 (N9084, N9076, N6067, N3498, N5577);
nand NAND2 (N9085, N9075, N298);
not NOT1 (N9086, N9077);
not NOT1 (N9087, N9074);
or OR2 (N9088, N9086, N806);
not NOT1 (N9089, N9088);
buf BUF1 (N9090, N9085);
nor NOR4 (N9091, N9083, N7233, N7478, N4323);
nor NOR3 (N9092, N9087, N3017, N6535);
nand NAND4 (N9093, N9082, N3171, N7821, N1435);
not NOT1 (N9094, N9093);
buf BUF1 (N9095, N9084);
or OR3 (N9096, N9095, N1999, N3741);
not NOT1 (N9097, N9091);
not NOT1 (N9098, N9096);
buf BUF1 (N9099, N9090);
not NOT1 (N9100, N9092);
or OR3 (N9101, N9100, N3833, N6112);
nand NAND4 (N9102, N9078, N7988, N1160, N4416);
or OR3 (N9103, N9079, N4271, N7546);
nor NOR2 (N9104, N9098, N3913);
buf BUF1 (N9105, N9067);
xor XOR2 (N9106, N9089, N663);
nand NAND3 (N9107, N9106, N2214, N5224);
buf BUF1 (N9108, N9105);
or OR4 (N9109, N9099, N3046, N5017, N2936);
not NOT1 (N9110, N9104);
xor XOR2 (N9111, N9094, N3930);
and AND2 (N9112, N9101, N5204);
or OR4 (N9113, N9097, N6898, N7336, N8486);
nor NOR4 (N9114, N9108, N328, N8265, N7844);
xor XOR2 (N9115, N9102, N412);
nand NAND3 (N9116, N9115, N5075, N7808);
and AND4 (N9117, N9112, N8029, N5339, N6862);
and AND3 (N9118, N9117, N7572, N3328);
nand NAND3 (N9119, N9109, N3986, N6853);
nand NAND4 (N9120, N9116, N6665, N4956, N7130);
nor NOR3 (N9121, N9073, N868, N6897);
nand NAND4 (N9122, N9110, N1195, N4821, N8187);
nor NOR2 (N9123, N9103, N2483);
and AND2 (N9124, N9120, N350);
or OR3 (N9125, N9123, N6479, N2880);
buf BUF1 (N9126, N9111);
buf BUF1 (N9127, N9119);
not NOT1 (N9128, N9127);
and AND4 (N9129, N9121, N8673, N3179, N881);
or OR4 (N9130, N9126, N6176, N1321, N1423);
and AND3 (N9131, N9128, N6528, N7535);
buf BUF1 (N9132, N9107);
buf BUF1 (N9133, N9113);
xor XOR2 (N9134, N9124, N4071);
nor NOR2 (N9135, N9125, N5679);
nand NAND4 (N9136, N9131, N1499, N1648, N1174);
and AND3 (N9137, N9129, N5996, N4266);
and AND3 (N9138, N9136, N8297, N1297);
nor NOR4 (N9139, N9133, N4555, N4459, N2149);
and AND3 (N9140, N9135, N3670, N3840);
nor NOR2 (N9141, N9137, N4733);
buf BUF1 (N9142, N9139);
xor XOR2 (N9143, N9122, N5764);
not NOT1 (N9144, N9118);
not NOT1 (N9145, N9114);
nor NOR4 (N9146, N9134, N6716, N6027, N5056);
nand NAND3 (N9147, N9132, N5842, N6739);
nor NOR4 (N9148, N9130, N6302, N4611, N6115);
nor NOR4 (N9149, N9141, N275, N3718, N1125);
xor XOR2 (N9150, N9142, N4335);
nor NOR4 (N9151, N9140, N4245, N1568, N3307);
not NOT1 (N9152, N9148);
and AND3 (N9153, N9150, N5496, N3708);
nor NOR4 (N9154, N9145, N8176, N3696, N8424);
buf BUF1 (N9155, N9153);
xor XOR2 (N9156, N9151, N4139);
nand NAND2 (N9157, N9155, N6109);
buf BUF1 (N9158, N9143);
or OR2 (N9159, N9156, N3091);
nand NAND3 (N9160, N9144, N2305, N5046);
nand NAND3 (N9161, N9146, N820, N801);
nor NOR2 (N9162, N9159, N943);
xor XOR2 (N9163, N9138, N7150);
or OR2 (N9164, N9163, N3323);
nand NAND3 (N9165, N9152, N327, N2184);
xor XOR2 (N9166, N9154, N6989);
or OR2 (N9167, N9161, N7402);
not NOT1 (N9168, N9164);
or OR3 (N9169, N9149, N1930, N1702);
nor NOR3 (N9170, N9157, N7975, N2334);
not NOT1 (N9171, N9158);
and AND2 (N9172, N9147, N4350);
or OR3 (N9173, N9168, N2261, N1965);
nand NAND3 (N9174, N9166, N736, N2477);
or OR3 (N9175, N9171, N9089, N2002);
not NOT1 (N9176, N9162);
nor NOR3 (N9177, N9169, N7772, N8331);
buf BUF1 (N9178, N9173);
not NOT1 (N9179, N9170);
not NOT1 (N9180, N9167);
not NOT1 (N9181, N9176);
buf BUF1 (N9182, N9165);
buf BUF1 (N9183, N9175);
nand NAND2 (N9184, N9182, N9111);
buf BUF1 (N9185, N9181);
not NOT1 (N9186, N9172);
buf BUF1 (N9187, N9186);
xor XOR2 (N9188, N9179, N5018);
nor NOR4 (N9189, N9177, N2588, N1369, N3838);
xor XOR2 (N9190, N9160, N2682);
nand NAND2 (N9191, N9190, N1311);
nand NAND4 (N9192, N9188, N6870, N3603, N3954);
or OR4 (N9193, N9180, N9000, N8419, N7752);
not NOT1 (N9194, N9191);
buf BUF1 (N9195, N9183);
or OR2 (N9196, N9187, N2204);
nand NAND3 (N9197, N9196, N4459, N8813);
nand NAND3 (N9198, N9174, N8952, N3700);
and AND3 (N9199, N9178, N5545, N4989);
nand NAND3 (N9200, N9192, N7130, N5395);
nand NAND3 (N9201, N9197, N8895, N8985);
nand NAND3 (N9202, N9199, N3026, N7981);
nand NAND3 (N9203, N9194, N3652, N1305);
not NOT1 (N9204, N9195);
not NOT1 (N9205, N9204);
nand NAND2 (N9206, N9202, N3766);
nor NOR2 (N9207, N9189, N1020);
buf BUF1 (N9208, N9193);
or OR4 (N9209, N9208, N7919, N7800, N8442);
buf BUF1 (N9210, N9203);
nand NAND2 (N9211, N9185, N5272);
buf BUF1 (N9212, N9184);
or OR4 (N9213, N9205, N9014, N2980, N5388);
nor NOR4 (N9214, N9212, N4564, N6274, N5328);
nand NAND4 (N9215, N9201, N6745, N4888, N4930);
xor XOR2 (N9216, N9200, N4877);
nor NOR2 (N9217, N9206, N7733);
not NOT1 (N9218, N9209);
buf BUF1 (N9219, N9211);
buf BUF1 (N9220, N9213);
not NOT1 (N9221, N9220);
and AND2 (N9222, N9221, N8890);
buf BUF1 (N9223, N9198);
and AND2 (N9224, N9217, N8208);
not NOT1 (N9225, N9210);
or OR3 (N9226, N9222, N1724, N5109);
nor NOR4 (N9227, N9225, N3254, N5101, N7221);
nor NOR2 (N9228, N9219, N1652);
and AND4 (N9229, N9215, N3563, N5199, N5493);
or OR3 (N9230, N9224, N8299, N7093);
not NOT1 (N9231, N9230);
buf BUF1 (N9232, N9231);
nand NAND4 (N9233, N9223, N2077, N4638, N4164);
and AND3 (N9234, N9229, N146, N7368);
nor NOR3 (N9235, N9218, N2793, N8188);
buf BUF1 (N9236, N9232);
nor NOR3 (N9237, N9233, N3915, N4748);
nor NOR2 (N9238, N9227, N914);
nor NOR3 (N9239, N9234, N8315, N2657);
xor XOR2 (N9240, N9235, N511);
not NOT1 (N9241, N9216);
nor NOR4 (N9242, N9236, N8180, N5514, N116);
nor NOR3 (N9243, N9207, N565, N9024);
buf BUF1 (N9244, N9228);
nand NAND4 (N9245, N9242, N3769, N3147, N214);
or OR2 (N9246, N9245, N7985);
xor XOR2 (N9247, N9243, N1904);
nand NAND3 (N9248, N9246, N5963, N8541);
buf BUF1 (N9249, N9239);
nor NOR2 (N9250, N9214, N4960);
xor XOR2 (N9251, N9238, N3917);
and AND2 (N9252, N9244, N8250);
not NOT1 (N9253, N9251);
xor XOR2 (N9254, N9247, N5343);
nor NOR4 (N9255, N9250, N5892, N7901, N4029);
and AND4 (N9256, N9241, N1913, N9183, N5628);
or OR2 (N9257, N9256, N6697);
or OR4 (N9258, N9253, N1179, N6930, N8655);
and AND4 (N9259, N9226, N742, N1951, N6297);
or OR2 (N9260, N9252, N2580);
nor NOR2 (N9261, N9249, N6517);
nor NOR3 (N9262, N9260, N562, N4030);
or OR2 (N9263, N9258, N536);
xor XOR2 (N9264, N9237, N2204);
xor XOR2 (N9265, N9248, N3303);
buf BUF1 (N9266, N9255);
nor NOR2 (N9267, N9262, N6683);
xor XOR2 (N9268, N9266, N7920);
buf BUF1 (N9269, N9254);
buf BUF1 (N9270, N9263);
nand NAND4 (N9271, N9265, N3366, N3675, N2185);
nor NOR2 (N9272, N9270, N6313);
xor XOR2 (N9273, N9257, N8387);
buf BUF1 (N9274, N9261);
xor XOR2 (N9275, N9269, N3759);
buf BUF1 (N9276, N9267);
nand NAND4 (N9277, N9271, N3451, N8370, N5647);
not NOT1 (N9278, N9264);
nand NAND4 (N9279, N9276, N3532, N1886, N2754);
not NOT1 (N9280, N9274);
buf BUF1 (N9281, N9277);
not NOT1 (N9282, N9272);
or OR3 (N9283, N9275, N4628, N522);
not NOT1 (N9284, N9281);
or OR3 (N9285, N9282, N1413, N7980);
nand NAND3 (N9286, N9278, N4864, N1077);
nor NOR3 (N9287, N9283, N1955, N6624);
and AND2 (N9288, N9284, N7719);
nor NOR4 (N9289, N9268, N1740, N5179, N1786);
nand NAND2 (N9290, N9240, N9008);
or OR4 (N9291, N9285, N3473, N5677, N9127);
or OR4 (N9292, N9289, N7888, N3784, N5013);
xor XOR2 (N9293, N9292, N4599);
nor NOR4 (N9294, N9273, N2740, N5926, N1586);
not NOT1 (N9295, N9290);
buf BUF1 (N9296, N9280);
xor XOR2 (N9297, N9279, N6880);
not NOT1 (N9298, N9293);
xor XOR2 (N9299, N9287, N8949);
nor NOR4 (N9300, N9294, N5670, N1639, N3212);
nor NOR4 (N9301, N9291, N1521, N3832, N8333);
or OR3 (N9302, N9298, N5465, N6990);
xor XOR2 (N9303, N9295, N7546);
nand NAND2 (N9304, N9299, N6213);
xor XOR2 (N9305, N9302, N3099);
nand NAND2 (N9306, N9301, N4009);
or OR3 (N9307, N9303, N6048, N9193);
and AND2 (N9308, N9307, N6080);
or OR3 (N9309, N9297, N6503, N8370);
buf BUF1 (N9310, N9309);
xor XOR2 (N9311, N9305, N9104);
xor XOR2 (N9312, N9304, N7478);
buf BUF1 (N9313, N9306);
nand NAND4 (N9314, N9313, N4326, N3946, N4391);
xor XOR2 (N9315, N9311, N2210);
nand NAND3 (N9316, N9286, N1155, N4717);
not NOT1 (N9317, N9288);
and AND4 (N9318, N9317, N4835, N6956, N4148);
xor XOR2 (N9319, N9315, N7808);
not NOT1 (N9320, N9296);
nor NOR4 (N9321, N9300, N2981, N873, N836);
or OR2 (N9322, N9310, N1514);
nand NAND4 (N9323, N9320, N4214, N8234, N6606);
nand NAND2 (N9324, N9314, N2848);
nor NOR4 (N9325, N9321, N3285, N4273, N2607);
or OR4 (N9326, N9323, N2988, N6051, N7441);
buf BUF1 (N9327, N9312);
or OR2 (N9328, N9324, N8060);
not NOT1 (N9329, N9327);
and AND3 (N9330, N9316, N1821, N7016);
buf BUF1 (N9331, N9319);
buf BUF1 (N9332, N9330);
nand NAND2 (N9333, N9328, N4172);
not NOT1 (N9334, N9325);
or OR4 (N9335, N9333, N5246, N7846, N5415);
xor XOR2 (N9336, N9322, N6041);
nor NOR3 (N9337, N9336, N3050, N7574);
not NOT1 (N9338, N9318);
xor XOR2 (N9339, N9326, N479);
buf BUF1 (N9340, N9338);
or OR3 (N9341, N9329, N7346, N7945);
nor NOR3 (N9342, N9341, N3187, N34);
buf BUF1 (N9343, N9332);
not NOT1 (N9344, N9335);
not NOT1 (N9345, N9334);
nor NOR3 (N9346, N9308, N189, N1818);
not NOT1 (N9347, N9343);
buf BUF1 (N9348, N9344);
or OR4 (N9349, N9342, N6215, N8669, N7984);
nor NOR3 (N9350, N9348, N5107, N1939);
buf BUF1 (N9351, N9345);
or OR3 (N9352, N9331, N2343, N982);
not NOT1 (N9353, N9352);
and AND2 (N9354, N9353, N8466);
and AND4 (N9355, N9347, N376, N1659, N1270);
nor NOR3 (N9356, N9349, N933, N9102);
xor XOR2 (N9357, N9355, N6483);
not NOT1 (N9358, N9337);
or OR2 (N9359, N9350, N3383);
not NOT1 (N9360, N9346);
and AND3 (N9361, N9357, N3558, N2364);
nand NAND4 (N9362, N9360, N3171, N5829, N4063);
and AND2 (N9363, N9356, N3320);
and AND2 (N9364, N9363, N8053);
or OR2 (N9365, N9364, N1077);
and AND4 (N9366, N9358, N7970, N3720, N7201);
and AND4 (N9367, N9259, N6388, N176, N4509);
not NOT1 (N9368, N9351);
or OR4 (N9369, N9361, N1465, N2383, N9020);
nor NOR4 (N9370, N9367, N3285, N2749, N5306);
or OR2 (N9371, N9366, N6641);
and AND3 (N9372, N9369, N8193, N490);
nand NAND3 (N9373, N9339, N8028, N3140);
nor NOR4 (N9374, N9372, N9132, N52, N4663);
and AND3 (N9375, N9371, N5357, N8631);
nand NAND4 (N9376, N9354, N5002, N7109, N1317);
or OR4 (N9377, N9362, N2556, N3810, N3642);
nor NOR3 (N9378, N9368, N1456, N4452);
xor XOR2 (N9379, N9373, N4520);
or OR3 (N9380, N9376, N6571, N2666);
buf BUF1 (N9381, N9380);
or OR3 (N9382, N9340, N7618, N3973);
or OR3 (N9383, N9359, N1764, N4694);
not NOT1 (N9384, N9381);
nor NOR3 (N9385, N9377, N4438, N1610);
nor NOR2 (N9386, N9385, N2829);
not NOT1 (N9387, N9379);
nor NOR2 (N9388, N9384, N4912);
or OR2 (N9389, N9387, N3743);
nand NAND3 (N9390, N9378, N370, N3106);
not NOT1 (N9391, N9374);
and AND3 (N9392, N9382, N1417, N5923);
xor XOR2 (N9393, N9391, N9138);
or OR3 (N9394, N9388, N9249, N5436);
and AND2 (N9395, N9390, N1400);
and AND3 (N9396, N9386, N4464, N7145);
nand NAND4 (N9397, N9392, N7541, N1923, N9203);
or OR3 (N9398, N9389, N1255, N5216);
or OR4 (N9399, N9370, N8148, N2440, N9012);
and AND2 (N9400, N9398, N5396);
nor NOR4 (N9401, N9399, N8531, N6423, N4595);
nor NOR4 (N9402, N9395, N8021, N8295, N2838);
nor NOR4 (N9403, N9383, N5668, N4895, N811);
buf BUF1 (N9404, N9400);
buf BUF1 (N9405, N9397);
xor XOR2 (N9406, N9402, N5057);
and AND4 (N9407, N9405, N3784, N9174, N8400);
not NOT1 (N9408, N9404);
not NOT1 (N9409, N9394);
nor NOR4 (N9410, N9365, N1320, N2009, N2541);
nor NOR2 (N9411, N9393, N8033);
buf BUF1 (N9412, N9408);
xor XOR2 (N9413, N9375, N783);
xor XOR2 (N9414, N9403, N2785);
xor XOR2 (N9415, N9407, N7907);
nand NAND3 (N9416, N9411, N1189, N5139);
nand NAND2 (N9417, N9415, N946);
nand NAND2 (N9418, N9412, N2527);
xor XOR2 (N9419, N9406, N6167);
or OR2 (N9420, N9414, N8697);
buf BUF1 (N9421, N9413);
or OR4 (N9422, N9409, N5856, N6891, N77);
buf BUF1 (N9423, N9419);
nand NAND3 (N9424, N9417, N5436, N8628);
not NOT1 (N9425, N9420);
not NOT1 (N9426, N9401);
and AND3 (N9427, N9421, N4920, N4247);
or OR2 (N9428, N9424, N8251);
xor XOR2 (N9429, N9410, N3418);
xor XOR2 (N9430, N9396, N5083);
xor XOR2 (N9431, N9418, N764);
and AND2 (N9432, N9416, N1097);
or OR3 (N9433, N9431, N3034, N8704);
not NOT1 (N9434, N9429);
not NOT1 (N9435, N9426);
xor XOR2 (N9436, N9428, N5793);
xor XOR2 (N9437, N9435, N6951);
not NOT1 (N9438, N9432);
not NOT1 (N9439, N9425);
nor NOR4 (N9440, N9423, N3527, N5706, N4459);
not NOT1 (N9441, N9440);
and AND4 (N9442, N9427, N9172, N9167, N6945);
not NOT1 (N9443, N9434);
not NOT1 (N9444, N9441);
xor XOR2 (N9445, N9433, N7557);
or OR3 (N9446, N9430, N3445, N3854);
buf BUF1 (N9447, N9445);
nand NAND2 (N9448, N9442, N6257);
nor NOR4 (N9449, N9422, N742, N5112, N7329);
not NOT1 (N9450, N9436);
buf BUF1 (N9451, N9449);
and AND3 (N9452, N9450, N7801, N9162);
nand NAND2 (N9453, N9451, N3779);
nor NOR2 (N9454, N9453, N5292);
xor XOR2 (N9455, N9454, N4029);
or OR2 (N9456, N9443, N1106);
and AND3 (N9457, N9444, N7604, N8623);
xor XOR2 (N9458, N9439, N8789);
and AND4 (N9459, N9446, N6060, N5519, N2349);
buf BUF1 (N9460, N9452);
xor XOR2 (N9461, N9438, N50);
nand NAND4 (N9462, N9460, N8471, N9021, N5785);
not NOT1 (N9463, N9456);
buf BUF1 (N9464, N9447);
or OR4 (N9465, N9437, N5400, N1725, N6427);
xor XOR2 (N9466, N9448, N750);
not NOT1 (N9467, N9457);
xor XOR2 (N9468, N9458, N8456);
not NOT1 (N9469, N9467);
xor XOR2 (N9470, N9461, N9062);
or OR3 (N9471, N9455, N4530, N6607);
nor NOR2 (N9472, N9468, N5148);
xor XOR2 (N9473, N9462, N7122);
and AND2 (N9474, N9472, N6992);
or OR2 (N9475, N9469, N6755);
and AND3 (N9476, N9470, N6077, N1239);
xor XOR2 (N9477, N9476, N8319);
or OR3 (N9478, N9473, N322, N1658);
nor NOR4 (N9479, N9471, N6679, N7349, N9287);
nand NAND3 (N9480, N9479, N4417, N5524);
or OR4 (N9481, N9477, N1729, N3919, N131);
xor XOR2 (N9482, N9459, N8971);
xor XOR2 (N9483, N9480, N2516);
buf BUF1 (N9484, N9464);
nand NAND2 (N9485, N9466, N7528);
nand NAND3 (N9486, N9481, N6998, N4914);
nor NOR3 (N9487, N9463, N1326, N5201);
nor NOR2 (N9488, N9483, N1136);
buf BUF1 (N9489, N9482);
and AND3 (N9490, N9478, N4999, N1737);
and AND3 (N9491, N9490, N3227, N2021);
and AND3 (N9492, N9485, N2068, N8998);
xor XOR2 (N9493, N9484, N3816);
or OR4 (N9494, N9486, N288, N2188, N6662);
nor NOR4 (N9495, N9474, N1541, N2001, N7617);
and AND3 (N9496, N9489, N6896, N1071);
nor NOR4 (N9497, N9487, N2402, N8319, N5000);
or OR4 (N9498, N9475, N2897, N4783, N7803);
or OR3 (N9499, N9497, N7980, N5576);
or OR3 (N9500, N9488, N7250, N2830);
and AND3 (N9501, N9498, N739, N1711);
xor XOR2 (N9502, N9491, N6734);
nand NAND3 (N9503, N9495, N1820, N5685);
nor NOR4 (N9504, N9499, N125, N6657, N8686);
nor NOR4 (N9505, N9494, N5252, N2507, N7672);
nor NOR3 (N9506, N9505, N3352, N6214);
nor NOR2 (N9507, N9506, N1471);
and AND3 (N9508, N9502, N147, N8796);
nor NOR2 (N9509, N9508, N7308);
nor NOR3 (N9510, N9496, N8219, N4460);
or OR4 (N9511, N9501, N5777, N2408, N1885);
buf BUF1 (N9512, N9507);
and AND4 (N9513, N9465, N3354, N1829, N1001);
nor NOR3 (N9514, N9510, N4215, N6900);
not NOT1 (N9515, N9513);
and AND4 (N9516, N9504, N6697, N1440, N6563);
not NOT1 (N9517, N9500);
not NOT1 (N9518, N9515);
buf BUF1 (N9519, N9503);
xor XOR2 (N9520, N9518, N935);
xor XOR2 (N9521, N9493, N7477);
xor XOR2 (N9522, N9512, N9132);
or OR4 (N9523, N9517, N7078, N6270, N4898);
not NOT1 (N9524, N9516);
xor XOR2 (N9525, N9509, N5814);
nor NOR3 (N9526, N9525, N2101, N8930);
nand NAND4 (N9527, N9511, N5994, N957, N6800);
and AND3 (N9528, N9521, N5297, N3587);
or OR2 (N9529, N9492, N4799);
or OR3 (N9530, N9528, N7906, N361);
nor NOR4 (N9531, N9519, N8046, N8711, N1863);
xor XOR2 (N9532, N9514, N2849);
xor XOR2 (N9533, N9530, N4519);
or OR3 (N9534, N9520, N8412, N5431);
xor XOR2 (N9535, N9522, N5330);
xor XOR2 (N9536, N9534, N4537);
nand NAND3 (N9537, N9524, N9326, N8236);
buf BUF1 (N9538, N9527);
buf BUF1 (N9539, N9523);
nand NAND3 (N9540, N9536, N5947, N102);
nand NAND4 (N9541, N9535, N3168, N9365, N7914);
or OR3 (N9542, N9540, N171, N5655);
and AND2 (N9543, N9538, N500);
nor NOR4 (N9544, N9541, N2850, N6854, N5106);
buf BUF1 (N9545, N9543);
nor NOR3 (N9546, N9531, N8209, N9078);
not NOT1 (N9547, N9542);
buf BUF1 (N9548, N9532);
nor NOR4 (N9549, N9544, N4994, N3384, N1151);
and AND3 (N9550, N9526, N8957, N7466);
nand NAND3 (N9551, N9547, N1729, N7611);
buf BUF1 (N9552, N9533);
nand NAND3 (N9553, N9550, N9217, N6069);
and AND4 (N9554, N9549, N2657, N2571, N6757);
nor NOR2 (N9555, N9546, N2218);
and AND4 (N9556, N9555, N2131, N4182, N7917);
buf BUF1 (N9557, N9553);
or OR3 (N9558, N9548, N4919, N258);
buf BUF1 (N9559, N9545);
nor NOR4 (N9560, N9539, N6615, N1437, N536);
and AND2 (N9561, N9537, N1679);
and AND3 (N9562, N9554, N8444, N2749);
and AND2 (N9563, N9561, N5202);
buf BUF1 (N9564, N9556);
not NOT1 (N9565, N9557);
not NOT1 (N9566, N9560);
and AND2 (N9567, N9566, N1791);
buf BUF1 (N9568, N9563);
nand NAND4 (N9569, N9529, N2361, N210, N3908);
nand NAND2 (N9570, N9568, N7832);
not NOT1 (N9571, N9551);
nand NAND4 (N9572, N9571, N7762, N4164, N4468);
or OR4 (N9573, N9558, N9256, N6259, N6557);
nand NAND4 (N9574, N9569, N7025, N8157, N4962);
buf BUF1 (N9575, N9564);
and AND2 (N9576, N9572, N8651);
and AND4 (N9577, N9562, N1628, N1285, N7605);
nand NAND4 (N9578, N9574, N1739, N3566, N4558);
not NOT1 (N9579, N9559);
buf BUF1 (N9580, N9578);
xor XOR2 (N9581, N9576, N9369);
or OR4 (N9582, N9552, N6986, N1117, N9092);
and AND2 (N9583, N9565, N2673);
and AND4 (N9584, N9579, N4020, N1151, N8667);
nand NAND3 (N9585, N9567, N550, N3068);
nor NOR3 (N9586, N9570, N7284, N1553);
and AND4 (N9587, N9581, N6104, N3488, N7814);
not NOT1 (N9588, N9582);
and AND2 (N9589, N9588, N2096);
nand NAND4 (N9590, N9587, N7567, N1593, N118);
buf BUF1 (N9591, N9580);
nor NOR3 (N9592, N9575, N3847, N9588);
not NOT1 (N9593, N9586);
not NOT1 (N9594, N9591);
buf BUF1 (N9595, N9590);
nand NAND2 (N9596, N9594, N7567);
nand NAND3 (N9597, N9583, N6160, N3448);
nor NOR2 (N9598, N9589, N4209);
and AND2 (N9599, N9598, N8886);
not NOT1 (N9600, N9597);
and AND2 (N9601, N9595, N5902);
nor NOR4 (N9602, N9593, N2698, N8411, N8680);
not NOT1 (N9603, N9602);
buf BUF1 (N9604, N9585);
xor XOR2 (N9605, N9601, N2327);
nand NAND3 (N9606, N9584, N7508, N2015);
nor NOR2 (N9607, N9577, N1584);
xor XOR2 (N9608, N9599, N5317);
not NOT1 (N9609, N9607);
xor XOR2 (N9610, N9609, N4873);
buf BUF1 (N9611, N9592);
buf BUF1 (N9612, N9596);
xor XOR2 (N9613, N9610, N6433);
and AND3 (N9614, N9604, N5703, N4005);
nor NOR4 (N9615, N9600, N5161, N9292, N7565);
and AND3 (N9616, N9606, N1186, N2494);
buf BUF1 (N9617, N9614);
nand NAND3 (N9618, N9612, N4418, N8723);
not NOT1 (N9619, N9608);
and AND2 (N9620, N9616, N8633);
or OR2 (N9621, N9611, N5439);
buf BUF1 (N9622, N9613);
or OR2 (N9623, N9573, N6901);
not NOT1 (N9624, N9615);
nand NAND2 (N9625, N9620, N652);
buf BUF1 (N9626, N9619);
not NOT1 (N9627, N9622);
nand NAND3 (N9628, N9618, N6951, N7248);
nor NOR3 (N9629, N9621, N1841, N2090);
and AND4 (N9630, N9626, N3617, N8499, N3981);
nand NAND3 (N9631, N9623, N6910, N7157);
or OR3 (N9632, N9627, N762, N1332);
nand NAND4 (N9633, N9631, N8183, N7289, N7893);
nand NAND3 (N9634, N9628, N9203, N6408);
xor XOR2 (N9635, N9624, N493);
buf BUF1 (N9636, N9625);
or OR4 (N9637, N9603, N8379, N9394, N1939);
nand NAND3 (N9638, N9634, N9539, N4281);
nand NAND2 (N9639, N9635, N8917);
and AND3 (N9640, N9630, N1775, N6012);
buf BUF1 (N9641, N9637);
nor NOR3 (N9642, N9639, N4485, N8400);
xor XOR2 (N9643, N9629, N2290);
xor XOR2 (N9644, N9636, N2809);
and AND4 (N9645, N9605, N6703, N8576, N5825);
nand NAND2 (N9646, N9641, N4088);
nand NAND2 (N9647, N9644, N2063);
nor NOR2 (N9648, N9638, N8495);
nand NAND2 (N9649, N9646, N2910);
nand NAND2 (N9650, N9643, N3292);
xor XOR2 (N9651, N9642, N5289);
buf BUF1 (N9652, N9651);
or OR2 (N9653, N9648, N7445);
or OR4 (N9654, N9652, N7043, N7868, N8649);
or OR4 (N9655, N9647, N9632, N9129, N3815);
or OR3 (N9656, N9384, N6008, N7630);
xor XOR2 (N9657, N9650, N8278);
and AND3 (N9658, N9655, N6503, N3807);
buf BUF1 (N9659, N9654);
xor XOR2 (N9660, N9653, N6566);
not NOT1 (N9661, N9645);
or OR3 (N9662, N9640, N9550, N7710);
or OR2 (N9663, N9656, N7088);
xor XOR2 (N9664, N9663, N138);
and AND2 (N9665, N9664, N204);
not NOT1 (N9666, N9662);
or OR2 (N9667, N9661, N9605);
and AND2 (N9668, N9659, N4095);
nor NOR3 (N9669, N9617, N901, N9065);
buf BUF1 (N9670, N9657);
and AND4 (N9671, N9658, N3149, N978, N7129);
not NOT1 (N9672, N9669);
or OR3 (N9673, N9671, N1702, N1177);
not NOT1 (N9674, N9660);
nand NAND3 (N9675, N9667, N1691, N1871);
xor XOR2 (N9676, N9674, N6031);
xor XOR2 (N9677, N9673, N5890);
not NOT1 (N9678, N9649);
nor NOR2 (N9679, N9666, N6757);
and AND2 (N9680, N9677, N2959);
xor XOR2 (N9681, N9665, N4464);
nand NAND2 (N9682, N9680, N5556);
xor XOR2 (N9683, N9681, N6492);
buf BUF1 (N9684, N9676);
nor NOR2 (N9685, N9633, N5185);
nor NOR3 (N9686, N9678, N8450, N2237);
nand NAND3 (N9687, N9672, N4109, N6802);
xor XOR2 (N9688, N9686, N91);
buf BUF1 (N9689, N9679);
nand NAND3 (N9690, N9687, N5208, N1539);
nor NOR4 (N9691, N9685, N4402, N4738, N1259);
not NOT1 (N9692, N9675);
buf BUF1 (N9693, N9684);
xor XOR2 (N9694, N9688, N3482);
not NOT1 (N9695, N9683);
nand NAND3 (N9696, N9689, N459, N8058);
xor XOR2 (N9697, N9691, N1425);
and AND3 (N9698, N9670, N4775, N1817);
and AND4 (N9699, N9697, N353, N4339, N4444);
not NOT1 (N9700, N9695);
and AND2 (N9701, N9668, N6194);
nor NOR2 (N9702, N9693, N8228);
or OR3 (N9703, N9698, N5307, N1999);
buf BUF1 (N9704, N9682);
nand NAND4 (N9705, N9699, N4071, N3761, N9095);
or OR4 (N9706, N9701, N5211, N7784, N9274);
xor XOR2 (N9707, N9706, N9528);
or OR4 (N9708, N9705, N6470, N3665, N2262);
nand NAND4 (N9709, N9694, N8371, N5341, N2351);
and AND3 (N9710, N9707, N8604, N5533);
xor XOR2 (N9711, N9703, N9116);
and AND4 (N9712, N9711, N985, N2673, N1430);
buf BUF1 (N9713, N9710);
nand NAND2 (N9714, N9696, N5268);
nor NOR4 (N9715, N9712, N1484, N9333, N6665);
and AND4 (N9716, N9708, N1224, N7817, N7572);
or OR2 (N9717, N9690, N5189);
xor XOR2 (N9718, N9704, N9572);
or OR2 (N9719, N9702, N2097);
nand NAND2 (N9720, N9715, N115);
nand NAND4 (N9721, N9709, N8683, N3124, N1256);
buf BUF1 (N9722, N9718);
buf BUF1 (N9723, N9716);
xor XOR2 (N9724, N9722, N9372);
xor XOR2 (N9725, N9719, N8292);
or OR4 (N9726, N9724, N5203, N9218, N77);
nand NAND3 (N9727, N9692, N8706, N9444);
buf BUF1 (N9728, N9721);
xor XOR2 (N9729, N9726, N1045);
and AND4 (N9730, N9720, N5139, N575, N5638);
xor XOR2 (N9731, N9729, N8771);
buf BUF1 (N9732, N9731);
not NOT1 (N9733, N9725);
and AND2 (N9734, N9727, N6949);
or OR4 (N9735, N9717, N1656, N1548, N8276);
or OR4 (N9736, N9730, N9135, N1977, N3618);
or OR2 (N9737, N9735, N3532);
nor NOR3 (N9738, N9700, N883, N5903);
xor XOR2 (N9739, N9736, N4553);
buf BUF1 (N9740, N9732);
buf BUF1 (N9741, N9738);
buf BUF1 (N9742, N9733);
and AND3 (N9743, N9723, N4453, N3242);
and AND3 (N9744, N9714, N270, N3904);
not NOT1 (N9745, N9741);
not NOT1 (N9746, N9740);
xor XOR2 (N9747, N9734, N1751);
nand NAND4 (N9748, N9745, N6468, N7902, N9352);
buf BUF1 (N9749, N9742);
xor XOR2 (N9750, N9743, N5329);
or OR3 (N9751, N9749, N3669, N9656);
nor NOR3 (N9752, N9744, N9583, N5394);
nand NAND2 (N9753, N9748, N5755);
nand NAND2 (N9754, N9746, N6014);
and AND3 (N9755, N9747, N9362, N3801);
not NOT1 (N9756, N9753);
or OR3 (N9757, N9756, N9358, N9414);
or OR4 (N9758, N9739, N8678, N8726, N5468);
and AND3 (N9759, N9754, N436, N6269);
and AND2 (N9760, N9757, N8081);
buf BUF1 (N9761, N9758);
and AND3 (N9762, N9728, N3000, N8202);
and AND3 (N9763, N9713, N3262, N2287);
nor NOR4 (N9764, N9752, N9363, N1957, N5579);
buf BUF1 (N9765, N9751);
nor NOR2 (N9766, N9737, N4080);
or OR2 (N9767, N9755, N5576);
nand NAND3 (N9768, N9762, N9245, N991);
buf BUF1 (N9769, N9765);
or OR2 (N9770, N9750, N4474);
buf BUF1 (N9771, N9770);
nor NOR2 (N9772, N9763, N95);
nor NOR2 (N9773, N9771, N6088);
buf BUF1 (N9774, N9768);
nor NOR4 (N9775, N9766, N8743, N1262, N8921);
xor XOR2 (N9776, N9764, N8371);
nor NOR4 (N9777, N9776, N7631, N6252, N7657);
and AND4 (N9778, N9772, N9768, N3027, N2323);
and AND4 (N9779, N9769, N1513, N2663, N7863);
buf BUF1 (N9780, N9779);
xor XOR2 (N9781, N9767, N4875);
nor NOR4 (N9782, N9759, N7767, N7381, N1917);
nand NAND4 (N9783, N9781, N2549, N2840, N6076);
nor NOR2 (N9784, N9778, N1271);
nand NAND3 (N9785, N9774, N4424, N1564);
xor XOR2 (N9786, N9760, N4155);
nor NOR2 (N9787, N9783, N5637);
and AND3 (N9788, N9782, N1324, N6141);
and AND4 (N9789, N9773, N3658, N1500, N4799);
xor XOR2 (N9790, N9775, N9067);
nand NAND2 (N9791, N9786, N580);
buf BUF1 (N9792, N9788);
nand NAND4 (N9793, N9761, N7844, N5795, N4969);
buf BUF1 (N9794, N9785);
buf BUF1 (N9795, N9784);
buf BUF1 (N9796, N9794);
xor XOR2 (N9797, N9793, N9021);
or OR2 (N9798, N9797, N5678);
not NOT1 (N9799, N9787);
not NOT1 (N9800, N9780);
and AND4 (N9801, N9789, N7354, N3809, N6253);
nor NOR2 (N9802, N9791, N7724);
nand NAND3 (N9803, N9795, N9053, N6460);
nor NOR2 (N9804, N9800, N9071);
and AND4 (N9805, N9798, N5268, N2398, N7047);
buf BUF1 (N9806, N9777);
or OR2 (N9807, N9790, N7568);
and AND2 (N9808, N9801, N1099);
not NOT1 (N9809, N9792);
or OR3 (N9810, N9796, N9749, N1132);
and AND2 (N9811, N9803, N7104);
or OR3 (N9812, N9804, N5648, N9591);
nor NOR2 (N9813, N9806, N6267);
and AND4 (N9814, N9808, N3260, N2631, N319);
or OR3 (N9815, N9813, N1725, N2341);
xor XOR2 (N9816, N9814, N9483);
xor XOR2 (N9817, N9809, N2323);
or OR4 (N9818, N9815, N9771, N7647, N5757);
or OR2 (N9819, N9816, N985);
or OR3 (N9820, N9799, N1445, N5597);
nor NOR4 (N9821, N9818, N2283, N5947, N8316);
and AND3 (N9822, N9811, N3061, N5012);
not NOT1 (N9823, N9810);
nor NOR3 (N9824, N9821, N721, N5898);
and AND3 (N9825, N9823, N5133, N3834);
and AND4 (N9826, N9802, N1693, N3834, N1742);
buf BUF1 (N9827, N9805);
nand NAND3 (N9828, N9826, N4128, N1090);
or OR2 (N9829, N9820, N1223);
and AND4 (N9830, N9817, N2939, N1201, N1028);
nand NAND3 (N9831, N9807, N3210, N267);
xor XOR2 (N9832, N9827, N4624);
and AND4 (N9833, N9829, N782, N6331, N2980);
buf BUF1 (N9834, N9828);
or OR2 (N9835, N9824, N7321);
nand NAND2 (N9836, N9833, N4407);
nor NOR2 (N9837, N9812, N391);
or OR2 (N9838, N9819, N6746);
not NOT1 (N9839, N9825);
nor NOR2 (N9840, N9835, N9612);
or OR2 (N9841, N9834, N206);
buf BUF1 (N9842, N9832);
buf BUF1 (N9843, N9837);
not NOT1 (N9844, N9830);
xor XOR2 (N9845, N9844, N8935);
and AND4 (N9846, N9838, N4021, N3062, N839);
buf BUF1 (N9847, N9822);
or OR3 (N9848, N9842, N5278, N6847);
or OR2 (N9849, N9848, N506);
buf BUF1 (N9850, N9841);
and AND4 (N9851, N9847, N1482, N5574, N117);
and AND3 (N9852, N9839, N3919, N4440);
buf BUF1 (N9853, N9840);
xor XOR2 (N9854, N9845, N3171);
or OR2 (N9855, N9846, N7915);
buf BUF1 (N9856, N9855);
not NOT1 (N9857, N9843);
nand NAND2 (N9858, N9851, N4954);
nor NOR4 (N9859, N9836, N4791, N6358, N7078);
or OR3 (N9860, N9856, N8799, N719);
or OR2 (N9861, N9859, N5911);
not NOT1 (N9862, N9831);
nand NAND2 (N9863, N9860, N2269);
nand NAND4 (N9864, N9858, N7000, N4304, N6781);
xor XOR2 (N9865, N9853, N70);
or OR2 (N9866, N9854, N2009);
and AND2 (N9867, N9849, N1997);
nand NAND2 (N9868, N9866, N7733);
nand NAND2 (N9869, N9852, N6427);
xor XOR2 (N9870, N9857, N4371);
nand NAND4 (N9871, N9862, N8205, N6844, N7756);
xor XOR2 (N9872, N9850, N5862);
or OR2 (N9873, N9865, N1443);
not NOT1 (N9874, N9864);
not NOT1 (N9875, N9869);
xor XOR2 (N9876, N9867, N444);
buf BUF1 (N9877, N9876);
buf BUF1 (N9878, N9861);
nand NAND4 (N9879, N9875, N3558, N7309, N7018);
and AND3 (N9880, N9873, N2280, N5037);
or OR4 (N9881, N9863, N9853, N8203, N2807);
and AND3 (N9882, N9872, N8698, N8650);
not NOT1 (N9883, N9882);
nand NAND2 (N9884, N9870, N7569);
nand NAND2 (N9885, N9883, N287);
nor NOR4 (N9886, N9871, N8744, N125, N5263);
nand NAND4 (N9887, N9868, N7681, N5338, N8693);
nand NAND4 (N9888, N9886, N2990, N6623, N694);
nor NOR4 (N9889, N9885, N5398, N1475, N2256);
buf BUF1 (N9890, N9887);
or OR3 (N9891, N9888, N414, N7979);
nor NOR4 (N9892, N9874, N3883, N723, N885);
or OR4 (N9893, N9879, N2890, N6451, N9280);
nor NOR4 (N9894, N9892, N656, N8607, N5459);
buf BUF1 (N9895, N9884);
or OR3 (N9896, N9890, N7705, N2348);
xor XOR2 (N9897, N9895, N3692);
not NOT1 (N9898, N9896);
nand NAND2 (N9899, N9881, N327);
or OR3 (N9900, N9893, N4126, N4075);
or OR4 (N9901, N9891, N9264, N3289, N6334);
nand NAND3 (N9902, N9880, N940, N932);
buf BUF1 (N9903, N9877);
not NOT1 (N9904, N9900);
nor NOR4 (N9905, N9889, N9338, N3265, N1539);
nand NAND4 (N9906, N9903, N8393, N9517, N371);
and AND4 (N9907, N9901, N2980, N2790, N4799);
nor NOR2 (N9908, N9905, N5737);
nand NAND4 (N9909, N9906, N7837, N3147, N2314);
nor NOR3 (N9910, N9878, N4395, N9506);
or OR4 (N9911, N9898, N6675, N4654, N6349);
or OR2 (N9912, N9908, N1071);
buf BUF1 (N9913, N9911);
or OR4 (N9914, N9894, N6473, N2457, N149);
and AND4 (N9915, N9910, N8372, N9037, N1296);
not NOT1 (N9916, N9914);
or OR2 (N9917, N9904, N4294);
and AND3 (N9918, N9907, N34, N6196);
buf BUF1 (N9919, N9902);
not NOT1 (N9920, N9899);
nor NOR2 (N9921, N9915, N8399);
xor XOR2 (N9922, N9909, N8774);
not NOT1 (N9923, N9921);
nand NAND4 (N9924, N9919, N7422, N7327, N2035);
nor NOR3 (N9925, N9923, N3350, N6487);
nand NAND4 (N9926, N9918, N9127, N3166, N6456);
nor NOR2 (N9927, N9920, N9160);
xor XOR2 (N9928, N9897, N982);
nand NAND3 (N9929, N9917, N1701, N7174);
not NOT1 (N9930, N9912);
xor XOR2 (N9931, N9930, N6806);
or OR3 (N9932, N9922, N5735, N7402);
and AND3 (N9933, N9927, N5593, N3711);
buf BUF1 (N9934, N9931);
buf BUF1 (N9935, N9925);
and AND3 (N9936, N9929, N4435, N9513);
or OR4 (N9937, N9913, N3470, N2244, N5146);
not NOT1 (N9938, N9936);
nor NOR2 (N9939, N9935, N7753);
not NOT1 (N9940, N9916);
or OR2 (N9941, N9934, N2389);
or OR2 (N9942, N9928, N6420);
buf BUF1 (N9943, N9937);
buf BUF1 (N9944, N9932);
or OR2 (N9945, N9926, N7800);
not NOT1 (N9946, N9933);
nand NAND2 (N9947, N9943, N3570);
nor NOR2 (N9948, N9945, N7582);
not NOT1 (N9949, N9948);
buf BUF1 (N9950, N9944);
not NOT1 (N9951, N9949);
nand NAND3 (N9952, N9938, N4991, N1382);
or OR4 (N9953, N9952, N9924, N946, N2232);
or OR2 (N9954, N5854, N1391);
nor NOR3 (N9955, N9939, N2984, N2114);
not NOT1 (N9956, N9954);
and AND4 (N9957, N9946, N5519, N6798, N4124);
and AND3 (N9958, N9942, N893, N223);
nand NAND4 (N9959, N9953, N6730, N5958, N6224);
nor NOR3 (N9960, N9955, N5743, N8474);
nor NOR4 (N9961, N9951, N8619, N8860, N3029);
xor XOR2 (N9962, N9961, N7558);
not NOT1 (N9963, N9947);
not NOT1 (N9964, N9958);
xor XOR2 (N9965, N9956, N1143);
or OR4 (N9966, N9965, N2584, N6595, N9040);
xor XOR2 (N9967, N9957, N5504);
buf BUF1 (N9968, N9960);
buf BUF1 (N9969, N9941);
or OR4 (N9970, N9962, N77, N7994, N1112);
xor XOR2 (N9971, N9968, N7538);
nor NOR4 (N9972, N9967, N816, N906, N482);
and AND3 (N9973, N9971, N1210, N6922);
xor XOR2 (N9974, N9972, N3871);
and AND4 (N9975, N9959, N514, N5574, N4319);
and AND3 (N9976, N9966, N106, N1790);
not NOT1 (N9977, N9969);
buf BUF1 (N9978, N9977);
xor XOR2 (N9979, N9978, N9561);
nor NOR3 (N9980, N9940, N2122, N1323);
not NOT1 (N9981, N9979);
or OR3 (N9982, N9970, N9525, N5580);
or OR4 (N9983, N9964, N7486, N1426, N6181);
buf BUF1 (N9984, N9975);
nor NOR4 (N9985, N9973, N6290, N7618, N335);
buf BUF1 (N9986, N9963);
buf BUF1 (N9987, N9974);
not NOT1 (N9988, N9950);
not NOT1 (N9989, N9981);
or OR4 (N9990, N9983, N9796, N566, N8803);
nand NAND4 (N9991, N9985, N1802, N5157, N7935);
and AND3 (N9992, N9986, N4607, N1444);
nor NOR3 (N9993, N9991, N937, N4037);
nor NOR4 (N9994, N9993, N8212, N9530, N1237);
not NOT1 (N9995, N9992);
or OR2 (N9996, N9988, N78);
not NOT1 (N9997, N9987);
nor NOR4 (N9998, N9984, N967, N6712, N7675);
nor NOR4 (N9999, N9998, N7807, N4597, N2139);
and AND3 (N10000, N9982, N8125, N2182);
xor XOR2 (N10001, N9990, N6464);
buf BUF1 (N10002, N9996);
nor NOR2 (N10003, N9999, N427);
not NOT1 (N10004, N10002);
xor XOR2 (N10005, N10004, N4294);
and AND2 (N10006, N9989, N8719);
buf BUF1 (N10007, N10006);
not NOT1 (N10008, N9976);
not NOT1 (N10009, N9994);
nor NOR2 (N10010, N10001, N6805);
not NOT1 (N10011, N9995);
nor NOR2 (N10012, N10009, N3978);
buf BUF1 (N10013, N10000);
nand NAND2 (N10014, N10013, N5373);
or OR4 (N10015, N10010, N3581, N3393, N2956);
or OR4 (N10016, N10015, N4614, N2622, N3608);
and AND3 (N10017, N9980, N6014, N5979);
nor NOR4 (N10018, N10007, N5832, N9463, N7745);
nand NAND2 (N10019, N9997, N8493);
or OR3 (N10020, N10016, N164, N1089);
not NOT1 (N10021, N10008);
not NOT1 (N10022, N10003);
not NOT1 (N10023, N10022);
and AND3 (N10024, N10011, N3471, N6221);
xor XOR2 (N10025, N10017, N4965);
xor XOR2 (N10026, N10020, N7788);
xor XOR2 (N10027, N10005, N6354);
buf BUF1 (N10028, N10023);
and AND3 (N10029, N10021, N5236, N2951);
nor NOR3 (N10030, N10019, N8836, N3081);
nor NOR4 (N10031, N10030, N5886, N2772, N6899);
or OR3 (N10032, N10027, N4853, N5867);
nor NOR4 (N10033, N10014, N5114, N8169, N7650);
and AND2 (N10034, N10028, N1119);
not NOT1 (N10035, N10012);
xor XOR2 (N10036, N10032, N3834);
nor NOR2 (N10037, N10034, N5439);
buf BUF1 (N10038, N10029);
or OR2 (N10039, N10026, N6739);
or OR4 (N10040, N10038, N6746, N1429, N5542);
or OR2 (N10041, N10033, N6041);
nand NAND4 (N10042, N10018, N7728, N5757, N850);
buf BUF1 (N10043, N10041);
or OR4 (N10044, N10024, N769, N5049, N97);
and AND4 (N10045, N10025, N7336, N2292, N4718);
nor NOR3 (N10046, N10037, N8708, N7716);
buf BUF1 (N10047, N10036);
and AND3 (N10048, N10042, N2434, N5335);
not NOT1 (N10049, N10043);
not NOT1 (N10050, N10035);
nand NAND4 (N10051, N10045, N5518, N2535, N7366);
nand NAND2 (N10052, N10031, N3324);
and AND3 (N10053, N10048, N1196, N985);
nand NAND4 (N10054, N10053, N9146, N8965, N4352);
and AND4 (N10055, N10050, N7888, N9525, N5746);
buf BUF1 (N10056, N10047);
and AND4 (N10057, N10046, N9365, N344, N5549);
nand NAND4 (N10058, N10055, N2622, N6268, N380);
xor XOR2 (N10059, N10058, N1002);
nand NAND2 (N10060, N10044, N9603);
and AND3 (N10061, N10052, N1228, N6199);
xor XOR2 (N10062, N10051, N3235);
nand NAND3 (N10063, N10057, N4601, N5102);
xor XOR2 (N10064, N10061, N3027);
buf BUF1 (N10065, N10064);
buf BUF1 (N10066, N10039);
and AND3 (N10067, N10054, N716, N5779);
xor XOR2 (N10068, N10067, N1304);
nand NAND3 (N10069, N10049, N7732, N5106);
not NOT1 (N10070, N10068);
and AND4 (N10071, N10040, N1502, N5466, N6663);
and AND3 (N10072, N10066, N9921, N2001);
or OR3 (N10073, N10065, N8016, N6353);
nand NAND3 (N10074, N10056, N6674, N760);
or OR3 (N10075, N10060, N3281, N5334);
nand NAND3 (N10076, N10062, N8849, N9716);
nor NOR2 (N10077, N10073, N1414);
or OR2 (N10078, N10077, N3711);
xor XOR2 (N10079, N10074, N7712);
nor NOR2 (N10080, N10063, N4273);
not NOT1 (N10081, N10071);
nor NOR2 (N10082, N10081, N3852);
xor XOR2 (N10083, N10070, N3169);
nor NOR3 (N10084, N10072, N170, N5406);
xor XOR2 (N10085, N10082, N280);
xor XOR2 (N10086, N10075, N486);
xor XOR2 (N10087, N10059, N3475);
not NOT1 (N10088, N10069);
nor NOR2 (N10089, N10079, N8096);
buf BUF1 (N10090, N10076);
and AND4 (N10091, N10088, N1045, N1378, N6994);
xor XOR2 (N10092, N10086, N678);
and AND4 (N10093, N10092, N9579, N8340, N6434);
buf BUF1 (N10094, N10087);
buf BUF1 (N10095, N10093);
buf BUF1 (N10096, N10084);
not NOT1 (N10097, N10078);
or OR4 (N10098, N10094, N5808, N5470, N184);
and AND2 (N10099, N10095, N7600);
buf BUF1 (N10100, N10099);
nor NOR3 (N10101, N10090, N1968, N9056);
and AND3 (N10102, N10097, N5140, N4123);
nand NAND3 (N10103, N10102, N3652, N8527);
buf BUF1 (N10104, N10091);
nor NOR2 (N10105, N10101, N8181);
nor NOR3 (N10106, N10096, N9845, N4002);
xor XOR2 (N10107, N10104, N2912);
and AND3 (N10108, N10103, N7394, N9896);
nor NOR4 (N10109, N10108, N1942, N4021, N5473);
not NOT1 (N10110, N10107);
or OR3 (N10111, N10085, N689, N4236);
nor NOR2 (N10112, N10106, N1413);
or OR4 (N10113, N10083, N6901, N812, N5682);
and AND4 (N10114, N10111, N8313, N3313, N7172);
and AND4 (N10115, N10105, N3924, N2532, N1359);
buf BUF1 (N10116, N10080);
not NOT1 (N10117, N10115);
nand NAND4 (N10118, N10113, N6576, N3753, N3646);
nand NAND3 (N10119, N10100, N4223, N5945);
nor NOR4 (N10120, N10109, N3427, N79, N2577);
nand NAND2 (N10121, N10118, N10035);
nand NAND3 (N10122, N10120, N6999, N6753);
or OR3 (N10123, N10089, N1104, N8145);
and AND4 (N10124, N10098, N8910, N5300, N3362);
not NOT1 (N10125, N10124);
xor XOR2 (N10126, N10125, N9371);
buf BUF1 (N10127, N10112);
xor XOR2 (N10128, N10126, N9879);
nand NAND4 (N10129, N10127, N10074, N6267, N2398);
and AND3 (N10130, N10129, N1681, N221);
nand NAND2 (N10131, N10123, N8400);
xor XOR2 (N10132, N10121, N3641);
nand NAND2 (N10133, N10110, N2815);
xor XOR2 (N10134, N10119, N7793);
buf BUF1 (N10135, N10134);
or OR4 (N10136, N10132, N5478, N6025, N3300);
and AND3 (N10137, N10135, N9049, N6239);
nand NAND4 (N10138, N10128, N7608, N5003, N2098);
and AND4 (N10139, N10122, N6211, N4120, N4308);
or OR3 (N10140, N10138, N5781, N3631);
buf BUF1 (N10141, N10114);
xor XOR2 (N10142, N10141, N2096);
and AND2 (N10143, N10136, N9240);
not NOT1 (N10144, N10117);
or OR3 (N10145, N10140, N9220, N5083);
xor XOR2 (N10146, N10144, N8113);
nor NOR2 (N10147, N10130, N465);
nand NAND3 (N10148, N10147, N640, N4025);
nand NAND2 (N10149, N10143, N8299);
nor NOR4 (N10150, N10148, N5078, N1310, N2412);
or OR3 (N10151, N10145, N2298, N5703);
not NOT1 (N10152, N10149);
xor XOR2 (N10153, N10139, N6555);
xor XOR2 (N10154, N10142, N372);
nand NAND3 (N10155, N10133, N4644, N7088);
or OR2 (N10156, N10152, N6485);
xor XOR2 (N10157, N10154, N1575);
or OR3 (N10158, N10150, N5053, N2789);
nor NOR4 (N10159, N10158, N2724, N1276, N6232);
not NOT1 (N10160, N10157);
not NOT1 (N10161, N10146);
buf BUF1 (N10162, N10160);
nor NOR4 (N10163, N10116, N2199, N9943, N7765);
not NOT1 (N10164, N10159);
or OR3 (N10165, N10161, N2989, N1059);
nor NOR4 (N10166, N10155, N7901, N8948, N1197);
or OR2 (N10167, N10156, N2750);
buf BUF1 (N10168, N10164);
or OR4 (N10169, N10167, N6541, N8642, N4436);
nand NAND3 (N10170, N10151, N2612, N2743);
nand NAND3 (N10171, N10153, N3302, N2220);
xor XOR2 (N10172, N10163, N8849);
nand NAND2 (N10173, N10165, N6179);
or OR4 (N10174, N10168, N158, N9802, N5599);
nand NAND2 (N10175, N10172, N1433);
nand NAND2 (N10176, N10169, N4120);
nand NAND2 (N10177, N10170, N7228);
nor NOR3 (N10178, N10162, N3752, N1601);
nand NAND3 (N10179, N10137, N713, N3654);
nand NAND2 (N10180, N10166, N606);
not NOT1 (N10181, N10131);
nand NAND2 (N10182, N10171, N6770);
or OR2 (N10183, N10174, N1341);
xor XOR2 (N10184, N10182, N2874);
buf BUF1 (N10185, N10184);
nand NAND3 (N10186, N10177, N9092, N4490);
not NOT1 (N10187, N10176);
and AND3 (N10188, N10179, N126, N7562);
xor XOR2 (N10189, N10186, N1348);
not NOT1 (N10190, N10173);
nand NAND2 (N10191, N10175, N8234);
and AND3 (N10192, N10181, N5682, N3734);
nand NAND4 (N10193, N10189, N6742, N2826, N1607);
nand NAND3 (N10194, N10188, N7489, N4076);
not NOT1 (N10195, N10191);
and AND3 (N10196, N10192, N2104, N221);
nor NOR2 (N10197, N10187, N6898);
nor NOR3 (N10198, N10180, N292, N3717);
buf BUF1 (N10199, N10183);
xor XOR2 (N10200, N10198, N6203);
buf BUF1 (N10201, N10178);
nor NOR3 (N10202, N10193, N6973, N8682);
xor XOR2 (N10203, N10202, N1864);
and AND2 (N10204, N10190, N5466);
buf BUF1 (N10205, N10185);
and AND3 (N10206, N10196, N9244, N8670);
buf BUF1 (N10207, N10197);
nand NAND2 (N10208, N10205, N9207);
not NOT1 (N10209, N10200);
xor XOR2 (N10210, N10194, N4701);
buf BUF1 (N10211, N10203);
buf BUF1 (N10212, N10204);
nand NAND3 (N10213, N10207, N3306, N8471);
or OR4 (N10214, N10213, N6722, N825, N2374);
or OR3 (N10215, N10212, N6489, N1278);
xor XOR2 (N10216, N10211, N3002);
xor XOR2 (N10217, N10206, N4818);
buf BUF1 (N10218, N10195);
nand NAND3 (N10219, N10215, N4691, N490);
buf BUF1 (N10220, N10209);
xor XOR2 (N10221, N10199, N3619);
or OR2 (N10222, N10210, N3398);
not NOT1 (N10223, N10221);
not NOT1 (N10224, N10208);
or OR4 (N10225, N10218, N1375, N1178, N7851);
and AND3 (N10226, N10216, N103, N5828);
nand NAND2 (N10227, N10224, N8701);
and AND3 (N10228, N10223, N2240, N6228);
nand NAND3 (N10229, N10222, N7688, N1172);
or OR3 (N10230, N10227, N4864, N6298);
nor NOR2 (N10231, N10219, N6266);
nor NOR3 (N10232, N10201, N755, N1275);
nor NOR2 (N10233, N10230, N1222);
buf BUF1 (N10234, N10217);
buf BUF1 (N10235, N10234);
and AND4 (N10236, N10226, N5779, N10055, N9751);
nor NOR4 (N10237, N10231, N4936, N9861, N3057);
not NOT1 (N10238, N10233);
nor NOR4 (N10239, N10232, N6263, N1521, N8677);
not NOT1 (N10240, N10228);
nor NOR4 (N10241, N10225, N3755, N1685, N53);
nor NOR2 (N10242, N10241, N4155);
nor NOR4 (N10243, N10220, N6303, N3351, N5310);
or OR2 (N10244, N10238, N7549);
or OR2 (N10245, N10229, N9241);
buf BUF1 (N10246, N10244);
nand NAND2 (N10247, N10242, N359);
and AND3 (N10248, N10237, N4634, N7776);
not NOT1 (N10249, N10239);
buf BUF1 (N10250, N10240);
nand NAND4 (N10251, N10249, N4083, N9454, N3264);
not NOT1 (N10252, N10243);
or OR4 (N10253, N10252, N5721, N7166, N1837);
or OR3 (N10254, N10248, N5667, N2394);
not NOT1 (N10255, N10253);
buf BUF1 (N10256, N10255);
or OR2 (N10257, N10247, N747);
and AND2 (N10258, N10256, N4004);
xor XOR2 (N10259, N10235, N9204);
nand NAND3 (N10260, N10258, N3857, N4077);
nor NOR3 (N10261, N10251, N7862, N2065);
nor NOR3 (N10262, N10250, N24, N10006);
nor NOR4 (N10263, N10257, N9825, N995, N6438);
nor NOR2 (N10264, N10261, N3436);
buf BUF1 (N10265, N10264);
and AND4 (N10266, N10263, N5381, N7168, N9785);
and AND2 (N10267, N10236, N8832);
not NOT1 (N10268, N10262);
not NOT1 (N10269, N10267);
nand NAND3 (N10270, N10260, N912, N9413);
nor NOR4 (N10271, N10214, N4367, N10017, N3238);
nand NAND4 (N10272, N10268, N8007, N5876, N10156);
xor XOR2 (N10273, N10246, N1253);
nand NAND2 (N10274, N10272, N6035);
and AND3 (N10275, N10245, N2187, N226);
or OR4 (N10276, N10273, N7652, N4424, N4819);
and AND2 (N10277, N10265, N2324);
buf BUF1 (N10278, N10274);
xor XOR2 (N10279, N10275, N3419);
and AND3 (N10280, N10278, N6189, N8421);
nor NOR4 (N10281, N10279, N632, N4527, N1154);
or OR2 (N10282, N10280, N1796);
buf BUF1 (N10283, N10270);
nand NAND3 (N10284, N10269, N1903, N9576);
nand NAND4 (N10285, N10281, N2949, N8163, N3674);
xor XOR2 (N10286, N10282, N916);
and AND4 (N10287, N10276, N9964, N2750, N272);
xor XOR2 (N10288, N10259, N3740);
nor NOR3 (N10289, N10286, N5051, N5505);
nor NOR4 (N10290, N10266, N108, N4939, N1877);
and AND4 (N10291, N10283, N2825, N6035, N3910);
and AND4 (N10292, N10285, N7225, N886, N2389);
nand NAND4 (N10293, N10254, N18, N4824, N7340);
nand NAND2 (N10294, N10292, N5228);
buf BUF1 (N10295, N10293);
and AND3 (N10296, N10289, N5905, N869);
nor NOR2 (N10297, N10291, N1197);
buf BUF1 (N10298, N10290);
nor NOR4 (N10299, N10297, N8526, N5562, N7169);
or OR3 (N10300, N10284, N2527, N4534);
xor XOR2 (N10301, N10287, N6042);
not NOT1 (N10302, N10301);
buf BUF1 (N10303, N10294);
not NOT1 (N10304, N10277);
xor XOR2 (N10305, N10299, N430);
nand NAND3 (N10306, N10303, N6681, N8843);
not NOT1 (N10307, N10304);
or OR3 (N10308, N10271, N1699, N7087);
or OR3 (N10309, N10306, N9619, N6518);
not NOT1 (N10310, N10298);
or OR4 (N10311, N10310, N10198, N3285, N6889);
or OR4 (N10312, N10302, N8608, N7451, N3760);
xor XOR2 (N10313, N10308, N4544);
nand NAND2 (N10314, N10300, N1848);
buf BUF1 (N10315, N10314);
nand NAND4 (N10316, N10313, N3150, N4798, N4703);
xor XOR2 (N10317, N10305, N4188);
nor NOR3 (N10318, N10288, N8009, N2270);
nand NAND4 (N10319, N10311, N7736, N1302, N7176);
xor XOR2 (N10320, N10309, N5117);
xor XOR2 (N10321, N10295, N3571);
buf BUF1 (N10322, N10296);
or OR4 (N10323, N10317, N8963, N8978, N3962);
or OR4 (N10324, N10307, N4847, N6592, N3217);
not NOT1 (N10325, N10320);
nor NOR3 (N10326, N10322, N7601, N1863);
not NOT1 (N10327, N10318);
nor NOR4 (N10328, N10315, N10041, N4499, N927);
and AND3 (N10329, N10328, N1964, N203);
buf BUF1 (N10330, N10321);
nand NAND4 (N10331, N10327, N6279, N10140, N5469);
or OR2 (N10332, N10326, N5035);
xor XOR2 (N10333, N10332, N7824);
not NOT1 (N10334, N10323);
nor NOR4 (N10335, N10325, N1594, N6276, N1934);
not NOT1 (N10336, N10329);
nand NAND2 (N10337, N10334, N2894);
not NOT1 (N10338, N10335);
buf BUF1 (N10339, N10319);
not NOT1 (N10340, N10312);
xor XOR2 (N10341, N10331, N1584);
or OR4 (N10342, N10339, N3015, N3781, N5902);
buf BUF1 (N10343, N10337);
xor XOR2 (N10344, N10342, N7618);
xor XOR2 (N10345, N10343, N5469);
not NOT1 (N10346, N10324);
buf BUF1 (N10347, N10338);
nor NOR4 (N10348, N10336, N5388, N5779, N9395);
not NOT1 (N10349, N10341);
nor NOR4 (N10350, N10346, N8653, N2172, N5703);
nor NOR2 (N10351, N10347, N3534);
or OR3 (N10352, N10316, N5703, N9162);
buf BUF1 (N10353, N10344);
not NOT1 (N10354, N10352);
and AND2 (N10355, N10353, N3763);
buf BUF1 (N10356, N10348);
nor NOR4 (N10357, N10333, N3933, N6576, N9139);
and AND2 (N10358, N10357, N1234);
xor XOR2 (N10359, N10358, N727);
or OR2 (N10360, N10359, N7638);
not NOT1 (N10361, N10354);
buf BUF1 (N10362, N10360);
or OR2 (N10363, N10330, N10186);
and AND2 (N10364, N10361, N10351);
or OR3 (N10365, N8091, N2930, N7302);
nand NAND4 (N10366, N10365, N3330, N4128, N5007);
nor NOR3 (N10367, N10356, N9239, N2582);
buf BUF1 (N10368, N10362);
xor XOR2 (N10369, N10355, N3463);
not NOT1 (N10370, N10369);
and AND3 (N10371, N10350, N1645, N596);
buf BUF1 (N10372, N10340);
buf BUF1 (N10373, N10370);
and AND2 (N10374, N10363, N387);
nand NAND3 (N10375, N10372, N6602, N4889);
buf BUF1 (N10376, N10366);
not NOT1 (N10377, N10376);
xor XOR2 (N10378, N10345, N8019);
xor XOR2 (N10379, N10378, N596);
nand NAND2 (N10380, N10373, N6811);
not NOT1 (N10381, N10380);
nor NOR3 (N10382, N10381, N7157, N6006);
and AND3 (N10383, N10382, N7780, N7320);
nor NOR3 (N10384, N10379, N10074, N781);
and AND2 (N10385, N10364, N5850);
buf BUF1 (N10386, N10367);
nor NOR3 (N10387, N10386, N7002, N4865);
or OR2 (N10388, N10384, N519);
nor NOR3 (N10389, N10383, N9239, N1522);
xor XOR2 (N10390, N10377, N3928);
and AND3 (N10391, N10389, N798, N9910);
or OR2 (N10392, N10390, N9375);
nor NOR2 (N10393, N10392, N6775);
or OR2 (N10394, N10385, N9467);
nor NOR2 (N10395, N10394, N1317);
xor XOR2 (N10396, N10395, N1734);
xor XOR2 (N10397, N10396, N47);
xor XOR2 (N10398, N10397, N5942);
buf BUF1 (N10399, N10371);
nand NAND4 (N10400, N10374, N8739, N1169, N4043);
and AND2 (N10401, N10393, N5313);
xor XOR2 (N10402, N10349, N10115);
or OR4 (N10403, N10387, N7115, N796, N7899);
buf BUF1 (N10404, N10399);
buf BUF1 (N10405, N10403);
nor NOR3 (N10406, N10404, N4767, N8627);
nand NAND2 (N10407, N10368, N10060);
buf BUF1 (N10408, N10391);
nor NOR3 (N10409, N10405, N3764, N6766);
nand NAND4 (N10410, N10388, N753, N9441, N6489);
xor XOR2 (N10411, N10375, N1247);
and AND2 (N10412, N10401, N7786);
buf BUF1 (N10413, N10408);
or OR4 (N10414, N10400, N9677, N8327, N2488);
nor NOR3 (N10415, N10410, N9494, N2780);
and AND4 (N10416, N10398, N8844, N1495, N9626);
buf BUF1 (N10417, N10415);
nor NOR3 (N10418, N10417, N5729, N2051);
not NOT1 (N10419, N10416);
or OR4 (N10420, N10407, N81, N13, N8349);
or OR4 (N10421, N10402, N3993, N1741, N1881);
xor XOR2 (N10422, N10413, N3190);
or OR3 (N10423, N10420, N2830, N3054);
nand NAND4 (N10424, N10419, N273, N431, N2204);
xor XOR2 (N10425, N10421, N10233);
nand NAND4 (N10426, N10411, N9713, N4444, N6228);
not NOT1 (N10427, N10418);
xor XOR2 (N10428, N10423, N9439);
nand NAND2 (N10429, N10406, N1689);
nor NOR2 (N10430, N10426, N892);
or OR4 (N10431, N10425, N7385, N8377, N8415);
not NOT1 (N10432, N10430);
not NOT1 (N10433, N10414);
or OR2 (N10434, N10429, N4630);
nor NOR4 (N10435, N10412, N2123, N5993, N10294);
xor XOR2 (N10436, N10428, N4933);
not NOT1 (N10437, N10435);
buf BUF1 (N10438, N10409);
not NOT1 (N10439, N10427);
or OR2 (N10440, N10431, N9946);
xor XOR2 (N10441, N10440, N793);
or OR4 (N10442, N10441, N5758, N1657, N6465);
nand NAND2 (N10443, N10438, N484);
nor NOR2 (N10444, N10436, N9073);
xor XOR2 (N10445, N10434, N36);
nand NAND4 (N10446, N10443, N9224, N5395, N5952);
nand NAND3 (N10447, N10432, N7624, N9062);
xor XOR2 (N10448, N10442, N10330);
nor NOR3 (N10449, N10439, N144, N10439);
nor NOR2 (N10450, N10447, N6408);
not NOT1 (N10451, N10437);
nand NAND2 (N10452, N10444, N76);
buf BUF1 (N10453, N10424);
or OR2 (N10454, N10448, N6334);
xor XOR2 (N10455, N10446, N7336);
and AND4 (N10456, N10449, N4724, N5214, N8297);
or OR3 (N10457, N10422, N4421, N8672);
not NOT1 (N10458, N10455);
nor NOR3 (N10459, N10458, N9771, N10120);
buf BUF1 (N10460, N10453);
xor XOR2 (N10461, N10459, N4719);
xor XOR2 (N10462, N10454, N4923);
buf BUF1 (N10463, N10452);
and AND4 (N10464, N10461, N7553, N3386, N2997);
and AND3 (N10465, N10433, N1534, N3684);
xor XOR2 (N10466, N10456, N6127);
or OR2 (N10467, N10451, N5752);
and AND4 (N10468, N10467, N8701, N10126, N1831);
not NOT1 (N10469, N10457);
nand NAND3 (N10470, N10460, N6621, N8555);
and AND3 (N10471, N10465, N460, N7576);
xor XOR2 (N10472, N10470, N3938);
buf BUF1 (N10473, N10472);
nor NOR2 (N10474, N10469, N6496);
and AND4 (N10475, N10466, N167, N5860, N6682);
or OR3 (N10476, N10473, N4728, N250);
xor XOR2 (N10477, N10450, N8064);
xor XOR2 (N10478, N10463, N10327);
xor XOR2 (N10479, N10474, N6302);
buf BUF1 (N10480, N10468);
nand NAND2 (N10481, N10479, N5288);
and AND3 (N10482, N10462, N3135, N5463);
buf BUF1 (N10483, N10481);
nand NAND2 (N10484, N10471, N10356);
xor XOR2 (N10485, N10484, N1962);
xor XOR2 (N10486, N10482, N9508);
buf BUF1 (N10487, N10478);
and AND4 (N10488, N10476, N6133, N8654, N1789);
xor XOR2 (N10489, N10483, N1192);
or OR2 (N10490, N10488, N7299);
nor NOR2 (N10491, N10464, N10165);
nand NAND3 (N10492, N10445, N3917, N10049);
or OR3 (N10493, N10486, N6717, N3148);
and AND2 (N10494, N10491, N2891);
not NOT1 (N10495, N10480);
not NOT1 (N10496, N10489);
xor XOR2 (N10497, N10493, N6214);
buf BUF1 (N10498, N10497);
nand NAND3 (N10499, N10490, N2193, N8489);
not NOT1 (N10500, N10498);
xor XOR2 (N10501, N10494, N9798);
nand NAND3 (N10502, N10500, N1078, N4839);
nand NAND3 (N10503, N10477, N21, N1857);
and AND3 (N10504, N10499, N9393, N5072);
xor XOR2 (N10505, N10503, N2765);
nand NAND2 (N10506, N10501, N4948);
not NOT1 (N10507, N10495);
xor XOR2 (N10508, N10502, N1891);
xor XOR2 (N10509, N10506, N2255);
or OR2 (N10510, N10504, N7053);
nand NAND3 (N10511, N10475, N6804, N2507);
buf BUF1 (N10512, N10505);
and AND3 (N10513, N10509, N5598, N5016);
or OR4 (N10514, N10512, N1002, N8028, N2034);
buf BUF1 (N10515, N10485);
xor XOR2 (N10516, N10508, N425);
or OR2 (N10517, N10515, N6434);
buf BUF1 (N10518, N10516);
and AND4 (N10519, N10507, N8779, N8578, N10102);
buf BUF1 (N10520, N10496);
or OR3 (N10521, N10518, N9579, N4625);
buf BUF1 (N10522, N10487);
and AND2 (N10523, N10510, N7961);
buf BUF1 (N10524, N10517);
xor XOR2 (N10525, N10514, N3852);
not NOT1 (N10526, N10511);
nor NOR3 (N10527, N10492, N7863, N4164);
not NOT1 (N10528, N10523);
and AND4 (N10529, N10519, N173, N230, N1613);
not NOT1 (N10530, N10513);
xor XOR2 (N10531, N10529, N1366);
or OR2 (N10532, N10524, N6022);
buf BUF1 (N10533, N10525);
buf BUF1 (N10534, N10530);
and AND2 (N10535, N10534, N7091);
not NOT1 (N10536, N10532);
buf BUF1 (N10537, N10521);
xor XOR2 (N10538, N10522, N6986);
xor XOR2 (N10539, N10537, N6903);
nand NAND3 (N10540, N10520, N10196, N6710);
nand NAND4 (N10541, N10536, N3762, N6858, N6652);
buf BUF1 (N10542, N10531);
or OR2 (N10543, N10528, N1149);
nand NAND3 (N10544, N10541, N4538, N9459);
nor NOR3 (N10545, N10527, N4905, N8155);
or OR3 (N10546, N10533, N7270, N4404);
nor NOR4 (N10547, N10538, N1413, N5809, N4558);
not NOT1 (N10548, N10546);
nor NOR2 (N10549, N10539, N7505);
nor NOR2 (N10550, N10547, N4392);
nor NOR2 (N10551, N10542, N9814);
xor XOR2 (N10552, N10549, N4504);
nor NOR3 (N10553, N10552, N9462, N3807);
xor XOR2 (N10554, N10553, N9997);
and AND3 (N10555, N10535, N9908, N10511);
xor XOR2 (N10556, N10543, N6745);
buf BUF1 (N10557, N10555);
and AND2 (N10558, N10556, N4226);
or OR3 (N10559, N10526, N7947, N30);
nand NAND4 (N10560, N10558, N1452, N8140, N5703);
nand NAND3 (N10561, N10544, N2260, N9396);
and AND4 (N10562, N10557, N9130, N3013, N1362);
and AND3 (N10563, N10560, N1792, N10142);
xor XOR2 (N10564, N10551, N3690);
nand NAND2 (N10565, N10559, N231);
not NOT1 (N10566, N10545);
xor XOR2 (N10567, N10564, N2675);
and AND2 (N10568, N10566, N3803);
and AND4 (N10569, N10567, N4009, N6491, N3707);
not NOT1 (N10570, N10554);
xor XOR2 (N10571, N10563, N9580);
nor NOR2 (N10572, N10561, N1660);
and AND3 (N10573, N10550, N9858, N10474);
nor NOR4 (N10574, N10562, N8918, N5746, N6816);
or OR4 (N10575, N10570, N10263, N9691, N3027);
and AND2 (N10576, N10573, N380);
and AND3 (N10577, N10576, N6780, N3205);
not NOT1 (N10578, N10574);
nand NAND3 (N10579, N10575, N6805, N7651);
not NOT1 (N10580, N10579);
xor XOR2 (N10581, N10548, N1748);
nand NAND4 (N10582, N10565, N393, N8339, N6000);
buf BUF1 (N10583, N10581);
not NOT1 (N10584, N10582);
nand NAND4 (N10585, N10569, N1444, N9915, N4602);
nand NAND4 (N10586, N10568, N10309, N4535, N313);
or OR3 (N10587, N10584, N9130, N5682);
not NOT1 (N10588, N10583);
buf BUF1 (N10589, N10587);
xor XOR2 (N10590, N10540, N7601);
or OR4 (N10591, N10572, N9657, N3135, N6134);
nand NAND2 (N10592, N10578, N10053);
buf BUF1 (N10593, N10585);
nand NAND3 (N10594, N10589, N3194, N6146);
or OR3 (N10595, N10590, N1627, N6533);
or OR2 (N10596, N10588, N3274);
or OR4 (N10597, N10593, N1235, N7718, N2918);
and AND4 (N10598, N10592, N3887, N3733, N1468);
xor XOR2 (N10599, N10595, N9470);
and AND4 (N10600, N10571, N3021, N6690, N2505);
and AND4 (N10601, N10597, N822, N9470, N8770);
nand NAND2 (N10602, N10577, N4299);
or OR3 (N10603, N10580, N4594, N9395);
buf BUF1 (N10604, N10591);
nor NOR3 (N10605, N10602, N1307, N6166);
xor XOR2 (N10606, N10586, N452);
or OR3 (N10607, N10603, N10449, N2925);
or OR2 (N10608, N10601, N2795);
nand NAND3 (N10609, N10600, N3185, N9222);
nor NOR2 (N10610, N10599, N8381);
nand NAND4 (N10611, N10604, N1551, N1458, N17);
nor NOR2 (N10612, N10598, N6429);
or OR3 (N10613, N10607, N5817, N7219);
not NOT1 (N10614, N10611);
not NOT1 (N10615, N10605);
nor NOR4 (N10616, N10612, N4264, N578, N4161);
and AND4 (N10617, N10609, N5407, N376, N2488);
buf BUF1 (N10618, N10594);
and AND4 (N10619, N10606, N6129, N4616, N3058);
or OR4 (N10620, N10608, N6764, N1889, N2091);
or OR2 (N10621, N10616, N6953);
nand NAND4 (N10622, N10618, N5881, N269, N7955);
nand NAND3 (N10623, N10614, N6551, N4724);
xor XOR2 (N10624, N10620, N7898);
buf BUF1 (N10625, N10622);
buf BUF1 (N10626, N10621);
not NOT1 (N10627, N10596);
xor XOR2 (N10628, N10619, N3952);
or OR3 (N10629, N10627, N5634, N4560);
or OR3 (N10630, N10610, N9303, N7375);
xor XOR2 (N10631, N10629, N9093);
or OR2 (N10632, N10624, N4430);
nand NAND3 (N10633, N10631, N3704, N7777);
and AND4 (N10634, N10613, N8541, N4687, N10410);
buf BUF1 (N10635, N10626);
buf BUF1 (N10636, N10623);
not NOT1 (N10637, N10633);
xor XOR2 (N10638, N10632, N7243);
buf BUF1 (N10639, N10628);
buf BUF1 (N10640, N10630);
or OR3 (N10641, N10640, N2813, N4530);
nor NOR2 (N10642, N10636, N4823);
nand NAND2 (N10643, N10638, N9609);
xor XOR2 (N10644, N10617, N10285);
nand NAND4 (N10645, N10639, N10454, N6137, N8048);
or OR2 (N10646, N10637, N4954);
buf BUF1 (N10647, N10646);
and AND4 (N10648, N10644, N1245, N10470, N10631);
xor XOR2 (N10649, N10642, N8853);
and AND3 (N10650, N10648, N10348, N2074);
nor NOR3 (N10651, N10645, N155, N420);
nand NAND3 (N10652, N10634, N4539, N5097);
buf BUF1 (N10653, N10641);
buf BUF1 (N10654, N10650);
nor NOR3 (N10655, N10653, N2753, N3046);
not NOT1 (N10656, N10655);
xor XOR2 (N10657, N10654, N4457);
or OR4 (N10658, N10657, N3584, N4068, N10568);
not NOT1 (N10659, N10643);
xor XOR2 (N10660, N10652, N8122);
xor XOR2 (N10661, N10659, N6769);
not NOT1 (N10662, N10625);
not NOT1 (N10663, N10656);
buf BUF1 (N10664, N10635);
nand NAND2 (N10665, N10661, N4370);
nor NOR2 (N10666, N10658, N3389);
nor NOR2 (N10667, N10665, N3612);
buf BUF1 (N10668, N10667);
not NOT1 (N10669, N10660);
nor NOR3 (N10670, N10669, N1882, N6531);
buf BUF1 (N10671, N10651);
xor XOR2 (N10672, N10647, N6470);
nand NAND4 (N10673, N10672, N10622, N3252, N442);
or OR3 (N10674, N10666, N5721, N8901);
or OR4 (N10675, N10674, N9740, N9810, N3338);
nand NAND3 (N10676, N10664, N3154, N3456);
nor NOR4 (N10677, N10662, N10319, N5824, N9500);
not NOT1 (N10678, N10663);
not NOT1 (N10679, N10668);
nand NAND2 (N10680, N10677, N5612);
and AND3 (N10681, N10615, N5022, N535);
nand NAND3 (N10682, N10671, N5411, N8608);
or OR2 (N10683, N10649, N6177);
nor NOR3 (N10684, N10681, N10313, N854);
or OR2 (N10685, N10670, N6711);
xor XOR2 (N10686, N10675, N6398);
or OR2 (N10687, N10678, N4608);
and AND2 (N10688, N10680, N2121);
and AND2 (N10689, N10673, N1970);
not NOT1 (N10690, N10684);
nor NOR3 (N10691, N10687, N4303, N8643);
buf BUF1 (N10692, N10679);
and AND4 (N10693, N10676, N3790, N101, N4586);
and AND3 (N10694, N10691, N3890, N7410);
nor NOR4 (N10695, N10693, N1174, N2455, N10246);
and AND4 (N10696, N10692, N9701, N9950, N6138);
buf BUF1 (N10697, N10686);
xor XOR2 (N10698, N10689, N6013);
or OR2 (N10699, N10688, N3730);
xor XOR2 (N10700, N10682, N493);
not NOT1 (N10701, N10694);
or OR3 (N10702, N10700, N5262, N1131);
nor NOR3 (N10703, N10696, N6138, N9013);
nor NOR4 (N10704, N10699, N4587, N5273, N2774);
nand NAND3 (N10705, N10701, N7876, N2313);
nor NOR3 (N10706, N10702, N1370, N284);
nor NOR2 (N10707, N10697, N5797);
xor XOR2 (N10708, N10706, N4780);
and AND3 (N10709, N10685, N7274, N6205);
or OR2 (N10710, N10709, N3464);
nand NAND2 (N10711, N10683, N988);
xor XOR2 (N10712, N10703, N275);
nand NAND3 (N10713, N10708, N6651, N6256);
or OR4 (N10714, N10704, N9568, N4551, N6275);
nor NOR3 (N10715, N10707, N9439, N7088);
xor XOR2 (N10716, N10711, N1230);
nand NAND2 (N10717, N10713, N5079);
or OR3 (N10718, N10717, N6854, N4998);
buf BUF1 (N10719, N10695);
buf BUF1 (N10720, N10712);
xor XOR2 (N10721, N10716, N7689);
not NOT1 (N10722, N10720);
and AND4 (N10723, N10705, N3698, N7166, N2584);
nor NOR4 (N10724, N10698, N132, N975, N94);
buf BUF1 (N10725, N10724);
and AND3 (N10726, N10719, N929, N1427);
nor NOR4 (N10727, N10715, N10138, N7322, N6495);
nor NOR3 (N10728, N10726, N7255, N7267);
nor NOR4 (N10729, N10690, N7292, N9214, N6696);
nand NAND3 (N10730, N10727, N4963, N10613);
xor XOR2 (N10731, N10730, N1002);
buf BUF1 (N10732, N10731);
not NOT1 (N10733, N10718);
buf BUF1 (N10734, N10732);
xor XOR2 (N10735, N10721, N10581);
or OR4 (N10736, N10728, N6743, N8928, N3513);
and AND2 (N10737, N10734, N5032);
and AND2 (N10738, N10729, N6509);
not NOT1 (N10739, N10737);
nand NAND4 (N10740, N10733, N3531, N5253, N3586);
not NOT1 (N10741, N10736);
nor NOR2 (N10742, N10714, N9505);
nor NOR4 (N10743, N10742, N2674, N10275, N9470);
nor NOR2 (N10744, N10722, N2561);
nor NOR4 (N10745, N10744, N3106, N1101, N3303);
buf BUF1 (N10746, N10743);
nand NAND4 (N10747, N10710, N2642, N1154, N1260);
or OR2 (N10748, N10738, N3829);
xor XOR2 (N10749, N10741, N2105);
nor NOR3 (N10750, N10745, N661, N6435);
or OR2 (N10751, N10748, N10181);
xor XOR2 (N10752, N10725, N5196);
and AND3 (N10753, N10740, N8536, N7695);
nand NAND3 (N10754, N10739, N5308, N10024);
nand NAND4 (N10755, N10749, N3437, N3476, N5584);
nor NOR3 (N10756, N10723, N7162, N4259);
and AND4 (N10757, N10754, N1315, N4337, N6037);
nor NOR3 (N10758, N10735, N4801, N4366);
buf BUF1 (N10759, N10751);
or OR4 (N10760, N10752, N2018, N7219, N4712);
and AND4 (N10761, N10760, N4880, N2679, N10733);
and AND4 (N10762, N10753, N3427, N6815, N5773);
not NOT1 (N10763, N10762);
or OR2 (N10764, N10763, N401);
nor NOR2 (N10765, N10757, N6812);
and AND3 (N10766, N10747, N10196, N8769);
and AND2 (N10767, N10766, N2009);
not NOT1 (N10768, N10758);
buf BUF1 (N10769, N10768);
xor XOR2 (N10770, N10767, N9898);
or OR4 (N10771, N10770, N3446, N2838, N8711);
nor NOR4 (N10772, N10769, N5995, N8566, N10389);
buf BUF1 (N10773, N10761);
or OR4 (N10774, N10750, N2789, N2385, N2247);
and AND4 (N10775, N10755, N2033, N2444, N5538);
nor NOR3 (N10776, N10771, N8371, N4549);
or OR3 (N10777, N10774, N8203, N1033);
not NOT1 (N10778, N10759);
nor NOR2 (N10779, N10778, N3646);
xor XOR2 (N10780, N10779, N9763);
nor NOR2 (N10781, N10777, N1767);
or OR4 (N10782, N10776, N973, N3212, N8513);
nor NOR3 (N10783, N10765, N2413, N1752);
buf BUF1 (N10784, N10783);
not NOT1 (N10785, N10784);
xor XOR2 (N10786, N10775, N9429);
or OR3 (N10787, N10785, N6084, N5709);
not NOT1 (N10788, N10782);
or OR3 (N10789, N10764, N9865, N1356);
nor NOR4 (N10790, N10787, N3628, N3398, N2623);
buf BUF1 (N10791, N10756);
buf BUF1 (N10792, N10786);
xor XOR2 (N10793, N10789, N7106);
xor XOR2 (N10794, N10790, N3729);
or OR3 (N10795, N10788, N10351, N4125);
xor XOR2 (N10796, N10793, N2136);
and AND4 (N10797, N10781, N4721, N1587, N6296);
buf BUF1 (N10798, N10795);
xor XOR2 (N10799, N10772, N3173);
nand NAND4 (N10800, N10746, N2282, N4075, N2201);
nor NOR3 (N10801, N10796, N6657, N8305);
not NOT1 (N10802, N10799);
nor NOR4 (N10803, N10797, N9107, N4446, N5388);
buf BUF1 (N10804, N10773);
nor NOR4 (N10805, N10780, N2935, N8495, N401);
not NOT1 (N10806, N10803);
buf BUF1 (N10807, N10805);
xor XOR2 (N10808, N10792, N1978);
not NOT1 (N10809, N10794);
and AND2 (N10810, N10801, N9699);
not NOT1 (N10811, N10809);
nor NOR4 (N10812, N10811, N2005, N10739, N9111);
nand NAND3 (N10813, N10798, N342, N4927);
not NOT1 (N10814, N10810);
not NOT1 (N10815, N10800);
and AND2 (N10816, N10808, N9140);
and AND4 (N10817, N10812, N1441, N8113, N10058);
nor NOR3 (N10818, N10815, N4241, N384);
or OR2 (N10819, N10791, N6324);
nor NOR3 (N10820, N10816, N3044, N10138);
xor XOR2 (N10821, N10807, N4126);
xor XOR2 (N10822, N10802, N3623);
nand NAND3 (N10823, N10820, N10678, N2557);
not NOT1 (N10824, N10814);
buf BUF1 (N10825, N10822);
nand NAND4 (N10826, N10825, N4242, N2230, N8041);
or OR4 (N10827, N10813, N3507, N983, N10511);
nor NOR3 (N10828, N10806, N10594, N2665);
xor XOR2 (N10829, N10818, N5983);
and AND4 (N10830, N10817, N8950, N7725, N5850);
nand NAND3 (N10831, N10823, N10052, N4002);
not NOT1 (N10832, N10826);
nand NAND4 (N10833, N10831, N9924, N22, N8792);
or OR2 (N10834, N10833, N10281);
not NOT1 (N10835, N10832);
xor XOR2 (N10836, N10830, N46);
xor XOR2 (N10837, N10834, N4767);
nand NAND4 (N10838, N10828, N5214, N8222, N2857);
and AND4 (N10839, N10835, N6164, N1900, N1679);
not NOT1 (N10840, N10804);
xor XOR2 (N10841, N10839, N3324);
nand NAND3 (N10842, N10836, N8034, N5691);
nand NAND3 (N10843, N10821, N7055, N7567);
nand NAND2 (N10844, N10829, N4863);
or OR2 (N10845, N10843, N9567);
nor NOR3 (N10846, N10838, N7528, N10414);
nand NAND2 (N10847, N10824, N10430);
buf BUF1 (N10848, N10837);
buf BUF1 (N10849, N10848);
nand NAND4 (N10850, N10844, N2368, N3977, N5561);
nor NOR3 (N10851, N10850, N7181, N3602);
not NOT1 (N10852, N10851);
or OR3 (N10853, N10847, N3654, N2981);
or OR3 (N10854, N10842, N9105, N9054);
and AND4 (N10855, N10852, N10670, N7123, N4957);
xor XOR2 (N10856, N10846, N8093);
and AND4 (N10857, N10853, N4176, N5246, N369);
nand NAND2 (N10858, N10849, N8498);
not NOT1 (N10859, N10845);
not NOT1 (N10860, N10856);
nor NOR3 (N10861, N10857, N622, N4665);
nand NAND3 (N10862, N10841, N7984, N1925);
and AND2 (N10863, N10854, N9186);
not NOT1 (N10864, N10819);
buf BUF1 (N10865, N10827);
not NOT1 (N10866, N10862);
nand NAND2 (N10867, N10860, N3098);
or OR4 (N10868, N10866, N10257, N2060, N2699);
or OR3 (N10869, N10865, N7544, N1704);
buf BUF1 (N10870, N10869);
nor NOR3 (N10871, N10859, N4390, N9083);
and AND3 (N10872, N10861, N2972, N6649);
nand NAND2 (N10873, N10868, N1211);
buf BUF1 (N10874, N10855);
nand NAND3 (N10875, N10840, N3754, N1719);
or OR4 (N10876, N10875, N10765, N7797, N1752);
nand NAND4 (N10877, N10858, N2936, N10251, N6871);
buf BUF1 (N10878, N10867);
nand NAND2 (N10879, N10874, N2486);
nor NOR3 (N10880, N10879, N6221, N3006);
and AND4 (N10881, N10880, N116, N6078, N1996);
not NOT1 (N10882, N10870);
nor NOR4 (N10883, N10877, N284, N9371, N9496);
buf BUF1 (N10884, N10871);
xor XOR2 (N10885, N10863, N9817);
and AND2 (N10886, N10884, N2462);
and AND4 (N10887, N10864, N631, N9518, N7004);
nand NAND4 (N10888, N10872, N2149, N6487, N1954);
nand NAND3 (N10889, N10886, N3897, N10312);
not NOT1 (N10890, N10876);
and AND2 (N10891, N10873, N2046);
and AND3 (N10892, N10891, N1118, N10520);
and AND2 (N10893, N10890, N5111);
nor NOR2 (N10894, N10889, N6751);
or OR2 (N10895, N10892, N7665);
nand NAND2 (N10896, N10885, N3638);
and AND2 (N10897, N10895, N3415);
not NOT1 (N10898, N10888);
nor NOR2 (N10899, N10882, N2516);
xor XOR2 (N10900, N10887, N8199);
not NOT1 (N10901, N10883);
nor NOR3 (N10902, N10898, N3318, N4877);
xor XOR2 (N10903, N10901, N1893);
not NOT1 (N10904, N10899);
nand NAND3 (N10905, N10900, N5534, N9845);
buf BUF1 (N10906, N10878);
or OR4 (N10907, N10903, N9367, N1787, N658);
not NOT1 (N10908, N10907);
or OR4 (N10909, N10881, N2731, N8092, N3710);
xor XOR2 (N10910, N10904, N3987);
nor NOR3 (N10911, N10897, N6737, N10236);
buf BUF1 (N10912, N10902);
xor XOR2 (N10913, N10908, N8614);
nand NAND2 (N10914, N10896, N6561);
or OR2 (N10915, N10905, N940);
nor NOR3 (N10916, N10906, N4270, N10667);
not NOT1 (N10917, N10893);
buf BUF1 (N10918, N10917);
and AND2 (N10919, N10915, N10769);
and AND3 (N10920, N10918, N7590, N7414);
nand NAND2 (N10921, N10912, N4288);
or OR2 (N10922, N10894, N2768);
or OR2 (N10923, N10921, N10074);
and AND3 (N10924, N10913, N10827, N9583);
not NOT1 (N10925, N10919);
not NOT1 (N10926, N10925);
nand NAND4 (N10927, N10920, N271, N9828, N347);
and AND2 (N10928, N10914, N1260);
or OR3 (N10929, N10916, N8524, N4332);
nor NOR4 (N10930, N10923, N9019, N6098, N3354);
nor NOR3 (N10931, N10910, N9858, N3987);
and AND2 (N10932, N10922, N7717);
nand NAND3 (N10933, N10924, N9678, N1151);
or OR3 (N10934, N10932, N6905, N7215);
not NOT1 (N10935, N10911);
nor NOR2 (N10936, N10928, N6008);
buf BUF1 (N10937, N10927);
not NOT1 (N10938, N10926);
nand NAND4 (N10939, N10937, N1014, N8158, N1493);
xor XOR2 (N10940, N10938, N8207);
or OR2 (N10941, N10935, N8842);
or OR2 (N10942, N10930, N2191);
or OR3 (N10943, N10933, N1990, N756);
xor XOR2 (N10944, N10929, N9254);
xor XOR2 (N10945, N10940, N3130);
nor NOR2 (N10946, N10941, N8828);
xor XOR2 (N10947, N10946, N6720);
xor XOR2 (N10948, N10934, N3371);
nor NOR2 (N10949, N10947, N8663);
not NOT1 (N10950, N10945);
buf BUF1 (N10951, N10936);
buf BUF1 (N10952, N10909);
not NOT1 (N10953, N10948);
xor XOR2 (N10954, N10953, N2377);
buf BUF1 (N10955, N10950);
xor XOR2 (N10956, N10931, N6856);
and AND4 (N10957, N10952, N5210, N3834, N10019);
nor NOR3 (N10958, N10954, N6458, N2245);
nand NAND4 (N10959, N10955, N5148, N2232, N2192);
or OR3 (N10960, N10949, N3225, N4707);
or OR4 (N10961, N10958, N10185, N3428, N543);
xor XOR2 (N10962, N10944, N6557);
buf BUF1 (N10963, N10959);
xor XOR2 (N10964, N10951, N3697);
or OR4 (N10965, N10963, N5876, N6749, N9563);
buf BUF1 (N10966, N10943);
buf BUF1 (N10967, N10939);
nand NAND4 (N10968, N10964, N5423, N5509, N941);
xor XOR2 (N10969, N10967, N8336);
buf BUF1 (N10970, N10956);
nand NAND3 (N10971, N10966, N6085, N3016);
nand NAND2 (N10972, N10942, N10704);
buf BUF1 (N10973, N10970);
xor XOR2 (N10974, N10973, N10615);
buf BUF1 (N10975, N10974);
nor NOR2 (N10976, N10962, N9863);
or OR4 (N10977, N10965, N9386, N3136, N10635);
not NOT1 (N10978, N10969);
or OR2 (N10979, N10978, N2130);
not NOT1 (N10980, N10971);
not NOT1 (N10981, N10972);
and AND2 (N10982, N10960, N5514);
xor XOR2 (N10983, N10981, N9952);
and AND3 (N10984, N10977, N9453, N472);
nor NOR3 (N10985, N10968, N4273, N9179);
or OR4 (N10986, N10984, N2773, N4200, N3579);
xor XOR2 (N10987, N10982, N7267);
buf BUF1 (N10988, N10983);
nor NOR2 (N10989, N10957, N4222);
not NOT1 (N10990, N10989);
buf BUF1 (N10991, N10988);
nor NOR3 (N10992, N10990, N10388, N6544);
nand NAND2 (N10993, N10976, N272);
not NOT1 (N10994, N10975);
or OR3 (N10995, N10993, N2530, N6188);
or OR3 (N10996, N10980, N2400, N6024);
and AND3 (N10997, N10992, N1232, N375);
xor XOR2 (N10998, N10994, N7589);
or OR2 (N10999, N10979, N5127);
nand NAND3 (N11000, N10987, N8996, N1017);
buf BUF1 (N11001, N10985);
nand NAND3 (N11002, N10998, N2993, N10636);
not NOT1 (N11003, N11000);
or OR4 (N11004, N10986, N1290, N7599, N10165);
buf BUF1 (N11005, N11004);
xor XOR2 (N11006, N11003, N1067);
nand NAND2 (N11007, N11006, N3474);
not NOT1 (N11008, N10997);
or OR2 (N11009, N10961, N9958);
not NOT1 (N11010, N11002);
nor NOR4 (N11011, N10999, N6862, N689, N4557);
nor NOR3 (N11012, N11010, N1195, N10386);
and AND2 (N11013, N11011, N9388);
nor NOR4 (N11014, N11012, N8228, N8763, N10122);
or OR2 (N11015, N11014, N5756);
and AND3 (N11016, N11013, N9951, N3827);
nand NAND4 (N11017, N10995, N6920, N4759, N1526);
or OR3 (N11018, N10996, N1282, N6023);
not NOT1 (N11019, N11009);
buf BUF1 (N11020, N11016);
buf BUF1 (N11021, N11008);
not NOT1 (N11022, N11019);
or OR4 (N11023, N11021, N2139, N5721, N3860);
or OR4 (N11024, N11007, N5685, N10470, N8146);
xor XOR2 (N11025, N11022, N3344);
buf BUF1 (N11026, N11005);
nand NAND3 (N11027, N11025, N7134, N4610);
nor NOR2 (N11028, N11017, N3549);
xor XOR2 (N11029, N11026, N7723);
nand NAND3 (N11030, N11024, N6301, N3988);
and AND4 (N11031, N11018, N5881, N902, N3495);
or OR2 (N11032, N11029, N2400);
not NOT1 (N11033, N11032);
not NOT1 (N11034, N10991);
and AND4 (N11035, N11034, N9653, N10509, N8970);
buf BUF1 (N11036, N11020);
nand NAND4 (N11037, N11035, N3387, N3100, N4717);
buf BUF1 (N11038, N11001);
nand NAND3 (N11039, N11031, N4549, N5747);
and AND2 (N11040, N11037, N6366);
buf BUF1 (N11041, N11036);
nor NOR4 (N11042, N11040, N7722, N3012, N4593);
and AND3 (N11043, N11028, N7413, N11005);
xor XOR2 (N11044, N11023, N5370);
nor NOR3 (N11045, N11027, N7613, N7337);
not NOT1 (N11046, N11030);
not NOT1 (N11047, N11043);
nand NAND4 (N11048, N11042, N2420, N6926, N9674);
not NOT1 (N11049, N11015);
not NOT1 (N11050, N11046);
buf BUF1 (N11051, N11039);
nand NAND3 (N11052, N11038, N8125, N7672);
not NOT1 (N11053, N11045);
nand NAND4 (N11054, N11041, N693, N7596, N2440);
nor NOR2 (N11055, N11051, N4981);
buf BUF1 (N11056, N11052);
not NOT1 (N11057, N11054);
nor NOR3 (N11058, N11053, N3325, N10175);
or OR4 (N11059, N11044, N1800, N9379, N9195);
or OR2 (N11060, N11033, N3501);
and AND3 (N11061, N11047, N1795, N1817);
nand NAND4 (N11062, N11055, N5459, N9676, N3923);
nand NAND4 (N11063, N11058, N8007, N1966, N7520);
or OR3 (N11064, N11049, N3628, N10587);
and AND2 (N11065, N11050, N9716);
not NOT1 (N11066, N11060);
and AND2 (N11067, N11064, N3773);
or OR3 (N11068, N11056, N11064, N6605);
or OR2 (N11069, N11061, N9604);
xor XOR2 (N11070, N11063, N3052);
nor NOR3 (N11071, N11068, N4230, N4302);
not NOT1 (N11072, N11065);
not NOT1 (N11073, N11057);
nor NOR3 (N11074, N11048, N2255, N175);
or OR3 (N11075, N11070, N2367, N779);
or OR3 (N11076, N11075, N7606, N3742);
nor NOR2 (N11077, N11074, N822);
or OR2 (N11078, N11062, N5996);
nand NAND4 (N11079, N11069, N3133, N10665, N6735);
nor NOR2 (N11080, N11073, N6409);
xor XOR2 (N11081, N11076, N6756);
not NOT1 (N11082, N11059);
xor XOR2 (N11083, N11078, N935);
not NOT1 (N11084, N11072);
xor XOR2 (N11085, N11077, N2394);
not NOT1 (N11086, N11066);
nor NOR3 (N11087, N11080, N1436, N6119);
nand NAND3 (N11088, N11087, N10317, N9102);
not NOT1 (N11089, N11079);
nand NAND4 (N11090, N11083, N2227, N7562, N8686);
nand NAND3 (N11091, N11090, N3367, N314);
and AND4 (N11092, N11084, N6812, N3690, N2487);
xor XOR2 (N11093, N11089, N6292);
buf BUF1 (N11094, N11081);
nor NOR4 (N11095, N11071, N6533, N9897, N923);
nor NOR2 (N11096, N11093, N1208);
nor NOR3 (N11097, N11085, N41, N6258);
nand NAND2 (N11098, N11091, N9632);
or OR4 (N11099, N11097, N5445, N9283, N6782);
and AND2 (N11100, N11082, N7994);
not NOT1 (N11101, N11100);
nand NAND4 (N11102, N11088, N6895, N2490, N9929);
or OR4 (N11103, N11095, N9552, N8617, N8039);
nand NAND2 (N11104, N11067, N1541);
nand NAND3 (N11105, N11104, N5255, N5358);
xor XOR2 (N11106, N11098, N4418);
and AND2 (N11107, N11092, N3661);
and AND4 (N11108, N11102, N5831, N842, N7380);
and AND3 (N11109, N11106, N6777, N79);
or OR2 (N11110, N11103, N231);
buf BUF1 (N11111, N11105);
nand NAND4 (N11112, N11086, N6313, N702, N3658);
buf BUF1 (N11113, N11101);
nor NOR2 (N11114, N11110, N5227);
not NOT1 (N11115, N11094);
or OR4 (N11116, N11112, N6469, N7450, N5840);
nand NAND3 (N11117, N11114, N5895, N9679);
and AND3 (N11118, N11116, N8242, N2114);
not NOT1 (N11119, N11099);
buf BUF1 (N11120, N11096);
nor NOR2 (N11121, N11115, N2553);
xor XOR2 (N11122, N11111, N4035);
buf BUF1 (N11123, N11120);
not NOT1 (N11124, N11121);
not NOT1 (N11125, N11109);
buf BUF1 (N11126, N11108);
not NOT1 (N11127, N11117);
or OR3 (N11128, N11126, N2739, N8103);
not NOT1 (N11129, N11122);
and AND3 (N11130, N11107, N2504, N3320);
nand NAND3 (N11131, N11113, N4910, N4584);
buf BUF1 (N11132, N11129);
or OR3 (N11133, N11130, N4833, N5636);
not NOT1 (N11134, N11119);
and AND4 (N11135, N11127, N2300, N3227, N1035);
nor NOR4 (N11136, N11133, N6347, N6784, N4355);
not NOT1 (N11137, N11131);
nor NOR4 (N11138, N11134, N3276, N6914, N1267);
nand NAND3 (N11139, N11137, N6365, N7324);
nor NOR4 (N11140, N11118, N3055, N759, N7738);
or OR4 (N11141, N11138, N836, N7111, N3906);
nand NAND2 (N11142, N11123, N456);
nor NOR2 (N11143, N11139, N10131);
nor NOR3 (N11144, N11124, N2277, N10010);
xor XOR2 (N11145, N11141, N5300);
nand NAND2 (N11146, N11143, N3895);
not NOT1 (N11147, N11146);
and AND2 (N11148, N11128, N8294);
or OR3 (N11149, N11136, N10809, N21);
xor XOR2 (N11150, N11140, N6251);
nor NOR2 (N11151, N11135, N8673);
or OR2 (N11152, N11147, N3746);
not NOT1 (N11153, N11142);
nand NAND2 (N11154, N11152, N10575);
not NOT1 (N11155, N11151);
not NOT1 (N11156, N11132);
and AND4 (N11157, N11149, N425, N5953, N8996);
nand NAND4 (N11158, N11150, N7821, N9757, N9733);
nand NAND3 (N11159, N11158, N7233, N4046);
nor NOR3 (N11160, N11145, N9183, N5787);
nor NOR3 (N11161, N11156, N4612, N639);
not NOT1 (N11162, N11144);
xor XOR2 (N11163, N11161, N10687);
xor XOR2 (N11164, N11162, N1111);
and AND2 (N11165, N11155, N4641);
buf BUF1 (N11166, N11125);
xor XOR2 (N11167, N11159, N3688);
nand NAND2 (N11168, N11164, N420);
buf BUF1 (N11169, N11168);
nand NAND3 (N11170, N11166, N10932, N8192);
buf BUF1 (N11171, N11165);
nor NOR4 (N11172, N11160, N3744, N5853, N3674);
and AND4 (N11173, N11153, N10951, N7777, N11021);
xor XOR2 (N11174, N11167, N4997);
and AND3 (N11175, N11174, N2857, N6592);
nand NAND2 (N11176, N11173, N5142);
or OR2 (N11177, N11154, N2627);
nor NOR2 (N11178, N11176, N467);
and AND4 (N11179, N11169, N8509, N9214, N7286);
nand NAND3 (N11180, N11175, N8109, N10033);
nand NAND3 (N11181, N11157, N2817, N5036);
not NOT1 (N11182, N11148);
xor XOR2 (N11183, N11170, N4920);
xor XOR2 (N11184, N11163, N7981);
and AND3 (N11185, N11178, N6968, N10581);
buf BUF1 (N11186, N11185);
nor NOR3 (N11187, N11186, N5430, N310);
xor XOR2 (N11188, N11171, N5706);
not NOT1 (N11189, N11181);
nor NOR3 (N11190, N11189, N7597, N5390);
and AND2 (N11191, N11172, N11035);
nor NOR4 (N11192, N11177, N7862, N2380, N773);
and AND4 (N11193, N11191, N4354, N4956, N4663);
buf BUF1 (N11194, N11182);
nand NAND3 (N11195, N11192, N5787, N9896);
nand NAND2 (N11196, N11184, N7740);
xor XOR2 (N11197, N11196, N1323);
and AND3 (N11198, N11194, N1496, N7154);
nor NOR2 (N11199, N11180, N6860);
not NOT1 (N11200, N11193);
buf BUF1 (N11201, N11188);
buf BUF1 (N11202, N11201);
or OR4 (N11203, N11195, N2887, N7356, N1292);
buf BUF1 (N11204, N11198);
not NOT1 (N11205, N11204);
buf BUF1 (N11206, N11199);
and AND3 (N11207, N11203, N1078, N863);
nand NAND2 (N11208, N11190, N7216);
nor NOR3 (N11209, N11208, N11164, N5850);
nand NAND3 (N11210, N11209, N2982, N8900);
buf BUF1 (N11211, N11202);
nand NAND3 (N11212, N11200, N10660, N6182);
nand NAND2 (N11213, N11205, N6332);
nor NOR2 (N11214, N11206, N6457);
nand NAND4 (N11215, N11187, N5714, N7995, N9877);
nor NOR4 (N11216, N11215, N3560, N3765, N5695);
and AND3 (N11217, N11213, N9268, N1135);
xor XOR2 (N11218, N11197, N4577);
or OR4 (N11219, N11218, N6663, N6979, N10882);
or OR2 (N11220, N11212, N3099);
and AND4 (N11221, N11214, N9550, N3927, N3132);
or OR3 (N11222, N11207, N1362, N10409);
and AND4 (N11223, N11222, N364, N236, N4898);
xor XOR2 (N11224, N11220, N3278);
nand NAND3 (N11225, N11219, N2078, N5328);
not NOT1 (N11226, N11216);
xor XOR2 (N11227, N11221, N8552);
and AND4 (N11228, N11227, N8829, N1767, N3190);
or OR2 (N11229, N11224, N8670);
xor XOR2 (N11230, N11211, N2543);
and AND2 (N11231, N11223, N1724);
buf BUF1 (N11232, N11228);
nor NOR3 (N11233, N11179, N44, N2991);
xor XOR2 (N11234, N11225, N9785);
nor NOR3 (N11235, N11210, N11012, N7144);
buf BUF1 (N11236, N11232);
nand NAND4 (N11237, N11236, N1491, N6302, N839);
or OR3 (N11238, N11237, N6585, N4620);
or OR3 (N11239, N11235, N10744, N2435);
xor XOR2 (N11240, N11226, N10111);
nor NOR2 (N11241, N11183, N573);
buf BUF1 (N11242, N11230);
or OR4 (N11243, N11239, N7794, N7337, N309);
or OR3 (N11244, N11241, N10533, N4190);
or OR2 (N11245, N11243, N4925);
nand NAND4 (N11246, N11231, N4707, N6849, N9524);
and AND4 (N11247, N11217, N5232, N2210, N4004);
or OR2 (N11248, N11229, N11125);
or OR2 (N11249, N11240, N10589);
nand NAND2 (N11250, N11245, N3136);
and AND4 (N11251, N11249, N6142, N9403, N2578);
or OR2 (N11252, N11246, N2032);
not NOT1 (N11253, N11242);
or OR4 (N11254, N11250, N866, N4088, N8355);
xor XOR2 (N11255, N11254, N9903);
xor XOR2 (N11256, N11233, N3096);
nor NOR2 (N11257, N11248, N7320);
or OR2 (N11258, N11238, N10668);
nor NOR2 (N11259, N11257, N1802);
nor NOR3 (N11260, N11247, N3258, N1238);
and AND3 (N11261, N11234, N6859, N2934);
nand NAND2 (N11262, N11258, N5520);
nor NOR4 (N11263, N11252, N10596, N297, N1047);
not NOT1 (N11264, N11253);
or OR3 (N11265, N11256, N6862, N5227);
buf BUF1 (N11266, N11259);
or OR2 (N11267, N11260, N7320);
xor XOR2 (N11268, N11265, N704);
buf BUF1 (N11269, N11251);
nand NAND2 (N11270, N11269, N9678);
not NOT1 (N11271, N11267);
nor NOR4 (N11272, N11261, N7772, N6371, N4377);
xor XOR2 (N11273, N11266, N7780);
or OR4 (N11274, N11270, N6317, N2528, N6194);
not NOT1 (N11275, N11274);
and AND2 (N11276, N11275, N2445);
nor NOR3 (N11277, N11271, N6451, N9216);
nand NAND2 (N11278, N11272, N10555);
not NOT1 (N11279, N11264);
and AND4 (N11280, N11278, N6498, N4089, N6986);
nand NAND3 (N11281, N11279, N8873, N9459);
nor NOR2 (N11282, N11263, N5510);
nor NOR2 (N11283, N11281, N6293);
xor XOR2 (N11284, N11273, N3002);
buf BUF1 (N11285, N11284);
nor NOR4 (N11286, N11282, N3090, N9817, N3441);
buf BUF1 (N11287, N11280);
xor XOR2 (N11288, N11255, N5470);
nand NAND4 (N11289, N11277, N8136, N3106, N9238);
buf BUF1 (N11290, N11287);
xor XOR2 (N11291, N11290, N9946);
and AND2 (N11292, N11244, N290);
nor NOR2 (N11293, N11289, N8402);
or OR4 (N11294, N11283, N5645, N8850, N9960);
buf BUF1 (N11295, N11292);
nor NOR3 (N11296, N11285, N3589, N8031);
and AND4 (N11297, N11286, N6611, N1108, N6663);
not NOT1 (N11298, N11268);
nand NAND2 (N11299, N11294, N6532);
or OR3 (N11300, N11299, N2715, N479);
buf BUF1 (N11301, N11288);
and AND3 (N11302, N11295, N7883, N820);
xor XOR2 (N11303, N11262, N8271);
or OR2 (N11304, N11300, N4907);
not NOT1 (N11305, N11293);
or OR2 (N11306, N11305, N9997);
nor NOR4 (N11307, N11304, N4115, N1162, N210);
not NOT1 (N11308, N11302);
or OR2 (N11309, N11276, N6491);
nor NOR2 (N11310, N11306, N1416);
not NOT1 (N11311, N11301);
or OR3 (N11312, N11309, N2215, N1281);
and AND2 (N11313, N11297, N1763);
nand NAND4 (N11314, N11296, N8825, N1184, N1852);
not NOT1 (N11315, N11314);
nand NAND2 (N11316, N11303, N8718);
xor XOR2 (N11317, N11316, N10255);
nor NOR3 (N11318, N11307, N10536, N6766);
and AND2 (N11319, N11308, N8128);
nor NOR4 (N11320, N11317, N10265, N10707, N201);
xor XOR2 (N11321, N11291, N2414);
nor NOR2 (N11322, N11298, N6278);
nor NOR3 (N11323, N11319, N9378, N7322);
not NOT1 (N11324, N11315);
nand NAND2 (N11325, N11312, N7572);
nor NOR2 (N11326, N11321, N1264);
nor NOR3 (N11327, N11310, N1521, N11009);
nor NOR3 (N11328, N11313, N2604, N9477);
xor XOR2 (N11329, N11322, N8561);
not NOT1 (N11330, N11320);
and AND4 (N11331, N11327, N739, N5233, N7454);
nor NOR2 (N11332, N11318, N6147);
buf BUF1 (N11333, N11326);
nand NAND4 (N11334, N11329, N204, N1524, N6790);
buf BUF1 (N11335, N11324);
and AND2 (N11336, N11332, N5079);
nand NAND4 (N11337, N11330, N7963, N9635, N7713);
or OR2 (N11338, N11336, N3578);
nand NAND3 (N11339, N11331, N1108, N9434);
xor XOR2 (N11340, N11328, N9732);
or OR3 (N11341, N11337, N6055, N8181);
not NOT1 (N11342, N11339);
and AND3 (N11343, N11340, N6007, N9235);
xor XOR2 (N11344, N11334, N6812);
xor XOR2 (N11345, N11343, N7165);
and AND4 (N11346, N11338, N731, N3414, N7472);
or OR3 (N11347, N11323, N4201, N2641);
xor XOR2 (N11348, N11333, N10168);
or OR4 (N11349, N11348, N5242, N2169, N8499);
or OR4 (N11350, N11346, N4723, N9810, N1220);
nand NAND3 (N11351, N11325, N1444, N2391);
or OR2 (N11352, N11349, N956);
buf BUF1 (N11353, N11311);
xor XOR2 (N11354, N11335, N2403);
xor XOR2 (N11355, N11341, N6010);
nor NOR4 (N11356, N11347, N11060, N11201, N10501);
nand NAND4 (N11357, N11342, N6146, N7015, N7065);
xor XOR2 (N11358, N11345, N7944);
or OR3 (N11359, N11353, N4925, N4821);
nor NOR2 (N11360, N11354, N5428);
xor XOR2 (N11361, N11352, N147);
and AND2 (N11362, N11351, N6123);
not NOT1 (N11363, N11350);
and AND4 (N11364, N11356, N7323, N8097, N3405);
nor NOR2 (N11365, N11358, N4494);
buf BUF1 (N11366, N11357);
nor NOR2 (N11367, N11365, N9557);
or OR2 (N11368, N11367, N6011);
nor NOR2 (N11369, N11359, N10365);
xor XOR2 (N11370, N11362, N8525);
and AND3 (N11371, N11344, N11084, N1002);
nor NOR3 (N11372, N11368, N10081, N2680);
and AND2 (N11373, N11364, N6640);
or OR3 (N11374, N11371, N9657, N7138);
buf BUF1 (N11375, N11369);
nand NAND4 (N11376, N11373, N9241, N2851, N9827);
and AND4 (N11377, N11363, N9849, N1352, N9599);
or OR4 (N11378, N11366, N6928, N10929, N1637);
not NOT1 (N11379, N11374);
nand NAND2 (N11380, N11375, N1315);
buf BUF1 (N11381, N11370);
nor NOR2 (N11382, N11377, N10436);
and AND4 (N11383, N11376, N6309, N10200, N3317);
not NOT1 (N11384, N11380);
not NOT1 (N11385, N11355);
and AND2 (N11386, N11384, N4366);
or OR4 (N11387, N11385, N7938, N1937, N3579);
and AND3 (N11388, N11372, N8807, N10122);
xor XOR2 (N11389, N11382, N6595);
xor XOR2 (N11390, N11383, N10647);
xor XOR2 (N11391, N11361, N4276);
buf BUF1 (N11392, N11390);
and AND3 (N11393, N11378, N2061, N11001);
not NOT1 (N11394, N11391);
not NOT1 (N11395, N11360);
nand NAND4 (N11396, N11388, N1239, N746, N10890);
and AND4 (N11397, N11393, N9654, N4621, N8917);
xor XOR2 (N11398, N11379, N3851);
and AND3 (N11399, N11398, N8088, N3468);
not NOT1 (N11400, N11392);
or OR4 (N11401, N11396, N3131, N9097, N9277);
and AND3 (N11402, N11399, N8519, N7268);
or OR2 (N11403, N11397, N7356);
not NOT1 (N11404, N11394);
nand NAND4 (N11405, N11381, N6849, N10354, N1040);
or OR2 (N11406, N11402, N1443);
or OR4 (N11407, N11395, N7599, N1789, N9431);
buf BUF1 (N11408, N11403);
nor NOR4 (N11409, N11404, N8050, N9481, N3534);
xor XOR2 (N11410, N11387, N10619);
buf BUF1 (N11411, N11406);
nand NAND4 (N11412, N11410, N11003, N5396, N1010);
buf BUF1 (N11413, N11386);
buf BUF1 (N11414, N11405);
nand NAND2 (N11415, N11409, N6366);
nor NOR3 (N11416, N11413, N8455, N9342);
xor XOR2 (N11417, N11415, N10675);
nand NAND3 (N11418, N11389, N6318, N6739);
xor XOR2 (N11419, N11412, N10362);
nor NOR2 (N11420, N11408, N9039);
and AND2 (N11421, N11407, N5141);
or OR3 (N11422, N11420, N5682, N7173);
and AND3 (N11423, N11401, N159, N550);
buf BUF1 (N11424, N11411);
and AND4 (N11425, N11400, N6020, N6034, N3439);
xor XOR2 (N11426, N11424, N750);
xor XOR2 (N11427, N11417, N9541);
xor XOR2 (N11428, N11425, N1828);
or OR2 (N11429, N11422, N5503);
buf BUF1 (N11430, N11419);
not NOT1 (N11431, N11421);
not NOT1 (N11432, N11418);
buf BUF1 (N11433, N11423);
xor XOR2 (N11434, N11427, N3027);
buf BUF1 (N11435, N11433);
nand NAND4 (N11436, N11431, N4489, N11077, N8828);
nand NAND3 (N11437, N11430, N6254, N6902);
nor NOR2 (N11438, N11432, N2894);
not NOT1 (N11439, N11438);
xor XOR2 (N11440, N11429, N2316);
and AND3 (N11441, N11434, N2790, N9841);
nor NOR4 (N11442, N11435, N1360, N3672, N3093);
buf BUF1 (N11443, N11442);
nor NOR4 (N11444, N11414, N9931, N8210, N2975);
nor NOR2 (N11445, N11443, N8849);
or OR4 (N11446, N11437, N10465, N7429, N5022);
and AND3 (N11447, N11416, N10192, N4226);
buf BUF1 (N11448, N11439);
buf BUF1 (N11449, N11426);
xor XOR2 (N11450, N11440, N3384);
nor NOR4 (N11451, N11447, N3518, N195, N2033);
and AND4 (N11452, N11444, N9292, N8150, N10000);
xor XOR2 (N11453, N11445, N10544);
not NOT1 (N11454, N11448);
and AND3 (N11455, N11436, N3781, N6994);
nor NOR3 (N11456, N11455, N5767, N7456);
xor XOR2 (N11457, N11454, N4578);
or OR4 (N11458, N11457, N8904, N3001, N6240);
nand NAND4 (N11459, N11428, N9145, N5776, N7789);
not NOT1 (N11460, N11452);
or OR3 (N11461, N11446, N3173, N6602);
nor NOR2 (N11462, N11449, N237);
nand NAND4 (N11463, N11461, N7835, N5520, N9237);
or OR3 (N11464, N11441, N5172, N6557);
or OR4 (N11465, N11460, N10663, N6387, N4677);
xor XOR2 (N11466, N11464, N3499);
nor NOR2 (N11467, N11465, N5377);
buf BUF1 (N11468, N11466);
not NOT1 (N11469, N11458);
nor NOR2 (N11470, N11462, N10948);
nand NAND2 (N11471, N11467, N7896);
nand NAND3 (N11472, N11450, N5976, N6626);
buf BUF1 (N11473, N11453);
not NOT1 (N11474, N11473);
not NOT1 (N11475, N11474);
or OR2 (N11476, N11459, N8574);
or OR2 (N11477, N11469, N3035);
nand NAND4 (N11478, N11451, N3678, N8689, N7143);
or OR3 (N11479, N11476, N11220, N9107);
and AND4 (N11480, N11456, N6153, N4908, N2184);
xor XOR2 (N11481, N11471, N259);
buf BUF1 (N11482, N11478);
or OR2 (N11483, N11477, N4116);
xor XOR2 (N11484, N11463, N714);
nand NAND4 (N11485, N11468, N6771, N8784, N2039);
not NOT1 (N11486, N11475);
nand NAND4 (N11487, N11470, N5640, N8762, N2708);
nor NOR4 (N11488, N11480, N5219, N5938, N6185);
nor NOR3 (N11489, N11472, N2931, N7146);
nor NOR4 (N11490, N11488, N340, N7526, N6860);
nand NAND3 (N11491, N11490, N7126, N1746);
nor NOR4 (N11492, N11482, N3912, N7127, N2756);
nand NAND3 (N11493, N11492, N10450, N5785);
and AND3 (N11494, N11487, N3706, N4063);
nor NOR2 (N11495, N11481, N3481);
buf BUF1 (N11496, N11494);
nor NOR2 (N11497, N11485, N9257);
xor XOR2 (N11498, N11489, N723);
or OR3 (N11499, N11479, N8566, N5337);
buf BUF1 (N11500, N11484);
or OR2 (N11501, N11497, N9951);
or OR3 (N11502, N11496, N5544, N814);
buf BUF1 (N11503, N11491);
and AND2 (N11504, N11500, N4615);
buf BUF1 (N11505, N11493);
nor NOR4 (N11506, N11503, N11192, N8036, N4438);
nor NOR2 (N11507, N11495, N6191);
not NOT1 (N11508, N11486);
and AND3 (N11509, N11499, N3531, N9107);
not NOT1 (N11510, N11498);
nor NOR3 (N11511, N11502, N8266, N4792);
and AND3 (N11512, N11510, N4614, N7818);
and AND3 (N11513, N11512, N1916, N320);
not NOT1 (N11514, N11507);
or OR2 (N11515, N11511, N2869);
nor NOR3 (N11516, N11501, N425, N10566);
nor NOR3 (N11517, N11513, N2750, N10193);
nor NOR2 (N11518, N11483, N2611);
xor XOR2 (N11519, N11516, N1641);
or OR2 (N11520, N11506, N741);
and AND3 (N11521, N11515, N6093, N6563);
not NOT1 (N11522, N11508);
xor XOR2 (N11523, N11521, N3658);
and AND3 (N11524, N11522, N3955, N5966);
nor NOR3 (N11525, N11520, N2696, N5894);
nand NAND4 (N11526, N11517, N1381, N9796, N6927);
nand NAND2 (N11527, N11509, N6709);
buf BUF1 (N11528, N11504);
not NOT1 (N11529, N11524);
or OR3 (N11530, N11527, N873, N10558);
nand NAND4 (N11531, N11523, N7329, N5766, N1020);
and AND4 (N11532, N11530, N1306, N11393, N4234);
nand NAND4 (N11533, N11505, N3015, N8231, N1);
nor NOR2 (N11534, N11532, N5790);
nand NAND3 (N11535, N11529, N1164, N2151);
buf BUF1 (N11536, N11533);
nand NAND2 (N11537, N11526, N10167);
nor NOR2 (N11538, N11514, N11222);
buf BUF1 (N11539, N11537);
nand NAND2 (N11540, N11534, N7793);
nor NOR4 (N11541, N11528, N3852, N2713, N8212);
and AND3 (N11542, N11531, N2548, N9320);
and AND2 (N11543, N11538, N11062);
nand NAND4 (N11544, N11518, N3401, N9231, N10838);
nor NOR3 (N11545, N11542, N4581, N857);
nand NAND2 (N11546, N11519, N3528);
nand NAND4 (N11547, N11545, N9861, N9276, N3513);
xor XOR2 (N11548, N11541, N1021);
nand NAND3 (N11549, N11535, N9034, N7399);
buf BUF1 (N11550, N11543);
nand NAND4 (N11551, N11540, N1524, N3347, N3578);
buf BUF1 (N11552, N11549);
buf BUF1 (N11553, N11525);
buf BUF1 (N11554, N11539);
not NOT1 (N11555, N11553);
nor NOR2 (N11556, N11552, N1989);
and AND3 (N11557, N11547, N9903, N4805);
not NOT1 (N11558, N11550);
nor NOR2 (N11559, N11536, N10351);
or OR4 (N11560, N11558, N5531, N8322, N3193);
not NOT1 (N11561, N11557);
nor NOR2 (N11562, N11555, N10985);
nand NAND2 (N11563, N11554, N6301);
nand NAND4 (N11564, N11563, N8901, N398, N6746);
xor XOR2 (N11565, N11548, N7607);
or OR3 (N11566, N11546, N5923, N11420);
nand NAND4 (N11567, N11565, N9570, N7581, N2644);
nor NOR4 (N11568, N11544, N9557, N6270, N5375);
nand NAND2 (N11569, N11562, N3389);
not NOT1 (N11570, N11561);
not NOT1 (N11571, N11566);
xor XOR2 (N11572, N11551, N10064);
nand NAND4 (N11573, N11559, N4573, N3378, N185);
and AND2 (N11574, N11556, N4348);
xor XOR2 (N11575, N11572, N8722);
nand NAND2 (N11576, N11574, N2575);
not NOT1 (N11577, N11569);
buf BUF1 (N11578, N11577);
and AND2 (N11579, N11568, N9212);
or OR3 (N11580, N11576, N10663, N11417);
buf BUF1 (N11581, N11579);
not NOT1 (N11582, N11571);
nand NAND3 (N11583, N11567, N8728, N334);
or OR3 (N11584, N11583, N3259, N10676);
nand NAND2 (N11585, N11570, N8137);
not NOT1 (N11586, N11584);
and AND2 (N11587, N11581, N8200);
or OR4 (N11588, N11580, N5170, N9937, N5937);
nand NAND4 (N11589, N11573, N1118, N2336, N1067);
not NOT1 (N11590, N11560);
xor XOR2 (N11591, N11588, N8655);
and AND2 (N11592, N11586, N9524);
nand NAND2 (N11593, N11564, N2776);
xor XOR2 (N11594, N11590, N2610);
not NOT1 (N11595, N11592);
nand NAND2 (N11596, N11593, N4651);
xor XOR2 (N11597, N11582, N10399);
and AND4 (N11598, N11594, N6726, N9147, N4582);
xor XOR2 (N11599, N11598, N5821);
nand NAND2 (N11600, N11578, N10125);
and AND4 (N11601, N11575, N553, N4693, N6160);
nor NOR2 (N11602, N11599, N5089);
xor XOR2 (N11603, N11596, N5122);
and AND3 (N11604, N11589, N5222, N268);
xor XOR2 (N11605, N11591, N10128);
not NOT1 (N11606, N11595);
xor XOR2 (N11607, N11600, N828);
nand NAND2 (N11608, N11587, N9674);
and AND2 (N11609, N11603, N8455);
not NOT1 (N11610, N11601);
nand NAND4 (N11611, N11609, N1962, N11346, N4149);
nor NOR2 (N11612, N11605, N6747);
not NOT1 (N11613, N11611);
buf BUF1 (N11614, N11610);
nor NOR2 (N11615, N11602, N3982);
not NOT1 (N11616, N11597);
nand NAND4 (N11617, N11616, N6119, N4462, N11005);
xor XOR2 (N11618, N11606, N9700);
buf BUF1 (N11619, N11614);
xor XOR2 (N11620, N11604, N4192);
and AND2 (N11621, N11607, N10809);
xor XOR2 (N11622, N11620, N2017);
nor NOR4 (N11623, N11621, N8148, N1528, N5508);
nand NAND4 (N11624, N11585, N2872, N9863, N9613);
nor NOR3 (N11625, N11613, N10595, N1534);
nor NOR4 (N11626, N11623, N4773, N8235, N5300);
xor XOR2 (N11627, N11618, N2492);
xor XOR2 (N11628, N11624, N94);
xor XOR2 (N11629, N11615, N3364);
nor NOR2 (N11630, N11612, N6633);
and AND2 (N11631, N11629, N10520);
or OR2 (N11632, N11625, N6542);
nor NOR4 (N11633, N11617, N582, N10820, N11020);
and AND4 (N11634, N11622, N5795, N6471, N722);
xor XOR2 (N11635, N11626, N1086);
or OR2 (N11636, N11634, N1005);
and AND2 (N11637, N11628, N2061);
and AND4 (N11638, N11627, N1810, N686, N1434);
buf BUF1 (N11639, N11635);
not NOT1 (N11640, N11633);
buf BUF1 (N11641, N11638);
or OR2 (N11642, N11619, N5425);
xor XOR2 (N11643, N11641, N8763);
nand NAND2 (N11644, N11643, N4196);
not NOT1 (N11645, N11640);
buf BUF1 (N11646, N11642);
and AND2 (N11647, N11636, N2972);
or OR3 (N11648, N11646, N8959, N11459);
nand NAND2 (N11649, N11632, N2340);
or OR3 (N11650, N11648, N10957, N3856);
and AND2 (N11651, N11637, N10532);
buf BUF1 (N11652, N11639);
not NOT1 (N11653, N11644);
and AND2 (N11654, N11653, N1539);
xor XOR2 (N11655, N11650, N1246);
not NOT1 (N11656, N11655);
nor NOR4 (N11657, N11608, N9069, N9634, N3028);
not NOT1 (N11658, N11656);
buf BUF1 (N11659, N11652);
xor XOR2 (N11660, N11657, N1154);
not NOT1 (N11661, N11645);
nand NAND4 (N11662, N11661, N5886, N2707, N7900);
nand NAND3 (N11663, N11662, N1841, N2129);
or OR4 (N11664, N11663, N2960, N7957, N2857);
xor XOR2 (N11665, N11651, N9156);
xor XOR2 (N11666, N11647, N4197);
and AND3 (N11667, N11665, N2808, N10207);
xor XOR2 (N11668, N11658, N6637);
nand NAND3 (N11669, N11654, N7754, N1878);
not NOT1 (N11670, N11669);
buf BUF1 (N11671, N11664);
buf BUF1 (N11672, N11630);
xor XOR2 (N11673, N11666, N3893);
and AND3 (N11674, N11670, N7739, N26);
buf BUF1 (N11675, N11672);
and AND2 (N11676, N11649, N9415);
nand NAND3 (N11677, N11675, N224, N5392);
buf BUF1 (N11678, N11668);
not NOT1 (N11679, N11677);
and AND3 (N11680, N11673, N7224, N4033);
nand NAND3 (N11681, N11679, N4530, N5718);
buf BUF1 (N11682, N11681);
and AND2 (N11683, N11660, N3213);
nand NAND4 (N11684, N11659, N3195, N434, N4483);
nand NAND2 (N11685, N11683, N8347);
nand NAND3 (N11686, N11682, N9728, N7420);
and AND3 (N11687, N11678, N1259, N11237);
buf BUF1 (N11688, N11676);
and AND3 (N11689, N11680, N7436, N5841);
nor NOR4 (N11690, N11689, N8765, N6129, N3528);
not NOT1 (N11691, N11687);
and AND4 (N11692, N11684, N7091, N4133, N8419);
and AND4 (N11693, N11671, N4651, N468, N5042);
buf BUF1 (N11694, N11686);
nand NAND3 (N11695, N11693, N753, N8635);
not NOT1 (N11696, N11690);
xor XOR2 (N11697, N11695, N670);
nor NOR2 (N11698, N11667, N9400);
buf BUF1 (N11699, N11698);
nand NAND2 (N11700, N11692, N7524);
and AND2 (N11701, N11700, N1966);
nand NAND2 (N11702, N11694, N9420);
xor XOR2 (N11703, N11691, N424);
buf BUF1 (N11704, N11701);
buf BUF1 (N11705, N11702);
xor XOR2 (N11706, N11631, N9218);
and AND3 (N11707, N11705, N2145, N6497);
and AND2 (N11708, N11688, N6091);
or OR2 (N11709, N11708, N4527);
nand NAND4 (N11710, N11709, N5248, N287, N10044);
nand NAND2 (N11711, N11696, N149);
nor NOR4 (N11712, N11711, N367, N9813, N5145);
nand NAND4 (N11713, N11706, N6470, N4296, N11207);
nand NAND4 (N11714, N11703, N6998, N132, N3228);
or OR4 (N11715, N11712, N8534, N4398, N8583);
not NOT1 (N11716, N11697);
xor XOR2 (N11717, N11716, N3864);
and AND3 (N11718, N11714, N3224, N4361);
not NOT1 (N11719, N11718);
not NOT1 (N11720, N11715);
and AND2 (N11721, N11713, N9140);
and AND3 (N11722, N11717, N944, N6421);
nor NOR2 (N11723, N11707, N1008);
and AND4 (N11724, N11720, N2471, N7813, N6161);
not NOT1 (N11725, N11704);
nand NAND3 (N11726, N11699, N7669, N185);
and AND2 (N11727, N11674, N154);
xor XOR2 (N11728, N11726, N10445);
and AND4 (N11729, N11685, N6780, N6547, N7818);
buf BUF1 (N11730, N11722);
buf BUF1 (N11731, N11723);
or OR2 (N11732, N11730, N1576);
xor XOR2 (N11733, N11731, N1209);
and AND2 (N11734, N11727, N6415);
not NOT1 (N11735, N11729);
and AND2 (N11736, N11724, N3023);
nand NAND4 (N11737, N11710, N1200, N10036, N7900);
nand NAND2 (N11738, N11736, N4740);
or OR2 (N11739, N11721, N2275);
not NOT1 (N11740, N11732);
not NOT1 (N11741, N11733);
xor XOR2 (N11742, N11740, N7860);
xor XOR2 (N11743, N11734, N5934);
nor NOR4 (N11744, N11741, N10015, N6246, N10524);
and AND4 (N11745, N11738, N1887, N6845, N11613);
xor XOR2 (N11746, N11742, N7531);
and AND2 (N11747, N11745, N2329);
xor XOR2 (N11748, N11744, N3223);
not NOT1 (N11749, N11719);
nand NAND4 (N11750, N11728, N11669, N11745, N4841);
not NOT1 (N11751, N11735);
buf BUF1 (N11752, N11725);
xor XOR2 (N11753, N11750, N7067);
nand NAND4 (N11754, N11752, N4711, N9778, N5012);
not NOT1 (N11755, N11753);
nand NAND3 (N11756, N11747, N11395, N6154);
nor NOR4 (N11757, N11737, N6681, N470, N11748);
and AND2 (N11758, N4365, N9602);
nand NAND2 (N11759, N11758, N810);
not NOT1 (N11760, N11755);
not NOT1 (N11761, N11743);
or OR3 (N11762, N11759, N5303, N8378);
or OR3 (N11763, N11746, N6644, N3885);
nand NAND4 (N11764, N11757, N7903, N8528, N2171);
xor XOR2 (N11765, N11764, N11248);
not NOT1 (N11766, N11760);
and AND2 (N11767, N11765, N4519);
and AND4 (N11768, N11767, N171, N9990, N8212);
xor XOR2 (N11769, N11739, N620);
or OR2 (N11770, N11761, N10941);
and AND4 (N11771, N11770, N5194, N9783, N10974);
buf BUF1 (N11772, N11754);
nor NOR2 (N11773, N11749, N7835);
nand NAND3 (N11774, N11771, N7281, N7222);
not NOT1 (N11775, N11762);
not NOT1 (N11776, N11766);
and AND2 (N11777, N11751, N2023);
not NOT1 (N11778, N11776);
or OR4 (N11779, N11774, N1228, N1335, N251);
buf BUF1 (N11780, N11756);
nand NAND3 (N11781, N11780, N5530, N3263);
xor XOR2 (N11782, N11769, N5925);
and AND3 (N11783, N11775, N2182, N8905);
or OR2 (N11784, N11772, N4214);
and AND2 (N11785, N11784, N3266);
nand NAND3 (N11786, N11768, N850, N3156);
and AND2 (N11787, N11783, N4543);
and AND4 (N11788, N11782, N3975, N4273, N2061);
nand NAND3 (N11789, N11785, N6219, N1982);
nand NAND4 (N11790, N11781, N4249, N6920, N9548);
and AND3 (N11791, N11786, N9842, N6199);
not NOT1 (N11792, N11788);
buf BUF1 (N11793, N11779);
not NOT1 (N11794, N11777);
nand NAND4 (N11795, N11793, N10061, N6917, N182);
xor XOR2 (N11796, N11778, N10338);
and AND3 (N11797, N11791, N8416, N6620);
or OR4 (N11798, N11763, N10953, N11603, N5711);
nor NOR3 (N11799, N11789, N9696, N5728);
buf BUF1 (N11800, N11799);
or OR3 (N11801, N11794, N2547, N6685);
not NOT1 (N11802, N11801);
xor XOR2 (N11803, N11797, N9983);
nand NAND4 (N11804, N11795, N3921, N11397, N6967);
nor NOR4 (N11805, N11792, N5300, N11404, N6621);
and AND4 (N11806, N11805, N7963, N9192, N10117);
not NOT1 (N11807, N11802);
nand NAND2 (N11808, N11787, N2925);
not NOT1 (N11809, N11804);
nor NOR3 (N11810, N11773, N949, N4705);
nor NOR4 (N11811, N11796, N4598, N10480, N1933);
or OR4 (N11812, N11806, N11171, N3826, N3379);
nand NAND2 (N11813, N11812, N11506);
xor XOR2 (N11814, N11811, N2924);
nand NAND4 (N11815, N11807, N7822, N6719, N11032);
not NOT1 (N11816, N11814);
or OR3 (N11817, N11800, N10556, N8096);
buf BUF1 (N11818, N11813);
nand NAND2 (N11819, N11818, N3823);
or OR4 (N11820, N11790, N8891, N2303, N1733);
and AND2 (N11821, N11816, N8709);
and AND4 (N11822, N11821, N11369, N5240, N184);
and AND3 (N11823, N11815, N7212, N11154);
and AND3 (N11824, N11823, N91, N6545);
nor NOR2 (N11825, N11810, N7507);
nand NAND4 (N11826, N11798, N8731, N330, N3246);
nor NOR3 (N11827, N11826, N4337, N2254);
nand NAND4 (N11828, N11820, N11192, N429, N5044);
xor XOR2 (N11829, N11825, N6264);
nand NAND2 (N11830, N11824, N11708);
buf BUF1 (N11831, N11819);
and AND3 (N11832, N11830, N504, N7533);
nand NAND3 (N11833, N11808, N8004, N4620);
not NOT1 (N11834, N11828);
nor NOR4 (N11835, N11803, N11483, N10489, N5812);
and AND4 (N11836, N11832, N11590, N1969, N1393);
xor XOR2 (N11837, N11822, N4623);
buf BUF1 (N11838, N11831);
nor NOR4 (N11839, N11835, N2328, N11683, N5858);
xor XOR2 (N11840, N11837, N7797);
nor NOR4 (N11841, N11833, N2565, N7890, N10342);
nor NOR3 (N11842, N11809, N2022, N5769);
buf BUF1 (N11843, N11842);
not NOT1 (N11844, N11840);
and AND3 (N11845, N11827, N7974, N7613);
not NOT1 (N11846, N11841);
xor XOR2 (N11847, N11843, N2774);
nand NAND2 (N11848, N11839, N9451);
xor XOR2 (N11849, N11834, N11113);
buf BUF1 (N11850, N11836);
nor NOR3 (N11851, N11846, N4941, N9279);
and AND3 (N11852, N11817, N5854, N2704);
buf BUF1 (N11853, N11851);
nor NOR3 (N11854, N11844, N6917, N610);
buf BUF1 (N11855, N11850);
xor XOR2 (N11856, N11838, N9267);
nand NAND3 (N11857, N11852, N1935, N1211);
or OR4 (N11858, N11847, N9224, N8064, N8321);
or OR4 (N11859, N11849, N7578, N4631, N4507);
buf BUF1 (N11860, N11853);
nand NAND3 (N11861, N11855, N5408, N9730);
or OR4 (N11862, N11845, N5518, N1089, N11201);
nand NAND4 (N11863, N11862, N6378, N10829, N7158);
xor XOR2 (N11864, N11860, N5134);
not NOT1 (N11865, N11829);
not NOT1 (N11866, N11859);
and AND4 (N11867, N11866, N5399, N1817, N110);
nor NOR4 (N11868, N11863, N8490, N8905, N909);
nor NOR2 (N11869, N11857, N9884);
nor NOR2 (N11870, N11867, N10354);
nand NAND4 (N11871, N11865, N8416, N7277, N2498);
not NOT1 (N11872, N11870);
nand NAND3 (N11873, N11872, N2912, N2234);
nor NOR4 (N11874, N11864, N11527, N5861, N4574);
nor NOR2 (N11875, N11869, N1649);
not NOT1 (N11876, N11875);
or OR2 (N11877, N11871, N9275);
buf BUF1 (N11878, N11848);
xor XOR2 (N11879, N11858, N11763);
and AND2 (N11880, N11878, N4852);
nor NOR2 (N11881, N11856, N3132);
xor XOR2 (N11882, N11880, N11274);
buf BUF1 (N11883, N11881);
and AND3 (N11884, N11879, N6604, N11482);
and AND4 (N11885, N11876, N3889, N2642, N11120);
nor NOR4 (N11886, N11883, N9776, N5112, N10337);
xor XOR2 (N11887, N11884, N2558);
xor XOR2 (N11888, N11885, N9864);
nand NAND4 (N11889, N11886, N2724, N2834, N11755);
xor XOR2 (N11890, N11861, N9705);
and AND4 (N11891, N11888, N5887, N6554, N6202);
or OR3 (N11892, N11874, N9503, N1959);
and AND3 (N11893, N11882, N3291, N1567);
and AND4 (N11894, N11891, N5224, N7111, N9619);
or OR4 (N11895, N11892, N385, N4172, N7993);
xor XOR2 (N11896, N11895, N3165);
nand NAND4 (N11897, N11896, N1586, N8743, N5900);
or OR3 (N11898, N11889, N10116, N1110);
and AND3 (N11899, N11893, N8764, N4675);
or OR3 (N11900, N11854, N10652, N4667);
and AND2 (N11901, N11900, N7221);
and AND4 (N11902, N11873, N9322, N7159, N3054);
or OR2 (N11903, N11897, N1271);
xor XOR2 (N11904, N11877, N9994);
and AND3 (N11905, N11868, N3374, N11589);
or OR3 (N11906, N11905, N10465, N7154);
buf BUF1 (N11907, N11898);
and AND3 (N11908, N11902, N11884, N1882);
nor NOR4 (N11909, N11904, N11322, N10020, N5108);
nand NAND4 (N11910, N11908, N5811, N9324, N8684);
or OR4 (N11911, N11910, N1534, N11139, N2407);
or OR4 (N11912, N11887, N1864, N3389, N90);
buf BUF1 (N11913, N11903);
nand NAND3 (N11914, N11912, N6108, N8061);
and AND3 (N11915, N11899, N5369, N538);
nand NAND2 (N11916, N11907, N3818);
or OR3 (N11917, N11911, N10168, N9683);
xor XOR2 (N11918, N11913, N11545);
nor NOR3 (N11919, N11894, N10437, N10623);
or OR2 (N11920, N11914, N3868);
buf BUF1 (N11921, N11918);
not NOT1 (N11922, N11890);
nand NAND4 (N11923, N11919, N8327, N10031, N9658);
and AND2 (N11924, N11909, N8811);
nor NOR2 (N11925, N11917, N8368);
not NOT1 (N11926, N11906);
buf BUF1 (N11927, N11924);
buf BUF1 (N11928, N11921);
xor XOR2 (N11929, N11920, N9547);
nand NAND3 (N11930, N11923, N6742, N380);
buf BUF1 (N11931, N11930);
or OR2 (N11932, N11916, N9680);
nor NOR3 (N11933, N11915, N8215, N4304);
buf BUF1 (N11934, N11932);
buf BUF1 (N11935, N11928);
xor XOR2 (N11936, N11934, N5622);
xor XOR2 (N11937, N11901, N7315);
nand NAND2 (N11938, N11927, N1340);
buf BUF1 (N11939, N11937);
buf BUF1 (N11940, N11925);
or OR4 (N11941, N11922, N11801, N10598, N665);
or OR2 (N11942, N11940, N5388);
not NOT1 (N11943, N11929);
or OR3 (N11944, N11938, N11324, N10383);
not NOT1 (N11945, N11936);
not NOT1 (N11946, N11935);
not NOT1 (N11947, N11944);
buf BUF1 (N11948, N11947);
nor NOR3 (N11949, N11939, N5224, N11472);
not NOT1 (N11950, N11941);
nand NAND2 (N11951, N11945, N3869);
nor NOR4 (N11952, N11926, N3621, N9570, N10731);
buf BUF1 (N11953, N11952);
or OR4 (N11954, N11951, N1987, N722, N9605);
not NOT1 (N11955, N11946);
and AND2 (N11956, N11949, N3165);
and AND4 (N11957, N11931, N2058, N3938, N2571);
or OR2 (N11958, N11953, N3573);
xor XOR2 (N11959, N11958, N6045);
buf BUF1 (N11960, N11942);
or OR4 (N11961, N11948, N7641, N4004, N9690);
xor XOR2 (N11962, N11961, N1918);
and AND4 (N11963, N11950, N905, N11321, N3680);
buf BUF1 (N11964, N11960);
buf BUF1 (N11965, N11943);
and AND2 (N11966, N11963, N6908);
xor XOR2 (N11967, N11962, N8270);
not NOT1 (N11968, N11966);
nand NAND4 (N11969, N11955, N11570, N4194, N7817);
nor NOR3 (N11970, N11959, N1273, N8527);
buf BUF1 (N11971, N11969);
nand NAND3 (N11972, N11970, N10394, N10821);
not NOT1 (N11973, N11933);
nor NOR3 (N11974, N11968, N6468, N8609);
xor XOR2 (N11975, N11964, N7852);
and AND3 (N11976, N11967, N9477, N5369);
buf BUF1 (N11977, N11973);
not NOT1 (N11978, N11974);
or OR2 (N11979, N11965, N7952);
xor XOR2 (N11980, N11977, N4707);
buf BUF1 (N11981, N11972);
xor XOR2 (N11982, N11976, N1165);
nor NOR3 (N11983, N11980, N2326, N714);
nand NAND2 (N11984, N11957, N3985);
or OR3 (N11985, N11956, N3090, N3142);
buf BUF1 (N11986, N11954);
and AND2 (N11987, N11978, N4025);
xor XOR2 (N11988, N11975, N11722);
xor XOR2 (N11989, N11985, N8117);
not NOT1 (N11990, N11971);
or OR3 (N11991, N11982, N307, N8422);
not NOT1 (N11992, N11990);
or OR2 (N11993, N11986, N209);
or OR3 (N11994, N11993, N3023, N6408);
or OR2 (N11995, N11984, N8141);
and AND2 (N11996, N11992, N1481);
nand NAND4 (N11997, N11991, N3672, N10164, N1407);
nand NAND4 (N11998, N11994, N10356, N11058, N6438);
or OR3 (N11999, N11989, N8607, N6763);
nor NOR4 (N12000, N11988, N11964, N5136, N7799);
not NOT1 (N12001, N12000);
nor NOR2 (N12002, N11987, N7624);
not NOT1 (N12003, N12002);
xor XOR2 (N12004, N11999, N2318);
nor NOR4 (N12005, N11983, N11135, N8824, N7894);
not NOT1 (N12006, N12004);
nor NOR4 (N12007, N11997, N2637, N9989, N9561);
and AND4 (N12008, N12003, N8979, N1643, N1489);
and AND3 (N12009, N11981, N9750, N9130);
or OR4 (N12010, N12006, N2254, N4688, N10055);
xor XOR2 (N12011, N12008, N9942);
or OR2 (N12012, N12009, N11674);
xor XOR2 (N12013, N11998, N797);
not NOT1 (N12014, N11996);
or OR3 (N12015, N12001, N1360, N9247);
xor XOR2 (N12016, N12010, N2055);
and AND3 (N12017, N12012, N11612, N8857);
not NOT1 (N12018, N12016);
buf BUF1 (N12019, N12013);
xor XOR2 (N12020, N12007, N2599);
not NOT1 (N12021, N12019);
nand NAND2 (N12022, N12021, N2253);
nor NOR3 (N12023, N12018, N9261, N9595);
and AND2 (N12024, N12023, N4908);
and AND3 (N12025, N12015, N11699, N10323);
not NOT1 (N12026, N12005);
buf BUF1 (N12027, N12011);
nor NOR2 (N12028, N12025, N3319);
xor XOR2 (N12029, N12020, N470);
buf BUF1 (N12030, N12022);
xor XOR2 (N12031, N12027, N6745);
nor NOR2 (N12032, N11995, N8398);
not NOT1 (N12033, N12032);
nand NAND4 (N12034, N12031, N8405, N1017, N339);
xor XOR2 (N12035, N12033, N2868);
buf BUF1 (N12036, N12034);
buf BUF1 (N12037, N12029);
not NOT1 (N12038, N12014);
nand NAND4 (N12039, N12030, N8941, N7381, N5688);
buf BUF1 (N12040, N12037);
nor NOR4 (N12041, N12036, N3598, N1476, N9370);
xor XOR2 (N12042, N12038, N8871);
xor XOR2 (N12043, N12035, N10664);
and AND2 (N12044, N12024, N7278);
nand NAND4 (N12045, N12039, N9194, N9925, N10745);
nor NOR2 (N12046, N12044, N11152);
buf BUF1 (N12047, N12017);
xor XOR2 (N12048, N12047, N7142);
buf BUF1 (N12049, N12043);
nor NOR4 (N12050, N12041, N8515, N3194, N1670);
not NOT1 (N12051, N12045);
xor XOR2 (N12052, N11979, N7153);
or OR4 (N12053, N12042, N4926, N3389, N6563);
buf BUF1 (N12054, N12046);
and AND3 (N12055, N12050, N7207, N1436);
or OR4 (N12056, N12054, N7542, N5458, N2466);
nand NAND3 (N12057, N12048, N5593, N3690);
nor NOR4 (N12058, N12053, N852, N4164, N9810);
not NOT1 (N12059, N12051);
nor NOR4 (N12060, N12052, N4468, N4769, N6482);
not NOT1 (N12061, N12059);
nand NAND2 (N12062, N12058, N2610);
nor NOR4 (N12063, N12055, N8394, N8110, N4690);
and AND2 (N12064, N12026, N3162);
xor XOR2 (N12065, N12063, N773);
xor XOR2 (N12066, N12057, N9752);
not NOT1 (N12067, N12028);
nor NOR2 (N12068, N12060, N6511);
not NOT1 (N12069, N12062);
or OR4 (N12070, N12068, N8114, N11497, N1028);
xor XOR2 (N12071, N12064, N10462);
or OR2 (N12072, N12071, N2595);
and AND3 (N12073, N12056, N4905, N9733);
or OR4 (N12074, N12040, N11224, N1280, N10215);
not NOT1 (N12075, N12066);
and AND2 (N12076, N12049, N3708);
xor XOR2 (N12077, N12067, N626);
nor NOR2 (N12078, N12061, N9964);
not NOT1 (N12079, N12078);
xor XOR2 (N12080, N12072, N4951);
or OR4 (N12081, N12080, N11859, N6917, N4332);
nand NAND3 (N12082, N12073, N10903, N10241);
xor XOR2 (N12083, N12074, N399);
or OR4 (N12084, N12076, N4193, N313, N10429);
not NOT1 (N12085, N12065);
or OR4 (N12086, N12082, N7283, N2062, N4315);
or OR4 (N12087, N12079, N3376, N11450, N11719);
or OR2 (N12088, N12077, N2973);
xor XOR2 (N12089, N12075, N4043);
xor XOR2 (N12090, N12081, N3629);
and AND2 (N12091, N12088, N1147);
and AND2 (N12092, N12069, N12078);
xor XOR2 (N12093, N12087, N11947);
buf BUF1 (N12094, N12070);
nand NAND2 (N12095, N12093, N8941);
buf BUF1 (N12096, N12086);
xor XOR2 (N12097, N12090, N2220);
nand NAND2 (N12098, N12089, N6616);
not NOT1 (N12099, N12084);
nor NOR4 (N12100, N12092, N406, N1529, N3671);
xor XOR2 (N12101, N12094, N5957);
xor XOR2 (N12102, N12096, N6512);
not NOT1 (N12103, N12100);
buf BUF1 (N12104, N12097);
xor XOR2 (N12105, N12103, N1768);
and AND4 (N12106, N12083, N9554, N2281, N169);
nand NAND2 (N12107, N12099, N9087);
nor NOR3 (N12108, N12095, N10347, N11561);
and AND4 (N12109, N12104, N7060, N11780, N4097);
and AND2 (N12110, N12109, N2510);
or OR2 (N12111, N12101, N8392);
not NOT1 (N12112, N12102);
nor NOR2 (N12113, N12085, N5897);
nand NAND3 (N12114, N12111, N7835, N9116);
xor XOR2 (N12115, N12107, N8295);
not NOT1 (N12116, N12112);
nor NOR2 (N12117, N12108, N7158);
nand NAND3 (N12118, N12115, N1580, N793);
and AND2 (N12119, N12091, N8592);
and AND3 (N12120, N12106, N11515, N5309);
not NOT1 (N12121, N12114);
not NOT1 (N12122, N12116);
buf BUF1 (N12123, N12121);
nor NOR2 (N12124, N12113, N1668);
buf BUF1 (N12125, N12124);
nor NOR2 (N12126, N12120, N160);
xor XOR2 (N12127, N12117, N11936);
not NOT1 (N12128, N12098);
or OR4 (N12129, N12119, N72, N1268, N11997);
or OR2 (N12130, N12129, N11994);
not NOT1 (N12131, N12118);
nor NOR3 (N12132, N12130, N2990, N10077);
xor XOR2 (N12133, N12123, N6059);
or OR2 (N12134, N12122, N8494);
nand NAND2 (N12135, N12132, N7332);
buf BUF1 (N12136, N12131);
or OR4 (N12137, N12110, N11957, N11987, N5861);
nor NOR4 (N12138, N12135, N8530, N7317, N6172);
xor XOR2 (N12139, N12128, N9223);
nor NOR3 (N12140, N12136, N5495, N6110);
xor XOR2 (N12141, N12125, N7665);
xor XOR2 (N12142, N12141, N6221);
or OR3 (N12143, N12138, N5130, N6706);
or OR4 (N12144, N12140, N3429, N2863, N9076);
or OR3 (N12145, N12133, N1521, N4578);
or OR2 (N12146, N12126, N7281);
and AND2 (N12147, N12127, N10841);
or OR4 (N12148, N12137, N2065, N8495, N10527);
and AND2 (N12149, N12105, N2790);
xor XOR2 (N12150, N12139, N8351);
nor NOR4 (N12151, N12149, N12048, N651, N422);
not NOT1 (N12152, N12142);
or OR3 (N12153, N12143, N10325, N10212);
nand NAND4 (N12154, N12147, N11622, N10154, N6041);
nand NAND4 (N12155, N12153, N7166, N5784, N5038);
nand NAND4 (N12156, N12148, N11547, N6973, N1652);
or OR4 (N12157, N12152, N3453, N1037, N904);
buf BUF1 (N12158, N12156);
not NOT1 (N12159, N12157);
buf BUF1 (N12160, N12145);
xor XOR2 (N12161, N12146, N11698);
not NOT1 (N12162, N12154);
and AND2 (N12163, N12158, N9332);
buf BUF1 (N12164, N12161);
and AND2 (N12165, N12155, N7920);
or OR4 (N12166, N12150, N46, N10830, N3368);
or OR2 (N12167, N12162, N7680);
or OR3 (N12168, N12164, N741, N10015);
or OR2 (N12169, N12160, N7168);
xor XOR2 (N12170, N12134, N5368);
and AND4 (N12171, N12169, N2795, N7286, N9516);
buf BUF1 (N12172, N12163);
xor XOR2 (N12173, N12165, N3805);
nor NOR2 (N12174, N12166, N9008);
xor XOR2 (N12175, N12159, N8288);
or OR3 (N12176, N12173, N8503, N4223);
not NOT1 (N12177, N12172);
xor XOR2 (N12178, N12175, N1307);
nand NAND2 (N12179, N12178, N4681);
nand NAND4 (N12180, N12167, N8554, N800, N10652);
not NOT1 (N12181, N12171);
nor NOR3 (N12182, N12180, N6274, N6691);
or OR2 (N12183, N12177, N1919);
not NOT1 (N12184, N12181);
or OR3 (N12185, N12144, N2396, N10702);
or OR2 (N12186, N12174, N8139);
and AND4 (N12187, N12184, N4698, N83, N10228);
not NOT1 (N12188, N12151);
buf BUF1 (N12189, N12185);
not NOT1 (N12190, N12176);
buf BUF1 (N12191, N12189);
and AND4 (N12192, N12191, N11046, N1622, N4183);
not NOT1 (N12193, N12183);
nor NOR3 (N12194, N12182, N8590, N3445);
nand NAND2 (N12195, N12190, N4969);
nor NOR4 (N12196, N12187, N6132, N1979, N11291);
buf BUF1 (N12197, N12168);
xor XOR2 (N12198, N12195, N5598);
buf BUF1 (N12199, N12197);
not NOT1 (N12200, N12170);
nand NAND4 (N12201, N12186, N8917, N2126, N10282);
nor NOR3 (N12202, N12198, N5326, N9847);
not NOT1 (N12203, N12179);
not NOT1 (N12204, N12193);
not NOT1 (N12205, N12192);
nand NAND4 (N12206, N12205, N7465, N8266, N3892);
not NOT1 (N12207, N12203);
buf BUF1 (N12208, N12200);
nand NAND2 (N12209, N12202, N1173);
and AND2 (N12210, N12196, N1482);
nand NAND2 (N12211, N12208, N369);
xor XOR2 (N12212, N12206, N2958);
nand NAND2 (N12213, N12207, N10838);
buf BUF1 (N12214, N12194);
nor NOR4 (N12215, N12201, N3002, N6651, N6875);
xor XOR2 (N12216, N12210, N432);
nand NAND4 (N12217, N12204, N8889, N2434, N8464);
and AND4 (N12218, N12199, N4355, N10251, N3675);
nor NOR4 (N12219, N12216, N6346, N2845, N4237);
not NOT1 (N12220, N12213);
or OR3 (N12221, N12211, N11799, N8640);
and AND4 (N12222, N12219, N6918, N9653, N11909);
nor NOR2 (N12223, N12209, N3772);
and AND4 (N12224, N12222, N6060, N10856, N3200);
nand NAND4 (N12225, N12221, N7179, N11789, N6768);
nand NAND2 (N12226, N12218, N11198);
nand NAND4 (N12227, N12214, N4365, N10492, N9759);
not NOT1 (N12228, N12212);
nand NAND2 (N12229, N12227, N6840);
and AND3 (N12230, N12188, N12155, N3496);
nand NAND2 (N12231, N12224, N6833);
not NOT1 (N12232, N12225);
and AND2 (N12233, N12226, N6375);
nand NAND2 (N12234, N12228, N10322);
nor NOR4 (N12235, N12215, N9752, N41, N8860);
nand NAND4 (N12236, N12217, N2513, N6413, N5802);
buf BUF1 (N12237, N12229);
nand NAND3 (N12238, N12232, N6466, N6252);
nand NAND2 (N12239, N12238, N9747);
nor NOR2 (N12240, N12236, N1070);
or OR3 (N12241, N12223, N9855, N8993);
xor XOR2 (N12242, N12239, N6799);
xor XOR2 (N12243, N12237, N7494);
xor XOR2 (N12244, N12220, N10789);
not NOT1 (N12245, N12243);
and AND3 (N12246, N12233, N11577, N12057);
xor XOR2 (N12247, N12241, N4805);
not NOT1 (N12248, N12234);
buf BUF1 (N12249, N12230);
xor XOR2 (N12250, N12240, N1114);
xor XOR2 (N12251, N12245, N9561);
xor XOR2 (N12252, N12247, N11155);
xor XOR2 (N12253, N12246, N2130);
xor XOR2 (N12254, N12244, N8632);
not NOT1 (N12255, N12248);
not NOT1 (N12256, N12242);
and AND2 (N12257, N12231, N3911);
and AND4 (N12258, N12253, N801, N2192, N3309);
and AND4 (N12259, N12249, N5027, N525, N12166);
and AND4 (N12260, N12235, N3640, N10152, N12190);
not NOT1 (N12261, N12258);
nor NOR4 (N12262, N12259, N8145, N12025, N9814);
buf BUF1 (N12263, N12257);
or OR3 (N12264, N12250, N8225, N1089);
and AND4 (N12265, N12256, N1346, N11542, N7194);
nor NOR4 (N12266, N12262, N2923, N4804, N12016);
nand NAND2 (N12267, N12264, N9862);
nor NOR2 (N12268, N12267, N8616);
not NOT1 (N12269, N12265);
or OR4 (N12270, N12255, N1932, N1750, N3134);
nand NAND3 (N12271, N12251, N1673, N4909);
not NOT1 (N12272, N12270);
not NOT1 (N12273, N12260);
and AND3 (N12274, N12252, N9823, N6567);
not NOT1 (N12275, N12268);
or OR4 (N12276, N12273, N8054, N6479, N890);
buf BUF1 (N12277, N12272);
nand NAND3 (N12278, N12254, N1268, N6934);
buf BUF1 (N12279, N12266);
buf BUF1 (N12280, N12275);
and AND3 (N12281, N12280, N3509, N1860);
nor NOR2 (N12282, N12277, N2277);
or OR2 (N12283, N12279, N2610);
nor NOR3 (N12284, N12278, N8583, N6309);
xor XOR2 (N12285, N12274, N8688);
not NOT1 (N12286, N12263);
nand NAND4 (N12287, N12285, N1773, N11492, N3911);
buf BUF1 (N12288, N12271);
xor XOR2 (N12289, N12281, N243);
nand NAND4 (N12290, N12287, N563, N9640, N7569);
and AND3 (N12291, N12290, N1242, N6615);
buf BUF1 (N12292, N12286);
xor XOR2 (N12293, N12291, N2042);
nand NAND4 (N12294, N12261, N6630, N8226, N9236);
xor XOR2 (N12295, N12294, N6624);
nor NOR4 (N12296, N12269, N10676, N4403, N8614);
nand NAND2 (N12297, N12289, N2147);
xor XOR2 (N12298, N12288, N10237);
and AND2 (N12299, N12284, N3205);
not NOT1 (N12300, N12283);
and AND4 (N12301, N12293, N7037, N9550, N5047);
not NOT1 (N12302, N12300);
or OR2 (N12303, N12282, N11787);
buf BUF1 (N12304, N12301);
and AND2 (N12305, N12296, N9118);
buf BUF1 (N12306, N12302);
xor XOR2 (N12307, N12305, N8664);
buf BUF1 (N12308, N12292);
buf BUF1 (N12309, N12295);
xor XOR2 (N12310, N12309, N7412);
not NOT1 (N12311, N12304);
nor NOR3 (N12312, N12303, N11354, N7669);
xor XOR2 (N12313, N12312, N7424);
buf BUF1 (N12314, N12299);
or OR3 (N12315, N12298, N2603, N10025);
nor NOR4 (N12316, N12311, N8308, N9059, N5070);
nand NAND4 (N12317, N12314, N7399, N7420, N4019);
buf BUF1 (N12318, N12306);
or OR4 (N12319, N12313, N10992, N11509, N11887);
xor XOR2 (N12320, N12318, N10786);
buf BUF1 (N12321, N12317);
buf BUF1 (N12322, N12307);
or OR4 (N12323, N12310, N6320, N12258, N729);
buf BUF1 (N12324, N12308);
xor XOR2 (N12325, N12321, N8498);
and AND3 (N12326, N12319, N7888, N12092);
xor XOR2 (N12327, N12297, N6686);
buf BUF1 (N12328, N12324);
or OR4 (N12329, N12315, N11435, N11516, N3556);
nand NAND3 (N12330, N12325, N4815, N6661);
or OR4 (N12331, N12328, N9512, N3414, N8878);
xor XOR2 (N12332, N12322, N7495);
buf BUF1 (N12333, N12276);
nor NOR4 (N12334, N12331, N5551, N5718, N1755);
and AND4 (N12335, N12329, N2399, N675, N9876);
nand NAND4 (N12336, N12327, N3262, N9064, N5781);
or OR3 (N12337, N12316, N2306, N8551);
or OR2 (N12338, N12323, N1332);
and AND4 (N12339, N12326, N3319, N2917, N3196);
not NOT1 (N12340, N12333);
or OR4 (N12341, N12334, N525, N4260, N7573);
nor NOR2 (N12342, N12332, N7995);
xor XOR2 (N12343, N12340, N9727);
or OR4 (N12344, N12343, N8135, N4497, N8857);
buf BUF1 (N12345, N12337);
nand NAND4 (N12346, N12320, N7400, N10294, N885);
and AND4 (N12347, N12335, N1779, N8153, N8280);
and AND2 (N12348, N12347, N6619);
nor NOR3 (N12349, N12341, N1471, N2585);
xor XOR2 (N12350, N12339, N1494);
nor NOR4 (N12351, N12350, N4578, N2894, N2819);
nand NAND3 (N12352, N12349, N4726, N10808);
xor XOR2 (N12353, N12330, N10690);
or OR2 (N12354, N12351, N6752);
buf BUF1 (N12355, N12345);
xor XOR2 (N12356, N12342, N7684);
buf BUF1 (N12357, N12336);
nor NOR2 (N12358, N12353, N2943);
nor NOR4 (N12359, N12348, N8006, N2472, N11793);
xor XOR2 (N12360, N12346, N6538);
or OR4 (N12361, N12356, N8894, N8888, N7537);
nor NOR2 (N12362, N12338, N2690);
and AND3 (N12363, N12361, N6831, N9967);
not NOT1 (N12364, N12362);
nand NAND2 (N12365, N12357, N10961);
or OR4 (N12366, N12352, N842, N10021, N9753);
nand NAND4 (N12367, N12366, N1063, N3093, N10796);
and AND2 (N12368, N12355, N10361);
not NOT1 (N12369, N12365);
not NOT1 (N12370, N12358);
not NOT1 (N12371, N12344);
xor XOR2 (N12372, N12367, N1213);
or OR3 (N12373, N12372, N7870, N9901);
buf BUF1 (N12374, N12369);
xor XOR2 (N12375, N12373, N572);
xor XOR2 (N12376, N12374, N1539);
or OR3 (N12377, N12364, N7566, N982);
buf BUF1 (N12378, N12376);
xor XOR2 (N12379, N12368, N7313);
and AND3 (N12380, N12371, N12277, N7518);
or OR2 (N12381, N12375, N9767);
buf BUF1 (N12382, N12380);
nor NOR2 (N12383, N12360, N7890);
not NOT1 (N12384, N12370);
not NOT1 (N12385, N12381);
buf BUF1 (N12386, N12354);
and AND2 (N12387, N12377, N1187);
and AND4 (N12388, N12386, N10787, N11583, N9986);
and AND2 (N12389, N12388, N9844);
xor XOR2 (N12390, N12379, N672);
not NOT1 (N12391, N12378);
and AND2 (N12392, N12391, N7617);
nand NAND2 (N12393, N12389, N2559);
and AND4 (N12394, N12390, N7180, N11982, N9370);
nand NAND3 (N12395, N12363, N12166, N10000);
buf BUF1 (N12396, N12395);
not NOT1 (N12397, N12392);
and AND4 (N12398, N12384, N8469, N6662, N1962);
or OR4 (N12399, N12393, N1837, N2817, N1578);
nor NOR4 (N12400, N12383, N2538, N3495, N9844);
xor XOR2 (N12401, N12385, N6786);
or OR3 (N12402, N12401, N6969, N11012);
xor XOR2 (N12403, N12402, N7972);
nand NAND2 (N12404, N12398, N2070);
nor NOR2 (N12405, N12400, N4063);
nand NAND3 (N12406, N12399, N9820, N10145);
buf BUF1 (N12407, N12403);
and AND2 (N12408, N12382, N7013);
or OR3 (N12409, N12407, N1113, N1723);
and AND3 (N12410, N12359, N8254, N9961);
xor XOR2 (N12411, N12397, N4646);
and AND2 (N12412, N12410, N5849);
buf BUF1 (N12413, N12404);
not NOT1 (N12414, N12406);
not NOT1 (N12415, N12411);
and AND4 (N12416, N12415, N10574, N7316, N4541);
nor NOR3 (N12417, N12413, N4512, N4921);
xor XOR2 (N12418, N12396, N3188);
buf BUF1 (N12419, N12409);
xor XOR2 (N12420, N12394, N9651);
or OR4 (N12421, N12416, N11016, N3122, N5665);
nor NOR4 (N12422, N12387, N9341, N975, N3744);
not NOT1 (N12423, N12422);
not NOT1 (N12424, N12423);
or OR4 (N12425, N12421, N11010, N1056, N8446);
or OR4 (N12426, N12424, N5892, N12077, N2660);
nand NAND2 (N12427, N12412, N1466);
and AND2 (N12428, N12419, N9771);
or OR4 (N12429, N12425, N5247, N10497, N9578);
nand NAND3 (N12430, N12405, N2975, N3471);
or OR3 (N12431, N12417, N6763, N11039);
nand NAND2 (N12432, N12420, N4587);
or OR3 (N12433, N12414, N10307, N6295);
or OR3 (N12434, N12432, N8388, N883);
and AND2 (N12435, N12429, N7585);
not NOT1 (N12436, N12433);
xor XOR2 (N12437, N12418, N1082);
not NOT1 (N12438, N12430);
nor NOR2 (N12439, N12436, N4369);
buf BUF1 (N12440, N12437);
nand NAND2 (N12441, N12438, N944);
xor XOR2 (N12442, N12434, N736);
nand NAND2 (N12443, N12426, N10496);
nand NAND4 (N12444, N12441, N1068, N7507, N3997);
nand NAND3 (N12445, N12440, N92, N7151);
not NOT1 (N12446, N12444);
buf BUF1 (N12447, N12427);
nand NAND3 (N12448, N12442, N12422, N7513);
and AND3 (N12449, N12408, N12044, N2758);
nor NOR4 (N12450, N12449, N214, N12278, N5140);
nand NAND2 (N12451, N12448, N11663);
not NOT1 (N12452, N12443);
and AND4 (N12453, N12447, N3712, N9809, N9670);
xor XOR2 (N12454, N12453, N4998);
or OR3 (N12455, N12428, N8782, N11685);
nor NOR4 (N12456, N12452, N5315, N11540, N8083);
buf BUF1 (N12457, N12455);
nor NOR2 (N12458, N12450, N3887);
nand NAND2 (N12459, N12439, N10960);
or OR3 (N12460, N12459, N11072, N11292);
xor XOR2 (N12461, N12431, N5509);
nand NAND2 (N12462, N12456, N836);
and AND4 (N12463, N12458, N6568, N6100, N3156);
nand NAND4 (N12464, N12454, N7973, N5758, N969);
and AND4 (N12465, N12461, N6904, N5778, N6552);
xor XOR2 (N12466, N12460, N8193);
nand NAND2 (N12467, N12463, N7909);
nand NAND2 (N12468, N12467, N7839);
nand NAND2 (N12469, N12465, N4951);
not NOT1 (N12470, N12446);
buf BUF1 (N12471, N12445);
and AND3 (N12472, N12469, N2087, N3497);
and AND2 (N12473, N12468, N11667);
not NOT1 (N12474, N12462);
buf BUF1 (N12475, N12451);
nor NOR4 (N12476, N12466, N271, N2273, N7433);
and AND4 (N12477, N12457, N11334, N11205, N1819);
xor XOR2 (N12478, N12473, N11434);
buf BUF1 (N12479, N12475);
nor NOR4 (N12480, N12435, N5706, N2564, N7798);
buf BUF1 (N12481, N12479);
not NOT1 (N12482, N12472);
not NOT1 (N12483, N12474);
nand NAND3 (N12484, N12482, N9985, N8531);
nor NOR2 (N12485, N12476, N5018);
not NOT1 (N12486, N12484);
nor NOR3 (N12487, N12480, N6911, N4728);
xor XOR2 (N12488, N12481, N9996);
buf BUF1 (N12489, N12485);
or OR2 (N12490, N12486, N313);
and AND4 (N12491, N12490, N11495, N6090, N206);
not NOT1 (N12492, N12489);
or OR2 (N12493, N12492, N7917);
or OR2 (N12494, N12477, N11544);
not NOT1 (N12495, N12488);
and AND4 (N12496, N12487, N8412, N3570, N11557);
nand NAND4 (N12497, N12483, N318, N11709, N4757);
nor NOR4 (N12498, N12493, N3903, N10661, N5680);
or OR3 (N12499, N12495, N2472, N4130);
and AND3 (N12500, N12470, N2682, N4764);
nor NOR3 (N12501, N12471, N1125, N4114);
or OR4 (N12502, N12499, N6935, N10835, N3404);
or OR3 (N12503, N12497, N1352, N9303);
nand NAND3 (N12504, N12491, N10764, N6784);
or OR4 (N12505, N12504, N8871, N4609, N1113);
or OR4 (N12506, N12502, N11860, N3285, N5308);
or OR4 (N12507, N12478, N8311, N3656, N3406);
not NOT1 (N12508, N12464);
or OR2 (N12509, N12503, N4758);
nand NAND4 (N12510, N12507, N8442, N5580, N2706);
nor NOR2 (N12511, N12509, N6444);
and AND3 (N12512, N12510, N8039, N11912);
nor NOR2 (N12513, N12494, N11441);
nand NAND4 (N12514, N12498, N9207, N8558, N8685);
xor XOR2 (N12515, N12514, N6410);
or OR2 (N12516, N12501, N697);
not NOT1 (N12517, N12515);
nor NOR3 (N12518, N12511, N7577, N10856);
buf BUF1 (N12519, N12500);
xor XOR2 (N12520, N12512, N10494);
nand NAND3 (N12521, N12496, N2678, N4015);
and AND2 (N12522, N12506, N7120);
and AND3 (N12523, N12508, N1170, N9336);
or OR3 (N12524, N12505, N6464, N4143);
not NOT1 (N12525, N12523);
or OR2 (N12526, N12520, N5872);
xor XOR2 (N12527, N12518, N7249);
or OR3 (N12528, N12521, N5118, N2446);
and AND2 (N12529, N12522, N5940);
buf BUF1 (N12530, N12517);
or OR3 (N12531, N12525, N640, N143);
nand NAND4 (N12532, N12527, N4257, N10249, N4209);
not NOT1 (N12533, N12519);
nand NAND4 (N12534, N12529, N12458, N1125, N5413);
buf BUF1 (N12535, N12516);
buf BUF1 (N12536, N12524);
or OR2 (N12537, N12532, N8178);
and AND4 (N12538, N12530, N2256, N11304, N7809);
xor XOR2 (N12539, N12528, N3664);
buf BUF1 (N12540, N12539);
not NOT1 (N12541, N12531);
nor NOR4 (N12542, N12537, N7621, N5747, N7696);
buf BUF1 (N12543, N12536);
nand NAND2 (N12544, N12535, N5395);
nor NOR2 (N12545, N12526, N11193);
nor NOR3 (N12546, N12541, N9268, N8866);
or OR4 (N12547, N12540, N3307, N11378, N12088);
xor XOR2 (N12548, N12538, N10909);
buf BUF1 (N12549, N12534);
or OR4 (N12550, N12543, N1903, N4555, N7244);
or OR2 (N12551, N12544, N9461);
or OR4 (N12552, N12548, N6734, N11999, N5300);
or OR2 (N12553, N12513, N1364);
not NOT1 (N12554, N12542);
nor NOR4 (N12555, N12554, N8376, N152, N5916);
buf BUF1 (N12556, N12546);
and AND4 (N12557, N12556, N2135, N412, N5057);
xor XOR2 (N12558, N12555, N3724);
nor NOR3 (N12559, N12552, N10705, N6879);
nand NAND4 (N12560, N12547, N7653, N210, N4777);
nand NAND2 (N12561, N12549, N5127);
and AND4 (N12562, N12550, N8735, N6282, N2975);
nand NAND3 (N12563, N12561, N1501, N12353);
and AND4 (N12564, N12545, N5949, N9889, N5723);
and AND4 (N12565, N12564, N8337, N4366, N2628);
xor XOR2 (N12566, N12557, N9023);
not NOT1 (N12567, N12565);
nor NOR2 (N12568, N12566, N8513);
and AND3 (N12569, N12558, N1466, N185);
not NOT1 (N12570, N12553);
nor NOR2 (N12571, N12533, N7807);
or OR3 (N12572, N12563, N1862, N236);
or OR4 (N12573, N12570, N7400, N6695, N4223);
xor XOR2 (N12574, N12567, N5940);
nand NAND3 (N12575, N12568, N10353, N8327);
or OR2 (N12576, N12574, N1243);
nor NOR2 (N12577, N12559, N2724);
not NOT1 (N12578, N12575);
nor NOR2 (N12579, N12576, N10132);
or OR2 (N12580, N12560, N3624);
or OR2 (N12581, N12562, N3398);
or OR2 (N12582, N12580, N12530);
or OR2 (N12583, N12569, N6463);
and AND4 (N12584, N12573, N598, N7279, N10488);
not NOT1 (N12585, N12582);
xor XOR2 (N12586, N12585, N10058);
and AND3 (N12587, N12579, N1911, N2221);
xor XOR2 (N12588, N12577, N5351);
not NOT1 (N12589, N12578);
xor XOR2 (N12590, N12571, N2157);
nand NAND3 (N12591, N12589, N3978, N7333);
or OR2 (N12592, N12590, N8795);
nand NAND2 (N12593, N12587, N4516);
buf BUF1 (N12594, N12591);
not NOT1 (N12595, N12572);
not NOT1 (N12596, N12595);
buf BUF1 (N12597, N12588);
xor XOR2 (N12598, N12594, N4481);
nor NOR4 (N12599, N12583, N2870, N227, N8899);
not NOT1 (N12600, N12599);
and AND2 (N12601, N12598, N4289);
or OR4 (N12602, N12551, N2864, N11511, N6169);
and AND3 (N12603, N12600, N4540, N832);
and AND4 (N12604, N12603, N4695, N12462, N7238);
nand NAND3 (N12605, N12601, N4063, N626);
xor XOR2 (N12606, N12586, N11582);
buf BUF1 (N12607, N12602);
buf BUF1 (N12608, N12597);
buf BUF1 (N12609, N12581);
nand NAND4 (N12610, N12596, N11200, N6974, N10645);
or OR2 (N12611, N12605, N3367);
buf BUF1 (N12612, N12607);
or OR4 (N12613, N12593, N623, N1294, N5377);
and AND2 (N12614, N12612, N9660);
buf BUF1 (N12615, N12606);
or OR4 (N12616, N12610, N362, N12090, N10029);
and AND2 (N12617, N12604, N910);
and AND3 (N12618, N12608, N11557, N8628);
xor XOR2 (N12619, N12613, N2167);
and AND3 (N12620, N12609, N7326, N9067);
or OR3 (N12621, N12611, N5085, N4606);
buf BUF1 (N12622, N12615);
buf BUF1 (N12623, N12614);
xor XOR2 (N12624, N12618, N5980);
buf BUF1 (N12625, N12624);
nor NOR3 (N12626, N12625, N3839, N11270);
nand NAND3 (N12627, N12592, N11584, N12232);
nand NAND4 (N12628, N12619, N4712, N3824, N5862);
nor NOR2 (N12629, N12616, N9392);
and AND3 (N12630, N12584, N7580, N4569);
nand NAND3 (N12631, N12623, N977, N1595);
or OR2 (N12632, N12626, N4107);
and AND3 (N12633, N12632, N9262, N12622);
nand NAND2 (N12634, N63, N7833);
nand NAND2 (N12635, N12633, N888);
not NOT1 (N12636, N12634);
nor NOR4 (N12637, N12621, N4693, N9710, N5828);
buf BUF1 (N12638, N12629);
nor NOR2 (N12639, N12630, N7064);
and AND3 (N12640, N12637, N6695, N148);
not NOT1 (N12641, N12639);
nand NAND4 (N12642, N12631, N10887, N12214, N5488);
and AND2 (N12643, N12638, N84);
xor XOR2 (N12644, N12617, N7945);
xor XOR2 (N12645, N12627, N724);
and AND2 (N12646, N12645, N2418);
or OR3 (N12647, N12635, N10493, N6753);
buf BUF1 (N12648, N12628);
nor NOR4 (N12649, N12646, N650, N432, N10672);
nor NOR2 (N12650, N12644, N6451);
nor NOR2 (N12651, N12643, N11285);
nand NAND3 (N12652, N12642, N4537, N6590);
nor NOR3 (N12653, N12641, N2734, N6839);
xor XOR2 (N12654, N12650, N7950);
or OR3 (N12655, N12647, N10138, N1446);
xor XOR2 (N12656, N12651, N1211);
and AND2 (N12657, N12648, N1413);
and AND2 (N12658, N12649, N10171);
nand NAND4 (N12659, N12656, N8975, N1307, N10069);
and AND4 (N12660, N12655, N10115, N8286, N5523);
buf BUF1 (N12661, N12636);
xor XOR2 (N12662, N12660, N3476);
or OR4 (N12663, N12652, N8637, N12089, N2124);
not NOT1 (N12664, N12653);
or OR4 (N12665, N12658, N4812, N11800, N7965);
nor NOR3 (N12666, N12620, N2796, N4632);
not NOT1 (N12667, N12665);
and AND3 (N12668, N12661, N270, N3529);
not NOT1 (N12669, N12666);
or OR4 (N12670, N12668, N7890, N2573, N8946);
or OR2 (N12671, N12670, N6127);
or OR3 (N12672, N12662, N10467, N494);
not NOT1 (N12673, N12654);
nand NAND3 (N12674, N12669, N10829, N8725);
and AND2 (N12675, N12671, N2010);
nor NOR2 (N12676, N12664, N4662);
or OR4 (N12677, N12674, N3352, N2994, N676);
nand NAND3 (N12678, N12675, N4241, N3392);
not NOT1 (N12679, N12673);
nand NAND2 (N12680, N12640, N11773);
nor NOR2 (N12681, N12657, N65);
and AND4 (N12682, N12672, N2245, N12463, N7541);
or OR2 (N12683, N12681, N1930);
xor XOR2 (N12684, N12680, N11501);
xor XOR2 (N12685, N12677, N286);
buf BUF1 (N12686, N12663);
and AND2 (N12687, N12667, N10845);
xor XOR2 (N12688, N12687, N5357);
or OR4 (N12689, N12659, N4891, N787, N6739);
nor NOR2 (N12690, N12689, N11795);
xor XOR2 (N12691, N12685, N7298);
nand NAND3 (N12692, N12683, N7561, N6847);
and AND4 (N12693, N12686, N2852, N10697, N10747);
buf BUF1 (N12694, N12679);
nand NAND3 (N12695, N12684, N554, N5390);
buf BUF1 (N12696, N12690);
nand NAND3 (N12697, N12692, N7896, N12176);
and AND3 (N12698, N12693, N4927, N10815);
and AND2 (N12699, N12691, N3670);
buf BUF1 (N12700, N12699);
nand NAND3 (N12701, N12696, N7103, N5439);
buf BUF1 (N12702, N12676);
nand NAND4 (N12703, N12694, N2327, N9431, N2602);
xor XOR2 (N12704, N12695, N7918);
nor NOR2 (N12705, N12704, N2760);
and AND2 (N12706, N12703, N3252);
not NOT1 (N12707, N12678);
nand NAND2 (N12708, N12697, N6217);
not NOT1 (N12709, N12706);
nor NOR3 (N12710, N12700, N10451, N841);
not NOT1 (N12711, N12710);
or OR3 (N12712, N12688, N10895, N10330);
xor XOR2 (N12713, N12682, N8749);
not NOT1 (N12714, N12713);
not NOT1 (N12715, N12708);
not NOT1 (N12716, N12712);
buf BUF1 (N12717, N12705);
or OR3 (N12718, N12711, N2639, N637);
or OR2 (N12719, N12718, N7238);
xor XOR2 (N12720, N12716, N11192);
xor XOR2 (N12721, N12709, N9460);
buf BUF1 (N12722, N12720);
not NOT1 (N12723, N12719);
not NOT1 (N12724, N12717);
nor NOR4 (N12725, N12721, N8054, N8593, N10285);
nand NAND4 (N12726, N12715, N11859, N10893, N7311);
buf BUF1 (N12727, N12722);
or OR4 (N12728, N12726, N1965, N4330, N10989);
nor NOR3 (N12729, N12728, N8248, N6681);
xor XOR2 (N12730, N12724, N7237);
buf BUF1 (N12731, N12701);
xor XOR2 (N12732, N12725, N8203);
not NOT1 (N12733, N12707);
nand NAND2 (N12734, N12698, N5366);
buf BUF1 (N12735, N12702);
or OR3 (N12736, N12723, N279, N10157);
xor XOR2 (N12737, N12714, N11404);
not NOT1 (N12738, N12729);
not NOT1 (N12739, N12727);
nand NAND2 (N12740, N12731, N9535);
and AND4 (N12741, N12732, N8035, N6068, N1228);
buf BUF1 (N12742, N12735);
not NOT1 (N12743, N12733);
nor NOR3 (N12744, N12741, N12588, N5579);
nor NOR4 (N12745, N12743, N5191, N8349, N11413);
nor NOR3 (N12746, N12737, N7093, N4256);
buf BUF1 (N12747, N12742);
and AND2 (N12748, N12736, N9171);
xor XOR2 (N12749, N12734, N8037);
not NOT1 (N12750, N12730);
nor NOR3 (N12751, N12745, N4891, N12611);
not NOT1 (N12752, N12744);
xor XOR2 (N12753, N12751, N11751);
nand NAND3 (N12754, N12750, N3837, N11484);
and AND3 (N12755, N12754, N8622, N10258);
nor NOR3 (N12756, N12753, N3031, N8302);
nor NOR3 (N12757, N12749, N1256, N11948);
nand NAND3 (N12758, N12757, N5021, N8087);
buf BUF1 (N12759, N12738);
buf BUF1 (N12760, N12756);
nor NOR4 (N12761, N12758, N8961, N7926, N4233);
buf BUF1 (N12762, N12740);
nor NOR3 (N12763, N12759, N11013, N689);
or OR2 (N12764, N12747, N4249);
not NOT1 (N12765, N12761);
xor XOR2 (N12766, N12765, N7112);
and AND4 (N12767, N12762, N6145, N1757, N730);
nand NAND4 (N12768, N12748, N12735, N8517, N9898);
buf BUF1 (N12769, N12739);
not NOT1 (N12770, N12746);
nand NAND2 (N12771, N12766, N758);
not NOT1 (N12772, N12767);
nor NOR2 (N12773, N12771, N3617);
and AND4 (N12774, N12764, N9674, N11666, N5840);
not NOT1 (N12775, N12755);
xor XOR2 (N12776, N12769, N8053);
or OR4 (N12777, N12773, N8720, N3693, N4404);
not NOT1 (N12778, N12768);
nand NAND3 (N12779, N12777, N10535, N4466);
not NOT1 (N12780, N12776);
or OR4 (N12781, N12778, N4863, N3828, N9842);
xor XOR2 (N12782, N12752, N9247);
or OR3 (N12783, N12760, N10057, N11695);
xor XOR2 (N12784, N12763, N7581);
xor XOR2 (N12785, N12774, N954);
nor NOR3 (N12786, N12779, N9795, N5876);
and AND4 (N12787, N12775, N12181, N2107, N7287);
or OR4 (N12788, N12783, N473, N7954, N4122);
nand NAND2 (N12789, N12786, N10966);
not NOT1 (N12790, N12780);
or OR4 (N12791, N12790, N12021, N8400, N7700);
not NOT1 (N12792, N12784);
or OR3 (N12793, N12791, N2637, N2221);
nor NOR4 (N12794, N12782, N7512, N5393, N6021);
not NOT1 (N12795, N12785);
xor XOR2 (N12796, N12781, N12784);
or OR4 (N12797, N12772, N8124, N6561, N4619);
not NOT1 (N12798, N12793);
nand NAND4 (N12799, N12788, N2094, N1249, N1961);
buf BUF1 (N12800, N12787);
xor XOR2 (N12801, N12797, N3792);
or OR4 (N12802, N12795, N11282, N3091, N5537);
not NOT1 (N12803, N12789);
not NOT1 (N12804, N12802);
nand NAND3 (N12805, N12799, N8487, N9562);
not NOT1 (N12806, N12804);
xor XOR2 (N12807, N12770, N11806);
buf BUF1 (N12808, N12794);
nor NOR2 (N12809, N12801, N9575);
xor XOR2 (N12810, N12796, N9348);
nor NOR4 (N12811, N12803, N10197, N8817, N12429);
xor XOR2 (N12812, N12806, N1894);
buf BUF1 (N12813, N12807);
not NOT1 (N12814, N12812);
xor XOR2 (N12815, N12792, N544);
not NOT1 (N12816, N12800);
not NOT1 (N12817, N12798);
nor NOR2 (N12818, N12817, N7116);
nand NAND4 (N12819, N12808, N9863, N4840, N977);
and AND4 (N12820, N12813, N589, N3439, N1239);
and AND3 (N12821, N12818, N9333, N5274);
endmodule