// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13;

output N8011,N7997,N8003,N7968,N8008,N8000,N7996,N8007,N8006,N8013;

not NOT1 (N14, N2);
xor XOR2 (N15, N2, N2);
and AND4 (N16, N7, N6, N15, N5);
nand NAND4 (N17, N2, N14, N6, N5);
nor NOR4 (N18, N7, N6, N15, N1);
nor NOR4 (N19, N6, N17, N5, N12);
and AND3 (N20, N2, N19, N2);
or OR3 (N21, N13, N5, N20);
and AND4 (N22, N4, N5, N14, N18);
nor NOR2 (N23, N1, N3);
and AND3 (N24, N17, N4, N15);
buf BUF1 (N25, N3);
and AND3 (N26, N13, N24, N10);
or OR2 (N27, N6, N12);
nor NOR4 (N28, N9, N15, N18, N3);
not NOT1 (N29, N23);
or OR2 (N30, N7, N20);
and AND4 (N31, N5, N5, N15, N3);
buf BUF1 (N32, N28);
or OR2 (N33, N25, N32);
nand NAND2 (N34, N32, N1);
xor XOR2 (N35, N34, N29);
and AND2 (N36, N6, N35);
not NOT1 (N37, N19);
not NOT1 (N38, N26);
nor NOR3 (N39, N37, N32, N34);
xor XOR2 (N40, N36, N8);
xor XOR2 (N41, N22, N34);
or OR3 (N42, N16, N35, N38);
not NOT1 (N43, N38);
buf BUF1 (N44, N30);
and AND3 (N45, N27, N16, N23);
nor NOR4 (N46, N44, N23, N24, N42);
nand NAND4 (N47, N10, N43, N19, N45);
not NOT1 (N48, N36);
not NOT1 (N49, N46);
or OR4 (N50, N24, N1, N34, N15);
and AND2 (N51, N31, N1);
xor XOR2 (N52, N50, N23);
nand NAND3 (N53, N39, N29, N14);
nand NAND4 (N54, N47, N38, N25, N16);
buf BUF1 (N55, N40);
not NOT1 (N56, N49);
and AND2 (N57, N51, N47);
xor XOR2 (N58, N56, N13);
nand NAND4 (N59, N57, N13, N21, N48);
nor NOR3 (N60, N9, N9, N40);
or OR2 (N61, N48, N56);
nor NOR2 (N62, N53, N13);
nor NOR2 (N63, N59, N62);
nor NOR2 (N64, N6, N20);
nor NOR4 (N65, N58, N34, N62, N30);
or OR2 (N66, N55, N39);
xor XOR2 (N67, N41, N58);
xor XOR2 (N68, N33, N13);
or OR3 (N69, N67, N15, N67);
buf BUF1 (N70, N65);
nor NOR4 (N71, N52, N40, N24, N33);
nand NAND3 (N72, N64, N57, N49);
and AND4 (N73, N71, N18, N11, N44);
and AND2 (N74, N66, N29);
not NOT1 (N75, N74);
nor NOR4 (N76, N73, N21, N51, N30);
buf BUF1 (N77, N75);
or OR2 (N78, N76, N1);
nor NOR4 (N79, N63, N50, N77, N25);
nor NOR4 (N80, N39, N38, N69, N37);
and AND4 (N81, N26, N68, N44, N6);
not NOT1 (N82, N68);
or OR2 (N83, N81, N18);
buf BUF1 (N84, N54);
nor NOR4 (N85, N70, N53, N57, N40);
buf BUF1 (N86, N83);
or OR2 (N87, N84, N59);
and AND2 (N88, N87, N47);
or OR2 (N89, N61, N51);
and AND4 (N90, N60, N6, N71, N78);
or OR4 (N91, N33, N36, N60, N37);
not NOT1 (N92, N72);
nor NOR3 (N93, N86, N21, N63);
xor XOR2 (N94, N92, N11);
buf BUF1 (N95, N82);
xor XOR2 (N96, N94, N22);
and AND2 (N97, N85, N25);
buf BUF1 (N98, N79);
or OR3 (N99, N88, N54, N60);
xor XOR2 (N100, N96, N75);
xor XOR2 (N101, N93, N11);
xor XOR2 (N102, N90, N49);
and AND2 (N103, N89, N10);
xor XOR2 (N104, N101, N36);
and AND4 (N105, N80, N2, N88, N50);
xor XOR2 (N106, N100, N20);
xor XOR2 (N107, N97, N85);
not NOT1 (N108, N98);
and AND3 (N109, N108, N18, N58);
buf BUF1 (N110, N104);
and AND4 (N111, N107, N91, N15, N48);
nand NAND3 (N112, N26, N70, N106);
and AND3 (N113, N33, N46, N35);
not NOT1 (N114, N113);
xor XOR2 (N115, N112, N79);
buf BUF1 (N116, N105);
xor XOR2 (N117, N109, N45);
xor XOR2 (N118, N116, N75);
and AND2 (N119, N103, N35);
not NOT1 (N120, N95);
and AND2 (N121, N110, N53);
or OR2 (N122, N115, N83);
and AND2 (N123, N114, N53);
and AND2 (N124, N111, N43);
not NOT1 (N125, N124);
not NOT1 (N126, N125);
nand NAND4 (N127, N118, N70, N98, N84);
and AND4 (N128, N119, N75, N69, N107);
xor XOR2 (N129, N102, N77);
nand NAND3 (N130, N129, N57, N21);
nand NAND3 (N131, N127, N47, N108);
or OR4 (N132, N126, N2, N97, N118);
buf BUF1 (N133, N123);
nand NAND4 (N134, N120, N116, N37, N84);
or OR4 (N135, N128, N56, N86, N95);
xor XOR2 (N136, N122, N60);
nand NAND3 (N137, N135, N107, N76);
nand NAND3 (N138, N130, N77, N62);
buf BUF1 (N139, N121);
or OR4 (N140, N132, N32, N137, N9);
not NOT1 (N141, N108);
or OR3 (N142, N134, N141, N67);
nand NAND4 (N143, N6, N22, N102, N112);
xor XOR2 (N144, N143, N81);
nor NOR3 (N145, N131, N36, N59);
nor NOR2 (N146, N145, N72);
and AND2 (N147, N146, N64);
xor XOR2 (N148, N139, N11);
not NOT1 (N149, N140);
not NOT1 (N150, N138);
nor NOR4 (N151, N150, N14, N77, N25);
nor NOR3 (N152, N148, N125, N51);
nand NAND3 (N153, N99, N12, N125);
not NOT1 (N154, N147);
nand NAND2 (N155, N117, N21);
xor XOR2 (N156, N133, N23);
or OR4 (N157, N156, N103, N26, N44);
buf BUF1 (N158, N155);
not NOT1 (N159, N158);
nand NAND2 (N160, N144, N16);
and AND3 (N161, N154, N80, N69);
nand NAND2 (N162, N151, N27);
buf BUF1 (N163, N136);
nor NOR2 (N164, N149, N28);
and AND3 (N165, N142, N118, N145);
nor NOR4 (N166, N163, N25, N141, N20);
not NOT1 (N167, N161);
buf BUF1 (N168, N157);
xor XOR2 (N169, N159, N92);
or OR3 (N170, N160, N94, N143);
nand NAND4 (N171, N165, N141, N77, N152);
or OR2 (N172, N170, N124);
not NOT1 (N173, N20);
not NOT1 (N174, N153);
not NOT1 (N175, N169);
not NOT1 (N176, N174);
xor XOR2 (N177, N172, N171);
xor XOR2 (N178, N106, N12);
and AND2 (N179, N177, N31);
and AND3 (N180, N178, N49, N6);
or OR2 (N181, N167, N80);
or OR2 (N182, N179, N114);
xor XOR2 (N183, N164, N72);
or OR4 (N184, N183, N80, N171, N50);
buf BUF1 (N185, N180);
nor NOR2 (N186, N185, N34);
not NOT1 (N187, N173);
buf BUF1 (N188, N168);
not NOT1 (N189, N176);
or OR4 (N190, N181, N2, N105, N163);
buf BUF1 (N191, N190);
buf BUF1 (N192, N162);
and AND3 (N193, N166, N67, N103);
nand NAND3 (N194, N191, N81, N24);
nand NAND3 (N195, N192, N95, N52);
not NOT1 (N196, N175);
nor NOR3 (N197, N194, N60, N21);
and AND3 (N198, N186, N155, N181);
buf BUF1 (N199, N184);
and AND3 (N200, N197, N157, N81);
or OR3 (N201, N198, N53, N55);
buf BUF1 (N202, N193);
nand NAND2 (N203, N201, N123);
not NOT1 (N204, N188);
not NOT1 (N205, N200);
or OR4 (N206, N187, N55, N94, N204);
and AND2 (N207, N178, N62);
or OR4 (N208, N203, N1, N168, N199);
and AND2 (N209, N191, N67);
nor NOR2 (N210, N195, N117);
xor XOR2 (N211, N205, N91);
buf BUF1 (N212, N206);
nor NOR3 (N213, N182, N205, N178);
xor XOR2 (N214, N196, N94);
buf BUF1 (N215, N202);
nand NAND4 (N216, N207, N149, N126, N36);
nand NAND4 (N217, N215, N87, N90, N51);
nor NOR4 (N218, N214, N80, N5, N75);
and AND4 (N219, N189, N33, N156, N211);
nand NAND3 (N220, N121, N133, N2);
nor NOR4 (N221, N220, N45, N10, N200);
buf BUF1 (N222, N219);
not NOT1 (N223, N210);
nor NOR2 (N224, N212, N64);
nand NAND2 (N225, N208, N89);
buf BUF1 (N226, N213);
buf BUF1 (N227, N226);
xor XOR2 (N228, N227, N192);
nor NOR2 (N229, N217, N226);
and AND4 (N230, N225, N5, N24, N134);
nand NAND4 (N231, N221, N121, N118, N51);
buf BUF1 (N232, N229);
nor NOR2 (N233, N224, N102);
nor NOR3 (N234, N216, N5, N117);
nor NOR2 (N235, N233, N178);
not NOT1 (N236, N218);
nor NOR3 (N237, N230, N138, N188);
xor XOR2 (N238, N228, N217);
or OR3 (N239, N237, N155, N152);
nor NOR4 (N240, N222, N122, N199, N89);
nor NOR2 (N241, N240, N73);
not NOT1 (N242, N223);
buf BUF1 (N243, N231);
and AND4 (N244, N238, N149, N97, N6);
xor XOR2 (N245, N232, N178);
nand NAND3 (N246, N234, N19, N48);
and AND3 (N247, N242, N198, N31);
nor NOR4 (N248, N245, N107, N124, N236);
nor NOR2 (N249, N22, N243);
buf BUF1 (N250, N48);
nor NOR3 (N251, N235, N54, N42);
nor NOR2 (N252, N247, N249);
or OR3 (N253, N80, N98, N32);
buf BUF1 (N254, N252);
nor NOR3 (N255, N248, N46, N22);
not NOT1 (N256, N253);
nand NAND2 (N257, N239, N226);
and AND3 (N258, N241, N74, N130);
buf BUF1 (N259, N254);
and AND3 (N260, N259, N174, N86);
buf BUF1 (N261, N256);
or OR2 (N262, N209, N177);
buf BUF1 (N263, N260);
and AND3 (N264, N258, N198, N155);
buf BUF1 (N265, N262);
and AND3 (N266, N257, N134, N204);
nand NAND2 (N267, N251, N193);
or OR4 (N268, N265, N153, N152, N246);
or OR4 (N269, N154, N211, N130, N12);
not NOT1 (N270, N266);
nor NOR3 (N271, N250, N43, N57);
nand NAND4 (N272, N244, N83, N17, N83);
nor NOR4 (N273, N271, N147, N155, N83);
not NOT1 (N274, N272);
not NOT1 (N275, N268);
or OR3 (N276, N273, N114, N209);
buf BUF1 (N277, N276);
not NOT1 (N278, N263);
buf BUF1 (N279, N275);
and AND2 (N280, N267, N27);
buf BUF1 (N281, N255);
not NOT1 (N282, N280);
nor NOR3 (N283, N279, N71, N170);
or OR4 (N284, N282, N53, N271, N89);
and AND2 (N285, N274, N268);
xor XOR2 (N286, N261, N55);
nand NAND2 (N287, N283, N18);
or OR2 (N288, N284, N137);
buf BUF1 (N289, N278);
not NOT1 (N290, N287);
nand NAND4 (N291, N290, N75, N204, N65);
or OR4 (N292, N277, N157, N203, N142);
not NOT1 (N293, N286);
nor NOR2 (N294, N264, N236);
nand NAND3 (N295, N293, N150, N255);
xor XOR2 (N296, N295, N63);
or OR4 (N297, N270, N259, N232, N117);
not NOT1 (N298, N296);
and AND3 (N299, N298, N231, N253);
buf BUF1 (N300, N285);
not NOT1 (N301, N291);
nor NOR4 (N302, N269, N186, N180, N265);
xor XOR2 (N303, N292, N42);
nand NAND2 (N304, N289, N51);
xor XOR2 (N305, N304, N44);
xor XOR2 (N306, N302, N204);
xor XOR2 (N307, N303, N2);
xor XOR2 (N308, N288, N199);
and AND2 (N309, N308, N234);
not NOT1 (N310, N281);
xor XOR2 (N311, N301, N220);
nand NAND2 (N312, N305, N123);
nor NOR4 (N313, N297, N209, N287, N83);
buf BUF1 (N314, N312);
or OR2 (N315, N307, N207);
xor XOR2 (N316, N299, N121);
and AND4 (N317, N306, N132, N200, N8);
and AND2 (N318, N313, N31);
buf BUF1 (N319, N294);
buf BUF1 (N320, N300);
nor NOR3 (N321, N317, N270, N291);
and AND4 (N322, N310, N198, N103, N172);
nand NAND2 (N323, N319, N63);
buf BUF1 (N324, N316);
nor NOR2 (N325, N324, N303);
xor XOR2 (N326, N323, N199);
buf BUF1 (N327, N320);
or OR2 (N328, N309, N95);
xor XOR2 (N329, N311, N327);
nand NAND2 (N330, N90, N259);
buf BUF1 (N331, N329);
buf BUF1 (N332, N321);
xor XOR2 (N333, N318, N63);
not NOT1 (N334, N314);
nand NAND2 (N335, N334, N329);
or OR3 (N336, N333, N96, N105);
xor XOR2 (N337, N315, N269);
not NOT1 (N338, N332);
and AND3 (N339, N338, N222, N16);
buf BUF1 (N340, N336);
or OR3 (N341, N331, N94, N168);
nor NOR2 (N342, N339, N69);
or OR4 (N343, N322, N230, N23, N290);
nor NOR2 (N344, N340, N119);
xor XOR2 (N345, N330, N96);
nor NOR4 (N346, N342, N280, N220, N155);
nand NAND3 (N347, N335, N199, N31);
nor NOR2 (N348, N346, N307);
not NOT1 (N349, N341);
buf BUF1 (N350, N344);
nor NOR3 (N351, N328, N56, N138);
nor NOR2 (N352, N348, N326);
or OR3 (N353, N340, N234, N135);
and AND3 (N354, N351, N108, N134);
nor NOR2 (N355, N325, N177);
nor NOR3 (N356, N352, N163, N42);
xor XOR2 (N357, N355, N330);
nor NOR3 (N358, N349, N111, N173);
and AND4 (N359, N343, N81, N215, N98);
or OR2 (N360, N347, N24);
and AND4 (N361, N358, N5, N179, N279);
and AND3 (N362, N337, N213, N268);
and AND2 (N363, N357, N234);
or OR4 (N364, N360, N358, N121, N269);
and AND3 (N365, N354, N57, N232);
xor XOR2 (N366, N359, N362);
buf BUF1 (N367, N46);
xor XOR2 (N368, N363, N56);
and AND3 (N369, N345, N223, N35);
nor NOR3 (N370, N367, N351, N59);
or OR3 (N371, N350, N366, N276);
nor NOR4 (N372, N324, N107, N323, N196);
buf BUF1 (N373, N369);
or OR2 (N374, N353, N252);
buf BUF1 (N375, N371);
or OR4 (N376, N361, N272, N139, N272);
or OR2 (N377, N368, N131);
not NOT1 (N378, N373);
and AND3 (N379, N376, N154, N261);
buf BUF1 (N380, N372);
nand NAND3 (N381, N374, N17, N81);
or OR4 (N382, N378, N88, N2, N75);
and AND3 (N383, N379, N295, N323);
and AND4 (N384, N365, N174, N288, N87);
buf BUF1 (N385, N381);
xor XOR2 (N386, N382, N209);
or OR3 (N387, N383, N154, N369);
and AND2 (N388, N370, N117);
xor XOR2 (N389, N364, N241);
xor XOR2 (N390, N380, N315);
or OR2 (N391, N390, N220);
nor NOR4 (N392, N356, N30, N8, N92);
buf BUF1 (N393, N391);
nand NAND4 (N394, N384, N19, N204, N241);
or OR3 (N395, N387, N137, N189);
nand NAND4 (N396, N377, N121, N137, N268);
buf BUF1 (N397, N388);
and AND2 (N398, N389, N377);
nor NOR3 (N399, N395, N232, N265);
xor XOR2 (N400, N386, N55);
nor NOR2 (N401, N396, N15);
xor XOR2 (N402, N393, N333);
buf BUF1 (N403, N375);
buf BUF1 (N404, N398);
xor XOR2 (N405, N399, N400);
buf BUF1 (N406, N177);
or OR3 (N407, N403, N42, N75);
not NOT1 (N408, N405);
buf BUF1 (N409, N401);
nand NAND2 (N410, N409, N55);
nand NAND2 (N411, N402, N400);
buf BUF1 (N412, N394);
nand NAND2 (N413, N410, N146);
and AND4 (N414, N397, N197, N241, N103);
xor XOR2 (N415, N407, N17);
not NOT1 (N416, N411);
buf BUF1 (N417, N415);
or OR2 (N418, N392, N17);
buf BUF1 (N419, N416);
buf BUF1 (N420, N419);
or OR4 (N421, N406, N186, N211, N266);
and AND3 (N422, N418, N323, N397);
xor XOR2 (N423, N420, N419);
buf BUF1 (N424, N412);
nor NOR4 (N425, N417, N410, N342, N238);
xor XOR2 (N426, N404, N351);
or OR4 (N427, N408, N204, N116, N186);
buf BUF1 (N428, N427);
buf BUF1 (N429, N423);
or OR3 (N430, N414, N6, N318);
nor NOR2 (N431, N428, N310);
nor NOR3 (N432, N430, N45, N422);
or OR3 (N433, N310, N322, N416);
xor XOR2 (N434, N385, N366);
not NOT1 (N435, N429);
buf BUF1 (N436, N424);
and AND3 (N437, N421, N146, N329);
xor XOR2 (N438, N425, N97);
nand NAND4 (N439, N431, N385, N106, N340);
and AND2 (N440, N433, N123);
xor XOR2 (N441, N426, N144);
xor XOR2 (N442, N438, N385);
not NOT1 (N443, N440);
xor XOR2 (N444, N442, N387);
not NOT1 (N445, N439);
or OR4 (N446, N413, N357, N256, N55);
xor XOR2 (N447, N441, N407);
xor XOR2 (N448, N437, N8);
nand NAND3 (N449, N447, N193, N80);
xor XOR2 (N450, N446, N447);
and AND4 (N451, N434, N412, N188, N292);
and AND4 (N452, N445, N75, N97, N444);
xor XOR2 (N453, N357, N98);
and AND3 (N454, N453, N387, N186);
not NOT1 (N455, N432);
xor XOR2 (N456, N435, N204);
xor XOR2 (N457, N456, N188);
nand NAND2 (N458, N451, N43);
not NOT1 (N459, N454);
and AND3 (N460, N459, N92, N113);
nand NAND2 (N461, N448, N59);
or OR4 (N462, N436, N385, N345, N263);
nand NAND4 (N463, N461, N40, N1, N241);
buf BUF1 (N464, N452);
nor NOR3 (N465, N462, N161, N5);
buf BUF1 (N466, N463);
nor NOR3 (N467, N460, N216, N145);
nand NAND4 (N468, N467, N381, N1, N213);
xor XOR2 (N469, N449, N163);
xor XOR2 (N470, N469, N242);
not NOT1 (N471, N450);
xor XOR2 (N472, N464, N117);
buf BUF1 (N473, N457);
xor XOR2 (N474, N458, N198);
or OR4 (N475, N473, N292, N251, N465);
or OR2 (N476, N357, N174);
and AND2 (N477, N474, N133);
and AND2 (N478, N471, N453);
and AND4 (N479, N472, N163, N373, N384);
nor NOR2 (N480, N475, N255);
not NOT1 (N481, N479);
nor NOR3 (N482, N480, N257, N326);
and AND4 (N483, N478, N223, N472, N418);
nand NAND4 (N484, N476, N102, N259, N114);
nor NOR4 (N485, N484, N255, N77, N294);
or OR2 (N486, N482, N196);
and AND4 (N487, N486, N272, N89, N409);
and AND4 (N488, N477, N193, N185, N24);
and AND4 (N489, N487, N146, N344, N156);
and AND2 (N490, N488, N328);
nor NOR3 (N491, N483, N329, N92);
not NOT1 (N492, N443);
buf BUF1 (N493, N489);
and AND2 (N494, N492, N248);
buf BUF1 (N495, N466);
nand NAND2 (N496, N468, N410);
not NOT1 (N497, N470);
nand NAND3 (N498, N493, N468, N404);
not NOT1 (N499, N485);
nand NAND4 (N500, N499, N413, N274, N311);
nor NOR3 (N501, N455, N5, N41);
nor NOR2 (N502, N497, N203);
buf BUF1 (N503, N502);
nor NOR2 (N504, N503, N412);
nor NOR2 (N505, N504, N386);
buf BUF1 (N506, N498);
or OR2 (N507, N496, N460);
not NOT1 (N508, N491);
nor NOR3 (N509, N490, N67, N121);
nand NAND2 (N510, N495, N459);
not NOT1 (N511, N500);
not NOT1 (N512, N481);
and AND3 (N513, N511, N168, N134);
not NOT1 (N514, N506);
nand NAND2 (N515, N505, N484);
nand NAND4 (N516, N513, N416, N11, N333);
not NOT1 (N517, N512);
and AND3 (N518, N501, N439, N311);
and AND3 (N519, N515, N95, N412);
buf BUF1 (N520, N509);
buf BUF1 (N521, N519);
nor NOR2 (N522, N516, N191);
nand NAND3 (N523, N510, N337, N506);
nor NOR2 (N524, N522, N128);
nand NAND4 (N525, N494, N253, N105, N102);
and AND2 (N526, N524, N402);
xor XOR2 (N527, N514, N320);
not NOT1 (N528, N508);
or OR3 (N529, N518, N335, N447);
nand NAND4 (N530, N527, N18, N491, N242);
nand NAND3 (N531, N529, N45, N370);
nand NAND4 (N532, N507, N441, N344, N450);
or OR2 (N533, N531, N462);
xor XOR2 (N534, N517, N415);
and AND4 (N535, N520, N519, N51, N331);
and AND3 (N536, N525, N450, N469);
xor XOR2 (N537, N534, N450);
nand NAND4 (N538, N536, N46, N122, N107);
or OR3 (N539, N521, N395, N189);
nor NOR3 (N540, N532, N2, N208);
nor NOR3 (N541, N526, N130, N102);
or OR3 (N542, N539, N283, N37);
nor NOR3 (N543, N535, N166, N266);
and AND4 (N544, N543, N112, N313, N310);
nand NAND2 (N545, N528, N134);
not NOT1 (N546, N542);
and AND4 (N547, N545, N77, N92, N243);
buf BUF1 (N548, N533);
nand NAND2 (N549, N544, N294);
nor NOR3 (N550, N546, N67, N359);
xor XOR2 (N551, N547, N524);
nand NAND4 (N552, N537, N358, N487, N386);
xor XOR2 (N553, N551, N98);
not NOT1 (N554, N549);
nor NOR2 (N555, N548, N348);
nand NAND3 (N556, N555, N247, N386);
nand NAND3 (N557, N552, N211, N362);
xor XOR2 (N558, N530, N402);
buf BUF1 (N559, N540);
xor XOR2 (N560, N538, N291);
xor XOR2 (N561, N554, N496);
nand NAND4 (N562, N561, N95, N361, N372);
not NOT1 (N563, N558);
nand NAND2 (N564, N563, N25);
nand NAND3 (N565, N557, N155, N529);
or OR4 (N566, N550, N318, N282, N300);
and AND2 (N567, N553, N468);
buf BUF1 (N568, N559);
or OR3 (N569, N564, N533, N361);
and AND3 (N570, N560, N198, N368);
or OR3 (N571, N541, N141, N176);
nand NAND4 (N572, N562, N379, N198, N362);
nand NAND2 (N573, N566, N92);
and AND2 (N574, N565, N65);
nand NAND3 (N575, N573, N225, N45);
not NOT1 (N576, N571);
and AND3 (N577, N572, N186, N244);
nor NOR4 (N578, N567, N377, N362, N426);
nor NOR4 (N579, N556, N449, N273, N271);
xor XOR2 (N580, N574, N203);
or OR3 (N581, N569, N230, N501);
xor XOR2 (N582, N523, N554);
xor XOR2 (N583, N578, N218);
not NOT1 (N584, N577);
nand NAND3 (N585, N576, N565, N391);
and AND2 (N586, N583, N370);
or OR4 (N587, N585, N38, N530, N73);
buf BUF1 (N588, N587);
and AND3 (N589, N586, N353, N226);
and AND3 (N590, N568, N247, N578);
or OR3 (N591, N590, N564, N7);
buf BUF1 (N592, N588);
nand NAND3 (N593, N581, N177, N578);
nor NOR2 (N594, N591, N37);
xor XOR2 (N595, N594, N354);
not NOT1 (N596, N579);
nand NAND4 (N597, N575, N148, N529, N198);
and AND4 (N598, N589, N175, N72, N90);
or OR4 (N599, N570, N332, N498, N562);
or OR4 (N600, N596, N374, N519, N189);
not NOT1 (N601, N597);
buf BUF1 (N602, N592);
and AND2 (N603, N602, N47);
nor NOR3 (N604, N601, N168, N536);
not NOT1 (N605, N604);
and AND4 (N606, N593, N372, N187, N426);
not NOT1 (N607, N603);
xor XOR2 (N608, N605, N7);
and AND3 (N609, N584, N46, N330);
or OR2 (N610, N580, N388);
and AND4 (N611, N607, N167, N474, N328);
buf BUF1 (N612, N598);
nor NOR4 (N613, N612, N419, N390, N170);
and AND3 (N614, N606, N123, N517);
and AND4 (N615, N610, N488, N452, N232);
nor NOR3 (N616, N614, N283, N587);
xor XOR2 (N617, N600, N86);
nor NOR2 (N618, N595, N570);
or OR4 (N619, N617, N570, N341, N185);
nor NOR3 (N620, N616, N178, N65);
and AND4 (N621, N620, N334, N277, N410);
not NOT1 (N622, N608);
or OR4 (N623, N615, N495, N605, N523);
and AND2 (N624, N622, N183);
not NOT1 (N625, N599);
and AND3 (N626, N619, N320, N209);
not NOT1 (N627, N611);
or OR3 (N628, N582, N66, N507);
xor XOR2 (N629, N625, N579);
nand NAND3 (N630, N623, N108, N469);
and AND3 (N631, N609, N154, N586);
nor NOR2 (N632, N628, N444);
or OR2 (N633, N626, N172);
and AND2 (N634, N627, N237);
xor XOR2 (N635, N632, N47);
or OR2 (N636, N618, N275);
xor XOR2 (N637, N633, N127);
xor XOR2 (N638, N635, N193);
and AND2 (N639, N637, N501);
or OR4 (N640, N613, N561, N546, N364);
buf BUF1 (N641, N630);
xor XOR2 (N642, N621, N120);
buf BUF1 (N643, N638);
and AND4 (N644, N642, N2, N471, N289);
or OR4 (N645, N641, N304, N252, N206);
buf BUF1 (N646, N643);
buf BUF1 (N647, N645);
or OR2 (N648, N631, N27);
not NOT1 (N649, N636);
nor NOR2 (N650, N639, N630);
nor NOR4 (N651, N624, N217, N70, N381);
not NOT1 (N652, N650);
buf BUF1 (N653, N629);
nor NOR2 (N654, N649, N382);
not NOT1 (N655, N640);
buf BUF1 (N656, N648);
nor NOR4 (N657, N654, N96, N594, N116);
xor XOR2 (N658, N656, N207);
not NOT1 (N659, N647);
buf BUF1 (N660, N644);
and AND3 (N661, N652, N130, N171);
nor NOR3 (N662, N651, N227, N123);
or OR3 (N663, N661, N188, N194);
and AND2 (N664, N658, N397);
buf BUF1 (N665, N664);
and AND4 (N666, N665, N208, N631, N622);
and AND3 (N667, N655, N453, N190);
or OR2 (N668, N660, N229);
nand NAND2 (N669, N657, N418);
xor XOR2 (N670, N634, N508);
nand NAND4 (N671, N670, N497, N182, N654);
nor NOR2 (N672, N666, N563);
not NOT1 (N673, N663);
or OR3 (N674, N667, N113, N251);
xor XOR2 (N675, N671, N521);
not NOT1 (N676, N674);
or OR4 (N677, N676, N158, N532, N160);
and AND3 (N678, N672, N444, N121);
and AND2 (N679, N668, N406);
and AND2 (N680, N673, N382);
nor NOR4 (N681, N662, N601, N413, N656);
buf BUF1 (N682, N677);
xor XOR2 (N683, N675, N127);
xor XOR2 (N684, N678, N371);
xor XOR2 (N685, N683, N677);
not NOT1 (N686, N681);
nor NOR2 (N687, N680, N165);
nand NAND3 (N688, N686, N254, N482);
nor NOR4 (N689, N688, N543, N78, N261);
buf BUF1 (N690, N653);
and AND4 (N691, N690, N379, N601, N421);
nor NOR4 (N692, N687, N645, N665, N615);
nor NOR3 (N693, N679, N630, N307);
and AND4 (N694, N692, N355, N644, N383);
and AND4 (N695, N669, N626, N596, N110);
nor NOR3 (N696, N646, N486, N277);
and AND3 (N697, N695, N688, N366);
buf BUF1 (N698, N684);
or OR4 (N699, N696, N476, N645, N604);
or OR4 (N700, N682, N14, N175, N167);
buf BUF1 (N701, N685);
xor XOR2 (N702, N691, N383);
not NOT1 (N703, N701);
or OR3 (N704, N694, N59, N512);
xor XOR2 (N705, N689, N511);
nor NOR3 (N706, N697, N540, N480);
xor XOR2 (N707, N698, N364);
and AND3 (N708, N705, N612, N228);
nor NOR2 (N709, N703, N304);
xor XOR2 (N710, N709, N288);
not NOT1 (N711, N710);
or OR3 (N712, N693, N230, N516);
or OR3 (N713, N708, N558, N108);
buf BUF1 (N714, N700);
buf BUF1 (N715, N713);
buf BUF1 (N716, N707);
and AND2 (N717, N714, N463);
or OR3 (N718, N715, N371, N237);
xor XOR2 (N719, N699, N558);
or OR4 (N720, N704, N638, N433, N4);
xor XOR2 (N721, N711, N528);
xor XOR2 (N722, N706, N190);
or OR4 (N723, N721, N241, N420, N649);
or OR3 (N724, N719, N347, N708);
buf BUF1 (N725, N722);
buf BUF1 (N726, N718);
and AND4 (N727, N659, N277, N337, N449);
and AND3 (N728, N725, N375, N270);
nand NAND4 (N729, N726, N659, N605, N48);
and AND3 (N730, N720, N12, N161);
buf BUF1 (N731, N728);
nand NAND4 (N732, N716, N224, N166, N421);
nor NOR2 (N733, N717, N706);
not NOT1 (N734, N733);
nor NOR3 (N735, N730, N228, N131);
buf BUF1 (N736, N712);
not NOT1 (N737, N724);
and AND2 (N738, N723, N476);
not NOT1 (N739, N734);
buf BUF1 (N740, N731);
xor XOR2 (N741, N736, N258);
nand NAND4 (N742, N741, N629, N518, N356);
or OR2 (N743, N739, N306);
not NOT1 (N744, N735);
nand NAND4 (N745, N737, N257, N65, N304);
not NOT1 (N746, N732);
or OR3 (N747, N727, N676, N14);
or OR4 (N748, N729, N106, N215, N127);
nand NAND3 (N749, N738, N586, N652);
buf BUF1 (N750, N743);
or OR2 (N751, N742, N521);
and AND4 (N752, N750, N382, N456, N214);
nand NAND2 (N753, N744, N660);
not NOT1 (N754, N753);
or OR3 (N755, N751, N328, N482);
not NOT1 (N756, N702);
not NOT1 (N757, N746);
or OR4 (N758, N740, N552, N221, N618);
nand NAND3 (N759, N749, N296, N717);
and AND2 (N760, N752, N419);
nand NAND3 (N761, N747, N279, N625);
nor NOR2 (N762, N748, N395);
nor NOR4 (N763, N762, N538, N474, N111);
and AND4 (N764, N745, N419, N203, N500);
or OR2 (N765, N756, N218);
nor NOR3 (N766, N765, N460, N602);
nand NAND2 (N767, N754, N552);
nand NAND4 (N768, N763, N275, N626, N13);
buf BUF1 (N769, N757);
and AND2 (N770, N767, N746);
or OR3 (N771, N761, N109, N631);
buf BUF1 (N772, N764);
xor XOR2 (N773, N759, N545);
or OR2 (N774, N771, N160);
or OR2 (N775, N766, N718);
nor NOR2 (N776, N768, N638);
nand NAND2 (N777, N774, N372);
nand NAND4 (N778, N770, N332, N341, N507);
not NOT1 (N779, N758);
and AND2 (N780, N755, N711);
xor XOR2 (N781, N779, N79);
nand NAND4 (N782, N776, N169, N550, N99);
or OR3 (N783, N782, N310, N48);
not NOT1 (N784, N780);
or OR3 (N785, N784, N532, N772);
buf BUF1 (N786, N515);
nand NAND2 (N787, N783, N369);
xor XOR2 (N788, N777, N137);
buf BUF1 (N789, N760);
nand NAND3 (N790, N787, N753, N424);
not NOT1 (N791, N773);
or OR4 (N792, N781, N674, N606, N147);
nand NAND2 (N793, N788, N554);
buf BUF1 (N794, N778);
not NOT1 (N795, N786);
buf BUF1 (N796, N795);
nand NAND2 (N797, N790, N234);
or OR4 (N798, N792, N758, N759, N785);
xor XOR2 (N799, N30, N236);
and AND4 (N800, N798, N41, N539, N7);
nand NAND4 (N801, N796, N196, N82, N385);
nand NAND3 (N802, N794, N360, N414);
or OR2 (N803, N802, N291);
and AND4 (N804, N793, N99, N567, N418);
not NOT1 (N805, N775);
nor NOR2 (N806, N769, N796);
nand NAND2 (N807, N789, N689);
and AND4 (N808, N799, N378, N541, N651);
not NOT1 (N809, N803);
xor XOR2 (N810, N804, N720);
not NOT1 (N811, N797);
not NOT1 (N812, N807);
and AND3 (N813, N801, N569, N626);
xor XOR2 (N814, N805, N270);
and AND3 (N815, N813, N738, N712);
nor NOR4 (N816, N800, N534, N424, N494);
not NOT1 (N817, N791);
buf BUF1 (N818, N806);
nand NAND3 (N819, N810, N430, N707);
nor NOR2 (N820, N809, N52);
and AND3 (N821, N816, N711, N34);
xor XOR2 (N822, N819, N561);
nor NOR4 (N823, N822, N782, N694, N268);
nand NAND2 (N824, N811, N447);
xor XOR2 (N825, N817, N559);
or OR2 (N826, N808, N773);
nand NAND2 (N827, N818, N648);
buf BUF1 (N828, N820);
not NOT1 (N829, N823);
and AND2 (N830, N828, N689);
nor NOR4 (N831, N814, N124, N94, N577);
nor NOR4 (N832, N815, N24, N231, N653);
nor NOR2 (N833, N827, N495);
nor NOR3 (N834, N830, N742, N461);
or OR2 (N835, N826, N45);
not NOT1 (N836, N824);
and AND3 (N837, N833, N750, N270);
nand NAND3 (N838, N821, N664, N159);
or OR3 (N839, N834, N697, N16);
xor XOR2 (N840, N825, N25);
xor XOR2 (N841, N829, N804);
not NOT1 (N842, N838);
and AND4 (N843, N842, N224, N561, N448);
nor NOR2 (N844, N840, N322);
buf BUF1 (N845, N836);
buf BUF1 (N846, N841);
buf BUF1 (N847, N846);
nand NAND4 (N848, N835, N143, N534, N208);
nand NAND2 (N849, N812, N516);
and AND2 (N850, N848, N421);
xor XOR2 (N851, N831, N586);
nand NAND2 (N852, N845, N342);
xor XOR2 (N853, N837, N464);
nand NAND4 (N854, N847, N581, N123, N101);
and AND2 (N855, N849, N87);
or OR3 (N856, N852, N76, N610);
nor NOR3 (N857, N844, N105, N143);
and AND4 (N858, N855, N204, N577, N293);
or OR2 (N859, N858, N86);
nor NOR2 (N860, N854, N513);
nor NOR4 (N861, N850, N345, N225, N266);
and AND4 (N862, N843, N215, N56, N344);
nand NAND3 (N863, N832, N64, N291);
and AND3 (N864, N857, N147, N448);
nand NAND2 (N865, N859, N67);
xor XOR2 (N866, N853, N845);
buf BUF1 (N867, N860);
nor NOR2 (N868, N856, N615);
not NOT1 (N869, N865);
or OR2 (N870, N861, N602);
and AND2 (N871, N839, N832);
and AND2 (N872, N864, N683);
xor XOR2 (N873, N863, N222);
and AND4 (N874, N851, N408, N227, N695);
nor NOR3 (N875, N873, N488, N248);
nand NAND4 (N876, N862, N678, N665, N347);
or OR4 (N877, N869, N237, N289, N201);
nor NOR2 (N878, N867, N358);
xor XOR2 (N879, N871, N408);
nor NOR3 (N880, N866, N294, N379);
or OR2 (N881, N876, N164);
not NOT1 (N882, N875);
nand NAND2 (N883, N872, N772);
not NOT1 (N884, N878);
not NOT1 (N885, N882);
nor NOR2 (N886, N877, N437);
not NOT1 (N887, N881);
nand NAND4 (N888, N868, N118, N869, N251);
or OR3 (N889, N874, N251, N649);
and AND3 (N890, N889, N50, N278);
xor XOR2 (N891, N890, N463);
xor XOR2 (N892, N870, N402);
nand NAND2 (N893, N879, N735);
and AND2 (N894, N888, N296);
or OR4 (N895, N894, N603, N885, N193);
and AND4 (N896, N558, N642, N827, N684);
xor XOR2 (N897, N886, N276);
nand NAND2 (N898, N896, N86);
or OR4 (N899, N880, N243, N841, N320);
nor NOR3 (N900, N895, N428, N700);
and AND4 (N901, N887, N347, N788, N58);
buf BUF1 (N902, N884);
nor NOR3 (N903, N891, N91, N367);
nor NOR4 (N904, N902, N176, N708, N504);
nand NAND4 (N905, N893, N893, N598, N226);
xor XOR2 (N906, N903, N546);
nor NOR2 (N907, N901, N197);
nor NOR2 (N908, N905, N281);
and AND3 (N909, N900, N249, N107);
not NOT1 (N910, N907);
and AND4 (N911, N910, N223, N25, N463);
and AND4 (N912, N899, N807, N617, N272);
nor NOR2 (N913, N906, N376);
and AND2 (N914, N909, N611);
not NOT1 (N915, N911);
or OR4 (N916, N913, N576, N101, N457);
or OR3 (N917, N898, N582, N615);
and AND3 (N918, N914, N437, N469);
not NOT1 (N919, N912);
and AND2 (N920, N917, N296);
nand NAND4 (N921, N920, N239, N532, N526);
or OR3 (N922, N921, N21, N36);
buf BUF1 (N923, N883);
or OR3 (N924, N897, N207, N622);
xor XOR2 (N925, N923, N713);
xor XOR2 (N926, N919, N271);
xor XOR2 (N927, N924, N797);
xor XOR2 (N928, N922, N564);
not NOT1 (N929, N904);
or OR3 (N930, N908, N888, N28);
not NOT1 (N931, N928);
nor NOR2 (N932, N926, N408);
xor XOR2 (N933, N929, N575);
or OR3 (N934, N918, N138, N735);
or OR4 (N935, N932, N93, N344, N798);
xor XOR2 (N936, N916, N544);
buf BUF1 (N937, N931);
nor NOR3 (N938, N925, N148, N771);
nand NAND4 (N939, N915, N860, N94, N842);
not NOT1 (N940, N930);
nor NOR2 (N941, N936, N106);
xor XOR2 (N942, N939, N15);
and AND3 (N943, N938, N638, N464);
nand NAND3 (N944, N892, N235, N682);
nor NOR3 (N945, N944, N912, N609);
buf BUF1 (N946, N933);
buf BUF1 (N947, N927);
nand NAND4 (N948, N947, N135, N790, N44);
not NOT1 (N949, N943);
buf BUF1 (N950, N946);
not NOT1 (N951, N934);
nand NAND4 (N952, N941, N929, N578, N799);
or OR3 (N953, N945, N36, N160);
nor NOR2 (N954, N940, N114);
not NOT1 (N955, N935);
nand NAND4 (N956, N950, N849, N290, N196);
nor NOR4 (N957, N953, N775, N901, N511);
xor XOR2 (N958, N952, N330);
nor NOR4 (N959, N954, N599, N721, N610);
not NOT1 (N960, N948);
nor NOR3 (N961, N956, N513, N692);
not NOT1 (N962, N937);
and AND2 (N963, N951, N282);
buf BUF1 (N964, N963);
xor XOR2 (N965, N960, N747);
and AND4 (N966, N942, N275, N298, N602);
buf BUF1 (N967, N957);
buf BUF1 (N968, N958);
nor NOR4 (N969, N962, N586, N898, N716);
not NOT1 (N970, N968);
xor XOR2 (N971, N955, N568);
nand NAND3 (N972, N949, N965, N577);
buf BUF1 (N973, N619);
buf BUF1 (N974, N973);
xor XOR2 (N975, N970, N794);
not NOT1 (N976, N975);
and AND4 (N977, N967, N722, N57, N606);
and AND3 (N978, N972, N974, N424);
nor NOR3 (N979, N30, N333, N662);
nand NAND4 (N980, N969, N477, N231, N947);
xor XOR2 (N981, N971, N808);
buf BUF1 (N982, N961);
buf BUF1 (N983, N978);
buf BUF1 (N984, N977);
xor XOR2 (N985, N959, N667);
xor XOR2 (N986, N979, N902);
not NOT1 (N987, N981);
buf BUF1 (N988, N980);
or OR2 (N989, N983, N527);
not NOT1 (N990, N984);
xor XOR2 (N991, N988, N6);
or OR2 (N992, N991, N772);
buf BUF1 (N993, N987);
nor NOR3 (N994, N966, N223, N262);
xor XOR2 (N995, N993, N758);
buf BUF1 (N996, N990);
not NOT1 (N997, N989);
xor XOR2 (N998, N976, N318);
and AND4 (N999, N986, N998, N860, N992);
and AND2 (N1000, N180, N418);
nand NAND2 (N1001, N152, N938);
and AND4 (N1002, N999, N137, N608, N595);
nand NAND3 (N1003, N996, N749, N38);
buf BUF1 (N1004, N985);
xor XOR2 (N1005, N997, N66);
not NOT1 (N1006, N1004);
and AND2 (N1007, N1006, N215);
and AND4 (N1008, N1005, N660, N92, N172);
nor NOR2 (N1009, N1001, N466);
and AND2 (N1010, N982, N480);
xor XOR2 (N1011, N994, N960);
nand NAND3 (N1012, N964, N988, N868);
xor XOR2 (N1013, N1002, N649);
xor XOR2 (N1014, N1010, N396);
xor XOR2 (N1015, N1008, N771);
buf BUF1 (N1016, N1003);
xor XOR2 (N1017, N1000, N903);
nor NOR2 (N1018, N1012, N315);
and AND2 (N1019, N1009, N519);
xor XOR2 (N1020, N1018, N5);
xor XOR2 (N1021, N1020, N569);
and AND4 (N1022, N1017, N934, N703, N138);
not NOT1 (N1023, N1019);
nor NOR2 (N1024, N1021, N317);
not NOT1 (N1025, N1015);
buf BUF1 (N1026, N1014);
buf BUF1 (N1027, N1022);
xor XOR2 (N1028, N995, N13);
nand NAND4 (N1029, N1007, N288, N632, N1010);
nor NOR4 (N1030, N1029, N963, N70, N1027);
nand NAND4 (N1031, N497, N392, N39, N900);
not NOT1 (N1032, N1026);
buf BUF1 (N1033, N1028);
nor NOR4 (N1034, N1032, N649, N854, N149);
xor XOR2 (N1035, N1025, N469);
not NOT1 (N1036, N1035);
not NOT1 (N1037, N1023);
and AND3 (N1038, N1034, N162, N184);
or OR3 (N1039, N1037, N679, N486);
buf BUF1 (N1040, N1031);
nand NAND2 (N1041, N1039, N876);
not NOT1 (N1042, N1030);
xor XOR2 (N1043, N1024, N504);
xor XOR2 (N1044, N1040, N198);
nor NOR3 (N1045, N1044, N475, N535);
and AND2 (N1046, N1041, N106);
buf BUF1 (N1047, N1013);
or OR4 (N1048, N1036, N240, N824, N256);
or OR3 (N1049, N1016, N944, N636);
nor NOR2 (N1050, N1038, N930);
nor NOR3 (N1051, N1048, N44, N909);
nor NOR4 (N1052, N1049, N1019, N635, N347);
nor NOR2 (N1053, N1052, N504);
buf BUF1 (N1054, N1046);
xor XOR2 (N1055, N1051, N1006);
or OR3 (N1056, N1047, N580, N782);
buf BUF1 (N1057, N1011);
or OR4 (N1058, N1053, N869, N420, N788);
nand NAND3 (N1059, N1043, N590, N686);
nor NOR4 (N1060, N1045, N933, N294, N1050);
not NOT1 (N1061, N201);
nor NOR2 (N1062, N1060, N249);
xor XOR2 (N1063, N1059, N904);
nor NOR4 (N1064, N1033, N672, N594, N834);
buf BUF1 (N1065, N1061);
or OR3 (N1066, N1054, N105, N434);
nor NOR2 (N1067, N1042, N866);
and AND2 (N1068, N1062, N513);
not NOT1 (N1069, N1068);
nand NAND2 (N1070, N1063, N751);
xor XOR2 (N1071, N1058, N86);
buf BUF1 (N1072, N1064);
not NOT1 (N1073, N1056);
nor NOR4 (N1074, N1066, N308, N328, N311);
buf BUF1 (N1075, N1065);
buf BUF1 (N1076, N1071);
and AND4 (N1077, N1070, N494, N604, N662);
not NOT1 (N1078, N1072);
and AND4 (N1079, N1075, N10, N454, N820);
nor NOR3 (N1080, N1076, N970, N194);
nor NOR3 (N1081, N1077, N399, N594);
and AND4 (N1082, N1081, N471, N258, N877);
buf BUF1 (N1083, N1055);
buf BUF1 (N1084, N1073);
xor XOR2 (N1085, N1074, N512);
or OR3 (N1086, N1080, N44, N863);
or OR2 (N1087, N1057, N1004);
buf BUF1 (N1088, N1082);
and AND4 (N1089, N1067, N978, N50, N851);
or OR4 (N1090, N1088, N573, N1074, N764);
or OR4 (N1091, N1085, N218, N100, N42);
nor NOR4 (N1092, N1069, N499, N619, N870);
not NOT1 (N1093, N1091);
nor NOR4 (N1094, N1089, N865, N506, N284);
nand NAND2 (N1095, N1078, N827);
not NOT1 (N1096, N1093);
xor XOR2 (N1097, N1087, N153);
buf BUF1 (N1098, N1084);
and AND3 (N1099, N1096, N480, N468);
and AND4 (N1100, N1090, N431, N414, N700);
xor XOR2 (N1101, N1079, N1010);
buf BUF1 (N1102, N1100);
or OR3 (N1103, N1097, N644, N644);
nand NAND4 (N1104, N1099, N268, N835, N294);
xor XOR2 (N1105, N1102, N303);
xor XOR2 (N1106, N1094, N606);
and AND4 (N1107, N1101, N804, N641, N182);
and AND2 (N1108, N1107, N406);
or OR3 (N1109, N1095, N163, N569);
or OR4 (N1110, N1108, N283, N714, N236);
nor NOR2 (N1111, N1106, N942);
nand NAND3 (N1112, N1105, N1045, N953);
not NOT1 (N1113, N1111);
nor NOR4 (N1114, N1113, N651, N74, N1039);
xor XOR2 (N1115, N1110, N677);
nand NAND2 (N1116, N1114, N578);
buf BUF1 (N1117, N1109);
nand NAND4 (N1118, N1104, N541, N665, N1073);
nand NAND2 (N1119, N1098, N362);
nor NOR2 (N1120, N1115, N219);
not NOT1 (N1121, N1092);
and AND4 (N1122, N1083, N583, N126, N102);
nand NAND3 (N1123, N1112, N926, N1081);
not NOT1 (N1124, N1116);
or OR4 (N1125, N1120, N288, N524, N975);
not NOT1 (N1126, N1123);
nor NOR2 (N1127, N1103, N292);
and AND4 (N1128, N1127, N465, N1020, N564);
or OR4 (N1129, N1119, N635, N753, N448);
buf BUF1 (N1130, N1126);
and AND3 (N1131, N1124, N1059, N265);
nor NOR4 (N1132, N1125, N1073, N443, N54);
not NOT1 (N1133, N1132);
xor XOR2 (N1134, N1121, N577);
and AND2 (N1135, N1134, N112);
nor NOR2 (N1136, N1130, N341);
nand NAND4 (N1137, N1131, N480, N746, N931);
nor NOR4 (N1138, N1122, N844, N9, N1050);
not NOT1 (N1139, N1128);
not NOT1 (N1140, N1136);
buf BUF1 (N1141, N1086);
xor XOR2 (N1142, N1117, N827);
not NOT1 (N1143, N1137);
and AND2 (N1144, N1142, N288);
and AND2 (N1145, N1133, N524);
buf BUF1 (N1146, N1141);
and AND3 (N1147, N1143, N262, N707);
not NOT1 (N1148, N1135);
and AND3 (N1149, N1144, N479, N725);
xor XOR2 (N1150, N1138, N556);
nor NOR4 (N1151, N1149, N78, N425, N1123);
nand NAND3 (N1152, N1148, N174, N194);
or OR3 (N1153, N1147, N322, N313);
nor NOR4 (N1154, N1145, N282, N1118, N1120);
xor XOR2 (N1155, N109, N841);
buf BUF1 (N1156, N1151);
or OR2 (N1157, N1129, N365);
nand NAND2 (N1158, N1154, N1104);
nor NOR2 (N1159, N1146, N935);
nand NAND2 (N1160, N1140, N740);
xor XOR2 (N1161, N1152, N919);
nor NOR3 (N1162, N1155, N505, N989);
not NOT1 (N1163, N1158);
or OR3 (N1164, N1162, N943, N718);
buf BUF1 (N1165, N1160);
nor NOR3 (N1166, N1163, N375, N410);
nand NAND3 (N1167, N1166, N334, N676);
or OR4 (N1168, N1157, N579, N400, N281);
nand NAND3 (N1169, N1139, N842, N306);
not NOT1 (N1170, N1156);
nor NOR2 (N1171, N1170, N1079);
nor NOR4 (N1172, N1167, N531, N203, N778);
buf BUF1 (N1173, N1161);
xor XOR2 (N1174, N1159, N257);
nor NOR3 (N1175, N1173, N692, N676);
xor XOR2 (N1176, N1150, N51);
nand NAND2 (N1177, N1175, N133);
and AND2 (N1178, N1165, N572);
nor NOR4 (N1179, N1178, N975, N1176, N211);
and AND2 (N1180, N670, N526);
xor XOR2 (N1181, N1153, N810);
nor NOR2 (N1182, N1179, N860);
nand NAND2 (N1183, N1174, N346);
buf BUF1 (N1184, N1164);
or OR3 (N1185, N1172, N90, N923);
or OR3 (N1186, N1183, N345, N645);
buf BUF1 (N1187, N1169);
not NOT1 (N1188, N1181);
buf BUF1 (N1189, N1177);
nand NAND4 (N1190, N1182, N649, N613, N115);
nand NAND2 (N1191, N1180, N1185);
or OR2 (N1192, N750, N754);
buf BUF1 (N1193, N1189);
nand NAND4 (N1194, N1192, N720, N1090, N845);
nor NOR4 (N1195, N1171, N682, N444, N439);
not NOT1 (N1196, N1188);
nand NAND2 (N1197, N1196, N231);
or OR4 (N1198, N1184, N301, N220, N491);
buf BUF1 (N1199, N1168);
nor NOR2 (N1200, N1190, N946);
or OR3 (N1201, N1187, N236, N723);
not NOT1 (N1202, N1193);
buf BUF1 (N1203, N1199);
nand NAND4 (N1204, N1186, N597, N835, N419);
xor XOR2 (N1205, N1198, N260);
nor NOR4 (N1206, N1204, N636, N377, N1203);
and AND4 (N1207, N67, N333, N425, N787);
not NOT1 (N1208, N1191);
and AND2 (N1209, N1195, N163);
buf BUF1 (N1210, N1207);
buf BUF1 (N1211, N1206);
nand NAND2 (N1212, N1201, N1202);
nor NOR4 (N1213, N19, N308, N916, N234);
xor XOR2 (N1214, N1209, N175);
or OR3 (N1215, N1214, N1076, N127);
buf BUF1 (N1216, N1211);
nand NAND4 (N1217, N1208, N709, N1017, N1150);
nor NOR4 (N1218, N1200, N505, N427, N746);
nor NOR3 (N1219, N1217, N576, N1047);
not NOT1 (N1220, N1215);
buf BUF1 (N1221, N1218);
or OR3 (N1222, N1197, N1132, N576);
nand NAND3 (N1223, N1213, N956, N44);
buf BUF1 (N1224, N1205);
not NOT1 (N1225, N1210);
buf BUF1 (N1226, N1222);
nand NAND4 (N1227, N1219, N532, N938, N664);
and AND2 (N1228, N1221, N403);
buf BUF1 (N1229, N1228);
buf BUF1 (N1230, N1227);
nand NAND3 (N1231, N1226, N1034, N948);
not NOT1 (N1232, N1229);
xor XOR2 (N1233, N1194, N912);
xor XOR2 (N1234, N1224, N248);
nor NOR3 (N1235, N1223, N55, N665);
or OR3 (N1236, N1233, N872, N903);
nor NOR4 (N1237, N1232, N330, N595, N552);
or OR3 (N1238, N1235, N282, N906);
or OR4 (N1239, N1231, N964, N902, N283);
nor NOR4 (N1240, N1220, N466, N1043, N505);
nor NOR4 (N1241, N1238, N137, N365, N592);
nand NAND2 (N1242, N1240, N1075);
not NOT1 (N1243, N1230);
nor NOR3 (N1244, N1212, N31, N743);
or OR3 (N1245, N1239, N1135, N771);
not NOT1 (N1246, N1244);
nand NAND3 (N1247, N1225, N1100, N185);
nand NAND3 (N1248, N1237, N760, N858);
xor XOR2 (N1249, N1216, N579);
or OR2 (N1250, N1247, N409);
nand NAND4 (N1251, N1234, N27, N860, N806);
not NOT1 (N1252, N1250);
xor XOR2 (N1253, N1251, N942);
buf BUF1 (N1254, N1248);
not NOT1 (N1255, N1252);
nor NOR4 (N1256, N1254, N557, N773, N987);
not NOT1 (N1257, N1256);
buf BUF1 (N1258, N1241);
nor NOR4 (N1259, N1258, N224, N721, N1244);
or OR4 (N1260, N1257, N479, N593, N1019);
nor NOR3 (N1261, N1255, N551, N308);
and AND2 (N1262, N1245, N877);
nand NAND3 (N1263, N1261, N668, N1122);
or OR3 (N1264, N1259, N640, N518);
nand NAND4 (N1265, N1260, N1130, N627, N1212);
nor NOR3 (N1266, N1242, N561, N77);
buf BUF1 (N1267, N1243);
not NOT1 (N1268, N1263);
nor NOR4 (N1269, N1236, N725, N1148, N1172);
or OR2 (N1270, N1264, N1266);
and AND2 (N1271, N1151, N900);
and AND4 (N1272, N1271, N575, N271, N335);
and AND3 (N1273, N1269, N181, N103);
or OR3 (N1274, N1262, N845, N987);
nand NAND2 (N1275, N1253, N75);
or OR4 (N1276, N1249, N1011, N435, N545);
nor NOR2 (N1277, N1276, N411);
nor NOR4 (N1278, N1268, N176, N864, N18);
and AND2 (N1279, N1274, N945);
not NOT1 (N1280, N1265);
or OR4 (N1281, N1270, N97, N283, N754);
xor XOR2 (N1282, N1273, N740);
or OR4 (N1283, N1267, N586, N1159, N184);
nand NAND3 (N1284, N1272, N369, N789);
not NOT1 (N1285, N1281);
not NOT1 (N1286, N1246);
nor NOR4 (N1287, N1284, N988, N1055, N34);
nand NAND4 (N1288, N1282, N609, N583, N329);
and AND2 (N1289, N1286, N452);
xor XOR2 (N1290, N1275, N634);
buf BUF1 (N1291, N1280);
nand NAND2 (N1292, N1278, N1106);
or OR2 (N1293, N1277, N108);
not NOT1 (N1294, N1279);
not NOT1 (N1295, N1293);
nand NAND3 (N1296, N1295, N930, N1177);
xor XOR2 (N1297, N1285, N785);
and AND3 (N1298, N1297, N417, N540);
nand NAND4 (N1299, N1287, N782, N474, N1256);
nand NAND2 (N1300, N1290, N1065);
buf BUF1 (N1301, N1289);
not NOT1 (N1302, N1291);
xor XOR2 (N1303, N1298, N841);
nor NOR4 (N1304, N1302, N516, N381, N545);
and AND3 (N1305, N1304, N1241, N946);
xor XOR2 (N1306, N1299, N1105);
and AND4 (N1307, N1301, N528, N688, N965);
or OR4 (N1308, N1292, N281, N910, N1056);
or OR2 (N1309, N1296, N591);
buf BUF1 (N1310, N1283);
buf BUF1 (N1311, N1305);
nor NOR3 (N1312, N1310, N678, N872);
or OR2 (N1313, N1306, N508);
not NOT1 (N1314, N1308);
nand NAND3 (N1315, N1303, N66, N1147);
nand NAND3 (N1316, N1313, N235, N701);
and AND3 (N1317, N1316, N905, N333);
and AND2 (N1318, N1307, N46);
not NOT1 (N1319, N1309);
buf BUF1 (N1320, N1300);
buf BUF1 (N1321, N1312);
buf BUF1 (N1322, N1294);
not NOT1 (N1323, N1319);
and AND2 (N1324, N1314, N1152);
nand NAND4 (N1325, N1315, N1003, N1088, N1318);
or OR3 (N1326, N359, N869, N50);
nand NAND4 (N1327, N1326, N222, N315, N391);
and AND4 (N1328, N1327, N1320, N287, N675);
nand NAND2 (N1329, N9, N1192);
xor XOR2 (N1330, N1311, N473);
nand NAND4 (N1331, N1324, N892, N559, N1092);
xor XOR2 (N1332, N1330, N1194);
nor NOR3 (N1333, N1288, N1068, N716);
nor NOR2 (N1334, N1329, N76);
nand NAND3 (N1335, N1328, N486, N480);
xor XOR2 (N1336, N1334, N559);
xor XOR2 (N1337, N1317, N985);
nand NAND4 (N1338, N1323, N789, N262, N679);
nor NOR2 (N1339, N1321, N1050);
nand NAND3 (N1340, N1325, N786, N41);
buf BUF1 (N1341, N1339);
nand NAND2 (N1342, N1338, N1186);
nand NAND4 (N1343, N1333, N339, N696, N1057);
and AND3 (N1344, N1332, N997, N26);
not NOT1 (N1345, N1340);
buf BUF1 (N1346, N1331);
or OR4 (N1347, N1342, N874, N756, N601);
or OR4 (N1348, N1346, N1142, N486, N270);
nor NOR2 (N1349, N1343, N747);
not NOT1 (N1350, N1348);
not NOT1 (N1351, N1344);
and AND2 (N1352, N1337, N1193);
not NOT1 (N1353, N1352);
nor NOR4 (N1354, N1349, N881, N736, N504);
and AND3 (N1355, N1354, N659, N434);
xor XOR2 (N1356, N1345, N177);
nor NOR3 (N1357, N1335, N99, N209);
and AND4 (N1358, N1336, N930, N976, N1005);
nand NAND3 (N1359, N1355, N891, N961);
buf BUF1 (N1360, N1347);
xor XOR2 (N1361, N1351, N310);
nand NAND2 (N1362, N1361, N941);
and AND2 (N1363, N1359, N1276);
or OR3 (N1364, N1356, N416, N1188);
nand NAND3 (N1365, N1322, N579, N939);
xor XOR2 (N1366, N1363, N1086);
nand NAND2 (N1367, N1358, N548);
nand NAND3 (N1368, N1364, N678, N543);
not NOT1 (N1369, N1362);
buf BUF1 (N1370, N1368);
xor XOR2 (N1371, N1366, N506);
and AND4 (N1372, N1341, N289, N181, N562);
not NOT1 (N1373, N1350);
nand NAND4 (N1374, N1373, N358, N556, N823);
not NOT1 (N1375, N1367);
nand NAND2 (N1376, N1374, N650);
xor XOR2 (N1377, N1353, N1119);
nor NOR2 (N1378, N1376, N327);
nand NAND3 (N1379, N1372, N94, N183);
nor NOR3 (N1380, N1375, N1340, N203);
or OR4 (N1381, N1357, N162, N245, N519);
not NOT1 (N1382, N1370);
xor XOR2 (N1383, N1381, N1115);
and AND3 (N1384, N1377, N440, N1005);
and AND2 (N1385, N1365, N1219);
and AND4 (N1386, N1360, N1302, N1261, N382);
xor XOR2 (N1387, N1379, N327);
or OR2 (N1388, N1387, N730);
nor NOR2 (N1389, N1369, N666);
nor NOR4 (N1390, N1384, N877, N11, N299);
buf BUF1 (N1391, N1388);
xor XOR2 (N1392, N1382, N506);
nor NOR4 (N1393, N1378, N303, N754, N1046);
buf BUF1 (N1394, N1393);
or OR3 (N1395, N1394, N564, N293);
or OR2 (N1396, N1391, N2);
nor NOR3 (N1397, N1380, N990, N659);
and AND3 (N1398, N1383, N231, N149);
nor NOR4 (N1399, N1395, N414, N804, N533);
and AND4 (N1400, N1398, N6, N1359, N1061);
nor NOR3 (N1401, N1389, N262, N1141);
buf BUF1 (N1402, N1396);
nor NOR4 (N1403, N1402, N388, N1171, N1385);
or OR4 (N1404, N1076, N428, N784, N672);
nand NAND4 (N1405, N1371, N574, N623, N643);
buf BUF1 (N1406, N1397);
and AND4 (N1407, N1392, N723, N868, N974);
buf BUF1 (N1408, N1407);
nor NOR4 (N1409, N1405, N565, N762, N421);
buf BUF1 (N1410, N1401);
or OR3 (N1411, N1406, N243, N418);
or OR3 (N1412, N1390, N986, N233);
buf BUF1 (N1413, N1400);
not NOT1 (N1414, N1403);
buf BUF1 (N1415, N1412);
xor XOR2 (N1416, N1408, N267);
or OR2 (N1417, N1415, N1396);
buf BUF1 (N1418, N1411);
xor XOR2 (N1419, N1404, N289);
and AND3 (N1420, N1410, N1339, N620);
not NOT1 (N1421, N1413);
or OR2 (N1422, N1416, N285);
not NOT1 (N1423, N1420);
or OR2 (N1424, N1418, N168);
buf BUF1 (N1425, N1386);
xor XOR2 (N1426, N1424, N368);
and AND4 (N1427, N1399, N648, N594, N244);
and AND3 (N1428, N1414, N1186, N1186);
buf BUF1 (N1429, N1425);
or OR2 (N1430, N1409, N994);
nor NOR3 (N1431, N1427, N288, N796);
not NOT1 (N1432, N1423);
or OR3 (N1433, N1429, N1279, N190);
nand NAND3 (N1434, N1431, N356, N1122);
nor NOR2 (N1435, N1422, N774);
xor XOR2 (N1436, N1432, N2);
nand NAND3 (N1437, N1430, N514, N1036);
nand NAND2 (N1438, N1433, N612);
and AND2 (N1439, N1428, N530);
buf BUF1 (N1440, N1419);
not NOT1 (N1441, N1417);
nand NAND3 (N1442, N1438, N170, N1288);
and AND3 (N1443, N1434, N850, N236);
xor XOR2 (N1444, N1441, N1154);
buf BUF1 (N1445, N1421);
or OR3 (N1446, N1436, N1283, N682);
buf BUF1 (N1447, N1446);
and AND2 (N1448, N1440, N1407);
and AND3 (N1449, N1444, N930, N505);
or OR3 (N1450, N1439, N449, N299);
nor NOR3 (N1451, N1448, N1292, N1071);
not NOT1 (N1452, N1449);
nor NOR4 (N1453, N1435, N53, N452, N893);
and AND3 (N1454, N1443, N821, N688);
not NOT1 (N1455, N1445);
nand NAND2 (N1456, N1454, N745);
or OR4 (N1457, N1450, N521, N897, N1169);
buf BUF1 (N1458, N1452);
xor XOR2 (N1459, N1453, N1354);
or OR3 (N1460, N1458, N1305, N1345);
xor XOR2 (N1461, N1457, N470);
not NOT1 (N1462, N1426);
not NOT1 (N1463, N1462);
nand NAND4 (N1464, N1442, N1159, N938, N685);
and AND4 (N1465, N1463, N569, N1100, N623);
nand NAND3 (N1466, N1456, N1376, N144);
nand NAND4 (N1467, N1451, N760, N1109, N772);
not NOT1 (N1468, N1465);
not NOT1 (N1469, N1447);
or OR4 (N1470, N1466, N269, N626, N190);
or OR3 (N1471, N1469, N1445, N1084);
xor XOR2 (N1472, N1470, N975);
or OR4 (N1473, N1472, N1264, N197, N1444);
nor NOR2 (N1474, N1461, N388);
buf BUF1 (N1475, N1474);
nand NAND3 (N1476, N1437, N578, N719);
not NOT1 (N1477, N1475);
nor NOR4 (N1478, N1467, N252, N603, N1226);
nor NOR4 (N1479, N1464, N344, N737, N658);
and AND4 (N1480, N1476, N173, N1312, N73);
and AND3 (N1481, N1480, N78, N1102);
buf BUF1 (N1482, N1459);
buf BUF1 (N1483, N1482);
xor XOR2 (N1484, N1479, N745);
or OR2 (N1485, N1460, N1088);
or OR4 (N1486, N1485, N228, N385, N1045);
and AND4 (N1487, N1486, N471, N792, N391);
not NOT1 (N1488, N1478);
nor NOR2 (N1489, N1455, N1114);
nor NOR3 (N1490, N1468, N245, N1429);
buf BUF1 (N1491, N1483);
xor XOR2 (N1492, N1488, N347);
buf BUF1 (N1493, N1473);
xor XOR2 (N1494, N1481, N279);
nand NAND2 (N1495, N1471, N592);
buf BUF1 (N1496, N1493);
nand NAND2 (N1497, N1491, N1050);
and AND4 (N1498, N1489, N1460, N472, N886);
xor XOR2 (N1499, N1487, N1122);
xor XOR2 (N1500, N1495, N890);
or OR3 (N1501, N1498, N839, N995);
and AND2 (N1502, N1501, N865);
xor XOR2 (N1503, N1502, N1449);
and AND2 (N1504, N1494, N879);
xor XOR2 (N1505, N1492, N645);
not NOT1 (N1506, N1505);
xor XOR2 (N1507, N1503, N299);
xor XOR2 (N1508, N1500, N481);
and AND2 (N1509, N1496, N1434);
xor XOR2 (N1510, N1504, N799);
xor XOR2 (N1511, N1508, N359);
nand NAND3 (N1512, N1499, N294, N1400);
and AND3 (N1513, N1509, N1311, N391);
xor XOR2 (N1514, N1490, N616);
not NOT1 (N1515, N1514);
or OR4 (N1516, N1515, N46, N1050, N118);
not NOT1 (N1517, N1497);
buf BUF1 (N1518, N1477);
xor XOR2 (N1519, N1511, N429);
or OR2 (N1520, N1510, N1134);
not NOT1 (N1521, N1484);
or OR3 (N1522, N1512, N1037, N244);
and AND2 (N1523, N1517, N904);
xor XOR2 (N1524, N1523, N426);
buf BUF1 (N1525, N1518);
not NOT1 (N1526, N1524);
not NOT1 (N1527, N1521);
buf BUF1 (N1528, N1519);
and AND3 (N1529, N1520, N1198, N1440);
xor XOR2 (N1530, N1527, N183);
and AND3 (N1531, N1513, N570, N898);
or OR4 (N1532, N1507, N46, N775, N680);
nor NOR3 (N1533, N1532, N1436, N449);
or OR3 (N1534, N1528, N405, N1084);
nand NAND4 (N1535, N1516, N304, N502, N686);
buf BUF1 (N1536, N1529);
nor NOR3 (N1537, N1526, N1032, N405);
nand NAND4 (N1538, N1535, N687, N1208, N528);
nand NAND4 (N1539, N1506, N909, N1330, N1026);
or OR2 (N1540, N1534, N135);
nor NOR3 (N1541, N1530, N23, N1);
buf BUF1 (N1542, N1531);
nand NAND3 (N1543, N1536, N1309, N952);
nor NOR3 (N1544, N1525, N948, N183);
or OR4 (N1545, N1541, N790, N1214, N947);
buf BUF1 (N1546, N1537);
nand NAND2 (N1547, N1522, N1190);
not NOT1 (N1548, N1547);
nand NAND2 (N1549, N1545, N527);
and AND3 (N1550, N1533, N1387, N489);
nand NAND3 (N1551, N1540, N261, N197);
not NOT1 (N1552, N1544);
xor XOR2 (N1553, N1542, N926);
nor NOR2 (N1554, N1546, N1030);
and AND3 (N1555, N1543, N1548, N1501);
nor NOR2 (N1556, N909, N1252);
nand NAND3 (N1557, N1550, N594, N778);
or OR3 (N1558, N1551, N976, N1469);
buf BUF1 (N1559, N1549);
nand NAND2 (N1560, N1539, N197);
or OR2 (N1561, N1554, N233);
and AND4 (N1562, N1560, N1050, N781, N320);
buf BUF1 (N1563, N1538);
buf BUF1 (N1564, N1562);
or OR2 (N1565, N1557, N260);
not NOT1 (N1566, N1559);
and AND4 (N1567, N1565, N1222, N1010, N796);
nand NAND4 (N1568, N1556, N1456, N349, N1360);
and AND2 (N1569, N1561, N738);
and AND3 (N1570, N1552, N35, N619);
xor XOR2 (N1571, N1570, N1014);
buf BUF1 (N1572, N1558);
nor NOR4 (N1573, N1567, N774, N967, N935);
not NOT1 (N1574, N1555);
or OR3 (N1575, N1574, N1218, N1165);
xor XOR2 (N1576, N1568, N1574);
and AND2 (N1577, N1563, N1293);
xor XOR2 (N1578, N1577, N1395);
nor NOR3 (N1579, N1576, N1519, N842);
not NOT1 (N1580, N1578);
nor NOR4 (N1581, N1569, N1152, N73, N1518);
and AND2 (N1582, N1575, N257);
not NOT1 (N1583, N1553);
and AND2 (N1584, N1573, N1442);
buf BUF1 (N1585, N1579);
nand NAND3 (N1586, N1583, N476, N1580);
not NOT1 (N1587, N841);
not NOT1 (N1588, N1572);
nor NOR4 (N1589, N1585, N378, N854, N561);
nor NOR4 (N1590, N1571, N962, N1050, N317);
not NOT1 (N1591, N1581);
not NOT1 (N1592, N1589);
not NOT1 (N1593, N1584);
nand NAND4 (N1594, N1588, N838, N47, N352);
or OR4 (N1595, N1591, N935, N480, N1396);
and AND3 (N1596, N1592, N459, N108);
nand NAND3 (N1597, N1594, N423, N563);
xor XOR2 (N1598, N1597, N1205);
nor NOR3 (N1599, N1593, N503, N322);
nand NAND4 (N1600, N1590, N933, N455, N45);
nand NAND4 (N1601, N1598, N631, N213, N705);
or OR3 (N1602, N1564, N252, N854);
xor XOR2 (N1603, N1601, N1353);
or OR3 (N1604, N1602, N24, N1113);
and AND3 (N1605, N1604, N295, N306);
buf BUF1 (N1606, N1587);
buf BUF1 (N1607, N1599);
nand NAND3 (N1608, N1600, N1149, N662);
buf BUF1 (N1609, N1586);
or OR4 (N1610, N1582, N1074, N190, N260);
nand NAND2 (N1611, N1603, N370);
or OR4 (N1612, N1611, N95, N392, N1180);
not NOT1 (N1613, N1566);
buf BUF1 (N1614, N1607);
or OR4 (N1615, N1596, N953, N1227, N1585);
xor XOR2 (N1616, N1610, N660);
xor XOR2 (N1617, N1606, N194);
nand NAND2 (N1618, N1617, N412);
buf BUF1 (N1619, N1616);
xor XOR2 (N1620, N1613, N50);
or OR2 (N1621, N1614, N1174);
xor XOR2 (N1622, N1595, N983);
or OR3 (N1623, N1608, N1209, N226);
not NOT1 (N1624, N1609);
nor NOR3 (N1625, N1620, N1179, N1607);
and AND3 (N1626, N1623, N554, N196);
or OR2 (N1627, N1612, N175);
not NOT1 (N1628, N1622);
and AND3 (N1629, N1621, N949, N57);
nand NAND4 (N1630, N1625, N1574, N1520, N913);
buf BUF1 (N1631, N1619);
not NOT1 (N1632, N1629);
xor XOR2 (N1633, N1618, N1277);
and AND4 (N1634, N1628, N567, N788, N1038);
not NOT1 (N1635, N1615);
buf BUF1 (N1636, N1627);
nor NOR2 (N1637, N1626, N1338);
and AND4 (N1638, N1634, N168, N1034, N1215);
not NOT1 (N1639, N1638);
xor XOR2 (N1640, N1639, N1491);
xor XOR2 (N1641, N1633, N520);
and AND3 (N1642, N1641, N1177, N1294);
not NOT1 (N1643, N1624);
xor XOR2 (N1644, N1632, N812);
nand NAND4 (N1645, N1631, N652, N306, N1605);
and AND2 (N1646, N695, N1329);
nand NAND3 (N1647, N1645, N16, N91);
and AND3 (N1648, N1643, N1049, N914);
and AND4 (N1649, N1642, N222, N665, N652);
not NOT1 (N1650, N1640);
buf BUF1 (N1651, N1635);
buf BUF1 (N1652, N1648);
buf BUF1 (N1653, N1650);
not NOT1 (N1654, N1646);
buf BUF1 (N1655, N1630);
not NOT1 (N1656, N1654);
or OR3 (N1657, N1652, N305, N1187);
xor XOR2 (N1658, N1653, N659);
or OR4 (N1659, N1658, N1313, N1387, N104);
nand NAND4 (N1660, N1649, N454, N670, N523);
and AND2 (N1661, N1655, N1601);
and AND4 (N1662, N1656, N1633, N626, N1253);
or OR3 (N1663, N1659, N69, N4);
not NOT1 (N1664, N1637);
not NOT1 (N1665, N1647);
and AND2 (N1666, N1662, N1440);
nand NAND3 (N1667, N1665, N1561, N872);
buf BUF1 (N1668, N1636);
buf BUF1 (N1669, N1651);
buf BUF1 (N1670, N1667);
nor NOR3 (N1671, N1644, N1104, N501);
nor NOR4 (N1672, N1666, N24, N1387, N1012);
and AND3 (N1673, N1672, N711, N412);
xor XOR2 (N1674, N1673, N1636);
not NOT1 (N1675, N1671);
xor XOR2 (N1676, N1663, N261);
xor XOR2 (N1677, N1660, N1655);
nor NOR3 (N1678, N1676, N49, N1005);
or OR3 (N1679, N1674, N584, N707);
xor XOR2 (N1680, N1675, N463);
xor XOR2 (N1681, N1669, N1192);
and AND4 (N1682, N1657, N1070, N924, N1537);
or OR3 (N1683, N1682, N1579, N1087);
nor NOR4 (N1684, N1680, N1201, N865, N1520);
xor XOR2 (N1685, N1684, N1385);
buf BUF1 (N1686, N1679);
nor NOR3 (N1687, N1686, N618, N930);
not NOT1 (N1688, N1677);
not NOT1 (N1689, N1668);
or OR4 (N1690, N1661, N805, N1374, N801);
nor NOR4 (N1691, N1690, N1174, N489, N695);
not NOT1 (N1692, N1687);
nand NAND3 (N1693, N1689, N1050, N1567);
and AND4 (N1694, N1681, N1253, N704, N403);
not NOT1 (N1695, N1693);
buf BUF1 (N1696, N1694);
or OR3 (N1697, N1683, N867, N329);
and AND4 (N1698, N1697, N873, N1242, N707);
nand NAND3 (N1699, N1696, N990, N1504);
xor XOR2 (N1700, N1664, N932);
nor NOR4 (N1701, N1685, N1688, N880, N639);
nand NAND2 (N1702, N550, N1461);
nand NAND3 (N1703, N1701, N790, N637);
xor XOR2 (N1704, N1703, N1252);
nor NOR2 (N1705, N1699, N820);
xor XOR2 (N1706, N1678, N588);
xor XOR2 (N1707, N1702, N416);
not NOT1 (N1708, N1698);
and AND4 (N1709, N1695, N1480, N265, N386);
or OR2 (N1710, N1705, N1505);
nand NAND2 (N1711, N1692, N674);
nand NAND3 (N1712, N1700, N1585, N107);
nand NAND4 (N1713, N1670, N253, N1628, N1411);
nor NOR3 (N1714, N1710, N1241, N1018);
and AND2 (N1715, N1713, N956);
nor NOR4 (N1716, N1708, N321, N404, N1592);
or OR2 (N1717, N1709, N179);
nand NAND2 (N1718, N1711, N1046);
and AND2 (N1719, N1717, N574);
nand NAND4 (N1720, N1712, N944, N1378, N633);
nor NOR4 (N1721, N1720, N1703, N1494, N1614);
xor XOR2 (N1722, N1718, N194);
and AND3 (N1723, N1721, N380, N570);
xor XOR2 (N1724, N1722, N562);
or OR2 (N1725, N1714, N1313);
nor NOR4 (N1726, N1691, N973, N737, N1425);
nor NOR4 (N1727, N1724, N246, N721, N1320);
and AND3 (N1728, N1727, N916, N421);
xor XOR2 (N1729, N1726, N541);
nor NOR4 (N1730, N1706, N846, N52, N462);
nand NAND3 (N1731, N1723, N1252, N422);
buf BUF1 (N1732, N1715);
and AND3 (N1733, N1732, N257, N1556);
not NOT1 (N1734, N1704);
and AND3 (N1735, N1730, N835, N647);
buf BUF1 (N1736, N1719);
xor XOR2 (N1737, N1716, N1195);
buf BUF1 (N1738, N1707);
buf BUF1 (N1739, N1738);
nor NOR2 (N1740, N1728, N1365);
and AND2 (N1741, N1733, N729);
nand NAND4 (N1742, N1737, N732, N1526, N1563);
nand NAND4 (N1743, N1739, N1250, N1473, N1666);
nand NAND4 (N1744, N1731, N494, N82, N1053);
and AND3 (N1745, N1742, N162, N678);
and AND2 (N1746, N1744, N1281);
nand NAND3 (N1747, N1729, N74, N710);
xor XOR2 (N1748, N1734, N1003);
and AND4 (N1749, N1743, N835, N1473, N646);
buf BUF1 (N1750, N1745);
not NOT1 (N1751, N1740);
nor NOR2 (N1752, N1747, N108);
or OR3 (N1753, N1741, N1536, N1684);
and AND4 (N1754, N1735, N162, N876, N1566);
buf BUF1 (N1755, N1753);
or OR2 (N1756, N1755, N615);
or OR3 (N1757, N1751, N1294, N489);
and AND2 (N1758, N1725, N1706);
nor NOR2 (N1759, N1754, N451);
nor NOR2 (N1760, N1736, N759);
nor NOR3 (N1761, N1759, N421, N80);
xor XOR2 (N1762, N1752, N477);
or OR3 (N1763, N1750, N848, N679);
or OR4 (N1764, N1761, N950, N896, N1606);
nor NOR4 (N1765, N1749, N1138, N687, N962);
nor NOR4 (N1766, N1756, N919, N1377, N57);
or OR2 (N1767, N1748, N442);
buf BUF1 (N1768, N1766);
not NOT1 (N1769, N1762);
not NOT1 (N1770, N1758);
xor XOR2 (N1771, N1746, N1220);
not NOT1 (N1772, N1765);
nand NAND3 (N1773, N1757, N1099, N332);
nand NAND3 (N1774, N1763, N1576, N1291);
nand NAND2 (N1775, N1760, N458);
buf BUF1 (N1776, N1764);
nand NAND2 (N1777, N1771, N1760);
or OR4 (N1778, N1767, N1064, N163, N823);
nand NAND4 (N1779, N1777, N153, N596, N361);
and AND3 (N1780, N1773, N347, N1698);
not NOT1 (N1781, N1779);
or OR2 (N1782, N1769, N643);
not NOT1 (N1783, N1770);
nand NAND3 (N1784, N1775, N750, N1018);
or OR3 (N1785, N1783, N853, N1115);
nand NAND4 (N1786, N1782, N1599, N331, N1769);
not NOT1 (N1787, N1786);
or OR2 (N1788, N1768, N454);
or OR4 (N1789, N1787, N1071, N746, N82);
nand NAND4 (N1790, N1781, N1505, N1534, N958);
nor NOR2 (N1791, N1784, N1246);
nor NOR4 (N1792, N1780, N1743, N826, N1659);
nor NOR4 (N1793, N1788, N1223, N223, N185);
not NOT1 (N1794, N1774);
xor XOR2 (N1795, N1776, N1054);
xor XOR2 (N1796, N1785, N159);
buf BUF1 (N1797, N1795);
not NOT1 (N1798, N1789);
nand NAND2 (N1799, N1794, N676);
and AND3 (N1800, N1792, N233, N405);
buf BUF1 (N1801, N1793);
or OR2 (N1802, N1800, N258);
nand NAND3 (N1803, N1799, N484, N1300);
and AND4 (N1804, N1791, N1235, N1235, N766);
xor XOR2 (N1805, N1801, N631);
nand NAND3 (N1806, N1778, N930, N432);
buf BUF1 (N1807, N1797);
or OR3 (N1808, N1798, N1781, N1221);
nand NAND2 (N1809, N1805, N1602);
and AND2 (N1810, N1803, N63);
nor NOR4 (N1811, N1790, N695, N1498, N286);
and AND3 (N1812, N1810, N752, N1318);
buf BUF1 (N1813, N1804);
buf BUF1 (N1814, N1813);
buf BUF1 (N1815, N1808);
nor NOR4 (N1816, N1807, N985, N665, N1543);
buf BUF1 (N1817, N1814);
buf BUF1 (N1818, N1816);
nand NAND2 (N1819, N1802, N1788);
not NOT1 (N1820, N1811);
or OR4 (N1821, N1806, N72, N284, N1265);
not NOT1 (N1822, N1819);
nor NOR4 (N1823, N1820, N788, N812, N721);
and AND4 (N1824, N1772, N1552, N250, N793);
xor XOR2 (N1825, N1823, N1409);
not NOT1 (N1826, N1824);
and AND3 (N1827, N1825, N371, N1378);
not NOT1 (N1828, N1809);
or OR3 (N1829, N1821, N732, N1662);
nor NOR2 (N1830, N1796, N1627);
not NOT1 (N1831, N1828);
not NOT1 (N1832, N1829);
buf BUF1 (N1833, N1832);
nor NOR4 (N1834, N1833, N126, N669, N291);
nand NAND2 (N1835, N1826, N609);
nand NAND2 (N1836, N1818, N841);
or OR4 (N1837, N1815, N1720, N271, N534);
buf BUF1 (N1838, N1822);
nand NAND3 (N1839, N1827, N106, N130);
not NOT1 (N1840, N1835);
or OR3 (N1841, N1831, N887, N1105);
not NOT1 (N1842, N1834);
buf BUF1 (N1843, N1837);
nand NAND2 (N1844, N1830, N1406);
xor XOR2 (N1845, N1817, N1018);
nor NOR2 (N1846, N1843, N982);
nand NAND4 (N1847, N1842, N1341, N1786, N658);
not NOT1 (N1848, N1846);
buf BUF1 (N1849, N1838);
and AND3 (N1850, N1848, N1646, N602);
and AND2 (N1851, N1845, N1016);
nor NOR4 (N1852, N1839, N16, N1851, N1004);
xor XOR2 (N1853, N1593, N1290);
not NOT1 (N1854, N1812);
or OR4 (N1855, N1854, N279, N899, N287);
and AND3 (N1856, N1853, N1592, N1281);
buf BUF1 (N1857, N1841);
nand NAND2 (N1858, N1849, N1003);
xor XOR2 (N1859, N1836, N210);
not NOT1 (N1860, N1840);
nand NAND4 (N1861, N1852, N517, N1757, N35);
xor XOR2 (N1862, N1844, N827);
nand NAND2 (N1863, N1847, N1430);
buf BUF1 (N1864, N1855);
nand NAND4 (N1865, N1860, N458, N1818, N1559);
and AND2 (N1866, N1858, N445);
buf BUF1 (N1867, N1861);
nand NAND4 (N1868, N1856, N1785, N432, N134);
or OR3 (N1869, N1868, N1441, N1300);
nand NAND4 (N1870, N1859, N651, N219, N500);
nand NAND4 (N1871, N1865, N1099, N1836, N407);
buf BUF1 (N1872, N1870);
not NOT1 (N1873, N1871);
not NOT1 (N1874, N1872);
not NOT1 (N1875, N1850);
xor XOR2 (N1876, N1869, N899);
xor XOR2 (N1877, N1863, N668);
nand NAND2 (N1878, N1876, N222);
buf BUF1 (N1879, N1857);
nand NAND2 (N1880, N1867, N930);
nor NOR4 (N1881, N1879, N674, N149, N1026);
nor NOR4 (N1882, N1864, N171, N1564, N686);
and AND4 (N1883, N1877, N1233, N1254, N805);
nor NOR4 (N1884, N1880, N618, N1565, N1362);
nor NOR2 (N1885, N1882, N914);
and AND4 (N1886, N1885, N79, N125, N928);
not NOT1 (N1887, N1874);
xor XOR2 (N1888, N1881, N1274);
nor NOR3 (N1889, N1862, N1813, N1212);
buf BUF1 (N1890, N1883);
xor XOR2 (N1891, N1884, N1868);
buf BUF1 (N1892, N1887);
xor XOR2 (N1893, N1888, N610);
and AND4 (N1894, N1889, N748, N124, N948);
buf BUF1 (N1895, N1894);
or OR4 (N1896, N1893, N733, N1116, N404);
or OR2 (N1897, N1878, N1048);
or OR4 (N1898, N1896, N1794, N603, N47);
nand NAND4 (N1899, N1886, N1595, N1186, N420);
or OR2 (N1900, N1866, N640);
nor NOR2 (N1901, N1897, N1570);
xor XOR2 (N1902, N1890, N1367);
xor XOR2 (N1903, N1875, N263);
or OR3 (N1904, N1873, N757, N853);
or OR2 (N1905, N1892, N1497);
xor XOR2 (N1906, N1905, N594);
nor NOR3 (N1907, N1899, N853, N1124);
buf BUF1 (N1908, N1895);
nand NAND3 (N1909, N1908, N86, N1373);
not NOT1 (N1910, N1906);
xor XOR2 (N1911, N1909, N1553);
and AND3 (N1912, N1900, N1091, N25);
buf BUF1 (N1913, N1907);
buf BUF1 (N1914, N1891);
not NOT1 (N1915, N1911);
nor NOR3 (N1916, N1915, N1779, N1339);
xor XOR2 (N1917, N1914, N84);
and AND4 (N1918, N1910, N1804, N1446, N50);
nor NOR2 (N1919, N1898, N1069);
not NOT1 (N1920, N1904);
buf BUF1 (N1921, N1913);
buf BUF1 (N1922, N1916);
nor NOR3 (N1923, N1912, N345, N1449);
buf BUF1 (N1924, N1917);
or OR4 (N1925, N1924, N1468, N1500, N23);
nor NOR2 (N1926, N1921, N693);
and AND3 (N1927, N1920, N1792, N486);
nand NAND3 (N1928, N1927, N879, N360);
and AND4 (N1929, N1901, N1605, N491, N760);
buf BUF1 (N1930, N1922);
and AND3 (N1931, N1926, N394, N1665);
and AND3 (N1932, N1929, N698, N901);
or OR3 (N1933, N1918, N1731, N1507);
nor NOR4 (N1934, N1903, N1600, N1586, N301);
or OR2 (N1935, N1902, N1262);
nor NOR3 (N1936, N1935, N361, N595);
and AND2 (N1937, N1923, N1817);
buf BUF1 (N1938, N1932);
nor NOR4 (N1939, N1938, N533, N1419, N702);
xor XOR2 (N1940, N1931, N1201);
xor XOR2 (N1941, N1936, N546);
not NOT1 (N1942, N1928);
or OR3 (N1943, N1934, N387, N988);
xor XOR2 (N1944, N1930, N1565);
nor NOR2 (N1945, N1919, N1221);
not NOT1 (N1946, N1933);
xor XOR2 (N1947, N1945, N410);
nand NAND3 (N1948, N1946, N1373, N635);
buf BUF1 (N1949, N1948);
nor NOR2 (N1950, N1937, N1337);
or OR2 (N1951, N1943, N1807);
nand NAND2 (N1952, N1925, N1675);
buf BUF1 (N1953, N1940);
nand NAND3 (N1954, N1941, N930, N1368);
and AND3 (N1955, N1949, N218, N912);
or OR3 (N1956, N1947, N941, N966);
nand NAND3 (N1957, N1939, N675, N292);
nand NAND4 (N1958, N1956, N1542, N1777, N1011);
not NOT1 (N1959, N1942);
nor NOR3 (N1960, N1958, N1518, N1934);
or OR4 (N1961, N1957, N1260, N449, N1352);
or OR2 (N1962, N1944, N1034);
not NOT1 (N1963, N1955);
xor XOR2 (N1964, N1953, N891);
buf BUF1 (N1965, N1959);
xor XOR2 (N1966, N1963, N1720);
buf BUF1 (N1967, N1961);
nor NOR4 (N1968, N1965, N751, N64, N1877);
xor XOR2 (N1969, N1967, N1735);
or OR3 (N1970, N1954, N1937, N1775);
nor NOR2 (N1971, N1966, N1768);
not NOT1 (N1972, N1951);
or OR4 (N1973, N1972, N67, N745, N1164);
nor NOR3 (N1974, N1973, N183, N1691);
nor NOR4 (N1975, N1952, N805, N1345, N24);
and AND4 (N1976, N1960, N798, N679, N1013);
not NOT1 (N1977, N1975);
xor XOR2 (N1978, N1968, N1671);
xor XOR2 (N1979, N1971, N1948);
xor XOR2 (N1980, N1979, N732);
buf BUF1 (N1981, N1950);
nand NAND3 (N1982, N1974, N39, N315);
or OR3 (N1983, N1981, N1471, N1252);
nor NOR2 (N1984, N1976, N160);
or OR2 (N1985, N1982, N1445);
nor NOR3 (N1986, N1970, N1761, N1361);
xor XOR2 (N1987, N1969, N787);
or OR3 (N1988, N1978, N938, N1961);
and AND2 (N1989, N1977, N254);
xor XOR2 (N1990, N1985, N294);
or OR2 (N1991, N1988, N564);
and AND2 (N1992, N1986, N1798);
and AND2 (N1993, N1984, N275);
and AND4 (N1994, N1983, N1342, N1835, N396);
buf BUF1 (N1995, N1993);
nor NOR2 (N1996, N1995, N382);
nand NAND3 (N1997, N1987, N1627, N309);
nor NOR3 (N1998, N1991, N567, N223);
or OR2 (N1999, N1998, N1025);
nor NOR4 (N2000, N1996, N657, N1375, N179);
buf BUF1 (N2001, N1999);
buf BUF1 (N2002, N1994);
not NOT1 (N2003, N1962);
and AND4 (N2004, N1980, N621, N1185, N277);
nor NOR4 (N2005, N2000, N142, N1200, N1005);
buf BUF1 (N2006, N2001);
xor XOR2 (N2007, N1997, N1532);
and AND3 (N2008, N2002, N1825, N1936);
nand NAND3 (N2009, N1992, N128, N1835);
or OR3 (N2010, N2003, N1072, N1425);
buf BUF1 (N2011, N1989);
nand NAND3 (N2012, N2011, N1987, N1139);
buf BUF1 (N2013, N2005);
or OR2 (N2014, N1990, N991);
or OR2 (N2015, N1964, N532);
and AND3 (N2016, N2009, N1132, N1956);
nor NOR2 (N2017, N2010, N114);
not NOT1 (N2018, N2015);
not NOT1 (N2019, N2014);
not NOT1 (N2020, N2013);
and AND2 (N2021, N2008, N903);
not NOT1 (N2022, N2016);
buf BUF1 (N2023, N2007);
nor NOR4 (N2024, N2022, N1946, N1903, N696);
xor XOR2 (N2025, N2012, N1155);
nand NAND3 (N2026, N2006, N1454, N1103);
nand NAND2 (N2027, N2021, N1005);
xor XOR2 (N2028, N2020, N1851);
not NOT1 (N2029, N2027);
xor XOR2 (N2030, N2017, N858);
xor XOR2 (N2031, N2004, N416);
and AND4 (N2032, N2029, N826, N240, N861);
or OR4 (N2033, N2025, N567, N1219, N1997);
nand NAND4 (N2034, N2024, N980, N331, N1359);
and AND3 (N2035, N2023, N1661, N1765);
and AND2 (N2036, N2019, N1494);
and AND4 (N2037, N2033, N1887, N1850, N563);
xor XOR2 (N2038, N2028, N414);
and AND3 (N2039, N2035, N780, N1828);
and AND4 (N2040, N2038, N1687, N1078, N1161);
nor NOR2 (N2041, N2036, N1884);
not NOT1 (N2042, N2040);
or OR2 (N2043, N2034, N1360);
nor NOR2 (N2044, N2030, N1632);
not NOT1 (N2045, N2041);
not NOT1 (N2046, N2032);
nand NAND3 (N2047, N2039, N342, N319);
nor NOR3 (N2048, N2026, N17, N376);
not NOT1 (N2049, N2043);
xor XOR2 (N2050, N2047, N1245);
nor NOR3 (N2051, N2048, N379, N109);
buf BUF1 (N2052, N2046);
nor NOR2 (N2053, N2051, N516);
buf BUF1 (N2054, N2049);
or OR2 (N2055, N2050, N1840);
or OR4 (N2056, N2018, N494, N948, N1703);
nand NAND2 (N2057, N2042, N1519);
buf BUF1 (N2058, N2055);
nor NOR2 (N2059, N2052, N911);
nor NOR2 (N2060, N2054, N674);
or OR4 (N2061, N2037, N1127, N1069, N1042);
or OR4 (N2062, N2059, N1262, N992, N1393);
or OR3 (N2063, N2058, N578, N280);
not NOT1 (N2064, N2053);
nand NAND3 (N2065, N2045, N1943, N101);
nor NOR4 (N2066, N2060, N1746, N1913, N1618);
nand NAND2 (N2067, N2061, N1838);
not NOT1 (N2068, N2066);
not NOT1 (N2069, N2068);
not NOT1 (N2070, N2057);
and AND2 (N2071, N2067, N1517);
nor NOR4 (N2072, N2056, N402, N915, N203);
buf BUF1 (N2073, N2070);
or OR3 (N2074, N2031, N1673, N1474);
not NOT1 (N2075, N2073);
xor XOR2 (N2076, N2069, N910);
not NOT1 (N2077, N2063);
xor XOR2 (N2078, N2071, N1046);
nand NAND4 (N2079, N2064, N1143, N1498, N1774);
buf BUF1 (N2080, N2074);
buf BUF1 (N2081, N2078);
xor XOR2 (N2082, N2077, N995);
nand NAND4 (N2083, N2062, N266, N1490, N644);
xor XOR2 (N2084, N2072, N1472);
nand NAND2 (N2085, N2075, N1696);
nor NOR2 (N2086, N2083, N1647);
not NOT1 (N2087, N2079);
xor XOR2 (N2088, N2065, N772);
not NOT1 (N2089, N2044);
nand NAND3 (N2090, N2076, N86, N1073);
nand NAND2 (N2091, N2089, N1421);
or OR4 (N2092, N2082, N472, N308, N2055);
not NOT1 (N2093, N2086);
and AND3 (N2094, N2088, N433, N253);
buf BUF1 (N2095, N2084);
nand NAND3 (N2096, N2091, N1300, N2028);
nand NAND2 (N2097, N2081, N1444);
buf BUF1 (N2098, N2095);
nand NAND3 (N2099, N2090, N1982, N727);
nand NAND4 (N2100, N2097, N1134, N874, N1695);
nand NAND4 (N2101, N2100, N494, N882, N914);
or OR4 (N2102, N2096, N500, N1473, N112);
not NOT1 (N2103, N2092);
or OR3 (N2104, N2087, N2060, N1961);
not NOT1 (N2105, N2103);
buf BUF1 (N2106, N2093);
nand NAND4 (N2107, N2094, N1455, N1526, N1598);
buf BUF1 (N2108, N2099);
xor XOR2 (N2109, N2085, N1338);
xor XOR2 (N2110, N2106, N1387);
nand NAND4 (N2111, N2102, N954, N1108, N806);
nand NAND3 (N2112, N2104, N275, N1806);
and AND4 (N2113, N2107, N581, N1789, N705);
nand NAND3 (N2114, N2105, N342, N391);
not NOT1 (N2115, N2080);
buf BUF1 (N2116, N2115);
not NOT1 (N2117, N2112);
nand NAND3 (N2118, N2113, N2076, N1336);
and AND2 (N2119, N2109, N1588);
and AND3 (N2120, N2116, N1432, N1275);
nand NAND4 (N2121, N2114, N734, N1870, N1102);
not NOT1 (N2122, N2120);
buf BUF1 (N2123, N2119);
xor XOR2 (N2124, N2101, N995);
buf BUF1 (N2125, N2118);
xor XOR2 (N2126, N2111, N350);
xor XOR2 (N2127, N2123, N1823);
nand NAND2 (N2128, N2110, N2016);
nand NAND2 (N2129, N2108, N1007);
nor NOR3 (N2130, N2121, N769, N1902);
xor XOR2 (N2131, N2122, N250);
not NOT1 (N2132, N2126);
and AND2 (N2133, N2125, N1154);
or OR4 (N2134, N2127, N78, N1006, N1364);
nand NAND2 (N2135, N2098, N306);
or OR2 (N2136, N2128, N1596);
xor XOR2 (N2137, N2117, N188);
nand NAND3 (N2138, N2136, N1453, N447);
xor XOR2 (N2139, N2138, N433);
xor XOR2 (N2140, N2124, N1424);
xor XOR2 (N2141, N2135, N2097);
nor NOR4 (N2142, N2141, N1740, N1127, N1450);
xor XOR2 (N2143, N2142, N1018);
nor NOR4 (N2144, N2130, N1623, N1958, N1613);
not NOT1 (N2145, N2137);
not NOT1 (N2146, N2131);
nor NOR3 (N2147, N2145, N1916, N681);
nand NAND2 (N2148, N2146, N1642);
and AND4 (N2149, N2143, N466, N851, N156);
nand NAND4 (N2150, N2129, N323, N276, N257);
nor NOR4 (N2151, N2150, N1821, N1642, N87);
buf BUF1 (N2152, N2151);
xor XOR2 (N2153, N2140, N614);
buf BUF1 (N2154, N2133);
or OR3 (N2155, N2132, N155, N1977);
buf BUF1 (N2156, N2152);
xor XOR2 (N2157, N2155, N23);
or OR4 (N2158, N2144, N546, N733, N1123);
xor XOR2 (N2159, N2156, N220);
not NOT1 (N2160, N2159);
xor XOR2 (N2161, N2149, N58);
xor XOR2 (N2162, N2147, N384);
or OR4 (N2163, N2148, N1813, N690, N1518);
and AND3 (N2164, N2160, N511, N372);
xor XOR2 (N2165, N2157, N1349);
buf BUF1 (N2166, N2158);
nand NAND2 (N2167, N2165, N825);
not NOT1 (N2168, N2139);
or OR3 (N2169, N2168, N2161, N654);
buf BUF1 (N2170, N982);
and AND2 (N2171, N2170, N1527);
xor XOR2 (N2172, N2154, N1387);
nand NAND4 (N2173, N2164, N1503, N1316, N1872);
or OR2 (N2174, N2172, N2104);
or OR2 (N2175, N2173, N1226);
buf BUF1 (N2176, N2169);
nand NAND4 (N2177, N2153, N2147, N208, N813);
xor XOR2 (N2178, N2166, N1144);
xor XOR2 (N2179, N2174, N2028);
nor NOR3 (N2180, N2178, N1824, N1840);
not NOT1 (N2181, N2176);
not NOT1 (N2182, N2181);
xor XOR2 (N2183, N2175, N2173);
nand NAND4 (N2184, N2182, N876, N966, N1179);
nor NOR3 (N2185, N2179, N1981, N634);
and AND3 (N2186, N2185, N1484, N1690);
xor XOR2 (N2187, N2183, N915);
xor XOR2 (N2188, N2186, N942);
xor XOR2 (N2189, N2187, N790);
nor NOR2 (N2190, N2188, N121);
xor XOR2 (N2191, N2134, N429);
or OR2 (N2192, N2167, N206);
not NOT1 (N2193, N2171);
buf BUF1 (N2194, N2162);
nor NOR4 (N2195, N2193, N817, N95, N146);
or OR3 (N2196, N2177, N1397, N1586);
buf BUF1 (N2197, N2196);
and AND3 (N2198, N2184, N1220, N1521);
and AND3 (N2199, N2192, N1318, N1023);
and AND2 (N2200, N2180, N999);
nor NOR3 (N2201, N2163, N2098, N1217);
or OR2 (N2202, N2190, N1469);
nor NOR2 (N2203, N2198, N877);
nand NAND3 (N2204, N2199, N203, N354);
xor XOR2 (N2205, N2204, N72);
and AND4 (N2206, N2189, N1485, N1508, N1166);
xor XOR2 (N2207, N2206, N307);
and AND3 (N2208, N2195, N581, N1651);
not NOT1 (N2209, N2205);
or OR4 (N2210, N2201, N1248, N1437, N578);
xor XOR2 (N2211, N2200, N1994);
buf BUF1 (N2212, N2211);
nor NOR2 (N2213, N2197, N948);
or OR2 (N2214, N2212, N1100);
and AND4 (N2215, N2207, N488, N1731, N1253);
buf BUF1 (N2216, N2194);
not NOT1 (N2217, N2210);
nor NOR4 (N2218, N2213, N937, N692, N2133);
xor XOR2 (N2219, N2209, N267);
nand NAND4 (N2220, N2203, N1161, N330, N1625);
xor XOR2 (N2221, N2217, N1544);
nor NOR2 (N2222, N2216, N1378);
nor NOR4 (N2223, N2208, N1666, N1366, N1090);
buf BUF1 (N2224, N2220);
buf BUF1 (N2225, N2218);
and AND2 (N2226, N2224, N908);
not NOT1 (N2227, N2226);
or OR3 (N2228, N2222, N499, N1229);
xor XOR2 (N2229, N2225, N176);
not NOT1 (N2230, N2214);
xor XOR2 (N2231, N2227, N2165);
nor NOR2 (N2232, N2223, N1379);
nor NOR2 (N2233, N2228, N1987);
nand NAND4 (N2234, N2215, N1886, N818, N334);
buf BUF1 (N2235, N2191);
buf BUF1 (N2236, N2231);
and AND3 (N2237, N2221, N1164, N2173);
nand NAND3 (N2238, N2219, N2140, N1394);
xor XOR2 (N2239, N2238, N552);
not NOT1 (N2240, N2237);
nand NAND3 (N2241, N2236, N1433, N598);
not NOT1 (N2242, N2235);
nor NOR4 (N2243, N2229, N319, N820, N898);
xor XOR2 (N2244, N2242, N1692);
buf BUF1 (N2245, N2239);
nand NAND2 (N2246, N2244, N1377);
or OR3 (N2247, N2245, N1672, N527);
not NOT1 (N2248, N2240);
or OR4 (N2249, N2234, N1034, N1548, N1996);
or OR2 (N2250, N2247, N139);
or OR2 (N2251, N2246, N1091);
nand NAND2 (N2252, N2248, N584);
or OR4 (N2253, N2202, N1818, N2207, N732);
not NOT1 (N2254, N2233);
nor NOR4 (N2255, N2254, N1474, N2109, N152);
and AND3 (N2256, N2253, N2054, N334);
nor NOR3 (N2257, N2232, N2009, N546);
nor NOR2 (N2258, N2230, N1293);
nand NAND2 (N2259, N2241, N2001);
nor NOR4 (N2260, N2251, N1332, N1517, N1111);
nand NAND4 (N2261, N2257, N2235, N1039, N1090);
nand NAND3 (N2262, N2252, N319, N191);
not NOT1 (N2263, N2255);
not NOT1 (N2264, N2243);
and AND4 (N2265, N2258, N1617, N1891, N707);
xor XOR2 (N2266, N2261, N1245);
or OR4 (N2267, N2256, N197, N1896, N440);
buf BUF1 (N2268, N2265);
nor NOR2 (N2269, N2250, N1317);
xor XOR2 (N2270, N2269, N2051);
xor XOR2 (N2271, N2268, N1401);
buf BUF1 (N2272, N2270);
or OR3 (N2273, N2259, N329, N1003);
or OR4 (N2274, N2272, N925, N475, N261);
nor NOR3 (N2275, N2263, N1095, N1736);
buf BUF1 (N2276, N2249);
and AND4 (N2277, N2262, N649, N1090, N1179);
nor NOR4 (N2278, N2260, N943, N591, N2083);
and AND4 (N2279, N2273, N983, N2161, N1735);
buf BUF1 (N2280, N2271);
and AND2 (N2281, N2274, N539);
nand NAND3 (N2282, N2277, N1465, N837);
buf BUF1 (N2283, N2280);
or OR4 (N2284, N2282, N748, N498, N1184);
buf BUF1 (N2285, N2284);
nand NAND2 (N2286, N2275, N2221);
not NOT1 (N2287, N2281);
xor XOR2 (N2288, N2286, N2015);
nor NOR4 (N2289, N2279, N461, N267, N43);
not NOT1 (N2290, N2289);
buf BUF1 (N2291, N2288);
and AND2 (N2292, N2285, N1421);
nand NAND2 (N2293, N2276, N592);
nand NAND4 (N2294, N2292, N1230, N2150, N1311);
not NOT1 (N2295, N2264);
nor NOR2 (N2296, N2266, N2220);
nand NAND4 (N2297, N2278, N1602, N1519, N409);
or OR4 (N2298, N2290, N1608, N1086, N1664);
or OR4 (N2299, N2294, N1454, N440, N1633);
nand NAND3 (N2300, N2291, N2228, N1356);
buf BUF1 (N2301, N2287);
or OR2 (N2302, N2298, N506);
and AND2 (N2303, N2302, N1338);
and AND2 (N2304, N2295, N2029);
nor NOR3 (N2305, N2296, N11, N1576);
nor NOR3 (N2306, N2305, N310, N1826);
or OR2 (N2307, N2301, N2259);
or OR2 (N2308, N2267, N647);
buf BUF1 (N2309, N2304);
or OR3 (N2310, N2300, N1610, N373);
buf BUF1 (N2311, N2293);
or OR3 (N2312, N2310, N1018, N2115);
xor XOR2 (N2313, N2309, N2215);
xor XOR2 (N2314, N2303, N2265);
not NOT1 (N2315, N2311);
or OR4 (N2316, N2299, N958, N823, N1416);
or OR3 (N2317, N2312, N2297, N1856);
not NOT1 (N2318, N1136);
and AND2 (N2319, N2308, N1483);
xor XOR2 (N2320, N2307, N228);
not NOT1 (N2321, N2306);
nand NAND4 (N2322, N2317, N332, N1042, N1402);
nor NOR2 (N2323, N2283, N2278);
not NOT1 (N2324, N2315);
nor NOR3 (N2325, N2313, N381, N1542);
and AND3 (N2326, N2325, N183, N1290);
nor NOR3 (N2327, N2320, N70, N25);
nor NOR3 (N2328, N2323, N217, N2095);
buf BUF1 (N2329, N2328);
nor NOR3 (N2330, N2327, N415, N1957);
nor NOR2 (N2331, N2318, N396);
or OR2 (N2332, N2324, N1826);
not NOT1 (N2333, N2332);
xor XOR2 (N2334, N2321, N2158);
xor XOR2 (N2335, N2316, N237);
and AND3 (N2336, N2330, N1392, N1964);
buf BUF1 (N2337, N2333);
not NOT1 (N2338, N2319);
nor NOR3 (N2339, N2334, N1835, N809);
buf BUF1 (N2340, N2331);
and AND2 (N2341, N2340, N830);
nor NOR3 (N2342, N2339, N1036, N495);
nand NAND3 (N2343, N2314, N410, N1448);
nor NOR2 (N2344, N2337, N5);
not NOT1 (N2345, N2343);
xor XOR2 (N2346, N2345, N2036);
nand NAND3 (N2347, N2335, N2323, N907);
nor NOR3 (N2348, N2344, N1259, N1913);
nand NAND4 (N2349, N2342, N1894, N1223, N1287);
xor XOR2 (N2350, N2346, N455);
nor NOR3 (N2351, N2349, N723, N1243);
or OR2 (N2352, N2350, N632);
nor NOR2 (N2353, N2329, N1746);
and AND4 (N2354, N2326, N1601, N1080, N1363);
and AND4 (N2355, N2352, N1424, N79, N141);
and AND2 (N2356, N2336, N1358);
not NOT1 (N2357, N2354);
nand NAND4 (N2358, N2357, N209, N237, N408);
not NOT1 (N2359, N2353);
or OR4 (N2360, N2358, N2156, N2020, N903);
nand NAND4 (N2361, N2347, N435, N1794, N2215);
nor NOR4 (N2362, N2361, N241, N1755, N1885);
xor XOR2 (N2363, N2341, N1522);
nand NAND2 (N2364, N2351, N32);
not NOT1 (N2365, N2363);
buf BUF1 (N2366, N2362);
nand NAND3 (N2367, N2338, N1566, N896);
xor XOR2 (N2368, N2348, N1664);
not NOT1 (N2369, N2366);
or OR3 (N2370, N2369, N1634, N2047);
nand NAND2 (N2371, N2360, N143);
xor XOR2 (N2372, N2367, N684);
xor XOR2 (N2373, N2364, N368);
and AND2 (N2374, N2373, N1222);
or OR4 (N2375, N2372, N995, N1996, N448);
nand NAND2 (N2376, N2322, N346);
xor XOR2 (N2377, N2374, N930);
buf BUF1 (N2378, N2370);
buf BUF1 (N2379, N2371);
not NOT1 (N2380, N2359);
nand NAND4 (N2381, N2379, N2021, N1704, N1150);
or OR4 (N2382, N2375, N209, N1254, N690);
buf BUF1 (N2383, N2365);
buf BUF1 (N2384, N2383);
nor NOR4 (N2385, N2378, N1024, N202, N618);
not NOT1 (N2386, N2377);
and AND3 (N2387, N2380, N1187, N880);
and AND4 (N2388, N2356, N1067, N2347, N1325);
not NOT1 (N2389, N2382);
nor NOR3 (N2390, N2368, N1210, N2080);
nor NOR3 (N2391, N2381, N2249, N2136);
buf BUF1 (N2392, N2355);
nand NAND3 (N2393, N2384, N1113, N2151);
nand NAND2 (N2394, N2388, N1120);
buf BUF1 (N2395, N2387);
nand NAND4 (N2396, N2389, N902, N2077, N275);
nand NAND4 (N2397, N2393, N2111, N1886, N139);
xor XOR2 (N2398, N2376, N1596);
and AND3 (N2399, N2397, N1438, N479);
buf BUF1 (N2400, N2395);
not NOT1 (N2401, N2400);
nand NAND4 (N2402, N2386, N704, N991, N1521);
nand NAND4 (N2403, N2394, N2262, N2023, N2099);
or OR3 (N2404, N2391, N5, N1537);
or OR4 (N2405, N2399, N1728, N1351, N1230);
or OR3 (N2406, N2402, N1884, N1931);
and AND2 (N2407, N2405, N122);
or OR3 (N2408, N2398, N894, N1307);
nand NAND3 (N2409, N2396, N926, N1407);
nor NOR2 (N2410, N2406, N1699);
or OR4 (N2411, N2408, N563, N349, N549);
xor XOR2 (N2412, N2390, N1732);
and AND3 (N2413, N2410, N2087, N859);
nor NOR3 (N2414, N2413, N5, N79);
not NOT1 (N2415, N2403);
nor NOR2 (N2416, N2414, N693);
xor XOR2 (N2417, N2401, N1226);
or OR4 (N2418, N2404, N455, N1666, N1593);
nor NOR2 (N2419, N2407, N699);
and AND3 (N2420, N2417, N168, N1670);
not NOT1 (N2421, N2415);
nor NOR3 (N2422, N2416, N1739, N117);
xor XOR2 (N2423, N2392, N57);
and AND2 (N2424, N2418, N1633);
nand NAND2 (N2425, N2424, N1348);
buf BUF1 (N2426, N2421);
not NOT1 (N2427, N2419);
or OR4 (N2428, N2412, N2338, N815, N121);
nand NAND4 (N2429, N2428, N1671, N1324, N1610);
and AND2 (N2430, N2426, N482);
not NOT1 (N2431, N2411);
buf BUF1 (N2432, N2423);
nand NAND4 (N2433, N2432, N254, N574, N1099);
or OR3 (N2434, N2433, N702, N792);
nand NAND4 (N2435, N2427, N1497, N4, N2066);
and AND3 (N2436, N2431, N877, N1189);
buf BUF1 (N2437, N2425);
and AND2 (N2438, N2429, N1111);
nand NAND3 (N2439, N2434, N666, N1527);
and AND3 (N2440, N2385, N2023, N1217);
not NOT1 (N2441, N2435);
xor XOR2 (N2442, N2439, N395);
and AND4 (N2443, N2409, N522, N181, N341);
buf BUF1 (N2444, N2440);
nor NOR3 (N2445, N2437, N2046, N96);
and AND3 (N2446, N2442, N873, N2332);
buf BUF1 (N2447, N2443);
buf BUF1 (N2448, N2446);
nor NOR2 (N2449, N2422, N1234);
and AND4 (N2450, N2449, N2143, N503, N902);
not NOT1 (N2451, N2448);
nor NOR3 (N2452, N2430, N1468, N1781);
or OR3 (N2453, N2436, N1401, N1376);
nand NAND3 (N2454, N2452, N577, N268);
and AND4 (N2455, N2441, N1165, N399, N2161);
not NOT1 (N2456, N2444);
not NOT1 (N2457, N2453);
or OR4 (N2458, N2447, N971, N1650, N1858);
nor NOR2 (N2459, N2455, N812);
nor NOR2 (N2460, N2450, N726);
and AND4 (N2461, N2438, N668, N1450, N2139);
or OR2 (N2462, N2420, N2437);
nand NAND3 (N2463, N2458, N1492, N31);
nand NAND2 (N2464, N2461, N732);
nand NAND4 (N2465, N2459, N1846, N2168, N165);
or OR2 (N2466, N2463, N1637);
not NOT1 (N2467, N2445);
and AND4 (N2468, N2454, N1884, N672, N1045);
nor NOR3 (N2469, N2451, N1621, N861);
or OR4 (N2470, N2457, N484, N1935, N476);
or OR2 (N2471, N2470, N1324);
not NOT1 (N2472, N2460);
not NOT1 (N2473, N2466);
or OR3 (N2474, N2462, N1813, N1089);
and AND2 (N2475, N2469, N2001);
xor XOR2 (N2476, N2473, N2259);
nor NOR4 (N2477, N2465, N1181, N1930, N41);
xor XOR2 (N2478, N2467, N962);
and AND4 (N2479, N2456, N383, N1265, N1213);
not NOT1 (N2480, N2474);
or OR3 (N2481, N2471, N1011, N2378);
not NOT1 (N2482, N2479);
buf BUF1 (N2483, N2478);
and AND4 (N2484, N2476, N1462, N100, N393);
or OR2 (N2485, N2477, N359);
nor NOR4 (N2486, N2481, N1691, N271, N2000);
nand NAND2 (N2487, N2480, N2256);
or OR3 (N2488, N2486, N2479, N1812);
not NOT1 (N2489, N2484);
or OR4 (N2490, N2472, N2029, N2075, N523);
xor XOR2 (N2491, N2483, N104);
buf BUF1 (N2492, N2482);
nand NAND3 (N2493, N2489, N4, N2371);
nand NAND2 (N2494, N2488, N414);
not NOT1 (N2495, N2475);
or OR3 (N2496, N2492, N1518, N1334);
xor XOR2 (N2497, N2496, N1530);
not NOT1 (N2498, N2490);
or OR3 (N2499, N2485, N1506, N832);
buf BUF1 (N2500, N2491);
or OR3 (N2501, N2494, N1564, N225);
nand NAND3 (N2502, N2501, N845, N264);
xor XOR2 (N2503, N2493, N99);
and AND3 (N2504, N2464, N1804, N2041);
and AND4 (N2505, N2498, N127, N2138, N1900);
or OR3 (N2506, N2502, N12, N312);
nand NAND3 (N2507, N2505, N2120, N1991);
and AND2 (N2508, N2500, N1980);
and AND4 (N2509, N2508, N700, N297, N2335);
or OR2 (N2510, N2509, N208);
or OR4 (N2511, N2487, N1745, N1090, N227);
xor XOR2 (N2512, N2506, N1705);
nand NAND2 (N2513, N2499, N847);
xor XOR2 (N2514, N2511, N820);
and AND3 (N2515, N2495, N2443, N821);
and AND2 (N2516, N2514, N486);
nor NOR4 (N2517, N2510, N884, N749, N2318);
nand NAND2 (N2518, N2516, N2284);
buf BUF1 (N2519, N2468);
and AND2 (N2520, N2504, N418);
and AND2 (N2521, N2503, N444);
nor NOR2 (N2522, N2507, N1228);
buf BUF1 (N2523, N2515);
or OR3 (N2524, N2518, N248, N2116);
not NOT1 (N2525, N2520);
or OR2 (N2526, N2512, N1440);
and AND2 (N2527, N2521, N822);
xor XOR2 (N2528, N2497, N291);
nor NOR4 (N2529, N2523, N817, N1546, N1700);
xor XOR2 (N2530, N2513, N214);
nor NOR3 (N2531, N2522, N1447, N702);
xor XOR2 (N2532, N2525, N1959);
not NOT1 (N2533, N2519);
nand NAND4 (N2534, N2530, N656, N649, N1431);
nand NAND4 (N2535, N2526, N2175, N1148, N271);
buf BUF1 (N2536, N2528);
nor NOR2 (N2537, N2524, N1093);
and AND2 (N2538, N2536, N2093);
or OR4 (N2539, N2537, N1515, N997, N850);
or OR3 (N2540, N2532, N1192, N979);
not NOT1 (N2541, N2534);
nand NAND3 (N2542, N2527, N1270, N1188);
and AND3 (N2543, N2535, N290, N1483);
nand NAND3 (N2544, N2541, N1971, N1947);
nand NAND2 (N2545, N2543, N2343);
not NOT1 (N2546, N2538);
buf BUF1 (N2547, N2517);
not NOT1 (N2548, N2545);
not NOT1 (N2549, N2544);
or OR4 (N2550, N2549, N633, N452, N526);
buf BUF1 (N2551, N2531);
xor XOR2 (N2552, N2533, N355);
or OR4 (N2553, N2552, N2470, N2503, N572);
not NOT1 (N2554, N2548);
or OR3 (N2555, N2550, N2241, N1710);
buf BUF1 (N2556, N2539);
buf BUF1 (N2557, N2542);
nand NAND3 (N2558, N2540, N581, N11);
buf BUF1 (N2559, N2553);
nor NOR2 (N2560, N2529, N394);
buf BUF1 (N2561, N2560);
nand NAND2 (N2562, N2551, N1195);
nor NOR3 (N2563, N2547, N450, N874);
xor XOR2 (N2564, N2562, N330);
xor XOR2 (N2565, N2558, N2469);
xor XOR2 (N2566, N2554, N1868);
or OR2 (N2567, N2557, N2351);
xor XOR2 (N2568, N2556, N2487);
xor XOR2 (N2569, N2565, N583);
or OR2 (N2570, N2563, N2366);
nor NOR2 (N2571, N2567, N1589);
nand NAND3 (N2572, N2569, N542, N329);
or OR3 (N2573, N2555, N2497, N181);
nand NAND4 (N2574, N2564, N154, N1978, N641);
and AND4 (N2575, N2573, N1758, N1421, N296);
xor XOR2 (N2576, N2574, N1677);
nor NOR2 (N2577, N2576, N1176);
buf BUF1 (N2578, N2572);
and AND2 (N2579, N2561, N51);
and AND2 (N2580, N2570, N1581);
nand NAND4 (N2581, N2571, N1724, N569, N568);
buf BUF1 (N2582, N2568);
nor NOR2 (N2583, N2577, N1632);
not NOT1 (N2584, N2566);
or OR3 (N2585, N2580, N2333, N335);
nand NAND4 (N2586, N2583, N358, N320, N919);
not NOT1 (N2587, N2575);
buf BUF1 (N2588, N2586);
nand NAND3 (N2589, N2582, N1673, N49);
or OR4 (N2590, N2559, N1123, N761, N122);
buf BUF1 (N2591, N2584);
or OR2 (N2592, N2591, N791);
and AND4 (N2593, N2587, N2481, N1209, N2099);
nor NOR4 (N2594, N2546, N1654, N303, N607);
xor XOR2 (N2595, N2594, N741);
buf BUF1 (N2596, N2588);
buf BUF1 (N2597, N2593);
xor XOR2 (N2598, N2585, N924);
nand NAND3 (N2599, N2590, N63, N2219);
xor XOR2 (N2600, N2581, N2358);
and AND2 (N2601, N2598, N628);
nand NAND4 (N2602, N2579, N1853, N1207, N606);
or OR4 (N2603, N2578, N1276, N766, N1690);
xor XOR2 (N2604, N2595, N307);
nor NOR3 (N2605, N2601, N1356, N2347);
or OR3 (N2606, N2605, N1558, N980);
buf BUF1 (N2607, N2596);
not NOT1 (N2608, N2607);
and AND2 (N2609, N2589, N924);
buf BUF1 (N2610, N2603);
buf BUF1 (N2611, N2610);
and AND2 (N2612, N2600, N2542);
not NOT1 (N2613, N2592);
nor NOR3 (N2614, N2604, N2473, N309);
buf BUF1 (N2615, N2597);
xor XOR2 (N2616, N2614, N1575);
nand NAND2 (N2617, N2602, N2282);
and AND4 (N2618, N2611, N492, N12, N26);
nand NAND3 (N2619, N2612, N223, N647);
buf BUF1 (N2620, N2616);
buf BUF1 (N2621, N2620);
not NOT1 (N2622, N2621);
not NOT1 (N2623, N2615);
nand NAND3 (N2624, N2606, N511, N2472);
nor NOR2 (N2625, N2623, N186);
xor XOR2 (N2626, N2599, N391);
and AND3 (N2627, N2608, N1510, N1539);
or OR4 (N2628, N2619, N1572, N2032, N1987);
and AND4 (N2629, N2624, N2611, N679, N1003);
nand NAND3 (N2630, N2628, N114, N2005);
and AND3 (N2631, N2613, N2073, N1442);
and AND3 (N2632, N2625, N2309, N1703);
xor XOR2 (N2633, N2627, N400);
and AND2 (N2634, N2630, N978);
and AND4 (N2635, N2634, N2252, N2188, N250);
xor XOR2 (N2636, N2622, N2380);
nand NAND4 (N2637, N2635, N2610, N1017, N2115);
and AND2 (N2638, N2626, N641);
nand NAND2 (N2639, N2637, N1045);
or OR3 (N2640, N2636, N1383, N113);
buf BUF1 (N2641, N2617);
buf BUF1 (N2642, N2618);
and AND4 (N2643, N2633, N878, N2362, N2627);
xor XOR2 (N2644, N2639, N1043);
not NOT1 (N2645, N2638);
or OR4 (N2646, N2645, N1514, N1665, N2095);
not NOT1 (N2647, N2609);
or OR4 (N2648, N2631, N1869, N1108, N2461);
and AND4 (N2649, N2629, N611, N1111, N1155);
nor NOR2 (N2650, N2640, N1543);
and AND2 (N2651, N2646, N1868);
buf BUF1 (N2652, N2632);
xor XOR2 (N2653, N2644, N308);
not NOT1 (N2654, N2647);
nor NOR2 (N2655, N2654, N698);
nor NOR3 (N2656, N2642, N954, N67);
not NOT1 (N2657, N2655);
or OR3 (N2658, N2653, N1289, N465);
buf BUF1 (N2659, N2652);
nor NOR3 (N2660, N2656, N1589, N2007);
and AND2 (N2661, N2643, N320);
or OR3 (N2662, N2641, N385, N1247);
or OR2 (N2663, N2658, N368);
buf BUF1 (N2664, N2650);
buf BUF1 (N2665, N2651);
not NOT1 (N2666, N2649);
and AND4 (N2667, N2665, N1872, N1627, N1599);
not NOT1 (N2668, N2657);
nand NAND4 (N2669, N2661, N941, N2284, N896);
or OR3 (N2670, N2669, N1840, N2431);
buf BUF1 (N2671, N2663);
xor XOR2 (N2672, N2671, N2414);
nand NAND2 (N2673, N2667, N1449);
nand NAND3 (N2674, N2672, N2125, N671);
or OR2 (N2675, N2660, N2098);
buf BUF1 (N2676, N2666);
nand NAND4 (N2677, N2675, N1918, N1193, N585);
not NOT1 (N2678, N2677);
and AND3 (N2679, N2674, N992, N2106);
or OR3 (N2680, N2676, N963, N895);
or OR4 (N2681, N2668, N590, N2167, N1941);
or OR2 (N2682, N2664, N410);
xor XOR2 (N2683, N2670, N16);
and AND3 (N2684, N2681, N1015, N1785);
xor XOR2 (N2685, N2682, N2143);
xor XOR2 (N2686, N2662, N246);
not NOT1 (N2687, N2648);
buf BUF1 (N2688, N2683);
buf BUF1 (N2689, N2673);
or OR4 (N2690, N2659, N1283, N455, N797);
buf BUF1 (N2691, N2678);
nor NOR3 (N2692, N2679, N909, N2150);
nor NOR3 (N2693, N2691, N1071, N228);
not NOT1 (N2694, N2690);
nor NOR4 (N2695, N2694, N366, N2047, N2558);
or OR3 (N2696, N2680, N2541, N2227);
and AND3 (N2697, N2692, N38, N830);
nand NAND3 (N2698, N2695, N1695, N1913);
or OR2 (N2699, N2693, N2121);
not NOT1 (N2700, N2698);
nand NAND2 (N2701, N2697, N889);
xor XOR2 (N2702, N2688, N1413);
and AND3 (N2703, N2687, N69, N867);
or OR4 (N2704, N2700, N621, N561, N1824);
buf BUF1 (N2705, N2696);
nor NOR4 (N2706, N2689, N790, N342, N373);
not NOT1 (N2707, N2701);
nand NAND3 (N2708, N2684, N568, N236);
buf BUF1 (N2709, N2707);
xor XOR2 (N2710, N2706, N2644);
nor NOR2 (N2711, N2709, N560);
or OR2 (N2712, N2710, N2395);
or OR4 (N2713, N2686, N533, N468, N2060);
and AND4 (N2714, N2703, N594, N1936, N1313);
nand NAND4 (N2715, N2704, N954, N1887, N2053);
not NOT1 (N2716, N2715);
nor NOR3 (N2717, N2711, N2126, N480);
nand NAND4 (N2718, N2705, N2625, N1282, N2266);
or OR4 (N2719, N2708, N1411, N724, N267);
xor XOR2 (N2720, N2713, N329);
and AND3 (N2721, N2712, N2710, N2188);
nor NOR3 (N2722, N2720, N939, N473);
nor NOR3 (N2723, N2719, N1849, N2472);
and AND2 (N2724, N2717, N520);
nand NAND4 (N2725, N2716, N1721, N1739, N855);
or OR4 (N2726, N2725, N2111, N1342, N1637);
not NOT1 (N2727, N2722);
and AND3 (N2728, N2714, N16, N505);
nor NOR2 (N2729, N2702, N1121);
and AND2 (N2730, N2726, N1885);
nand NAND3 (N2731, N2724, N2479, N1671);
nor NOR4 (N2732, N2731, N336, N723, N2438);
xor XOR2 (N2733, N2699, N2087);
or OR4 (N2734, N2732, N62, N130, N2258);
nand NAND2 (N2735, N2730, N2468);
xor XOR2 (N2736, N2735, N1786);
nand NAND3 (N2737, N2736, N2695, N356);
or OR4 (N2738, N2718, N2025, N517, N1589);
buf BUF1 (N2739, N2721);
and AND4 (N2740, N2729, N1896, N817, N2081);
nor NOR3 (N2741, N2723, N308, N239);
xor XOR2 (N2742, N2685, N1556);
nor NOR3 (N2743, N2733, N2272, N471);
not NOT1 (N2744, N2743);
nor NOR4 (N2745, N2739, N979, N2664, N475);
or OR2 (N2746, N2728, N1847);
not NOT1 (N2747, N2745);
not NOT1 (N2748, N2738);
nor NOR3 (N2749, N2741, N1847, N1894);
not NOT1 (N2750, N2740);
and AND4 (N2751, N2750, N2492, N1515, N63);
not NOT1 (N2752, N2744);
or OR4 (N2753, N2742, N1349, N2689, N1915);
xor XOR2 (N2754, N2746, N1479);
nand NAND3 (N2755, N2737, N1922, N2363);
nand NAND3 (N2756, N2734, N1221, N1237);
and AND4 (N2757, N2748, N564, N953, N529);
nor NOR3 (N2758, N2757, N740, N787);
not NOT1 (N2759, N2752);
xor XOR2 (N2760, N2754, N433);
not NOT1 (N2761, N2759);
buf BUF1 (N2762, N2751);
nand NAND4 (N2763, N2727, N1132, N890, N726);
buf BUF1 (N2764, N2760);
or OR3 (N2765, N2763, N2281, N1834);
not NOT1 (N2766, N2755);
buf BUF1 (N2767, N2747);
or OR2 (N2768, N2762, N2359);
nand NAND2 (N2769, N2758, N2453);
nand NAND4 (N2770, N2749, N2343, N487, N2592);
nand NAND3 (N2771, N2766, N2005, N2364);
xor XOR2 (N2772, N2753, N433);
not NOT1 (N2773, N2772);
nand NAND4 (N2774, N2768, N2613, N967, N2438);
nor NOR4 (N2775, N2761, N1518, N463, N682);
or OR3 (N2776, N2767, N1424, N1483);
xor XOR2 (N2777, N2756, N1676);
xor XOR2 (N2778, N2765, N2572);
xor XOR2 (N2779, N2776, N1114);
nor NOR3 (N2780, N2770, N1108, N36);
buf BUF1 (N2781, N2773);
buf BUF1 (N2782, N2764);
not NOT1 (N2783, N2777);
not NOT1 (N2784, N2783);
buf BUF1 (N2785, N2769);
xor XOR2 (N2786, N2781, N2220);
nor NOR3 (N2787, N2779, N1057, N75);
buf BUF1 (N2788, N2782);
buf BUF1 (N2789, N2788);
or OR3 (N2790, N2789, N964, N1328);
or OR2 (N2791, N2787, N199);
not NOT1 (N2792, N2774);
or OR3 (N2793, N2771, N985, N1926);
buf BUF1 (N2794, N2780);
not NOT1 (N2795, N2775);
nor NOR4 (N2796, N2793, N645, N537, N2308);
xor XOR2 (N2797, N2794, N1796);
or OR3 (N2798, N2778, N2253, N610);
nand NAND2 (N2799, N2784, N2532);
buf BUF1 (N2800, N2796);
buf BUF1 (N2801, N2785);
xor XOR2 (N2802, N2798, N580);
or OR4 (N2803, N2802, N2428, N1496, N273);
buf BUF1 (N2804, N2786);
nor NOR3 (N2805, N2799, N1933, N1226);
buf BUF1 (N2806, N2803);
nor NOR4 (N2807, N2800, N993, N327, N164);
buf BUF1 (N2808, N2806);
xor XOR2 (N2809, N2797, N1069);
xor XOR2 (N2810, N2804, N754);
or OR4 (N2811, N2790, N2219, N1500, N1667);
and AND2 (N2812, N2805, N1415);
buf BUF1 (N2813, N2812);
xor XOR2 (N2814, N2807, N2382);
buf BUF1 (N2815, N2801);
buf BUF1 (N2816, N2811);
and AND2 (N2817, N2814, N1895);
and AND3 (N2818, N2808, N2622, N890);
or OR4 (N2819, N2809, N1364, N2222, N1923);
and AND2 (N2820, N2795, N1474);
not NOT1 (N2821, N2819);
or OR3 (N2822, N2821, N2184, N711);
and AND2 (N2823, N2817, N1368);
xor XOR2 (N2824, N2823, N355);
and AND3 (N2825, N2792, N1383, N2396);
buf BUF1 (N2826, N2816);
nor NOR2 (N2827, N2825, N2183);
and AND3 (N2828, N2824, N251, N1306);
buf BUF1 (N2829, N2828);
nor NOR2 (N2830, N2822, N1411);
buf BUF1 (N2831, N2820);
xor XOR2 (N2832, N2830, N1435);
buf BUF1 (N2833, N2829);
and AND3 (N2834, N2833, N2151, N926);
nor NOR4 (N2835, N2827, N560, N436, N575);
not NOT1 (N2836, N2835);
xor XOR2 (N2837, N2826, N866);
not NOT1 (N2838, N2818);
and AND4 (N2839, N2836, N450, N193, N1729);
buf BUF1 (N2840, N2831);
or OR2 (N2841, N2839, N991);
nor NOR4 (N2842, N2834, N1092, N1644, N410);
and AND2 (N2843, N2837, N2403);
or OR2 (N2844, N2842, N2208);
nor NOR4 (N2845, N2810, N792, N1454, N2641);
nor NOR4 (N2846, N2841, N646, N285, N2829);
not NOT1 (N2847, N2845);
buf BUF1 (N2848, N2843);
and AND4 (N2849, N2813, N1758, N453, N858);
nand NAND2 (N2850, N2846, N1651);
and AND3 (N2851, N2838, N1441, N111);
not NOT1 (N2852, N2847);
buf BUF1 (N2853, N2852);
buf BUF1 (N2854, N2844);
buf BUF1 (N2855, N2840);
or OR2 (N2856, N2851, N1251);
xor XOR2 (N2857, N2853, N103);
not NOT1 (N2858, N2832);
buf BUF1 (N2859, N2815);
buf BUF1 (N2860, N2858);
and AND3 (N2861, N2857, N1695, N2063);
or OR2 (N2862, N2791, N769);
and AND3 (N2863, N2856, N2344, N259);
nor NOR2 (N2864, N2855, N553);
or OR4 (N2865, N2854, N1805, N2296, N97);
buf BUF1 (N2866, N2861);
xor XOR2 (N2867, N2865, N548);
and AND2 (N2868, N2849, N1720);
xor XOR2 (N2869, N2860, N2050);
xor XOR2 (N2870, N2869, N780);
nand NAND4 (N2871, N2864, N717, N796, N1496);
nor NOR4 (N2872, N2863, N957, N2726, N774);
and AND3 (N2873, N2848, N1721, N286);
nor NOR4 (N2874, N2868, N2773, N2161, N1342);
not NOT1 (N2875, N2871);
or OR2 (N2876, N2850, N2302);
xor XOR2 (N2877, N2862, N2793);
nand NAND4 (N2878, N2876, N2569, N172, N2002);
xor XOR2 (N2879, N2873, N2286);
xor XOR2 (N2880, N2879, N1312);
and AND3 (N2881, N2877, N1042, N751);
and AND4 (N2882, N2859, N1245, N1263, N2758);
nand NAND2 (N2883, N2874, N452);
buf BUF1 (N2884, N2880);
or OR3 (N2885, N2881, N160, N2721);
not NOT1 (N2886, N2866);
nor NOR4 (N2887, N2882, N2221, N456, N2428);
nor NOR3 (N2888, N2885, N1080, N2062);
buf BUF1 (N2889, N2875);
buf BUF1 (N2890, N2886);
nand NAND2 (N2891, N2888, N542);
and AND4 (N2892, N2872, N81, N323, N605);
buf BUF1 (N2893, N2883);
or OR3 (N2894, N2891, N1938, N49);
nor NOR2 (N2895, N2878, N994);
and AND4 (N2896, N2895, N1228, N2686, N2158);
or OR3 (N2897, N2892, N11, N678);
or OR4 (N2898, N2870, N1979, N2357, N1316);
nor NOR4 (N2899, N2893, N2540, N2398, N620);
or OR3 (N2900, N2894, N1064, N324);
nor NOR3 (N2901, N2898, N1227, N473);
nand NAND2 (N2902, N2900, N453);
not NOT1 (N2903, N2897);
not NOT1 (N2904, N2899);
xor XOR2 (N2905, N2887, N954);
and AND2 (N2906, N2889, N1283);
nor NOR2 (N2907, N2867, N2817);
nor NOR2 (N2908, N2901, N82);
nand NAND2 (N2909, N2908, N619);
and AND2 (N2910, N2905, N749);
and AND3 (N2911, N2909, N361, N2680);
not NOT1 (N2912, N2903);
or OR3 (N2913, N2890, N1025, N2861);
nand NAND4 (N2914, N2907, N12, N1153, N651);
xor XOR2 (N2915, N2913, N2401);
buf BUF1 (N2916, N2902);
buf BUF1 (N2917, N2906);
nand NAND4 (N2918, N2917, N356, N2050, N2323);
nor NOR4 (N2919, N2915, N2065, N2184, N1225);
nand NAND2 (N2920, N2896, N2449);
and AND4 (N2921, N2914, N875, N2869, N2036);
nor NOR4 (N2922, N2911, N1836, N386, N317);
nor NOR3 (N2923, N2922, N286, N148);
xor XOR2 (N2924, N2920, N1525);
buf BUF1 (N2925, N2918);
nor NOR3 (N2926, N2921, N175, N1052);
and AND2 (N2927, N2924, N1334);
not NOT1 (N2928, N2884);
or OR3 (N2929, N2916, N491, N906);
or OR3 (N2930, N2910, N2691, N2921);
xor XOR2 (N2931, N2926, N1129);
or OR2 (N2932, N2912, N2142);
buf BUF1 (N2933, N2919);
or OR2 (N2934, N2928, N2920);
not NOT1 (N2935, N2904);
nor NOR4 (N2936, N2935, N2148, N2374, N1840);
not NOT1 (N2937, N2934);
xor XOR2 (N2938, N2936, N2228);
or OR3 (N2939, N2932, N804, N1703);
or OR4 (N2940, N2930, N1674, N2911, N1678);
buf BUF1 (N2941, N2925);
nand NAND4 (N2942, N2927, N2336, N425, N159);
xor XOR2 (N2943, N2938, N1188);
buf BUF1 (N2944, N2933);
buf BUF1 (N2945, N2942);
buf BUF1 (N2946, N2940);
not NOT1 (N2947, N2939);
nor NOR3 (N2948, N2929, N1870, N874);
nor NOR4 (N2949, N2946, N1275, N684, N383);
buf BUF1 (N2950, N2941);
or OR3 (N2951, N2944, N1428, N2730);
buf BUF1 (N2952, N2950);
buf BUF1 (N2953, N2948);
and AND2 (N2954, N2953, N739);
xor XOR2 (N2955, N2954, N107);
xor XOR2 (N2956, N2955, N2190);
xor XOR2 (N2957, N2947, N324);
and AND2 (N2958, N2943, N2795);
or OR4 (N2959, N2956, N586, N1548, N1084);
not NOT1 (N2960, N2945);
or OR4 (N2961, N2960, N1935, N1083, N2087);
xor XOR2 (N2962, N2949, N1434);
not NOT1 (N2963, N2959);
buf BUF1 (N2964, N2923);
or OR3 (N2965, N2958, N1308, N2277);
nand NAND4 (N2966, N2957, N1630, N326, N381);
nand NAND3 (N2967, N2951, N1925, N614);
xor XOR2 (N2968, N2965, N1440);
nor NOR2 (N2969, N2952, N1325);
nor NOR2 (N2970, N2931, N2172);
nand NAND3 (N2971, N2966, N931, N774);
buf BUF1 (N2972, N2937);
not NOT1 (N2973, N2971);
nor NOR4 (N2974, N2967, N1878, N973, N1372);
not NOT1 (N2975, N2972);
buf BUF1 (N2976, N2968);
xor XOR2 (N2977, N2970, N2820);
xor XOR2 (N2978, N2961, N2232);
nor NOR2 (N2979, N2977, N282);
nor NOR2 (N2980, N2963, N1675);
not NOT1 (N2981, N2976);
buf BUF1 (N2982, N2979);
buf BUF1 (N2983, N2964);
and AND4 (N2984, N2982, N1719, N284, N2040);
nor NOR2 (N2985, N2980, N1263);
xor XOR2 (N2986, N2981, N1658);
not NOT1 (N2987, N2973);
buf BUF1 (N2988, N2983);
buf BUF1 (N2989, N2987);
or OR2 (N2990, N2988, N2707);
nand NAND4 (N2991, N2989, N2385, N2970, N899);
nand NAND4 (N2992, N2991, N917, N1240, N2838);
xor XOR2 (N2993, N2990, N763);
buf BUF1 (N2994, N2978);
not NOT1 (N2995, N2985);
xor XOR2 (N2996, N2992, N1109);
xor XOR2 (N2997, N2993, N1990);
not NOT1 (N2998, N2984);
or OR2 (N2999, N2969, N2425);
not NOT1 (N3000, N2997);
xor XOR2 (N3001, N2995, N2366);
not NOT1 (N3002, N2986);
xor XOR2 (N3003, N2998, N961);
buf BUF1 (N3004, N3002);
nor NOR3 (N3005, N3001, N2444, N1686);
buf BUF1 (N3006, N2999);
or OR3 (N3007, N2975, N2589, N1679);
xor XOR2 (N3008, N2974, N2082);
or OR4 (N3009, N3005, N1244, N2801, N348);
or OR3 (N3010, N3006, N2276, N644);
not NOT1 (N3011, N3009);
buf BUF1 (N3012, N3010);
not NOT1 (N3013, N3011);
and AND3 (N3014, N3008, N732, N860);
nand NAND2 (N3015, N2962, N545);
or OR3 (N3016, N3004, N3008, N1112);
not NOT1 (N3017, N3000);
nand NAND4 (N3018, N3017, N1912, N2407, N1769);
nand NAND4 (N3019, N3013, N2538, N516, N2206);
nand NAND4 (N3020, N3019, N824, N25, N262);
and AND3 (N3021, N2994, N1833, N1335);
buf BUF1 (N3022, N3007);
nor NOR3 (N3023, N3003, N2217, N2832);
not NOT1 (N3024, N3021);
not NOT1 (N3025, N3018);
and AND3 (N3026, N3024, N573, N1607);
nand NAND4 (N3027, N3026, N1611, N2717, N201);
buf BUF1 (N3028, N3012);
not NOT1 (N3029, N3014);
nand NAND2 (N3030, N3020, N2329);
xor XOR2 (N3031, N3029, N2778);
not NOT1 (N3032, N3031);
nand NAND2 (N3033, N3022, N2671);
or OR4 (N3034, N2996, N1595, N759, N123);
not NOT1 (N3035, N3025);
xor XOR2 (N3036, N3034, N438);
xor XOR2 (N3037, N3036, N2223);
and AND3 (N3038, N3028, N2315, N1361);
buf BUF1 (N3039, N3033);
xor XOR2 (N3040, N3015, N2079);
or OR2 (N3041, N3023, N2550);
nor NOR4 (N3042, N3040, N2646, N2673, N1949);
nor NOR2 (N3043, N3027, N1210);
nor NOR4 (N3044, N3042, N2787, N436, N584);
not NOT1 (N3045, N3043);
nand NAND4 (N3046, N3039, N1980, N1199, N1501);
not NOT1 (N3047, N3041);
nor NOR3 (N3048, N3037, N2435, N1189);
and AND2 (N3049, N3048, N1432);
and AND2 (N3050, N3038, N695);
nand NAND3 (N3051, N3032, N2628, N983);
or OR2 (N3052, N3050, N1580);
and AND3 (N3053, N3049, N1738, N641);
not NOT1 (N3054, N3052);
nand NAND4 (N3055, N3051, N2799, N2787, N1553);
not NOT1 (N3056, N3054);
nand NAND3 (N3057, N3046, N602, N1499);
nand NAND2 (N3058, N3055, N1420);
not NOT1 (N3059, N3057);
nand NAND2 (N3060, N3059, N2880);
or OR2 (N3061, N3060, N20);
nor NOR2 (N3062, N3058, N18);
or OR3 (N3063, N3061, N1338, N1625);
buf BUF1 (N3064, N3053);
and AND4 (N3065, N3044, N1047, N1978, N2360);
xor XOR2 (N3066, N3030, N853);
nand NAND3 (N3067, N3063, N1749, N3014);
buf BUF1 (N3068, N3056);
nor NOR2 (N3069, N3016, N2240);
nor NOR3 (N3070, N3035, N1629, N2377);
not NOT1 (N3071, N3064);
nand NAND3 (N3072, N3068, N375, N1135);
not NOT1 (N3073, N3066);
nand NAND4 (N3074, N3067, N3046, N511, N1190);
nand NAND3 (N3075, N3072, N2163, N2317);
nor NOR3 (N3076, N3047, N2395, N691);
not NOT1 (N3077, N3062);
buf BUF1 (N3078, N3073);
and AND3 (N3079, N3045, N2520, N2636);
or OR3 (N3080, N3075, N2325, N1663);
and AND3 (N3081, N3079, N1995, N1756);
and AND2 (N3082, N3070, N440);
nand NAND3 (N3083, N3065, N755, N60);
and AND3 (N3084, N3082, N473, N1153);
and AND2 (N3085, N3081, N2029);
or OR4 (N3086, N3074, N2169, N2605, N2672);
xor XOR2 (N3087, N3071, N1999);
buf BUF1 (N3088, N3080);
nor NOR4 (N3089, N3083, N2752, N2627, N2979);
nor NOR4 (N3090, N3084, N689, N517, N2724);
nand NAND4 (N3091, N3088, N589, N2622, N1533);
buf BUF1 (N3092, N3091);
nor NOR4 (N3093, N3092, N1912, N619, N1788);
nor NOR3 (N3094, N3093, N2681, N592);
nand NAND3 (N3095, N3089, N109, N1162);
not NOT1 (N3096, N3077);
xor XOR2 (N3097, N3085, N1527);
not NOT1 (N3098, N3086);
nand NAND4 (N3099, N3095, N667, N1332, N2791);
nor NOR4 (N3100, N3087, N1343, N1755, N2220);
xor XOR2 (N3101, N3100, N149);
not NOT1 (N3102, N3097);
nor NOR2 (N3103, N3102, N243);
nor NOR4 (N3104, N3090, N2447, N1591, N2183);
or OR4 (N3105, N3103, N1818, N2162, N2639);
and AND3 (N3106, N3069, N2334, N852);
not NOT1 (N3107, N3101);
or OR2 (N3108, N3104, N446);
and AND4 (N3109, N3099, N2581, N634, N2776);
nor NOR3 (N3110, N3078, N73, N42);
xor XOR2 (N3111, N3110, N138);
and AND4 (N3112, N3105, N2793, N523, N184);
not NOT1 (N3113, N3098);
not NOT1 (N3114, N3112);
nand NAND4 (N3115, N3094, N2541, N1562, N514);
nor NOR2 (N3116, N3111, N565);
buf BUF1 (N3117, N3115);
or OR4 (N3118, N3116, N1128, N1277, N3052);
or OR4 (N3119, N3107, N2276, N697, N1891);
nor NOR4 (N3120, N3109, N3017, N158, N169);
xor XOR2 (N3121, N3114, N1909);
buf BUF1 (N3122, N3096);
nor NOR3 (N3123, N3120, N2498, N1727);
and AND2 (N3124, N3106, N901);
nor NOR3 (N3125, N3122, N1081, N1479);
and AND3 (N3126, N3076, N452, N1);
nand NAND3 (N3127, N3126, N892, N39);
and AND4 (N3128, N3118, N1167, N1153, N3073);
nor NOR3 (N3129, N3108, N474, N1353);
xor XOR2 (N3130, N3128, N1285);
xor XOR2 (N3131, N3124, N1598);
nor NOR4 (N3132, N3130, N1238, N1518, N477);
nor NOR3 (N3133, N3117, N1502, N1505);
and AND2 (N3134, N3127, N2608);
nand NAND4 (N3135, N3125, N1500, N2912, N3077);
buf BUF1 (N3136, N3134);
or OR3 (N3137, N3129, N673, N323);
buf BUF1 (N3138, N3113);
not NOT1 (N3139, N3138);
not NOT1 (N3140, N3139);
nor NOR2 (N3141, N3132, N1049);
buf BUF1 (N3142, N3137);
buf BUF1 (N3143, N3119);
nand NAND4 (N3144, N3123, N2815, N1279, N1111);
not NOT1 (N3145, N3140);
xor XOR2 (N3146, N3136, N1051);
nand NAND3 (N3147, N3142, N2, N2444);
and AND3 (N3148, N3135, N1466, N616);
nand NAND4 (N3149, N3133, N3050, N2060, N3040);
nor NOR3 (N3150, N3146, N1929, N2794);
buf BUF1 (N3151, N3121);
or OR4 (N3152, N3148, N2869, N524, N1198);
not NOT1 (N3153, N3151);
xor XOR2 (N3154, N3153, N86);
not NOT1 (N3155, N3145);
nand NAND2 (N3156, N3155, N2048);
nor NOR4 (N3157, N3156, N1852, N400, N880);
xor XOR2 (N3158, N3157, N2825);
and AND3 (N3159, N3149, N73, N1859);
buf BUF1 (N3160, N3152);
xor XOR2 (N3161, N3147, N1505);
xor XOR2 (N3162, N3131, N2193);
nand NAND2 (N3163, N3144, N954);
nand NAND2 (N3164, N3160, N455);
xor XOR2 (N3165, N3161, N1074);
nor NOR4 (N3166, N3141, N1677, N2836, N2849);
xor XOR2 (N3167, N3163, N678);
or OR2 (N3168, N3164, N2372);
and AND4 (N3169, N3167, N2112, N1892, N962);
and AND4 (N3170, N3150, N2975, N2385, N2571);
nand NAND3 (N3171, N3169, N1388, N1031);
and AND3 (N3172, N3154, N1294, N634);
xor XOR2 (N3173, N3166, N2449);
not NOT1 (N3174, N3159);
and AND4 (N3175, N3143, N1485, N3083, N245);
nand NAND2 (N3176, N3162, N2747);
buf BUF1 (N3177, N3168);
xor XOR2 (N3178, N3175, N2396);
nor NOR4 (N3179, N3171, N2008, N2996, N321);
buf BUF1 (N3180, N3174);
nand NAND4 (N3181, N3165, N1923, N2285, N2419);
and AND2 (N3182, N3176, N1769);
buf BUF1 (N3183, N3173);
and AND3 (N3184, N3181, N2764, N1961);
nand NAND2 (N3185, N3184, N1802);
nor NOR2 (N3186, N3185, N2979);
nand NAND2 (N3187, N3186, N1916);
not NOT1 (N3188, N3180);
nand NAND2 (N3189, N3177, N233);
not NOT1 (N3190, N3183);
or OR3 (N3191, N3158, N2920, N1961);
and AND4 (N3192, N3179, N1733, N1778, N852);
and AND3 (N3193, N3188, N1055, N378);
and AND2 (N3194, N3191, N1058);
or OR3 (N3195, N3178, N1102, N523);
xor XOR2 (N3196, N3193, N1462);
and AND3 (N3197, N3190, N2752, N1643);
and AND4 (N3198, N3172, N2726, N1879, N3030);
nor NOR3 (N3199, N3197, N1754, N1029);
nor NOR4 (N3200, N3196, N2302, N1117, N529);
xor XOR2 (N3201, N3194, N1324);
buf BUF1 (N3202, N3198);
not NOT1 (N3203, N3182);
xor XOR2 (N3204, N3189, N2513);
xor XOR2 (N3205, N3203, N584);
nor NOR2 (N3206, N3192, N2485);
not NOT1 (N3207, N3206);
nor NOR4 (N3208, N3199, N2781, N1798, N1210);
nor NOR2 (N3209, N3205, N291);
nand NAND3 (N3210, N3204, N719, N2058);
nor NOR4 (N3211, N3208, N2125, N1006, N3200);
xor XOR2 (N3212, N933, N2778);
xor XOR2 (N3213, N3209, N1658);
nand NAND2 (N3214, N3195, N1959);
nor NOR3 (N3215, N3211, N2194, N264);
xor XOR2 (N3216, N3207, N1129);
xor XOR2 (N3217, N3215, N958);
or OR4 (N3218, N3217, N3090, N426, N1896);
nor NOR2 (N3219, N3170, N2011);
buf BUF1 (N3220, N3212);
nor NOR4 (N3221, N3187, N73, N1980, N212);
or OR2 (N3222, N3221, N2862);
or OR4 (N3223, N3210, N1066, N847, N542);
buf BUF1 (N3224, N3216);
not NOT1 (N3225, N3219);
not NOT1 (N3226, N3201);
nor NOR4 (N3227, N3202, N635, N3159, N791);
buf BUF1 (N3228, N3226);
not NOT1 (N3229, N3227);
nor NOR2 (N3230, N3220, N1561);
or OR4 (N3231, N3229, N738, N1426, N2700);
nor NOR3 (N3232, N3222, N640, N2447);
nor NOR4 (N3233, N3231, N873, N965, N3176);
not NOT1 (N3234, N3213);
and AND3 (N3235, N3230, N2085, N2149);
and AND2 (N3236, N3232, N199);
or OR2 (N3237, N3235, N2573);
and AND2 (N3238, N3234, N961);
nand NAND3 (N3239, N3224, N1248, N3127);
nand NAND4 (N3240, N3233, N73, N1038, N981);
xor XOR2 (N3241, N3238, N1885);
and AND2 (N3242, N3240, N729);
xor XOR2 (N3243, N3228, N867);
xor XOR2 (N3244, N3239, N2267);
and AND4 (N3245, N3236, N2998, N616, N479);
xor XOR2 (N3246, N3225, N1574);
or OR2 (N3247, N3241, N2429);
nor NOR3 (N3248, N3214, N1902, N523);
xor XOR2 (N3249, N3242, N946);
or OR2 (N3250, N3243, N2329);
and AND3 (N3251, N3248, N558, N298);
nor NOR3 (N3252, N3249, N722, N462);
xor XOR2 (N3253, N3247, N2767);
xor XOR2 (N3254, N3251, N2329);
nor NOR4 (N3255, N3244, N3119, N1844, N462);
buf BUF1 (N3256, N3218);
buf BUF1 (N3257, N3237);
or OR2 (N3258, N3257, N1819);
buf BUF1 (N3259, N3246);
nand NAND3 (N3260, N3253, N3185, N114);
xor XOR2 (N3261, N3250, N2821);
nor NOR4 (N3262, N3261, N2447, N1124, N2452);
or OR2 (N3263, N3256, N97);
buf BUF1 (N3264, N3260);
or OR4 (N3265, N3255, N1816, N1689, N529);
and AND3 (N3266, N3263, N1504, N2121);
nand NAND4 (N3267, N3262, N353, N2493, N836);
buf BUF1 (N3268, N3252);
nor NOR3 (N3269, N3254, N352, N401);
buf BUF1 (N3270, N3269);
xor XOR2 (N3271, N3267, N2409);
and AND3 (N3272, N3271, N2877, N2130);
and AND3 (N3273, N3266, N1762, N450);
buf BUF1 (N3274, N3265);
not NOT1 (N3275, N3259);
nor NOR3 (N3276, N3258, N2849, N1074);
not NOT1 (N3277, N3264);
not NOT1 (N3278, N3276);
nand NAND4 (N3279, N3272, N2578, N2463, N879);
buf BUF1 (N3280, N3279);
or OR2 (N3281, N3277, N1897);
nor NOR2 (N3282, N3274, N1258);
and AND4 (N3283, N3280, N3237, N676, N501);
nor NOR3 (N3284, N3245, N1179, N529);
buf BUF1 (N3285, N3275);
buf BUF1 (N3286, N3270);
xor XOR2 (N3287, N3278, N1360);
and AND2 (N3288, N3284, N1332);
nor NOR2 (N3289, N3281, N1731);
nand NAND3 (N3290, N3287, N1445, N2137);
xor XOR2 (N3291, N3223, N113);
not NOT1 (N3292, N3289);
and AND2 (N3293, N3290, N2109);
buf BUF1 (N3294, N3283);
not NOT1 (N3295, N3294);
xor XOR2 (N3296, N3291, N2182);
and AND2 (N3297, N3286, N496);
nand NAND2 (N3298, N3268, N630);
xor XOR2 (N3299, N3293, N372);
and AND4 (N3300, N3292, N2839, N1656, N1532);
nor NOR3 (N3301, N3296, N2470, N1623);
not NOT1 (N3302, N3300);
nor NOR4 (N3303, N3301, N315, N985, N847);
nand NAND2 (N3304, N3303, N201);
or OR3 (N3305, N3285, N565, N570);
xor XOR2 (N3306, N3304, N576);
buf BUF1 (N3307, N3297);
nand NAND2 (N3308, N3273, N3109);
or OR4 (N3309, N3308, N1492, N2992, N801);
or OR2 (N3310, N3309, N700);
or OR3 (N3311, N3305, N2932, N1606);
xor XOR2 (N3312, N3295, N416);
or OR3 (N3313, N3298, N3291, N2778);
not NOT1 (N3314, N3299);
not NOT1 (N3315, N3306);
and AND2 (N3316, N3314, N84);
nand NAND3 (N3317, N3288, N759, N3311);
not NOT1 (N3318, N3220);
nand NAND2 (N3319, N3313, N110);
or OR3 (N3320, N3318, N1679, N269);
xor XOR2 (N3321, N3317, N3040);
xor XOR2 (N3322, N3315, N1511);
not NOT1 (N3323, N3320);
nand NAND4 (N3324, N3310, N2291, N1910, N3262);
xor XOR2 (N3325, N3307, N3007);
xor XOR2 (N3326, N3319, N111);
nor NOR3 (N3327, N3324, N1225, N1829);
nor NOR2 (N3328, N3302, N204);
buf BUF1 (N3329, N3322);
nand NAND4 (N3330, N3282, N327, N307, N2011);
nand NAND2 (N3331, N3328, N2928);
and AND4 (N3332, N3323, N363, N2997, N3180);
nand NAND3 (N3333, N3326, N3134, N2996);
nor NOR2 (N3334, N3331, N1660);
nand NAND4 (N3335, N3332, N1233, N2037, N1625);
and AND2 (N3336, N3327, N1024);
and AND3 (N3337, N3312, N2382, N2291);
nor NOR2 (N3338, N3337, N3089);
buf BUF1 (N3339, N3330);
nand NAND2 (N3340, N3333, N2089);
xor XOR2 (N3341, N3316, N2223);
xor XOR2 (N3342, N3340, N2362);
and AND3 (N3343, N3321, N146, N295);
xor XOR2 (N3344, N3336, N2980);
nor NOR4 (N3345, N3343, N850, N2240, N308);
nand NAND2 (N3346, N3339, N902);
or OR3 (N3347, N3335, N293, N1098);
not NOT1 (N3348, N3334);
nand NAND4 (N3349, N3346, N1152, N3234, N2965);
not NOT1 (N3350, N3329);
not NOT1 (N3351, N3325);
xor XOR2 (N3352, N3344, N582);
not NOT1 (N3353, N3349);
nand NAND3 (N3354, N3338, N330, N2043);
buf BUF1 (N3355, N3342);
xor XOR2 (N3356, N3350, N1863);
or OR4 (N3357, N3345, N1853, N1735, N512);
and AND4 (N3358, N3341, N844, N736, N387);
nor NOR3 (N3359, N3356, N690, N1007);
or OR3 (N3360, N3347, N3015, N2941);
or OR4 (N3361, N3351, N2879, N2434, N1122);
nand NAND4 (N3362, N3353, N1930, N980, N604);
nand NAND2 (N3363, N3352, N296);
not NOT1 (N3364, N3363);
not NOT1 (N3365, N3355);
not NOT1 (N3366, N3362);
xor XOR2 (N3367, N3358, N1389);
xor XOR2 (N3368, N3360, N2169);
nor NOR4 (N3369, N3361, N2365, N2182, N560);
nand NAND3 (N3370, N3354, N2396, N1623);
buf BUF1 (N3371, N3364);
or OR3 (N3372, N3357, N3322, N1907);
xor XOR2 (N3373, N3368, N2692);
nand NAND4 (N3374, N3370, N3107, N762, N3101);
or OR2 (N3375, N3374, N960);
not NOT1 (N3376, N3372);
buf BUF1 (N3377, N3376);
buf BUF1 (N3378, N3371);
not NOT1 (N3379, N3377);
xor XOR2 (N3380, N3348, N2722);
buf BUF1 (N3381, N3373);
or OR3 (N3382, N3366, N2242, N423);
buf BUF1 (N3383, N3375);
not NOT1 (N3384, N3382);
not NOT1 (N3385, N3379);
buf BUF1 (N3386, N3365);
not NOT1 (N3387, N3367);
or OR4 (N3388, N3369, N31, N752, N2322);
not NOT1 (N3389, N3381);
not NOT1 (N3390, N3389);
or OR4 (N3391, N3380, N2228, N2992, N1153);
not NOT1 (N3392, N3384);
and AND2 (N3393, N3385, N734);
or OR3 (N3394, N3393, N716, N2899);
nand NAND2 (N3395, N3387, N3073);
nand NAND3 (N3396, N3359, N828, N1406);
buf BUF1 (N3397, N3395);
and AND4 (N3398, N3388, N2949, N26, N1868);
nand NAND4 (N3399, N3396, N2546, N2800, N1496);
nor NOR4 (N3400, N3378, N2044, N935, N923);
nand NAND2 (N3401, N3386, N3031);
buf BUF1 (N3402, N3398);
xor XOR2 (N3403, N3394, N743);
nor NOR4 (N3404, N3392, N1528, N2685, N281);
not NOT1 (N3405, N3403);
not NOT1 (N3406, N3397);
or OR3 (N3407, N3400, N2016, N781);
nor NOR3 (N3408, N3407, N1606, N678);
nor NOR4 (N3409, N3401, N1950, N2986, N2456);
nand NAND3 (N3410, N3405, N2733, N2841);
xor XOR2 (N3411, N3399, N656);
buf BUF1 (N3412, N3409);
not NOT1 (N3413, N3402);
or OR4 (N3414, N3412, N1215, N423, N3218);
or OR4 (N3415, N3404, N3232, N2621, N3194);
or OR3 (N3416, N3414, N3337, N1488);
not NOT1 (N3417, N3390);
and AND3 (N3418, N3406, N3417, N2912);
or OR2 (N3419, N2776, N2884);
and AND2 (N3420, N3408, N1920);
xor XOR2 (N3421, N3419, N2662);
and AND4 (N3422, N3420, N1441, N825, N51);
nand NAND4 (N3423, N3418, N983, N2603, N1733);
nand NAND3 (N3424, N3410, N442, N2939);
xor XOR2 (N3425, N3383, N2695);
nor NOR2 (N3426, N3424, N1864);
xor XOR2 (N3427, N3416, N810);
xor XOR2 (N3428, N3422, N1460);
not NOT1 (N3429, N3426);
xor XOR2 (N3430, N3413, N2359);
and AND4 (N3431, N3423, N781, N3107, N35);
not NOT1 (N3432, N3429);
not NOT1 (N3433, N3432);
buf BUF1 (N3434, N3415);
buf BUF1 (N3435, N3411);
xor XOR2 (N3436, N3391, N879);
and AND4 (N3437, N3434, N488, N309, N2564);
xor XOR2 (N3438, N3435, N2060);
xor XOR2 (N3439, N3425, N1046);
nand NAND2 (N3440, N3431, N2066);
and AND4 (N3441, N3421, N2469, N133, N1595);
not NOT1 (N3442, N3430);
not NOT1 (N3443, N3436);
nand NAND2 (N3444, N3441, N1929);
nand NAND3 (N3445, N3440, N3296, N104);
not NOT1 (N3446, N3442);
xor XOR2 (N3447, N3427, N2249);
not NOT1 (N3448, N3443);
not NOT1 (N3449, N3437);
nor NOR4 (N3450, N3447, N2789, N261, N729);
xor XOR2 (N3451, N3445, N97);
nand NAND2 (N3452, N3439, N1519);
xor XOR2 (N3453, N3433, N2706);
and AND2 (N3454, N3450, N2193);
xor XOR2 (N3455, N3446, N2989);
or OR3 (N3456, N3454, N2833, N1000);
nor NOR3 (N3457, N3448, N2197, N1771);
not NOT1 (N3458, N3444);
buf BUF1 (N3459, N3457);
xor XOR2 (N3460, N3458, N3227);
not NOT1 (N3461, N3460);
or OR2 (N3462, N3451, N209);
nand NAND2 (N3463, N3459, N2651);
or OR2 (N3464, N3455, N1966);
or OR3 (N3465, N3462, N270, N2587);
xor XOR2 (N3466, N3438, N3398);
nand NAND2 (N3467, N3461, N941);
xor XOR2 (N3468, N3456, N788);
not NOT1 (N3469, N3467);
buf BUF1 (N3470, N3469);
or OR3 (N3471, N3449, N2696, N493);
nor NOR2 (N3472, N3466, N2083);
buf BUF1 (N3473, N3453);
buf BUF1 (N3474, N3463);
nand NAND4 (N3475, N3474, N2967, N2563, N538);
nand NAND2 (N3476, N3470, N3106);
buf BUF1 (N3477, N3428);
nand NAND4 (N3478, N3472, N3114, N1316, N1035);
or OR4 (N3479, N3465, N1409, N3143, N3266);
nand NAND3 (N3480, N3478, N66, N2442);
nand NAND3 (N3481, N3479, N261, N1707);
and AND2 (N3482, N3480, N2316);
xor XOR2 (N3483, N3476, N2144);
nand NAND3 (N3484, N3483, N229, N1422);
buf BUF1 (N3485, N3484);
nand NAND3 (N3486, N3481, N767, N739);
nor NOR3 (N3487, N3475, N361, N2461);
and AND2 (N3488, N3487, N1555);
xor XOR2 (N3489, N3468, N648);
or OR4 (N3490, N3452, N2994, N1033, N1192);
not NOT1 (N3491, N3486);
or OR2 (N3492, N3490, N753);
and AND4 (N3493, N3471, N1596, N734, N2765);
not NOT1 (N3494, N3493);
nand NAND3 (N3495, N3491, N2275, N674);
xor XOR2 (N3496, N3488, N1357);
xor XOR2 (N3497, N3494, N3017);
xor XOR2 (N3498, N3482, N1367);
nor NOR3 (N3499, N3498, N305, N2538);
nand NAND3 (N3500, N3496, N3148, N1271);
not NOT1 (N3501, N3495);
not NOT1 (N3502, N3499);
not NOT1 (N3503, N3492);
nand NAND2 (N3504, N3497, N2925);
or OR3 (N3505, N3500, N2813, N3500);
buf BUF1 (N3506, N3477);
nor NOR4 (N3507, N3503, N853, N2760, N1947);
xor XOR2 (N3508, N3504, N2604);
nand NAND4 (N3509, N3506, N344, N361, N1804);
xor XOR2 (N3510, N3464, N606);
or OR4 (N3511, N3485, N368, N2073, N1122);
and AND3 (N3512, N3489, N1133, N2459);
xor XOR2 (N3513, N3512, N3310);
and AND2 (N3514, N3507, N1400);
not NOT1 (N3515, N3509);
not NOT1 (N3516, N3513);
and AND3 (N3517, N3514, N2649, N1629);
nand NAND2 (N3518, N3517, N124);
nor NOR4 (N3519, N3473, N3189, N3049, N1462);
nand NAND3 (N3520, N3519, N1301, N1844);
nand NAND3 (N3521, N3505, N1743, N2714);
nor NOR3 (N3522, N3515, N1203, N3343);
xor XOR2 (N3523, N3502, N1482);
not NOT1 (N3524, N3516);
buf BUF1 (N3525, N3521);
not NOT1 (N3526, N3510);
not NOT1 (N3527, N3501);
or OR3 (N3528, N3511, N1093, N1860);
not NOT1 (N3529, N3527);
buf BUF1 (N3530, N3508);
not NOT1 (N3531, N3528);
nor NOR4 (N3532, N3530, N1414, N1658, N1085);
not NOT1 (N3533, N3523);
xor XOR2 (N3534, N3520, N3334);
not NOT1 (N3535, N3524);
or OR3 (N3536, N3531, N3143, N65);
or OR2 (N3537, N3533, N2419);
buf BUF1 (N3538, N3536);
nand NAND4 (N3539, N3535, N448, N1774, N2247);
nand NAND2 (N3540, N3529, N16);
buf BUF1 (N3541, N3525);
buf BUF1 (N3542, N3540);
nor NOR4 (N3543, N3518, N830, N86, N2976);
nor NOR3 (N3544, N3539, N1885, N2535);
nor NOR4 (N3545, N3522, N2721, N3513, N2925);
not NOT1 (N3546, N3537);
xor XOR2 (N3547, N3526, N1836);
and AND4 (N3548, N3546, N483, N1999, N2738);
and AND4 (N3549, N3548, N1009, N1051, N3125);
buf BUF1 (N3550, N3549);
nand NAND2 (N3551, N3541, N3486);
nand NAND4 (N3552, N3551, N872, N330, N918);
not NOT1 (N3553, N3542);
xor XOR2 (N3554, N3538, N2787);
or OR3 (N3555, N3553, N2447, N2213);
nor NOR2 (N3556, N3552, N3120);
nor NOR3 (N3557, N3554, N2304, N1787);
or OR2 (N3558, N3555, N3049);
or OR4 (N3559, N3556, N242, N1370, N2762);
buf BUF1 (N3560, N3558);
or OR2 (N3561, N3545, N367);
buf BUF1 (N3562, N3547);
xor XOR2 (N3563, N3561, N2566);
xor XOR2 (N3564, N3534, N426);
and AND3 (N3565, N3563, N1620, N715);
buf BUF1 (N3566, N3544);
or OR4 (N3567, N3543, N2533, N2352, N1292);
or OR4 (N3568, N3562, N3206, N1476, N141);
buf BUF1 (N3569, N3568);
nand NAND2 (N3570, N3532, N39);
nand NAND3 (N3571, N3570, N2491, N1256);
not NOT1 (N3572, N3564);
buf BUF1 (N3573, N3565);
not NOT1 (N3574, N3557);
and AND3 (N3575, N3571, N592, N1916);
or OR3 (N3576, N3575, N918, N3151);
and AND2 (N3577, N3572, N3155);
nor NOR3 (N3578, N3574, N500, N3041);
not NOT1 (N3579, N3560);
not NOT1 (N3580, N3559);
nor NOR3 (N3581, N3566, N554, N245);
or OR4 (N3582, N3577, N1645, N3568, N2365);
nand NAND2 (N3583, N3569, N1678);
buf BUF1 (N3584, N3582);
and AND4 (N3585, N3578, N2226, N1284, N338);
xor XOR2 (N3586, N3550, N1605);
not NOT1 (N3587, N3580);
xor XOR2 (N3588, N3567, N185);
buf BUF1 (N3589, N3573);
xor XOR2 (N3590, N3589, N2004);
not NOT1 (N3591, N3576);
nand NAND3 (N3592, N3590, N1984, N3326);
or OR4 (N3593, N3587, N3348, N633, N1941);
buf BUF1 (N3594, N3583);
and AND2 (N3595, N3588, N2810);
and AND4 (N3596, N3585, N3590, N3547, N1502);
nand NAND2 (N3597, N3594, N1569);
nand NAND4 (N3598, N3597, N1931, N2367, N1109);
nand NAND4 (N3599, N3595, N2086, N37, N3475);
xor XOR2 (N3600, N3596, N119);
nand NAND4 (N3601, N3592, N3153, N3474, N1837);
not NOT1 (N3602, N3591);
xor XOR2 (N3603, N3600, N552);
nand NAND4 (N3604, N3603, N2783, N740, N358);
not NOT1 (N3605, N3604);
nor NOR2 (N3606, N3602, N2249);
or OR4 (N3607, N3599, N1187, N3595, N3197);
and AND4 (N3608, N3579, N2311, N1725, N1914);
nor NOR2 (N3609, N3593, N440);
and AND4 (N3610, N3608, N341, N1070, N165);
buf BUF1 (N3611, N3606);
or OR2 (N3612, N3607, N3138);
nand NAND4 (N3613, N3611, N1533, N3108, N3527);
xor XOR2 (N3614, N3581, N93);
buf BUF1 (N3615, N3613);
xor XOR2 (N3616, N3615, N2564);
xor XOR2 (N3617, N3598, N1182);
nor NOR2 (N3618, N3605, N1921);
or OR2 (N3619, N3616, N777);
nand NAND4 (N3620, N3614, N2062, N557, N2254);
or OR2 (N3621, N3609, N539);
nand NAND4 (N3622, N3620, N1093, N2191, N2706);
or OR2 (N3623, N3617, N2004);
or OR2 (N3624, N3584, N2038);
not NOT1 (N3625, N3623);
and AND3 (N3626, N3586, N2316, N497);
buf BUF1 (N3627, N3619);
nor NOR2 (N3628, N3610, N1267);
and AND2 (N3629, N3625, N2067);
nand NAND3 (N3630, N3627, N568, N1395);
or OR2 (N3631, N3626, N607);
or OR2 (N3632, N3631, N1364);
nand NAND2 (N3633, N3612, N2853);
nand NAND3 (N3634, N3622, N2752, N3113);
not NOT1 (N3635, N3632);
buf BUF1 (N3636, N3635);
not NOT1 (N3637, N3634);
xor XOR2 (N3638, N3618, N2490);
or OR3 (N3639, N3628, N935, N1493);
and AND3 (N3640, N3621, N3272, N2261);
buf BUF1 (N3641, N3629);
or OR3 (N3642, N3624, N2731, N2668);
or OR3 (N3643, N3633, N2977, N61);
not NOT1 (N3644, N3636);
nor NOR4 (N3645, N3644, N607, N2003, N1296);
nor NOR2 (N3646, N3643, N2525);
xor XOR2 (N3647, N3638, N58);
xor XOR2 (N3648, N3637, N546);
not NOT1 (N3649, N3601);
not NOT1 (N3650, N3646);
xor XOR2 (N3651, N3645, N2267);
not NOT1 (N3652, N3642);
or OR2 (N3653, N3651, N2566);
xor XOR2 (N3654, N3630, N2209);
not NOT1 (N3655, N3648);
nand NAND2 (N3656, N3652, N1946);
not NOT1 (N3657, N3655);
nand NAND2 (N3658, N3657, N517);
and AND3 (N3659, N3639, N2090, N1766);
or OR2 (N3660, N3649, N1252);
buf BUF1 (N3661, N3647);
buf BUF1 (N3662, N3659);
and AND2 (N3663, N3640, N1361);
buf BUF1 (N3664, N3653);
nand NAND3 (N3665, N3650, N3538, N1106);
nand NAND4 (N3666, N3641, N651, N1281, N3485);
and AND4 (N3667, N3656, N307, N2237, N1034);
nor NOR3 (N3668, N3664, N3546, N3563);
nor NOR3 (N3669, N3668, N2115, N1721);
nand NAND3 (N3670, N3667, N3250, N686);
not NOT1 (N3671, N3661);
and AND3 (N3672, N3669, N86, N2612);
nor NOR2 (N3673, N3670, N1689);
and AND3 (N3674, N3673, N963, N2080);
not NOT1 (N3675, N3674);
nand NAND3 (N3676, N3663, N1254, N2459);
xor XOR2 (N3677, N3671, N3586);
and AND4 (N3678, N3676, N1373, N1476, N907);
xor XOR2 (N3679, N3660, N2098);
nor NOR4 (N3680, N3679, N2077, N1144, N2540);
xor XOR2 (N3681, N3675, N3037);
and AND4 (N3682, N3662, N431, N2167, N234);
buf BUF1 (N3683, N3665);
nor NOR4 (N3684, N3666, N1993, N2468, N975);
xor XOR2 (N3685, N3682, N79);
or OR4 (N3686, N3654, N1575, N2361, N3571);
and AND3 (N3687, N3683, N3500, N3133);
and AND2 (N3688, N3681, N252);
nor NOR2 (N3689, N3687, N2275);
nand NAND3 (N3690, N3658, N3060, N3673);
and AND2 (N3691, N3690, N3497);
and AND4 (N3692, N3685, N2772, N68, N372);
and AND4 (N3693, N3678, N527, N2859, N2496);
or OR3 (N3694, N3677, N2366, N976);
buf BUF1 (N3695, N3691);
xor XOR2 (N3696, N3692, N616);
not NOT1 (N3697, N3693);
xor XOR2 (N3698, N3672, N1442);
nand NAND4 (N3699, N3698, N1182, N2245, N1302);
and AND3 (N3700, N3694, N1546, N3056);
and AND4 (N3701, N3699, N3034, N456, N423);
and AND4 (N3702, N3688, N1119, N3693, N614);
xor XOR2 (N3703, N3702, N143);
buf BUF1 (N3704, N3684);
and AND4 (N3705, N3695, N2362, N104, N1530);
buf BUF1 (N3706, N3701);
and AND4 (N3707, N3705, N1417, N1124, N290);
buf BUF1 (N3708, N3703);
or OR4 (N3709, N3689, N75, N342, N1397);
and AND4 (N3710, N3680, N1336, N26, N2678);
nor NOR3 (N3711, N3697, N3533, N519);
buf BUF1 (N3712, N3700);
nor NOR2 (N3713, N3704, N3608);
xor XOR2 (N3714, N3712, N2832);
or OR3 (N3715, N3696, N1305, N2141);
buf BUF1 (N3716, N3714);
or OR4 (N3717, N3713, N3221, N1737, N2382);
buf BUF1 (N3718, N3706);
nand NAND4 (N3719, N3707, N1542, N711, N3708);
not NOT1 (N3720, N2023);
nand NAND3 (N3721, N3709, N3081, N834);
not NOT1 (N3722, N3715);
not NOT1 (N3723, N3716);
and AND3 (N3724, N3717, N1945, N506);
nand NAND3 (N3725, N3711, N2284, N2595);
buf BUF1 (N3726, N3724);
xor XOR2 (N3727, N3718, N3136);
and AND4 (N3728, N3725, N3684, N244, N1875);
xor XOR2 (N3729, N3721, N2995);
buf BUF1 (N3730, N3710);
xor XOR2 (N3731, N3726, N2166);
nor NOR4 (N3732, N3729, N1759, N1524, N2933);
nor NOR4 (N3733, N3731, N1285, N1512, N3670);
nand NAND2 (N3734, N3730, N3246);
nor NOR3 (N3735, N3686, N880, N973);
nor NOR4 (N3736, N3734, N2098, N3219, N2702);
buf BUF1 (N3737, N3728);
or OR4 (N3738, N3736, N3477, N3136, N2439);
or OR2 (N3739, N3719, N441);
xor XOR2 (N3740, N3735, N1901);
or OR3 (N3741, N3720, N769, N2709);
nor NOR3 (N3742, N3723, N882, N2273);
xor XOR2 (N3743, N3740, N3272);
or OR4 (N3744, N3741, N3358, N1597, N1360);
nand NAND3 (N3745, N3743, N1797, N2766);
or OR4 (N3746, N3722, N1881, N2011, N1655);
xor XOR2 (N3747, N3737, N3395);
buf BUF1 (N3748, N3738);
or OR4 (N3749, N3748, N1959, N1121, N804);
buf BUF1 (N3750, N3749);
xor XOR2 (N3751, N3739, N3150);
not NOT1 (N3752, N3742);
and AND2 (N3753, N3752, N2776);
and AND2 (N3754, N3753, N893);
nor NOR4 (N3755, N3744, N2574, N3639, N2702);
nor NOR2 (N3756, N3732, N2419);
nand NAND2 (N3757, N3750, N423);
or OR3 (N3758, N3755, N1508, N142);
not NOT1 (N3759, N3727);
not NOT1 (N3760, N3759);
buf BUF1 (N3761, N3760);
buf BUF1 (N3762, N3754);
and AND3 (N3763, N3733, N829, N3171);
or OR4 (N3764, N3758, N1523, N820, N1230);
xor XOR2 (N3765, N3762, N2833);
and AND3 (N3766, N3751, N3401, N301);
not NOT1 (N3767, N3761);
nand NAND2 (N3768, N3765, N2831);
not NOT1 (N3769, N3745);
buf BUF1 (N3770, N3756);
or OR2 (N3771, N3764, N3571);
nand NAND2 (N3772, N3747, N2144);
nand NAND3 (N3773, N3766, N2554, N1688);
or OR3 (N3774, N3763, N222, N2105);
nand NAND4 (N3775, N3772, N2996, N1346, N674);
xor XOR2 (N3776, N3769, N758);
buf BUF1 (N3777, N3771);
not NOT1 (N3778, N3768);
xor XOR2 (N3779, N3774, N890);
buf BUF1 (N3780, N3777);
and AND2 (N3781, N3767, N3089);
xor XOR2 (N3782, N3746, N1184);
and AND2 (N3783, N3782, N3154);
xor XOR2 (N3784, N3783, N2871);
or OR4 (N3785, N3770, N815, N283, N3698);
nor NOR3 (N3786, N3779, N3056, N1372);
or OR3 (N3787, N3785, N3336, N3306);
not NOT1 (N3788, N3780);
xor XOR2 (N3789, N3757, N2342);
or OR2 (N3790, N3786, N2207);
buf BUF1 (N3791, N3788);
or OR2 (N3792, N3791, N372);
nor NOR3 (N3793, N3781, N3374, N777);
nor NOR4 (N3794, N3773, N2795, N956, N2729);
nand NAND2 (N3795, N3778, N9);
nand NAND4 (N3796, N3793, N3556, N3594, N1616);
xor XOR2 (N3797, N3796, N1446);
xor XOR2 (N3798, N3776, N345);
not NOT1 (N3799, N3775);
nand NAND4 (N3800, N3799, N2984, N260, N3764);
xor XOR2 (N3801, N3789, N1119);
xor XOR2 (N3802, N3784, N2897);
nor NOR2 (N3803, N3795, N1819);
nor NOR4 (N3804, N3801, N2415, N602, N733);
or OR3 (N3805, N3798, N611, N3146);
nor NOR4 (N3806, N3790, N2973, N2885, N3402);
buf BUF1 (N3807, N3802);
or OR3 (N3808, N3792, N1303, N3327);
or OR3 (N3809, N3800, N3086, N3573);
not NOT1 (N3810, N3787);
or OR3 (N3811, N3797, N2114, N1217);
or OR4 (N3812, N3803, N70, N537, N622);
buf BUF1 (N3813, N3805);
xor XOR2 (N3814, N3809, N62);
and AND4 (N3815, N3814, N3358, N1945, N2663);
nand NAND3 (N3816, N3794, N1748, N1116);
and AND3 (N3817, N3807, N3594, N2791);
buf BUF1 (N3818, N3811);
xor XOR2 (N3819, N3815, N2511);
buf BUF1 (N3820, N3816);
nor NOR4 (N3821, N3817, N3110, N2843, N1443);
xor XOR2 (N3822, N3806, N593);
and AND3 (N3823, N3808, N3188, N3609);
nor NOR4 (N3824, N3822, N2928, N2638, N2662);
not NOT1 (N3825, N3820);
xor XOR2 (N3826, N3810, N962);
buf BUF1 (N3827, N3824);
nor NOR4 (N3828, N3825, N2324, N804, N3648);
nand NAND3 (N3829, N3813, N3210, N3517);
or OR2 (N3830, N3828, N3613);
nor NOR2 (N3831, N3826, N247);
xor XOR2 (N3832, N3831, N569);
and AND2 (N3833, N3823, N2632);
nand NAND3 (N3834, N3833, N3531, N113);
nor NOR4 (N3835, N3818, N2801, N378, N3019);
and AND2 (N3836, N3804, N1818);
or OR4 (N3837, N3827, N1608, N26, N3080);
not NOT1 (N3838, N3829);
nand NAND3 (N3839, N3819, N1170, N104);
xor XOR2 (N3840, N3830, N1743);
xor XOR2 (N3841, N3812, N2559);
nand NAND2 (N3842, N3821, N2113);
nor NOR3 (N3843, N3839, N1395, N564);
xor XOR2 (N3844, N3838, N2078);
or OR3 (N3845, N3835, N260, N3576);
xor XOR2 (N3846, N3837, N184);
nand NAND2 (N3847, N3836, N1192);
nor NOR2 (N3848, N3842, N2147);
nand NAND3 (N3849, N3834, N1884, N3599);
and AND2 (N3850, N3832, N1863);
xor XOR2 (N3851, N3850, N1909);
nor NOR4 (N3852, N3846, N2944, N2268, N3707);
or OR4 (N3853, N3852, N1513, N3813, N1658);
and AND3 (N3854, N3847, N3190, N708);
and AND3 (N3855, N3841, N1608, N2735);
xor XOR2 (N3856, N3851, N2623);
not NOT1 (N3857, N3845);
nor NOR2 (N3858, N3848, N339);
nor NOR2 (N3859, N3843, N241);
nand NAND3 (N3860, N3855, N3485, N2487);
buf BUF1 (N3861, N3854);
buf BUF1 (N3862, N3860);
xor XOR2 (N3863, N3862, N1036);
or OR2 (N3864, N3853, N388);
buf BUF1 (N3865, N3863);
nor NOR2 (N3866, N3864, N3415);
xor XOR2 (N3867, N3858, N264);
xor XOR2 (N3868, N3856, N2324);
not NOT1 (N3869, N3867);
nand NAND3 (N3870, N3861, N2243, N1923);
nor NOR2 (N3871, N3844, N187);
xor XOR2 (N3872, N3857, N2577);
and AND3 (N3873, N3868, N2494, N2155);
buf BUF1 (N3874, N3872);
buf BUF1 (N3875, N3866);
not NOT1 (N3876, N3865);
not NOT1 (N3877, N3876);
buf BUF1 (N3878, N3875);
xor XOR2 (N3879, N3869, N895);
nand NAND4 (N3880, N3871, N1279, N84, N781);
or OR3 (N3881, N3840, N1366, N3518);
buf BUF1 (N3882, N3878);
or OR4 (N3883, N3882, N638, N3554, N30);
buf BUF1 (N3884, N3877);
or OR3 (N3885, N3873, N50, N2964);
and AND3 (N3886, N3870, N937, N1049);
nor NOR3 (N3887, N3874, N3701, N1621);
buf BUF1 (N3888, N3887);
buf BUF1 (N3889, N3881);
nand NAND2 (N3890, N3888, N1430);
and AND4 (N3891, N3849, N1167, N231, N136);
nor NOR4 (N3892, N3891, N1461, N1451, N1593);
and AND3 (N3893, N3886, N3508, N3090);
xor XOR2 (N3894, N3889, N2168);
and AND3 (N3895, N3885, N3759, N3038);
nand NAND2 (N3896, N3890, N1449);
and AND2 (N3897, N3896, N1541);
or OR2 (N3898, N3859, N1759);
buf BUF1 (N3899, N3894);
not NOT1 (N3900, N3883);
buf BUF1 (N3901, N3893);
or OR3 (N3902, N3879, N2512, N768);
or OR4 (N3903, N3880, N719, N629, N1294);
and AND2 (N3904, N3884, N3713);
not NOT1 (N3905, N3897);
buf BUF1 (N3906, N3901);
nand NAND2 (N3907, N3904, N2453);
nor NOR2 (N3908, N3906, N127);
not NOT1 (N3909, N3902);
or OR4 (N3910, N3892, N2128, N213, N2330);
nand NAND2 (N3911, N3908, N2940);
not NOT1 (N3912, N3907);
nand NAND3 (N3913, N3903, N2765, N1545);
xor XOR2 (N3914, N3905, N2933);
or OR4 (N3915, N3914, N1343, N3647, N1163);
nor NOR3 (N3916, N3900, N1906, N715);
xor XOR2 (N3917, N3895, N2321);
or OR2 (N3918, N3909, N499);
nand NAND4 (N3919, N3916, N3246, N1202, N2644);
nand NAND4 (N3920, N3911, N2775, N3248, N2232);
xor XOR2 (N3921, N3918, N2888);
and AND2 (N3922, N3899, N3047);
not NOT1 (N3923, N3922);
nor NOR3 (N3924, N3920, N2182, N1117);
or OR4 (N3925, N3919, N3509, N1974, N2109);
xor XOR2 (N3926, N3923, N920);
nor NOR4 (N3927, N3925, N151, N2416, N3248);
not NOT1 (N3928, N3924);
not NOT1 (N3929, N3927);
and AND3 (N3930, N3912, N2605, N1998);
not NOT1 (N3931, N3930);
nor NOR4 (N3932, N3913, N2903, N3886, N3096);
nor NOR2 (N3933, N3929, N2024);
nand NAND2 (N3934, N3910, N2507);
not NOT1 (N3935, N3915);
or OR3 (N3936, N3928, N802, N2691);
not NOT1 (N3937, N3926);
nor NOR4 (N3938, N3935, N3060, N309, N2148);
xor XOR2 (N3939, N3936, N2402);
xor XOR2 (N3940, N3898, N1530);
and AND3 (N3941, N3938, N2521, N264);
and AND3 (N3942, N3932, N2954, N940);
nor NOR4 (N3943, N3939, N726, N3095, N3289);
nand NAND4 (N3944, N3917, N1373, N1417, N3181);
xor XOR2 (N3945, N3940, N2200);
or OR4 (N3946, N3944, N2440, N739, N2444);
and AND2 (N3947, N3945, N592);
buf BUF1 (N3948, N3946);
nor NOR2 (N3949, N3948, N619);
not NOT1 (N3950, N3947);
nor NOR4 (N3951, N3943, N2052, N56, N290);
nor NOR3 (N3952, N3937, N1424, N3734);
and AND3 (N3953, N3949, N3305, N3410);
buf BUF1 (N3954, N3953);
and AND3 (N3955, N3942, N1324, N1398);
nor NOR3 (N3956, N3950, N3588, N873);
nand NAND3 (N3957, N3933, N855, N3329);
buf BUF1 (N3958, N3956);
nand NAND4 (N3959, N3957, N3786, N3497, N1052);
nand NAND2 (N3960, N3934, N3848);
and AND2 (N3961, N3952, N900);
nand NAND3 (N3962, N3955, N446, N3241);
not NOT1 (N3963, N3941);
buf BUF1 (N3964, N3959);
or OR3 (N3965, N3963, N1717, N3677);
or OR3 (N3966, N3962, N193, N1555);
buf BUF1 (N3967, N3960);
or OR4 (N3968, N3931, N2973, N2872, N1963);
nor NOR2 (N3969, N3954, N1968);
and AND4 (N3970, N3969, N3480, N3780, N1948);
buf BUF1 (N3971, N3951);
and AND2 (N3972, N3967, N1447);
buf BUF1 (N3973, N3972);
xor XOR2 (N3974, N3961, N127);
xor XOR2 (N3975, N3968, N1998);
xor XOR2 (N3976, N3965, N611);
nor NOR4 (N3977, N3921, N3371, N1796, N12);
and AND4 (N3978, N3977, N3382, N2368, N565);
nor NOR4 (N3979, N3973, N815, N1509, N3123);
xor XOR2 (N3980, N3971, N1733);
not NOT1 (N3981, N3958);
buf BUF1 (N3982, N3980);
nand NAND2 (N3983, N3976, N2414);
or OR4 (N3984, N3978, N2374, N2023, N3981);
xor XOR2 (N3985, N26, N2237);
nor NOR4 (N3986, N3982, N749, N276, N802);
and AND2 (N3987, N3984, N3796);
xor XOR2 (N3988, N3985, N1834);
buf BUF1 (N3989, N3979);
buf BUF1 (N3990, N3964);
and AND2 (N3991, N3983, N1290);
not NOT1 (N3992, N3987);
and AND3 (N3993, N3988, N2834, N3961);
or OR3 (N3994, N3966, N2318, N1235);
and AND3 (N3995, N3986, N2716, N3034);
nand NAND3 (N3996, N3975, N1169, N135);
buf BUF1 (N3997, N3996);
not NOT1 (N3998, N3995);
buf BUF1 (N3999, N3997);
nand NAND3 (N4000, N3990, N476, N3183);
not NOT1 (N4001, N3974);
buf BUF1 (N4002, N3970);
nor NOR2 (N4003, N3991, N2097);
nor NOR4 (N4004, N3998, N3191, N204, N3743);
or OR2 (N4005, N3992, N2092);
or OR4 (N4006, N4002, N2329, N3891, N1529);
not NOT1 (N4007, N3994);
xor XOR2 (N4008, N4001, N3339);
not NOT1 (N4009, N4006);
or OR3 (N4010, N4008, N2772, N1578);
or OR2 (N4011, N3999, N3697);
nand NAND3 (N4012, N4005, N3482, N2929);
not NOT1 (N4013, N4009);
nor NOR2 (N4014, N4000, N2504);
and AND4 (N4015, N3993, N909, N3822, N2980);
and AND3 (N4016, N4014, N2388, N1124);
nor NOR3 (N4017, N4004, N140, N973);
or OR4 (N4018, N4003, N1077, N2764, N2997);
nand NAND2 (N4019, N4017, N2911);
or OR2 (N4020, N4018, N2748);
xor XOR2 (N4021, N4020, N1321);
xor XOR2 (N4022, N4010, N1548);
and AND4 (N4023, N4016, N2849, N649, N646);
and AND3 (N4024, N3989, N1622, N530);
and AND3 (N4025, N4015, N3970, N2592);
xor XOR2 (N4026, N4007, N3192);
or OR4 (N4027, N4024, N2018, N1468, N1214);
nand NAND2 (N4028, N4012, N3348);
not NOT1 (N4029, N4021);
xor XOR2 (N4030, N4026, N3474);
buf BUF1 (N4031, N4013);
xor XOR2 (N4032, N4028, N2768);
or OR4 (N4033, N4025, N729, N1224, N3750);
or OR2 (N4034, N4032, N3869);
xor XOR2 (N4035, N4027, N2456);
nand NAND4 (N4036, N4022, N852, N2783, N457);
nand NAND4 (N4037, N4033, N3337, N2013, N2384);
not NOT1 (N4038, N4029);
xor XOR2 (N4039, N4038, N1393);
xor XOR2 (N4040, N4031, N1084);
or OR2 (N4041, N4019, N31);
or OR2 (N4042, N4035, N298);
buf BUF1 (N4043, N4040);
buf BUF1 (N4044, N4042);
not NOT1 (N4045, N4039);
nor NOR2 (N4046, N4036, N3186);
buf BUF1 (N4047, N4023);
or OR3 (N4048, N4045, N3543, N3943);
not NOT1 (N4049, N4046);
not NOT1 (N4050, N4048);
or OR2 (N4051, N4050, N2667);
or OR2 (N4052, N4037, N52);
nor NOR4 (N4053, N4011, N548, N182, N677);
xor XOR2 (N4054, N4047, N3631);
and AND4 (N4055, N4030, N3323, N2003, N2974);
and AND2 (N4056, N4055, N2009);
and AND3 (N4057, N4043, N2368, N2223);
buf BUF1 (N4058, N4052);
or OR2 (N4059, N4041, N394);
xor XOR2 (N4060, N4057, N1808);
xor XOR2 (N4061, N4049, N708);
or OR3 (N4062, N4059, N122, N693);
not NOT1 (N4063, N4062);
nand NAND4 (N4064, N4053, N1274, N1201, N1111);
not NOT1 (N4065, N4058);
nand NAND4 (N4066, N4054, N994, N1234, N3382);
not NOT1 (N4067, N4060);
or OR4 (N4068, N4066, N3322, N2345, N1542);
xor XOR2 (N4069, N4061, N2184);
nor NOR3 (N4070, N4064, N860, N1358);
nor NOR2 (N4071, N4065, N1619);
and AND2 (N4072, N4063, N54);
or OR2 (N4073, N4071, N3220);
and AND2 (N4074, N4073, N3482);
and AND2 (N4075, N4068, N992);
buf BUF1 (N4076, N4034);
not NOT1 (N4077, N4056);
nand NAND3 (N4078, N4076, N807, N2392);
or OR2 (N4079, N4051, N2523);
nor NOR2 (N4080, N4070, N567);
buf BUF1 (N4081, N4067);
buf BUF1 (N4082, N4069);
nand NAND2 (N4083, N4072, N1658);
and AND2 (N4084, N4074, N1250);
xor XOR2 (N4085, N4075, N3202);
not NOT1 (N4086, N4081);
not NOT1 (N4087, N4077);
not NOT1 (N4088, N4087);
or OR2 (N4089, N4082, N2023);
not NOT1 (N4090, N4086);
buf BUF1 (N4091, N4090);
nand NAND2 (N4092, N4084, N1644);
not NOT1 (N4093, N4083);
and AND4 (N4094, N4080, N368, N777, N1486);
and AND4 (N4095, N4091, N3370, N1690, N533);
and AND3 (N4096, N4078, N3812, N230);
nand NAND3 (N4097, N4079, N3610, N1525);
nor NOR2 (N4098, N4094, N3433);
xor XOR2 (N4099, N4095, N1810);
nor NOR4 (N4100, N4098, N867, N902, N2900);
xor XOR2 (N4101, N4088, N2123);
not NOT1 (N4102, N4089);
and AND3 (N4103, N4096, N2788, N1427);
buf BUF1 (N4104, N4100);
and AND4 (N4105, N4092, N168, N441, N3521);
not NOT1 (N4106, N4102);
xor XOR2 (N4107, N4104, N2192);
nor NOR2 (N4108, N4106, N1860);
nor NOR2 (N4109, N4099, N4033);
and AND3 (N4110, N4097, N3670, N2835);
not NOT1 (N4111, N4107);
and AND4 (N4112, N4044, N434, N3912, N2306);
and AND2 (N4113, N4085, N281);
nor NOR4 (N4114, N4112, N2486, N2763, N2278);
buf BUF1 (N4115, N4105);
xor XOR2 (N4116, N4103, N606);
buf BUF1 (N4117, N4109);
and AND4 (N4118, N4116, N191, N3412, N1362);
not NOT1 (N4119, N4115);
xor XOR2 (N4120, N4110, N388);
nand NAND2 (N4121, N4108, N844);
xor XOR2 (N4122, N4111, N3900);
and AND4 (N4123, N4093, N3058, N1671, N965);
or OR3 (N4124, N4122, N423, N515);
and AND3 (N4125, N4101, N2422, N239);
buf BUF1 (N4126, N4125);
buf BUF1 (N4127, N4120);
and AND3 (N4128, N4124, N3120, N4102);
or OR2 (N4129, N4114, N773);
nor NOR4 (N4130, N4118, N425, N2669, N905);
xor XOR2 (N4131, N4128, N1964);
or OR2 (N4132, N4121, N482);
or OR2 (N4133, N4132, N3915);
or OR4 (N4134, N4127, N1045, N3214, N1231);
and AND4 (N4135, N4119, N3169, N4084, N1083);
and AND4 (N4136, N4134, N2647, N3664, N229);
buf BUF1 (N4137, N4136);
buf BUF1 (N4138, N4133);
and AND2 (N4139, N4126, N3199);
nand NAND3 (N4140, N4130, N3925, N2998);
nand NAND2 (N4141, N4123, N753);
nor NOR2 (N4142, N4131, N1029);
or OR3 (N4143, N4113, N3098, N996);
nand NAND3 (N4144, N4135, N4085, N3662);
not NOT1 (N4145, N4129);
and AND4 (N4146, N4140, N956, N2937, N2180);
or OR2 (N4147, N4141, N1543);
nor NOR2 (N4148, N4142, N3761);
not NOT1 (N4149, N4138);
xor XOR2 (N4150, N4117, N925);
buf BUF1 (N4151, N4146);
xor XOR2 (N4152, N4143, N1558);
or OR4 (N4153, N4148, N3568, N486, N82);
nor NOR2 (N4154, N4149, N4033);
nand NAND3 (N4155, N4152, N2972, N382);
nor NOR3 (N4156, N4145, N3317, N1254);
and AND4 (N4157, N4154, N3153, N2832, N2704);
nand NAND2 (N4158, N4151, N1309);
buf BUF1 (N4159, N4157);
or OR2 (N4160, N4158, N1990);
xor XOR2 (N4161, N4160, N593);
nor NOR2 (N4162, N4153, N3147);
or OR4 (N4163, N4150, N369, N604, N3877);
buf BUF1 (N4164, N4163);
and AND2 (N4165, N4162, N3737);
nand NAND3 (N4166, N4165, N1905, N1253);
not NOT1 (N4167, N4155);
buf BUF1 (N4168, N4164);
nand NAND4 (N4169, N4167, N2979, N3, N3046);
buf BUF1 (N4170, N4168);
buf BUF1 (N4171, N4159);
not NOT1 (N4172, N4171);
nand NAND4 (N4173, N4170, N3948, N2643, N3099);
not NOT1 (N4174, N4147);
and AND4 (N4175, N4144, N344, N2395, N1398);
xor XOR2 (N4176, N4137, N102);
and AND4 (N4177, N4176, N1167, N3854, N2871);
and AND4 (N4178, N4174, N3163, N2001, N890);
buf BUF1 (N4179, N4172);
not NOT1 (N4180, N4166);
buf BUF1 (N4181, N4161);
or OR2 (N4182, N4178, N1085);
nand NAND2 (N4183, N4177, N1661);
or OR3 (N4184, N4139, N3241, N1562);
not NOT1 (N4185, N4180);
or OR4 (N4186, N4184, N1899, N536, N1923);
nor NOR2 (N4187, N4186, N4159);
nand NAND4 (N4188, N4156, N4099, N1679, N2414);
and AND2 (N4189, N4179, N2425);
xor XOR2 (N4190, N4181, N2752);
xor XOR2 (N4191, N4188, N4143);
buf BUF1 (N4192, N4190);
xor XOR2 (N4193, N4173, N835);
xor XOR2 (N4194, N4183, N147);
nand NAND4 (N4195, N4187, N259, N2141, N2908);
buf BUF1 (N4196, N4194);
buf BUF1 (N4197, N4193);
xor XOR2 (N4198, N4169, N4060);
nor NOR4 (N4199, N4197, N2446, N1600, N431);
buf BUF1 (N4200, N4196);
xor XOR2 (N4201, N4189, N1962);
not NOT1 (N4202, N4199);
nor NOR4 (N4203, N4201, N484, N1501, N772);
xor XOR2 (N4204, N4182, N3572);
nand NAND2 (N4205, N4200, N580);
nor NOR2 (N4206, N4198, N2814);
or OR3 (N4207, N4203, N1463, N2873);
nand NAND3 (N4208, N4175, N3755, N3730);
nand NAND2 (N4209, N4195, N2969);
xor XOR2 (N4210, N4191, N731);
xor XOR2 (N4211, N4206, N932);
nand NAND3 (N4212, N4211, N184, N2797);
nand NAND3 (N4213, N4202, N1554, N386);
or OR2 (N4214, N4185, N3881);
xor XOR2 (N4215, N4214, N894);
buf BUF1 (N4216, N4207);
or OR2 (N4217, N4209, N2505);
or OR3 (N4218, N4216, N2354, N2300);
xor XOR2 (N4219, N4218, N1070);
not NOT1 (N4220, N4205);
nand NAND4 (N4221, N4212, N3727, N1590, N2448);
buf BUF1 (N4222, N4215);
not NOT1 (N4223, N4210);
xor XOR2 (N4224, N4223, N1512);
and AND2 (N4225, N4204, N3154);
and AND2 (N4226, N4217, N230);
nor NOR2 (N4227, N4222, N641);
and AND3 (N4228, N4208, N3137, N3667);
nand NAND2 (N4229, N4219, N3020);
nor NOR2 (N4230, N4224, N2108);
nand NAND3 (N4231, N4192, N2482, N2375);
not NOT1 (N4232, N4230);
and AND3 (N4233, N4225, N1906, N1581);
buf BUF1 (N4234, N4233);
nor NOR3 (N4235, N4221, N1579, N282);
xor XOR2 (N4236, N4235, N3616);
nor NOR4 (N4237, N4213, N2031, N1553, N3842);
xor XOR2 (N4238, N4231, N138);
nand NAND3 (N4239, N4227, N1081, N1027);
and AND4 (N4240, N4236, N2072, N2914, N3214);
not NOT1 (N4241, N4232);
or OR3 (N4242, N4237, N382, N1501);
and AND2 (N4243, N4229, N1933);
nor NOR3 (N4244, N4240, N1839, N1855);
buf BUF1 (N4245, N4243);
or OR2 (N4246, N4228, N1092);
not NOT1 (N4247, N4234);
xor XOR2 (N4248, N4247, N927);
xor XOR2 (N4249, N4238, N2630);
xor XOR2 (N4250, N4249, N1621);
nor NOR3 (N4251, N4242, N3046, N556);
nor NOR4 (N4252, N4250, N450, N2268, N80);
or OR3 (N4253, N4244, N2010, N1913);
and AND4 (N4254, N4220, N101, N3894, N1213);
nand NAND3 (N4255, N4252, N172, N1473);
nor NOR3 (N4256, N4239, N809, N3536);
buf BUF1 (N4257, N4241);
buf BUF1 (N4258, N4246);
or OR3 (N4259, N4245, N923, N2398);
or OR2 (N4260, N4254, N570);
nand NAND3 (N4261, N4258, N1652, N505);
nor NOR4 (N4262, N4260, N1107, N2682, N1690);
xor XOR2 (N4263, N4248, N2154);
and AND4 (N4264, N4257, N1688, N949, N1359);
or OR4 (N4265, N4264, N4025, N2826, N112);
nand NAND4 (N4266, N4256, N3886, N1246, N534);
nor NOR2 (N4267, N4259, N4208);
nand NAND2 (N4268, N4261, N2297);
nand NAND4 (N4269, N4253, N3893, N2166, N481);
not NOT1 (N4270, N4267);
not NOT1 (N4271, N4255);
or OR2 (N4272, N4263, N2830);
or OR2 (N4273, N4266, N2794);
not NOT1 (N4274, N4270);
nand NAND4 (N4275, N4269, N4183, N1094, N275);
not NOT1 (N4276, N4265);
or OR2 (N4277, N4274, N1497);
and AND3 (N4278, N4273, N509, N3841);
xor XOR2 (N4279, N4277, N872);
buf BUF1 (N4280, N4226);
and AND2 (N4281, N4268, N2411);
and AND3 (N4282, N4280, N3248, N2601);
nor NOR4 (N4283, N4278, N2296, N1529, N713);
buf BUF1 (N4284, N4282);
nand NAND4 (N4285, N4251, N2860, N2690, N2203);
buf BUF1 (N4286, N4284);
nor NOR2 (N4287, N4262, N38);
nor NOR3 (N4288, N4283, N3332, N2395);
nand NAND4 (N4289, N4272, N3643, N2477, N3817);
buf BUF1 (N4290, N4275);
xor XOR2 (N4291, N4287, N11);
buf BUF1 (N4292, N4271);
not NOT1 (N4293, N4289);
nor NOR3 (N4294, N4285, N1590, N3119);
nor NOR4 (N4295, N4290, N2798, N2556, N1153);
nor NOR4 (N4296, N4294, N2724, N268, N4066);
nand NAND4 (N4297, N4286, N3596, N1716, N1766);
not NOT1 (N4298, N4288);
buf BUF1 (N4299, N4276);
not NOT1 (N4300, N4291);
nor NOR4 (N4301, N4298, N3949, N645, N1222);
nand NAND4 (N4302, N4300, N2856, N1443, N4069);
and AND3 (N4303, N4297, N93, N426);
and AND4 (N4304, N4295, N4231, N597, N3454);
xor XOR2 (N4305, N4279, N1124);
xor XOR2 (N4306, N4292, N1670);
not NOT1 (N4307, N4303);
buf BUF1 (N4308, N4293);
buf BUF1 (N4309, N4307);
nand NAND2 (N4310, N4305, N356);
nor NOR4 (N4311, N4296, N3513, N1819, N2496);
nor NOR4 (N4312, N4310, N1515, N2970, N2861);
nand NAND3 (N4313, N4302, N973, N139);
xor XOR2 (N4314, N4308, N2894);
not NOT1 (N4315, N4304);
nand NAND4 (N4316, N4311, N1574, N2746, N710);
xor XOR2 (N4317, N4316, N3710);
and AND3 (N4318, N4314, N513, N1039);
and AND4 (N4319, N4317, N2800, N4010, N1036);
nand NAND3 (N4320, N4306, N2441, N3452);
xor XOR2 (N4321, N4312, N2923);
and AND4 (N4322, N4301, N2268, N3374, N4185);
xor XOR2 (N4323, N4321, N3654);
or OR2 (N4324, N4309, N3754);
xor XOR2 (N4325, N4319, N1360);
buf BUF1 (N4326, N4322);
nand NAND2 (N4327, N4281, N3984);
xor XOR2 (N4328, N4326, N415);
xor XOR2 (N4329, N4299, N1578);
buf BUF1 (N4330, N4324);
buf BUF1 (N4331, N4330);
and AND3 (N4332, N4327, N1931, N2670);
xor XOR2 (N4333, N4332, N2093);
and AND4 (N4334, N4331, N3214, N2212, N4274);
not NOT1 (N4335, N4334);
not NOT1 (N4336, N4313);
not NOT1 (N4337, N4323);
and AND3 (N4338, N4337, N675, N3038);
nor NOR3 (N4339, N4315, N3070, N4118);
nor NOR3 (N4340, N4320, N2756, N4301);
xor XOR2 (N4341, N4333, N3094);
not NOT1 (N4342, N4340);
and AND4 (N4343, N4318, N3538, N745, N1253);
and AND4 (N4344, N4335, N3683, N3751, N2579);
buf BUF1 (N4345, N4336);
nand NAND4 (N4346, N4344, N1257, N554, N2515);
nand NAND3 (N4347, N4328, N35, N259);
or OR3 (N4348, N4325, N1067, N1597);
nor NOR3 (N4349, N4346, N2349, N2500);
xor XOR2 (N4350, N4349, N571);
not NOT1 (N4351, N4345);
xor XOR2 (N4352, N4350, N2221);
nor NOR3 (N4353, N4352, N3806, N477);
not NOT1 (N4354, N4353);
buf BUF1 (N4355, N4348);
xor XOR2 (N4356, N4341, N2949);
nand NAND2 (N4357, N4329, N810);
nand NAND2 (N4358, N4339, N299);
buf BUF1 (N4359, N4342);
nand NAND3 (N4360, N4354, N2811, N3910);
nor NOR3 (N4361, N4358, N4135, N1057);
nor NOR3 (N4362, N4355, N2447, N2493);
or OR3 (N4363, N4357, N3407, N3071);
xor XOR2 (N4364, N4359, N27);
nor NOR2 (N4365, N4363, N4028);
and AND4 (N4366, N4364, N1834, N2412, N3815);
not NOT1 (N4367, N4366);
or OR3 (N4368, N4347, N263, N1602);
nand NAND2 (N4369, N4338, N271);
and AND3 (N4370, N4369, N1605, N3227);
xor XOR2 (N4371, N4370, N2345);
nor NOR2 (N4372, N4367, N702);
xor XOR2 (N4373, N4365, N2861);
nand NAND4 (N4374, N4368, N1506, N3539, N2408);
buf BUF1 (N4375, N4356);
xor XOR2 (N4376, N4362, N553);
and AND3 (N4377, N4360, N2042, N487);
and AND2 (N4378, N4376, N3989);
nand NAND2 (N4379, N4378, N1257);
nand NAND3 (N4380, N4379, N4249, N4002);
buf BUF1 (N4381, N4371);
nor NOR3 (N4382, N4372, N2808, N278);
xor XOR2 (N4383, N4343, N1968);
and AND4 (N4384, N4351, N4038, N3328, N1286);
nor NOR3 (N4385, N4383, N1426, N2131);
buf BUF1 (N4386, N4385);
xor XOR2 (N4387, N4375, N1821);
xor XOR2 (N4388, N4373, N3109);
or OR3 (N4389, N4380, N1837, N772);
and AND4 (N4390, N4377, N3261, N3722, N2434);
or OR4 (N4391, N4384, N1930, N2529, N3623);
or OR2 (N4392, N4387, N4159);
not NOT1 (N4393, N4388);
or OR2 (N4394, N4382, N4334);
xor XOR2 (N4395, N4392, N2364);
nor NOR3 (N4396, N4389, N3971, N81);
buf BUF1 (N4397, N4395);
xor XOR2 (N4398, N4396, N2736);
and AND4 (N4399, N4391, N1888, N1598, N2620);
nor NOR2 (N4400, N4390, N2049);
xor XOR2 (N4401, N4399, N580);
and AND2 (N4402, N4386, N2192);
and AND2 (N4403, N4401, N121);
not NOT1 (N4404, N4381);
or OR3 (N4405, N4404, N3786, N4180);
and AND4 (N4406, N4394, N2116, N3500, N2235);
xor XOR2 (N4407, N4403, N2253);
and AND3 (N4408, N4407, N1597, N2681);
not NOT1 (N4409, N4406);
nor NOR3 (N4410, N4361, N2344, N4345);
nor NOR4 (N4411, N4393, N2631, N1520, N3169);
or OR4 (N4412, N4408, N4286, N2133, N2016);
buf BUF1 (N4413, N4400);
or OR4 (N4414, N4374, N1941, N1922, N2354);
nor NOR2 (N4415, N4398, N1270);
nand NAND3 (N4416, N4413, N4282, N3105);
nor NOR4 (N4417, N4405, N3443, N961, N781);
nor NOR4 (N4418, N4415, N974, N1698, N670);
buf BUF1 (N4419, N4409);
and AND2 (N4420, N4418, N3961);
nand NAND2 (N4421, N4397, N1377);
or OR2 (N4422, N4412, N2570);
nand NAND4 (N4423, N4410, N696, N1057, N3023);
nand NAND3 (N4424, N4419, N2540, N2783);
not NOT1 (N4425, N4414);
nand NAND2 (N4426, N4416, N4243);
buf BUF1 (N4427, N4423);
xor XOR2 (N4428, N4424, N3351);
nor NOR3 (N4429, N4420, N1181, N3808);
nor NOR4 (N4430, N4421, N4000, N4345, N2110);
not NOT1 (N4431, N4427);
or OR4 (N4432, N4429, N3968, N3700, N4186);
not NOT1 (N4433, N4417);
xor XOR2 (N4434, N4411, N2164);
or OR2 (N4435, N4428, N135);
nor NOR2 (N4436, N4426, N3722);
not NOT1 (N4437, N4402);
buf BUF1 (N4438, N4435);
xor XOR2 (N4439, N4425, N2919);
xor XOR2 (N4440, N4439, N465);
nand NAND4 (N4441, N4422, N2373, N2786, N697);
or OR2 (N4442, N4430, N3713);
buf BUF1 (N4443, N4432);
xor XOR2 (N4444, N4441, N838);
or OR2 (N4445, N4438, N2713);
and AND2 (N4446, N4442, N3665);
not NOT1 (N4447, N4434);
nand NAND2 (N4448, N4446, N824);
or OR4 (N4449, N4448, N592, N2627, N2);
nor NOR4 (N4450, N4436, N595, N1983, N2084);
nor NOR3 (N4451, N4450, N163, N1977);
and AND2 (N4452, N4437, N3378);
nor NOR2 (N4453, N4433, N2524);
and AND3 (N4454, N4449, N3856, N3153);
buf BUF1 (N4455, N4445);
not NOT1 (N4456, N4454);
not NOT1 (N4457, N4455);
nor NOR4 (N4458, N4453, N3541, N3912, N2155);
not NOT1 (N4459, N4457);
xor XOR2 (N4460, N4451, N854);
xor XOR2 (N4461, N4452, N12);
not NOT1 (N4462, N4444);
nor NOR2 (N4463, N4460, N356);
nand NAND2 (N4464, N4431, N2013);
xor XOR2 (N4465, N4464, N707);
xor XOR2 (N4466, N4447, N3095);
not NOT1 (N4467, N4443);
or OR4 (N4468, N4440, N2230, N67, N2548);
xor XOR2 (N4469, N4462, N332);
buf BUF1 (N4470, N4467);
nand NAND4 (N4471, N4465, N2934, N2794, N1212);
nor NOR3 (N4472, N4471, N3457, N1855);
xor XOR2 (N4473, N4463, N4142);
buf BUF1 (N4474, N4470);
or OR2 (N4475, N4461, N2030);
nor NOR3 (N4476, N4456, N2433, N1018);
buf BUF1 (N4477, N4473);
or OR3 (N4478, N4474, N2247, N4236);
buf BUF1 (N4479, N4468);
or OR4 (N4480, N4476, N2933, N163, N3789);
xor XOR2 (N4481, N4480, N4117);
buf BUF1 (N4482, N4475);
xor XOR2 (N4483, N4459, N1293);
or OR3 (N4484, N4483, N1280, N1410);
buf BUF1 (N4485, N4481);
and AND2 (N4486, N4466, N2223);
and AND3 (N4487, N4486, N4373, N1778);
nor NOR4 (N4488, N4479, N2844, N384, N2911);
nor NOR4 (N4489, N4472, N2076, N4339, N1059);
or OR3 (N4490, N4482, N3464, N1612);
and AND2 (N4491, N4478, N2706);
nand NAND2 (N4492, N4491, N2757);
and AND3 (N4493, N4484, N4138, N1224);
nand NAND4 (N4494, N4490, N953, N1574, N994);
not NOT1 (N4495, N4487);
nor NOR3 (N4496, N4488, N3862, N543);
xor XOR2 (N4497, N4494, N823);
not NOT1 (N4498, N4497);
buf BUF1 (N4499, N4498);
and AND2 (N4500, N4496, N520);
nor NOR2 (N4501, N4500, N1821);
nor NOR2 (N4502, N4469, N2893);
nand NAND4 (N4503, N4495, N2852, N3543, N1855);
nor NOR3 (N4504, N4492, N2986, N2318);
and AND4 (N4505, N4502, N1401, N3993, N1915);
nor NOR2 (N4506, N4485, N1144);
nand NAND4 (N4507, N4506, N4166, N2834, N2981);
not NOT1 (N4508, N4504);
or OR3 (N4509, N4501, N2700, N3753);
buf BUF1 (N4510, N4509);
and AND2 (N4511, N4507, N1122);
xor XOR2 (N4512, N4489, N907);
not NOT1 (N4513, N4503);
xor XOR2 (N4514, N4508, N2678);
nand NAND4 (N4515, N4493, N3994, N1354, N1617);
and AND2 (N4516, N4499, N1181);
buf BUF1 (N4517, N4515);
nand NAND4 (N4518, N4477, N3037, N2220, N690);
nor NOR2 (N4519, N4514, N1611);
nor NOR3 (N4520, N4510, N3830, N413);
nor NOR2 (N4521, N4520, N695);
or OR3 (N4522, N4521, N3270, N2);
nand NAND3 (N4523, N4513, N533, N4432);
and AND4 (N4524, N4511, N2337, N3469, N306);
buf BUF1 (N4525, N4518);
nor NOR4 (N4526, N4524, N2831, N4145, N2953);
or OR2 (N4527, N4519, N2041);
xor XOR2 (N4528, N4526, N4113);
buf BUF1 (N4529, N4517);
buf BUF1 (N4530, N4522);
buf BUF1 (N4531, N4530);
nor NOR3 (N4532, N4531, N810, N3583);
xor XOR2 (N4533, N4532, N3380);
or OR3 (N4534, N4528, N305, N4015);
buf BUF1 (N4535, N4533);
not NOT1 (N4536, N4534);
xor XOR2 (N4537, N4512, N3464);
not NOT1 (N4538, N4527);
not NOT1 (N4539, N4516);
buf BUF1 (N4540, N4525);
not NOT1 (N4541, N4537);
nor NOR3 (N4542, N4523, N3992, N2126);
nor NOR4 (N4543, N4541, N4482, N3515, N317);
buf BUF1 (N4544, N4505);
or OR3 (N4545, N4538, N3881, N1313);
buf BUF1 (N4546, N4539);
or OR4 (N4547, N4544, N2286, N4518, N1791);
or OR4 (N4548, N4545, N2735, N1920, N1115);
nor NOR2 (N4549, N4548, N4263);
buf BUF1 (N4550, N4529);
nor NOR3 (N4551, N4547, N4157, N2060);
xor XOR2 (N4552, N4535, N2235);
not NOT1 (N4553, N4536);
not NOT1 (N4554, N4552);
not NOT1 (N4555, N4458);
or OR3 (N4556, N4550, N1835, N3241);
not NOT1 (N4557, N4549);
not NOT1 (N4558, N4543);
xor XOR2 (N4559, N4555, N3355);
nand NAND3 (N4560, N4554, N3616, N3866);
xor XOR2 (N4561, N4558, N849);
nand NAND4 (N4562, N4551, N3056, N2482, N799);
or OR3 (N4563, N4560, N510, N3149);
or OR2 (N4564, N4540, N1410);
or OR3 (N4565, N4559, N2374, N1857);
or OR4 (N4566, N4563, N1670, N3581, N3893);
not NOT1 (N4567, N4553);
buf BUF1 (N4568, N4561);
nor NOR4 (N4569, N4542, N2900, N1942, N3464);
xor XOR2 (N4570, N4564, N753);
and AND3 (N4571, N4568, N117, N3967);
xor XOR2 (N4572, N4571, N3747);
not NOT1 (N4573, N4567);
xor XOR2 (N4574, N4556, N3619);
buf BUF1 (N4575, N4562);
nor NOR4 (N4576, N4572, N2822, N517, N420);
and AND2 (N4577, N4574, N910);
nor NOR3 (N4578, N4575, N2612, N3107);
nand NAND3 (N4579, N4573, N2779, N4148);
not NOT1 (N4580, N4566);
nor NOR2 (N4581, N4570, N982);
not NOT1 (N4582, N4580);
xor XOR2 (N4583, N4569, N605);
and AND2 (N4584, N4565, N2914);
or OR3 (N4585, N4577, N1331, N3475);
and AND4 (N4586, N4581, N1763, N1906, N589);
xor XOR2 (N4587, N4586, N4137);
nor NOR2 (N4588, N4578, N2002);
xor XOR2 (N4589, N4584, N1049);
or OR4 (N4590, N4589, N4505, N2280, N1225);
buf BUF1 (N4591, N4590);
nand NAND2 (N4592, N4591, N4343);
or OR3 (N4593, N4582, N3336, N2909);
or OR4 (N4594, N4587, N2807, N3976, N3273);
not NOT1 (N4595, N4588);
not NOT1 (N4596, N4592);
xor XOR2 (N4597, N4585, N878);
and AND3 (N4598, N4597, N1305, N125);
nor NOR3 (N4599, N4579, N4153, N4401);
xor XOR2 (N4600, N4598, N2979);
xor XOR2 (N4601, N4593, N2560);
and AND2 (N4602, N4546, N3340);
buf BUF1 (N4603, N4583);
buf BUF1 (N4604, N4602);
xor XOR2 (N4605, N4596, N1663);
and AND3 (N4606, N4595, N960, N2344);
nand NAND3 (N4607, N4603, N3313, N1623);
buf BUF1 (N4608, N4576);
not NOT1 (N4609, N4601);
not NOT1 (N4610, N4608);
nor NOR2 (N4611, N4599, N669);
and AND2 (N4612, N4606, N407);
nor NOR2 (N4613, N4607, N3489);
or OR4 (N4614, N4613, N265, N2612, N4596);
and AND2 (N4615, N4557, N2870);
buf BUF1 (N4616, N4605);
nor NOR2 (N4617, N4615, N3405);
not NOT1 (N4618, N4611);
xor XOR2 (N4619, N4614, N1572);
nand NAND3 (N4620, N4610, N1870, N2943);
nand NAND4 (N4621, N4609, N865, N962, N1522);
buf BUF1 (N4622, N4616);
nand NAND3 (N4623, N4600, N3656, N4023);
nand NAND2 (N4624, N4620, N2979);
not NOT1 (N4625, N4618);
nor NOR3 (N4626, N4612, N2434, N2280);
xor XOR2 (N4627, N4604, N3573);
nand NAND4 (N4628, N4617, N2587, N1538, N944);
or OR4 (N4629, N4624, N3054, N1030, N3833);
xor XOR2 (N4630, N4625, N3306);
xor XOR2 (N4631, N4627, N1614);
not NOT1 (N4632, N4630);
not NOT1 (N4633, N4626);
and AND2 (N4634, N4628, N2528);
buf BUF1 (N4635, N4632);
buf BUF1 (N4636, N4623);
buf BUF1 (N4637, N4636);
not NOT1 (N4638, N4633);
nand NAND3 (N4639, N4619, N1392, N3542);
xor XOR2 (N4640, N4639, N1260);
or OR3 (N4641, N4629, N2757, N2530);
and AND4 (N4642, N4594, N2442, N1189, N1890);
buf BUF1 (N4643, N4640);
or OR3 (N4644, N4634, N3347, N270);
xor XOR2 (N4645, N4631, N2611);
buf BUF1 (N4646, N4642);
nor NOR4 (N4647, N4635, N3478, N664, N1397);
and AND4 (N4648, N4645, N1077, N2687, N213);
buf BUF1 (N4649, N4622);
not NOT1 (N4650, N4644);
and AND2 (N4651, N4650, N2904);
or OR3 (N4652, N4641, N4196, N1169);
not NOT1 (N4653, N4646);
and AND3 (N4654, N4653, N4540, N696);
buf BUF1 (N4655, N4647);
buf BUF1 (N4656, N4654);
or OR3 (N4657, N4649, N4346, N2022);
and AND3 (N4658, N4637, N1189, N3605);
or OR2 (N4659, N4648, N2983);
and AND3 (N4660, N4658, N1756, N1366);
xor XOR2 (N4661, N4652, N4429);
xor XOR2 (N4662, N4651, N1431);
or OR4 (N4663, N4662, N2778, N1648, N1149);
or OR2 (N4664, N4643, N4454);
nor NOR3 (N4665, N4655, N2080, N3449);
or OR4 (N4666, N4663, N1164, N39, N1524);
nand NAND2 (N4667, N4621, N1914);
xor XOR2 (N4668, N4664, N2716);
buf BUF1 (N4669, N4660);
nor NOR2 (N4670, N4669, N2595);
nor NOR2 (N4671, N4661, N3325);
and AND4 (N4672, N4665, N4311, N1738, N501);
or OR2 (N4673, N4667, N4557);
buf BUF1 (N4674, N4659);
nand NAND3 (N4675, N4670, N805, N162);
or OR3 (N4676, N4673, N240, N3899);
nor NOR2 (N4677, N4668, N2887);
nor NOR3 (N4678, N4674, N476, N1020);
or OR3 (N4679, N4677, N1417, N3531);
or OR3 (N4680, N4656, N4635, N4034);
xor XOR2 (N4681, N4638, N3589);
xor XOR2 (N4682, N4676, N4543);
not NOT1 (N4683, N4675);
nor NOR3 (N4684, N4683, N3944, N1445);
xor XOR2 (N4685, N4680, N2282);
not NOT1 (N4686, N4671);
buf BUF1 (N4687, N4682);
or OR2 (N4688, N4685, N4282);
or OR3 (N4689, N4678, N2274, N1064);
nor NOR3 (N4690, N4687, N2560, N3168);
or OR4 (N4691, N4690, N2682, N3783, N588);
xor XOR2 (N4692, N4686, N3596);
xor XOR2 (N4693, N4666, N904);
buf BUF1 (N4694, N4681);
buf BUF1 (N4695, N4679);
or OR2 (N4696, N4657, N1632);
nor NOR4 (N4697, N4691, N1683, N443, N2565);
buf BUF1 (N4698, N4684);
or OR4 (N4699, N4688, N1263, N2696, N2304);
nor NOR3 (N4700, N4696, N1310, N1140);
and AND4 (N4701, N4698, N3567, N3535, N1232);
nand NAND3 (N4702, N4701, N3651, N744);
not NOT1 (N4703, N4672);
nor NOR4 (N4704, N4693, N3964, N4173, N3955);
and AND3 (N4705, N4697, N4090, N3994);
not NOT1 (N4706, N4692);
and AND3 (N4707, N4706, N3315, N2721);
nand NAND3 (N4708, N4699, N2146, N576);
nand NAND3 (N4709, N4707, N3856, N298);
nor NOR3 (N4710, N4689, N4091, N2277);
nand NAND2 (N4711, N4695, N4495);
not NOT1 (N4712, N4700);
nand NAND3 (N4713, N4709, N2285, N3681);
buf BUF1 (N4714, N4712);
buf BUF1 (N4715, N4713);
or OR4 (N4716, N4708, N2022, N4510, N1854);
not NOT1 (N4717, N4702);
or OR4 (N4718, N4717, N3347, N1251, N4375);
buf BUF1 (N4719, N4718);
nand NAND3 (N4720, N4711, N1495, N393);
nor NOR2 (N4721, N4714, N2241);
and AND2 (N4722, N4705, N1476);
nor NOR2 (N4723, N4720, N1359);
nor NOR3 (N4724, N4694, N3375, N653);
nor NOR2 (N4725, N4704, N83);
buf BUF1 (N4726, N4719);
and AND2 (N4727, N4710, N630);
buf BUF1 (N4728, N4726);
buf BUF1 (N4729, N4716);
buf BUF1 (N4730, N4703);
not NOT1 (N4731, N4715);
nand NAND2 (N4732, N4729, N1773);
buf BUF1 (N4733, N4731);
nand NAND3 (N4734, N4723, N4461, N2649);
or OR4 (N4735, N4722, N2101, N163, N1319);
xor XOR2 (N4736, N4733, N2345);
nor NOR4 (N4737, N4725, N1852, N3631, N4714);
buf BUF1 (N4738, N4728);
xor XOR2 (N4739, N4737, N1214);
not NOT1 (N4740, N4736);
xor XOR2 (N4741, N4727, N3045);
and AND4 (N4742, N4734, N273, N2290, N683);
nor NOR2 (N4743, N4735, N206);
or OR4 (N4744, N4738, N3813, N4127, N3846);
and AND4 (N4745, N4742, N1070, N3169, N4120);
nand NAND2 (N4746, N4724, N2902);
not NOT1 (N4747, N4740);
xor XOR2 (N4748, N4743, N444);
xor XOR2 (N4749, N4721, N1068);
nor NOR4 (N4750, N4730, N267, N1207, N1896);
xor XOR2 (N4751, N4749, N410);
buf BUF1 (N4752, N4744);
or OR4 (N4753, N4752, N55, N3504, N1932);
nand NAND2 (N4754, N4751, N180);
or OR4 (N4755, N4732, N1779, N743, N4251);
nor NOR2 (N4756, N4747, N3054);
and AND2 (N4757, N4748, N3167);
or OR2 (N4758, N4753, N4097);
nor NOR2 (N4759, N4746, N4581);
and AND4 (N4760, N4750, N520, N1993, N318);
buf BUF1 (N4761, N4757);
buf BUF1 (N4762, N4739);
nor NOR4 (N4763, N4754, N2105, N3939, N2998);
nor NOR2 (N4764, N4745, N519);
or OR2 (N4765, N4762, N3391);
nor NOR2 (N4766, N4763, N4640);
or OR4 (N4767, N4741, N1682, N3084, N4157);
buf BUF1 (N4768, N4764);
nor NOR4 (N4769, N4765, N427, N2212, N3875);
not NOT1 (N4770, N4759);
xor XOR2 (N4771, N4760, N1389);
nor NOR2 (N4772, N4756, N2328);
xor XOR2 (N4773, N4766, N695);
xor XOR2 (N4774, N4769, N2668);
not NOT1 (N4775, N4767);
nand NAND2 (N4776, N4761, N124);
nand NAND4 (N4777, N4776, N2591, N2274, N43);
and AND2 (N4778, N4772, N2701);
nor NOR4 (N4779, N4768, N38, N3673, N2603);
or OR4 (N4780, N4771, N2918, N3983, N475);
nor NOR4 (N4781, N4780, N2189, N499, N3070);
nand NAND4 (N4782, N4775, N3488, N693, N4686);
buf BUF1 (N4783, N4777);
nor NOR2 (N4784, N4778, N875);
or OR2 (N4785, N4784, N4465);
not NOT1 (N4786, N4782);
or OR4 (N4787, N4770, N463, N3981, N4224);
and AND4 (N4788, N4787, N2796, N3471, N3439);
not NOT1 (N4789, N4773);
xor XOR2 (N4790, N4755, N471);
nor NOR2 (N4791, N4785, N1635);
nor NOR4 (N4792, N4758, N290, N3384, N2305);
and AND3 (N4793, N4774, N1272, N961);
nor NOR3 (N4794, N4789, N2619, N2936);
not NOT1 (N4795, N4781);
nor NOR2 (N4796, N4786, N2635);
buf BUF1 (N4797, N4793);
xor XOR2 (N4798, N4788, N3448);
or OR3 (N4799, N4791, N4660, N1079);
nor NOR4 (N4800, N4795, N3574, N4578, N4673);
or OR2 (N4801, N4779, N4132);
and AND2 (N4802, N4799, N3370);
and AND4 (N4803, N4794, N572, N1291, N2001);
not NOT1 (N4804, N4783);
or OR3 (N4805, N4797, N1204, N4685);
not NOT1 (N4806, N4804);
and AND2 (N4807, N4806, N3601);
nand NAND3 (N4808, N4801, N2681, N1732);
or OR2 (N4809, N4807, N1201);
buf BUF1 (N4810, N4798);
nor NOR2 (N4811, N4796, N4528);
not NOT1 (N4812, N4802);
nand NAND2 (N4813, N4803, N1122);
not NOT1 (N4814, N4811);
xor XOR2 (N4815, N4808, N4497);
or OR2 (N4816, N4812, N4260);
xor XOR2 (N4817, N4814, N2561);
and AND2 (N4818, N4813, N1701);
and AND2 (N4819, N4818, N3859);
or OR4 (N4820, N4819, N1530, N3459, N4342);
buf BUF1 (N4821, N4816);
buf BUF1 (N4822, N4809);
buf BUF1 (N4823, N4821);
and AND4 (N4824, N4810, N1108, N276, N1351);
or OR3 (N4825, N4822, N202, N3674);
or OR3 (N4826, N4824, N1126, N3640);
nand NAND3 (N4827, N4790, N1547, N3002);
nand NAND2 (N4828, N4823, N2773);
not NOT1 (N4829, N4817);
or OR2 (N4830, N4792, N1222);
and AND2 (N4831, N4805, N4565);
and AND2 (N4832, N4827, N2382);
nand NAND3 (N4833, N4832, N4579, N1170);
not NOT1 (N4834, N4800);
nand NAND2 (N4835, N4831, N2129);
and AND2 (N4836, N4815, N1250);
or OR4 (N4837, N4830, N2543, N955, N910);
or OR3 (N4838, N4835, N1264, N2795);
xor XOR2 (N4839, N4833, N1726);
and AND2 (N4840, N4826, N1006);
buf BUF1 (N4841, N4838);
buf BUF1 (N4842, N4839);
nor NOR3 (N4843, N4842, N2578, N1591);
not NOT1 (N4844, N4837);
nand NAND2 (N4845, N4829, N1296);
and AND2 (N4846, N4844, N4320);
xor XOR2 (N4847, N4828, N4452);
buf BUF1 (N4848, N4846);
buf BUF1 (N4849, N4847);
nor NOR2 (N4850, N4841, N2665);
nand NAND4 (N4851, N4834, N2276, N4644, N1783);
or OR3 (N4852, N4840, N3017, N3941);
not NOT1 (N4853, N4852);
not NOT1 (N4854, N4848);
nand NAND3 (N4855, N4845, N736, N3023);
buf BUF1 (N4856, N4853);
buf BUF1 (N4857, N4856);
not NOT1 (N4858, N4843);
nand NAND2 (N4859, N4857, N3199);
and AND4 (N4860, N4854, N3059, N1962, N2606);
not NOT1 (N4861, N4860);
buf BUF1 (N4862, N4849);
buf BUF1 (N4863, N4862);
not NOT1 (N4864, N4851);
or OR3 (N4865, N4861, N2929, N1386);
not NOT1 (N4866, N4864);
not NOT1 (N4867, N4865);
nand NAND3 (N4868, N4855, N388, N2824);
and AND3 (N4869, N4820, N796, N1958);
xor XOR2 (N4870, N4869, N4507);
buf BUF1 (N4871, N4836);
xor XOR2 (N4872, N4863, N3041);
not NOT1 (N4873, N4868);
nand NAND2 (N4874, N4859, N1413);
or OR3 (N4875, N4871, N2636, N3396);
xor XOR2 (N4876, N4870, N2955);
and AND3 (N4877, N4875, N1381, N773);
not NOT1 (N4878, N4850);
or OR4 (N4879, N4873, N217, N1056, N2564);
xor XOR2 (N4880, N4872, N2915);
not NOT1 (N4881, N4877);
and AND2 (N4882, N4878, N82);
and AND2 (N4883, N4879, N1553);
or OR4 (N4884, N4883, N1373, N313, N116);
not NOT1 (N4885, N4881);
nand NAND4 (N4886, N4885, N4342, N3756, N4085);
xor XOR2 (N4887, N4884, N4623);
or OR4 (N4888, N4880, N1124, N4505, N2817);
and AND2 (N4889, N4858, N820);
nand NAND3 (N4890, N4874, N414, N3188);
not NOT1 (N4891, N4825);
buf BUF1 (N4892, N4886);
nor NOR4 (N4893, N4887, N1404, N2900, N2657);
and AND2 (N4894, N4888, N1462);
xor XOR2 (N4895, N4892, N2795);
xor XOR2 (N4896, N4876, N3129);
nand NAND4 (N4897, N4867, N1784, N1613, N4074);
and AND2 (N4898, N4896, N471);
and AND3 (N4899, N4898, N3074, N3869);
not NOT1 (N4900, N4882);
xor XOR2 (N4901, N4893, N1876);
and AND2 (N4902, N4897, N2008);
not NOT1 (N4903, N4889);
nor NOR3 (N4904, N4903, N1401, N774);
nand NAND3 (N4905, N4901, N2614, N2739);
nor NOR3 (N4906, N4905, N2443, N1118);
nor NOR4 (N4907, N4906, N1770, N4453, N4570);
nand NAND3 (N4908, N4899, N647, N3796);
or OR4 (N4909, N4907, N4829, N3711, N3027);
nor NOR4 (N4910, N4902, N1659, N2208, N162);
xor XOR2 (N4911, N4890, N2351);
not NOT1 (N4912, N4904);
buf BUF1 (N4913, N4894);
or OR4 (N4914, N4866, N3074, N1809, N4164);
or OR3 (N4915, N4900, N1495, N2784);
or OR3 (N4916, N4895, N4813, N4402);
not NOT1 (N4917, N4914);
nor NOR2 (N4918, N4915, N3930);
buf BUF1 (N4919, N4891);
and AND4 (N4920, N4913, N1206, N4116, N1181);
or OR4 (N4921, N4911, N1329, N1954, N1192);
or OR2 (N4922, N4919, N4550);
buf BUF1 (N4923, N4910);
nor NOR3 (N4924, N4921, N1785, N1694);
buf BUF1 (N4925, N4916);
nor NOR2 (N4926, N4923, N1077);
and AND4 (N4927, N4924, N1489, N3388, N4652);
not NOT1 (N4928, N4927);
buf BUF1 (N4929, N4928);
and AND3 (N4930, N4918, N2945, N4190);
xor XOR2 (N4931, N4917, N1172);
or OR2 (N4932, N4931, N2193);
xor XOR2 (N4933, N4926, N3292);
and AND3 (N4934, N4909, N309, N4158);
not NOT1 (N4935, N4933);
nor NOR4 (N4936, N4908, N2942, N4262, N2413);
buf BUF1 (N4937, N4936);
and AND4 (N4938, N4930, N2166, N3232, N3046);
nor NOR4 (N4939, N4912, N3019, N396, N2985);
xor XOR2 (N4940, N4939, N1412);
nor NOR3 (N4941, N4932, N3491, N1884);
not NOT1 (N4942, N4929);
and AND2 (N4943, N4922, N3695);
nand NAND4 (N4944, N4943, N2189, N4511, N4211);
not NOT1 (N4945, N4935);
not NOT1 (N4946, N4934);
nand NAND3 (N4947, N4937, N1689, N2577);
nand NAND4 (N4948, N4925, N4835, N378, N1145);
not NOT1 (N4949, N4941);
xor XOR2 (N4950, N4942, N2308);
buf BUF1 (N4951, N4950);
nor NOR3 (N4952, N4938, N649, N3917);
or OR2 (N4953, N4951, N4598);
nor NOR3 (N4954, N4945, N3822, N4098);
nand NAND3 (N4955, N4954, N565, N4457);
not NOT1 (N4956, N4953);
or OR4 (N4957, N4948, N2491, N3667, N3591);
or OR4 (N4958, N4946, N803, N941, N3139);
not NOT1 (N4959, N4956);
and AND4 (N4960, N4958, N4370, N1333, N3670);
buf BUF1 (N4961, N4955);
nand NAND2 (N4962, N4959, N95);
not NOT1 (N4963, N4944);
or OR4 (N4964, N4963, N3620, N2107, N3889);
xor XOR2 (N4965, N4957, N2595);
nand NAND4 (N4966, N4964, N4537, N1678, N1448);
buf BUF1 (N4967, N4949);
nor NOR3 (N4968, N4966, N3934, N3442);
or OR4 (N4969, N4960, N4559, N2405, N1015);
xor XOR2 (N4970, N4969, N126);
buf BUF1 (N4971, N4947);
xor XOR2 (N4972, N4952, N3749);
buf BUF1 (N4973, N4968);
nand NAND3 (N4974, N4962, N3898, N1103);
or OR3 (N4975, N4940, N1257, N4711);
not NOT1 (N4976, N4965);
xor XOR2 (N4977, N4970, N1167);
not NOT1 (N4978, N4973);
and AND4 (N4979, N4977, N258, N3065, N2441);
not NOT1 (N4980, N4961);
xor XOR2 (N4981, N4980, N3453);
nor NOR4 (N4982, N4979, N3372, N2794, N2991);
xor XOR2 (N4983, N4976, N703);
not NOT1 (N4984, N4972);
buf BUF1 (N4985, N4984);
not NOT1 (N4986, N4983);
nand NAND3 (N4987, N4978, N2891, N4084);
not NOT1 (N4988, N4986);
nand NAND4 (N4989, N4982, N1178, N2137, N1933);
not NOT1 (N4990, N4974);
and AND4 (N4991, N4981, N2940, N191, N1786);
nor NOR3 (N4992, N4988, N1292, N1697);
buf BUF1 (N4993, N4985);
xor XOR2 (N4994, N4987, N1182);
xor XOR2 (N4995, N4992, N4719);
and AND3 (N4996, N4975, N2934, N3682);
or OR2 (N4997, N4994, N4542);
nand NAND4 (N4998, N4920, N4467, N3315, N3000);
nand NAND4 (N4999, N4990, N3484, N1833, N175);
nor NOR4 (N5000, N4996, N2226, N27, N1495);
or OR4 (N5001, N4971, N2399, N3979, N3053);
nand NAND2 (N5002, N4991, N2885);
nand NAND4 (N5003, N5001, N2711, N826, N2558);
nand NAND2 (N5004, N4967, N574);
or OR4 (N5005, N4995, N1888, N2486, N1717);
nor NOR3 (N5006, N5003, N3471, N219);
not NOT1 (N5007, N4999);
not NOT1 (N5008, N5002);
not NOT1 (N5009, N5008);
or OR4 (N5010, N5009, N4720, N3614, N3469);
nand NAND4 (N5011, N4998, N281, N577, N4294);
not NOT1 (N5012, N5005);
not NOT1 (N5013, N5006);
or OR4 (N5014, N5012, N3273, N2803, N3849);
nand NAND2 (N5015, N4989, N680);
not NOT1 (N5016, N5015);
and AND3 (N5017, N5010, N2692, N1237);
not NOT1 (N5018, N5017);
and AND2 (N5019, N5000, N2558);
nor NOR3 (N5020, N5004, N1073, N1113);
not NOT1 (N5021, N4997);
and AND4 (N5022, N5013, N4147, N3239, N2283);
nand NAND2 (N5023, N5022, N4815);
buf BUF1 (N5024, N5020);
nor NOR3 (N5025, N4993, N1272, N4282);
nor NOR2 (N5026, N5007, N1724);
not NOT1 (N5027, N5021);
nor NOR2 (N5028, N5016, N1595);
nand NAND3 (N5029, N5014, N3768, N2293);
xor XOR2 (N5030, N5019, N4497);
buf BUF1 (N5031, N5026);
buf BUF1 (N5032, N5023);
xor XOR2 (N5033, N5030, N1279);
and AND3 (N5034, N5032, N406, N2206);
and AND2 (N5035, N5011, N3908);
nor NOR2 (N5036, N5031, N336);
not NOT1 (N5037, N5036);
xor XOR2 (N5038, N5025, N3995);
xor XOR2 (N5039, N5038, N1102);
xor XOR2 (N5040, N5018, N3674);
and AND3 (N5041, N5027, N662, N1901);
nor NOR2 (N5042, N5034, N3108);
nor NOR2 (N5043, N5042, N1974);
not NOT1 (N5044, N5040);
nand NAND4 (N5045, N5044, N288, N3587, N3553);
xor XOR2 (N5046, N5033, N2245);
xor XOR2 (N5047, N5024, N1778);
buf BUF1 (N5048, N5043);
not NOT1 (N5049, N5029);
xor XOR2 (N5050, N5048, N500);
buf BUF1 (N5051, N5047);
buf BUF1 (N5052, N5050);
nor NOR3 (N5053, N5051, N3627, N1666);
xor XOR2 (N5054, N5028, N4031);
xor XOR2 (N5055, N5035, N2054);
buf BUF1 (N5056, N5045);
or OR4 (N5057, N5054, N4571, N33, N4925);
xor XOR2 (N5058, N5049, N599);
nor NOR3 (N5059, N5056, N3117, N1155);
and AND2 (N5060, N5041, N3233);
nand NAND4 (N5061, N5052, N4986, N886, N2939);
buf BUF1 (N5062, N5061);
and AND3 (N5063, N5057, N3411, N3124);
nand NAND3 (N5064, N5039, N2752, N3894);
nor NOR2 (N5065, N5064, N1059);
xor XOR2 (N5066, N5058, N3964);
nor NOR3 (N5067, N5053, N1037, N945);
buf BUF1 (N5068, N5066);
nand NAND2 (N5069, N5055, N3847);
and AND4 (N5070, N5068, N665, N4414, N2688);
or OR3 (N5071, N5059, N2143, N5036);
or OR3 (N5072, N5063, N3221, N1589);
xor XOR2 (N5073, N5037, N681);
not NOT1 (N5074, N5046);
and AND2 (N5075, N5073, N2427);
nand NAND2 (N5076, N5067, N2882);
not NOT1 (N5077, N5076);
nor NOR3 (N5078, N5077, N2786, N2871);
nand NAND3 (N5079, N5074, N828, N1713);
nand NAND2 (N5080, N5079, N775);
not NOT1 (N5081, N5070);
xor XOR2 (N5082, N5065, N580);
and AND4 (N5083, N5060, N2400, N3539, N1282);
buf BUF1 (N5084, N5083);
buf BUF1 (N5085, N5071);
and AND2 (N5086, N5072, N3956);
not NOT1 (N5087, N5086);
nand NAND2 (N5088, N5080, N1410);
or OR3 (N5089, N5085, N5037, N2962);
or OR3 (N5090, N5075, N4110, N274);
nand NAND2 (N5091, N5078, N2425);
and AND3 (N5092, N5081, N2975, N4337);
buf BUF1 (N5093, N5088);
nor NOR4 (N5094, N5093, N3531, N3071, N146);
not NOT1 (N5095, N5089);
and AND2 (N5096, N5062, N4764);
or OR4 (N5097, N5084, N3943, N2392, N2826);
or OR3 (N5098, N5090, N4598, N2275);
xor XOR2 (N5099, N5069, N3459);
nor NOR3 (N5100, N5092, N487, N4234);
buf BUF1 (N5101, N5087);
and AND2 (N5102, N5099, N921);
nand NAND3 (N5103, N5101, N917, N1783);
nand NAND3 (N5104, N5095, N2404, N3496);
nand NAND2 (N5105, N5094, N4003);
or OR3 (N5106, N5103, N3085, N3114);
buf BUF1 (N5107, N5100);
nor NOR4 (N5108, N5082, N330, N2969, N326);
nand NAND2 (N5109, N5108, N1988);
nor NOR3 (N5110, N5107, N3506, N2847);
xor XOR2 (N5111, N5097, N4979);
nand NAND2 (N5112, N5111, N3401);
or OR4 (N5113, N5110, N4872, N273, N1487);
xor XOR2 (N5114, N5096, N1277);
buf BUF1 (N5115, N5112);
or OR4 (N5116, N5098, N122, N3520, N3013);
and AND3 (N5117, N5115, N2001, N2314);
and AND4 (N5118, N5105, N2894, N2407, N24);
not NOT1 (N5119, N5102);
or OR3 (N5120, N5109, N4564, N1437);
not NOT1 (N5121, N5114);
or OR4 (N5122, N5118, N4231, N4658, N357);
buf BUF1 (N5123, N5113);
nor NOR2 (N5124, N5120, N4666);
or OR2 (N5125, N5104, N624);
nand NAND4 (N5126, N5121, N3939, N5031, N4041);
or OR3 (N5127, N5125, N1713, N2408);
or OR2 (N5128, N5119, N2028);
nand NAND4 (N5129, N5106, N1059, N4155, N4132);
or OR2 (N5130, N5091, N970);
or OR4 (N5131, N5126, N4677, N3158, N3246);
and AND3 (N5132, N5116, N4299, N3094);
nor NOR4 (N5133, N5131, N2007, N3325, N2381);
nand NAND3 (N5134, N5129, N3140, N1678);
nand NAND4 (N5135, N5117, N867, N733, N1673);
not NOT1 (N5136, N5130);
nor NOR4 (N5137, N5135, N557, N2102, N1363);
not NOT1 (N5138, N5123);
or OR2 (N5139, N5132, N59);
nor NOR2 (N5140, N5138, N3614);
not NOT1 (N5141, N5124);
or OR2 (N5142, N5139, N5007);
not NOT1 (N5143, N5133);
nand NAND4 (N5144, N5122, N1329, N4799, N4698);
nor NOR3 (N5145, N5128, N4724, N2606);
nand NAND3 (N5146, N5142, N1602, N2593);
nor NOR3 (N5147, N5140, N3422, N3105);
not NOT1 (N5148, N5144);
nor NOR2 (N5149, N5146, N2243);
nor NOR2 (N5150, N5127, N2167);
and AND2 (N5151, N5134, N3390);
or OR3 (N5152, N5149, N2544, N3798);
buf BUF1 (N5153, N5143);
or OR4 (N5154, N5141, N202, N3262, N94);
and AND2 (N5155, N5154, N4601);
and AND3 (N5156, N5148, N1984, N2925);
buf BUF1 (N5157, N5137);
buf BUF1 (N5158, N5156);
buf BUF1 (N5159, N5158);
nand NAND4 (N5160, N5155, N2123, N949, N1571);
or OR3 (N5161, N5160, N2750, N1837);
nor NOR4 (N5162, N5152, N4687, N2648, N4951);
nand NAND3 (N5163, N5153, N738, N4798);
and AND4 (N5164, N5151, N1758, N1249, N3143);
nor NOR3 (N5165, N5147, N4130, N4421);
buf BUF1 (N5166, N5165);
or OR2 (N5167, N5136, N4439);
xor XOR2 (N5168, N5167, N4657);
xor XOR2 (N5169, N5162, N2911);
and AND4 (N5170, N5157, N2720, N1695, N3085);
nor NOR3 (N5171, N5145, N707, N3435);
nor NOR2 (N5172, N5159, N4072);
and AND4 (N5173, N5170, N1538, N2020, N3218);
and AND2 (N5174, N5161, N3367);
nor NOR3 (N5175, N5174, N3238, N1070);
xor XOR2 (N5176, N5175, N3701);
not NOT1 (N5177, N5163);
nand NAND3 (N5178, N5176, N1831, N4553);
or OR2 (N5179, N5173, N1352);
not NOT1 (N5180, N5179);
xor XOR2 (N5181, N5178, N1258);
nand NAND4 (N5182, N5177, N3835, N1751, N1913);
xor XOR2 (N5183, N5182, N3953);
not NOT1 (N5184, N5164);
buf BUF1 (N5185, N5169);
nor NOR4 (N5186, N5168, N183, N3733, N1751);
or OR4 (N5187, N5172, N3185, N2047, N4409);
or OR4 (N5188, N5185, N1480, N733, N203);
and AND2 (N5189, N5184, N1432);
and AND2 (N5190, N5166, N3120);
nand NAND2 (N5191, N5190, N5032);
xor XOR2 (N5192, N5187, N1880);
and AND2 (N5193, N5186, N2617);
not NOT1 (N5194, N5181);
buf BUF1 (N5195, N5188);
or OR2 (N5196, N5192, N4627);
or OR4 (N5197, N5196, N2350, N1380, N4616);
buf BUF1 (N5198, N5194);
xor XOR2 (N5199, N5171, N4178);
not NOT1 (N5200, N5189);
or OR4 (N5201, N5198, N1834, N2637, N3897);
nor NOR2 (N5202, N5201, N3393);
or OR2 (N5203, N5195, N2477);
buf BUF1 (N5204, N5183);
xor XOR2 (N5205, N5199, N1555);
not NOT1 (N5206, N5200);
buf BUF1 (N5207, N5193);
or OR4 (N5208, N5202, N4487, N447, N3876);
xor XOR2 (N5209, N5207, N713);
xor XOR2 (N5210, N5206, N2441);
nand NAND2 (N5211, N5208, N4225);
xor XOR2 (N5212, N5204, N2785);
nand NAND4 (N5213, N5180, N2866, N2785, N2558);
not NOT1 (N5214, N5203);
buf BUF1 (N5215, N5197);
or OR4 (N5216, N5211, N4195, N3876, N4141);
or OR4 (N5217, N5209, N4684, N1971, N4898);
xor XOR2 (N5218, N5210, N4843);
buf BUF1 (N5219, N5205);
or OR2 (N5220, N5191, N4455);
nand NAND4 (N5221, N5213, N4631, N88, N1011);
nor NOR2 (N5222, N5216, N4782);
buf BUF1 (N5223, N5220);
not NOT1 (N5224, N5218);
buf BUF1 (N5225, N5222);
not NOT1 (N5226, N5223);
and AND3 (N5227, N5226, N3277, N4492);
or OR4 (N5228, N5219, N1577, N4788, N22);
or OR4 (N5229, N5150, N446, N1879, N2539);
buf BUF1 (N5230, N5217);
nor NOR4 (N5231, N5228, N201, N4845, N2687);
not NOT1 (N5232, N5225);
nor NOR4 (N5233, N5227, N4087, N981, N1235);
xor XOR2 (N5234, N5230, N4817);
nor NOR2 (N5235, N5231, N2100);
nand NAND3 (N5236, N5234, N3419, N4083);
buf BUF1 (N5237, N5235);
nor NOR3 (N5238, N5229, N1194, N585);
nor NOR2 (N5239, N5238, N3512);
and AND2 (N5240, N5236, N1244);
or OR3 (N5241, N5214, N4102, N470);
not NOT1 (N5242, N5233);
and AND4 (N5243, N5241, N1186, N5198, N3404);
nand NAND3 (N5244, N5240, N1749, N1871);
not NOT1 (N5245, N5239);
nand NAND3 (N5246, N5232, N4403, N1445);
or OR4 (N5247, N5242, N3319, N1219, N4586);
and AND4 (N5248, N5212, N1624, N3252, N1455);
nor NOR4 (N5249, N5244, N1615, N3892, N5145);
nor NOR3 (N5250, N5215, N4960, N3968);
buf BUF1 (N5251, N5249);
or OR3 (N5252, N5250, N4774, N1961);
nor NOR2 (N5253, N5252, N4352);
or OR2 (N5254, N5243, N4955);
nor NOR4 (N5255, N5248, N1305, N3094, N603);
and AND4 (N5256, N5246, N3613, N4628, N138);
buf BUF1 (N5257, N5224);
buf BUF1 (N5258, N5254);
nand NAND3 (N5259, N5245, N4516, N2147);
xor XOR2 (N5260, N5237, N312);
and AND2 (N5261, N5256, N281);
nor NOR3 (N5262, N5255, N234, N2460);
xor XOR2 (N5263, N5258, N425);
and AND4 (N5264, N5260, N5183, N23, N383);
not NOT1 (N5265, N5259);
nand NAND4 (N5266, N5264, N4149, N5224, N2897);
not NOT1 (N5267, N5247);
not NOT1 (N5268, N5266);
not NOT1 (N5269, N5261);
nand NAND4 (N5270, N5257, N3297, N555, N4907);
or OR4 (N5271, N5268, N3173, N3646, N597);
xor XOR2 (N5272, N5253, N1512);
or OR2 (N5273, N5262, N640);
buf BUF1 (N5274, N5251);
buf BUF1 (N5275, N5272);
nand NAND4 (N5276, N5265, N2375, N4894, N1282);
not NOT1 (N5277, N5276);
nor NOR3 (N5278, N5221, N4683, N4040);
or OR4 (N5279, N5275, N442, N4789, N5029);
not NOT1 (N5280, N5274);
xor XOR2 (N5281, N5280, N5242);
nand NAND2 (N5282, N5278, N1070);
buf BUF1 (N5283, N5277);
buf BUF1 (N5284, N5267);
or OR2 (N5285, N5270, N2723);
xor XOR2 (N5286, N5282, N566);
nand NAND4 (N5287, N5284, N2791, N4176, N301);
xor XOR2 (N5288, N5287, N2627);
nor NOR3 (N5289, N5273, N83, N2412);
or OR4 (N5290, N5289, N2790, N328, N10);
nor NOR2 (N5291, N5288, N1404);
not NOT1 (N5292, N5290);
buf BUF1 (N5293, N5263);
or OR4 (N5294, N5285, N2279, N928, N3192);
xor XOR2 (N5295, N5293, N5036);
nand NAND3 (N5296, N5295, N2929, N413);
nand NAND2 (N5297, N5292, N2257);
not NOT1 (N5298, N5269);
nand NAND3 (N5299, N5281, N4258, N2789);
xor XOR2 (N5300, N5299, N3128);
xor XOR2 (N5301, N5279, N2937);
not NOT1 (N5302, N5296);
not NOT1 (N5303, N5297);
and AND4 (N5304, N5301, N339, N1500, N1282);
nand NAND2 (N5305, N5303, N2029);
buf BUF1 (N5306, N5305);
and AND3 (N5307, N5304, N849, N5246);
or OR2 (N5308, N5291, N1830);
nor NOR2 (N5309, N5306, N3197);
nor NOR3 (N5310, N5286, N1487, N4573);
not NOT1 (N5311, N5271);
nand NAND3 (N5312, N5309, N3519, N1085);
not NOT1 (N5313, N5312);
buf BUF1 (N5314, N5298);
nor NOR4 (N5315, N5310, N356, N2384, N401);
nor NOR4 (N5316, N5308, N3741, N2209, N2414);
not NOT1 (N5317, N5294);
nor NOR2 (N5318, N5313, N5279);
xor XOR2 (N5319, N5315, N3542);
nand NAND4 (N5320, N5316, N4517, N2653, N5296);
nor NOR3 (N5321, N5314, N338, N401);
buf BUF1 (N5322, N5317);
xor XOR2 (N5323, N5319, N1679);
buf BUF1 (N5324, N5283);
buf BUF1 (N5325, N5320);
or OR4 (N5326, N5323, N2054, N2669, N3667);
not NOT1 (N5327, N5302);
nor NOR2 (N5328, N5307, N5327);
or OR3 (N5329, N862, N1904, N1885);
not NOT1 (N5330, N5326);
and AND2 (N5331, N5325, N3665);
and AND4 (N5332, N5300, N674, N3552, N3149);
or OR4 (N5333, N5324, N5244, N985, N973);
nand NAND3 (N5334, N5321, N2650, N4163);
or OR3 (N5335, N5322, N2881, N2603);
xor XOR2 (N5336, N5329, N3716);
or OR4 (N5337, N5331, N2057, N379, N52);
not NOT1 (N5338, N5333);
not NOT1 (N5339, N5328);
nor NOR3 (N5340, N5332, N11, N2213);
and AND4 (N5341, N5339, N4859, N792, N417);
or OR4 (N5342, N5330, N2972, N2854, N1602);
and AND2 (N5343, N5318, N4727);
not NOT1 (N5344, N5343);
and AND3 (N5345, N5337, N1442, N4346);
buf BUF1 (N5346, N5336);
or OR3 (N5347, N5345, N2374, N592);
nand NAND3 (N5348, N5342, N4858, N2536);
or OR2 (N5349, N5348, N132);
nor NOR4 (N5350, N5346, N580, N2580, N584);
not NOT1 (N5351, N5338);
buf BUF1 (N5352, N5344);
buf BUF1 (N5353, N5352);
nand NAND3 (N5354, N5340, N1977, N750);
and AND2 (N5355, N5351, N2822);
xor XOR2 (N5356, N5347, N1391);
nor NOR4 (N5357, N5354, N3894, N2249, N4177);
nor NOR3 (N5358, N5335, N4970, N4827);
not NOT1 (N5359, N5350);
xor XOR2 (N5360, N5359, N4855);
buf BUF1 (N5361, N5356);
buf BUF1 (N5362, N5360);
nor NOR2 (N5363, N5361, N3990);
nor NOR2 (N5364, N5341, N2554);
nor NOR2 (N5365, N5358, N1939);
or OR3 (N5366, N5355, N3422, N4529);
buf BUF1 (N5367, N5357);
xor XOR2 (N5368, N5367, N3688);
and AND2 (N5369, N5349, N1395);
not NOT1 (N5370, N5364);
and AND4 (N5371, N5334, N4671, N2888, N4618);
not NOT1 (N5372, N5366);
nand NAND3 (N5373, N5353, N2515, N1548);
nor NOR3 (N5374, N5370, N3012, N1988);
or OR3 (N5375, N5371, N1282, N3651);
buf BUF1 (N5376, N5311);
nor NOR3 (N5377, N5369, N3085, N3501);
not NOT1 (N5378, N5372);
or OR3 (N5379, N5368, N4992, N5069);
nor NOR3 (N5380, N5376, N327, N2061);
not NOT1 (N5381, N5374);
or OR4 (N5382, N5380, N1223, N3323, N1086);
or OR3 (N5383, N5382, N659, N1013);
or OR3 (N5384, N5362, N2119, N2444);
and AND4 (N5385, N5365, N248, N1338, N288);
buf BUF1 (N5386, N5384);
not NOT1 (N5387, N5383);
and AND4 (N5388, N5381, N3744, N1621, N289);
nand NAND2 (N5389, N5377, N179);
xor XOR2 (N5390, N5378, N2911);
buf BUF1 (N5391, N5375);
or OR3 (N5392, N5390, N723, N4451);
and AND3 (N5393, N5379, N687, N473);
buf BUF1 (N5394, N5389);
nand NAND2 (N5395, N5387, N2055);
or OR3 (N5396, N5386, N3546, N953);
or OR2 (N5397, N5363, N5112);
or OR2 (N5398, N5388, N743);
nor NOR2 (N5399, N5385, N340);
or OR3 (N5400, N5373, N5265, N1810);
not NOT1 (N5401, N5392);
or OR3 (N5402, N5394, N4400, N585);
xor XOR2 (N5403, N5402, N4603);
not NOT1 (N5404, N5401);
and AND2 (N5405, N5397, N352);
and AND3 (N5406, N5399, N4298, N480);
and AND4 (N5407, N5395, N3227, N2253, N3037);
nand NAND2 (N5408, N5403, N205);
nand NAND2 (N5409, N5400, N2098);
and AND2 (N5410, N5398, N2403);
not NOT1 (N5411, N5406);
nand NAND3 (N5412, N5393, N688, N4091);
nor NOR2 (N5413, N5407, N4282);
buf BUF1 (N5414, N5408);
not NOT1 (N5415, N5396);
buf BUF1 (N5416, N5404);
and AND2 (N5417, N5405, N5404);
nor NOR4 (N5418, N5416, N3256, N3678, N2358);
xor XOR2 (N5419, N5391, N3537);
nor NOR3 (N5420, N5415, N613, N3832);
nor NOR3 (N5421, N5412, N126, N1155);
or OR2 (N5422, N5409, N3557);
nor NOR2 (N5423, N5422, N4823);
xor XOR2 (N5424, N5421, N2523);
nor NOR4 (N5425, N5410, N3413, N2525, N3257);
nand NAND3 (N5426, N5419, N4576, N2308);
nand NAND3 (N5427, N5413, N4738, N4499);
not NOT1 (N5428, N5427);
and AND2 (N5429, N5411, N5026);
not NOT1 (N5430, N5418);
or OR3 (N5431, N5430, N230, N2860);
or OR4 (N5432, N5423, N1959, N836, N5114);
nor NOR3 (N5433, N5431, N2963, N2489);
xor XOR2 (N5434, N5429, N3937);
xor XOR2 (N5435, N5420, N294);
nor NOR3 (N5436, N5425, N858, N428);
nor NOR3 (N5437, N5435, N2975, N1773);
nor NOR2 (N5438, N5426, N2401);
and AND3 (N5439, N5433, N129, N1093);
nor NOR2 (N5440, N5436, N322);
and AND4 (N5441, N5424, N1553, N1225, N5055);
not NOT1 (N5442, N5439);
nand NAND2 (N5443, N5438, N1713);
buf BUF1 (N5444, N5441);
nor NOR3 (N5445, N5414, N4110, N1648);
xor XOR2 (N5446, N5428, N4570);
nor NOR3 (N5447, N5417, N3296, N1990);
and AND4 (N5448, N5443, N4821, N2666, N2582);
not NOT1 (N5449, N5434);
nor NOR4 (N5450, N5440, N2638, N3843, N3923);
not NOT1 (N5451, N5432);
nor NOR4 (N5452, N5437, N2596, N274, N5198);
nand NAND3 (N5453, N5452, N2093, N1120);
buf BUF1 (N5454, N5449);
or OR3 (N5455, N5442, N3801, N2112);
nor NOR4 (N5456, N5445, N3774, N392, N4523);
nor NOR3 (N5457, N5448, N3815, N1572);
xor XOR2 (N5458, N5456, N1507);
or OR3 (N5459, N5444, N2890, N3139);
xor XOR2 (N5460, N5453, N1247);
nand NAND4 (N5461, N5451, N3072, N2448, N1443);
and AND2 (N5462, N5457, N2880);
and AND2 (N5463, N5455, N4103);
nand NAND2 (N5464, N5461, N2486);
xor XOR2 (N5465, N5462, N4766);
xor XOR2 (N5466, N5460, N1644);
nand NAND4 (N5467, N5466, N871, N1991, N3418);
xor XOR2 (N5468, N5454, N1536);
buf BUF1 (N5469, N5463);
not NOT1 (N5470, N5467);
and AND4 (N5471, N5459, N2502, N1965, N1278);
not NOT1 (N5472, N5468);
or OR4 (N5473, N5464, N2819, N2804, N887);
xor XOR2 (N5474, N5450, N1465);
nand NAND3 (N5475, N5465, N390, N117);
buf BUF1 (N5476, N5447);
or OR3 (N5477, N5474, N1237, N1428);
and AND4 (N5478, N5458, N4478, N138, N4372);
xor XOR2 (N5479, N5469, N832);
and AND3 (N5480, N5473, N1904, N1032);
nor NOR4 (N5481, N5446, N1989, N5191, N2742);
or OR4 (N5482, N5472, N489, N559, N21);
nor NOR3 (N5483, N5479, N597, N417);
buf BUF1 (N5484, N5482);
or OR3 (N5485, N5476, N403, N2210);
nor NOR4 (N5486, N5483, N4603, N3880, N2560);
or OR3 (N5487, N5478, N2570, N1168);
nand NAND4 (N5488, N5470, N1185, N5299, N549);
or OR2 (N5489, N5487, N3258);
or OR4 (N5490, N5489, N5161, N2284, N2444);
nor NOR4 (N5491, N5488, N1132, N1712, N4042);
and AND2 (N5492, N5485, N721);
buf BUF1 (N5493, N5471);
not NOT1 (N5494, N5492);
or OR4 (N5495, N5486, N4061, N4654, N5254);
nor NOR2 (N5496, N5493, N978);
buf BUF1 (N5497, N5496);
not NOT1 (N5498, N5491);
buf BUF1 (N5499, N5475);
xor XOR2 (N5500, N5477, N3332);
xor XOR2 (N5501, N5498, N3858);
nand NAND3 (N5502, N5480, N5404, N3422);
xor XOR2 (N5503, N5490, N2015);
xor XOR2 (N5504, N5495, N1435);
nor NOR2 (N5505, N5484, N1294);
or OR4 (N5506, N5500, N1952, N4060, N3184);
not NOT1 (N5507, N5499);
nor NOR2 (N5508, N5506, N2145);
not NOT1 (N5509, N5504);
or OR3 (N5510, N5509, N1403, N2724);
nand NAND3 (N5511, N5494, N1907, N4247);
nor NOR3 (N5512, N5507, N4790, N1994);
nand NAND4 (N5513, N5501, N436, N4684, N1600);
buf BUF1 (N5514, N5481);
xor XOR2 (N5515, N5514, N4536);
and AND3 (N5516, N5505, N59, N2879);
nand NAND2 (N5517, N5516, N5355);
nand NAND4 (N5518, N5511, N1397, N2996, N1520);
and AND4 (N5519, N5510, N610, N1026, N2892);
not NOT1 (N5520, N5513);
nand NAND3 (N5521, N5502, N4392, N2759);
buf BUF1 (N5522, N5517);
nor NOR3 (N5523, N5522, N2249, N1311);
and AND4 (N5524, N5508, N4597, N1860, N5180);
not NOT1 (N5525, N5520);
and AND2 (N5526, N5503, N639);
buf BUF1 (N5527, N5526);
and AND3 (N5528, N5518, N135, N1457);
nand NAND3 (N5529, N5519, N4779, N2592);
not NOT1 (N5530, N5527);
nand NAND4 (N5531, N5528, N2923, N2151, N762);
nand NAND3 (N5532, N5530, N1495, N191);
and AND2 (N5533, N5525, N4161);
buf BUF1 (N5534, N5533);
buf BUF1 (N5535, N5524);
buf BUF1 (N5536, N5521);
nand NAND3 (N5537, N5515, N1831, N458);
not NOT1 (N5538, N5536);
buf BUF1 (N5539, N5537);
buf BUF1 (N5540, N5538);
xor XOR2 (N5541, N5534, N5188);
nor NOR4 (N5542, N5539, N5392, N5127, N3292);
or OR3 (N5543, N5512, N1968, N2909);
buf BUF1 (N5544, N5542);
or OR4 (N5545, N5541, N1221, N3805, N122);
xor XOR2 (N5546, N5545, N4530);
nor NOR4 (N5547, N5523, N2699, N792, N4168);
nor NOR2 (N5548, N5529, N2526);
or OR2 (N5549, N5547, N4978);
nand NAND4 (N5550, N5543, N369, N1943, N3752);
and AND2 (N5551, N5540, N3192);
not NOT1 (N5552, N5544);
nor NOR3 (N5553, N5546, N1938, N4855);
not NOT1 (N5554, N5531);
not NOT1 (N5555, N5535);
buf BUF1 (N5556, N5548);
or OR4 (N5557, N5497, N505, N4930, N3445);
xor XOR2 (N5558, N5556, N3327);
nand NAND3 (N5559, N5557, N5338, N4119);
nor NOR2 (N5560, N5558, N4163);
nor NOR2 (N5561, N5532, N5401);
and AND4 (N5562, N5554, N4075, N5210, N2480);
xor XOR2 (N5563, N5549, N5195);
xor XOR2 (N5564, N5559, N3593);
and AND4 (N5565, N5552, N3211, N1884, N125);
buf BUF1 (N5566, N5561);
not NOT1 (N5567, N5551);
and AND3 (N5568, N5562, N1249, N5399);
buf BUF1 (N5569, N5564);
and AND3 (N5570, N5568, N191, N4671);
not NOT1 (N5571, N5553);
nand NAND2 (N5572, N5567, N2729);
not NOT1 (N5573, N5570);
xor XOR2 (N5574, N5563, N1388);
buf BUF1 (N5575, N5560);
or OR4 (N5576, N5571, N3537, N3074, N1879);
or OR4 (N5577, N5566, N2372, N1084, N3157);
and AND4 (N5578, N5569, N4436, N2861, N4114);
nor NOR3 (N5579, N5576, N352, N492);
nand NAND4 (N5580, N5577, N3845, N408, N5291);
not NOT1 (N5581, N5580);
or OR2 (N5582, N5575, N926);
and AND4 (N5583, N5572, N1252, N949, N5116);
nand NAND3 (N5584, N5579, N2212, N2046);
nand NAND3 (N5585, N5573, N2169, N2143);
nor NOR3 (N5586, N5550, N1481, N2606);
not NOT1 (N5587, N5583);
nor NOR4 (N5588, N5586, N1809, N5008, N701);
and AND2 (N5589, N5587, N1993);
xor XOR2 (N5590, N5589, N1028);
and AND3 (N5591, N5585, N3931, N4677);
xor XOR2 (N5592, N5574, N5);
nand NAND3 (N5593, N5582, N1959, N4423);
buf BUF1 (N5594, N5593);
and AND2 (N5595, N5588, N5248);
not NOT1 (N5596, N5590);
nand NAND3 (N5597, N5578, N2126, N4725);
and AND4 (N5598, N5584, N45, N2506, N4953);
not NOT1 (N5599, N5594);
and AND4 (N5600, N5565, N1941, N2798, N1301);
nor NOR4 (N5601, N5592, N2441, N4147, N624);
nor NOR4 (N5602, N5555, N5483, N3650, N5394);
buf BUF1 (N5603, N5591);
nand NAND4 (N5604, N5595, N4519, N4943, N2510);
not NOT1 (N5605, N5581);
not NOT1 (N5606, N5597);
buf BUF1 (N5607, N5601);
or OR2 (N5608, N5606, N274);
and AND4 (N5609, N5607, N2223, N3406, N2128);
or OR3 (N5610, N5603, N3670, N1512);
xor XOR2 (N5611, N5602, N450);
nor NOR4 (N5612, N5605, N3655, N868, N285);
xor XOR2 (N5613, N5610, N3741);
or OR4 (N5614, N5612, N2871, N3321, N5593);
and AND4 (N5615, N5599, N5458, N1322, N4499);
nand NAND4 (N5616, N5615, N1714, N5517, N5348);
and AND4 (N5617, N5611, N5445, N5154, N603);
or OR3 (N5618, N5616, N4598, N4581);
or OR4 (N5619, N5609, N2215, N2775, N1201);
or OR3 (N5620, N5614, N999, N1694);
not NOT1 (N5621, N5598);
and AND2 (N5622, N5608, N4182);
nor NOR4 (N5623, N5604, N2732, N3564, N474);
buf BUF1 (N5624, N5623);
and AND2 (N5625, N5621, N3728);
and AND2 (N5626, N5596, N3413);
xor XOR2 (N5627, N5613, N3867);
nor NOR4 (N5628, N5626, N2429, N4435, N351);
nor NOR3 (N5629, N5622, N835, N3736);
nor NOR4 (N5630, N5625, N3083, N2035, N4868);
xor XOR2 (N5631, N5628, N4903);
and AND4 (N5632, N5617, N1018, N3635, N4081);
not NOT1 (N5633, N5632);
xor XOR2 (N5634, N5620, N242);
xor XOR2 (N5635, N5631, N5491);
buf BUF1 (N5636, N5629);
nor NOR4 (N5637, N5634, N4524, N4207, N772);
xor XOR2 (N5638, N5630, N1120);
nor NOR2 (N5639, N5635, N2898);
and AND3 (N5640, N5633, N4318, N1748);
nor NOR4 (N5641, N5639, N2754, N4180, N4375);
not NOT1 (N5642, N5640);
or OR3 (N5643, N5642, N110, N5373);
nor NOR3 (N5644, N5619, N3666, N5107);
or OR4 (N5645, N5600, N5074, N240, N4724);
and AND2 (N5646, N5641, N2545);
buf BUF1 (N5647, N5636);
and AND4 (N5648, N5647, N3424, N663, N3737);
and AND3 (N5649, N5645, N777, N72);
nor NOR3 (N5650, N5627, N3787, N4134);
not NOT1 (N5651, N5649);
or OR3 (N5652, N5638, N954, N2429);
buf BUF1 (N5653, N5652);
or OR2 (N5654, N5648, N4885);
and AND2 (N5655, N5653, N946);
not NOT1 (N5656, N5654);
buf BUF1 (N5657, N5646);
and AND4 (N5658, N5651, N837, N987, N2505);
xor XOR2 (N5659, N5656, N1435);
not NOT1 (N5660, N5657);
or OR2 (N5661, N5660, N2840);
xor XOR2 (N5662, N5637, N2876);
xor XOR2 (N5663, N5643, N830);
nor NOR4 (N5664, N5644, N1035, N3470, N4221);
not NOT1 (N5665, N5661);
not NOT1 (N5666, N5618);
nor NOR4 (N5667, N5664, N2237, N99, N1006);
and AND2 (N5668, N5665, N4933);
nand NAND3 (N5669, N5667, N2954, N3064);
or OR3 (N5670, N5658, N3758, N2476);
buf BUF1 (N5671, N5624);
nor NOR2 (N5672, N5669, N3790);
xor XOR2 (N5673, N5670, N5439);
not NOT1 (N5674, N5659);
or OR2 (N5675, N5674, N1399);
xor XOR2 (N5676, N5650, N2538);
nor NOR4 (N5677, N5666, N2635, N545, N4341);
and AND2 (N5678, N5668, N4012);
nand NAND4 (N5679, N5662, N5641, N2829, N94);
nor NOR2 (N5680, N5676, N4381);
xor XOR2 (N5681, N5671, N4246);
nand NAND3 (N5682, N5678, N4055, N1891);
not NOT1 (N5683, N5672);
nor NOR2 (N5684, N5683, N897);
or OR3 (N5685, N5673, N5652, N1214);
not NOT1 (N5686, N5684);
and AND3 (N5687, N5682, N3686, N4792);
buf BUF1 (N5688, N5687);
nor NOR2 (N5689, N5688, N1545);
not NOT1 (N5690, N5677);
not NOT1 (N5691, N5690);
nand NAND3 (N5692, N5686, N1558, N4429);
not NOT1 (N5693, N5680);
nand NAND4 (N5694, N5693, N3378, N209, N4896);
buf BUF1 (N5695, N5679);
nand NAND3 (N5696, N5675, N700, N2250);
xor XOR2 (N5697, N5694, N3343);
nand NAND4 (N5698, N5695, N590, N3703, N94);
or OR3 (N5699, N5698, N2696, N4513);
nand NAND4 (N5700, N5681, N2651, N3292, N1464);
buf BUF1 (N5701, N5699);
or OR2 (N5702, N5691, N5147);
and AND3 (N5703, N5702, N2000, N4483);
buf BUF1 (N5704, N5701);
not NOT1 (N5705, N5655);
and AND3 (N5706, N5663, N5319, N4460);
buf BUF1 (N5707, N5706);
and AND2 (N5708, N5685, N3138);
and AND2 (N5709, N5696, N1841);
nor NOR3 (N5710, N5692, N831, N5069);
nand NAND3 (N5711, N5704, N3431, N5374);
xor XOR2 (N5712, N5708, N5139);
buf BUF1 (N5713, N5703);
nor NOR2 (N5714, N5713, N3335);
not NOT1 (N5715, N5707);
and AND2 (N5716, N5689, N1422);
not NOT1 (N5717, N5716);
or OR4 (N5718, N5711, N3301, N108, N3662);
nor NOR3 (N5719, N5705, N4225, N1315);
or OR4 (N5720, N5710, N4171, N3256, N3162);
not NOT1 (N5721, N5700);
buf BUF1 (N5722, N5717);
not NOT1 (N5723, N5720);
or OR4 (N5724, N5714, N2126, N5278, N5231);
buf BUF1 (N5725, N5712);
nand NAND2 (N5726, N5723, N1071);
or OR4 (N5727, N5718, N1369, N520, N3507);
buf BUF1 (N5728, N5726);
nand NAND4 (N5729, N5725, N2266, N3666, N2196);
nand NAND3 (N5730, N5728, N4893, N3413);
buf BUF1 (N5731, N5722);
xor XOR2 (N5732, N5715, N2208);
buf BUF1 (N5733, N5730);
not NOT1 (N5734, N5697);
nor NOR2 (N5735, N5732, N240);
xor XOR2 (N5736, N5735, N4536);
nor NOR2 (N5737, N5731, N5463);
nand NAND2 (N5738, N5727, N1208);
not NOT1 (N5739, N5736);
nor NOR4 (N5740, N5709, N3342, N3958, N1330);
or OR3 (N5741, N5729, N2065, N1676);
nand NAND3 (N5742, N5737, N4608, N4504);
nor NOR2 (N5743, N5741, N423);
nor NOR3 (N5744, N5719, N1348, N2192);
xor XOR2 (N5745, N5740, N5441);
buf BUF1 (N5746, N5742);
or OR3 (N5747, N5746, N1826, N3558);
or OR2 (N5748, N5734, N2682);
or OR3 (N5749, N5738, N825, N3320);
nor NOR4 (N5750, N5747, N3735, N726, N2142);
and AND4 (N5751, N5748, N3227, N4821, N4419);
nor NOR4 (N5752, N5721, N4621, N2005, N504);
and AND3 (N5753, N5745, N3598, N2012);
or OR3 (N5754, N5749, N5088, N3387);
buf BUF1 (N5755, N5753);
or OR4 (N5756, N5744, N5293, N3750, N664);
nand NAND4 (N5757, N5750, N5263, N375, N1152);
and AND3 (N5758, N5743, N1816, N2447);
not NOT1 (N5759, N5757);
not NOT1 (N5760, N5754);
xor XOR2 (N5761, N5756, N3061);
not NOT1 (N5762, N5755);
nor NOR4 (N5763, N5760, N1602, N3328, N2569);
or OR3 (N5764, N5762, N2284, N804);
not NOT1 (N5765, N5733);
and AND4 (N5766, N5758, N2376, N3049, N2615);
nor NOR3 (N5767, N5752, N4615, N2140);
buf BUF1 (N5768, N5751);
and AND2 (N5769, N5724, N5256);
nor NOR4 (N5770, N5765, N2024, N1503, N2824);
nor NOR2 (N5771, N5768, N2218);
buf BUF1 (N5772, N5771);
buf BUF1 (N5773, N5767);
buf BUF1 (N5774, N5761);
and AND2 (N5775, N5763, N5076);
nor NOR3 (N5776, N5766, N5203, N5008);
buf BUF1 (N5777, N5775);
not NOT1 (N5778, N5759);
not NOT1 (N5779, N5772);
not NOT1 (N5780, N5739);
nor NOR4 (N5781, N5769, N1863, N4645, N5725);
nor NOR4 (N5782, N5770, N3812, N4770, N5069);
or OR2 (N5783, N5779, N2527);
and AND3 (N5784, N5780, N4281, N2405);
buf BUF1 (N5785, N5778);
nor NOR4 (N5786, N5777, N2286, N4054, N2455);
nor NOR3 (N5787, N5782, N1486, N889);
or OR4 (N5788, N5774, N1859, N3686, N2375);
xor XOR2 (N5789, N5786, N2269);
xor XOR2 (N5790, N5784, N825);
or OR4 (N5791, N5781, N4173, N245, N1666);
nand NAND4 (N5792, N5764, N3829, N1289, N5763);
nand NAND4 (N5793, N5788, N1350, N5268, N5777);
not NOT1 (N5794, N5785);
nand NAND3 (N5795, N5794, N1695, N5361);
xor XOR2 (N5796, N5791, N127);
buf BUF1 (N5797, N5783);
not NOT1 (N5798, N5776);
and AND3 (N5799, N5773, N4778, N2161);
buf BUF1 (N5800, N5790);
nor NOR3 (N5801, N5793, N3851, N1576);
or OR4 (N5802, N5797, N669, N4949, N1956);
not NOT1 (N5803, N5800);
buf BUF1 (N5804, N5792);
buf BUF1 (N5805, N5798);
nor NOR2 (N5806, N5796, N3268);
xor XOR2 (N5807, N5802, N5595);
nand NAND3 (N5808, N5803, N3966, N508);
or OR2 (N5809, N5799, N4347);
not NOT1 (N5810, N5807);
buf BUF1 (N5811, N5804);
nand NAND4 (N5812, N5806, N4259, N1317, N4643);
nor NOR4 (N5813, N5809, N5043, N1467, N2893);
nor NOR2 (N5814, N5805, N1744);
nand NAND4 (N5815, N5813, N1345, N1994, N3441);
and AND3 (N5816, N5801, N4632, N633);
nand NAND3 (N5817, N5816, N303, N5746);
or OR3 (N5818, N5787, N1902, N4887);
buf BUF1 (N5819, N5818);
not NOT1 (N5820, N5814);
nor NOR3 (N5821, N5808, N2687, N2917);
nand NAND2 (N5822, N5817, N5054);
not NOT1 (N5823, N5795);
or OR4 (N5824, N5789, N461, N4388, N1143);
or OR4 (N5825, N5822, N2327, N4431, N2760);
nand NAND4 (N5826, N5810, N4564, N74, N1718);
buf BUF1 (N5827, N5824);
nor NOR4 (N5828, N5826, N724, N4117, N7);
buf BUF1 (N5829, N5823);
nand NAND4 (N5830, N5812, N5428, N4064, N2886);
xor XOR2 (N5831, N5815, N1412);
nor NOR3 (N5832, N5830, N5819, N4186);
nor NOR3 (N5833, N1907, N4658, N2153);
nand NAND3 (N5834, N5829, N2049, N5647);
nor NOR2 (N5835, N5832, N3348);
buf BUF1 (N5836, N5827);
and AND2 (N5837, N5835, N2526);
or OR2 (N5838, N5820, N5627);
nand NAND4 (N5839, N5838, N2914, N1463, N2152);
nand NAND4 (N5840, N5811, N1565, N2654, N3686);
nor NOR2 (N5841, N5831, N4279);
and AND4 (N5842, N5833, N1181, N4176, N499);
and AND3 (N5843, N5834, N1328, N5643);
xor XOR2 (N5844, N5836, N4405);
and AND4 (N5845, N5842, N5365, N5640, N5496);
not NOT1 (N5846, N5825);
or OR4 (N5847, N5845, N999, N4259, N3384);
buf BUF1 (N5848, N5837);
buf BUF1 (N5849, N5840);
nand NAND4 (N5850, N5847, N2609, N2861, N5485);
nand NAND3 (N5851, N5849, N1953, N935);
and AND2 (N5852, N5841, N1793);
or OR3 (N5853, N5850, N2971, N1762);
buf BUF1 (N5854, N5852);
nor NOR2 (N5855, N5853, N5738);
buf BUF1 (N5856, N5846);
and AND4 (N5857, N5851, N3057, N3821, N151);
not NOT1 (N5858, N5839);
and AND4 (N5859, N5858, N3456, N3848, N4806);
or OR2 (N5860, N5854, N3179);
xor XOR2 (N5861, N5860, N138);
or OR4 (N5862, N5855, N89, N5628, N3531);
not NOT1 (N5863, N5857);
xor XOR2 (N5864, N5828, N2804);
nand NAND2 (N5865, N5848, N2366);
and AND4 (N5866, N5821, N1913, N2131, N3185);
not NOT1 (N5867, N5862);
nor NOR4 (N5868, N5864, N2522, N437, N3849);
xor XOR2 (N5869, N5865, N4153);
and AND4 (N5870, N5856, N3761, N983, N3505);
nand NAND2 (N5871, N5844, N2497);
or OR2 (N5872, N5843, N3090);
nor NOR3 (N5873, N5868, N110, N4250);
and AND2 (N5874, N5867, N2062);
or OR4 (N5875, N5859, N1100, N2749, N2923);
buf BUF1 (N5876, N5874);
buf BUF1 (N5877, N5869);
nand NAND4 (N5878, N5872, N4424, N5867, N187);
xor XOR2 (N5879, N5870, N391);
xor XOR2 (N5880, N5861, N5801);
not NOT1 (N5881, N5866);
buf BUF1 (N5882, N5871);
nor NOR4 (N5883, N5878, N1324, N1052, N5609);
and AND4 (N5884, N5877, N2054, N2514, N2767);
buf BUF1 (N5885, N5882);
not NOT1 (N5886, N5873);
or OR4 (N5887, N5883, N4187, N2628, N2137);
and AND3 (N5888, N5879, N2050, N1171);
not NOT1 (N5889, N5863);
xor XOR2 (N5890, N5887, N5558);
buf BUF1 (N5891, N5890);
not NOT1 (N5892, N5891);
xor XOR2 (N5893, N5880, N2920);
buf BUF1 (N5894, N5881);
nand NAND3 (N5895, N5884, N4188, N4284);
or OR3 (N5896, N5886, N809, N2504);
and AND2 (N5897, N5892, N2253);
xor XOR2 (N5898, N5889, N4983);
and AND4 (N5899, N5894, N115, N4143, N5339);
nand NAND4 (N5900, N5896, N3760, N4832, N2318);
nor NOR2 (N5901, N5897, N5500);
not NOT1 (N5902, N5901);
nand NAND3 (N5903, N5885, N1383, N5683);
buf BUF1 (N5904, N5903);
or OR3 (N5905, N5902, N763, N3210);
or OR2 (N5906, N5899, N2722);
and AND3 (N5907, N5895, N5044, N3745);
and AND2 (N5908, N5898, N4973);
not NOT1 (N5909, N5888);
nor NOR3 (N5910, N5904, N3326, N521);
buf BUF1 (N5911, N5893);
buf BUF1 (N5912, N5875);
xor XOR2 (N5913, N5907, N1216);
nor NOR3 (N5914, N5909, N184, N5264);
xor XOR2 (N5915, N5914, N5054);
not NOT1 (N5916, N5912);
buf BUF1 (N5917, N5913);
or OR4 (N5918, N5917, N1, N859, N19);
nand NAND4 (N5919, N5905, N3184, N5042, N1486);
xor XOR2 (N5920, N5919, N5828);
buf BUF1 (N5921, N5911);
xor XOR2 (N5922, N5900, N5067);
or OR2 (N5923, N5921, N2550);
or OR2 (N5924, N5908, N3045);
and AND4 (N5925, N5922, N484, N5036, N3832);
or OR4 (N5926, N5915, N1513, N3667, N733);
xor XOR2 (N5927, N5910, N1021);
or OR3 (N5928, N5923, N1870, N518);
buf BUF1 (N5929, N5927);
not NOT1 (N5930, N5924);
and AND4 (N5931, N5918, N3058, N2412, N382);
not NOT1 (N5932, N5930);
or OR4 (N5933, N5906, N3287, N4382, N1910);
nand NAND3 (N5934, N5876, N73, N5120);
xor XOR2 (N5935, N5925, N3317);
nand NAND2 (N5936, N5920, N1805);
and AND4 (N5937, N5934, N169, N2529, N1377);
nor NOR2 (N5938, N5929, N1090);
or OR4 (N5939, N5928, N4057, N1894, N5084);
nor NOR4 (N5940, N5936, N1191, N4876, N730);
or OR4 (N5941, N5926, N1732, N4144, N360);
or OR3 (N5942, N5931, N2357, N768);
not NOT1 (N5943, N5938);
buf BUF1 (N5944, N5937);
nor NOR3 (N5945, N5940, N1478, N3974);
not NOT1 (N5946, N5932);
and AND3 (N5947, N5933, N2418, N40);
and AND2 (N5948, N5941, N2017);
nor NOR4 (N5949, N5945, N4719, N4330, N5445);
nand NAND2 (N5950, N5939, N4442);
nor NOR4 (N5951, N5948, N1874, N3549, N5682);
and AND4 (N5952, N5946, N2384, N900, N1215);
nor NOR2 (N5953, N5947, N1574);
and AND2 (N5954, N5944, N633);
nand NAND2 (N5955, N5935, N5330);
or OR2 (N5956, N5943, N1973);
or OR4 (N5957, N5955, N5438, N2872, N1455);
or OR3 (N5958, N5956, N1161, N40);
nand NAND4 (N5959, N5957, N5709, N3764, N4603);
or OR2 (N5960, N5953, N331);
not NOT1 (N5961, N5916);
xor XOR2 (N5962, N5950, N736);
not NOT1 (N5963, N5954);
buf BUF1 (N5964, N5952);
nand NAND3 (N5965, N5960, N2683, N4465);
not NOT1 (N5966, N5962);
buf BUF1 (N5967, N5964);
nor NOR3 (N5968, N5949, N2016, N485);
buf BUF1 (N5969, N5967);
nand NAND4 (N5970, N5968, N3107, N5308, N5517);
nor NOR3 (N5971, N5958, N4766, N875);
buf BUF1 (N5972, N5951);
and AND4 (N5973, N5972, N1566, N4327, N2698);
xor XOR2 (N5974, N5963, N2148);
buf BUF1 (N5975, N5942);
buf BUF1 (N5976, N5970);
nand NAND3 (N5977, N5974, N3463, N711);
nor NOR3 (N5978, N5971, N2989, N1482);
nand NAND3 (N5979, N5978, N2991, N5830);
not NOT1 (N5980, N5977);
and AND3 (N5981, N5966, N4494, N3048);
nand NAND3 (N5982, N5975, N1305, N2629);
nor NOR3 (N5983, N5959, N1541, N4035);
not NOT1 (N5984, N5980);
or OR3 (N5985, N5961, N3451, N5915);
nand NAND3 (N5986, N5976, N499, N4035);
buf BUF1 (N5987, N5979);
nor NOR3 (N5988, N5981, N5052, N5282);
xor XOR2 (N5989, N5965, N3289);
nor NOR3 (N5990, N5983, N5256, N4939);
or OR3 (N5991, N5988, N5242, N2028);
or OR2 (N5992, N5987, N2858);
not NOT1 (N5993, N5990);
xor XOR2 (N5994, N5985, N1001);
nand NAND4 (N5995, N5984, N4811, N5296, N4806);
not NOT1 (N5996, N5992);
or OR3 (N5997, N5982, N876, N3991);
or OR3 (N5998, N5973, N1588, N2412);
buf BUF1 (N5999, N5991);
not NOT1 (N6000, N5989);
nand NAND2 (N6001, N5995, N2801);
and AND2 (N6002, N5994, N3334);
buf BUF1 (N6003, N5997);
nor NOR4 (N6004, N6003, N4716, N959, N2912);
or OR4 (N6005, N6000, N2185, N1376, N3855);
and AND3 (N6006, N6002, N3537, N2383);
nor NOR4 (N6007, N5993, N4365, N1240, N1788);
buf BUF1 (N6008, N6004);
not NOT1 (N6009, N6005);
buf BUF1 (N6010, N5998);
nor NOR3 (N6011, N6001, N5456, N1220);
buf BUF1 (N6012, N5969);
buf BUF1 (N6013, N6006);
nor NOR2 (N6014, N6012, N729);
xor XOR2 (N6015, N6014, N3592);
nand NAND2 (N6016, N6011, N4891);
nand NAND3 (N6017, N6013, N3981, N3153);
not NOT1 (N6018, N6010);
and AND2 (N6019, N6009, N4281);
not NOT1 (N6020, N5996);
and AND3 (N6021, N6008, N6016, N829);
nor NOR2 (N6022, N1124, N774);
not NOT1 (N6023, N6018);
xor XOR2 (N6024, N6007, N5429);
nor NOR4 (N6025, N6015, N2610, N1711, N3027);
xor XOR2 (N6026, N6025, N462);
xor XOR2 (N6027, N6019, N3775);
nor NOR3 (N6028, N6017, N3047, N160);
not NOT1 (N6029, N6022);
nand NAND3 (N6030, N6021, N3182, N2462);
buf BUF1 (N6031, N6029);
buf BUF1 (N6032, N6024);
or OR4 (N6033, N6027, N2977, N5589, N935);
nand NAND4 (N6034, N6028, N5755, N4855, N3992);
not NOT1 (N6035, N6020);
nand NAND3 (N6036, N6026, N1406, N1419);
nor NOR3 (N6037, N6032, N562, N4477);
and AND4 (N6038, N6035, N3991, N1110, N4745);
nand NAND2 (N6039, N6038, N2179);
xor XOR2 (N6040, N6023, N633);
nor NOR3 (N6041, N6037, N263, N3260);
or OR2 (N6042, N6031, N5420);
buf BUF1 (N6043, N6036);
or OR4 (N6044, N6042, N1427, N4532, N4136);
nand NAND2 (N6045, N6034, N5026);
not NOT1 (N6046, N6045);
not NOT1 (N6047, N6039);
nor NOR4 (N6048, N6041, N91, N2293, N1609);
and AND4 (N6049, N5999, N5039, N2044, N4431);
buf BUF1 (N6050, N6043);
not NOT1 (N6051, N6030);
not NOT1 (N6052, N6044);
and AND3 (N6053, N6050, N1587, N3078);
xor XOR2 (N6054, N6033, N1352);
and AND2 (N6055, N6053, N2551);
nor NOR2 (N6056, N6054, N3640);
and AND4 (N6057, N6056, N4068, N1346, N1709);
not NOT1 (N6058, N6055);
or OR4 (N6059, N6048, N5655, N1469, N4698);
nor NOR4 (N6060, N6057, N3747, N2511, N5386);
nor NOR2 (N6061, N6047, N4050);
not NOT1 (N6062, N6061);
xor XOR2 (N6063, N6040, N1690);
nand NAND2 (N6064, N6059, N2965);
xor XOR2 (N6065, N6063, N5629);
buf BUF1 (N6066, N6060);
xor XOR2 (N6067, N6058, N5188);
xor XOR2 (N6068, N6052, N1853);
and AND3 (N6069, N6065, N2154, N1385);
and AND3 (N6070, N6051, N4179, N1470);
buf BUF1 (N6071, N6046);
nand NAND2 (N6072, N6062, N3462);
buf BUF1 (N6073, N6064);
buf BUF1 (N6074, N6069);
or OR2 (N6075, N6049, N3583);
not NOT1 (N6076, N6070);
nor NOR4 (N6077, N6071, N5561, N5723, N2113);
not NOT1 (N6078, N6073);
and AND4 (N6079, N6066, N1387, N3646, N3478);
not NOT1 (N6080, N6068);
xor XOR2 (N6081, N6076, N801);
buf BUF1 (N6082, N6072);
and AND3 (N6083, N6080, N4742, N2265);
buf BUF1 (N6084, N6075);
and AND3 (N6085, N6082, N762, N4598);
xor XOR2 (N6086, N6074, N700);
or OR3 (N6087, N6083, N1217, N1612);
and AND4 (N6088, N6078, N264, N4175, N1385);
nor NOR4 (N6089, N6086, N963, N5510, N2881);
or OR2 (N6090, N6084, N1065);
not NOT1 (N6091, N6088);
nor NOR2 (N6092, N6067, N4173);
nor NOR3 (N6093, N6091, N556, N513);
nor NOR3 (N6094, N6085, N1700, N4242);
or OR2 (N6095, N5986, N3422);
or OR3 (N6096, N6087, N4772, N4299);
or OR3 (N6097, N6096, N2475, N2211);
not NOT1 (N6098, N6079);
and AND2 (N6099, N6089, N3905);
or OR3 (N6100, N6090, N3101, N4814);
nor NOR2 (N6101, N6099, N5715);
nor NOR2 (N6102, N6095, N2178);
buf BUF1 (N6103, N6102);
not NOT1 (N6104, N6103);
and AND4 (N6105, N6092, N1545, N5331, N487);
and AND2 (N6106, N6098, N5174);
nand NAND3 (N6107, N6106, N2677, N3608);
xor XOR2 (N6108, N6100, N1421);
not NOT1 (N6109, N6104);
and AND3 (N6110, N6101, N4468, N5617);
nand NAND2 (N6111, N6093, N1369);
nor NOR3 (N6112, N6097, N2894, N366);
xor XOR2 (N6113, N6077, N3188);
and AND2 (N6114, N6107, N4812);
not NOT1 (N6115, N6081);
or OR3 (N6116, N6109, N5742, N2227);
and AND2 (N6117, N6111, N374);
buf BUF1 (N6118, N6108);
and AND4 (N6119, N6117, N1957, N3625, N5601);
nand NAND3 (N6120, N6105, N4164, N6018);
nor NOR2 (N6121, N6116, N1991);
buf BUF1 (N6122, N6115);
nor NOR2 (N6123, N6121, N4776);
nor NOR3 (N6124, N6120, N3351, N44);
nand NAND2 (N6125, N6123, N3433);
xor XOR2 (N6126, N6124, N4064);
or OR2 (N6127, N6110, N916);
not NOT1 (N6128, N6125);
not NOT1 (N6129, N6118);
nand NAND3 (N6130, N6114, N4149, N2469);
not NOT1 (N6131, N6094);
xor XOR2 (N6132, N6119, N2416);
xor XOR2 (N6133, N6132, N3031);
nor NOR3 (N6134, N6122, N3166, N3147);
not NOT1 (N6135, N6128);
buf BUF1 (N6136, N6126);
xor XOR2 (N6137, N6112, N3876);
not NOT1 (N6138, N6131);
or OR4 (N6139, N6138, N3187, N1636, N4646);
xor XOR2 (N6140, N6113, N5132);
nor NOR4 (N6141, N6127, N4829, N4356, N5480);
nand NAND4 (N6142, N6139, N2454, N1288, N5930);
and AND4 (N6143, N6142, N4141, N5196, N41);
and AND3 (N6144, N6140, N2798, N716);
buf BUF1 (N6145, N6137);
xor XOR2 (N6146, N6134, N5520);
nor NOR2 (N6147, N6133, N5476);
or OR2 (N6148, N6129, N1927);
nand NAND3 (N6149, N6147, N5309, N1735);
not NOT1 (N6150, N6135);
xor XOR2 (N6151, N6136, N3651);
buf BUF1 (N6152, N6151);
and AND2 (N6153, N6141, N2366);
xor XOR2 (N6154, N6145, N1585);
nor NOR3 (N6155, N6150, N918, N2592);
nor NOR2 (N6156, N6154, N5386);
or OR4 (N6157, N6153, N1333, N491, N1260);
not NOT1 (N6158, N6130);
or OR4 (N6159, N6148, N3814, N4794, N4546);
nor NOR3 (N6160, N6152, N5892, N701);
and AND3 (N6161, N6157, N1846, N5566);
not NOT1 (N6162, N6146);
nor NOR3 (N6163, N6155, N5888, N3188);
xor XOR2 (N6164, N6161, N5350);
buf BUF1 (N6165, N6158);
nor NOR2 (N6166, N6159, N2002);
and AND4 (N6167, N6163, N1122, N2354, N2190);
nor NOR4 (N6168, N6162, N727, N3570, N4657);
and AND4 (N6169, N6168, N5905, N3842, N3640);
nor NOR4 (N6170, N6169, N1039, N2404, N1688);
not NOT1 (N6171, N6170);
not NOT1 (N6172, N6143);
and AND2 (N6173, N6167, N4992);
or OR3 (N6174, N6160, N5371, N2000);
nor NOR4 (N6175, N6172, N5503, N1974, N3355);
buf BUF1 (N6176, N6171);
nand NAND3 (N6177, N6156, N3446, N1338);
nand NAND2 (N6178, N6164, N2133);
buf BUF1 (N6179, N6144);
or OR4 (N6180, N6165, N4871, N4702, N3756);
nor NOR2 (N6181, N6178, N578);
xor XOR2 (N6182, N6175, N3724);
xor XOR2 (N6183, N6149, N3343);
not NOT1 (N6184, N6177);
and AND3 (N6185, N6179, N1196, N3538);
xor XOR2 (N6186, N6181, N2541);
nor NOR2 (N6187, N6166, N877);
buf BUF1 (N6188, N6180);
and AND4 (N6189, N6183, N1271, N2639, N4216);
nor NOR3 (N6190, N6173, N2025, N2922);
or OR4 (N6191, N6176, N5944, N5208, N4845);
nor NOR4 (N6192, N6186, N2808, N2413, N2094);
and AND4 (N6193, N6182, N575, N2780, N6043);
nand NAND2 (N6194, N6191, N3601);
nand NAND2 (N6195, N6187, N5967);
xor XOR2 (N6196, N6190, N4897);
nor NOR3 (N6197, N6194, N4010, N4673);
or OR3 (N6198, N6189, N3035, N5284);
and AND2 (N6199, N6195, N3984);
and AND3 (N6200, N6199, N4244, N4726);
nor NOR3 (N6201, N6174, N5922, N637);
nor NOR2 (N6202, N6184, N3110);
and AND4 (N6203, N6202, N5808, N3121, N5820);
xor XOR2 (N6204, N6200, N4492);
and AND4 (N6205, N6203, N1419, N3034, N3626);
not NOT1 (N6206, N6197);
buf BUF1 (N6207, N6205);
and AND3 (N6208, N6185, N1583, N5487);
nor NOR4 (N6209, N6206, N3890, N5011, N4482);
nor NOR2 (N6210, N6193, N3594);
buf BUF1 (N6211, N6209);
buf BUF1 (N6212, N6210);
or OR2 (N6213, N6208, N2350);
nand NAND3 (N6214, N6212, N4754, N1175);
buf BUF1 (N6215, N6211);
and AND4 (N6216, N6214, N3344, N3872, N4567);
or OR2 (N6217, N6207, N1222);
or OR3 (N6218, N6204, N4336, N4005);
xor XOR2 (N6219, N6213, N88);
nand NAND2 (N6220, N6219, N830);
xor XOR2 (N6221, N6217, N1278);
xor XOR2 (N6222, N6192, N420);
nand NAND4 (N6223, N6188, N3639, N4345, N2671);
buf BUF1 (N6224, N6198);
and AND3 (N6225, N6222, N676, N157);
nor NOR3 (N6226, N6223, N591, N4493);
and AND4 (N6227, N6216, N1903, N2682, N2846);
not NOT1 (N6228, N6215);
or OR4 (N6229, N6225, N4361, N6076, N386);
buf BUF1 (N6230, N6226);
and AND4 (N6231, N6228, N6085, N6188, N2527);
and AND2 (N6232, N6229, N5750);
xor XOR2 (N6233, N6230, N731);
nor NOR2 (N6234, N6201, N2605);
buf BUF1 (N6235, N6221);
buf BUF1 (N6236, N6235);
buf BUF1 (N6237, N6234);
not NOT1 (N6238, N6218);
nor NOR2 (N6239, N6220, N4999);
nand NAND3 (N6240, N6196, N148, N6230);
or OR2 (N6241, N6224, N3288);
buf BUF1 (N6242, N6238);
not NOT1 (N6243, N6242);
xor XOR2 (N6244, N6233, N1585);
buf BUF1 (N6245, N6244);
and AND3 (N6246, N6240, N5070, N5216);
or OR4 (N6247, N6231, N820, N3140, N2488);
and AND3 (N6248, N6239, N3087, N442);
xor XOR2 (N6249, N6237, N2813);
and AND2 (N6250, N6232, N5007);
buf BUF1 (N6251, N6249);
and AND2 (N6252, N6250, N1749);
xor XOR2 (N6253, N6248, N5450);
xor XOR2 (N6254, N6246, N4319);
nand NAND3 (N6255, N6227, N501, N3615);
nand NAND3 (N6256, N6241, N2986, N916);
xor XOR2 (N6257, N6245, N1992);
and AND4 (N6258, N6253, N2645, N3007, N1063);
or OR4 (N6259, N6258, N1333, N3363, N1705);
buf BUF1 (N6260, N6256);
nand NAND4 (N6261, N6259, N2629, N370, N1129);
xor XOR2 (N6262, N6236, N5494);
not NOT1 (N6263, N6251);
nor NOR2 (N6264, N6254, N5282);
and AND4 (N6265, N6261, N21, N1704, N4270);
buf BUF1 (N6266, N6265);
nand NAND2 (N6267, N6266, N362);
or OR4 (N6268, N6262, N2830, N4258, N5131);
nand NAND2 (N6269, N6260, N5222);
xor XOR2 (N6270, N6263, N2187);
not NOT1 (N6271, N6252);
nor NOR4 (N6272, N6271, N768, N4742, N358);
and AND2 (N6273, N6255, N4590);
not NOT1 (N6274, N6272);
nor NOR2 (N6275, N6247, N2649);
nand NAND4 (N6276, N6243, N4572, N98, N2569);
nand NAND4 (N6277, N6270, N3105, N5404, N5488);
buf BUF1 (N6278, N6267);
buf BUF1 (N6279, N6269);
nor NOR4 (N6280, N6279, N5718, N1495, N1566);
nand NAND4 (N6281, N6257, N2497, N1757, N530);
not NOT1 (N6282, N6276);
not NOT1 (N6283, N6277);
nor NOR2 (N6284, N6282, N3354);
nor NOR3 (N6285, N6274, N4659, N5206);
buf BUF1 (N6286, N6275);
buf BUF1 (N6287, N6281);
xor XOR2 (N6288, N6283, N3916);
nand NAND4 (N6289, N6268, N1288, N4323, N6059);
not NOT1 (N6290, N6278);
not NOT1 (N6291, N6290);
nand NAND2 (N6292, N6287, N4083);
or OR4 (N6293, N6264, N4545, N2809, N4761);
or OR4 (N6294, N6289, N5418, N3853, N2659);
nor NOR2 (N6295, N6288, N3324);
and AND2 (N6296, N6294, N5784);
not NOT1 (N6297, N6291);
buf BUF1 (N6298, N6273);
nor NOR3 (N6299, N6286, N4309, N2001);
nand NAND4 (N6300, N6299, N4040, N2405, N2710);
nor NOR2 (N6301, N6292, N5963);
not NOT1 (N6302, N6293);
not NOT1 (N6303, N6280);
buf BUF1 (N6304, N6298);
nand NAND2 (N6305, N6303, N136);
buf BUF1 (N6306, N6301);
xor XOR2 (N6307, N6296, N885);
and AND4 (N6308, N6304, N1022, N939, N5466);
and AND2 (N6309, N6284, N1300);
nor NOR2 (N6310, N6285, N3781);
or OR2 (N6311, N6300, N4827);
xor XOR2 (N6312, N6308, N3858);
nand NAND4 (N6313, N6297, N5051, N1849, N512);
or OR2 (N6314, N6302, N3479);
buf BUF1 (N6315, N6309);
xor XOR2 (N6316, N6313, N67);
buf BUF1 (N6317, N6312);
or OR4 (N6318, N6305, N843, N5108, N3839);
not NOT1 (N6319, N6318);
nor NOR4 (N6320, N6310, N2757, N5508, N4807);
nand NAND3 (N6321, N6315, N2231, N2993);
nand NAND4 (N6322, N6319, N4013, N3865, N3313);
or OR2 (N6323, N6321, N823);
not NOT1 (N6324, N6320);
or OR3 (N6325, N6323, N3156, N3124);
or OR2 (N6326, N6316, N5299);
nor NOR4 (N6327, N6324, N4908, N467, N3391);
buf BUF1 (N6328, N6327);
nand NAND4 (N6329, N6314, N4777, N18, N5912);
and AND2 (N6330, N6311, N4056);
not NOT1 (N6331, N6330);
nand NAND2 (N6332, N6326, N695);
and AND4 (N6333, N6332, N1750, N717, N1879);
buf BUF1 (N6334, N6325);
or OR3 (N6335, N6307, N2920, N4732);
nor NOR4 (N6336, N6317, N4701, N4360, N2362);
buf BUF1 (N6337, N6329);
nor NOR2 (N6338, N6331, N4256);
and AND2 (N6339, N6322, N5217);
nand NAND3 (N6340, N6328, N5413, N5844);
and AND4 (N6341, N6335, N6034, N4576, N1927);
and AND3 (N6342, N6341, N1935, N4769);
buf BUF1 (N6343, N6295);
xor XOR2 (N6344, N6338, N231);
not NOT1 (N6345, N6333);
and AND4 (N6346, N6344, N2574, N1535, N3274);
or OR4 (N6347, N6337, N3963, N5763, N1);
not NOT1 (N6348, N6334);
xor XOR2 (N6349, N6336, N1257);
not NOT1 (N6350, N6306);
buf BUF1 (N6351, N6349);
nand NAND2 (N6352, N6350, N1199);
buf BUF1 (N6353, N6347);
not NOT1 (N6354, N6342);
buf BUF1 (N6355, N6354);
not NOT1 (N6356, N6353);
and AND3 (N6357, N6348, N3247, N3203);
xor XOR2 (N6358, N6339, N3630);
buf BUF1 (N6359, N6346);
or OR2 (N6360, N6351, N4902);
or OR3 (N6361, N6355, N3041, N5168);
not NOT1 (N6362, N6358);
and AND2 (N6363, N6340, N1334);
nor NOR3 (N6364, N6357, N2021, N4658);
or OR4 (N6365, N6352, N2987, N5427, N5921);
or OR3 (N6366, N6345, N3819, N863);
and AND3 (N6367, N6359, N1657, N332);
xor XOR2 (N6368, N6365, N5189);
or OR2 (N6369, N6366, N3454);
buf BUF1 (N6370, N6368);
xor XOR2 (N6371, N6363, N2541);
buf BUF1 (N6372, N6360);
nand NAND2 (N6373, N6364, N2672);
buf BUF1 (N6374, N6361);
nand NAND2 (N6375, N6374, N1039);
not NOT1 (N6376, N6371);
xor XOR2 (N6377, N6343, N4110);
nand NAND4 (N6378, N6369, N6080, N2169, N1692);
xor XOR2 (N6379, N6370, N1528);
nand NAND4 (N6380, N6376, N112, N1170, N4795);
buf BUF1 (N6381, N6367);
nor NOR3 (N6382, N6362, N5410, N1568);
and AND2 (N6383, N6379, N5189);
nor NOR2 (N6384, N6375, N1786);
xor XOR2 (N6385, N6383, N3734);
or OR4 (N6386, N6380, N6035, N423, N5544);
or OR3 (N6387, N6381, N151, N3198);
or OR4 (N6388, N6372, N1754, N3868, N1485);
and AND4 (N6389, N6378, N4959, N5677, N252);
not NOT1 (N6390, N6388);
buf BUF1 (N6391, N6356);
nand NAND2 (N6392, N6386, N3471);
or OR4 (N6393, N6382, N4521, N5192, N6286);
and AND2 (N6394, N6390, N1545);
buf BUF1 (N6395, N6394);
xor XOR2 (N6396, N6393, N297);
and AND4 (N6397, N6392, N5500, N1936, N804);
nand NAND3 (N6398, N6373, N168, N2454);
or OR2 (N6399, N6397, N6290);
buf BUF1 (N6400, N6377);
xor XOR2 (N6401, N6396, N79);
nand NAND3 (N6402, N6395, N3906, N2921);
or OR3 (N6403, N6402, N4581, N814);
and AND2 (N6404, N6387, N1567);
nand NAND2 (N6405, N6384, N1715);
not NOT1 (N6406, N6385);
xor XOR2 (N6407, N6401, N6292);
and AND4 (N6408, N6398, N3187, N906, N466);
or OR4 (N6409, N6408, N3944, N1008, N3333);
xor XOR2 (N6410, N6403, N1999);
nand NAND2 (N6411, N6391, N6204);
not NOT1 (N6412, N6406);
nor NOR3 (N6413, N6404, N4791, N2440);
xor XOR2 (N6414, N6412, N3889);
and AND3 (N6415, N6413, N2917, N5279);
and AND3 (N6416, N6411, N3138, N4516);
not NOT1 (N6417, N6399);
not NOT1 (N6418, N6409);
xor XOR2 (N6419, N6417, N4295);
xor XOR2 (N6420, N6416, N1961);
not NOT1 (N6421, N6400);
or OR2 (N6422, N6405, N907);
xor XOR2 (N6423, N6410, N4344);
not NOT1 (N6424, N6415);
or OR4 (N6425, N6423, N1018, N4145, N4825);
nand NAND4 (N6426, N6422, N5703, N1933, N2426);
buf BUF1 (N6427, N6419);
nand NAND4 (N6428, N6418, N5681, N1985, N1387);
nand NAND3 (N6429, N6389, N4153, N1046);
nor NOR4 (N6430, N6425, N2697, N2340, N5947);
nand NAND3 (N6431, N6427, N2495, N2093);
nand NAND2 (N6432, N6428, N1635);
xor XOR2 (N6433, N6430, N2613);
buf BUF1 (N6434, N6426);
buf BUF1 (N6435, N6429);
xor XOR2 (N6436, N6433, N3250);
xor XOR2 (N6437, N6414, N3300);
not NOT1 (N6438, N6421);
nor NOR3 (N6439, N6436, N6246, N5567);
buf BUF1 (N6440, N6407);
not NOT1 (N6441, N6437);
and AND2 (N6442, N6439, N4374);
xor XOR2 (N6443, N6438, N4066);
buf BUF1 (N6444, N6432);
nand NAND3 (N6445, N6434, N3265, N848);
not NOT1 (N6446, N6444);
nor NOR2 (N6447, N6420, N5149);
or OR4 (N6448, N6424, N5749, N3776, N679);
nor NOR3 (N6449, N6445, N1003, N1234);
or OR3 (N6450, N6446, N414, N1211);
xor XOR2 (N6451, N6440, N5472);
nor NOR2 (N6452, N6431, N3857);
and AND3 (N6453, N6441, N2201, N2542);
nand NAND2 (N6454, N6447, N3526);
buf BUF1 (N6455, N6450);
buf BUF1 (N6456, N6442);
nand NAND2 (N6457, N6456, N6194);
and AND3 (N6458, N6454, N324, N1425);
xor XOR2 (N6459, N6448, N1464);
not NOT1 (N6460, N6457);
buf BUF1 (N6461, N6458);
and AND2 (N6462, N6443, N5677);
xor XOR2 (N6463, N6462, N2001);
not NOT1 (N6464, N6452);
xor XOR2 (N6465, N6461, N1451);
not NOT1 (N6466, N6455);
not NOT1 (N6467, N6459);
buf BUF1 (N6468, N6435);
or OR2 (N6469, N6451, N4412);
nor NOR4 (N6470, N6467, N4656, N1276, N4256);
buf BUF1 (N6471, N6468);
not NOT1 (N6472, N6469);
buf BUF1 (N6473, N6449);
xor XOR2 (N6474, N6471, N4247);
and AND3 (N6475, N6470, N2931, N5924);
xor XOR2 (N6476, N6472, N3092);
buf BUF1 (N6477, N6476);
or OR4 (N6478, N6475, N6109, N3856, N3340);
and AND3 (N6479, N6478, N4974, N4026);
nor NOR4 (N6480, N6464, N1667, N2701, N4978);
nand NAND2 (N6481, N6453, N2137);
xor XOR2 (N6482, N6480, N4251);
buf BUF1 (N6483, N6479);
not NOT1 (N6484, N6474);
or OR4 (N6485, N6483, N2630, N4594, N5220);
and AND4 (N6486, N6465, N6267, N908, N4455);
or OR4 (N6487, N6485, N2372, N853, N4961);
not NOT1 (N6488, N6460);
nand NAND2 (N6489, N6488, N1516);
buf BUF1 (N6490, N6482);
or OR3 (N6491, N6473, N4824, N4515);
nand NAND4 (N6492, N6477, N795, N2307, N5808);
not NOT1 (N6493, N6481);
not NOT1 (N6494, N6490);
nand NAND3 (N6495, N6492, N686, N1275);
or OR3 (N6496, N6495, N5054, N2534);
buf BUF1 (N6497, N6489);
and AND3 (N6498, N6466, N85, N2714);
xor XOR2 (N6499, N6486, N2287);
or OR4 (N6500, N6484, N4876, N5035, N5199);
buf BUF1 (N6501, N6493);
buf BUF1 (N6502, N6487);
nand NAND3 (N6503, N6497, N2886, N948);
nor NOR2 (N6504, N6499, N4402);
buf BUF1 (N6505, N6501);
nor NOR3 (N6506, N6463, N2824, N4056);
and AND4 (N6507, N6500, N2954, N1495, N5598);
or OR3 (N6508, N6502, N673, N4510);
and AND4 (N6509, N6507, N4761, N806, N2166);
and AND4 (N6510, N6506, N2137, N553, N5929);
nand NAND3 (N6511, N6498, N932, N274);
or OR2 (N6512, N6511, N613);
nand NAND3 (N6513, N6508, N531, N372);
nor NOR2 (N6514, N6509, N4684);
nor NOR2 (N6515, N6510, N2416);
or OR3 (N6516, N6503, N2168, N2589);
nand NAND2 (N6517, N6516, N5939);
not NOT1 (N6518, N6515);
xor XOR2 (N6519, N6496, N166);
xor XOR2 (N6520, N6504, N3148);
buf BUF1 (N6521, N6514);
and AND4 (N6522, N6505, N150, N4710, N1845);
nor NOR2 (N6523, N6491, N4117);
nor NOR2 (N6524, N6520, N1110);
nand NAND4 (N6525, N6518, N436, N3376, N5578);
not NOT1 (N6526, N6512);
nor NOR3 (N6527, N6522, N4260, N2568);
or OR4 (N6528, N6519, N1747, N6263, N1308);
nor NOR2 (N6529, N6521, N4269);
or OR4 (N6530, N6517, N347, N3892, N86);
and AND4 (N6531, N6524, N935, N5644, N4260);
not NOT1 (N6532, N6513);
nand NAND4 (N6533, N6528, N2008, N3001, N3568);
and AND4 (N6534, N6527, N2068, N4646, N1374);
xor XOR2 (N6535, N6523, N1427);
xor XOR2 (N6536, N6531, N5581);
not NOT1 (N6537, N6534);
nand NAND3 (N6538, N6536, N3817, N48);
buf BUF1 (N6539, N6525);
or OR4 (N6540, N6529, N2183, N5801, N616);
xor XOR2 (N6541, N6530, N2033);
nand NAND2 (N6542, N6539, N3450);
and AND4 (N6543, N6538, N332, N6523, N933);
nor NOR2 (N6544, N6532, N5373);
not NOT1 (N6545, N6541);
nor NOR2 (N6546, N6545, N4653);
not NOT1 (N6547, N6494);
buf BUF1 (N6548, N6540);
xor XOR2 (N6549, N6526, N5507);
or OR4 (N6550, N6533, N1058, N6306, N4792);
nand NAND4 (N6551, N6548, N2859, N4098, N1168);
not NOT1 (N6552, N6543);
or OR2 (N6553, N6542, N1084);
xor XOR2 (N6554, N6549, N4510);
nand NAND3 (N6555, N6537, N328, N4428);
buf BUF1 (N6556, N6535);
buf BUF1 (N6557, N6555);
nand NAND4 (N6558, N6556, N6058, N4527, N2621);
xor XOR2 (N6559, N6544, N2536);
xor XOR2 (N6560, N6551, N4801);
xor XOR2 (N6561, N6554, N5995);
or OR2 (N6562, N6560, N6054);
nand NAND2 (N6563, N6562, N5720);
buf BUF1 (N6564, N6547);
or OR4 (N6565, N6561, N1673, N103, N4509);
or OR3 (N6566, N6553, N3501, N2351);
xor XOR2 (N6567, N6558, N4252);
xor XOR2 (N6568, N6567, N4862);
nor NOR3 (N6569, N6552, N2570, N3927);
xor XOR2 (N6570, N6568, N420);
and AND4 (N6571, N6563, N1595, N5743, N5322);
not NOT1 (N6572, N6559);
not NOT1 (N6573, N6569);
nor NOR3 (N6574, N6566, N1107, N190);
nor NOR2 (N6575, N6570, N2555);
xor XOR2 (N6576, N6574, N1773);
or OR3 (N6577, N6564, N2616, N2131);
xor XOR2 (N6578, N6571, N6495);
buf BUF1 (N6579, N6546);
nand NAND2 (N6580, N6573, N178);
nor NOR4 (N6581, N6557, N2976, N5624, N3523);
nand NAND2 (N6582, N6550, N4451);
nand NAND2 (N6583, N6579, N3489);
not NOT1 (N6584, N6583);
not NOT1 (N6585, N6581);
nor NOR4 (N6586, N6585, N3414, N6575, N5522);
or OR3 (N6587, N1296, N875, N6052);
xor XOR2 (N6588, N6587, N3632);
buf BUF1 (N6589, N6577);
or OR4 (N6590, N6588, N1850, N3186, N4925);
not NOT1 (N6591, N6582);
or OR3 (N6592, N6589, N6530, N2141);
not NOT1 (N6593, N6576);
or OR2 (N6594, N6584, N4561);
or OR4 (N6595, N6586, N4870, N278, N4213);
buf BUF1 (N6596, N6591);
or OR4 (N6597, N6578, N4202, N4515, N5060);
and AND2 (N6598, N6594, N1826);
buf BUF1 (N6599, N6596);
and AND4 (N6600, N6592, N4562, N2756, N6050);
buf BUF1 (N6601, N6580);
nor NOR4 (N6602, N6595, N2127, N3425, N5389);
nor NOR4 (N6603, N6565, N2495, N4077, N730);
nor NOR4 (N6604, N6599, N439, N255, N5417);
buf BUF1 (N6605, N6600);
not NOT1 (N6606, N6572);
and AND3 (N6607, N6604, N6582, N2400);
nor NOR3 (N6608, N6606, N2369, N3927);
nor NOR4 (N6609, N6607, N1704, N5082, N6134);
and AND2 (N6610, N6603, N5376);
or OR3 (N6611, N6610, N6320, N6337);
xor XOR2 (N6612, N6602, N5497);
and AND3 (N6613, N6609, N5755, N2665);
nand NAND4 (N6614, N6597, N3029, N3040, N6436);
nor NOR4 (N6615, N6614, N1877, N1193, N6487);
and AND3 (N6616, N6593, N2218, N4933);
xor XOR2 (N6617, N6601, N1449);
xor XOR2 (N6618, N6608, N4510);
or OR4 (N6619, N6618, N3336, N1005, N5946);
not NOT1 (N6620, N6613);
xor XOR2 (N6621, N6598, N2482);
xor XOR2 (N6622, N6590, N5948);
nand NAND2 (N6623, N6615, N6038);
xor XOR2 (N6624, N6616, N3672);
xor XOR2 (N6625, N6624, N2060);
or OR3 (N6626, N6625, N2632, N6111);
not NOT1 (N6627, N6619);
xor XOR2 (N6628, N6627, N484);
nor NOR2 (N6629, N6617, N5099);
xor XOR2 (N6630, N6626, N2638);
or OR2 (N6631, N6611, N3580);
buf BUF1 (N6632, N6629);
buf BUF1 (N6633, N6621);
nor NOR3 (N6634, N6628, N2598, N5404);
nor NOR2 (N6635, N6623, N976);
xor XOR2 (N6636, N6622, N6603);
xor XOR2 (N6637, N6632, N4075);
nand NAND2 (N6638, N6620, N3181);
buf BUF1 (N6639, N6633);
nor NOR3 (N6640, N6605, N6364, N834);
buf BUF1 (N6641, N6640);
buf BUF1 (N6642, N6635);
xor XOR2 (N6643, N6612, N6506);
buf BUF1 (N6644, N6643);
or OR3 (N6645, N6642, N5739, N5741);
buf BUF1 (N6646, N6638);
or OR4 (N6647, N6630, N5728, N1697, N134);
or OR2 (N6648, N6646, N6631);
nor NOR4 (N6649, N3612, N4253, N3751, N3427);
not NOT1 (N6650, N6641);
and AND3 (N6651, N6636, N2566, N745);
xor XOR2 (N6652, N6647, N101);
not NOT1 (N6653, N6651);
buf BUF1 (N6654, N6650);
nor NOR4 (N6655, N6648, N4048, N2108, N231);
nand NAND4 (N6656, N6652, N1562, N2905, N3527);
and AND4 (N6657, N6634, N102, N4446, N5533);
xor XOR2 (N6658, N6639, N5106);
nor NOR4 (N6659, N6656, N6477, N2164, N4291);
or OR4 (N6660, N6659, N5165, N4268, N2837);
nor NOR4 (N6661, N6644, N569, N3308, N5531);
xor XOR2 (N6662, N6658, N3323);
buf BUF1 (N6663, N6645);
xor XOR2 (N6664, N6655, N4637);
and AND4 (N6665, N6649, N2697, N5124, N4015);
buf BUF1 (N6666, N6665);
or OR4 (N6667, N6666, N2740, N567, N1207);
xor XOR2 (N6668, N6654, N215);
nand NAND3 (N6669, N6667, N1541, N3059);
or OR3 (N6670, N6669, N2781, N4201);
buf BUF1 (N6671, N6670);
nor NOR3 (N6672, N6653, N1573, N6318);
and AND2 (N6673, N6660, N1477);
and AND3 (N6674, N6673, N4464, N1014);
buf BUF1 (N6675, N6662);
and AND3 (N6676, N6674, N2027, N3591);
nor NOR3 (N6677, N6661, N794, N4154);
and AND2 (N6678, N6657, N248);
xor XOR2 (N6679, N6677, N635);
xor XOR2 (N6680, N6671, N746);
or OR3 (N6681, N6678, N6204, N1414);
or OR3 (N6682, N6672, N4570, N1517);
or OR4 (N6683, N6681, N1204, N4958, N3042);
or OR3 (N6684, N6676, N3364, N3905);
nand NAND4 (N6685, N6682, N218, N1038, N6455);
xor XOR2 (N6686, N6679, N2951);
buf BUF1 (N6687, N6637);
buf BUF1 (N6688, N6684);
buf BUF1 (N6689, N6683);
xor XOR2 (N6690, N6685, N6232);
buf BUF1 (N6691, N6689);
nand NAND2 (N6692, N6687, N3889);
and AND2 (N6693, N6663, N4498);
nand NAND4 (N6694, N6680, N6245, N3940, N3688);
or OR3 (N6695, N6664, N5013, N4080);
buf BUF1 (N6696, N6690);
nand NAND4 (N6697, N6692, N194, N4307, N2526);
and AND4 (N6698, N6693, N1179, N1886, N2331);
not NOT1 (N6699, N6686);
xor XOR2 (N6700, N6675, N1021);
not NOT1 (N6701, N6696);
and AND4 (N6702, N6700, N5007, N5106, N1847);
nand NAND4 (N6703, N6688, N5325, N6323, N2731);
and AND2 (N6704, N6691, N2936);
nor NOR3 (N6705, N6694, N452, N4466);
not NOT1 (N6706, N6699);
buf BUF1 (N6707, N6701);
and AND4 (N6708, N6668, N917, N3225, N5719);
buf BUF1 (N6709, N6706);
nor NOR3 (N6710, N6698, N1825, N406);
xor XOR2 (N6711, N6703, N1908);
xor XOR2 (N6712, N6704, N2525);
xor XOR2 (N6713, N6705, N6547);
or OR3 (N6714, N6708, N1288, N6060);
buf BUF1 (N6715, N6710);
buf BUF1 (N6716, N6707);
xor XOR2 (N6717, N6715, N4759);
or OR3 (N6718, N6717, N3799, N1481);
nand NAND4 (N6719, N6713, N4782, N4696, N6107);
buf BUF1 (N6720, N6712);
and AND3 (N6721, N6709, N4370, N3608);
buf BUF1 (N6722, N6702);
buf BUF1 (N6723, N6721);
or OR2 (N6724, N6714, N6055);
buf BUF1 (N6725, N6720);
nor NOR2 (N6726, N6711, N548);
nand NAND3 (N6727, N6723, N3211, N5597);
and AND4 (N6728, N6719, N5564, N2578, N2504);
and AND3 (N6729, N6716, N4531, N686);
xor XOR2 (N6730, N6722, N1809);
buf BUF1 (N6731, N6718);
nor NOR2 (N6732, N6695, N6249);
or OR4 (N6733, N6731, N1701, N3822, N4502);
buf BUF1 (N6734, N6726);
xor XOR2 (N6735, N6734, N6674);
or OR2 (N6736, N6727, N4774);
buf BUF1 (N6737, N6729);
not NOT1 (N6738, N6697);
not NOT1 (N6739, N6732);
or OR4 (N6740, N6724, N4604, N3550, N2229);
or OR4 (N6741, N6737, N2112, N5689, N5519);
nand NAND4 (N6742, N6730, N5699, N2780, N2397);
not NOT1 (N6743, N6739);
buf BUF1 (N6744, N6738);
not NOT1 (N6745, N6735);
buf BUF1 (N6746, N6725);
not NOT1 (N6747, N6743);
and AND2 (N6748, N6736, N2137);
nor NOR3 (N6749, N6742, N5138, N409);
xor XOR2 (N6750, N6740, N2229);
nor NOR4 (N6751, N6745, N660, N3459, N3420);
and AND4 (N6752, N6746, N1195, N3993, N1098);
nand NAND2 (N6753, N6741, N5939);
nand NAND2 (N6754, N6728, N2726);
nor NOR2 (N6755, N6753, N442);
nor NOR3 (N6756, N6747, N5445, N6545);
nor NOR3 (N6757, N6733, N1915, N4015);
nor NOR4 (N6758, N6757, N5651, N2489, N2514);
nand NAND3 (N6759, N6751, N2045, N927);
buf BUF1 (N6760, N6750);
or OR2 (N6761, N6749, N3517);
nor NOR2 (N6762, N6755, N3044);
and AND4 (N6763, N6754, N4326, N5590, N4836);
not NOT1 (N6764, N6744);
xor XOR2 (N6765, N6756, N3479);
not NOT1 (N6766, N6765);
nand NAND4 (N6767, N6766, N4063, N5712, N705);
buf BUF1 (N6768, N6752);
or OR4 (N6769, N6759, N4269, N1584, N5385);
or OR3 (N6770, N6761, N2254, N3335);
and AND2 (N6771, N6763, N3500);
xor XOR2 (N6772, N6770, N676);
nor NOR2 (N6773, N6760, N566);
buf BUF1 (N6774, N6764);
not NOT1 (N6775, N6767);
nor NOR2 (N6776, N6769, N6756);
or OR4 (N6777, N6772, N5399, N6691, N5395);
or OR2 (N6778, N6768, N6258);
not NOT1 (N6779, N6775);
nand NAND3 (N6780, N6774, N4366, N6483);
nor NOR4 (N6781, N6748, N1433, N1213, N6274);
not NOT1 (N6782, N6771);
nand NAND4 (N6783, N6758, N5021, N30, N1327);
or OR4 (N6784, N6777, N4314, N2688, N4187);
and AND3 (N6785, N6781, N3317, N120);
not NOT1 (N6786, N6778);
nor NOR4 (N6787, N6776, N1746, N1108, N2363);
xor XOR2 (N6788, N6779, N6720);
nor NOR3 (N6789, N6784, N3244, N6305);
or OR4 (N6790, N6780, N2999, N887, N3319);
buf BUF1 (N6791, N6762);
nor NOR4 (N6792, N6785, N1137, N1338, N4965);
and AND2 (N6793, N6782, N700);
nand NAND3 (N6794, N6793, N6161, N3261);
nand NAND3 (N6795, N6789, N2029, N6090);
not NOT1 (N6796, N6773);
nor NOR2 (N6797, N6796, N774);
and AND3 (N6798, N6786, N3581, N3324);
nor NOR2 (N6799, N6798, N327);
and AND2 (N6800, N6790, N3041);
buf BUF1 (N6801, N6800);
nand NAND4 (N6802, N6797, N2735, N6315, N3812);
not NOT1 (N6803, N6788);
not NOT1 (N6804, N6803);
not NOT1 (N6805, N6799);
nor NOR2 (N6806, N6795, N1462);
not NOT1 (N6807, N6804);
nor NOR2 (N6808, N6794, N1760);
not NOT1 (N6809, N6806);
buf BUF1 (N6810, N6801);
nor NOR2 (N6811, N6802, N203);
not NOT1 (N6812, N6787);
buf BUF1 (N6813, N6810);
xor XOR2 (N6814, N6783, N3262);
xor XOR2 (N6815, N6814, N5388);
not NOT1 (N6816, N6811);
and AND3 (N6817, N6815, N521, N3742);
nor NOR3 (N6818, N6805, N5323, N3818);
nand NAND4 (N6819, N6813, N3032, N1527, N2461);
buf BUF1 (N6820, N6791);
or OR3 (N6821, N6817, N4092, N5930);
or OR2 (N6822, N6819, N822);
and AND3 (N6823, N6809, N6388, N6001);
not NOT1 (N6824, N6818);
nand NAND2 (N6825, N6824, N1708);
or OR2 (N6826, N6823, N4032);
nor NOR2 (N6827, N6826, N3792);
xor XOR2 (N6828, N6822, N294);
xor XOR2 (N6829, N6825, N758);
buf BUF1 (N6830, N6829);
and AND2 (N6831, N6820, N3778);
buf BUF1 (N6832, N6828);
and AND4 (N6833, N6816, N3409, N2212, N2053);
or OR2 (N6834, N6832, N2918);
or OR2 (N6835, N6833, N2778);
and AND4 (N6836, N6792, N2581, N1295, N110);
or OR4 (N6837, N6834, N6365, N6379, N2098);
nand NAND2 (N6838, N6808, N4548);
or OR3 (N6839, N6837, N3294, N5712);
nor NOR3 (N6840, N6821, N917, N5135);
xor XOR2 (N6841, N6840, N3516);
nor NOR4 (N6842, N6807, N5449, N3984, N2032);
xor XOR2 (N6843, N6831, N440);
nor NOR4 (N6844, N6835, N5249, N1977, N3036);
and AND2 (N6845, N6830, N339);
or OR3 (N6846, N6845, N6358, N5165);
and AND3 (N6847, N6827, N3597, N1903);
xor XOR2 (N6848, N6844, N313);
not NOT1 (N6849, N6838);
and AND2 (N6850, N6839, N5555);
and AND4 (N6851, N6846, N5673, N4722, N3310);
nor NOR2 (N6852, N6850, N6747);
nand NAND3 (N6853, N6812, N4204, N4196);
xor XOR2 (N6854, N6849, N4027);
nor NOR4 (N6855, N6852, N1220, N414, N505);
not NOT1 (N6856, N6855);
not NOT1 (N6857, N6848);
nand NAND2 (N6858, N6854, N5682);
or OR4 (N6859, N6851, N4728, N2660, N2689);
and AND3 (N6860, N6836, N6689, N5209);
buf BUF1 (N6861, N6856);
or OR3 (N6862, N6853, N1667, N5100);
and AND2 (N6863, N6841, N261);
or OR3 (N6864, N6842, N4535, N1744);
and AND4 (N6865, N6857, N3788, N5680, N4956);
nand NAND3 (N6866, N6865, N3986, N6779);
xor XOR2 (N6867, N6858, N5255);
not NOT1 (N6868, N6847);
buf BUF1 (N6869, N6861);
or OR4 (N6870, N6864, N711, N4590, N6424);
and AND2 (N6871, N6869, N1317);
buf BUF1 (N6872, N6843);
xor XOR2 (N6873, N6866, N2629);
nand NAND4 (N6874, N6870, N4231, N1558, N3375);
or OR2 (N6875, N6863, N3164);
not NOT1 (N6876, N6867);
or OR2 (N6877, N6874, N4993);
xor XOR2 (N6878, N6873, N2033);
or OR4 (N6879, N6876, N361, N1994, N3348);
and AND2 (N6880, N6871, N723);
xor XOR2 (N6881, N6880, N2217);
and AND2 (N6882, N6877, N4550);
xor XOR2 (N6883, N6878, N5074);
nor NOR4 (N6884, N6879, N3240, N525, N5379);
or OR2 (N6885, N6859, N4234);
not NOT1 (N6886, N6872);
nor NOR4 (N6887, N6882, N4373, N4896, N4562);
nor NOR4 (N6888, N6883, N4497, N3463, N6445);
buf BUF1 (N6889, N6888);
or OR4 (N6890, N6886, N138, N1057, N3954);
nor NOR3 (N6891, N6881, N1140, N101);
not NOT1 (N6892, N6889);
nand NAND4 (N6893, N6891, N3568, N3892, N2938);
nor NOR2 (N6894, N6887, N2549);
buf BUF1 (N6895, N6868);
xor XOR2 (N6896, N6892, N1896);
or OR2 (N6897, N6862, N330);
xor XOR2 (N6898, N6894, N2569);
buf BUF1 (N6899, N6896);
xor XOR2 (N6900, N6884, N5116);
xor XOR2 (N6901, N6890, N292);
and AND2 (N6902, N6875, N3985);
xor XOR2 (N6903, N6901, N630);
and AND4 (N6904, N6899, N2493, N202, N1548);
nor NOR3 (N6905, N6897, N5594, N5415);
buf BUF1 (N6906, N6905);
xor XOR2 (N6907, N6904, N373);
not NOT1 (N6908, N6900);
xor XOR2 (N6909, N6903, N750);
and AND3 (N6910, N6885, N1243, N1172);
nand NAND2 (N6911, N6898, N4596);
xor XOR2 (N6912, N6902, N3948);
xor XOR2 (N6913, N6893, N3672);
or OR2 (N6914, N6909, N1236);
buf BUF1 (N6915, N6907);
nand NAND4 (N6916, N6895, N5317, N3072, N3509);
nor NOR3 (N6917, N6914, N3525, N6497);
or OR3 (N6918, N6906, N4512, N3172);
buf BUF1 (N6919, N6910);
buf BUF1 (N6920, N6911);
not NOT1 (N6921, N6860);
and AND3 (N6922, N6915, N2680, N1511);
and AND2 (N6923, N6922, N6864);
nor NOR4 (N6924, N6921, N4351, N2562, N1827);
xor XOR2 (N6925, N6923, N1478);
xor XOR2 (N6926, N6925, N2411);
or OR2 (N6927, N6918, N4713);
nand NAND4 (N6928, N6908, N4027, N2261, N3608);
not NOT1 (N6929, N6926);
buf BUF1 (N6930, N6927);
nand NAND2 (N6931, N6929, N3226);
xor XOR2 (N6932, N6931, N6113);
nand NAND2 (N6933, N6920, N541);
nor NOR4 (N6934, N6928, N2683, N836, N6824);
nand NAND3 (N6935, N6912, N6557, N1980);
buf BUF1 (N6936, N6935);
or OR3 (N6937, N6917, N6574, N1374);
not NOT1 (N6938, N6933);
not NOT1 (N6939, N6932);
xor XOR2 (N6940, N6938, N889);
and AND4 (N6941, N6919, N36, N5456, N2129);
buf BUF1 (N6942, N6934);
and AND2 (N6943, N6916, N4966);
xor XOR2 (N6944, N6937, N5047);
or OR4 (N6945, N6936, N2964, N3898, N1389);
not NOT1 (N6946, N6924);
and AND3 (N6947, N6945, N3749, N5265);
nor NOR4 (N6948, N6930, N4646, N2429, N6904);
or OR4 (N6949, N6947, N2552, N6812, N2970);
xor XOR2 (N6950, N6941, N6584);
or OR2 (N6951, N6940, N1559);
and AND2 (N6952, N6950, N2512);
xor XOR2 (N6953, N6948, N1156);
nand NAND2 (N6954, N6952, N2046);
or OR2 (N6955, N6953, N6420);
nand NAND4 (N6956, N6946, N1244, N2930, N2478);
nor NOR3 (N6957, N6956, N4603, N1034);
not NOT1 (N6958, N6949);
nor NOR2 (N6959, N6942, N2440);
or OR4 (N6960, N6951, N4692, N421, N4779);
not NOT1 (N6961, N6954);
or OR3 (N6962, N6943, N4260, N3821);
not NOT1 (N6963, N6955);
and AND3 (N6964, N6963, N5073, N132);
xor XOR2 (N6965, N6961, N5428);
nand NAND4 (N6966, N6958, N935, N5711, N3465);
not NOT1 (N6967, N6964);
nor NOR3 (N6968, N6944, N4674, N5811);
nand NAND4 (N6969, N6967, N2930, N5873, N4444);
or OR3 (N6970, N6969, N1017, N1274);
nand NAND3 (N6971, N6939, N5506, N4695);
and AND3 (N6972, N6965, N3601, N2989);
nand NAND2 (N6973, N6966, N2853);
nand NAND4 (N6974, N6960, N3649, N393, N2265);
or OR3 (N6975, N6974, N2725, N6331);
not NOT1 (N6976, N6971);
not NOT1 (N6977, N6957);
nand NAND4 (N6978, N6973, N2071, N3297, N4118);
and AND4 (N6979, N6975, N1698, N5601, N942);
nand NAND2 (N6980, N6978, N3892);
nor NOR3 (N6981, N6959, N1169, N856);
buf BUF1 (N6982, N6981);
and AND2 (N6983, N6972, N5424);
xor XOR2 (N6984, N6976, N5648);
xor XOR2 (N6985, N6979, N2173);
nor NOR4 (N6986, N6977, N4504, N1632, N5309);
not NOT1 (N6987, N6980);
nand NAND3 (N6988, N6913, N684, N503);
and AND3 (N6989, N6983, N2214, N4965);
xor XOR2 (N6990, N6985, N4130);
xor XOR2 (N6991, N6986, N4002);
not NOT1 (N6992, N6982);
nand NAND2 (N6993, N6970, N3698);
or OR2 (N6994, N6989, N3493);
xor XOR2 (N6995, N6992, N2165);
xor XOR2 (N6996, N6990, N2898);
xor XOR2 (N6997, N6994, N2488);
or OR4 (N6998, N6984, N551, N5137, N514);
or OR4 (N6999, N6991, N73, N1853, N462);
and AND2 (N7000, N6968, N6107);
buf BUF1 (N7001, N6997);
not NOT1 (N7002, N6987);
xor XOR2 (N7003, N6995, N2310);
nand NAND2 (N7004, N6993, N1718);
not NOT1 (N7005, N6998);
xor XOR2 (N7006, N7000, N1111);
buf BUF1 (N7007, N7002);
buf BUF1 (N7008, N7007);
buf BUF1 (N7009, N7004);
or OR2 (N7010, N7003, N3466);
nor NOR2 (N7011, N6996, N5413);
xor XOR2 (N7012, N7010, N2711);
and AND4 (N7013, N7009, N379, N710, N2185);
nand NAND3 (N7014, N6999, N1257, N6888);
nand NAND2 (N7015, N6962, N6178);
nand NAND3 (N7016, N7015, N6817, N6716);
buf BUF1 (N7017, N7011);
xor XOR2 (N7018, N7005, N6839);
and AND3 (N7019, N7018, N3010, N2426);
or OR4 (N7020, N6988, N2698, N2025, N849);
xor XOR2 (N7021, N7017, N5488);
xor XOR2 (N7022, N7019, N1681);
buf BUF1 (N7023, N7021);
xor XOR2 (N7024, N7006, N4492);
nor NOR2 (N7025, N7020, N468);
nand NAND3 (N7026, N7001, N5609, N2242);
buf BUF1 (N7027, N7013);
or OR4 (N7028, N7008, N6499, N6580, N1610);
buf BUF1 (N7029, N7022);
xor XOR2 (N7030, N7014, N3703);
buf BUF1 (N7031, N7029);
nor NOR3 (N7032, N7028, N6522, N448);
nor NOR2 (N7033, N7030, N228);
or OR4 (N7034, N7016, N1732, N6553, N1633);
nand NAND4 (N7035, N7033, N3057, N6599, N799);
nand NAND2 (N7036, N7027, N1863);
or OR3 (N7037, N7031, N3725, N5328);
nor NOR3 (N7038, N7032, N7026, N5737);
nor NOR2 (N7039, N3607, N904);
buf BUF1 (N7040, N7024);
not NOT1 (N7041, N7012);
buf BUF1 (N7042, N7034);
xor XOR2 (N7043, N7040, N270);
and AND4 (N7044, N7037, N3721, N3376, N4998);
not NOT1 (N7045, N7036);
nor NOR4 (N7046, N7044, N1404, N2362, N3503);
xor XOR2 (N7047, N7038, N5928);
and AND2 (N7048, N7023, N4989);
buf BUF1 (N7049, N7043);
and AND3 (N7050, N7049, N4714, N4179);
nand NAND3 (N7051, N7046, N3575, N4056);
and AND3 (N7052, N7048, N3009, N2199);
xor XOR2 (N7053, N7041, N899);
not NOT1 (N7054, N7052);
nor NOR3 (N7055, N7035, N457, N1109);
xor XOR2 (N7056, N7050, N6291);
nand NAND3 (N7057, N7056, N748, N2336);
nor NOR3 (N7058, N7045, N1227, N6919);
xor XOR2 (N7059, N7053, N1822);
nand NAND4 (N7060, N7058, N3529, N5855, N3418);
buf BUF1 (N7061, N7057);
or OR4 (N7062, N7061, N3315, N4629, N1313);
not NOT1 (N7063, N7051);
nand NAND2 (N7064, N7062, N4859);
not NOT1 (N7065, N7059);
not NOT1 (N7066, N7047);
and AND2 (N7067, N7055, N2891);
nand NAND3 (N7068, N7025, N2978, N6674);
xor XOR2 (N7069, N7063, N2066);
nand NAND3 (N7070, N7054, N6215, N6952);
or OR4 (N7071, N7039, N5586, N4201, N5707);
xor XOR2 (N7072, N7068, N3409);
nor NOR4 (N7073, N7069, N3353, N2986, N4979);
and AND4 (N7074, N7071, N6227, N1872, N5261);
and AND3 (N7075, N7042, N6590, N4264);
nand NAND2 (N7076, N7074, N3604);
xor XOR2 (N7077, N7072, N5390);
and AND3 (N7078, N7073, N5245, N6238);
or OR4 (N7079, N7064, N4098, N1676, N1037);
and AND2 (N7080, N7079, N502);
and AND2 (N7081, N7070, N4343);
xor XOR2 (N7082, N7081, N6477);
buf BUF1 (N7083, N7075);
buf BUF1 (N7084, N7083);
nor NOR2 (N7085, N7077, N878);
buf BUF1 (N7086, N7066);
buf BUF1 (N7087, N7078);
buf BUF1 (N7088, N7060);
or OR2 (N7089, N7082, N3512);
xor XOR2 (N7090, N7088, N502);
xor XOR2 (N7091, N7065, N1207);
or OR3 (N7092, N7089, N7063, N6323);
or OR4 (N7093, N7090, N6285, N2108, N6408);
or OR4 (N7094, N7076, N1422, N4110, N5521);
not NOT1 (N7095, N7080);
xor XOR2 (N7096, N7091, N4182);
and AND2 (N7097, N7067, N3630);
xor XOR2 (N7098, N7095, N505);
nor NOR3 (N7099, N7098, N6564, N970);
xor XOR2 (N7100, N7084, N3774);
nor NOR4 (N7101, N7097, N5280, N2950, N7025);
not NOT1 (N7102, N7099);
nor NOR3 (N7103, N7087, N1356, N7027);
or OR3 (N7104, N7102, N568, N4309);
xor XOR2 (N7105, N7096, N951);
nor NOR3 (N7106, N7094, N6765, N4600);
and AND2 (N7107, N7103, N2040);
nand NAND4 (N7108, N7100, N4803, N3510, N5247);
nor NOR4 (N7109, N7107, N2953, N1673, N655);
and AND2 (N7110, N7105, N5881);
buf BUF1 (N7111, N7093);
buf BUF1 (N7112, N7110);
nor NOR3 (N7113, N7101, N1348, N6084);
or OR2 (N7114, N7086, N4132);
buf BUF1 (N7115, N7104);
not NOT1 (N7116, N7092);
and AND2 (N7117, N7111, N876);
buf BUF1 (N7118, N7115);
nor NOR2 (N7119, N7117, N5305);
xor XOR2 (N7120, N7085, N4219);
not NOT1 (N7121, N7120);
nand NAND2 (N7122, N7116, N3797);
and AND2 (N7123, N7118, N203);
xor XOR2 (N7124, N7113, N6293);
nor NOR3 (N7125, N7112, N2142, N4357);
or OR3 (N7126, N7106, N6766, N2454);
nand NAND4 (N7127, N7122, N3326, N89, N2758);
nand NAND4 (N7128, N7126, N3585, N7035, N4336);
buf BUF1 (N7129, N7121);
nand NAND3 (N7130, N7127, N786, N2760);
not NOT1 (N7131, N7114);
xor XOR2 (N7132, N7119, N5054);
and AND2 (N7133, N7123, N777);
buf BUF1 (N7134, N7133);
or OR2 (N7135, N7129, N6878);
not NOT1 (N7136, N7124);
and AND4 (N7137, N7131, N5178, N3209, N7010);
nand NAND3 (N7138, N7132, N4727, N1591);
xor XOR2 (N7139, N7136, N612);
and AND4 (N7140, N7135, N2836, N6500, N734);
buf BUF1 (N7141, N7138);
xor XOR2 (N7142, N7134, N2753);
and AND3 (N7143, N7140, N2713, N6723);
not NOT1 (N7144, N7139);
xor XOR2 (N7145, N7144, N4769);
not NOT1 (N7146, N7142);
buf BUF1 (N7147, N7141);
and AND2 (N7148, N7146, N806);
nor NOR2 (N7149, N7148, N3900);
nand NAND3 (N7150, N7149, N6102, N3391);
and AND3 (N7151, N7150, N4596, N2561);
nor NOR4 (N7152, N7145, N1707, N5376, N480);
xor XOR2 (N7153, N7130, N3020);
nor NOR2 (N7154, N7109, N6814);
nor NOR2 (N7155, N7151, N3223);
buf BUF1 (N7156, N7108);
not NOT1 (N7157, N7137);
not NOT1 (N7158, N7147);
buf BUF1 (N7159, N7154);
and AND2 (N7160, N7155, N5034);
buf BUF1 (N7161, N7158);
or OR2 (N7162, N7152, N4248);
nor NOR3 (N7163, N7157, N3096, N2952);
xor XOR2 (N7164, N7125, N6146);
xor XOR2 (N7165, N7162, N608);
or OR2 (N7166, N7165, N1203);
xor XOR2 (N7167, N7166, N2042);
buf BUF1 (N7168, N7161);
not NOT1 (N7169, N7164);
and AND2 (N7170, N7160, N7068);
nor NOR2 (N7171, N7159, N3361);
buf BUF1 (N7172, N7143);
buf BUF1 (N7173, N7153);
or OR4 (N7174, N7128, N6226, N5865, N1583);
xor XOR2 (N7175, N7171, N5224);
and AND4 (N7176, N7173, N5682, N196, N5296);
not NOT1 (N7177, N7167);
xor XOR2 (N7178, N7176, N1804);
and AND3 (N7179, N7172, N4865, N1693);
nand NAND3 (N7180, N7169, N6445, N1874);
buf BUF1 (N7181, N7156);
xor XOR2 (N7182, N7174, N4283);
nor NOR2 (N7183, N7163, N788);
or OR3 (N7184, N7179, N1731, N4539);
not NOT1 (N7185, N7184);
or OR3 (N7186, N7185, N3996, N2040);
or OR2 (N7187, N7175, N4772);
xor XOR2 (N7188, N7178, N2243);
and AND3 (N7189, N7168, N2255, N1105);
or OR4 (N7190, N7183, N4421, N6756, N1053);
buf BUF1 (N7191, N7189);
or OR3 (N7192, N7191, N802, N5168);
nor NOR2 (N7193, N7180, N3488);
not NOT1 (N7194, N7182);
nor NOR2 (N7195, N7192, N3845);
xor XOR2 (N7196, N7188, N7107);
nand NAND4 (N7197, N7170, N6497, N4992, N4532);
nand NAND2 (N7198, N7187, N3481);
and AND4 (N7199, N7186, N6594, N4304, N4479);
xor XOR2 (N7200, N7198, N3500);
xor XOR2 (N7201, N7197, N2145);
nand NAND2 (N7202, N7199, N1900);
nor NOR4 (N7203, N7190, N6244, N2795, N7193);
buf BUF1 (N7204, N3481);
or OR4 (N7205, N7203, N125, N4178, N5292);
and AND2 (N7206, N7205, N2679);
or OR2 (N7207, N7177, N4638);
and AND4 (N7208, N7206, N4615, N367, N3704);
xor XOR2 (N7209, N7202, N6620);
buf BUF1 (N7210, N7181);
buf BUF1 (N7211, N7210);
nand NAND2 (N7212, N7207, N3837);
not NOT1 (N7213, N7196);
not NOT1 (N7214, N7208);
nor NOR4 (N7215, N7200, N4228, N571, N4037);
and AND4 (N7216, N7211, N1185, N2406, N3633);
or OR2 (N7217, N7195, N2626);
nor NOR4 (N7218, N7213, N5299, N830, N505);
not NOT1 (N7219, N7204);
nand NAND4 (N7220, N7216, N5407, N3764, N6661);
buf BUF1 (N7221, N7217);
buf BUF1 (N7222, N7221);
and AND4 (N7223, N7214, N1904, N943, N2507);
nand NAND4 (N7224, N7218, N5155, N3316, N2089);
or OR4 (N7225, N7220, N2416, N1865, N6250);
xor XOR2 (N7226, N7201, N1010);
buf BUF1 (N7227, N7212);
not NOT1 (N7228, N7225);
buf BUF1 (N7229, N7223);
buf BUF1 (N7230, N7194);
and AND3 (N7231, N7215, N1002, N5074);
xor XOR2 (N7232, N7231, N5127);
or OR3 (N7233, N7224, N2278, N5098);
buf BUF1 (N7234, N7232);
nor NOR2 (N7235, N7209, N6553);
and AND3 (N7236, N7226, N3772, N4238);
not NOT1 (N7237, N7219);
not NOT1 (N7238, N7227);
and AND3 (N7239, N7222, N4858, N5433);
buf BUF1 (N7240, N7239);
nand NAND2 (N7241, N7228, N4537);
nand NAND4 (N7242, N7230, N6752, N4551, N2996);
not NOT1 (N7243, N7236);
or OR3 (N7244, N7229, N165, N2932);
buf BUF1 (N7245, N7244);
xor XOR2 (N7246, N7235, N2044);
and AND3 (N7247, N7246, N1418, N5674);
xor XOR2 (N7248, N7233, N1382);
xor XOR2 (N7249, N7248, N6099);
nor NOR2 (N7250, N7242, N4254);
or OR3 (N7251, N7247, N4915, N3664);
not NOT1 (N7252, N7241);
nor NOR3 (N7253, N7240, N6259, N3119);
nor NOR3 (N7254, N7249, N5886, N2088);
buf BUF1 (N7255, N7251);
nand NAND2 (N7256, N7255, N2262);
or OR2 (N7257, N7238, N5048);
xor XOR2 (N7258, N7245, N2408);
xor XOR2 (N7259, N7250, N2256);
nand NAND3 (N7260, N7254, N2408, N1792);
not NOT1 (N7261, N7234);
nor NOR3 (N7262, N7253, N3051, N6942);
nand NAND4 (N7263, N7261, N3936, N2089, N2807);
xor XOR2 (N7264, N7263, N4273);
buf BUF1 (N7265, N7256);
not NOT1 (N7266, N7265);
or OR3 (N7267, N7259, N715, N4568);
or OR3 (N7268, N7266, N5270, N6994);
nand NAND2 (N7269, N7260, N1238);
not NOT1 (N7270, N7269);
xor XOR2 (N7271, N7258, N4983);
nor NOR2 (N7272, N7267, N1802);
nor NOR4 (N7273, N7272, N4002, N6066, N5931);
nor NOR4 (N7274, N7237, N6788, N1444, N3518);
not NOT1 (N7275, N7271);
not NOT1 (N7276, N7257);
nand NAND2 (N7277, N7243, N3336);
xor XOR2 (N7278, N7270, N2333);
nand NAND2 (N7279, N7252, N68);
nand NAND3 (N7280, N7264, N4934, N2207);
buf BUF1 (N7281, N7273);
nand NAND2 (N7282, N7279, N6237);
nor NOR3 (N7283, N7278, N1305, N1653);
nand NAND3 (N7284, N7281, N3104, N1652);
nor NOR4 (N7285, N7277, N480, N5314, N3460);
not NOT1 (N7286, N7280);
or OR3 (N7287, N7283, N2403, N5299);
and AND3 (N7288, N7284, N2209, N3493);
or OR2 (N7289, N7275, N7275);
not NOT1 (N7290, N7276);
not NOT1 (N7291, N7268);
xor XOR2 (N7292, N7287, N2425);
xor XOR2 (N7293, N7274, N3776);
nor NOR3 (N7294, N7291, N6024, N1621);
and AND4 (N7295, N7262, N3319, N1935, N6160);
buf BUF1 (N7296, N7289);
or OR3 (N7297, N7295, N834, N3241);
xor XOR2 (N7298, N7282, N2315);
not NOT1 (N7299, N7298);
or OR3 (N7300, N7286, N5596, N454);
not NOT1 (N7301, N7297);
not NOT1 (N7302, N7296);
not NOT1 (N7303, N7299);
xor XOR2 (N7304, N7288, N3402);
and AND3 (N7305, N7301, N2031, N6666);
nor NOR2 (N7306, N7303, N4706);
or OR2 (N7307, N7304, N6450);
and AND4 (N7308, N7285, N5120, N4919, N6722);
or OR2 (N7309, N7307, N1277);
not NOT1 (N7310, N7294);
not NOT1 (N7311, N7300);
or OR3 (N7312, N7306, N4488, N4305);
buf BUF1 (N7313, N7292);
xor XOR2 (N7314, N7308, N1311);
nand NAND4 (N7315, N7310, N6428, N3899, N4985);
or OR2 (N7316, N7302, N2777);
and AND3 (N7317, N7312, N3793, N5917);
nand NAND3 (N7318, N7311, N1357, N4064);
nor NOR3 (N7319, N7317, N1860, N7141);
buf BUF1 (N7320, N7293);
buf BUF1 (N7321, N7290);
nor NOR2 (N7322, N7305, N6050);
nand NAND4 (N7323, N7318, N2644, N5262, N7189);
nand NAND4 (N7324, N7323, N2427, N4073, N5140);
or OR3 (N7325, N7321, N2496, N3065);
not NOT1 (N7326, N7319);
xor XOR2 (N7327, N7313, N3200);
and AND3 (N7328, N7322, N6800, N2860);
nor NOR3 (N7329, N7320, N2779, N251);
xor XOR2 (N7330, N7325, N5306);
and AND3 (N7331, N7309, N1899, N6162);
xor XOR2 (N7332, N7326, N2110);
or OR4 (N7333, N7329, N4017, N4343, N4327);
or OR3 (N7334, N7315, N3437, N1658);
not NOT1 (N7335, N7316);
not NOT1 (N7336, N7331);
buf BUF1 (N7337, N7333);
nand NAND4 (N7338, N7330, N1411, N5583, N2793);
and AND4 (N7339, N7314, N5452, N6190, N1217);
and AND4 (N7340, N7339, N6326, N7220, N4907);
and AND3 (N7341, N7336, N5009, N6245);
buf BUF1 (N7342, N7337);
xor XOR2 (N7343, N7328, N1715);
nor NOR4 (N7344, N7334, N380, N332, N7133);
nor NOR3 (N7345, N7338, N6370, N6115);
nor NOR3 (N7346, N7343, N4431, N3561);
buf BUF1 (N7347, N7332);
nand NAND2 (N7348, N7342, N6720);
nand NAND3 (N7349, N7341, N930, N632);
buf BUF1 (N7350, N7346);
or OR2 (N7351, N7345, N1651);
nand NAND4 (N7352, N7351, N3779, N1605, N2113);
xor XOR2 (N7353, N7347, N2610);
not NOT1 (N7354, N7324);
not NOT1 (N7355, N7348);
buf BUF1 (N7356, N7355);
buf BUF1 (N7357, N7340);
nand NAND2 (N7358, N7350, N1097);
buf BUF1 (N7359, N7353);
and AND4 (N7360, N7358, N1062, N3925, N7316);
nor NOR4 (N7361, N7335, N7194, N5260, N4289);
and AND3 (N7362, N7360, N4663, N3227);
or OR4 (N7363, N7362, N4328, N6138, N5393);
or OR2 (N7364, N7349, N2452);
nor NOR3 (N7365, N7352, N5277, N6678);
buf BUF1 (N7366, N7363);
or OR4 (N7367, N7327, N4759, N5215, N2900);
buf BUF1 (N7368, N7366);
or OR4 (N7369, N7354, N5177, N3309, N5896);
nor NOR3 (N7370, N7369, N5780, N3565);
xor XOR2 (N7371, N7359, N2181);
or OR2 (N7372, N7371, N5185);
nor NOR3 (N7373, N7361, N1187, N624);
buf BUF1 (N7374, N7367);
buf BUF1 (N7375, N7373);
nor NOR2 (N7376, N7374, N5941);
not NOT1 (N7377, N7375);
buf BUF1 (N7378, N7370);
buf BUF1 (N7379, N7364);
or OR4 (N7380, N7344, N1271, N4505, N4950);
and AND2 (N7381, N7380, N3700);
buf BUF1 (N7382, N7378);
not NOT1 (N7383, N7376);
and AND3 (N7384, N7372, N3317, N3094);
not NOT1 (N7385, N7381);
nor NOR2 (N7386, N7365, N5962);
nand NAND2 (N7387, N7382, N7258);
and AND3 (N7388, N7384, N3290, N396);
or OR3 (N7389, N7383, N6542, N6350);
and AND3 (N7390, N7385, N1954, N696);
or OR3 (N7391, N7389, N3900, N976);
xor XOR2 (N7392, N7388, N3662);
and AND4 (N7393, N7390, N2363, N5518, N3799);
buf BUF1 (N7394, N7387);
not NOT1 (N7395, N7393);
nor NOR4 (N7396, N7356, N2401, N6678, N687);
xor XOR2 (N7397, N7379, N6883);
and AND4 (N7398, N7396, N6906, N5196, N430);
or OR3 (N7399, N7398, N4833, N1057);
xor XOR2 (N7400, N7357, N1942);
buf BUF1 (N7401, N7368);
nor NOR2 (N7402, N7400, N4083);
nor NOR3 (N7403, N7391, N5344, N4067);
nor NOR2 (N7404, N7386, N5079);
nor NOR3 (N7405, N7397, N4173, N6115);
xor XOR2 (N7406, N7399, N1868);
nand NAND4 (N7407, N7377, N2020, N3248, N6952);
xor XOR2 (N7408, N7402, N6014);
not NOT1 (N7409, N7407);
or OR4 (N7410, N7394, N4305, N2218, N4004);
not NOT1 (N7411, N7404);
buf BUF1 (N7412, N7405);
not NOT1 (N7413, N7395);
buf BUF1 (N7414, N7406);
xor XOR2 (N7415, N7403, N60);
and AND3 (N7416, N7408, N3130, N1177);
xor XOR2 (N7417, N7412, N1786);
and AND3 (N7418, N7392, N1598, N251);
buf BUF1 (N7419, N7414);
buf BUF1 (N7420, N7416);
buf BUF1 (N7421, N7419);
buf BUF1 (N7422, N7415);
xor XOR2 (N7423, N7422, N7351);
or OR2 (N7424, N7410, N323);
xor XOR2 (N7425, N7421, N6359);
or OR4 (N7426, N7409, N4660, N5357, N2168);
xor XOR2 (N7427, N7413, N3031);
buf BUF1 (N7428, N7423);
not NOT1 (N7429, N7426);
not NOT1 (N7430, N7418);
nor NOR2 (N7431, N7424, N2153);
nand NAND4 (N7432, N7411, N5502, N1972, N4635);
nand NAND2 (N7433, N7428, N4301);
and AND4 (N7434, N7432, N2524, N5069, N3106);
and AND3 (N7435, N7429, N6174, N4381);
xor XOR2 (N7436, N7435, N109);
or OR2 (N7437, N7417, N7131);
or OR3 (N7438, N7420, N7389, N1145);
nor NOR2 (N7439, N7438, N2353);
not NOT1 (N7440, N7431);
or OR2 (N7441, N7437, N1277);
not NOT1 (N7442, N7441);
nor NOR2 (N7443, N7427, N2423);
nand NAND4 (N7444, N7433, N2912, N7242, N3169);
nand NAND2 (N7445, N7444, N7263);
nand NAND4 (N7446, N7440, N7275, N3, N5487);
or OR3 (N7447, N7436, N3684, N6296);
not NOT1 (N7448, N7434);
nor NOR2 (N7449, N7446, N44);
xor XOR2 (N7450, N7448, N4319);
nor NOR2 (N7451, N7401, N5305);
xor XOR2 (N7452, N7451, N7087);
nand NAND3 (N7453, N7445, N2125, N1506);
nor NOR4 (N7454, N7452, N5305, N287, N2578);
and AND4 (N7455, N7453, N2657, N3710, N5762);
buf BUF1 (N7456, N7454);
xor XOR2 (N7457, N7430, N333);
nand NAND3 (N7458, N7455, N3955, N3824);
nand NAND3 (N7459, N7425, N4906, N2543);
nand NAND2 (N7460, N7442, N792);
or OR3 (N7461, N7443, N4682, N295);
nand NAND3 (N7462, N7460, N2716, N5372);
nand NAND4 (N7463, N7457, N6508, N1214, N5333);
nand NAND3 (N7464, N7458, N6915, N3591);
nor NOR4 (N7465, N7462, N3477, N3245, N6327);
or OR3 (N7466, N7459, N1467, N6818);
nand NAND2 (N7467, N7461, N526);
and AND2 (N7468, N7439, N3193);
or OR2 (N7469, N7468, N714);
not NOT1 (N7470, N7449);
buf BUF1 (N7471, N7469);
nand NAND3 (N7472, N7447, N854, N1322);
xor XOR2 (N7473, N7467, N4676);
xor XOR2 (N7474, N7470, N1592);
buf BUF1 (N7475, N7450);
xor XOR2 (N7476, N7475, N925);
or OR3 (N7477, N7463, N2615, N1015);
xor XOR2 (N7478, N7476, N3273);
nand NAND4 (N7479, N7478, N3483, N553, N1454);
and AND2 (N7480, N7479, N7024);
not NOT1 (N7481, N7465);
and AND2 (N7482, N7464, N704);
and AND2 (N7483, N7471, N2309);
nor NOR2 (N7484, N7472, N1118);
or OR2 (N7485, N7482, N2089);
buf BUF1 (N7486, N7456);
xor XOR2 (N7487, N7483, N6914);
nand NAND2 (N7488, N7480, N1642);
and AND3 (N7489, N7487, N5414, N6542);
and AND2 (N7490, N7481, N7038);
xor XOR2 (N7491, N7474, N383);
nand NAND4 (N7492, N7488, N1318, N168, N6616);
xor XOR2 (N7493, N7486, N3279);
not NOT1 (N7494, N7490);
and AND2 (N7495, N7485, N7464);
nand NAND2 (N7496, N7473, N6289);
or OR3 (N7497, N7491, N2050, N6712);
or OR2 (N7498, N7496, N2962);
nand NAND3 (N7499, N7492, N5, N3202);
nand NAND4 (N7500, N7494, N7499, N5060, N1211);
or OR4 (N7501, N6415, N803, N437, N2570);
and AND2 (N7502, N7500, N6892);
nand NAND4 (N7503, N7493, N2149, N2985, N43);
buf BUF1 (N7504, N7466);
nor NOR3 (N7505, N7504, N5650, N855);
and AND3 (N7506, N7495, N2103, N3561);
nand NAND4 (N7507, N7502, N3931, N5543, N1160);
xor XOR2 (N7508, N7477, N2142);
not NOT1 (N7509, N7497);
not NOT1 (N7510, N7484);
and AND4 (N7511, N7489, N4549, N6249, N3918);
not NOT1 (N7512, N7503);
not NOT1 (N7513, N7505);
buf BUF1 (N7514, N7513);
nand NAND2 (N7515, N7512, N5983);
not NOT1 (N7516, N7508);
nor NOR2 (N7517, N7510, N5298);
or OR2 (N7518, N7498, N3436);
buf BUF1 (N7519, N7518);
nor NOR2 (N7520, N7517, N740);
or OR3 (N7521, N7519, N1720, N6694);
and AND2 (N7522, N7506, N5326);
xor XOR2 (N7523, N7511, N629);
buf BUF1 (N7524, N7520);
nor NOR3 (N7525, N7523, N239, N4498);
and AND4 (N7526, N7522, N7385, N4014, N4615);
not NOT1 (N7527, N7521);
nor NOR2 (N7528, N7525, N7410);
not NOT1 (N7529, N7509);
nand NAND3 (N7530, N7529, N2079, N3290);
nand NAND4 (N7531, N7526, N5246, N6972, N504);
nand NAND2 (N7532, N7516, N400);
nor NOR2 (N7533, N7531, N3961);
and AND2 (N7534, N7524, N2192);
or OR3 (N7535, N7534, N3273, N4575);
nor NOR4 (N7536, N7507, N2512, N3693, N6814);
nand NAND2 (N7537, N7530, N1391);
xor XOR2 (N7538, N7514, N6527);
nand NAND4 (N7539, N7538, N291, N7263, N3526);
or OR3 (N7540, N7539, N3444, N5019);
nor NOR4 (N7541, N7527, N4862, N3301, N5855);
xor XOR2 (N7542, N7536, N2676);
nor NOR4 (N7543, N7532, N3366, N6224, N3798);
and AND2 (N7544, N7533, N2704);
or OR4 (N7545, N7544, N3480, N526, N1306);
nand NAND2 (N7546, N7542, N7205);
or OR2 (N7547, N7541, N6008);
buf BUF1 (N7548, N7515);
nand NAND3 (N7549, N7540, N7146, N7066);
and AND3 (N7550, N7501, N4246, N6251);
nor NOR4 (N7551, N7547, N7481, N171, N1734);
xor XOR2 (N7552, N7550, N431);
nand NAND3 (N7553, N7552, N5012, N5225);
xor XOR2 (N7554, N7537, N4509);
xor XOR2 (N7555, N7528, N1278);
buf BUF1 (N7556, N7553);
nor NOR2 (N7557, N7555, N2604);
xor XOR2 (N7558, N7557, N799);
nor NOR3 (N7559, N7548, N2413, N2960);
and AND2 (N7560, N7556, N5641);
nor NOR3 (N7561, N7560, N2995, N332);
not NOT1 (N7562, N7559);
not NOT1 (N7563, N7543);
and AND2 (N7564, N7535, N6423);
nor NOR3 (N7565, N7564, N6887, N5673);
nand NAND3 (N7566, N7545, N6122, N6335);
nor NOR2 (N7567, N7554, N5363);
xor XOR2 (N7568, N7562, N6775);
nor NOR2 (N7569, N7549, N2372);
and AND3 (N7570, N7565, N3298, N4552);
buf BUF1 (N7571, N7569);
xor XOR2 (N7572, N7546, N1773);
or OR2 (N7573, N7558, N7425);
buf BUF1 (N7574, N7561);
or OR3 (N7575, N7571, N6833, N853);
nand NAND2 (N7576, N7566, N2627);
buf BUF1 (N7577, N7551);
xor XOR2 (N7578, N7563, N1753);
xor XOR2 (N7579, N7568, N2847);
buf BUF1 (N7580, N7577);
buf BUF1 (N7581, N7574);
and AND3 (N7582, N7580, N285, N5235);
xor XOR2 (N7583, N7582, N3060);
not NOT1 (N7584, N7576);
and AND3 (N7585, N7581, N3907, N952);
not NOT1 (N7586, N7572);
or OR4 (N7587, N7584, N375, N1721, N267);
or OR2 (N7588, N7587, N6261);
xor XOR2 (N7589, N7575, N6694);
or OR4 (N7590, N7579, N6627, N3242, N1860);
nor NOR2 (N7591, N7589, N4493);
xor XOR2 (N7592, N7578, N3670);
and AND3 (N7593, N7592, N3993, N6477);
nor NOR3 (N7594, N7588, N4888, N810);
xor XOR2 (N7595, N7573, N5771);
buf BUF1 (N7596, N7591);
nand NAND4 (N7597, N7570, N6474, N4059, N3712);
buf BUF1 (N7598, N7594);
and AND2 (N7599, N7590, N1646);
and AND2 (N7600, N7596, N3660);
and AND4 (N7601, N7599, N4535, N5732, N7205);
not NOT1 (N7602, N7586);
nor NOR3 (N7603, N7597, N6668, N4440);
nand NAND3 (N7604, N7585, N5547, N997);
buf BUF1 (N7605, N7603);
nor NOR2 (N7606, N7601, N822);
not NOT1 (N7607, N7567);
buf BUF1 (N7608, N7593);
buf BUF1 (N7609, N7583);
and AND3 (N7610, N7600, N3593, N1806);
or OR3 (N7611, N7605, N3181, N1603);
and AND3 (N7612, N7602, N7305, N1675);
and AND2 (N7613, N7598, N2779);
not NOT1 (N7614, N7610);
buf BUF1 (N7615, N7614);
nor NOR3 (N7616, N7609, N7400, N382);
nor NOR3 (N7617, N7611, N922, N1147);
or OR4 (N7618, N7613, N1067, N3197, N6042);
nor NOR2 (N7619, N7612, N5360);
nor NOR4 (N7620, N7617, N703, N1187, N2901);
not NOT1 (N7621, N7606);
buf BUF1 (N7622, N7621);
or OR2 (N7623, N7604, N4463);
xor XOR2 (N7624, N7619, N3928);
xor XOR2 (N7625, N7618, N5504);
buf BUF1 (N7626, N7622);
nor NOR4 (N7627, N7625, N5150, N4610, N5486);
and AND4 (N7628, N7615, N5548, N1112, N6158);
xor XOR2 (N7629, N7607, N7485);
nand NAND2 (N7630, N7629, N833);
nand NAND2 (N7631, N7623, N5258);
xor XOR2 (N7632, N7616, N3306);
nor NOR4 (N7633, N7632, N2059, N7161, N7600);
and AND3 (N7634, N7633, N7308, N7467);
nand NAND3 (N7635, N7634, N1779, N963);
buf BUF1 (N7636, N7635);
nor NOR2 (N7637, N7608, N3555);
and AND2 (N7638, N7624, N855);
or OR3 (N7639, N7636, N4519, N4859);
buf BUF1 (N7640, N7631);
xor XOR2 (N7641, N7627, N3259);
xor XOR2 (N7642, N7626, N5847);
buf BUF1 (N7643, N7630);
nand NAND3 (N7644, N7639, N2882, N716);
nor NOR3 (N7645, N7595, N7198, N240);
xor XOR2 (N7646, N7620, N716);
nor NOR3 (N7647, N7642, N3487, N2734);
nand NAND2 (N7648, N7644, N4862);
or OR2 (N7649, N7647, N3845);
nand NAND4 (N7650, N7646, N326, N3471, N1259);
nor NOR2 (N7651, N7641, N5775);
and AND2 (N7652, N7628, N2555);
buf BUF1 (N7653, N7645);
nand NAND2 (N7654, N7638, N1363);
nand NAND3 (N7655, N7651, N3268, N4638);
xor XOR2 (N7656, N7653, N339);
not NOT1 (N7657, N7637);
nand NAND2 (N7658, N7649, N1454);
nand NAND2 (N7659, N7658, N749);
and AND3 (N7660, N7654, N1104, N3983);
nor NOR3 (N7661, N7659, N2182, N7072);
xor XOR2 (N7662, N7650, N682);
not NOT1 (N7663, N7662);
buf BUF1 (N7664, N7657);
not NOT1 (N7665, N7661);
buf BUF1 (N7666, N7643);
nand NAND3 (N7667, N7665, N4320, N3755);
nor NOR3 (N7668, N7666, N6357, N780);
and AND2 (N7669, N7668, N6400);
or OR4 (N7670, N7656, N1097, N5277, N1376);
not NOT1 (N7671, N7670);
nand NAND3 (N7672, N7648, N3292, N3605);
and AND3 (N7673, N7655, N1532, N178);
nand NAND4 (N7674, N7673, N4686, N736, N4237);
buf BUF1 (N7675, N7671);
and AND3 (N7676, N7672, N6650, N1798);
or OR4 (N7677, N7675, N501, N4895, N6744);
and AND4 (N7678, N7640, N2545, N1986, N5942);
xor XOR2 (N7679, N7677, N7408);
not NOT1 (N7680, N7652);
nor NOR2 (N7681, N7664, N1609);
and AND2 (N7682, N7676, N726);
and AND4 (N7683, N7678, N5279, N6968, N1581);
not NOT1 (N7684, N7663);
and AND2 (N7685, N7684, N1345);
buf BUF1 (N7686, N7679);
not NOT1 (N7687, N7674);
not NOT1 (N7688, N7683);
xor XOR2 (N7689, N7688, N5279);
and AND4 (N7690, N7681, N5499, N3058, N2330);
and AND2 (N7691, N7680, N1075);
not NOT1 (N7692, N7691);
buf BUF1 (N7693, N7669);
nand NAND4 (N7694, N7682, N2109, N6911, N3597);
and AND3 (N7695, N7693, N6736, N7123);
nand NAND3 (N7696, N7695, N5487, N876);
nand NAND4 (N7697, N7685, N2350, N7499, N4606);
nor NOR4 (N7698, N7697, N453, N2671, N4470);
nor NOR2 (N7699, N7686, N2107);
buf BUF1 (N7700, N7699);
and AND2 (N7701, N7667, N5472);
or OR2 (N7702, N7700, N1599);
xor XOR2 (N7703, N7687, N5751);
and AND2 (N7704, N7692, N623);
and AND4 (N7705, N7690, N5431, N1239, N3923);
buf BUF1 (N7706, N7704);
or OR2 (N7707, N7694, N281);
xor XOR2 (N7708, N7705, N3595);
buf BUF1 (N7709, N7703);
not NOT1 (N7710, N7689);
and AND4 (N7711, N7709, N6930, N578, N1517);
nand NAND2 (N7712, N7711, N3368);
xor XOR2 (N7713, N7708, N4004);
buf BUF1 (N7714, N7710);
or OR3 (N7715, N7698, N7685, N2455);
nor NOR3 (N7716, N7707, N323, N4304);
not NOT1 (N7717, N7696);
nor NOR2 (N7718, N7716, N2307);
buf BUF1 (N7719, N7706);
not NOT1 (N7720, N7715);
xor XOR2 (N7721, N7713, N3621);
or OR4 (N7722, N7721, N3225, N1121, N4442);
buf BUF1 (N7723, N7720);
not NOT1 (N7724, N7712);
and AND4 (N7725, N7701, N7223, N1540, N7303);
xor XOR2 (N7726, N7719, N5997);
xor XOR2 (N7727, N7702, N4488);
buf BUF1 (N7728, N7725);
nand NAND3 (N7729, N7727, N4578, N1090);
not NOT1 (N7730, N7729);
and AND4 (N7731, N7726, N5426, N1720, N6946);
and AND2 (N7732, N7660, N6173);
not NOT1 (N7733, N7730);
or OR4 (N7734, N7732, N1628, N4617, N747);
and AND4 (N7735, N7734, N920, N4717, N4588);
or OR3 (N7736, N7735, N2663, N5024);
nand NAND4 (N7737, N7736, N3342, N2917, N4085);
nand NAND4 (N7738, N7718, N6514, N3224, N2324);
xor XOR2 (N7739, N7737, N4656);
buf BUF1 (N7740, N7733);
and AND3 (N7741, N7739, N5560, N2294);
buf BUF1 (N7742, N7724);
and AND4 (N7743, N7714, N1245, N6402, N5442);
nand NAND2 (N7744, N7723, N1610);
buf BUF1 (N7745, N7744);
nor NOR4 (N7746, N7728, N3745, N4150, N3893);
buf BUF1 (N7747, N7743);
not NOT1 (N7748, N7740);
and AND4 (N7749, N7722, N6272, N1399, N1748);
buf BUF1 (N7750, N7742);
not NOT1 (N7751, N7717);
not NOT1 (N7752, N7750);
nor NOR2 (N7753, N7747, N5736);
nand NAND3 (N7754, N7749, N3018, N5116);
nand NAND2 (N7755, N7746, N1533);
or OR2 (N7756, N7753, N4907);
nor NOR2 (N7757, N7741, N6935);
nand NAND4 (N7758, N7757, N7544, N7536, N1494);
nor NOR4 (N7759, N7748, N4042, N4588, N5414);
not NOT1 (N7760, N7756);
not NOT1 (N7761, N7754);
nor NOR2 (N7762, N7761, N5596);
or OR2 (N7763, N7738, N875);
xor XOR2 (N7764, N7751, N909);
not NOT1 (N7765, N7745);
xor XOR2 (N7766, N7760, N5138);
or OR3 (N7767, N7765, N5580, N3451);
not NOT1 (N7768, N7731);
buf BUF1 (N7769, N7764);
buf BUF1 (N7770, N7755);
buf BUF1 (N7771, N7752);
nand NAND4 (N7772, N7769, N1799, N3974, N6660);
not NOT1 (N7773, N7763);
buf BUF1 (N7774, N7759);
nor NOR4 (N7775, N7772, N6658, N2065, N2344);
nand NAND4 (N7776, N7775, N4924, N2771, N6417);
xor XOR2 (N7777, N7770, N468);
buf BUF1 (N7778, N7777);
or OR2 (N7779, N7758, N2929);
and AND4 (N7780, N7768, N528, N2012, N3791);
xor XOR2 (N7781, N7773, N3204);
xor XOR2 (N7782, N7778, N1676);
buf BUF1 (N7783, N7774);
xor XOR2 (N7784, N7762, N604);
nand NAND4 (N7785, N7767, N3522, N5271, N6055);
nand NAND3 (N7786, N7766, N1682, N6927);
nor NOR3 (N7787, N7785, N1858, N5768);
or OR4 (N7788, N7781, N3955, N2232, N213);
and AND4 (N7789, N7782, N4676, N3595, N1176);
or OR4 (N7790, N7783, N2400, N5587, N7213);
and AND4 (N7791, N7788, N5949, N1768, N254);
not NOT1 (N7792, N7786);
xor XOR2 (N7793, N7776, N951);
xor XOR2 (N7794, N7792, N5133);
buf BUF1 (N7795, N7780);
buf BUF1 (N7796, N7795);
or OR4 (N7797, N7793, N2859, N3681, N5639);
buf BUF1 (N7798, N7787);
buf BUF1 (N7799, N7771);
buf BUF1 (N7800, N7789);
or OR2 (N7801, N7798, N5915);
and AND2 (N7802, N7779, N1403);
nor NOR2 (N7803, N7799, N2794);
xor XOR2 (N7804, N7803, N3942);
and AND3 (N7805, N7784, N5349, N7770);
buf BUF1 (N7806, N7802);
buf BUF1 (N7807, N7800);
xor XOR2 (N7808, N7791, N5459);
and AND3 (N7809, N7796, N6244, N4543);
not NOT1 (N7810, N7808);
nand NAND3 (N7811, N7806, N4852, N1314);
xor XOR2 (N7812, N7797, N6719);
buf BUF1 (N7813, N7801);
and AND3 (N7814, N7807, N4844, N6657);
or OR3 (N7815, N7812, N1565, N353);
and AND2 (N7816, N7813, N6944);
nor NOR3 (N7817, N7816, N251, N6643);
not NOT1 (N7818, N7790);
or OR2 (N7819, N7804, N6893);
buf BUF1 (N7820, N7805);
buf BUF1 (N7821, N7814);
or OR2 (N7822, N7820, N5846);
nand NAND3 (N7823, N7819, N3170, N4174);
buf BUF1 (N7824, N7817);
xor XOR2 (N7825, N7822, N5323);
nand NAND3 (N7826, N7809, N4672, N3001);
nand NAND2 (N7827, N7815, N5299);
buf BUF1 (N7828, N7821);
or OR2 (N7829, N7825, N7644);
or OR3 (N7830, N7823, N1544, N4079);
nand NAND2 (N7831, N7811, N3432);
nor NOR4 (N7832, N7831, N7432, N7320, N4151);
and AND2 (N7833, N7829, N6150);
xor XOR2 (N7834, N7794, N1114);
and AND4 (N7835, N7832, N5824, N4744, N181);
and AND2 (N7836, N7828, N218);
xor XOR2 (N7837, N7826, N4044);
and AND3 (N7838, N7818, N71, N7726);
nor NOR2 (N7839, N7837, N4974);
not NOT1 (N7840, N7810);
not NOT1 (N7841, N7833);
xor XOR2 (N7842, N7834, N5227);
nand NAND3 (N7843, N7838, N895, N1346);
and AND2 (N7844, N7840, N4938);
and AND2 (N7845, N7827, N5382);
or OR4 (N7846, N7830, N1067, N5137, N4994);
and AND2 (N7847, N7844, N423);
nand NAND2 (N7848, N7842, N7533);
and AND4 (N7849, N7836, N419, N6946, N5028);
nand NAND4 (N7850, N7824, N208, N4601, N95);
buf BUF1 (N7851, N7848);
or OR2 (N7852, N7847, N6439);
nand NAND3 (N7853, N7835, N1741, N544);
not NOT1 (N7854, N7852);
nor NOR4 (N7855, N7843, N4383, N3041, N3206);
not NOT1 (N7856, N7850);
xor XOR2 (N7857, N7839, N3966);
nand NAND2 (N7858, N7857, N3511);
buf BUF1 (N7859, N7851);
nor NOR3 (N7860, N7854, N480, N7798);
or OR4 (N7861, N7846, N1703, N3790, N7476);
or OR4 (N7862, N7853, N6493, N6034, N6489);
or OR3 (N7863, N7858, N5980, N4637);
nand NAND4 (N7864, N7856, N6812, N1917, N175);
nand NAND2 (N7865, N7860, N6401);
buf BUF1 (N7866, N7864);
and AND4 (N7867, N7862, N3301, N7446, N2069);
or OR3 (N7868, N7866, N2421, N424);
and AND4 (N7869, N7865, N638, N6074, N3789);
or OR3 (N7870, N7849, N3179, N1308);
nand NAND2 (N7871, N7859, N1510);
buf BUF1 (N7872, N7870);
xor XOR2 (N7873, N7872, N1034);
not NOT1 (N7874, N7841);
xor XOR2 (N7875, N7873, N7024);
buf BUF1 (N7876, N7871);
buf BUF1 (N7877, N7863);
xor XOR2 (N7878, N7875, N6131);
xor XOR2 (N7879, N7869, N569);
buf BUF1 (N7880, N7867);
not NOT1 (N7881, N7880);
nor NOR4 (N7882, N7878, N7559, N1096, N5007);
not NOT1 (N7883, N7879);
and AND2 (N7884, N7876, N4966);
not NOT1 (N7885, N7861);
nor NOR2 (N7886, N7868, N423);
not NOT1 (N7887, N7886);
and AND4 (N7888, N7855, N2423, N5297, N3068);
not NOT1 (N7889, N7888);
xor XOR2 (N7890, N7877, N819);
not NOT1 (N7891, N7881);
xor XOR2 (N7892, N7874, N3307);
or OR2 (N7893, N7883, N6475);
nand NAND3 (N7894, N7890, N7193, N7506);
nor NOR4 (N7895, N7884, N4654, N3472, N1769);
not NOT1 (N7896, N7885);
nand NAND4 (N7897, N7882, N7643, N1934, N6529);
nand NAND4 (N7898, N7892, N4319, N5438, N4685);
buf BUF1 (N7899, N7891);
nor NOR2 (N7900, N7896, N5377);
nand NAND2 (N7901, N7900, N6095);
nor NOR4 (N7902, N7899, N5973, N5934, N3154);
nor NOR2 (N7903, N7894, N4195);
nand NAND4 (N7904, N7898, N3641, N6437, N751);
or OR2 (N7905, N7893, N35);
nor NOR3 (N7906, N7903, N2753, N6762);
buf BUF1 (N7907, N7897);
nor NOR2 (N7908, N7904, N5942);
nor NOR2 (N7909, N7908, N6502);
or OR2 (N7910, N7901, N2290);
or OR2 (N7911, N7902, N218);
xor XOR2 (N7912, N7905, N3683);
xor XOR2 (N7913, N7889, N4305);
not NOT1 (N7914, N7906);
nand NAND3 (N7915, N7912, N2935, N4444);
xor XOR2 (N7916, N7887, N3282);
nand NAND4 (N7917, N7914, N5778, N4084, N586);
xor XOR2 (N7918, N7917, N5285);
buf BUF1 (N7919, N7916);
and AND3 (N7920, N7895, N3335, N6591);
or OR3 (N7921, N7918, N3566, N2212);
and AND3 (N7922, N7911, N822, N4903);
or OR3 (N7923, N7909, N3721, N6062);
and AND2 (N7924, N7907, N7893);
xor XOR2 (N7925, N7923, N4868);
nand NAND4 (N7926, N7919, N4225, N5689, N5988);
and AND2 (N7927, N7920, N136);
or OR2 (N7928, N7845, N2264);
not NOT1 (N7929, N7921);
and AND2 (N7930, N7915, N1044);
nand NAND2 (N7931, N7926, N3721);
nand NAND3 (N7932, N7910, N4587, N594);
nor NOR2 (N7933, N7927, N7173);
xor XOR2 (N7934, N7931, N3490);
and AND3 (N7935, N7929, N3259, N7495);
xor XOR2 (N7936, N7930, N3516);
or OR3 (N7937, N7928, N508, N1213);
nand NAND3 (N7938, N7937, N2436, N5179);
nand NAND4 (N7939, N7936, N6103, N3368, N1061);
nand NAND4 (N7940, N7938, N7554, N2484, N7690);
or OR4 (N7941, N7924, N3669, N7057, N6153);
or OR2 (N7942, N7934, N4600);
xor XOR2 (N7943, N7925, N4202);
xor XOR2 (N7944, N7940, N5695);
xor XOR2 (N7945, N7935, N589);
and AND3 (N7946, N7941, N5798, N7238);
buf BUF1 (N7947, N7932);
not NOT1 (N7948, N7942);
and AND4 (N7949, N7922, N5604, N2439, N237);
nand NAND4 (N7950, N7949, N891, N2156, N342);
nor NOR2 (N7951, N7939, N4032);
not NOT1 (N7952, N7943);
or OR4 (N7953, N7948, N4782, N3446, N1175);
buf BUF1 (N7954, N7950);
xor XOR2 (N7955, N7947, N3078);
or OR2 (N7956, N7955, N3419);
nand NAND4 (N7957, N7953, N7690, N6417, N5913);
xor XOR2 (N7958, N7956, N7591);
buf BUF1 (N7959, N7944);
and AND2 (N7960, N7945, N851);
nor NOR4 (N7961, N7958, N865, N7610, N206);
buf BUF1 (N7962, N7959);
not NOT1 (N7963, N7961);
nor NOR4 (N7964, N7962, N7284, N2908, N602);
xor XOR2 (N7965, N7951, N6958);
nand NAND3 (N7966, N7954, N7428, N3653);
xor XOR2 (N7967, N7933, N3090);
nor NOR3 (N7968, N7967, N2575, N184);
buf BUF1 (N7969, N7913);
not NOT1 (N7970, N7969);
and AND2 (N7971, N7960, N340);
nor NOR3 (N7972, N7963, N784, N7320);
not NOT1 (N7973, N7971);
not NOT1 (N7974, N7966);
nor NOR4 (N7975, N7970, N1894, N3077, N7788);
buf BUF1 (N7976, N7957);
and AND3 (N7977, N7952, N6580, N1476);
nor NOR2 (N7978, N7973, N3038);
buf BUF1 (N7979, N7974);
buf BUF1 (N7980, N7964);
and AND4 (N7981, N7980, N4947, N2709, N6697);
and AND3 (N7982, N7979, N2586, N2407);
and AND3 (N7983, N7965, N2233, N2552);
nor NOR4 (N7984, N7972, N554, N2849, N5031);
not NOT1 (N7985, N7975);
nand NAND3 (N7986, N7981, N4264, N101);
nand NAND2 (N7987, N7986, N1190);
not NOT1 (N7988, N7946);
buf BUF1 (N7989, N7987);
nor NOR3 (N7990, N7989, N6392, N4349);
xor XOR2 (N7991, N7990, N7894);
xor XOR2 (N7992, N7988, N5022);
or OR4 (N7993, N7992, N5427, N7182, N5548);
or OR2 (N7994, N7983, N1034);
not NOT1 (N7995, N7984);
not NOT1 (N7996, N7977);
not NOT1 (N7997, N7978);
nor NOR4 (N7998, N7985, N943, N3610, N4853);
or OR2 (N7999, N7993, N6173);
not NOT1 (N8000, N7976);
or OR3 (N8001, N7994, N6530, N7422);
nand NAND4 (N8002, N7999, N154, N6679, N6907);
nor NOR3 (N8003, N7991, N2772, N7678);
or OR3 (N8004, N7982, N490, N6830);
xor XOR2 (N8005, N8001, N2005);
nand NAND3 (N8006, N8002, N3843, N6224);
nor NOR3 (N8007, N7998, N7414, N6801);
nor NOR2 (N8008, N7995, N4219);
nor NOR3 (N8009, N8005, N1163, N1946);
nand NAND2 (N8010, N8004, N1636);
buf BUF1 (N8011, N8009);
not NOT1 (N8012, N8010);
nor NOR2 (N8013, N8012, N1130);
endmodule