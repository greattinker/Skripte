// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14;

output N895,N898,N910,N891,N908,N899,N909,N913,N911,N914;

and AND4 (N15, N12, N11, N1, N14);
nor NOR4 (N16, N3, N10, N13, N11);
nand NAND4 (N17, N10, N2, N9, N15);
nor NOR3 (N18, N16, N17, N13);
nor NOR2 (N19, N12, N1);
nor NOR3 (N20, N10, N14, N9);
nor NOR3 (N21, N9, N10, N14);
not NOT1 (N22, N18);
nand NAND2 (N23, N16, N19);
nand NAND3 (N24, N6, N7, N18);
nand NAND2 (N25, N14, N23);
or OR4 (N26, N13, N12, N4, N8);
nor NOR2 (N27, N25, N6);
xor XOR2 (N28, N4, N19);
nor NOR2 (N29, N5, N14);
nor NOR2 (N30, N26, N17);
nand NAND3 (N31, N15, N11, N17);
not NOT1 (N32, N23);
buf BUF1 (N33, N29);
and AND4 (N34, N31, N24, N18, N27);
not NOT1 (N35, N23);
nand NAND3 (N36, N8, N28, N18);
nand NAND2 (N37, N31, N1);
nor NOR2 (N38, N20, N35);
nor NOR4 (N39, N38, N33, N29, N8);
nand NAND3 (N40, N13, N23, N15);
buf BUF1 (N41, N12);
not NOT1 (N42, N30);
and AND2 (N43, N42, N22);
and AND4 (N44, N23, N29, N19, N26);
xor XOR2 (N45, N40, N44);
nor NOR4 (N46, N15, N21, N7, N5);
nand NAND3 (N47, N45, N2, N33);
not NOT1 (N48, N43);
and AND3 (N49, N44, N9, N14);
nand NAND4 (N50, N37, N12, N10, N39);
and AND4 (N51, N1, N38, N28, N12);
nor NOR4 (N52, N51, N46, N36, N4);
not NOT1 (N53, N20);
and AND4 (N54, N47, N21, N18, N7);
buf BUF1 (N55, N48);
buf BUF1 (N56, N28);
not NOT1 (N57, N41);
nor NOR3 (N58, N49, N57, N22);
buf BUF1 (N59, N5);
xor XOR2 (N60, N50, N16);
nand NAND4 (N61, N32, N52, N40, N29);
nand NAND2 (N62, N9, N34);
buf BUF1 (N63, N5);
not NOT1 (N64, N59);
xor XOR2 (N65, N53, N42);
nor NOR3 (N66, N63, N56, N20);
or OR2 (N67, N45, N43);
not NOT1 (N68, N67);
or OR3 (N69, N65, N14, N28);
buf BUF1 (N70, N69);
and AND4 (N71, N64, N18, N8, N5);
xor XOR2 (N72, N70, N30);
and AND2 (N73, N66, N54);
or OR2 (N74, N10, N35);
buf BUF1 (N75, N55);
not NOT1 (N76, N75);
not NOT1 (N77, N72);
nand NAND3 (N78, N68, N54, N63);
xor XOR2 (N79, N58, N14);
nor NOR2 (N80, N62, N37);
not NOT1 (N81, N77);
or OR3 (N82, N78, N17, N61);
xor XOR2 (N83, N24, N66);
not NOT1 (N84, N76);
and AND4 (N85, N83, N38, N15, N42);
and AND4 (N86, N71, N25, N72, N45);
and AND4 (N87, N80, N85, N61, N20);
xor XOR2 (N88, N86, N36);
not NOT1 (N89, N74);
xor XOR2 (N90, N83, N16);
or OR2 (N91, N88, N39);
and AND2 (N92, N82, N67);
buf BUF1 (N93, N90);
nor NOR3 (N94, N79, N91, N91);
nand NAND2 (N95, N87, N30);
not NOT1 (N96, N54);
and AND4 (N97, N73, N96, N41, N35);
nand NAND4 (N98, N78, N86, N77, N56);
xor XOR2 (N99, N60, N12);
and AND4 (N100, N93, N21, N81, N68);
xor XOR2 (N101, N64, N22);
buf BUF1 (N102, N92);
or OR4 (N103, N98, N43, N33, N66);
buf BUF1 (N104, N100);
xor XOR2 (N105, N102, N45);
buf BUF1 (N106, N89);
nand NAND3 (N107, N95, N42, N79);
not NOT1 (N108, N106);
buf BUF1 (N109, N107);
and AND2 (N110, N108, N46);
nor NOR3 (N111, N109, N64, N27);
nor NOR3 (N112, N103, N97, N100);
buf BUF1 (N113, N62);
nor NOR2 (N114, N112, N65);
buf BUF1 (N115, N105);
nand NAND3 (N116, N99, N19, N101);
or OR3 (N117, N6, N104, N108);
buf BUF1 (N118, N86);
or OR2 (N119, N113, N62);
or OR2 (N120, N116, N47);
not NOT1 (N121, N111);
nand NAND2 (N122, N84, N119);
not NOT1 (N123, N26);
nand NAND4 (N124, N123, N85, N84, N77);
not NOT1 (N125, N118);
xor XOR2 (N126, N121, N112);
xor XOR2 (N127, N117, N67);
and AND3 (N128, N126, N36, N10);
nand NAND4 (N129, N122, N120, N127, N44);
or OR3 (N130, N19, N70, N126);
not NOT1 (N131, N84);
nor NOR4 (N132, N110, N114, N110, N119);
not NOT1 (N133, N3);
and AND2 (N134, N128, N8);
xor XOR2 (N135, N131, N80);
xor XOR2 (N136, N125, N44);
and AND4 (N137, N134, N9, N37, N110);
nor NOR2 (N138, N115, N46);
nand NAND3 (N139, N133, N25, N90);
or OR4 (N140, N136, N117, N94, N39);
not NOT1 (N141, N85);
and AND4 (N142, N129, N44, N86, N120);
xor XOR2 (N143, N137, N128);
buf BUF1 (N144, N142);
or OR2 (N145, N135, N119);
nand NAND4 (N146, N144, N46, N134, N26);
not NOT1 (N147, N130);
nand NAND2 (N148, N145, N131);
and AND2 (N149, N124, N51);
and AND4 (N150, N140, N119, N2, N95);
buf BUF1 (N151, N141);
buf BUF1 (N152, N132);
nand NAND2 (N153, N143, N43);
and AND4 (N154, N152, N31, N58, N74);
nand NAND2 (N155, N150, N117);
nand NAND3 (N156, N151, N73, N38);
or OR4 (N157, N138, N87, N126, N27);
not NOT1 (N158, N154);
xor XOR2 (N159, N153, N89);
nor NOR2 (N160, N156, N6);
not NOT1 (N161, N160);
nand NAND4 (N162, N139, N86, N130, N49);
nand NAND4 (N163, N147, N123, N121, N44);
nor NOR2 (N164, N162, N148);
nor NOR2 (N165, N153, N23);
xor XOR2 (N166, N157, N103);
buf BUF1 (N167, N166);
buf BUF1 (N168, N155);
not NOT1 (N169, N159);
not NOT1 (N170, N169);
nor NOR3 (N171, N168, N93, N59);
xor XOR2 (N172, N171, N168);
buf BUF1 (N173, N146);
buf BUF1 (N174, N167);
nand NAND3 (N175, N172, N155, N78);
and AND4 (N176, N163, N142, N43, N41);
nor NOR3 (N177, N161, N145, N174);
and AND4 (N178, N117, N95, N155, N109);
xor XOR2 (N179, N175, N46);
not NOT1 (N180, N165);
buf BUF1 (N181, N176);
xor XOR2 (N182, N149, N148);
and AND3 (N183, N173, N5, N105);
or OR4 (N184, N181, N48, N146, N13);
nand NAND3 (N185, N177, N11, N122);
nor NOR4 (N186, N183, N10, N40, N150);
nand NAND2 (N187, N184, N142);
buf BUF1 (N188, N179);
nor NOR4 (N189, N164, N164, N146, N179);
or OR4 (N190, N189, N15, N177, N156);
nand NAND4 (N191, N187, N13, N154, N183);
and AND4 (N192, N158, N75, N40, N139);
not NOT1 (N193, N180);
nor NOR2 (N194, N188, N148);
buf BUF1 (N195, N182);
nand NAND3 (N196, N192, N82, N136);
nor NOR3 (N197, N185, N12, N94);
buf BUF1 (N198, N194);
buf BUF1 (N199, N195);
nand NAND2 (N200, N186, N59);
nand NAND4 (N201, N196, N105, N86, N115);
not NOT1 (N202, N197);
or OR4 (N203, N199, N105, N129, N100);
buf BUF1 (N204, N200);
xor XOR2 (N205, N202, N90);
not NOT1 (N206, N178);
or OR2 (N207, N203, N138);
not NOT1 (N208, N190);
xor XOR2 (N209, N206, N149);
buf BUF1 (N210, N201);
nor NOR4 (N211, N170, N101, N175, N17);
nand NAND2 (N212, N193, N179);
nand NAND3 (N213, N204, N31, N12);
buf BUF1 (N214, N208);
and AND4 (N215, N213, N92, N102, N157);
xor XOR2 (N216, N198, N3);
or OR4 (N217, N207, N211, N32, N136);
and AND2 (N218, N112, N143);
not NOT1 (N219, N216);
and AND3 (N220, N218, N4, N207);
nand NAND4 (N221, N210, N204, N78, N219);
or OR3 (N222, N70, N95, N79);
buf BUF1 (N223, N214);
nor NOR3 (N224, N220, N187, N91);
and AND2 (N225, N205, N64);
not NOT1 (N226, N225);
nor NOR3 (N227, N221, N121, N169);
nor NOR4 (N228, N215, N149, N119, N74);
nor NOR2 (N229, N224, N114);
buf BUF1 (N230, N227);
xor XOR2 (N231, N226, N78);
nand NAND2 (N232, N217, N51);
buf BUF1 (N233, N223);
or OR2 (N234, N212, N1);
nand NAND2 (N235, N229, N99);
xor XOR2 (N236, N222, N26);
and AND2 (N237, N231, N112);
xor XOR2 (N238, N233, N195);
nor NOR2 (N239, N238, N114);
buf BUF1 (N240, N230);
nor NOR4 (N241, N236, N62, N107, N48);
not NOT1 (N242, N232);
xor XOR2 (N243, N239, N49);
buf BUF1 (N244, N243);
not NOT1 (N245, N241);
nand NAND4 (N246, N244, N222, N139, N180);
not NOT1 (N247, N191);
or OR3 (N248, N234, N229, N103);
nor NOR3 (N249, N237, N81, N122);
nor NOR4 (N250, N249, N8, N238, N141);
nor NOR4 (N251, N248, N62, N240, N57);
buf BUF1 (N252, N158);
nor NOR3 (N253, N250, N6, N201);
xor XOR2 (N254, N235, N198);
and AND2 (N255, N228, N192);
xor XOR2 (N256, N209, N77);
buf BUF1 (N257, N255);
xor XOR2 (N258, N254, N66);
buf BUF1 (N259, N246);
nand NAND4 (N260, N251, N125, N184, N255);
xor XOR2 (N261, N242, N213);
and AND4 (N262, N252, N62, N161, N123);
buf BUF1 (N263, N256);
buf BUF1 (N264, N257);
and AND4 (N265, N259, N242, N207, N191);
or OR2 (N266, N263, N84);
and AND4 (N267, N253, N181, N171, N199);
or OR2 (N268, N261, N232);
nor NOR2 (N269, N266, N54);
buf BUF1 (N270, N265);
xor XOR2 (N271, N264, N7);
and AND4 (N272, N262, N28, N78, N77);
buf BUF1 (N273, N269);
not NOT1 (N274, N260);
or OR2 (N275, N274, N263);
nand NAND3 (N276, N258, N144, N193);
nand NAND3 (N277, N273, N147, N192);
xor XOR2 (N278, N275, N172);
or OR3 (N279, N277, N148, N12);
nor NOR3 (N280, N268, N131, N104);
buf BUF1 (N281, N279);
nand NAND3 (N282, N270, N49, N189);
not NOT1 (N283, N247);
or OR2 (N284, N283, N110);
not NOT1 (N285, N278);
buf BUF1 (N286, N276);
or OR3 (N287, N282, N194, N96);
and AND2 (N288, N287, N141);
and AND4 (N289, N286, N32, N262, N106);
nand NAND4 (N290, N272, N46, N184, N205);
nand NAND4 (N291, N290, N275, N179, N268);
buf BUF1 (N292, N289);
not NOT1 (N293, N291);
nor NOR2 (N294, N245, N22);
buf BUF1 (N295, N293);
nor NOR4 (N296, N280, N133, N47, N232);
buf BUF1 (N297, N295);
xor XOR2 (N298, N294, N252);
not NOT1 (N299, N284);
xor XOR2 (N300, N271, N286);
and AND4 (N301, N297, N167, N79, N152);
buf BUF1 (N302, N300);
xor XOR2 (N303, N267, N136);
xor XOR2 (N304, N301, N73);
or OR3 (N305, N303, N199, N191);
or OR3 (N306, N296, N55, N80);
xor XOR2 (N307, N281, N268);
xor XOR2 (N308, N299, N262);
or OR4 (N309, N292, N192, N214, N185);
nor NOR3 (N310, N298, N97, N239);
not NOT1 (N311, N305);
buf BUF1 (N312, N308);
xor XOR2 (N313, N288, N86);
nor NOR3 (N314, N313, N102, N158);
buf BUF1 (N315, N309);
and AND3 (N316, N307, N19, N196);
xor XOR2 (N317, N311, N147);
buf BUF1 (N318, N306);
xor XOR2 (N319, N318, N182);
and AND2 (N320, N285, N10);
and AND3 (N321, N312, N108, N67);
buf BUF1 (N322, N321);
or OR4 (N323, N316, N263, N290, N179);
nand NAND2 (N324, N322, N253);
nand NAND4 (N325, N324, N44, N80, N130);
buf BUF1 (N326, N315);
buf BUF1 (N327, N314);
xor XOR2 (N328, N320, N146);
buf BUF1 (N329, N323);
buf BUF1 (N330, N319);
not NOT1 (N331, N328);
not NOT1 (N332, N302);
not NOT1 (N333, N326);
nor NOR4 (N334, N330, N210, N269, N205);
or OR3 (N335, N325, N291, N222);
xor XOR2 (N336, N304, N283);
and AND3 (N337, N332, N75, N95);
nor NOR4 (N338, N335, N165, N10, N119);
xor XOR2 (N339, N338, N298);
and AND3 (N340, N310, N26, N285);
not NOT1 (N341, N339);
xor XOR2 (N342, N337, N137);
nor NOR2 (N343, N342, N17);
nand NAND3 (N344, N329, N65, N9);
xor XOR2 (N345, N331, N319);
and AND3 (N346, N344, N277, N128);
nor NOR3 (N347, N317, N142, N240);
nand NAND4 (N348, N336, N162, N145, N97);
or OR4 (N349, N343, N67, N68, N225);
nand NAND4 (N350, N347, N349, N110, N101);
xor XOR2 (N351, N19, N186);
buf BUF1 (N352, N340);
nor NOR3 (N353, N334, N36, N232);
or OR3 (N354, N351, N64, N50);
nand NAND2 (N355, N327, N338);
not NOT1 (N356, N350);
buf BUF1 (N357, N345);
and AND2 (N358, N355, N351);
and AND3 (N359, N358, N309, N150);
or OR4 (N360, N359, N350, N159, N145);
and AND3 (N361, N354, N295, N209);
nor NOR3 (N362, N346, N80, N115);
xor XOR2 (N363, N353, N231);
nor NOR4 (N364, N348, N131, N16, N300);
xor XOR2 (N365, N363, N178);
nor NOR4 (N366, N341, N44, N46, N289);
xor XOR2 (N367, N352, N47);
nor NOR3 (N368, N362, N144, N234);
not NOT1 (N369, N366);
xor XOR2 (N370, N369, N254);
nand NAND3 (N371, N365, N63, N274);
nand NAND2 (N372, N361, N366);
buf BUF1 (N373, N370);
and AND2 (N374, N367, N161);
and AND4 (N375, N374, N57, N92, N274);
xor XOR2 (N376, N357, N315);
nand NAND3 (N377, N360, N212, N341);
nand NAND2 (N378, N375, N35);
xor XOR2 (N379, N371, N236);
and AND3 (N380, N376, N351, N190);
not NOT1 (N381, N373);
nor NOR4 (N382, N356, N1, N46, N379);
nand NAND4 (N383, N190, N99, N260, N66);
or OR4 (N384, N382, N342, N288, N338);
nand NAND4 (N385, N377, N378, N193, N154);
buf BUF1 (N386, N186);
nand NAND4 (N387, N385, N341, N221, N285);
not NOT1 (N388, N381);
nor NOR3 (N389, N368, N268, N46);
buf BUF1 (N390, N383);
not NOT1 (N391, N372);
not NOT1 (N392, N384);
or OR3 (N393, N388, N39, N155);
nand NAND4 (N394, N389, N65, N6, N141);
and AND4 (N395, N380, N115, N22, N143);
xor XOR2 (N396, N386, N243);
buf BUF1 (N397, N333);
not NOT1 (N398, N392);
and AND2 (N399, N398, N289);
nand NAND2 (N400, N399, N74);
or OR4 (N401, N393, N291, N105, N272);
nand NAND4 (N402, N395, N43, N174, N251);
and AND4 (N403, N387, N396, N107, N339);
nor NOR2 (N404, N7, N284);
buf BUF1 (N405, N390);
and AND4 (N406, N403, N156, N335, N116);
xor XOR2 (N407, N404, N368);
xor XOR2 (N408, N405, N330);
nand NAND2 (N409, N397, N271);
not NOT1 (N410, N394);
nand NAND2 (N411, N391, N153);
not NOT1 (N412, N406);
or OR2 (N413, N412, N287);
xor XOR2 (N414, N409, N113);
or OR3 (N415, N410, N295, N84);
nand NAND3 (N416, N407, N259, N345);
and AND3 (N417, N402, N93, N168);
nor NOR3 (N418, N411, N135, N34);
buf BUF1 (N419, N414);
nor NOR2 (N420, N419, N232);
not NOT1 (N421, N417);
buf BUF1 (N422, N421);
not NOT1 (N423, N408);
not NOT1 (N424, N420);
and AND3 (N425, N364, N151, N125);
or OR4 (N426, N425, N81, N150, N137);
buf BUF1 (N427, N413);
and AND3 (N428, N418, N265, N184);
or OR2 (N429, N422, N106);
or OR3 (N430, N428, N94, N320);
buf BUF1 (N431, N430);
nand NAND2 (N432, N423, N102);
xor XOR2 (N433, N429, N136);
nor NOR4 (N434, N401, N232, N284, N287);
not NOT1 (N435, N426);
or OR2 (N436, N432, N149);
nor NOR3 (N437, N433, N158, N137);
buf BUF1 (N438, N431);
nor NOR4 (N439, N400, N230, N266, N239);
nor NOR2 (N440, N415, N236);
nor NOR3 (N441, N424, N354, N272);
buf BUF1 (N442, N436);
not NOT1 (N443, N427);
nor NOR3 (N444, N434, N431, N277);
xor XOR2 (N445, N437, N439);
nand NAND2 (N446, N197, N441);
not NOT1 (N447, N139);
nand NAND4 (N448, N445, N398, N28, N116);
not NOT1 (N449, N435);
or OR2 (N450, N447, N197);
and AND3 (N451, N440, N266, N425);
nand NAND2 (N452, N446, N48);
or OR2 (N453, N443, N368);
not NOT1 (N454, N448);
buf BUF1 (N455, N416);
buf BUF1 (N456, N442);
nor NOR3 (N457, N438, N385, N386);
buf BUF1 (N458, N444);
xor XOR2 (N459, N455, N456);
nor NOR2 (N460, N231, N314);
nor NOR2 (N461, N450, N78);
nor NOR2 (N462, N458, N326);
nand NAND4 (N463, N451, N209, N166, N440);
or OR2 (N464, N449, N238);
not NOT1 (N465, N459);
buf BUF1 (N466, N460);
and AND2 (N467, N454, N207);
buf BUF1 (N468, N452);
or OR2 (N469, N466, N189);
nor NOR3 (N470, N457, N76, N40);
nor NOR4 (N471, N470, N404, N4, N108);
nand NAND4 (N472, N463, N427, N320, N71);
and AND4 (N473, N471, N410, N171, N243);
buf BUF1 (N474, N453);
buf BUF1 (N475, N472);
not NOT1 (N476, N467);
buf BUF1 (N477, N462);
nor NOR4 (N478, N465, N24, N393, N249);
nand NAND4 (N479, N478, N36, N281, N174);
nand NAND3 (N480, N468, N114, N468);
nor NOR3 (N481, N477, N209, N394);
or OR3 (N482, N474, N477, N381);
not NOT1 (N483, N481);
or OR3 (N484, N473, N47, N164);
and AND3 (N485, N483, N228, N359);
or OR4 (N486, N476, N263, N315, N456);
nor NOR2 (N487, N464, N79);
or OR2 (N488, N487, N419);
buf BUF1 (N489, N484);
not NOT1 (N490, N488);
not NOT1 (N491, N480);
nor NOR3 (N492, N485, N150, N276);
nor NOR4 (N493, N461, N137, N447, N42);
xor XOR2 (N494, N469, N21);
buf BUF1 (N495, N482);
xor XOR2 (N496, N492, N207);
not NOT1 (N497, N491);
nor NOR3 (N498, N490, N326, N148);
nand NAND3 (N499, N496, N229, N22);
or OR2 (N500, N486, N322);
xor XOR2 (N501, N500, N371);
nor NOR4 (N502, N499, N14, N237, N223);
nand NAND2 (N503, N495, N278);
or OR3 (N504, N493, N22, N194);
or OR4 (N505, N497, N87, N186, N334);
nand NAND4 (N506, N502, N203, N267, N412);
nor NOR3 (N507, N503, N263, N128);
nor NOR4 (N508, N505, N339, N132, N301);
nor NOR4 (N509, N508, N22, N465, N227);
nand NAND4 (N510, N494, N396, N112, N430);
xor XOR2 (N511, N510, N163);
not NOT1 (N512, N489);
nand NAND4 (N513, N498, N313, N330, N164);
nor NOR4 (N514, N511, N477, N341, N374);
and AND4 (N515, N509, N324, N125, N419);
and AND4 (N516, N506, N16, N173, N19);
not NOT1 (N517, N501);
nand NAND3 (N518, N516, N301, N83);
and AND4 (N519, N507, N2, N411, N319);
and AND4 (N520, N517, N262, N69, N298);
buf BUF1 (N521, N479);
and AND2 (N522, N521, N448);
xor XOR2 (N523, N520, N192);
not NOT1 (N524, N523);
not NOT1 (N525, N522);
not NOT1 (N526, N504);
nor NOR3 (N527, N475, N313, N154);
buf BUF1 (N528, N527);
buf BUF1 (N529, N514);
nand NAND2 (N530, N526, N418);
xor XOR2 (N531, N515, N367);
and AND2 (N532, N530, N31);
buf BUF1 (N533, N519);
and AND2 (N534, N533, N431);
xor XOR2 (N535, N525, N54);
not NOT1 (N536, N531);
xor XOR2 (N537, N524, N408);
and AND4 (N538, N537, N298, N270, N428);
xor XOR2 (N539, N534, N221);
xor XOR2 (N540, N532, N27);
or OR4 (N541, N513, N374, N176, N176);
buf BUF1 (N542, N528);
not NOT1 (N543, N542);
or OR4 (N544, N539, N350, N147, N175);
nor NOR4 (N545, N543, N434, N389, N356);
not NOT1 (N546, N545);
or OR2 (N547, N546, N266);
nand NAND3 (N548, N540, N224, N399);
or OR2 (N549, N547, N529);
and AND3 (N550, N9, N4, N144);
or OR4 (N551, N541, N292, N520, N77);
or OR2 (N552, N548, N370);
and AND3 (N553, N544, N173, N56);
nor NOR3 (N554, N551, N447, N6);
not NOT1 (N555, N538);
and AND3 (N556, N518, N501, N205);
and AND2 (N557, N555, N308);
buf BUF1 (N558, N554);
nand NAND4 (N559, N558, N221, N4, N164);
or OR3 (N560, N550, N307, N474);
not NOT1 (N561, N552);
nor NOR3 (N562, N536, N333, N505);
nand NAND2 (N563, N562, N427);
and AND3 (N564, N557, N271, N297);
or OR3 (N565, N553, N379, N74);
xor XOR2 (N566, N535, N324);
not NOT1 (N567, N549);
buf BUF1 (N568, N560);
and AND4 (N569, N565, N517, N157, N40);
nand NAND2 (N570, N561, N118);
nand NAND3 (N571, N566, N500, N289);
or OR4 (N572, N559, N117, N174, N340);
not NOT1 (N573, N570);
buf BUF1 (N574, N567);
or OR2 (N575, N574, N49);
buf BUF1 (N576, N563);
not NOT1 (N577, N556);
and AND4 (N578, N512, N142, N486, N186);
and AND3 (N579, N575, N46, N117);
nor NOR4 (N580, N578, N408, N337, N562);
not NOT1 (N581, N569);
not NOT1 (N582, N573);
xor XOR2 (N583, N564, N299);
or OR4 (N584, N577, N168, N169, N3);
not NOT1 (N585, N572);
or OR3 (N586, N576, N396, N281);
buf BUF1 (N587, N568);
nor NOR3 (N588, N585, N537, N95);
buf BUF1 (N589, N583);
buf BUF1 (N590, N586);
or OR4 (N591, N579, N130, N6, N518);
and AND4 (N592, N589, N545, N390, N175);
not NOT1 (N593, N592);
and AND2 (N594, N588, N5);
nand NAND4 (N595, N582, N171, N514, N319);
nand NAND4 (N596, N584, N59, N238, N497);
nand NAND3 (N597, N571, N409, N149);
xor XOR2 (N598, N593, N142);
nand NAND2 (N599, N590, N558);
xor XOR2 (N600, N581, N344);
buf BUF1 (N601, N595);
and AND4 (N602, N600, N72, N531, N297);
xor XOR2 (N603, N602, N70);
not NOT1 (N604, N598);
or OR3 (N605, N603, N497, N454);
nand NAND4 (N606, N605, N19, N429, N176);
or OR4 (N607, N599, N344, N530, N372);
and AND2 (N608, N606, N220);
or OR2 (N609, N591, N103);
or OR4 (N610, N587, N579, N561, N247);
xor XOR2 (N611, N607, N67);
or OR4 (N612, N601, N132, N420, N165);
and AND3 (N613, N594, N440, N441);
xor XOR2 (N614, N611, N465);
nand NAND4 (N615, N614, N373, N74, N322);
and AND3 (N616, N604, N119, N211);
or OR2 (N617, N609, N31);
not NOT1 (N618, N613);
not NOT1 (N619, N608);
or OR2 (N620, N617, N84);
not NOT1 (N621, N620);
nor NOR3 (N622, N618, N39, N587);
not NOT1 (N623, N580);
and AND3 (N624, N619, N206, N76);
and AND2 (N625, N616, N352);
xor XOR2 (N626, N597, N388);
buf BUF1 (N627, N624);
not NOT1 (N628, N612);
buf BUF1 (N629, N615);
nor NOR4 (N630, N625, N354, N111, N28);
and AND2 (N631, N623, N408);
not NOT1 (N632, N628);
xor XOR2 (N633, N621, N105);
or OR4 (N634, N627, N60, N114, N231);
not NOT1 (N635, N631);
buf BUF1 (N636, N635);
nand NAND2 (N637, N634, N587);
not NOT1 (N638, N636);
nor NOR3 (N639, N626, N584, N476);
xor XOR2 (N640, N638, N606);
or OR2 (N641, N629, N595);
and AND2 (N642, N637, N500);
not NOT1 (N643, N633);
buf BUF1 (N644, N642);
nor NOR4 (N645, N596, N32, N550, N357);
nor NOR4 (N646, N643, N437, N282, N489);
not NOT1 (N647, N640);
or OR4 (N648, N647, N563, N404, N319);
buf BUF1 (N649, N622);
nand NAND3 (N650, N639, N124, N214);
buf BUF1 (N651, N641);
buf BUF1 (N652, N649);
or OR3 (N653, N644, N112, N495);
xor XOR2 (N654, N651, N281);
xor XOR2 (N655, N610, N424);
buf BUF1 (N656, N650);
buf BUF1 (N657, N656);
nand NAND3 (N658, N657, N572, N493);
or OR3 (N659, N655, N171, N101);
buf BUF1 (N660, N648);
xor XOR2 (N661, N654, N382);
buf BUF1 (N662, N660);
buf BUF1 (N663, N658);
nor NOR4 (N664, N659, N455, N618, N522);
not NOT1 (N665, N630);
and AND3 (N666, N663, N372, N397);
nand NAND2 (N667, N646, N198);
not NOT1 (N668, N645);
nand NAND3 (N669, N632, N291, N330);
buf BUF1 (N670, N666);
and AND3 (N671, N670, N19, N169);
and AND4 (N672, N661, N296, N272, N219);
and AND4 (N673, N669, N569, N503, N628);
and AND3 (N674, N662, N221, N355);
nand NAND3 (N675, N652, N157, N404);
xor XOR2 (N676, N668, N498);
nand NAND2 (N677, N672, N287);
xor XOR2 (N678, N673, N505);
nor NOR3 (N679, N653, N434, N532);
not NOT1 (N680, N679);
buf BUF1 (N681, N671);
nand NAND4 (N682, N664, N382, N607, N175);
buf BUF1 (N683, N680);
xor XOR2 (N684, N667, N376);
buf BUF1 (N685, N677);
nand NAND2 (N686, N674, N352);
and AND3 (N687, N684, N83, N551);
nor NOR4 (N688, N687, N138, N155, N357);
not NOT1 (N689, N686);
nor NOR4 (N690, N676, N36, N205, N119);
or OR4 (N691, N678, N194, N160, N206);
nor NOR3 (N692, N675, N145, N85);
nor NOR3 (N693, N665, N428, N49);
or OR3 (N694, N688, N79, N679);
xor XOR2 (N695, N693, N498);
not NOT1 (N696, N689);
not NOT1 (N697, N683);
or OR3 (N698, N692, N480, N242);
or OR2 (N699, N698, N407);
nand NAND4 (N700, N682, N220, N79, N647);
buf BUF1 (N701, N690);
buf BUF1 (N702, N691);
nor NOR4 (N703, N695, N503, N79, N242);
xor XOR2 (N704, N702, N260);
nor NOR2 (N705, N704, N336);
xor XOR2 (N706, N700, N429);
or OR4 (N707, N699, N314, N69, N258);
nor NOR4 (N708, N701, N680, N133, N162);
or OR3 (N709, N685, N391, N318);
nand NAND2 (N710, N696, N30);
not NOT1 (N711, N681);
buf BUF1 (N712, N694);
not NOT1 (N713, N697);
not NOT1 (N714, N709);
not NOT1 (N715, N711);
nor NOR4 (N716, N706, N193, N245, N310);
nand NAND3 (N717, N707, N82, N169);
nor NOR4 (N718, N717, N168, N180, N535);
buf BUF1 (N719, N708);
xor XOR2 (N720, N710, N372);
nor NOR2 (N721, N714, N532);
and AND3 (N722, N705, N670, N67);
nand NAND3 (N723, N715, N465, N605);
xor XOR2 (N724, N718, N292);
nand NAND4 (N725, N716, N383, N54, N69);
and AND3 (N726, N722, N11, N610);
and AND4 (N727, N720, N467, N717, N174);
buf BUF1 (N728, N713);
xor XOR2 (N729, N721, N26);
not NOT1 (N730, N725);
xor XOR2 (N731, N723, N526);
and AND3 (N732, N719, N577, N595);
xor XOR2 (N733, N726, N732);
buf BUF1 (N734, N171);
or OR2 (N735, N712, N504);
not NOT1 (N736, N724);
nand NAND2 (N737, N729, N569);
xor XOR2 (N738, N731, N686);
nand NAND4 (N739, N733, N578, N6, N55);
not NOT1 (N740, N703);
nor NOR4 (N741, N738, N207, N672, N330);
buf BUF1 (N742, N734);
not NOT1 (N743, N730);
xor XOR2 (N744, N728, N23);
nor NOR2 (N745, N727, N345);
or OR3 (N746, N744, N712, N349);
and AND3 (N747, N745, N649, N152);
nand NAND4 (N748, N737, N607, N566, N509);
xor XOR2 (N749, N748, N97);
or OR2 (N750, N740, N451);
nor NOR4 (N751, N743, N250, N401, N345);
buf BUF1 (N752, N750);
nand NAND2 (N753, N747, N555);
not NOT1 (N754, N753);
or OR3 (N755, N742, N744, N393);
and AND4 (N756, N739, N171, N740, N219);
or OR4 (N757, N755, N8, N591, N671);
xor XOR2 (N758, N749, N28);
buf BUF1 (N759, N746);
xor XOR2 (N760, N735, N698);
not NOT1 (N761, N756);
nand NAND2 (N762, N751, N327);
nor NOR3 (N763, N741, N187, N41);
buf BUF1 (N764, N762);
buf BUF1 (N765, N761);
nand NAND3 (N766, N758, N707, N540);
or OR4 (N767, N764, N362, N705, N580);
nand NAND2 (N768, N754, N603);
nor NOR4 (N769, N763, N30, N250, N405);
and AND4 (N770, N759, N489, N385, N23);
nor NOR4 (N771, N765, N33, N28, N386);
xor XOR2 (N772, N760, N605);
nor NOR2 (N773, N736, N473);
nor NOR3 (N774, N752, N525, N649);
nand NAND2 (N775, N774, N609);
or OR2 (N776, N772, N699);
or OR3 (N777, N770, N572, N18);
not NOT1 (N778, N771);
nor NOR4 (N779, N775, N80, N707, N750);
and AND3 (N780, N776, N519, N144);
nor NOR2 (N781, N766, N23);
or OR2 (N782, N757, N318);
buf BUF1 (N783, N773);
not NOT1 (N784, N778);
nand NAND4 (N785, N781, N214, N17, N242);
nor NOR3 (N786, N782, N603, N634);
and AND3 (N787, N777, N279, N583);
or OR3 (N788, N785, N227, N282);
or OR4 (N789, N767, N421, N512, N222);
nand NAND3 (N790, N787, N416, N653);
not NOT1 (N791, N779);
nor NOR4 (N792, N784, N480, N51, N426);
or OR4 (N793, N789, N208, N792, N541);
nand NAND3 (N794, N129, N49, N735);
xor XOR2 (N795, N783, N560);
xor XOR2 (N796, N768, N67);
and AND3 (N797, N793, N60, N586);
nand NAND3 (N798, N795, N213, N731);
buf BUF1 (N799, N797);
buf BUF1 (N800, N786);
xor XOR2 (N801, N800, N439);
nand NAND3 (N802, N791, N258, N613);
and AND2 (N803, N790, N74);
or OR4 (N804, N788, N121, N371, N350);
and AND3 (N805, N796, N253, N591);
xor XOR2 (N806, N798, N686);
buf BUF1 (N807, N803);
nand NAND4 (N808, N807, N432, N332, N269);
and AND2 (N809, N808, N220);
xor XOR2 (N810, N801, N454);
and AND3 (N811, N804, N219, N319);
buf BUF1 (N812, N769);
nor NOR2 (N813, N780, N408);
xor XOR2 (N814, N813, N47);
xor XOR2 (N815, N811, N35);
and AND3 (N816, N794, N685, N643);
not NOT1 (N817, N806);
buf BUF1 (N818, N810);
nand NAND4 (N819, N799, N458, N600, N689);
not NOT1 (N820, N802);
xor XOR2 (N821, N820, N589);
nand NAND3 (N822, N809, N792, N314);
or OR3 (N823, N814, N239, N295);
not NOT1 (N824, N821);
nor NOR4 (N825, N822, N574, N29, N144);
or OR3 (N826, N815, N142, N679);
buf BUF1 (N827, N819);
nand NAND4 (N828, N825, N682, N820, N790);
not NOT1 (N829, N827);
xor XOR2 (N830, N826, N228);
nor NOR4 (N831, N830, N465, N395, N113);
nor NOR3 (N832, N831, N459, N325);
xor XOR2 (N833, N828, N528);
buf BUF1 (N834, N818);
not NOT1 (N835, N832);
nor NOR4 (N836, N805, N158, N806, N474);
nand NAND3 (N837, N836, N5, N633);
xor XOR2 (N838, N833, N157);
xor XOR2 (N839, N812, N779);
not NOT1 (N840, N823);
xor XOR2 (N841, N824, N802);
and AND4 (N842, N816, N759, N760, N819);
not NOT1 (N843, N817);
not NOT1 (N844, N841);
and AND2 (N845, N840, N545);
or OR4 (N846, N845, N732, N255, N842);
and AND4 (N847, N738, N267, N733, N18);
xor XOR2 (N848, N844, N293);
buf BUF1 (N849, N847);
not NOT1 (N850, N848);
not NOT1 (N851, N829);
not NOT1 (N852, N835);
not NOT1 (N853, N838);
nand NAND3 (N854, N849, N634, N846);
and AND2 (N855, N415, N139);
xor XOR2 (N856, N852, N203);
buf BUF1 (N857, N850);
nand NAND4 (N858, N857, N812, N669, N641);
xor XOR2 (N859, N854, N851);
xor XOR2 (N860, N439, N817);
not NOT1 (N861, N859);
or OR3 (N862, N837, N489, N602);
xor XOR2 (N863, N862, N320);
and AND2 (N864, N858, N491);
and AND3 (N865, N864, N235, N841);
and AND4 (N866, N865, N844, N628, N547);
xor XOR2 (N867, N839, N826);
nand NAND4 (N868, N855, N439, N317, N603);
not NOT1 (N869, N843);
xor XOR2 (N870, N869, N77);
and AND4 (N871, N866, N358, N618, N649);
and AND4 (N872, N860, N120, N47, N744);
and AND4 (N873, N863, N478, N28, N60);
nor NOR2 (N874, N834, N350);
nor NOR2 (N875, N867, N288);
xor XOR2 (N876, N875, N81);
or OR2 (N877, N856, N201);
and AND4 (N878, N874, N151, N67, N875);
and AND3 (N879, N870, N21, N5);
nand NAND4 (N880, N876, N174, N182, N867);
and AND4 (N881, N871, N694, N668, N157);
xor XOR2 (N882, N881, N382);
nand NAND4 (N883, N872, N38, N541, N60);
not NOT1 (N884, N880);
nor NOR2 (N885, N884, N357);
xor XOR2 (N886, N879, N573);
buf BUF1 (N887, N868);
not NOT1 (N888, N887);
nand NAND2 (N889, N882, N278);
not NOT1 (N890, N889);
buf BUF1 (N891, N853);
or OR4 (N892, N888, N47, N50, N889);
nor NOR3 (N893, N883, N778, N422);
nand NAND3 (N894, N892, N386, N614);
not NOT1 (N895, N894);
and AND2 (N896, N886, N372);
xor XOR2 (N897, N877, N761);
nand NAND3 (N898, N878, N66, N189);
nand NAND3 (N899, N896, N442, N522);
nand NAND4 (N900, N890, N888, N804, N853);
not NOT1 (N901, N900);
and AND3 (N902, N901, N536, N540);
buf BUF1 (N903, N902);
and AND4 (N904, N861, N189, N861, N374);
not NOT1 (N905, N873);
nor NOR4 (N906, N905, N726, N154, N243);
buf BUF1 (N907, N897);
or OR2 (N908, N904, N863);
or OR3 (N909, N906, N550, N104);
nor NOR3 (N910, N893, N812, N579);
not NOT1 (N911, N885);
nand NAND2 (N912, N903, N615);
or OR3 (N913, N907, N905, N453);
buf BUF1 (N914, N912);
endmodule