// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22;

output N113,N119,N89,N108,N109,N115,N117,N120,N121,N122;

nand NAND4 (N23, N13, N19, N18, N10);
xor XOR2 (N24, N19, N8);
nand NAND2 (N25, N12, N19);
not NOT1 (N26, N17);
not NOT1 (N27, N3);
and AND3 (N28, N21, N21, N22);
buf BUF1 (N29, N25);
nand NAND2 (N30, N9, N3);
buf BUF1 (N31, N30);
nor NOR4 (N32, N2, N1, N30, N20);
or OR4 (N33, N30, N22, N11, N14);
or OR2 (N34, N1, N2);
xor XOR2 (N35, N32, N22);
and AND4 (N36, N35, N28, N7, N11);
nor NOR2 (N37, N21, N36);
xor XOR2 (N38, N22, N28);
xor XOR2 (N39, N23, N28);
nor NOR3 (N40, N38, N31, N11);
xor XOR2 (N41, N5, N12);
and AND4 (N42, N26, N17, N12, N28);
xor XOR2 (N43, N27, N23);
and AND3 (N44, N43, N34, N7);
and AND3 (N45, N5, N40, N37);
buf BUF1 (N46, N12);
or OR2 (N47, N38, N12);
nand NAND3 (N48, N46, N27, N36);
nor NOR3 (N49, N41, N13, N9);
or OR4 (N50, N33, N19, N4, N11);
nand NAND4 (N51, N24, N19, N13, N16);
or OR3 (N52, N50, N10, N15);
buf BUF1 (N53, N39);
xor XOR2 (N54, N42, N45);
and AND4 (N55, N11, N8, N31, N10);
xor XOR2 (N56, N49, N7);
nor NOR3 (N57, N44, N40, N33);
nand NAND2 (N58, N52, N25);
and AND4 (N59, N56, N44, N58, N19);
and AND2 (N60, N57, N47);
not NOT1 (N61, N8);
not NOT1 (N62, N42);
buf BUF1 (N63, N60);
not NOT1 (N64, N62);
nand NAND2 (N65, N51, N5);
buf BUF1 (N66, N29);
or OR2 (N67, N61, N53);
not NOT1 (N68, N41);
and AND4 (N69, N63, N4, N29, N54);
or OR2 (N70, N69, N6);
or OR4 (N71, N21, N28, N68, N58);
and AND4 (N72, N32, N32, N45, N48);
not NOT1 (N73, N14);
not NOT1 (N74, N72);
buf BUF1 (N75, N64);
or OR4 (N76, N55, N2, N74, N69);
nand NAND3 (N77, N10, N58, N18);
and AND3 (N78, N75, N61, N40);
or OR4 (N79, N76, N34, N56, N59);
and AND2 (N80, N20, N45);
or OR4 (N81, N73, N33, N51, N67);
xor XOR2 (N82, N78, N7);
not NOT1 (N83, N69);
nor NOR2 (N84, N81, N64);
xor XOR2 (N85, N84, N81);
nand NAND3 (N86, N80, N61, N58);
nor NOR2 (N87, N66, N23);
not NOT1 (N88, N86);
or OR3 (N89, N83, N9, N46);
or OR4 (N90, N85, N64, N59, N75);
not NOT1 (N91, N79);
nand NAND2 (N92, N91, N44);
buf BUF1 (N93, N65);
nand NAND2 (N94, N70, N71);
not NOT1 (N95, N92);
not NOT1 (N96, N90);
xor XOR2 (N97, N24, N6);
and AND4 (N98, N97, N28, N28, N14);
or OR2 (N99, N95, N57);
nand NAND3 (N100, N96, N95, N60);
nor NOR3 (N101, N88, N41, N48);
or OR4 (N102, N93, N54, N69, N101);
nand NAND3 (N103, N81, N82, N53);
or OR3 (N104, N10, N30, N61);
buf BUF1 (N105, N77);
or OR2 (N106, N98, N71);
xor XOR2 (N107, N94, N20);
buf BUF1 (N108, N107);
and AND4 (N109, N105, N103, N28, N10);
or OR2 (N110, N87, N86);
or OR3 (N111, N3, N27, N76);
nor NOR2 (N112, N111, N13);
xor XOR2 (N113, N104, N1);
not NOT1 (N114, N110);
xor XOR2 (N115, N112, N95);
xor XOR2 (N116, N102, N74);
nor NOR4 (N117, N99, N44, N26, N81);
not NOT1 (N118, N116);
buf BUF1 (N119, N100);
or OR4 (N120, N118, N53, N114, N47);
nand NAND4 (N121, N106, N45, N40, N26);
nand NAND2 (N122, N66, N8);
endmodule