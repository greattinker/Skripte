// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24;

output N3223,N3189,N3221,N3218,N3219,N3222,N3215,N3200,N3197,N3224;

nand NAND3 (N25, N11, N23, N14);
and AND4 (N26, N9, N2, N6, N13);
xor XOR2 (N27, N11, N16);
nand NAND3 (N28, N6, N3, N13);
xor XOR2 (N29, N11, N27);
or OR2 (N30, N19, N27);
not NOT1 (N31, N22);
nor NOR3 (N32, N4, N17, N5);
not NOT1 (N33, N14);
and AND3 (N34, N24, N24, N31);
nor NOR4 (N35, N9, N15, N7, N28);
and AND3 (N36, N15, N10, N31);
and AND2 (N37, N15, N17);
xor XOR2 (N38, N37, N2);
and AND3 (N39, N36, N25, N38);
nand NAND2 (N40, N37, N38);
not NOT1 (N41, N6);
and AND4 (N42, N35, N24, N25, N14);
or OR4 (N43, N39, N16, N10, N15);
nor NOR4 (N44, N34, N21, N27, N12);
nand NAND4 (N45, N30, N18, N12, N8);
and AND2 (N46, N32, N40);
nand NAND3 (N47, N37, N16, N39);
and AND2 (N48, N46, N2);
nand NAND4 (N49, N29, N27, N42, N1);
buf BUF1 (N50, N42);
nand NAND2 (N51, N48, N24);
or OR3 (N52, N43, N1, N27);
or OR4 (N53, N33, N9, N51, N30);
nand NAND4 (N54, N32, N48, N27, N31);
xor XOR2 (N55, N50, N11);
nor NOR4 (N56, N55, N29, N46, N4);
not NOT1 (N57, N45);
nor NOR2 (N58, N26, N53);
buf BUF1 (N59, N41);
or OR2 (N60, N14, N19);
xor XOR2 (N61, N56, N54);
or OR3 (N62, N56, N13, N37);
or OR2 (N63, N62, N41);
nand NAND4 (N64, N60, N19, N61, N34);
nand NAND4 (N65, N54, N51, N11, N53);
not NOT1 (N66, N44);
buf BUF1 (N67, N52);
and AND3 (N68, N59, N10, N15);
and AND4 (N69, N68, N55, N35, N33);
buf BUF1 (N70, N58);
or OR3 (N71, N49, N30, N44);
and AND4 (N72, N64, N13, N54, N2);
nor NOR4 (N73, N57, N6, N58, N4);
nand NAND3 (N74, N70, N15, N55);
nand NAND3 (N75, N65, N58, N56);
buf BUF1 (N76, N47);
not NOT1 (N77, N63);
xor XOR2 (N78, N76, N20);
nor NOR4 (N79, N75, N22, N51, N34);
buf BUF1 (N80, N66);
xor XOR2 (N81, N79, N34);
xor XOR2 (N82, N69, N29);
not NOT1 (N83, N72);
nor NOR2 (N84, N81, N62);
or OR2 (N85, N82, N74);
and AND3 (N86, N51, N61, N72);
buf BUF1 (N87, N73);
nand NAND3 (N88, N85, N14, N40);
nor NOR4 (N89, N78, N20, N7, N32);
xor XOR2 (N90, N67, N31);
nor NOR3 (N91, N80, N12, N52);
buf BUF1 (N92, N77);
buf BUF1 (N93, N89);
or OR3 (N94, N93, N87, N47);
nor NOR3 (N95, N16, N63, N61);
or OR4 (N96, N94, N5, N1, N67);
and AND3 (N97, N84, N85, N1);
and AND4 (N98, N92, N26, N51, N67);
nand NAND3 (N99, N97, N43, N19);
nor NOR4 (N100, N95, N55, N46, N22);
nand NAND2 (N101, N100, N39);
and AND2 (N102, N88, N54);
nand NAND3 (N103, N96, N101, N58);
xor XOR2 (N104, N13, N8);
not NOT1 (N105, N99);
nor NOR3 (N106, N86, N89, N14);
or OR3 (N107, N103, N24, N42);
not NOT1 (N108, N104);
not NOT1 (N109, N108);
xor XOR2 (N110, N71, N93);
xor XOR2 (N111, N106, N65);
xor XOR2 (N112, N90, N55);
nor NOR4 (N113, N112, N18, N22, N112);
nor NOR4 (N114, N111, N11, N10, N28);
or OR2 (N115, N91, N92);
and AND4 (N116, N109, N88, N84, N3);
or OR4 (N117, N115, N83, N63, N50);
not NOT1 (N118, N57);
buf BUF1 (N119, N98);
nand NAND4 (N120, N116, N47, N7, N37);
or OR3 (N121, N117, N58, N27);
xor XOR2 (N122, N118, N83);
xor XOR2 (N123, N105, N76);
xor XOR2 (N124, N110, N89);
nor NOR4 (N125, N121, N25, N5, N88);
or OR2 (N126, N107, N58);
or OR4 (N127, N124, N8, N41, N23);
nor NOR3 (N128, N114, N36, N20);
nor NOR2 (N129, N113, N113);
nand NAND2 (N130, N129, N125);
buf BUF1 (N131, N21);
nand NAND3 (N132, N122, N79, N8);
nor NOR4 (N133, N119, N17, N110, N9);
buf BUF1 (N134, N130);
xor XOR2 (N135, N127, N64);
or OR4 (N136, N128, N73, N12, N24);
nor NOR3 (N137, N134, N117, N136);
and AND3 (N138, N82, N20, N78);
nand NAND2 (N139, N126, N129);
buf BUF1 (N140, N133);
xor XOR2 (N141, N140, N68);
nor NOR3 (N142, N135, N42, N90);
xor XOR2 (N143, N139, N1);
or OR2 (N144, N138, N107);
not NOT1 (N145, N120);
and AND3 (N146, N141, N113, N43);
nor NOR2 (N147, N144, N43);
nand NAND4 (N148, N132, N1, N108, N69);
or OR2 (N149, N143, N4);
nand NAND3 (N150, N142, N119, N88);
xor XOR2 (N151, N147, N138);
or OR4 (N152, N151, N136, N88, N56);
and AND4 (N153, N123, N100, N104, N21);
xor XOR2 (N154, N146, N36);
buf BUF1 (N155, N137);
not NOT1 (N156, N131);
nor NOR2 (N157, N102, N104);
and AND3 (N158, N148, N34, N68);
buf BUF1 (N159, N154);
and AND2 (N160, N158, N137);
nand NAND3 (N161, N156, N48, N74);
and AND4 (N162, N160, N102, N61, N42);
or OR3 (N163, N145, N129, N23);
buf BUF1 (N164, N153);
buf BUF1 (N165, N152);
xor XOR2 (N166, N159, N14);
not NOT1 (N167, N161);
and AND4 (N168, N167, N156, N85, N97);
buf BUF1 (N169, N165);
buf BUF1 (N170, N164);
and AND4 (N171, N169, N128, N102, N121);
buf BUF1 (N172, N163);
nor NOR2 (N173, N168, N85);
buf BUF1 (N174, N149);
and AND2 (N175, N150, N145);
nand NAND3 (N176, N175, N52, N151);
xor XOR2 (N177, N174, N44);
or OR4 (N178, N170, N19, N67, N73);
nand NAND2 (N179, N173, N162);
and AND2 (N180, N67, N60);
not NOT1 (N181, N177);
nor NOR4 (N182, N179, N177, N43, N161);
nand NAND2 (N183, N171, N170);
not NOT1 (N184, N178);
nor NOR3 (N185, N176, N72, N169);
xor XOR2 (N186, N183, N31);
nand NAND2 (N187, N155, N180);
nand NAND2 (N188, N69, N135);
not NOT1 (N189, N185);
not NOT1 (N190, N157);
or OR3 (N191, N182, N190, N167);
and AND3 (N192, N134, N86, N125);
xor XOR2 (N193, N184, N35);
and AND3 (N194, N188, N64, N120);
xor XOR2 (N195, N172, N152);
and AND2 (N196, N195, N182);
xor XOR2 (N197, N193, N85);
nor NOR3 (N198, N194, N19, N159);
xor XOR2 (N199, N192, N22);
nor NOR2 (N200, N196, N183);
nor NOR3 (N201, N191, N84, N161);
not NOT1 (N202, N197);
nand NAND2 (N203, N202, N80);
or OR3 (N204, N199, N10, N71);
nand NAND3 (N205, N189, N38, N165);
and AND3 (N206, N204, N44, N159);
not NOT1 (N207, N200);
nor NOR2 (N208, N198, N91);
nand NAND3 (N209, N206, N167, N79);
xor XOR2 (N210, N166, N116);
nor NOR3 (N211, N209, N144, N77);
and AND4 (N212, N201, N91, N66, N121);
buf BUF1 (N213, N203);
or OR2 (N214, N205, N74);
not NOT1 (N215, N213);
nand NAND3 (N216, N212, N65, N95);
or OR3 (N217, N208, N13, N156);
nand NAND4 (N218, N217, N113, N130, N202);
nand NAND2 (N219, N187, N61);
xor XOR2 (N220, N216, N97);
not NOT1 (N221, N210);
not NOT1 (N222, N221);
not NOT1 (N223, N211);
and AND4 (N224, N214, N88, N63, N47);
nand NAND4 (N225, N223, N106, N97, N110);
xor XOR2 (N226, N218, N206);
and AND4 (N227, N220, N133, N144, N15);
and AND3 (N228, N215, N93, N16);
not NOT1 (N229, N186);
nand NAND2 (N230, N228, N69);
xor XOR2 (N231, N207, N186);
or OR4 (N232, N229, N77, N138, N208);
xor XOR2 (N233, N222, N81);
and AND2 (N234, N226, N33);
buf BUF1 (N235, N225);
not NOT1 (N236, N227);
nor NOR4 (N237, N230, N207, N121, N61);
nand NAND3 (N238, N234, N155, N176);
nor NOR2 (N239, N224, N18);
and AND4 (N240, N238, N169, N234, N183);
nand NAND4 (N241, N181, N58, N16, N18);
nor NOR4 (N242, N233, N26, N32, N32);
xor XOR2 (N243, N241, N137);
buf BUF1 (N244, N236);
and AND2 (N245, N239, N104);
and AND3 (N246, N242, N176, N161);
buf BUF1 (N247, N243);
buf BUF1 (N248, N219);
buf BUF1 (N249, N248);
nand NAND3 (N250, N244, N225, N185);
or OR4 (N251, N247, N148, N199, N149);
or OR4 (N252, N240, N43, N133, N105);
nand NAND2 (N253, N251, N73);
buf BUF1 (N254, N252);
or OR4 (N255, N237, N25, N247, N76);
and AND3 (N256, N245, N223, N136);
nor NOR2 (N257, N231, N186);
nand NAND4 (N258, N254, N89, N202, N109);
nor NOR2 (N259, N249, N38);
xor XOR2 (N260, N235, N6);
xor XOR2 (N261, N258, N216);
nand NAND2 (N262, N246, N75);
nor NOR2 (N263, N232, N102);
not NOT1 (N264, N256);
not NOT1 (N265, N257);
and AND4 (N266, N259, N15, N175, N124);
buf BUF1 (N267, N264);
nand NAND3 (N268, N255, N209, N28);
not NOT1 (N269, N253);
buf BUF1 (N270, N266);
not NOT1 (N271, N250);
xor XOR2 (N272, N260, N135);
not NOT1 (N273, N272);
xor XOR2 (N274, N273, N80);
xor XOR2 (N275, N262, N182);
buf BUF1 (N276, N265);
and AND2 (N277, N276, N180);
nand NAND2 (N278, N275, N23);
xor XOR2 (N279, N271, N182);
buf BUF1 (N280, N277);
buf BUF1 (N281, N279);
xor XOR2 (N282, N263, N121);
xor XOR2 (N283, N282, N218);
nor NOR4 (N284, N268, N119, N65, N117);
not NOT1 (N285, N269);
nor NOR3 (N286, N270, N202, N6);
nor NOR2 (N287, N274, N201);
nor NOR4 (N288, N285, N258, N64, N172);
nand NAND4 (N289, N288, N247, N31, N255);
and AND3 (N290, N261, N17, N204);
not NOT1 (N291, N284);
not NOT1 (N292, N278);
buf BUF1 (N293, N283);
and AND2 (N294, N291, N176);
xor XOR2 (N295, N281, N107);
nand NAND2 (N296, N287, N141);
or OR2 (N297, N295, N53);
xor XOR2 (N298, N290, N107);
xor XOR2 (N299, N267, N249);
or OR3 (N300, N280, N267, N6);
and AND3 (N301, N297, N134, N233);
nand NAND4 (N302, N286, N48, N240, N211);
and AND3 (N303, N296, N102, N249);
xor XOR2 (N304, N303, N59);
or OR4 (N305, N293, N140, N272, N211);
buf BUF1 (N306, N301);
not NOT1 (N307, N302);
buf BUF1 (N308, N300);
nor NOR2 (N309, N308, N284);
buf BUF1 (N310, N289);
nand NAND2 (N311, N305, N130);
nor NOR4 (N312, N310, N33, N48, N201);
or OR2 (N313, N306, N263);
not NOT1 (N314, N307);
buf BUF1 (N315, N292);
or OR4 (N316, N309, N163, N169, N156);
buf BUF1 (N317, N312);
xor XOR2 (N318, N298, N152);
not NOT1 (N319, N318);
nor NOR4 (N320, N311, N161, N23, N242);
xor XOR2 (N321, N320, N119);
or OR4 (N322, N321, N53, N121, N280);
not NOT1 (N323, N316);
buf BUF1 (N324, N319);
xor XOR2 (N325, N314, N232);
and AND3 (N326, N322, N169, N307);
nand NAND3 (N327, N323, N106, N117);
xor XOR2 (N328, N326, N125);
and AND2 (N329, N324, N285);
or OR2 (N330, N313, N215);
xor XOR2 (N331, N328, N113);
or OR3 (N332, N315, N155, N276);
nand NAND4 (N333, N299, N277, N275, N148);
or OR4 (N334, N332, N192, N261, N5);
buf BUF1 (N335, N325);
xor XOR2 (N336, N304, N269);
or OR4 (N337, N330, N81, N29, N106);
and AND2 (N338, N335, N112);
not NOT1 (N339, N338);
nand NAND3 (N340, N329, N47, N175);
xor XOR2 (N341, N339, N95);
or OR2 (N342, N340, N233);
and AND3 (N343, N331, N281, N117);
or OR3 (N344, N294, N167, N121);
nand NAND4 (N345, N344, N136, N312, N117);
nor NOR3 (N346, N333, N270, N110);
and AND2 (N347, N317, N242);
xor XOR2 (N348, N345, N141);
xor XOR2 (N349, N348, N273);
nor NOR2 (N350, N349, N163);
not NOT1 (N351, N336);
buf BUF1 (N352, N342);
or OR3 (N353, N351, N234, N142);
nor NOR3 (N354, N337, N227, N303);
or OR3 (N355, N352, N314, N110);
not NOT1 (N356, N353);
not NOT1 (N357, N327);
and AND3 (N358, N347, N194, N158);
nand NAND4 (N359, N341, N329, N88, N241);
xor XOR2 (N360, N358, N242);
and AND3 (N361, N354, N229, N41);
not NOT1 (N362, N355);
nand NAND4 (N363, N334, N165, N161, N224);
or OR4 (N364, N359, N243, N361, N248);
nor NOR2 (N365, N121, N275);
nor NOR4 (N366, N343, N329, N85, N309);
nand NAND3 (N367, N350, N91, N188);
nor NOR2 (N368, N357, N316);
nand NAND2 (N369, N356, N46);
buf BUF1 (N370, N366);
and AND4 (N371, N370, N73, N199, N210);
nor NOR3 (N372, N364, N134, N298);
not NOT1 (N373, N362);
and AND3 (N374, N360, N351, N294);
not NOT1 (N375, N368);
nor NOR3 (N376, N375, N71, N126);
xor XOR2 (N377, N374, N278);
buf BUF1 (N378, N372);
buf BUF1 (N379, N376);
and AND4 (N380, N365, N337, N24, N164);
not NOT1 (N381, N369);
nand NAND3 (N382, N367, N123, N278);
or OR3 (N383, N382, N77, N262);
xor XOR2 (N384, N377, N325);
nand NAND2 (N385, N363, N373);
buf BUF1 (N386, N56);
buf BUF1 (N387, N380);
buf BUF1 (N388, N378);
xor XOR2 (N389, N385, N323);
or OR2 (N390, N389, N294);
or OR4 (N391, N386, N183, N43, N204);
nand NAND2 (N392, N346, N340);
not NOT1 (N393, N383);
buf BUF1 (N394, N390);
or OR2 (N395, N394, N319);
buf BUF1 (N396, N395);
nor NOR4 (N397, N371, N92, N236, N219);
not NOT1 (N398, N381);
nor NOR3 (N399, N396, N398, N380);
or OR3 (N400, N381, N223, N362);
nand NAND2 (N401, N384, N34);
buf BUF1 (N402, N399);
or OR4 (N403, N391, N24, N175, N127);
not NOT1 (N404, N400);
buf BUF1 (N405, N404);
nand NAND4 (N406, N402, N351, N114, N190);
buf BUF1 (N407, N397);
not NOT1 (N408, N392);
buf BUF1 (N409, N405);
nand NAND3 (N410, N387, N262, N201);
nor NOR4 (N411, N409, N285, N216, N295);
not NOT1 (N412, N408);
and AND4 (N413, N388, N380, N31, N115);
not NOT1 (N414, N410);
nand NAND3 (N415, N413, N313, N107);
buf BUF1 (N416, N412);
or OR4 (N417, N407, N193, N47, N365);
buf BUF1 (N418, N401);
or OR2 (N419, N403, N153);
not NOT1 (N420, N415);
xor XOR2 (N421, N416, N59);
buf BUF1 (N422, N414);
buf BUF1 (N423, N418);
nand NAND4 (N424, N423, N46, N352, N41);
not NOT1 (N425, N379);
nand NAND2 (N426, N424, N245);
or OR2 (N427, N419, N107);
xor XOR2 (N428, N427, N71);
and AND2 (N429, N406, N99);
nand NAND4 (N430, N393, N22, N150, N175);
and AND4 (N431, N417, N307, N385, N153);
and AND4 (N432, N422, N341, N168, N251);
or OR4 (N433, N432, N134, N49, N2);
buf BUF1 (N434, N430);
xor XOR2 (N435, N420, N254);
nand NAND2 (N436, N426, N358);
and AND4 (N437, N429, N350, N14, N166);
nand NAND4 (N438, N421, N199, N387, N79);
and AND2 (N439, N437, N323);
and AND3 (N440, N436, N362, N125);
buf BUF1 (N441, N428);
and AND2 (N442, N434, N371);
buf BUF1 (N443, N425);
and AND4 (N444, N431, N57, N260, N381);
not NOT1 (N445, N442);
not NOT1 (N446, N439);
or OR2 (N447, N435, N288);
nor NOR4 (N448, N411, N123, N236, N325);
nand NAND2 (N449, N444, N402);
and AND4 (N450, N449, N214, N350, N62);
xor XOR2 (N451, N440, N374);
nor NOR2 (N452, N441, N436);
or OR3 (N453, N443, N283, N112);
nor NOR3 (N454, N446, N258, N363);
nor NOR4 (N455, N453, N72, N384, N76);
nand NAND2 (N456, N438, N406);
nor NOR2 (N457, N454, N98);
not NOT1 (N458, N450);
nor NOR2 (N459, N447, N457);
not NOT1 (N460, N272);
nor NOR3 (N461, N451, N179, N429);
nor NOR2 (N462, N461, N365);
nor NOR2 (N463, N456, N346);
nand NAND3 (N464, N463, N166, N210);
nand NAND3 (N465, N458, N144, N141);
or OR2 (N466, N464, N232);
buf BUF1 (N467, N466);
or OR3 (N468, N433, N3, N329);
and AND3 (N469, N455, N328, N69);
nor NOR2 (N470, N468, N382);
or OR4 (N471, N452, N364, N93, N449);
not NOT1 (N472, N460);
or OR2 (N473, N459, N91);
not NOT1 (N474, N472);
buf BUF1 (N475, N467);
and AND4 (N476, N471, N83, N177, N302);
nor NOR4 (N477, N469, N19, N272, N149);
or OR2 (N478, N445, N27);
buf BUF1 (N479, N478);
and AND3 (N480, N462, N322, N184);
and AND4 (N481, N475, N126, N318, N459);
or OR4 (N482, N474, N346, N343, N203);
nor NOR2 (N483, N482, N275);
and AND2 (N484, N480, N403);
not NOT1 (N485, N479);
and AND4 (N486, N476, N328, N389, N215);
and AND3 (N487, N465, N411, N422);
nor NOR3 (N488, N473, N367, N310);
and AND3 (N489, N483, N313, N276);
buf BUF1 (N490, N484);
or OR4 (N491, N489, N10, N451, N421);
or OR2 (N492, N487, N416);
xor XOR2 (N493, N490, N207);
xor XOR2 (N494, N481, N319);
and AND2 (N495, N470, N153);
and AND4 (N496, N491, N246, N206, N487);
nor NOR3 (N497, N485, N303, N414);
nand NAND3 (N498, N486, N441, N141);
and AND2 (N499, N494, N435);
and AND4 (N500, N448, N277, N248, N312);
buf BUF1 (N501, N495);
xor XOR2 (N502, N501, N472);
buf BUF1 (N503, N477);
or OR3 (N504, N492, N222, N351);
not NOT1 (N505, N493);
not NOT1 (N506, N502);
nand NAND4 (N507, N499, N194, N469, N264);
xor XOR2 (N508, N507, N90);
and AND4 (N509, N505, N347, N254, N364);
not NOT1 (N510, N506);
nand NAND3 (N511, N488, N178, N158);
xor XOR2 (N512, N508, N339);
xor XOR2 (N513, N497, N34);
not NOT1 (N514, N503);
nand NAND2 (N515, N498, N425);
and AND2 (N516, N509, N509);
buf BUF1 (N517, N510);
nand NAND2 (N518, N513, N116);
buf BUF1 (N519, N512);
or OR4 (N520, N511, N359, N454, N49);
nor NOR4 (N521, N520, N225, N160, N18);
or OR2 (N522, N516, N43);
and AND2 (N523, N519, N454);
nor NOR2 (N524, N515, N143);
not NOT1 (N525, N514);
not NOT1 (N526, N521);
nand NAND2 (N527, N526, N33);
nor NOR2 (N528, N500, N363);
and AND3 (N529, N496, N64, N212);
or OR4 (N530, N528, N327, N370, N333);
not NOT1 (N531, N522);
and AND4 (N532, N524, N74, N353, N193);
buf BUF1 (N533, N517);
and AND4 (N534, N527, N314, N371, N338);
nand NAND4 (N535, N532, N531, N379, N364);
nor NOR4 (N536, N230, N460, N408, N317);
buf BUF1 (N537, N518);
not NOT1 (N538, N530);
not NOT1 (N539, N538);
xor XOR2 (N540, N539, N526);
xor XOR2 (N541, N533, N162);
or OR4 (N542, N540, N464, N272, N494);
nor NOR3 (N543, N525, N369, N320);
not NOT1 (N544, N534);
nor NOR2 (N545, N542, N107);
and AND3 (N546, N543, N103, N60);
and AND3 (N547, N544, N524, N251);
buf BUF1 (N548, N535);
nand NAND2 (N549, N545, N87);
xor XOR2 (N550, N547, N350);
xor XOR2 (N551, N549, N92);
or OR4 (N552, N550, N363, N38, N418);
nor NOR3 (N553, N523, N314, N137);
or OR3 (N554, N546, N26, N342);
or OR2 (N555, N504, N107);
and AND4 (N556, N541, N538, N540, N320);
and AND4 (N557, N536, N313, N330, N332);
or OR4 (N558, N556, N217, N526, N192);
nor NOR2 (N559, N537, N415);
buf BUF1 (N560, N557);
and AND3 (N561, N553, N468, N38);
and AND2 (N562, N548, N479);
or OR2 (N563, N551, N90);
or OR2 (N564, N554, N549);
nand NAND3 (N565, N559, N176, N8);
or OR4 (N566, N561, N554, N446, N447);
not NOT1 (N567, N565);
or OR2 (N568, N560, N90);
or OR2 (N569, N552, N315);
or OR2 (N570, N562, N234);
nand NAND3 (N571, N567, N334, N282);
not NOT1 (N572, N566);
nor NOR3 (N573, N570, N24, N453);
not NOT1 (N574, N572);
not NOT1 (N575, N571);
buf BUF1 (N576, N568);
nand NAND3 (N577, N573, N402, N231);
nand NAND3 (N578, N569, N233, N520);
xor XOR2 (N579, N577, N451);
or OR4 (N580, N578, N224, N204, N313);
and AND2 (N581, N555, N53);
nor NOR3 (N582, N581, N160, N205);
and AND3 (N583, N576, N290, N368);
nand NAND3 (N584, N579, N7, N549);
nand NAND2 (N585, N558, N348);
nor NOR3 (N586, N564, N159, N125);
not NOT1 (N587, N582);
nor NOR4 (N588, N574, N468, N321, N118);
not NOT1 (N589, N575);
xor XOR2 (N590, N587, N109);
nand NAND2 (N591, N580, N576);
and AND4 (N592, N529, N153, N118, N484);
nand NAND2 (N593, N563, N273);
buf BUF1 (N594, N584);
nor NOR4 (N595, N590, N125, N315, N333);
buf BUF1 (N596, N586);
xor XOR2 (N597, N589, N258);
nand NAND2 (N598, N596, N568);
xor XOR2 (N599, N598, N268);
or OR4 (N600, N595, N38, N511, N117);
or OR3 (N601, N588, N499, N45);
and AND4 (N602, N591, N554, N589, N457);
or OR4 (N603, N594, N133, N255, N548);
nor NOR3 (N604, N599, N161, N80);
xor XOR2 (N605, N601, N296);
xor XOR2 (N606, N605, N359);
or OR2 (N607, N592, N346);
not NOT1 (N608, N607);
not NOT1 (N609, N593);
or OR2 (N610, N609, N159);
nand NAND4 (N611, N600, N385, N307, N584);
xor XOR2 (N612, N606, N246);
and AND2 (N613, N608, N155);
buf BUF1 (N614, N602);
nand NAND4 (N615, N613, N590, N410, N296);
nor NOR3 (N616, N612, N565, N162);
nor NOR3 (N617, N610, N217, N550);
buf BUF1 (N618, N585);
xor XOR2 (N619, N614, N577);
xor XOR2 (N620, N617, N458);
and AND3 (N621, N615, N219, N123);
nand NAND2 (N622, N603, N177);
or OR2 (N623, N597, N218);
nor NOR4 (N624, N619, N206, N300, N489);
not NOT1 (N625, N622);
nand NAND2 (N626, N616, N94);
or OR4 (N627, N625, N237, N608, N82);
xor XOR2 (N628, N621, N345);
not NOT1 (N629, N611);
nand NAND2 (N630, N583, N272);
xor XOR2 (N631, N629, N134);
not NOT1 (N632, N620);
xor XOR2 (N633, N604, N10);
not NOT1 (N634, N631);
and AND2 (N635, N632, N236);
nand NAND4 (N636, N624, N310, N626, N206);
or OR2 (N637, N44, N77);
and AND2 (N638, N634, N452);
xor XOR2 (N639, N638, N349);
or OR3 (N640, N627, N70, N460);
not NOT1 (N641, N640);
buf BUF1 (N642, N639);
and AND4 (N643, N630, N41, N623, N508);
buf BUF1 (N644, N246);
xor XOR2 (N645, N633, N557);
or OR2 (N646, N641, N619);
xor XOR2 (N647, N635, N421);
nor NOR3 (N648, N643, N599, N644);
xor XOR2 (N649, N542, N458);
nor NOR4 (N650, N637, N6, N341, N265);
not NOT1 (N651, N645);
xor XOR2 (N652, N650, N200);
and AND3 (N653, N618, N152, N132);
buf BUF1 (N654, N646);
and AND4 (N655, N642, N513, N504, N566);
nand NAND3 (N656, N655, N572, N615);
xor XOR2 (N657, N653, N508);
nand NAND4 (N658, N648, N441, N11, N336);
nand NAND4 (N659, N636, N267, N434, N377);
buf BUF1 (N660, N659);
buf BUF1 (N661, N647);
buf BUF1 (N662, N652);
nor NOR4 (N663, N658, N77, N291, N80);
xor XOR2 (N664, N649, N37);
nand NAND3 (N665, N628, N426, N590);
nand NAND4 (N666, N656, N547, N650, N635);
nand NAND4 (N667, N663, N385, N99, N657);
nand NAND4 (N668, N566, N277, N455, N15);
not NOT1 (N669, N666);
and AND2 (N670, N665, N68);
nor NOR2 (N671, N662, N619);
or OR4 (N672, N667, N50, N574, N591);
buf BUF1 (N673, N670);
not NOT1 (N674, N664);
and AND2 (N675, N669, N128);
nor NOR4 (N676, N675, N580, N98, N365);
nor NOR4 (N677, N674, N586, N283, N27);
buf BUF1 (N678, N673);
or OR4 (N679, N651, N466, N219, N663);
not NOT1 (N680, N661);
and AND2 (N681, N672, N514);
and AND2 (N682, N668, N524);
nor NOR2 (N683, N654, N411);
xor XOR2 (N684, N660, N609);
nor NOR4 (N685, N679, N334, N344, N3);
and AND3 (N686, N676, N191, N52);
or OR3 (N687, N671, N651, N620);
nor NOR2 (N688, N687, N520);
not NOT1 (N689, N684);
and AND4 (N690, N688, N463, N368, N574);
nand NAND2 (N691, N681, N174);
and AND3 (N692, N690, N162, N565);
and AND2 (N693, N683, N526);
and AND2 (N694, N693, N157);
or OR4 (N695, N677, N562, N535, N89);
xor XOR2 (N696, N695, N157);
and AND3 (N697, N692, N145, N503);
and AND3 (N698, N686, N358, N511);
not NOT1 (N699, N696);
nor NOR4 (N700, N680, N147, N477, N170);
nor NOR2 (N701, N691, N124);
nand NAND3 (N702, N700, N611, N504);
nor NOR4 (N703, N699, N489, N27, N574);
not NOT1 (N704, N701);
not NOT1 (N705, N703);
not NOT1 (N706, N702);
buf BUF1 (N707, N685);
buf BUF1 (N708, N707);
and AND2 (N709, N698, N200);
or OR4 (N710, N682, N81, N21, N420);
nand NAND2 (N711, N689, N43);
nand NAND4 (N712, N694, N344, N128, N245);
xor XOR2 (N713, N697, N356);
and AND4 (N714, N713, N138, N77, N231);
buf BUF1 (N715, N706);
nand NAND3 (N716, N710, N35, N699);
and AND3 (N717, N704, N503, N3);
and AND2 (N718, N715, N602);
buf BUF1 (N719, N714);
nand NAND4 (N720, N678, N597, N318, N192);
or OR2 (N721, N716, N319);
nand NAND4 (N722, N719, N417, N553, N260);
or OR3 (N723, N720, N266, N438);
nand NAND3 (N724, N723, N428, N257);
nand NAND3 (N725, N722, N579, N209);
or OR2 (N726, N708, N705);
or OR4 (N727, N152, N103, N514, N123);
not NOT1 (N728, N709);
nand NAND3 (N729, N727, N408, N639);
not NOT1 (N730, N724);
nand NAND4 (N731, N711, N714, N550, N205);
or OR3 (N732, N725, N93, N658);
or OR2 (N733, N712, N97);
buf BUF1 (N734, N718);
or OR3 (N735, N728, N688, N667);
or OR3 (N736, N732, N102, N675);
buf BUF1 (N737, N721);
xor XOR2 (N738, N726, N497);
buf BUF1 (N739, N729);
not NOT1 (N740, N730);
xor XOR2 (N741, N735, N446);
nor NOR4 (N742, N739, N98, N640, N261);
buf BUF1 (N743, N717);
nor NOR4 (N744, N736, N347, N149, N419);
buf BUF1 (N745, N742);
xor XOR2 (N746, N745, N385);
not NOT1 (N747, N731);
nor NOR2 (N748, N743, N532);
xor XOR2 (N749, N734, N705);
not NOT1 (N750, N747);
not NOT1 (N751, N733);
buf BUF1 (N752, N740);
xor XOR2 (N753, N738, N706);
xor XOR2 (N754, N753, N431);
not NOT1 (N755, N750);
xor XOR2 (N756, N754, N214);
xor XOR2 (N757, N751, N198);
not NOT1 (N758, N748);
nor NOR4 (N759, N749, N410, N415, N502);
not NOT1 (N760, N741);
buf BUF1 (N761, N752);
not NOT1 (N762, N757);
or OR3 (N763, N756, N550, N141);
not NOT1 (N764, N737);
and AND2 (N765, N758, N570);
not NOT1 (N766, N746);
nor NOR4 (N767, N763, N592, N436, N207);
xor XOR2 (N768, N767, N369);
nor NOR4 (N769, N761, N588, N69, N256);
nor NOR2 (N770, N759, N441);
and AND4 (N771, N760, N529, N334, N44);
and AND2 (N772, N764, N651);
nor NOR4 (N773, N766, N744, N354, N443);
xor XOR2 (N774, N125, N141);
and AND3 (N775, N755, N76, N710);
nor NOR3 (N776, N771, N217, N51);
xor XOR2 (N777, N774, N702);
xor XOR2 (N778, N769, N662);
nand NAND2 (N779, N772, N735);
not NOT1 (N780, N779);
nand NAND3 (N781, N780, N708, N669);
xor XOR2 (N782, N781, N470);
or OR2 (N783, N765, N681);
nand NAND2 (N784, N782, N215);
buf BUF1 (N785, N778);
xor XOR2 (N786, N776, N576);
and AND2 (N787, N762, N307);
not NOT1 (N788, N787);
not NOT1 (N789, N786);
buf BUF1 (N790, N789);
xor XOR2 (N791, N788, N698);
nand NAND3 (N792, N768, N118, N150);
not NOT1 (N793, N783);
and AND4 (N794, N770, N566, N470, N668);
buf BUF1 (N795, N791);
and AND2 (N796, N777, N790);
nand NAND2 (N797, N253, N767);
and AND2 (N798, N797, N168);
not NOT1 (N799, N795);
and AND3 (N800, N785, N706, N26);
buf BUF1 (N801, N793);
and AND2 (N802, N773, N411);
buf BUF1 (N803, N802);
nand NAND2 (N804, N792, N774);
buf BUF1 (N805, N798);
not NOT1 (N806, N799);
and AND4 (N807, N801, N534, N755, N145);
nor NOR3 (N808, N775, N395, N362);
or OR2 (N809, N807, N389);
nand NAND2 (N810, N796, N123);
not NOT1 (N811, N794);
nor NOR3 (N812, N809, N70, N301);
or OR4 (N813, N806, N405, N205, N338);
not NOT1 (N814, N804);
buf BUF1 (N815, N805);
not NOT1 (N816, N800);
buf BUF1 (N817, N811);
not NOT1 (N818, N808);
not NOT1 (N819, N813);
xor XOR2 (N820, N819, N558);
nor NOR4 (N821, N812, N554, N621, N542);
nand NAND4 (N822, N814, N557, N587, N682);
nand NAND3 (N823, N815, N10, N449);
nand NAND3 (N824, N784, N86, N106);
buf BUF1 (N825, N817);
nand NAND3 (N826, N824, N600, N166);
not NOT1 (N827, N810);
nand NAND3 (N828, N818, N745, N664);
or OR3 (N829, N821, N683, N95);
nand NAND2 (N830, N826, N388);
buf BUF1 (N831, N827);
xor XOR2 (N832, N820, N381);
not NOT1 (N833, N831);
not NOT1 (N834, N830);
nand NAND4 (N835, N822, N124, N6, N673);
nor NOR4 (N836, N828, N456, N352, N554);
nor NOR2 (N837, N836, N54);
nor NOR2 (N838, N803, N677);
buf BUF1 (N839, N823);
nand NAND2 (N840, N835, N631);
xor XOR2 (N841, N829, N351);
buf BUF1 (N842, N834);
or OR4 (N843, N842, N284, N518, N442);
buf BUF1 (N844, N843);
xor XOR2 (N845, N840, N742);
not NOT1 (N846, N825);
nand NAND2 (N847, N832, N154);
not NOT1 (N848, N841);
and AND4 (N849, N845, N387, N63, N238);
buf BUF1 (N850, N849);
or OR3 (N851, N850, N466, N123);
nand NAND3 (N852, N846, N817, N721);
xor XOR2 (N853, N847, N58);
buf BUF1 (N854, N816);
or OR4 (N855, N839, N460, N596, N535);
or OR2 (N856, N854, N714);
buf BUF1 (N857, N853);
nor NOR3 (N858, N856, N826, N363);
not NOT1 (N859, N855);
not NOT1 (N860, N837);
not NOT1 (N861, N858);
and AND3 (N862, N848, N742, N578);
xor XOR2 (N863, N859, N830);
nand NAND3 (N864, N862, N615, N759);
xor XOR2 (N865, N863, N704);
not NOT1 (N866, N851);
nand NAND3 (N867, N857, N437, N277);
xor XOR2 (N868, N861, N133);
or OR4 (N869, N865, N163, N91, N590);
and AND3 (N870, N833, N198, N454);
or OR4 (N871, N860, N228, N126, N16);
nand NAND4 (N872, N871, N541, N756, N365);
nand NAND4 (N873, N838, N18, N345, N678);
or OR2 (N874, N873, N306);
nor NOR3 (N875, N869, N721, N240);
nor NOR2 (N876, N868, N255);
buf BUF1 (N877, N867);
not NOT1 (N878, N872);
nand NAND3 (N879, N870, N579, N560);
buf BUF1 (N880, N864);
not NOT1 (N881, N875);
and AND3 (N882, N852, N106, N245);
not NOT1 (N883, N866);
and AND4 (N884, N876, N253, N153, N417);
and AND4 (N885, N878, N831, N780, N243);
nand NAND4 (N886, N877, N162, N867, N54);
buf BUF1 (N887, N886);
nor NOR3 (N888, N887, N342, N428);
or OR3 (N889, N881, N392, N186);
or OR4 (N890, N882, N90, N547, N716);
buf BUF1 (N891, N888);
buf BUF1 (N892, N885);
and AND2 (N893, N892, N841);
nor NOR4 (N894, N893, N719, N230, N488);
or OR3 (N895, N879, N700, N123);
and AND3 (N896, N880, N376, N882);
and AND3 (N897, N891, N216, N586);
nor NOR4 (N898, N889, N791, N472, N86);
not NOT1 (N899, N897);
buf BUF1 (N900, N896);
or OR4 (N901, N874, N387, N698, N485);
and AND2 (N902, N901, N529);
xor XOR2 (N903, N895, N193);
and AND4 (N904, N890, N437, N550, N798);
buf BUF1 (N905, N898);
buf BUF1 (N906, N899);
or OR2 (N907, N883, N100);
not NOT1 (N908, N902);
buf BUF1 (N909, N900);
buf BUF1 (N910, N844);
and AND3 (N911, N906, N655, N783);
not NOT1 (N912, N911);
not NOT1 (N913, N912);
xor XOR2 (N914, N894, N697);
not NOT1 (N915, N913);
buf BUF1 (N916, N903);
or OR4 (N917, N904, N726, N91, N22);
buf BUF1 (N918, N905);
nor NOR3 (N919, N884, N626, N486);
and AND4 (N920, N908, N445, N215, N722);
not NOT1 (N921, N909);
buf BUF1 (N922, N920);
nand NAND2 (N923, N915, N243);
xor XOR2 (N924, N919, N443);
nand NAND4 (N925, N921, N713, N253, N114);
buf BUF1 (N926, N923);
not NOT1 (N927, N916);
or OR4 (N928, N917, N438, N482, N602);
or OR3 (N929, N924, N70, N157);
and AND3 (N930, N926, N858, N15);
buf BUF1 (N931, N928);
nand NAND4 (N932, N914, N806, N586, N165);
buf BUF1 (N933, N918);
and AND3 (N934, N929, N762, N134);
nor NOR4 (N935, N925, N10, N912, N889);
nor NOR3 (N936, N934, N682, N857);
xor XOR2 (N937, N922, N68);
or OR3 (N938, N907, N526, N878);
buf BUF1 (N939, N910);
nand NAND2 (N940, N937, N540);
or OR2 (N941, N939, N332);
nor NOR4 (N942, N931, N524, N88, N459);
and AND4 (N943, N935, N736, N374, N838);
and AND4 (N944, N943, N27, N457, N641);
nand NAND3 (N945, N938, N793, N925);
and AND3 (N946, N940, N367, N260);
buf BUF1 (N947, N946);
xor XOR2 (N948, N942, N142);
and AND2 (N949, N930, N704);
nor NOR4 (N950, N949, N579, N210, N189);
not NOT1 (N951, N947);
nor NOR2 (N952, N951, N262);
not NOT1 (N953, N944);
nor NOR4 (N954, N936, N538, N880, N680);
xor XOR2 (N955, N941, N903);
xor XOR2 (N956, N952, N638);
not NOT1 (N957, N932);
not NOT1 (N958, N927);
buf BUF1 (N959, N954);
or OR2 (N960, N948, N951);
nor NOR3 (N961, N958, N701, N11);
nand NAND2 (N962, N957, N311);
buf BUF1 (N963, N950);
nor NOR4 (N964, N963, N224, N101, N953);
not NOT1 (N965, N283);
and AND3 (N966, N960, N87, N346);
xor XOR2 (N967, N959, N764);
nand NAND3 (N968, N962, N271, N773);
buf BUF1 (N969, N956);
or OR3 (N970, N964, N731, N812);
nor NOR2 (N971, N961, N133);
xor XOR2 (N972, N970, N674);
or OR3 (N973, N955, N250, N99);
buf BUF1 (N974, N965);
or OR3 (N975, N967, N257, N679);
not NOT1 (N976, N968);
buf BUF1 (N977, N973);
not NOT1 (N978, N969);
buf BUF1 (N979, N974);
and AND4 (N980, N966, N561, N480, N528);
nand NAND4 (N981, N972, N278, N884, N708);
nand NAND3 (N982, N979, N757, N538);
and AND2 (N983, N945, N677);
buf BUF1 (N984, N975);
buf BUF1 (N985, N978);
and AND2 (N986, N976, N750);
nand NAND4 (N987, N933, N146, N80, N560);
not NOT1 (N988, N985);
buf BUF1 (N989, N986);
xor XOR2 (N990, N981, N549);
nand NAND2 (N991, N977, N276);
and AND2 (N992, N991, N877);
or OR3 (N993, N984, N205, N225);
buf BUF1 (N994, N983);
nor NOR4 (N995, N980, N491, N111, N470);
or OR4 (N996, N987, N739, N828, N235);
or OR3 (N997, N995, N29, N405);
nor NOR4 (N998, N982, N813, N688, N253);
and AND3 (N999, N992, N486, N761);
buf BUF1 (N1000, N997);
nor NOR4 (N1001, N996, N750, N438, N590);
xor XOR2 (N1002, N988, N662);
nor NOR4 (N1003, N1000, N585, N248, N456);
and AND2 (N1004, N971, N925);
or OR2 (N1005, N993, N812);
nor NOR3 (N1006, N999, N379, N947);
buf BUF1 (N1007, N1003);
or OR2 (N1008, N990, N670);
not NOT1 (N1009, N998);
nor NOR2 (N1010, N989, N396);
and AND2 (N1011, N1007, N300);
buf BUF1 (N1012, N1002);
buf BUF1 (N1013, N1005);
and AND3 (N1014, N1009, N365, N475);
buf BUF1 (N1015, N1012);
and AND3 (N1016, N1010, N533, N605);
not NOT1 (N1017, N1001);
xor XOR2 (N1018, N1014, N1009);
or OR2 (N1019, N1008, N583);
and AND4 (N1020, N1011, N683, N366, N241);
nor NOR3 (N1021, N994, N578, N937);
nand NAND4 (N1022, N1013, N27, N506, N731);
buf BUF1 (N1023, N1018);
nand NAND3 (N1024, N1016, N756, N39);
or OR3 (N1025, N1024, N242, N344);
xor XOR2 (N1026, N1015, N809);
nor NOR2 (N1027, N1025, N914);
xor XOR2 (N1028, N1019, N48);
and AND2 (N1029, N1004, N843);
xor XOR2 (N1030, N1023, N588);
nand NAND2 (N1031, N1021, N844);
xor XOR2 (N1032, N1029, N606);
buf BUF1 (N1033, N1017);
xor XOR2 (N1034, N1033, N139);
nand NAND3 (N1035, N1027, N85, N309);
or OR2 (N1036, N1031, N571);
not NOT1 (N1037, N1022);
or OR3 (N1038, N1035, N825, N408);
not NOT1 (N1039, N1032);
not NOT1 (N1040, N1020);
or OR4 (N1041, N1036, N79, N548, N329);
and AND4 (N1042, N1034, N217, N839, N875);
not NOT1 (N1043, N1028);
and AND3 (N1044, N1026, N65, N549);
nand NAND4 (N1045, N1039, N131, N857, N499);
xor XOR2 (N1046, N1030, N290);
not NOT1 (N1047, N1043);
and AND2 (N1048, N1041, N1040);
not NOT1 (N1049, N16);
xor XOR2 (N1050, N1042, N463);
buf BUF1 (N1051, N1006);
xor XOR2 (N1052, N1037, N1038);
and AND3 (N1053, N936, N3, N560);
xor XOR2 (N1054, N1052, N327);
and AND3 (N1055, N1046, N393, N99);
or OR3 (N1056, N1044, N1000, N951);
xor XOR2 (N1057, N1054, N221);
nand NAND4 (N1058, N1051, N1009, N1022, N79);
nor NOR3 (N1059, N1048, N237, N511);
xor XOR2 (N1060, N1047, N506);
nand NAND3 (N1061, N1055, N605, N930);
not NOT1 (N1062, N1060);
not NOT1 (N1063, N1053);
xor XOR2 (N1064, N1059, N413);
or OR3 (N1065, N1050, N654, N662);
or OR2 (N1066, N1056, N884);
xor XOR2 (N1067, N1049, N821);
or OR2 (N1068, N1065, N766);
nand NAND2 (N1069, N1061, N1046);
buf BUF1 (N1070, N1064);
nor NOR4 (N1071, N1062, N44, N982, N612);
or OR4 (N1072, N1067, N233, N164, N80);
or OR2 (N1073, N1058, N356);
nor NOR3 (N1074, N1071, N192, N236);
and AND3 (N1075, N1073, N851, N714);
not NOT1 (N1076, N1066);
nand NAND4 (N1077, N1063, N825, N185, N622);
and AND2 (N1078, N1075, N137);
nor NOR4 (N1079, N1070, N252, N912, N750);
buf BUF1 (N1080, N1078);
not NOT1 (N1081, N1069);
or OR3 (N1082, N1079, N774, N416);
or OR2 (N1083, N1068, N643);
nor NOR2 (N1084, N1045, N208);
nor NOR3 (N1085, N1077, N492, N889);
or OR4 (N1086, N1057, N466, N795, N887);
nor NOR2 (N1087, N1080, N648);
or OR4 (N1088, N1082, N224, N605, N815);
not NOT1 (N1089, N1083);
xor XOR2 (N1090, N1087, N765);
buf BUF1 (N1091, N1085);
nand NAND4 (N1092, N1086, N956, N924, N787);
buf BUF1 (N1093, N1081);
xor XOR2 (N1094, N1091, N645);
xor XOR2 (N1095, N1093, N231);
nor NOR2 (N1096, N1076, N243);
buf BUF1 (N1097, N1092);
not NOT1 (N1098, N1096);
nor NOR3 (N1099, N1084, N142, N640);
and AND4 (N1100, N1095, N373, N407, N145);
or OR2 (N1101, N1074, N74);
nor NOR2 (N1102, N1098, N287);
and AND4 (N1103, N1102, N720, N38, N1043);
nor NOR2 (N1104, N1097, N333);
nand NAND4 (N1105, N1090, N692, N171, N952);
or OR3 (N1106, N1100, N196, N95);
not NOT1 (N1107, N1103);
nor NOR3 (N1108, N1104, N754, N521);
xor XOR2 (N1109, N1108, N322);
and AND3 (N1110, N1088, N496, N411);
nand NAND4 (N1111, N1101, N285, N580, N854);
xor XOR2 (N1112, N1111, N321);
and AND2 (N1113, N1107, N1023);
nor NOR2 (N1114, N1072, N476);
and AND3 (N1115, N1105, N1069, N67);
not NOT1 (N1116, N1114);
buf BUF1 (N1117, N1113);
buf BUF1 (N1118, N1109);
nand NAND2 (N1119, N1117, N627);
buf BUF1 (N1120, N1115);
or OR3 (N1121, N1110, N1069, N478);
or OR2 (N1122, N1118, N978);
or OR3 (N1123, N1099, N675, N742);
nand NAND3 (N1124, N1112, N255, N175);
or OR4 (N1125, N1121, N764, N910, N608);
nor NOR4 (N1126, N1094, N142, N36, N589);
nor NOR2 (N1127, N1119, N854);
nor NOR2 (N1128, N1089, N539);
not NOT1 (N1129, N1127);
or OR2 (N1130, N1122, N256);
buf BUF1 (N1131, N1106);
nor NOR3 (N1132, N1129, N250, N771);
not NOT1 (N1133, N1130);
or OR4 (N1134, N1123, N831, N1080, N275);
nand NAND4 (N1135, N1128, N408, N510, N420);
nor NOR2 (N1136, N1124, N771);
nor NOR3 (N1137, N1132, N226, N256);
xor XOR2 (N1138, N1120, N623);
or OR3 (N1139, N1136, N476, N542);
and AND4 (N1140, N1125, N929, N157, N344);
not NOT1 (N1141, N1137);
not NOT1 (N1142, N1135);
buf BUF1 (N1143, N1116);
nor NOR2 (N1144, N1133, N701);
nor NOR4 (N1145, N1138, N155, N503, N591);
and AND4 (N1146, N1144, N742, N493, N1128);
xor XOR2 (N1147, N1126, N247);
xor XOR2 (N1148, N1146, N396);
or OR3 (N1149, N1139, N288, N314);
xor XOR2 (N1150, N1147, N546);
or OR3 (N1151, N1150, N900, N576);
not NOT1 (N1152, N1142);
buf BUF1 (N1153, N1145);
nor NOR4 (N1154, N1151, N201, N373, N442);
nor NOR3 (N1155, N1140, N770, N519);
nand NAND4 (N1156, N1155, N763, N471, N31);
nand NAND2 (N1157, N1148, N284);
xor XOR2 (N1158, N1154, N372);
or OR3 (N1159, N1131, N294, N830);
nand NAND4 (N1160, N1159, N966, N798, N1060);
nand NAND4 (N1161, N1149, N626, N156, N247);
or OR2 (N1162, N1141, N36);
not NOT1 (N1163, N1160);
buf BUF1 (N1164, N1157);
and AND4 (N1165, N1152, N406, N507, N823);
buf BUF1 (N1166, N1158);
buf BUF1 (N1167, N1163);
nor NOR3 (N1168, N1153, N751, N106);
not NOT1 (N1169, N1161);
or OR2 (N1170, N1143, N311);
and AND2 (N1171, N1167, N160);
nand NAND2 (N1172, N1168, N617);
nand NAND3 (N1173, N1172, N706, N153);
and AND4 (N1174, N1173, N2, N967, N698);
nor NOR4 (N1175, N1170, N739, N75, N307);
nor NOR2 (N1176, N1175, N469);
or OR3 (N1177, N1169, N949, N955);
or OR2 (N1178, N1162, N877);
nand NAND4 (N1179, N1178, N726, N362, N411);
buf BUF1 (N1180, N1165);
or OR2 (N1181, N1164, N689);
and AND2 (N1182, N1181, N987);
buf BUF1 (N1183, N1134);
and AND3 (N1184, N1171, N7, N688);
buf BUF1 (N1185, N1156);
nand NAND3 (N1186, N1179, N1126, N769);
and AND2 (N1187, N1185, N295);
nand NAND3 (N1188, N1176, N729, N1080);
not NOT1 (N1189, N1177);
and AND4 (N1190, N1180, N420, N801, N445);
buf BUF1 (N1191, N1189);
xor XOR2 (N1192, N1183, N1082);
or OR3 (N1193, N1182, N17, N983);
not NOT1 (N1194, N1188);
nor NOR4 (N1195, N1186, N934, N1091, N699);
nor NOR4 (N1196, N1187, N360, N247, N265);
not NOT1 (N1197, N1184);
nor NOR2 (N1198, N1192, N562);
and AND4 (N1199, N1190, N1195, N721, N466);
xor XOR2 (N1200, N259, N889);
and AND3 (N1201, N1194, N78, N1194);
nor NOR4 (N1202, N1199, N4, N1116, N350);
buf BUF1 (N1203, N1193);
xor XOR2 (N1204, N1191, N84);
not NOT1 (N1205, N1197);
or OR4 (N1206, N1198, N73, N971, N404);
not NOT1 (N1207, N1205);
nand NAND2 (N1208, N1196, N176);
not NOT1 (N1209, N1174);
and AND4 (N1210, N1204, N330, N673, N708);
nand NAND3 (N1211, N1208, N151, N251);
buf BUF1 (N1212, N1209);
or OR3 (N1213, N1211, N662, N701);
and AND4 (N1214, N1210, N473, N68, N628);
nand NAND4 (N1215, N1214, N363, N128, N1117);
buf BUF1 (N1216, N1212);
nor NOR2 (N1217, N1203, N128);
nand NAND2 (N1218, N1215, N756);
and AND2 (N1219, N1206, N963);
not NOT1 (N1220, N1219);
nand NAND2 (N1221, N1216, N601);
and AND4 (N1222, N1202, N78, N282, N629);
or OR2 (N1223, N1200, N675);
and AND4 (N1224, N1217, N1136, N711, N27);
xor XOR2 (N1225, N1224, N1029);
and AND2 (N1226, N1222, N333);
and AND2 (N1227, N1166, N677);
buf BUF1 (N1228, N1225);
not NOT1 (N1229, N1220);
nand NAND4 (N1230, N1221, N513, N1137, N697);
or OR2 (N1231, N1230, N461);
xor XOR2 (N1232, N1213, N326);
buf BUF1 (N1233, N1228);
and AND3 (N1234, N1201, N1107, N1195);
not NOT1 (N1235, N1227);
and AND4 (N1236, N1226, N1230, N214, N42);
xor XOR2 (N1237, N1235, N71);
not NOT1 (N1238, N1229);
buf BUF1 (N1239, N1218);
nor NOR4 (N1240, N1236, N123, N434, N652);
not NOT1 (N1241, N1223);
and AND2 (N1242, N1241, N288);
or OR2 (N1243, N1231, N1124);
not NOT1 (N1244, N1242);
buf BUF1 (N1245, N1238);
or OR4 (N1246, N1234, N467, N865, N1104);
nor NOR3 (N1247, N1243, N1057, N1027);
buf BUF1 (N1248, N1247);
buf BUF1 (N1249, N1237);
nand NAND3 (N1250, N1249, N1083, N27);
nor NOR4 (N1251, N1248, N104, N875, N1148);
and AND4 (N1252, N1251, N949, N342, N1135);
and AND2 (N1253, N1240, N68);
nor NOR3 (N1254, N1232, N1154, N795);
or OR4 (N1255, N1246, N603, N781, N110);
nor NOR4 (N1256, N1255, N1062, N48, N475);
or OR2 (N1257, N1250, N618);
and AND3 (N1258, N1244, N150, N461);
xor XOR2 (N1259, N1254, N449);
xor XOR2 (N1260, N1239, N82);
nor NOR4 (N1261, N1259, N11, N1227, N113);
and AND2 (N1262, N1252, N384);
not NOT1 (N1263, N1261);
nand NAND2 (N1264, N1262, N719);
buf BUF1 (N1265, N1263);
not NOT1 (N1266, N1256);
and AND4 (N1267, N1264, N1186, N814, N731);
nor NOR4 (N1268, N1245, N1219, N688, N253);
nand NAND4 (N1269, N1233, N212, N309, N97);
and AND3 (N1270, N1260, N946, N129);
xor XOR2 (N1271, N1257, N22);
or OR2 (N1272, N1269, N163);
or OR3 (N1273, N1265, N338, N15);
and AND3 (N1274, N1267, N606, N1018);
and AND2 (N1275, N1258, N102);
nand NAND3 (N1276, N1207, N186, N542);
and AND2 (N1277, N1275, N239);
not NOT1 (N1278, N1253);
and AND4 (N1279, N1270, N362, N427, N590);
buf BUF1 (N1280, N1277);
xor XOR2 (N1281, N1268, N567);
xor XOR2 (N1282, N1272, N308);
or OR4 (N1283, N1281, N79, N1215, N571);
nor NOR2 (N1284, N1276, N876);
and AND3 (N1285, N1273, N312, N335);
not NOT1 (N1286, N1279);
not NOT1 (N1287, N1286);
nand NAND2 (N1288, N1287, N561);
buf BUF1 (N1289, N1285);
buf BUF1 (N1290, N1274);
and AND2 (N1291, N1266, N167);
buf BUF1 (N1292, N1284);
xor XOR2 (N1293, N1290, N1113);
nor NOR4 (N1294, N1292, N462, N504, N223);
and AND4 (N1295, N1288, N533, N26, N437);
not NOT1 (N1296, N1291);
or OR2 (N1297, N1296, N1136);
xor XOR2 (N1298, N1297, N260);
and AND4 (N1299, N1295, N571, N1044, N215);
not NOT1 (N1300, N1293);
nand NAND3 (N1301, N1294, N321, N592);
nand NAND4 (N1302, N1299, N1167, N634, N1137);
or OR2 (N1303, N1300, N32);
and AND2 (N1304, N1278, N1048);
buf BUF1 (N1305, N1298);
or OR2 (N1306, N1271, N320);
and AND2 (N1307, N1306, N930);
and AND2 (N1308, N1301, N1167);
or OR2 (N1309, N1282, N60);
nor NOR4 (N1310, N1289, N1264, N52, N930);
and AND4 (N1311, N1305, N380, N497, N1009);
and AND2 (N1312, N1311, N1077);
buf BUF1 (N1313, N1304);
nor NOR3 (N1314, N1303, N274, N1078);
xor XOR2 (N1315, N1307, N482);
not NOT1 (N1316, N1309);
and AND4 (N1317, N1313, N234, N147, N1159);
xor XOR2 (N1318, N1312, N1178);
or OR4 (N1319, N1302, N1184, N529, N207);
xor XOR2 (N1320, N1318, N554);
or OR3 (N1321, N1283, N168, N603);
or OR3 (N1322, N1310, N367, N425);
nor NOR3 (N1323, N1280, N169, N669);
or OR3 (N1324, N1320, N1158, N260);
xor XOR2 (N1325, N1319, N773);
buf BUF1 (N1326, N1317);
nor NOR2 (N1327, N1324, N894);
buf BUF1 (N1328, N1323);
xor XOR2 (N1329, N1325, N602);
nand NAND3 (N1330, N1322, N511, N173);
xor XOR2 (N1331, N1321, N127);
or OR2 (N1332, N1316, N749);
and AND4 (N1333, N1329, N1094, N120, N322);
nand NAND2 (N1334, N1314, N976);
or OR4 (N1335, N1334, N191, N647, N1063);
not NOT1 (N1336, N1331);
nor NOR4 (N1337, N1315, N346, N1332, N18);
buf BUF1 (N1338, N293);
and AND4 (N1339, N1335, N153, N240, N673);
nand NAND4 (N1340, N1337, N609, N810, N976);
and AND3 (N1341, N1336, N234, N145);
not NOT1 (N1342, N1308);
or OR3 (N1343, N1326, N501, N12);
nor NOR4 (N1344, N1342, N463, N355, N204);
and AND2 (N1345, N1341, N393);
xor XOR2 (N1346, N1343, N1150);
nand NAND2 (N1347, N1340, N1189);
and AND4 (N1348, N1344, N440, N1169, N1148);
nor NOR3 (N1349, N1345, N1217, N926);
buf BUF1 (N1350, N1347);
buf BUF1 (N1351, N1349);
not NOT1 (N1352, N1339);
or OR2 (N1353, N1328, N25);
nor NOR2 (N1354, N1350, N775);
or OR3 (N1355, N1351, N946, N1083);
and AND4 (N1356, N1327, N97, N1125, N1252);
nand NAND4 (N1357, N1346, N1103, N921, N750);
nand NAND4 (N1358, N1353, N1099, N1138, N197);
not NOT1 (N1359, N1330);
nand NAND4 (N1360, N1359, N283, N623, N352);
xor XOR2 (N1361, N1352, N672);
and AND4 (N1362, N1357, N975, N763, N758);
not NOT1 (N1363, N1358);
not NOT1 (N1364, N1356);
xor XOR2 (N1365, N1354, N75);
nor NOR3 (N1366, N1363, N838, N558);
nand NAND2 (N1367, N1361, N1146);
nor NOR4 (N1368, N1333, N311, N1196, N998);
or OR4 (N1369, N1355, N1338, N911, N697);
nand NAND3 (N1370, N144, N272, N211);
nor NOR4 (N1371, N1369, N347, N76, N488);
buf BUF1 (N1372, N1360);
xor XOR2 (N1373, N1348, N1251);
not NOT1 (N1374, N1371);
or OR3 (N1375, N1366, N488, N415);
nand NAND3 (N1376, N1375, N1088, N464);
not NOT1 (N1377, N1367);
nand NAND4 (N1378, N1362, N117, N216, N1087);
nand NAND2 (N1379, N1365, N1063);
not NOT1 (N1380, N1376);
nor NOR4 (N1381, N1370, N32, N881, N930);
xor XOR2 (N1382, N1378, N636);
nor NOR2 (N1383, N1372, N1330);
not NOT1 (N1384, N1373);
buf BUF1 (N1385, N1364);
xor XOR2 (N1386, N1379, N274);
nand NAND3 (N1387, N1383, N575, N528);
buf BUF1 (N1388, N1374);
not NOT1 (N1389, N1385);
nor NOR3 (N1390, N1389, N868, N457);
and AND3 (N1391, N1380, N72, N91);
and AND4 (N1392, N1387, N86, N154, N997);
nand NAND3 (N1393, N1386, N1158, N1149);
and AND2 (N1394, N1368, N826);
and AND2 (N1395, N1392, N577);
nor NOR2 (N1396, N1377, N810);
not NOT1 (N1397, N1393);
nand NAND2 (N1398, N1395, N1209);
or OR2 (N1399, N1396, N716);
nand NAND2 (N1400, N1398, N108);
xor XOR2 (N1401, N1400, N474);
or OR4 (N1402, N1388, N960, N1195, N1307);
buf BUF1 (N1403, N1382);
nand NAND4 (N1404, N1403, N671, N857, N207);
buf BUF1 (N1405, N1390);
nor NOR3 (N1406, N1397, N146, N867);
and AND4 (N1407, N1381, N770, N1029, N207);
and AND3 (N1408, N1407, N401, N52);
and AND4 (N1409, N1401, N754, N188, N327);
xor XOR2 (N1410, N1408, N842);
or OR2 (N1411, N1404, N789);
nor NOR3 (N1412, N1402, N735, N84);
and AND2 (N1413, N1391, N1361);
nor NOR2 (N1414, N1405, N913);
nor NOR3 (N1415, N1412, N918, N1224);
buf BUF1 (N1416, N1415);
not NOT1 (N1417, N1416);
buf BUF1 (N1418, N1414);
buf BUF1 (N1419, N1417);
not NOT1 (N1420, N1409);
not NOT1 (N1421, N1413);
not NOT1 (N1422, N1410);
and AND3 (N1423, N1421, N36, N137);
nand NAND2 (N1424, N1394, N357);
nor NOR2 (N1425, N1406, N1301);
buf BUF1 (N1426, N1420);
not NOT1 (N1427, N1422);
nand NAND4 (N1428, N1423, N452, N167, N960);
or OR3 (N1429, N1411, N439, N337);
not NOT1 (N1430, N1429);
or OR4 (N1431, N1384, N1144, N272, N201);
not NOT1 (N1432, N1427);
not NOT1 (N1433, N1430);
not NOT1 (N1434, N1424);
not NOT1 (N1435, N1434);
nand NAND2 (N1436, N1435, N280);
buf BUF1 (N1437, N1432);
buf BUF1 (N1438, N1437);
or OR2 (N1439, N1431, N468);
nand NAND2 (N1440, N1436, N779);
nand NAND2 (N1441, N1399, N210);
xor XOR2 (N1442, N1428, N336);
buf BUF1 (N1443, N1433);
not NOT1 (N1444, N1442);
not NOT1 (N1445, N1426);
and AND2 (N1446, N1438, N453);
and AND2 (N1447, N1444, N1159);
xor XOR2 (N1448, N1447, N1032);
or OR2 (N1449, N1446, N424);
not NOT1 (N1450, N1449);
xor XOR2 (N1451, N1450, N298);
or OR2 (N1452, N1451, N383);
xor XOR2 (N1453, N1448, N599);
nor NOR2 (N1454, N1419, N855);
not NOT1 (N1455, N1440);
nand NAND3 (N1456, N1454, N300, N223);
xor XOR2 (N1457, N1441, N810);
nor NOR3 (N1458, N1425, N1132, N966);
nand NAND4 (N1459, N1456, N382, N175, N633);
xor XOR2 (N1460, N1459, N829);
xor XOR2 (N1461, N1418, N565);
or OR2 (N1462, N1453, N1111);
nand NAND4 (N1463, N1445, N925, N959, N721);
and AND4 (N1464, N1455, N153, N1277, N196);
not NOT1 (N1465, N1457);
and AND3 (N1466, N1462, N942, N747);
and AND2 (N1467, N1439, N138);
xor XOR2 (N1468, N1467, N702);
xor XOR2 (N1469, N1464, N242);
nand NAND2 (N1470, N1468, N341);
and AND4 (N1471, N1463, N601, N1290, N223);
xor XOR2 (N1472, N1461, N167);
not NOT1 (N1473, N1470);
or OR4 (N1474, N1465, N750, N369, N1206);
buf BUF1 (N1475, N1471);
buf BUF1 (N1476, N1443);
nand NAND2 (N1477, N1452, N19);
nand NAND4 (N1478, N1473, N1394, N104, N399);
not NOT1 (N1479, N1469);
buf BUF1 (N1480, N1479);
not NOT1 (N1481, N1458);
buf BUF1 (N1482, N1460);
and AND4 (N1483, N1477, N591, N1291, N1120);
or OR3 (N1484, N1481, N1137, N1331);
and AND4 (N1485, N1466, N893, N502, N989);
buf BUF1 (N1486, N1475);
xor XOR2 (N1487, N1478, N88);
nor NOR3 (N1488, N1485, N970, N6);
nand NAND4 (N1489, N1487, N970, N48, N266);
not NOT1 (N1490, N1474);
xor XOR2 (N1491, N1490, N1150);
and AND3 (N1492, N1482, N519, N690);
nor NOR4 (N1493, N1476, N215, N1123, N698);
buf BUF1 (N1494, N1493);
nand NAND4 (N1495, N1494, N289, N105, N187);
nand NAND4 (N1496, N1483, N931, N827, N207);
nand NAND4 (N1497, N1489, N948, N1037, N947);
and AND2 (N1498, N1484, N1402);
nand NAND4 (N1499, N1495, N1069, N713, N145);
nand NAND2 (N1500, N1496, N1117);
and AND3 (N1501, N1486, N907, N766);
nand NAND3 (N1502, N1491, N1151, N1352);
not NOT1 (N1503, N1499);
xor XOR2 (N1504, N1472, N625);
and AND3 (N1505, N1492, N1359, N101);
or OR2 (N1506, N1498, N548);
nor NOR2 (N1507, N1503, N361);
and AND3 (N1508, N1504, N134, N899);
buf BUF1 (N1509, N1508);
xor XOR2 (N1510, N1501, N359);
buf BUF1 (N1511, N1505);
not NOT1 (N1512, N1500);
nor NOR3 (N1513, N1488, N105, N1164);
buf BUF1 (N1514, N1512);
xor XOR2 (N1515, N1480, N696);
not NOT1 (N1516, N1511);
xor XOR2 (N1517, N1514, N605);
not NOT1 (N1518, N1497);
not NOT1 (N1519, N1513);
nor NOR4 (N1520, N1510, N443, N941, N669);
xor XOR2 (N1521, N1520, N176);
nor NOR4 (N1522, N1515, N993, N700, N1246);
and AND3 (N1523, N1506, N158, N1265);
xor XOR2 (N1524, N1522, N991);
not NOT1 (N1525, N1518);
xor XOR2 (N1526, N1524, N795);
or OR4 (N1527, N1523, N1153, N31, N903);
xor XOR2 (N1528, N1516, N119);
xor XOR2 (N1529, N1528, N778);
nor NOR4 (N1530, N1507, N250, N687, N467);
and AND4 (N1531, N1527, N1017, N104, N187);
xor XOR2 (N1532, N1509, N23);
buf BUF1 (N1533, N1519);
nand NAND3 (N1534, N1532, N1304, N1311);
or OR4 (N1535, N1531, N1479, N376, N1089);
buf BUF1 (N1536, N1530);
not NOT1 (N1537, N1521);
not NOT1 (N1538, N1534);
and AND2 (N1539, N1538, N977);
or OR3 (N1540, N1536, N853, N550);
or OR4 (N1541, N1502, N1537, N1277, N80);
buf BUF1 (N1542, N690);
buf BUF1 (N1543, N1525);
or OR4 (N1544, N1529, N457, N207, N1230);
and AND4 (N1545, N1535, N401, N1020, N712);
and AND4 (N1546, N1541, N837, N852, N73);
nor NOR4 (N1547, N1546, N1507, N1447, N1083);
or OR3 (N1548, N1547, N353, N1129);
nor NOR2 (N1549, N1545, N1041);
and AND2 (N1550, N1526, N981);
or OR3 (N1551, N1549, N1336, N1104);
xor XOR2 (N1552, N1539, N1424);
not NOT1 (N1553, N1517);
not NOT1 (N1554, N1551);
and AND4 (N1555, N1548, N1512, N1047, N1490);
nor NOR4 (N1556, N1555, N1110, N1144, N1127);
not NOT1 (N1557, N1540);
nor NOR4 (N1558, N1554, N780, N9, N899);
buf BUF1 (N1559, N1556);
buf BUF1 (N1560, N1558);
nand NAND3 (N1561, N1550, N598, N1420);
buf BUF1 (N1562, N1542);
not NOT1 (N1563, N1552);
xor XOR2 (N1564, N1533, N626);
not NOT1 (N1565, N1564);
xor XOR2 (N1566, N1565, N724);
not NOT1 (N1567, N1561);
buf BUF1 (N1568, N1562);
buf BUF1 (N1569, N1553);
xor XOR2 (N1570, N1557, N144);
xor XOR2 (N1571, N1567, N421);
and AND3 (N1572, N1566, N75, N1245);
and AND4 (N1573, N1544, N19, N135, N618);
and AND4 (N1574, N1568, N217, N1192, N138);
nor NOR4 (N1575, N1573, N1092, N805, N134);
not NOT1 (N1576, N1563);
xor XOR2 (N1577, N1574, N627);
nand NAND2 (N1578, N1572, N19);
nor NOR4 (N1579, N1570, N1352, N747, N38);
xor XOR2 (N1580, N1559, N780);
buf BUF1 (N1581, N1579);
not NOT1 (N1582, N1576);
xor XOR2 (N1583, N1569, N383);
and AND4 (N1584, N1577, N1254, N400, N1351);
buf BUF1 (N1585, N1575);
nor NOR4 (N1586, N1581, N1380, N789, N303);
and AND2 (N1587, N1583, N956);
nand NAND4 (N1588, N1587, N341, N970, N584);
nor NOR3 (N1589, N1543, N1237, N616);
not NOT1 (N1590, N1571);
or OR4 (N1591, N1590, N1429, N1537, N487);
nand NAND3 (N1592, N1580, N34, N56);
or OR4 (N1593, N1588, N1165, N1371, N139);
buf BUF1 (N1594, N1591);
not NOT1 (N1595, N1585);
xor XOR2 (N1596, N1582, N1272);
xor XOR2 (N1597, N1593, N1446);
nand NAND3 (N1598, N1560, N70, N926);
buf BUF1 (N1599, N1596);
or OR4 (N1600, N1595, N1394, N1148, N498);
nor NOR3 (N1601, N1586, N115, N670);
and AND4 (N1602, N1600, N568, N1533, N1155);
not NOT1 (N1603, N1602);
not NOT1 (N1604, N1594);
and AND2 (N1605, N1603, N184);
xor XOR2 (N1606, N1584, N37);
or OR3 (N1607, N1601, N367, N1569);
or OR4 (N1608, N1606, N777, N1602, N1273);
not NOT1 (N1609, N1598);
nand NAND2 (N1610, N1604, N698);
or OR3 (N1611, N1609, N606, N867);
not NOT1 (N1612, N1611);
not NOT1 (N1613, N1607);
buf BUF1 (N1614, N1613);
not NOT1 (N1615, N1578);
nand NAND3 (N1616, N1608, N1587, N1615);
nand NAND4 (N1617, N1348, N163, N4, N397);
nand NAND3 (N1618, N1605, N972, N1138);
or OR4 (N1619, N1618, N624, N963, N1390);
xor XOR2 (N1620, N1597, N1032);
buf BUF1 (N1621, N1614);
nor NOR4 (N1622, N1592, N1206, N811, N1417);
nand NAND2 (N1623, N1616, N1520);
and AND2 (N1624, N1620, N681);
buf BUF1 (N1625, N1617);
buf BUF1 (N1626, N1599);
buf BUF1 (N1627, N1619);
not NOT1 (N1628, N1627);
nor NOR2 (N1629, N1612, N917);
nor NOR3 (N1630, N1626, N581, N528);
nand NAND4 (N1631, N1622, N534, N362, N1083);
not NOT1 (N1632, N1623);
and AND3 (N1633, N1589, N646, N1063);
buf BUF1 (N1634, N1633);
buf BUF1 (N1635, N1628);
not NOT1 (N1636, N1632);
and AND2 (N1637, N1621, N1144);
nor NOR3 (N1638, N1610, N1106, N784);
and AND2 (N1639, N1638, N1049);
not NOT1 (N1640, N1639);
nor NOR4 (N1641, N1629, N863, N1632, N201);
buf BUF1 (N1642, N1630);
not NOT1 (N1643, N1635);
nor NOR3 (N1644, N1643, N745, N760);
not NOT1 (N1645, N1637);
or OR4 (N1646, N1634, N1287, N351, N1228);
nand NAND4 (N1647, N1645, N625, N412, N1398);
or OR4 (N1648, N1631, N508, N1595, N543);
buf BUF1 (N1649, N1647);
not NOT1 (N1650, N1642);
nor NOR3 (N1651, N1649, N1052, N350);
and AND3 (N1652, N1636, N638, N1129);
xor XOR2 (N1653, N1644, N1095);
and AND4 (N1654, N1624, N146, N1621, N1232);
not NOT1 (N1655, N1648);
buf BUF1 (N1656, N1655);
nand NAND4 (N1657, N1652, N1539, N1176, N1086);
not NOT1 (N1658, N1650);
and AND3 (N1659, N1657, N556, N1487);
not NOT1 (N1660, N1640);
nand NAND3 (N1661, N1658, N1577, N307);
and AND4 (N1662, N1661, N210, N1636, N288);
or OR4 (N1663, N1654, N832, N1221, N1247);
and AND4 (N1664, N1663, N1021, N715, N14);
nand NAND3 (N1665, N1660, N716, N1111);
or OR3 (N1666, N1662, N281, N1014);
buf BUF1 (N1667, N1665);
nor NOR4 (N1668, N1666, N1645, N22, N1052);
nand NAND3 (N1669, N1625, N409, N1432);
and AND2 (N1670, N1646, N27);
buf BUF1 (N1671, N1641);
not NOT1 (N1672, N1653);
nand NAND4 (N1673, N1651, N1098, N1049, N998);
and AND4 (N1674, N1664, N976, N1446, N631);
not NOT1 (N1675, N1670);
not NOT1 (N1676, N1668);
nor NOR2 (N1677, N1669, N161);
and AND3 (N1678, N1656, N191, N1158);
or OR4 (N1679, N1677, N1363, N314, N648);
xor XOR2 (N1680, N1679, N765);
xor XOR2 (N1681, N1671, N1138);
nand NAND3 (N1682, N1674, N777, N621);
nor NOR2 (N1683, N1675, N1);
nor NOR4 (N1684, N1673, N1625, N1271, N728);
nand NAND4 (N1685, N1659, N1530, N1436, N502);
or OR2 (N1686, N1678, N1463);
buf BUF1 (N1687, N1685);
nand NAND4 (N1688, N1682, N482, N242, N1554);
or OR4 (N1689, N1667, N761, N509, N480);
xor XOR2 (N1690, N1686, N83);
and AND3 (N1691, N1689, N434, N1553);
xor XOR2 (N1692, N1691, N616);
xor XOR2 (N1693, N1676, N1173);
or OR4 (N1694, N1680, N1315, N762, N1647);
buf BUF1 (N1695, N1694);
nor NOR2 (N1696, N1693, N69);
not NOT1 (N1697, N1681);
buf BUF1 (N1698, N1695);
buf BUF1 (N1699, N1696);
xor XOR2 (N1700, N1699, N380);
not NOT1 (N1701, N1684);
xor XOR2 (N1702, N1687, N49);
nand NAND2 (N1703, N1698, N1255);
not NOT1 (N1704, N1672);
and AND4 (N1705, N1690, N9, N82, N977);
xor XOR2 (N1706, N1688, N1395);
not NOT1 (N1707, N1701);
nand NAND4 (N1708, N1697, N1537, N1366, N805);
and AND4 (N1709, N1706, N50, N1147, N294);
xor XOR2 (N1710, N1707, N510);
buf BUF1 (N1711, N1692);
xor XOR2 (N1712, N1702, N1606);
not NOT1 (N1713, N1709);
or OR3 (N1714, N1683, N16, N574);
nand NAND2 (N1715, N1700, N1227);
not NOT1 (N1716, N1714);
nor NOR2 (N1717, N1715, N980);
xor XOR2 (N1718, N1705, N71);
nand NAND4 (N1719, N1716, N1233, N1202, N527);
buf BUF1 (N1720, N1710);
not NOT1 (N1721, N1704);
buf BUF1 (N1722, N1721);
and AND4 (N1723, N1722, N734, N1371, N289);
not NOT1 (N1724, N1712);
nand NAND3 (N1725, N1713, N727, N757);
xor XOR2 (N1726, N1717, N89);
buf BUF1 (N1727, N1724);
buf BUF1 (N1728, N1726);
nand NAND3 (N1729, N1723, N381, N914);
buf BUF1 (N1730, N1729);
nor NOR3 (N1731, N1728, N983, N334);
buf BUF1 (N1732, N1727);
nand NAND3 (N1733, N1732, N1731, N447);
nor NOR4 (N1734, N1644, N1649, N1019, N1428);
and AND2 (N1735, N1725, N292);
nor NOR3 (N1736, N1730, N623, N1682);
not NOT1 (N1737, N1703);
nand NAND4 (N1738, N1708, N1604, N1171, N647);
nor NOR2 (N1739, N1719, N1531);
xor XOR2 (N1740, N1737, N860);
buf BUF1 (N1741, N1736);
and AND4 (N1742, N1711, N393, N657, N338);
not NOT1 (N1743, N1741);
xor XOR2 (N1744, N1739, N871);
or OR3 (N1745, N1735, N1738, N1004);
or OR4 (N1746, N718, N16, N902, N118);
not NOT1 (N1747, N1733);
xor XOR2 (N1748, N1746, N1089);
nand NAND2 (N1749, N1718, N158);
nor NOR4 (N1750, N1747, N945, N647, N317);
buf BUF1 (N1751, N1744);
nand NAND2 (N1752, N1743, N513);
buf BUF1 (N1753, N1742);
buf BUF1 (N1754, N1749);
nor NOR3 (N1755, N1720, N749, N340);
buf BUF1 (N1756, N1734);
and AND2 (N1757, N1751, N1748);
or OR4 (N1758, N391, N1609, N1561, N493);
not NOT1 (N1759, N1745);
and AND4 (N1760, N1754, N1682, N1406, N274);
nand NAND3 (N1761, N1756, N583, N828);
nor NOR2 (N1762, N1760, N655);
or OR3 (N1763, N1762, N799, N115);
not NOT1 (N1764, N1752);
nor NOR2 (N1765, N1755, N154);
xor XOR2 (N1766, N1750, N279);
and AND4 (N1767, N1761, N512, N1545, N157);
buf BUF1 (N1768, N1753);
buf BUF1 (N1769, N1740);
buf BUF1 (N1770, N1765);
not NOT1 (N1771, N1759);
and AND4 (N1772, N1771, N1397, N68, N289);
buf BUF1 (N1773, N1766);
xor XOR2 (N1774, N1773, N984);
nor NOR4 (N1775, N1763, N490, N819, N1006);
xor XOR2 (N1776, N1770, N1663);
buf BUF1 (N1777, N1764);
or OR2 (N1778, N1772, N718);
or OR3 (N1779, N1778, N762, N1037);
not NOT1 (N1780, N1767);
or OR4 (N1781, N1757, N191, N1510, N1227);
nand NAND2 (N1782, N1768, N1351);
nand NAND4 (N1783, N1780, N1413, N1351, N964);
or OR3 (N1784, N1774, N177, N1570);
or OR3 (N1785, N1775, N1661, N718);
nand NAND4 (N1786, N1781, N75, N970, N110);
nand NAND4 (N1787, N1769, N397, N10, N78);
nor NOR4 (N1788, N1783, N478, N832, N75);
nor NOR4 (N1789, N1777, N66, N479, N674);
or OR2 (N1790, N1787, N1248);
buf BUF1 (N1791, N1779);
nor NOR4 (N1792, N1790, N1475, N31, N1194);
nor NOR2 (N1793, N1792, N28);
or OR4 (N1794, N1793, N1359, N1001, N1030);
or OR4 (N1795, N1788, N1463, N1317, N409);
not NOT1 (N1796, N1785);
nand NAND3 (N1797, N1782, N68, N1173);
nand NAND4 (N1798, N1794, N398, N577, N46);
xor XOR2 (N1799, N1776, N1252);
xor XOR2 (N1800, N1799, N1441);
not NOT1 (N1801, N1758);
nand NAND3 (N1802, N1786, N878, N95);
buf BUF1 (N1803, N1791);
xor XOR2 (N1804, N1797, N1069);
nor NOR3 (N1805, N1804, N1251, N1582);
nor NOR2 (N1806, N1789, N1285);
xor XOR2 (N1807, N1805, N1112);
xor XOR2 (N1808, N1798, N1261);
and AND4 (N1809, N1808, N165, N169, N65);
nand NAND4 (N1810, N1806, N937, N327, N544);
buf BUF1 (N1811, N1784);
nand NAND4 (N1812, N1811, N27, N1276, N666);
and AND2 (N1813, N1801, N154);
and AND2 (N1814, N1807, N226);
not NOT1 (N1815, N1812);
nor NOR3 (N1816, N1815, N1192, N1565);
buf BUF1 (N1817, N1814);
or OR3 (N1818, N1796, N1576, N1533);
nor NOR3 (N1819, N1800, N598, N402);
or OR3 (N1820, N1810, N367, N820);
not NOT1 (N1821, N1813);
not NOT1 (N1822, N1818);
nor NOR3 (N1823, N1795, N333, N1008);
nor NOR2 (N1824, N1802, N1388);
xor XOR2 (N1825, N1819, N178);
buf BUF1 (N1826, N1821);
and AND4 (N1827, N1820, N386, N132, N378);
not NOT1 (N1828, N1823);
not NOT1 (N1829, N1826);
or OR2 (N1830, N1809, N1507);
or OR4 (N1831, N1829, N1759, N585, N887);
not NOT1 (N1832, N1822);
not NOT1 (N1833, N1816);
not NOT1 (N1834, N1817);
nor NOR3 (N1835, N1833, N431, N1028);
nand NAND4 (N1836, N1824, N816, N1253, N1006);
or OR2 (N1837, N1828, N539);
xor XOR2 (N1838, N1803, N132);
and AND3 (N1839, N1835, N1273, N618);
and AND3 (N1840, N1838, N1162, N267);
buf BUF1 (N1841, N1832);
xor XOR2 (N1842, N1841, N94);
xor XOR2 (N1843, N1830, N134);
xor XOR2 (N1844, N1831, N1362);
and AND4 (N1845, N1840, N1193, N1204, N652);
nor NOR2 (N1846, N1834, N130);
not NOT1 (N1847, N1846);
nor NOR2 (N1848, N1836, N1079);
and AND2 (N1849, N1843, N257);
nand NAND3 (N1850, N1845, N1587, N1004);
xor XOR2 (N1851, N1844, N745);
nand NAND3 (N1852, N1851, N282, N279);
or OR2 (N1853, N1842, N561);
buf BUF1 (N1854, N1837);
nand NAND2 (N1855, N1850, N1804);
or OR3 (N1856, N1853, N1637, N1497);
buf BUF1 (N1857, N1854);
buf BUF1 (N1858, N1857);
not NOT1 (N1859, N1839);
buf BUF1 (N1860, N1855);
xor XOR2 (N1861, N1858, N570);
not NOT1 (N1862, N1861);
nand NAND3 (N1863, N1859, N1732, N20);
nand NAND3 (N1864, N1848, N600, N1810);
or OR3 (N1865, N1856, N1233, N280);
or OR4 (N1866, N1852, N1248, N689, N217);
or OR3 (N1867, N1862, N592, N408);
nor NOR4 (N1868, N1864, N629, N1643, N1264);
nand NAND3 (N1869, N1867, N377, N161);
nor NOR4 (N1870, N1863, N790, N1478, N1712);
or OR4 (N1871, N1866, N1172, N847, N816);
xor XOR2 (N1872, N1849, N927);
not NOT1 (N1873, N1847);
and AND3 (N1874, N1825, N644, N1733);
xor XOR2 (N1875, N1865, N1690);
nand NAND2 (N1876, N1875, N1873);
nor NOR2 (N1877, N65, N394);
and AND3 (N1878, N1874, N1745, N707);
or OR3 (N1879, N1870, N1553, N706);
buf BUF1 (N1880, N1860);
not NOT1 (N1881, N1877);
and AND4 (N1882, N1869, N1384, N136, N674);
not NOT1 (N1883, N1868);
buf BUF1 (N1884, N1879);
and AND3 (N1885, N1883, N304, N236);
and AND3 (N1886, N1871, N673, N945);
or OR3 (N1887, N1876, N448, N90);
and AND4 (N1888, N1887, N395, N1441, N143);
xor XOR2 (N1889, N1886, N836);
and AND2 (N1890, N1885, N145);
buf BUF1 (N1891, N1872);
not NOT1 (N1892, N1880);
and AND4 (N1893, N1884, N853, N1875, N491);
xor XOR2 (N1894, N1893, N490);
and AND3 (N1895, N1888, N821, N1768);
xor XOR2 (N1896, N1890, N1554);
or OR3 (N1897, N1891, N1679, N499);
buf BUF1 (N1898, N1878);
buf BUF1 (N1899, N1895);
or OR3 (N1900, N1889, N1049, N396);
xor XOR2 (N1901, N1892, N1540);
or OR3 (N1902, N1827, N1537, N1066);
not NOT1 (N1903, N1897);
buf BUF1 (N1904, N1900);
buf BUF1 (N1905, N1899);
not NOT1 (N1906, N1882);
not NOT1 (N1907, N1906);
buf BUF1 (N1908, N1898);
not NOT1 (N1909, N1904);
buf BUF1 (N1910, N1901);
nand NAND4 (N1911, N1907, N798, N879, N1268);
buf BUF1 (N1912, N1902);
nor NOR3 (N1913, N1910, N1200, N1767);
not NOT1 (N1914, N1912);
xor XOR2 (N1915, N1914, N1511);
and AND4 (N1916, N1915, N1711, N1327, N1453);
or OR3 (N1917, N1896, N554, N609);
buf BUF1 (N1918, N1894);
or OR4 (N1919, N1903, N310, N977, N1222);
and AND3 (N1920, N1917, N1780, N10);
xor XOR2 (N1921, N1881, N1612);
and AND2 (N1922, N1916, N1419);
or OR3 (N1923, N1911, N1793, N393);
or OR3 (N1924, N1920, N1393, N620);
nand NAND3 (N1925, N1922, N1143, N1685);
buf BUF1 (N1926, N1905);
buf BUF1 (N1927, N1918);
or OR4 (N1928, N1925, N1057, N1818, N202);
or OR3 (N1929, N1927, N875, N1395);
and AND3 (N1930, N1926, N376, N1414);
nor NOR3 (N1931, N1930, N627, N85);
buf BUF1 (N1932, N1929);
buf BUF1 (N1933, N1909);
nand NAND3 (N1934, N1932, N55, N3);
nand NAND3 (N1935, N1913, N1112, N1798);
nor NOR2 (N1936, N1924, N518);
buf BUF1 (N1937, N1935);
xor XOR2 (N1938, N1908, N1918);
or OR2 (N1939, N1921, N1828);
nor NOR4 (N1940, N1934, N622, N286, N551);
xor XOR2 (N1941, N1931, N478);
xor XOR2 (N1942, N1928, N1392);
buf BUF1 (N1943, N1936);
not NOT1 (N1944, N1923);
nand NAND4 (N1945, N1942, N1928, N863, N365);
not NOT1 (N1946, N1941);
and AND2 (N1947, N1937, N1338);
nand NAND2 (N1948, N1933, N1333);
not NOT1 (N1949, N1945);
xor XOR2 (N1950, N1943, N41);
nand NAND2 (N1951, N1946, N1339);
nor NOR4 (N1952, N1944, N557, N1183, N1540);
nor NOR4 (N1953, N1952, N1381, N37, N1398);
nor NOR3 (N1954, N1940, N870, N1279);
nand NAND3 (N1955, N1953, N1686, N1788);
or OR4 (N1956, N1919, N1906, N412, N1514);
nand NAND3 (N1957, N1956, N785, N334);
and AND3 (N1958, N1939, N781, N1798);
or OR3 (N1959, N1957, N242, N1860);
and AND4 (N1960, N1955, N1062, N464, N1651);
buf BUF1 (N1961, N1954);
not NOT1 (N1962, N1958);
nor NOR3 (N1963, N1959, N1792, N936);
nor NOR4 (N1964, N1963, N525, N1055, N1616);
or OR2 (N1965, N1950, N1309);
nor NOR2 (N1966, N1965, N480);
or OR3 (N1967, N1951, N200, N1170);
nor NOR2 (N1968, N1938, N213);
xor XOR2 (N1969, N1947, N1688);
and AND3 (N1970, N1969, N361, N1967);
xor XOR2 (N1971, N1808, N1104);
buf BUF1 (N1972, N1960);
or OR4 (N1973, N1964, N511, N1898, N1341);
and AND3 (N1974, N1949, N1482, N1347);
not NOT1 (N1975, N1973);
xor XOR2 (N1976, N1971, N1939);
or OR4 (N1977, N1962, N1210, N1126, N652);
not NOT1 (N1978, N1961);
xor XOR2 (N1979, N1976, N223);
not NOT1 (N1980, N1972);
buf BUF1 (N1981, N1948);
buf BUF1 (N1982, N1981);
xor XOR2 (N1983, N1978, N725);
or OR2 (N1984, N1983, N1872);
and AND2 (N1985, N1980, N1656);
not NOT1 (N1986, N1979);
not NOT1 (N1987, N1985);
and AND3 (N1988, N1970, N1231, N995);
and AND2 (N1989, N1966, N322);
nand NAND2 (N1990, N1968, N1535);
nor NOR2 (N1991, N1984, N1448);
or OR3 (N1992, N1977, N643, N1544);
and AND3 (N1993, N1975, N1195, N1916);
nand NAND4 (N1994, N1982, N115, N1681, N933);
buf BUF1 (N1995, N1974);
or OR3 (N1996, N1991, N682, N811);
buf BUF1 (N1997, N1987);
xor XOR2 (N1998, N1992, N1003);
nor NOR2 (N1999, N1994, N1520);
not NOT1 (N2000, N1998);
not NOT1 (N2001, N1986);
xor XOR2 (N2002, N1995, N1276);
or OR3 (N2003, N1999, N1618, N41);
nor NOR2 (N2004, N1988, N1320);
buf BUF1 (N2005, N1996);
and AND2 (N2006, N2002, N1828);
buf BUF1 (N2007, N1993);
not NOT1 (N2008, N2000);
and AND4 (N2009, N2003, N802, N446, N1629);
xor XOR2 (N2010, N1989, N338);
nand NAND4 (N2011, N2001, N896, N954, N739);
and AND2 (N2012, N2007, N1505);
xor XOR2 (N2013, N2008, N1343);
nand NAND4 (N2014, N2004, N1156, N1448, N1164);
nand NAND2 (N2015, N2006, N1982);
nand NAND4 (N2016, N2005, N1733, N389, N901);
not NOT1 (N2017, N2013);
xor XOR2 (N2018, N2012, N1379);
and AND4 (N2019, N2016, N262, N982, N7);
buf BUF1 (N2020, N2015);
nand NAND3 (N2021, N2019, N1873, N1189);
buf BUF1 (N2022, N2014);
nor NOR2 (N2023, N1997, N1884);
buf BUF1 (N2024, N1990);
xor XOR2 (N2025, N2020, N29);
nor NOR4 (N2026, N2023, N21, N614, N700);
and AND4 (N2027, N2021, N395, N1858, N1222);
and AND2 (N2028, N2018, N1972);
xor XOR2 (N2029, N2011, N1364);
and AND3 (N2030, N2025, N452, N491);
not NOT1 (N2031, N2010);
and AND2 (N2032, N2029, N271);
nand NAND3 (N2033, N2026, N701, N1975);
nor NOR2 (N2034, N2030, N391);
nor NOR4 (N2035, N2028, N2034, N233, N351);
xor XOR2 (N2036, N1927, N1541);
nor NOR2 (N2037, N2036, N1367);
or OR2 (N2038, N2031, N1659);
buf BUF1 (N2039, N2022);
and AND4 (N2040, N2017, N1769, N573, N1219);
nor NOR3 (N2041, N2035, N380, N320);
xor XOR2 (N2042, N2032, N252);
or OR3 (N2043, N2024, N1904, N511);
xor XOR2 (N2044, N2037, N1503);
xor XOR2 (N2045, N2044, N1243);
not NOT1 (N2046, N2033);
buf BUF1 (N2047, N2040);
not NOT1 (N2048, N2041);
nand NAND4 (N2049, N2009, N181, N71, N635);
or OR4 (N2050, N2049, N1815, N1512, N946);
or OR2 (N2051, N2043, N427);
buf BUF1 (N2052, N2050);
nand NAND4 (N2053, N2046, N1085, N736, N1162);
xor XOR2 (N2054, N2047, N393);
buf BUF1 (N2055, N2052);
or OR3 (N2056, N2042, N196, N408);
nor NOR2 (N2057, N2038, N1212);
buf BUF1 (N2058, N2027);
and AND2 (N2059, N2048, N1531);
or OR3 (N2060, N2053, N396, N1172);
buf BUF1 (N2061, N2060);
and AND3 (N2062, N2061, N639, N211);
xor XOR2 (N2063, N2039, N1216);
buf BUF1 (N2064, N2056);
xor XOR2 (N2065, N2058, N260);
not NOT1 (N2066, N2065);
nor NOR2 (N2067, N2057, N1543);
nor NOR2 (N2068, N2059, N1561);
or OR2 (N2069, N2063, N958);
buf BUF1 (N2070, N2068);
not NOT1 (N2071, N2067);
not NOT1 (N2072, N2066);
buf BUF1 (N2073, N2055);
not NOT1 (N2074, N2051);
nor NOR2 (N2075, N2062, N1942);
nand NAND3 (N2076, N2064, N390, N1645);
xor XOR2 (N2077, N2045, N334);
nor NOR4 (N2078, N2076, N445, N2000, N508);
and AND4 (N2079, N2078, N1966, N488, N1689);
not NOT1 (N2080, N2077);
xor XOR2 (N2081, N2070, N44);
not NOT1 (N2082, N2075);
nor NOR4 (N2083, N2082, N1656, N16, N544);
not NOT1 (N2084, N2079);
nor NOR4 (N2085, N2054, N870, N241, N789);
and AND2 (N2086, N2080, N289);
not NOT1 (N2087, N2069);
not NOT1 (N2088, N2081);
not NOT1 (N2089, N2072);
xor XOR2 (N2090, N2085, N1530);
xor XOR2 (N2091, N2071, N845);
buf BUF1 (N2092, N2087);
nand NAND4 (N2093, N2092, N457, N618, N1000);
nor NOR2 (N2094, N2083, N138);
or OR4 (N2095, N2088, N764, N759, N2080);
and AND3 (N2096, N2091, N844, N1605);
nor NOR2 (N2097, N2084, N1129);
xor XOR2 (N2098, N2094, N1481);
nand NAND4 (N2099, N2096, N1805, N1235, N928);
or OR3 (N2100, N2099, N550, N1078);
buf BUF1 (N2101, N2086);
not NOT1 (N2102, N2093);
not NOT1 (N2103, N2073);
not NOT1 (N2104, N2074);
or OR2 (N2105, N2101, N382);
not NOT1 (N2106, N2098);
xor XOR2 (N2107, N2103, N1439);
and AND4 (N2108, N2090, N1449, N571, N1052);
nor NOR4 (N2109, N2107, N43, N1152, N2064);
nor NOR4 (N2110, N2089, N31, N264, N1955);
nor NOR4 (N2111, N2108, N1440, N1018, N1772);
nor NOR4 (N2112, N2109, N229, N1007, N176);
buf BUF1 (N2113, N2102);
nand NAND4 (N2114, N2113, N1162, N52, N358);
not NOT1 (N2115, N2104);
buf BUF1 (N2116, N2112);
nand NAND4 (N2117, N2106, N1666, N351, N1356);
and AND2 (N2118, N2097, N988);
nor NOR4 (N2119, N2110, N142, N298, N1671);
or OR2 (N2120, N2116, N1335);
or OR3 (N2121, N2111, N724, N620);
not NOT1 (N2122, N2114);
or OR3 (N2123, N2117, N124, N352);
not NOT1 (N2124, N2095);
buf BUF1 (N2125, N2122);
not NOT1 (N2126, N2119);
xor XOR2 (N2127, N2118, N87);
and AND3 (N2128, N2127, N1277, N1532);
nor NOR2 (N2129, N2115, N275);
nor NOR3 (N2130, N2121, N1427, N1004);
not NOT1 (N2131, N2100);
nand NAND4 (N2132, N2130, N1418, N996, N74);
or OR3 (N2133, N2128, N860, N2073);
buf BUF1 (N2134, N2133);
buf BUF1 (N2135, N2132);
nand NAND2 (N2136, N2126, N1119);
not NOT1 (N2137, N2125);
buf BUF1 (N2138, N2123);
nand NAND4 (N2139, N2134, N20, N1659, N1920);
nand NAND3 (N2140, N2124, N1078, N1218);
and AND3 (N2141, N2140, N891, N239);
nor NOR3 (N2142, N2139, N1764, N1456);
xor XOR2 (N2143, N2129, N1363);
nor NOR3 (N2144, N2120, N693, N928);
or OR2 (N2145, N2143, N825);
not NOT1 (N2146, N2142);
xor XOR2 (N2147, N2144, N233);
xor XOR2 (N2148, N2146, N114);
and AND4 (N2149, N2148, N805, N619, N1548);
xor XOR2 (N2150, N2137, N507);
not NOT1 (N2151, N2150);
not NOT1 (N2152, N2141);
not NOT1 (N2153, N2152);
and AND4 (N2154, N2131, N1471, N1076, N130);
xor XOR2 (N2155, N2154, N264);
buf BUF1 (N2156, N2147);
or OR2 (N2157, N2105, N869);
buf BUF1 (N2158, N2151);
and AND4 (N2159, N2153, N1054, N679, N1838);
and AND4 (N2160, N2136, N1108, N1001, N1254);
nor NOR3 (N2161, N2135, N151, N1792);
buf BUF1 (N2162, N2138);
nand NAND2 (N2163, N2160, N878);
not NOT1 (N2164, N2157);
and AND3 (N2165, N2162, N1800, N1410);
xor XOR2 (N2166, N2163, N2071);
nand NAND2 (N2167, N2159, N849);
xor XOR2 (N2168, N2145, N2041);
not NOT1 (N2169, N2164);
buf BUF1 (N2170, N2168);
and AND4 (N2171, N2165, N1931, N1627, N1702);
and AND2 (N2172, N2149, N2081);
nand NAND2 (N2173, N2158, N2117);
not NOT1 (N2174, N2161);
nand NAND3 (N2175, N2169, N125, N294);
nand NAND3 (N2176, N2166, N1680, N594);
buf BUF1 (N2177, N2156);
or OR2 (N2178, N2172, N2128);
xor XOR2 (N2179, N2170, N2099);
xor XOR2 (N2180, N2155, N657);
or OR3 (N2181, N2179, N521, N1576);
not NOT1 (N2182, N2174);
xor XOR2 (N2183, N2171, N1955);
nand NAND4 (N2184, N2173, N1601, N91, N1671);
or OR4 (N2185, N2182, N243, N812, N223);
xor XOR2 (N2186, N2177, N62);
xor XOR2 (N2187, N2178, N1185);
and AND3 (N2188, N2181, N147, N1974);
nand NAND2 (N2189, N2175, N993);
nor NOR4 (N2190, N2187, N698, N1428, N467);
buf BUF1 (N2191, N2167);
nor NOR2 (N2192, N2186, N1185);
and AND3 (N2193, N2180, N1615, N1970);
nand NAND2 (N2194, N2192, N2161);
or OR2 (N2195, N2194, N1437);
not NOT1 (N2196, N2185);
or OR4 (N2197, N2189, N1564, N2193, N16);
not NOT1 (N2198, N1149);
not NOT1 (N2199, N2190);
buf BUF1 (N2200, N2176);
xor XOR2 (N2201, N2196, N160);
or OR4 (N2202, N2188, N222, N1308, N1316);
or OR3 (N2203, N2184, N1276, N263);
nand NAND2 (N2204, N2200, N200);
not NOT1 (N2205, N2197);
nand NAND4 (N2206, N2203, N274, N1124, N1728);
nand NAND3 (N2207, N2204, N1048, N1227);
and AND2 (N2208, N2195, N1451);
or OR4 (N2209, N2205, N1607, N98, N124);
nand NAND4 (N2210, N2209, N120, N88, N717);
xor XOR2 (N2211, N2206, N796);
buf BUF1 (N2212, N2208);
and AND4 (N2213, N2191, N1784, N2151, N97);
and AND4 (N2214, N2198, N500, N1043, N1802);
or OR2 (N2215, N2201, N927);
and AND3 (N2216, N2213, N1891, N1805);
nor NOR2 (N2217, N2210, N271);
nor NOR4 (N2218, N2217, N1790, N276, N2076);
not NOT1 (N2219, N2183);
buf BUF1 (N2220, N2214);
not NOT1 (N2221, N2199);
not NOT1 (N2222, N2219);
nor NOR3 (N2223, N2212, N1079, N1515);
nor NOR3 (N2224, N2222, N1565, N474);
buf BUF1 (N2225, N2202);
or OR3 (N2226, N2216, N1482, N2145);
or OR4 (N2227, N2215, N800, N824, N537);
buf BUF1 (N2228, N2221);
nor NOR3 (N2229, N2207, N1585, N722);
not NOT1 (N2230, N2211);
nor NOR2 (N2231, N2230, N916);
or OR4 (N2232, N2218, N1782, N927, N1382);
nand NAND3 (N2233, N2220, N478, N156);
xor XOR2 (N2234, N2229, N438);
and AND4 (N2235, N2228, N4, N2138, N1872);
buf BUF1 (N2236, N2225);
not NOT1 (N2237, N2223);
not NOT1 (N2238, N2237);
buf BUF1 (N2239, N2236);
or OR4 (N2240, N2232, N1070, N1955, N897);
nand NAND3 (N2241, N2238, N1036, N83);
and AND2 (N2242, N2241, N1100);
nor NOR2 (N2243, N2233, N936);
or OR3 (N2244, N2231, N1451, N1017);
xor XOR2 (N2245, N2244, N1736);
buf BUF1 (N2246, N2234);
or OR3 (N2247, N2243, N426, N265);
and AND2 (N2248, N2239, N409);
nand NAND3 (N2249, N2240, N132, N1334);
buf BUF1 (N2250, N2242);
xor XOR2 (N2251, N2247, N541);
or OR3 (N2252, N2224, N844, N2218);
nand NAND2 (N2253, N2251, N171);
xor XOR2 (N2254, N2227, N1212);
nand NAND4 (N2255, N2248, N934, N174, N1353);
nand NAND4 (N2256, N2235, N1664, N547, N793);
and AND2 (N2257, N2249, N1038);
nor NOR4 (N2258, N2246, N897, N1866, N2179);
and AND3 (N2259, N2256, N424, N648);
xor XOR2 (N2260, N2245, N1376);
not NOT1 (N2261, N2258);
or OR3 (N2262, N2252, N777, N1652);
buf BUF1 (N2263, N2261);
not NOT1 (N2264, N2262);
nor NOR4 (N2265, N2226, N1332, N1844, N1601);
and AND2 (N2266, N2257, N1207);
xor XOR2 (N2267, N2265, N1579);
buf BUF1 (N2268, N2267);
and AND2 (N2269, N2266, N102);
and AND3 (N2270, N2263, N851, N1830);
buf BUF1 (N2271, N2269);
or OR4 (N2272, N2264, N1697, N1068, N597);
xor XOR2 (N2273, N2271, N1180);
not NOT1 (N2274, N2272);
or OR4 (N2275, N2273, N1302, N760, N1150);
buf BUF1 (N2276, N2270);
or OR3 (N2277, N2276, N362, N2244);
nor NOR2 (N2278, N2250, N687);
and AND3 (N2279, N2255, N1772, N600);
buf BUF1 (N2280, N2277);
and AND2 (N2281, N2279, N1150);
and AND3 (N2282, N2260, N129, N1380);
not NOT1 (N2283, N2254);
not NOT1 (N2284, N2281);
and AND4 (N2285, N2284, N1358, N1913, N1160);
buf BUF1 (N2286, N2275);
and AND2 (N2287, N2285, N581);
or OR2 (N2288, N2274, N1438);
and AND3 (N2289, N2280, N76, N185);
xor XOR2 (N2290, N2287, N83);
and AND4 (N2291, N2290, N2171, N526, N127);
nand NAND4 (N2292, N2282, N917, N222, N2161);
xor XOR2 (N2293, N2268, N2172);
or OR2 (N2294, N2288, N132);
nor NOR2 (N2295, N2259, N399);
and AND4 (N2296, N2294, N393, N754, N2035);
nand NAND3 (N2297, N2278, N1067, N1929);
nor NOR2 (N2298, N2286, N1575);
nor NOR3 (N2299, N2298, N1793, N984);
buf BUF1 (N2300, N2253);
xor XOR2 (N2301, N2292, N973);
not NOT1 (N2302, N2283);
nor NOR4 (N2303, N2299, N716, N701, N1544);
nor NOR2 (N2304, N2297, N440);
nor NOR3 (N2305, N2300, N1174, N928);
nand NAND3 (N2306, N2302, N432, N2261);
buf BUF1 (N2307, N2304);
nor NOR3 (N2308, N2291, N414, N210);
not NOT1 (N2309, N2303);
nor NOR2 (N2310, N2295, N1176);
nor NOR2 (N2311, N2289, N999);
not NOT1 (N2312, N2309);
and AND2 (N2313, N2305, N736);
nand NAND2 (N2314, N2312, N1884);
and AND4 (N2315, N2308, N20, N1984, N1230);
buf BUF1 (N2316, N2311);
xor XOR2 (N2317, N2307, N1171);
xor XOR2 (N2318, N2296, N1658);
buf BUF1 (N2319, N2318);
and AND2 (N2320, N2315, N1969);
or OR4 (N2321, N2314, N915, N555, N1153);
not NOT1 (N2322, N2301);
and AND3 (N2323, N2317, N835, N1674);
and AND3 (N2324, N2316, N845, N591);
buf BUF1 (N2325, N2313);
buf BUF1 (N2326, N2310);
or OR2 (N2327, N2323, N624);
and AND3 (N2328, N2327, N2025, N1749);
nor NOR3 (N2329, N2306, N1315, N992);
nand NAND4 (N2330, N2326, N1834, N2097, N1951);
nor NOR3 (N2331, N2328, N525, N308);
nor NOR3 (N2332, N2329, N554, N301);
and AND3 (N2333, N2320, N1092, N782);
buf BUF1 (N2334, N2333);
nor NOR2 (N2335, N2330, N2294);
or OR2 (N2336, N2334, N980);
buf BUF1 (N2337, N2331);
xor XOR2 (N2338, N2324, N1730);
and AND2 (N2339, N2338, N2270);
nand NAND3 (N2340, N2332, N2249, N373);
and AND2 (N2341, N2325, N1440);
or OR2 (N2342, N2319, N1199);
or OR3 (N2343, N2339, N508, N1304);
and AND2 (N2344, N2337, N1992);
xor XOR2 (N2345, N2293, N958);
not NOT1 (N2346, N2340);
and AND2 (N2347, N2346, N173);
xor XOR2 (N2348, N2341, N688);
and AND3 (N2349, N2347, N2185, N1864);
nand NAND4 (N2350, N2343, N1804, N1561, N695);
nor NOR3 (N2351, N2349, N1913, N383);
not NOT1 (N2352, N2345);
and AND2 (N2353, N2348, N757);
and AND2 (N2354, N2321, N2192);
nor NOR2 (N2355, N2335, N1615);
and AND3 (N2356, N2342, N998, N2078);
buf BUF1 (N2357, N2355);
or OR4 (N2358, N2356, N1393, N2038, N802);
buf BUF1 (N2359, N2357);
or OR2 (N2360, N2359, N1114);
and AND4 (N2361, N2350, N699, N1215, N721);
nand NAND3 (N2362, N2344, N1679, N1692);
buf BUF1 (N2363, N2362);
not NOT1 (N2364, N2322);
not NOT1 (N2365, N2336);
xor XOR2 (N2366, N2354, N2037);
not NOT1 (N2367, N2363);
and AND3 (N2368, N2361, N276, N1785);
not NOT1 (N2369, N2353);
xor XOR2 (N2370, N2360, N1244);
not NOT1 (N2371, N2351);
or OR4 (N2372, N2366, N933, N1883, N2094);
buf BUF1 (N2373, N2368);
xor XOR2 (N2374, N2373, N2227);
buf BUF1 (N2375, N2371);
nand NAND4 (N2376, N2369, N213, N1130, N2015);
xor XOR2 (N2377, N2375, N2164);
xor XOR2 (N2378, N2352, N2325);
or OR2 (N2379, N2376, N2331);
or OR2 (N2380, N2364, N421);
not NOT1 (N2381, N2372);
nand NAND2 (N2382, N2378, N970);
xor XOR2 (N2383, N2358, N880);
not NOT1 (N2384, N2383);
not NOT1 (N2385, N2384);
nor NOR3 (N2386, N2380, N741, N2182);
not NOT1 (N2387, N2377);
nor NOR2 (N2388, N2379, N546);
buf BUF1 (N2389, N2365);
not NOT1 (N2390, N2386);
or OR4 (N2391, N2367, N614, N77, N1352);
nand NAND3 (N2392, N2382, N557, N350);
buf BUF1 (N2393, N2374);
nand NAND3 (N2394, N2387, N60, N180);
or OR3 (N2395, N2370, N2091, N940);
and AND4 (N2396, N2393, N560, N974, N1998);
and AND2 (N2397, N2385, N172);
or OR3 (N2398, N2390, N1987, N2377);
or OR4 (N2399, N2391, N5, N1112, N1224);
nand NAND3 (N2400, N2392, N1116, N2042);
and AND2 (N2401, N2388, N870);
or OR4 (N2402, N2398, N1021, N40, N578);
or OR4 (N2403, N2400, N1580, N1424, N1529);
or OR2 (N2404, N2401, N987);
or OR3 (N2405, N2397, N1182, N920);
or OR4 (N2406, N2403, N143, N1160, N228);
buf BUF1 (N2407, N2396);
or OR2 (N2408, N2389, N146);
buf BUF1 (N2409, N2407);
not NOT1 (N2410, N2405);
not NOT1 (N2411, N2395);
nor NOR3 (N2412, N2408, N1364, N1479);
and AND4 (N2413, N2399, N610, N1318, N1309);
not NOT1 (N2414, N2406);
xor XOR2 (N2415, N2412, N1944);
nand NAND2 (N2416, N2415, N2272);
buf BUF1 (N2417, N2414);
not NOT1 (N2418, N2409);
and AND3 (N2419, N2402, N807, N1578);
not NOT1 (N2420, N2413);
xor XOR2 (N2421, N2419, N1085);
or OR3 (N2422, N2381, N1546, N1787);
nand NAND2 (N2423, N2394, N1175);
nor NOR4 (N2424, N2421, N1155, N645, N2092);
xor XOR2 (N2425, N2423, N1695);
buf BUF1 (N2426, N2404);
nand NAND2 (N2427, N2411, N1725);
xor XOR2 (N2428, N2424, N250);
buf BUF1 (N2429, N2417);
nor NOR4 (N2430, N2416, N1692, N1210, N1765);
nand NAND2 (N2431, N2429, N2063);
and AND3 (N2432, N2420, N496, N1169);
xor XOR2 (N2433, N2422, N242);
xor XOR2 (N2434, N2426, N775);
and AND4 (N2435, N2432, N1571, N2224, N2221);
not NOT1 (N2436, N2434);
buf BUF1 (N2437, N2425);
nand NAND3 (N2438, N2410, N1125, N312);
nand NAND4 (N2439, N2435, N1011, N883, N1154);
not NOT1 (N2440, N2438);
not NOT1 (N2441, N2430);
buf BUF1 (N2442, N2431);
not NOT1 (N2443, N2441);
buf BUF1 (N2444, N2437);
nand NAND4 (N2445, N2439, N1848, N654, N2285);
and AND2 (N2446, N2427, N2126);
xor XOR2 (N2447, N2442, N214);
buf BUF1 (N2448, N2447);
and AND3 (N2449, N2445, N1632, N768);
nand NAND4 (N2450, N2436, N696, N1201, N1458);
and AND3 (N2451, N2446, N434, N804);
buf BUF1 (N2452, N2428);
not NOT1 (N2453, N2452);
nor NOR4 (N2454, N2444, N2334, N987, N1236);
or OR4 (N2455, N2440, N775, N1499, N763);
not NOT1 (N2456, N2448);
nand NAND2 (N2457, N2453, N1901);
not NOT1 (N2458, N2450);
or OR4 (N2459, N2449, N1744, N118, N1300);
buf BUF1 (N2460, N2455);
buf BUF1 (N2461, N2418);
nand NAND4 (N2462, N2459, N1758, N155, N1075);
xor XOR2 (N2463, N2462, N912);
not NOT1 (N2464, N2463);
xor XOR2 (N2465, N2458, N1780);
or OR4 (N2466, N2457, N738, N2429, N1216);
xor XOR2 (N2467, N2465, N1550);
xor XOR2 (N2468, N2451, N181);
or OR2 (N2469, N2443, N389);
nand NAND4 (N2470, N2464, N298, N274, N2257);
nand NAND2 (N2471, N2433, N1113);
or OR4 (N2472, N2470, N941, N1539, N200);
nand NAND3 (N2473, N2467, N383, N1066);
nor NOR2 (N2474, N2472, N1296);
not NOT1 (N2475, N2471);
nand NAND4 (N2476, N2475, N1968, N1403, N2302);
nor NOR2 (N2477, N2460, N1586);
and AND3 (N2478, N2474, N202, N724);
buf BUF1 (N2479, N2478);
nand NAND2 (N2480, N2479, N2197);
nand NAND2 (N2481, N2480, N1584);
buf BUF1 (N2482, N2456);
and AND4 (N2483, N2468, N17, N564, N603);
and AND3 (N2484, N2469, N1787, N2138);
not NOT1 (N2485, N2477);
nand NAND4 (N2486, N2473, N1259, N520, N1711);
and AND2 (N2487, N2486, N1172);
not NOT1 (N2488, N2485);
buf BUF1 (N2489, N2461);
nor NOR3 (N2490, N2489, N1097, N771);
and AND2 (N2491, N2482, N809);
nor NOR4 (N2492, N2491, N627, N2271, N307);
or OR4 (N2493, N2481, N1470, N1914, N2179);
xor XOR2 (N2494, N2466, N530);
nand NAND4 (N2495, N2493, N297, N145, N983);
nand NAND2 (N2496, N2490, N622);
nand NAND3 (N2497, N2476, N1410, N1381);
or OR2 (N2498, N2487, N1856);
nand NAND4 (N2499, N2492, N1255, N1391, N311);
buf BUF1 (N2500, N2484);
nand NAND3 (N2501, N2454, N891, N40);
not NOT1 (N2502, N2501);
or OR2 (N2503, N2496, N1869);
and AND4 (N2504, N2500, N383, N1344, N915);
nand NAND4 (N2505, N2494, N2286, N791, N325);
or OR3 (N2506, N2505, N1656, N2197);
not NOT1 (N2507, N2488);
buf BUF1 (N2508, N2499);
buf BUF1 (N2509, N2497);
nor NOR3 (N2510, N2503, N271, N858);
not NOT1 (N2511, N2510);
and AND4 (N2512, N2507, N1810, N842, N1654);
xor XOR2 (N2513, N2511, N1629);
and AND2 (N2514, N2495, N2369);
nand NAND2 (N2515, N2513, N222);
or OR3 (N2516, N2512, N313, N111);
nand NAND3 (N2517, N2515, N1105, N228);
and AND4 (N2518, N2502, N1188, N1476, N2484);
and AND3 (N2519, N2514, N619, N55);
buf BUF1 (N2520, N2504);
not NOT1 (N2521, N2506);
buf BUF1 (N2522, N2521);
or OR2 (N2523, N2508, N1827);
or OR3 (N2524, N2498, N1571, N2055);
not NOT1 (N2525, N2518);
buf BUF1 (N2526, N2517);
or OR4 (N2527, N2520, N2335, N148, N1441);
and AND4 (N2528, N2519, N2296, N1829, N1600);
buf BUF1 (N2529, N2509);
not NOT1 (N2530, N2526);
nor NOR3 (N2531, N2528, N352, N1511);
not NOT1 (N2532, N2525);
not NOT1 (N2533, N2483);
not NOT1 (N2534, N2533);
and AND2 (N2535, N2534, N1275);
or OR4 (N2536, N2524, N1449, N674, N1354);
nand NAND2 (N2537, N2530, N140);
and AND2 (N2538, N2516, N1614);
xor XOR2 (N2539, N2537, N2160);
and AND4 (N2540, N2522, N1383, N1298, N755);
or OR3 (N2541, N2531, N1685, N1208);
nand NAND2 (N2542, N2540, N632);
nand NAND2 (N2543, N2535, N257);
buf BUF1 (N2544, N2523);
not NOT1 (N2545, N2544);
not NOT1 (N2546, N2529);
or OR2 (N2547, N2536, N1900);
not NOT1 (N2548, N2547);
and AND3 (N2549, N2539, N516, N356);
nor NOR4 (N2550, N2527, N929, N1770, N2227);
nor NOR3 (N2551, N2541, N1706, N1737);
nor NOR2 (N2552, N2532, N328);
buf BUF1 (N2553, N2543);
xor XOR2 (N2554, N2548, N387);
or OR3 (N2555, N2549, N371, N2235);
buf BUF1 (N2556, N2546);
buf BUF1 (N2557, N2545);
not NOT1 (N2558, N2555);
or OR4 (N2559, N2550, N2447, N2358, N428);
and AND2 (N2560, N2556, N1086);
and AND4 (N2561, N2551, N1402, N842, N868);
or OR2 (N2562, N2560, N386);
and AND3 (N2563, N2559, N69, N488);
buf BUF1 (N2564, N2563);
not NOT1 (N2565, N2554);
xor XOR2 (N2566, N2552, N589);
xor XOR2 (N2567, N2558, N1314);
and AND2 (N2568, N2542, N1964);
not NOT1 (N2569, N2557);
not NOT1 (N2570, N2569);
nand NAND2 (N2571, N2570, N9);
nand NAND3 (N2572, N2571, N752, N1906);
not NOT1 (N2573, N2568);
not NOT1 (N2574, N2565);
xor XOR2 (N2575, N2572, N342);
nand NAND3 (N2576, N2573, N1791, N1670);
nor NOR2 (N2577, N2538, N1349);
not NOT1 (N2578, N2562);
xor XOR2 (N2579, N2578, N710);
buf BUF1 (N2580, N2564);
xor XOR2 (N2581, N2574, N280);
nor NOR3 (N2582, N2553, N677, N1481);
not NOT1 (N2583, N2561);
or OR4 (N2584, N2576, N1074, N1882, N661);
or OR2 (N2585, N2579, N384);
and AND2 (N2586, N2567, N1782);
and AND2 (N2587, N2586, N828);
xor XOR2 (N2588, N2575, N10);
or OR2 (N2589, N2566, N1040);
nor NOR2 (N2590, N2581, N1342);
and AND4 (N2591, N2577, N506, N1804, N17);
and AND4 (N2592, N2580, N1603, N1786, N1172);
xor XOR2 (N2593, N2589, N1659);
buf BUF1 (N2594, N2590);
nand NAND4 (N2595, N2588, N289, N2080, N1078);
buf BUF1 (N2596, N2587);
buf BUF1 (N2597, N2584);
buf BUF1 (N2598, N2583);
buf BUF1 (N2599, N2593);
or OR3 (N2600, N2591, N2337, N538);
buf BUF1 (N2601, N2595);
or OR2 (N2602, N2592, N2051);
or OR2 (N2603, N2601, N1494);
and AND2 (N2604, N2585, N2107);
buf BUF1 (N2605, N2600);
or OR4 (N2606, N2582, N1932, N2406, N126);
nor NOR4 (N2607, N2605, N550, N1819, N458);
not NOT1 (N2608, N2599);
nand NAND2 (N2609, N2596, N493);
and AND3 (N2610, N2603, N2437, N1210);
and AND4 (N2611, N2604, N2107, N1095, N1792);
buf BUF1 (N2612, N2611);
xor XOR2 (N2613, N2594, N1984);
or OR2 (N2614, N2612, N1793);
xor XOR2 (N2615, N2606, N2015);
nor NOR3 (N2616, N2598, N2337, N2318);
not NOT1 (N2617, N2597);
not NOT1 (N2618, N2607);
buf BUF1 (N2619, N2608);
or OR2 (N2620, N2615, N2083);
buf BUF1 (N2621, N2620);
and AND4 (N2622, N2617, N751, N917, N2490);
xor XOR2 (N2623, N2613, N2006);
nor NOR2 (N2624, N2619, N2280);
nand NAND3 (N2625, N2624, N1052, N1106);
or OR3 (N2626, N2602, N773, N467);
buf BUF1 (N2627, N2622);
nor NOR2 (N2628, N2623, N1680);
and AND2 (N2629, N2610, N756);
nor NOR4 (N2630, N2626, N546, N479, N1580);
buf BUF1 (N2631, N2630);
and AND4 (N2632, N2614, N235, N2490, N418);
buf BUF1 (N2633, N2609);
or OR3 (N2634, N2631, N2033, N1916);
nor NOR2 (N2635, N2627, N1591);
or OR2 (N2636, N2616, N2466);
or OR2 (N2637, N2628, N1518);
buf BUF1 (N2638, N2634);
and AND4 (N2639, N2637, N1756, N4, N459);
buf BUF1 (N2640, N2625);
or OR4 (N2641, N2635, N2163, N2538, N1874);
not NOT1 (N2642, N2632);
buf BUF1 (N2643, N2640);
nor NOR3 (N2644, N2629, N1484, N141);
xor XOR2 (N2645, N2642, N2118);
or OR4 (N2646, N2643, N2272, N277, N2618);
nand NAND4 (N2647, N876, N2220, N2521, N2361);
or OR2 (N2648, N2639, N2122);
xor XOR2 (N2649, N2646, N862);
and AND2 (N2650, N2648, N11);
and AND4 (N2651, N2650, N1667, N28, N48);
xor XOR2 (N2652, N2649, N340);
buf BUF1 (N2653, N2645);
xor XOR2 (N2654, N2652, N535);
xor XOR2 (N2655, N2644, N1721);
not NOT1 (N2656, N2633);
or OR3 (N2657, N2653, N1418, N717);
buf BUF1 (N2658, N2655);
or OR3 (N2659, N2658, N2390, N1078);
nand NAND2 (N2660, N2641, N2141);
nor NOR3 (N2661, N2638, N179, N1804);
buf BUF1 (N2662, N2654);
not NOT1 (N2663, N2656);
buf BUF1 (N2664, N2657);
buf BUF1 (N2665, N2636);
nor NOR3 (N2666, N2663, N572, N154);
nand NAND2 (N2667, N2662, N1169);
buf BUF1 (N2668, N2661);
not NOT1 (N2669, N2666);
nand NAND3 (N2670, N2621, N2534, N844);
xor XOR2 (N2671, N2664, N50);
xor XOR2 (N2672, N2667, N863);
and AND2 (N2673, N2660, N1458);
or OR4 (N2674, N2669, N1264, N1493, N492);
nand NAND2 (N2675, N2671, N273);
xor XOR2 (N2676, N2674, N505);
xor XOR2 (N2677, N2651, N289);
nor NOR2 (N2678, N2659, N1047);
nor NOR3 (N2679, N2678, N591, N656);
xor XOR2 (N2680, N2665, N92);
not NOT1 (N2681, N2670);
xor XOR2 (N2682, N2647, N1917);
and AND2 (N2683, N2680, N712);
not NOT1 (N2684, N2682);
or OR2 (N2685, N2684, N2499);
not NOT1 (N2686, N2668);
nor NOR4 (N2687, N2683, N1604, N1562, N1208);
and AND3 (N2688, N2673, N446, N554);
or OR3 (N2689, N2672, N2126, N2079);
nor NOR4 (N2690, N2675, N2339, N2135, N2607);
nor NOR4 (N2691, N2687, N668, N1943, N2330);
nand NAND4 (N2692, N2689, N2310, N1360, N917);
and AND4 (N2693, N2681, N1974, N1411, N1706);
xor XOR2 (N2694, N2679, N2332);
or OR4 (N2695, N2677, N399, N1268, N2496);
nand NAND3 (N2696, N2685, N29, N1776);
xor XOR2 (N2697, N2691, N2547);
and AND3 (N2698, N2697, N1555, N1882);
and AND3 (N2699, N2692, N1450, N2082);
xor XOR2 (N2700, N2688, N1419);
and AND4 (N2701, N2693, N900, N1445, N30);
xor XOR2 (N2702, N2701, N1526);
xor XOR2 (N2703, N2686, N1650);
or OR2 (N2704, N2695, N561);
nand NAND2 (N2705, N2696, N1741);
buf BUF1 (N2706, N2703);
nor NOR4 (N2707, N2700, N885, N1218, N814);
nor NOR2 (N2708, N2702, N1212);
nand NAND2 (N2709, N2704, N2644);
and AND2 (N2710, N2706, N460);
not NOT1 (N2711, N2708);
buf BUF1 (N2712, N2694);
or OR3 (N2713, N2712, N405, N2251);
nand NAND2 (N2714, N2698, N1580);
or OR3 (N2715, N2690, N372, N1984);
xor XOR2 (N2716, N2707, N2416);
buf BUF1 (N2717, N2713);
nor NOR2 (N2718, N2717, N1726);
nor NOR3 (N2719, N2718, N1317, N1059);
or OR3 (N2720, N2711, N2524, N717);
and AND4 (N2721, N2705, N537, N120, N1125);
or OR3 (N2722, N2721, N694, N1551);
nand NAND2 (N2723, N2710, N435);
and AND4 (N2724, N2719, N739, N350, N42);
and AND4 (N2725, N2724, N1979, N590, N779);
not NOT1 (N2726, N2714);
xor XOR2 (N2727, N2699, N1360);
nor NOR4 (N2728, N2725, N63, N593, N2082);
buf BUF1 (N2729, N2715);
and AND4 (N2730, N2720, N199, N1333, N2663);
buf BUF1 (N2731, N2727);
buf BUF1 (N2732, N2726);
buf BUF1 (N2733, N2722);
buf BUF1 (N2734, N2728);
or OR4 (N2735, N2734, N1995, N716, N1422);
or OR4 (N2736, N2732, N187, N1922, N843);
and AND3 (N2737, N2709, N1176, N385);
xor XOR2 (N2738, N2733, N1757);
and AND4 (N2739, N2730, N215, N2715, N2543);
nor NOR2 (N2740, N2716, N2359);
and AND4 (N2741, N2739, N1254, N1974, N2138);
not NOT1 (N2742, N2736);
and AND4 (N2743, N2676, N24, N2727, N2185);
not NOT1 (N2744, N2740);
or OR3 (N2745, N2737, N249, N2384);
xor XOR2 (N2746, N2735, N1182);
buf BUF1 (N2747, N2731);
or OR3 (N2748, N2742, N48, N314);
not NOT1 (N2749, N2738);
nand NAND2 (N2750, N2745, N1180);
xor XOR2 (N2751, N2748, N953);
not NOT1 (N2752, N2749);
or OR3 (N2753, N2752, N1842, N1991);
nand NAND3 (N2754, N2751, N461, N2172);
nand NAND4 (N2755, N2743, N1818, N1750, N2033);
xor XOR2 (N2756, N2723, N1903);
buf BUF1 (N2757, N2754);
nor NOR4 (N2758, N2753, N2474, N399, N1584);
or OR3 (N2759, N2744, N291, N2392);
nor NOR2 (N2760, N2755, N774);
buf BUF1 (N2761, N2750);
not NOT1 (N2762, N2759);
not NOT1 (N2763, N2757);
nand NAND3 (N2764, N2741, N1680, N406);
nor NOR3 (N2765, N2747, N319, N2003);
nor NOR4 (N2766, N2761, N1659, N1644, N1115);
buf BUF1 (N2767, N2764);
xor XOR2 (N2768, N2760, N2408);
not NOT1 (N2769, N2763);
buf BUF1 (N2770, N2767);
and AND2 (N2771, N2765, N1904);
nand NAND4 (N2772, N2762, N1657, N667, N2637);
xor XOR2 (N2773, N2746, N480);
and AND4 (N2774, N2770, N765, N585, N2320);
nor NOR3 (N2775, N2773, N2653, N2063);
nand NAND2 (N2776, N2775, N1953);
not NOT1 (N2777, N2766);
nand NAND3 (N2778, N2777, N2291, N2030);
buf BUF1 (N2779, N2729);
nor NOR4 (N2780, N2776, N1414, N2066, N1762);
or OR3 (N2781, N2772, N549, N1523);
or OR4 (N2782, N2758, N130, N889, N1487);
and AND3 (N2783, N2782, N726, N2177);
xor XOR2 (N2784, N2771, N2755);
or OR3 (N2785, N2774, N1959, N2102);
or OR4 (N2786, N2783, N2404, N1328, N818);
xor XOR2 (N2787, N2769, N1028);
not NOT1 (N2788, N2780);
nand NAND3 (N2789, N2779, N2710, N1811);
or OR4 (N2790, N2789, N1522, N749, N2719);
buf BUF1 (N2791, N2784);
and AND4 (N2792, N2768, N731, N1932, N1683);
buf BUF1 (N2793, N2787);
xor XOR2 (N2794, N2788, N2603);
or OR3 (N2795, N2778, N1062, N656);
xor XOR2 (N2796, N2794, N1491);
nand NAND4 (N2797, N2785, N132, N761, N2314);
buf BUF1 (N2798, N2792);
nor NOR2 (N2799, N2795, N169);
or OR2 (N2800, N2791, N1581);
buf BUF1 (N2801, N2793);
or OR3 (N2802, N2799, N2230, N433);
not NOT1 (N2803, N2797);
or OR2 (N2804, N2800, N2384);
nand NAND4 (N2805, N2803, N1494, N2337, N1606);
nor NOR4 (N2806, N2802, N1794, N1462, N849);
and AND3 (N2807, N2801, N1634, N2107);
nand NAND4 (N2808, N2756, N1033, N2215, N2273);
nor NOR2 (N2809, N2808, N825);
nor NOR2 (N2810, N2798, N1901);
and AND3 (N2811, N2786, N338, N833);
or OR4 (N2812, N2809, N1398, N310, N1773);
nand NAND3 (N2813, N2810, N975, N314);
buf BUF1 (N2814, N2790);
xor XOR2 (N2815, N2813, N2625);
nand NAND4 (N2816, N2781, N826, N2680, N2382);
nor NOR4 (N2817, N2811, N119, N2059, N952);
nand NAND4 (N2818, N2807, N1497, N2609, N1474);
and AND3 (N2819, N2815, N1650, N1645);
xor XOR2 (N2820, N2818, N1082);
xor XOR2 (N2821, N2804, N984);
not NOT1 (N2822, N2814);
not NOT1 (N2823, N2819);
nor NOR4 (N2824, N2805, N613, N1556, N225);
or OR3 (N2825, N2796, N307, N1347);
buf BUF1 (N2826, N2820);
and AND3 (N2827, N2806, N947, N2455);
or OR3 (N2828, N2822, N2713, N1566);
buf BUF1 (N2829, N2812);
xor XOR2 (N2830, N2824, N1053);
nand NAND2 (N2831, N2826, N2360);
or OR2 (N2832, N2831, N1092);
nor NOR3 (N2833, N2830, N166, N404);
or OR3 (N2834, N2827, N2786, N1685);
nand NAND2 (N2835, N2832, N155);
buf BUF1 (N2836, N2816);
nor NOR3 (N2837, N2821, N658, N1370);
xor XOR2 (N2838, N2829, N1351);
xor XOR2 (N2839, N2825, N1358);
and AND2 (N2840, N2833, N10);
xor XOR2 (N2841, N2840, N1558);
not NOT1 (N2842, N2834);
nor NOR3 (N2843, N2823, N2335, N1287);
buf BUF1 (N2844, N2837);
buf BUF1 (N2845, N2841);
and AND4 (N2846, N2839, N827, N2315, N2444);
buf BUF1 (N2847, N2836);
buf BUF1 (N2848, N2828);
and AND2 (N2849, N2843, N2464);
or OR3 (N2850, N2844, N1967, N2537);
nor NOR3 (N2851, N2849, N1554, N1352);
or OR3 (N2852, N2850, N2031, N2366);
xor XOR2 (N2853, N2852, N463);
and AND2 (N2854, N2817, N513);
nand NAND4 (N2855, N2838, N2777, N1690, N215);
nor NOR2 (N2856, N2848, N791);
nor NOR3 (N2857, N2855, N815, N876);
buf BUF1 (N2858, N2851);
or OR4 (N2859, N2846, N1312, N1112, N1725);
nor NOR2 (N2860, N2853, N2308);
buf BUF1 (N2861, N2857);
xor XOR2 (N2862, N2842, N870);
nor NOR4 (N2863, N2862, N1212, N1569, N2504);
buf BUF1 (N2864, N2835);
and AND3 (N2865, N2845, N1169, N863);
nor NOR4 (N2866, N2856, N1641, N1136, N1920);
nand NAND4 (N2867, N2861, N1498, N1826, N1308);
not NOT1 (N2868, N2858);
or OR3 (N2869, N2864, N649, N2329);
or OR4 (N2870, N2860, N2695, N2160, N469);
buf BUF1 (N2871, N2863);
or OR4 (N2872, N2868, N2583, N354, N858);
nand NAND4 (N2873, N2872, N1794, N2472, N1289);
and AND4 (N2874, N2867, N2634, N56, N596);
xor XOR2 (N2875, N2859, N496);
buf BUF1 (N2876, N2854);
nand NAND4 (N2877, N2869, N1533, N1856, N2603);
buf BUF1 (N2878, N2847);
nand NAND4 (N2879, N2875, N315, N198, N1704);
xor XOR2 (N2880, N2871, N1769);
and AND3 (N2881, N2880, N2481, N1141);
nor NOR3 (N2882, N2876, N1482, N2165);
or OR3 (N2883, N2870, N1014, N2681);
xor XOR2 (N2884, N2873, N2642);
nand NAND3 (N2885, N2881, N789, N2848);
buf BUF1 (N2886, N2882);
buf BUF1 (N2887, N2874);
xor XOR2 (N2888, N2884, N1250);
nand NAND3 (N2889, N2885, N2626, N1725);
not NOT1 (N2890, N2879);
xor XOR2 (N2891, N2886, N419);
nand NAND2 (N2892, N2889, N1102);
and AND3 (N2893, N2877, N1126, N1858);
xor XOR2 (N2894, N2887, N2584);
and AND3 (N2895, N2891, N1397, N2085);
nand NAND2 (N2896, N2893, N913);
xor XOR2 (N2897, N2883, N1934);
buf BUF1 (N2898, N2888);
or OR2 (N2899, N2897, N2737);
xor XOR2 (N2900, N2896, N1455);
buf BUF1 (N2901, N2866);
or OR2 (N2902, N2865, N395);
or OR2 (N2903, N2902, N1104);
or OR2 (N2904, N2901, N336);
xor XOR2 (N2905, N2898, N1518);
nor NOR3 (N2906, N2904, N1453, N1218);
or OR4 (N2907, N2899, N729, N1884, N1464);
xor XOR2 (N2908, N2900, N2023);
xor XOR2 (N2909, N2907, N2506);
and AND3 (N2910, N2906, N2663, N643);
nor NOR3 (N2911, N2905, N1580, N580);
and AND2 (N2912, N2890, N1858);
or OR2 (N2913, N2909, N1636);
nor NOR3 (N2914, N2911, N2259, N2745);
buf BUF1 (N2915, N2913);
or OR3 (N2916, N2895, N2902, N733);
not NOT1 (N2917, N2916);
buf BUF1 (N2918, N2894);
nor NOR4 (N2919, N2918, N2166, N2577, N2736);
not NOT1 (N2920, N2915);
not NOT1 (N2921, N2892);
nor NOR2 (N2922, N2903, N865);
and AND2 (N2923, N2919, N1596);
nor NOR2 (N2924, N2878, N1470);
xor XOR2 (N2925, N2923, N2730);
buf BUF1 (N2926, N2910);
and AND4 (N2927, N2926, N2051, N2230, N1263);
and AND2 (N2928, N2927, N2704);
or OR2 (N2929, N2924, N1344);
xor XOR2 (N2930, N2908, N1453);
xor XOR2 (N2931, N2930, N279);
xor XOR2 (N2932, N2931, N2108);
nor NOR2 (N2933, N2917, N1932);
and AND4 (N2934, N2929, N2443, N1768, N2337);
and AND2 (N2935, N2920, N908);
not NOT1 (N2936, N2935);
not NOT1 (N2937, N2914);
and AND4 (N2938, N2921, N2009, N197, N2009);
and AND2 (N2939, N2912, N2713);
xor XOR2 (N2940, N2922, N1838);
nand NAND3 (N2941, N2938, N1222, N1717);
nand NAND4 (N2942, N2932, N1502, N1484, N353);
and AND2 (N2943, N2937, N34);
or OR2 (N2944, N2939, N1926);
and AND2 (N2945, N2925, N18);
nand NAND3 (N2946, N2933, N1525, N888);
or OR2 (N2947, N2934, N2050);
xor XOR2 (N2948, N2945, N146);
not NOT1 (N2949, N2946);
nor NOR4 (N2950, N2948, N2034, N2691, N1018);
nand NAND4 (N2951, N2949, N257, N397, N484);
buf BUF1 (N2952, N2947);
nor NOR2 (N2953, N2943, N1571);
buf BUF1 (N2954, N2940);
and AND2 (N2955, N2936, N1691);
not NOT1 (N2956, N2941);
nand NAND2 (N2957, N2950, N2015);
buf BUF1 (N2958, N2944);
or OR2 (N2959, N2956, N1218);
and AND3 (N2960, N2959, N1636, N1775);
and AND2 (N2961, N2952, N797);
nor NOR2 (N2962, N2928, N1544);
xor XOR2 (N2963, N2958, N1020);
or OR2 (N2964, N2961, N482);
buf BUF1 (N2965, N2955);
buf BUF1 (N2966, N2942);
nand NAND2 (N2967, N2953, N1364);
buf BUF1 (N2968, N2960);
or OR4 (N2969, N2962, N2480, N2254, N2137);
nand NAND2 (N2970, N2964, N2168);
xor XOR2 (N2971, N2965, N2024);
or OR3 (N2972, N2969, N1955, N1670);
nand NAND4 (N2973, N2970, N327, N2836, N2607);
buf BUF1 (N2974, N2951);
and AND4 (N2975, N2957, N2164, N1233, N2724);
nand NAND3 (N2976, N2971, N2427, N744);
nand NAND2 (N2977, N2974, N1776);
or OR3 (N2978, N2975, N171, N1415);
or OR2 (N2979, N2963, N2377);
xor XOR2 (N2980, N2976, N2435);
nand NAND3 (N2981, N2979, N2019, N619);
and AND4 (N2982, N2977, N502, N797, N2862);
and AND3 (N2983, N2967, N2976, N2965);
xor XOR2 (N2984, N2972, N433);
buf BUF1 (N2985, N2973);
buf BUF1 (N2986, N2981);
and AND4 (N2987, N2954, N2866, N1161, N185);
and AND4 (N2988, N2982, N846, N2089, N330);
buf BUF1 (N2989, N2966);
not NOT1 (N2990, N2987);
buf BUF1 (N2991, N2978);
xor XOR2 (N2992, N2985, N224);
and AND3 (N2993, N2986, N225, N1660);
buf BUF1 (N2994, N2984);
or OR2 (N2995, N2980, N2166);
not NOT1 (N2996, N2989);
nand NAND4 (N2997, N2994, N2071, N1839, N1181);
not NOT1 (N2998, N2991);
or OR3 (N2999, N2988, N2115, N259);
or OR3 (N3000, N2993, N766, N2794);
not NOT1 (N3001, N2968);
xor XOR2 (N3002, N2998, N585);
buf BUF1 (N3003, N3002);
buf BUF1 (N3004, N2997);
nand NAND3 (N3005, N3003, N2874, N2776);
or OR3 (N3006, N2995, N1970, N615);
or OR3 (N3007, N3000, N1325, N1677);
nor NOR2 (N3008, N3005, N475);
and AND2 (N3009, N3001, N2833);
buf BUF1 (N3010, N2983);
not NOT1 (N3011, N3007);
xor XOR2 (N3012, N2990, N241);
or OR3 (N3013, N3008, N797, N1467);
buf BUF1 (N3014, N3011);
not NOT1 (N3015, N3010);
nor NOR3 (N3016, N3015, N647, N1890);
xor XOR2 (N3017, N3012, N2867);
and AND4 (N3018, N2999, N1290, N238, N1278);
nand NAND2 (N3019, N3006, N718);
not NOT1 (N3020, N3017);
or OR4 (N3021, N3020, N2926, N2417, N867);
buf BUF1 (N3022, N2992);
nand NAND3 (N3023, N3013, N2779, N158);
or OR3 (N3024, N3016, N13, N2224);
not NOT1 (N3025, N3004);
and AND3 (N3026, N3019, N479, N869);
xor XOR2 (N3027, N3018, N218);
and AND2 (N3028, N3024, N2818);
buf BUF1 (N3029, N3025);
nor NOR4 (N3030, N3014, N2727, N2955, N1731);
xor XOR2 (N3031, N3022, N1849);
xor XOR2 (N3032, N2996, N1622);
nor NOR2 (N3033, N3027, N460);
and AND2 (N3034, N3032, N617);
xor XOR2 (N3035, N3030, N2272);
not NOT1 (N3036, N3031);
not NOT1 (N3037, N3034);
nor NOR3 (N3038, N3026, N2714, N549);
buf BUF1 (N3039, N3033);
buf BUF1 (N3040, N3035);
nand NAND4 (N3041, N3039, N149, N1651, N2195);
not NOT1 (N3042, N3040);
or OR2 (N3043, N3009, N2076);
nand NAND2 (N3044, N3029, N152);
xor XOR2 (N3045, N3044, N1557);
nor NOR2 (N3046, N3045, N2781);
nor NOR2 (N3047, N3046, N1580);
not NOT1 (N3048, N3043);
not NOT1 (N3049, N3041);
buf BUF1 (N3050, N3036);
nand NAND4 (N3051, N3050, N1318, N2325, N2121);
xor XOR2 (N3052, N3037, N2537);
nand NAND2 (N3053, N3042, N1652);
nor NOR3 (N3054, N3028, N2610, N1388);
not NOT1 (N3055, N3048);
or OR3 (N3056, N3023, N937, N2131);
nor NOR2 (N3057, N3021, N1931);
xor XOR2 (N3058, N3056, N2019);
xor XOR2 (N3059, N3049, N2781);
not NOT1 (N3060, N3054);
nor NOR4 (N3061, N3057, N932, N433, N254);
nand NAND4 (N3062, N3060, N2041, N2596, N2817);
not NOT1 (N3063, N3055);
and AND2 (N3064, N3052, N2829);
xor XOR2 (N3065, N3051, N2744);
nor NOR3 (N3066, N3038, N2970, N823);
or OR3 (N3067, N3063, N144, N1097);
nor NOR4 (N3068, N3065, N389, N528, N1076);
and AND2 (N3069, N3064, N139);
not NOT1 (N3070, N3067);
xor XOR2 (N3071, N3068, N262);
buf BUF1 (N3072, N3069);
and AND4 (N3073, N3070, N2139, N47, N995);
not NOT1 (N3074, N3061);
and AND2 (N3075, N3047, N1491);
nor NOR3 (N3076, N3058, N1914, N2);
nand NAND2 (N3077, N3073, N2712);
not NOT1 (N3078, N3053);
buf BUF1 (N3079, N3075);
or OR4 (N3080, N3078, N2033, N97, N468);
or OR3 (N3081, N3074, N2957, N328);
or OR4 (N3082, N3079, N1171, N1670, N2041);
xor XOR2 (N3083, N3077, N176);
nand NAND4 (N3084, N3076, N1096, N2542, N243);
nand NAND2 (N3085, N3082, N1497);
not NOT1 (N3086, N3072);
buf BUF1 (N3087, N3081);
nand NAND3 (N3088, N3062, N726, N2481);
buf BUF1 (N3089, N3059);
nand NAND4 (N3090, N3080, N3067, N2229, N876);
not NOT1 (N3091, N3090);
not NOT1 (N3092, N3088);
not NOT1 (N3093, N3092);
nor NOR2 (N3094, N3087, N2345);
nand NAND2 (N3095, N3093, N2705);
or OR4 (N3096, N3095, N2990, N1536, N3067);
and AND3 (N3097, N3085, N536, N2521);
or OR4 (N3098, N3094, N2096, N2227, N1526);
xor XOR2 (N3099, N3091, N342);
not NOT1 (N3100, N3096);
xor XOR2 (N3101, N3089, N1315);
nand NAND3 (N3102, N3101, N1704, N867);
or OR4 (N3103, N3099, N1649, N2710, N1979);
not NOT1 (N3104, N3103);
nor NOR2 (N3105, N3098, N1475);
nor NOR2 (N3106, N3071, N2249);
not NOT1 (N3107, N3105);
or OR2 (N3108, N3107, N753);
xor XOR2 (N3109, N3066, N774);
or OR3 (N3110, N3109, N1747, N3020);
xor XOR2 (N3111, N3106, N1507);
xor XOR2 (N3112, N3084, N384);
not NOT1 (N3113, N3100);
not NOT1 (N3114, N3111);
nand NAND3 (N3115, N3104, N1314, N2619);
not NOT1 (N3116, N3114);
and AND3 (N3117, N3112, N2488, N2325);
xor XOR2 (N3118, N3086, N1576);
nand NAND3 (N3119, N3113, N1681, N1846);
nor NOR2 (N3120, N3118, N1371);
and AND4 (N3121, N3120, N1402, N531, N2722);
not NOT1 (N3122, N3117);
nor NOR4 (N3123, N3121, N1846, N762, N2731);
nor NOR4 (N3124, N3122, N613, N1468, N2433);
not NOT1 (N3125, N3108);
xor XOR2 (N3126, N3116, N2716);
or OR4 (N3127, N3126, N2917, N1472, N2423);
not NOT1 (N3128, N3119);
nand NAND3 (N3129, N3083, N1247, N111);
not NOT1 (N3130, N3128);
or OR3 (N3131, N3097, N1163, N1158);
buf BUF1 (N3132, N3102);
buf BUF1 (N3133, N3131);
nor NOR4 (N3134, N3130, N2053, N1807, N710);
or OR2 (N3135, N3134, N2967);
or OR2 (N3136, N3125, N214);
or OR2 (N3137, N3127, N1479);
not NOT1 (N3138, N3135);
and AND3 (N3139, N3137, N273, N500);
buf BUF1 (N3140, N3123);
nand NAND4 (N3141, N3136, N1612, N2203, N58);
buf BUF1 (N3142, N3110);
and AND2 (N3143, N3132, N1587);
nor NOR3 (N3144, N3140, N686, N2781);
and AND3 (N3145, N3115, N481, N676);
buf BUF1 (N3146, N3144);
xor XOR2 (N3147, N3141, N2392);
buf BUF1 (N3148, N3147);
nor NOR3 (N3149, N3139, N3011, N1116);
buf BUF1 (N3150, N3129);
and AND4 (N3151, N3124, N1972, N1268, N883);
or OR3 (N3152, N3151, N502, N323);
and AND4 (N3153, N3146, N807, N2313, N781);
buf BUF1 (N3154, N3150);
not NOT1 (N3155, N3145);
xor XOR2 (N3156, N3152, N2184);
not NOT1 (N3157, N3148);
and AND3 (N3158, N3142, N1810, N2600);
not NOT1 (N3159, N3153);
nor NOR4 (N3160, N3157, N501, N1050, N2622);
or OR4 (N3161, N3156, N1691, N1831, N2574);
or OR4 (N3162, N3149, N3134, N1915, N2538);
or OR2 (N3163, N3138, N459);
nand NAND4 (N3164, N3160, N714, N2683, N2346);
or OR2 (N3165, N3162, N2741);
nor NOR2 (N3166, N3165, N1314);
buf BUF1 (N3167, N3159);
buf BUF1 (N3168, N3167);
or OR3 (N3169, N3166, N2130, N2499);
nand NAND2 (N3170, N3168, N2910);
nor NOR3 (N3171, N3133, N300, N1771);
not NOT1 (N3172, N3161);
buf BUF1 (N3173, N3172);
nand NAND4 (N3174, N3171, N1825, N2771, N2363);
nand NAND4 (N3175, N3155, N440, N1902, N1695);
or OR2 (N3176, N3169, N176);
not NOT1 (N3177, N3143);
nand NAND4 (N3178, N3174, N517, N1409, N763);
not NOT1 (N3179, N3173);
xor XOR2 (N3180, N3154, N2140);
or OR3 (N3181, N3158, N2095, N885);
nand NAND4 (N3182, N3177, N3087, N2359, N839);
or OR4 (N3183, N3176, N2705, N3037, N2000);
buf BUF1 (N3184, N3178);
nand NAND2 (N3185, N3182, N2290);
and AND3 (N3186, N3164, N2293, N92);
nor NOR2 (N3187, N3185, N186);
not NOT1 (N3188, N3184);
nor NOR2 (N3189, N3170, N638);
nand NAND2 (N3190, N3175, N1816);
not NOT1 (N3191, N3163);
and AND2 (N3192, N3187, N16);
nand NAND2 (N3193, N3190, N562);
and AND3 (N3194, N3192, N1037, N2683);
nor NOR4 (N3195, N3194, N2350, N1868, N2564);
or OR3 (N3196, N3180, N2214, N1494);
and AND3 (N3197, N3196, N2399, N2604);
or OR2 (N3198, N3188, N1658);
buf BUF1 (N3199, N3181);
buf BUF1 (N3200, N3191);
buf BUF1 (N3201, N3195);
nor NOR3 (N3202, N3186, N1186, N2525);
or OR4 (N3203, N3198, N2165, N2260, N2349);
nor NOR4 (N3204, N3203, N1629, N1600, N687);
not NOT1 (N3205, N3204);
nor NOR4 (N3206, N3183, N2191, N1250, N2834);
and AND4 (N3207, N3201, N548, N2712, N1163);
nor NOR4 (N3208, N3193, N1097, N1614, N826);
xor XOR2 (N3209, N3206, N565);
and AND3 (N3210, N3208, N216, N608);
or OR2 (N3211, N3199, N1037);
and AND3 (N3212, N3207, N2985, N1597);
nand NAND2 (N3213, N3211, N1731);
not NOT1 (N3214, N3209);
and AND2 (N3215, N3214, N666);
xor XOR2 (N3216, N3202, N460);
not NOT1 (N3217, N3210);
xor XOR2 (N3218, N3179, N2055);
nand NAND3 (N3219, N3205, N2091, N890);
nand NAND4 (N3220, N3213, N1763, N3129, N3099);
and AND2 (N3221, N3212, N934);
and AND2 (N3222, N3217, N2399);
nor NOR3 (N3223, N3220, N3030, N2941);
nor NOR2 (N3224, N3216, N2339);
endmodule