// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12;

output N16003,N16009,N16008,N16010,N16001,N15995,N16005,N15999,N15994,N16012;

buf BUF1 (N13, N3);
xor XOR2 (N14, N13, N10);
not NOT1 (N15, N1);
or OR3 (N16, N4, N8, N15);
buf BUF1 (N17, N15);
or OR4 (N18, N8, N5, N10, N1);
not NOT1 (N19, N7);
not NOT1 (N20, N17);
nor NOR4 (N21, N18, N11, N5, N3);
or OR4 (N22, N13, N1, N17, N3);
not NOT1 (N23, N4);
buf BUF1 (N24, N23);
not NOT1 (N25, N20);
nor NOR3 (N26, N6, N2, N6);
buf BUF1 (N27, N12);
or OR2 (N28, N1, N8);
not NOT1 (N29, N14);
and AND2 (N30, N24, N22);
and AND3 (N31, N13, N20, N13);
buf BUF1 (N32, N27);
nand NAND2 (N33, N19, N27);
or OR3 (N34, N16, N31, N6);
not NOT1 (N35, N5);
not NOT1 (N36, N32);
and AND4 (N37, N21, N29, N17, N20);
or OR2 (N38, N12, N34);
nor NOR3 (N39, N35, N15, N38);
and AND3 (N40, N20, N7, N6);
not NOT1 (N41, N26);
xor XOR2 (N42, N20, N29);
and AND2 (N43, N41, N27);
or OR4 (N44, N40, N35, N8, N15);
buf BUF1 (N45, N33);
nor NOR3 (N46, N43, N41, N1);
nor NOR3 (N47, N37, N27, N35);
xor XOR2 (N48, N39, N22);
nor NOR4 (N49, N48, N48, N10, N27);
nor NOR4 (N50, N47, N5, N8, N14);
nor NOR2 (N51, N42, N22);
nand NAND2 (N52, N51, N2);
nor NOR2 (N53, N36, N14);
nand NAND4 (N54, N44, N1, N15, N5);
or OR2 (N55, N28, N32);
or OR4 (N56, N30, N54, N2, N28);
not NOT1 (N57, N45);
xor XOR2 (N58, N17, N20);
nand NAND2 (N59, N57, N9);
not NOT1 (N60, N56);
buf BUF1 (N61, N52);
nand NAND3 (N62, N55, N18, N11);
not NOT1 (N63, N62);
buf BUF1 (N64, N60);
nor NOR2 (N65, N50, N31);
or OR4 (N66, N59, N53, N19, N41);
and AND4 (N67, N57, N56, N37, N3);
or OR4 (N68, N61, N25, N34, N64);
nand NAND2 (N69, N65, N42);
or OR2 (N70, N9, N41);
xor XOR2 (N71, N55, N26);
not NOT1 (N72, N63);
nor NOR3 (N73, N49, N11, N72);
not NOT1 (N74, N53);
and AND2 (N75, N68, N48);
nand NAND2 (N76, N71, N44);
not NOT1 (N77, N58);
buf BUF1 (N78, N75);
xor XOR2 (N79, N69, N20);
and AND4 (N80, N66, N19, N36, N63);
nor NOR4 (N81, N70, N70, N15, N7);
nand NAND2 (N82, N77, N32);
nor NOR4 (N83, N74, N61, N46, N62);
not NOT1 (N84, N42);
xor XOR2 (N85, N83, N82);
xor XOR2 (N86, N10, N37);
and AND2 (N87, N81, N51);
or OR4 (N88, N78, N24, N71, N36);
nand NAND4 (N89, N76, N87, N49, N22);
nand NAND3 (N90, N13, N32, N50);
nand NAND2 (N91, N79, N73);
buf BUF1 (N92, N8);
or OR2 (N93, N91, N82);
nor NOR2 (N94, N90, N45);
nand NAND4 (N95, N84, N47, N9, N74);
not NOT1 (N96, N89);
nand NAND2 (N97, N80, N8);
and AND4 (N98, N88, N16, N61, N64);
nor NOR2 (N99, N95, N10);
nand NAND4 (N100, N85, N76, N67, N10);
xor XOR2 (N101, N62, N27);
nand NAND2 (N102, N86, N51);
nor NOR4 (N103, N98, N82, N77, N55);
buf BUF1 (N104, N94);
nand NAND2 (N105, N101, N11);
nand NAND3 (N106, N92, N14, N43);
nor NOR4 (N107, N100, N76, N36, N98);
xor XOR2 (N108, N103, N14);
buf BUF1 (N109, N108);
nor NOR3 (N110, N102, N31, N54);
buf BUF1 (N111, N97);
nor NOR3 (N112, N99, N6, N35);
xor XOR2 (N113, N96, N20);
not NOT1 (N114, N111);
buf BUF1 (N115, N106);
and AND3 (N116, N113, N76, N70);
nand NAND4 (N117, N114, N34, N75, N45);
and AND2 (N118, N115, N62);
buf BUF1 (N119, N112);
nand NAND4 (N120, N119, N43, N118, N24);
or OR2 (N121, N32, N89);
or OR3 (N122, N120, N42, N12);
and AND4 (N123, N121, N60, N39, N49);
nand NAND3 (N124, N104, N38, N107);
nor NOR2 (N125, N58, N6);
not NOT1 (N126, N124);
and AND2 (N127, N125, N93);
or OR4 (N128, N114, N62, N32, N15);
nand NAND2 (N129, N116, N98);
or OR4 (N130, N105, N97, N64, N31);
not NOT1 (N131, N123);
buf BUF1 (N132, N127);
or OR3 (N133, N129, N11, N26);
nor NOR3 (N134, N132, N25, N56);
nand NAND4 (N135, N133, N57, N121, N68);
buf BUF1 (N136, N122);
and AND2 (N137, N110, N109);
not NOT1 (N138, N37);
nand NAND2 (N139, N136, N125);
nor NOR4 (N140, N137, N32, N5, N30);
buf BUF1 (N141, N139);
or OR4 (N142, N131, N133, N138, N33);
and AND2 (N143, N17, N122);
not NOT1 (N144, N142);
xor XOR2 (N145, N140, N108);
xor XOR2 (N146, N117, N43);
nor NOR4 (N147, N128, N17, N113, N101);
or OR4 (N148, N147, N147, N111, N11);
buf BUF1 (N149, N144);
nor NOR4 (N150, N130, N88, N70, N54);
or OR2 (N151, N135, N97);
nand NAND3 (N152, N143, N53, N79);
or OR2 (N153, N148, N22);
and AND4 (N154, N153, N87, N83, N14);
not NOT1 (N155, N154);
buf BUF1 (N156, N150);
and AND3 (N157, N126, N48, N152);
not NOT1 (N158, N156);
and AND4 (N159, N112, N87, N31, N32);
nor NOR4 (N160, N134, N37, N39, N92);
and AND2 (N161, N146, N103);
buf BUF1 (N162, N161);
xor XOR2 (N163, N160, N116);
and AND4 (N164, N158, N109, N116, N124);
not NOT1 (N165, N157);
or OR3 (N166, N162, N118, N45);
not NOT1 (N167, N159);
nor NOR3 (N168, N141, N83, N52);
and AND2 (N169, N168, N25);
and AND2 (N170, N169, N5);
or OR3 (N171, N167, N8, N152);
or OR3 (N172, N165, N72, N90);
or OR2 (N173, N155, N101);
not NOT1 (N174, N173);
or OR3 (N175, N170, N104, N61);
nand NAND4 (N176, N172, N71, N78, N47);
buf BUF1 (N177, N149);
buf BUF1 (N178, N176);
or OR4 (N179, N145, N10, N162, N134);
buf BUF1 (N180, N177);
or OR3 (N181, N171, N106, N46);
or OR4 (N182, N174, N178, N31, N74);
nor NOR3 (N183, N119, N178, N162);
xor XOR2 (N184, N166, N155);
nand NAND2 (N185, N164, N85);
nor NOR2 (N186, N151, N24);
nor NOR3 (N187, N180, N15, N29);
nand NAND2 (N188, N186, N56);
not NOT1 (N189, N183);
or OR4 (N190, N179, N61, N84, N108);
buf BUF1 (N191, N187);
and AND2 (N192, N184, N179);
buf BUF1 (N193, N163);
or OR3 (N194, N185, N153, N177);
and AND4 (N195, N181, N85, N64, N133);
not NOT1 (N196, N191);
and AND2 (N197, N195, N87);
buf BUF1 (N198, N193);
not NOT1 (N199, N197);
nand NAND4 (N200, N182, N10, N164, N45);
buf BUF1 (N201, N190);
or OR2 (N202, N192, N139);
or OR2 (N203, N202, N88);
nand NAND2 (N204, N203, N166);
nor NOR4 (N205, N201, N112, N103, N180);
not NOT1 (N206, N204);
and AND4 (N207, N189, N157, N24, N133);
nand NAND2 (N208, N175, N150);
nand NAND4 (N209, N198, N55, N120, N70);
or OR3 (N210, N206, N72, N168);
nor NOR2 (N211, N210, N77);
nor NOR3 (N212, N209, N101, N48);
not NOT1 (N213, N200);
nand NAND4 (N214, N194, N110, N178, N199);
nand NAND4 (N215, N207, N71, N207, N182);
buf BUF1 (N216, N145);
not NOT1 (N217, N211);
nor NOR3 (N218, N208, N60, N130);
or OR3 (N219, N215, N194, N101);
nor NOR3 (N220, N213, N198, N186);
nand NAND4 (N221, N212, N135, N80, N184);
and AND3 (N222, N221, N208, N210);
nand NAND2 (N223, N205, N215);
not NOT1 (N224, N220);
nor NOR3 (N225, N223, N149, N90);
xor XOR2 (N226, N188, N10);
nor NOR4 (N227, N226, N110, N90, N5);
nand NAND2 (N228, N218, N147);
not NOT1 (N229, N222);
buf BUF1 (N230, N228);
buf BUF1 (N231, N217);
or OR3 (N232, N230, N224, N60);
nand NAND3 (N233, N132, N5, N210);
buf BUF1 (N234, N232);
or OR4 (N235, N233, N73, N190, N165);
xor XOR2 (N236, N227, N234);
nand NAND3 (N237, N124, N165, N196);
not NOT1 (N238, N34);
nand NAND2 (N239, N238, N206);
or OR4 (N240, N239, N47, N106, N181);
and AND3 (N241, N214, N82, N178);
nor NOR2 (N242, N240, N73);
nor NOR2 (N243, N231, N65);
and AND3 (N244, N242, N205, N113);
or OR4 (N245, N229, N69, N21, N16);
xor XOR2 (N246, N244, N39);
xor XOR2 (N247, N216, N1);
and AND2 (N248, N236, N176);
nand NAND3 (N249, N248, N84, N231);
not NOT1 (N250, N249);
and AND4 (N251, N237, N40, N98, N215);
not NOT1 (N252, N235);
buf BUF1 (N253, N246);
or OR3 (N254, N253, N141, N107);
buf BUF1 (N255, N254);
buf BUF1 (N256, N252);
xor XOR2 (N257, N250, N109);
buf BUF1 (N258, N255);
buf BUF1 (N259, N241);
and AND4 (N260, N251, N185, N116, N167);
xor XOR2 (N261, N247, N106);
buf BUF1 (N262, N245);
nand NAND3 (N263, N256, N133, N131);
or OR4 (N264, N262, N211, N128, N235);
xor XOR2 (N265, N258, N87);
or OR4 (N266, N257, N158, N215, N30);
and AND3 (N267, N265, N72, N183);
or OR4 (N268, N219, N78, N38, N129);
buf BUF1 (N269, N261);
nor NOR2 (N270, N259, N60);
buf BUF1 (N271, N243);
nor NOR3 (N272, N269, N162, N119);
not NOT1 (N273, N225);
not NOT1 (N274, N271);
not NOT1 (N275, N272);
nand NAND2 (N276, N264, N250);
or OR4 (N277, N263, N239, N133, N51);
xor XOR2 (N278, N274, N222);
or OR2 (N279, N270, N199);
xor XOR2 (N280, N266, N68);
not NOT1 (N281, N278);
buf BUF1 (N282, N260);
or OR4 (N283, N280, N272, N208, N75);
nand NAND4 (N284, N282, N25, N46, N48);
nor NOR4 (N285, N284, N134, N283, N30);
and AND4 (N286, N66, N111, N244, N283);
nand NAND3 (N287, N277, N74, N107);
xor XOR2 (N288, N285, N189);
buf BUF1 (N289, N286);
buf BUF1 (N290, N267);
xor XOR2 (N291, N288, N121);
xor XOR2 (N292, N279, N136);
or OR3 (N293, N281, N154, N18);
xor XOR2 (N294, N293, N64);
nand NAND3 (N295, N294, N4, N46);
xor XOR2 (N296, N275, N176);
and AND3 (N297, N292, N79, N174);
xor XOR2 (N298, N296, N227);
nand NAND2 (N299, N268, N277);
nor NOR3 (N300, N295, N80, N206);
nand NAND3 (N301, N291, N28, N239);
nand NAND2 (N302, N301, N272);
xor XOR2 (N303, N273, N24);
or OR2 (N304, N276, N13);
not NOT1 (N305, N300);
not NOT1 (N306, N289);
and AND2 (N307, N303, N201);
nand NAND2 (N308, N297, N237);
buf BUF1 (N309, N290);
nor NOR4 (N310, N298, N18, N26, N301);
not NOT1 (N311, N310);
not NOT1 (N312, N299);
or OR3 (N313, N308, N178, N23);
not NOT1 (N314, N302);
buf BUF1 (N315, N313);
nand NAND3 (N316, N305, N73, N31);
or OR3 (N317, N315, N99, N147);
or OR4 (N318, N304, N45, N152, N196);
and AND3 (N319, N316, N244, N225);
not NOT1 (N320, N311);
not NOT1 (N321, N312);
and AND3 (N322, N287, N180, N264);
and AND4 (N323, N321, N35, N149, N297);
and AND2 (N324, N320, N251);
buf BUF1 (N325, N317);
buf BUF1 (N326, N325);
xor XOR2 (N327, N307, N126);
buf BUF1 (N328, N327);
not NOT1 (N329, N306);
not NOT1 (N330, N328);
and AND4 (N331, N319, N49, N152, N106);
buf BUF1 (N332, N314);
and AND4 (N333, N326, N210, N47, N209);
not NOT1 (N334, N329);
nand NAND2 (N335, N333, N9);
nor NOR3 (N336, N334, N65, N253);
buf BUF1 (N337, N336);
buf BUF1 (N338, N309);
and AND2 (N339, N335, N261);
nand NAND3 (N340, N323, N78, N94);
not NOT1 (N341, N337);
xor XOR2 (N342, N341, N230);
or OR2 (N343, N322, N14);
not NOT1 (N344, N342);
and AND3 (N345, N318, N301, N41);
buf BUF1 (N346, N324);
and AND2 (N347, N346, N301);
buf BUF1 (N348, N338);
not NOT1 (N349, N339);
buf BUF1 (N350, N347);
nand NAND2 (N351, N332, N319);
buf BUF1 (N352, N348);
buf BUF1 (N353, N331);
xor XOR2 (N354, N353, N90);
not NOT1 (N355, N349);
or OR4 (N356, N351, N353, N15, N226);
nand NAND3 (N357, N345, N74, N266);
nand NAND2 (N358, N344, N141);
buf BUF1 (N359, N354);
and AND3 (N360, N343, N69, N12);
nor NOR3 (N361, N355, N8, N114);
nor NOR2 (N362, N358, N226);
not NOT1 (N363, N361);
or OR3 (N364, N362, N267, N186);
not NOT1 (N365, N363);
nand NAND3 (N366, N359, N265, N84);
and AND4 (N367, N340, N299, N71, N38);
xor XOR2 (N368, N330, N238);
and AND3 (N369, N352, N250, N127);
xor XOR2 (N370, N365, N247);
not NOT1 (N371, N360);
buf BUF1 (N372, N357);
buf BUF1 (N373, N356);
not NOT1 (N374, N370);
buf BUF1 (N375, N367);
and AND2 (N376, N373, N225);
xor XOR2 (N377, N368, N121);
or OR4 (N378, N366, N46, N132, N151);
or OR2 (N379, N350, N80);
or OR3 (N380, N375, N150, N59);
and AND2 (N381, N377, N358);
xor XOR2 (N382, N369, N318);
nor NOR3 (N383, N382, N219, N233);
and AND4 (N384, N372, N88, N329, N205);
nor NOR4 (N385, N378, N351, N380, N376);
nor NOR2 (N386, N314, N153);
buf BUF1 (N387, N264);
nand NAND3 (N388, N386, N64, N385);
nand NAND2 (N389, N247, N17);
or OR4 (N390, N383, N113, N236, N157);
buf BUF1 (N391, N390);
and AND3 (N392, N389, N358, N346);
and AND2 (N393, N371, N225);
not NOT1 (N394, N379);
xor XOR2 (N395, N364, N289);
nand NAND2 (N396, N374, N271);
xor XOR2 (N397, N396, N202);
or OR4 (N398, N381, N189, N53, N91);
not NOT1 (N399, N394);
buf BUF1 (N400, N387);
not NOT1 (N401, N397);
not NOT1 (N402, N401);
nor NOR2 (N403, N391, N329);
buf BUF1 (N404, N384);
or OR3 (N405, N388, N66, N308);
buf BUF1 (N406, N399);
and AND2 (N407, N405, N150);
nand NAND4 (N408, N398, N158, N370, N46);
xor XOR2 (N409, N406, N362);
xor XOR2 (N410, N404, N380);
not NOT1 (N411, N403);
nand NAND4 (N412, N392, N18, N109, N103);
or OR3 (N413, N410, N30, N107);
and AND3 (N414, N409, N309, N94);
nor NOR2 (N415, N412, N104);
nand NAND2 (N416, N395, N88);
or OR3 (N417, N415, N164, N122);
and AND2 (N418, N393, N275);
or OR4 (N419, N400, N50, N361, N136);
buf BUF1 (N420, N417);
nor NOR3 (N421, N418, N303, N388);
or OR4 (N422, N402, N161, N352, N307);
or OR4 (N423, N419, N282, N86, N104);
nor NOR2 (N424, N408, N396);
nand NAND4 (N425, N422, N335, N297, N222);
or OR2 (N426, N425, N132);
and AND4 (N427, N426, N233, N310, N26);
not NOT1 (N428, N421);
or OR4 (N429, N427, N301, N177, N410);
nor NOR4 (N430, N411, N366, N160, N96);
or OR2 (N431, N413, N84);
and AND2 (N432, N431, N286);
not NOT1 (N433, N414);
and AND4 (N434, N433, N299, N37, N193);
nand NAND3 (N435, N429, N399, N292);
not NOT1 (N436, N435);
xor XOR2 (N437, N432, N414);
nand NAND4 (N438, N436, N175, N339, N268);
and AND2 (N439, N407, N161);
nor NOR2 (N440, N416, N50);
and AND3 (N441, N434, N224, N397);
nand NAND3 (N442, N438, N382, N219);
xor XOR2 (N443, N430, N98);
and AND2 (N444, N442, N314);
not NOT1 (N445, N444);
nand NAND4 (N446, N443, N288, N285, N336);
nor NOR4 (N447, N423, N250, N305, N168);
buf BUF1 (N448, N447);
or OR4 (N449, N420, N385, N248, N356);
nor NOR2 (N450, N441, N9);
buf BUF1 (N451, N448);
nand NAND2 (N452, N446, N83);
not NOT1 (N453, N424);
or OR3 (N454, N452, N276, N108);
not NOT1 (N455, N451);
not NOT1 (N456, N437);
not NOT1 (N457, N440);
nand NAND4 (N458, N455, N336, N257, N322);
buf BUF1 (N459, N449);
or OR2 (N460, N454, N272);
xor XOR2 (N461, N439, N229);
or OR2 (N462, N459, N434);
buf BUF1 (N463, N450);
buf BUF1 (N464, N461);
nor NOR3 (N465, N456, N107, N270);
and AND2 (N466, N465, N111);
buf BUF1 (N467, N457);
or OR4 (N468, N463, N174, N56, N266);
buf BUF1 (N469, N458);
or OR3 (N470, N462, N243, N317);
xor XOR2 (N471, N428, N305);
or OR2 (N472, N460, N169);
xor XOR2 (N473, N471, N132);
nand NAND2 (N474, N464, N459);
and AND4 (N475, N468, N410, N257, N103);
nand NAND3 (N476, N469, N221, N210);
nand NAND2 (N477, N467, N414);
and AND3 (N478, N475, N434, N226);
not NOT1 (N479, N477);
and AND3 (N480, N470, N429, N156);
or OR2 (N481, N480, N97);
nand NAND4 (N482, N472, N194, N37, N456);
nand NAND2 (N483, N478, N185);
nor NOR3 (N484, N483, N4, N212);
nand NAND4 (N485, N466, N393, N9, N46);
buf BUF1 (N486, N482);
or OR3 (N487, N473, N418, N399);
not NOT1 (N488, N474);
buf BUF1 (N489, N484);
nand NAND2 (N490, N453, N388);
buf BUF1 (N491, N445);
and AND3 (N492, N486, N226, N478);
not NOT1 (N493, N488);
or OR4 (N494, N481, N248, N158, N143);
nor NOR3 (N495, N479, N206, N158);
nor NOR3 (N496, N487, N86, N438);
nand NAND3 (N497, N495, N397, N69);
nand NAND2 (N498, N476, N346);
xor XOR2 (N499, N493, N17);
nand NAND4 (N500, N491, N45, N187, N251);
xor XOR2 (N501, N494, N241);
or OR2 (N502, N500, N70);
buf BUF1 (N503, N490);
xor XOR2 (N504, N485, N389);
or OR3 (N505, N496, N109, N138);
buf BUF1 (N506, N502);
xor XOR2 (N507, N506, N233);
nor NOR4 (N508, N492, N96, N395, N356);
nor NOR4 (N509, N504, N441, N389, N174);
nor NOR2 (N510, N509, N500);
not NOT1 (N511, N497);
buf BUF1 (N512, N505);
xor XOR2 (N513, N510, N348);
nand NAND2 (N514, N507, N194);
or OR2 (N515, N503, N301);
or OR4 (N516, N513, N385, N491, N442);
nor NOR2 (N517, N498, N286);
xor XOR2 (N518, N501, N226);
buf BUF1 (N519, N516);
or OR3 (N520, N517, N179, N36);
nor NOR4 (N521, N512, N383, N114, N228);
nand NAND3 (N522, N519, N115, N60);
nand NAND3 (N523, N521, N385, N5);
nor NOR4 (N524, N518, N57, N134, N177);
and AND4 (N525, N499, N466, N504, N190);
nand NAND2 (N526, N525, N75);
and AND3 (N527, N489, N272, N141);
and AND3 (N528, N515, N414, N214);
and AND3 (N529, N523, N447, N40);
xor XOR2 (N530, N528, N409);
or OR4 (N531, N529, N154, N303, N381);
not NOT1 (N532, N514);
and AND3 (N533, N522, N244, N373);
nor NOR3 (N534, N532, N266, N102);
xor XOR2 (N535, N524, N9);
nand NAND4 (N536, N531, N166, N311, N159);
nand NAND2 (N537, N533, N90);
not NOT1 (N538, N536);
not NOT1 (N539, N537);
buf BUF1 (N540, N535);
or OR4 (N541, N539, N129, N501, N213);
not NOT1 (N542, N538);
and AND4 (N543, N511, N460, N311, N456);
or OR2 (N544, N541, N233);
nand NAND4 (N545, N527, N29, N364, N102);
nor NOR4 (N546, N520, N147, N225, N459);
nor NOR3 (N547, N545, N460, N302);
not NOT1 (N548, N542);
or OR4 (N549, N544, N258, N22, N510);
xor XOR2 (N550, N548, N226);
and AND3 (N551, N540, N218, N344);
xor XOR2 (N552, N547, N247);
not NOT1 (N553, N552);
and AND3 (N554, N508, N502, N314);
buf BUF1 (N555, N526);
nor NOR3 (N556, N549, N197, N400);
or OR2 (N557, N530, N444);
xor XOR2 (N558, N553, N190);
nor NOR3 (N559, N546, N419, N434);
xor XOR2 (N560, N558, N240);
nor NOR4 (N561, N554, N401, N90, N288);
not NOT1 (N562, N559);
or OR3 (N563, N560, N123, N40);
not NOT1 (N564, N561);
and AND4 (N565, N534, N142, N298, N282);
and AND2 (N566, N555, N200);
nor NOR2 (N567, N563, N460);
and AND2 (N568, N565, N8);
or OR3 (N569, N543, N415, N34);
and AND4 (N570, N551, N27, N439, N247);
nand NAND4 (N571, N556, N152, N241, N4);
nor NOR4 (N572, N569, N197, N225, N256);
and AND4 (N573, N562, N218, N321, N346);
nand NAND4 (N574, N567, N343, N133, N138);
and AND2 (N575, N568, N543);
nor NOR4 (N576, N566, N423, N395, N224);
not NOT1 (N577, N571);
buf BUF1 (N578, N576);
nor NOR4 (N579, N550, N300, N166, N31);
xor XOR2 (N580, N579, N177);
not NOT1 (N581, N574);
and AND2 (N582, N557, N296);
xor XOR2 (N583, N564, N485);
and AND4 (N584, N577, N381, N182, N380);
or OR3 (N585, N573, N73, N246);
buf BUF1 (N586, N583);
not NOT1 (N587, N581);
nor NOR3 (N588, N570, N530, N155);
nand NAND3 (N589, N572, N578, N53);
xor XOR2 (N590, N139, N252);
xor XOR2 (N591, N586, N92);
or OR4 (N592, N582, N134, N169, N483);
nand NAND4 (N593, N580, N347, N578, N169);
buf BUF1 (N594, N585);
or OR2 (N595, N590, N555);
nor NOR2 (N596, N584, N251);
xor XOR2 (N597, N587, N438);
or OR3 (N598, N588, N189, N500);
nand NAND3 (N599, N598, N120, N534);
nand NAND4 (N600, N594, N59, N58, N255);
and AND4 (N601, N595, N85, N170, N332);
not NOT1 (N602, N575);
xor XOR2 (N603, N591, N153);
not NOT1 (N604, N592);
or OR2 (N605, N603, N502);
buf BUF1 (N606, N599);
nor NOR3 (N607, N602, N569, N243);
or OR2 (N608, N600, N324);
xor XOR2 (N609, N608, N75);
nor NOR4 (N610, N589, N331, N341, N26);
nand NAND3 (N611, N597, N325, N22);
xor XOR2 (N612, N609, N141);
xor XOR2 (N613, N612, N439);
or OR4 (N614, N601, N423, N598, N200);
or OR4 (N615, N593, N399, N413, N48);
nor NOR4 (N616, N606, N229, N331, N221);
or OR4 (N617, N610, N564, N446, N598);
or OR3 (N618, N596, N507, N602);
and AND2 (N619, N611, N574);
xor XOR2 (N620, N618, N504);
buf BUF1 (N621, N616);
xor XOR2 (N622, N619, N103);
xor XOR2 (N623, N622, N216);
xor XOR2 (N624, N617, N169);
nand NAND2 (N625, N621, N533);
buf BUF1 (N626, N607);
not NOT1 (N627, N604);
xor XOR2 (N628, N627, N383);
buf BUF1 (N629, N620);
nor NOR4 (N630, N615, N576, N466, N354);
or OR4 (N631, N625, N572, N270, N149);
nand NAND2 (N632, N605, N298);
buf BUF1 (N633, N624);
buf BUF1 (N634, N613);
or OR2 (N635, N634, N586);
and AND3 (N636, N630, N407, N379);
not NOT1 (N637, N626);
not NOT1 (N638, N637);
not NOT1 (N639, N633);
nor NOR4 (N640, N638, N401, N448, N223);
not NOT1 (N641, N628);
buf BUF1 (N642, N614);
nor NOR3 (N643, N641, N152, N157);
nand NAND2 (N644, N623, N117);
not NOT1 (N645, N642);
or OR4 (N646, N631, N527, N289, N413);
and AND3 (N647, N639, N644, N269);
not NOT1 (N648, N57);
and AND3 (N649, N643, N346, N620);
and AND3 (N650, N649, N586, N50);
nand NAND4 (N651, N648, N72, N116, N237);
and AND4 (N652, N632, N621, N263, N334);
nor NOR2 (N653, N635, N86);
buf BUF1 (N654, N651);
nand NAND3 (N655, N650, N300, N570);
or OR3 (N656, N654, N377, N294);
xor XOR2 (N657, N640, N333);
or OR4 (N658, N652, N369, N268, N279);
nand NAND3 (N659, N657, N589, N66);
and AND2 (N660, N656, N141);
buf BUF1 (N661, N629);
not NOT1 (N662, N653);
xor XOR2 (N663, N662, N351);
xor XOR2 (N664, N645, N251);
nor NOR4 (N665, N659, N401, N100, N104);
nor NOR3 (N666, N665, N456, N26);
buf BUF1 (N667, N646);
or OR3 (N668, N660, N241, N362);
and AND3 (N669, N661, N97, N503);
and AND2 (N670, N636, N158);
and AND4 (N671, N666, N24, N455, N549);
and AND4 (N672, N670, N595, N300, N45);
and AND4 (N673, N672, N36, N228, N240);
and AND3 (N674, N663, N338, N52);
nor NOR3 (N675, N667, N392, N382);
or OR3 (N676, N674, N305, N573);
not NOT1 (N677, N647);
not NOT1 (N678, N655);
xor XOR2 (N679, N664, N539);
not NOT1 (N680, N668);
xor XOR2 (N681, N680, N376);
or OR3 (N682, N675, N564, N125);
not NOT1 (N683, N681);
not NOT1 (N684, N677);
or OR4 (N685, N669, N378, N557, N377);
or OR2 (N686, N679, N66);
xor XOR2 (N687, N673, N462);
nand NAND3 (N688, N686, N172, N505);
and AND4 (N689, N678, N278, N48, N640);
not NOT1 (N690, N689);
nor NOR3 (N691, N685, N61, N498);
and AND3 (N692, N658, N189, N306);
nand NAND4 (N693, N671, N13, N441, N648);
not NOT1 (N694, N691);
and AND3 (N695, N688, N466, N90);
and AND3 (N696, N692, N398, N468);
xor XOR2 (N697, N684, N513);
nand NAND2 (N698, N695, N567);
buf BUF1 (N699, N683);
nand NAND2 (N700, N682, N545);
xor XOR2 (N701, N697, N558);
buf BUF1 (N702, N696);
buf BUF1 (N703, N690);
nand NAND2 (N704, N701, N328);
nand NAND4 (N705, N700, N203, N675, N297);
buf BUF1 (N706, N694);
buf BUF1 (N707, N706);
nand NAND3 (N708, N699, N175, N410);
or OR3 (N709, N703, N684, N403);
nand NAND3 (N710, N705, N248, N501);
buf BUF1 (N711, N710);
buf BUF1 (N712, N687);
not NOT1 (N713, N704);
nand NAND3 (N714, N708, N191, N491);
buf BUF1 (N715, N676);
nand NAND3 (N716, N711, N290, N624);
buf BUF1 (N717, N693);
nor NOR2 (N718, N709, N535);
buf BUF1 (N719, N712);
nand NAND4 (N720, N707, N1, N449, N622);
and AND4 (N721, N717, N436, N304, N196);
nand NAND2 (N722, N718, N649);
not NOT1 (N723, N702);
xor XOR2 (N724, N698, N92);
not NOT1 (N725, N714);
nand NAND2 (N726, N721, N670);
or OR2 (N727, N726, N23);
nand NAND2 (N728, N720, N609);
nor NOR4 (N729, N723, N566, N433, N694);
not NOT1 (N730, N728);
and AND2 (N731, N727, N180);
xor XOR2 (N732, N715, N547);
nor NOR3 (N733, N713, N322, N359);
buf BUF1 (N734, N733);
or OR2 (N735, N729, N588);
nor NOR3 (N736, N734, N159, N277);
nand NAND4 (N737, N735, N500, N705, N630);
or OR3 (N738, N724, N135, N452);
nor NOR2 (N739, N725, N119);
not NOT1 (N740, N730);
xor XOR2 (N741, N722, N562);
nand NAND3 (N742, N732, N63, N508);
nand NAND4 (N743, N719, N209, N455, N261);
and AND4 (N744, N738, N511, N375, N384);
and AND2 (N745, N740, N635);
or OR2 (N746, N716, N516);
nand NAND2 (N747, N743, N717);
and AND2 (N748, N739, N624);
nand NAND2 (N749, N745, N701);
not NOT1 (N750, N749);
or OR2 (N751, N747, N57);
or OR3 (N752, N731, N42, N607);
buf BUF1 (N753, N748);
nor NOR4 (N754, N744, N381, N629, N77);
xor XOR2 (N755, N754, N388);
not NOT1 (N756, N752);
or OR3 (N757, N741, N428, N55);
and AND3 (N758, N755, N365, N581);
and AND4 (N759, N757, N82, N388, N76);
nand NAND3 (N760, N751, N354, N367);
xor XOR2 (N761, N746, N621);
xor XOR2 (N762, N756, N371);
or OR4 (N763, N750, N421, N619, N471);
nand NAND4 (N764, N761, N536, N605, N706);
not NOT1 (N765, N764);
and AND3 (N766, N765, N145, N642);
buf BUF1 (N767, N760);
nand NAND2 (N768, N758, N154);
nor NOR2 (N769, N768, N737);
xor XOR2 (N770, N661, N120);
not NOT1 (N771, N753);
nor NOR2 (N772, N736, N552);
nand NAND4 (N773, N767, N387, N230, N650);
and AND4 (N774, N762, N419, N685, N191);
or OR4 (N775, N769, N319, N93, N583);
buf BUF1 (N776, N773);
xor XOR2 (N777, N759, N127);
nand NAND2 (N778, N775, N600);
and AND3 (N779, N770, N369, N519);
buf BUF1 (N780, N778);
buf BUF1 (N781, N774);
nor NOR4 (N782, N776, N134, N736, N394);
not NOT1 (N783, N781);
buf BUF1 (N784, N782);
buf BUF1 (N785, N784);
buf BUF1 (N786, N766);
and AND3 (N787, N786, N298, N318);
nor NOR2 (N788, N772, N347);
and AND4 (N789, N777, N702, N60, N174);
nor NOR4 (N790, N763, N379, N400, N16);
not NOT1 (N791, N779);
or OR2 (N792, N791, N9);
not NOT1 (N793, N790);
buf BUF1 (N794, N785);
and AND3 (N795, N792, N2, N719);
buf BUF1 (N796, N795);
not NOT1 (N797, N789);
nand NAND3 (N798, N796, N517, N699);
not NOT1 (N799, N742);
buf BUF1 (N800, N771);
buf BUF1 (N801, N780);
or OR2 (N802, N797, N492);
nand NAND2 (N803, N800, N696);
nor NOR2 (N804, N803, N558);
nand NAND2 (N805, N793, N550);
nor NOR2 (N806, N788, N467);
xor XOR2 (N807, N801, N57);
nand NAND2 (N808, N805, N503);
nand NAND4 (N809, N806, N498, N174, N707);
not NOT1 (N810, N807);
or OR4 (N811, N809, N83, N445, N226);
nand NAND4 (N812, N794, N272, N140, N717);
xor XOR2 (N813, N802, N39);
xor XOR2 (N814, N787, N26);
not NOT1 (N815, N813);
and AND2 (N816, N814, N108);
and AND2 (N817, N815, N793);
not NOT1 (N818, N804);
nor NOR2 (N819, N818, N391);
and AND2 (N820, N817, N527);
nor NOR2 (N821, N783, N347);
buf BUF1 (N822, N798);
or OR4 (N823, N810, N678, N697, N288);
xor XOR2 (N824, N799, N285);
nand NAND2 (N825, N816, N785);
nor NOR3 (N826, N823, N410, N620);
or OR3 (N827, N812, N691, N207);
nand NAND2 (N828, N811, N91);
nand NAND3 (N829, N808, N94, N10);
buf BUF1 (N830, N824);
or OR4 (N831, N821, N500, N480, N517);
buf BUF1 (N832, N828);
nand NAND2 (N833, N820, N572);
and AND3 (N834, N832, N163, N96);
and AND3 (N835, N833, N441, N733);
not NOT1 (N836, N834);
not NOT1 (N837, N830);
nor NOR3 (N838, N827, N404, N678);
buf BUF1 (N839, N829);
nor NOR3 (N840, N825, N99, N114);
or OR2 (N841, N826, N421);
and AND3 (N842, N822, N524, N558);
nor NOR4 (N843, N841, N550, N689, N528);
buf BUF1 (N844, N819);
nand NAND2 (N845, N837, N502);
not NOT1 (N846, N845);
and AND2 (N847, N840, N613);
and AND4 (N848, N847, N284, N265, N447);
and AND2 (N849, N846, N765);
xor XOR2 (N850, N842, N835);
and AND3 (N851, N489, N739, N11);
or OR2 (N852, N848, N799);
nor NOR4 (N853, N843, N105, N604, N51);
and AND3 (N854, N851, N272, N460);
nand NAND3 (N855, N853, N747, N175);
not NOT1 (N856, N839);
not NOT1 (N857, N855);
nand NAND4 (N858, N849, N249, N113, N721);
buf BUF1 (N859, N858);
not NOT1 (N860, N850);
xor XOR2 (N861, N838, N592);
xor XOR2 (N862, N831, N102);
and AND3 (N863, N861, N186, N482);
nor NOR3 (N864, N862, N225, N593);
buf BUF1 (N865, N859);
xor XOR2 (N866, N856, N436);
xor XOR2 (N867, N852, N455);
xor XOR2 (N868, N866, N800);
not NOT1 (N869, N844);
xor XOR2 (N870, N867, N208);
and AND2 (N871, N863, N348);
or OR2 (N872, N869, N363);
and AND4 (N873, N872, N848, N148, N828);
not NOT1 (N874, N871);
buf BUF1 (N875, N870);
xor XOR2 (N876, N873, N836);
not NOT1 (N877, N760);
buf BUF1 (N878, N864);
buf BUF1 (N879, N865);
nor NOR2 (N880, N877, N325);
nand NAND2 (N881, N878, N636);
nor NOR2 (N882, N860, N130);
nor NOR3 (N883, N868, N224, N763);
and AND3 (N884, N879, N409, N435);
nand NAND4 (N885, N883, N790, N423, N631);
nor NOR4 (N886, N874, N582, N522, N409);
nand NAND3 (N887, N880, N100, N481);
xor XOR2 (N888, N881, N399);
or OR3 (N889, N886, N168, N720);
nor NOR2 (N890, N885, N733);
or OR3 (N891, N854, N435, N862);
or OR4 (N892, N887, N850, N737, N340);
nor NOR4 (N893, N875, N655, N694, N696);
buf BUF1 (N894, N888);
not NOT1 (N895, N857);
or OR2 (N896, N884, N568);
buf BUF1 (N897, N893);
buf BUF1 (N898, N890);
xor XOR2 (N899, N895, N21);
or OR3 (N900, N892, N720, N85);
buf BUF1 (N901, N876);
xor XOR2 (N902, N900, N97);
not NOT1 (N903, N891);
nor NOR2 (N904, N897, N209);
nand NAND4 (N905, N901, N160, N512, N344);
and AND2 (N906, N896, N227);
buf BUF1 (N907, N905);
nor NOR3 (N908, N889, N322, N567);
xor XOR2 (N909, N898, N758);
nand NAND4 (N910, N906, N79, N259, N243);
or OR4 (N911, N908, N392, N222, N795);
and AND2 (N912, N894, N90);
nand NAND3 (N913, N907, N192, N373);
or OR4 (N914, N903, N438, N819, N224);
and AND2 (N915, N882, N734);
nand NAND4 (N916, N902, N331, N865, N577);
xor XOR2 (N917, N914, N870);
and AND3 (N918, N912, N588, N623);
nand NAND3 (N919, N918, N512, N563);
not NOT1 (N920, N916);
buf BUF1 (N921, N911);
buf BUF1 (N922, N919);
buf BUF1 (N923, N920);
nand NAND4 (N924, N915, N873, N431, N131);
nor NOR3 (N925, N923, N108, N180);
and AND2 (N926, N917, N796);
or OR4 (N927, N926, N859, N659, N149);
xor XOR2 (N928, N904, N143);
and AND3 (N929, N913, N529, N756);
not NOT1 (N930, N929);
nand NAND3 (N931, N922, N930, N212);
nand NAND3 (N932, N782, N767, N900);
buf BUF1 (N933, N931);
and AND4 (N934, N910, N3, N746, N390);
xor XOR2 (N935, N909, N501);
buf BUF1 (N936, N899);
or OR2 (N937, N928, N244);
xor XOR2 (N938, N934, N147);
xor XOR2 (N939, N932, N204);
nor NOR2 (N940, N921, N472);
and AND2 (N941, N938, N625);
xor XOR2 (N942, N940, N486);
not NOT1 (N943, N935);
xor XOR2 (N944, N942, N782);
and AND3 (N945, N941, N420, N173);
not NOT1 (N946, N937);
or OR4 (N947, N945, N14, N226, N457);
not NOT1 (N948, N947);
buf BUF1 (N949, N939);
not NOT1 (N950, N943);
and AND2 (N951, N948, N355);
and AND4 (N952, N924, N609, N252, N621);
not NOT1 (N953, N946);
nand NAND2 (N954, N944, N943);
or OR4 (N955, N953, N61, N63, N726);
nor NOR4 (N956, N955, N476, N669, N576);
or OR4 (N957, N951, N264, N563, N191);
xor XOR2 (N958, N950, N688);
and AND4 (N959, N925, N354, N258, N23);
nand NAND4 (N960, N959, N516, N101, N293);
nor NOR4 (N961, N952, N866, N106, N598);
xor XOR2 (N962, N954, N182);
nor NOR4 (N963, N962, N492, N928, N404);
and AND2 (N964, N961, N328);
and AND2 (N965, N964, N803);
xor XOR2 (N966, N933, N594);
buf BUF1 (N967, N927);
nor NOR2 (N968, N958, N728);
not NOT1 (N969, N936);
not NOT1 (N970, N957);
xor XOR2 (N971, N968, N770);
or OR4 (N972, N970, N660, N479, N64);
xor XOR2 (N973, N963, N812);
and AND4 (N974, N966, N419, N238, N21);
not NOT1 (N975, N960);
buf BUF1 (N976, N956);
nor NOR3 (N977, N974, N919, N749);
buf BUF1 (N978, N967);
or OR2 (N979, N972, N67);
not NOT1 (N980, N975);
xor XOR2 (N981, N965, N47);
buf BUF1 (N982, N969);
not NOT1 (N983, N982);
nand NAND4 (N984, N983, N192, N595, N679);
buf BUF1 (N985, N981);
not NOT1 (N986, N985);
buf BUF1 (N987, N949);
buf BUF1 (N988, N980);
or OR4 (N989, N977, N75, N306, N395);
nor NOR3 (N990, N986, N738, N236);
or OR2 (N991, N973, N451);
nor NOR3 (N992, N990, N769, N284);
not NOT1 (N993, N979);
and AND4 (N994, N988, N856, N158, N483);
nand NAND4 (N995, N993, N748, N614, N692);
nor NOR3 (N996, N971, N202, N86);
buf BUF1 (N997, N976);
or OR3 (N998, N978, N616, N624);
and AND4 (N999, N994, N506, N492, N525);
xor XOR2 (N1000, N996, N702);
nand NAND4 (N1001, N992, N190, N921, N982);
nor NOR4 (N1002, N995, N305, N543, N767);
nor NOR2 (N1003, N1000, N913);
xor XOR2 (N1004, N987, N645);
and AND3 (N1005, N997, N980, N594);
nand NAND3 (N1006, N991, N452, N268);
xor XOR2 (N1007, N1004, N706);
nand NAND3 (N1008, N1005, N67, N223);
nor NOR3 (N1009, N1008, N446, N632);
nand NAND2 (N1010, N999, N408);
or OR2 (N1011, N998, N23);
nor NOR3 (N1012, N1010, N851, N323);
buf BUF1 (N1013, N1009);
xor XOR2 (N1014, N1003, N175);
buf BUF1 (N1015, N984);
not NOT1 (N1016, N1006);
xor XOR2 (N1017, N1014, N289);
or OR4 (N1018, N1017, N742, N734, N170);
or OR3 (N1019, N1007, N1003, N323);
nor NOR4 (N1020, N1016, N132, N194, N78);
xor XOR2 (N1021, N1019, N496);
nand NAND3 (N1022, N1013, N527, N661);
not NOT1 (N1023, N1001);
nor NOR2 (N1024, N1015, N240);
xor XOR2 (N1025, N1020, N159);
or OR2 (N1026, N1024, N838);
xor XOR2 (N1027, N1026, N935);
nand NAND2 (N1028, N1023, N690);
or OR4 (N1029, N1028, N953, N403, N424);
nor NOR3 (N1030, N1002, N639, N763);
not NOT1 (N1031, N989);
or OR4 (N1032, N1022, N776, N61, N196);
not NOT1 (N1033, N1018);
not NOT1 (N1034, N1012);
nor NOR2 (N1035, N1030, N923);
not NOT1 (N1036, N1027);
xor XOR2 (N1037, N1029, N938);
or OR4 (N1038, N1033, N1033, N118, N637);
nor NOR3 (N1039, N1011, N963, N405);
nor NOR3 (N1040, N1032, N114, N774);
buf BUF1 (N1041, N1035);
not NOT1 (N1042, N1040);
nor NOR3 (N1043, N1021, N297, N824);
not NOT1 (N1044, N1037);
nor NOR3 (N1045, N1036, N346, N420);
nor NOR2 (N1046, N1044, N643);
nand NAND2 (N1047, N1031, N32);
or OR2 (N1048, N1041, N598);
nor NOR3 (N1049, N1045, N276, N432);
not NOT1 (N1050, N1039);
xor XOR2 (N1051, N1038, N780);
buf BUF1 (N1052, N1051);
not NOT1 (N1053, N1034);
nand NAND2 (N1054, N1050, N509);
nor NOR2 (N1055, N1054, N236);
xor XOR2 (N1056, N1055, N389);
xor XOR2 (N1057, N1046, N298);
buf BUF1 (N1058, N1047);
and AND3 (N1059, N1057, N427, N60);
xor XOR2 (N1060, N1042, N584);
buf BUF1 (N1061, N1056);
or OR2 (N1062, N1043, N108);
buf BUF1 (N1063, N1049);
nor NOR3 (N1064, N1061, N56, N493);
and AND3 (N1065, N1064, N178, N159);
xor XOR2 (N1066, N1065, N561);
nand NAND2 (N1067, N1025, N742);
xor XOR2 (N1068, N1063, N956);
and AND2 (N1069, N1068, N438);
or OR4 (N1070, N1058, N90, N837, N127);
xor XOR2 (N1071, N1067, N861);
nand NAND3 (N1072, N1053, N412, N847);
or OR3 (N1073, N1071, N196, N57);
or OR4 (N1074, N1070, N317, N742, N897);
not NOT1 (N1075, N1069);
xor XOR2 (N1076, N1048, N1008);
xor XOR2 (N1077, N1060, N865);
and AND4 (N1078, N1076, N78, N1063, N592);
not NOT1 (N1079, N1075);
not NOT1 (N1080, N1072);
xor XOR2 (N1081, N1079, N166);
nor NOR4 (N1082, N1080, N671, N986, N966);
nor NOR2 (N1083, N1059, N696);
or OR2 (N1084, N1052, N988);
buf BUF1 (N1085, N1062);
or OR3 (N1086, N1081, N803, N171);
xor XOR2 (N1087, N1085, N660);
nand NAND2 (N1088, N1073, N241);
nand NAND3 (N1089, N1088, N720, N798);
or OR4 (N1090, N1084, N893, N1033, N327);
nand NAND4 (N1091, N1077, N98, N725, N47);
or OR2 (N1092, N1083, N779);
or OR3 (N1093, N1092, N260, N305);
or OR4 (N1094, N1090, N595, N74, N129);
buf BUF1 (N1095, N1087);
or OR2 (N1096, N1091, N111);
nor NOR3 (N1097, N1093, N352, N350);
not NOT1 (N1098, N1096);
buf BUF1 (N1099, N1095);
or OR2 (N1100, N1086, N941);
nand NAND2 (N1101, N1094, N899);
xor XOR2 (N1102, N1099, N59);
and AND4 (N1103, N1101, N424, N483, N485);
nand NAND3 (N1104, N1078, N556, N102);
and AND2 (N1105, N1089, N141);
or OR3 (N1106, N1100, N229, N879);
xor XOR2 (N1107, N1097, N1104);
xor XOR2 (N1108, N184, N967);
not NOT1 (N1109, N1102);
nor NOR2 (N1110, N1074, N262);
or OR4 (N1111, N1098, N496, N1072, N1080);
xor XOR2 (N1112, N1066, N738);
xor XOR2 (N1113, N1110, N319);
buf BUF1 (N1114, N1107);
nand NAND2 (N1115, N1108, N148);
nor NOR2 (N1116, N1106, N921);
xor XOR2 (N1117, N1111, N324);
and AND4 (N1118, N1116, N863, N905, N368);
not NOT1 (N1119, N1114);
xor XOR2 (N1120, N1113, N978);
nor NOR2 (N1121, N1118, N6);
nand NAND3 (N1122, N1115, N169, N1062);
not NOT1 (N1123, N1117);
nor NOR3 (N1124, N1123, N943, N275);
or OR4 (N1125, N1122, N748, N341, N483);
nand NAND2 (N1126, N1105, N714);
buf BUF1 (N1127, N1125);
buf BUF1 (N1128, N1124);
xor XOR2 (N1129, N1109, N324);
or OR3 (N1130, N1082, N87, N678);
nor NOR2 (N1131, N1121, N403);
not NOT1 (N1132, N1120);
and AND2 (N1133, N1128, N705);
nor NOR4 (N1134, N1119, N454, N878, N75);
and AND2 (N1135, N1129, N599);
and AND2 (N1136, N1131, N280);
nand NAND3 (N1137, N1130, N414, N231);
xor XOR2 (N1138, N1137, N1122);
buf BUF1 (N1139, N1126);
buf BUF1 (N1140, N1133);
not NOT1 (N1141, N1138);
buf BUF1 (N1142, N1127);
xor XOR2 (N1143, N1135, N610);
nand NAND4 (N1144, N1112, N265, N618, N315);
nor NOR2 (N1145, N1139, N247);
buf BUF1 (N1146, N1140);
and AND2 (N1147, N1144, N964);
not NOT1 (N1148, N1132);
xor XOR2 (N1149, N1143, N742);
nand NAND2 (N1150, N1141, N108);
or OR4 (N1151, N1142, N961, N162, N708);
nand NAND3 (N1152, N1149, N1095, N321);
xor XOR2 (N1153, N1150, N1108);
nor NOR4 (N1154, N1153, N582, N584, N870);
or OR2 (N1155, N1148, N48);
not NOT1 (N1156, N1155);
or OR4 (N1157, N1147, N63, N185, N639);
nand NAND3 (N1158, N1136, N635, N188);
buf BUF1 (N1159, N1158);
buf BUF1 (N1160, N1145);
nor NOR2 (N1161, N1146, N1014);
xor XOR2 (N1162, N1157, N1099);
and AND2 (N1163, N1151, N411);
xor XOR2 (N1164, N1156, N949);
and AND2 (N1165, N1163, N713);
not NOT1 (N1166, N1154);
xor XOR2 (N1167, N1164, N939);
nor NOR4 (N1168, N1165, N697, N651, N105);
nor NOR2 (N1169, N1161, N1129);
nand NAND3 (N1170, N1168, N582, N257);
xor XOR2 (N1171, N1159, N657);
xor XOR2 (N1172, N1167, N674);
not NOT1 (N1173, N1170);
and AND4 (N1174, N1169, N79, N1128, N892);
and AND4 (N1175, N1103, N1154, N884, N509);
not NOT1 (N1176, N1134);
xor XOR2 (N1177, N1162, N336);
nand NAND3 (N1178, N1177, N290, N571);
not NOT1 (N1179, N1172);
not NOT1 (N1180, N1179);
xor XOR2 (N1181, N1178, N476);
xor XOR2 (N1182, N1166, N619);
or OR3 (N1183, N1175, N159, N757);
and AND2 (N1184, N1152, N920);
not NOT1 (N1185, N1176);
not NOT1 (N1186, N1171);
nand NAND4 (N1187, N1184, N262, N515, N72);
nand NAND3 (N1188, N1181, N1020, N645);
nand NAND4 (N1189, N1188, N952, N1113, N405);
or OR2 (N1190, N1183, N421);
xor XOR2 (N1191, N1187, N614);
xor XOR2 (N1192, N1189, N501);
xor XOR2 (N1193, N1186, N290);
and AND4 (N1194, N1185, N489, N670, N990);
nand NAND3 (N1195, N1190, N787, N541);
and AND3 (N1196, N1194, N304, N680);
xor XOR2 (N1197, N1174, N543);
not NOT1 (N1198, N1191);
and AND3 (N1199, N1196, N11, N367);
not NOT1 (N1200, N1182);
and AND4 (N1201, N1160, N602, N404, N1168);
or OR2 (N1202, N1193, N621);
buf BUF1 (N1203, N1198);
nand NAND3 (N1204, N1199, N107, N201);
not NOT1 (N1205, N1180);
nor NOR3 (N1206, N1197, N1204, N664);
and AND2 (N1207, N871, N1039);
and AND4 (N1208, N1192, N617, N539, N891);
xor XOR2 (N1209, N1201, N884);
not NOT1 (N1210, N1203);
nor NOR2 (N1211, N1206, N36);
buf BUF1 (N1212, N1211);
and AND4 (N1213, N1208, N1024, N399, N791);
and AND3 (N1214, N1202, N342, N867);
not NOT1 (N1215, N1213);
xor XOR2 (N1216, N1210, N1168);
or OR2 (N1217, N1215, N301);
or OR3 (N1218, N1200, N824, N471);
buf BUF1 (N1219, N1173);
or OR2 (N1220, N1205, N348);
not NOT1 (N1221, N1217);
buf BUF1 (N1222, N1214);
and AND3 (N1223, N1218, N1104, N371);
not NOT1 (N1224, N1195);
nor NOR4 (N1225, N1216, N540, N509, N41);
xor XOR2 (N1226, N1222, N1158);
and AND3 (N1227, N1219, N454, N209);
nor NOR2 (N1228, N1221, N37);
not NOT1 (N1229, N1225);
and AND3 (N1230, N1226, N555, N613);
buf BUF1 (N1231, N1212);
xor XOR2 (N1232, N1228, N950);
xor XOR2 (N1233, N1220, N7);
nor NOR4 (N1234, N1207, N1122, N1188, N740);
not NOT1 (N1235, N1230);
nand NAND2 (N1236, N1227, N802);
not NOT1 (N1237, N1229);
or OR4 (N1238, N1209, N204, N135, N282);
nand NAND3 (N1239, N1224, N622, N96);
not NOT1 (N1240, N1238);
or OR3 (N1241, N1236, N26, N766);
nor NOR4 (N1242, N1234, N1004, N806, N783);
and AND2 (N1243, N1239, N823);
nor NOR3 (N1244, N1240, N1133, N162);
nand NAND4 (N1245, N1223, N1104, N1014, N527);
nor NOR3 (N1246, N1237, N410, N59);
buf BUF1 (N1247, N1241);
xor XOR2 (N1248, N1233, N119);
buf BUF1 (N1249, N1247);
nor NOR4 (N1250, N1235, N1144, N959, N930);
or OR4 (N1251, N1231, N521, N726, N526);
nand NAND2 (N1252, N1244, N863);
buf BUF1 (N1253, N1243);
not NOT1 (N1254, N1250);
and AND3 (N1255, N1245, N336, N11);
xor XOR2 (N1256, N1242, N18);
nor NOR4 (N1257, N1251, N719, N181, N536);
xor XOR2 (N1258, N1256, N595);
nand NAND3 (N1259, N1258, N816, N538);
not NOT1 (N1260, N1254);
not NOT1 (N1261, N1255);
xor XOR2 (N1262, N1260, N159);
and AND3 (N1263, N1253, N799, N1170);
or OR4 (N1264, N1263, N436, N677, N782);
not NOT1 (N1265, N1264);
buf BUF1 (N1266, N1249);
xor XOR2 (N1267, N1262, N865);
and AND3 (N1268, N1257, N467, N1061);
or OR3 (N1269, N1265, N734, N1156);
nand NAND4 (N1270, N1232, N1185, N1254, N118);
and AND4 (N1271, N1267, N1071, N185, N276);
nand NAND4 (N1272, N1248, N739, N1209, N387);
or OR4 (N1273, N1252, N837, N419, N1204);
nor NOR4 (N1274, N1266, N1132, N943, N350);
and AND3 (N1275, N1259, N596, N855);
and AND2 (N1276, N1274, N1019);
and AND2 (N1277, N1272, N6);
xor XOR2 (N1278, N1275, N179);
buf BUF1 (N1279, N1269);
and AND3 (N1280, N1270, N920, N487);
xor XOR2 (N1281, N1280, N1050);
nand NAND2 (N1282, N1246, N594);
buf BUF1 (N1283, N1277);
nand NAND3 (N1284, N1281, N491, N1234);
and AND2 (N1285, N1284, N1209);
buf BUF1 (N1286, N1276);
not NOT1 (N1287, N1279);
not NOT1 (N1288, N1261);
xor XOR2 (N1289, N1271, N107);
nor NOR2 (N1290, N1278, N1105);
or OR2 (N1291, N1287, N710);
or OR4 (N1292, N1285, N547, N558, N505);
nor NOR4 (N1293, N1290, N1137, N360, N249);
nor NOR4 (N1294, N1289, N132, N1157, N1025);
and AND3 (N1295, N1288, N605, N308);
and AND3 (N1296, N1268, N360, N66);
not NOT1 (N1297, N1283);
xor XOR2 (N1298, N1297, N1273);
buf BUF1 (N1299, N1105);
xor XOR2 (N1300, N1296, N1197);
nand NAND3 (N1301, N1293, N1158, N277);
buf BUF1 (N1302, N1298);
or OR4 (N1303, N1302, N525, N214, N350);
or OR2 (N1304, N1291, N354);
and AND4 (N1305, N1304, N1122, N474, N140);
nor NOR2 (N1306, N1299, N137);
or OR2 (N1307, N1306, N327);
and AND3 (N1308, N1301, N696, N430);
and AND4 (N1309, N1307, N1082, N453, N271);
or OR2 (N1310, N1292, N1181);
buf BUF1 (N1311, N1310);
xor XOR2 (N1312, N1311, N178);
nor NOR2 (N1313, N1282, N970);
nor NOR2 (N1314, N1300, N297);
not NOT1 (N1315, N1286);
buf BUF1 (N1316, N1313);
xor XOR2 (N1317, N1308, N227);
buf BUF1 (N1318, N1303);
xor XOR2 (N1319, N1316, N715);
and AND3 (N1320, N1317, N32, N95);
not NOT1 (N1321, N1305);
nand NAND3 (N1322, N1294, N464, N168);
not NOT1 (N1323, N1312);
and AND3 (N1324, N1321, N1155, N714);
and AND4 (N1325, N1319, N336, N981, N151);
nand NAND4 (N1326, N1323, N1038, N414, N247);
not NOT1 (N1327, N1295);
nand NAND4 (N1328, N1325, N192, N701, N533);
buf BUF1 (N1329, N1326);
not NOT1 (N1330, N1324);
nor NOR2 (N1331, N1327, N564);
xor XOR2 (N1332, N1330, N391);
and AND3 (N1333, N1328, N441, N160);
not NOT1 (N1334, N1314);
or OR4 (N1335, N1329, N82, N886, N346);
nand NAND4 (N1336, N1331, N1037, N873, N429);
xor XOR2 (N1337, N1322, N529);
and AND3 (N1338, N1334, N1297, N1031);
or OR2 (N1339, N1337, N510);
and AND2 (N1340, N1333, N1183);
not NOT1 (N1341, N1338);
xor XOR2 (N1342, N1340, N1043);
buf BUF1 (N1343, N1336);
not NOT1 (N1344, N1309);
nand NAND3 (N1345, N1339, N663, N1109);
not NOT1 (N1346, N1342);
buf BUF1 (N1347, N1343);
or OR4 (N1348, N1315, N516, N1113, N101);
buf BUF1 (N1349, N1348);
nand NAND2 (N1350, N1341, N1215);
or OR4 (N1351, N1349, N1349, N644, N284);
nor NOR3 (N1352, N1335, N151, N261);
nor NOR2 (N1353, N1352, N772);
nor NOR4 (N1354, N1350, N669, N1285, N519);
xor XOR2 (N1355, N1347, N447);
and AND4 (N1356, N1346, N552, N1352, N717);
and AND2 (N1357, N1320, N1262);
not NOT1 (N1358, N1357);
xor XOR2 (N1359, N1344, N526);
xor XOR2 (N1360, N1358, N525);
or OR2 (N1361, N1332, N821);
and AND3 (N1362, N1353, N1300, N97);
nor NOR4 (N1363, N1351, N652, N1142, N868);
nand NAND4 (N1364, N1318, N956, N138, N824);
nand NAND2 (N1365, N1364, N582);
and AND4 (N1366, N1365, N558, N31, N477);
xor XOR2 (N1367, N1356, N1365);
nor NOR4 (N1368, N1362, N807, N943, N1324);
buf BUF1 (N1369, N1355);
and AND4 (N1370, N1363, N395, N405, N576);
and AND4 (N1371, N1368, N730, N146, N243);
buf BUF1 (N1372, N1354);
nand NAND2 (N1373, N1371, N898);
nor NOR4 (N1374, N1367, N642, N40, N289);
xor XOR2 (N1375, N1372, N464);
not NOT1 (N1376, N1359);
nand NAND3 (N1377, N1361, N1256, N85);
or OR2 (N1378, N1345, N1037);
or OR2 (N1379, N1374, N489);
not NOT1 (N1380, N1373);
nand NAND2 (N1381, N1376, N705);
buf BUF1 (N1382, N1370);
and AND2 (N1383, N1369, N1050);
not NOT1 (N1384, N1366);
not NOT1 (N1385, N1380);
nand NAND3 (N1386, N1377, N116, N169);
or OR2 (N1387, N1383, N1215);
xor XOR2 (N1388, N1382, N408);
xor XOR2 (N1389, N1378, N858);
not NOT1 (N1390, N1360);
nor NOR2 (N1391, N1386, N1082);
xor XOR2 (N1392, N1384, N358);
not NOT1 (N1393, N1389);
nand NAND4 (N1394, N1379, N668, N1224, N1311);
and AND4 (N1395, N1388, N248, N997, N437);
nand NAND4 (N1396, N1390, N1371, N309, N11);
not NOT1 (N1397, N1395);
xor XOR2 (N1398, N1396, N877);
not NOT1 (N1399, N1397);
not NOT1 (N1400, N1375);
or OR4 (N1401, N1399, N744, N831, N1387);
and AND3 (N1402, N799, N1175, N411);
and AND2 (N1403, N1394, N1191);
or OR4 (N1404, N1393, N157, N1074, N1368);
xor XOR2 (N1405, N1404, N604);
nor NOR3 (N1406, N1400, N1033, N1329);
nor NOR3 (N1407, N1405, N1127, N60);
nor NOR2 (N1408, N1407, N821);
nor NOR2 (N1409, N1385, N283);
xor XOR2 (N1410, N1392, N853);
and AND2 (N1411, N1410, N685);
not NOT1 (N1412, N1401);
not NOT1 (N1413, N1391);
nor NOR2 (N1414, N1381, N992);
and AND2 (N1415, N1411, N949);
buf BUF1 (N1416, N1415);
nor NOR3 (N1417, N1403, N1228, N1119);
buf BUF1 (N1418, N1414);
nand NAND3 (N1419, N1398, N786, N156);
nand NAND4 (N1420, N1402, N78, N429, N1119);
and AND3 (N1421, N1406, N747, N1068);
and AND2 (N1422, N1417, N595);
xor XOR2 (N1423, N1419, N913);
not NOT1 (N1424, N1422);
or OR4 (N1425, N1420, N1136, N351, N293);
buf BUF1 (N1426, N1424);
not NOT1 (N1427, N1418);
buf BUF1 (N1428, N1421);
not NOT1 (N1429, N1416);
or OR2 (N1430, N1408, N1423);
xor XOR2 (N1431, N354, N900);
nor NOR3 (N1432, N1431, N410, N769);
and AND3 (N1433, N1432, N1035, N344);
not NOT1 (N1434, N1409);
nor NOR2 (N1435, N1425, N528);
or OR4 (N1436, N1433, N184, N1248, N19);
nand NAND4 (N1437, N1428, N795, N600, N480);
xor XOR2 (N1438, N1435, N873);
not NOT1 (N1439, N1429);
and AND4 (N1440, N1438, N594, N232, N1299);
and AND3 (N1441, N1436, N592, N1406);
nor NOR4 (N1442, N1441, N908, N773, N915);
buf BUF1 (N1443, N1434);
not NOT1 (N1444, N1427);
not NOT1 (N1445, N1413);
nor NOR3 (N1446, N1430, N1058, N1105);
or OR4 (N1447, N1426, N1097, N436, N945);
buf BUF1 (N1448, N1412);
xor XOR2 (N1449, N1439, N1116);
and AND2 (N1450, N1447, N846);
not NOT1 (N1451, N1437);
nor NOR2 (N1452, N1445, N165);
buf BUF1 (N1453, N1448);
xor XOR2 (N1454, N1453, N471);
xor XOR2 (N1455, N1443, N1171);
nor NOR2 (N1456, N1449, N137);
buf BUF1 (N1457, N1446);
nor NOR3 (N1458, N1452, N279, N203);
or OR2 (N1459, N1454, N459);
not NOT1 (N1460, N1442);
nand NAND2 (N1461, N1457, N14);
and AND4 (N1462, N1461, N972, N1166, N1033);
and AND4 (N1463, N1440, N430, N72, N118);
not NOT1 (N1464, N1450);
buf BUF1 (N1465, N1460);
nand NAND4 (N1466, N1459, N1298, N544, N1445);
not NOT1 (N1467, N1466);
xor XOR2 (N1468, N1465, N831);
not NOT1 (N1469, N1462);
buf BUF1 (N1470, N1444);
nand NAND4 (N1471, N1469, N642, N861, N413);
or OR2 (N1472, N1471, N420);
nor NOR2 (N1473, N1472, N399);
nand NAND2 (N1474, N1456, N1254);
not NOT1 (N1475, N1451);
nor NOR2 (N1476, N1474, N921);
nand NAND3 (N1477, N1476, N886, N385);
nor NOR4 (N1478, N1477, N400, N818, N1456);
and AND3 (N1479, N1458, N844, N53);
or OR3 (N1480, N1464, N1024, N139);
or OR3 (N1481, N1467, N1264, N1235);
xor XOR2 (N1482, N1468, N1124);
nand NAND3 (N1483, N1480, N607, N968);
or OR4 (N1484, N1473, N291, N391, N1415);
nand NAND2 (N1485, N1481, N750);
nor NOR4 (N1486, N1484, N1409, N295, N1029);
or OR3 (N1487, N1483, N451, N1434);
nor NOR3 (N1488, N1455, N1273, N1400);
xor XOR2 (N1489, N1486, N1404);
xor XOR2 (N1490, N1475, N1114);
and AND3 (N1491, N1487, N1312, N906);
xor XOR2 (N1492, N1489, N275);
xor XOR2 (N1493, N1478, N1420);
nor NOR2 (N1494, N1470, N1107);
xor XOR2 (N1495, N1463, N638);
buf BUF1 (N1496, N1482);
xor XOR2 (N1497, N1495, N115);
or OR2 (N1498, N1488, N699);
buf BUF1 (N1499, N1494);
not NOT1 (N1500, N1498);
and AND2 (N1501, N1499, N184);
buf BUF1 (N1502, N1501);
nand NAND3 (N1503, N1500, N209, N447);
buf BUF1 (N1504, N1503);
and AND3 (N1505, N1504, N1230, N862);
and AND3 (N1506, N1502, N1421, N882);
nor NOR2 (N1507, N1493, N1222);
not NOT1 (N1508, N1505);
or OR3 (N1509, N1492, N391, N181);
nand NAND4 (N1510, N1490, N1132, N1155, N226);
buf BUF1 (N1511, N1497);
buf BUF1 (N1512, N1511);
nor NOR2 (N1513, N1491, N739);
xor XOR2 (N1514, N1479, N1439);
xor XOR2 (N1515, N1512, N1442);
nand NAND4 (N1516, N1514, N246, N899, N67);
or OR3 (N1517, N1509, N968, N1487);
buf BUF1 (N1518, N1517);
not NOT1 (N1519, N1510);
buf BUF1 (N1520, N1508);
buf BUF1 (N1521, N1516);
buf BUF1 (N1522, N1520);
and AND3 (N1523, N1519, N153, N36);
nor NOR2 (N1524, N1506, N869);
buf BUF1 (N1525, N1518);
buf BUF1 (N1526, N1525);
xor XOR2 (N1527, N1513, N775);
nand NAND3 (N1528, N1522, N587, N656);
and AND2 (N1529, N1485, N1284);
not NOT1 (N1530, N1507);
xor XOR2 (N1531, N1524, N1284);
and AND4 (N1532, N1528, N1365, N1381, N222);
not NOT1 (N1533, N1530);
or OR4 (N1534, N1533, N12, N167, N933);
or OR2 (N1535, N1526, N642);
and AND2 (N1536, N1531, N718);
xor XOR2 (N1537, N1532, N306);
nand NAND2 (N1538, N1521, N1527);
xor XOR2 (N1539, N678, N492);
nor NOR3 (N1540, N1523, N1437, N309);
nor NOR3 (N1541, N1537, N288, N1033);
and AND3 (N1542, N1515, N969, N1322);
nor NOR2 (N1543, N1535, N853);
xor XOR2 (N1544, N1539, N214);
buf BUF1 (N1545, N1541);
buf BUF1 (N1546, N1542);
buf BUF1 (N1547, N1538);
and AND4 (N1548, N1543, N662, N699, N501);
xor XOR2 (N1549, N1545, N1212);
nor NOR4 (N1550, N1548, N775, N500, N895);
nand NAND4 (N1551, N1544, N531, N1335, N1031);
xor XOR2 (N1552, N1529, N1476);
and AND4 (N1553, N1534, N555, N1290, N846);
nor NOR2 (N1554, N1550, N608);
buf BUF1 (N1555, N1540);
not NOT1 (N1556, N1547);
not NOT1 (N1557, N1552);
xor XOR2 (N1558, N1554, N711);
xor XOR2 (N1559, N1553, N1051);
nor NOR4 (N1560, N1549, N746, N1039, N972);
nand NAND4 (N1561, N1551, N1132, N655, N1228);
xor XOR2 (N1562, N1536, N115);
xor XOR2 (N1563, N1496, N148);
buf BUF1 (N1564, N1562);
nor NOR4 (N1565, N1563, N52, N1354, N160);
and AND2 (N1566, N1559, N1144);
buf BUF1 (N1567, N1561);
and AND4 (N1568, N1555, N354, N1238, N270);
or OR2 (N1569, N1546, N554);
buf BUF1 (N1570, N1560);
xor XOR2 (N1571, N1569, N1555);
buf BUF1 (N1572, N1566);
buf BUF1 (N1573, N1570);
and AND3 (N1574, N1567, N1462, N1078);
or OR2 (N1575, N1574, N55);
buf BUF1 (N1576, N1573);
buf BUF1 (N1577, N1565);
or OR3 (N1578, N1575, N1087, N458);
or OR2 (N1579, N1568, N29);
or OR4 (N1580, N1558, N1299, N785, N1395);
or OR3 (N1581, N1577, N1318, N5);
or OR3 (N1582, N1576, N520, N756);
not NOT1 (N1583, N1582);
nor NOR3 (N1584, N1556, N285, N1123);
and AND4 (N1585, N1557, N20, N1069, N1033);
buf BUF1 (N1586, N1581);
not NOT1 (N1587, N1585);
or OR4 (N1588, N1564, N1279, N1167, N1005);
and AND4 (N1589, N1580, N1093, N1420, N326);
or OR2 (N1590, N1572, N1056);
xor XOR2 (N1591, N1578, N127);
and AND4 (N1592, N1588, N631, N978, N617);
or OR4 (N1593, N1589, N1549, N1213, N696);
not NOT1 (N1594, N1590);
or OR4 (N1595, N1591, N1237, N1527, N694);
and AND4 (N1596, N1593, N816, N19, N1514);
nand NAND2 (N1597, N1594, N377);
not NOT1 (N1598, N1584);
buf BUF1 (N1599, N1583);
buf BUF1 (N1600, N1592);
buf BUF1 (N1601, N1595);
xor XOR2 (N1602, N1598, N854);
not NOT1 (N1603, N1596);
not NOT1 (N1604, N1579);
and AND4 (N1605, N1599, N1268, N239, N1163);
nor NOR4 (N1606, N1601, N35, N1100, N296);
not NOT1 (N1607, N1571);
buf BUF1 (N1608, N1606);
or OR4 (N1609, N1586, N930, N1081, N1288);
or OR4 (N1610, N1597, N1366, N983, N128);
xor XOR2 (N1611, N1605, N242);
nor NOR3 (N1612, N1604, N118, N817);
nor NOR2 (N1613, N1609, N11);
or OR3 (N1614, N1602, N981, N16);
nand NAND2 (N1615, N1607, N734);
not NOT1 (N1616, N1610);
not NOT1 (N1617, N1600);
nand NAND2 (N1618, N1613, N295);
buf BUF1 (N1619, N1603);
nand NAND2 (N1620, N1612, N1034);
nor NOR2 (N1621, N1616, N370);
and AND3 (N1622, N1611, N849, N1575);
buf BUF1 (N1623, N1587);
or OR2 (N1624, N1622, N1618);
nand NAND2 (N1625, N95, N397);
nor NOR3 (N1626, N1608, N879, N124);
nor NOR3 (N1627, N1614, N628, N1433);
not NOT1 (N1628, N1627);
buf BUF1 (N1629, N1619);
xor XOR2 (N1630, N1617, N915);
buf BUF1 (N1631, N1623);
and AND2 (N1632, N1624, N369);
and AND2 (N1633, N1620, N1255);
or OR2 (N1634, N1631, N368);
buf BUF1 (N1635, N1626);
and AND3 (N1636, N1634, N1430, N1507);
buf BUF1 (N1637, N1628);
nor NOR3 (N1638, N1625, N1592, N529);
nor NOR2 (N1639, N1638, N1563);
nand NAND4 (N1640, N1633, N1115, N300, N448);
not NOT1 (N1641, N1640);
and AND2 (N1642, N1635, N314);
not NOT1 (N1643, N1641);
buf BUF1 (N1644, N1642);
and AND2 (N1645, N1621, N68);
or OR2 (N1646, N1644, N1345);
xor XOR2 (N1647, N1645, N78);
nor NOR4 (N1648, N1639, N1342, N717, N57);
xor XOR2 (N1649, N1629, N630);
buf BUF1 (N1650, N1648);
xor XOR2 (N1651, N1636, N1530);
buf BUF1 (N1652, N1615);
xor XOR2 (N1653, N1632, N258);
or OR2 (N1654, N1647, N1197);
nand NAND2 (N1655, N1646, N1396);
buf BUF1 (N1656, N1643);
not NOT1 (N1657, N1656);
nand NAND3 (N1658, N1652, N1391, N96);
buf BUF1 (N1659, N1658);
not NOT1 (N1660, N1649);
not NOT1 (N1661, N1657);
and AND3 (N1662, N1660, N896, N1337);
xor XOR2 (N1663, N1637, N1428);
nand NAND2 (N1664, N1630, N5);
or OR4 (N1665, N1661, N1509, N82, N1077);
nor NOR3 (N1666, N1654, N1442, N1549);
nor NOR2 (N1667, N1659, N392);
buf BUF1 (N1668, N1666);
and AND3 (N1669, N1650, N509, N1656);
not NOT1 (N1670, N1665);
or OR3 (N1671, N1662, N727, N1329);
or OR2 (N1672, N1671, N449);
and AND2 (N1673, N1672, N35);
not NOT1 (N1674, N1667);
xor XOR2 (N1675, N1655, N1538);
nand NAND3 (N1676, N1673, N1651, N619);
xor XOR2 (N1677, N211, N1420);
and AND2 (N1678, N1670, N856);
and AND4 (N1679, N1675, N866, N383, N1374);
buf BUF1 (N1680, N1678);
or OR4 (N1681, N1664, N1347, N1612, N437);
buf BUF1 (N1682, N1680);
and AND3 (N1683, N1669, N776, N1117);
xor XOR2 (N1684, N1676, N150);
not NOT1 (N1685, N1674);
not NOT1 (N1686, N1653);
xor XOR2 (N1687, N1668, N1566);
or OR2 (N1688, N1686, N342);
buf BUF1 (N1689, N1683);
xor XOR2 (N1690, N1677, N836);
not NOT1 (N1691, N1690);
not NOT1 (N1692, N1685);
not NOT1 (N1693, N1684);
or OR4 (N1694, N1691, N1552, N9, N1669);
xor XOR2 (N1695, N1694, N49);
and AND3 (N1696, N1688, N291, N484);
and AND2 (N1697, N1682, N202);
buf BUF1 (N1698, N1663);
nor NOR4 (N1699, N1692, N467, N990, N895);
or OR4 (N1700, N1698, N1083, N1143, N1552);
nor NOR4 (N1701, N1693, N508, N276, N628);
nand NAND2 (N1702, N1697, N136);
not NOT1 (N1703, N1689);
or OR2 (N1704, N1702, N207);
or OR4 (N1705, N1700, N918, N154, N609);
xor XOR2 (N1706, N1695, N1352);
xor XOR2 (N1707, N1705, N1370);
not NOT1 (N1708, N1696);
nand NAND3 (N1709, N1708, N942, N44);
xor XOR2 (N1710, N1709, N267);
not NOT1 (N1711, N1706);
nor NOR3 (N1712, N1703, N1183, N264);
or OR2 (N1713, N1679, N1497);
and AND2 (N1714, N1699, N1349);
and AND3 (N1715, N1687, N1164, N1398);
not NOT1 (N1716, N1712);
nor NOR3 (N1717, N1681, N143, N934);
or OR4 (N1718, N1713, N394, N855, N1715);
not NOT1 (N1719, N231);
nand NAND3 (N1720, N1714, N38, N651);
nand NAND4 (N1721, N1716, N804, N1251, N26);
buf BUF1 (N1722, N1721);
buf BUF1 (N1723, N1704);
and AND4 (N1724, N1718, N1213, N1646, N1323);
nand NAND2 (N1725, N1719, N1633);
and AND4 (N1726, N1724, N309, N1590, N216);
or OR4 (N1727, N1720, N849, N376, N1685);
or OR4 (N1728, N1723, N1296, N480, N1204);
xor XOR2 (N1729, N1725, N1476);
buf BUF1 (N1730, N1711);
nand NAND2 (N1731, N1722, N433);
nand NAND4 (N1732, N1730, N474, N980, N1719);
or OR2 (N1733, N1728, N1219);
nand NAND4 (N1734, N1733, N841, N1164, N910);
nand NAND4 (N1735, N1731, N519, N1356, N1265);
buf BUF1 (N1736, N1727);
or OR2 (N1737, N1732, N355);
xor XOR2 (N1738, N1717, N496);
xor XOR2 (N1739, N1707, N1459);
nor NOR4 (N1740, N1710, N1616, N1041, N438);
buf BUF1 (N1741, N1729);
xor XOR2 (N1742, N1737, N917);
nand NAND4 (N1743, N1726, N646, N1127, N915);
or OR2 (N1744, N1738, N442);
buf BUF1 (N1745, N1740);
xor XOR2 (N1746, N1742, N78);
not NOT1 (N1747, N1741);
buf BUF1 (N1748, N1736);
not NOT1 (N1749, N1746);
nor NOR4 (N1750, N1743, N927, N1724, N1007);
buf BUF1 (N1751, N1748);
nand NAND3 (N1752, N1749, N786, N281);
and AND3 (N1753, N1751, N934, N1109);
nor NOR2 (N1754, N1752, N184);
buf BUF1 (N1755, N1735);
nor NOR3 (N1756, N1753, N1750, N1525);
or OR3 (N1757, N1686, N1265, N900);
not NOT1 (N1758, N1744);
nand NAND4 (N1759, N1745, N1023, N457, N144);
not NOT1 (N1760, N1701);
buf BUF1 (N1761, N1757);
or OR4 (N1762, N1739, N1396, N1072, N1274);
and AND2 (N1763, N1755, N1550);
and AND4 (N1764, N1756, N286, N1305, N1335);
nand NAND2 (N1765, N1760, N274);
buf BUF1 (N1766, N1761);
nor NOR4 (N1767, N1734, N1206, N294, N590);
buf BUF1 (N1768, N1763);
xor XOR2 (N1769, N1765, N377);
xor XOR2 (N1770, N1762, N1558);
buf BUF1 (N1771, N1768);
buf BUF1 (N1772, N1769);
and AND3 (N1773, N1758, N757, N1687);
and AND3 (N1774, N1771, N173, N765);
nand NAND4 (N1775, N1773, N1571, N862, N405);
and AND2 (N1776, N1766, N1462);
or OR4 (N1777, N1759, N941, N622, N854);
nor NOR2 (N1778, N1747, N1297);
nor NOR3 (N1779, N1774, N100, N1774);
nor NOR2 (N1780, N1767, N1703);
nand NAND4 (N1781, N1772, N332, N1680, N1090);
and AND2 (N1782, N1770, N1037);
and AND4 (N1783, N1775, N642, N1750, N1754);
buf BUF1 (N1784, N573);
xor XOR2 (N1785, N1776, N114);
and AND3 (N1786, N1780, N480, N1144);
buf BUF1 (N1787, N1781);
xor XOR2 (N1788, N1778, N1677);
nor NOR2 (N1789, N1777, N738);
and AND3 (N1790, N1785, N457, N117);
buf BUF1 (N1791, N1764);
or OR3 (N1792, N1787, N175, N1770);
nand NAND2 (N1793, N1789, N1425);
buf BUF1 (N1794, N1784);
nor NOR4 (N1795, N1788, N279, N424, N1573);
nor NOR3 (N1796, N1794, N1231, N577);
nand NAND4 (N1797, N1783, N682, N1653, N666);
and AND2 (N1798, N1791, N806);
xor XOR2 (N1799, N1798, N1666);
nor NOR4 (N1800, N1797, N757, N176, N451);
buf BUF1 (N1801, N1790);
nor NOR3 (N1802, N1800, N290, N168);
or OR2 (N1803, N1779, N748);
and AND3 (N1804, N1799, N12, N1171);
and AND2 (N1805, N1792, N603);
not NOT1 (N1806, N1801);
nor NOR4 (N1807, N1803, N1704, N957, N63);
buf BUF1 (N1808, N1802);
xor XOR2 (N1809, N1804, N384);
xor XOR2 (N1810, N1808, N964);
or OR4 (N1811, N1809, N700, N390, N1414);
and AND2 (N1812, N1806, N1447);
or OR3 (N1813, N1805, N855, N323);
buf BUF1 (N1814, N1795);
not NOT1 (N1815, N1810);
and AND2 (N1816, N1796, N852);
nand NAND3 (N1817, N1811, N1719, N783);
or OR4 (N1818, N1816, N1440, N1299, N54);
buf BUF1 (N1819, N1807);
not NOT1 (N1820, N1793);
buf BUF1 (N1821, N1818);
nand NAND2 (N1822, N1786, N712);
and AND4 (N1823, N1813, N965, N1071, N45);
nor NOR3 (N1824, N1814, N1023, N354);
not NOT1 (N1825, N1817);
or OR2 (N1826, N1819, N1223);
nor NOR4 (N1827, N1822, N211, N1788, N42);
xor XOR2 (N1828, N1821, N1623);
or OR3 (N1829, N1825, N1640, N404);
xor XOR2 (N1830, N1827, N495);
nand NAND2 (N1831, N1823, N1286);
xor XOR2 (N1832, N1820, N1013);
and AND2 (N1833, N1831, N340);
or OR2 (N1834, N1833, N1407);
buf BUF1 (N1835, N1824);
nor NOR4 (N1836, N1832, N1560, N581, N991);
or OR4 (N1837, N1829, N1047, N190, N1719);
not NOT1 (N1838, N1815);
and AND4 (N1839, N1826, N1087, N744, N53);
not NOT1 (N1840, N1838);
buf BUF1 (N1841, N1830);
or OR2 (N1842, N1837, N929);
xor XOR2 (N1843, N1782, N298);
xor XOR2 (N1844, N1840, N61);
nor NOR4 (N1845, N1835, N1467, N1515, N1682);
or OR2 (N1846, N1842, N2);
nor NOR4 (N1847, N1828, N794, N1707, N1039);
not NOT1 (N1848, N1836);
nor NOR4 (N1849, N1839, N517, N815, N469);
xor XOR2 (N1850, N1848, N918);
xor XOR2 (N1851, N1834, N1206);
nand NAND2 (N1852, N1846, N1479);
nand NAND3 (N1853, N1845, N1701, N430);
nand NAND4 (N1854, N1844, N24, N575, N742);
not NOT1 (N1855, N1854);
buf BUF1 (N1856, N1853);
xor XOR2 (N1857, N1850, N633);
not NOT1 (N1858, N1856);
nand NAND3 (N1859, N1855, N771, N1782);
or OR4 (N1860, N1812, N764, N833, N1500);
or OR4 (N1861, N1847, N1820, N121, N1813);
nand NAND3 (N1862, N1861, N355, N41);
nor NOR2 (N1863, N1858, N1330);
buf BUF1 (N1864, N1857);
not NOT1 (N1865, N1849);
xor XOR2 (N1866, N1864, N818);
or OR4 (N1867, N1866, N239, N1711, N15);
nor NOR2 (N1868, N1860, N1648);
xor XOR2 (N1869, N1862, N597);
and AND4 (N1870, N1869, N454, N559, N1271);
buf BUF1 (N1871, N1859);
buf BUF1 (N1872, N1851);
or OR4 (N1873, N1841, N654, N1312, N1715);
nand NAND2 (N1874, N1868, N311);
and AND2 (N1875, N1863, N1643);
xor XOR2 (N1876, N1865, N1285);
nor NOR2 (N1877, N1872, N140);
nor NOR2 (N1878, N1870, N1316);
or OR2 (N1879, N1874, N1126);
and AND4 (N1880, N1867, N157, N1811, N316);
and AND4 (N1881, N1843, N134, N650, N1119);
buf BUF1 (N1882, N1881);
or OR3 (N1883, N1880, N1433, N1014);
not NOT1 (N1884, N1883);
nor NOR2 (N1885, N1873, N282);
nor NOR3 (N1886, N1879, N1271, N1702);
not NOT1 (N1887, N1876);
not NOT1 (N1888, N1877);
buf BUF1 (N1889, N1878);
nor NOR4 (N1890, N1884, N821, N781, N1045);
nand NAND2 (N1891, N1886, N570);
and AND2 (N1892, N1891, N1675);
buf BUF1 (N1893, N1889);
nand NAND3 (N1894, N1882, N922, N1473);
not NOT1 (N1895, N1852);
or OR3 (N1896, N1885, N1124, N682);
nor NOR4 (N1897, N1871, N244, N593, N1093);
nand NAND3 (N1898, N1887, N225, N1269);
nor NOR4 (N1899, N1898, N1645, N274, N1561);
nor NOR2 (N1900, N1895, N1065);
or OR4 (N1901, N1875, N423, N381, N487);
nor NOR2 (N1902, N1896, N788);
buf BUF1 (N1903, N1890);
nand NAND2 (N1904, N1894, N1064);
buf BUF1 (N1905, N1902);
xor XOR2 (N1906, N1900, N1851);
nand NAND3 (N1907, N1892, N1901, N171);
xor XOR2 (N1908, N394, N878);
nor NOR4 (N1909, N1888, N1566, N376, N986);
nor NOR3 (N1910, N1903, N973, N1148);
xor XOR2 (N1911, N1893, N776);
not NOT1 (N1912, N1909);
nor NOR4 (N1913, N1904, N1584, N127, N260);
nor NOR4 (N1914, N1912, N378, N1034, N31);
not NOT1 (N1915, N1908);
buf BUF1 (N1916, N1915);
nand NAND4 (N1917, N1916, N1470, N41, N1226);
nand NAND3 (N1918, N1913, N1582, N1300);
or OR3 (N1919, N1910, N372, N862);
and AND3 (N1920, N1917, N306, N1904);
nand NAND2 (N1921, N1920, N884);
xor XOR2 (N1922, N1921, N285);
and AND3 (N1923, N1899, N1451, N1071);
nor NOR4 (N1924, N1922, N458, N303, N611);
buf BUF1 (N1925, N1897);
not NOT1 (N1926, N1924);
nor NOR2 (N1927, N1926, N1375);
xor XOR2 (N1928, N1914, N668);
nand NAND3 (N1929, N1911, N1584, N1051);
buf BUF1 (N1930, N1923);
and AND3 (N1931, N1905, N1267, N895);
buf BUF1 (N1932, N1930);
or OR3 (N1933, N1925, N1688, N451);
xor XOR2 (N1934, N1907, N110);
xor XOR2 (N1935, N1928, N779);
not NOT1 (N1936, N1919);
not NOT1 (N1937, N1929);
nand NAND3 (N1938, N1931, N536, N360);
not NOT1 (N1939, N1935);
and AND2 (N1940, N1938, N1800);
and AND2 (N1941, N1936, N1000);
or OR4 (N1942, N1940, N1200, N1666, N1750);
nand NAND3 (N1943, N1941, N1266, N1788);
not NOT1 (N1944, N1906);
or OR2 (N1945, N1927, N241);
buf BUF1 (N1946, N1933);
and AND2 (N1947, N1918, N1840);
buf BUF1 (N1948, N1946);
xor XOR2 (N1949, N1937, N616);
buf BUF1 (N1950, N1945);
and AND4 (N1951, N1949, N328, N912, N1315);
buf BUF1 (N1952, N1951);
or OR3 (N1953, N1948, N1872, N1560);
or OR2 (N1954, N1942, N47);
nor NOR2 (N1955, N1952, N861);
and AND4 (N1956, N1953, N1192, N365, N1638);
nand NAND2 (N1957, N1950, N836);
or OR3 (N1958, N1954, N22, N48);
and AND3 (N1959, N1944, N1762, N1265);
nor NOR4 (N1960, N1934, N410, N745, N1522);
nor NOR2 (N1961, N1956, N193);
xor XOR2 (N1962, N1943, N1876);
buf BUF1 (N1963, N1961);
or OR3 (N1964, N1959, N1148, N1388);
nand NAND2 (N1965, N1947, N1524);
nor NOR4 (N1966, N1957, N1302, N1351, N994);
not NOT1 (N1967, N1965);
xor XOR2 (N1968, N1955, N1525);
not NOT1 (N1969, N1968);
nand NAND2 (N1970, N1939, N1402);
buf BUF1 (N1971, N1969);
nor NOR2 (N1972, N1958, N1894);
not NOT1 (N1973, N1964);
xor XOR2 (N1974, N1966, N1129);
not NOT1 (N1975, N1960);
not NOT1 (N1976, N1971);
nand NAND3 (N1977, N1972, N518, N407);
and AND4 (N1978, N1973, N200, N543, N747);
nor NOR3 (N1979, N1962, N1079, N1399);
xor XOR2 (N1980, N1975, N1782);
nand NAND2 (N1981, N1977, N1393);
not NOT1 (N1982, N1967);
or OR4 (N1983, N1932, N1622, N820, N245);
nand NAND2 (N1984, N1970, N995);
nand NAND4 (N1985, N1974, N1094, N580, N1453);
nand NAND2 (N1986, N1978, N1157);
nor NOR3 (N1987, N1986, N1683, N1729);
nor NOR3 (N1988, N1980, N1935, N991);
or OR2 (N1989, N1985, N1653);
and AND4 (N1990, N1987, N1450, N876, N1530);
or OR4 (N1991, N1982, N943, N928, N145);
and AND3 (N1992, N1989, N798, N42);
xor XOR2 (N1993, N1979, N1223);
not NOT1 (N1994, N1990);
or OR2 (N1995, N1991, N928);
and AND4 (N1996, N1994, N102, N1645, N299);
not NOT1 (N1997, N1993);
nand NAND2 (N1998, N1997, N1416);
nor NOR2 (N1999, N1995, N1767);
buf BUF1 (N2000, N1988);
not NOT1 (N2001, N2000);
nor NOR2 (N2002, N1981, N18);
nor NOR3 (N2003, N1984, N26, N805);
or OR2 (N2004, N1992, N1055);
not NOT1 (N2005, N1976);
nand NAND4 (N2006, N1983, N979, N1731, N1789);
xor XOR2 (N2007, N1996, N1714);
nor NOR4 (N2008, N2004, N354, N427, N1254);
nand NAND4 (N2009, N2006, N1768, N1753, N279);
or OR3 (N2010, N2001, N1597, N411);
buf BUF1 (N2011, N2007);
nand NAND2 (N2012, N2011, N1543);
xor XOR2 (N2013, N1999, N762);
and AND4 (N2014, N1998, N732, N436, N1480);
xor XOR2 (N2015, N2014, N1859);
buf BUF1 (N2016, N2008);
buf BUF1 (N2017, N2016);
nand NAND3 (N2018, N2012, N491, N911);
and AND4 (N2019, N2018, N1800, N1268, N1089);
and AND4 (N2020, N2015, N965, N878, N1325);
nand NAND2 (N2021, N1963, N237);
buf BUF1 (N2022, N2017);
and AND3 (N2023, N2005, N164, N1558);
xor XOR2 (N2024, N2023, N1189);
buf BUF1 (N2025, N2002);
buf BUF1 (N2026, N2003);
not NOT1 (N2027, N2022);
and AND2 (N2028, N2013, N1871);
nand NAND3 (N2029, N2009, N606, N1602);
nand NAND2 (N2030, N2019, N1115);
not NOT1 (N2031, N2010);
or OR2 (N2032, N2026, N403);
not NOT1 (N2033, N2031);
and AND2 (N2034, N2029, N418);
nor NOR3 (N2035, N2027, N293, N87);
xor XOR2 (N2036, N2020, N508);
not NOT1 (N2037, N2034);
nor NOR4 (N2038, N2021, N803, N378, N1659);
nor NOR2 (N2039, N2036, N801);
nand NAND2 (N2040, N2035, N652);
and AND3 (N2041, N2025, N687, N27);
buf BUF1 (N2042, N2038);
not NOT1 (N2043, N2030);
buf BUF1 (N2044, N2033);
xor XOR2 (N2045, N2032, N1343);
not NOT1 (N2046, N2044);
buf BUF1 (N2047, N2028);
xor XOR2 (N2048, N2047, N896);
buf BUF1 (N2049, N2041);
nand NAND3 (N2050, N2042, N672, N89);
nand NAND4 (N2051, N2046, N678, N743, N781);
and AND4 (N2052, N2037, N288, N1122, N467);
buf BUF1 (N2053, N2049);
buf BUF1 (N2054, N2045);
nand NAND3 (N2055, N2053, N1148, N1060);
buf BUF1 (N2056, N2039);
xor XOR2 (N2057, N2054, N1810);
buf BUF1 (N2058, N2051);
nand NAND4 (N2059, N2040, N828, N1998, N1246);
nor NOR2 (N2060, N2052, N2038);
xor XOR2 (N2061, N2043, N718);
or OR3 (N2062, N2050, N1274, N1117);
nand NAND2 (N2063, N2024, N1720);
or OR3 (N2064, N2057, N730, N834);
buf BUF1 (N2065, N2062);
or OR2 (N2066, N2065, N660);
nor NOR2 (N2067, N2066, N2022);
buf BUF1 (N2068, N2061);
nand NAND4 (N2069, N2059, N1134, N1072, N1990);
buf BUF1 (N2070, N2048);
or OR4 (N2071, N2056, N21, N142, N851);
nor NOR2 (N2072, N2071, N1999);
xor XOR2 (N2073, N2060, N1972);
and AND3 (N2074, N2055, N1268, N1727);
nor NOR2 (N2075, N2069, N1285);
not NOT1 (N2076, N2074);
xor XOR2 (N2077, N2068, N1340);
nand NAND4 (N2078, N2073, N91, N798, N752);
nand NAND2 (N2079, N2078, N1958);
nor NOR3 (N2080, N2076, N1286, N1722);
and AND3 (N2081, N2070, N397, N457);
nand NAND3 (N2082, N2063, N1138, N1829);
nand NAND2 (N2083, N2081, N1833);
and AND2 (N2084, N2067, N234);
nor NOR3 (N2085, N2082, N245, N181);
nor NOR2 (N2086, N2064, N1896);
nor NOR3 (N2087, N2084, N330, N1886);
or OR2 (N2088, N2080, N1696);
xor XOR2 (N2089, N2077, N154);
buf BUF1 (N2090, N2085);
or OR3 (N2091, N2072, N1760, N614);
and AND4 (N2092, N2079, N223, N1369, N429);
buf BUF1 (N2093, N2090);
or OR2 (N2094, N2058, N173);
or OR4 (N2095, N2088, N2040, N1891, N1765);
nand NAND3 (N2096, N2095, N1451, N431);
nand NAND3 (N2097, N2091, N740, N119);
or OR4 (N2098, N2093, N906, N638, N183);
not NOT1 (N2099, N2089);
and AND2 (N2100, N2099, N1613);
not NOT1 (N2101, N2075);
and AND3 (N2102, N2087, N1025, N752);
or OR2 (N2103, N2100, N333);
buf BUF1 (N2104, N2101);
and AND3 (N2105, N2097, N1866, N1978);
xor XOR2 (N2106, N2104, N892);
not NOT1 (N2107, N2096);
nand NAND4 (N2108, N2103, N502, N46, N1928);
nor NOR2 (N2109, N2083, N1705);
or OR2 (N2110, N2102, N1049);
xor XOR2 (N2111, N2094, N1334);
or OR2 (N2112, N2098, N197);
not NOT1 (N2113, N2110);
not NOT1 (N2114, N2108);
buf BUF1 (N2115, N2086);
nor NOR2 (N2116, N2092, N1354);
buf BUF1 (N2117, N2111);
nand NAND3 (N2118, N2114, N455, N1229);
nand NAND4 (N2119, N2112, N943, N158, N1725);
nor NOR3 (N2120, N2115, N2016, N1092);
xor XOR2 (N2121, N2117, N1335);
nor NOR3 (N2122, N2109, N1747, N68);
nand NAND2 (N2123, N2121, N416);
not NOT1 (N2124, N2119);
xor XOR2 (N2125, N2120, N1794);
or OR3 (N2126, N2116, N1856, N1184);
nor NOR3 (N2127, N2123, N1071, N1151);
or OR2 (N2128, N2125, N1158);
nand NAND4 (N2129, N2118, N1108, N1786, N509);
or OR4 (N2130, N2129, N1509, N1957, N1621);
and AND3 (N2131, N2126, N1865, N2075);
nand NAND4 (N2132, N2131, N647, N232, N624);
nand NAND4 (N2133, N2130, N1967, N1355, N1149);
nor NOR3 (N2134, N2122, N961, N1779);
nand NAND2 (N2135, N2107, N1906);
buf BUF1 (N2136, N2105);
and AND3 (N2137, N2128, N443, N552);
xor XOR2 (N2138, N2106, N757);
nor NOR4 (N2139, N2133, N188, N1669, N550);
nor NOR3 (N2140, N2113, N1227, N1235);
or OR3 (N2141, N2140, N729, N1175);
nand NAND4 (N2142, N2127, N1610, N725, N127);
and AND2 (N2143, N2139, N975);
and AND2 (N2144, N2142, N315);
or OR3 (N2145, N2138, N1037, N1560);
nor NOR3 (N2146, N2141, N1280, N726);
xor XOR2 (N2147, N2132, N1500);
or OR4 (N2148, N2135, N865, N731, N1643);
and AND2 (N2149, N2143, N239);
or OR3 (N2150, N2147, N1126, N245);
not NOT1 (N2151, N2134);
buf BUF1 (N2152, N2137);
xor XOR2 (N2153, N2152, N967);
nand NAND4 (N2154, N2149, N920, N1243, N1973);
not NOT1 (N2155, N2124);
nor NOR4 (N2156, N2148, N1589, N1377, N963);
not NOT1 (N2157, N2145);
and AND2 (N2158, N2155, N481);
nor NOR3 (N2159, N2146, N457, N1970);
and AND3 (N2160, N2150, N204, N1643);
buf BUF1 (N2161, N2153);
and AND4 (N2162, N2160, N938, N1693, N563);
nand NAND3 (N2163, N2151, N181, N326);
and AND4 (N2164, N2136, N1349, N1685, N2145);
xor XOR2 (N2165, N2163, N331);
or OR2 (N2166, N2161, N1362);
nand NAND3 (N2167, N2144, N334, N1772);
xor XOR2 (N2168, N2166, N2027);
or OR2 (N2169, N2165, N779);
nand NAND4 (N2170, N2156, N2101, N1692, N1882);
xor XOR2 (N2171, N2157, N62);
or OR4 (N2172, N2158, N369, N8, N433);
or OR4 (N2173, N2171, N1500, N1048, N381);
not NOT1 (N2174, N2164);
buf BUF1 (N2175, N2174);
buf BUF1 (N2176, N2154);
nor NOR2 (N2177, N2170, N108);
xor XOR2 (N2178, N2176, N353);
not NOT1 (N2179, N2167);
buf BUF1 (N2180, N2177);
or OR2 (N2181, N2180, N738);
buf BUF1 (N2182, N2159);
xor XOR2 (N2183, N2181, N172);
nor NOR3 (N2184, N2183, N1358, N519);
or OR4 (N2185, N2173, N335, N1132, N1937);
or OR4 (N2186, N2175, N1598, N1482, N1125);
not NOT1 (N2187, N2182);
xor XOR2 (N2188, N2178, N611);
or OR2 (N2189, N2186, N1395);
xor XOR2 (N2190, N2168, N1151);
and AND2 (N2191, N2189, N1830);
xor XOR2 (N2192, N2185, N609);
nor NOR2 (N2193, N2184, N235);
or OR3 (N2194, N2162, N31, N1031);
and AND4 (N2195, N2188, N1420, N1259, N1980);
nor NOR4 (N2196, N2172, N1286, N1047, N937);
xor XOR2 (N2197, N2190, N930);
and AND2 (N2198, N2196, N1193);
buf BUF1 (N2199, N2194);
and AND4 (N2200, N2191, N1196, N1070, N1819);
buf BUF1 (N2201, N2179);
not NOT1 (N2202, N2195);
or OR4 (N2203, N2202, N972, N1557, N146);
not NOT1 (N2204, N2187);
not NOT1 (N2205, N2192);
nor NOR3 (N2206, N2201, N1421, N536);
xor XOR2 (N2207, N2198, N1042);
buf BUF1 (N2208, N2193);
xor XOR2 (N2209, N2197, N299);
buf BUF1 (N2210, N2205);
nand NAND3 (N2211, N2208, N1993, N1598);
nor NOR4 (N2212, N2207, N923, N125, N88);
nand NAND4 (N2213, N2211, N546, N879, N2064);
and AND3 (N2214, N2209, N1088, N1263);
nor NOR3 (N2215, N2213, N53, N195);
buf BUF1 (N2216, N2169);
nand NAND2 (N2217, N2206, N1130);
nand NAND4 (N2218, N2215, N1425, N916, N1336);
nand NAND4 (N2219, N2199, N613, N2008, N1033);
and AND4 (N2220, N2204, N1720, N343, N1912);
xor XOR2 (N2221, N2200, N205);
or OR4 (N2222, N2210, N2152, N380, N1258);
xor XOR2 (N2223, N2214, N532);
nor NOR3 (N2224, N2203, N561, N1997);
and AND2 (N2225, N2220, N2054);
nand NAND3 (N2226, N2218, N257, N2007);
not NOT1 (N2227, N2219);
buf BUF1 (N2228, N2216);
buf BUF1 (N2229, N2212);
and AND4 (N2230, N2217, N1996, N1138, N2157);
xor XOR2 (N2231, N2230, N1715);
and AND2 (N2232, N2226, N312);
buf BUF1 (N2233, N2222);
xor XOR2 (N2234, N2225, N47);
xor XOR2 (N2235, N2234, N1152);
not NOT1 (N2236, N2235);
xor XOR2 (N2237, N2236, N101);
or OR3 (N2238, N2224, N2037, N2084);
or OR3 (N2239, N2237, N250, N261);
nand NAND3 (N2240, N2229, N1665, N478);
xor XOR2 (N2241, N2227, N1364);
xor XOR2 (N2242, N2241, N1222);
buf BUF1 (N2243, N2223);
nand NAND2 (N2244, N2232, N1401);
or OR4 (N2245, N2233, N246, N1849, N616);
not NOT1 (N2246, N2231);
buf BUF1 (N2247, N2221);
not NOT1 (N2248, N2243);
buf BUF1 (N2249, N2247);
nand NAND4 (N2250, N2245, N1751, N982, N1278);
or OR2 (N2251, N2250, N659);
nor NOR4 (N2252, N2238, N364, N1050, N1536);
not NOT1 (N2253, N2251);
buf BUF1 (N2254, N2242);
nand NAND4 (N2255, N2248, N1882, N265, N1361);
nand NAND4 (N2256, N2244, N407, N1058, N936);
nand NAND2 (N2257, N2246, N1879);
buf BUF1 (N2258, N2253);
xor XOR2 (N2259, N2258, N836);
or OR2 (N2260, N2256, N689);
or OR4 (N2261, N2260, N352, N31, N929);
nor NOR2 (N2262, N2249, N1784);
not NOT1 (N2263, N2252);
not NOT1 (N2264, N2254);
buf BUF1 (N2265, N2257);
buf BUF1 (N2266, N2259);
not NOT1 (N2267, N2261);
nor NOR3 (N2268, N2266, N107, N1802);
not NOT1 (N2269, N2255);
buf BUF1 (N2270, N2269);
nor NOR3 (N2271, N2240, N1673, N666);
and AND2 (N2272, N2267, N582);
and AND2 (N2273, N2228, N2122);
nand NAND2 (N2274, N2262, N1760);
nand NAND3 (N2275, N2263, N457, N2249);
and AND3 (N2276, N2239, N1543, N1315);
buf BUF1 (N2277, N2274);
and AND4 (N2278, N2276, N8, N2134, N1436);
nand NAND2 (N2279, N2277, N349);
nand NAND4 (N2280, N2268, N563, N1200, N1965);
not NOT1 (N2281, N2272);
and AND3 (N2282, N2280, N986, N1631);
nor NOR4 (N2283, N2273, N1436, N556, N2255);
nand NAND3 (N2284, N2279, N2065, N2047);
and AND2 (N2285, N2271, N233);
or OR2 (N2286, N2264, N2101);
or OR2 (N2287, N2275, N580);
or OR2 (N2288, N2281, N2220);
and AND2 (N2289, N2265, N2219);
xor XOR2 (N2290, N2284, N187);
nand NAND2 (N2291, N2288, N1172);
buf BUF1 (N2292, N2282);
nor NOR4 (N2293, N2283, N2081, N1908, N427);
xor XOR2 (N2294, N2270, N1739);
buf BUF1 (N2295, N2286);
xor XOR2 (N2296, N2287, N1834);
buf BUF1 (N2297, N2285);
and AND3 (N2298, N2290, N1578, N249);
not NOT1 (N2299, N2295);
or OR4 (N2300, N2299, N1351, N1913, N488);
nor NOR3 (N2301, N2278, N1867, N1218);
and AND2 (N2302, N2291, N452);
not NOT1 (N2303, N2300);
buf BUF1 (N2304, N2302);
nand NAND2 (N2305, N2303, N227);
nor NOR4 (N2306, N2296, N1033, N840, N269);
xor XOR2 (N2307, N2298, N1113);
or OR3 (N2308, N2297, N1287, N619);
and AND3 (N2309, N2306, N530, N2093);
or OR2 (N2310, N2292, N828);
buf BUF1 (N2311, N2304);
and AND4 (N2312, N2308, N1112, N149, N360);
buf BUF1 (N2313, N2307);
nor NOR4 (N2314, N2293, N1160, N2102, N1016);
nor NOR4 (N2315, N2305, N294, N1010, N1205);
nand NAND3 (N2316, N2314, N2158, N1241);
and AND2 (N2317, N2312, N1909);
and AND3 (N2318, N2294, N382, N1791);
not NOT1 (N2319, N2301);
nor NOR3 (N2320, N2311, N1971, N1591);
not NOT1 (N2321, N2309);
buf BUF1 (N2322, N2313);
not NOT1 (N2323, N2317);
xor XOR2 (N2324, N2323, N1665);
buf BUF1 (N2325, N2322);
not NOT1 (N2326, N2320);
and AND3 (N2327, N2321, N843, N1401);
not NOT1 (N2328, N2310);
and AND4 (N2329, N2289, N579, N906, N1176);
xor XOR2 (N2330, N2324, N1561);
nand NAND2 (N2331, N2316, N2107);
xor XOR2 (N2332, N2328, N644);
not NOT1 (N2333, N2326);
buf BUF1 (N2334, N2327);
nor NOR3 (N2335, N2319, N217, N1412);
or OR2 (N2336, N2331, N746);
nand NAND4 (N2337, N2334, N614, N1406, N1171);
not NOT1 (N2338, N2336);
or OR3 (N2339, N2315, N1842, N1633);
or OR2 (N2340, N2337, N63);
or OR2 (N2341, N2325, N694);
buf BUF1 (N2342, N2340);
xor XOR2 (N2343, N2338, N453);
nor NOR4 (N2344, N2330, N660, N854, N454);
and AND4 (N2345, N2335, N1642, N1785, N690);
and AND4 (N2346, N2339, N1776, N1479, N1265);
not NOT1 (N2347, N2318);
or OR2 (N2348, N2345, N2107);
nand NAND2 (N2349, N2332, N183);
and AND3 (N2350, N2347, N514, N2292);
nor NOR2 (N2351, N2349, N1840);
buf BUF1 (N2352, N2344);
and AND2 (N2353, N2342, N724);
nand NAND2 (N2354, N2333, N179);
xor XOR2 (N2355, N2343, N1371);
or OR4 (N2356, N2354, N1442, N1508, N801);
not NOT1 (N2357, N2341);
nand NAND3 (N2358, N2357, N782, N1762);
not NOT1 (N2359, N2355);
buf BUF1 (N2360, N2353);
and AND3 (N2361, N2356, N1516, N704);
or OR4 (N2362, N2348, N601, N1583, N1800);
and AND4 (N2363, N2329, N681, N820, N541);
xor XOR2 (N2364, N2351, N1772);
nand NAND2 (N2365, N2363, N2317);
or OR4 (N2366, N2346, N1343, N318, N918);
buf BUF1 (N2367, N2365);
buf BUF1 (N2368, N2364);
nand NAND4 (N2369, N2350, N827, N423, N1932);
and AND4 (N2370, N2358, N690, N962, N409);
not NOT1 (N2371, N2362);
not NOT1 (N2372, N2359);
not NOT1 (N2373, N2361);
buf BUF1 (N2374, N2372);
buf BUF1 (N2375, N2367);
xor XOR2 (N2376, N2360, N709);
not NOT1 (N2377, N2375);
not NOT1 (N2378, N2368);
buf BUF1 (N2379, N2371);
or OR3 (N2380, N2376, N329, N1475);
nor NOR4 (N2381, N2369, N1784, N1447, N450);
and AND4 (N2382, N2381, N2046, N862, N435);
nand NAND3 (N2383, N2352, N187, N1504);
and AND3 (N2384, N2380, N1329, N1049);
xor XOR2 (N2385, N2384, N416);
xor XOR2 (N2386, N2383, N1939);
buf BUF1 (N2387, N2378);
xor XOR2 (N2388, N2387, N2358);
or OR2 (N2389, N2382, N332);
nand NAND2 (N2390, N2370, N1835);
buf BUF1 (N2391, N2377);
not NOT1 (N2392, N2385);
not NOT1 (N2393, N2386);
buf BUF1 (N2394, N2374);
nor NOR2 (N2395, N2389, N1973);
not NOT1 (N2396, N2392);
nor NOR4 (N2397, N2391, N1605, N63, N1181);
nand NAND3 (N2398, N2366, N723, N2085);
xor XOR2 (N2399, N2390, N277);
nor NOR3 (N2400, N2373, N160, N400);
nor NOR3 (N2401, N2397, N483, N1662);
buf BUF1 (N2402, N2401);
buf BUF1 (N2403, N2379);
or OR3 (N2404, N2394, N2042, N1284);
xor XOR2 (N2405, N2404, N508);
buf BUF1 (N2406, N2395);
nand NAND2 (N2407, N2398, N117);
nand NAND3 (N2408, N2388, N1907, N1768);
and AND4 (N2409, N2403, N1541, N1223, N360);
not NOT1 (N2410, N2396);
xor XOR2 (N2411, N2400, N1106);
nand NAND3 (N2412, N2406, N393, N2157);
xor XOR2 (N2413, N2409, N311);
buf BUF1 (N2414, N2399);
nand NAND3 (N2415, N2407, N1, N723);
nor NOR3 (N2416, N2414, N1209, N986);
and AND2 (N2417, N2412, N2381);
xor XOR2 (N2418, N2405, N1449);
not NOT1 (N2419, N2413);
nor NOR4 (N2420, N2411, N2042, N972, N355);
nand NAND2 (N2421, N2418, N1316);
nand NAND3 (N2422, N2419, N1705, N2158);
and AND4 (N2423, N2393, N505, N1656, N1505);
xor XOR2 (N2424, N2402, N1675);
nand NAND4 (N2425, N2416, N616, N310, N1411);
nand NAND3 (N2426, N2417, N1379, N206);
or OR3 (N2427, N2424, N74, N2143);
not NOT1 (N2428, N2425);
or OR3 (N2429, N2427, N415, N2193);
or OR4 (N2430, N2415, N863, N923, N2295);
nor NOR4 (N2431, N2428, N2175, N2128, N2203);
xor XOR2 (N2432, N2431, N1519);
not NOT1 (N2433, N2410);
or OR4 (N2434, N2430, N1337, N1460, N332);
not NOT1 (N2435, N2426);
not NOT1 (N2436, N2433);
nand NAND2 (N2437, N2423, N552);
not NOT1 (N2438, N2432);
xor XOR2 (N2439, N2436, N197);
buf BUF1 (N2440, N2434);
not NOT1 (N2441, N2420);
xor XOR2 (N2442, N2408, N349);
buf BUF1 (N2443, N2439);
nor NOR2 (N2444, N2422, N566);
not NOT1 (N2445, N2441);
buf BUF1 (N2446, N2442);
xor XOR2 (N2447, N2440, N1639);
or OR4 (N2448, N2437, N2154, N606, N542);
xor XOR2 (N2449, N2445, N39);
buf BUF1 (N2450, N2421);
nor NOR4 (N2451, N2446, N390, N2104, N2061);
and AND4 (N2452, N2447, N2313, N1396, N651);
nor NOR4 (N2453, N2429, N1808, N1291, N779);
and AND3 (N2454, N2449, N2061, N1144);
xor XOR2 (N2455, N2443, N2169);
and AND2 (N2456, N2454, N1741);
or OR4 (N2457, N2444, N360, N2454, N1911);
nand NAND4 (N2458, N2448, N1746, N1175, N1544);
and AND3 (N2459, N2435, N437, N2225);
xor XOR2 (N2460, N2455, N794);
xor XOR2 (N2461, N2456, N21);
nand NAND4 (N2462, N2458, N2010, N674, N121);
or OR2 (N2463, N2438, N868);
and AND2 (N2464, N2451, N731);
not NOT1 (N2465, N2464);
nand NAND2 (N2466, N2463, N687);
not NOT1 (N2467, N2452);
xor XOR2 (N2468, N2453, N835);
and AND2 (N2469, N2457, N391);
not NOT1 (N2470, N2462);
or OR2 (N2471, N2450, N255);
and AND4 (N2472, N2460, N607, N394, N1073);
buf BUF1 (N2473, N2468);
or OR3 (N2474, N2469, N2459, N1586);
xor XOR2 (N2475, N2066, N1688);
or OR4 (N2476, N2465, N269, N225, N1441);
buf BUF1 (N2477, N2474);
or OR4 (N2478, N2461, N44, N767, N119);
or OR3 (N2479, N2473, N2294, N1196);
xor XOR2 (N2480, N2476, N2386);
and AND2 (N2481, N2471, N1060);
and AND4 (N2482, N2472, N1244, N2118, N1122);
or OR2 (N2483, N2481, N493);
and AND4 (N2484, N2466, N227, N1452, N1838);
or OR4 (N2485, N2482, N1518, N1954, N613);
xor XOR2 (N2486, N2467, N1802);
xor XOR2 (N2487, N2484, N2415);
nor NOR4 (N2488, N2475, N979, N230, N1647);
or OR2 (N2489, N2488, N1870);
or OR4 (N2490, N2477, N2032, N923, N1163);
buf BUF1 (N2491, N2470);
xor XOR2 (N2492, N2480, N2154);
nand NAND3 (N2493, N2489, N2081, N202);
buf BUF1 (N2494, N2493);
xor XOR2 (N2495, N2494, N1498);
buf BUF1 (N2496, N2490);
nand NAND3 (N2497, N2486, N200, N2357);
nand NAND3 (N2498, N2485, N2110, N504);
or OR4 (N2499, N2496, N2126, N1895, N1274);
or OR2 (N2500, N2497, N2416);
xor XOR2 (N2501, N2499, N1722);
buf BUF1 (N2502, N2491);
or OR3 (N2503, N2479, N853, N264);
nor NOR4 (N2504, N2495, N2189, N8, N1014);
not NOT1 (N2505, N2498);
and AND2 (N2506, N2502, N922);
or OR3 (N2507, N2492, N1252, N914);
xor XOR2 (N2508, N2501, N853);
xor XOR2 (N2509, N2506, N103);
not NOT1 (N2510, N2483);
nor NOR3 (N2511, N2504, N1710, N148);
nand NAND2 (N2512, N2508, N1039);
xor XOR2 (N2513, N2500, N1386);
nor NOR2 (N2514, N2510, N400);
not NOT1 (N2515, N2509);
buf BUF1 (N2516, N2478);
not NOT1 (N2517, N2515);
xor XOR2 (N2518, N2516, N1087);
buf BUF1 (N2519, N2511);
xor XOR2 (N2520, N2487, N1458);
or OR3 (N2521, N2512, N282, N2093);
buf BUF1 (N2522, N2519);
nor NOR3 (N2523, N2518, N957, N412);
not NOT1 (N2524, N2520);
nand NAND4 (N2525, N2517, N1711, N1528, N329);
buf BUF1 (N2526, N2522);
not NOT1 (N2527, N2525);
xor XOR2 (N2528, N2521, N1977);
or OR2 (N2529, N2526, N350);
xor XOR2 (N2530, N2505, N548);
and AND3 (N2531, N2528, N1275, N1193);
xor XOR2 (N2532, N2527, N997);
and AND3 (N2533, N2529, N2317, N724);
nand NAND3 (N2534, N2532, N2514, N1355);
nor NOR4 (N2535, N1788, N1917, N411, N2457);
nor NOR3 (N2536, N2524, N322, N1598);
nor NOR3 (N2537, N2535, N257, N767);
nand NAND4 (N2538, N2537, N986, N1936, N2199);
nand NAND3 (N2539, N2503, N2248, N1037);
xor XOR2 (N2540, N2536, N1347);
nand NAND2 (N2541, N2531, N2103);
nand NAND4 (N2542, N2539, N10, N1860, N1071);
or OR4 (N2543, N2530, N1047, N402, N1239);
xor XOR2 (N2544, N2513, N744);
and AND3 (N2545, N2542, N1013, N2022);
buf BUF1 (N2546, N2507);
or OR4 (N2547, N2523, N926, N738, N2098);
not NOT1 (N2548, N2538);
and AND3 (N2549, N2547, N229, N1809);
xor XOR2 (N2550, N2541, N794);
buf BUF1 (N2551, N2548);
or OR3 (N2552, N2546, N1389, N851);
or OR4 (N2553, N2540, N1559, N237, N2518);
xor XOR2 (N2554, N2549, N1400);
xor XOR2 (N2555, N2553, N1363);
buf BUF1 (N2556, N2551);
nor NOR4 (N2557, N2550, N1319, N1081, N2416);
xor XOR2 (N2558, N2543, N2347);
or OR2 (N2559, N2557, N667);
nor NOR4 (N2560, N2555, N1742, N373, N1297);
and AND4 (N2561, N2552, N2103, N166, N1645);
buf BUF1 (N2562, N2545);
buf BUF1 (N2563, N2533);
and AND4 (N2564, N2544, N181, N367, N1579);
xor XOR2 (N2565, N2561, N2114);
nor NOR2 (N2566, N2559, N136);
and AND3 (N2567, N2566, N859, N1379);
nand NAND4 (N2568, N2556, N794, N982, N344);
and AND2 (N2569, N2564, N564);
and AND3 (N2570, N2569, N2038, N1880);
xor XOR2 (N2571, N2558, N2531);
and AND4 (N2572, N2568, N1908, N1305, N2185);
and AND2 (N2573, N2565, N922);
or OR4 (N2574, N2572, N758, N102, N1082);
nand NAND4 (N2575, N2571, N342, N607, N848);
and AND2 (N2576, N2554, N924);
or OR2 (N2577, N2570, N1072);
nor NOR2 (N2578, N2562, N569);
and AND4 (N2579, N2560, N978, N1311, N1397);
nand NAND2 (N2580, N2534, N2292);
not NOT1 (N2581, N2580);
nand NAND4 (N2582, N2575, N2440, N1470, N183);
xor XOR2 (N2583, N2573, N1325);
not NOT1 (N2584, N2583);
and AND4 (N2585, N2576, N2429, N881, N309);
nand NAND3 (N2586, N2585, N2227, N1930);
xor XOR2 (N2587, N2578, N1506);
not NOT1 (N2588, N2577);
buf BUF1 (N2589, N2588);
nand NAND2 (N2590, N2567, N1229);
buf BUF1 (N2591, N2579);
not NOT1 (N2592, N2563);
xor XOR2 (N2593, N2582, N1327);
nor NOR4 (N2594, N2574, N2355, N1214, N528);
and AND4 (N2595, N2591, N2047, N836, N2230);
or OR4 (N2596, N2595, N2009, N1011, N1037);
xor XOR2 (N2597, N2593, N120);
and AND4 (N2598, N2597, N500, N1045, N1049);
and AND4 (N2599, N2592, N641, N931, N2234);
buf BUF1 (N2600, N2587);
or OR4 (N2601, N2590, N757, N43, N1337);
xor XOR2 (N2602, N2598, N2166);
xor XOR2 (N2603, N2599, N483);
buf BUF1 (N2604, N2601);
nand NAND2 (N2605, N2600, N1433);
nand NAND2 (N2606, N2594, N2136);
nor NOR4 (N2607, N2603, N1184, N1887, N1694);
xor XOR2 (N2608, N2604, N1746);
not NOT1 (N2609, N2605);
and AND3 (N2610, N2586, N767, N952);
nand NAND2 (N2611, N2607, N4);
buf BUF1 (N2612, N2608);
not NOT1 (N2613, N2606);
xor XOR2 (N2614, N2581, N732);
buf BUF1 (N2615, N2584);
not NOT1 (N2616, N2589);
xor XOR2 (N2617, N2612, N1443);
xor XOR2 (N2618, N2609, N120);
buf BUF1 (N2619, N2596);
xor XOR2 (N2620, N2613, N704);
or OR2 (N2621, N2611, N157);
and AND2 (N2622, N2619, N2087);
nor NOR4 (N2623, N2614, N960, N1896, N774);
or OR3 (N2624, N2622, N817, N1633);
nand NAND2 (N2625, N2621, N1102);
xor XOR2 (N2626, N2617, N2440);
nand NAND2 (N2627, N2623, N944);
xor XOR2 (N2628, N2602, N1582);
xor XOR2 (N2629, N2610, N2026);
or OR3 (N2630, N2629, N1822, N1525);
xor XOR2 (N2631, N2616, N2365);
not NOT1 (N2632, N2615);
nor NOR4 (N2633, N2632, N318, N2441, N1134);
or OR3 (N2634, N2620, N998, N659);
xor XOR2 (N2635, N2627, N1277);
nor NOR4 (N2636, N2630, N1982, N2541, N1485);
and AND3 (N2637, N2628, N2461, N1905);
buf BUF1 (N2638, N2624);
nor NOR3 (N2639, N2631, N320, N1939);
xor XOR2 (N2640, N2625, N1344);
and AND4 (N2641, N2618, N164, N2484, N1760);
not NOT1 (N2642, N2639);
or OR4 (N2643, N2635, N830, N2116, N1477);
nor NOR4 (N2644, N2633, N1097, N1228, N24);
nor NOR2 (N2645, N2642, N1065);
and AND3 (N2646, N2644, N2380, N1804);
xor XOR2 (N2647, N2641, N446);
xor XOR2 (N2648, N2645, N1407);
not NOT1 (N2649, N2648);
buf BUF1 (N2650, N2638);
nor NOR2 (N2651, N2647, N1870);
nor NOR4 (N2652, N2646, N700, N352, N698);
not NOT1 (N2653, N2626);
or OR3 (N2654, N2652, N1562, N2169);
not NOT1 (N2655, N2637);
xor XOR2 (N2656, N2649, N1641);
nand NAND4 (N2657, N2640, N1182, N1360, N1863);
buf BUF1 (N2658, N2651);
or OR3 (N2659, N2656, N1024, N540);
nand NAND2 (N2660, N2659, N1087);
and AND3 (N2661, N2636, N1634, N661);
xor XOR2 (N2662, N2657, N932);
nor NOR3 (N2663, N2655, N693, N1030);
nand NAND3 (N2664, N2663, N1580, N1938);
not NOT1 (N2665, N2661);
xor XOR2 (N2666, N2664, N108);
or OR4 (N2667, N2665, N1967, N921, N1721);
xor XOR2 (N2668, N2667, N980);
nor NOR2 (N2669, N2654, N2296);
buf BUF1 (N2670, N2643);
nand NAND4 (N2671, N2668, N1084, N2492, N527);
not NOT1 (N2672, N2650);
and AND3 (N2673, N2658, N582, N674);
nand NAND2 (N2674, N2671, N372);
buf BUF1 (N2675, N2662);
nor NOR4 (N2676, N2653, N1766, N2187, N2545);
buf BUF1 (N2677, N2675);
not NOT1 (N2678, N2677);
nor NOR2 (N2679, N2634, N734);
nand NAND3 (N2680, N2678, N2156, N2018);
nor NOR3 (N2681, N2669, N1757, N1767);
or OR4 (N2682, N2670, N1486, N36, N1379);
not NOT1 (N2683, N2681);
not NOT1 (N2684, N2672);
buf BUF1 (N2685, N2679);
nand NAND3 (N2686, N2676, N535, N1580);
or OR2 (N2687, N2682, N1979);
nand NAND4 (N2688, N2673, N577, N796, N1420);
not NOT1 (N2689, N2660);
nand NAND2 (N2690, N2687, N1147);
buf BUF1 (N2691, N2688);
or OR2 (N2692, N2686, N1713);
or OR4 (N2693, N2674, N2170, N662, N672);
buf BUF1 (N2694, N2691);
and AND3 (N2695, N2692, N503, N1635);
xor XOR2 (N2696, N2689, N2099);
or OR4 (N2697, N2684, N2492, N1363, N1059);
and AND4 (N2698, N2697, N1448, N1691, N2403);
or OR2 (N2699, N2693, N1152);
or OR3 (N2700, N2698, N575, N28);
buf BUF1 (N2701, N2696);
buf BUF1 (N2702, N2690);
not NOT1 (N2703, N2699);
not NOT1 (N2704, N2685);
xor XOR2 (N2705, N2680, N1637);
nand NAND4 (N2706, N2700, N900, N1177, N2165);
buf BUF1 (N2707, N2695);
nor NOR3 (N2708, N2705, N627, N998);
buf BUF1 (N2709, N2704);
nand NAND4 (N2710, N2702, N2282, N863, N2541);
nor NOR3 (N2711, N2666, N2007, N695);
and AND3 (N2712, N2701, N657, N1130);
not NOT1 (N2713, N2683);
or OR3 (N2714, N2706, N2294, N829);
xor XOR2 (N2715, N2712, N2014);
buf BUF1 (N2716, N2703);
and AND3 (N2717, N2694, N1717, N274);
xor XOR2 (N2718, N2711, N1338);
nand NAND3 (N2719, N2714, N759, N1189);
and AND3 (N2720, N2717, N2308, N1715);
or OR3 (N2721, N2707, N2438, N2491);
nor NOR2 (N2722, N2708, N1289);
and AND4 (N2723, N2718, N1241, N2634, N60);
xor XOR2 (N2724, N2720, N2681);
nor NOR4 (N2725, N2722, N1271, N923, N1303);
buf BUF1 (N2726, N2710);
and AND4 (N2727, N2719, N1956, N485, N1857);
not NOT1 (N2728, N2721);
buf BUF1 (N2729, N2726);
not NOT1 (N2730, N2724);
xor XOR2 (N2731, N2730, N1347);
or OR4 (N2732, N2723, N622, N249, N1090);
buf BUF1 (N2733, N2732);
buf BUF1 (N2734, N2731);
nor NOR4 (N2735, N2729, N1684, N2555, N75);
or OR2 (N2736, N2716, N911);
or OR3 (N2737, N2713, N647, N858);
nand NAND2 (N2738, N2735, N1580);
and AND4 (N2739, N2736, N1314, N1634, N2600);
xor XOR2 (N2740, N2733, N1325);
nand NAND2 (N2741, N2727, N1188);
xor XOR2 (N2742, N2739, N1602);
nand NAND2 (N2743, N2715, N1916);
buf BUF1 (N2744, N2738);
not NOT1 (N2745, N2734);
or OR3 (N2746, N2745, N964, N1873);
nor NOR2 (N2747, N2737, N1348);
buf BUF1 (N2748, N2744);
nor NOR4 (N2749, N2746, N94, N1650, N2093);
not NOT1 (N2750, N2725);
nor NOR2 (N2751, N2750, N46);
xor XOR2 (N2752, N2741, N1093);
and AND2 (N2753, N2747, N714);
buf BUF1 (N2754, N2751);
nor NOR2 (N2755, N2743, N870);
xor XOR2 (N2756, N2754, N676);
xor XOR2 (N2757, N2752, N1534);
nor NOR4 (N2758, N2742, N2256, N238, N1429);
not NOT1 (N2759, N2753);
not NOT1 (N2760, N2759);
or OR3 (N2761, N2728, N1840, N232);
or OR2 (N2762, N2709, N121);
not NOT1 (N2763, N2762);
xor XOR2 (N2764, N2740, N1003);
xor XOR2 (N2765, N2764, N2429);
nor NOR4 (N2766, N2760, N2219, N1526, N1394);
and AND4 (N2767, N2766, N2689, N1012, N1018);
nor NOR4 (N2768, N2755, N1999, N962, N836);
xor XOR2 (N2769, N2763, N2152);
and AND4 (N2770, N2767, N693, N43, N2692);
or OR4 (N2771, N2769, N1350, N2305, N2662);
buf BUF1 (N2772, N2748);
nor NOR4 (N2773, N2771, N1272, N2135, N557);
nor NOR3 (N2774, N2765, N2222, N873);
nand NAND2 (N2775, N2768, N1660);
xor XOR2 (N2776, N2758, N154);
not NOT1 (N2777, N2775);
or OR2 (N2778, N2773, N2674);
or OR3 (N2779, N2776, N421, N792);
not NOT1 (N2780, N2757);
nand NAND3 (N2781, N2756, N1950, N1653);
and AND3 (N2782, N2774, N85, N1840);
nor NOR4 (N2783, N2782, N1908, N2177, N621);
not NOT1 (N2784, N2779);
buf BUF1 (N2785, N2770);
nand NAND3 (N2786, N2784, N1690, N2268);
xor XOR2 (N2787, N2780, N509);
or OR4 (N2788, N2786, N1051, N1054, N142);
nand NAND4 (N2789, N2772, N1072, N2186, N1459);
xor XOR2 (N2790, N2789, N1964);
xor XOR2 (N2791, N2777, N757);
and AND4 (N2792, N2778, N1043, N1520, N786);
and AND3 (N2793, N2783, N2743, N88);
and AND2 (N2794, N2793, N2362);
nor NOR2 (N2795, N2761, N1074);
nand NAND4 (N2796, N2790, N2133, N648, N1181);
nand NAND2 (N2797, N2794, N1483);
and AND4 (N2798, N2795, N963, N359, N1484);
or OR3 (N2799, N2787, N1435, N381);
nor NOR4 (N2800, N2781, N1696, N2381, N1541);
nor NOR3 (N2801, N2798, N1098, N1421);
and AND2 (N2802, N2788, N191);
buf BUF1 (N2803, N2797);
and AND4 (N2804, N2802, N2183, N2681, N1798);
nand NAND2 (N2805, N2792, N2340);
or OR3 (N2806, N2803, N1537, N765);
nor NOR4 (N2807, N2806, N1268, N1027, N656);
or OR4 (N2808, N2804, N1172, N1574, N355);
and AND2 (N2809, N2800, N221);
xor XOR2 (N2810, N2796, N2748);
buf BUF1 (N2811, N2805);
nand NAND3 (N2812, N2785, N112, N141);
not NOT1 (N2813, N2809);
xor XOR2 (N2814, N2799, N2763);
xor XOR2 (N2815, N2811, N2685);
and AND3 (N2816, N2791, N1310, N20);
xor XOR2 (N2817, N2815, N2269);
xor XOR2 (N2818, N2807, N2018);
not NOT1 (N2819, N2810);
or OR4 (N2820, N2749, N1380, N2062, N1791);
and AND2 (N2821, N2814, N829);
or OR3 (N2822, N2818, N2041, N2262);
not NOT1 (N2823, N2813);
buf BUF1 (N2824, N2822);
xor XOR2 (N2825, N2808, N800);
and AND4 (N2826, N2820, N2749, N1455, N695);
not NOT1 (N2827, N2823);
nor NOR2 (N2828, N2801, N1419);
and AND4 (N2829, N2827, N2646, N1594, N2366);
buf BUF1 (N2830, N2817);
or OR3 (N2831, N2819, N2019, N913);
nor NOR3 (N2832, N2824, N1837, N236);
not NOT1 (N2833, N2828);
or OR4 (N2834, N2816, N683, N2241, N1032);
nand NAND3 (N2835, N2821, N864, N1646);
or OR3 (N2836, N2833, N1178, N2649);
xor XOR2 (N2837, N2832, N705);
buf BUF1 (N2838, N2837);
not NOT1 (N2839, N2838);
and AND2 (N2840, N2829, N1993);
buf BUF1 (N2841, N2826);
nand NAND3 (N2842, N2841, N1958, N2774);
nand NAND4 (N2843, N2836, N355, N2017, N596);
buf BUF1 (N2844, N2840);
and AND2 (N2845, N2844, N1242);
xor XOR2 (N2846, N2843, N2162);
buf BUF1 (N2847, N2830);
nand NAND3 (N2848, N2845, N535, N1687);
buf BUF1 (N2849, N2834);
xor XOR2 (N2850, N2812, N2497);
nor NOR4 (N2851, N2839, N1347, N1751, N1245);
nor NOR2 (N2852, N2850, N296);
nor NOR4 (N2853, N2825, N230, N1706, N471);
buf BUF1 (N2854, N2835);
buf BUF1 (N2855, N2853);
not NOT1 (N2856, N2851);
xor XOR2 (N2857, N2847, N201);
xor XOR2 (N2858, N2846, N1539);
or OR3 (N2859, N2848, N2348, N899);
buf BUF1 (N2860, N2854);
buf BUF1 (N2861, N2857);
nor NOR2 (N2862, N2852, N2333);
or OR4 (N2863, N2861, N1915, N1030, N1241);
not NOT1 (N2864, N2862);
and AND2 (N2865, N2858, N2000);
xor XOR2 (N2866, N2863, N2183);
nand NAND4 (N2867, N2855, N204, N2522, N26);
and AND3 (N2868, N2864, N1157, N2470);
not NOT1 (N2869, N2842);
nor NOR4 (N2870, N2856, N945, N2536, N2664);
nor NOR3 (N2871, N2867, N1511, N2561);
nor NOR4 (N2872, N2870, N1550, N1493, N399);
and AND4 (N2873, N2865, N1508, N1410, N503);
xor XOR2 (N2874, N2873, N2424);
xor XOR2 (N2875, N2868, N1303);
xor XOR2 (N2876, N2859, N366);
nand NAND3 (N2877, N2872, N2622, N2819);
and AND4 (N2878, N2866, N2326, N1652, N500);
and AND4 (N2879, N2871, N2470, N1540, N2133);
nor NOR2 (N2880, N2879, N2420);
nand NAND2 (N2881, N2880, N870);
nor NOR4 (N2882, N2877, N1734, N1129, N2501);
xor XOR2 (N2883, N2869, N1264);
buf BUF1 (N2884, N2876);
buf BUF1 (N2885, N2884);
nand NAND2 (N2886, N2831, N1743);
nand NAND3 (N2887, N2881, N2684, N1462);
nand NAND2 (N2888, N2860, N1591);
not NOT1 (N2889, N2883);
not NOT1 (N2890, N2889);
not NOT1 (N2891, N2890);
or OR4 (N2892, N2849, N2215, N448, N1143);
nor NOR3 (N2893, N2891, N2450, N1569);
nor NOR2 (N2894, N2874, N2103);
nand NAND2 (N2895, N2885, N51);
not NOT1 (N2896, N2882);
nand NAND4 (N2897, N2893, N1356, N10, N2681);
and AND2 (N2898, N2886, N2222);
and AND3 (N2899, N2875, N2121, N247);
xor XOR2 (N2900, N2898, N811);
not NOT1 (N2901, N2887);
xor XOR2 (N2902, N2897, N703);
nor NOR3 (N2903, N2878, N2830, N2728);
xor XOR2 (N2904, N2894, N1715);
not NOT1 (N2905, N2901);
or OR2 (N2906, N2892, N193);
xor XOR2 (N2907, N2899, N2644);
nand NAND3 (N2908, N2907, N1720, N591);
nor NOR4 (N2909, N2904, N1070, N1870, N1094);
nand NAND4 (N2910, N2906, N1276, N225, N785);
not NOT1 (N2911, N2888);
not NOT1 (N2912, N2895);
nand NAND2 (N2913, N2909, N109);
buf BUF1 (N2914, N2910);
and AND4 (N2915, N2896, N2708, N838, N810);
and AND2 (N2916, N2914, N1779);
nor NOR3 (N2917, N2912, N2554, N561);
and AND4 (N2918, N2915, N2549, N1069, N1011);
and AND4 (N2919, N2903, N1030, N865, N2514);
and AND4 (N2920, N2919, N326, N966, N1276);
buf BUF1 (N2921, N2920);
or OR4 (N2922, N2911, N1741, N820, N2800);
and AND3 (N2923, N2916, N1900, N1828);
nand NAND4 (N2924, N2900, N2417, N1601, N264);
nand NAND3 (N2925, N2918, N1085, N1981);
and AND2 (N2926, N2921, N120);
or OR3 (N2927, N2905, N1667, N68);
nor NOR3 (N2928, N2927, N2396, N1176);
nand NAND3 (N2929, N2926, N2699, N2273);
nor NOR3 (N2930, N2928, N1452, N797);
nand NAND4 (N2931, N2930, N1585, N2045, N2113);
xor XOR2 (N2932, N2923, N1450);
buf BUF1 (N2933, N2922);
nand NAND2 (N2934, N2931, N2915);
xor XOR2 (N2935, N2933, N1781);
not NOT1 (N2936, N2929);
not NOT1 (N2937, N2908);
nor NOR2 (N2938, N2917, N2810);
and AND4 (N2939, N2932, N2437, N2210, N914);
buf BUF1 (N2940, N2937);
buf BUF1 (N2941, N2925);
xor XOR2 (N2942, N2935, N2559);
and AND3 (N2943, N2924, N1947, N159);
or OR3 (N2944, N2941, N890, N1147);
nor NOR4 (N2945, N2939, N1584, N2546, N722);
nor NOR2 (N2946, N2945, N177);
buf BUF1 (N2947, N2944);
and AND4 (N2948, N2913, N160, N1055, N1678);
not NOT1 (N2949, N2948);
nand NAND2 (N2950, N2943, N1079);
nand NAND3 (N2951, N2946, N302, N113);
or OR3 (N2952, N2902, N51, N1973);
nor NOR3 (N2953, N2938, N1499, N43);
nor NOR4 (N2954, N2951, N1046, N2587, N192);
or OR3 (N2955, N2942, N569, N2739);
and AND3 (N2956, N2936, N1597, N1201);
xor XOR2 (N2957, N2950, N238);
and AND2 (N2958, N2955, N799);
nand NAND3 (N2959, N2953, N2086, N61);
nor NOR4 (N2960, N2949, N250, N2002, N542);
buf BUF1 (N2961, N2934);
and AND2 (N2962, N2954, N1487);
nand NAND2 (N2963, N2961, N1719);
xor XOR2 (N2964, N2957, N824);
xor XOR2 (N2965, N2962, N1509);
nor NOR2 (N2966, N2964, N1655);
nand NAND3 (N2967, N2966, N708, N536);
not NOT1 (N2968, N2940);
or OR3 (N2969, N2968, N2586, N81);
xor XOR2 (N2970, N2947, N648);
xor XOR2 (N2971, N2969, N515);
and AND3 (N2972, N2965, N2715, N1767);
and AND2 (N2973, N2960, N2925);
nor NOR2 (N2974, N2970, N2619);
nand NAND4 (N2975, N2952, N11, N2267, N1658);
or OR3 (N2976, N2956, N2053, N2528);
buf BUF1 (N2977, N2976);
nor NOR4 (N2978, N2967, N2613, N1573, N466);
not NOT1 (N2979, N2973);
not NOT1 (N2980, N2978);
not NOT1 (N2981, N2979);
nor NOR2 (N2982, N2972, N2021);
nor NOR4 (N2983, N2959, N1982, N703, N1967);
not NOT1 (N2984, N2982);
nand NAND4 (N2985, N2980, N1728, N1894, N811);
xor XOR2 (N2986, N2974, N388);
nor NOR3 (N2987, N2984, N2886, N1534);
xor XOR2 (N2988, N2958, N221);
buf BUF1 (N2989, N2971);
xor XOR2 (N2990, N2988, N824);
nand NAND4 (N2991, N2975, N1288, N2035, N678);
or OR3 (N2992, N2987, N1825, N1910);
xor XOR2 (N2993, N2985, N1460);
nand NAND3 (N2994, N2983, N1168, N2497);
nand NAND2 (N2995, N2990, N1390);
buf BUF1 (N2996, N2991);
nand NAND2 (N2997, N2995, N359);
nand NAND2 (N2998, N2997, N2950);
buf BUF1 (N2999, N2986);
nand NAND4 (N3000, N2992, N1167, N1544, N287);
nand NAND4 (N3001, N2981, N1623, N2453, N173);
buf BUF1 (N3002, N2977);
or OR4 (N3003, N3002, N2819, N253, N2576);
xor XOR2 (N3004, N2999, N2575);
nor NOR4 (N3005, N2993, N2087, N2159, N656);
nand NAND3 (N3006, N3003, N2489, N1522);
buf BUF1 (N3007, N3005);
and AND3 (N3008, N2989, N1765, N1801);
xor XOR2 (N3009, N2996, N2692);
nand NAND2 (N3010, N3008, N1945);
buf BUF1 (N3011, N3010);
not NOT1 (N3012, N3011);
buf BUF1 (N3013, N2998);
buf BUF1 (N3014, N3007);
buf BUF1 (N3015, N2963);
nor NOR3 (N3016, N3009, N1766, N1908);
xor XOR2 (N3017, N3001, N2243);
xor XOR2 (N3018, N2994, N900);
nand NAND3 (N3019, N3016, N1078, N465);
nand NAND4 (N3020, N3012, N1555, N2076, N2976);
buf BUF1 (N3021, N3017);
buf BUF1 (N3022, N3004);
nand NAND2 (N3023, N3022, N2906);
not NOT1 (N3024, N3020);
buf BUF1 (N3025, N3000);
nand NAND3 (N3026, N3006, N2595, N465);
nand NAND4 (N3027, N3021, N692, N2225, N592);
not NOT1 (N3028, N3024);
nor NOR2 (N3029, N3027, N472);
or OR3 (N3030, N3019, N592, N2466);
nand NAND2 (N3031, N3023, N819);
nand NAND2 (N3032, N3030, N2899);
nor NOR2 (N3033, N3031, N2706);
or OR4 (N3034, N3015, N770, N1055, N1899);
xor XOR2 (N3035, N3025, N2076);
nor NOR2 (N3036, N3034, N2526);
buf BUF1 (N3037, N3035);
nand NAND3 (N3038, N3036, N2977, N2650);
not NOT1 (N3039, N3033);
not NOT1 (N3040, N3018);
and AND3 (N3041, N3029, N131, N251);
nor NOR2 (N3042, N3013, N1030);
and AND2 (N3043, N3032, N1136);
and AND4 (N3044, N3043, N2011, N1871, N990);
and AND2 (N3045, N3042, N2900);
buf BUF1 (N3046, N3026);
not NOT1 (N3047, N3037);
nor NOR3 (N3048, N3014, N1070, N968);
xor XOR2 (N3049, N3044, N2061);
or OR2 (N3050, N3047, N2667);
or OR3 (N3051, N3039, N2607, N1436);
nand NAND3 (N3052, N3051, N1240, N756);
and AND3 (N3053, N3038, N2782, N1208);
xor XOR2 (N3054, N3046, N1540);
nand NAND3 (N3055, N3053, N104, N905);
nor NOR4 (N3056, N3045, N768, N649, N2903);
nor NOR4 (N3057, N3040, N1407, N1775, N467);
and AND3 (N3058, N3049, N1565, N2345);
buf BUF1 (N3059, N3052);
nand NAND2 (N3060, N3050, N2871);
not NOT1 (N3061, N3055);
or OR3 (N3062, N3041, N1991, N1528);
not NOT1 (N3063, N3059);
xor XOR2 (N3064, N3062, N493);
nor NOR2 (N3065, N3064, N2682);
or OR4 (N3066, N3057, N2902, N2504, N523);
nor NOR3 (N3067, N3058, N1350, N907);
or OR2 (N3068, N3056, N1198);
buf BUF1 (N3069, N3028);
nor NOR4 (N3070, N3065, N579, N1332, N2436);
nor NOR3 (N3071, N3054, N2358, N2341);
nand NAND2 (N3072, N3067, N2647);
xor XOR2 (N3073, N3066, N2984);
nand NAND2 (N3074, N3072, N26);
nor NOR2 (N3075, N3060, N510);
not NOT1 (N3076, N3071);
not NOT1 (N3077, N3074);
or OR2 (N3078, N3068, N1470);
not NOT1 (N3079, N3048);
nand NAND2 (N3080, N3078, N1894);
or OR4 (N3081, N3077, N1373, N1259, N94);
buf BUF1 (N3082, N3069);
nor NOR2 (N3083, N3075, N401);
nor NOR4 (N3084, N3081, N1332, N403, N234);
not NOT1 (N3085, N3080);
and AND2 (N3086, N3085, N371);
nor NOR3 (N3087, N3063, N2399, N535);
or OR4 (N3088, N3084, N993, N1892, N69);
xor XOR2 (N3089, N3087, N1333);
not NOT1 (N3090, N3088);
or OR3 (N3091, N3073, N2740, N1488);
or OR3 (N3092, N3061, N2991, N1224);
not NOT1 (N3093, N3086);
buf BUF1 (N3094, N3092);
nand NAND4 (N3095, N3082, N620, N2233, N951);
nor NOR2 (N3096, N3076, N1743);
or OR4 (N3097, N3079, N790, N758, N2858);
xor XOR2 (N3098, N3091, N3055);
not NOT1 (N3099, N3090);
not NOT1 (N3100, N3089);
buf BUF1 (N3101, N3100);
buf BUF1 (N3102, N3070);
not NOT1 (N3103, N3094);
xor XOR2 (N3104, N3083, N481);
nand NAND2 (N3105, N3093, N250);
nor NOR4 (N3106, N3102, N260, N2876, N1274);
nand NAND2 (N3107, N3098, N2884);
or OR4 (N3108, N3103, N897, N2271, N524);
nand NAND2 (N3109, N3108, N2560);
or OR3 (N3110, N3109, N1086, N575);
nand NAND2 (N3111, N3101, N1891);
nor NOR3 (N3112, N3104, N2513, N2179);
or OR4 (N3113, N3106, N2038, N1188, N2491);
nor NOR3 (N3114, N3111, N135, N2109);
nand NAND3 (N3115, N3097, N506, N1113);
nand NAND4 (N3116, N3112, N2028, N764, N39);
nand NAND4 (N3117, N3099, N1343, N1409, N1759);
buf BUF1 (N3118, N3117);
xor XOR2 (N3119, N3096, N1496);
or OR4 (N3120, N3114, N779, N100, N2307);
or OR2 (N3121, N3119, N2388);
and AND3 (N3122, N3105, N1536, N1393);
and AND4 (N3123, N3116, N2118, N2438, N631);
not NOT1 (N3124, N3120);
and AND3 (N3125, N3095, N2346, N1325);
or OR3 (N3126, N3125, N890, N537);
nor NOR2 (N3127, N3107, N2700);
xor XOR2 (N3128, N3126, N2994);
nor NOR4 (N3129, N3122, N42, N845, N2837);
nor NOR4 (N3130, N3124, N2681, N2952, N398);
buf BUF1 (N3131, N3121);
and AND4 (N3132, N3110, N1010, N1312, N2347);
not NOT1 (N3133, N3129);
xor XOR2 (N3134, N3130, N440);
not NOT1 (N3135, N3127);
or OR2 (N3136, N3115, N2618);
and AND3 (N3137, N3118, N2330, N2);
or OR2 (N3138, N3136, N182);
xor XOR2 (N3139, N3133, N2856);
nor NOR4 (N3140, N3137, N1166, N1290, N2856);
nand NAND3 (N3141, N3131, N2362, N821);
xor XOR2 (N3142, N3132, N2030);
not NOT1 (N3143, N3123);
nor NOR3 (N3144, N3140, N1881, N2679);
and AND2 (N3145, N3113, N1874);
not NOT1 (N3146, N3134);
nor NOR2 (N3147, N3135, N2009);
nor NOR4 (N3148, N3145, N290, N2108, N283);
or OR2 (N3149, N3141, N739);
or OR3 (N3150, N3143, N3042, N2756);
nand NAND2 (N3151, N3142, N799);
not NOT1 (N3152, N3138);
xor XOR2 (N3153, N3147, N1604);
not NOT1 (N3154, N3146);
and AND2 (N3155, N3153, N755);
and AND4 (N3156, N3149, N679, N2436, N990);
buf BUF1 (N3157, N3154);
and AND2 (N3158, N3128, N1297);
xor XOR2 (N3159, N3155, N2584);
and AND4 (N3160, N3159, N175, N1246, N1372);
or OR2 (N3161, N3156, N1139);
or OR4 (N3162, N3161, N237, N2421, N2969);
not NOT1 (N3163, N3152);
nand NAND4 (N3164, N3160, N604, N1934, N2176);
nor NOR2 (N3165, N3139, N2074);
buf BUF1 (N3166, N3162);
buf BUF1 (N3167, N3157);
buf BUF1 (N3168, N3167);
not NOT1 (N3169, N3148);
xor XOR2 (N3170, N3158, N1909);
not NOT1 (N3171, N3165);
not NOT1 (N3172, N3168);
and AND4 (N3173, N3169, N3143, N2755, N785);
or OR4 (N3174, N3172, N3000, N2243, N2498);
buf BUF1 (N3175, N3174);
not NOT1 (N3176, N3144);
or OR4 (N3177, N3163, N2920, N2067, N858);
and AND3 (N3178, N3176, N40, N144);
buf BUF1 (N3179, N3171);
nand NAND2 (N3180, N3179, N2858);
nor NOR4 (N3181, N3173, N1455, N2099, N2319);
and AND2 (N3182, N3166, N218);
buf BUF1 (N3183, N3178);
buf BUF1 (N3184, N3182);
nand NAND2 (N3185, N3150, N1873);
xor XOR2 (N3186, N3181, N2866);
not NOT1 (N3187, N3184);
not NOT1 (N3188, N3187);
buf BUF1 (N3189, N3183);
nand NAND3 (N3190, N3186, N2066, N1613);
nand NAND3 (N3191, N3190, N2779, N527);
buf BUF1 (N3192, N3175);
or OR2 (N3193, N3185, N671);
nor NOR2 (N3194, N3151, N3054);
not NOT1 (N3195, N3193);
buf BUF1 (N3196, N3189);
buf BUF1 (N3197, N3180);
nor NOR2 (N3198, N3188, N1930);
not NOT1 (N3199, N3197);
or OR2 (N3200, N3195, N1259);
buf BUF1 (N3201, N3198);
nand NAND4 (N3202, N3164, N3011, N2702, N608);
not NOT1 (N3203, N3200);
or OR3 (N3204, N3196, N1251, N1220);
buf BUF1 (N3205, N3204);
nand NAND3 (N3206, N3199, N1927, N1409);
nand NAND3 (N3207, N3206, N3075, N2614);
and AND2 (N3208, N3177, N1327);
xor XOR2 (N3209, N3207, N2098);
not NOT1 (N3210, N3208);
and AND3 (N3211, N3202, N2546, N1682);
not NOT1 (N3212, N3170);
buf BUF1 (N3213, N3194);
nor NOR2 (N3214, N3191, N2712);
and AND4 (N3215, N3210, N1271, N121, N403);
buf BUF1 (N3216, N3205);
buf BUF1 (N3217, N3211);
nand NAND4 (N3218, N3217, N2574, N3117, N2027);
and AND2 (N3219, N3212, N482);
not NOT1 (N3220, N3209);
nand NAND3 (N3221, N3201, N2108, N321);
nor NOR3 (N3222, N3215, N3013, N1770);
nor NOR3 (N3223, N3213, N2218, N2585);
or OR4 (N3224, N3222, N2666, N2263, N2050);
or OR2 (N3225, N3218, N539);
nand NAND2 (N3226, N3220, N2245);
nor NOR4 (N3227, N3223, N197, N850, N2348);
and AND4 (N3228, N3224, N544, N2784, N2096);
or OR4 (N3229, N3192, N1582, N1370, N1416);
nand NAND4 (N3230, N3203, N725, N3137, N2659);
nor NOR3 (N3231, N3230, N932, N3021);
not NOT1 (N3232, N3225);
nor NOR2 (N3233, N3214, N3045);
xor XOR2 (N3234, N3221, N313);
nand NAND2 (N3235, N3231, N141);
xor XOR2 (N3236, N3226, N2461);
and AND3 (N3237, N3229, N2370, N2592);
and AND2 (N3238, N3216, N409);
nor NOR4 (N3239, N3227, N2498, N397, N2803);
nand NAND4 (N3240, N3234, N1166, N1806, N3008);
nand NAND3 (N3241, N3237, N1303, N338);
xor XOR2 (N3242, N3236, N2229);
not NOT1 (N3243, N3219);
nor NOR2 (N3244, N3242, N975);
nand NAND3 (N3245, N3240, N2942, N1940);
nor NOR2 (N3246, N3235, N2656);
buf BUF1 (N3247, N3233);
and AND3 (N3248, N3245, N2904, N2146);
or OR2 (N3249, N3244, N2361);
and AND4 (N3250, N3239, N1988, N1827, N2257);
not NOT1 (N3251, N3249);
nand NAND3 (N3252, N3241, N1634, N2115);
nor NOR3 (N3253, N3251, N2601, N2352);
or OR2 (N3254, N3228, N1191);
and AND4 (N3255, N3254, N489, N1798, N914);
buf BUF1 (N3256, N3243);
nand NAND2 (N3257, N3248, N1022);
not NOT1 (N3258, N3252);
nand NAND4 (N3259, N3250, N3127, N1290, N90);
or OR2 (N3260, N3246, N1384);
xor XOR2 (N3261, N3257, N3001);
or OR4 (N3262, N3258, N1581, N1073, N962);
xor XOR2 (N3263, N3247, N2780);
and AND4 (N3264, N3263, N1384, N2071, N2759);
or OR3 (N3265, N3261, N3125, N1621);
or OR4 (N3266, N3262, N2737, N1047, N2472);
buf BUF1 (N3267, N3255);
not NOT1 (N3268, N3259);
or OR3 (N3269, N3264, N777, N621);
buf BUF1 (N3270, N3268);
nand NAND3 (N3271, N3253, N2739, N1933);
buf BUF1 (N3272, N3238);
nor NOR2 (N3273, N3270, N2573);
buf BUF1 (N3274, N3260);
or OR2 (N3275, N3269, N2459);
buf BUF1 (N3276, N3256);
not NOT1 (N3277, N3276);
buf BUF1 (N3278, N3275);
nor NOR2 (N3279, N3266, N1155);
not NOT1 (N3280, N3272);
buf BUF1 (N3281, N3232);
nor NOR3 (N3282, N3280, N1640, N2504);
nand NAND2 (N3283, N3274, N1602);
buf BUF1 (N3284, N3265);
buf BUF1 (N3285, N3271);
and AND3 (N3286, N3283, N1768, N690);
xor XOR2 (N3287, N3273, N170);
not NOT1 (N3288, N3277);
nor NOR3 (N3289, N3267, N831, N2341);
xor XOR2 (N3290, N3289, N542);
nor NOR2 (N3291, N3282, N538);
nor NOR2 (N3292, N3288, N2473);
and AND4 (N3293, N3281, N955, N973, N1831);
and AND4 (N3294, N3278, N3165, N832, N2894);
buf BUF1 (N3295, N3286);
or OR2 (N3296, N3279, N392);
nand NAND2 (N3297, N3296, N3227);
nor NOR4 (N3298, N3292, N1087, N3017, N2686);
nor NOR4 (N3299, N3285, N7, N1220, N116);
or OR2 (N3300, N3298, N1412);
nor NOR4 (N3301, N3300, N41, N2172, N1549);
not NOT1 (N3302, N3297);
buf BUF1 (N3303, N3295);
xor XOR2 (N3304, N3301, N1070);
and AND3 (N3305, N3293, N504, N2810);
nand NAND3 (N3306, N3305, N3134, N988);
xor XOR2 (N3307, N3284, N788);
not NOT1 (N3308, N3291);
xor XOR2 (N3309, N3308, N89);
nor NOR2 (N3310, N3294, N1880);
xor XOR2 (N3311, N3304, N1230);
or OR4 (N3312, N3306, N3246, N2445, N2224);
or OR2 (N3313, N3307, N2771);
and AND3 (N3314, N3309, N58, N968);
or OR3 (N3315, N3312, N1102, N2516);
not NOT1 (N3316, N3315);
xor XOR2 (N3317, N3310, N1257);
and AND3 (N3318, N3287, N187, N3176);
and AND3 (N3319, N3317, N987, N397);
or OR2 (N3320, N3311, N807);
not NOT1 (N3321, N3303);
or OR4 (N3322, N3302, N1119, N1624, N3265);
nor NOR2 (N3323, N3321, N2724);
and AND4 (N3324, N3299, N1919, N3049, N946);
nor NOR3 (N3325, N3314, N2358, N1119);
buf BUF1 (N3326, N3325);
nor NOR2 (N3327, N3322, N859);
and AND2 (N3328, N3316, N3063);
nand NAND4 (N3329, N3323, N1758, N254, N2327);
nand NAND4 (N3330, N3326, N3315, N1115, N2595);
nor NOR3 (N3331, N3327, N3048, N1390);
or OR2 (N3332, N3313, N98);
not NOT1 (N3333, N3319);
xor XOR2 (N3334, N3331, N134);
nand NAND4 (N3335, N3332, N597, N1356, N959);
nor NOR3 (N3336, N3324, N2850, N389);
xor XOR2 (N3337, N3335, N2313);
and AND2 (N3338, N3318, N2033);
or OR2 (N3339, N3333, N1595);
nand NAND2 (N3340, N3337, N2628);
nor NOR3 (N3341, N3334, N186, N2205);
buf BUF1 (N3342, N3290);
and AND4 (N3343, N3342, N2158, N771, N1939);
or OR2 (N3344, N3330, N48);
and AND4 (N3345, N3343, N3210, N1347, N3297);
not NOT1 (N3346, N3338);
buf BUF1 (N3347, N3341);
xor XOR2 (N3348, N3339, N1969);
or OR4 (N3349, N3328, N282, N3154, N2506);
nor NOR3 (N3350, N3347, N909, N3266);
or OR4 (N3351, N3344, N833, N62, N633);
xor XOR2 (N3352, N3346, N2731);
or OR2 (N3353, N3345, N357);
xor XOR2 (N3354, N3351, N3074);
buf BUF1 (N3355, N3329);
buf BUF1 (N3356, N3348);
not NOT1 (N3357, N3340);
nor NOR3 (N3358, N3355, N1446, N302);
buf BUF1 (N3359, N3336);
nand NAND4 (N3360, N3350, N2979, N1851, N1287);
nand NAND4 (N3361, N3360, N1481, N2312, N3080);
nor NOR2 (N3362, N3354, N1813);
nor NOR3 (N3363, N3320, N1422, N1530);
buf BUF1 (N3364, N3362);
nand NAND2 (N3365, N3358, N745);
xor XOR2 (N3366, N3359, N1445);
buf BUF1 (N3367, N3361);
nand NAND4 (N3368, N3357, N2050, N818, N1928);
nor NOR2 (N3369, N3365, N774);
nor NOR2 (N3370, N3352, N2946);
buf BUF1 (N3371, N3367);
not NOT1 (N3372, N3363);
buf BUF1 (N3373, N3356);
or OR4 (N3374, N3370, N226, N543, N411);
nor NOR4 (N3375, N3366, N1610, N2902, N3142);
or OR4 (N3376, N3373, N2235, N321, N1997);
not NOT1 (N3377, N3375);
not NOT1 (N3378, N3377);
buf BUF1 (N3379, N3364);
and AND4 (N3380, N3371, N3337, N3328, N1049);
and AND4 (N3381, N3380, N1878, N2707, N2383);
and AND3 (N3382, N3374, N962, N2712);
or OR4 (N3383, N3349, N2621, N929, N2067);
or OR3 (N3384, N3372, N1775, N736);
or OR2 (N3385, N3369, N1707);
buf BUF1 (N3386, N3378);
and AND4 (N3387, N3384, N3012, N1225, N2630);
and AND2 (N3388, N3385, N3210);
buf BUF1 (N3389, N3383);
not NOT1 (N3390, N3387);
xor XOR2 (N3391, N3368, N481);
nor NOR3 (N3392, N3353, N1300, N1029);
and AND3 (N3393, N3391, N1074, N2909);
and AND3 (N3394, N3379, N1620, N464);
not NOT1 (N3395, N3394);
or OR3 (N3396, N3390, N757, N903);
and AND3 (N3397, N3396, N2454, N2597);
xor XOR2 (N3398, N3392, N735);
xor XOR2 (N3399, N3393, N3116);
nor NOR3 (N3400, N3399, N2976, N1015);
nor NOR3 (N3401, N3381, N3380, N440);
not NOT1 (N3402, N3397);
not NOT1 (N3403, N3398);
not NOT1 (N3404, N3388);
not NOT1 (N3405, N3404);
nand NAND3 (N3406, N3386, N193, N1940);
or OR4 (N3407, N3402, N1754, N2796, N2020);
nand NAND3 (N3408, N3405, N11, N1076);
xor XOR2 (N3409, N3408, N881);
nand NAND4 (N3410, N3406, N2405, N3144, N1960);
nand NAND2 (N3411, N3407, N3333);
or OR2 (N3412, N3382, N923);
xor XOR2 (N3413, N3389, N324);
nor NOR3 (N3414, N3401, N1612, N2279);
not NOT1 (N3415, N3376);
and AND2 (N3416, N3395, N944);
nor NOR3 (N3417, N3413, N2298, N1162);
xor XOR2 (N3418, N3410, N1413);
not NOT1 (N3419, N3416);
and AND4 (N3420, N3403, N2611, N3321, N1977);
nand NAND3 (N3421, N3411, N1611, N2500);
and AND2 (N3422, N3417, N290);
or OR2 (N3423, N3420, N1067);
and AND3 (N3424, N3400, N2531, N691);
and AND2 (N3425, N3418, N2096);
and AND3 (N3426, N3414, N2464, N1220);
not NOT1 (N3427, N3412);
buf BUF1 (N3428, N3423);
nand NAND3 (N3429, N3428, N1236, N2111);
or OR3 (N3430, N3424, N2688, N670);
or OR3 (N3431, N3415, N181, N935);
nor NOR3 (N3432, N3421, N831, N539);
buf BUF1 (N3433, N3432);
or OR4 (N3434, N3430, N3237, N31, N1249);
xor XOR2 (N3435, N3425, N2908);
xor XOR2 (N3436, N3429, N2471);
and AND2 (N3437, N3422, N1885);
buf BUF1 (N3438, N3437);
buf BUF1 (N3439, N3409);
nor NOR3 (N3440, N3427, N2634, N1016);
xor XOR2 (N3441, N3435, N1586);
nand NAND4 (N3442, N3426, N3146, N2258, N2913);
xor XOR2 (N3443, N3442, N2490);
xor XOR2 (N3444, N3434, N3418);
nand NAND2 (N3445, N3440, N1655);
or OR3 (N3446, N3419, N3271, N1179);
nor NOR2 (N3447, N3431, N2938);
and AND3 (N3448, N3445, N3378, N725);
and AND4 (N3449, N3446, N1520, N297, N1785);
or OR2 (N3450, N3448, N3091);
nand NAND3 (N3451, N3450, N2358, N1648);
nor NOR2 (N3452, N3439, N16);
xor XOR2 (N3453, N3443, N1234);
buf BUF1 (N3454, N3447);
buf BUF1 (N3455, N3451);
buf BUF1 (N3456, N3455);
and AND3 (N3457, N3441, N897, N716);
or OR2 (N3458, N3449, N2918);
and AND2 (N3459, N3456, N656);
or OR2 (N3460, N3433, N2078);
nor NOR2 (N3461, N3457, N2030);
xor XOR2 (N3462, N3436, N2871);
or OR2 (N3463, N3460, N683);
not NOT1 (N3464, N3461);
and AND2 (N3465, N3452, N714);
buf BUF1 (N3466, N3465);
xor XOR2 (N3467, N3464, N3461);
xor XOR2 (N3468, N3467, N1591);
and AND2 (N3469, N3453, N2774);
nor NOR3 (N3470, N3438, N891, N3274);
and AND2 (N3471, N3459, N2425);
nand NAND3 (N3472, N3463, N1382, N114);
xor XOR2 (N3473, N3458, N1814);
nand NAND3 (N3474, N3466, N863, N1479);
nor NOR2 (N3475, N3472, N1716);
or OR4 (N3476, N3470, N2612, N1458, N1272);
not NOT1 (N3477, N3475);
or OR2 (N3478, N3474, N2701);
xor XOR2 (N3479, N3478, N1696);
buf BUF1 (N3480, N3469);
or OR3 (N3481, N3454, N2771, N834);
nor NOR4 (N3482, N3471, N3242, N1713, N989);
not NOT1 (N3483, N3468);
xor XOR2 (N3484, N3473, N2586);
nand NAND2 (N3485, N3481, N3127);
or OR4 (N3486, N3477, N53, N1854, N791);
and AND4 (N3487, N3444, N2962, N1329, N2493);
or OR3 (N3488, N3480, N1093, N34);
buf BUF1 (N3489, N3484);
nand NAND4 (N3490, N3487, N2599, N2173, N1211);
buf BUF1 (N3491, N3476);
and AND2 (N3492, N3489, N525);
buf BUF1 (N3493, N3479);
or OR4 (N3494, N3493, N2419, N2109, N2183);
nand NAND2 (N3495, N3485, N2031);
xor XOR2 (N3496, N3492, N141);
not NOT1 (N3497, N3488);
xor XOR2 (N3498, N3462, N1029);
or OR2 (N3499, N3494, N1795);
buf BUF1 (N3500, N3490);
nor NOR3 (N3501, N3498, N1614, N2263);
and AND3 (N3502, N3500, N2953, N507);
nand NAND4 (N3503, N3499, N805, N316, N2342);
xor XOR2 (N3504, N3503, N2697);
nand NAND4 (N3505, N3502, N1963, N1686, N850);
not NOT1 (N3506, N3497);
nand NAND2 (N3507, N3506, N2461);
buf BUF1 (N3508, N3501);
xor XOR2 (N3509, N3486, N2865);
and AND2 (N3510, N3495, N784);
or OR4 (N3511, N3483, N2143, N754, N3131);
and AND4 (N3512, N3508, N1238, N1851, N666);
or OR3 (N3513, N3482, N358, N2893);
not NOT1 (N3514, N3504);
buf BUF1 (N3515, N3510);
xor XOR2 (N3516, N3496, N1261);
xor XOR2 (N3517, N3491, N878);
nor NOR3 (N3518, N3507, N629, N3010);
nor NOR3 (N3519, N3513, N1703, N1796);
or OR4 (N3520, N3505, N2214, N2781, N67);
xor XOR2 (N3521, N3511, N2896);
xor XOR2 (N3522, N3517, N497);
or OR3 (N3523, N3519, N2012, N435);
xor XOR2 (N3524, N3521, N3144);
and AND2 (N3525, N3523, N2283);
not NOT1 (N3526, N3518);
or OR2 (N3527, N3516, N951);
buf BUF1 (N3528, N3524);
buf BUF1 (N3529, N3515);
or OR3 (N3530, N3514, N1429, N2708);
buf BUF1 (N3531, N3522);
xor XOR2 (N3532, N3520, N993);
nand NAND4 (N3533, N3531, N36, N250, N261);
nor NOR2 (N3534, N3530, N665);
nand NAND3 (N3535, N3512, N1857, N2245);
or OR3 (N3536, N3527, N2914, N103);
and AND4 (N3537, N3529, N468, N3254, N3171);
buf BUF1 (N3538, N3537);
nor NOR3 (N3539, N3535, N1196, N2842);
nand NAND2 (N3540, N3533, N1918);
and AND2 (N3541, N3539, N1901);
nand NAND2 (N3542, N3540, N3337);
xor XOR2 (N3543, N3528, N587);
or OR4 (N3544, N3532, N2423, N149, N969);
not NOT1 (N3545, N3541);
xor XOR2 (N3546, N3538, N161);
or OR3 (N3547, N3536, N3488, N692);
not NOT1 (N3548, N3546);
nand NAND4 (N3549, N3526, N3144, N1351, N1460);
or OR4 (N3550, N3509, N1676, N131, N1895);
nand NAND4 (N3551, N3534, N2704, N2424, N2414);
buf BUF1 (N3552, N3547);
and AND2 (N3553, N3542, N3128);
nand NAND4 (N3554, N3548, N2804, N2790, N1864);
buf BUF1 (N3555, N3549);
xor XOR2 (N3556, N3551, N960);
nand NAND4 (N3557, N3525, N1999, N3375, N3550);
nand NAND2 (N3558, N2269, N1885);
and AND2 (N3559, N3554, N33);
nor NOR2 (N3560, N3558, N2743);
not NOT1 (N3561, N3557);
nand NAND3 (N3562, N3543, N2065, N1693);
nor NOR2 (N3563, N3556, N964);
xor XOR2 (N3564, N3545, N574);
nor NOR3 (N3565, N3555, N3377, N354);
or OR3 (N3566, N3564, N360, N2671);
nand NAND4 (N3567, N3559, N3351, N297, N2332);
not NOT1 (N3568, N3560);
not NOT1 (N3569, N3563);
xor XOR2 (N3570, N3562, N1676);
nand NAND4 (N3571, N3565, N1420, N3014, N1042);
xor XOR2 (N3572, N3553, N2972);
nor NOR2 (N3573, N3544, N828);
buf BUF1 (N3574, N3567);
nand NAND3 (N3575, N3573, N3534, N3256);
nand NAND2 (N3576, N3552, N3219);
nor NOR2 (N3577, N3569, N4);
nor NOR2 (N3578, N3571, N2915);
buf BUF1 (N3579, N3574);
nor NOR3 (N3580, N3568, N51, N89);
and AND3 (N3581, N3577, N542, N2056);
and AND4 (N3582, N3561, N1194, N1675, N1231);
nor NOR4 (N3583, N3576, N1515, N3276, N1499);
xor XOR2 (N3584, N3582, N2536);
nand NAND4 (N3585, N3572, N224, N300, N1990);
or OR4 (N3586, N3575, N3241, N1779, N3173);
xor XOR2 (N3587, N3586, N1502);
nor NOR3 (N3588, N3585, N278, N3547);
or OR3 (N3589, N3566, N2648, N2166);
and AND4 (N3590, N3578, N1717, N1849, N3526);
xor XOR2 (N3591, N3589, N143);
or OR3 (N3592, N3570, N3161, N3026);
nand NAND4 (N3593, N3584, N715, N3068, N2292);
nand NAND2 (N3594, N3593, N139);
nor NOR2 (N3595, N3591, N1422);
xor XOR2 (N3596, N3580, N2346);
not NOT1 (N3597, N3590);
buf BUF1 (N3598, N3596);
xor XOR2 (N3599, N3579, N1619);
nand NAND4 (N3600, N3595, N3432, N1839, N3153);
xor XOR2 (N3601, N3598, N1984);
buf BUF1 (N3602, N3597);
nand NAND3 (N3603, N3602, N3534, N2601);
not NOT1 (N3604, N3594);
not NOT1 (N3605, N3592);
nor NOR2 (N3606, N3600, N2150);
and AND4 (N3607, N3606, N22, N1443, N2495);
nand NAND4 (N3608, N3599, N140, N2232, N1052);
nand NAND4 (N3609, N3608, N3107, N1827, N3087);
nor NOR3 (N3610, N3604, N1655, N1174);
nor NOR2 (N3611, N3583, N3475);
nand NAND3 (N3612, N3581, N64, N220);
and AND2 (N3613, N3610, N3031);
xor XOR2 (N3614, N3613, N200);
nand NAND2 (N3615, N3611, N415);
nand NAND4 (N3616, N3588, N1946, N6, N386);
nand NAND4 (N3617, N3587, N1855, N133, N795);
xor XOR2 (N3618, N3605, N810);
buf BUF1 (N3619, N3615);
xor XOR2 (N3620, N3617, N2661);
xor XOR2 (N3621, N3601, N31);
and AND3 (N3622, N3621, N311, N1109);
or OR4 (N3623, N3609, N1551, N1918, N633);
and AND3 (N3624, N3614, N3516, N363);
not NOT1 (N3625, N3612);
and AND3 (N3626, N3623, N3000, N572);
xor XOR2 (N3627, N3603, N2378);
not NOT1 (N3628, N3616);
not NOT1 (N3629, N3628);
buf BUF1 (N3630, N3629);
or OR4 (N3631, N3626, N2289, N1814, N1671);
or OR4 (N3632, N3624, N1985, N725, N1505);
not NOT1 (N3633, N3631);
and AND4 (N3634, N3633, N1718, N2161, N1637);
buf BUF1 (N3635, N3630);
xor XOR2 (N3636, N3619, N1004);
and AND2 (N3637, N3636, N1271);
or OR3 (N3638, N3635, N899, N2466);
buf BUF1 (N3639, N3618);
not NOT1 (N3640, N3639);
and AND2 (N3641, N3622, N2135);
and AND3 (N3642, N3625, N3430, N2591);
and AND2 (N3643, N3640, N2986);
and AND3 (N3644, N3620, N2185, N2703);
or OR4 (N3645, N3607, N2147, N3179, N1574);
not NOT1 (N3646, N3643);
xor XOR2 (N3647, N3642, N3155);
or OR2 (N3648, N3632, N522);
xor XOR2 (N3649, N3647, N362);
not NOT1 (N3650, N3644);
or OR3 (N3651, N3627, N438, N582);
nand NAND3 (N3652, N3645, N2715, N1538);
not NOT1 (N3653, N3638);
and AND4 (N3654, N3634, N1635, N63, N2045);
or OR3 (N3655, N3653, N458, N2848);
nand NAND3 (N3656, N3646, N3448, N940);
and AND2 (N3657, N3649, N682);
xor XOR2 (N3658, N3637, N1636);
nor NOR2 (N3659, N3658, N578);
buf BUF1 (N3660, N3650);
nor NOR4 (N3661, N3657, N142, N517, N480);
buf BUF1 (N3662, N3656);
not NOT1 (N3663, N3660);
not NOT1 (N3664, N3652);
xor XOR2 (N3665, N3663, N2004);
buf BUF1 (N3666, N3654);
nand NAND4 (N3667, N3641, N1801, N1624, N1133);
xor XOR2 (N3668, N3648, N475);
and AND4 (N3669, N3668, N3530, N3567, N2590);
buf BUF1 (N3670, N3655);
nor NOR3 (N3671, N3667, N76, N316);
not NOT1 (N3672, N3665);
or OR3 (N3673, N3662, N2, N1795);
nor NOR4 (N3674, N3669, N1897, N815, N3574);
or OR4 (N3675, N3651, N1356, N3112, N1177);
and AND3 (N3676, N3673, N801, N1921);
nand NAND2 (N3677, N3674, N80);
and AND3 (N3678, N3677, N464, N2927);
not NOT1 (N3679, N3664);
not NOT1 (N3680, N3676);
not NOT1 (N3681, N3675);
or OR3 (N3682, N3678, N1884, N1571);
xor XOR2 (N3683, N3680, N3641);
or OR3 (N3684, N3671, N2489, N2160);
nor NOR4 (N3685, N3670, N1812, N1586, N1482);
xor XOR2 (N3686, N3666, N1568);
buf BUF1 (N3687, N3681);
not NOT1 (N3688, N3659);
nand NAND2 (N3689, N3679, N3657);
not NOT1 (N3690, N3686);
buf BUF1 (N3691, N3685);
buf BUF1 (N3692, N3689);
not NOT1 (N3693, N3688);
or OR2 (N3694, N3683, N1594);
xor XOR2 (N3695, N3684, N556);
nor NOR4 (N3696, N3690, N1057, N2237, N2360);
or OR2 (N3697, N3696, N3198);
nor NOR4 (N3698, N3692, N2370, N3278, N1864);
xor XOR2 (N3699, N3687, N2116);
or OR3 (N3700, N3694, N3037, N1880);
or OR4 (N3701, N3691, N2098, N2004, N316);
not NOT1 (N3702, N3661);
and AND2 (N3703, N3695, N3420);
and AND2 (N3704, N3700, N1530);
buf BUF1 (N3705, N3672);
or OR4 (N3706, N3697, N2717, N1116, N226);
nand NAND3 (N3707, N3702, N1222, N1504);
nor NOR2 (N3708, N3693, N1078);
or OR3 (N3709, N3682, N448, N3136);
nor NOR3 (N3710, N3708, N9, N1046);
nor NOR4 (N3711, N3703, N822, N1527, N885);
and AND3 (N3712, N3711, N1234, N2167);
nor NOR4 (N3713, N3712, N514, N2188, N1771);
buf BUF1 (N3714, N3709);
nor NOR3 (N3715, N3699, N98, N285);
not NOT1 (N3716, N3706);
nor NOR3 (N3717, N3707, N1982, N1271);
buf BUF1 (N3718, N3714);
and AND2 (N3719, N3716, N2867);
nor NOR3 (N3720, N3718, N2478, N610);
not NOT1 (N3721, N3719);
nor NOR4 (N3722, N3701, N2248, N1261, N2393);
and AND4 (N3723, N3698, N1095, N1621, N3121);
not NOT1 (N3724, N3720);
and AND3 (N3725, N3710, N1363, N1502);
and AND2 (N3726, N3722, N2190);
xor XOR2 (N3727, N3704, N3095);
and AND2 (N3728, N3727, N3365);
buf BUF1 (N3729, N3725);
and AND3 (N3730, N3721, N1361, N1665);
nand NAND4 (N3731, N3705, N1237, N3624, N3713);
nand NAND4 (N3732, N2251, N3269, N1410, N3699);
not NOT1 (N3733, N3715);
or OR4 (N3734, N3717, N1803, N905, N580);
not NOT1 (N3735, N3732);
buf BUF1 (N3736, N3734);
and AND2 (N3737, N3730, N263);
and AND2 (N3738, N3728, N1269);
buf BUF1 (N3739, N3738);
nand NAND4 (N3740, N3736, N390, N1962, N2789);
nor NOR2 (N3741, N3739, N484);
and AND3 (N3742, N3729, N3152, N3063);
xor XOR2 (N3743, N3740, N39);
nand NAND3 (N3744, N3742, N2670, N684);
nand NAND3 (N3745, N3741, N2841, N1316);
xor XOR2 (N3746, N3724, N914);
xor XOR2 (N3747, N3735, N1834);
not NOT1 (N3748, N3745);
nand NAND2 (N3749, N3746, N43);
not NOT1 (N3750, N3744);
nand NAND2 (N3751, N3748, N945);
not NOT1 (N3752, N3737);
and AND2 (N3753, N3733, N2992);
or OR4 (N3754, N3750, N161, N3728, N2713);
and AND3 (N3755, N3751, N974, N1593);
nand NAND4 (N3756, N3755, N1607, N1126, N2625);
buf BUF1 (N3757, N3752);
not NOT1 (N3758, N3749);
or OR4 (N3759, N3747, N386, N3399, N2318);
xor XOR2 (N3760, N3754, N194);
buf BUF1 (N3761, N3756);
or OR2 (N3762, N3731, N3031);
and AND4 (N3763, N3757, N2917, N2246, N1265);
or OR3 (N3764, N3759, N1569, N1301);
or OR2 (N3765, N3723, N497);
nand NAND3 (N3766, N3765, N1220, N870);
buf BUF1 (N3767, N3760);
buf BUF1 (N3768, N3726);
nand NAND2 (N3769, N3762, N148);
buf BUF1 (N3770, N3743);
or OR3 (N3771, N3766, N3282, N2701);
buf BUF1 (N3772, N3758);
xor XOR2 (N3773, N3764, N1689);
not NOT1 (N3774, N3771);
buf BUF1 (N3775, N3761);
or OR3 (N3776, N3763, N3469, N84);
not NOT1 (N3777, N3768);
not NOT1 (N3778, N3773);
not NOT1 (N3779, N3769);
or OR3 (N3780, N3753, N544, N2210);
and AND3 (N3781, N3778, N312, N1702);
and AND4 (N3782, N3779, N2266, N2148, N1790);
nand NAND4 (N3783, N3767, N3444, N2965, N680);
nor NOR4 (N3784, N3777, N3187, N128, N2247);
and AND4 (N3785, N3772, N733, N2396, N1754);
nand NAND4 (N3786, N3783, N2891, N817, N273);
or OR3 (N3787, N3774, N178, N3333);
nor NOR2 (N3788, N3776, N2604);
nor NOR3 (N3789, N3786, N2639, N3104);
nor NOR2 (N3790, N3789, N714);
nand NAND4 (N3791, N3770, N2270, N1787, N2195);
not NOT1 (N3792, N3781);
xor XOR2 (N3793, N3788, N25);
nand NAND2 (N3794, N3782, N1353);
nor NOR2 (N3795, N3790, N2157);
buf BUF1 (N3796, N3775);
or OR3 (N3797, N3794, N42, N811);
or OR2 (N3798, N3793, N1447);
buf BUF1 (N3799, N3797);
nand NAND2 (N3800, N3796, N1015);
or OR2 (N3801, N3791, N2939);
nand NAND2 (N3802, N3801, N822);
and AND2 (N3803, N3785, N3315);
and AND2 (N3804, N3784, N3641);
and AND2 (N3805, N3780, N2720);
not NOT1 (N3806, N3800);
or OR3 (N3807, N3802, N397, N3445);
and AND2 (N3808, N3806, N602);
and AND2 (N3809, N3807, N2890);
nor NOR3 (N3810, N3798, N1878, N2796);
buf BUF1 (N3811, N3808);
or OR3 (N3812, N3805, N3433, N3802);
nor NOR2 (N3813, N3809, N2706);
xor XOR2 (N3814, N3792, N2323);
not NOT1 (N3815, N3799);
nor NOR2 (N3816, N3787, N1132);
or OR3 (N3817, N3816, N1009, N788);
buf BUF1 (N3818, N3804);
xor XOR2 (N3819, N3795, N1644);
or OR4 (N3820, N3810, N1834, N2325, N1357);
or OR3 (N3821, N3818, N283, N2779);
or OR4 (N3822, N3813, N1715, N59, N3718);
nor NOR2 (N3823, N3822, N1222);
and AND3 (N3824, N3820, N3613, N1430);
nand NAND2 (N3825, N3821, N1111);
and AND4 (N3826, N3815, N2265, N1466, N1032);
xor XOR2 (N3827, N3819, N1450);
not NOT1 (N3828, N3812);
nor NOR2 (N3829, N3828, N3746);
xor XOR2 (N3830, N3825, N1395);
nor NOR4 (N3831, N3823, N1774, N2382, N3372);
buf BUF1 (N3832, N3824);
not NOT1 (N3833, N3814);
xor XOR2 (N3834, N3831, N1863);
buf BUF1 (N3835, N3833);
or OR3 (N3836, N3832, N2632, N1618);
buf BUF1 (N3837, N3830);
not NOT1 (N3838, N3837);
not NOT1 (N3839, N3829);
buf BUF1 (N3840, N3836);
buf BUF1 (N3841, N3839);
xor XOR2 (N3842, N3838, N3409);
xor XOR2 (N3843, N3842, N3764);
buf BUF1 (N3844, N3841);
xor XOR2 (N3845, N3803, N3254);
buf BUF1 (N3846, N3845);
or OR4 (N3847, N3843, N982, N3537, N2396);
not NOT1 (N3848, N3817);
nand NAND3 (N3849, N3834, N1614, N1400);
nand NAND3 (N3850, N3849, N1966, N521);
or OR2 (N3851, N3840, N1481);
nor NOR2 (N3852, N3851, N2578);
xor XOR2 (N3853, N3852, N962);
nor NOR3 (N3854, N3853, N1223, N139);
nor NOR3 (N3855, N3844, N484, N1437);
nand NAND4 (N3856, N3854, N3162, N2984, N2000);
nand NAND4 (N3857, N3826, N3502, N335, N549);
nor NOR3 (N3858, N3857, N1537, N2009);
nor NOR4 (N3859, N3856, N182, N34, N2652);
nor NOR4 (N3860, N3827, N3310, N614, N3764);
xor XOR2 (N3861, N3859, N2000);
and AND3 (N3862, N3860, N85, N1712);
not NOT1 (N3863, N3811);
xor XOR2 (N3864, N3835, N2575);
and AND4 (N3865, N3864, N1019, N3394, N3334);
xor XOR2 (N3866, N3861, N2473);
nor NOR3 (N3867, N3862, N3844, N1768);
not NOT1 (N3868, N3846);
not NOT1 (N3869, N3848);
xor XOR2 (N3870, N3866, N3508);
not NOT1 (N3871, N3865);
and AND3 (N3872, N3871, N1379, N2860);
xor XOR2 (N3873, N3850, N1189);
nor NOR4 (N3874, N3847, N3659, N2970, N10);
nor NOR3 (N3875, N3867, N1141, N1474);
nor NOR3 (N3876, N3868, N2250, N2790);
buf BUF1 (N3877, N3869);
nor NOR2 (N3878, N3863, N1518);
xor XOR2 (N3879, N3855, N721);
and AND2 (N3880, N3870, N3756);
nand NAND4 (N3881, N3876, N99, N616, N1825);
or OR4 (N3882, N3858, N2730, N1433, N1271);
nand NAND4 (N3883, N3881, N3701, N957, N2593);
not NOT1 (N3884, N3878);
nor NOR4 (N3885, N3875, N1355, N693, N2824);
nand NAND3 (N3886, N3884, N2055, N1965);
or OR3 (N3887, N3873, N2430, N1674);
not NOT1 (N3888, N3882);
buf BUF1 (N3889, N3874);
buf BUF1 (N3890, N3880);
xor XOR2 (N3891, N3885, N61);
and AND4 (N3892, N3879, N3044, N3803, N2844);
or OR2 (N3893, N3891, N474);
nor NOR2 (N3894, N3893, N405);
xor XOR2 (N3895, N3883, N2091);
nand NAND4 (N3896, N3877, N3317, N2498, N2249);
and AND2 (N3897, N3890, N2441);
buf BUF1 (N3898, N3897);
nand NAND4 (N3899, N3894, N2817, N3148, N1390);
xor XOR2 (N3900, N3899, N3869);
or OR3 (N3901, N3886, N1135, N547);
not NOT1 (N3902, N3887);
not NOT1 (N3903, N3900);
buf BUF1 (N3904, N3896);
or OR2 (N3905, N3904, N2128);
buf BUF1 (N3906, N3903);
nor NOR3 (N3907, N3901, N2373, N3220);
buf BUF1 (N3908, N3905);
and AND4 (N3909, N3908, N1738, N2267, N1532);
and AND3 (N3910, N3892, N3040, N3039);
xor XOR2 (N3911, N3898, N2878);
buf BUF1 (N3912, N3889);
buf BUF1 (N3913, N3906);
and AND4 (N3914, N3912, N311, N350, N3077);
and AND3 (N3915, N3895, N3730, N2232);
nor NOR4 (N3916, N3872, N2721, N2118, N409);
nand NAND3 (N3917, N3911, N746, N3789);
nor NOR2 (N3918, N3888, N1938);
not NOT1 (N3919, N3907);
not NOT1 (N3920, N3914);
and AND3 (N3921, N3915, N1826, N1643);
not NOT1 (N3922, N3910);
and AND4 (N3923, N3920, N2999, N3768, N2468);
not NOT1 (N3924, N3922);
not NOT1 (N3925, N3921);
or OR3 (N3926, N3917, N2861, N910);
or OR2 (N3927, N3913, N1971);
not NOT1 (N3928, N3925);
nor NOR3 (N3929, N3918, N2989, N2262);
nor NOR3 (N3930, N3916, N3428, N1512);
nand NAND2 (N3931, N3924, N1132);
and AND3 (N3932, N3930, N239, N2764);
or OR4 (N3933, N3931, N2196, N3286, N276);
buf BUF1 (N3934, N3933);
not NOT1 (N3935, N3919);
buf BUF1 (N3936, N3932);
or OR2 (N3937, N3936, N741);
not NOT1 (N3938, N3902);
nand NAND2 (N3939, N3928, N3270);
nor NOR3 (N3940, N3926, N3459, N2281);
not NOT1 (N3941, N3923);
nor NOR4 (N3942, N3927, N3086, N2544, N2906);
xor XOR2 (N3943, N3937, N162);
not NOT1 (N3944, N3943);
not NOT1 (N3945, N3939);
not NOT1 (N3946, N3944);
nand NAND2 (N3947, N3938, N275);
not NOT1 (N3948, N3947);
and AND3 (N3949, N3942, N2713, N1776);
buf BUF1 (N3950, N3929);
not NOT1 (N3951, N3949);
or OR3 (N3952, N3948, N1371, N367);
nand NAND2 (N3953, N3934, N47);
or OR2 (N3954, N3952, N2028);
xor XOR2 (N3955, N3954, N3433);
or OR2 (N3956, N3909, N62);
xor XOR2 (N3957, N3951, N1783);
or OR4 (N3958, N3945, N3744, N2587, N1738);
or OR4 (N3959, N3940, N2439, N1448, N1296);
nor NOR4 (N3960, N3941, N3290, N1760, N1294);
not NOT1 (N3961, N3935);
nor NOR4 (N3962, N3946, N550, N3340, N2820);
nor NOR2 (N3963, N3953, N3101);
and AND4 (N3964, N3957, N990, N894, N1414);
not NOT1 (N3965, N3963);
and AND3 (N3966, N3950, N190, N3525);
buf BUF1 (N3967, N3955);
xor XOR2 (N3968, N3966, N3380);
nand NAND3 (N3969, N3964, N2312, N825);
xor XOR2 (N3970, N3959, N393);
and AND3 (N3971, N3968, N203, N664);
xor XOR2 (N3972, N3958, N519);
and AND2 (N3973, N3965, N1052);
nor NOR4 (N3974, N3960, N1527, N3098, N637);
buf BUF1 (N3975, N3974);
not NOT1 (N3976, N3975);
and AND2 (N3977, N3971, N3731);
xor XOR2 (N3978, N3956, N1932);
buf BUF1 (N3979, N3977);
xor XOR2 (N3980, N3961, N1853);
xor XOR2 (N3981, N3976, N219);
nand NAND4 (N3982, N3973, N3903, N2556, N3343);
not NOT1 (N3983, N3969);
buf BUF1 (N3984, N3962);
not NOT1 (N3985, N3972);
nand NAND2 (N3986, N3985, N3130);
not NOT1 (N3987, N3979);
buf BUF1 (N3988, N3983);
not NOT1 (N3989, N3970);
nor NOR2 (N3990, N3987, N3921);
and AND4 (N3991, N3990, N3929, N1688, N1333);
and AND3 (N3992, N3967, N1396, N2831);
nand NAND3 (N3993, N3980, N2396, N1746);
not NOT1 (N3994, N3993);
and AND2 (N3995, N3988, N3994);
nor NOR2 (N3996, N820, N1140);
buf BUF1 (N3997, N3978);
nor NOR2 (N3998, N3986, N3987);
and AND2 (N3999, N3997, N987);
xor XOR2 (N4000, N3984, N1107);
xor XOR2 (N4001, N3999, N2207);
and AND2 (N4002, N3998, N539);
nand NAND4 (N4003, N4002, N2183, N1986, N2924);
nand NAND3 (N4004, N4003, N823, N961);
nor NOR3 (N4005, N4000, N372, N2749);
or OR3 (N4006, N4001, N2503, N3693);
and AND3 (N4007, N3982, N3628, N849);
and AND3 (N4008, N3991, N2469, N955);
nor NOR4 (N4009, N4006, N1158, N3004, N2307);
buf BUF1 (N4010, N4005);
xor XOR2 (N4011, N3992, N2752);
nor NOR3 (N4012, N4009, N29, N501);
or OR2 (N4013, N4011, N619);
buf BUF1 (N4014, N3995);
xor XOR2 (N4015, N4012, N1096);
and AND2 (N4016, N4013, N505);
buf BUF1 (N4017, N4008);
buf BUF1 (N4018, N4014);
not NOT1 (N4019, N4015);
xor XOR2 (N4020, N3996, N3531);
xor XOR2 (N4021, N4010, N1280);
or OR3 (N4022, N3989, N3764, N1936);
xor XOR2 (N4023, N4020, N1797);
nor NOR3 (N4024, N4016, N2676, N3361);
nor NOR3 (N4025, N4019, N805, N1663);
and AND4 (N4026, N4024, N1034, N3237, N2375);
or OR3 (N4027, N4026, N3680, N986);
xor XOR2 (N4028, N4027, N3789);
nor NOR3 (N4029, N3981, N2077, N2791);
not NOT1 (N4030, N4022);
or OR4 (N4031, N4021, N690, N1514, N2520);
nand NAND3 (N4032, N4007, N3217, N3110);
or OR3 (N4033, N4004, N2625, N1177);
or OR3 (N4034, N4033, N3041, N3155);
and AND4 (N4035, N4032, N18, N372, N1909);
and AND3 (N4036, N4028, N3426, N767);
not NOT1 (N4037, N4025);
and AND3 (N4038, N4035, N3721, N413);
or OR2 (N4039, N4029, N2317);
not NOT1 (N4040, N4030);
not NOT1 (N4041, N4031);
buf BUF1 (N4042, N4036);
and AND3 (N4043, N4037, N1715, N104);
or OR2 (N4044, N4039, N481);
and AND3 (N4045, N4017, N1898, N2839);
not NOT1 (N4046, N4041);
and AND4 (N4047, N4018, N3620, N506, N2287);
nand NAND4 (N4048, N4043, N1567, N2159, N703);
nand NAND4 (N4049, N4034, N458, N2789, N1006);
nor NOR4 (N4050, N4042, N1675, N1338, N1442);
nand NAND4 (N4051, N4045, N2259, N375, N3268);
or OR2 (N4052, N4048, N878);
nor NOR2 (N4053, N4040, N2495);
nor NOR3 (N4054, N4050, N1490, N4036);
and AND2 (N4055, N4023, N3142);
and AND3 (N4056, N4047, N877, N1893);
nor NOR2 (N4057, N4046, N2424);
and AND3 (N4058, N4055, N1063, N1571);
xor XOR2 (N4059, N4054, N1812);
nand NAND2 (N4060, N4056, N1297);
and AND3 (N4061, N4060, N2060, N3437);
nand NAND4 (N4062, N4044, N1524, N3853, N2298);
nand NAND4 (N4063, N4061, N96, N2790, N2674);
xor XOR2 (N4064, N4057, N1471);
nand NAND3 (N4065, N4062, N3548, N1321);
buf BUF1 (N4066, N4053);
buf BUF1 (N4067, N4049);
and AND3 (N4068, N4038, N1118, N2848);
xor XOR2 (N4069, N4064, N2143);
not NOT1 (N4070, N4063);
nor NOR2 (N4071, N4067, N2712);
buf BUF1 (N4072, N4058);
nor NOR4 (N4073, N4072, N3171, N1192, N1129);
nor NOR3 (N4074, N4059, N390, N546);
and AND2 (N4075, N4052, N2826);
nor NOR3 (N4076, N4066, N3699, N1855);
nand NAND3 (N4077, N4071, N3187, N3635);
nand NAND2 (N4078, N4065, N3207);
or OR3 (N4079, N4068, N2740, N3170);
or OR2 (N4080, N4074, N658);
buf BUF1 (N4081, N4076);
or OR4 (N4082, N4077, N3721, N2868, N2448);
buf BUF1 (N4083, N4080);
buf BUF1 (N4084, N4079);
or OR4 (N4085, N4081, N784, N300, N1015);
and AND3 (N4086, N4069, N2186, N3646);
or OR4 (N4087, N4083, N3411, N1341, N3008);
buf BUF1 (N4088, N4087);
xor XOR2 (N4089, N4086, N425);
and AND2 (N4090, N4085, N2993);
xor XOR2 (N4091, N4075, N3134);
nor NOR3 (N4092, N4091, N1735, N4059);
xor XOR2 (N4093, N4092, N1639);
not NOT1 (N4094, N4073);
xor XOR2 (N4095, N4088, N3367);
not NOT1 (N4096, N4090);
nor NOR2 (N4097, N4094, N2134);
nor NOR4 (N4098, N4096, N3067, N2410, N3285);
xor XOR2 (N4099, N4089, N924);
nor NOR3 (N4100, N4070, N2729, N2795);
nand NAND4 (N4101, N4082, N3982, N3321, N1298);
not NOT1 (N4102, N4100);
buf BUF1 (N4103, N4051);
xor XOR2 (N4104, N4099, N3349);
buf BUF1 (N4105, N4103);
nor NOR4 (N4106, N4101, N679, N2768, N1704);
nor NOR4 (N4107, N4097, N1094, N3836, N3527);
and AND3 (N4108, N4098, N1320, N3195);
not NOT1 (N4109, N4084);
buf BUF1 (N4110, N4078);
nor NOR2 (N4111, N4108, N2080);
xor XOR2 (N4112, N4106, N693);
nor NOR3 (N4113, N4107, N110, N2066);
nand NAND3 (N4114, N4093, N1136, N979);
nor NOR3 (N4115, N4102, N3994, N232);
xor XOR2 (N4116, N4112, N1944);
not NOT1 (N4117, N4105);
and AND4 (N4118, N4110, N3090, N2095, N1845);
and AND2 (N4119, N4115, N2554);
and AND4 (N4120, N4114, N3012, N185, N2319);
or OR3 (N4121, N4095, N3939, N2505);
buf BUF1 (N4122, N4120);
not NOT1 (N4123, N4111);
not NOT1 (N4124, N4109);
buf BUF1 (N4125, N4104);
nor NOR4 (N4126, N4122, N2314, N4049, N1590);
nand NAND2 (N4127, N4121, N949);
and AND2 (N4128, N4118, N3533);
nor NOR4 (N4129, N4127, N719, N739, N2843);
not NOT1 (N4130, N4116);
nor NOR2 (N4131, N4128, N2917);
nor NOR2 (N4132, N4117, N148);
buf BUF1 (N4133, N4125);
xor XOR2 (N4134, N4126, N3034);
nor NOR2 (N4135, N4131, N1769);
xor XOR2 (N4136, N4119, N4133);
or OR2 (N4137, N2838, N1963);
and AND2 (N4138, N4136, N1505);
buf BUF1 (N4139, N4137);
xor XOR2 (N4140, N4130, N2617);
nand NAND4 (N4141, N4124, N3081, N2271, N3468);
nand NAND3 (N4142, N4134, N827, N3944);
buf BUF1 (N4143, N4129);
nor NOR4 (N4144, N4141, N1376, N2123, N2831);
nand NAND3 (N4145, N4144, N1617, N113);
xor XOR2 (N4146, N4138, N2394);
xor XOR2 (N4147, N4140, N1660);
nor NOR2 (N4148, N4139, N1291);
xor XOR2 (N4149, N4143, N3367);
or OR4 (N4150, N4145, N3546, N3289, N3706);
nor NOR4 (N4151, N4113, N3428, N2109, N753);
or OR2 (N4152, N4123, N1024);
xor XOR2 (N4153, N4148, N4118);
xor XOR2 (N4154, N4152, N3271);
xor XOR2 (N4155, N4149, N1812);
and AND2 (N4156, N4150, N2430);
buf BUF1 (N4157, N4146);
and AND2 (N4158, N4147, N3777);
xor XOR2 (N4159, N4151, N2184);
nand NAND3 (N4160, N4153, N2029, N3198);
or OR2 (N4161, N4135, N3895);
nor NOR2 (N4162, N4154, N3443);
nand NAND3 (N4163, N4156, N2928, N1360);
and AND4 (N4164, N4163, N3599, N3021, N1044);
nor NOR3 (N4165, N4162, N2234, N3821);
or OR2 (N4166, N4164, N2720);
not NOT1 (N4167, N4159);
or OR2 (N4168, N4155, N3737);
not NOT1 (N4169, N4165);
nand NAND4 (N4170, N4166, N2475, N2219, N1877);
xor XOR2 (N4171, N4161, N947);
or OR3 (N4172, N4158, N597, N1658);
not NOT1 (N4173, N4168);
not NOT1 (N4174, N4171);
xor XOR2 (N4175, N4170, N1534);
nand NAND4 (N4176, N4132, N1557, N2672, N311);
nor NOR2 (N4177, N4142, N97);
nor NOR2 (N4178, N4176, N4056);
nand NAND2 (N4179, N4173, N806);
and AND4 (N4180, N4175, N2421, N1499, N1488);
nor NOR3 (N4181, N4167, N3734, N2083);
or OR3 (N4182, N4178, N1293, N1809);
xor XOR2 (N4183, N4172, N3100);
nand NAND2 (N4184, N4177, N1022);
nor NOR2 (N4185, N4179, N1836);
not NOT1 (N4186, N4185);
not NOT1 (N4187, N4157);
nor NOR2 (N4188, N4186, N2071);
nor NOR2 (N4189, N4187, N670);
or OR2 (N4190, N4184, N1669);
nand NAND2 (N4191, N4160, N3253);
xor XOR2 (N4192, N4188, N1269);
xor XOR2 (N4193, N4191, N355);
nor NOR3 (N4194, N4169, N2731, N3060);
nor NOR4 (N4195, N4189, N3260, N451, N4175);
nand NAND4 (N4196, N4182, N1042, N1127, N3681);
or OR4 (N4197, N4181, N3812, N3221, N1411);
xor XOR2 (N4198, N4174, N3530);
xor XOR2 (N4199, N4193, N3397);
and AND2 (N4200, N4190, N3614);
buf BUF1 (N4201, N4196);
or OR3 (N4202, N4195, N577, N3579);
not NOT1 (N4203, N4194);
xor XOR2 (N4204, N4192, N2211);
nand NAND2 (N4205, N4202, N2779);
nor NOR2 (N4206, N4199, N1082);
nand NAND3 (N4207, N4197, N2647, N1328);
nor NOR2 (N4208, N4206, N2244);
buf BUF1 (N4209, N4203);
or OR3 (N4210, N4201, N363, N1526);
and AND4 (N4211, N4210, N2234, N1495, N2800);
buf BUF1 (N4212, N4209);
buf BUF1 (N4213, N4198);
and AND4 (N4214, N4211, N3236, N464, N1793);
nor NOR2 (N4215, N4208, N423);
and AND3 (N4216, N4205, N1165, N1851);
xor XOR2 (N4217, N4180, N2048);
not NOT1 (N4218, N4212);
nand NAND3 (N4219, N4213, N4118, N3116);
nor NOR2 (N4220, N4215, N311);
nand NAND4 (N4221, N4217, N3977, N3919, N1273);
not NOT1 (N4222, N4183);
xor XOR2 (N4223, N4221, N409);
xor XOR2 (N4224, N4223, N775);
not NOT1 (N4225, N4214);
nand NAND2 (N4226, N4224, N3589);
and AND2 (N4227, N4219, N864);
nand NAND4 (N4228, N4225, N376, N3566, N1146);
buf BUF1 (N4229, N4222);
and AND3 (N4230, N4200, N3578, N4054);
and AND2 (N4231, N4218, N4174);
and AND4 (N4232, N4204, N3403, N1928, N1353);
nand NAND3 (N4233, N4230, N69, N705);
not NOT1 (N4234, N4226);
not NOT1 (N4235, N4233);
and AND3 (N4236, N4228, N2000, N3779);
nand NAND4 (N4237, N4216, N1424, N1457, N3920);
nor NOR3 (N4238, N4229, N114, N3073);
nor NOR3 (N4239, N4227, N2583, N1546);
not NOT1 (N4240, N4238);
buf BUF1 (N4241, N4239);
buf BUF1 (N4242, N4240);
nor NOR4 (N4243, N4242, N3341, N2370, N3729);
nand NAND3 (N4244, N4234, N3408, N1941);
nor NOR4 (N4245, N4231, N3148, N590, N1714);
and AND4 (N4246, N4220, N552, N942, N2894);
and AND4 (N4247, N4243, N4057, N34, N2544);
and AND3 (N4248, N4247, N4204, N2872);
buf BUF1 (N4249, N4241);
or OR3 (N4250, N4244, N2003, N232);
xor XOR2 (N4251, N4207, N390);
not NOT1 (N4252, N4249);
and AND3 (N4253, N4232, N413, N2734);
xor XOR2 (N4254, N4245, N1296);
nor NOR3 (N4255, N4251, N1870, N3570);
xor XOR2 (N4256, N4237, N1983);
buf BUF1 (N4257, N4235);
not NOT1 (N4258, N4254);
not NOT1 (N4259, N4252);
nor NOR2 (N4260, N4248, N45);
nor NOR3 (N4261, N4250, N2882, N2269);
nand NAND4 (N4262, N4259, N1347, N2260, N291);
and AND4 (N4263, N4258, N2469, N1093, N2535);
and AND2 (N4264, N4246, N2884);
not NOT1 (N4265, N4263);
not NOT1 (N4266, N4257);
nand NAND3 (N4267, N4260, N2975, N3183);
and AND2 (N4268, N4255, N1964);
buf BUF1 (N4269, N4268);
or OR3 (N4270, N4265, N3482, N3116);
xor XOR2 (N4271, N4256, N3765);
and AND2 (N4272, N4269, N3169);
buf BUF1 (N4273, N4267);
xor XOR2 (N4274, N4272, N3292);
and AND3 (N4275, N4264, N3670, N2242);
xor XOR2 (N4276, N4275, N291);
and AND2 (N4277, N4253, N693);
nor NOR2 (N4278, N4236, N1137);
nand NAND2 (N4279, N4278, N4160);
and AND4 (N4280, N4271, N3894, N2280, N3526);
and AND3 (N4281, N4274, N774, N1958);
xor XOR2 (N4282, N4277, N914);
buf BUF1 (N4283, N4266);
xor XOR2 (N4284, N4276, N3437);
and AND4 (N4285, N4281, N2323, N3819, N3656);
and AND4 (N4286, N4282, N3390, N2702, N3254);
or OR3 (N4287, N4283, N1026, N3940);
nor NOR2 (N4288, N4261, N2450);
not NOT1 (N4289, N4286);
not NOT1 (N4290, N4273);
nand NAND2 (N4291, N4279, N1177);
xor XOR2 (N4292, N4270, N1326);
or OR4 (N4293, N4287, N3198, N4063, N597);
nor NOR4 (N4294, N4288, N3015, N2937, N2135);
not NOT1 (N4295, N4291);
buf BUF1 (N4296, N4290);
buf BUF1 (N4297, N4285);
buf BUF1 (N4298, N4280);
nand NAND2 (N4299, N4295, N215);
or OR2 (N4300, N4293, N1950);
and AND3 (N4301, N4300, N1859, N2378);
xor XOR2 (N4302, N4301, N2607);
or OR4 (N4303, N4292, N769, N1276, N2382);
nor NOR3 (N4304, N4296, N2989, N3549);
buf BUF1 (N4305, N4302);
or OR4 (N4306, N4304, N10, N2578, N3726);
or OR3 (N4307, N4303, N1770, N2478);
xor XOR2 (N4308, N4305, N3264);
and AND4 (N4309, N4307, N1928, N1809, N2915);
or OR4 (N4310, N4299, N4238, N737, N4129);
buf BUF1 (N4311, N4309);
buf BUF1 (N4312, N4284);
or OR3 (N4313, N4306, N998, N261);
or OR3 (N4314, N4289, N3080, N1540);
buf BUF1 (N4315, N4310);
not NOT1 (N4316, N4312);
xor XOR2 (N4317, N4308, N2889);
and AND3 (N4318, N4315, N2444, N3238);
buf BUF1 (N4319, N4311);
and AND2 (N4320, N4319, N2465);
nand NAND2 (N4321, N4262, N1441);
nand NAND4 (N4322, N4313, N1095, N2657, N738);
buf BUF1 (N4323, N4297);
or OR4 (N4324, N4323, N3352, N4200, N4245);
nor NOR3 (N4325, N4318, N1703, N2348);
nand NAND2 (N4326, N4324, N4052);
and AND3 (N4327, N4326, N1422, N479);
xor XOR2 (N4328, N4327, N2318);
not NOT1 (N4329, N4314);
or OR3 (N4330, N4329, N200, N3050);
xor XOR2 (N4331, N4317, N4058);
and AND3 (N4332, N4294, N3766, N2885);
and AND4 (N4333, N4331, N3287, N3534, N4084);
and AND4 (N4334, N4332, N1358, N2350, N3483);
or OR3 (N4335, N4328, N2936, N4161);
nor NOR4 (N4336, N4333, N1412, N3070, N3550);
nor NOR4 (N4337, N4325, N3871, N1611, N1494);
or OR3 (N4338, N4322, N1645, N4077);
nand NAND3 (N4339, N4334, N929, N4280);
xor XOR2 (N4340, N4330, N1843);
or OR3 (N4341, N4338, N1309, N3101);
nand NAND4 (N4342, N4339, N525, N3353, N1528);
nand NAND3 (N4343, N4336, N3194, N4076);
or OR3 (N4344, N4321, N3190, N220);
or OR3 (N4345, N4341, N2855, N1654);
nor NOR4 (N4346, N4320, N2917, N554, N2979);
or OR2 (N4347, N4346, N1857);
nor NOR2 (N4348, N4344, N3918);
not NOT1 (N4349, N4345);
nor NOR2 (N4350, N4298, N407);
nand NAND3 (N4351, N4347, N3013, N261);
not NOT1 (N4352, N4337);
and AND4 (N4353, N4351, N2932, N3820, N291);
nor NOR3 (N4354, N4349, N621, N4169);
or OR3 (N4355, N4353, N248, N259);
not NOT1 (N4356, N4340);
nor NOR4 (N4357, N4335, N1868, N1716, N29);
not NOT1 (N4358, N4355);
or OR2 (N4359, N4357, N3811);
buf BUF1 (N4360, N4316);
not NOT1 (N4361, N4352);
buf BUF1 (N4362, N4358);
or OR3 (N4363, N4343, N190, N638);
nor NOR4 (N4364, N4359, N2682, N2266, N3103);
buf BUF1 (N4365, N4354);
and AND4 (N4366, N4350, N1101, N1642, N2404);
xor XOR2 (N4367, N4342, N3779);
not NOT1 (N4368, N4365);
nor NOR2 (N4369, N4364, N3820);
and AND4 (N4370, N4366, N3624, N4172, N2094);
xor XOR2 (N4371, N4356, N2479);
not NOT1 (N4372, N4360);
and AND3 (N4373, N4370, N1594, N2142);
nor NOR3 (N4374, N4367, N1178, N3940);
xor XOR2 (N4375, N4374, N2011);
or OR4 (N4376, N4369, N1053, N2112, N602);
not NOT1 (N4377, N4363);
nor NOR3 (N4378, N4377, N1981, N2324);
and AND4 (N4379, N4368, N779, N3568, N2372);
xor XOR2 (N4380, N4373, N4252);
not NOT1 (N4381, N4376);
and AND2 (N4382, N4381, N1123);
not NOT1 (N4383, N4372);
and AND3 (N4384, N4378, N4306, N1611);
or OR2 (N4385, N4348, N242);
xor XOR2 (N4386, N4384, N4042);
nand NAND2 (N4387, N4386, N3530);
not NOT1 (N4388, N4375);
nand NAND3 (N4389, N4380, N3004, N3831);
or OR3 (N4390, N4387, N3451, N2482);
nand NAND4 (N4391, N4389, N757, N299, N4191);
and AND2 (N4392, N4362, N2064);
xor XOR2 (N4393, N4392, N209);
xor XOR2 (N4394, N4388, N1643);
xor XOR2 (N4395, N4385, N2789);
nor NOR3 (N4396, N4383, N4356, N1263);
and AND4 (N4397, N4382, N4167, N4086, N2716);
nand NAND2 (N4398, N4393, N3440);
nand NAND4 (N4399, N4398, N3981, N4205, N873);
or OR3 (N4400, N4379, N3464, N1553);
and AND4 (N4401, N4391, N3874, N3454, N2251);
nor NOR3 (N4402, N4390, N2606, N2673);
buf BUF1 (N4403, N4400);
xor XOR2 (N4404, N4371, N3474);
not NOT1 (N4405, N4394);
or OR3 (N4406, N4403, N602, N2712);
or OR4 (N4407, N4361, N1928, N320, N4320);
and AND3 (N4408, N4401, N1480, N3597);
not NOT1 (N4409, N4402);
nand NAND4 (N4410, N4399, N793, N605, N2608);
buf BUF1 (N4411, N4404);
or OR2 (N4412, N4410, N2926);
xor XOR2 (N4413, N4411, N199);
nor NOR4 (N4414, N4395, N3396, N3092, N2134);
not NOT1 (N4415, N4405);
buf BUF1 (N4416, N4396);
nand NAND3 (N4417, N4412, N2925, N1396);
or OR3 (N4418, N4407, N2832, N829);
or OR2 (N4419, N4406, N4035);
nor NOR3 (N4420, N4408, N1979, N3961);
not NOT1 (N4421, N4416);
buf BUF1 (N4422, N4409);
buf BUF1 (N4423, N4414);
and AND3 (N4424, N4397, N3297, N1446);
and AND2 (N4425, N4423, N2173);
xor XOR2 (N4426, N4419, N800);
not NOT1 (N4427, N4425);
and AND4 (N4428, N4415, N118, N1871, N2060);
nor NOR4 (N4429, N4422, N4397, N2540, N2499);
buf BUF1 (N4430, N4428);
and AND3 (N4431, N4420, N433, N1430);
xor XOR2 (N4432, N4430, N4335);
xor XOR2 (N4433, N4413, N363);
buf BUF1 (N4434, N4417);
or OR2 (N4435, N4424, N511);
not NOT1 (N4436, N4421);
xor XOR2 (N4437, N4426, N1056);
buf BUF1 (N4438, N4431);
and AND3 (N4439, N4427, N1890, N708);
and AND4 (N4440, N4435, N3605, N1443, N4422);
xor XOR2 (N4441, N4439, N1532);
nor NOR2 (N4442, N4437, N3939);
not NOT1 (N4443, N4433);
and AND4 (N4444, N4440, N2589, N830, N189);
and AND4 (N4445, N4438, N1805, N3948, N436);
nor NOR3 (N4446, N4444, N2905, N2010);
and AND2 (N4447, N4442, N520);
nor NOR4 (N4448, N4445, N3515, N3370, N3804);
buf BUF1 (N4449, N4436);
nand NAND4 (N4450, N4418, N4395, N1021, N1536);
buf BUF1 (N4451, N4450);
not NOT1 (N4452, N4447);
nor NOR3 (N4453, N4441, N2750, N804);
nand NAND4 (N4454, N4451, N1587, N794, N3680);
buf BUF1 (N4455, N4446);
and AND4 (N4456, N4454, N4135, N1175, N3523);
xor XOR2 (N4457, N4443, N3127);
nand NAND3 (N4458, N4452, N3778, N1722);
or OR3 (N4459, N4448, N3486, N3992);
nor NOR4 (N4460, N4457, N1747, N3260, N623);
or OR3 (N4461, N4455, N787, N2285);
buf BUF1 (N4462, N4458);
and AND3 (N4463, N4456, N3965, N746);
buf BUF1 (N4464, N4434);
not NOT1 (N4465, N4461);
xor XOR2 (N4466, N4429, N284);
buf BUF1 (N4467, N4453);
buf BUF1 (N4468, N4463);
nand NAND4 (N4469, N4459, N3713, N3409, N2242);
or OR4 (N4470, N4469, N3632, N2608, N3138);
buf BUF1 (N4471, N4468);
not NOT1 (N4472, N4466);
nand NAND2 (N4473, N4462, N1380);
not NOT1 (N4474, N4460);
not NOT1 (N4475, N4472);
xor XOR2 (N4476, N4467, N4072);
nor NOR2 (N4477, N4465, N1163);
not NOT1 (N4478, N4449);
nor NOR4 (N4479, N4477, N1963, N366, N833);
not NOT1 (N4480, N4471);
and AND3 (N4481, N4475, N2233, N83);
or OR4 (N4482, N4476, N1679, N2268, N4089);
nor NOR2 (N4483, N4470, N58);
buf BUF1 (N4484, N4432);
and AND4 (N4485, N4478, N2446, N3658, N3054);
nand NAND4 (N4486, N4479, N3560, N1077, N1336);
not NOT1 (N4487, N4473);
nor NOR3 (N4488, N4485, N2128, N1194);
not NOT1 (N4489, N4483);
xor XOR2 (N4490, N4486, N2419);
nor NOR2 (N4491, N4482, N3463);
not NOT1 (N4492, N4464);
and AND3 (N4493, N4484, N1565, N16);
buf BUF1 (N4494, N4488);
not NOT1 (N4495, N4487);
buf BUF1 (N4496, N4489);
and AND3 (N4497, N4492, N1847, N3862);
xor XOR2 (N4498, N4497, N3997);
not NOT1 (N4499, N4490);
not NOT1 (N4500, N4491);
xor XOR2 (N4501, N4480, N3055);
nor NOR3 (N4502, N4493, N897, N3082);
nor NOR3 (N4503, N4474, N4244, N885);
buf BUF1 (N4504, N4501);
not NOT1 (N4505, N4502);
buf BUF1 (N4506, N4496);
not NOT1 (N4507, N4500);
xor XOR2 (N4508, N4495, N2857);
and AND2 (N4509, N4481, N1296);
nand NAND2 (N4510, N4498, N3700);
buf BUF1 (N4511, N4509);
nand NAND4 (N4512, N4505, N4024, N1851, N3346);
and AND4 (N4513, N4504, N321, N1751, N2353);
not NOT1 (N4514, N4503);
buf BUF1 (N4515, N4512);
not NOT1 (N4516, N4510);
nor NOR4 (N4517, N4513, N3064, N4038, N3755);
and AND2 (N4518, N4494, N4219);
or OR3 (N4519, N4508, N4328, N1206);
nor NOR3 (N4520, N4519, N1599, N4142);
xor XOR2 (N4521, N4511, N391);
buf BUF1 (N4522, N4499);
or OR2 (N4523, N4515, N2642);
buf BUF1 (N4524, N4523);
or OR3 (N4525, N4521, N2878, N1418);
not NOT1 (N4526, N4507);
or OR3 (N4527, N4518, N4152, N1863);
xor XOR2 (N4528, N4525, N762);
or OR3 (N4529, N4524, N2826, N1569);
nand NAND3 (N4530, N4516, N2896, N350);
not NOT1 (N4531, N4529);
xor XOR2 (N4532, N4517, N2719);
nand NAND3 (N4533, N4522, N1078, N2560);
or OR4 (N4534, N4533, N4265, N1028, N4143);
buf BUF1 (N4535, N4531);
nor NOR4 (N4536, N4528, N1344, N2317, N3818);
not NOT1 (N4537, N4532);
and AND2 (N4538, N4527, N3468);
xor XOR2 (N4539, N4538, N2346);
buf BUF1 (N4540, N4514);
nor NOR2 (N4541, N4534, N3634);
and AND3 (N4542, N4540, N901, N3088);
not NOT1 (N4543, N4530);
nor NOR3 (N4544, N4526, N4480, N3449);
nand NAND2 (N4545, N4542, N3051);
nor NOR4 (N4546, N4543, N286, N1595, N1702);
not NOT1 (N4547, N4539);
nand NAND4 (N4548, N4520, N1083, N1262, N475);
buf BUF1 (N4549, N4541);
and AND4 (N4550, N4535, N4205, N1243, N4132);
not NOT1 (N4551, N4537);
and AND2 (N4552, N4544, N1733);
buf BUF1 (N4553, N4552);
and AND4 (N4554, N4549, N2993, N4278, N4062);
buf BUF1 (N4555, N4548);
and AND4 (N4556, N4550, N132, N452, N977);
nor NOR2 (N4557, N4551, N1120);
not NOT1 (N4558, N4536);
and AND4 (N4559, N4554, N4013, N2679, N1781);
xor XOR2 (N4560, N4555, N2967);
not NOT1 (N4561, N4547);
and AND4 (N4562, N4545, N2542, N3964, N208);
and AND3 (N4563, N4558, N3185, N3091);
nand NAND3 (N4564, N4546, N285, N1341);
or OR3 (N4565, N4559, N2014, N909);
buf BUF1 (N4566, N4561);
and AND2 (N4567, N4563, N871);
nor NOR3 (N4568, N4564, N4182, N846);
not NOT1 (N4569, N4557);
nor NOR4 (N4570, N4506, N210, N562, N1060);
nand NAND2 (N4571, N4556, N548);
nand NAND4 (N4572, N4565, N3343, N4545, N25);
xor XOR2 (N4573, N4571, N736);
buf BUF1 (N4574, N4553);
nor NOR2 (N4575, N4562, N4224);
and AND3 (N4576, N4560, N4175, N1562);
nor NOR2 (N4577, N4572, N859);
or OR4 (N4578, N4570, N2573, N3900, N2205);
nand NAND2 (N4579, N4574, N4130);
and AND3 (N4580, N4573, N636, N1411);
nand NAND3 (N4581, N4576, N2374, N3386);
or OR2 (N4582, N4580, N2812);
or OR2 (N4583, N4575, N3209);
buf BUF1 (N4584, N4583);
nor NOR4 (N4585, N4584, N4191, N2200, N2079);
nor NOR4 (N4586, N4579, N3116, N272, N349);
buf BUF1 (N4587, N4566);
nand NAND2 (N4588, N4578, N85);
or OR2 (N4589, N4587, N4492);
not NOT1 (N4590, N4569);
buf BUF1 (N4591, N4588);
not NOT1 (N4592, N4582);
xor XOR2 (N4593, N4567, N3217);
buf BUF1 (N4594, N4593);
nand NAND3 (N4595, N4581, N2825, N639);
buf BUF1 (N4596, N4585);
nand NAND4 (N4597, N4586, N791, N2239, N1263);
or OR4 (N4598, N4568, N4052, N3822, N4579);
and AND2 (N4599, N4590, N810);
nor NOR4 (N4600, N4592, N4216, N4162, N81);
not NOT1 (N4601, N4596);
or OR2 (N4602, N4600, N221);
not NOT1 (N4603, N4599);
xor XOR2 (N4604, N4603, N2268);
or OR4 (N4605, N4601, N233, N366, N3290);
nand NAND2 (N4606, N4591, N2385);
buf BUF1 (N4607, N4594);
or OR2 (N4608, N4595, N429);
xor XOR2 (N4609, N4605, N3261);
and AND3 (N4610, N4607, N3898, N2833);
or OR4 (N4611, N4602, N40, N3842, N3475);
nand NAND3 (N4612, N4604, N2566, N351);
xor XOR2 (N4613, N4608, N776);
nand NAND2 (N4614, N4612, N1381);
buf BUF1 (N4615, N4597);
buf BUF1 (N4616, N4609);
nand NAND2 (N4617, N4606, N2671);
nand NAND3 (N4618, N4611, N2647, N1065);
xor XOR2 (N4619, N4577, N1057);
buf BUF1 (N4620, N4610);
nor NOR3 (N4621, N4616, N1692, N4237);
nor NOR3 (N4622, N4619, N4121, N3931);
nor NOR3 (N4623, N4615, N2445, N3704);
nor NOR3 (N4624, N4621, N1695, N1453);
not NOT1 (N4625, N4617);
not NOT1 (N4626, N4624);
buf BUF1 (N4627, N4589);
or OR3 (N4628, N4614, N1494, N1473);
nand NAND4 (N4629, N4618, N2779, N898, N426);
or OR2 (N4630, N4622, N4578);
buf BUF1 (N4631, N4627);
xor XOR2 (N4632, N4629, N4275);
xor XOR2 (N4633, N4623, N367);
not NOT1 (N4634, N4625);
not NOT1 (N4635, N4633);
and AND3 (N4636, N4598, N990, N2066);
nor NOR3 (N4637, N4636, N3791, N3924);
and AND2 (N4638, N4620, N1204);
nor NOR4 (N4639, N4613, N4254, N1587, N2465);
buf BUF1 (N4640, N4632);
nand NAND4 (N4641, N4640, N2068, N2869, N1410);
not NOT1 (N4642, N4637);
buf BUF1 (N4643, N4626);
and AND4 (N4644, N4631, N4630, N3622, N4574);
not NOT1 (N4645, N2405);
buf BUF1 (N4646, N4638);
or OR2 (N4647, N4628, N3666);
nor NOR4 (N4648, N4635, N82, N773, N3071);
nand NAND3 (N4649, N4645, N907, N2298);
or OR2 (N4650, N4643, N3362);
xor XOR2 (N4651, N4641, N1055);
or OR2 (N4652, N4647, N430);
and AND2 (N4653, N4639, N2470);
nand NAND4 (N4654, N4634, N3719, N2552, N451);
not NOT1 (N4655, N4651);
xor XOR2 (N4656, N4654, N2885);
nand NAND2 (N4657, N4652, N1775);
or OR3 (N4658, N4657, N1855, N2031);
nand NAND3 (N4659, N4653, N264, N2945);
buf BUF1 (N4660, N4646);
nand NAND3 (N4661, N4660, N4264, N1755);
not NOT1 (N4662, N4648);
buf BUF1 (N4663, N4662);
nor NOR2 (N4664, N4649, N4188);
and AND4 (N4665, N4644, N1815, N3485, N4445);
not NOT1 (N4666, N4664);
or OR3 (N4667, N4656, N675, N4408);
or OR2 (N4668, N4650, N2580);
buf BUF1 (N4669, N4665);
and AND2 (N4670, N4667, N2554);
or OR4 (N4671, N4663, N1055, N2234, N2376);
or OR4 (N4672, N4655, N2245, N619, N2095);
buf BUF1 (N4673, N4670);
nor NOR4 (N4674, N4659, N4594, N3065, N1331);
not NOT1 (N4675, N4661);
not NOT1 (N4676, N4674);
and AND2 (N4677, N4672, N2576);
and AND4 (N4678, N4642, N499, N1846, N17);
or OR3 (N4679, N4671, N4591, N4334);
nor NOR2 (N4680, N4676, N2722);
nand NAND2 (N4681, N4669, N1984);
or OR4 (N4682, N4678, N1806, N1428, N4259);
nor NOR2 (N4683, N4675, N790);
xor XOR2 (N4684, N4683, N3559);
nand NAND2 (N4685, N4684, N4334);
and AND2 (N4686, N4673, N1178);
nor NOR3 (N4687, N4686, N3236, N2402);
and AND2 (N4688, N4680, N265);
xor XOR2 (N4689, N4687, N3624);
not NOT1 (N4690, N4689);
and AND4 (N4691, N4681, N599, N3480, N4044);
and AND3 (N4692, N4685, N2000, N2259);
nor NOR2 (N4693, N4682, N2850);
nand NAND2 (N4694, N4690, N4364);
and AND4 (N4695, N4679, N2001, N4364, N1551);
or OR4 (N4696, N4695, N3498, N442, N2214);
not NOT1 (N4697, N4688);
buf BUF1 (N4698, N4696);
nor NOR2 (N4699, N4658, N958);
or OR3 (N4700, N4692, N1923, N424);
or OR3 (N4701, N4698, N812, N188);
nand NAND4 (N4702, N4691, N512, N379, N2387);
buf BUF1 (N4703, N4668);
xor XOR2 (N4704, N4699, N1700);
buf BUF1 (N4705, N4703);
xor XOR2 (N4706, N4704, N3834);
nand NAND2 (N4707, N4701, N792);
and AND3 (N4708, N4666, N1381, N3840);
buf BUF1 (N4709, N4702);
xor XOR2 (N4710, N4707, N973);
buf BUF1 (N4711, N4700);
xor XOR2 (N4712, N4710, N790);
nor NOR4 (N4713, N4706, N3965, N1536, N148);
not NOT1 (N4714, N4713);
buf BUF1 (N4715, N4677);
xor XOR2 (N4716, N4711, N3508);
buf BUF1 (N4717, N4712);
xor XOR2 (N4718, N4714, N1209);
buf BUF1 (N4719, N4697);
and AND2 (N4720, N4717, N544);
nor NOR3 (N4721, N4719, N3385, N4108);
and AND3 (N4722, N4721, N1437, N4065);
or OR3 (N4723, N4708, N3331, N3044);
and AND2 (N4724, N4716, N1064);
or OR2 (N4725, N4694, N3872);
and AND3 (N4726, N4724, N767, N592);
nand NAND2 (N4727, N4709, N2856);
or OR4 (N4728, N4715, N3872, N4415, N3690);
buf BUF1 (N4729, N4727);
buf BUF1 (N4730, N4726);
nor NOR4 (N4731, N4729, N3021, N4052, N3722);
xor XOR2 (N4732, N4730, N1564);
not NOT1 (N4733, N4722);
not NOT1 (N4734, N4693);
nor NOR4 (N4735, N4723, N4066, N3043, N147);
or OR2 (N4736, N4728, N2378);
xor XOR2 (N4737, N4731, N3657);
nand NAND3 (N4738, N4718, N3873, N2884);
not NOT1 (N4739, N4734);
nand NAND3 (N4740, N4735, N383, N531);
or OR3 (N4741, N4705, N2338, N3843);
or OR2 (N4742, N4738, N2675);
and AND3 (N4743, N4742, N3323, N3863);
xor XOR2 (N4744, N4741, N4458);
not NOT1 (N4745, N4732);
xor XOR2 (N4746, N4736, N1147);
buf BUF1 (N4747, N4739);
xor XOR2 (N4748, N4737, N3429);
nand NAND4 (N4749, N4744, N182, N1416, N4020);
and AND2 (N4750, N4740, N742);
and AND4 (N4751, N4747, N1713, N1888, N3387);
nor NOR3 (N4752, N4749, N4581, N1698);
not NOT1 (N4753, N4746);
or OR4 (N4754, N4752, N1509, N4558, N3988);
and AND2 (N4755, N4745, N305);
nand NAND2 (N4756, N4720, N798);
not NOT1 (N4757, N4733);
and AND4 (N4758, N4725, N875, N1155, N378);
xor XOR2 (N4759, N4753, N3022);
nor NOR3 (N4760, N4757, N3495, N2183);
and AND4 (N4761, N4759, N2582, N4161, N4392);
or OR2 (N4762, N4758, N2222);
xor XOR2 (N4763, N4761, N3440);
nand NAND2 (N4764, N4763, N2358);
or OR2 (N4765, N4755, N4312);
nor NOR2 (N4766, N4743, N2445);
buf BUF1 (N4767, N4766);
buf BUF1 (N4768, N4765);
nand NAND2 (N4769, N4760, N2908);
or OR2 (N4770, N4754, N3341);
and AND4 (N4771, N4756, N2696, N1859, N1057);
not NOT1 (N4772, N4768);
nor NOR3 (N4773, N4751, N2596, N33);
nor NOR2 (N4774, N4767, N3105);
and AND3 (N4775, N4762, N2424, N3728);
nor NOR3 (N4776, N4764, N3844, N2920);
or OR3 (N4777, N4750, N1253, N564);
xor XOR2 (N4778, N4769, N1668);
nor NOR4 (N4779, N4774, N1396, N755, N363);
not NOT1 (N4780, N4776);
or OR4 (N4781, N4780, N3976, N4247, N232);
and AND4 (N4782, N4778, N2785, N2123, N452);
buf BUF1 (N4783, N4772);
nand NAND3 (N4784, N4779, N3665, N1803);
nor NOR2 (N4785, N4784, N474);
or OR4 (N4786, N4771, N4058, N2379, N4195);
not NOT1 (N4787, N4777);
nor NOR2 (N4788, N4775, N589);
and AND4 (N4789, N4783, N3074, N3889, N4651);
nor NOR3 (N4790, N4770, N942, N983);
xor XOR2 (N4791, N4787, N4510);
or OR4 (N4792, N4748, N3287, N3259, N3340);
buf BUF1 (N4793, N4788);
nor NOR3 (N4794, N4793, N1645, N4497);
not NOT1 (N4795, N4786);
or OR4 (N4796, N4773, N4738, N3950, N4420);
or OR4 (N4797, N4794, N4515, N3474, N2894);
and AND3 (N4798, N4789, N3607, N3730);
and AND4 (N4799, N4791, N2865, N282, N944);
nand NAND3 (N4800, N4785, N1643, N1793);
or OR2 (N4801, N4799, N4437);
buf BUF1 (N4802, N4792);
nand NAND2 (N4803, N4801, N647);
or OR4 (N4804, N4802, N1328, N860, N4749);
nor NOR3 (N4805, N4804, N696, N4244);
nor NOR3 (N4806, N4795, N2511, N4543);
not NOT1 (N4807, N4798);
nor NOR4 (N4808, N4796, N2383, N399, N361);
and AND3 (N4809, N4790, N3912, N2353);
nor NOR3 (N4810, N4803, N3321, N188);
or OR3 (N4811, N4797, N2070, N3544);
or OR3 (N4812, N4808, N1682, N3090);
nand NAND2 (N4813, N4781, N300);
nor NOR2 (N4814, N4810, N1248);
xor XOR2 (N4815, N4814, N3548);
and AND2 (N4816, N4809, N4771);
nand NAND3 (N4817, N4806, N3587, N2915);
buf BUF1 (N4818, N4813);
and AND4 (N4819, N4816, N4108, N4691, N1197);
nor NOR2 (N4820, N4817, N1300);
nor NOR4 (N4821, N4818, N2566, N4807, N3185);
xor XOR2 (N4822, N618, N2364);
buf BUF1 (N4823, N4822);
nor NOR3 (N4824, N4782, N3589, N1966);
and AND3 (N4825, N4800, N4792, N3372);
buf BUF1 (N4826, N4820);
not NOT1 (N4827, N4821);
or OR3 (N4828, N4805, N4326, N4004);
or OR2 (N4829, N4811, N4825);
xor XOR2 (N4830, N4590, N3173);
not NOT1 (N4831, N4827);
xor XOR2 (N4832, N4823, N3499);
xor XOR2 (N4833, N4824, N1294);
or OR4 (N4834, N4833, N4327, N1630, N2229);
or OR2 (N4835, N4812, N1612);
not NOT1 (N4836, N4819);
nor NOR2 (N4837, N4815, N4669);
buf BUF1 (N4838, N4828);
xor XOR2 (N4839, N4829, N2012);
xor XOR2 (N4840, N4831, N224);
not NOT1 (N4841, N4830);
and AND2 (N4842, N4837, N424);
nor NOR3 (N4843, N4832, N1503, N4658);
nor NOR2 (N4844, N4838, N1966);
and AND4 (N4845, N4834, N1715, N3338, N2065);
nand NAND2 (N4846, N4839, N634);
nor NOR4 (N4847, N4845, N1115, N118, N3103);
nand NAND3 (N4848, N4846, N2016, N1001);
not NOT1 (N4849, N4836);
or OR4 (N4850, N4826, N2829, N3657, N2999);
nand NAND4 (N4851, N4835, N3962, N4512, N1746);
nor NOR2 (N4852, N4848, N1153);
not NOT1 (N4853, N4849);
nand NAND4 (N4854, N4850, N500, N1398, N2257);
nor NOR2 (N4855, N4842, N2141);
buf BUF1 (N4856, N4844);
xor XOR2 (N4857, N4853, N52);
and AND2 (N4858, N4854, N2878);
xor XOR2 (N4859, N4840, N4465);
and AND2 (N4860, N4851, N1164);
not NOT1 (N4861, N4860);
nor NOR3 (N4862, N4859, N1590, N1314);
and AND4 (N4863, N4843, N2696, N4098, N3725);
xor XOR2 (N4864, N4861, N4779);
nor NOR4 (N4865, N4864, N3478, N605, N2779);
nor NOR3 (N4866, N4841, N2333, N3954);
and AND4 (N4867, N4847, N291, N2316, N3988);
not NOT1 (N4868, N4857);
xor XOR2 (N4869, N4868, N3655);
xor XOR2 (N4870, N4852, N1719);
not NOT1 (N4871, N4867);
nor NOR3 (N4872, N4855, N2607, N477);
nor NOR4 (N4873, N4866, N289, N4255, N3986);
not NOT1 (N4874, N4872);
nor NOR2 (N4875, N4862, N1084);
and AND4 (N4876, N4865, N1806, N1319, N4293);
and AND4 (N4877, N4869, N3162, N3770, N1812);
nand NAND3 (N4878, N4870, N3882, N1077);
xor XOR2 (N4879, N4874, N4252);
nor NOR3 (N4880, N4871, N2517, N1334);
and AND4 (N4881, N4875, N1941, N1263, N2168);
not NOT1 (N4882, N4877);
xor XOR2 (N4883, N4880, N531);
not NOT1 (N4884, N4878);
xor XOR2 (N4885, N4879, N651);
or OR3 (N4886, N4885, N1746, N708);
buf BUF1 (N4887, N4884);
xor XOR2 (N4888, N4873, N416);
nand NAND3 (N4889, N4876, N2021, N4637);
buf BUF1 (N4890, N4886);
nand NAND4 (N4891, N4856, N4279, N968, N1729);
nand NAND3 (N4892, N4889, N102, N670);
and AND2 (N4893, N4858, N2436);
buf BUF1 (N4894, N4890);
nand NAND4 (N4895, N4882, N2053, N2453, N2459);
buf BUF1 (N4896, N4863);
xor XOR2 (N4897, N4888, N4304);
and AND2 (N4898, N4892, N1306);
and AND3 (N4899, N4891, N3688, N585);
nand NAND3 (N4900, N4893, N945, N74);
and AND3 (N4901, N4883, N1692, N3008);
nor NOR2 (N4902, N4899, N3545);
and AND4 (N4903, N4887, N3330, N3637, N4383);
nor NOR4 (N4904, N4903, N477, N1268, N3060);
nor NOR4 (N4905, N4881, N842, N3129, N1461);
nand NAND2 (N4906, N4897, N2783);
nand NAND4 (N4907, N4902, N112, N3479, N2672);
and AND3 (N4908, N4900, N1566, N3043);
nand NAND4 (N4909, N4907, N3524, N307, N4291);
nand NAND2 (N4910, N4901, N3590);
and AND4 (N4911, N4895, N636, N2835, N2550);
nand NAND4 (N4912, N4911, N3285, N2719, N1660);
nand NAND4 (N4913, N4910, N527, N590, N980);
not NOT1 (N4914, N4906);
xor XOR2 (N4915, N4912, N2228);
buf BUF1 (N4916, N4914);
nor NOR4 (N4917, N4904, N707, N1770, N2660);
nor NOR2 (N4918, N4913, N839);
or OR3 (N4919, N4896, N2680, N4322);
and AND2 (N4920, N4905, N1);
nand NAND3 (N4921, N4918, N3547, N105);
nand NAND2 (N4922, N4919, N3997);
or OR3 (N4923, N4921, N1074, N1096);
nand NAND2 (N4924, N4916, N1939);
not NOT1 (N4925, N4924);
or OR2 (N4926, N4894, N2264);
not NOT1 (N4927, N4908);
and AND4 (N4928, N4917, N4696, N1722, N3198);
nand NAND2 (N4929, N4925, N4218);
xor XOR2 (N4930, N4927, N2956);
nand NAND4 (N4931, N4926, N3485, N3996, N1398);
or OR2 (N4932, N4922, N4851);
xor XOR2 (N4933, N4931, N3384);
not NOT1 (N4934, N4928);
nor NOR4 (N4935, N4898, N3678, N4420, N542);
and AND2 (N4936, N4934, N2430);
nor NOR4 (N4937, N4936, N4738, N4733, N3885);
not NOT1 (N4938, N4929);
and AND3 (N4939, N4920, N3282, N3389);
not NOT1 (N4940, N4923);
and AND4 (N4941, N4933, N454, N2097, N1242);
not NOT1 (N4942, N4941);
and AND2 (N4943, N4930, N2164);
nor NOR3 (N4944, N4939, N801, N3910);
not NOT1 (N4945, N4944);
nor NOR4 (N4946, N4945, N3910, N4798, N281);
buf BUF1 (N4947, N4942);
xor XOR2 (N4948, N4943, N188);
or OR4 (N4949, N4947, N4271, N479, N2428);
buf BUF1 (N4950, N4940);
and AND3 (N4951, N4932, N2320, N4816);
not NOT1 (N4952, N4949);
xor XOR2 (N4953, N4946, N834);
and AND3 (N4954, N4915, N4933, N2237);
nor NOR3 (N4955, N4951, N4880, N2277);
buf BUF1 (N4956, N4953);
not NOT1 (N4957, N4948);
not NOT1 (N4958, N4909);
not NOT1 (N4959, N4958);
buf BUF1 (N4960, N4955);
xor XOR2 (N4961, N4959, N4815);
or OR2 (N4962, N4961, N466);
or OR3 (N4963, N4950, N3733, N4639);
or OR2 (N4964, N4960, N2320);
and AND3 (N4965, N4962, N4713, N1828);
nand NAND2 (N4966, N4957, N1797);
or OR2 (N4967, N4964, N2682);
nand NAND3 (N4968, N4956, N4379, N4485);
or OR2 (N4969, N4963, N4922);
and AND2 (N4970, N4952, N3850);
nand NAND3 (N4971, N4965, N3108, N4153);
buf BUF1 (N4972, N4970);
or OR4 (N4973, N4937, N2916, N834, N4494);
nand NAND2 (N4974, N4966, N3543);
nand NAND2 (N4975, N4954, N2197);
buf BUF1 (N4976, N4969);
or OR3 (N4977, N4973, N1642, N4267);
xor XOR2 (N4978, N4974, N1921);
nor NOR4 (N4979, N4971, N3408, N561, N4548);
not NOT1 (N4980, N4938);
nor NOR2 (N4981, N4980, N4238);
buf BUF1 (N4982, N4977);
not NOT1 (N4983, N4979);
or OR3 (N4984, N4972, N2774, N634);
buf BUF1 (N4985, N4968);
and AND2 (N4986, N4967, N4300);
nand NAND2 (N4987, N4985, N398);
nor NOR4 (N4988, N4935, N142, N522, N1537);
nand NAND2 (N4989, N4975, N3579);
nor NOR3 (N4990, N4981, N4966, N1608);
or OR2 (N4991, N4990, N2620);
nor NOR3 (N4992, N4989, N2803, N3196);
not NOT1 (N4993, N4982);
nand NAND2 (N4994, N4991, N2953);
nand NAND3 (N4995, N4986, N3758, N4952);
nand NAND2 (N4996, N4983, N4215);
xor XOR2 (N4997, N4995, N544);
or OR2 (N4998, N4988, N4372);
xor XOR2 (N4999, N4993, N3733);
not NOT1 (N5000, N4997);
nand NAND4 (N5001, N4976, N3549, N459, N3324);
nand NAND2 (N5002, N4978, N4925);
or OR2 (N5003, N4992, N711);
not NOT1 (N5004, N4984);
and AND2 (N5005, N4999, N2272);
and AND3 (N5006, N5001, N3870, N628);
or OR2 (N5007, N4998, N2048);
nand NAND4 (N5008, N5005, N2637, N4817, N2979);
and AND3 (N5009, N5002, N4880, N376);
buf BUF1 (N5010, N5006);
or OR2 (N5011, N4996, N3291);
or OR4 (N5012, N4987, N1988, N410, N1652);
and AND2 (N5013, N5008, N3975);
buf BUF1 (N5014, N4994);
or OR2 (N5015, N5010, N2336);
not NOT1 (N5016, N5003);
nor NOR3 (N5017, N5009, N1645, N229);
buf BUF1 (N5018, N5007);
nand NAND3 (N5019, N5012, N164, N4591);
not NOT1 (N5020, N5015);
or OR2 (N5021, N5004, N793);
xor XOR2 (N5022, N5019, N1824);
nand NAND2 (N5023, N5013, N1178);
xor XOR2 (N5024, N5022, N4702);
xor XOR2 (N5025, N5020, N2434);
xor XOR2 (N5026, N5021, N4823);
or OR3 (N5027, N5017, N479, N464);
xor XOR2 (N5028, N5011, N914);
nor NOR3 (N5029, N5026, N397, N2286);
nor NOR4 (N5030, N5025, N2283, N1064, N4785);
and AND4 (N5031, N5029, N1647, N1312, N3596);
nand NAND2 (N5032, N5000, N3100);
xor XOR2 (N5033, N5027, N3470);
or OR4 (N5034, N5032, N1897, N3043, N4489);
and AND3 (N5035, N5033, N3542, N3183);
buf BUF1 (N5036, N5034);
nor NOR4 (N5037, N5016, N2042, N3556, N3617);
buf BUF1 (N5038, N5035);
buf BUF1 (N5039, N5028);
nand NAND2 (N5040, N5030, N4499);
xor XOR2 (N5041, N5036, N3841);
and AND3 (N5042, N5031, N1674, N661);
nand NAND2 (N5043, N5014, N4972);
buf BUF1 (N5044, N5018);
xor XOR2 (N5045, N5024, N169);
xor XOR2 (N5046, N5042, N3053);
or OR3 (N5047, N5043, N4630, N4342);
xor XOR2 (N5048, N5040, N2132);
and AND3 (N5049, N5041, N1403, N2360);
or OR3 (N5050, N5047, N3153, N3408);
xor XOR2 (N5051, N5049, N4981);
nand NAND4 (N5052, N5050, N1824, N3653, N506);
xor XOR2 (N5053, N5051, N4138);
not NOT1 (N5054, N5038);
buf BUF1 (N5055, N5023);
not NOT1 (N5056, N5054);
nor NOR3 (N5057, N5056, N3277, N4520);
nand NAND2 (N5058, N5057, N4569);
xor XOR2 (N5059, N5048, N4348);
nor NOR4 (N5060, N5055, N1783, N717, N1707);
nand NAND2 (N5061, N5053, N3413);
nor NOR2 (N5062, N5037, N4051);
xor XOR2 (N5063, N5046, N2133);
nor NOR2 (N5064, N5044, N2647);
not NOT1 (N5065, N5060);
nor NOR3 (N5066, N5052, N58, N2260);
and AND4 (N5067, N5063, N2355, N670, N3968);
nor NOR3 (N5068, N5065, N3382, N3382);
nand NAND4 (N5069, N5062, N165, N3910, N4703);
not NOT1 (N5070, N5039);
or OR3 (N5071, N5069, N4946, N1638);
xor XOR2 (N5072, N5068, N4058);
not NOT1 (N5073, N5061);
or OR4 (N5074, N5064, N1735, N1190, N3438);
and AND2 (N5075, N5066, N908);
nor NOR3 (N5076, N5075, N610, N4374);
buf BUF1 (N5077, N5059);
and AND2 (N5078, N5067, N2495);
buf BUF1 (N5079, N5072);
and AND4 (N5080, N5074, N894, N3250, N1224);
and AND2 (N5081, N5079, N2496);
not NOT1 (N5082, N5078);
buf BUF1 (N5083, N5077);
xor XOR2 (N5084, N5070, N1518);
not NOT1 (N5085, N5045);
xor XOR2 (N5086, N5080, N2684);
buf BUF1 (N5087, N5071);
nand NAND3 (N5088, N5084, N110, N413);
and AND3 (N5089, N5081, N1709, N5062);
nand NAND4 (N5090, N5082, N1859, N2233, N1443);
and AND2 (N5091, N5085, N2354);
nand NAND3 (N5092, N5090, N1251, N1634);
xor XOR2 (N5093, N5087, N563);
nand NAND3 (N5094, N5088, N500, N3915);
xor XOR2 (N5095, N5094, N4010);
not NOT1 (N5096, N5083);
not NOT1 (N5097, N5058);
or OR4 (N5098, N5093, N3458, N4871, N1123);
nand NAND2 (N5099, N5091, N4002);
not NOT1 (N5100, N5095);
nor NOR2 (N5101, N5099, N1125);
or OR4 (N5102, N5092, N67, N1868, N2768);
or OR3 (N5103, N5086, N2472, N1171);
nor NOR3 (N5104, N5102, N4170, N1666);
nand NAND4 (N5105, N5076, N3727, N2504, N4618);
buf BUF1 (N5106, N5104);
nand NAND2 (N5107, N5106, N3433);
buf BUF1 (N5108, N5073);
nand NAND2 (N5109, N5096, N2759);
buf BUF1 (N5110, N5089);
not NOT1 (N5111, N5108);
xor XOR2 (N5112, N5100, N2512);
not NOT1 (N5113, N5103);
buf BUF1 (N5114, N5111);
xor XOR2 (N5115, N5114, N110);
or OR4 (N5116, N5109, N1473, N569, N2351);
buf BUF1 (N5117, N5115);
buf BUF1 (N5118, N5105);
nand NAND3 (N5119, N5113, N3216, N1980);
nor NOR4 (N5120, N5116, N595, N2421, N1616);
nand NAND4 (N5121, N5118, N1872, N4249, N4860);
and AND4 (N5122, N5098, N4140, N2933, N4778);
or OR2 (N5123, N5122, N1990);
xor XOR2 (N5124, N5120, N2107);
not NOT1 (N5125, N5101);
xor XOR2 (N5126, N5097, N1719);
nand NAND3 (N5127, N5123, N955, N1989);
and AND2 (N5128, N5125, N3534);
not NOT1 (N5129, N5112);
or OR2 (N5130, N5127, N940);
nand NAND4 (N5131, N5130, N4954, N460, N2820);
xor XOR2 (N5132, N5128, N2044);
xor XOR2 (N5133, N5119, N4415);
nand NAND3 (N5134, N5133, N2469, N1755);
or OR2 (N5135, N5121, N440);
buf BUF1 (N5136, N5126);
xor XOR2 (N5137, N5124, N3261);
nand NAND3 (N5138, N5134, N1228, N1711);
nand NAND2 (N5139, N5135, N4843);
nand NAND3 (N5140, N5132, N3303, N408);
nor NOR3 (N5141, N5117, N5005, N2057);
xor XOR2 (N5142, N5107, N2809);
and AND2 (N5143, N5140, N691);
buf BUF1 (N5144, N5143);
xor XOR2 (N5145, N5144, N3273);
nand NAND4 (N5146, N5145, N4978, N951, N2735);
or OR3 (N5147, N5139, N2680, N805);
or OR2 (N5148, N5147, N1992);
nor NOR4 (N5149, N5131, N2931, N873, N1658);
xor XOR2 (N5150, N5142, N532);
buf BUF1 (N5151, N5146);
and AND4 (N5152, N5151, N1659, N1626, N4310);
nand NAND2 (N5153, N5148, N4948);
buf BUF1 (N5154, N5152);
and AND3 (N5155, N5137, N3155, N3566);
nor NOR4 (N5156, N5155, N3061, N65, N902);
buf BUF1 (N5157, N5129);
xor XOR2 (N5158, N5156, N2146);
nand NAND3 (N5159, N5158, N1232, N1947);
and AND4 (N5160, N5157, N1959, N4921, N1346);
or OR2 (N5161, N5141, N1758);
nor NOR2 (N5162, N5150, N1993);
xor XOR2 (N5163, N5159, N3605);
and AND4 (N5164, N5153, N191, N1468, N4070);
xor XOR2 (N5165, N5163, N1926);
nor NOR2 (N5166, N5110, N2114);
nand NAND4 (N5167, N5164, N2347, N4336, N4402);
nand NAND3 (N5168, N5160, N1051, N3512);
xor XOR2 (N5169, N5138, N3338);
nand NAND2 (N5170, N5161, N1417);
not NOT1 (N5171, N5149);
nor NOR4 (N5172, N5136, N3129, N90, N1649);
buf BUF1 (N5173, N5166);
nand NAND2 (N5174, N5170, N919);
buf BUF1 (N5175, N5174);
xor XOR2 (N5176, N5175, N675);
nor NOR4 (N5177, N5176, N4346, N752, N2093);
buf BUF1 (N5178, N5165);
buf BUF1 (N5179, N5154);
buf BUF1 (N5180, N5169);
and AND3 (N5181, N5167, N1906, N3472);
nor NOR3 (N5182, N5179, N3367, N3506);
and AND4 (N5183, N5181, N1871, N487, N2289);
xor XOR2 (N5184, N5162, N3015);
xor XOR2 (N5185, N5182, N72);
or OR2 (N5186, N5171, N3089);
or OR2 (N5187, N5184, N3385);
and AND3 (N5188, N5183, N4490, N752);
not NOT1 (N5189, N5180);
nand NAND2 (N5190, N5186, N965);
nor NOR3 (N5191, N5178, N2127, N5083);
buf BUF1 (N5192, N5187);
nor NOR3 (N5193, N5185, N4615, N4640);
and AND3 (N5194, N5177, N1428, N891);
buf BUF1 (N5195, N5168);
not NOT1 (N5196, N5173);
not NOT1 (N5197, N5188);
buf BUF1 (N5198, N5190);
nor NOR2 (N5199, N5198, N3677);
buf BUF1 (N5200, N5194);
not NOT1 (N5201, N5192);
nand NAND4 (N5202, N5191, N53, N2713, N5031);
xor XOR2 (N5203, N5199, N3416);
or OR2 (N5204, N5193, N690);
or OR4 (N5205, N5200, N3517, N967, N128);
nor NOR4 (N5206, N5204, N879, N2574, N3150);
nand NAND2 (N5207, N5172, N909);
buf BUF1 (N5208, N5196);
buf BUF1 (N5209, N5203);
not NOT1 (N5210, N5207);
or OR4 (N5211, N5205, N4813, N2698, N1539);
or OR2 (N5212, N5209, N4649);
nand NAND3 (N5213, N5189, N3243, N2699);
not NOT1 (N5214, N5201);
xor XOR2 (N5215, N5213, N5093);
and AND3 (N5216, N5202, N2293, N4735);
not NOT1 (N5217, N5206);
xor XOR2 (N5218, N5208, N3291);
xor XOR2 (N5219, N5210, N1148);
buf BUF1 (N5220, N5217);
or OR4 (N5221, N5195, N4642, N4472, N742);
nand NAND3 (N5222, N5216, N3902, N5125);
xor XOR2 (N5223, N5222, N4839);
or OR2 (N5224, N5211, N3155);
nand NAND3 (N5225, N5223, N1505, N4726);
buf BUF1 (N5226, N5219);
buf BUF1 (N5227, N5212);
or OR3 (N5228, N5197, N4905, N4119);
and AND2 (N5229, N5226, N663);
not NOT1 (N5230, N5221);
nor NOR2 (N5231, N5230, N4975);
nand NAND3 (N5232, N5224, N45, N4943);
buf BUF1 (N5233, N5229);
nor NOR3 (N5234, N5215, N2361, N4714);
nand NAND3 (N5235, N5214, N2497, N3384);
nand NAND3 (N5236, N5232, N3300, N1521);
and AND3 (N5237, N5236, N4457, N3353);
not NOT1 (N5238, N5218);
nand NAND4 (N5239, N5234, N2991, N2723, N4269);
not NOT1 (N5240, N5235);
nor NOR3 (N5241, N5225, N1499, N4641);
buf BUF1 (N5242, N5239);
or OR2 (N5243, N5227, N5027);
nand NAND2 (N5244, N5231, N2123);
nand NAND3 (N5245, N5228, N142, N2467);
nor NOR3 (N5246, N5238, N5120, N2401);
nand NAND4 (N5247, N5244, N3727, N1845, N4173);
and AND4 (N5248, N5241, N588, N300, N2758);
xor XOR2 (N5249, N5248, N3478);
nand NAND3 (N5250, N5243, N3168, N4237);
buf BUF1 (N5251, N5220);
buf BUF1 (N5252, N5246);
xor XOR2 (N5253, N5252, N1938);
not NOT1 (N5254, N5240);
xor XOR2 (N5255, N5242, N24);
xor XOR2 (N5256, N5253, N1333);
xor XOR2 (N5257, N5233, N2822);
buf BUF1 (N5258, N5251);
or OR2 (N5259, N5249, N1579);
not NOT1 (N5260, N5247);
xor XOR2 (N5261, N5245, N3903);
buf BUF1 (N5262, N5257);
nor NOR4 (N5263, N5256, N980, N3477, N4552);
nor NOR2 (N5264, N5259, N2950);
xor XOR2 (N5265, N5264, N432);
and AND2 (N5266, N5261, N3199);
buf BUF1 (N5267, N5262);
not NOT1 (N5268, N5250);
nand NAND3 (N5269, N5255, N2370, N2951);
and AND3 (N5270, N5266, N4224, N3543);
not NOT1 (N5271, N5269);
and AND2 (N5272, N5270, N1668);
nand NAND2 (N5273, N5267, N4623);
nor NOR4 (N5274, N5272, N3657, N5087, N41);
nand NAND2 (N5275, N5263, N1285);
nor NOR4 (N5276, N5254, N3215, N3425, N2443);
nand NAND3 (N5277, N5268, N3301, N3165);
buf BUF1 (N5278, N5275);
not NOT1 (N5279, N5276);
buf BUF1 (N5280, N5265);
not NOT1 (N5281, N5237);
buf BUF1 (N5282, N5278);
xor XOR2 (N5283, N5260, N1089);
nand NAND2 (N5284, N5281, N1137);
nand NAND4 (N5285, N5282, N3884, N2552, N2650);
buf BUF1 (N5286, N5271);
nand NAND3 (N5287, N5277, N1469, N3143);
nand NAND3 (N5288, N5283, N1151, N1749);
or OR4 (N5289, N5285, N4558, N3052, N2694);
xor XOR2 (N5290, N5279, N3841);
buf BUF1 (N5291, N5274);
xor XOR2 (N5292, N5287, N4834);
nand NAND4 (N5293, N5273, N717, N4366, N2213);
nand NAND4 (N5294, N5290, N2202, N3253, N1268);
xor XOR2 (N5295, N5292, N1315);
and AND4 (N5296, N5280, N478, N535, N3118);
nand NAND4 (N5297, N5295, N5183, N2653, N1508);
and AND4 (N5298, N5286, N4433, N2894, N4284);
nor NOR3 (N5299, N5297, N989, N4943);
buf BUF1 (N5300, N5284);
xor XOR2 (N5301, N5288, N1820);
nor NOR3 (N5302, N5293, N3630, N257);
buf BUF1 (N5303, N5294);
xor XOR2 (N5304, N5301, N1007);
buf BUF1 (N5305, N5300);
and AND3 (N5306, N5258, N1157, N2091);
nor NOR4 (N5307, N5306, N1059, N2419, N4726);
not NOT1 (N5308, N5303);
or OR2 (N5309, N5289, N3255);
nor NOR2 (N5310, N5291, N1324);
xor XOR2 (N5311, N5304, N1837);
buf BUF1 (N5312, N5296);
and AND4 (N5313, N5298, N2534, N2175, N5147);
nor NOR4 (N5314, N5312, N3013, N575, N2176);
and AND4 (N5315, N5307, N1665, N3894, N166);
or OR2 (N5316, N5305, N694);
nor NOR3 (N5317, N5309, N157, N1598);
nand NAND2 (N5318, N5317, N1019);
nor NOR2 (N5319, N5310, N1972);
buf BUF1 (N5320, N5302);
and AND3 (N5321, N5315, N3361, N341);
buf BUF1 (N5322, N5321);
nor NOR2 (N5323, N5318, N3659);
and AND3 (N5324, N5311, N487, N2702);
not NOT1 (N5325, N5299);
and AND3 (N5326, N5323, N3104, N597);
buf BUF1 (N5327, N5326);
not NOT1 (N5328, N5324);
nor NOR2 (N5329, N5314, N2229);
and AND2 (N5330, N5316, N305);
xor XOR2 (N5331, N5327, N2367);
nor NOR4 (N5332, N5325, N3602, N3120, N2025);
not NOT1 (N5333, N5328);
nor NOR2 (N5334, N5322, N5044);
nor NOR4 (N5335, N5331, N2253, N3144, N2521);
buf BUF1 (N5336, N5334);
or OR3 (N5337, N5320, N2654, N4866);
nand NAND2 (N5338, N5308, N1856);
xor XOR2 (N5339, N5333, N4418);
nand NAND4 (N5340, N5319, N432, N2303, N3894);
buf BUF1 (N5341, N5340);
and AND2 (N5342, N5330, N1976);
or OR2 (N5343, N5335, N2319);
or OR3 (N5344, N5329, N1613, N944);
not NOT1 (N5345, N5339);
not NOT1 (N5346, N5337);
nor NOR2 (N5347, N5336, N2295);
nor NOR2 (N5348, N5342, N2168);
or OR4 (N5349, N5341, N3798, N1542, N2610);
xor XOR2 (N5350, N5343, N5177);
or OR2 (N5351, N5347, N453);
xor XOR2 (N5352, N5313, N2331);
not NOT1 (N5353, N5349);
not NOT1 (N5354, N5345);
nand NAND2 (N5355, N5352, N3374);
and AND4 (N5356, N5350, N1707, N1687, N493);
nand NAND4 (N5357, N5332, N2618, N1364, N4939);
not NOT1 (N5358, N5348);
or OR4 (N5359, N5354, N4535, N222, N2073);
buf BUF1 (N5360, N5359);
not NOT1 (N5361, N5353);
buf BUF1 (N5362, N5351);
not NOT1 (N5363, N5358);
buf BUF1 (N5364, N5362);
not NOT1 (N5365, N5346);
nor NOR2 (N5366, N5363, N3427);
buf BUF1 (N5367, N5360);
xor XOR2 (N5368, N5361, N283);
nor NOR2 (N5369, N5338, N1602);
and AND4 (N5370, N5368, N4931, N3346, N412);
nand NAND2 (N5371, N5366, N4681);
nor NOR2 (N5372, N5369, N1115);
nor NOR3 (N5373, N5356, N300, N4796);
not NOT1 (N5374, N5370);
buf BUF1 (N5375, N5344);
buf BUF1 (N5376, N5371);
buf BUF1 (N5377, N5357);
nand NAND4 (N5378, N5367, N3780, N2788, N318);
buf BUF1 (N5379, N5378);
not NOT1 (N5380, N5375);
and AND4 (N5381, N5373, N4269, N820, N4583);
or OR4 (N5382, N5364, N2315, N3338, N3855);
not NOT1 (N5383, N5355);
not NOT1 (N5384, N5380);
xor XOR2 (N5385, N5384, N3391);
not NOT1 (N5386, N5365);
nand NAND2 (N5387, N5382, N194);
nor NOR3 (N5388, N5374, N380, N1012);
or OR3 (N5389, N5379, N3805, N4561);
nor NOR4 (N5390, N5388, N2708, N3381, N1725);
xor XOR2 (N5391, N5385, N202);
not NOT1 (N5392, N5383);
nand NAND4 (N5393, N5389, N5246, N5055, N5367);
xor XOR2 (N5394, N5391, N391);
buf BUF1 (N5395, N5387);
nand NAND3 (N5396, N5377, N3431, N2759);
nor NOR3 (N5397, N5386, N3911, N1945);
nand NAND3 (N5398, N5395, N2677, N1990);
not NOT1 (N5399, N5397);
buf BUF1 (N5400, N5396);
nand NAND2 (N5401, N5376, N2208);
nor NOR2 (N5402, N5390, N4004);
xor XOR2 (N5403, N5399, N1404);
not NOT1 (N5404, N5381);
nor NOR4 (N5405, N5400, N2100, N4471, N511);
nor NOR4 (N5406, N5402, N745, N1111, N4419);
or OR3 (N5407, N5393, N4575, N4536);
buf BUF1 (N5408, N5392);
nor NOR2 (N5409, N5408, N11);
not NOT1 (N5410, N5405);
or OR4 (N5411, N5401, N3091, N97, N1916);
not NOT1 (N5412, N5394);
not NOT1 (N5413, N5407);
nand NAND3 (N5414, N5398, N284, N1173);
nor NOR2 (N5415, N5404, N69);
buf BUF1 (N5416, N5412);
and AND2 (N5417, N5372, N1564);
nor NOR2 (N5418, N5411, N3220);
xor XOR2 (N5419, N5416, N1341);
nand NAND4 (N5420, N5417, N207, N663, N916);
not NOT1 (N5421, N5419);
nand NAND2 (N5422, N5414, N3459);
not NOT1 (N5423, N5406);
or OR3 (N5424, N5413, N99, N1565);
nor NOR4 (N5425, N5423, N3462, N4846, N5078);
xor XOR2 (N5426, N5410, N2200);
not NOT1 (N5427, N5421);
nand NAND3 (N5428, N5427, N3614, N2445);
and AND4 (N5429, N5409, N2964, N1765, N1561);
nand NAND3 (N5430, N5429, N5263, N2917);
not NOT1 (N5431, N5403);
nor NOR3 (N5432, N5415, N3584, N2214);
or OR3 (N5433, N5428, N2885, N117);
nor NOR4 (N5434, N5431, N2179, N2364, N4410);
not NOT1 (N5435, N5433);
and AND2 (N5436, N5430, N3793);
and AND2 (N5437, N5420, N2595);
and AND2 (N5438, N5434, N2319);
xor XOR2 (N5439, N5438, N2231);
nor NOR2 (N5440, N5436, N2645);
xor XOR2 (N5441, N5439, N2452);
buf BUF1 (N5442, N5422);
and AND2 (N5443, N5432, N2063);
not NOT1 (N5444, N5443);
and AND2 (N5445, N5424, N4590);
nor NOR4 (N5446, N5426, N1474, N5362, N1339);
not NOT1 (N5447, N5446);
xor XOR2 (N5448, N5437, N5056);
and AND4 (N5449, N5447, N1218, N3394, N3700);
or OR4 (N5450, N5445, N4954, N3699, N4040);
nand NAND4 (N5451, N5425, N4890, N1801, N2849);
or OR3 (N5452, N5451, N3000, N2508);
nand NAND4 (N5453, N5435, N5135, N2365, N3596);
nand NAND4 (N5454, N5418, N4919, N5130, N1833);
or OR2 (N5455, N5449, N2748);
not NOT1 (N5456, N5452);
nand NAND2 (N5457, N5448, N2949);
and AND4 (N5458, N5455, N2316, N3847, N2574);
buf BUF1 (N5459, N5441);
nand NAND4 (N5460, N5457, N1236, N2082, N4283);
buf BUF1 (N5461, N5459);
nor NOR2 (N5462, N5444, N3502);
xor XOR2 (N5463, N5454, N1179);
buf BUF1 (N5464, N5458);
or OR4 (N5465, N5453, N2589, N2667, N1782);
xor XOR2 (N5466, N5465, N1404);
nand NAND3 (N5467, N5460, N5466, N2710);
nand NAND3 (N5468, N1859, N2226, N3409);
buf BUF1 (N5469, N5464);
and AND4 (N5470, N5468, N3103, N3524, N213);
or OR4 (N5471, N5467, N502, N1906, N3863);
nand NAND2 (N5472, N5462, N3784);
not NOT1 (N5473, N5471);
nor NOR4 (N5474, N5456, N2258, N3191, N4310);
or OR2 (N5475, N5442, N4813);
buf BUF1 (N5476, N5475);
not NOT1 (N5477, N5474);
xor XOR2 (N5478, N5440, N1824);
xor XOR2 (N5479, N5478, N1133);
xor XOR2 (N5480, N5472, N3634);
nand NAND2 (N5481, N5477, N217);
buf BUF1 (N5482, N5461);
and AND3 (N5483, N5450, N3905, N3457);
not NOT1 (N5484, N5479);
nor NOR4 (N5485, N5469, N3751, N5371, N1231);
nor NOR4 (N5486, N5463, N4544, N2501, N5264);
not NOT1 (N5487, N5482);
or OR3 (N5488, N5470, N1851, N1327);
nor NOR4 (N5489, N5484, N5233, N2063, N1327);
buf BUF1 (N5490, N5476);
xor XOR2 (N5491, N5481, N3395);
nand NAND2 (N5492, N5489, N1316);
or OR4 (N5493, N5490, N974, N575, N1183);
or OR4 (N5494, N5493, N2015, N4698, N1704);
nand NAND2 (N5495, N5494, N3631);
xor XOR2 (N5496, N5486, N2414);
nor NOR3 (N5497, N5488, N3384, N4470);
nor NOR4 (N5498, N5473, N235, N738, N725);
xor XOR2 (N5499, N5483, N2980);
buf BUF1 (N5500, N5496);
and AND4 (N5501, N5495, N2956, N411, N4424);
or OR2 (N5502, N5499, N3378);
xor XOR2 (N5503, N5502, N934);
nor NOR3 (N5504, N5492, N798, N819);
and AND2 (N5505, N5491, N3307);
xor XOR2 (N5506, N5480, N3124);
xor XOR2 (N5507, N5505, N902);
or OR2 (N5508, N5485, N1055);
not NOT1 (N5509, N5501);
nor NOR2 (N5510, N5506, N1348);
nand NAND4 (N5511, N5500, N2659, N5380, N3350);
buf BUF1 (N5512, N5504);
not NOT1 (N5513, N5503);
buf BUF1 (N5514, N5498);
and AND3 (N5515, N5508, N2325, N2297);
not NOT1 (N5516, N5512);
or OR2 (N5517, N5511, N761);
and AND2 (N5518, N5497, N1133);
buf BUF1 (N5519, N5513);
or OR3 (N5520, N5509, N2721, N979);
xor XOR2 (N5521, N5487, N4384);
not NOT1 (N5522, N5516);
or OR2 (N5523, N5518, N953);
xor XOR2 (N5524, N5507, N722);
nand NAND4 (N5525, N5510, N2214, N2561, N1532);
not NOT1 (N5526, N5524);
xor XOR2 (N5527, N5514, N4521);
not NOT1 (N5528, N5526);
xor XOR2 (N5529, N5527, N4893);
nand NAND4 (N5530, N5515, N4595, N4526, N395);
and AND4 (N5531, N5528, N2585, N917, N1979);
xor XOR2 (N5532, N5520, N399);
not NOT1 (N5533, N5521);
or OR2 (N5534, N5530, N262);
xor XOR2 (N5535, N5517, N288);
xor XOR2 (N5536, N5533, N2641);
xor XOR2 (N5537, N5531, N46);
nand NAND4 (N5538, N5532, N1423, N412, N4418);
nand NAND4 (N5539, N5523, N514, N1707, N1599);
or OR2 (N5540, N5536, N1299);
xor XOR2 (N5541, N5525, N3366);
nand NAND3 (N5542, N5529, N917, N4815);
not NOT1 (N5543, N5535);
nor NOR3 (N5544, N5519, N1355, N3307);
or OR3 (N5545, N5540, N3729, N3132);
buf BUF1 (N5546, N5543);
nand NAND4 (N5547, N5534, N875, N2225, N1535);
or OR4 (N5548, N5537, N4222, N620, N4386);
buf BUF1 (N5549, N5539);
not NOT1 (N5550, N5545);
buf BUF1 (N5551, N5522);
nor NOR3 (N5552, N5551, N2528, N1913);
nor NOR3 (N5553, N5549, N656, N5090);
xor XOR2 (N5554, N5547, N2323);
nand NAND4 (N5555, N5546, N4841, N2453, N3559);
not NOT1 (N5556, N5544);
and AND2 (N5557, N5542, N2099);
xor XOR2 (N5558, N5556, N3845);
xor XOR2 (N5559, N5557, N2892);
and AND4 (N5560, N5553, N3237, N2131, N1908);
or OR4 (N5561, N5555, N1096, N1119, N2600);
xor XOR2 (N5562, N5560, N3848);
and AND2 (N5563, N5558, N3882);
buf BUF1 (N5564, N5552);
or OR3 (N5565, N5541, N4402, N3574);
xor XOR2 (N5566, N5554, N5036);
nor NOR4 (N5567, N5564, N1158, N5244, N353);
nor NOR4 (N5568, N5548, N4402, N865, N3355);
nand NAND3 (N5569, N5550, N3358, N5304);
xor XOR2 (N5570, N5563, N2843);
and AND3 (N5571, N5570, N4863, N546);
nand NAND4 (N5572, N5565, N949, N3205, N4793);
buf BUF1 (N5573, N5568);
buf BUF1 (N5574, N5572);
and AND2 (N5575, N5573, N4909);
buf BUF1 (N5576, N5562);
xor XOR2 (N5577, N5574, N3644);
not NOT1 (N5578, N5575);
xor XOR2 (N5579, N5559, N2976);
nor NOR2 (N5580, N5569, N3533);
buf BUF1 (N5581, N5567);
not NOT1 (N5582, N5571);
or OR4 (N5583, N5576, N2024, N1007, N2604);
and AND2 (N5584, N5579, N1208);
nor NOR3 (N5585, N5577, N5496, N876);
not NOT1 (N5586, N5581);
not NOT1 (N5587, N5578);
xor XOR2 (N5588, N5566, N3787);
buf BUF1 (N5589, N5588);
buf BUF1 (N5590, N5584);
or OR4 (N5591, N5589, N153, N832, N1836);
xor XOR2 (N5592, N5580, N576);
buf BUF1 (N5593, N5582);
nor NOR4 (N5594, N5587, N5230, N681, N70);
xor XOR2 (N5595, N5591, N7);
nor NOR4 (N5596, N5583, N2252, N287, N2176);
and AND3 (N5597, N5593, N2754, N4850);
buf BUF1 (N5598, N5586);
nand NAND4 (N5599, N5561, N3078, N4493, N2164);
or OR2 (N5600, N5538, N1381);
or OR2 (N5601, N5596, N4926);
nor NOR2 (N5602, N5595, N2266);
buf BUF1 (N5603, N5600);
and AND4 (N5604, N5592, N724, N5518, N5120);
xor XOR2 (N5605, N5594, N5392);
nand NAND2 (N5606, N5585, N4562);
nor NOR2 (N5607, N5602, N167);
nor NOR3 (N5608, N5606, N3230, N1414);
or OR2 (N5609, N5597, N1039);
or OR4 (N5610, N5590, N1614, N737, N5132);
and AND4 (N5611, N5610, N2515, N5093, N1012);
buf BUF1 (N5612, N5599);
and AND2 (N5613, N5609, N3096);
xor XOR2 (N5614, N5607, N481);
buf BUF1 (N5615, N5604);
nor NOR4 (N5616, N5598, N2133, N608, N800);
buf BUF1 (N5617, N5613);
and AND4 (N5618, N5605, N3911, N3486, N4013);
not NOT1 (N5619, N5608);
nand NAND2 (N5620, N5603, N4870);
nand NAND3 (N5621, N5611, N2515, N3474);
buf BUF1 (N5622, N5617);
and AND4 (N5623, N5612, N935, N4396, N999);
or OR4 (N5624, N5601, N2552, N4697, N5045);
nand NAND3 (N5625, N5622, N2081, N5153);
and AND3 (N5626, N5625, N1941, N2326);
xor XOR2 (N5627, N5618, N4997);
and AND2 (N5628, N5627, N2919);
or OR3 (N5629, N5619, N5011, N4529);
and AND4 (N5630, N5615, N3389, N2229, N4030);
nand NAND2 (N5631, N5621, N2000);
buf BUF1 (N5632, N5628);
or OR2 (N5633, N5629, N2548);
or OR2 (N5634, N5630, N1188);
or OR3 (N5635, N5614, N4592, N1024);
nand NAND4 (N5636, N5631, N426, N4944, N3731);
buf BUF1 (N5637, N5624);
not NOT1 (N5638, N5633);
or OR4 (N5639, N5634, N4706, N5544, N3476);
buf BUF1 (N5640, N5626);
or OR2 (N5641, N5616, N3947);
nand NAND3 (N5642, N5639, N2401, N3875);
and AND4 (N5643, N5636, N1748, N5220, N2808);
or OR3 (N5644, N5632, N4763, N4360);
not NOT1 (N5645, N5623);
not NOT1 (N5646, N5640);
or OR4 (N5647, N5642, N1916, N4378, N946);
not NOT1 (N5648, N5644);
nor NOR4 (N5649, N5638, N2370, N598, N101);
xor XOR2 (N5650, N5620, N5536);
buf BUF1 (N5651, N5635);
buf BUF1 (N5652, N5646);
nor NOR4 (N5653, N5649, N2901, N994, N2029);
buf BUF1 (N5654, N5651);
and AND3 (N5655, N5654, N4364, N703);
nand NAND3 (N5656, N5647, N3235, N1057);
nor NOR4 (N5657, N5637, N4340, N5423, N443);
not NOT1 (N5658, N5641);
buf BUF1 (N5659, N5658);
buf BUF1 (N5660, N5652);
not NOT1 (N5661, N5657);
nand NAND3 (N5662, N5645, N1604, N253);
xor XOR2 (N5663, N5653, N4960);
nor NOR4 (N5664, N5656, N1315, N1169, N5628);
buf BUF1 (N5665, N5664);
or OR4 (N5666, N5665, N5622, N154, N2246);
and AND2 (N5667, N5655, N2934);
nor NOR2 (N5668, N5666, N4074);
buf BUF1 (N5669, N5660);
and AND2 (N5670, N5662, N803);
or OR4 (N5671, N5650, N3698, N1873, N3892);
or OR4 (N5672, N5668, N3632, N1815, N42);
nor NOR2 (N5673, N5667, N683);
or OR2 (N5674, N5661, N4169);
buf BUF1 (N5675, N5643);
xor XOR2 (N5676, N5659, N5061);
or OR4 (N5677, N5671, N317, N1354, N2499);
buf BUF1 (N5678, N5673);
and AND3 (N5679, N5678, N4222, N3599);
not NOT1 (N5680, N5648);
or OR2 (N5681, N5672, N3444);
buf BUF1 (N5682, N5675);
and AND3 (N5683, N5670, N319, N1608);
nand NAND2 (N5684, N5676, N5424);
not NOT1 (N5685, N5684);
xor XOR2 (N5686, N5663, N1283);
xor XOR2 (N5687, N5681, N410);
or OR4 (N5688, N5686, N3398, N149, N3408);
and AND3 (N5689, N5677, N1486, N3240);
xor XOR2 (N5690, N5685, N4191);
or OR4 (N5691, N5680, N422, N118, N1957);
nand NAND3 (N5692, N5679, N343, N102);
and AND4 (N5693, N5688, N481, N2689, N2001);
nand NAND4 (N5694, N5674, N2595, N3675, N68);
buf BUF1 (N5695, N5691);
not NOT1 (N5696, N5694);
xor XOR2 (N5697, N5682, N1607);
xor XOR2 (N5698, N5687, N3015);
xor XOR2 (N5699, N5696, N5123);
nand NAND4 (N5700, N5683, N2744, N3890, N541);
buf BUF1 (N5701, N5698);
or OR2 (N5702, N5699, N3478);
not NOT1 (N5703, N5700);
not NOT1 (N5704, N5703);
nand NAND4 (N5705, N5689, N5504, N3806, N4796);
buf BUF1 (N5706, N5690);
nand NAND2 (N5707, N5706, N1956);
xor XOR2 (N5708, N5695, N29);
xor XOR2 (N5709, N5669, N3942);
or OR3 (N5710, N5702, N3032, N4254);
or OR4 (N5711, N5705, N3768, N26, N1976);
not NOT1 (N5712, N5709);
or OR4 (N5713, N5693, N2775, N3369, N2014);
buf BUF1 (N5714, N5713);
nor NOR2 (N5715, N5708, N2818);
xor XOR2 (N5716, N5701, N659);
not NOT1 (N5717, N5704);
and AND4 (N5718, N5717, N2136, N951, N4679);
not NOT1 (N5719, N5712);
nand NAND4 (N5720, N5719, N4443, N1367, N226);
nand NAND4 (N5721, N5715, N4621, N2317, N1344);
buf BUF1 (N5722, N5720);
nand NAND4 (N5723, N5707, N4902, N550, N1159);
or OR2 (N5724, N5711, N4769);
nor NOR2 (N5725, N5692, N2801);
and AND4 (N5726, N5714, N110, N3540, N65);
and AND3 (N5727, N5718, N1910, N4564);
not NOT1 (N5728, N5727);
nor NOR3 (N5729, N5710, N293, N453);
xor XOR2 (N5730, N5722, N1680);
nor NOR2 (N5731, N5721, N1665);
and AND3 (N5732, N5730, N1252, N4606);
not NOT1 (N5733, N5728);
xor XOR2 (N5734, N5723, N5616);
nor NOR3 (N5735, N5734, N5098, N4953);
nand NAND2 (N5736, N5724, N5050);
xor XOR2 (N5737, N5716, N3482);
nor NOR3 (N5738, N5697, N4547, N3980);
not NOT1 (N5739, N5738);
and AND3 (N5740, N5731, N1859, N231);
or OR4 (N5741, N5725, N5389, N2937, N2969);
and AND2 (N5742, N5739, N3581);
and AND4 (N5743, N5733, N5573, N1687, N1076);
nor NOR4 (N5744, N5742, N3871, N2168, N2176);
buf BUF1 (N5745, N5744);
and AND2 (N5746, N5732, N738);
and AND3 (N5747, N5735, N5552, N1185);
not NOT1 (N5748, N5746);
and AND4 (N5749, N5741, N5711, N3051, N3673);
or OR2 (N5750, N5726, N1850);
and AND3 (N5751, N5729, N4484, N2641);
nor NOR4 (N5752, N5747, N3215, N828, N4855);
or OR2 (N5753, N5751, N4868);
and AND4 (N5754, N5743, N3918, N1143, N3932);
nor NOR3 (N5755, N5745, N44, N2737);
not NOT1 (N5756, N5736);
and AND2 (N5757, N5755, N3860);
buf BUF1 (N5758, N5749);
and AND2 (N5759, N5737, N3406);
buf BUF1 (N5760, N5752);
buf BUF1 (N5761, N5758);
nor NOR4 (N5762, N5750, N3308, N5613, N166);
nor NOR3 (N5763, N5754, N302, N4501);
buf BUF1 (N5764, N5748);
not NOT1 (N5765, N5760);
or OR2 (N5766, N5763, N2204);
and AND2 (N5767, N5740, N1977);
buf BUF1 (N5768, N5765);
buf BUF1 (N5769, N5753);
xor XOR2 (N5770, N5756, N4771);
nor NOR3 (N5771, N5767, N1202, N5765);
buf BUF1 (N5772, N5769);
nand NAND4 (N5773, N5766, N3883, N12, N1469);
and AND3 (N5774, N5757, N690, N2470);
nand NAND3 (N5775, N5773, N1433, N574);
and AND4 (N5776, N5775, N2866, N4419, N3042);
or OR2 (N5777, N5770, N489);
nor NOR4 (N5778, N5762, N1684, N3380, N3529);
or OR3 (N5779, N5776, N5685, N756);
xor XOR2 (N5780, N5761, N5587);
nor NOR3 (N5781, N5777, N3948, N5671);
not NOT1 (N5782, N5778);
nand NAND2 (N5783, N5772, N2078);
buf BUF1 (N5784, N5768);
and AND3 (N5785, N5783, N3189, N4152);
xor XOR2 (N5786, N5771, N4356);
not NOT1 (N5787, N5785);
not NOT1 (N5788, N5786);
not NOT1 (N5789, N5779);
buf BUF1 (N5790, N5764);
buf BUF1 (N5791, N5790);
not NOT1 (N5792, N5789);
buf BUF1 (N5793, N5782);
not NOT1 (N5794, N5784);
xor XOR2 (N5795, N5788, N5364);
xor XOR2 (N5796, N5793, N3533);
not NOT1 (N5797, N5791);
xor XOR2 (N5798, N5795, N3419);
nor NOR3 (N5799, N5794, N3263, N2422);
nand NAND4 (N5800, N5798, N2387, N5408, N695);
and AND3 (N5801, N5780, N4175, N2336);
buf BUF1 (N5802, N5774);
xor XOR2 (N5803, N5799, N3841);
nor NOR4 (N5804, N5787, N1983, N2226, N2988);
and AND4 (N5805, N5792, N1266, N1621, N3083);
not NOT1 (N5806, N5802);
and AND2 (N5807, N5805, N3762);
nor NOR4 (N5808, N5759, N1941, N4091, N1165);
nand NAND3 (N5809, N5797, N1306, N5525);
nor NOR4 (N5810, N5804, N1779, N4478, N4458);
nor NOR2 (N5811, N5808, N2324);
xor XOR2 (N5812, N5806, N1083);
not NOT1 (N5813, N5810);
and AND2 (N5814, N5781, N495);
xor XOR2 (N5815, N5813, N317);
not NOT1 (N5816, N5803);
not NOT1 (N5817, N5809);
buf BUF1 (N5818, N5817);
buf BUF1 (N5819, N5812);
or OR4 (N5820, N5800, N4907, N709, N4178);
buf BUF1 (N5821, N5801);
or OR2 (N5822, N5821, N2806);
or OR3 (N5823, N5816, N4040, N5536);
not NOT1 (N5824, N5815);
and AND4 (N5825, N5818, N3967, N4949, N3753);
not NOT1 (N5826, N5824);
xor XOR2 (N5827, N5826, N2597);
nand NAND2 (N5828, N5822, N1805);
nor NOR2 (N5829, N5823, N5077);
not NOT1 (N5830, N5811);
xor XOR2 (N5831, N5796, N1878);
and AND3 (N5832, N5828, N4209, N2151);
buf BUF1 (N5833, N5831);
buf BUF1 (N5834, N5827);
not NOT1 (N5835, N5820);
xor XOR2 (N5836, N5807, N2637);
nand NAND4 (N5837, N5829, N3738, N5005, N5782);
nor NOR3 (N5838, N5832, N4736, N4905);
and AND4 (N5839, N5837, N1184, N3447, N2614);
buf BUF1 (N5840, N5825);
nor NOR3 (N5841, N5836, N1516, N4848);
xor XOR2 (N5842, N5841, N3309);
and AND3 (N5843, N5839, N5752, N997);
nand NAND2 (N5844, N5833, N2839);
buf BUF1 (N5845, N5842);
nand NAND3 (N5846, N5838, N475, N918);
buf BUF1 (N5847, N5814);
buf BUF1 (N5848, N5845);
and AND3 (N5849, N5840, N526, N240);
xor XOR2 (N5850, N5847, N335);
nor NOR3 (N5851, N5849, N1774, N3408);
nor NOR2 (N5852, N5835, N3579);
nand NAND2 (N5853, N5846, N1267);
and AND2 (N5854, N5844, N2333);
buf BUF1 (N5855, N5852);
and AND2 (N5856, N5853, N82);
nand NAND4 (N5857, N5850, N5049, N3205, N1017);
xor XOR2 (N5858, N5830, N1279);
and AND3 (N5859, N5851, N3867, N3852);
or OR3 (N5860, N5858, N427, N399);
not NOT1 (N5861, N5857);
nand NAND4 (N5862, N5834, N1292, N3817, N4985);
and AND2 (N5863, N5861, N4621);
not NOT1 (N5864, N5848);
xor XOR2 (N5865, N5843, N3435);
nand NAND2 (N5866, N5819, N4942);
not NOT1 (N5867, N5855);
xor XOR2 (N5868, N5867, N5508);
not NOT1 (N5869, N5862);
and AND2 (N5870, N5856, N1125);
xor XOR2 (N5871, N5860, N5642);
and AND4 (N5872, N5865, N4286, N1816, N4675);
not NOT1 (N5873, N5869);
or OR2 (N5874, N5870, N2202);
buf BUF1 (N5875, N5871);
and AND2 (N5876, N5864, N2058);
nand NAND4 (N5877, N5874, N623, N2114, N2044);
not NOT1 (N5878, N5875);
xor XOR2 (N5879, N5854, N4511);
or OR2 (N5880, N5877, N1526);
or OR4 (N5881, N5872, N4602, N2699, N1075);
xor XOR2 (N5882, N5866, N5114);
or OR4 (N5883, N5863, N3410, N4600, N5652);
nand NAND3 (N5884, N5873, N3569, N3880);
buf BUF1 (N5885, N5882);
not NOT1 (N5886, N5884);
nor NOR2 (N5887, N5868, N5267);
nor NOR3 (N5888, N5878, N4649, N731);
buf BUF1 (N5889, N5887);
not NOT1 (N5890, N5881);
and AND3 (N5891, N5879, N3060, N1668);
buf BUF1 (N5892, N5859);
not NOT1 (N5893, N5889);
nand NAND3 (N5894, N5876, N695, N4805);
or OR3 (N5895, N5885, N4697, N4245);
xor XOR2 (N5896, N5893, N2062);
nor NOR2 (N5897, N5883, N2278);
not NOT1 (N5898, N5892);
buf BUF1 (N5899, N5895);
buf BUF1 (N5900, N5886);
not NOT1 (N5901, N5899);
nand NAND4 (N5902, N5888, N4380, N1771, N2831);
not NOT1 (N5903, N5900);
buf BUF1 (N5904, N5902);
and AND3 (N5905, N5880, N5002, N1488);
buf BUF1 (N5906, N5905);
and AND4 (N5907, N5894, N971, N363, N2419);
or OR2 (N5908, N5901, N2638);
not NOT1 (N5909, N5903);
xor XOR2 (N5910, N5908, N5191);
nand NAND3 (N5911, N5890, N333, N2268);
or OR2 (N5912, N5910, N572);
buf BUF1 (N5913, N5909);
not NOT1 (N5914, N5911);
nor NOR2 (N5915, N5914, N3842);
and AND4 (N5916, N5915, N4394, N3920, N2713);
buf BUF1 (N5917, N5896);
not NOT1 (N5918, N5898);
nand NAND4 (N5919, N5891, N274, N3122, N3952);
not NOT1 (N5920, N5904);
xor XOR2 (N5921, N5906, N5069);
not NOT1 (N5922, N5912);
and AND3 (N5923, N5918, N4645, N2535);
or OR2 (N5924, N5919, N3487);
xor XOR2 (N5925, N5923, N1355);
nand NAND2 (N5926, N5916, N5694);
buf BUF1 (N5927, N5917);
and AND4 (N5928, N5897, N3126, N5849, N5401);
xor XOR2 (N5929, N5920, N1759);
not NOT1 (N5930, N5929);
or OR3 (N5931, N5924, N3869, N2781);
nor NOR2 (N5932, N5931, N2055);
xor XOR2 (N5933, N5907, N105);
or OR4 (N5934, N5921, N657, N784, N2544);
buf BUF1 (N5935, N5927);
nand NAND2 (N5936, N5932, N5139);
xor XOR2 (N5937, N5930, N2157);
or OR3 (N5938, N5913, N2117, N2548);
buf BUF1 (N5939, N5925);
xor XOR2 (N5940, N5939, N3454);
or OR2 (N5941, N5933, N4838);
not NOT1 (N5942, N5926);
buf BUF1 (N5943, N5934);
nand NAND3 (N5944, N5936, N5364, N349);
not NOT1 (N5945, N5928);
nor NOR3 (N5946, N5938, N4628, N348);
nor NOR4 (N5947, N5941, N4305, N4154, N3641);
buf BUF1 (N5948, N5947);
buf BUF1 (N5949, N5944);
buf BUF1 (N5950, N5942);
not NOT1 (N5951, N5945);
and AND3 (N5952, N5949, N4334, N560);
buf BUF1 (N5953, N5948);
buf BUF1 (N5954, N5950);
xor XOR2 (N5955, N5937, N4173);
nor NOR4 (N5956, N5953, N1611, N799, N2833);
or OR3 (N5957, N5922, N1031, N5777);
xor XOR2 (N5958, N5957, N1422);
nor NOR4 (N5959, N5954, N3481, N5554, N1758);
nor NOR4 (N5960, N5955, N1236, N2340, N1078);
buf BUF1 (N5961, N5956);
and AND2 (N5962, N5961, N840);
xor XOR2 (N5963, N5962, N4644);
xor XOR2 (N5964, N5943, N1681);
and AND2 (N5965, N5952, N3250);
and AND2 (N5966, N5959, N2160);
buf BUF1 (N5967, N5951);
and AND4 (N5968, N5935, N2034, N4357, N1798);
xor XOR2 (N5969, N5958, N4629);
and AND3 (N5970, N5965, N927, N4545);
nand NAND2 (N5971, N5964, N2424);
not NOT1 (N5972, N5970);
buf BUF1 (N5973, N5963);
xor XOR2 (N5974, N5973, N1579);
buf BUF1 (N5975, N5960);
and AND3 (N5976, N5967, N3126, N3673);
and AND2 (N5977, N5972, N1276);
and AND4 (N5978, N5966, N275, N2114, N5395);
or OR2 (N5979, N5976, N3243);
nand NAND4 (N5980, N5968, N5275, N5853, N4639);
nand NAND3 (N5981, N5946, N2512, N892);
buf BUF1 (N5982, N5971);
buf BUF1 (N5983, N5975);
or OR3 (N5984, N5977, N938, N2972);
and AND3 (N5985, N5969, N264, N4761);
or OR2 (N5986, N5974, N1442);
nor NOR2 (N5987, N5978, N3114);
and AND3 (N5988, N5982, N4965, N2565);
or OR2 (N5989, N5981, N4753);
xor XOR2 (N5990, N5980, N2585);
not NOT1 (N5991, N5989);
xor XOR2 (N5992, N5986, N894);
buf BUF1 (N5993, N5979);
xor XOR2 (N5994, N5991, N5079);
nand NAND3 (N5995, N5940, N5057, N4175);
or OR2 (N5996, N5984, N4408);
or OR3 (N5997, N5988, N4825, N1610);
nand NAND3 (N5998, N5993, N4339, N3695);
nand NAND4 (N5999, N5997, N4395, N2924, N5476);
buf BUF1 (N6000, N5990);
or OR4 (N6001, N5987, N2073, N2612, N177);
and AND4 (N6002, N5998, N5246, N254, N1893);
buf BUF1 (N6003, N5985);
buf BUF1 (N6004, N6000);
and AND4 (N6005, N6004, N793, N5958, N2820);
and AND3 (N6006, N6005, N3304, N2350);
nor NOR3 (N6007, N5992, N234, N3585);
or OR2 (N6008, N6001, N3261);
nand NAND4 (N6009, N5994, N3525, N4034, N4825);
and AND2 (N6010, N6002, N908);
nor NOR2 (N6011, N5983, N3147);
nor NOR3 (N6012, N5996, N3302, N204);
not NOT1 (N6013, N6003);
not NOT1 (N6014, N6013);
not NOT1 (N6015, N6010);
buf BUF1 (N6016, N6007);
xor XOR2 (N6017, N6009, N3373);
not NOT1 (N6018, N5995);
xor XOR2 (N6019, N6011, N2601);
xor XOR2 (N6020, N6008, N3926);
or OR4 (N6021, N6016, N2331, N2556, N4418);
and AND2 (N6022, N6019, N3137);
or OR4 (N6023, N6014, N5005, N5345, N5548);
xor XOR2 (N6024, N6023, N2603);
nand NAND2 (N6025, N6021, N2540);
buf BUF1 (N6026, N6018);
xor XOR2 (N6027, N6020, N637);
not NOT1 (N6028, N6027);
xor XOR2 (N6029, N6012, N1230);
nor NOR4 (N6030, N6024, N2512, N5986, N4779);
nand NAND2 (N6031, N6006, N2542);
xor XOR2 (N6032, N6025, N2768);
not NOT1 (N6033, N5999);
or OR3 (N6034, N6032, N4157, N2651);
not NOT1 (N6035, N6033);
nor NOR3 (N6036, N6015, N3906, N3106);
xor XOR2 (N6037, N6030, N4383);
or OR4 (N6038, N6017, N1875, N3838, N926);
and AND2 (N6039, N6029, N341);
nand NAND4 (N6040, N6028, N4407, N4997, N3656);
and AND3 (N6041, N6031, N5492, N4217);
nand NAND4 (N6042, N6022, N4272, N1904, N1877);
nor NOR2 (N6043, N6041, N5779);
nor NOR3 (N6044, N6042, N5545, N2416);
xor XOR2 (N6045, N6038, N1276);
nand NAND3 (N6046, N6045, N1407, N1396);
nor NOR4 (N6047, N6034, N2222, N3623, N3119);
buf BUF1 (N6048, N6026);
nor NOR2 (N6049, N6048, N5085);
buf BUF1 (N6050, N6046);
or OR2 (N6051, N6037, N701);
and AND4 (N6052, N6035, N472, N741, N2820);
or OR3 (N6053, N6047, N4410, N3758);
buf BUF1 (N6054, N6036);
not NOT1 (N6055, N6039);
or OR2 (N6056, N6049, N2858);
buf BUF1 (N6057, N6050);
nor NOR2 (N6058, N6044, N5579);
and AND2 (N6059, N6040, N3640);
and AND3 (N6060, N6051, N494, N1904);
nand NAND4 (N6061, N6058, N3308, N1491, N4321);
xor XOR2 (N6062, N6060, N1046);
buf BUF1 (N6063, N6057);
xor XOR2 (N6064, N6063, N2461);
buf BUF1 (N6065, N6053);
buf BUF1 (N6066, N6054);
xor XOR2 (N6067, N6064, N5890);
nor NOR3 (N6068, N6065, N3293, N1290);
and AND3 (N6069, N6061, N726, N4236);
and AND3 (N6070, N6066, N3674, N5932);
buf BUF1 (N6071, N6068);
nand NAND2 (N6072, N6056, N2076);
and AND2 (N6073, N6043, N1998);
xor XOR2 (N6074, N6073, N480);
or OR3 (N6075, N6055, N5037, N3366);
not NOT1 (N6076, N6062);
nand NAND2 (N6077, N6067, N3378);
and AND3 (N6078, N6059, N3149, N2304);
nand NAND3 (N6079, N6075, N1639, N1644);
nand NAND4 (N6080, N6078, N6068, N4722, N5024);
nor NOR2 (N6081, N6074, N2527);
nand NAND2 (N6082, N6052, N1726);
nor NOR3 (N6083, N6069, N3617, N2074);
or OR2 (N6084, N6080, N1873);
buf BUF1 (N6085, N6070);
nor NOR3 (N6086, N6083, N840, N5248);
buf BUF1 (N6087, N6072);
buf BUF1 (N6088, N6077);
not NOT1 (N6089, N6085);
or OR4 (N6090, N6071, N4520, N146, N741);
xor XOR2 (N6091, N6090, N821);
xor XOR2 (N6092, N6088, N3642);
nand NAND4 (N6093, N6081, N1416, N538, N5069);
nand NAND3 (N6094, N6079, N4155, N1044);
nor NOR2 (N6095, N6084, N4687);
xor XOR2 (N6096, N6095, N2141);
xor XOR2 (N6097, N6092, N4553);
nand NAND4 (N6098, N6093, N4387, N5905, N9);
or OR3 (N6099, N6097, N4119, N3557);
nand NAND2 (N6100, N6096, N4599);
not NOT1 (N6101, N6089);
buf BUF1 (N6102, N6082);
xor XOR2 (N6103, N6101, N709);
and AND4 (N6104, N6098, N1872, N2417, N1702);
nand NAND3 (N6105, N6102, N5267, N3790);
nand NAND2 (N6106, N6086, N144);
xor XOR2 (N6107, N6106, N2391);
xor XOR2 (N6108, N6100, N3289);
and AND2 (N6109, N6108, N2604);
xor XOR2 (N6110, N6104, N4482);
and AND4 (N6111, N6105, N5961, N4720, N1158);
nand NAND3 (N6112, N6111, N541, N3195);
or OR2 (N6113, N6110, N3802);
and AND2 (N6114, N6094, N6058);
and AND2 (N6115, N6091, N569);
xor XOR2 (N6116, N6114, N541);
or OR2 (N6117, N6115, N4667);
nor NOR3 (N6118, N6116, N2779, N1192);
nor NOR3 (N6119, N6109, N53, N5218);
or OR2 (N6120, N6119, N4126);
nand NAND4 (N6121, N6099, N3934, N1600, N4672);
or OR2 (N6122, N6076, N5646);
or OR4 (N6123, N6122, N5904, N4497, N5708);
and AND2 (N6124, N6118, N5752);
nor NOR2 (N6125, N6103, N2595);
and AND2 (N6126, N6087, N3704);
or OR3 (N6127, N6117, N4698, N5367);
xor XOR2 (N6128, N6113, N2832);
xor XOR2 (N6129, N6123, N1837);
and AND4 (N6130, N6124, N4001, N5379, N2760);
buf BUF1 (N6131, N6121);
xor XOR2 (N6132, N6129, N2727);
not NOT1 (N6133, N6132);
nand NAND2 (N6134, N6127, N1496);
or OR3 (N6135, N6131, N2438, N5531);
buf BUF1 (N6136, N6107);
xor XOR2 (N6137, N6120, N4561);
not NOT1 (N6138, N6133);
xor XOR2 (N6139, N6135, N3597);
not NOT1 (N6140, N6136);
nor NOR2 (N6141, N6128, N3788);
not NOT1 (N6142, N6130);
nand NAND4 (N6143, N6139, N872, N5461, N4016);
nor NOR2 (N6144, N6126, N2613);
and AND2 (N6145, N6144, N1663);
buf BUF1 (N6146, N6138);
nor NOR3 (N6147, N6143, N627, N3046);
not NOT1 (N6148, N6145);
nor NOR4 (N6149, N6137, N5544, N340, N814);
nor NOR3 (N6150, N6147, N568, N2771);
buf BUF1 (N6151, N6148);
or OR3 (N6152, N6140, N3007, N3025);
buf BUF1 (N6153, N6152);
not NOT1 (N6154, N6134);
buf BUF1 (N6155, N6153);
nor NOR3 (N6156, N6112, N1047, N5420);
and AND3 (N6157, N6141, N2419, N3079);
not NOT1 (N6158, N6150);
nand NAND2 (N6159, N6154, N2098);
and AND2 (N6160, N6149, N309);
xor XOR2 (N6161, N6156, N397);
nand NAND4 (N6162, N6160, N1570, N5757, N2580);
not NOT1 (N6163, N6142);
nand NAND3 (N6164, N6146, N3953, N379);
or OR2 (N6165, N6158, N5178);
nor NOR2 (N6166, N6161, N1748);
xor XOR2 (N6167, N6125, N991);
xor XOR2 (N6168, N6167, N2998);
or OR2 (N6169, N6157, N5150);
or OR3 (N6170, N6155, N4706, N5050);
nor NOR2 (N6171, N6170, N811);
xor XOR2 (N6172, N6162, N2985);
xor XOR2 (N6173, N6163, N424);
nor NOR2 (N6174, N6165, N2521);
and AND4 (N6175, N6168, N5617, N4428, N2864);
not NOT1 (N6176, N6151);
buf BUF1 (N6177, N6159);
and AND3 (N6178, N6171, N146, N1117);
not NOT1 (N6179, N6173);
buf BUF1 (N6180, N6169);
nor NOR2 (N6181, N6178, N5241);
and AND4 (N6182, N6177, N426, N4806, N5578);
or OR3 (N6183, N6175, N412, N3297);
buf BUF1 (N6184, N6179);
nand NAND2 (N6185, N6166, N2326);
or OR2 (N6186, N6172, N5848);
nand NAND2 (N6187, N6183, N3310);
buf BUF1 (N6188, N6187);
not NOT1 (N6189, N6186);
or OR2 (N6190, N6184, N3165);
xor XOR2 (N6191, N6164, N5082);
and AND4 (N6192, N6190, N4642, N4400, N871);
and AND3 (N6193, N6181, N3671, N4945);
not NOT1 (N6194, N6182);
or OR3 (N6195, N6188, N4971, N1932);
buf BUF1 (N6196, N6174);
and AND2 (N6197, N6180, N577);
or OR3 (N6198, N6176, N4956, N3796);
and AND3 (N6199, N6193, N5285, N4526);
nor NOR3 (N6200, N6194, N4146, N4798);
nand NAND2 (N6201, N6192, N1415);
or OR4 (N6202, N6197, N4158, N5376, N394);
nor NOR2 (N6203, N6201, N4537);
nand NAND3 (N6204, N6198, N1553, N877);
nor NOR3 (N6205, N6189, N2759, N4349);
nand NAND2 (N6206, N6185, N1262);
xor XOR2 (N6207, N6204, N5491);
buf BUF1 (N6208, N6207);
nor NOR4 (N6209, N6191, N4929, N5862, N290);
nand NAND3 (N6210, N6196, N1995, N1445);
not NOT1 (N6211, N6208);
nor NOR3 (N6212, N6199, N3830, N1487);
xor XOR2 (N6213, N6206, N4895);
buf BUF1 (N6214, N6200);
not NOT1 (N6215, N6211);
or OR3 (N6216, N6214, N3113, N1553);
or OR3 (N6217, N6215, N5958, N2170);
nor NOR2 (N6218, N6213, N3654);
or OR3 (N6219, N6205, N2900, N4739);
or OR4 (N6220, N6217, N790, N1082, N2739);
nand NAND3 (N6221, N6220, N6093, N1837);
or OR3 (N6222, N6219, N701, N4352);
not NOT1 (N6223, N6222);
and AND3 (N6224, N6210, N3746, N4188);
or OR3 (N6225, N6221, N341, N3454);
xor XOR2 (N6226, N6212, N5498);
buf BUF1 (N6227, N6216);
nor NOR3 (N6228, N6227, N4611, N2763);
or OR4 (N6229, N6203, N3375, N3849, N1399);
and AND2 (N6230, N6209, N533);
buf BUF1 (N6231, N6225);
and AND4 (N6232, N6202, N1660, N1153, N3518);
buf BUF1 (N6233, N6232);
or OR2 (N6234, N6226, N4093);
nor NOR2 (N6235, N6233, N5688);
and AND3 (N6236, N6234, N5029, N3835);
and AND2 (N6237, N6228, N5638);
nor NOR3 (N6238, N6218, N4799, N158);
not NOT1 (N6239, N6231);
nor NOR2 (N6240, N6229, N5770);
and AND3 (N6241, N6237, N6153, N4431);
or OR3 (N6242, N6223, N5449, N1038);
not NOT1 (N6243, N6240);
or OR2 (N6244, N6235, N5599);
xor XOR2 (N6245, N6239, N168);
or OR4 (N6246, N6195, N5644, N3941, N5950);
and AND2 (N6247, N6236, N1990);
xor XOR2 (N6248, N6245, N984);
nor NOR4 (N6249, N6242, N5489, N4359, N4226);
nor NOR4 (N6250, N6224, N5224, N3561, N429);
nor NOR2 (N6251, N6250, N1614);
xor XOR2 (N6252, N6244, N1955);
nand NAND2 (N6253, N6251, N3251);
xor XOR2 (N6254, N6230, N1923);
nor NOR2 (N6255, N6243, N3538);
xor XOR2 (N6256, N6248, N3407);
or OR4 (N6257, N6256, N5812, N2194, N650);
and AND4 (N6258, N6238, N3931, N2972, N4258);
and AND2 (N6259, N6252, N1894);
xor XOR2 (N6260, N6258, N6160);
nand NAND2 (N6261, N6257, N299);
or OR4 (N6262, N6260, N2290, N4556, N6002);
not NOT1 (N6263, N6249);
not NOT1 (N6264, N6247);
buf BUF1 (N6265, N6261);
not NOT1 (N6266, N6254);
nand NAND3 (N6267, N6264, N352, N4358);
nand NAND3 (N6268, N6265, N4468, N5021);
buf BUF1 (N6269, N6246);
or OR4 (N6270, N6255, N1380, N3619, N6237);
or OR3 (N6271, N6269, N159, N3849);
or OR2 (N6272, N6268, N2526);
nor NOR2 (N6273, N6263, N723);
and AND3 (N6274, N6272, N1233, N4696);
nand NAND3 (N6275, N6241, N5085, N5727);
and AND2 (N6276, N6253, N2872);
buf BUF1 (N6277, N6259);
xor XOR2 (N6278, N6277, N223);
or OR4 (N6279, N6275, N6266, N3746, N2851);
or OR4 (N6280, N1793, N4967, N5662, N1493);
nand NAND2 (N6281, N6280, N723);
not NOT1 (N6282, N6271);
or OR3 (N6283, N6279, N2106, N4951);
and AND2 (N6284, N6274, N900);
and AND3 (N6285, N6281, N221, N2382);
nor NOR4 (N6286, N6278, N2016, N1507, N178);
xor XOR2 (N6287, N6282, N4072);
and AND3 (N6288, N6286, N1051, N226);
nor NOR4 (N6289, N6273, N2907, N5618, N3123);
not NOT1 (N6290, N6283);
and AND2 (N6291, N6270, N2402);
not NOT1 (N6292, N6267);
xor XOR2 (N6293, N6287, N3755);
xor XOR2 (N6294, N6290, N5840);
nand NAND3 (N6295, N6285, N5929, N2393);
and AND2 (N6296, N6262, N2980);
nor NOR3 (N6297, N6289, N2834, N3450);
nand NAND2 (N6298, N6291, N869);
and AND2 (N6299, N6297, N5144);
nand NAND2 (N6300, N6295, N5028);
or OR4 (N6301, N6288, N361, N4191, N3881);
xor XOR2 (N6302, N6298, N4772);
and AND2 (N6303, N6293, N154);
xor XOR2 (N6304, N6302, N2476);
and AND3 (N6305, N6276, N5147, N5416);
buf BUF1 (N6306, N6304);
xor XOR2 (N6307, N6301, N2691);
buf BUF1 (N6308, N6284);
buf BUF1 (N6309, N6299);
and AND2 (N6310, N6305, N6297);
and AND4 (N6311, N6296, N2719, N5978, N6308);
not NOT1 (N6312, N4611);
not NOT1 (N6313, N6306);
and AND3 (N6314, N6300, N4500, N2606);
not NOT1 (N6315, N6294);
buf BUF1 (N6316, N6303);
buf BUF1 (N6317, N6310);
nand NAND2 (N6318, N6311, N2952);
and AND4 (N6319, N6317, N3723, N475, N1893);
nand NAND4 (N6320, N6314, N1554, N2489, N3331);
and AND3 (N6321, N6315, N58, N1965);
buf BUF1 (N6322, N6318);
or OR2 (N6323, N6322, N456);
xor XOR2 (N6324, N6321, N1191);
nor NOR3 (N6325, N6316, N4577, N3535);
not NOT1 (N6326, N6324);
nor NOR2 (N6327, N6323, N755);
and AND2 (N6328, N6326, N576);
nand NAND2 (N6329, N6313, N5965);
nor NOR3 (N6330, N6319, N1218, N312);
and AND4 (N6331, N6325, N4250, N4818, N5907);
not NOT1 (N6332, N6320);
nand NAND2 (N6333, N6327, N2799);
not NOT1 (N6334, N6312);
not NOT1 (N6335, N6328);
nor NOR3 (N6336, N6292, N223, N5427);
and AND2 (N6337, N6334, N4220);
nor NOR4 (N6338, N6330, N4833, N2304, N3289);
nand NAND3 (N6339, N6309, N3498, N4619);
nor NOR3 (N6340, N6336, N2363, N6027);
nand NAND4 (N6341, N6333, N2056, N6307, N4997);
not NOT1 (N6342, N4497);
xor XOR2 (N6343, N6332, N3672);
nand NAND4 (N6344, N6338, N4801, N2283, N680);
not NOT1 (N6345, N6340);
or OR4 (N6346, N6341, N4880, N5611, N61);
buf BUF1 (N6347, N6342);
not NOT1 (N6348, N6347);
xor XOR2 (N6349, N6331, N3792);
nor NOR3 (N6350, N6343, N190, N6244);
not NOT1 (N6351, N6346);
nor NOR3 (N6352, N6349, N5493, N4462);
or OR3 (N6353, N6344, N1933, N4527);
nand NAND4 (N6354, N6352, N190, N5886, N2626);
and AND4 (N6355, N6354, N4321, N205, N730);
or OR2 (N6356, N6353, N1611);
or OR2 (N6357, N6356, N5755);
and AND2 (N6358, N6335, N4449);
nor NOR2 (N6359, N6337, N2035);
not NOT1 (N6360, N6355);
xor XOR2 (N6361, N6357, N25);
nand NAND4 (N6362, N6360, N919, N2147, N3975);
nand NAND3 (N6363, N6358, N326, N817);
or OR4 (N6364, N6361, N874, N5847, N1729);
and AND4 (N6365, N6348, N2047, N278, N5572);
and AND3 (N6366, N6364, N124, N4276);
xor XOR2 (N6367, N6363, N449);
or OR2 (N6368, N6362, N314);
nor NOR2 (N6369, N6345, N4562);
or OR3 (N6370, N6351, N389, N5173);
or OR3 (N6371, N6339, N1566, N3000);
or OR2 (N6372, N6350, N1714);
or OR4 (N6373, N6367, N1325, N4417, N3749);
and AND4 (N6374, N6371, N5724, N5466, N4453);
or OR3 (N6375, N6372, N1216, N5379);
or OR3 (N6376, N6370, N4007, N124);
buf BUF1 (N6377, N6329);
nand NAND3 (N6378, N6359, N2243, N3787);
nand NAND4 (N6379, N6374, N5797, N194, N829);
buf BUF1 (N6380, N6376);
not NOT1 (N6381, N6378);
not NOT1 (N6382, N6366);
or OR4 (N6383, N6382, N4784, N4361, N2756);
nor NOR3 (N6384, N6373, N3816, N1159);
and AND3 (N6385, N6375, N5763, N25);
nand NAND3 (N6386, N6380, N4918, N5145);
buf BUF1 (N6387, N6377);
buf BUF1 (N6388, N6383);
and AND4 (N6389, N6379, N3746, N1667, N3354);
xor XOR2 (N6390, N6369, N3359);
or OR4 (N6391, N6387, N1566, N5780, N3470);
nand NAND2 (N6392, N6368, N578);
buf BUF1 (N6393, N6389);
not NOT1 (N6394, N6384);
nor NOR3 (N6395, N6393, N3330, N2969);
and AND3 (N6396, N6388, N3751, N71);
nand NAND3 (N6397, N6395, N1619, N4828);
and AND3 (N6398, N6396, N947, N512);
nor NOR4 (N6399, N6385, N3686, N6237, N4317);
not NOT1 (N6400, N6398);
nor NOR2 (N6401, N6391, N5719);
not NOT1 (N6402, N6399);
xor XOR2 (N6403, N6401, N1542);
xor XOR2 (N6404, N6400, N1512);
xor XOR2 (N6405, N6403, N5977);
nor NOR2 (N6406, N6405, N5983);
nor NOR3 (N6407, N6381, N3787, N3352);
nor NOR3 (N6408, N6406, N5280, N3268);
and AND4 (N6409, N6386, N254, N4577, N1176);
or OR2 (N6410, N6392, N474);
not NOT1 (N6411, N6402);
buf BUF1 (N6412, N6390);
and AND2 (N6413, N6394, N5125);
or OR2 (N6414, N6413, N6409);
nor NOR4 (N6415, N3033, N2148, N682, N6289);
buf BUF1 (N6416, N6411);
nand NAND4 (N6417, N6410, N5095, N545, N3302);
xor XOR2 (N6418, N6365, N3745);
nand NAND3 (N6419, N6414, N3798, N3859);
buf BUF1 (N6420, N6415);
nand NAND2 (N6421, N6404, N2584);
or OR4 (N6422, N6421, N6370, N5359, N4785);
xor XOR2 (N6423, N6418, N1815);
nand NAND2 (N6424, N6422, N6257);
or OR3 (N6425, N6419, N4814, N5033);
xor XOR2 (N6426, N6417, N3206);
or OR3 (N6427, N6423, N6288, N5207);
and AND4 (N6428, N6408, N2546, N1635, N1561);
not NOT1 (N6429, N6397);
or OR4 (N6430, N6412, N4677, N4964, N788);
or OR2 (N6431, N6420, N238);
not NOT1 (N6432, N6425);
not NOT1 (N6433, N6428);
nor NOR3 (N6434, N6433, N247, N5458);
nor NOR4 (N6435, N6430, N257, N1544, N4116);
and AND2 (N6436, N6435, N695);
nand NAND4 (N6437, N6429, N3307, N405, N3814);
or OR3 (N6438, N6427, N636, N1932);
nand NAND3 (N6439, N6437, N3121, N277);
buf BUF1 (N6440, N6438);
buf BUF1 (N6441, N6440);
nor NOR4 (N6442, N6439, N691, N3569, N4559);
xor XOR2 (N6443, N6436, N2463);
nand NAND3 (N6444, N6416, N3955, N6349);
xor XOR2 (N6445, N6434, N5371);
not NOT1 (N6446, N6441);
or OR2 (N6447, N6442, N86);
nand NAND3 (N6448, N6444, N6294, N5923);
nand NAND2 (N6449, N6445, N2334);
and AND2 (N6450, N6447, N3611);
nand NAND3 (N6451, N6443, N223, N522);
not NOT1 (N6452, N6450);
not NOT1 (N6453, N6451);
not NOT1 (N6454, N6453);
buf BUF1 (N6455, N6452);
nand NAND4 (N6456, N6454, N5039, N105, N4633);
and AND3 (N6457, N6448, N5752, N2074);
nor NOR3 (N6458, N6455, N3672, N56);
and AND2 (N6459, N6426, N138);
nor NOR3 (N6460, N6459, N3173, N889);
xor XOR2 (N6461, N6458, N4984);
nor NOR4 (N6462, N6407, N2264, N2071, N4521);
buf BUF1 (N6463, N6431);
buf BUF1 (N6464, N6446);
not NOT1 (N6465, N6449);
buf BUF1 (N6466, N6460);
nor NOR4 (N6467, N6466, N2749, N1917, N6296);
buf BUF1 (N6468, N6462);
nor NOR3 (N6469, N6465, N1707, N2163);
or OR4 (N6470, N6469, N3602, N5990, N370);
and AND2 (N6471, N6464, N1443);
xor XOR2 (N6472, N6424, N895);
not NOT1 (N6473, N6470);
buf BUF1 (N6474, N6473);
nor NOR4 (N6475, N6432, N302, N5496, N4042);
not NOT1 (N6476, N6471);
nor NOR2 (N6477, N6457, N1712);
nor NOR2 (N6478, N6461, N1762);
buf BUF1 (N6479, N6475);
or OR2 (N6480, N6472, N3425);
or OR2 (N6481, N6476, N3986);
buf BUF1 (N6482, N6479);
buf BUF1 (N6483, N6481);
and AND4 (N6484, N6483, N5635, N4381, N4883);
xor XOR2 (N6485, N6474, N2395);
nor NOR4 (N6486, N6467, N2622, N105, N3119);
or OR4 (N6487, N6485, N3221, N4353, N543);
nor NOR2 (N6488, N6478, N2880);
or OR2 (N6489, N6480, N4227);
nand NAND2 (N6490, N6489, N3644);
and AND4 (N6491, N6487, N6387, N1143, N6082);
and AND2 (N6492, N6490, N840);
buf BUF1 (N6493, N6486);
and AND2 (N6494, N6492, N5960);
buf BUF1 (N6495, N6491);
nor NOR4 (N6496, N6495, N4269, N1587, N3247);
buf BUF1 (N6497, N6468);
xor XOR2 (N6498, N6456, N2925);
nand NAND3 (N6499, N6496, N4479, N1999);
not NOT1 (N6500, N6477);
nor NOR2 (N6501, N6493, N3994);
nor NOR3 (N6502, N6484, N1839, N5618);
nor NOR4 (N6503, N6482, N2992, N1404, N1937);
or OR4 (N6504, N6500, N616, N4540, N4415);
xor XOR2 (N6505, N6463, N5564);
nand NAND3 (N6506, N6499, N2316, N1546);
nand NAND4 (N6507, N6505, N5558, N4577, N1347);
nand NAND4 (N6508, N6494, N3225, N3075, N6108);
nand NAND3 (N6509, N6504, N5804, N2248);
nor NOR4 (N6510, N6502, N1749, N3929, N2934);
not NOT1 (N6511, N6488);
buf BUF1 (N6512, N6503);
buf BUF1 (N6513, N6510);
not NOT1 (N6514, N6498);
nand NAND3 (N6515, N6509, N5892, N1245);
and AND3 (N6516, N6512, N2854, N1164);
not NOT1 (N6517, N6514);
nor NOR2 (N6518, N6497, N4420);
not NOT1 (N6519, N6507);
nand NAND4 (N6520, N6518, N5878, N675, N5224);
nor NOR3 (N6521, N6517, N2907, N4558);
xor XOR2 (N6522, N6508, N5310);
buf BUF1 (N6523, N6501);
nor NOR3 (N6524, N6513, N5545, N1868);
nand NAND4 (N6525, N6511, N4616, N3564, N6043);
or OR3 (N6526, N6516, N5076, N5796);
not NOT1 (N6527, N6519);
or OR4 (N6528, N6525, N4358, N5091, N5747);
and AND2 (N6529, N6526, N286);
not NOT1 (N6530, N6521);
nand NAND4 (N6531, N6515, N4536, N2597, N1587);
buf BUF1 (N6532, N6523);
xor XOR2 (N6533, N6532, N2447);
or OR3 (N6534, N6524, N1921, N896);
and AND4 (N6535, N6529, N4880, N2268, N6410);
not NOT1 (N6536, N6528);
nand NAND4 (N6537, N6535, N4516, N121, N3798);
nor NOR4 (N6538, N6533, N3486, N5282, N80);
nor NOR3 (N6539, N6531, N2237, N3166);
nand NAND2 (N6540, N6506, N5774);
nand NAND4 (N6541, N6527, N4772, N1532, N1002);
buf BUF1 (N6542, N6538);
buf BUF1 (N6543, N6522);
nor NOR2 (N6544, N6542, N340);
buf BUF1 (N6545, N6541);
or OR3 (N6546, N6537, N3347, N5856);
nand NAND3 (N6547, N6544, N3911, N4618);
not NOT1 (N6548, N6520);
or OR4 (N6549, N6548, N6047, N3348, N5805);
not NOT1 (N6550, N6546);
and AND2 (N6551, N6536, N1427);
or OR4 (N6552, N6530, N3629, N4352, N2747);
buf BUF1 (N6553, N6534);
or OR2 (N6554, N6551, N962);
nor NOR2 (N6555, N6552, N3555);
nor NOR4 (N6556, N6547, N2560, N1848, N1894);
buf BUF1 (N6557, N6556);
not NOT1 (N6558, N6549);
nor NOR2 (N6559, N6545, N636);
or OR2 (N6560, N6539, N78);
buf BUF1 (N6561, N6554);
nand NAND2 (N6562, N6557, N4929);
nand NAND4 (N6563, N6558, N3022, N3822, N6323);
or OR4 (N6564, N6543, N5773, N6188, N2560);
buf BUF1 (N6565, N6540);
not NOT1 (N6566, N6560);
not NOT1 (N6567, N6559);
nor NOR3 (N6568, N6564, N5098, N4841);
not NOT1 (N6569, N6550);
buf BUF1 (N6570, N6553);
xor XOR2 (N6571, N6563, N1097);
or OR3 (N6572, N6555, N3481, N6367);
not NOT1 (N6573, N6567);
xor XOR2 (N6574, N6572, N4027);
nor NOR2 (N6575, N6566, N5368);
not NOT1 (N6576, N6575);
and AND4 (N6577, N6576, N1290, N1736, N2614);
not NOT1 (N6578, N6574);
xor XOR2 (N6579, N6565, N1021);
not NOT1 (N6580, N6561);
buf BUF1 (N6581, N6569);
nand NAND4 (N6582, N6578, N914, N3453, N1960);
xor XOR2 (N6583, N6570, N3878);
and AND2 (N6584, N6577, N1533);
nor NOR3 (N6585, N6568, N2231, N5087);
nor NOR2 (N6586, N6562, N1622);
and AND4 (N6587, N6583, N969, N434, N5838);
buf BUF1 (N6588, N6573);
not NOT1 (N6589, N6585);
and AND3 (N6590, N6587, N1094, N2857);
xor XOR2 (N6591, N6571, N2905);
nand NAND2 (N6592, N6591, N4586);
or OR2 (N6593, N6586, N3477);
nand NAND2 (N6594, N6582, N1564);
and AND4 (N6595, N6593, N978, N1739, N5184);
and AND3 (N6596, N6580, N985, N4537);
not NOT1 (N6597, N6579);
and AND3 (N6598, N6597, N5089, N837);
buf BUF1 (N6599, N6595);
nand NAND4 (N6600, N6594, N5181, N6473, N262);
or OR4 (N6601, N6590, N2659, N3123, N1673);
nor NOR4 (N6602, N6581, N2516, N2128, N4766);
buf BUF1 (N6603, N6600);
xor XOR2 (N6604, N6584, N484);
xor XOR2 (N6605, N6596, N6324);
and AND3 (N6606, N6602, N6262, N1888);
buf BUF1 (N6607, N6604);
and AND4 (N6608, N6606, N4483, N4115, N3473);
xor XOR2 (N6609, N6592, N4785);
buf BUF1 (N6610, N6605);
or OR2 (N6611, N6598, N1094);
buf BUF1 (N6612, N6601);
xor XOR2 (N6613, N6599, N2238);
or OR4 (N6614, N6603, N4324, N6335, N5397);
not NOT1 (N6615, N6613);
or OR3 (N6616, N6609, N6402, N4293);
buf BUF1 (N6617, N6610);
nand NAND2 (N6618, N6616, N5946);
nand NAND4 (N6619, N6589, N4062, N3408, N5450);
or OR4 (N6620, N6608, N2028, N1036, N4534);
not NOT1 (N6621, N6614);
or OR3 (N6622, N6611, N2153, N5597);
buf BUF1 (N6623, N6620);
nor NOR3 (N6624, N6621, N6286, N1246);
not NOT1 (N6625, N6615);
xor XOR2 (N6626, N6625, N4792);
nor NOR3 (N6627, N6619, N6544, N165);
and AND3 (N6628, N6626, N5670, N4603);
xor XOR2 (N6629, N6618, N4045);
not NOT1 (N6630, N6617);
buf BUF1 (N6631, N6612);
xor XOR2 (N6632, N6624, N1297);
xor XOR2 (N6633, N6629, N3440);
not NOT1 (N6634, N6627);
buf BUF1 (N6635, N6622);
nor NOR3 (N6636, N6631, N1969, N6192);
nor NOR4 (N6637, N6635, N5663, N5381, N5486);
and AND3 (N6638, N6623, N1716, N1676);
and AND4 (N6639, N6630, N3707, N5036, N166);
not NOT1 (N6640, N6634);
nor NOR2 (N6641, N6628, N4872);
buf BUF1 (N6642, N6638);
and AND3 (N6643, N6641, N5405, N2675);
and AND2 (N6644, N6636, N205);
not NOT1 (N6645, N6642);
nand NAND3 (N6646, N6643, N1718, N2386);
not NOT1 (N6647, N6639);
xor XOR2 (N6648, N6632, N2427);
xor XOR2 (N6649, N6644, N5726);
not NOT1 (N6650, N6637);
xor XOR2 (N6651, N6633, N4709);
or OR2 (N6652, N6649, N5725);
or OR4 (N6653, N6588, N3330, N316, N2130);
nand NAND2 (N6654, N6607, N651);
xor XOR2 (N6655, N6654, N2791);
not NOT1 (N6656, N6651);
and AND2 (N6657, N6640, N1539);
nor NOR3 (N6658, N6648, N6009, N3824);
buf BUF1 (N6659, N6650);
and AND2 (N6660, N6645, N5592);
and AND4 (N6661, N6659, N3601, N6462, N3314);
buf BUF1 (N6662, N6652);
not NOT1 (N6663, N6662);
nor NOR4 (N6664, N6663, N2783, N1066, N5379);
or OR4 (N6665, N6653, N6176, N3625, N960);
or OR2 (N6666, N6661, N3515);
and AND2 (N6667, N6655, N2950);
buf BUF1 (N6668, N6647);
or OR4 (N6669, N6664, N1892, N3470, N4233);
xor XOR2 (N6670, N6658, N455);
not NOT1 (N6671, N6665);
buf BUF1 (N6672, N6660);
not NOT1 (N6673, N6666);
buf BUF1 (N6674, N6670);
and AND3 (N6675, N6657, N1315, N2893);
nor NOR4 (N6676, N6667, N2466, N4448, N5197);
xor XOR2 (N6677, N6673, N5837);
xor XOR2 (N6678, N6677, N5559);
buf BUF1 (N6679, N6668);
and AND2 (N6680, N6674, N491);
xor XOR2 (N6681, N6672, N3660);
not NOT1 (N6682, N6671);
not NOT1 (N6683, N6656);
buf BUF1 (N6684, N6681);
nor NOR3 (N6685, N6678, N5559, N4130);
not NOT1 (N6686, N6669);
xor XOR2 (N6687, N6679, N6553);
xor XOR2 (N6688, N6684, N6389);
not NOT1 (N6689, N6682);
nand NAND3 (N6690, N6646, N3946, N1349);
not NOT1 (N6691, N6683);
nand NAND2 (N6692, N6675, N4423);
nor NOR2 (N6693, N6689, N2390);
nand NAND4 (N6694, N6680, N3197, N5080, N129);
or OR3 (N6695, N6694, N4828, N1985);
buf BUF1 (N6696, N6692);
nand NAND4 (N6697, N6685, N5769, N5368, N6241);
or OR3 (N6698, N6696, N5421, N3663);
and AND3 (N6699, N6690, N695, N6505);
and AND2 (N6700, N6691, N66);
nand NAND4 (N6701, N6700, N6352, N529, N3220);
xor XOR2 (N6702, N6687, N1625);
xor XOR2 (N6703, N6697, N3880);
nand NAND4 (N6704, N6676, N1470, N4618, N528);
nor NOR3 (N6705, N6704, N3891, N3844);
xor XOR2 (N6706, N6701, N6312);
nor NOR4 (N6707, N6693, N2227, N5989, N6480);
nor NOR3 (N6708, N6686, N3714, N2661);
xor XOR2 (N6709, N6708, N5373);
xor XOR2 (N6710, N6705, N467);
not NOT1 (N6711, N6699);
not NOT1 (N6712, N6706);
xor XOR2 (N6713, N6710, N5258);
xor XOR2 (N6714, N6711, N1194);
nor NOR4 (N6715, N6688, N492, N1214, N1178);
not NOT1 (N6716, N6698);
not NOT1 (N6717, N6695);
xor XOR2 (N6718, N6707, N3343);
or OR2 (N6719, N6703, N6021);
nor NOR4 (N6720, N6714, N3704, N5778, N2548);
nand NAND2 (N6721, N6718, N1972);
not NOT1 (N6722, N6716);
xor XOR2 (N6723, N6715, N4927);
nand NAND2 (N6724, N6720, N980);
or OR2 (N6725, N6723, N6197);
nor NOR3 (N6726, N6724, N786, N2857);
nand NAND4 (N6727, N6719, N3886, N3386, N6702);
and AND2 (N6728, N3427, N1061);
or OR4 (N6729, N6725, N1420, N2214, N4107);
not NOT1 (N6730, N6722);
nand NAND2 (N6731, N6726, N5563);
nand NAND2 (N6732, N6717, N3786);
nor NOR4 (N6733, N6712, N3119, N712, N4929);
nor NOR3 (N6734, N6713, N1134, N1399);
not NOT1 (N6735, N6730);
or OR3 (N6736, N6729, N6259, N4811);
buf BUF1 (N6737, N6734);
nand NAND2 (N6738, N6736, N5214);
nand NAND4 (N6739, N6738, N616, N6524, N2607);
xor XOR2 (N6740, N6739, N5898);
or OR3 (N6741, N6733, N140, N2734);
nand NAND3 (N6742, N6732, N5813, N3711);
and AND3 (N6743, N6740, N137, N2312);
nand NAND4 (N6744, N6731, N1586, N4680, N546);
or OR2 (N6745, N6728, N3035);
and AND2 (N6746, N6741, N5771);
and AND4 (N6747, N6744, N2009, N1255, N5937);
xor XOR2 (N6748, N6709, N878);
or OR3 (N6749, N6727, N5598, N3497);
not NOT1 (N6750, N6748);
nand NAND2 (N6751, N6735, N2847);
not NOT1 (N6752, N6721);
xor XOR2 (N6753, N6743, N4628);
xor XOR2 (N6754, N6742, N3138);
buf BUF1 (N6755, N6746);
or OR2 (N6756, N6754, N4919);
nor NOR2 (N6757, N6737, N6601);
or OR3 (N6758, N6753, N3629, N5593);
not NOT1 (N6759, N6749);
buf BUF1 (N6760, N6752);
or OR4 (N6761, N6747, N4036, N150, N6453);
nand NAND4 (N6762, N6761, N972, N3868, N5008);
not NOT1 (N6763, N6759);
buf BUF1 (N6764, N6757);
xor XOR2 (N6765, N6762, N3607);
buf BUF1 (N6766, N6765);
xor XOR2 (N6767, N6751, N2490);
nand NAND3 (N6768, N6756, N5221, N6263);
nand NAND3 (N6769, N6766, N1133, N1171);
buf BUF1 (N6770, N6767);
or OR2 (N6771, N6770, N5601);
buf BUF1 (N6772, N6750);
buf BUF1 (N6773, N6768);
nor NOR2 (N6774, N6763, N4779);
buf BUF1 (N6775, N6769);
nor NOR2 (N6776, N6764, N5862);
nand NAND2 (N6777, N6776, N2850);
or OR2 (N6778, N6745, N2557);
not NOT1 (N6779, N6758);
or OR3 (N6780, N6775, N1364, N5403);
nand NAND4 (N6781, N6774, N3, N4508, N2642);
or OR3 (N6782, N6777, N330, N6184);
and AND2 (N6783, N6771, N2474);
nor NOR4 (N6784, N6780, N509, N5708, N2021);
xor XOR2 (N6785, N6781, N124);
nor NOR3 (N6786, N6772, N5374, N389);
buf BUF1 (N6787, N6784);
nor NOR4 (N6788, N6782, N3660, N4325, N3554);
not NOT1 (N6789, N6755);
and AND3 (N6790, N6788, N3621, N1183);
not NOT1 (N6791, N6779);
nor NOR4 (N6792, N6789, N2338, N1992, N5216);
not NOT1 (N6793, N6786);
nor NOR2 (N6794, N6791, N862);
nor NOR3 (N6795, N6793, N4312, N3312);
or OR2 (N6796, N6783, N4869);
not NOT1 (N6797, N6794);
not NOT1 (N6798, N6797);
or OR3 (N6799, N6785, N4245, N5943);
not NOT1 (N6800, N6799);
or OR4 (N6801, N6787, N6492, N3959, N2771);
xor XOR2 (N6802, N6796, N917);
and AND4 (N6803, N6773, N5553, N5348, N3336);
buf BUF1 (N6804, N6778);
not NOT1 (N6805, N6798);
nand NAND2 (N6806, N6760, N1943);
nand NAND4 (N6807, N6805, N4251, N1214, N4936);
buf BUF1 (N6808, N6792);
and AND2 (N6809, N6802, N3877);
or OR3 (N6810, N6790, N2151, N6457);
not NOT1 (N6811, N6809);
or OR2 (N6812, N6810, N20);
buf BUF1 (N6813, N6812);
xor XOR2 (N6814, N6811, N290);
or OR3 (N6815, N6807, N4328, N791);
not NOT1 (N6816, N6804);
not NOT1 (N6817, N6816);
nor NOR4 (N6818, N6800, N5715, N1989, N4100);
nand NAND2 (N6819, N6813, N6458);
buf BUF1 (N6820, N6819);
xor XOR2 (N6821, N6818, N1869);
nand NAND2 (N6822, N6820, N1154);
nor NOR2 (N6823, N6814, N910);
and AND3 (N6824, N6823, N105, N2365);
nor NOR4 (N6825, N6795, N2834, N3597, N5434);
nand NAND2 (N6826, N6815, N1017);
or OR2 (N6827, N6826, N2798);
not NOT1 (N6828, N6821);
xor XOR2 (N6829, N6825, N6135);
xor XOR2 (N6830, N6803, N482);
nand NAND2 (N6831, N6806, N3339);
xor XOR2 (N6832, N6831, N54);
and AND4 (N6833, N6824, N1180, N3786, N2986);
nor NOR3 (N6834, N6822, N5432, N4345);
not NOT1 (N6835, N6832);
and AND4 (N6836, N6830, N5318, N3643, N3374);
buf BUF1 (N6837, N6808);
not NOT1 (N6838, N6833);
not NOT1 (N6839, N6835);
or OR4 (N6840, N6827, N1950, N888, N4617);
or OR3 (N6841, N6840, N4105, N6233);
nor NOR3 (N6842, N6817, N193, N5632);
not NOT1 (N6843, N6842);
nor NOR3 (N6844, N6834, N3503, N2428);
and AND2 (N6845, N6829, N6281);
buf BUF1 (N6846, N6843);
buf BUF1 (N6847, N6838);
xor XOR2 (N6848, N6828, N925);
and AND3 (N6849, N6845, N6674, N1922);
xor XOR2 (N6850, N6839, N1374);
nand NAND4 (N6851, N6849, N5989, N5834, N3875);
buf BUF1 (N6852, N6850);
not NOT1 (N6853, N6851);
nand NAND2 (N6854, N6846, N5128);
or OR4 (N6855, N6853, N845, N2390, N6621);
xor XOR2 (N6856, N6837, N4083);
not NOT1 (N6857, N6836);
and AND2 (N6858, N6841, N4595);
buf BUF1 (N6859, N6856);
xor XOR2 (N6860, N6858, N4838);
buf BUF1 (N6861, N6859);
xor XOR2 (N6862, N6861, N2426);
xor XOR2 (N6863, N6854, N2812);
and AND3 (N6864, N6863, N2275, N953);
xor XOR2 (N6865, N6852, N5475);
or OR2 (N6866, N6862, N6758);
not NOT1 (N6867, N6844);
xor XOR2 (N6868, N6864, N2303);
not NOT1 (N6869, N6860);
buf BUF1 (N6870, N6868);
not NOT1 (N6871, N6848);
buf BUF1 (N6872, N6866);
xor XOR2 (N6873, N6801, N1484);
or OR2 (N6874, N6869, N5617);
not NOT1 (N6875, N6867);
xor XOR2 (N6876, N6855, N695);
nor NOR4 (N6877, N6857, N3195, N2208, N4659);
or OR3 (N6878, N6874, N3916, N188);
buf BUF1 (N6879, N6877);
not NOT1 (N6880, N6870);
nand NAND4 (N6881, N6872, N1735, N3059, N3622);
xor XOR2 (N6882, N6878, N868);
nor NOR4 (N6883, N6847, N18, N3335, N3519);
xor XOR2 (N6884, N6881, N3965);
buf BUF1 (N6885, N6882);
nor NOR4 (N6886, N6879, N1794, N3999, N605);
xor XOR2 (N6887, N6876, N2139);
xor XOR2 (N6888, N6884, N2850);
nand NAND4 (N6889, N6880, N5357, N4438, N6578);
xor XOR2 (N6890, N6886, N40);
nand NAND3 (N6891, N6888, N2513, N3498);
nand NAND3 (N6892, N6889, N4411, N751);
not NOT1 (N6893, N6875);
and AND2 (N6894, N6865, N1657);
and AND2 (N6895, N6892, N5800);
nor NOR4 (N6896, N6893, N4989, N4653, N2890);
not NOT1 (N6897, N6887);
xor XOR2 (N6898, N6890, N340);
and AND4 (N6899, N6873, N541, N6185, N5897);
nor NOR2 (N6900, N6883, N2385);
not NOT1 (N6901, N6891);
xor XOR2 (N6902, N6871, N4665);
xor XOR2 (N6903, N6896, N2425);
or OR4 (N6904, N6894, N471, N2207, N2697);
not NOT1 (N6905, N6899);
nor NOR2 (N6906, N6902, N6084);
nor NOR3 (N6907, N6895, N1860, N4059);
nand NAND3 (N6908, N6906, N4124, N6119);
nor NOR4 (N6909, N6904, N5649, N3209, N3668);
nand NAND2 (N6910, N6885, N6352);
xor XOR2 (N6911, N6908, N3878);
buf BUF1 (N6912, N6903);
xor XOR2 (N6913, N6898, N3623);
nor NOR4 (N6914, N6910, N3650, N3388, N5440);
not NOT1 (N6915, N6905);
buf BUF1 (N6916, N6907);
or OR3 (N6917, N6913, N1128, N4882);
and AND3 (N6918, N6909, N1549, N4228);
nand NAND3 (N6919, N6901, N1640, N2629);
nand NAND2 (N6920, N6914, N6256);
xor XOR2 (N6921, N6919, N6672);
xor XOR2 (N6922, N6900, N4143);
and AND3 (N6923, N6915, N5488, N6698);
or OR3 (N6924, N6918, N5785, N641);
nand NAND3 (N6925, N6911, N1307, N3550);
not NOT1 (N6926, N6922);
xor XOR2 (N6927, N6920, N1460);
nand NAND2 (N6928, N6925, N1125);
or OR4 (N6929, N6916, N3356, N1539, N1897);
not NOT1 (N6930, N6928);
or OR2 (N6931, N6926, N2985);
not NOT1 (N6932, N6927);
or OR2 (N6933, N6912, N4754);
buf BUF1 (N6934, N6931);
or OR2 (N6935, N6917, N1065);
nor NOR4 (N6936, N6933, N5808, N4025, N3803);
nand NAND4 (N6937, N6897, N5750, N4426, N262);
nor NOR2 (N6938, N6929, N463);
and AND2 (N6939, N6937, N5691);
and AND4 (N6940, N6923, N6102, N1755, N5354);
buf BUF1 (N6941, N6940);
or OR2 (N6942, N6930, N3311);
buf BUF1 (N6943, N6941);
or OR4 (N6944, N6935, N3641, N5608, N6805);
buf BUF1 (N6945, N6924);
nand NAND3 (N6946, N6945, N6139, N1856);
or OR3 (N6947, N6932, N6052, N2659);
xor XOR2 (N6948, N6946, N1385);
and AND3 (N6949, N6921, N1929, N3629);
not NOT1 (N6950, N6944);
buf BUF1 (N6951, N6950);
buf BUF1 (N6952, N6951);
nand NAND4 (N6953, N6939, N2984, N5190, N5520);
xor XOR2 (N6954, N6953, N672);
buf BUF1 (N6955, N6948);
xor XOR2 (N6956, N6947, N3187);
not NOT1 (N6957, N6952);
xor XOR2 (N6958, N6956, N4000);
not NOT1 (N6959, N6954);
xor XOR2 (N6960, N6943, N2426);
buf BUF1 (N6961, N6959);
xor XOR2 (N6962, N6949, N2125);
buf BUF1 (N6963, N6962);
and AND4 (N6964, N6957, N3850, N2442, N7);
not NOT1 (N6965, N6961);
or OR4 (N6966, N6955, N5921, N4295, N939);
or OR2 (N6967, N6960, N2875);
buf BUF1 (N6968, N6936);
or OR4 (N6969, N6934, N5329, N4130, N717);
buf BUF1 (N6970, N6963);
and AND2 (N6971, N6958, N6330);
buf BUF1 (N6972, N6942);
or OR3 (N6973, N6966, N955, N6893);
nor NOR2 (N6974, N6968, N25);
not NOT1 (N6975, N6971);
xor XOR2 (N6976, N6965, N3876);
xor XOR2 (N6977, N6973, N6546);
xor XOR2 (N6978, N6967, N336);
xor XOR2 (N6979, N6969, N119);
nand NAND2 (N6980, N6938, N3875);
not NOT1 (N6981, N6980);
not NOT1 (N6982, N6974);
and AND4 (N6983, N6976, N5148, N1014, N2971);
and AND3 (N6984, N6972, N1338, N1182);
nor NOR4 (N6985, N6975, N5524, N128, N5410);
buf BUF1 (N6986, N6964);
or OR4 (N6987, N6977, N894, N1867, N2183);
and AND3 (N6988, N6981, N1283, N659);
nand NAND2 (N6989, N6982, N4814);
nor NOR3 (N6990, N6986, N980, N5232);
not NOT1 (N6991, N6988);
buf BUF1 (N6992, N6987);
nand NAND4 (N6993, N6992, N3411, N5164, N6900);
or OR2 (N6994, N6983, N2213);
or OR3 (N6995, N6994, N5727, N2692);
not NOT1 (N6996, N6991);
or OR4 (N6997, N6984, N1077, N5698, N6708);
or OR3 (N6998, N6997, N1301, N4939);
and AND2 (N6999, N6996, N606);
and AND3 (N7000, N6998, N4951, N3918);
not NOT1 (N7001, N6993);
nand NAND3 (N7002, N6990, N5074, N5802);
buf BUF1 (N7003, N6989);
and AND2 (N7004, N6979, N5892);
xor XOR2 (N7005, N7003, N1091);
xor XOR2 (N7006, N7002, N6145);
nand NAND2 (N7007, N7001, N3521);
or OR4 (N7008, N7000, N3199, N3774, N6111);
or OR3 (N7009, N7004, N196, N6040);
and AND4 (N7010, N6999, N1147, N6104, N6339);
or OR3 (N7011, N7010, N3538, N1678);
and AND4 (N7012, N7009, N1736, N6848, N6439);
xor XOR2 (N7013, N7006, N5597);
nand NAND2 (N7014, N7005, N6890);
or OR4 (N7015, N7013, N5584, N2791, N4105);
buf BUF1 (N7016, N6995);
nand NAND4 (N7017, N7016, N4597, N3776, N3167);
nor NOR4 (N7018, N7012, N5864, N2761, N236);
buf BUF1 (N7019, N7007);
nor NOR3 (N7020, N7014, N159, N1974);
buf BUF1 (N7021, N7015);
not NOT1 (N7022, N7017);
nand NAND3 (N7023, N6985, N2645, N863);
not NOT1 (N7024, N7019);
buf BUF1 (N7025, N7021);
xor XOR2 (N7026, N7011, N3406);
buf BUF1 (N7027, N6978);
xor XOR2 (N7028, N7024, N6214);
or OR2 (N7029, N7020, N941);
or OR2 (N7030, N7022, N4946);
nand NAND4 (N7031, N7030, N3338, N4912, N6462);
or OR4 (N7032, N7028, N4434, N315, N5712);
and AND3 (N7033, N7031, N1427, N2054);
xor XOR2 (N7034, N7033, N5217);
xor XOR2 (N7035, N7034, N4930);
nor NOR2 (N7036, N7035, N5876);
or OR2 (N7037, N7023, N2980);
or OR2 (N7038, N7029, N727);
nor NOR3 (N7039, N7018, N6160, N5762);
not NOT1 (N7040, N7027);
xor XOR2 (N7041, N7040, N3199);
buf BUF1 (N7042, N7036);
xor XOR2 (N7043, N7038, N4638);
buf BUF1 (N7044, N7039);
and AND4 (N7045, N7044, N694, N704, N4397);
buf BUF1 (N7046, N7041);
buf BUF1 (N7047, N7008);
nand NAND4 (N7048, N7046, N4601, N5360, N6231);
buf BUF1 (N7049, N7025);
and AND3 (N7050, N7047, N6514, N5096);
and AND3 (N7051, N7049, N7008, N2746);
not NOT1 (N7052, N6970);
buf BUF1 (N7053, N7026);
buf BUF1 (N7054, N7048);
and AND2 (N7055, N7051, N737);
xor XOR2 (N7056, N7053, N4912);
xor XOR2 (N7057, N7056, N2467);
not NOT1 (N7058, N7042);
buf BUF1 (N7059, N7032);
nor NOR3 (N7060, N7055, N2391, N2069);
xor XOR2 (N7061, N7057, N4282);
or OR2 (N7062, N7043, N6089);
buf BUF1 (N7063, N7054);
xor XOR2 (N7064, N7045, N2183);
xor XOR2 (N7065, N7060, N2369);
or OR2 (N7066, N7062, N2330);
nor NOR2 (N7067, N7058, N4168);
nand NAND3 (N7068, N7052, N5149, N3238);
buf BUF1 (N7069, N7064);
nor NOR2 (N7070, N7067, N593);
nand NAND3 (N7071, N7066, N3505, N3609);
buf BUF1 (N7072, N7050);
nand NAND4 (N7073, N7037, N5232, N2439, N1449);
nor NOR2 (N7074, N7071, N5458);
xor XOR2 (N7075, N7059, N5358);
xor XOR2 (N7076, N7069, N2304);
not NOT1 (N7077, N7063);
nand NAND4 (N7078, N7072, N3370, N3620, N1444);
xor XOR2 (N7079, N7073, N6934);
nor NOR4 (N7080, N7065, N3142, N6282, N2622);
nand NAND2 (N7081, N7080, N1726);
buf BUF1 (N7082, N7076);
and AND2 (N7083, N7061, N2938);
or OR2 (N7084, N7070, N1385);
not NOT1 (N7085, N7077);
not NOT1 (N7086, N7084);
and AND3 (N7087, N7081, N1436, N4321);
not NOT1 (N7088, N7087);
or OR4 (N7089, N7088, N4680, N2154, N4320);
buf BUF1 (N7090, N7079);
not NOT1 (N7091, N7082);
nand NAND3 (N7092, N7083, N6179, N1952);
and AND3 (N7093, N7075, N1835, N3907);
nand NAND4 (N7094, N7091, N1541, N3320, N3008);
xor XOR2 (N7095, N7094, N4133);
not NOT1 (N7096, N7078);
and AND4 (N7097, N7095, N4432, N3027, N1813);
nand NAND4 (N7098, N7096, N1022, N4512, N126);
and AND3 (N7099, N7074, N2701, N5376);
or OR3 (N7100, N7086, N3492, N857);
xor XOR2 (N7101, N7099, N4799);
nand NAND3 (N7102, N7085, N6138, N3593);
buf BUF1 (N7103, N7097);
buf BUF1 (N7104, N7102);
nor NOR4 (N7105, N7101, N129, N3134, N7048);
buf BUF1 (N7106, N7105);
or OR4 (N7107, N7106, N3681, N4142, N2087);
or OR3 (N7108, N7092, N2368, N4917);
not NOT1 (N7109, N7103);
xor XOR2 (N7110, N7089, N1399);
not NOT1 (N7111, N7109);
buf BUF1 (N7112, N7107);
and AND2 (N7113, N7110, N1603);
not NOT1 (N7114, N7098);
xor XOR2 (N7115, N7114, N6652);
and AND3 (N7116, N7115, N578, N1816);
not NOT1 (N7117, N7116);
buf BUF1 (N7118, N7111);
nor NOR3 (N7119, N7100, N6708, N4136);
xor XOR2 (N7120, N7104, N6455);
not NOT1 (N7121, N7112);
and AND4 (N7122, N7117, N4989, N721, N4745);
not NOT1 (N7123, N7121);
not NOT1 (N7124, N7108);
nand NAND4 (N7125, N7090, N7082, N3139, N2501);
and AND4 (N7126, N7068, N4591, N6677, N5866);
nand NAND2 (N7127, N7124, N6978);
xor XOR2 (N7128, N7125, N725);
nor NOR3 (N7129, N7128, N898, N5332);
xor XOR2 (N7130, N7093, N484);
xor XOR2 (N7131, N7118, N2170);
nand NAND2 (N7132, N7127, N6354);
nor NOR2 (N7133, N7131, N2133);
buf BUF1 (N7134, N7132);
not NOT1 (N7135, N7119);
or OR4 (N7136, N7126, N6682, N4915, N6973);
not NOT1 (N7137, N7122);
buf BUF1 (N7138, N7130);
xor XOR2 (N7139, N7136, N1928);
and AND3 (N7140, N7129, N5508, N6578);
buf BUF1 (N7141, N7120);
nor NOR2 (N7142, N7113, N6026);
nand NAND4 (N7143, N7123, N5699, N5561, N359);
or OR3 (N7144, N7138, N6530, N1108);
nor NOR2 (N7145, N7144, N2372);
or OR4 (N7146, N7137, N5048, N6820, N3494);
and AND4 (N7147, N7133, N360, N6129, N3042);
xor XOR2 (N7148, N7140, N5104);
nor NOR4 (N7149, N7134, N6515, N3108, N6185);
nor NOR4 (N7150, N7139, N38, N1247, N5140);
or OR2 (N7151, N7142, N3286);
nand NAND3 (N7152, N7146, N6518, N4156);
or OR4 (N7153, N7135, N5324, N5253, N3574);
or OR3 (N7154, N7143, N6506, N2645);
buf BUF1 (N7155, N7150);
and AND2 (N7156, N7154, N687);
not NOT1 (N7157, N7152);
and AND2 (N7158, N7155, N3417);
not NOT1 (N7159, N7148);
and AND4 (N7160, N7153, N3018, N5835, N5553);
or OR3 (N7161, N7158, N3142, N2452);
buf BUF1 (N7162, N7141);
nor NOR3 (N7163, N7160, N1161, N3530);
or OR4 (N7164, N7163, N3962, N5468, N1177);
buf BUF1 (N7165, N7145);
nand NAND2 (N7166, N7159, N833);
nor NOR4 (N7167, N7161, N5708, N1064, N1330);
nor NOR4 (N7168, N7164, N236, N6709, N3147);
nor NOR4 (N7169, N7168, N7019, N4629, N3288);
nor NOR3 (N7170, N7165, N5024, N3463);
xor XOR2 (N7171, N7157, N1899);
or OR3 (N7172, N7156, N753, N5650);
or OR3 (N7173, N7171, N4067, N190);
and AND4 (N7174, N7170, N4886, N2465, N3517);
not NOT1 (N7175, N7147);
xor XOR2 (N7176, N7167, N4286);
xor XOR2 (N7177, N7162, N607);
nand NAND4 (N7178, N7175, N4023, N2705, N1214);
nand NAND3 (N7179, N7173, N449, N29);
and AND3 (N7180, N7166, N910, N6826);
not NOT1 (N7181, N7180);
and AND3 (N7182, N7169, N5918, N1839);
nand NAND2 (N7183, N7181, N2325);
and AND3 (N7184, N7151, N7107, N3506);
or OR2 (N7185, N7149, N5189);
and AND4 (N7186, N7182, N6218, N6962, N2162);
nand NAND4 (N7187, N7179, N1949, N674, N4486);
not NOT1 (N7188, N7184);
xor XOR2 (N7189, N7177, N3689);
buf BUF1 (N7190, N7183);
xor XOR2 (N7191, N7190, N3809);
or OR2 (N7192, N7188, N7191);
or OR4 (N7193, N5493, N6994, N221, N5493);
and AND3 (N7194, N7176, N5046, N1046);
and AND4 (N7195, N7192, N4658, N4072, N7170);
buf BUF1 (N7196, N7172);
nand NAND4 (N7197, N7194, N655, N3101, N3093);
or OR2 (N7198, N7174, N4181);
xor XOR2 (N7199, N7178, N6720);
not NOT1 (N7200, N7187);
or OR4 (N7201, N7200, N2632, N6906, N1586);
or OR4 (N7202, N7186, N4629, N3239, N5621);
or OR4 (N7203, N7193, N1165, N3955, N1177);
buf BUF1 (N7204, N7199);
buf BUF1 (N7205, N7204);
not NOT1 (N7206, N7201);
xor XOR2 (N7207, N7197, N2234);
not NOT1 (N7208, N7206);
nor NOR3 (N7209, N7189, N711, N6095);
xor XOR2 (N7210, N7205, N5855);
nand NAND3 (N7211, N7195, N6324, N5432);
not NOT1 (N7212, N7208);
and AND2 (N7213, N7198, N2300);
or OR3 (N7214, N7213, N7021, N7116);
buf BUF1 (N7215, N7210);
xor XOR2 (N7216, N7207, N6125);
or OR4 (N7217, N7203, N3464, N1030, N5199);
xor XOR2 (N7218, N7212, N4216);
or OR4 (N7219, N7218, N1293, N5192, N4351);
nor NOR3 (N7220, N7196, N1103, N5460);
xor XOR2 (N7221, N7215, N353);
xor XOR2 (N7222, N7217, N3238);
nor NOR2 (N7223, N7211, N3986);
nand NAND3 (N7224, N7185, N6985, N2299);
or OR4 (N7225, N7220, N6084, N6801, N2490);
and AND3 (N7226, N7216, N2272, N803);
and AND4 (N7227, N7202, N4231, N6099, N4940);
and AND2 (N7228, N7222, N5715);
and AND2 (N7229, N7209, N6710);
and AND4 (N7230, N7223, N253, N6294, N2231);
xor XOR2 (N7231, N7226, N2406);
not NOT1 (N7232, N7229);
nand NAND4 (N7233, N7224, N6642, N1194, N3211);
and AND2 (N7234, N7214, N2012);
nand NAND4 (N7235, N7227, N2224, N4171, N267);
or OR3 (N7236, N7221, N7147, N5863);
nor NOR4 (N7237, N7219, N1007, N3915, N685);
xor XOR2 (N7238, N7235, N1342);
xor XOR2 (N7239, N7237, N5981);
or OR2 (N7240, N7225, N1995);
or OR4 (N7241, N7228, N3506, N5633, N6204);
nor NOR3 (N7242, N7232, N6466, N5382);
xor XOR2 (N7243, N7231, N7074);
nand NAND2 (N7244, N7243, N1681);
not NOT1 (N7245, N7240);
or OR2 (N7246, N7244, N5327);
and AND4 (N7247, N7236, N6667, N3877, N3058);
buf BUF1 (N7248, N7247);
nand NAND2 (N7249, N7239, N7196);
and AND3 (N7250, N7242, N2715, N2778);
nor NOR2 (N7251, N7246, N4127);
or OR3 (N7252, N7230, N5295, N3191);
not NOT1 (N7253, N7251);
not NOT1 (N7254, N7252);
or OR3 (N7255, N7248, N5557, N2694);
nor NOR3 (N7256, N7249, N1586, N1846);
or OR4 (N7257, N7238, N4365, N4392, N2664);
not NOT1 (N7258, N7253);
or OR3 (N7259, N7234, N2790, N3023);
or OR3 (N7260, N7241, N4251, N3385);
not NOT1 (N7261, N7259);
buf BUF1 (N7262, N7250);
nor NOR3 (N7263, N7256, N5330, N2782);
nor NOR2 (N7264, N7258, N2358);
or OR2 (N7265, N7245, N6066);
nand NAND4 (N7266, N7233, N1733, N4265, N6039);
buf BUF1 (N7267, N7263);
and AND2 (N7268, N7257, N4820);
and AND2 (N7269, N7260, N4453);
xor XOR2 (N7270, N7266, N2705);
xor XOR2 (N7271, N7262, N3554);
xor XOR2 (N7272, N7254, N2702);
nor NOR2 (N7273, N7265, N1879);
not NOT1 (N7274, N7269);
nor NOR2 (N7275, N7255, N7074);
xor XOR2 (N7276, N7271, N5285);
nand NAND4 (N7277, N7264, N4515, N3247, N4587);
nor NOR3 (N7278, N7274, N6211, N7152);
xor XOR2 (N7279, N7273, N7018);
nor NOR2 (N7280, N7276, N2478);
nand NAND4 (N7281, N7278, N7167, N2280, N6267);
buf BUF1 (N7282, N7281);
and AND3 (N7283, N7270, N5739, N3123);
xor XOR2 (N7284, N7279, N3907);
buf BUF1 (N7285, N7275);
or OR3 (N7286, N7272, N7038, N772);
nand NAND3 (N7287, N7261, N2132, N3498);
not NOT1 (N7288, N7267);
or OR3 (N7289, N7288, N3241, N1341);
nand NAND4 (N7290, N7289, N3503, N1539, N5143);
and AND2 (N7291, N7282, N336);
and AND3 (N7292, N7287, N1859, N2858);
buf BUF1 (N7293, N7277);
xor XOR2 (N7294, N7284, N1043);
nand NAND4 (N7295, N7285, N2032, N4936, N6639);
not NOT1 (N7296, N7293);
buf BUF1 (N7297, N7286);
nor NOR2 (N7298, N7280, N2591);
not NOT1 (N7299, N7295);
or OR2 (N7300, N7296, N2225);
buf BUF1 (N7301, N7298);
and AND3 (N7302, N7297, N176, N4037);
and AND3 (N7303, N7302, N1234, N400);
and AND3 (N7304, N7291, N4492, N1685);
nor NOR2 (N7305, N7283, N1648);
xor XOR2 (N7306, N7304, N2452);
nor NOR4 (N7307, N7290, N2098, N5758, N3999);
or OR3 (N7308, N7299, N586, N7188);
xor XOR2 (N7309, N7305, N4538);
buf BUF1 (N7310, N7300);
nand NAND4 (N7311, N7306, N1923, N4114, N5225);
xor XOR2 (N7312, N7311, N5259);
or OR2 (N7313, N7309, N2291);
xor XOR2 (N7314, N7312, N1738);
nand NAND2 (N7315, N7308, N6218);
xor XOR2 (N7316, N7294, N4671);
not NOT1 (N7317, N7301);
buf BUF1 (N7318, N7317);
nand NAND2 (N7319, N7268, N3723);
not NOT1 (N7320, N7314);
nand NAND4 (N7321, N7319, N2880, N3880, N3068);
and AND4 (N7322, N7307, N426, N599, N3935);
or OR3 (N7323, N7320, N2249, N3237);
buf BUF1 (N7324, N7315);
not NOT1 (N7325, N7323);
or OR3 (N7326, N7325, N2109, N7119);
not NOT1 (N7327, N7326);
not NOT1 (N7328, N7316);
xor XOR2 (N7329, N7327, N4879);
not NOT1 (N7330, N7329);
buf BUF1 (N7331, N7292);
buf BUF1 (N7332, N7328);
not NOT1 (N7333, N7321);
and AND2 (N7334, N7322, N5799);
or OR4 (N7335, N7310, N7296, N895, N2915);
nor NOR3 (N7336, N7331, N1398, N4156);
not NOT1 (N7337, N7313);
xor XOR2 (N7338, N7337, N299);
or OR4 (N7339, N7334, N3485, N3629, N7135);
buf BUF1 (N7340, N7335);
or OR4 (N7341, N7333, N1490, N398, N6387);
and AND2 (N7342, N7330, N67);
and AND3 (N7343, N7324, N1065, N5474);
or OR3 (N7344, N7332, N3170, N7331);
buf BUF1 (N7345, N7342);
nor NOR3 (N7346, N7341, N5412, N1417);
or OR4 (N7347, N7345, N2139, N1075, N4390);
nor NOR3 (N7348, N7343, N7096, N2165);
buf BUF1 (N7349, N7318);
nor NOR3 (N7350, N7346, N2222, N3690);
and AND3 (N7351, N7350, N3182, N4785);
or OR3 (N7352, N7349, N4486, N6249);
and AND2 (N7353, N7340, N576);
xor XOR2 (N7354, N7303, N3155);
not NOT1 (N7355, N7344);
not NOT1 (N7356, N7338);
buf BUF1 (N7357, N7336);
nand NAND3 (N7358, N7348, N4935, N6393);
not NOT1 (N7359, N7358);
and AND4 (N7360, N7359, N980, N2911, N5958);
not NOT1 (N7361, N7355);
and AND4 (N7362, N7347, N1846, N136, N5182);
nand NAND3 (N7363, N7352, N1232, N4757);
buf BUF1 (N7364, N7360);
buf BUF1 (N7365, N7339);
nor NOR3 (N7366, N7356, N1635, N6836);
and AND2 (N7367, N7366, N5363);
nor NOR4 (N7368, N7367, N3482, N1171, N4898);
nand NAND4 (N7369, N7357, N2203, N1964, N5910);
xor XOR2 (N7370, N7364, N6293);
nor NOR2 (N7371, N7365, N6418);
not NOT1 (N7372, N7363);
not NOT1 (N7373, N7369);
or OR2 (N7374, N7362, N1049);
nand NAND2 (N7375, N7351, N1283);
buf BUF1 (N7376, N7371);
not NOT1 (N7377, N7374);
nor NOR3 (N7378, N7373, N7278, N1460);
xor XOR2 (N7379, N7354, N3021);
or OR2 (N7380, N7368, N3383);
or OR2 (N7381, N7370, N372);
nand NAND3 (N7382, N7378, N967, N6450);
xor XOR2 (N7383, N7353, N2566);
and AND3 (N7384, N7380, N7059, N4604);
nor NOR3 (N7385, N7379, N5564, N552);
not NOT1 (N7386, N7381);
or OR4 (N7387, N7375, N712, N3512, N3526);
nor NOR3 (N7388, N7387, N894, N2321);
xor XOR2 (N7389, N7372, N6989);
and AND3 (N7390, N7383, N5404, N6793);
buf BUF1 (N7391, N7361);
xor XOR2 (N7392, N7391, N4622);
or OR2 (N7393, N7388, N209);
xor XOR2 (N7394, N7384, N216);
buf BUF1 (N7395, N7382);
xor XOR2 (N7396, N7389, N470);
xor XOR2 (N7397, N7393, N5497);
buf BUF1 (N7398, N7385);
xor XOR2 (N7399, N7390, N963);
and AND2 (N7400, N7395, N1278);
not NOT1 (N7401, N7400);
and AND2 (N7402, N7398, N7083);
not NOT1 (N7403, N7377);
and AND4 (N7404, N7403, N1504, N7223, N6781);
nand NAND2 (N7405, N7404, N2786);
buf BUF1 (N7406, N7386);
nand NAND4 (N7407, N7396, N2942, N6049, N6937);
and AND3 (N7408, N7405, N6289, N4151);
buf BUF1 (N7409, N7399);
nand NAND2 (N7410, N7394, N4535);
not NOT1 (N7411, N7402);
not NOT1 (N7412, N7410);
buf BUF1 (N7413, N7401);
and AND4 (N7414, N7409, N3675, N1253, N4910);
nand NAND3 (N7415, N7413, N3103, N5554);
xor XOR2 (N7416, N7376, N2009);
or OR3 (N7417, N7406, N3879, N2176);
or OR3 (N7418, N7412, N2261, N4709);
nor NOR4 (N7419, N7408, N111, N6694, N6030);
nor NOR2 (N7420, N7414, N3088);
nor NOR3 (N7421, N7415, N7059, N7411);
buf BUF1 (N7422, N2381);
not NOT1 (N7423, N7418);
xor XOR2 (N7424, N7416, N6077);
or OR2 (N7425, N7423, N279);
nand NAND2 (N7426, N7392, N503);
and AND3 (N7427, N7424, N3145, N3899);
buf BUF1 (N7428, N7427);
nand NAND3 (N7429, N7421, N6308, N6935);
nor NOR2 (N7430, N7429, N5670);
xor XOR2 (N7431, N7428, N7030);
and AND2 (N7432, N7426, N2080);
or OR3 (N7433, N7422, N3312, N4461);
xor XOR2 (N7434, N7420, N6665);
nand NAND4 (N7435, N7432, N1531, N6346, N2595);
buf BUF1 (N7436, N7407);
nor NOR3 (N7437, N7430, N4251, N3400);
nor NOR4 (N7438, N7436, N2397, N5648, N1678);
buf BUF1 (N7439, N7397);
and AND3 (N7440, N7437, N5476, N1379);
or OR2 (N7441, N7417, N2200);
or OR2 (N7442, N7419, N6920);
nor NOR3 (N7443, N7435, N1532, N2466);
buf BUF1 (N7444, N7434);
not NOT1 (N7445, N7439);
buf BUF1 (N7446, N7438);
nand NAND4 (N7447, N7446, N5760, N2694, N5035);
nand NAND2 (N7448, N7431, N1464);
nor NOR4 (N7449, N7445, N86, N6093, N888);
or OR3 (N7450, N7441, N5360, N1354);
not NOT1 (N7451, N7440);
buf BUF1 (N7452, N7448);
not NOT1 (N7453, N7450);
not NOT1 (N7454, N7447);
xor XOR2 (N7455, N7452, N6213);
nor NOR4 (N7456, N7454, N6191, N5803, N6123);
and AND3 (N7457, N7453, N6826, N3477);
or OR3 (N7458, N7433, N1521, N2035);
xor XOR2 (N7459, N7449, N2530);
xor XOR2 (N7460, N7455, N606);
xor XOR2 (N7461, N7460, N4675);
nand NAND3 (N7462, N7459, N4112, N1117);
or OR3 (N7463, N7461, N858, N157);
or OR4 (N7464, N7442, N6749, N3786, N353);
xor XOR2 (N7465, N7451, N4760);
xor XOR2 (N7466, N7465, N7324);
xor XOR2 (N7467, N7464, N4003);
and AND3 (N7468, N7458, N1903, N2469);
or OR2 (N7469, N7443, N4691);
nand NAND3 (N7470, N7425, N213, N4061);
or OR2 (N7471, N7470, N3017);
buf BUF1 (N7472, N7468);
xor XOR2 (N7473, N7467, N1201);
not NOT1 (N7474, N7456);
nor NOR2 (N7475, N7469, N6860);
xor XOR2 (N7476, N7471, N4099);
not NOT1 (N7477, N7462);
or OR3 (N7478, N7477, N2608, N3279);
not NOT1 (N7479, N7478);
nor NOR4 (N7480, N7475, N3081, N3135, N7119);
nor NOR4 (N7481, N7444, N3284, N3002, N3683);
buf BUF1 (N7482, N7466);
buf BUF1 (N7483, N7474);
nand NAND2 (N7484, N7476, N5030);
xor XOR2 (N7485, N7463, N5673);
nor NOR2 (N7486, N7480, N3178);
not NOT1 (N7487, N7486);
not NOT1 (N7488, N7472);
or OR3 (N7489, N7482, N4957, N1004);
or OR3 (N7490, N7489, N2370, N1467);
nor NOR3 (N7491, N7457, N3018, N3418);
and AND3 (N7492, N7488, N6102, N5048);
not NOT1 (N7493, N7491);
and AND3 (N7494, N7492, N1030, N3908);
and AND4 (N7495, N7485, N202, N3149, N6008);
and AND4 (N7496, N7487, N917, N2515, N6273);
or OR4 (N7497, N7481, N5316, N5528, N2274);
buf BUF1 (N7498, N7493);
nor NOR2 (N7499, N7497, N2359);
nand NAND3 (N7500, N7490, N1370, N4653);
nor NOR3 (N7501, N7499, N1029, N5837);
buf BUF1 (N7502, N7500);
nand NAND4 (N7503, N7498, N6233, N3920, N5853);
or OR2 (N7504, N7496, N6802);
not NOT1 (N7505, N7484);
not NOT1 (N7506, N7504);
nor NOR2 (N7507, N7505, N4089);
nor NOR2 (N7508, N7483, N5970);
nor NOR3 (N7509, N7479, N4874, N7013);
nand NAND2 (N7510, N7508, N3893);
and AND2 (N7511, N7501, N5470);
or OR4 (N7512, N7507, N6285, N7192, N2669);
and AND4 (N7513, N7473, N5573, N6393, N4552);
nand NAND3 (N7514, N7502, N2426, N6764);
buf BUF1 (N7515, N7511);
nand NAND3 (N7516, N7506, N2269, N2690);
and AND4 (N7517, N7494, N3363, N7292, N6879);
and AND2 (N7518, N7503, N3543);
nor NOR4 (N7519, N7517, N6359, N2457, N1164);
xor XOR2 (N7520, N7516, N1507);
xor XOR2 (N7521, N7495, N6598);
and AND3 (N7522, N7518, N7355, N3512);
and AND2 (N7523, N7522, N3819);
not NOT1 (N7524, N7513);
or OR2 (N7525, N7512, N1447);
buf BUF1 (N7526, N7514);
buf BUF1 (N7527, N7524);
not NOT1 (N7528, N7509);
xor XOR2 (N7529, N7525, N6998);
and AND4 (N7530, N7528, N2646, N7364, N6798);
xor XOR2 (N7531, N7527, N1304);
nor NOR4 (N7532, N7523, N5335, N2616, N480);
xor XOR2 (N7533, N7530, N1810);
or OR4 (N7534, N7521, N3746, N4455, N7044);
or OR2 (N7535, N7531, N2344);
xor XOR2 (N7536, N7515, N2563);
nand NAND2 (N7537, N7526, N3414);
nand NAND4 (N7538, N7532, N1750, N7067, N6376);
buf BUF1 (N7539, N7529);
or OR2 (N7540, N7537, N2482);
buf BUF1 (N7541, N7519);
or OR4 (N7542, N7510, N5853, N1472, N3167);
and AND2 (N7543, N7520, N7445);
and AND2 (N7544, N7533, N4761);
or OR2 (N7545, N7538, N4060);
or OR2 (N7546, N7536, N4256);
buf BUF1 (N7547, N7534);
nand NAND3 (N7548, N7543, N5311, N5825);
xor XOR2 (N7549, N7542, N656);
buf BUF1 (N7550, N7549);
not NOT1 (N7551, N7539);
and AND4 (N7552, N7541, N4729, N6370, N7462);
buf BUF1 (N7553, N7552);
buf BUF1 (N7554, N7546);
not NOT1 (N7555, N7554);
and AND3 (N7556, N7545, N5708, N4233);
or OR3 (N7557, N7556, N7505, N6489);
and AND3 (N7558, N7555, N3072, N1620);
not NOT1 (N7559, N7535);
nor NOR3 (N7560, N7544, N7471, N5275);
xor XOR2 (N7561, N7540, N6532);
nand NAND2 (N7562, N7557, N6275);
nor NOR4 (N7563, N7548, N5803, N315, N2464);
and AND3 (N7564, N7553, N560, N4760);
or OR2 (N7565, N7560, N2593);
not NOT1 (N7566, N7547);
or OR2 (N7567, N7563, N2895);
xor XOR2 (N7568, N7566, N866);
xor XOR2 (N7569, N7559, N7093);
buf BUF1 (N7570, N7562);
nor NOR3 (N7571, N7569, N4754, N2228);
nand NAND4 (N7572, N7570, N2077, N5215, N4198);
or OR3 (N7573, N7565, N149, N4857);
or OR2 (N7574, N7568, N5981);
nand NAND3 (N7575, N7551, N1101, N5163);
or OR3 (N7576, N7573, N4527, N3272);
xor XOR2 (N7577, N7561, N7060);
buf BUF1 (N7578, N7577);
buf BUF1 (N7579, N7576);
nor NOR3 (N7580, N7564, N1500, N4067);
not NOT1 (N7581, N7558);
xor XOR2 (N7582, N7571, N3494);
nor NOR3 (N7583, N7579, N6704, N116);
not NOT1 (N7584, N7574);
nand NAND2 (N7585, N7550, N7359);
nor NOR3 (N7586, N7583, N5224, N4083);
not NOT1 (N7587, N7580);
xor XOR2 (N7588, N7567, N6760);
nor NOR2 (N7589, N7587, N3729);
buf BUF1 (N7590, N7584);
buf BUF1 (N7591, N7581);
buf BUF1 (N7592, N7572);
xor XOR2 (N7593, N7588, N4258);
xor XOR2 (N7594, N7591, N5674);
xor XOR2 (N7595, N7575, N5528);
xor XOR2 (N7596, N7589, N4591);
or OR2 (N7597, N7593, N394);
not NOT1 (N7598, N7596);
nor NOR4 (N7599, N7582, N1661, N7521, N2974);
nor NOR2 (N7600, N7595, N2224);
xor XOR2 (N7601, N7600, N6251);
and AND2 (N7602, N7586, N2238);
xor XOR2 (N7603, N7602, N6093);
xor XOR2 (N7604, N7578, N2195);
nor NOR4 (N7605, N7598, N692, N4535, N768);
nor NOR3 (N7606, N7594, N908, N4366);
nor NOR4 (N7607, N7585, N4308, N3766, N212);
and AND4 (N7608, N7604, N6174, N7008, N6987);
and AND3 (N7609, N7603, N6515, N327);
buf BUF1 (N7610, N7597);
nor NOR3 (N7611, N7610, N5371, N2746);
buf BUF1 (N7612, N7601);
buf BUF1 (N7613, N7608);
nand NAND2 (N7614, N7606, N966);
and AND4 (N7615, N7592, N6823, N4771, N2107);
buf BUF1 (N7616, N7612);
nor NOR3 (N7617, N7611, N2439, N5949);
and AND3 (N7618, N7614, N6357, N5306);
xor XOR2 (N7619, N7599, N3569);
nor NOR3 (N7620, N7609, N5810, N2478);
or OR2 (N7621, N7605, N4002);
nor NOR3 (N7622, N7619, N935, N2248);
not NOT1 (N7623, N7615);
xor XOR2 (N7624, N7616, N4833);
nand NAND4 (N7625, N7590, N4201, N4381, N5220);
or OR3 (N7626, N7622, N1781, N5301);
nand NAND3 (N7627, N7623, N7511, N4658);
nand NAND3 (N7628, N7607, N1226, N1539);
and AND3 (N7629, N7624, N2849, N2697);
xor XOR2 (N7630, N7625, N5713);
buf BUF1 (N7631, N7617);
buf BUF1 (N7632, N7628);
xor XOR2 (N7633, N7627, N2574);
xor XOR2 (N7634, N7633, N6161);
nand NAND2 (N7635, N7634, N2107);
nor NOR2 (N7636, N7626, N1878);
buf BUF1 (N7637, N7636);
nor NOR4 (N7638, N7637, N2131, N4469, N5888);
not NOT1 (N7639, N7635);
or OR2 (N7640, N7630, N3242);
buf BUF1 (N7641, N7629);
and AND2 (N7642, N7618, N5005);
and AND2 (N7643, N7638, N6178);
or OR4 (N7644, N7631, N6008, N1694, N4163);
or OR3 (N7645, N7640, N5968, N1090);
or OR3 (N7646, N7621, N3808, N6191);
or OR4 (N7647, N7645, N6882, N166, N2139);
xor XOR2 (N7648, N7646, N959);
nor NOR2 (N7649, N7613, N5464);
nor NOR3 (N7650, N7639, N6305, N2717);
and AND4 (N7651, N7620, N1302, N6544, N6908);
not NOT1 (N7652, N7647);
not NOT1 (N7653, N7644);
nor NOR2 (N7654, N7642, N6455);
buf BUF1 (N7655, N7632);
and AND2 (N7656, N7652, N7493);
or OR3 (N7657, N7654, N5315, N3516);
xor XOR2 (N7658, N7655, N4124);
xor XOR2 (N7659, N7657, N7173);
xor XOR2 (N7660, N7641, N109);
buf BUF1 (N7661, N7658);
xor XOR2 (N7662, N7653, N6027);
not NOT1 (N7663, N7656);
and AND2 (N7664, N7648, N7329);
nand NAND2 (N7665, N7663, N3850);
and AND4 (N7666, N7662, N6599, N2023, N6274);
not NOT1 (N7667, N7665);
nor NOR2 (N7668, N7664, N5269);
nand NAND4 (N7669, N7660, N4419, N7505, N343);
buf BUF1 (N7670, N7661);
buf BUF1 (N7671, N7643);
or OR4 (N7672, N7667, N5053, N6208, N5813);
nor NOR4 (N7673, N7651, N7127, N3509, N872);
nand NAND2 (N7674, N7650, N267);
or OR4 (N7675, N7674, N5515, N7639, N5065);
xor XOR2 (N7676, N7673, N5169);
xor XOR2 (N7677, N7669, N2818);
and AND3 (N7678, N7670, N1662, N3934);
and AND3 (N7679, N7678, N2319, N4308);
buf BUF1 (N7680, N7672);
buf BUF1 (N7681, N7649);
buf BUF1 (N7682, N7666);
nor NOR2 (N7683, N7682, N6816);
xor XOR2 (N7684, N7677, N2358);
nor NOR4 (N7685, N7679, N2525, N5165, N4967);
and AND2 (N7686, N7676, N6730);
or OR2 (N7687, N7686, N4624);
and AND2 (N7688, N7668, N5464);
xor XOR2 (N7689, N7688, N2288);
or OR4 (N7690, N7671, N2898, N7440, N3028);
buf BUF1 (N7691, N7684);
buf BUF1 (N7692, N7685);
not NOT1 (N7693, N7675);
buf BUF1 (N7694, N7687);
and AND3 (N7695, N7680, N3087, N5404);
nand NAND4 (N7696, N7683, N1450, N3573, N6101);
nor NOR4 (N7697, N7691, N1213, N5410, N7683);
or OR4 (N7698, N7695, N6804, N4224, N2997);
nand NAND3 (N7699, N7689, N3636, N7167);
nor NOR4 (N7700, N7692, N2933, N3111, N4663);
nand NAND4 (N7701, N7690, N6318, N6836, N174);
not NOT1 (N7702, N7681);
nand NAND2 (N7703, N7702, N3349);
nand NAND3 (N7704, N7703, N203, N6171);
not NOT1 (N7705, N7700);
nand NAND4 (N7706, N7693, N1767, N7577, N2661);
buf BUF1 (N7707, N7694);
not NOT1 (N7708, N7696);
buf BUF1 (N7709, N7697);
or OR2 (N7710, N7708, N2090);
or OR2 (N7711, N7698, N7354);
nand NAND2 (N7712, N7704, N6695);
nor NOR2 (N7713, N7701, N1827);
xor XOR2 (N7714, N7710, N5559);
buf BUF1 (N7715, N7659);
nand NAND3 (N7716, N7713, N4571, N5054);
not NOT1 (N7717, N7711);
nor NOR2 (N7718, N7709, N6929);
buf BUF1 (N7719, N7712);
nor NOR4 (N7720, N7705, N3550, N3342, N7281);
or OR3 (N7721, N7718, N5667, N4587);
nand NAND3 (N7722, N7715, N4334, N891);
or OR3 (N7723, N7720, N6967, N6003);
nor NOR2 (N7724, N7707, N7344);
and AND2 (N7725, N7723, N2891);
buf BUF1 (N7726, N7725);
and AND3 (N7727, N7724, N4603, N2044);
buf BUF1 (N7728, N7706);
nand NAND3 (N7729, N7727, N417, N1971);
nand NAND2 (N7730, N7719, N7006);
or OR2 (N7731, N7716, N4148);
xor XOR2 (N7732, N7726, N2728);
and AND2 (N7733, N7714, N81);
and AND3 (N7734, N7733, N7092, N4633);
not NOT1 (N7735, N7731);
or OR2 (N7736, N7735, N1955);
nand NAND4 (N7737, N7722, N5589, N623, N360);
nand NAND3 (N7738, N7736, N719, N5987);
nor NOR4 (N7739, N7737, N2199, N6202, N368);
nor NOR3 (N7740, N7730, N5618, N5188);
nand NAND2 (N7741, N7734, N3063);
xor XOR2 (N7742, N7741, N2250);
or OR2 (N7743, N7738, N3493);
nand NAND3 (N7744, N7742, N4617, N2626);
xor XOR2 (N7745, N7699, N5712);
not NOT1 (N7746, N7717);
or OR2 (N7747, N7732, N1168);
buf BUF1 (N7748, N7747);
not NOT1 (N7749, N7721);
nand NAND4 (N7750, N7748, N3292, N7087, N7719);
nand NAND3 (N7751, N7746, N7249, N6787);
nor NOR3 (N7752, N7749, N617, N7000);
or OR3 (N7753, N7744, N2988, N3789);
xor XOR2 (N7754, N7750, N544);
not NOT1 (N7755, N7743);
buf BUF1 (N7756, N7751);
nand NAND2 (N7757, N7739, N6756);
nor NOR3 (N7758, N7754, N4737, N4807);
or OR2 (N7759, N7745, N2897);
and AND2 (N7760, N7759, N949);
buf BUF1 (N7761, N7758);
or OR4 (N7762, N7761, N6205, N4389, N2878);
nor NOR4 (N7763, N7752, N4169, N5192, N5635);
and AND4 (N7764, N7728, N6947, N3513, N4433);
and AND4 (N7765, N7755, N6014, N4817, N4085);
nand NAND2 (N7766, N7765, N7074);
buf BUF1 (N7767, N7740);
nor NOR2 (N7768, N7753, N410);
nand NAND3 (N7769, N7764, N4305, N3324);
nor NOR2 (N7770, N7762, N2045);
not NOT1 (N7771, N7756);
buf BUF1 (N7772, N7769);
xor XOR2 (N7773, N7757, N2336);
not NOT1 (N7774, N7767);
buf BUF1 (N7775, N7773);
nor NOR2 (N7776, N7768, N6382);
nor NOR3 (N7777, N7763, N4525, N882);
xor XOR2 (N7778, N7766, N630);
nand NAND4 (N7779, N7772, N6901, N5306, N6541);
and AND3 (N7780, N7760, N731, N1421);
nor NOR3 (N7781, N7771, N6057, N3119);
buf BUF1 (N7782, N7776);
buf BUF1 (N7783, N7782);
nor NOR4 (N7784, N7770, N2787, N5113, N870);
nand NAND4 (N7785, N7780, N642, N3900, N2313);
not NOT1 (N7786, N7777);
and AND3 (N7787, N7779, N347, N3559);
not NOT1 (N7788, N7783);
nor NOR2 (N7789, N7778, N2821);
and AND4 (N7790, N7781, N7094, N3802, N1354);
nand NAND4 (N7791, N7789, N3051, N4159, N5895);
xor XOR2 (N7792, N7784, N3482);
buf BUF1 (N7793, N7790);
not NOT1 (N7794, N7785);
buf BUF1 (N7795, N7775);
not NOT1 (N7796, N7792);
and AND3 (N7797, N7794, N2984, N3959);
xor XOR2 (N7798, N7729, N4211);
xor XOR2 (N7799, N7788, N2690);
buf BUF1 (N7800, N7786);
or OR4 (N7801, N7798, N5415, N2683, N4366);
not NOT1 (N7802, N7787);
and AND3 (N7803, N7797, N4636, N7181);
nor NOR3 (N7804, N7799, N3683, N6344);
nor NOR4 (N7805, N7800, N2073, N3161, N7340);
buf BUF1 (N7806, N7791);
or OR4 (N7807, N7804, N423, N1326, N7685);
nand NAND2 (N7808, N7805, N2720);
not NOT1 (N7809, N7795);
nand NAND3 (N7810, N7801, N2505, N6722);
nor NOR3 (N7811, N7808, N5447, N1315);
or OR3 (N7812, N7774, N1814, N3466);
not NOT1 (N7813, N7793);
buf BUF1 (N7814, N7811);
nor NOR2 (N7815, N7810, N3352);
nor NOR4 (N7816, N7796, N146, N5527, N1247);
or OR3 (N7817, N7809, N3100, N6323);
nand NAND3 (N7818, N7802, N2460, N5058);
nand NAND4 (N7819, N7814, N861, N4515, N3482);
nor NOR4 (N7820, N7817, N22, N4411, N4229);
and AND2 (N7821, N7819, N7720);
buf BUF1 (N7822, N7807);
xor XOR2 (N7823, N7806, N4430);
or OR2 (N7824, N7812, N99);
buf BUF1 (N7825, N7824);
not NOT1 (N7826, N7825);
nor NOR4 (N7827, N7818, N714, N7314, N6492);
nand NAND3 (N7828, N7820, N1128, N5476);
or OR2 (N7829, N7821, N5773);
nand NAND4 (N7830, N7823, N1139, N1014, N6384);
nand NAND2 (N7831, N7803, N3225);
buf BUF1 (N7832, N7816);
nand NAND2 (N7833, N7826, N5801);
nand NAND3 (N7834, N7831, N1928, N717);
nor NOR4 (N7835, N7827, N5403, N7279, N5398);
not NOT1 (N7836, N7833);
nor NOR4 (N7837, N7830, N487, N4458, N3375);
xor XOR2 (N7838, N7822, N3176);
buf BUF1 (N7839, N7828);
or OR3 (N7840, N7813, N4618, N7628);
xor XOR2 (N7841, N7840, N3120);
nor NOR4 (N7842, N7839, N6552, N5037, N3171);
xor XOR2 (N7843, N7835, N6320);
not NOT1 (N7844, N7837);
not NOT1 (N7845, N7815);
nand NAND4 (N7846, N7834, N413, N6427, N7546);
and AND3 (N7847, N7841, N623, N5200);
xor XOR2 (N7848, N7846, N553);
nand NAND4 (N7849, N7842, N2828, N5031, N6847);
buf BUF1 (N7850, N7849);
nor NOR2 (N7851, N7843, N7427);
not NOT1 (N7852, N7845);
nor NOR4 (N7853, N7848, N125, N1957, N3388);
or OR2 (N7854, N7836, N4232);
nor NOR3 (N7855, N7850, N4111, N7631);
or OR3 (N7856, N7854, N4728, N3402);
not NOT1 (N7857, N7838);
nand NAND4 (N7858, N7844, N5846, N3139, N3977);
nor NOR2 (N7859, N7856, N1177);
nor NOR4 (N7860, N7847, N1259, N2587, N6854);
not NOT1 (N7861, N7853);
and AND2 (N7862, N7860, N3994);
xor XOR2 (N7863, N7851, N5182);
or OR2 (N7864, N7857, N805);
buf BUF1 (N7865, N7852);
xor XOR2 (N7866, N7862, N6122);
or OR2 (N7867, N7858, N437);
or OR3 (N7868, N7866, N1794, N7016);
xor XOR2 (N7869, N7864, N1153);
nand NAND3 (N7870, N7863, N7514, N412);
buf BUF1 (N7871, N7869);
nand NAND4 (N7872, N7871, N7548, N5770, N7547);
buf BUF1 (N7873, N7865);
xor XOR2 (N7874, N7829, N7278);
not NOT1 (N7875, N7861);
xor XOR2 (N7876, N7855, N6123);
nor NOR4 (N7877, N7868, N2803, N6818, N2792);
xor XOR2 (N7878, N7873, N3538);
or OR2 (N7879, N7875, N6985);
xor XOR2 (N7880, N7870, N3739);
or OR4 (N7881, N7877, N3557, N3775, N5338);
xor XOR2 (N7882, N7859, N6937);
xor XOR2 (N7883, N7874, N5568);
xor XOR2 (N7884, N7879, N378);
not NOT1 (N7885, N7882);
nor NOR3 (N7886, N7867, N4959, N4695);
not NOT1 (N7887, N7832);
nor NOR3 (N7888, N7883, N5231, N3096);
xor XOR2 (N7889, N7888, N7328);
or OR4 (N7890, N7876, N2068, N1914, N7729);
nor NOR3 (N7891, N7880, N7204, N5006);
and AND2 (N7892, N7884, N7418);
and AND4 (N7893, N7881, N7596, N5723, N5789);
not NOT1 (N7894, N7893);
not NOT1 (N7895, N7890);
not NOT1 (N7896, N7892);
or OR3 (N7897, N7889, N1867, N7063);
nor NOR3 (N7898, N7887, N6053, N7578);
xor XOR2 (N7899, N7897, N13);
nor NOR4 (N7900, N7886, N4348, N4871, N1629);
buf BUF1 (N7901, N7891);
buf BUF1 (N7902, N7901);
buf BUF1 (N7903, N7902);
and AND4 (N7904, N7898, N1293, N7192, N1457);
buf BUF1 (N7905, N7900);
nor NOR3 (N7906, N7872, N7445, N4142);
or OR3 (N7907, N7899, N2153, N2266);
not NOT1 (N7908, N7894);
not NOT1 (N7909, N7905);
nor NOR3 (N7910, N7908, N4149, N7005);
nand NAND3 (N7911, N7907, N1225, N4479);
xor XOR2 (N7912, N7896, N407);
xor XOR2 (N7913, N7878, N5394);
or OR3 (N7914, N7885, N6212, N1978);
not NOT1 (N7915, N7904);
xor XOR2 (N7916, N7915, N2654);
nand NAND4 (N7917, N7913, N4382, N63, N2175);
nor NOR3 (N7918, N7917, N1739, N2567);
xor XOR2 (N7919, N7912, N6152);
or OR2 (N7920, N7916, N1043);
xor XOR2 (N7921, N7914, N189);
and AND4 (N7922, N7918, N3019, N212, N3661);
and AND2 (N7923, N7922, N5948);
not NOT1 (N7924, N7910);
buf BUF1 (N7925, N7919);
nand NAND4 (N7926, N7909, N1390, N6510, N3494);
not NOT1 (N7927, N7923);
not NOT1 (N7928, N7906);
and AND3 (N7929, N7926, N5780, N2416);
or OR2 (N7930, N7924, N5381);
xor XOR2 (N7931, N7921, N1670);
xor XOR2 (N7932, N7925, N4634);
xor XOR2 (N7933, N7928, N4854);
and AND3 (N7934, N7931, N4769, N1266);
not NOT1 (N7935, N7929);
xor XOR2 (N7936, N7920, N6499);
nor NOR3 (N7937, N7930, N3967, N2928);
xor XOR2 (N7938, N7932, N2422);
nor NOR3 (N7939, N7938, N5241, N3204);
or OR3 (N7940, N7939, N3336, N2567);
nor NOR2 (N7941, N7940, N7841);
buf BUF1 (N7942, N7941);
xor XOR2 (N7943, N7937, N4993);
nor NOR4 (N7944, N7911, N4152, N635, N6453);
or OR3 (N7945, N7895, N6990, N1670);
xor XOR2 (N7946, N7903, N3697);
not NOT1 (N7947, N7944);
and AND2 (N7948, N7943, N7161);
nand NAND2 (N7949, N7934, N3702);
or OR3 (N7950, N7936, N1983, N199);
or OR4 (N7951, N7946, N3953, N6515, N7450);
xor XOR2 (N7952, N7949, N2317);
and AND3 (N7953, N7948, N7331, N4949);
or OR2 (N7954, N7933, N1889);
and AND3 (N7955, N7947, N2952, N223);
not NOT1 (N7956, N7935);
or OR4 (N7957, N7950, N153, N318, N1359);
and AND4 (N7958, N7954, N6950, N5237, N4834);
nor NOR2 (N7959, N7945, N4878);
not NOT1 (N7960, N7956);
nand NAND3 (N7961, N7960, N3049, N7318);
nand NAND3 (N7962, N7942, N7612, N2540);
buf BUF1 (N7963, N7962);
nor NOR3 (N7964, N7953, N7846, N1221);
nor NOR2 (N7965, N7961, N4876);
buf BUF1 (N7966, N7965);
nand NAND2 (N7967, N7966, N5795);
and AND4 (N7968, N7959, N1717, N1261, N3557);
nand NAND2 (N7969, N7964, N4066);
nand NAND3 (N7970, N7955, N1354, N4105);
nand NAND3 (N7971, N7970, N3048, N3415);
xor XOR2 (N7972, N7952, N1946);
not NOT1 (N7973, N7971);
xor XOR2 (N7974, N7968, N4624);
not NOT1 (N7975, N7963);
xor XOR2 (N7976, N7975, N4806);
or OR3 (N7977, N7974, N6203, N223);
or OR3 (N7978, N7967, N6417, N6395);
xor XOR2 (N7979, N7957, N3657);
or OR4 (N7980, N7958, N6906, N519, N2676);
buf BUF1 (N7981, N7973);
xor XOR2 (N7982, N7972, N5021);
nor NOR2 (N7983, N7969, N7057);
buf BUF1 (N7984, N7979);
xor XOR2 (N7985, N7977, N2673);
buf BUF1 (N7986, N7983);
and AND2 (N7987, N7978, N4131);
buf BUF1 (N7988, N7986);
nand NAND3 (N7989, N7981, N6662, N3373);
xor XOR2 (N7990, N7951, N6931);
buf BUF1 (N7991, N7990);
or OR2 (N7992, N7980, N1345);
xor XOR2 (N7993, N7976, N3542);
buf BUF1 (N7994, N7987);
and AND4 (N7995, N7994, N4181, N6458, N4476);
or OR3 (N7996, N7989, N4026, N4774);
and AND2 (N7997, N7984, N4259);
nand NAND3 (N7998, N7988, N1482, N4776);
buf BUF1 (N7999, N7995);
nand NAND2 (N8000, N7991, N5066);
and AND2 (N8001, N7992, N1034);
buf BUF1 (N8002, N7927);
nand NAND2 (N8003, N7999, N5804);
not NOT1 (N8004, N8002);
and AND3 (N8005, N7997, N4531, N2594);
nand NAND4 (N8006, N8004, N3052, N1819, N5843);
or OR4 (N8007, N8003, N6132, N7427, N5045);
nand NAND4 (N8008, N8007, N3873, N7333, N2990);
buf BUF1 (N8009, N7993);
buf BUF1 (N8010, N7998);
not NOT1 (N8011, N8009);
nor NOR2 (N8012, N8006, N7876);
nor NOR2 (N8013, N7982, N5231);
nor NOR2 (N8014, N8008, N3640);
xor XOR2 (N8015, N8005, N6995);
nor NOR4 (N8016, N7985, N6289, N3668, N90);
nor NOR2 (N8017, N8001, N1216);
buf BUF1 (N8018, N8015);
nor NOR3 (N8019, N8017, N5110, N4192);
and AND4 (N8020, N8013, N4188, N4230, N2309);
or OR3 (N8021, N8012, N5495, N3344);
nand NAND2 (N8022, N8010, N2050);
or OR3 (N8023, N8020, N5283, N298);
nand NAND4 (N8024, N8011, N2987, N5217, N1328);
and AND2 (N8025, N8016, N7475);
or OR2 (N8026, N8019, N276);
xor XOR2 (N8027, N8026, N3512);
nor NOR2 (N8028, N8025, N632);
not NOT1 (N8029, N8000);
buf BUF1 (N8030, N8018);
and AND3 (N8031, N8023, N5684, N3949);
nand NAND2 (N8032, N8030, N2275);
nor NOR3 (N8033, N7996, N582, N3045);
buf BUF1 (N8034, N8028);
xor XOR2 (N8035, N8031, N4559);
or OR4 (N8036, N8014, N7079, N2595, N632);
not NOT1 (N8037, N8032);
nand NAND2 (N8038, N8033, N7980);
nand NAND4 (N8039, N8037, N3205, N2779, N1554);
xor XOR2 (N8040, N8035, N1859);
nand NAND4 (N8041, N8040, N5039, N5283, N5825);
or OR3 (N8042, N8041, N4525, N4473);
not NOT1 (N8043, N8034);
buf BUF1 (N8044, N8039);
not NOT1 (N8045, N8029);
xor XOR2 (N8046, N8022, N3977);
and AND4 (N8047, N8043, N5444, N7304, N667);
nor NOR4 (N8048, N8024, N7070, N8034, N5508);
and AND4 (N8049, N8038, N4956, N2842, N5209);
not NOT1 (N8050, N8045);
xor XOR2 (N8051, N8036, N4102);
nand NAND2 (N8052, N8021, N6742);
or OR3 (N8053, N8044, N5200, N1850);
or OR4 (N8054, N8042, N3261, N6218, N7395);
nand NAND4 (N8055, N8051, N1262, N7530, N3847);
and AND3 (N8056, N8046, N3247, N7274);
buf BUF1 (N8057, N8053);
and AND3 (N8058, N8050, N8007, N4976);
buf BUF1 (N8059, N8056);
nor NOR4 (N8060, N8027, N2374, N5286, N3551);
not NOT1 (N8061, N8059);
xor XOR2 (N8062, N8055, N6044);
xor XOR2 (N8063, N8057, N907);
or OR4 (N8064, N8049, N3808, N6775, N1534);
and AND3 (N8065, N8054, N4047, N211);
buf BUF1 (N8066, N8064);
xor XOR2 (N8067, N8061, N1992);
nor NOR4 (N8068, N8066, N4108, N7547, N7498);
and AND3 (N8069, N8052, N7174, N6275);
or OR4 (N8070, N8047, N6271, N3151, N6478);
and AND2 (N8071, N8069, N6089);
xor XOR2 (N8072, N8048, N1864);
nor NOR2 (N8073, N8062, N4167);
and AND3 (N8074, N8060, N4645, N1678);
buf BUF1 (N8075, N8073);
buf BUF1 (N8076, N8058);
nor NOR2 (N8077, N8072, N540);
xor XOR2 (N8078, N8067, N4463);
nand NAND2 (N8079, N8074, N6836);
not NOT1 (N8080, N8076);
or OR4 (N8081, N8071, N6166, N7255, N4335);
xor XOR2 (N8082, N8068, N5087);
xor XOR2 (N8083, N8063, N1406);
xor XOR2 (N8084, N8075, N18);
or OR3 (N8085, N8080, N933, N2009);
nor NOR2 (N8086, N8083, N133);
nand NAND2 (N8087, N8086, N2837);
buf BUF1 (N8088, N8079);
and AND4 (N8089, N8088, N1509, N1120, N4917);
not NOT1 (N8090, N8087);
buf BUF1 (N8091, N8078);
or OR3 (N8092, N8081, N3838, N3217);
xor XOR2 (N8093, N8092, N4717);
and AND3 (N8094, N8065, N596, N4822);
buf BUF1 (N8095, N8089);
nand NAND2 (N8096, N8090, N4586);
buf BUF1 (N8097, N8093);
xor XOR2 (N8098, N8095, N2015);
or OR3 (N8099, N8091, N2685, N2998);
xor XOR2 (N8100, N8084, N5123);
and AND3 (N8101, N8085, N4600, N6935);
and AND3 (N8102, N8101, N6288, N5065);
or OR3 (N8103, N8077, N2009, N6317);
or OR2 (N8104, N8082, N4319);
buf BUF1 (N8105, N8094);
and AND2 (N8106, N8098, N2232);
buf BUF1 (N8107, N8096);
xor XOR2 (N8108, N8104, N5784);
or OR4 (N8109, N8100, N174, N6996, N796);
xor XOR2 (N8110, N8107, N3249);
and AND4 (N8111, N8103, N7363, N4948, N5940);
xor XOR2 (N8112, N8108, N4203);
not NOT1 (N8113, N8070);
buf BUF1 (N8114, N8109);
not NOT1 (N8115, N8105);
not NOT1 (N8116, N8106);
xor XOR2 (N8117, N8097, N987);
or OR4 (N8118, N8114, N662, N3776, N7252);
and AND2 (N8119, N8102, N455);
not NOT1 (N8120, N8116);
xor XOR2 (N8121, N8120, N2920);
buf BUF1 (N8122, N8119);
buf BUF1 (N8123, N8122);
or OR4 (N8124, N8118, N7746, N535, N7847);
or OR4 (N8125, N8111, N3009, N5761, N7670);
buf BUF1 (N8126, N8099);
nor NOR4 (N8127, N8123, N352, N7721, N6589);
or OR3 (N8128, N8115, N3551, N6094);
buf BUF1 (N8129, N8112);
and AND3 (N8130, N8113, N5396, N1227);
nor NOR3 (N8131, N8124, N6101, N746);
buf BUF1 (N8132, N8121);
xor XOR2 (N8133, N8117, N2595);
nor NOR4 (N8134, N8128, N2767, N2476, N7480);
or OR4 (N8135, N8127, N2563, N7801, N6463);
nand NAND4 (N8136, N8132, N7324, N2375, N901);
nor NOR3 (N8137, N8126, N6505, N7526);
not NOT1 (N8138, N8129);
or OR3 (N8139, N8138, N5595, N2888);
and AND2 (N8140, N8135, N5917);
nor NOR4 (N8141, N8134, N2142, N8043, N5363);
or OR2 (N8142, N8110, N3603);
or OR2 (N8143, N8137, N4247);
xor XOR2 (N8144, N8139, N6636);
and AND3 (N8145, N8130, N5262, N1528);
buf BUF1 (N8146, N8131);
xor XOR2 (N8147, N8136, N2308);
not NOT1 (N8148, N8143);
nor NOR3 (N8149, N8144, N5085, N6070);
or OR3 (N8150, N8148, N4153, N1692);
nor NOR3 (N8151, N8146, N1845, N1487);
nor NOR3 (N8152, N8149, N4221, N3219);
buf BUF1 (N8153, N8152);
and AND3 (N8154, N8153, N4855, N970);
nor NOR4 (N8155, N8154, N7098, N750, N2438);
xor XOR2 (N8156, N8140, N4496);
buf BUF1 (N8157, N8142);
buf BUF1 (N8158, N8145);
or OR4 (N8159, N8133, N4083, N1362, N347);
or OR4 (N8160, N8155, N6686, N766, N125);
or OR2 (N8161, N8151, N484);
nand NAND2 (N8162, N8157, N2854);
not NOT1 (N8163, N8162);
xor XOR2 (N8164, N8161, N2567);
or OR4 (N8165, N8150, N864, N1304, N2419);
xor XOR2 (N8166, N8141, N2806);
nor NOR4 (N8167, N8125, N3601, N4876, N920);
not NOT1 (N8168, N8159);
and AND4 (N8169, N8158, N4162, N4104, N4097);
nor NOR3 (N8170, N8160, N4627, N7614);
and AND2 (N8171, N8166, N260);
not NOT1 (N8172, N8168);
not NOT1 (N8173, N8170);
or OR3 (N8174, N8167, N4903, N1019);
nand NAND2 (N8175, N8163, N7326);
not NOT1 (N8176, N8165);
nor NOR4 (N8177, N8156, N909, N3551, N3468);
xor XOR2 (N8178, N8147, N3755);
xor XOR2 (N8179, N8175, N6345);
or OR3 (N8180, N8164, N8153, N5156);
nand NAND3 (N8181, N8174, N3573, N2340);
nand NAND4 (N8182, N8176, N4550, N3288, N6057);
xor XOR2 (N8183, N8179, N7748);
and AND3 (N8184, N8178, N2023, N1821);
nor NOR4 (N8185, N8172, N2501, N3923, N3038);
xor XOR2 (N8186, N8173, N4295);
xor XOR2 (N8187, N8183, N8169);
buf BUF1 (N8188, N6503);
xor XOR2 (N8189, N8188, N1855);
buf BUF1 (N8190, N8177);
not NOT1 (N8191, N8189);
and AND4 (N8192, N8171, N2931, N6755, N112);
nand NAND3 (N8193, N8187, N7973, N7027);
nor NOR2 (N8194, N8191, N7739);
or OR4 (N8195, N8194, N4159, N560, N7009);
nor NOR2 (N8196, N8182, N2362);
nand NAND2 (N8197, N8196, N2574);
nand NAND4 (N8198, N8193, N1265, N6922, N7236);
and AND3 (N8199, N8186, N6617, N4409);
or OR2 (N8200, N8184, N6355);
or OR4 (N8201, N8192, N8050, N7437, N3247);
buf BUF1 (N8202, N8180);
not NOT1 (N8203, N8198);
nor NOR4 (N8204, N8190, N7454, N2758, N6106);
and AND2 (N8205, N8199, N2763);
nand NAND2 (N8206, N8203, N7265);
xor XOR2 (N8207, N8197, N3724);
nor NOR3 (N8208, N8207, N6577, N3075);
or OR3 (N8209, N8204, N2932, N2031);
not NOT1 (N8210, N8209);
not NOT1 (N8211, N8210);
or OR2 (N8212, N8206, N5260);
xor XOR2 (N8213, N8181, N6962);
and AND4 (N8214, N8201, N5146, N2943, N1789);
nand NAND2 (N8215, N8214, N1697);
and AND2 (N8216, N8195, N6069);
not NOT1 (N8217, N8205);
or OR4 (N8218, N8216, N7103, N2972, N3861);
nor NOR4 (N8219, N8208, N305, N7725, N5661);
nand NAND4 (N8220, N8217, N3606, N1176, N3216);
or OR4 (N8221, N8185, N6582, N4456, N3429);
and AND3 (N8222, N8221, N4843, N4116);
xor XOR2 (N8223, N8218, N5739);
xor XOR2 (N8224, N8219, N3677);
and AND4 (N8225, N8212, N3678, N6569, N1551);
not NOT1 (N8226, N8213);
nor NOR4 (N8227, N8211, N466, N4389, N519);
or OR3 (N8228, N8223, N6816, N2405);
or OR3 (N8229, N8228, N214, N4564);
nor NOR4 (N8230, N8222, N5033, N2877, N4032);
nor NOR2 (N8231, N8202, N1851);
not NOT1 (N8232, N8230);
buf BUF1 (N8233, N8227);
not NOT1 (N8234, N8200);
and AND4 (N8235, N8232, N5706, N1173, N3044);
buf BUF1 (N8236, N8225);
nand NAND4 (N8237, N8234, N1666, N1736, N3110);
not NOT1 (N8238, N8233);
buf BUF1 (N8239, N8224);
nor NOR2 (N8240, N8235, N1088);
not NOT1 (N8241, N8220);
buf BUF1 (N8242, N8241);
nand NAND4 (N8243, N8240, N4581, N7754, N552);
or OR2 (N8244, N8231, N1061);
not NOT1 (N8245, N8242);
nand NAND2 (N8246, N8245, N4746);
xor XOR2 (N8247, N8226, N599);
buf BUF1 (N8248, N8229);
nor NOR3 (N8249, N8247, N5392, N5192);
or OR4 (N8250, N8237, N7714, N7682, N3611);
or OR2 (N8251, N8238, N5024);
nor NOR3 (N8252, N8243, N1504, N1624);
buf BUF1 (N8253, N8246);
and AND2 (N8254, N8253, N4432);
nor NOR4 (N8255, N8236, N5278, N1123, N741);
or OR3 (N8256, N8215, N3824, N440);
buf BUF1 (N8257, N8250);
nand NAND4 (N8258, N8257, N7542, N6221, N7872);
nand NAND4 (N8259, N8239, N7271, N3410, N5789);
nand NAND3 (N8260, N8256, N6360, N7785);
nor NOR4 (N8261, N8251, N4676, N5847, N4676);
or OR2 (N8262, N8244, N5460);
nand NAND4 (N8263, N8262, N1600, N2011, N3799);
xor XOR2 (N8264, N8263, N5862);
nand NAND2 (N8265, N8249, N7804);
buf BUF1 (N8266, N8259);
or OR2 (N8267, N8264, N4554);
not NOT1 (N8268, N8258);
xor XOR2 (N8269, N8254, N998);
buf BUF1 (N8270, N8261);
or OR2 (N8271, N8268, N6068);
nand NAND4 (N8272, N8255, N6143, N5919, N1214);
not NOT1 (N8273, N8269);
or OR3 (N8274, N8248, N4590, N2709);
nor NOR3 (N8275, N8270, N2017, N8049);
nand NAND2 (N8276, N8260, N708);
not NOT1 (N8277, N8252);
or OR2 (N8278, N8266, N5029);
or OR4 (N8279, N8265, N2359, N7745, N7162);
nand NAND4 (N8280, N8277, N595, N1681, N465);
and AND3 (N8281, N8267, N4227, N5709);
nor NOR2 (N8282, N8275, N3136);
and AND4 (N8283, N8272, N4667, N4343, N5617);
buf BUF1 (N8284, N8282);
nand NAND3 (N8285, N8273, N5572, N82);
xor XOR2 (N8286, N8280, N1694);
and AND2 (N8287, N8274, N8230);
not NOT1 (N8288, N8286);
or OR3 (N8289, N8281, N6658, N3871);
nor NOR3 (N8290, N8284, N5844, N7794);
not NOT1 (N8291, N8279);
nor NOR4 (N8292, N8289, N6422, N6615, N5831);
xor XOR2 (N8293, N8278, N8163);
buf BUF1 (N8294, N8291);
xor XOR2 (N8295, N8293, N165);
not NOT1 (N8296, N8285);
or OR3 (N8297, N8283, N1499, N7577);
not NOT1 (N8298, N8288);
nand NAND4 (N8299, N8271, N6564, N6235, N1550);
and AND3 (N8300, N8294, N8022, N3125);
or OR3 (N8301, N8276, N190, N7036);
buf BUF1 (N8302, N8301);
nand NAND4 (N8303, N8297, N7445, N6579, N6403);
xor XOR2 (N8304, N8298, N6173);
xor XOR2 (N8305, N8302, N4510);
buf BUF1 (N8306, N8287);
nand NAND4 (N8307, N8295, N541, N5015, N7739);
not NOT1 (N8308, N8296);
xor XOR2 (N8309, N8290, N466);
xor XOR2 (N8310, N8305, N5495);
or OR2 (N8311, N8307, N7785);
and AND3 (N8312, N8303, N431, N3889);
nor NOR3 (N8313, N8308, N26, N5845);
not NOT1 (N8314, N8300);
and AND2 (N8315, N8311, N1118);
or OR2 (N8316, N8314, N5239);
and AND3 (N8317, N8312, N5723, N2630);
nand NAND4 (N8318, N8304, N6483, N1932, N1364);
or OR3 (N8319, N8310, N395, N3783);
nor NOR3 (N8320, N8316, N3901, N593);
not NOT1 (N8321, N8317);
not NOT1 (N8322, N8319);
and AND3 (N8323, N8306, N3780, N2543);
nand NAND3 (N8324, N8320, N5693, N5334);
nor NOR2 (N8325, N8315, N3041);
and AND3 (N8326, N8321, N4288, N1423);
or OR4 (N8327, N8313, N3334, N7294, N5562);
buf BUF1 (N8328, N8322);
or OR2 (N8329, N8309, N3283);
nand NAND3 (N8330, N8327, N47, N6512);
buf BUF1 (N8331, N8318);
nand NAND4 (N8332, N8325, N825, N934, N1586);
and AND2 (N8333, N8323, N853);
and AND4 (N8334, N8329, N3449, N3411, N1035);
xor XOR2 (N8335, N8331, N4666);
nand NAND3 (N8336, N8328, N8159, N468);
xor XOR2 (N8337, N8299, N4831);
or OR2 (N8338, N8330, N5956);
buf BUF1 (N8339, N8326);
xor XOR2 (N8340, N8324, N6133);
xor XOR2 (N8341, N8338, N1104);
nand NAND4 (N8342, N8340, N1609, N4232, N4293);
nor NOR3 (N8343, N8341, N2561, N11);
not NOT1 (N8344, N8333);
buf BUF1 (N8345, N8337);
and AND3 (N8346, N8343, N257, N2027);
or OR4 (N8347, N8345, N6024, N4796, N4561);
and AND4 (N8348, N8292, N5897, N5289, N2060);
buf BUF1 (N8349, N8339);
nand NAND4 (N8350, N8334, N7173, N3130, N3422);
nand NAND2 (N8351, N8350, N4212);
and AND2 (N8352, N8336, N1089);
nor NOR3 (N8353, N8346, N3768, N4380);
buf BUF1 (N8354, N8332);
nand NAND4 (N8355, N8351, N7257, N171, N6722);
nand NAND4 (N8356, N8353, N2314, N709, N5137);
buf BUF1 (N8357, N8356);
or OR2 (N8358, N8349, N8009);
buf BUF1 (N8359, N8335);
xor XOR2 (N8360, N8342, N4459);
nand NAND4 (N8361, N8359, N2326, N2460, N7639);
and AND2 (N8362, N8361, N6786);
nand NAND4 (N8363, N8354, N2088, N2011, N144);
buf BUF1 (N8364, N8363);
not NOT1 (N8365, N8357);
buf BUF1 (N8366, N8352);
xor XOR2 (N8367, N8348, N1973);
xor XOR2 (N8368, N8347, N4461);
nor NOR3 (N8369, N8344, N6377, N5575);
or OR2 (N8370, N8362, N156);
not NOT1 (N8371, N8370);
nor NOR3 (N8372, N8360, N7943, N2324);
nor NOR3 (N8373, N8366, N638, N1300);
nand NAND4 (N8374, N8369, N2764, N5348, N3033);
nor NOR3 (N8375, N8365, N1200, N1925);
nor NOR2 (N8376, N8358, N1836);
and AND2 (N8377, N8371, N4535);
nand NAND4 (N8378, N8377, N1022, N4261, N676);
xor XOR2 (N8379, N8373, N8205);
buf BUF1 (N8380, N8379);
not NOT1 (N8381, N8375);
nor NOR2 (N8382, N8374, N3339);
nor NOR3 (N8383, N8367, N8196, N5087);
nand NAND3 (N8384, N8383, N6932, N5729);
not NOT1 (N8385, N8384);
xor XOR2 (N8386, N8368, N3130);
or OR4 (N8387, N8385, N1143, N1564, N8205);
buf BUF1 (N8388, N8387);
or OR3 (N8389, N8388, N814, N2149);
buf BUF1 (N8390, N8382);
not NOT1 (N8391, N8372);
nand NAND3 (N8392, N8364, N6319, N4641);
or OR3 (N8393, N8376, N7081, N7380);
buf BUF1 (N8394, N8380);
and AND3 (N8395, N8355, N2743, N3793);
and AND3 (N8396, N8393, N4036, N7571);
xor XOR2 (N8397, N8390, N8317);
nand NAND2 (N8398, N8386, N4337);
nand NAND2 (N8399, N8391, N7421);
nand NAND4 (N8400, N8397, N6056, N273, N5538);
or OR4 (N8401, N8378, N8053, N4602, N3051);
or OR3 (N8402, N8381, N5949, N5627);
nand NAND3 (N8403, N8398, N4909, N2797);
not NOT1 (N8404, N8392);
and AND3 (N8405, N8394, N1575, N6942);
buf BUF1 (N8406, N8402);
and AND4 (N8407, N8403, N7561, N1168, N6763);
and AND2 (N8408, N8389, N4184);
xor XOR2 (N8409, N8401, N7435);
xor XOR2 (N8410, N8408, N533);
xor XOR2 (N8411, N8395, N1131);
not NOT1 (N8412, N8409);
xor XOR2 (N8413, N8407, N290);
nand NAND4 (N8414, N8399, N3103, N5310, N1700);
xor XOR2 (N8415, N8406, N612);
and AND2 (N8416, N8412, N4651);
buf BUF1 (N8417, N8416);
not NOT1 (N8418, N8417);
nand NAND2 (N8419, N8404, N7955);
not NOT1 (N8420, N8415);
and AND2 (N8421, N8410, N5295);
or OR4 (N8422, N8413, N7312, N7768, N6700);
xor XOR2 (N8423, N8396, N339);
buf BUF1 (N8424, N8421);
buf BUF1 (N8425, N8424);
nor NOR2 (N8426, N8423, N132);
not NOT1 (N8427, N8422);
nor NOR2 (N8428, N8411, N8205);
or OR2 (N8429, N8419, N3561);
nand NAND4 (N8430, N8429, N3106, N6832, N3728);
or OR2 (N8431, N8418, N2710);
not NOT1 (N8432, N8430);
not NOT1 (N8433, N8425);
nand NAND4 (N8434, N8426, N7096, N6224, N7331);
nand NAND4 (N8435, N8431, N5825, N6911, N1374);
or OR2 (N8436, N8427, N5606);
nand NAND2 (N8437, N8400, N2343);
buf BUF1 (N8438, N8437);
buf BUF1 (N8439, N8433);
nand NAND4 (N8440, N8420, N6580, N1271, N2386);
and AND4 (N8441, N8435, N254, N5550, N1011);
nand NAND3 (N8442, N8441, N1063, N6232);
buf BUF1 (N8443, N8434);
and AND4 (N8444, N8405, N3117, N7829, N8167);
buf BUF1 (N8445, N8432);
nor NOR2 (N8446, N8443, N1849);
or OR2 (N8447, N8444, N4853);
and AND4 (N8448, N8442, N5319, N6226, N3859);
or OR3 (N8449, N8446, N2059, N4264);
buf BUF1 (N8450, N8449);
nand NAND4 (N8451, N8448, N7091, N6351, N3538);
nand NAND3 (N8452, N8436, N640, N3087);
and AND3 (N8453, N8439, N3020, N712);
not NOT1 (N8454, N8450);
not NOT1 (N8455, N8438);
and AND3 (N8456, N8445, N1799, N2313);
nand NAND2 (N8457, N8454, N2176);
not NOT1 (N8458, N8451);
nand NAND2 (N8459, N8440, N495);
buf BUF1 (N8460, N8447);
and AND4 (N8461, N8457, N2948, N3719, N8373);
or OR3 (N8462, N8414, N1797, N1731);
buf BUF1 (N8463, N8428);
nand NAND2 (N8464, N8452, N7592);
not NOT1 (N8465, N8458);
not NOT1 (N8466, N8455);
buf BUF1 (N8467, N8463);
and AND3 (N8468, N8453, N524, N7816);
nor NOR2 (N8469, N8468, N2432);
not NOT1 (N8470, N8464);
nand NAND2 (N8471, N8462, N7134);
or OR4 (N8472, N8471, N6253, N2627, N1944);
and AND2 (N8473, N8472, N321);
and AND3 (N8474, N8466, N3068, N1459);
nand NAND2 (N8475, N8474, N1502);
nand NAND2 (N8476, N8460, N8324);
or OR2 (N8477, N8465, N2139);
xor XOR2 (N8478, N8476, N7326);
xor XOR2 (N8479, N8475, N5277);
buf BUF1 (N8480, N8461);
not NOT1 (N8481, N8480);
buf BUF1 (N8482, N8477);
xor XOR2 (N8483, N8459, N5467);
nand NAND2 (N8484, N8467, N632);
nor NOR4 (N8485, N8484, N5464, N1084, N3649);
not NOT1 (N8486, N8456);
nand NAND2 (N8487, N8470, N3171);
buf BUF1 (N8488, N8478);
nand NAND3 (N8489, N8485, N6268, N5000);
or OR4 (N8490, N8488, N6113, N1073, N7444);
nand NAND4 (N8491, N8479, N7293, N1555, N3209);
nand NAND3 (N8492, N8483, N8132, N2895);
and AND3 (N8493, N8491, N7351, N7155);
nor NOR4 (N8494, N8487, N4309, N8032, N2260);
nor NOR2 (N8495, N8482, N2436);
not NOT1 (N8496, N8473);
buf BUF1 (N8497, N8492);
nand NAND3 (N8498, N8494, N5314, N6204);
nor NOR2 (N8499, N8495, N1145);
xor XOR2 (N8500, N8498, N4405);
not NOT1 (N8501, N8489);
nand NAND3 (N8502, N8486, N1892, N3968);
nor NOR3 (N8503, N8501, N4530, N2862);
nand NAND4 (N8504, N8502, N1290, N721, N6429);
and AND4 (N8505, N8481, N4483, N4204, N4092);
or OR3 (N8506, N8497, N5361, N8165);
nor NOR2 (N8507, N8504, N7154);
xor XOR2 (N8508, N8503, N4367);
or OR2 (N8509, N8490, N996);
or OR4 (N8510, N8496, N4027, N672, N5767);
buf BUF1 (N8511, N8499);
or OR3 (N8512, N8505, N1072, N3680);
nand NAND4 (N8513, N8493, N2313, N3835, N3975);
or OR4 (N8514, N8506, N1209, N3653, N7109);
and AND3 (N8515, N8514, N3308, N5457);
xor XOR2 (N8516, N8513, N7966);
nand NAND4 (N8517, N8509, N6920, N2426, N1132);
nand NAND3 (N8518, N8511, N6554, N1208);
and AND4 (N8519, N8508, N1847, N6834, N7801);
and AND3 (N8520, N8516, N1502, N2005);
or OR2 (N8521, N8507, N8160);
nand NAND4 (N8522, N8521, N1202, N49, N6215);
nor NOR2 (N8523, N8519, N1603);
nor NOR4 (N8524, N8520, N3129, N3210, N4077);
nor NOR2 (N8525, N8469, N2758);
and AND4 (N8526, N8512, N6193, N5749, N8018);
nand NAND3 (N8527, N8525, N6693, N2002);
and AND2 (N8528, N8510, N8461);
buf BUF1 (N8529, N8500);
nor NOR2 (N8530, N8526, N907);
not NOT1 (N8531, N8527);
nor NOR2 (N8532, N8524, N2630);
nor NOR2 (N8533, N8518, N1472);
or OR4 (N8534, N8530, N6301, N2163, N1344);
nand NAND2 (N8535, N8517, N814);
nand NAND3 (N8536, N8523, N241, N8308);
not NOT1 (N8537, N8536);
buf BUF1 (N8538, N8515);
or OR4 (N8539, N8522, N2771, N3925, N5505);
or OR2 (N8540, N8534, N3474);
xor XOR2 (N8541, N8538, N2987);
and AND3 (N8542, N8528, N7738, N1903);
buf BUF1 (N8543, N8542);
buf BUF1 (N8544, N8543);
nand NAND3 (N8545, N8541, N3868, N4343);
xor XOR2 (N8546, N8539, N1977);
xor XOR2 (N8547, N8531, N356);
buf BUF1 (N8548, N8547);
buf BUF1 (N8549, N8546);
nor NOR4 (N8550, N8540, N642, N3864, N1395);
nor NOR2 (N8551, N8529, N1597);
or OR4 (N8552, N8548, N3666, N3837, N3989);
xor XOR2 (N8553, N8550, N7081);
nand NAND4 (N8554, N8545, N782, N538, N7242);
buf BUF1 (N8555, N8533);
and AND2 (N8556, N8544, N7977);
not NOT1 (N8557, N8551);
or OR2 (N8558, N8552, N1856);
not NOT1 (N8559, N8554);
or OR3 (N8560, N8556, N3027, N3525);
nand NAND4 (N8561, N8537, N622, N6218, N3918);
or OR2 (N8562, N8559, N6818);
or OR2 (N8563, N8549, N6857);
not NOT1 (N8564, N8535);
nor NOR3 (N8565, N8564, N48, N76);
or OR3 (N8566, N8565, N5967, N2862);
xor XOR2 (N8567, N8563, N8085);
and AND2 (N8568, N8532, N6704);
xor XOR2 (N8569, N8560, N6961);
nor NOR4 (N8570, N8558, N1084, N4495, N8369);
nand NAND2 (N8571, N8562, N5432);
not NOT1 (N8572, N8553);
xor XOR2 (N8573, N8567, N5911);
or OR3 (N8574, N8573, N6649, N4086);
xor XOR2 (N8575, N8574, N8524);
buf BUF1 (N8576, N8570);
nand NAND2 (N8577, N8569, N7886);
not NOT1 (N8578, N8555);
nor NOR3 (N8579, N8575, N1164, N1290);
or OR4 (N8580, N8579, N143, N1408, N822);
nor NOR2 (N8581, N8578, N2537);
buf BUF1 (N8582, N8557);
or OR3 (N8583, N8568, N6658, N7807);
not NOT1 (N8584, N8571);
nand NAND2 (N8585, N8582, N2748);
xor XOR2 (N8586, N8581, N7856);
xor XOR2 (N8587, N8576, N4860);
xor XOR2 (N8588, N8566, N7745);
and AND2 (N8589, N8585, N4199);
or OR2 (N8590, N8588, N6939);
or OR2 (N8591, N8580, N4430);
or OR3 (N8592, N8586, N1261, N2336);
and AND3 (N8593, N8589, N4323, N2737);
not NOT1 (N8594, N8577);
xor XOR2 (N8595, N8592, N4952);
buf BUF1 (N8596, N8572);
buf BUF1 (N8597, N8583);
nor NOR4 (N8598, N8561, N7355, N6947, N7553);
or OR2 (N8599, N8594, N4374);
xor XOR2 (N8600, N8591, N5537);
xor XOR2 (N8601, N8587, N6343);
buf BUF1 (N8602, N8590);
buf BUF1 (N8603, N8596);
nand NAND4 (N8604, N8598, N7249, N7963, N1838);
buf BUF1 (N8605, N8600);
buf BUF1 (N8606, N8604);
xor XOR2 (N8607, N8595, N3171);
nor NOR3 (N8608, N8593, N7058, N2944);
buf BUF1 (N8609, N8599);
nor NOR2 (N8610, N8609, N1201);
not NOT1 (N8611, N8603);
not NOT1 (N8612, N8610);
xor XOR2 (N8613, N8602, N4547);
buf BUF1 (N8614, N8584);
buf BUF1 (N8615, N8597);
nand NAND2 (N8616, N8608, N71);
buf BUF1 (N8617, N8614);
buf BUF1 (N8618, N8617);
and AND2 (N8619, N8605, N6723);
not NOT1 (N8620, N8619);
and AND3 (N8621, N8611, N2028, N7684);
nand NAND4 (N8622, N8616, N5792, N4359, N3275);
buf BUF1 (N8623, N8621);
nand NAND4 (N8624, N8612, N4022, N7408, N6020);
not NOT1 (N8625, N8620);
nor NOR2 (N8626, N8625, N3161);
nor NOR3 (N8627, N8624, N6667, N8191);
nand NAND2 (N8628, N8601, N8475);
and AND4 (N8629, N8626, N7504, N741, N8139);
xor XOR2 (N8630, N8623, N2732);
or OR2 (N8631, N8607, N4314);
nor NOR3 (N8632, N8622, N1396, N1129);
nand NAND4 (N8633, N8632, N5862, N6174, N3810);
nor NOR3 (N8634, N8631, N6350, N7506);
buf BUF1 (N8635, N8633);
not NOT1 (N8636, N8635);
or OR3 (N8637, N8629, N5500, N7817);
nand NAND3 (N8638, N8613, N5234, N1995);
nand NAND3 (N8639, N8630, N1257, N6540);
or OR2 (N8640, N8636, N6122);
or OR3 (N8641, N8618, N7731, N588);
xor XOR2 (N8642, N8606, N6428);
buf BUF1 (N8643, N8627);
buf BUF1 (N8644, N8638);
nand NAND4 (N8645, N8644, N7301, N4307, N4375);
xor XOR2 (N8646, N8645, N7032);
and AND3 (N8647, N8641, N6513, N8508);
nor NOR3 (N8648, N8615, N4207, N5451);
xor XOR2 (N8649, N8643, N201);
and AND4 (N8650, N8649, N5675, N7083, N4576);
nor NOR3 (N8651, N8639, N1331, N35);
or OR2 (N8652, N8640, N8146);
not NOT1 (N8653, N8628);
or OR3 (N8654, N8653, N1906, N6038);
buf BUF1 (N8655, N8646);
or OR3 (N8656, N8651, N7908, N3479);
or OR4 (N8657, N8652, N1246, N2796, N293);
buf BUF1 (N8658, N8634);
nor NOR4 (N8659, N8650, N7196, N3353, N3809);
nand NAND2 (N8660, N8637, N6863);
buf BUF1 (N8661, N8656);
nor NOR2 (N8662, N8658, N3331);
nor NOR2 (N8663, N8642, N6883);
nor NOR2 (N8664, N8648, N1555);
nor NOR2 (N8665, N8662, N4358);
and AND4 (N8666, N8660, N766, N4111, N5740);
and AND3 (N8667, N8665, N6843, N8452);
not NOT1 (N8668, N8663);
nor NOR3 (N8669, N8666, N597, N7796);
nor NOR2 (N8670, N8664, N33);
buf BUF1 (N8671, N8670);
nor NOR3 (N8672, N8671, N608, N3244);
and AND3 (N8673, N8647, N1169, N8076);
nor NOR4 (N8674, N8673, N2320, N5813, N6588);
and AND4 (N8675, N8674, N3583, N957, N6529);
xor XOR2 (N8676, N8655, N484);
and AND4 (N8677, N8657, N3416, N6105, N685);
and AND2 (N8678, N8668, N3206);
xor XOR2 (N8679, N8659, N5863);
nand NAND2 (N8680, N8676, N3248);
nand NAND4 (N8681, N8661, N7962, N517, N1457);
nor NOR4 (N8682, N8672, N6295, N452, N2891);
not NOT1 (N8683, N8682);
xor XOR2 (N8684, N8667, N3643);
nor NOR2 (N8685, N8679, N7606);
and AND2 (N8686, N8675, N7136);
xor XOR2 (N8687, N8684, N7892);
nor NOR3 (N8688, N8683, N6628, N1033);
nor NOR3 (N8689, N8680, N2971, N5334);
nand NAND3 (N8690, N8688, N3380, N910);
nor NOR4 (N8691, N8681, N1337, N591, N7279);
nor NOR3 (N8692, N8686, N1515, N7121);
nor NOR4 (N8693, N8677, N1928, N4238, N5722);
xor XOR2 (N8694, N8678, N5309);
nor NOR4 (N8695, N8691, N3695, N1040, N8219);
nand NAND4 (N8696, N8692, N2136, N4121, N1490);
or OR3 (N8697, N8689, N4487, N4240);
buf BUF1 (N8698, N8685);
and AND2 (N8699, N8696, N6961);
nand NAND2 (N8700, N8690, N5369);
nor NOR2 (N8701, N8699, N4573);
buf BUF1 (N8702, N8700);
nand NAND4 (N8703, N8701, N204, N2860, N1417);
and AND2 (N8704, N8703, N4630);
not NOT1 (N8705, N8693);
nor NOR3 (N8706, N8704, N8667, N2806);
nand NAND3 (N8707, N8694, N8419, N4680);
or OR4 (N8708, N8695, N8138, N8632, N7918);
not NOT1 (N8709, N8697);
or OR3 (N8710, N8709, N4274, N824);
and AND4 (N8711, N8698, N5733, N1242, N6553);
buf BUF1 (N8712, N8706);
xor XOR2 (N8713, N8669, N3961);
xor XOR2 (N8714, N8713, N4179);
or OR3 (N8715, N8705, N1163, N6475);
nand NAND2 (N8716, N8710, N5564);
buf BUF1 (N8717, N8687);
and AND3 (N8718, N8711, N1531, N3272);
buf BUF1 (N8719, N8708);
nor NOR4 (N8720, N8712, N5880, N6192, N1096);
nand NAND3 (N8721, N8702, N4370, N4809);
not NOT1 (N8722, N8714);
nand NAND3 (N8723, N8707, N7277, N7903);
buf BUF1 (N8724, N8715);
buf BUF1 (N8725, N8723);
nand NAND3 (N8726, N8722, N1976, N9);
nor NOR2 (N8727, N8717, N8281);
not NOT1 (N8728, N8727);
xor XOR2 (N8729, N8719, N3575);
xor XOR2 (N8730, N8716, N8698);
buf BUF1 (N8731, N8726);
buf BUF1 (N8732, N8718);
or OR4 (N8733, N8720, N7519, N2433, N60);
buf BUF1 (N8734, N8733);
not NOT1 (N8735, N8728);
nand NAND3 (N8736, N8730, N3608, N1972);
and AND3 (N8737, N8725, N2364, N7896);
and AND2 (N8738, N8654, N5969);
not NOT1 (N8739, N8738);
not NOT1 (N8740, N8737);
buf BUF1 (N8741, N8732);
and AND2 (N8742, N8736, N155);
nor NOR3 (N8743, N8735, N6560, N3712);
not NOT1 (N8744, N8724);
or OR2 (N8745, N8731, N6159);
not NOT1 (N8746, N8734);
or OR4 (N8747, N8742, N6158, N7507, N2755);
not NOT1 (N8748, N8746);
xor XOR2 (N8749, N8739, N6002);
or OR3 (N8750, N8721, N5200, N6870);
or OR2 (N8751, N8743, N7185);
or OR2 (N8752, N8740, N7111);
and AND2 (N8753, N8744, N792);
not NOT1 (N8754, N8751);
and AND2 (N8755, N8750, N3216);
buf BUF1 (N8756, N8747);
or OR3 (N8757, N8756, N7909, N7240);
and AND2 (N8758, N8754, N2411);
nor NOR2 (N8759, N8745, N8090);
xor XOR2 (N8760, N8753, N2798);
nor NOR3 (N8761, N8752, N4237, N5803);
and AND4 (N8762, N8741, N4738, N4818, N6990);
buf BUF1 (N8763, N8759);
or OR2 (N8764, N8760, N8335);
and AND2 (N8765, N8762, N1560);
buf BUF1 (N8766, N8765);
nand NAND3 (N8767, N8748, N1886, N7496);
nor NOR2 (N8768, N8729, N2003);
xor XOR2 (N8769, N8764, N1925);
nand NAND4 (N8770, N8757, N3732, N7480, N4672);
nand NAND2 (N8771, N8749, N379);
not NOT1 (N8772, N8761);
buf BUF1 (N8773, N8758);
or OR4 (N8774, N8755, N4814, N4689, N77);
nor NOR3 (N8775, N8769, N342, N8413);
nand NAND4 (N8776, N8774, N8480, N1305, N8404);
buf BUF1 (N8777, N8772);
xor XOR2 (N8778, N8777, N5588);
xor XOR2 (N8779, N8763, N5683);
nand NAND2 (N8780, N8773, N2284);
and AND3 (N8781, N8775, N4594, N6362);
xor XOR2 (N8782, N8778, N1150);
or OR2 (N8783, N8770, N5109);
and AND3 (N8784, N8781, N2817, N6722);
xor XOR2 (N8785, N8768, N3310);
nand NAND4 (N8786, N8783, N6539, N5752, N7423);
not NOT1 (N8787, N8771);
and AND3 (N8788, N8786, N4446, N5660);
xor XOR2 (N8789, N8780, N1496);
nand NAND4 (N8790, N8787, N3140, N1325, N1848);
nor NOR4 (N8791, N8784, N6861, N6945, N5943);
nor NOR3 (N8792, N8766, N5459, N7390);
or OR4 (N8793, N8792, N7533, N1547, N6694);
nor NOR4 (N8794, N8779, N101, N26, N7425);
and AND2 (N8795, N8790, N200);
not NOT1 (N8796, N8789);
buf BUF1 (N8797, N8785);
nor NOR2 (N8798, N8797, N4659);
xor XOR2 (N8799, N8794, N5717);
buf BUF1 (N8800, N8799);
or OR4 (N8801, N8776, N1223, N1451, N2064);
xor XOR2 (N8802, N8800, N4232);
buf BUF1 (N8803, N8801);
nand NAND2 (N8804, N8791, N2156);
or OR4 (N8805, N8793, N6624, N427, N5764);
or OR3 (N8806, N8802, N570, N7567);
nor NOR3 (N8807, N8798, N2800, N8692);
and AND4 (N8808, N8782, N5123, N2696, N7550);
nand NAND2 (N8809, N8788, N4718);
nand NAND4 (N8810, N8795, N919, N2814, N11);
nor NOR3 (N8811, N8809, N87, N2093);
nor NOR3 (N8812, N8810, N6739, N5420);
or OR3 (N8813, N8804, N3445, N5138);
nand NAND2 (N8814, N8808, N6651);
and AND3 (N8815, N8803, N4458, N2391);
not NOT1 (N8816, N8807);
or OR4 (N8817, N8796, N3527, N5054, N5914);
not NOT1 (N8818, N8815);
and AND3 (N8819, N8818, N5117, N7766);
or OR3 (N8820, N8811, N5122, N8059);
xor XOR2 (N8821, N8812, N5595);
not NOT1 (N8822, N8816);
buf BUF1 (N8823, N8805);
and AND3 (N8824, N8814, N3626, N3020);
nand NAND3 (N8825, N8819, N6207, N6172);
nand NAND3 (N8826, N8821, N4553, N7439);
nand NAND3 (N8827, N8826, N8788, N5893);
or OR4 (N8828, N8767, N4479, N8121, N4258);
or OR3 (N8829, N8828, N4151, N5049);
nand NAND4 (N8830, N8829, N7769, N7009, N219);
nor NOR4 (N8831, N8806, N3092, N6385, N4915);
nand NAND2 (N8832, N8824, N397);
nand NAND4 (N8833, N8813, N2450, N1871, N8810);
not NOT1 (N8834, N8820);
buf BUF1 (N8835, N8834);
xor XOR2 (N8836, N8835, N1385);
nor NOR3 (N8837, N8823, N1698, N4685);
not NOT1 (N8838, N8817);
buf BUF1 (N8839, N8833);
not NOT1 (N8840, N8831);
nor NOR2 (N8841, N8838, N8745);
not NOT1 (N8842, N8840);
not NOT1 (N8843, N8830);
and AND4 (N8844, N8843, N6332, N5147, N1781);
xor XOR2 (N8845, N8832, N8402);
xor XOR2 (N8846, N8845, N6448);
not NOT1 (N8847, N8839);
buf BUF1 (N8848, N8844);
xor XOR2 (N8849, N8837, N6749);
nor NOR3 (N8850, N8836, N5027, N4226);
xor XOR2 (N8851, N8827, N7888);
buf BUF1 (N8852, N8842);
xor XOR2 (N8853, N8850, N3681);
or OR2 (N8854, N8825, N7656);
buf BUF1 (N8855, N8853);
buf BUF1 (N8856, N8854);
or OR3 (N8857, N8846, N6926, N375);
nor NOR4 (N8858, N8856, N1485, N5845, N5139);
and AND2 (N8859, N8822, N3048);
or OR4 (N8860, N8848, N2548, N6400, N1405);
nand NAND3 (N8861, N8841, N1939, N8375);
and AND2 (N8862, N8855, N5777);
nor NOR4 (N8863, N8852, N1064, N2222, N7980);
nor NOR2 (N8864, N8862, N8119);
or OR3 (N8865, N8858, N6772, N5638);
and AND2 (N8866, N8860, N5098);
nand NAND2 (N8867, N8861, N2873);
buf BUF1 (N8868, N8865);
nor NOR3 (N8869, N8857, N7384, N8538);
xor XOR2 (N8870, N8868, N7970);
or OR4 (N8871, N8859, N4213, N1675, N6170);
xor XOR2 (N8872, N8864, N686);
not NOT1 (N8873, N8871);
nor NOR4 (N8874, N8863, N4620, N7489, N84);
or OR3 (N8875, N8849, N6329, N2281);
buf BUF1 (N8876, N8873);
buf BUF1 (N8877, N8851);
xor XOR2 (N8878, N8867, N2905);
not NOT1 (N8879, N8878);
nor NOR3 (N8880, N8866, N3351, N7613);
not NOT1 (N8881, N8847);
buf BUF1 (N8882, N8870);
or OR2 (N8883, N8880, N491);
or OR4 (N8884, N8879, N4305, N1289, N7185);
nand NAND3 (N8885, N8869, N3769, N8138);
buf BUF1 (N8886, N8872);
nor NOR3 (N8887, N8886, N2084, N5111);
xor XOR2 (N8888, N8885, N1264);
and AND4 (N8889, N8881, N6025, N130, N7707);
and AND3 (N8890, N8888, N3719, N8804);
not NOT1 (N8891, N8877);
or OR4 (N8892, N8882, N3750, N3180, N6815);
or OR3 (N8893, N8887, N1161, N8140);
and AND3 (N8894, N8892, N4735, N4726);
nor NOR2 (N8895, N8874, N3466);
nand NAND3 (N8896, N8876, N3373, N5445);
xor XOR2 (N8897, N8895, N4657);
nor NOR2 (N8898, N8896, N3695);
nor NOR4 (N8899, N8889, N6051, N4872, N3613);
and AND2 (N8900, N8893, N398);
nor NOR3 (N8901, N8899, N1775, N7316);
xor XOR2 (N8902, N8897, N8312);
xor XOR2 (N8903, N8891, N8748);
buf BUF1 (N8904, N8900);
or OR2 (N8905, N8883, N2085);
or OR2 (N8906, N8890, N4926);
xor XOR2 (N8907, N8884, N1478);
and AND3 (N8908, N8907, N5171, N8825);
nand NAND2 (N8909, N8894, N3881);
nor NOR4 (N8910, N8905, N2652, N1377, N5550);
nand NAND4 (N8911, N8909, N8457, N3770, N5307);
buf BUF1 (N8912, N8904);
xor XOR2 (N8913, N8906, N1293);
or OR2 (N8914, N8911, N7728);
nand NAND4 (N8915, N8875, N827, N4447, N6384);
and AND2 (N8916, N8901, N6070);
nand NAND2 (N8917, N8915, N7382);
nor NOR2 (N8918, N8914, N5935);
xor XOR2 (N8919, N8898, N6544);
xor XOR2 (N8920, N8918, N50);
nor NOR2 (N8921, N8916, N7409);
and AND3 (N8922, N8917, N8463, N4425);
or OR2 (N8923, N8922, N6032);
or OR4 (N8924, N8923, N7354, N7160, N2148);
nor NOR3 (N8925, N8919, N427, N3887);
and AND4 (N8926, N8910, N8623, N2047, N216);
nor NOR4 (N8927, N8902, N7189, N4346, N6074);
xor XOR2 (N8928, N8927, N1379);
nor NOR4 (N8929, N8928, N4357, N2834, N2736);
xor XOR2 (N8930, N8921, N3798);
or OR2 (N8931, N8912, N3504);
nor NOR4 (N8932, N8903, N5261, N2817, N3732);
nor NOR3 (N8933, N8924, N57, N4906);
nor NOR2 (N8934, N8929, N1627);
xor XOR2 (N8935, N8930, N5472);
nor NOR3 (N8936, N8931, N2622, N4293);
nand NAND3 (N8937, N8925, N7486, N5548);
buf BUF1 (N8938, N8926);
and AND4 (N8939, N8934, N284, N5438, N4194);
not NOT1 (N8940, N8908);
not NOT1 (N8941, N8938);
not NOT1 (N8942, N8935);
nand NAND2 (N8943, N8913, N1606);
xor XOR2 (N8944, N8939, N4590);
not NOT1 (N8945, N8942);
or OR4 (N8946, N8945, N6088, N4006, N3363);
or OR3 (N8947, N8932, N2293, N8790);
nor NOR4 (N8948, N8941, N1103, N7240, N1550);
nand NAND4 (N8949, N8936, N8567, N709, N8407);
nor NOR4 (N8950, N8946, N8249, N2794, N864);
nor NOR4 (N8951, N8943, N1211, N3902, N1311);
xor XOR2 (N8952, N8947, N600);
or OR4 (N8953, N8920, N4730, N1861, N1955);
xor XOR2 (N8954, N8940, N8363);
not NOT1 (N8955, N8950);
and AND3 (N8956, N8952, N7889, N4062);
or OR3 (N8957, N8937, N2565, N1177);
xor XOR2 (N8958, N8954, N1066);
nor NOR4 (N8959, N8957, N1546, N692, N25);
nand NAND3 (N8960, N8948, N6542, N1946);
buf BUF1 (N8961, N8958);
nand NAND2 (N8962, N8949, N618);
and AND3 (N8963, N8933, N2336, N5341);
and AND4 (N8964, N8944, N5202, N5498, N1436);
and AND2 (N8965, N8961, N5978);
or OR4 (N8966, N8964, N8644, N4178, N6442);
nor NOR4 (N8967, N8962, N7564, N7534, N4329);
buf BUF1 (N8968, N8966);
or OR3 (N8969, N8968, N4906, N635);
nand NAND3 (N8970, N8969, N5811, N5384);
buf BUF1 (N8971, N8967);
not NOT1 (N8972, N8960);
or OR2 (N8973, N8956, N8302);
xor XOR2 (N8974, N8973, N6706);
and AND4 (N8975, N8974, N8124, N6003, N564);
xor XOR2 (N8976, N8965, N8089);
and AND4 (N8977, N8971, N5209, N6178, N5151);
and AND3 (N8978, N8976, N6461, N6719);
nand NAND2 (N8979, N8977, N2895);
or OR3 (N8980, N8951, N7368, N62);
nand NAND4 (N8981, N8978, N4042, N8026, N819);
not NOT1 (N8982, N8980);
buf BUF1 (N8983, N8959);
nor NOR2 (N8984, N8963, N1009);
buf BUF1 (N8985, N8972);
nand NAND2 (N8986, N8982, N7083);
xor XOR2 (N8987, N8979, N3855);
nand NAND3 (N8988, N8955, N207, N3050);
and AND4 (N8989, N8988, N4436, N3362, N885);
or OR4 (N8990, N8989, N8324, N8128, N6371);
xor XOR2 (N8991, N8984, N7528);
buf BUF1 (N8992, N8987);
buf BUF1 (N8993, N8983);
buf BUF1 (N8994, N8991);
xor XOR2 (N8995, N8981, N1125);
nor NOR3 (N8996, N8994, N4080, N962);
nand NAND3 (N8997, N8953, N4972, N4227);
nand NAND2 (N8998, N8992, N710);
or OR4 (N8999, N8985, N8397, N3972, N5918);
and AND3 (N9000, N8975, N7816, N5290);
xor XOR2 (N9001, N8995, N5813);
not NOT1 (N9002, N8998);
and AND2 (N9003, N8999, N2609);
or OR2 (N9004, N8993, N6834);
and AND3 (N9005, N9002, N5164, N3321);
xor XOR2 (N9006, N8970, N8974);
not NOT1 (N9007, N9005);
buf BUF1 (N9008, N9001);
nor NOR2 (N9009, N9004, N459);
nor NOR4 (N9010, N9009, N2233, N3557, N4070);
not NOT1 (N9011, N9006);
not NOT1 (N9012, N9000);
buf BUF1 (N9013, N9012);
not NOT1 (N9014, N8996);
not NOT1 (N9015, N9013);
xor XOR2 (N9016, N9003, N7044);
buf BUF1 (N9017, N8997);
not NOT1 (N9018, N8986);
nand NAND2 (N9019, N9016, N7047);
xor XOR2 (N9020, N9008, N6760);
buf BUF1 (N9021, N9020);
or OR3 (N9022, N8990, N1481, N4669);
not NOT1 (N9023, N9011);
buf BUF1 (N9024, N9010);
nand NAND4 (N9025, N9015, N5476, N1219, N7381);
or OR3 (N9026, N9022, N256, N1634);
not NOT1 (N9027, N9019);
or OR3 (N9028, N9027, N1870, N5390);
not NOT1 (N9029, N9025);
nor NOR4 (N9030, N9017, N2293, N6802, N3199);
and AND2 (N9031, N9007, N1559);
and AND2 (N9032, N9030, N3922);
nand NAND4 (N9033, N9024, N3552, N7990, N4261);
and AND4 (N9034, N9018, N4293, N4016, N2228);
or OR2 (N9035, N9031, N342);
nand NAND2 (N9036, N9026, N3773);
and AND4 (N9037, N9021, N1410, N5684, N3210);
xor XOR2 (N9038, N9029, N8506);
and AND4 (N9039, N9035, N318, N999, N4270);
nand NAND4 (N9040, N9028, N4834, N2745, N2167);
buf BUF1 (N9041, N9023);
xor XOR2 (N9042, N9039, N8778);
and AND3 (N9043, N9038, N2869, N4355);
or OR4 (N9044, N9033, N2336, N3949, N5554);
nor NOR2 (N9045, N9043, N6841);
not NOT1 (N9046, N9044);
or OR2 (N9047, N9014, N3088);
and AND3 (N9048, N9041, N4722, N8715);
buf BUF1 (N9049, N9032);
and AND4 (N9050, N9046, N2528, N9032, N3552);
or OR3 (N9051, N9036, N6359, N502);
not NOT1 (N9052, N9049);
nand NAND2 (N9053, N9052, N4185);
or OR3 (N9054, N9050, N633, N8896);
xor XOR2 (N9055, N9047, N4047);
xor XOR2 (N9056, N9053, N143);
xor XOR2 (N9057, N9040, N3027);
nand NAND4 (N9058, N9048, N2567, N6762, N3049);
nor NOR3 (N9059, N9045, N8381, N6153);
nor NOR2 (N9060, N9058, N6324);
or OR2 (N9061, N9055, N6523);
or OR2 (N9062, N9037, N1681);
not NOT1 (N9063, N9051);
nor NOR3 (N9064, N9062, N381, N5267);
nor NOR3 (N9065, N9057, N1093, N1794);
nor NOR2 (N9066, N9034, N7846);
buf BUF1 (N9067, N9042);
xor XOR2 (N9068, N9059, N2873);
or OR2 (N9069, N9068, N7957);
buf BUF1 (N9070, N9054);
or OR4 (N9071, N9069, N3755, N6213, N2547);
and AND4 (N9072, N9061, N953, N1200, N8300);
xor XOR2 (N9073, N9072, N5247);
or OR4 (N9074, N9067, N928, N8754, N6131);
not NOT1 (N9075, N9071);
nand NAND3 (N9076, N9056, N7039, N3199);
buf BUF1 (N9077, N9066);
nor NOR3 (N9078, N9070, N2800, N8331);
nand NAND3 (N9079, N9063, N929, N8889);
nor NOR2 (N9080, N9060, N6004);
not NOT1 (N9081, N9073);
nand NAND3 (N9082, N9078, N861, N1195);
nand NAND4 (N9083, N9079, N127, N4318, N8615);
not NOT1 (N9084, N9080);
xor XOR2 (N9085, N9076, N5569);
nand NAND3 (N9086, N9065, N5372, N6493);
not NOT1 (N9087, N9084);
xor XOR2 (N9088, N9082, N6767);
nand NAND3 (N9089, N9087, N5459, N7410);
and AND3 (N9090, N9086, N3118, N3151);
and AND2 (N9091, N9089, N8911);
xor XOR2 (N9092, N9091, N6922);
or OR4 (N9093, N9090, N541, N8923, N2538);
nand NAND4 (N9094, N9081, N565, N5285, N5833);
nor NOR4 (N9095, N9074, N6157, N5923, N9080);
or OR2 (N9096, N9083, N2530);
nand NAND2 (N9097, N9092, N5311);
and AND2 (N9098, N9094, N4046);
and AND2 (N9099, N9095, N2007);
and AND3 (N9100, N9085, N1668, N7087);
or OR3 (N9101, N9099, N8520, N2393);
nor NOR2 (N9102, N9101, N957);
and AND3 (N9103, N9077, N1962, N4605);
not NOT1 (N9104, N9093);
and AND3 (N9105, N9102, N4058, N3004);
xor XOR2 (N9106, N9103, N5050);
buf BUF1 (N9107, N9096);
nand NAND2 (N9108, N9097, N5753);
not NOT1 (N9109, N9106);
nor NOR2 (N9110, N9108, N2612);
and AND3 (N9111, N9064, N2285, N8204);
nand NAND2 (N9112, N9100, N6748);
and AND3 (N9113, N9088, N4602, N6369);
nand NAND4 (N9114, N9105, N8591, N3313, N8848);
xor XOR2 (N9115, N9098, N5468);
or OR3 (N9116, N9107, N2245, N6446);
not NOT1 (N9117, N9075);
or OR3 (N9118, N9109, N1187, N3226);
xor XOR2 (N9119, N9111, N5493);
nor NOR3 (N9120, N9110, N3665, N1620);
buf BUF1 (N9121, N9104);
xor XOR2 (N9122, N9116, N5949);
xor XOR2 (N9123, N9118, N3321);
and AND3 (N9124, N9115, N7537, N411);
buf BUF1 (N9125, N9120);
or OR3 (N9126, N9122, N1110, N3838);
or OR2 (N9127, N9125, N6596);
and AND2 (N9128, N9121, N7556);
buf BUF1 (N9129, N9126);
or OR4 (N9130, N9119, N7248, N3263, N7959);
nand NAND3 (N9131, N9127, N16, N9088);
buf BUF1 (N9132, N9128);
buf BUF1 (N9133, N9129);
nor NOR2 (N9134, N9132, N8623);
xor XOR2 (N9135, N9133, N8431);
nand NAND3 (N9136, N9135, N2881, N6141);
nor NOR2 (N9137, N9134, N8724);
not NOT1 (N9138, N9131);
or OR3 (N9139, N9123, N3174, N5851);
and AND2 (N9140, N9124, N5626);
buf BUF1 (N9141, N9130);
buf BUF1 (N9142, N9136);
nor NOR4 (N9143, N9139, N6050, N1442, N3402);
buf BUF1 (N9144, N9112);
and AND2 (N9145, N9138, N2009);
and AND4 (N9146, N9144, N2646, N4579, N1570);
nor NOR2 (N9147, N9117, N2411);
not NOT1 (N9148, N9114);
xor XOR2 (N9149, N9147, N8163);
and AND4 (N9150, N9148, N1049, N2746, N8895);
or OR3 (N9151, N9150, N115, N3454);
nand NAND3 (N9152, N9149, N6347, N4149);
nor NOR2 (N9153, N9143, N1972);
nor NOR4 (N9154, N9141, N796, N7114, N4070);
or OR2 (N9155, N9154, N4353);
not NOT1 (N9156, N9140);
and AND4 (N9157, N9153, N1170, N212, N217);
buf BUF1 (N9158, N9157);
nand NAND4 (N9159, N9146, N5792, N4840, N4024);
or OR4 (N9160, N9137, N8432, N9094, N1977);
buf BUF1 (N9161, N9160);
buf BUF1 (N9162, N9145);
nand NAND4 (N9163, N9113, N3697, N1584, N6753);
not NOT1 (N9164, N9155);
xor XOR2 (N9165, N9158, N2498);
and AND2 (N9166, N9159, N3112);
or OR4 (N9167, N9156, N5917, N1950, N1590);
nand NAND2 (N9168, N9165, N8939);
and AND3 (N9169, N9167, N1615, N9167);
buf BUF1 (N9170, N9166);
nor NOR4 (N9171, N9163, N3591, N277, N3708);
nand NAND3 (N9172, N9151, N1883, N3685);
or OR4 (N9173, N9162, N2166, N4496, N7492);
nor NOR2 (N9174, N9161, N7031);
not NOT1 (N9175, N9168);
and AND3 (N9176, N9164, N3313, N4622);
buf BUF1 (N9177, N9171);
xor XOR2 (N9178, N9172, N8682);
nand NAND2 (N9179, N9142, N4258);
nor NOR3 (N9180, N9179, N8302, N509);
nand NAND2 (N9181, N9177, N5183);
and AND2 (N9182, N9181, N1807);
and AND4 (N9183, N9174, N5316, N3255, N1187);
buf BUF1 (N9184, N9180);
and AND3 (N9185, N9173, N990, N1548);
and AND3 (N9186, N9176, N7223, N2868);
nand NAND4 (N9187, N9184, N4032, N3209, N7536);
buf BUF1 (N9188, N9178);
buf BUF1 (N9189, N9175);
or OR2 (N9190, N9183, N613);
or OR2 (N9191, N9190, N6580);
or OR3 (N9192, N9182, N9182, N1118);
or OR2 (N9193, N9191, N2264);
or OR2 (N9194, N9189, N1044);
xor XOR2 (N9195, N9169, N1663);
and AND2 (N9196, N9188, N7187);
xor XOR2 (N9197, N9193, N8649);
nand NAND2 (N9198, N9185, N3090);
buf BUF1 (N9199, N9196);
not NOT1 (N9200, N9192);
xor XOR2 (N9201, N9187, N2260);
or OR3 (N9202, N9197, N5603, N9195);
nand NAND3 (N9203, N2253, N7352, N5919);
or OR2 (N9204, N9152, N5985);
and AND3 (N9205, N9203, N4291, N7883);
buf BUF1 (N9206, N9202);
xor XOR2 (N9207, N9186, N2310);
nor NOR2 (N9208, N9206, N1466);
xor XOR2 (N9209, N9208, N2456);
not NOT1 (N9210, N9201);
and AND4 (N9211, N9205, N4491, N278, N1930);
not NOT1 (N9212, N9207);
nand NAND2 (N9213, N9212, N7249);
nor NOR4 (N9214, N9209, N9162, N3249, N3561);
or OR4 (N9215, N9204, N1011, N3443, N2398);
buf BUF1 (N9216, N9214);
or OR4 (N9217, N9210, N303, N3848, N1829);
not NOT1 (N9218, N9217);
nor NOR4 (N9219, N9200, N6191, N5461, N6772);
or OR3 (N9220, N9218, N2362, N4470);
buf BUF1 (N9221, N9213);
not NOT1 (N9222, N9170);
xor XOR2 (N9223, N9221, N1574);
and AND2 (N9224, N9219, N3905);
nor NOR4 (N9225, N9199, N6591, N8146, N6257);
or OR3 (N9226, N9211, N6575, N2112);
nand NAND4 (N9227, N9198, N7301, N6812, N1735);
nand NAND3 (N9228, N9216, N1221, N3872);
buf BUF1 (N9229, N9226);
xor XOR2 (N9230, N9227, N3602);
nor NOR3 (N9231, N9225, N435, N5932);
xor XOR2 (N9232, N9223, N6625);
buf BUF1 (N9233, N9194);
xor XOR2 (N9234, N9231, N7386);
or OR2 (N9235, N9229, N3823);
xor XOR2 (N9236, N9215, N1144);
nor NOR2 (N9237, N9236, N9042);
and AND3 (N9238, N9228, N9098, N3843);
or OR4 (N9239, N9235, N708, N3103, N81);
xor XOR2 (N9240, N9224, N604);
not NOT1 (N9241, N9230);
buf BUF1 (N9242, N9237);
and AND2 (N9243, N9239, N489);
or OR4 (N9244, N9242, N8305, N7412, N6961);
not NOT1 (N9245, N9244);
xor XOR2 (N9246, N9220, N103);
xor XOR2 (N9247, N9234, N3015);
or OR3 (N9248, N9243, N7407, N1641);
and AND3 (N9249, N9238, N9199, N227);
or OR4 (N9250, N9232, N5963, N5886, N4824);
and AND3 (N9251, N9245, N7608, N2715);
xor XOR2 (N9252, N9246, N7668);
or OR2 (N9253, N9233, N7243);
not NOT1 (N9254, N9248);
nor NOR4 (N9255, N9247, N8269, N4072, N2491);
not NOT1 (N9256, N9249);
or OR2 (N9257, N9252, N5585);
or OR3 (N9258, N9222, N8179, N1173);
nor NOR2 (N9259, N9241, N1379);
nor NOR3 (N9260, N9253, N3979, N6254);
and AND3 (N9261, N9255, N6528, N6415);
and AND2 (N9262, N9251, N7939);
and AND2 (N9263, N9256, N8240);
and AND3 (N9264, N9250, N8950, N2069);
not NOT1 (N9265, N9263);
nor NOR4 (N9266, N9257, N5725, N6544, N6785);
not NOT1 (N9267, N9265);
buf BUF1 (N9268, N9266);
buf BUF1 (N9269, N9260);
and AND2 (N9270, N9258, N185);
or OR4 (N9271, N9269, N5207, N2795, N319);
buf BUF1 (N9272, N9271);
xor XOR2 (N9273, N9254, N3032);
not NOT1 (N9274, N9259);
xor XOR2 (N9275, N9262, N8796);
or OR4 (N9276, N9273, N5910, N4022, N226);
nor NOR4 (N9277, N9268, N3641, N1221, N7500);
and AND2 (N9278, N9267, N57);
nand NAND2 (N9279, N9274, N7334);
or OR2 (N9280, N9276, N5143);
xor XOR2 (N9281, N9272, N6683);
nand NAND2 (N9282, N9270, N4379);
nand NAND4 (N9283, N9240, N6944, N4220, N2464);
not NOT1 (N9284, N9264);
xor XOR2 (N9285, N9278, N3312);
buf BUF1 (N9286, N9261);
nand NAND2 (N9287, N9279, N8607);
buf BUF1 (N9288, N9284);
and AND2 (N9289, N9288, N5564);
nor NOR3 (N9290, N9289, N6603, N8384);
or OR3 (N9291, N9282, N1274, N1192);
and AND2 (N9292, N9275, N3736);
xor XOR2 (N9293, N9291, N8520);
not NOT1 (N9294, N9286);
xor XOR2 (N9295, N9293, N5921);
nor NOR3 (N9296, N9285, N4464, N1748);
not NOT1 (N9297, N9283);
not NOT1 (N9298, N9281);
or OR4 (N9299, N9277, N5818, N7135, N7989);
and AND4 (N9300, N9299, N6593, N8220, N1253);
nand NAND3 (N9301, N9287, N992, N1964);
nand NAND4 (N9302, N9300, N6917, N2562, N881);
and AND2 (N9303, N9292, N5604);
nor NOR3 (N9304, N9290, N951, N1204);
nand NAND3 (N9305, N9296, N6448, N5728);
nand NAND2 (N9306, N9304, N5316);
not NOT1 (N9307, N9295);
buf BUF1 (N9308, N9303);
xor XOR2 (N9309, N9302, N2069);
nor NOR2 (N9310, N9309, N2563);
nor NOR3 (N9311, N9305, N5975, N3902);
nor NOR4 (N9312, N9311, N2565, N2801, N5697);
nand NAND4 (N9313, N9310, N137, N6484, N512);
xor XOR2 (N9314, N9307, N5794);
and AND2 (N9315, N9312, N790);
nand NAND3 (N9316, N9301, N310, N9273);
or OR2 (N9317, N9314, N3152);
not NOT1 (N9318, N9315);
xor XOR2 (N9319, N9294, N2457);
xor XOR2 (N9320, N9313, N6194);
and AND2 (N9321, N9308, N6722);
xor XOR2 (N9322, N9317, N1578);
xor XOR2 (N9323, N9320, N3129);
or OR2 (N9324, N9316, N2606);
buf BUF1 (N9325, N9323);
nor NOR2 (N9326, N9298, N7094);
xor XOR2 (N9327, N9280, N9261);
and AND2 (N9328, N9322, N3678);
and AND2 (N9329, N9325, N7378);
not NOT1 (N9330, N9321);
nand NAND2 (N9331, N9318, N254);
buf BUF1 (N9332, N9331);
and AND3 (N9333, N9332, N1612, N844);
and AND4 (N9334, N9297, N3886, N4760, N5024);
not NOT1 (N9335, N9334);
or OR4 (N9336, N9319, N7672, N3970, N2253);
buf BUF1 (N9337, N9327);
not NOT1 (N9338, N9326);
not NOT1 (N9339, N9329);
buf BUF1 (N9340, N9338);
nand NAND3 (N9341, N9333, N8149, N6897);
buf BUF1 (N9342, N9341);
xor XOR2 (N9343, N9324, N5482);
xor XOR2 (N9344, N9339, N9098);
xor XOR2 (N9345, N9342, N5913);
buf BUF1 (N9346, N9337);
nor NOR2 (N9347, N9328, N477);
nand NAND2 (N9348, N9346, N3264);
or OR3 (N9349, N9345, N5853, N3094);
not NOT1 (N9350, N9349);
xor XOR2 (N9351, N9306, N2588);
nor NOR4 (N9352, N9335, N618, N7622, N5439);
not NOT1 (N9353, N9336);
nand NAND3 (N9354, N9348, N17, N3351);
not NOT1 (N9355, N9343);
nor NOR2 (N9356, N9347, N4424);
not NOT1 (N9357, N9330);
not NOT1 (N9358, N9357);
nand NAND2 (N9359, N9352, N8294);
xor XOR2 (N9360, N9344, N2194);
not NOT1 (N9361, N9353);
and AND2 (N9362, N9340, N9104);
not NOT1 (N9363, N9355);
buf BUF1 (N9364, N9363);
not NOT1 (N9365, N9358);
nor NOR4 (N9366, N9362, N2176, N6782, N9094);
and AND2 (N9367, N9359, N8080);
not NOT1 (N9368, N9367);
buf BUF1 (N9369, N9365);
nor NOR3 (N9370, N9354, N8729, N5346);
nor NOR4 (N9371, N9370, N5997, N250, N8259);
and AND4 (N9372, N9361, N5777, N8877, N4880);
or OR4 (N9373, N9369, N9321, N1316, N2455);
xor XOR2 (N9374, N9372, N4703);
and AND3 (N9375, N9371, N5376, N1428);
or OR2 (N9376, N9374, N2339);
nand NAND2 (N9377, N9356, N4567);
nand NAND2 (N9378, N9366, N5238);
xor XOR2 (N9379, N9351, N2563);
nand NAND4 (N9380, N9377, N5532, N4295, N2220);
not NOT1 (N9381, N9364);
or OR4 (N9382, N9360, N3717, N6837, N1170);
buf BUF1 (N9383, N9380);
and AND3 (N9384, N9375, N7467, N7410);
xor XOR2 (N9385, N9350, N5228);
nand NAND2 (N9386, N9373, N7488);
nand NAND2 (N9387, N9382, N7316);
nor NOR4 (N9388, N9383, N230, N2316, N8887);
nand NAND2 (N9389, N9387, N1536);
or OR2 (N9390, N9389, N1416);
xor XOR2 (N9391, N9384, N5656);
and AND2 (N9392, N9378, N4901);
xor XOR2 (N9393, N9388, N8327);
or OR4 (N9394, N9379, N7834, N3429, N6129);
nand NAND4 (N9395, N9394, N4351, N8444, N3181);
and AND4 (N9396, N9395, N7067, N3304, N1085);
nand NAND3 (N9397, N9393, N4610, N5333);
or OR3 (N9398, N9392, N230, N7738);
nor NOR4 (N9399, N9386, N3351, N7977, N8053);
buf BUF1 (N9400, N9399);
nand NAND4 (N9401, N9376, N982, N315, N8047);
not NOT1 (N9402, N9390);
nand NAND3 (N9403, N9385, N8578, N6238);
buf BUF1 (N9404, N9403);
nor NOR2 (N9405, N9404, N1997);
and AND2 (N9406, N9401, N6789);
xor XOR2 (N9407, N9405, N3202);
or OR3 (N9408, N9391, N2431, N5656);
not NOT1 (N9409, N9406);
or OR4 (N9410, N9407, N5239, N5551, N8328);
xor XOR2 (N9411, N9410, N5853);
buf BUF1 (N9412, N9398);
or OR2 (N9413, N9409, N2678);
and AND2 (N9414, N9400, N2017);
nor NOR4 (N9415, N9412, N3963, N4677, N1473);
or OR2 (N9416, N9402, N4947);
not NOT1 (N9417, N9368);
nor NOR2 (N9418, N9415, N8481);
nor NOR2 (N9419, N9411, N7135);
buf BUF1 (N9420, N9396);
not NOT1 (N9421, N9420);
or OR2 (N9422, N9419, N4023);
or OR4 (N9423, N9417, N8289, N2703, N5899);
nor NOR4 (N9424, N9413, N6973, N8265, N2526);
xor XOR2 (N9425, N9416, N4039);
not NOT1 (N9426, N9408);
xor XOR2 (N9427, N9397, N1086);
not NOT1 (N9428, N9427);
not NOT1 (N9429, N9381);
and AND2 (N9430, N9425, N8424);
xor XOR2 (N9431, N9418, N8901);
xor XOR2 (N9432, N9414, N7292);
and AND4 (N9433, N9430, N2564, N425, N5209);
and AND2 (N9434, N9426, N5770);
nand NAND3 (N9435, N9423, N4391, N6518);
or OR4 (N9436, N9433, N7211, N9067, N854);
not NOT1 (N9437, N9424);
not NOT1 (N9438, N9437);
not NOT1 (N9439, N9428);
xor XOR2 (N9440, N9421, N7051);
nand NAND4 (N9441, N9431, N8437, N1075, N6379);
xor XOR2 (N9442, N9429, N3033);
nor NOR3 (N9443, N9439, N7081, N4351);
nand NAND4 (N9444, N9436, N7388, N6963, N2383);
nand NAND3 (N9445, N9440, N8707, N4225);
or OR2 (N9446, N9441, N2763);
not NOT1 (N9447, N9442);
and AND3 (N9448, N9432, N6223, N676);
or OR4 (N9449, N9445, N1912, N5581, N5908);
or OR4 (N9450, N9444, N363, N674, N328);
or OR3 (N9451, N9435, N3268, N9224);
nand NAND4 (N9452, N9449, N3140, N5439, N8307);
nor NOR3 (N9453, N9434, N6489, N7677);
or OR2 (N9454, N9447, N296);
xor XOR2 (N9455, N9452, N5931);
and AND3 (N9456, N9451, N1030, N5688);
not NOT1 (N9457, N9438);
not NOT1 (N9458, N9448);
nand NAND2 (N9459, N9457, N3475);
not NOT1 (N9460, N9456);
xor XOR2 (N9461, N9455, N8645);
and AND4 (N9462, N9454, N2847, N8316, N2980);
xor XOR2 (N9463, N9458, N4999);
xor XOR2 (N9464, N9461, N5505);
nand NAND4 (N9465, N9463, N690, N5293, N7423);
and AND3 (N9466, N9460, N1389, N2094);
xor XOR2 (N9467, N9422, N5638);
not NOT1 (N9468, N9464);
nor NOR2 (N9469, N9466, N5337);
or OR4 (N9470, N9453, N5551, N3701, N9308);
or OR4 (N9471, N9469, N3582, N4703, N1844);
and AND4 (N9472, N9459, N6933, N4888, N6185);
buf BUF1 (N9473, N9472);
and AND2 (N9474, N9473, N3179);
not NOT1 (N9475, N9467);
nand NAND4 (N9476, N9470, N9309, N5528, N5814);
and AND4 (N9477, N9465, N9265, N5765, N5808);
and AND2 (N9478, N9471, N1695);
nand NAND4 (N9479, N9446, N2479, N4426, N1295);
and AND2 (N9480, N9476, N7309);
not NOT1 (N9481, N9477);
xor XOR2 (N9482, N9479, N1951);
or OR4 (N9483, N9443, N8174, N7433, N5709);
and AND3 (N9484, N9474, N4363, N872);
and AND3 (N9485, N9484, N4970, N3179);
nor NOR2 (N9486, N9478, N619);
buf BUF1 (N9487, N9481);
nor NOR3 (N9488, N9450, N4512, N6262);
xor XOR2 (N9489, N9485, N7887);
and AND2 (N9490, N9482, N1726);
not NOT1 (N9491, N9487);
nor NOR2 (N9492, N9483, N4772);
buf BUF1 (N9493, N9475);
buf BUF1 (N9494, N9468);
buf BUF1 (N9495, N9462);
or OR3 (N9496, N9494, N376, N6106);
nand NAND3 (N9497, N9486, N5058, N3982);
nor NOR3 (N9498, N9497, N6107, N3335);
or OR2 (N9499, N9480, N802);
nor NOR2 (N9500, N9492, N5484);
not NOT1 (N9501, N9489);
and AND3 (N9502, N9495, N9309, N5919);
nor NOR4 (N9503, N9499, N6183, N8667, N1840);
not NOT1 (N9504, N9496);
nand NAND3 (N9505, N9491, N1879, N264);
xor XOR2 (N9506, N9504, N4178);
or OR2 (N9507, N9500, N5033);
xor XOR2 (N9508, N9505, N2982);
nor NOR2 (N9509, N9502, N3942);
not NOT1 (N9510, N9509);
or OR3 (N9511, N9508, N20, N8707);
and AND2 (N9512, N9490, N2928);
buf BUF1 (N9513, N9506);
buf BUF1 (N9514, N9498);
and AND3 (N9515, N9501, N5096, N8941);
not NOT1 (N9516, N9510);
xor XOR2 (N9517, N9516, N9023);
or OR3 (N9518, N9507, N4559, N4770);
nand NAND3 (N9519, N9513, N6367, N8372);
not NOT1 (N9520, N9493);
or OR3 (N9521, N9503, N56, N419);
or OR2 (N9522, N9517, N4941);
buf BUF1 (N9523, N9515);
nor NOR2 (N9524, N9512, N1075);
nor NOR2 (N9525, N9521, N34);
buf BUF1 (N9526, N9514);
and AND2 (N9527, N9525, N2913);
not NOT1 (N9528, N9524);
nand NAND2 (N9529, N9518, N8678);
buf BUF1 (N9530, N9526);
not NOT1 (N9531, N9529);
and AND3 (N9532, N9527, N519, N6034);
nor NOR2 (N9533, N9530, N2142);
xor XOR2 (N9534, N9532, N1412);
nor NOR2 (N9535, N9511, N1176);
or OR2 (N9536, N9534, N4469);
or OR2 (N9537, N9488, N5903);
buf BUF1 (N9538, N9536);
not NOT1 (N9539, N9533);
xor XOR2 (N9540, N9537, N7800);
and AND3 (N9541, N9528, N5189, N898);
not NOT1 (N9542, N9540);
and AND3 (N9543, N9538, N1289, N7299);
xor XOR2 (N9544, N9522, N7318);
not NOT1 (N9545, N9523);
not NOT1 (N9546, N9544);
and AND2 (N9547, N9546, N7182);
nor NOR4 (N9548, N9539, N2614, N844, N7585);
nand NAND4 (N9549, N9535, N5193, N6146, N2438);
and AND3 (N9550, N9520, N8112, N1375);
nand NAND2 (N9551, N9541, N2845);
nor NOR4 (N9552, N9545, N7386, N340, N929);
not NOT1 (N9553, N9552);
nand NAND3 (N9554, N9543, N4845, N3569);
or OR4 (N9555, N9549, N8086, N805, N9384);
buf BUF1 (N9556, N9555);
buf BUF1 (N9557, N9531);
nor NOR3 (N9558, N9554, N3739, N3487);
not NOT1 (N9559, N9551);
or OR3 (N9560, N9547, N3971, N8912);
nand NAND3 (N9561, N9553, N5440, N116);
xor XOR2 (N9562, N9560, N9505);
not NOT1 (N9563, N9556);
xor XOR2 (N9564, N9561, N9363);
nor NOR4 (N9565, N9557, N1244, N3277, N5550);
xor XOR2 (N9566, N9550, N9006);
and AND4 (N9567, N9562, N8776, N3933, N2602);
or OR3 (N9568, N9566, N2917, N6134);
xor XOR2 (N9569, N9563, N6390);
nor NOR2 (N9570, N9558, N8612);
xor XOR2 (N9571, N9564, N7960);
and AND3 (N9572, N9568, N4501, N7023);
and AND2 (N9573, N9519, N3471);
xor XOR2 (N9574, N9565, N4825);
not NOT1 (N9575, N9571);
nor NOR4 (N9576, N9559, N3808, N3082, N6636);
xor XOR2 (N9577, N9548, N2684);
xor XOR2 (N9578, N9542, N4784);
or OR4 (N9579, N9574, N1645, N5295, N502);
or OR2 (N9580, N9575, N1658);
not NOT1 (N9581, N9567);
or OR2 (N9582, N9572, N6781);
nor NOR3 (N9583, N9582, N3432, N2115);
buf BUF1 (N9584, N9569);
not NOT1 (N9585, N9580);
buf BUF1 (N9586, N9585);
nand NAND4 (N9587, N9581, N4431, N3853, N781);
nand NAND4 (N9588, N9584, N1211, N2412, N3512);
xor XOR2 (N9589, N9588, N1265);
xor XOR2 (N9590, N9573, N2172);
xor XOR2 (N9591, N9570, N388);
or OR2 (N9592, N9577, N4296);
not NOT1 (N9593, N9591);
or OR2 (N9594, N9587, N2671);
and AND4 (N9595, N9578, N8268, N1378, N3056);
nor NOR4 (N9596, N9589, N3698, N6376, N9270);
buf BUF1 (N9597, N9593);
not NOT1 (N9598, N9576);
nor NOR3 (N9599, N9592, N4828, N4803);
nor NOR3 (N9600, N9594, N9228, N3913);
xor XOR2 (N9601, N9583, N4980);
and AND3 (N9602, N9579, N8839, N4743);
xor XOR2 (N9603, N9598, N3236);
xor XOR2 (N9604, N9595, N6475);
nand NAND4 (N9605, N9590, N7008, N799, N1734);
and AND2 (N9606, N9602, N1873);
nand NAND2 (N9607, N9586, N6515);
not NOT1 (N9608, N9603);
not NOT1 (N9609, N9604);
not NOT1 (N9610, N9609);
buf BUF1 (N9611, N9601);
buf BUF1 (N9612, N9600);
and AND4 (N9613, N9608, N2193, N2918, N4822);
not NOT1 (N9614, N9605);
and AND4 (N9615, N9610, N4446, N6115, N4980);
xor XOR2 (N9616, N9606, N2137);
and AND3 (N9617, N9614, N1787, N1456);
or OR4 (N9618, N9611, N1766, N1358, N49);
and AND3 (N9619, N9599, N2581, N8555);
not NOT1 (N9620, N9617);
nor NOR2 (N9621, N9607, N4031);
or OR2 (N9622, N9619, N4410);
buf BUF1 (N9623, N9612);
buf BUF1 (N9624, N9621);
nor NOR2 (N9625, N9615, N2008);
nand NAND2 (N9626, N9618, N5582);
and AND2 (N9627, N9597, N9601);
and AND3 (N9628, N9596, N2928, N9115);
buf BUF1 (N9629, N9625);
buf BUF1 (N9630, N9620);
nand NAND4 (N9631, N9630, N6497, N496, N6749);
not NOT1 (N9632, N9616);
and AND3 (N9633, N9629, N7659, N1199);
nand NAND4 (N9634, N9626, N4495, N8809, N5160);
not NOT1 (N9635, N9634);
not NOT1 (N9636, N9624);
not NOT1 (N9637, N9613);
buf BUF1 (N9638, N9636);
buf BUF1 (N9639, N9632);
not NOT1 (N9640, N9622);
nor NOR2 (N9641, N9639, N2575);
xor XOR2 (N9642, N9628, N4136);
nand NAND2 (N9643, N9623, N9613);
not NOT1 (N9644, N9637);
xor XOR2 (N9645, N9641, N3241);
or OR3 (N9646, N9640, N1640, N9574);
not NOT1 (N9647, N9627);
or OR4 (N9648, N9647, N9250, N8687, N9563);
xor XOR2 (N9649, N9643, N1098);
nor NOR2 (N9650, N9645, N9401);
buf BUF1 (N9651, N9638);
not NOT1 (N9652, N9635);
and AND3 (N9653, N9650, N5329, N569);
not NOT1 (N9654, N9633);
and AND2 (N9655, N9654, N6314);
nor NOR4 (N9656, N9642, N599, N4122, N5557);
not NOT1 (N9657, N9644);
nor NOR2 (N9658, N9646, N1544);
or OR4 (N9659, N9648, N2543, N5364, N3084);
not NOT1 (N9660, N9651);
nor NOR3 (N9661, N9649, N4451, N2324);
or OR4 (N9662, N9655, N5858, N2182, N1856);
nor NOR3 (N9663, N9657, N5183, N4701);
or OR4 (N9664, N9631, N7677, N3850, N1671);
xor XOR2 (N9665, N9661, N8449);
not NOT1 (N9666, N9664);
or OR4 (N9667, N9665, N1949, N6435, N9425);
nor NOR2 (N9668, N9652, N3261);
xor XOR2 (N9669, N9666, N5704);
or OR2 (N9670, N9659, N7058);
nand NAND2 (N9671, N9668, N8180);
xor XOR2 (N9672, N9667, N5821);
xor XOR2 (N9673, N9656, N8173);
or OR3 (N9674, N9669, N993, N2566);
nor NOR2 (N9675, N9653, N4770);
buf BUF1 (N9676, N9674);
nor NOR4 (N9677, N9672, N1925, N7519, N5156);
nor NOR4 (N9678, N9670, N6547, N6472, N7246);
nor NOR2 (N9679, N9663, N8560);
not NOT1 (N9680, N9671);
not NOT1 (N9681, N9660);
or OR3 (N9682, N9681, N5383, N3006);
xor XOR2 (N9683, N9676, N3627);
xor XOR2 (N9684, N9677, N5527);
xor XOR2 (N9685, N9673, N7706);
xor XOR2 (N9686, N9685, N1987);
and AND4 (N9687, N9658, N1770, N642, N3301);
and AND3 (N9688, N9684, N792, N6255);
not NOT1 (N9689, N9662);
or OR3 (N9690, N9683, N7015, N4682);
xor XOR2 (N9691, N9686, N6252);
nand NAND4 (N9692, N9679, N6768, N2841, N4761);
nor NOR2 (N9693, N9692, N6481);
nor NOR3 (N9694, N9687, N3905, N6474);
nand NAND3 (N9695, N9694, N7701, N6725);
or OR3 (N9696, N9678, N3519, N5431);
or OR4 (N9697, N9689, N3949, N8288, N830);
or OR4 (N9698, N9695, N5779, N8603, N946);
not NOT1 (N9699, N9675);
buf BUF1 (N9700, N9699);
nor NOR3 (N9701, N9697, N2624, N7846);
and AND4 (N9702, N9690, N2786, N4962, N165);
nor NOR3 (N9703, N9700, N7789, N5512);
and AND4 (N9704, N9702, N4059, N3298, N4515);
nor NOR4 (N9705, N9704, N2465, N2398, N6015);
or OR3 (N9706, N9705, N7779, N9130);
buf BUF1 (N9707, N9703);
or OR2 (N9708, N9693, N7664);
nand NAND4 (N9709, N9708, N472, N9640, N6819);
nor NOR4 (N9710, N9701, N6527, N6658, N113);
or OR2 (N9711, N9696, N6496);
and AND2 (N9712, N9706, N6958);
nor NOR3 (N9713, N9682, N6894, N2973);
and AND4 (N9714, N9712, N3539, N3827, N8185);
not NOT1 (N9715, N9711);
and AND4 (N9716, N9710, N1126, N8828, N4379);
and AND3 (N9717, N9714, N4821, N2618);
buf BUF1 (N9718, N9691);
nand NAND4 (N9719, N9688, N282, N4903, N6792);
or OR3 (N9720, N9717, N1194, N4061);
and AND4 (N9721, N9719, N1144, N4213, N6467);
nand NAND3 (N9722, N9709, N7192, N5757);
nor NOR4 (N9723, N9716, N7273, N2279, N4659);
nand NAND3 (N9724, N9720, N7897, N1682);
xor XOR2 (N9725, N9698, N7620);
or OR2 (N9726, N9725, N1433);
buf BUF1 (N9727, N9724);
xor XOR2 (N9728, N9715, N92);
or OR3 (N9729, N9728, N2095, N6397);
buf BUF1 (N9730, N9722);
nor NOR2 (N9731, N9713, N970);
buf BUF1 (N9732, N9727);
nor NOR3 (N9733, N9729, N5513, N7655);
buf BUF1 (N9734, N9731);
xor XOR2 (N9735, N9732, N353);
nand NAND2 (N9736, N9723, N7479);
and AND2 (N9737, N9733, N1532);
buf BUF1 (N9738, N9726);
nor NOR2 (N9739, N9721, N619);
nor NOR3 (N9740, N9736, N3287, N122);
nor NOR4 (N9741, N9707, N6254, N843, N2577);
xor XOR2 (N9742, N9734, N1282);
xor XOR2 (N9743, N9680, N1268);
nor NOR3 (N9744, N9743, N7935, N9371);
xor XOR2 (N9745, N9718, N3372);
xor XOR2 (N9746, N9738, N4003);
nor NOR3 (N9747, N9739, N4594, N3526);
or OR4 (N9748, N9741, N8516, N2065, N1630);
xor XOR2 (N9749, N9740, N8731);
buf BUF1 (N9750, N9737);
not NOT1 (N9751, N9745);
and AND3 (N9752, N9749, N1639, N7533);
buf BUF1 (N9753, N9742);
or OR3 (N9754, N9730, N6651, N3533);
or OR2 (N9755, N9752, N2286);
and AND2 (N9756, N9751, N4111);
nor NOR4 (N9757, N9754, N8123, N7296, N3093);
buf BUF1 (N9758, N9744);
or OR2 (N9759, N9735, N6677);
nand NAND2 (N9760, N9750, N2236);
buf BUF1 (N9761, N9748);
or OR3 (N9762, N9759, N1028, N1130);
nor NOR3 (N9763, N9758, N9217, N5435);
not NOT1 (N9764, N9761);
xor XOR2 (N9765, N9760, N598);
or OR2 (N9766, N9757, N5374);
not NOT1 (N9767, N9756);
and AND2 (N9768, N9747, N3589);
and AND2 (N9769, N9753, N3365);
nor NOR3 (N9770, N9768, N1044, N94);
and AND2 (N9771, N9765, N6566);
not NOT1 (N9772, N9770);
not NOT1 (N9773, N9771);
or OR3 (N9774, N9764, N7086, N4980);
buf BUF1 (N9775, N9773);
and AND2 (N9776, N9762, N940);
and AND4 (N9777, N9775, N4151, N2247, N7791);
buf BUF1 (N9778, N9766);
xor XOR2 (N9779, N9767, N5849);
or OR3 (N9780, N9777, N664, N4969);
buf BUF1 (N9781, N9778);
xor XOR2 (N9782, N9774, N9338);
nand NAND3 (N9783, N9746, N8516, N5793);
or OR2 (N9784, N9769, N5965);
or OR4 (N9785, N9784, N3319, N2619, N3106);
nor NOR4 (N9786, N9782, N3121, N9523, N1492);
and AND4 (N9787, N9776, N9658, N9335, N7913);
xor XOR2 (N9788, N9783, N304);
nand NAND4 (N9789, N9779, N6371, N201, N9547);
and AND4 (N9790, N9786, N8180, N2855, N6251);
nand NAND4 (N9791, N9788, N4454, N4717, N273);
or OR2 (N9792, N9785, N3947);
buf BUF1 (N9793, N9792);
and AND3 (N9794, N9763, N4130, N7800);
nor NOR4 (N9795, N9781, N2696, N2506, N951);
xor XOR2 (N9796, N9772, N6124);
and AND3 (N9797, N9787, N3885, N5704);
buf BUF1 (N9798, N9789);
nor NOR2 (N9799, N9798, N1014);
not NOT1 (N9800, N9795);
or OR4 (N9801, N9780, N1466, N7515, N5885);
not NOT1 (N9802, N9796);
nor NOR4 (N9803, N9801, N7538, N6372, N4221);
and AND4 (N9804, N9797, N2868, N4742, N7997);
xor XOR2 (N9805, N9791, N7905);
not NOT1 (N9806, N9794);
nand NAND2 (N9807, N9804, N2779);
nand NAND3 (N9808, N9802, N9394, N2359);
or OR4 (N9809, N9805, N8513, N5820, N2399);
buf BUF1 (N9810, N9799);
buf BUF1 (N9811, N9803);
and AND2 (N9812, N9811, N7908);
buf BUF1 (N9813, N9806);
not NOT1 (N9814, N9793);
and AND3 (N9815, N9810, N2742, N8176);
or OR3 (N9816, N9755, N3366, N9389);
nand NAND2 (N9817, N9814, N1851);
xor XOR2 (N9818, N9800, N1965);
not NOT1 (N9819, N9808);
not NOT1 (N9820, N9816);
nand NAND4 (N9821, N9812, N7756, N204, N9553);
and AND2 (N9822, N9815, N9454);
or OR4 (N9823, N9822, N7904, N9783, N2190);
nand NAND2 (N9824, N9809, N7118);
nor NOR4 (N9825, N9819, N2341, N2255, N8317);
and AND4 (N9826, N9824, N7125, N7767, N7247);
and AND3 (N9827, N9813, N8652, N2718);
and AND4 (N9828, N9820, N6286, N5231, N1806);
buf BUF1 (N9829, N9827);
nand NAND2 (N9830, N9818, N5198);
not NOT1 (N9831, N9829);
nor NOR2 (N9832, N9790, N9410);
not NOT1 (N9833, N9830);
nor NOR4 (N9834, N9823, N5508, N1158, N9450);
xor XOR2 (N9835, N9821, N5828);
nand NAND4 (N9836, N9835, N8423, N4337, N8382);
nand NAND4 (N9837, N9833, N759, N5085, N2247);
or OR3 (N9838, N9832, N18, N9580);
or OR3 (N9839, N9834, N8780, N1015);
buf BUF1 (N9840, N9837);
buf BUF1 (N9841, N9839);
and AND2 (N9842, N9831, N5372);
or OR4 (N9843, N9842, N8042, N4650, N5608);
nand NAND3 (N9844, N9838, N8370, N428);
xor XOR2 (N9845, N9826, N693);
nand NAND3 (N9846, N9807, N8730, N5683);
and AND2 (N9847, N9825, N9580);
or OR2 (N9848, N9846, N7710);
not NOT1 (N9849, N9828);
xor XOR2 (N9850, N9843, N5653);
nand NAND4 (N9851, N9845, N3901, N4057, N7610);
or OR3 (N9852, N9851, N6570, N2452);
nand NAND3 (N9853, N9840, N1014, N1723);
nor NOR3 (N9854, N9817, N7388, N7398);
or OR4 (N9855, N9852, N4884, N3380, N6918);
nor NOR3 (N9856, N9844, N3856, N2105);
nand NAND4 (N9857, N9854, N2330, N8413, N1397);
nor NOR4 (N9858, N9857, N8030, N3565, N6545);
nor NOR3 (N9859, N9855, N3338, N6226);
nor NOR4 (N9860, N9836, N9706, N1992, N5806);
nor NOR4 (N9861, N9853, N2789, N2178, N9544);
and AND3 (N9862, N9858, N5519, N5858);
or OR3 (N9863, N9860, N2452, N511);
nand NAND4 (N9864, N9861, N3825, N2693, N3940);
or OR4 (N9865, N9864, N594, N5948, N4449);
nor NOR2 (N9866, N9862, N3061);
nor NOR3 (N9867, N9863, N1191, N4220);
nand NAND4 (N9868, N9867, N7427, N3971, N9791);
nand NAND3 (N9869, N9856, N4936, N3754);
nor NOR2 (N9870, N9859, N2306);
nand NAND4 (N9871, N9870, N3211, N230, N3936);
and AND4 (N9872, N9869, N747, N3356, N4166);
not NOT1 (N9873, N9871);
nor NOR2 (N9874, N9841, N212);
nand NAND2 (N9875, N9866, N4601);
xor XOR2 (N9876, N9868, N2909);
buf BUF1 (N9877, N9874);
xor XOR2 (N9878, N9849, N9747);
xor XOR2 (N9879, N9865, N3043);
nor NOR3 (N9880, N9877, N3787, N1828);
xor XOR2 (N9881, N9872, N2487);
nor NOR4 (N9882, N9878, N4194, N583, N8808);
buf BUF1 (N9883, N9873);
not NOT1 (N9884, N9881);
xor XOR2 (N9885, N9876, N8412);
and AND2 (N9886, N9880, N1764);
and AND4 (N9887, N9884, N7445, N9337, N2774);
nand NAND4 (N9888, N9885, N5321, N3172, N6840);
xor XOR2 (N9889, N9882, N5064);
and AND4 (N9890, N9847, N4825, N403, N2043);
nand NAND3 (N9891, N9890, N1549, N5129);
nor NOR3 (N9892, N9889, N131, N561);
or OR3 (N9893, N9891, N3360, N7443);
xor XOR2 (N9894, N9850, N4859);
nor NOR4 (N9895, N9894, N226, N5969, N5424);
and AND3 (N9896, N9848, N2686, N6404);
not NOT1 (N9897, N9888);
and AND3 (N9898, N9887, N9540, N6700);
nand NAND3 (N9899, N9897, N1909, N6820);
buf BUF1 (N9900, N9883);
not NOT1 (N9901, N9875);
nand NAND3 (N9902, N9879, N9647, N6963);
buf BUF1 (N9903, N9902);
nor NOR4 (N9904, N9901, N1717, N4590, N925);
or OR3 (N9905, N9899, N2771, N4102);
nor NOR4 (N9906, N9893, N1063, N3280, N3955);
xor XOR2 (N9907, N9896, N9383);
buf BUF1 (N9908, N9907);
nor NOR4 (N9909, N9904, N5556, N9296, N771);
nand NAND4 (N9910, N9886, N6606, N6078, N4614);
and AND2 (N9911, N9905, N522);
buf BUF1 (N9912, N9900);
not NOT1 (N9913, N9912);
buf BUF1 (N9914, N9913);
nor NOR4 (N9915, N9906, N1239, N8642, N9458);
nand NAND4 (N9916, N9908, N1096, N3648, N7243);
nand NAND2 (N9917, N9916, N6508);
not NOT1 (N9918, N9903);
and AND4 (N9919, N9909, N8209, N8523, N781);
or OR3 (N9920, N9914, N2839, N124);
and AND3 (N9921, N9910, N4499, N4823);
not NOT1 (N9922, N9915);
nand NAND4 (N9923, N9918, N4584, N8568, N2359);
xor XOR2 (N9924, N9923, N5232);
buf BUF1 (N9925, N9892);
nand NAND2 (N9926, N9917, N8704);
nor NOR4 (N9927, N9922, N712, N616, N7203);
nand NAND2 (N9928, N9926, N5558);
xor XOR2 (N9929, N9919, N7067);
nor NOR3 (N9930, N9920, N5962, N8302);
nor NOR3 (N9931, N9924, N1715, N4464);
not NOT1 (N9932, N9930);
nor NOR3 (N9933, N9895, N925, N6160);
and AND4 (N9934, N9931, N7264, N7398, N8047);
buf BUF1 (N9935, N9921);
or OR4 (N9936, N9929, N31, N5658, N8985);
not NOT1 (N9937, N9927);
buf BUF1 (N9938, N9935);
not NOT1 (N9939, N9932);
and AND2 (N9940, N9936, N8952);
and AND4 (N9941, N9940, N4388, N6755, N1038);
nor NOR3 (N9942, N9934, N1615, N2095);
nor NOR3 (N9943, N9942, N9668, N312);
buf BUF1 (N9944, N9933);
buf BUF1 (N9945, N9944);
and AND3 (N9946, N9941, N1477, N2027);
nand NAND3 (N9947, N9943, N6295, N6312);
nand NAND3 (N9948, N9945, N2376, N6770);
nand NAND3 (N9949, N9928, N8695, N1762);
xor XOR2 (N9950, N9911, N427);
nand NAND3 (N9951, N9938, N489, N5471);
nor NOR2 (N9952, N9947, N7136);
or OR2 (N9953, N9950, N6439);
buf BUF1 (N9954, N9951);
buf BUF1 (N9955, N9954);
xor XOR2 (N9956, N9939, N2153);
nor NOR4 (N9957, N9955, N4733, N9102, N5581);
or OR2 (N9958, N9937, N1035);
and AND2 (N9959, N9952, N5066);
and AND3 (N9960, N9957, N6217, N9751);
or OR2 (N9961, N9949, N3455);
and AND3 (N9962, N9946, N907, N6809);
or OR2 (N9963, N9959, N4212);
nand NAND2 (N9964, N9925, N2401);
or OR3 (N9965, N9963, N7194, N7000);
not NOT1 (N9966, N9965);
and AND2 (N9967, N9948, N2199);
buf BUF1 (N9968, N9962);
nor NOR3 (N9969, N9898, N6753, N4792);
not NOT1 (N9970, N9953);
nor NOR4 (N9971, N9961, N3436, N8603, N7720);
or OR4 (N9972, N9958, N1913, N5137, N5693);
nand NAND2 (N9973, N9971, N7056);
buf BUF1 (N9974, N9969);
xor XOR2 (N9975, N9972, N4057);
nor NOR4 (N9976, N9975, N8071, N7860, N7003);
and AND2 (N9977, N9973, N9715);
nand NAND3 (N9978, N9970, N3549, N8853);
xor XOR2 (N9979, N9960, N1699);
buf BUF1 (N9980, N9956);
and AND2 (N9981, N9978, N7375);
nand NAND3 (N9982, N9976, N9628, N2935);
nand NAND3 (N9983, N9982, N5477, N8942);
nor NOR4 (N9984, N9981, N1776, N7118, N1527);
buf BUF1 (N9985, N9983);
and AND3 (N9986, N9977, N1703, N9943);
and AND2 (N9987, N9979, N4624);
nor NOR3 (N9988, N9968, N8114, N3902);
xor XOR2 (N9989, N9980, N5460);
buf BUF1 (N9990, N9985);
and AND3 (N9991, N9964, N91, N5441);
nand NAND3 (N9992, N9991, N4915, N7171);
nor NOR3 (N9993, N9987, N3883, N4199);
nand NAND4 (N9994, N9988, N8906, N9215, N9732);
not NOT1 (N9995, N9993);
nor NOR3 (N9996, N9990, N494, N801);
or OR3 (N9997, N9974, N2944, N1252);
nand NAND2 (N9998, N9996, N7483);
buf BUF1 (N9999, N9966);
or OR2 (N10000, N9998, N3595);
xor XOR2 (N10001, N9967, N9562);
nand NAND3 (N10002, N9999, N1802, N1375);
and AND2 (N10003, N9994, N4113);
xor XOR2 (N10004, N9986, N4280);
nand NAND2 (N10005, N10003, N5740);
nor NOR3 (N10006, N10004, N5538, N9007);
and AND4 (N10007, N10005, N5027, N4306, N9299);
nor NOR2 (N10008, N9984, N2604);
xor XOR2 (N10009, N10007, N3332);
nand NAND4 (N10010, N10006, N7924, N9336, N3837);
or OR4 (N10011, N10002, N5316, N9394, N6770);
xor XOR2 (N10012, N10009, N2493);
nor NOR2 (N10013, N10000, N2173);
and AND3 (N10014, N10008, N9988, N3602);
nand NAND2 (N10015, N10010, N596);
nor NOR4 (N10016, N10011, N9281, N7101, N5807);
nand NAND4 (N10017, N9989, N891, N5120, N5006);
or OR4 (N10018, N10012, N6728, N6247, N3135);
and AND2 (N10019, N10014, N3310);
nor NOR3 (N10020, N10019, N2871, N1587);
and AND4 (N10021, N9997, N6641, N4033, N1257);
and AND3 (N10022, N10001, N567, N788);
and AND4 (N10023, N10015, N6885, N3940, N4547);
or OR2 (N10024, N10016, N1671);
nand NAND4 (N10025, N10020, N2308, N8917, N1260);
xor XOR2 (N10026, N10017, N6200);
and AND3 (N10027, N10024, N7756, N5690);
xor XOR2 (N10028, N9995, N1852);
buf BUF1 (N10029, N10027);
nor NOR4 (N10030, N10018, N131, N9655, N181);
and AND3 (N10031, N10023, N5675, N824);
buf BUF1 (N10032, N10026);
not NOT1 (N10033, N10013);
buf BUF1 (N10034, N10025);
nand NAND4 (N10035, N10028, N8896, N3809, N7597);
and AND2 (N10036, N10022, N4999);
xor XOR2 (N10037, N10033, N6356);
nor NOR3 (N10038, N10031, N3637, N4288);
nor NOR2 (N10039, N10038, N5673);
or OR4 (N10040, N10039, N8345, N7705, N5046);
and AND2 (N10041, N10032, N8006);
nor NOR3 (N10042, N10041, N9355, N3587);
nor NOR2 (N10043, N9992, N8808);
nand NAND2 (N10044, N10040, N7067);
nor NOR2 (N10045, N10021, N8669);
not NOT1 (N10046, N10044);
nor NOR3 (N10047, N10036, N4924, N9575);
xor XOR2 (N10048, N10045, N3273);
not NOT1 (N10049, N10029);
and AND3 (N10050, N10043, N8470, N677);
xor XOR2 (N10051, N10030, N5817);
nand NAND2 (N10052, N10050, N1183);
buf BUF1 (N10053, N10037);
not NOT1 (N10054, N10048);
or OR4 (N10055, N10054, N3504, N2933, N2193);
xor XOR2 (N10056, N10046, N294);
xor XOR2 (N10057, N10034, N3028);
nand NAND3 (N10058, N10047, N9226, N308);
xor XOR2 (N10059, N10051, N7655);
not NOT1 (N10060, N10055);
and AND4 (N10061, N10053, N6763, N6212, N9724);
and AND4 (N10062, N10042, N9495, N6759, N7928);
nor NOR2 (N10063, N10061, N9562);
xor XOR2 (N10064, N10059, N5639);
or OR4 (N10065, N10063, N4586, N1671, N7995);
and AND4 (N10066, N10052, N2772, N5675, N3973);
nand NAND3 (N10067, N10060, N7018, N6845);
not NOT1 (N10068, N10064);
or OR2 (N10069, N10067, N5520);
not NOT1 (N10070, N10069);
or OR2 (N10071, N10035, N2124);
or OR3 (N10072, N10068, N223, N3892);
not NOT1 (N10073, N10065);
nand NAND3 (N10074, N10073, N9959, N659);
nand NAND2 (N10075, N10062, N9186);
nand NAND4 (N10076, N10075, N7744, N4702, N2969);
xor XOR2 (N10077, N10056, N9113);
xor XOR2 (N10078, N10057, N7338);
buf BUF1 (N10079, N10058);
buf BUF1 (N10080, N10049);
and AND4 (N10081, N10070, N7083, N1723, N1365);
or OR4 (N10082, N10079, N8935, N3444, N9548);
and AND2 (N10083, N10074, N2440);
not NOT1 (N10084, N10083);
or OR2 (N10085, N10066, N6548);
xor XOR2 (N10086, N10082, N4102);
xor XOR2 (N10087, N10086, N128);
nand NAND2 (N10088, N10072, N4002);
nor NOR4 (N10089, N10078, N9818, N4937, N3802);
nand NAND2 (N10090, N10081, N2347);
nand NAND4 (N10091, N10085, N1129, N3925, N6870);
and AND3 (N10092, N10089, N2236, N6684);
buf BUF1 (N10093, N10090);
nand NAND2 (N10094, N10071, N351);
buf BUF1 (N10095, N10088);
not NOT1 (N10096, N10093);
buf BUF1 (N10097, N10077);
xor XOR2 (N10098, N10087, N2477);
nand NAND4 (N10099, N10094, N2513, N1358, N1302);
buf BUF1 (N10100, N10091);
nor NOR2 (N10101, N10099, N8571);
buf BUF1 (N10102, N10076);
not NOT1 (N10103, N10102);
nor NOR3 (N10104, N10084, N10057, N6723);
nand NAND2 (N10105, N10104, N8631);
nor NOR4 (N10106, N10098, N5631, N328, N3371);
buf BUF1 (N10107, N10080);
nor NOR2 (N10108, N10096, N3248);
or OR3 (N10109, N10095, N5223, N6648);
and AND4 (N10110, N10107, N10085, N6110, N8697);
nor NOR3 (N10111, N10097, N9312, N7028);
nor NOR2 (N10112, N10109, N4656);
buf BUF1 (N10113, N10110);
nor NOR2 (N10114, N10108, N3517);
or OR2 (N10115, N10101, N5158);
nor NOR2 (N10116, N10114, N1654);
nor NOR3 (N10117, N10100, N6030, N8283);
and AND3 (N10118, N10103, N5780, N6708);
buf BUF1 (N10119, N10112);
nor NOR2 (N10120, N10111, N8701);
not NOT1 (N10121, N10106);
buf BUF1 (N10122, N10092);
nand NAND2 (N10123, N10116, N7519);
or OR4 (N10124, N10123, N7126, N8898, N8588);
or OR4 (N10125, N10122, N547, N8343, N2975);
or OR3 (N10126, N10120, N738, N3201);
or OR3 (N10127, N10105, N6343, N230);
and AND3 (N10128, N10127, N5853, N8284);
buf BUF1 (N10129, N10113);
not NOT1 (N10130, N10125);
nor NOR4 (N10131, N10126, N2161, N3958, N3027);
or OR3 (N10132, N10121, N9587, N7528);
not NOT1 (N10133, N10119);
xor XOR2 (N10134, N10133, N3500);
nand NAND2 (N10135, N10129, N6746);
nand NAND2 (N10136, N10117, N3245);
and AND2 (N10137, N10124, N3070);
or OR3 (N10138, N10130, N4876, N1558);
nor NOR2 (N10139, N10138, N7417);
buf BUF1 (N10140, N10139);
nand NAND3 (N10141, N10140, N1920, N7418);
or OR2 (N10142, N10132, N652);
or OR2 (N10143, N10137, N639);
nand NAND3 (N10144, N10118, N8707, N3307);
xor XOR2 (N10145, N10115, N3224);
nor NOR3 (N10146, N10136, N585, N125);
xor XOR2 (N10147, N10144, N4745);
or OR4 (N10148, N10134, N9439, N4487, N9945);
buf BUF1 (N10149, N10143);
or OR3 (N10150, N10128, N6660, N1060);
nor NOR4 (N10151, N10146, N335, N9785, N4274);
xor XOR2 (N10152, N10151, N740);
xor XOR2 (N10153, N10142, N7376);
buf BUF1 (N10154, N10148);
nand NAND2 (N10155, N10154, N2375);
buf BUF1 (N10156, N10141);
not NOT1 (N10157, N10156);
buf BUF1 (N10158, N10152);
or OR3 (N10159, N10135, N3748, N9646);
nor NOR4 (N10160, N10155, N7721, N7581, N2819);
nand NAND3 (N10161, N10149, N9032, N8011);
buf BUF1 (N10162, N10147);
nand NAND4 (N10163, N10161, N3696, N6288, N4726);
nor NOR4 (N10164, N10150, N2293, N1025, N9868);
and AND2 (N10165, N10159, N1499);
or OR3 (N10166, N10153, N4820, N7828);
or OR2 (N10167, N10160, N174);
not NOT1 (N10168, N10167);
and AND2 (N10169, N10157, N2444);
or OR2 (N10170, N10164, N8838);
not NOT1 (N10171, N10145);
or OR2 (N10172, N10170, N948);
buf BUF1 (N10173, N10166);
not NOT1 (N10174, N10162);
or OR2 (N10175, N10173, N166);
and AND2 (N10176, N10168, N10160);
and AND2 (N10177, N10163, N6766);
xor XOR2 (N10178, N10171, N5309);
nor NOR2 (N10179, N10174, N6458);
and AND3 (N10180, N10177, N5851, N10006);
and AND2 (N10181, N10179, N5886);
nor NOR2 (N10182, N10165, N1957);
not NOT1 (N10183, N10158);
and AND2 (N10184, N10172, N6258);
and AND4 (N10185, N10178, N6911, N4491, N7684);
not NOT1 (N10186, N10131);
and AND3 (N10187, N10169, N11, N3836);
not NOT1 (N10188, N10183);
nor NOR2 (N10189, N10188, N6181);
not NOT1 (N10190, N10176);
and AND4 (N10191, N10186, N9086, N7842, N6828);
nor NOR4 (N10192, N10190, N7218, N9342, N859);
buf BUF1 (N10193, N10182);
or OR2 (N10194, N10185, N8824);
and AND3 (N10195, N10193, N2099, N2417);
xor XOR2 (N10196, N10180, N6377);
not NOT1 (N10197, N10187);
xor XOR2 (N10198, N10197, N7079);
nor NOR4 (N10199, N10194, N10026, N8095, N7804);
buf BUF1 (N10200, N10198);
nor NOR4 (N10201, N10195, N1753, N2552, N4850);
and AND2 (N10202, N10175, N7145);
xor XOR2 (N10203, N10181, N889);
nor NOR2 (N10204, N10189, N6620);
and AND2 (N10205, N10201, N9533);
not NOT1 (N10206, N10202);
or OR3 (N10207, N10196, N6587, N8278);
nor NOR2 (N10208, N10206, N7166);
nor NOR2 (N10209, N10208, N2029);
buf BUF1 (N10210, N10192);
buf BUF1 (N10211, N10200);
nor NOR4 (N10212, N10199, N4515, N3486, N7207);
xor XOR2 (N10213, N10210, N10202);
and AND2 (N10214, N10205, N1415);
nor NOR3 (N10215, N10211, N6892, N883);
xor XOR2 (N10216, N10213, N167);
or OR4 (N10217, N10204, N8346, N368, N9367);
nand NAND3 (N10218, N10207, N7867, N4054);
or OR3 (N10219, N10191, N4840, N10110);
nor NOR3 (N10220, N10219, N4572, N2712);
and AND3 (N10221, N10203, N9725, N1792);
nor NOR2 (N10222, N10214, N1149);
or OR3 (N10223, N10218, N4490, N1833);
and AND3 (N10224, N10215, N10212, N6885);
xor XOR2 (N10225, N7624, N533);
xor XOR2 (N10226, N10184, N5946);
nor NOR2 (N10227, N10224, N4111);
xor XOR2 (N10228, N10216, N4496);
buf BUF1 (N10229, N10228);
or OR4 (N10230, N10226, N2926, N3831, N4742);
and AND3 (N10231, N10217, N9625, N4533);
buf BUF1 (N10232, N10223);
buf BUF1 (N10233, N10229);
nor NOR3 (N10234, N10220, N644, N8060);
xor XOR2 (N10235, N10230, N4391);
or OR4 (N10236, N10209, N2658, N7493, N6951);
buf BUF1 (N10237, N10233);
and AND4 (N10238, N10231, N7788, N1833, N6160);
not NOT1 (N10239, N10234);
not NOT1 (N10240, N10239);
nor NOR4 (N10241, N10221, N1455, N6890, N2163);
xor XOR2 (N10242, N10225, N9487);
buf BUF1 (N10243, N10227);
buf BUF1 (N10244, N10237);
xor XOR2 (N10245, N10238, N4208);
not NOT1 (N10246, N10241);
not NOT1 (N10247, N10243);
not NOT1 (N10248, N10245);
nor NOR4 (N10249, N10247, N6456, N7937, N5296);
nor NOR2 (N10250, N10222, N4715);
nand NAND2 (N10251, N10232, N3607);
and AND3 (N10252, N10242, N5773, N1870);
not NOT1 (N10253, N10248);
buf BUF1 (N10254, N10235);
nand NAND2 (N10255, N10244, N8318);
nor NOR3 (N10256, N10252, N72, N9550);
nand NAND2 (N10257, N10250, N8864);
not NOT1 (N10258, N10255);
buf BUF1 (N10259, N10257);
nor NOR3 (N10260, N10253, N6086, N749);
or OR2 (N10261, N10240, N2284);
xor XOR2 (N10262, N10260, N4268);
and AND3 (N10263, N10261, N6629, N6836);
not NOT1 (N10264, N10256);
and AND4 (N10265, N10259, N1057, N6853, N361);
xor XOR2 (N10266, N10264, N5631);
xor XOR2 (N10267, N10263, N9089);
or OR2 (N10268, N10265, N7751);
xor XOR2 (N10269, N10258, N1697);
nor NOR2 (N10270, N10262, N1485);
nor NOR2 (N10271, N10236, N3979);
xor XOR2 (N10272, N10271, N2483);
and AND4 (N10273, N10266, N6416, N8974, N4553);
nand NAND2 (N10274, N10254, N6750);
buf BUF1 (N10275, N10274);
xor XOR2 (N10276, N10268, N2878);
and AND4 (N10277, N10246, N7235, N8585, N3120);
or OR2 (N10278, N10251, N2244);
not NOT1 (N10279, N10276);
not NOT1 (N10280, N10275);
and AND3 (N10281, N10277, N5733, N7184);
nand NAND2 (N10282, N10278, N8003);
or OR2 (N10283, N10273, N1069);
nand NAND2 (N10284, N10272, N3142);
not NOT1 (N10285, N10267);
buf BUF1 (N10286, N10269);
or OR3 (N10287, N10283, N1233, N5566);
not NOT1 (N10288, N10249);
and AND2 (N10289, N10286, N8044);
or OR4 (N10290, N10284, N3012, N797, N4615);
not NOT1 (N10291, N10290);
buf BUF1 (N10292, N10287);
nor NOR4 (N10293, N10288, N9494, N526, N3686);
not NOT1 (N10294, N10280);
nand NAND2 (N10295, N10292, N9218);
nor NOR4 (N10296, N10294, N4771, N7595, N9479);
or OR2 (N10297, N10285, N7386);
xor XOR2 (N10298, N10297, N7104);
or OR2 (N10299, N10289, N7633);
xor XOR2 (N10300, N10279, N1203);
buf BUF1 (N10301, N10270);
buf BUF1 (N10302, N10296);
and AND4 (N10303, N10293, N3442, N4144, N7208);
and AND4 (N10304, N10291, N7345, N717, N2569);
xor XOR2 (N10305, N10299, N4147);
and AND2 (N10306, N10295, N1373);
nor NOR4 (N10307, N10306, N5925, N3507, N514);
buf BUF1 (N10308, N10304);
nor NOR4 (N10309, N10300, N4552, N2604, N4773);
buf BUF1 (N10310, N10305);
and AND4 (N10311, N10309, N2251, N925, N3343);
nor NOR3 (N10312, N10311, N4611, N4167);
buf BUF1 (N10313, N10310);
not NOT1 (N10314, N10312);
or OR4 (N10315, N10313, N5764, N4994, N3917);
nor NOR4 (N10316, N10282, N4343, N529, N10084);
not NOT1 (N10317, N10281);
or OR4 (N10318, N10315, N3850, N5778, N582);
buf BUF1 (N10319, N10301);
buf BUF1 (N10320, N10314);
or OR2 (N10321, N10318, N7938);
nor NOR2 (N10322, N10308, N2084);
and AND3 (N10323, N10302, N9565, N7955);
nand NAND4 (N10324, N10317, N4911, N4517, N2);
or OR2 (N10325, N10321, N10075);
xor XOR2 (N10326, N10303, N10254);
and AND3 (N10327, N10323, N4379, N6524);
buf BUF1 (N10328, N10327);
and AND2 (N10329, N10322, N5914);
buf BUF1 (N10330, N10326);
and AND2 (N10331, N10319, N3622);
or OR2 (N10332, N10298, N1106);
or OR2 (N10333, N10332, N10067);
buf BUF1 (N10334, N10320);
buf BUF1 (N10335, N10325);
nand NAND2 (N10336, N10329, N7733);
or OR3 (N10337, N10316, N2116, N1550);
xor XOR2 (N10338, N10336, N9001);
nor NOR4 (N10339, N10333, N3766, N6451, N9428);
not NOT1 (N10340, N10338);
and AND4 (N10341, N10328, N7792, N1705, N3547);
buf BUF1 (N10342, N10337);
or OR3 (N10343, N10341, N9662, N5169);
not NOT1 (N10344, N10335);
not NOT1 (N10345, N10331);
buf BUF1 (N10346, N10330);
buf BUF1 (N10347, N10307);
buf BUF1 (N10348, N10324);
or OR3 (N10349, N10348, N7182, N5955);
nor NOR2 (N10350, N10334, N316);
buf BUF1 (N10351, N10340);
and AND2 (N10352, N10339, N9752);
nand NAND3 (N10353, N10352, N9292, N287);
buf BUF1 (N10354, N10350);
nor NOR4 (N10355, N10351, N5779, N7971, N3237);
xor XOR2 (N10356, N10345, N7365);
nor NOR2 (N10357, N10344, N9142);
and AND2 (N10358, N10347, N4981);
and AND3 (N10359, N10343, N9083, N803);
and AND4 (N10360, N10342, N8011, N6418, N10168);
xor XOR2 (N10361, N10357, N4711);
nand NAND3 (N10362, N10354, N6186, N6519);
buf BUF1 (N10363, N10358);
nand NAND4 (N10364, N10359, N8502, N6111, N6787);
or OR2 (N10365, N10349, N3004);
buf BUF1 (N10366, N10364);
or OR3 (N10367, N10363, N5048, N3100);
or OR2 (N10368, N10355, N1327);
not NOT1 (N10369, N10365);
and AND2 (N10370, N10346, N7066);
buf BUF1 (N10371, N10370);
or OR4 (N10372, N10369, N9025, N3519, N8090);
and AND3 (N10373, N10362, N2997, N7699);
or OR4 (N10374, N10366, N4968, N7481, N6424);
or OR4 (N10375, N10372, N7813, N3480, N8719);
xor XOR2 (N10376, N10367, N8474);
nor NOR3 (N10377, N10373, N5039, N6145);
buf BUF1 (N10378, N10356);
or OR3 (N10379, N10377, N9618, N4252);
not NOT1 (N10380, N10374);
buf BUF1 (N10381, N10379);
not NOT1 (N10382, N10360);
or OR2 (N10383, N10368, N5088);
buf BUF1 (N10384, N10361);
buf BUF1 (N10385, N10384);
buf BUF1 (N10386, N10353);
not NOT1 (N10387, N10385);
xor XOR2 (N10388, N10381, N8960);
or OR4 (N10389, N10378, N2181, N5752, N2063);
nor NOR3 (N10390, N10371, N5991, N2160);
xor XOR2 (N10391, N10390, N8904);
buf BUF1 (N10392, N10376);
nor NOR2 (N10393, N10391, N5846);
not NOT1 (N10394, N10386);
nand NAND3 (N10395, N10389, N5601, N7865);
and AND4 (N10396, N10383, N4923, N7984, N1071);
or OR3 (N10397, N10382, N619, N7949);
or OR3 (N10398, N10395, N5768, N6743);
xor XOR2 (N10399, N10398, N2348);
nor NOR3 (N10400, N10375, N2540, N5207);
not NOT1 (N10401, N10397);
buf BUF1 (N10402, N10401);
or OR3 (N10403, N10396, N3231, N4272);
xor XOR2 (N10404, N10393, N7492);
not NOT1 (N10405, N10400);
buf BUF1 (N10406, N10404);
xor XOR2 (N10407, N10388, N3067);
and AND2 (N10408, N10380, N1352);
and AND4 (N10409, N10406, N10336, N989, N10242);
xor XOR2 (N10410, N10402, N9526);
not NOT1 (N10411, N10410);
buf BUF1 (N10412, N10387);
nor NOR2 (N10413, N10409, N7266);
xor XOR2 (N10414, N10394, N3509);
nand NAND4 (N10415, N10412, N8904, N1870, N2760);
nand NAND4 (N10416, N10415, N2626, N7270, N609);
buf BUF1 (N10417, N10403);
nand NAND2 (N10418, N10407, N2045);
and AND3 (N10419, N10405, N7807, N4741);
nor NOR2 (N10420, N10418, N8583);
not NOT1 (N10421, N10414);
and AND4 (N10422, N10417, N9214, N10238, N8070);
not NOT1 (N10423, N10399);
nand NAND4 (N10424, N10392, N7621, N4968, N257);
xor XOR2 (N10425, N10413, N3293);
buf BUF1 (N10426, N10421);
xor XOR2 (N10427, N10416, N686);
and AND4 (N10428, N10408, N5081, N4516, N5896);
xor XOR2 (N10429, N10428, N4066);
nor NOR2 (N10430, N10422, N692);
xor XOR2 (N10431, N10427, N9705);
xor XOR2 (N10432, N10431, N6437);
nor NOR4 (N10433, N10429, N1513, N4220, N3591);
xor XOR2 (N10434, N10425, N9310);
or OR2 (N10435, N10419, N5956);
or OR3 (N10436, N10433, N1347, N498);
not NOT1 (N10437, N10423);
or OR4 (N10438, N10426, N3708, N1781, N7514);
nand NAND4 (N10439, N10432, N9078, N2680, N4266);
buf BUF1 (N10440, N10430);
buf BUF1 (N10441, N10434);
buf BUF1 (N10442, N10441);
buf BUF1 (N10443, N10435);
buf BUF1 (N10444, N10420);
nor NOR3 (N10445, N10439, N4868, N2129);
not NOT1 (N10446, N10442);
nor NOR2 (N10447, N10411, N7406);
xor XOR2 (N10448, N10436, N963);
xor XOR2 (N10449, N10445, N4730);
xor XOR2 (N10450, N10440, N3269);
nand NAND3 (N10451, N10438, N5932, N9934);
nor NOR3 (N10452, N10444, N1490, N3952);
and AND4 (N10453, N10449, N3378, N2909, N4262);
or OR4 (N10454, N10450, N3636, N6164, N4651);
nor NOR3 (N10455, N10424, N5100, N9140);
or OR3 (N10456, N10453, N5673, N7430);
buf BUF1 (N10457, N10451);
nand NAND2 (N10458, N10443, N1240);
and AND4 (N10459, N10458, N3810, N8246, N4821);
and AND2 (N10460, N10446, N2479);
or OR2 (N10461, N10456, N7481);
not NOT1 (N10462, N10448);
nand NAND4 (N10463, N10460, N9880, N1356, N4940);
nand NAND3 (N10464, N10462, N5005, N5458);
nand NAND2 (N10465, N10447, N10199);
or OR3 (N10466, N10459, N4630, N8518);
buf BUF1 (N10467, N10454);
nand NAND2 (N10468, N10457, N2843);
nor NOR2 (N10469, N10452, N9891);
nand NAND2 (N10470, N10466, N3352);
and AND2 (N10471, N10463, N7502);
or OR2 (N10472, N10461, N1504);
and AND4 (N10473, N10455, N6505, N6990, N6833);
not NOT1 (N10474, N10472);
and AND2 (N10475, N10437, N3623);
buf BUF1 (N10476, N10464);
nand NAND4 (N10477, N10473, N4272, N6088, N4178);
nor NOR4 (N10478, N10468, N10187, N6343, N7513);
nor NOR2 (N10479, N10476, N162);
and AND2 (N10480, N10477, N1510);
or OR2 (N10481, N10467, N8050);
not NOT1 (N10482, N10469);
buf BUF1 (N10483, N10465);
buf BUF1 (N10484, N10471);
or OR4 (N10485, N10478, N7027, N5162, N1328);
not NOT1 (N10486, N10470);
or OR2 (N10487, N10480, N8998);
or OR4 (N10488, N10484, N6011, N952, N6115);
and AND2 (N10489, N10482, N9226);
xor XOR2 (N10490, N10483, N6313);
or OR3 (N10491, N10490, N2883, N4232);
or OR2 (N10492, N10475, N3723);
buf BUF1 (N10493, N10489);
buf BUF1 (N10494, N10481);
buf BUF1 (N10495, N10479);
xor XOR2 (N10496, N10494, N9514);
and AND3 (N10497, N10493, N4387, N1185);
nand NAND4 (N10498, N10492, N1080, N9994, N8947);
nor NOR4 (N10499, N10497, N2587, N8816, N2895);
not NOT1 (N10500, N10487);
not NOT1 (N10501, N10488);
or OR2 (N10502, N10500, N3759);
and AND3 (N10503, N10502, N6905, N8854);
and AND2 (N10504, N10474, N1627);
not NOT1 (N10505, N10496);
or OR3 (N10506, N10499, N3261, N9687);
nand NAND2 (N10507, N10486, N6789);
or OR2 (N10508, N10485, N9967);
or OR3 (N10509, N10503, N4072, N1716);
nor NOR4 (N10510, N10507, N6822, N9010, N2031);
nand NAND2 (N10511, N10509, N8433);
buf BUF1 (N10512, N10495);
nand NAND3 (N10513, N10505, N10197, N3841);
xor XOR2 (N10514, N10491, N10175);
buf BUF1 (N10515, N10513);
nand NAND4 (N10516, N10515, N7408, N8789, N1781);
not NOT1 (N10517, N10514);
nand NAND4 (N10518, N10498, N4520, N3130, N1043);
not NOT1 (N10519, N10512);
or OR4 (N10520, N10510, N8124, N502, N7191);
nor NOR4 (N10521, N10518, N907, N1577, N5695);
or OR4 (N10522, N10508, N6633, N4674, N8353);
not NOT1 (N10523, N10501);
nor NOR2 (N10524, N10516, N1241);
xor XOR2 (N10525, N10504, N4183);
not NOT1 (N10526, N10523);
and AND4 (N10527, N10525, N4605, N6181, N9533);
not NOT1 (N10528, N10526);
nor NOR3 (N10529, N10519, N5786, N9650);
buf BUF1 (N10530, N10511);
and AND3 (N10531, N10528, N9672, N9711);
or OR3 (N10532, N10522, N4774, N4604);
and AND3 (N10533, N10521, N9615, N9204);
nand NAND4 (N10534, N10524, N4306, N6256, N10123);
buf BUF1 (N10535, N10533);
nor NOR4 (N10536, N10535, N3386, N5889, N923);
not NOT1 (N10537, N10527);
or OR3 (N10538, N10531, N4517, N1536);
nand NAND2 (N10539, N10520, N5171);
nand NAND3 (N10540, N10529, N6696, N8679);
buf BUF1 (N10541, N10532);
nor NOR4 (N10542, N10517, N4025, N656, N2940);
nor NOR4 (N10543, N10537, N8649, N6599, N9789);
xor XOR2 (N10544, N10506, N8459);
or OR3 (N10545, N10543, N7557, N5781);
nor NOR2 (N10546, N10540, N2099);
and AND4 (N10547, N10544, N628, N1779, N305);
xor XOR2 (N10548, N10534, N7514);
and AND3 (N10549, N10545, N9473, N2696);
and AND2 (N10550, N10539, N1536);
xor XOR2 (N10551, N10550, N2423);
not NOT1 (N10552, N10551);
buf BUF1 (N10553, N10542);
not NOT1 (N10554, N10546);
or OR2 (N10555, N10541, N4521);
or OR4 (N10556, N10554, N8101, N1773, N2336);
xor XOR2 (N10557, N10530, N8443);
xor XOR2 (N10558, N10553, N4271);
or OR2 (N10559, N10549, N5354);
or OR4 (N10560, N10559, N1992, N9499, N6927);
nor NOR3 (N10561, N10536, N2731, N4745);
xor XOR2 (N10562, N10548, N7556);
nand NAND2 (N10563, N10557, N5383);
not NOT1 (N10564, N10560);
nand NAND2 (N10565, N10547, N6129);
buf BUF1 (N10566, N10564);
xor XOR2 (N10567, N10538, N6081);
not NOT1 (N10568, N10565);
not NOT1 (N10569, N10555);
nor NOR2 (N10570, N10562, N679);
xor XOR2 (N10571, N10569, N7513);
not NOT1 (N10572, N10568);
buf BUF1 (N10573, N10558);
not NOT1 (N10574, N10561);
and AND3 (N10575, N10573, N4177, N5652);
buf BUF1 (N10576, N10567);
nand NAND4 (N10577, N10571, N7615, N8202, N7957);
nor NOR3 (N10578, N10556, N2421, N5223);
nand NAND2 (N10579, N10572, N5671);
nor NOR3 (N10580, N10574, N8348, N7757);
nand NAND2 (N10581, N10566, N9182);
xor XOR2 (N10582, N10576, N8565);
not NOT1 (N10583, N10578);
xor XOR2 (N10584, N10552, N1011);
nor NOR3 (N10585, N10581, N7353, N6901);
or OR2 (N10586, N10582, N6440);
not NOT1 (N10587, N10563);
nor NOR2 (N10588, N10580, N3895);
not NOT1 (N10589, N10584);
buf BUF1 (N10590, N10575);
or OR3 (N10591, N10585, N491, N6806);
xor XOR2 (N10592, N10586, N6098);
or OR2 (N10593, N10589, N5389);
nor NOR4 (N10594, N10591, N5999, N4444, N8309);
nand NAND4 (N10595, N10590, N3192, N650, N6077);
buf BUF1 (N10596, N10577);
xor XOR2 (N10597, N10579, N7525);
and AND3 (N10598, N10595, N2621, N1957);
nand NAND3 (N10599, N10570, N1034, N7018);
and AND4 (N10600, N10598, N850, N5344, N207);
nand NAND2 (N10601, N10588, N7483);
nand NAND4 (N10602, N10600, N9553, N3126, N9435);
xor XOR2 (N10603, N10596, N6756);
nand NAND4 (N10604, N10603, N9967, N9503, N8739);
nor NOR3 (N10605, N10602, N2317, N3174);
and AND2 (N10606, N10599, N4294);
not NOT1 (N10607, N10587);
buf BUF1 (N10608, N10606);
and AND3 (N10609, N10605, N8559, N10371);
and AND4 (N10610, N10607, N8661, N9836, N1482);
buf BUF1 (N10611, N10597);
nand NAND2 (N10612, N10583, N6909);
nand NAND2 (N10613, N10612, N870);
xor XOR2 (N10614, N10609, N1645);
or OR4 (N10615, N10604, N1137, N7342, N1989);
xor XOR2 (N10616, N10610, N4408);
and AND4 (N10617, N10615, N8974, N8587, N263);
buf BUF1 (N10618, N10593);
buf BUF1 (N10619, N10608);
buf BUF1 (N10620, N10594);
nor NOR3 (N10621, N10617, N10570, N5235);
nor NOR3 (N10622, N10592, N5811, N9983);
buf BUF1 (N10623, N10620);
buf BUF1 (N10624, N10601);
not NOT1 (N10625, N10613);
not NOT1 (N10626, N10624);
not NOT1 (N10627, N10611);
and AND3 (N10628, N10619, N6012, N6796);
or OR3 (N10629, N10627, N7709, N426);
xor XOR2 (N10630, N10618, N5816);
or OR3 (N10631, N10616, N8865, N7145);
not NOT1 (N10632, N10623);
nor NOR2 (N10633, N10628, N970);
nor NOR2 (N10634, N10631, N6806);
nand NAND4 (N10635, N10622, N7626, N4360, N3218);
buf BUF1 (N10636, N10635);
nor NOR3 (N10637, N10633, N2069, N5246);
buf BUF1 (N10638, N10621);
buf BUF1 (N10639, N10614);
buf BUF1 (N10640, N10630);
nor NOR4 (N10641, N10638, N3713, N4511, N29);
not NOT1 (N10642, N10641);
nand NAND2 (N10643, N10642, N6414);
nand NAND3 (N10644, N10639, N6662, N10199);
or OR3 (N10645, N10629, N5309, N1488);
buf BUF1 (N10646, N10626);
nor NOR2 (N10647, N10640, N9157);
buf BUF1 (N10648, N10645);
and AND3 (N10649, N10637, N10151, N964);
and AND2 (N10650, N10634, N2890);
and AND2 (N10651, N10647, N629);
buf BUF1 (N10652, N10650);
xor XOR2 (N10653, N10636, N1521);
xor XOR2 (N10654, N10625, N3477);
or OR3 (N10655, N10649, N2584, N1077);
or OR3 (N10656, N10648, N5818, N1071);
nand NAND3 (N10657, N10651, N6046, N7716);
xor XOR2 (N10658, N10646, N2828);
or OR2 (N10659, N10655, N6275);
nor NOR3 (N10660, N10654, N9166, N847);
not NOT1 (N10661, N10660);
nand NAND3 (N10662, N10652, N6382, N5659);
and AND4 (N10663, N10632, N364, N2968, N4285);
xor XOR2 (N10664, N10653, N7126);
nand NAND3 (N10665, N10664, N6191, N5965);
nor NOR4 (N10666, N10644, N4742, N3189, N3358);
and AND3 (N10667, N10656, N4479, N2519);
and AND4 (N10668, N10658, N10135, N6511, N4292);
xor XOR2 (N10669, N10643, N3970);
or OR2 (N10670, N10657, N3836);
and AND4 (N10671, N10666, N9768, N1147, N2645);
xor XOR2 (N10672, N10662, N10275);
or OR2 (N10673, N10671, N5257);
nor NOR2 (N10674, N10673, N6606);
and AND2 (N10675, N10674, N6127);
nor NOR2 (N10676, N10667, N4654);
or OR3 (N10677, N10675, N6035, N6576);
not NOT1 (N10678, N10669);
xor XOR2 (N10679, N10659, N10034);
nor NOR2 (N10680, N10678, N9167);
nand NAND2 (N10681, N10672, N5409);
nand NAND4 (N10682, N10663, N8483, N7126, N5963);
and AND4 (N10683, N10677, N6750, N8320, N2391);
or OR4 (N10684, N10681, N4181, N3010, N552);
nor NOR4 (N10685, N10680, N9865, N3621, N8830);
xor XOR2 (N10686, N10665, N2279);
or OR4 (N10687, N10676, N6782, N9118, N9816);
not NOT1 (N10688, N10661);
or OR2 (N10689, N10682, N39);
not NOT1 (N10690, N10683);
nor NOR4 (N10691, N10685, N9122, N10043, N4069);
nand NAND4 (N10692, N10684, N1726, N2113, N1283);
and AND4 (N10693, N10688, N9571, N1707, N9413);
xor XOR2 (N10694, N10690, N3497);
xor XOR2 (N10695, N10686, N7094);
or OR2 (N10696, N10687, N4644);
and AND4 (N10697, N10692, N6126, N2296, N1639);
nor NOR2 (N10698, N10691, N1976);
nand NAND2 (N10699, N10668, N286);
and AND2 (N10700, N10693, N9042);
or OR3 (N10701, N10696, N302, N1870);
nand NAND2 (N10702, N10701, N9321);
nand NAND4 (N10703, N10679, N117, N3902, N9067);
xor XOR2 (N10704, N10695, N10264);
buf BUF1 (N10705, N10694);
not NOT1 (N10706, N10700);
and AND4 (N10707, N10703, N6272, N9616, N7319);
not NOT1 (N10708, N10698);
buf BUF1 (N10709, N10670);
and AND3 (N10710, N10699, N898, N9179);
or OR4 (N10711, N10697, N1826, N2692, N1351);
and AND3 (N10712, N10709, N620, N1983);
or OR2 (N10713, N10704, N8987);
nor NOR3 (N10714, N10711, N5785, N3909);
not NOT1 (N10715, N10710);
not NOT1 (N10716, N10715);
nor NOR3 (N10717, N10689, N41, N7607);
or OR4 (N10718, N10713, N8901, N10257, N9994);
nand NAND4 (N10719, N10702, N10060, N2659, N10169);
xor XOR2 (N10720, N10705, N9445);
not NOT1 (N10721, N10708);
not NOT1 (N10722, N10707);
xor XOR2 (N10723, N10721, N3607);
not NOT1 (N10724, N10720);
or OR2 (N10725, N10719, N9580);
nand NAND4 (N10726, N10706, N7233, N5280, N4482);
xor XOR2 (N10727, N10722, N3744);
not NOT1 (N10728, N10726);
and AND2 (N10729, N10723, N2508);
buf BUF1 (N10730, N10724);
or OR2 (N10731, N10725, N4625);
nor NOR4 (N10732, N10714, N10382, N7480, N7960);
and AND3 (N10733, N10732, N10474, N5323);
buf BUF1 (N10734, N10733);
nand NAND2 (N10735, N10727, N8829);
nor NOR3 (N10736, N10716, N9475, N8480);
and AND3 (N10737, N10734, N1551, N1113);
nor NOR3 (N10738, N10735, N2147, N10388);
xor XOR2 (N10739, N10728, N2732);
nand NAND4 (N10740, N10717, N3598, N3225, N7311);
nand NAND3 (N10741, N10718, N5315, N10657);
nor NOR2 (N10742, N10729, N9922);
nor NOR4 (N10743, N10731, N306, N2685, N9685);
and AND2 (N10744, N10738, N10528);
xor XOR2 (N10745, N10743, N5687);
not NOT1 (N10746, N10742);
xor XOR2 (N10747, N10736, N564);
buf BUF1 (N10748, N10746);
xor XOR2 (N10749, N10712, N7110);
buf BUF1 (N10750, N10737);
and AND3 (N10751, N10740, N8500, N1754);
or OR2 (N10752, N10748, N245);
nand NAND3 (N10753, N10751, N1941, N829);
buf BUF1 (N10754, N10752);
xor XOR2 (N10755, N10745, N9402);
or OR2 (N10756, N10754, N8486);
and AND4 (N10757, N10753, N3753, N4625, N8150);
and AND3 (N10758, N10757, N5063, N973);
and AND2 (N10759, N10750, N2782);
or OR4 (N10760, N10741, N4124, N7965, N6620);
buf BUF1 (N10761, N10739);
not NOT1 (N10762, N10756);
nor NOR3 (N10763, N10747, N6309, N3927);
and AND4 (N10764, N10760, N10312, N10507, N6618);
not NOT1 (N10765, N10762);
nand NAND3 (N10766, N10744, N5970, N9567);
xor XOR2 (N10767, N10761, N4224);
and AND4 (N10768, N10730, N3157, N4949, N5563);
and AND2 (N10769, N10749, N3560);
or OR2 (N10770, N10755, N4533);
nor NOR4 (N10771, N10766, N7721, N2902, N9358);
or OR2 (N10772, N10768, N3722);
or OR2 (N10773, N10758, N6944);
and AND3 (N10774, N10764, N10472, N2861);
and AND2 (N10775, N10769, N254);
nand NAND4 (N10776, N10773, N7116, N278, N6900);
and AND3 (N10777, N10767, N5798, N3758);
and AND2 (N10778, N10770, N3424);
and AND4 (N10779, N10778, N647, N3118, N7144);
buf BUF1 (N10780, N10779);
nand NAND3 (N10781, N10774, N5736, N7570);
buf BUF1 (N10782, N10763);
nor NOR2 (N10783, N10782, N2121);
buf BUF1 (N10784, N10772);
and AND2 (N10785, N10783, N778);
xor XOR2 (N10786, N10785, N9398);
not NOT1 (N10787, N10771);
and AND3 (N10788, N10765, N4525, N6150);
or OR4 (N10789, N10781, N7588, N9404, N1132);
or OR2 (N10790, N10759, N8910);
xor XOR2 (N10791, N10780, N3601);
xor XOR2 (N10792, N10791, N5945);
and AND4 (N10793, N10775, N5555, N5681, N9673);
and AND2 (N10794, N10789, N9190);
buf BUF1 (N10795, N10786);
and AND2 (N10796, N10794, N1534);
and AND2 (N10797, N10792, N9511);
buf BUF1 (N10798, N10776);
xor XOR2 (N10799, N10798, N312);
xor XOR2 (N10800, N10795, N1023);
nor NOR4 (N10801, N10797, N1248, N9975, N10313);
nor NOR2 (N10802, N10784, N5207);
and AND4 (N10803, N10787, N5018, N488, N7764);
and AND2 (N10804, N10793, N3460);
nand NAND2 (N10805, N10790, N1299);
or OR4 (N10806, N10800, N8709, N4221, N6963);
xor XOR2 (N10807, N10788, N10610);
buf BUF1 (N10808, N10805);
nor NOR4 (N10809, N10807, N8083, N6773, N8097);
or OR3 (N10810, N10809, N6338, N10557);
and AND4 (N10811, N10806, N4181, N8075, N8305);
or OR3 (N10812, N10808, N4430, N8022);
buf BUF1 (N10813, N10802);
xor XOR2 (N10814, N10796, N7874);
or OR4 (N10815, N10803, N8679, N6068, N5929);
not NOT1 (N10816, N10777);
and AND2 (N10817, N10801, N7248);
or OR4 (N10818, N10804, N10553, N9056, N8610);
and AND2 (N10819, N10799, N7875);
xor XOR2 (N10820, N10815, N1683);
and AND2 (N10821, N10816, N537);
not NOT1 (N10822, N10813);
or OR2 (N10823, N10819, N8577);
nand NAND4 (N10824, N10821, N1015, N2381, N6390);
and AND3 (N10825, N10814, N3987, N3426);
xor XOR2 (N10826, N10823, N9269);
buf BUF1 (N10827, N10826);
not NOT1 (N10828, N10811);
not NOT1 (N10829, N10812);
nand NAND3 (N10830, N10825, N8154, N10704);
or OR4 (N10831, N10822, N10615, N3691, N9653);
or OR4 (N10832, N10810, N9352, N3511, N5394);
not NOT1 (N10833, N10830);
or OR4 (N10834, N10833, N6260, N2061, N8092);
xor XOR2 (N10835, N10824, N9666);
not NOT1 (N10836, N10817);
nand NAND2 (N10837, N10829, N3429);
not NOT1 (N10838, N10837);
nor NOR2 (N10839, N10834, N1250);
nand NAND2 (N10840, N10838, N3374);
buf BUF1 (N10841, N10836);
nor NOR4 (N10842, N10820, N347, N5369, N5358);
nand NAND3 (N10843, N10841, N6827, N892);
buf BUF1 (N10844, N10840);
buf BUF1 (N10845, N10827);
buf BUF1 (N10846, N10839);
or OR3 (N10847, N10835, N8443, N4672);
buf BUF1 (N10848, N10832);
not NOT1 (N10849, N10828);
buf BUF1 (N10850, N10842);
nor NOR4 (N10851, N10831, N6111, N3417, N10268);
or OR3 (N10852, N10818, N3737, N4934);
nand NAND3 (N10853, N10844, N3089, N1932);
or OR3 (N10854, N10853, N2040, N3659);
or OR4 (N10855, N10848, N5995, N414, N7284);
buf BUF1 (N10856, N10855);
and AND4 (N10857, N10854, N3944, N599, N7661);
nand NAND3 (N10858, N10849, N5409, N8674);
buf BUF1 (N10859, N10851);
or OR3 (N10860, N10850, N4190, N703);
and AND3 (N10861, N10847, N3943, N9344);
not NOT1 (N10862, N10857);
and AND2 (N10863, N10858, N8588);
not NOT1 (N10864, N10863);
nor NOR2 (N10865, N10846, N7465);
xor XOR2 (N10866, N10861, N9460);
or OR4 (N10867, N10845, N3720, N5813, N3225);
xor XOR2 (N10868, N10859, N2456);
xor XOR2 (N10869, N10864, N3082);
nor NOR3 (N10870, N10869, N6374, N4261);
xor XOR2 (N10871, N10843, N5862);
and AND2 (N10872, N10862, N2947);
buf BUF1 (N10873, N10866);
nor NOR4 (N10874, N10860, N2696, N8153, N6779);
not NOT1 (N10875, N10865);
or OR3 (N10876, N10856, N9547, N5880);
buf BUF1 (N10877, N10876);
buf BUF1 (N10878, N10874);
xor XOR2 (N10879, N10852, N4400);
nand NAND3 (N10880, N10871, N9662, N2568);
nor NOR2 (N10881, N10877, N4442);
or OR4 (N10882, N10875, N5177, N1468, N7096);
xor XOR2 (N10883, N10868, N1915);
xor XOR2 (N10884, N10873, N6539);
or OR2 (N10885, N10879, N2177);
nor NOR2 (N10886, N10872, N258);
nor NOR2 (N10887, N10880, N1927);
or OR4 (N10888, N10885, N6857, N3944, N2694);
or OR3 (N10889, N10883, N6641, N9313);
not NOT1 (N10890, N10878);
xor XOR2 (N10891, N10884, N6886);
not NOT1 (N10892, N10886);
buf BUF1 (N10893, N10892);
xor XOR2 (N10894, N10889, N10223);
nor NOR2 (N10895, N10887, N2497);
or OR3 (N10896, N10894, N4052, N9109);
and AND2 (N10897, N10890, N9504);
or OR4 (N10898, N10882, N5489, N6238, N5530);
and AND2 (N10899, N10870, N8009);
not NOT1 (N10900, N10897);
xor XOR2 (N10901, N10888, N4606);
nor NOR4 (N10902, N10901, N1685, N5158, N3196);
or OR2 (N10903, N10891, N7189);
xor XOR2 (N10904, N10881, N9880);
and AND3 (N10905, N10904, N4713, N4193);
buf BUF1 (N10906, N10898);
xor XOR2 (N10907, N10903, N4436);
and AND2 (N10908, N10896, N6356);
xor XOR2 (N10909, N10902, N1389);
not NOT1 (N10910, N10909);
nand NAND2 (N10911, N10900, N8856);
xor XOR2 (N10912, N10907, N8421);
buf BUF1 (N10913, N10906);
or OR3 (N10914, N10910, N10111, N5717);
or OR2 (N10915, N10899, N2617);
buf BUF1 (N10916, N10895);
not NOT1 (N10917, N10893);
nand NAND2 (N10918, N10905, N7571);
not NOT1 (N10919, N10867);
nand NAND3 (N10920, N10916, N8541, N4839);
nor NOR4 (N10921, N10914, N4158, N1862, N4037);
buf BUF1 (N10922, N10913);
nand NAND4 (N10923, N10915, N6764, N1823, N3122);
xor XOR2 (N10924, N10921, N3155);
xor XOR2 (N10925, N10918, N2179);
nor NOR3 (N10926, N10922, N9998, N6009);
nor NOR3 (N10927, N10925, N7668, N5488);
and AND3 (N10928, N10912, N7026, N3908);
xor XOR2 (N10929, N10923, N3127);
or OR4 (N10930, N10929, N3558, N6146, N8124);
or OR4 (N10931, N10908, N1864, N313, N1832);
or OR2 (N10932, N10927, N8697);
nor NOR3 (N10933, N10911, N2459, N4211);
and AND4 (N10934, N10931, N9614, N2307, N8045);
not NOT1 (N10935, N10934);
or OR3 (N10936, N10933, N1021, N1582);
nand NAND4 (N10937, N10935, N9502, N2317, N10882);
buf BUF1 (N10938, N10919);
nand NAND3 (N10939, N10932, N710, N124);
xor XOR2 (N10940, N10924, N1068);
or OR3 (N10941, N10937, N5607, N1332);
nand NAND4 (N10942, N10926, N6984, N134, N4606);
or OR3 (N10943, N10940, N2701, N7777);
or OR2 (N10944, N10917, N3541);
nand NAND4 (N10945, N10941, N5610, N8347, N7984);
and AND3 (N10946, N10938, N3587, N3261);
nand NAND4 (N10947, N10930, N1980, N1941, N6177);
or OR2 (N10948, N10947, N6337);
nand NAND3 (N10949, N10936, N826, N1761);
xor XOR2 (N10950, N10948, N5572);
nor NOR2 (N10951, N10950, N366);
buf BUF1 (N10952, N10951);
xor XOR2 (N10953, N10945, N5228);
nor NOR3 (N10954, N10928, N8558, N4511);
nand NAND4 (N10955, N10944, N6883, N10809, N8246);
or OR2 (N10956, N10953, N2053);
and AND4 (N10957, N10920, N8393, N8314, N6652);
and AND3 (N10958, N10949, N5974, N4270);
xor XOR2 (N10959, N10946, N7950);
xor XOR2 (N10960, N10939, N250);
xor XOR2 (N10961, N10955, N8842);
buf BUF1 (N10962, N10961);
nor NOR4 (N10963, N10942, N3600, N3765, N2990);
not NOT1 (N10964, N10943);
not NOT1 (N10965, N10964);
xor XOR2 (N10966, N10959, N5392);
nor NOR3 (N10967, N10963, N3545, N10871);
nor NOR3 (N10968, N10966, N3236, N8278);
and AND2 (N10969, N10957, N8406);
not NOT1 (N10970, N10968);
not NOT1 (N10971, N10965);
or OR4 (N10972, N10960, N639, N6475, N6030);
nor NOR3 (N10973, N10952, N3363, N6961);
and AND3 (N10974, N10969, N7236, N10832);
buf BUF1 (N10975, N10972);
nor NOR2 (N10976, N10973, N6216);
xor XOR2 (N10977, N10971, N10437);
buf BUF1 (N10978, N10975);
nand NAND4 (N10979, N10962, N5838, N1515, N5489);
and AND4 (N10980, N10970, N5700, N4123, N5430);
not NOT1 (N10981, N10978);
and AND2 (N10982, N10974, N2095);
not NOT1 (N10983, N10976);
nor NOR2 (N10984, N10980, N1618);
not NOT1 (N10985, N10984);
and AND4 (N10986, N10979, N7142, N3179, N8789);
not NOT1 (N10987, N10981);
buf BUF1 (N10988, N10986);
nor NOR3 (N10989, N10985, N965, N10436);
nor NOR4 (N10990, N10954, N7525, N4928, N1431);
and AND3 (N10991, N10982, N8299, N6472);
buf BUF1 (N10992, N10991);
or OR4 (N10993, N10992, N10310, N9612, N31);
nor NOR3 (N10994, N10956, N5366, N10686);
xor XOR2 (N10995, N10990, N2996);
xor XOR2 (N10996, N10967, N2879);
buf BUF1 (N10997, N10977);
or OR3 (N10998, N10989, N3731, N8210);
nor NOR4 (N10999, N10997, N9550, N3211, N6553);
xor XOR2 (N11000, N10999, N8029);
not NOT1 (N11001, N10996);
nand NAND2 (N11002, N10987, N9411);
not NOT1 (N11003, N10998);
or OR2 (N11004, N10995, N10406);
and AND2 (N11005, N11003, N9886);
nand NAND3 (N11006, N11005, N4452, N6159);
buf BUF1 (N11007, N10958);
and AND3 (N11008, N10988, N5353, N9022);
nor NOR4 (N11009, N11006, N9728, N5339, N191);
or OR3 (N11010, N11004, N3371, N10823);
nand NAND4 (N11011, N11000, N457, N4061, N8351);
buf BUF1 (N11012, N10983);
nor NOR2 (N11013, N11002, N8807);
nand NAND4 (N11014, N11008, N1114, N6063, N7794);
nand NAND2 (N11015, N11011, N8916);
and AND2 (N11016, N10993, N2689);
buf BUF1 (N11017, N11014);
buf BUF1 (N11018, N11009);
xor XOR2 (N11019, N11013, N777);
xor XOR2 (N11020, N11012, N10058);
buf BUF1 (N11021, N11018);
xor XOR2 (N11022, N11007, N947);
xor XOR2 (N11023, N11001, N826);
xor XOR2 (N11024, N11015, N9649);
and AND2 (N11025, N11019, N9250);
nand NAND3 (N11026, N11023, N4960, N3530);
nand NAND4 (N11027, N11024, N2336, N1329, N1596);
nand NAND4 (N11028, N11020, N133, N10100, N9726);
buf BUF1 (N11029, N11026);
xor XOR2 (N11030, N11027, N5062);
or OR2 (N11031, N11010, N10709);
and AND2 (N11032, N11030, N3745);
nor NOR2 (N11033, N11025, N7796);
and AND4 (N11034, N11032, N6278, N3828, N4524);
buf BUF1 (N11035, N11017);
xor XOR2 (N11036, N11033, N5958);
xor XOR2 (N11037, N11021, N8881);
xor XOR2 (N11038, N11022, N4500);
xor XOR2 (N11039, N11034, N2254);
or OR2 (N11040, N11035, N6688);
not NOT1 (N11041, N11036);
nand NAND4 (N11042, N10994, N2961, N6466, N8192);
nand NAND2 (N11043, N11039, N4957);
or OR3 (N11044, N11029, N1073, N798);
nand NAND2 (N11045, N11031, N6737);
or OR2 (N11046, N11028, N868);
or OR2 (N11047, N11016, N11017);
not NOT1 (N11048, N11044);
or OR2 (N11049, N11038, N1);
and AND2 (N11050, N11041, N1369);
buf BUF1 (N11051, N11037);
and AND3 (N11052, N11040, N9597, N4942);
xor XOR2 (N11053, N11049, N2944);
xor XOR2 (N11054, N11050, N1591);
nand NAND4 (N11055, N11046, N3780, N3973, N9144);
nor NOR3 (N11056, N11048, N9568, N2098);
buf BUF1 (N11057, N11056);
buf BUF1 (N11058, N11042);
nor NOR3 (N11059, N11045, N7830, N5927);
or OR3 (N11060, N11057, N7474, N2100);
and AND2 (N11061, N11059, N698);
or OR4 (N11062, N11051, N5937, N6122, N4652);
not NOT1 (N11063, N11053);
nand NAND3 (N11064, N11043, N6788, N10500);
nor NOR2 (N11065, N11058, N8631);
buf BUF1 (N11066, N11060);
nand NAND3 (N11067, N11054, N10398, N5992);
or OR3 (N11068, N11064, N2782, N1542);
xor XOR2 (N11069, N11068, N9292);
nor NOR3 (N11070, N11065, N10550, N3966);
nand NAND2 (N11071, N11047, N8027);
and AND3 (N11072, N11062, N6927, N10515);
not NOT1 (N11073, N11071);
buf BUF1 (N11074, N11066);
nand NAND4 (N11075, N11074, N6133, N10569, N10398);
nor NOR4 (N11076, N11055, N7854, N10935, N6522);
xor XOR2 (N11077, N11067, N2154);
or OR2 (N11078, N11069, N3464);
nor NOR3 (N11079, N11078, N1938, N5866);
buf BUF1 (N11080, N11070);
not NOT1 (N11081, N11076);
not NOT1 (N11082, N11079);
nor NOR3 (N11083, N11075, N4020, N2578);
xor XOR2 (N11084, N11063, N6581);
nand NAND2 (N11085, N11052, N7461);
nand NAND4 (N11086, N11082, N3513, N627, N6468);
nor NOR3 (N11087, N11061, N9321, N10654);
buf BUF1 (N11088, N11073);
xor XOR2 (N11089, N11088, N4036);
or OR2 (N11090, N11081, N6327);
xor XOR2 (N11091, N11083, N4752);
or OR3 (N11092, N11085, N4591, N690);
and AND2 (N11093, N11087, N10907);
not NOT1 (N11094, N11077);
nor NOR3 (N11095, N11084, N3307, N9565);
xor XOR2 (N11096, N11094, N10688);
buf BUF1 (N11097, N11080);
or OR2 (N11098, N11091, N5625);
not NOT1 (N11099, N11096);
not NOT1 (N11100, N11092);
xor XOR2 (N11101, N11099, N6263);
nand NAND4 (N11102, N11090, N794, N378, N8854);
nand NAND3 (N11103, N11101, N7924, N5207);
nor NOR3 (N11104, N11102, N8581, N7396);
nor NOR2 (N11105, N11086, N4687);
or OR4 (N11106, N11095, N5331, N2813, N2027);
nor NOR3 (N11107, N11097, N8644, N9271);
or OR2 (N11108, N11103, N4104);
and AND3 (N11109, N11107, N3809, N923);
or OR4 (N11110, N11100, N3434, N6968, N3215);
buf BUF1 (N11111, N11106);
nand NAND3 (N11112, N11093, N8146, N5816);
nand NAND4 (N11113, N11110, N9671, N501, N9962);
or OR3 (N11114, N11105, N7994, N8135);
buf BUF1 (N11115, N11072);
or OR4 (N11116, N11108, N6247, N9736, N6043);
not NOT1 (N11117, N11113);
nand NAND3 (N11118, N11115, N10463, N7877);
and AND4 (N11119, N11116, N3382, N5618, N1467);
nor NOR2 (N11120, N11111, N7659);
not NOT1 (N11121, N11112);
nor NOR3 (N11122, N11109, N6495, N5930);
buf BUF1 (N11123, N11089);
nor NOR3 (N11124, N11119, N10113, N7349);
nand NAND4 (N11125, N11123, N10598, N8170, N4208);
buf BUF1 (N11126, N11117);
nor NOR4 (N11127, N11122, N3991, N6960, N7103);
not NOT1 (N11128, N11114);
not NOT1 (N11129, N11128);
or OR2 (N11130, N11125, N8072);
buf BUF1 (N11131, N11118);
buf BUF1 (N11132, N11130);
buf BUF1 (N11133, N11126);
or OR2 (N11134, N11131, N6876);
xor XOR2 (N11135, N11132, N7804);
nor NOR4 (N11136, N11134, N1179, N6786, N5373);
or OR2 (N11137, N11129, N2511);
not NOT1 (N11138, N11127);
xor XOR2 (N11139, N11135, N999);
not NOT1 (N11140, N11137);
nand NAND2 (N11141, N11139, N8540);
xor XOR2 (N11142, N11138, N9136);
xor XOR2 (N11143, N11140, N596);
or OR3 (N11144, N11098, N7165, N2140);
nand NAND3 (N11145, N11121, N2749, N7129);
xor XOR2 (N11146, N11124, N1611);
nand NAND3 (N11147, N11136, N1729, N2653);
buf BUF1 (N11148, N11147);
not NOT1 (N11149, N11144);
nand NAND3 (N11150, N11146, N4679, N3649);
nor NOR4 (N11151, N11149, N10729, N760, N5037);
or OR2 (N11152, N11145, N2748);
or OR3 (N11153, N11150, N7518, N5959);
nor NOR2 (N11154, N11151, N10825);
not NOT1 (N11155, N11148);
not NOT1 (N11156, N11155);
xor XOR2 (N11157, N11153, N8363);
or OR4 (N11158, N11152, N4870, N2967, N5016);
buf BUF1 (N11159, N11133);
nor NOR3 (N11160, N11159, N3511, N6963);
nand NAND4 (N11161, N11154, N8202, N5585, N9836);
or OR3 (N11162, N11143, N3291, N11108);
nor NOR2 (N11163, N11104, N9614);
nor NOR3 (N11164, N11163, N6029, N5370);
and AND4 (N11165, N11156, N3771, N10470, N3639);
or OR2 (N11166, N11141, N1384);
nand NAND4 (N11167, N11165, N5366, N1701, N1644);
buf BUF1 (N11168, N11120);
nor NOR4 (N11169, N11164, N10861, N7331, N9311);
xor XOR2 (N11170, N11157, N7528);
and AND2 (N11171, N11170, N7727);
buf BUF1 (N11172, N11161);
not NOT1 (N11173, N11168);
not NOT1 (N11174, N11167);
and AND2 (N11175, N11142, N4433);
nor NOR3 (N11176, N11173, N3109, N507);
not NOT1 (N11177, N11174);
nand NAND3 (N11178, N11177, N4109, N1888);
nand NAND3 (N11179, N11162, N3137, N1538);
xor XOR2 (N11180, N11166, N2576);
buf BUF1 (N11181, N11175);
nand NAND2 (N11182, N11160, N5660);
buf BUF1 (N11183, N11182);
nor NOR3 (N11184, N11183, N7810, N5139);
buf BUF1 (N11185, N11172);
not NOT1 (N11186, N11176);
and AND3 (N11187, N11185, N9903, N4541);
not NOT1 (N11188, N11171);
and AND2 (N11189, N11188, N7010);
nand NAND2 (N11190, N11184, N1286);
not NOT1 (N11191, N11180);
nand NAND3 (N11192, N11187, N3983, N1167);
nor NOR3 (N11193, N11186, N2397, N3397);
nor NOR4 (N11194, N11192, N2304, N9378, N4160);
nor NOR2 (N11195, N11178, N9087);
buf BUF1 (N11196, N11193);
buf BUF1 (N11197, N11194);
or OR2 (N11198, N11181, N2871);
or OR3 (N11199, N11189, N5925, N3097);
nand NAND3 (N11200, N11197, N9089, N1547);
buf BUF1 (N11201, N11199);
nand NAND3 (N11202, N11190, N1322, N6659);
nand NAND3 (N11203, N11191, N4040, N9961);
buf BUF1 (N11204, N11196);
buf BUF1 (N11205, N11158);
nor NOR3 (N11206, N11205, N8768, N9285);
nand NAND3 (N11207, N11198, N7432, N637);
nor NOR4 (N11208, N11206, N3777, N259, N3619);
not NOT1 (N11209, N11204);
xor XOR2 (N11210, N11207, N4136);
or OR4 (N11211, N11209, N6645, N6860, N2284);
nand NAND4 (N11212, N11195, N2109, N2058, N7637);
buf BUF1 (N11213, N11202);
xor XOR2 (N11214, N11208, N3193);
and AND2 (N11215, N11200, N2626);
buf BUF1 (N11216, N11211);
and AND4 (N11217, N11203, N491, N1769, N1249);
nor NOR2 (N11218, N11213, N2944);
nor NOR4 (N11219, N11218, N7363, N7815, N2451);
not NOT1 (N11220, N11210);
or OR2 (N11221, N11215, N2563);
xor XOR2 (N11222, N11214, N987);
nand NAND4 (N11223, N11221, N2416, N3825, N6615);
not NOT1 (N11224, N11222);
not NOT1 (N11225, N11219);
and AND3 (N11226, N11216, N7522, N6024);
nor NOR4 (N11227, N11169, N9489, N9231, N5661);
xor XOR2 (N11228, N11212, N786);
not NOT1 (N11229, N11179);
not NOT1 (N11230, N11217);
and AND2 (N11231, N11229, N4383);
xor XOR2 (N11232, N11230, N4527);
buf BUF1 (N11233, N11228);
nor NOR4 (N11234, N11231, N11212, N3380, N6623);
and AND3 (N11235, N11225, N3450, N6015);
not NOT1 (N11236, N11227);
or OR3 (N11237, N11235, N2469, N1428);
and AND2 (N11238, N11233, N8503);
or OR4 (N11239, N11224, N10570, N362, N10812);
xor XOR2 (N11240, N11232, N8731);
nand NAND2 (N11241, N11237, N2010);
and AND3 (N11242, N11241, N9571, N4886);
nand NAND2 (N11243, N11220, N592);
nand NAND4 (N11244, N11234, N8022, N3162, N8260);
buf BUF1 (N11245, N11242);
nor NOR3 (N11246, N11245, N6461, N3488);
buf BUF1 (N11247, N11243);
nand NAND2 (N11248, N11247, N7760);
nor NOR2 (N11249, N11244, N10481);
nand NAND4 (N11250, N11240, N606, N10918, N5442);
and AND4 (N11251, N11239, N2901, N6058, N7606);
buf BUF1 (N11252, N11248);
and AND4 (N11253, N11201, N8076, N2949, N4034);
xor XOR2 (N11254, N11246, N11072);
and AND3 (N11255, N11253, N3564, N5959);
xor XOR2 (N11256, N11250, N5541);
not NOT1 (N11257, N11254);
or OR4 (N11258, N11238, N810, N10612, N6222);
buf BUF1 (N11259, N11236);
nor NOR3 (N11260, N11258, N4156, N9648);
xor XOR2 (N11261, N11251, N249);
nand NAND3 (N11262, N11261, N6073, N277);
nor NOR4 (N11263, N11223, N3533, N8271, N8696);
xor XOR2 (N11264, N11256, N6712);
not NOT1 (N11265, N11249);
buf BUF1 (N11266, N11257);
or OR3 (N11267, N11265, N1467, N7034);
xor XOR2 (N11268, N11264, N3032);
not NOT1 (N11269, N11262);
not NOT1 (N11270, N11260);
or OR2 (N11271, N11259, N4396);
nand NAND2 (N11272, N11267, N5273);
and AND2 (N11273, N11266, N3703);
or OR3 (N11274, N11272, N994, N7646);
nand NAND4 (N11275, N11271, N2759, N10979, N10908);
or OR4 (N11276, N11226, N9287, N520, N7976);
nor NOR4 (N11277, N11270, N6970, N4154, N7826);
not NOT1 (N11278, N11277);
nand NAND4 (N11279, N11263, N10925, N7992, N3979);
xor XOR2 (N11280, N11268, N4403);
nand NAND3 (N11281, N11279, N6183, N7181);
or OR4 (N11282, N11252, N2985, N2624, N9599);
nor NOR3 (N11283, N11269, N3841, N4194);
or OR4 (N11284, N11275, N9517, N8329, N627);
not NOT1 (N11285, N11274);
not NOT1 (N11286, N11255);
or OR3 (N11287, N11281, N10901, N3197);
nand NAND4 (N11288, N11286, N2786, N482, N3477);
xor XOR2 (N11289, N11288, N9048);
nand NAND4 (N11290, N11276, N2500, N5455, N6984);
not NOT1 (N11291, N11285);
nand NAND3 (N11292, N11290, N5419, N8778);
xor XOR2 (N11293, N11280, N3883);
xor XOR2 (N11294, N11284, N5599);
xor XOR2 (N11295, N11291, N6336);
and AND2 (N11296, N11293, N3431);
and AND3 (N11297, N11282, N1461, N5322);
nor NOR2 (N11298, N11297, N6591);
nor NOR3 (N11299, N11294, N2517, N8551);
buf BUF1 (N11300, N11273);
or OR3 (N11301, N11300, N4777, N5625);
and AND4 (N11302, N11301, N505, N8446, N1152);
xor XOR2 (N11303, N11292, N3856);
not NOT1 (N11304, N11303);
buf BUF1 (N11305, N11298);
nor NOR4 (N11306, N11295, N4950, N10424, N10999);
not NOT1 (N11307, N11299);
nor NOR3 (N11308, N11283, N6956, N959);
nand NAND3 (N11309, N11305, N3286, N4936);
or OR4 (N11310, N11306, N6062, N8661, N1664);
and AND3 (N11311, N11296, N9684, N2035);
nor NOR4 (N11312, N11308, N2515, N1055, N6898);
xor XOR2 (N11313, N11287, N9010);
and AND4 (N11314, N11310, N750, N3525, N220);
not NOT1 (N11315, N11311);
nand NAND2 (N11316, N11302, N6274);
nor NOR4 (N11317, N11309, N6595, N3146, N6838);
xor XOR2 (N11318, N11312, N176);
buf BUF1 (N11319, N11316);
not NOT1 (N11320, N11278);
nand NAND4 (N11321, N11319, N988, N2023, N6512);
and AND2 (N11322, N11320, N3818);
xor XOR2 (N11323, N11321, N4429);
not NOT1 (N11324, N11307);
nand NAND4 (N11325, N11314, N6432, N1632, N1006);
or OR4 (N11326, N11318, N2121, N10979, N9767);
and AND2 (N11327, N11322, N4866);
not NOT1 (N11328, N11327);
not NOT1 (N11329, N11313);
not NOT1 (N11330, N11289);
and AND2 (N11331, N11324, N654);
or OR2 (N11332, N11326, N3806);
xor XOR2 (N11333, N11304, N2403);
xor XOR2 (N11334, N11328, N7214);
nand NAND3 (N11335, N11323, N7236, N1124);
xor XOR2 (N11336, N11315, N6627);
buf BUF1 (N11337, N11335);
not NOT1 (N11338, N11336);
not NOT1 (N11339, N11325);
or OR2 (N11340, N11339, N9534);
nor NOR4 (N11341, N11317, N6158, N7019, N4048);
or OR4 (N11342, N11329, N7465, N9589, N2598);
or OR2 (N11343, N11334, N6213);
nor NOR2 (N11344, N11331, N10470);
xor XOR2 (N11345, N11344, N4045);
nor NOR4 (N11346, N11338, N5061, N749, N10144);
nand NAND2 (N11347, N11332, N3070);
and AND3 (N11348, N11330, N4323, N4305);
nor NOR2 (N11349, N11343, N3179);
and AND3 (N11350, N11345, N5068, N6873);
nor NOR2 (N11351, N11340, N10120);
not NOT1 (N11352, N11349);
nand NAND4 (N11353, N11342, N5766, N5525, N8495);
nand NAND2 (N11354, N11333, N7965);
not NOT1 (N11355, N11354);
or OR3 (N11356, N11350, N10411, N8628);
not NOT1 (N11357, N11337);
and AND2 (N11358, N11355, N175);
or OR2 (N11359, N11358, N4696);
or OR2 (N11360, N11347, N3431);
nor NOR3 (N11361, N11357, N6329, N941);
nor NOR4 (N11362, N11353, N10542, N3591, N6810);
and AND2 (N11363, N11359, N1054);
nand NAND2 (N11364, N11352, N1163);
and AND4 (N11365, N11341, N5750, N5672, N7473);
buf BUF1 (N11366, N11361);
or OR3 (N11367, N11362, N3253, N1665);
nor NOR4 (N11368, N11366, N10439, N7720, N7962);
nor NOR3 (N11369, N11348, N8019, N2912);
or OR4 (N11370, N11368, N7131, N509, N3725);
xor XOR2 (N11371, N11363, N133);
or OR3 (N11372, N11364, N448, N3895);
or OR3 (N11373, N11356, N5965, N8751);
and AND2 (N11374, N11365, N11000);
nor NOR3 (N11375, N11369, N8213, N10797);
nand NAND4 (N11376, N11372, N7321, N9107, N5040);
buf BUF1 (N11377, N11367);
buf BUF1 (N11378, N11377);
or OR4 (N11379, N11351, N10568, N8690, N6950);
xor XOR2 (N11380, N11360, N579);
and AND4 (N11381, N11373, N11152, N1503, N436);
not NOT1 (N11382, N11379);
buf BUF1 (N11383, N11375);
not NOT1 (N11384, N11378);
buf BUF1 (N11385, N11374);
nand NAND4 (N11386, N11383, N9024, N7710, N7626);
xor XOR2 (N11387, N11385, N10287);
and AND4 (N11388, N11384, N669, N1708, N10035);
nand NAND4 (N11389, N11380, N10760, N10648, N2826);
nand NAND2 (N11390, N11382, N10987);
nand NAND3 (N11391, N11381, N6030, N8087);
and AND3 (N11392, N11388, N9601, N11238);
nand NAND4 (N11393, N11346, N169, N2166, N6728);
xor XOR2 (N11394, N11390, N3760);
nand NAND4 (N11395, N11371, N8414, N7210, N8233);
xor XOR2 (N11396, N11389, N4371);
nor NOR3 (N11397, N11394, N7859, N34);
not NOT1 (N11398, N11393);
and AND2 (N11399, N11387, N8376);
xor XOR2 (N11400, N11370, N6527);
nand NAND2 (N11401, N11391, N6798);
nand NAND2 (N11402, N11401, N2684);
and AND4 (N11403, N11386, N6606, N5684, N5929);
and AND3 (N11404, N11402, N11075, N136);
nand NAND2 (N11405, N11392, N8242);
nor NOR3 (N11406, N11396, N1944, N9384);
nor NOR4 (N11407, N11406, N3290, N7481, N1659);
buf BUF1 (N11408, N11395);
buf BUF1 (N11409, N11404);
and AND3 (N11410, N11408, N5154, N6406);
not NOT1 (N11411, N11410);
not NOT1 (N11412, N11376);
buf BUF1 (N11413, N11400);
nand NAND4 (N11414, N11413, N11272, N7755, N3614);
nor NOR4 (N11415, N11407, N38, N9479, N1727);
nor NOR2 (N11416, N11398, N10499);
and AND4 (N11417, N11403, N1107, N9006, N7746);
nor NOR3 (N11418, N11411, N10219, N10520);
buf BUF1 (N11419, N11412);
buf BUF1 (N11420, N11399);
or OR3 (N11421, N11419, N3284, N9599);
xor XOR2 (N11422, N11418, N43);
xor XOR2 (N11423, N11409, N6968);
and AND2 (N11424, N11416, N2188);
nor NOR2 (N11425, N11424, N6406);
nand NAND4 (N11426, N11415, N4610, N10388, N9841);
nor NOR3 (N11427, N11414, N2079, N8080);
not NOT1 (N11428, N11425);
nand NAND3 (N11429, N11428, N8983, N7178);
buf BUF1 (N11430, N11397);
nand NAND2 (N11431, N11422, N8669);
buf BUF1 (N11432, N11429);
xor XOR2 (N11433, N11426, N6363);
and AND3 (N11434, N11433, N7665, N173);
or OR3 (N11435, N11405, N8345, N2942);
buf BUF1 (N11436, N11417);
or OR2 (N11437, N11432, N5004);
not NOT1 (N11438, N11430);
or OR3 (N11439, N11437, N6471, N9950);
xor XOR2 (N11440, N11431, N10885);
or OR2 (N11441, N11439, N8418);
not NOT1 (N11442, N11435);
buf BUF1 (N11443, N11434);
nor NOR4 (N11444, N11443, N7181, N5347, N10257);
buf BUF1 (N11445, N11440);
buf BUF1 (N11446, N11423);
and AND2 (N11447, N11441, N7197);
and AND4 (N11448, N11445, N9851, N1573, N10147);
buf BUF1 (N11449, N11446);
xor XOR2 (N11450, N11420, N6950);
not NOT1 (N11451, N11436);
or OR4 (N11452, N11442, N10464, N4130, N8961);
buf BUF1 (N11453, N11438);
or OR2 (N11454, N11453, N554);
or OR2 (N11455, N11427, N7329);
xor XOR2 (N11456, N11449, N8699);
not NOT1 (N11457, N11447);
not NOT1 (N11458, N11451);
buf BUF1 (N11459, N11455);
nor NOR2 (N11460, N11452, N5841);
nand NAND3 (N11461, N11458, N4616, N2971);
xor XOR2 (N11462, N11454, N10786);
and AND3 (N11463, N11456, N5965, N10104);
nand NAND4 (N11464, N11463, N11228, N2732, N10077);
nor NOR2 (N11465, N11448, N7140);
buf BUF1 (N11466, N11444);
nand NAND2 (N11467, N11421, N4324);
xor XOR2 (N11468, N11460, N1689);
and AND3 (N11469, N11450, N8744, N3405);
xor XOR2 (N11470, N11468, N447);
xor XOR2 (N11471, N11467, N7522);
xor XOR2 (N11472, N11462, N3399);
buf BUF1 (N11473, N11470);
nand NAND3 (N11474, N11466, N9981, N7823);
buf BUF1 (N11475, N11474);
or OR4 (N11476, N11472, N1405, N7449, N6723);
buf BUF1 (N11477, N11476);
and AND2 (N11478, N11475, N11041);
or OR3 (N11479, N11459, N10067, N9141);
or OR3 (N11480, N11471, N11053, N4378);
nor NOR3 (N11481, N11465, N1666, N4490);
or OR2 (N11482, N11477, N9211);
or OR4 (N11483, N11457, N10183, N299, N1522);
and AND4 (N11484, N11481, N10348, N10985, N1936);
xor XOR2 (N11485, N11479, N1441);
and AND3 (N11486, N11484, N3561, N8969);
buf BUF1 (N11487, N11473);
nor NOR3 (N11488, N11485, N3400, N4252);
xor XOR2 (N11489, N11478, N3533);
nor NOR4 (N11490, N11489, N8443, N3378, N10976);
and AND4 (N11491, N11482, N1739, N11124, N5491);
xor XOR2 (N11492, N11480, N5018);
or OR4 (N11493, N11492, N1684, N4661, N6950);
nor NOR3 (N11494, N11488, N8761, N3096);
or OR2 (N11495, N11493, N6544);
nand NAND2 (N11496, N11487, N9030);
or OR2 (N11497, N11469, N4055);
and AND2 (N11498, N11491, N7961);
and AND2 (N11499, N11486, N9755);
nor NOR3 (N11500, N11496, N9611, N11099);
nor NOR4 (N11501, N11483, N5012, N4154, N1422);
not NOT1 (N11502, N11494);
nand NAND4 (N11503, N11490, N3598, N213, N8445);
buf BUF1 (N11504, N11498);
not NOT1 (N11505, N11461);
buf BUF1 (N11506, N11499);
not NOT1 (N11507, N11497);
nand NAND3 (N11508, N11464, N10945, N4285);
buf BUF1 (N11509, N11504);
buf BUF1 (N11510, N11507);
and AND2 (N11511, N11509, N7399);
xor XOR2 (N11512, N11506, N9163);
or OR2 (N11513, N11512, N6098);
not NOT1 (N11514, N11495);
buf BUF1 (N11515, N11513);
not NOT1 (N11516, N11503);
or OR3 (N11517, N11505, N11505, N6944);
or OR2 (N11518, N11510, N2286);
xor XOR2 (N11519, N11511, N10679);
xor XOR2 (N11520, N11501, N5252);
buf BUF1 (N11521, N11514);
and AND2 (N11522, N11520, N10521);
buf BUF1 (N11523, N11521);
or OR4 (N11524, N11515, N3192, N3106, N9602);
buf BUF1 (N11525, N11502);
xor XOR2 (N11526, N11517, N5197);
not NOT1 (N11527, N11526);
not NOT1 (N11528, N11527);
and AND3 (N11529, N11522, N8493, N4845);
nor NOR2 (N11530, N11518, N8591);
buf BUF1 (N11531, N11519);
and AND4 (N11532, N11516, N4627, N2938, N1117);
nand NAND4 (N11533, N11523, N4196, N2293, N383);
buf BUF1 (N11534, N11530);
not NOT1 (N11535, N11534);
not NOT1 (N11536, N11528);
or OR3 (N11537, N11525, N2274, N8490);
xor XOR2 (N11538, N11500, N1149);
nand NAND3 (N11539, N11538, N8825, N4082);
and AND2 (N11540, N11533, N7802);
or OR2 (N11541, N11535, N6892);
nor NOR3 (N11542, N11540, N5131, N790);
or OR4 (N11543, N11508, N7692, N9773, N3270);
nor NOR3 (N11544, N11531, N9504, N11484);
xor XOR2 (N11545, N11544, N10533);
buf BUF1 (N11546, N11542);
or OR4 (N11547, N11545, N6699, N981, N6569);
xor XOR2 (N11548, N11537, N10736);
nand NAND4 (N11549, N11529, N10625, N7150, N3113);
or OR4 (N11550, N11546, N8248, N4243, N5230);
or OR3 (N11551, N11550, N5755, N6714);
nor NOR2 (N11552, N11541, N4741);
buf BUF1 (N11553, N11552);
xor XOR2 (N11554, N11549, N6851);
not NOT1 (N11555, N11524);
nand NAND2 (N11556, N11551, N1956);
xor XOR2 (N11557, N11548, N216);
xor XOR2 (N11558, N11554, N7793);
or OR4 (N11559, N11558, N4729, N5189, N8686);
or OR4 (N11560, N11557, N8532, N9930, N3387);
nor NOR3 (N11561, N11560, N10683, N2615);
buf BUF1 (N11562, N11553);
not NOT1 (N11563, N11543);
or OR4 (N11564, N11555, N7780, N5733, N3503);
and AND3 (N11565, N11564, N6670, N5971);
or OR3 (N11566, N11561, N5958, N9841);
buf BUF1 (N11567, N11566);
buf BUF1 (N11568, N11563);
and AND2 (N11569, N11536, N1764);
buf BUF1 (N11570, N11565);
nor NOR2 (N11571, N11539, N3692);
and AND4 (N11572, N11547, N1437, N275, N5960);
and AND3 (N11573, N11567, N11060, N3639);
buf BUF1 (N11574, N11573);
buf BUF1 (N11575, N11572);
buf BUF1 (N11576, N11532);
nand NAND2 (N11577, N11571, N6099);
nor NOR3 (N11578, N11575, N9873, N7027);
not NOT1 (N11579, N11556);
buf BUF1 (N11580, N11562);
not NOT1 (N11581, N11574);
xor XOR2 (N11582, N11559, N10129);
nand NAND3 (N11583, N11576, N809, N10728);
buf BUF1 (N11584, N11583);
nor NOR4 (N11585, N11584, N8958, N6704, N8996);
nand NAND3 (N11586, N11577, N1373, N2132);
not NOT1 (N11587, N11586);
nor NOR4 (N11588, N11578, N8174, N6307, N11452);
not NOT1 (N11589, N11588);
and AND3 (N11590, N11570, N4578, N4026);
nor NOR2 (N11591, N11590, N9464);
not NOT1 (N11592, N11589);
nor NOR4 (N11593, N11591, N3931, N8030, N5324);
or OR3 (N11594, N11592, N11115, N8272);
nand NAND4 (N11595, N11587, N4956, N3645, N10487);
nor NOR3 (N11596, N11581, N6379, N4915);
buf BUF1 (N11597, N11593);
or OR3 (N11598, N11579, N8423, N9290);
or OR2 (N11599, N11594, N9195);
xor XOR2 (N11600, N11568, N4433);
nand NAND2 (N11601, N11596, N7994);
and AND2 (N11602, N11600, N6505);
nand NAND4 (N11603, N11598, N1663, N10206, N5937);
nand NAND2 (N11604, N11585, N11296);
nand NAND4 (N11605, N11569, N3579, N95, N5455);
and AND4 (N11606, N11602, N111, N5061, N817);
or OR2 (N11607, N11599, N3471);
xor XOR2 (N11608, N11595, N11607);
and AND3 (N11609, N180, N2960, N1512);
not NOT1 (N11610, N11604);
and AND2 (N11611, N11582, N4143);
and AND3 (N11612, N11603, N3106, N78);
buf BUF1 (N11613, N11612);
nor NOR2 (N11614, N11610, N7497);
and AND4 (N11615, N11613, N1698, N156, N9269);
xor XOR2 (N11616, N11601, N2624);
nand NAND3 (N11617, N11616, N5290, N1126);
buf BUF1 (N11618, N11597);
nand NAND2 (N11619, N11614, N7869);
not NOT1 (N11620, N11605);
nand NAND4 (N11621, N11615, N9109, N3025, N3829);
buf BUF1 (N11622, N11620);
not NOT1 (N11623, N11609);
or OR2 (N11624, N11621, N4748);
not NOT1 (N11625, N11617);
nor NOR3 (N11626, N11580, N11475, N1916);
or OR4 (N11627, N11606, N4974, N3961, N10345);
and AND3 (N11628, N11622, N8548, N1558);
or OR4 (N11629, N11618, N9138, N1103, N8236);
nor NOR3 (N11630, N11629, N865, N8906);
and AND3 (N11631, N11608, N576, N228);
buf BUF1 (N11632, N11627);
buf BUF1 (N11633, N11631);
nor NOR4 (N11634, N11619, N6120, N1787, N659);
xor XOR2 (N11635, N11633, N6650);
not NOT1 (N11636, N11611);
nor NOR2 (N11637, N11636, N9956);
nor NOR2 (N11638, N11626, N5580);
nor NOR4 (N11639, N11637, N800, N8612, N6320);
not NOT1 (N11640, N11639);
nor NOR3 (N11641, N11628, N3960, N2117);
nor NOR2 (N11642, N11625, N5554);
nand NAND4 (N11643, N11640, N11536, N10428, N4327);
nor NOR3 (N11644, N11635, N8369, N325);
and AND4 (N11645, N11632, N1632, N10130, N8490);
not NOT1 (N11646, N11634);
nor NOR4 (N11647, N11645, N4868, N606, N10295);
nand NAND2 (N11648, N11638, N8271);
not NOT1 (N11649, N11644);
buf BUF1 (N11650, N11642);
nor NOR2 (N11651, N11643, N9788);
buf BUF1 (N11652, N11646);
or OR3 (N11653, N11649, N11449, N532);
nand NAND2 (N11654, N11652, N4380);
and AND2 (N11655, N11641, N9898);
and AND2 (N11656, N11651, N4690);
and AND3 (N11657, N11647, N8902, N9988);
or OR3 (N11658, N11650, N5561, N10261);
nand NAND3 (N11659, N11657, N4724, N4771);
nand NAND4 (N11660, N11624, N10171, N10203, N9715);
nand NAND3 (N11661, N11655, N1623, N4881);
nor NOR4 (N11662, N11654, N3998, N2384, N5038);
nor NOR3 (N11663, N11653, N2531, N10160);
not NOT1 (N11664, N11630);
and AND3 (N11665, N11663, N2835, N10393);
xor XOR2 (N11666, N11658, N9160);
not NOT1 (N11667, N11659);
xor XOR2 (N11668, N11648, N5020);
nand NAND3 (N11669, N11662, N8911, N9651);
nor NOR3 (N11670, N11623, N9535, N3852);
buf BUF1 (N11671, N11656);
not NOT1 (N11672, N11661);
xor XOR2 (N11673, N11669, N3083);
nor NOR3 (N11674, N11664, N841, N11204);
buf BUF1 (N11675, N11672);
buf BUF1 (N11676, N11665);
and AND3 (N11677, N11670, N10058, N4115);
nor NOR4 (N11678, N11671, N5892, N9497, N3798);
nor NOR2 (N11679, N11666, N1043);
nand NAND3 (N11680, N11679, N9692, N3428);
nor NOR4 (N11681, N11675, N7229, N8569, N2662);
nand NAND3 (N11682, N11668, N3370, N2197);
buf BUF1 (N11683, N11673);
nor NOR2 (N11684, N11677, N9581);
buf BUF1 (N11685, N11682);
buf BUF1 (N11686, N11667);
nor NOR2 (N11687, N11683, N5898);
xor XOR2 (N11688, N11680, N1102);
and AND3 (N11689, N11684, N6186, N6325);
xor XOR2 (N11690, N11678, N7063);
buf BUF1 (N11691, N11687);
and AND2 (N11692, N11681, N5080);
or OR3 (N11693, N11689, N5405, N4042);
xor XOR2 (N11694, N11692, N9282);
not NOT1 (N11695, N11693);
and AND3 (N11696, N11676, N10694, N7236);
or OR4 (N11697, N11688, N4053, N6690, N1647);
and AND4 (N11698, N11694, N9919, N10396, N7541);
nor NOR3 (N11699, N11697, N3647, N2848);
nand NAND2 (N11700, N11685, N2508);
nor NOR2 (N11701, N11690, N3991);
xor XOR2 (N11702, N11695, N9162);
and AND2 (N11703, N11699, N8587);
xor XOR2 (N11704, N11698, N1226);
and AND2 (N11705, N11700, N11636);
xor XOR2 (N11706, N11674, N7817);
or OR2 (N11707, N11701, N11243);
or OR4 (N11708, N11704, N9124, N2910, N11292);
nand NAND3 (N11709, N11703, N44, N10538);
or OR2 (N11710, N11696, N1621);
not NOT1 (N11711, N11710);
nand NAND3 (N11712, N11707, N2269, N10807);
nand NAND4 (N11713, N11686, N9718, N5018, N4529);
nor NOR2 (N11714, N11705, N5446);
nor NOR3 (N11715, N11709, N6431, N9956);
nand NAND2 (N11716, N11660, N11252);
nand NAND3 (N11717, N11713, N11458, N5590);
xor XOR2 (N11718, N11715, N960);
xor XOR2 (N11719, N11718, N10812);
not NOT1 (N11720, N11702);
not NOT1 (N11721, N11714);
or OR4 (N11722, N11706, N10381, N3095, N2438);
and AND2 (N11723, N11711, N9390);
xor XOR2 (N11724, N11708, N6979);
not NOT1 (N11725, N11721);
not NOT1 (N11726, N11724);
or OR2 (N11727, N11719, N7952);
and AND4 (N11728, N11727, N9509, N1995, N5303);
and AND3 (N11729, N11720, N5059, N749);
buf BUF1 (N11730, N11691);
and AND2 (N11731, N11730, N9806);
and AND3 (N11732, N11723, N103, N1854);
buf BUF1 (N11733, N11726);
xor XOR2 (N11734, N11732, N5867);
xor XOR2 (N11735, N11725, N11590);
and AND3 (N11736, N11722, N9514, N4690);
nand NAND4 (N11737, N11728, N9087, N38, N8910);
nand NAND4 (N11738, N11712, N4398, N6316, N8587);
nor NOR3 (N11739, N11717, N4847, N4243);
nor NOR3 (N11740, N11739, N2794, N8153);
not NOT1 (N11741, N11735);
nor NOR3 (N11742, N11731, N9550, N1064);
nand NAND4 (N11743, N11729, N3592, N7980, N4333);
and AND2 (N11744, N11741, N2343);
nor NOR4 (N11745, N11738, N5978, N10891, N73);
or OR4 (N11746, N11745, N8860, N2802, N9167);
and AND3 (N11747, N11744, N2957, N6210);
and AND2 (N11748, N11737, N1437);
xor XOR2 (N11749, N11747, N10727);
or OR3 (N11750, N11746, N226, N1034);
not NOT1 (N11751, N11736);
nand NAND3 (N11752, N11743, N7444, N6664);
buf BUF1 (N11753, N11734);
not NOT1 (N11754, N11750);
nor NOR4 (N11755, N11748, N5987, N7648, N2918);
not NOT1 (N11756, N11740);
nand NAND3 (N11757, N11756, N3145, N1972);
buf BUF1 (N11758, N11751);
and AND4 (N11759, N11754, N1422, N5538, N8367);
nand NAND2 (N11760, N11758, N1124);
xor XOR2 (N11761, N11753, N8392);
nand NAND3 (N11762, N11761, N4223, N6789);
not NOT1 (N11763, N11757);
nand NAND4 (N11764, N11762, N188, N5291, N3514);
and AND3 (N11765, N11716, N4859, N1061);
nand NAND4 (N11766, N11763, N4001, N9952, N1242);
xor XOR2 (N11767, N11749, N10839);
xor XOR2 (N11768, N11764, N9926);
and AND4 (N11769, N11755, N931, N6548, N2088);
buf BUF1 (N11770, N11766);
not NOT1 (N11771, N11770);
xor XOR2 (N11772, N11760, N10823);
not NOT1 (N11773, N11759);
not NOT1 (N11774, N11752);
nand NAND2 (N11775, N11772, N815);
xor XOR2 (N11776, N11773, N6494);
not NOT1 (N11777, N11776);
and AND4 (N11778, N11742, N7047, N7318, N83);
nor NOR3 (N11779, N11769, N11074, N4433);
not NOT1 (N11780, N11767);
nor NOR4 (N11781, N11777, N11627, N8190, N4399);
nand NAND4 (N11782, N11778, N733, N8839, N1462);
nor NOR4 (N11783, N11779, N6581, N9757, N9905);
nand NAND2 (N11784, N11780, N5567);
nand NAND3 (N11785, N11783, N5954, N245);
nand NAND3 (N11786, N11771, N11227, N9732);
nand NAND4 (N11787, N11781, N9227, N5983, N3096);
and AND2 (N11788, N11733, N10144);
or OR2 (N11789, N11775, N11438);
xor XOR2 (N11790, N11765, N11058);
not NOT1 (N11791, N11790);
and AND4 (N11792, N11784, N5556, N3258, N9672);
not NOT1 (N11793, N11791);
not NOT1 (N11794, N11774);
or OR4 (N11795, N11786, N270, N11619, N9427);
or OR2 (N11796, N11789, N5701);
nand NAND4 (N11797, N11796, N6149, N1146, N9898);
and AND3 (N11798, N11787, N704, N8254);
not NOT1 (N11799, N11797);
nor NOR2 (N11800, N11795, N8439);
or OR2 (N11801, N11794, N7599);
xor XOR2 (N11802, N11785, N7268);
or OR4 (N11803, N11788, N6666, N11754, N3836);
buf BUF1 (N11804, N11802);
nor NOR4 (N11805, N11803, N6856, N2550, N6121);
nand NAND3 (N11806, N11801, N10824, N3942);
and AND3 (N11807, N11798, N1500, N3244);
or OR3 (N11808, N11806, N1924, N5514);
and AND4 (N11809, N11807, N5259, N3091, N2439);
nor NOR3 (N11810, N11799, N4140, N1050);
nand NAND2 (N11811, N11782, N8071);
nor NOR4 (N11812, N11793, N1545, N9385, N8301);
nand NAND4 (N11813, N11792, N4875, N5664, N2313);
buf BUF1 (N11814, N11809);
xor XOR2 (N11815, N11813, N1552);
nor NOR2 (N11816, N11805, N7268);
or OR4 (N11817, N11810, N7003, N2427, N431);
and AND3 (N11818, N11817, N4341, N5313);
nor NOR2 (N11819, N11800, N4923);
nand NAND4 (N11820, N11814, N6207, N6853, N828);
and AND4 (N11821, N11808, N2325, N2167, N9375);
not NOT1 (N11822, N11816);
and AND4 (N11823, N11819, N5774, N7950, N7329);
xor XOR2 (N11824, N11818, N3960);
not NOT1 (N11825, N11811);
nand NAND2 (N11826, N11812, N9037);
buf BUF1 (N11827, N11823);
not NOT1 (N11828, N11768);
nor NOR3 (N11829, N11821, N3592, N11625);
buf BUF1 (N11830, N11820);
not NOT1 (N11831, N11815);
nor NOR3 (N11832, N11827, N8253, N9941);
and AND2 (N11833, N11829, N9819);
xor XOR2 (N11834, N11832, N7548);
not NOT1 (N11835, N11826);
nor NOR4 (N11836, N11825, N4921, N10676, N9882);
buf BUF1 (N11837, N11834);
nand NAND2 (N11838, N11822, N5224);
xor XOR2 (N11839, N11838, N3021);
or OR3 (N11840, N11828, N11365, N1126);
and AND2 (N11841, N11836, N454);
not NOT1 (N11842, N11830);
not NOT1 (N11843, N11842);
buf BUF1 (N11844, N11835);
and AND4 (N11845, N11843, N7279, N4707, N1041);
nor NOR3 (N11846, N11837, N1261, N9067);
nand NAND3 (N11847, N11841, N465, N3142);
not NOT1 (N11848, N11844);
nor NOR3 (N11849, N11847, N3965, N11306);
buf BUF1 (N11850, N11848);
buf BUF1 (N11851, N11849);
and AND4 (N11852, N11839, N7961, N7870, N3809);
not NOT1 (N11853, N11804);
or OR2 (N11854, N11850, N419);
and AND4 (N11855, N11824, N8244, N4485, N7979);
and AND2 (N11856, N11846, N1671);
and AND4 (N11857, N11853, N4218, N4695, N5873);
nand NAND4 (N11858, N11833, N7807, N11821, N3706);
not NOT1 (N11859, N11845);
xor XOR2 (N11860, N11852, N4403);
buf BUF1 (N11861, N11857);
nand NAND4 (N11862, N11856, N5814, N8550, N6616);
not NOT1 (N11863, N11851);
not NOT1 (N11864, N11854);
not NOT1 (N11865, N11864);
buf BUF1 (N11866, N11860);
nor NOR2 (N11867, N11840, N2206);
nand NAND4 (N11868, N11863, N4637, N5046, N10867);
buf BUF1 (N11869, N11862);
or OR3 (N11870, N11868, N7469, N2104);
nor NOR4 (N11871, N11867, N6503, N8629, N9529);
not NOT1 (N11872, N11831);
xor XOR2 (N11873, N11871, N830);
buf BUF1 (N11874, N11870);
xor XOR2 (N11875, N11873, N6359);
nor NOR3 (N11876, N11866, N3220, N3540);
or OR2 (N11877, N11859, N4020);
xor XOR2 (N11878, N11877, N10507);
nor NOR2 (N11879, N11874, N744);
not NOT1 (N11880, N11861);
not NOT1 (N11881, N11865);
nand NAND3 (N11882, N11872, N3398, N2871);
buf BUF1 (N11883, N11875);
buf BUF1 (N11884, N11858);
xor XOR2 (N11885, N11878, N331);
not NOT1 (N11886, N11883);
nor NOR2 (N11887, N11881, N2285);
and AND3 (N11888, N11879, N5217, N6183);
nor NOR3 (N11889, N11876, N5576, N11076);
xor XOR2 (N11890, N11885, N8742);
buf BUF1 (N11891, N11889);
or OR3 (N11892, N11882, N9588, N4338);
or OR3 (N11893, N11880, N7436, N5566);
nand NAND3 (N11894, N11884, N6167, N153);
and AND3 (N11895, N11855, N5501, N2675);
xor XOR2 (N11896, N11894, N10740);
or OR3 (N11897, N11893, N7965, N3626);
buf BUF1 (N11898, N11886);
nor NOR2 (N11899, N11892, N5091);
and AND2 (N11900, N11897, N2715);
and AND4 (N11901, N11890, N3455, N10001, N11780);
nand NAND2 (N11902, N11869, N2972);
nor NOR2 (N11903, N11900, N11445);
not NOT1 (N11904, N11891);
buf BUF1 (N11905, N11901);
or OR4 (N11906, N11887, N9283, N3365, N6007);
or OR3 (N11907, N11903, N5672, N234);
not NOT1 (N11908, N11896);
nor NOR4 (N11909, N11907, N11423, N8255, N2381);
and AND2 (N11910, N11904, N80);
xor XOR2 (N11911, N11898, N9005);
nor NOR4 (N11912, N11911, N21, N5188, N7771);
nand NAND4 (N11913, N11912, N3301, N7046, N1748);
buf BUF1 (N11914, N11910);
and AND2 (N11915, N11914, N10706);
xor XOR2 (N11916, N11895, N2666);
not NOT1 (N11917, N11909);
nand NAND2 (N11918, N11888, N3094);
or OR2 (N11919, N11913, N11857);
or OR4 (N11920, N11906, N5731, N8591, N6258);
nand NAND3 (N11921, N11918, N6960, N4451);
nor NOR2 (N11922, N11899, N8242);
nand NAND4 (N11923, N11922, N1708, N3311, N5956);
or OR4 (N11924, N11921, N5312, N3005, N10097);
nand NAND4 (N11925, N11916, N11335, N9571, N6164);
not NOT1 (N11926, N11919);
or OR4 (N11927, N11902, N208, N10122, N8234);
not NOT1 (N11928, N11926);
nand NAND3 (N11929, N11925, N6981, N3480);
nor NOR4 (N11930, N11928, N3034, N3344, N4547);
buf BUF1 (N11931, N11923);
not NOT1 (N11932, N11920);
xor XOR2 (N11933, N11924, N6909);
xor XOR2 (N11934, N11908, N3614);
buf BUF1 (N11935, N11930);
buf BUF1 (N11936, N11934);
xor XOR2 (N11937, N11936, N10609);
buf BUF1 (N11938, N11932);
or OR2 (N11939, N11935, N5870);
and AND2 (N11940, N11937, N6514);
or OR3 (N11941, N11929, N8564, N9490);
nor NOR2 (N11942, N11938, N1913);
nor NOR4 (N11943, N11941, N8316, N1394, N277);
or OR3 (N11944, N11940, N6642, N1839);
or OR2 (N11945, N11915, N1275);
nand NAND3 (N11946, N11931, N4417, N8008);
not NOT1 (N11947, N11933);
nor NOR4 (N11948, N11945, N3174, N3476, N11004);
not NOT1 (N11949, N11944);
nand NAND4 (N11950, N11943, N7433, N2171, N10760);
buf BUF1 (N11951, N11946);
xor XOR2 (N11952, N11951, N1524);
nand NAND4 (N11953, N11952, N2927, N129, N4471);
nor NOR2 (N11954, N11939, N8194);
not NOT1 (N11955, N11905);
and AND3 (N11956, N11950, N3731, N5519);
or OR2 (N11957, N11927, N7552);
nor NOR4 (N11958, N11957, N7098, N4475, N3343);
or OR3 (N11959, N11954, N2210, N1085);
buf BUF1 (N11960, N11942);
nand NAND4 (N11961, N11917, N1192, N10276, N6124);
nor NOR3 (N11962, N11959, N7665, N2780);
buf BUF1 (N11963, N11960);
not NOT1 (N11964, N11956);
and AND2 (N11965, N11947, N9698);
and AND2 (N11966, N11948, N2762);
not NOT1 (N11967, N11965);
xor XOR2 (N11968, N11964, N4806);
buf BUF1 (N11969, N11955);
or OR2 (N11970, N11963, N10016);
not NOT1 (N11971, N11958);
buf BUF1 (N11972, N11966);
not NOT1 (N11973, N11969);
xor XOR2 (N11974, N11968, N10499);
not NOT1 (N11975, N11962);
buf BUF1 (N11976, N11975);
or OR2 (N11977, N11961, N10932);
and AND4 (N11978, N11970, N9432, N3538, N1877);
nand NAND4 (N11979, N11976, N4747, N8850, N3059);
not NOT1 (N11980, N11967);
nand NAND4 (N11981, N11980, N2879, N182, N4410);
nand NAND3 (N11982, N11979, N4922, N2630);
and AND3 (N11983, N11971, N7531, N8268);
not NOT1 (N11984, N11973);
and AND4 (N11985, N11981, N2768, N1451, N8391);
and AND4 (N11986, N11985, N11310, N11296, N5347);
or OR4 (N11987, N11978, N7218, N11046, N10267);
or OR4 (N11988, N11982, N5074, N6057, N7930);
or OR4 (N11989, N11974, N6192, N8221, N11229);
and AND2 (N11990, N11949, N9420);
nor NOR2 (N11991, N11984, N7360);
and AND2 (N11992, N11988, N6556);
buf BUF1 (N11993, N11953);
nor NOR3 (N11994, N11993, N10538, N11375);
not NOT1 (N11995, N11990);
or OR3 (N11996, N11986, N2837, N3514);
xor XOR2 (N11997, N11991, N8071);
nor NOR3 (N11998, N11972, N352, N10487);
xor XOR2 (N11999, N11994, N11820);
or OR3 (N12000, N11987, N9895, N5536);
or OR4 (N12001, N11995, N5359, N1792, N11386);
nand NAND2 (N12002, N11989, N7367);
xor XOR2 (N12003, N11992, N9586);
nand NAND3 (N12004, N12001, N11877, N6651);
nor NOR3 (N12005, N11996, N3011, N5089);
not NOT1 (N12006, N11998);
nor NOR2 (N12007, N11997, N5664);
nor NOR2 (N12008, N12004, N8452);
nor NOR3 (N12009, N12005, N11726, N870);
and AND3 (N12010, N12008, N4203, N7412);
buf BUF1 (N12011, N11983);
xor XOR2 (N12012, N12000, N10990);
not NOT1 (N12013, N12009);
nor NOR3 (N12014, N12011, N4981, N7961);
xor XOR2 (N12015, N12006, N8768);
nor NOR4 (N12016, N12007, N8684, N10855, N10190);
xor XOR2 (N12017, N12014, N2414);
nor NOR3 (N12018, N12017, N7384, N8390);
or OR3 (N12019, N12010, N7431, N1763);
xor XOR2 (N12020, N12002, N5792);
nor NOR2 (N12021, N12020, N11158);
xor XOR2 (N12022, N12019, N9623);
nand NAND4 (N12023, N12021, N7158, N4062, N4268);
and AND2 (N12024, N12012, N2278);
nor NOR3 (N12025, N12013, N9515, N7579);
xor XOR2 (N12026, N12018, N11357);
xor XOR2 (N12027, N12015, N11436);
buf BUF1 (N12028, N12016);
xor XOR2 (N12029, N12026, N3462);
and AND4 (N12030, N12022, N2750, N9361, N9649);
and AND2 (N12031, N12030, N7219);
not NOT1 (N12032, N12027);
nor NOR2 (N12033, N12032, N9964);
nand NAND3 (N12034, N12028, N2617, N5635);
buf BUF1 (N12035, N11977);
nor NOR2 (N12036, N12025, N419);
xor XOR2 (N12037, N12023, N3916);
or OR2 (N12038, N12029, N9295);
not NOT1 (N12039, N12031);
nand NAND2 (N12040, N12038, N7425);
buf BUF1 (N12041, N12040);
buf BUF1 (N12042, N12036);
buf BUF1 (N12043, N11999);
and AND2 (N12044, N12024, N8873);
xor XOR2 (N12045, N12035, N1747);
nand NAND4 (N12046, N12034, N8833, N8267, N3601);
nand NAND4 (N12047, N12044, N3464, N9513, N5040);
nand NAND3 (N12048, N12039, N1384, N1781);
and AND3 (N12049, N12003, N1818, N9672);
xor XOR2 (N12050, N12046, N6222);
not NOT1 (N12051, N12042);
buf BUF1 (N12052, N12049);
xor XOR2 (N12053, N12045, N9478);
not NOT1 (N12054, N12048);
or OR3 (N12055, N12043, N2316, N1528);
and AND4 (N12056, N12033, N8609, N3406, N2263);
buf BUF1 (N12057, N12041);
nor NOR3 (N12058, N12051, N1986, N3531);
not NOT1 (N12059, N12055);
buf BUF1 (N12060, N12059);
and AND3 (N12061, N12053, N10967, N3772);
buf BUF1 (N12062, N12060);
not NOT1 (N12063, N12056);
buf BUF1 (N12064, N12052);
not NOT1 (N12065, N12050);
not NOT1 (N12066, N12057);
or OR2 (N12067, N12063, N3957);
buf BUF1 (N12068, N12061);
or OR3 (N12069, N12067, N4282, N9953);
or OR3 (N12070, N12062, N4560, N2200);
or OR4 (N12071, N12069, N10232, N6931, N8818);
or OR2 (N12072, N12037, N521);
or OR2 (N12073, N12066, N11942);
nor NOR2 (N12074, N12064, N1503);
nor NOR3 (N12075, N12074, N4697, N1367);
and AND4 (N12076, N12072, N5925, N10595, N10161);
buf BUF1 (N12077, N12073);
and AND2 (N12078, N12075, N529);
nor NOR2 (N12079, N12078, N3635);
nand NAND3 (N12080, N12076, N10276, N8032);
not NOT1 (N12081, N12079);
not NOT1 (N12082, N12054);
and AND4 (N12083, N12047, N1364, N12023, N1848);
buf BUF1 (N12084, N12068);
and AND3 (N12085, N12070, N6872, N551);
nor NOR2 (N12086, N12071, N5078);
xor XOR2 (N12087, N12082, N94);
buf BUF1 (N12088, N12086);
not NOT1 (N12089, N12087);
nand NAND2 (N12090, N12088, N9395);
xor XOR2 (N12091, N12058, N5729);
buf BUF1 (N12092, N12065);
buf BUF1 (N12093, N12090);
nor NOR2 (N12094, N12083, N11196);
buf BUF1 (N12095, N12091);
nor NOR4 (N12096, N12089, N6825, N1176, N5702);
xor XOR2 (N12097, N12094, N1862);
nor NOR4 (N12098, N12095, N4001, N3635, N10082);
nor NOR4 (N12099, N12085, N4007, N10096, N11831);
not NOT1 (N12100, N12077);
not NOT1 (N12101, N12093);
nand NAND3 (N12102, N12099, N2675, N11195);
nor NOR2 (N12103, N12100, N3681);
nor NOR2 (N12104, N12103, N4066);
or OR4 (N12105, N12104, N7167, N5096, N3107);
or OR4 (N12106, N12080, N6189, N7504, N2143);
nor NOR3 (N12107, N12098, N5920, N3839);
nor NOR3 (N12108, N12102, N4552, N5058);
not NOT1 (N12109, N12105);
buf BUF1 (N12110, N12107);
buf BUF1 (N12111, N12084);
or OR3 (N12112, N12110, N836, N6489);
nand NAND4 (N12113, N12106, N6438, N6087, N8531);
or OR4 (N12114, N12109, N3799, N7210, N9079);
or OR3 (N12115, N12081, N9771, N5711);
or OR2 (N12116, N12101, N837);
not NOT1 (N12117, N12113);
nor NOR4 (N12118, N12115, N9036, N11514, N732);
xor XOR2 (N12119, N12112, N8507);
buf BUF1 (N12120, N12114);
nor NOR4 (N12121, N12111, N5728, N6907, N5384);
or OR4 (N12122, N12121, N941, N208, N3390);
nor NOR4 (N12123, N12108, N1676, N7524, N7098);
buf BUF1 (N12124, N12120);
nor NOR4 (N12125, N12117, N9805, N1678, N11114);
nand NAND4 (N12126, N12097, N4006, N5654, N8873);
nand NAND2 (N12127, N12116, N10166);
not NOT1 (N12128, N12125);
not NOT1 (N12129, N12128);
or OR4 (N12130, N12124, N7970, N10826, N885);
xor XOR2 (N12131, N12127, N9220);
nor NOR3 (N12132, N12096, N2777, N4632);
nand NAND3 (N12133, N12126, N9739, N5418);
nor NOR4 (N12134, N12132, N3492, N3356, N11547);
and AND2 (N12135, N12129, N9808);
and AND3 (N12136, N12092, N8162, N7904);
nor NOR4 (N12137, N12133, N1986, N9476, N1572);
not NOT1 (N12138, N12123);
xor XOR2 (N12139, N12119, N10620);
or OR2 (N12140, N12139, N4319);
and AND2 (N12141, N12137, N7695);
not NOT1 (N12142, N12134);
nor NOR4 (N12143, N12131, N6645, N6317, N2375);
buf BUF1 (N12144, N12140);
xor XOR2 (N12145, N12130, N10920);
or OR4 (N12146, N12118, N2722, N11275, N6834);
buf BUF1 (N12147, N12143);
nor NOR4 (N12148, N12147, N1320, N243, N1584);
or OR4 (N12149, N12142, N5816, N5959, N11126);
buf BUF1 (N12150, N12145);
xor XOR2 (N12151, N12149, N11300);
and AND2 (N12152, N12148, N2428);
buf BUF1 (N12153, N12150);
buf BUF1 (N12154, N12146);
nand NAND3 (N12155, N12144, N3706, N10118);
not NOT1 (N12156, N12136);
and AND4 (N12157, N12155, N8759, N520, N7885);
buf BUF1 (N12158, N12153);
and AND2 (N12159, N12122, N474);
not NOT1 (N12160, N12156);
not NOT1 (N12161, N12157);
not NOT1 (N12162, N12158);
buf BUF1 (N12163, N12162);
buf BUF1 (N12164, N12154);
buf BUF1 (N12165, N12152);
or OR4 (N12166, N12135, N11548, N9821, N3950);
buf BUF1 (N12167, N12163);
buf BUF1 (N12168, N12159);
and AND4 (N12169, N12168, N3683, N6278, N9451);
not NOT1 (N12170, N12141);
and AND3 (N12171, N12164, N8086, N3061);
nand NAND4 (N12172, N12166, N6904, N9555, N6553);
not NOT1 (N12173, N12170);
and AND3 (N12174, N12151, N2351, N2018);
or OR4 (N12175, N12174, N5503, N10208, N1073);
nand NAND4 (N12176, N12173, N5209, N4169, N11497);
nor NOR4 (N12177, N12160, N8988, N4205, N11644);
and AND3 (N12178, N12177, N1203, N10185);
nand NAND3 (N12179, N12175, N11693, N3606);
not NOT1 (N12180, N12171);
not NOT1 (N12181, N12165);
buf BUF1 (N12182, N12181);
buf BUF1 (N12183, N12138);
nand NAND4 (N12184, N12180, N11412, N9456, N4597);
not NOT1 (N12185, N12167);
nand NAND4 (N12186, N12178, N5301, N11304, N6858);
and AND2 (N12187, N12179, N10292);
not NOT1 (N12188, N12184);
or OR4 (N12189, N12185, N4526, N9762, N2470);
nand NAND4 (N12190, N12161, N8589, N5990, N1047);
buf BUF1 (N12191, N12182);
or OR2 (N12192, N12189, N3051);
nor NOR4 (N12193, N12183, N4613, N11973, N11171);
not NOT1 (N12194, N12190);
nor NOR2 (N12195, N12191, N5134);
nor NOR3 (N12196, N12176, N8577, N9657);
nand NAND4 (N12197, N12169, N4839, N2407, N9322);
not NOT1 (N12198, N12196);
buf BUF1 (N12199, N12172);
buf BUF1 (N12200, N12195);
nor NOR3 (N12201, N12198, N3366, N12021);
nor NOR2 (N12202, N12188, N10986);
or OR4 (N12203, N12200, N3154, N6539, N11570);
xor XOR2 (N12204, N12187, N990);
nor NOR4 (N12205, N12202, N7175, N2217, N6290);
nor NOR4 (N12206, N12197, N7511, N4895, N2349);
nand NAND4 (N12207, N12201, N10652, N11422, N4051);
or OR2 (N12208, N12193, N9520);
buf BUF1 (N12209, N12205);
xor XOR2 (N12210, N12206, N7050);
nand NAND4 (N12211, N12203, N4823, N10612, N2274);
and AND3 (N12212, N12208, N5036, N1363);
and AND3 (N12213, N12194, N5697, N2526);
buf BUF1 (N12214, N12199);
buf BUF1 (N12215, N12209);
xor XOR2 (N12216, N12214, N3807);
xor XOR2 (N12217, N12213, N7750);
xor XOR2 (N12218, N12186, N1204);
nand NAND2 (N12219, N12218, N9257);
and AND4 (N12220, N12192, N523, N5070, N3984);
nor NOR3 (N12221, N12212, N4913, N2450);
nand NAND4 (N12222, N12217, N11840, N3670, N2613);
nor NOR2 (N12223, N12216, N4583);
nand NAND4 (N12224, N12222, N3095, N4595, N2796);
and AND3 (N12225, N12219, N9004, N9630);
or OR2 (N12226, N12211, N1544);
nand NAND4 (N12227, N12210, N6110, N5658, N7231);
not NOT1 (N12228, N12215);
buf BUF1 (N12229, N12220);
xor XOR2 (N12230, N12225, N2459);
xor XOR2 (N12231, N12221, N10070);
xor XOR2 (N12232, N12224, N672);
or OR4 (N12233, N12229, N10781, N9481, N2962);
not NOT1 (N12234, N12230);
nor NOR2 (N12235, N12204, N2825);
buf BUF1 (N12236, N12233);
nand NAND3 (N12237, N12227, N4982, N10591);
buf BUF1 (N12238, N12236);
not NOT1 (N12239, N12238);
and AND3 (N12240, N12226, N227, N1936);
xor XOR2 (N12241, N12239, N824);
not NOT1 (N12242, N12223);
nand NAND2 (N12243, N12241, N11890);
and AND4 (N12244, N12207, N5992, N8266, N7416);
and AND4 (N12245, N12240, N997, N5356, N9056);
not NOT1 (N12246, N12245);
or OR4 (N12247, N12246, N11246, N7464, N4044);
and AND4 (N12248, N12237, N1678, N5009, N1980);
buf BUF1 (N12249, N12234);
or OR3 (N12250, N12243, N5419, N3799);
nor NOR4 (N12251, N12228, N7281, N10885, N7585);
and AND4 (N12252, N12232, N12113, N7814, N3421);
nand NAND2 (N12253, N12248, N6822);
nor NOR4 (N12254, N12250, N10877, N4381, N10416);
buf BUF1 (N12255, N12253);
and AND3 (N12256, N12242, N11507, N7699);
xor XOR2 (N12257, N12244, N7793);
not NOT1 (N12258, N12247);
and AND4 (N12259, N12258, N8833, N1983, N1524);
not NOT1 (N12260, N12255);
or OR3 (N12261, N12251, N1032, N1843);
and AND3 (N12262, N12252, N10191, N10934);
nor NOR2 (N12263, N12262, N1685);
and AND2 (N12264, N12249, N10819);
xor XOR2 (N12265, N12264, N3733);
nor NOR3 (N12266, N12263, N7538, N10946);
buf BUF1 (N12267, N12235);
nand NAND4 (N12268, N12231, N7755, N7296, N8759);
buf BUF1 (N12269, N12259);
not NOT1 (N12270, N12267);
or OR3 (N12271, N12256, N3020, N213);
nand NAND3 (N12272, N12266, N5064, N8218);
xor XOR2 (N12273, N12271, N2958);
and AND2 (N12274, N12270, N565);
not NOT1 (N12275, N12261);
buf BUF1 (N12276, N12254);
xor XOR2 (N12277, N12265, N2809);
not NOT1 (N12278, N12273);
xor XOR2 (N12279, N12268, N8434);
not NOT1 (N12280, N12275);
not NOT1 (N12281, N12269);
or OR3 (N12282, N12272, N8268, N3244);
xor XOR2 (N12283, N12257, N9188);
and AND2 (N12284, N12276, N11483);
and AND2 (N12285, N12283, N5027);
and AND3 (N12286, N12278, N6806, N3488);
or OR3 (N12287, N12285, N6360, N1335);
nor NOR3 (N12288, N12260, N2475, N3930);
not NOT1 (N12289, N12282);
nand NAND2 (N12290, N12287, N4176);
or OR4 (N12291, N12290, N9692, N1849, N9889);
or OR3 (N12292, N12288, N4125, N3947);
and AND3 (N12293, N12274, N8380, N10408);
buf BUF1 (N12294, N12284);
or OR4 (N12295, N12286, N7392, N80, N3821);
and AND4 (N12296, N12277, N1660, N11460, N7980);
or OR2 (N12297, N12296, N7250);
buf BUF1 (N12298, N12279);
xor XOR2 (N12299, N12295, N5819);
nand NAND4 (N12300, N12291, N8417, N3071, N1487);
xor XOR2 (N12301, N12300, N8161);
nand NAND4 (N12302, N12299, N7660, N1059, N8381);
not NOT1 (N12303, N12281);
nor NOR4 (N12304, N12298, N7157, N8836, N10182);
buf BUF1 (N12305, N12294);
nand NAND3 (N12306, N12303, N8889, N9295);
nor NOR3 (N12307, N12297, N1222, N6565);
nand NAND4 (N12308, N12301, N912, N4789, N9585);
or OR4 (N12309, N12306, N7824, N288, N3836);
nor NOR3 (N12310, N12305, N11203, N12065);
buf BUF1 (N12311, N12310);
xor XOR2 (N12312, N12304, N5120);
not NOT1 (N12313, N12308);
buf BUF1 (N12314, N12292);
buf BUF1 (N12315, N12312);
nand NAND4 (N12316, N12280, N5917, N3360, N4426);
nand NAND2 (N12317, N12307, N5017);
nand NAND4 (N12318, N12314, N3857, N12075, N9549);
nor NOR2 (N12319, N12289, N5975);
not NOT1 (N12320, N12318);
and AND2 (N12321, N12317, N11515);
nand NAND3 (N12322, N12293, N11189, N3636);
and AND3 (N12323, N12313, N3890, N3402);
nor NOR4 (N12324, N12322, N3198, N2442, N522);
not NOT1 (N12325, N12316);
xor XOR2 (N12326, N12321, N5946);
nand NAND4 (N12327, N12326, N7648, N4292, N12320);
nand NAND3 (N12328, N3126, N8352, N9874);
not NOT1 (N12329, N12324);
nand NAND3 (N12330, N12325, N2352, N528);
nand NAND3 (N12331, N12329, N6337, N12106);
xor XOR2 (N12332, N12327, N437);
or OR4 (N12333, N12319, N3876, N1114, N7695);
buf BUF1 (N12334, N12323);
or OR4 (N12335, N12302, N1375, N9534, N9154);
buf BUF1 (N12336, N12309);
nand NAND2 (N12337, N12315, N4537);
not NOT1 (N12338, N12331);
nand NAND2 (N12339, N12332, N6168);
nand NAND4 (N12340, N12334, N9157, N6166, N6754);
buf BUF1 (N12341, N12339);
or OR4 (N12342, N12333, N1675, N1783, N9405);
nand NAND3 (N12343, N12336, N2348, N11270);
and AND2 (N12344, N12340, N3450);
xor XOR2 (N12345, N12342, N4981);
xor XOR2 (N12346, N12337, N2906);
buf BUF1 (N12347, N12344);
xor XOR2 (N12348, N12345, N9116);
xor XOR2 (N12349, N12343, N8559);
or OR4 (N12350, N12311, N1249, N2621, N1671);
buf BUF1 (N12351, N12338);
buf BUF1 (N12352, N12349);
xor XOR2 (N12353, N12351, N6880);
nand NAND4 (N12354, N12346, N1989, N8136, N10436);
xor XOR2 (N12355, N12352, N3677);
xor XOR2 (N12356, N12348, N1802);
nand NAND3 (N12357, N12328, N11086, N11282);
nor NOR2 (N12358, N12335, N258);
or OR2 (N12359, N12358, N7002);
or OR2 (N12360, N12350, N9286);
nor NOR4 (N12361, N12330, N10609, N9326, N2558);
xor XOR2 (N12362, N12356, N1773);
and AND3 (N12363, N12347, N3756, N2551);
xor XOR2 (N12364, N12363, N8995);
and AND3 (N12365, N12364, N3796, N9433);
nor NOR3 (N12366, N12365, N8428, N11287);
nor NOR4 (N12367, N12357, N10618, N1385, N703);
not NOT1 (N12368, N12362);
not NOT1 (N12369, N12368);
not NOT1 (N12370, N12359);
and AND4 (N12371, N12354, N5120, N11690, N11315);
nor NOR3 (N12372, N12371, N6108, N10625);
or OR2 (N12373, N12361, N11801);
xor XOR2 (N12374, N12355, N9003);
and AND4 (N12375, N12367, N9078, N442, N9166);
and AND3 (N12376, N12341, N8112, N10865);
and AND3 (N12377, N12366, N7892, N1631);
xor XOR2 (N12378, N12369, N135);
xor XOR2 (N12379, N12374, N1545);
nand NAND4 (N12380, N12372, N6488, N9540, N6588);
not NOT1 (N12381, N12379);
buf BUF1 (N12382, N12381);
nand NAND3 (N12383, N12370, N10986, N1062);
buf BUF1 (N12384, N12353);
and AND4 (N12385, N12380, N12177, N7132, N1261);
nand NAND3 (N12386, N12382, N6023, N1253);
buf BUF1 (N12387, N12375);
or OR3 (N12388, N12377, N11201, N2372);
nor NOR3 (N12389, N12385, N12057, N5819);
or OR3 (N12390, N12384, N11303, N6292);
nand NAND2 (N12391, N12389, N3737);
nor NOR2 (N12392, N12378, N2944);
not NOT1 (N12393, N12387);
or OR3 (N12394, N12391, N4606, N2489);
buf BUF1 (N12395, N12373);
xor XOR2 (N12396, N12395, N9674);
xor XOR2 (N12397, N12394, N4395);
and AND4 (N12398, N12392, N1443, N9857, N7464);
or OR2 (N12399, N12386, N11919);
xor XOR2 (N12400, N12398, N2993);
nor NOR4 (N12401, N12376, N9431, N12156, N11628);
buf BUF1 (N12402, N12360);
nor NOR3 (N12403, N12399, N6127, N1196);
not NOT1 (N12404, N12383);
nand NAND4 (N12405, N12404, N3578, N9560, N5390);
nand NAND4 (N12406, N12400, N10774, N778, N3152);
or OR2 (N12407, N12401, N7105);
or OR4 (N12408, N12396, N1701, N8584, N4887);
or OR3 (N12409, N12402, N4716, N5200);
buf BUF1 (N12410, N12388);
nand NAND4 (N12411, N12408, N9561, N2569, N5746);
nand NAND3 (N12412, N12397, N3279, N1646);
buf BUF1 (N12413, N12412);
nor NOR4 (N12414, N12409, N11980, N9659, N3995);
xor XOR2 (N12415, N12390, N8187);
nor NOR3 (N12416, N12407, N10438, N2624);
buf BUF1 (N12417, N12410);
and AND2 (N12418, N12411, N431);
not NOT1 (N12419, N12416);
nor NOR3 (N12420, N12417, N11316, N4076);
nand NAND2 (N12421, N12419, N9650);
not NOT1 (N12422, N12421);
buf BUF1 (N12423, N12413);
nand NAND2 (N12424, N12418, N1767);
xor XOR2 (N12425, N12415, N28);
or OR2 (N12426, N12424, N2026);
buf BUF1 (N12427, N12422);
and AND4 (N12428, N12406, N2600, N5050, N8314);
nor NOR4 (N12429, N12414, N1066, N1457, N8044);
nand NAND2 (N12430, N12425, N3298);
not NOT1 (N12431, N12420);
not NOT1 (N12432, N12393);
nand NAND2 (N12433, N12405, N11763);
buf BUF1 (N12434, N12433);
xor XOR2 (N12435, N12423, N142);
and AND4 (N12436, N12434, N2824, N4090, N5423);
nand NAND4 (N12437, N12427, N1113, N10125, N8266);
and AND2 (N12438, N12428, N7047);
buf BUF1 (N12439, N12435);
buf BUF1 (N12440, N12430);
not NOT1 (N12441, N12403);
nor NOR4 (N12442, N12429, N8308, N7061, N6486);
not NOT1 (N12443, N12441);
not NOT1 (N12444, N12438);
nor NOR3 (N12445, N12442, N6217, N2596);
and AND2 (N12446, N12443, N4865);
not NOT1 (N12447, N12431);
not NOT1 (N12448, N12447);
not NOT1 (N12449, N12448);
nand NAND4 (N12450, N12446, N6305, N5867, N8918);
nor NOR2 (N12451, N12440, N10209);
nand NAND2 (N12452, N12432, N4);
buf BUF1 (N12453, N12437);
or OR2 (N12454, N12445, N3591);
buf BUF1 (N12455, N12453);
xor XOR2 (N12456, N12455, N12249);
or OR4 (N12457, N12451, N6952, N2916, N7531);
nand NAND2 (N12458, N12449, N11428);
nand NAND2 (N12459, N12450, N4597);
xor XOR2 (N12460, N12459, N1396);
nor NOR2 (N12461, N12456, N4515);
buf BUF1 (N12462, N12454);
not NOT1 (N12463, N12460);
nand NAND3 (N12464, N12461, N9197, N11939);
or OR2 (N12465, N12464, N7075);
xor XOR2 (N12466, N12463, N11592);
not NOT1 (N12467, N12426);
nand NAND2 (N12468, N12465, N6982);
and AND4 (N12469, N12457, N8257, N4886, N1719);
nor NOR2 (N12470, N12452, N3159);
nand NAND2 (N12471, N12436, N6427);
buf BUF1 (N12472, N12444);
nand NAND3 (N12473, N12471, N4246, N11955);
nor NOR3 (N12474, N12472, N7314, N1290);
nor NOR3 (N12475, N12458, N8926, N8546);
buf BUF1 (N12476, N12466);
nor NOR4 (N12477, N12468, N7773, N5925, N9061);
not NOT1 (N12478, N12473);
buf BUF1 (N12479, N12477);
nand NAND4 (N12480, N12469, N9946, N11320, N9307);
nor NOR3 (N12481, N12467, N6043, N5892);
xor XOR2 (N12482, N12475, N6328);
nor NOR2 (N12483, N12470, N9601);
not NOT1 (N12484, N12439);
and AND3 (N12485, N12462, N808, N10174);
nor NOR2 (N12486, N12476, N10264);
nor NOR3 (N12487, N12483, N9089, N5764);
buf BUF1 (N12488, N12482);
nor NOR2 (N12489, N12474, N9608);
not NOT1 (N12490, N12480);
nor NOR2 (N12491, N12484, N6360);
xor XOR2 (N12492, N12485, N7414);
buf BUF1 (N12493, N12488);
nand NAND2 (N12494, N12492, N5222);
not NOT1 (N12495, N12491);
not NOT1 (N12496, N12494);
xor XOR2 (N12497, N12479, N6622);
nand NAND4 (N12498, N12478, N8613, N11409, N3153);
nand NAND4 (N12499, N12498, N8377, N11326, N3392);
not NOT1 (N12500, N12495);
or OR2 (N12501, N12493, N8698);
and AND4 (N12502, N12490, N4139, N1474, N6583);
not NOT1 (N12503, N12481);
nor NOR3 (N12504, N12487, N3865, N7936);
nand NAND2 (N12505, N12496, N99);
xor XOR2 (N12506, N12502, N12174);
nor NOR3 (N12507, N12506, N5050, N7254);
and AND3 (N12508, N12507, N7443, N7941);
nand NAND3 (N12509, N12486, N9403, N8144);
nor NOR3 (N12510, N12500, N4284, N6252);
nand NAND4 (N12511, N12504, N4493, N10532, N5418);
buf BUF1 (N12512, N12505);
not NOT1 (N12513, N12497);
and AND4 (N12514, N12503, N12069, N11019, N5421);
nor NOR4 (N12515, N12512, N6636, N2622, N4176);
not NOT1 (N12516, N12499);
not NOT1 (N12517, N12509);
nand NAND2 (N12518, N12517, N8564);
buf BUF1 (N12519, N12501);
or OR2 (N12520, N12518, N12089);
or OR4 (N12521, N12520, N3871, N9476, N4786);
or OR3 (N12522, N12516, N770, N11416);
nand NAND2 (N12523, N12513, N11786);
buf BUF1 (N12524, N12508);
and AND2 (N12525, N12524, N7812);
or OR2 (N12526, N12510, N5144);
not NOT1 (N12527, N12514);
not NOT1 (N12528, N12523);
nand NAND4 (N12529, N12515, N6362, N411, N8374);
or OR3 (N12530, N12528, N2581, N2721);
xor XOR2 (N12531, N12525, N4880);
nand NAND3 (N12532, N12529, N8176, N159);
nand NAND3 (N12533, N12526, N9221, N4133);
and AND3 (N12534, N12519, N11882, N8722);
nor NOR2 (N12535, N12527, N5363);
and AND4 (N12536, N12522, N2891, N8383, N2473);
not NOT1 (N12537, N12521);
nor NOR4 (N12538, N12532, N8662, N11008, N1888);
xor XOR2 (N12539, N12533, N11681);
nor NOR3 (N12540, N12534, N881, N242);
or OR2 (N12541, N12537, N7432);
or OR4 (N12542, N12540, N6448, N7156, N9744);
nor NOR3 (N12543, N12541, N10618, N1858);
or OR3 (N12544, N12511, N672, N7264);
not NOT1 (N12545, N12543);
xor XOR2 (N12546, N12542, N6907);
nand NAND2 (N12547, N12530, N5381);
xor XOR2 (N12548, N12536, N1677);
buf BUF1 (N12549, N12547);
nand NAND3 (N12550, N12538, N4937, N9856);
and AND2 (N12551, N12548, N7888);
not NOT1 (N12552, N12531);
buf BUF1 (N12553, N12551);
not NOT1 (N12554, N12549);
buf BUF1 (N12555, N12489);
xor XOR2 (N12556, N12544, N11142);
not NOT1 (N12557, N12554);
or OR4 (N12558, N12545, N10529, N7076, N10388);
not NOT1 (N12559, N12546);
nor NOR4 (N12560, N12552, N5647, N251, N1266);
xor XOR2 (N12561, N12555, N1384);
and AND3 (N12562, N12558, N595, N5746);
nor NOR3 (N12563, N12559, N2029, N9749);
nand NAND3 (N12564, N12539, N12162, N11882);
nor NOR3 (N12565, N12561, N8042, N5077);
nand NAND2 (N12566, N12565, N11909);
nand NAND2 (N12567, N12535, N506);
or OR3 (N12568, N12563, N4009, N12535);
nand NAND4 (N12569, N12567, N4604, N2339, N10866);
nand NAND3 (N12570, N12553, N7908, N5058);
and AND3 (N12571, N12556, N12099, N9209);
or OR3 (N12572, N12571, N12567, N11506);
buf BUF1 (N12573, N12550);
and AND4 (N12574, N12566, N7401, N2655, N6740);
or OR3 (N12575, N12557, N7336, N11410);
buf BUF1 (N12576, N12569);
or OR4 (N12577, N12568, N8607, N10165, N10118);
nor NOR2 (N12578, N12572, N8916);
nor NOR3 (N12579, N12562, N4229, N11221);
and AND2 (N12580, N12576, N6683);
and AND2 (N12581, N12580, N3525);
xor XOR2 (N12582, N12581, N4351);
xor XOR2 (N12583, N12560, N4870);
nand NAND3 (N12584, N12577, N9646, N2538);
not NOT1 (N12585, N12575);
nor NOR4 (N12586, N12570, N2924, N3287, N7540);
and AND2 (N12587, N12586, N4303);
xor XOR2 (N12588, N12585, N9259);
not NOT1 (N12589, N12578);
nand NAND4 (N12590, N12582, N8219, N5562, N11686);
nor NOR4 (N12591, N12579, N7289, N6149, N12421);
nor NOR2 (N12592, N12589, N455);
buf BUF1 (N12593, N12592);
nand NAND3 (N12594, N12564, N7334, N3581);
or OR2 (N12595, N12588, N1743);
xor XOR2 (N12596, N12584, N10632);
and AND2 (N12597, N12595, N9386);
xor XOR2 (N12598, N12574, N963);
xor XOR2 (N12599, N12583, N10943);
nand NAND4 (N12600, N12587, N2636, N5, N12056);
buf BUF1 (N12601, N12590);
buf BUF1 (N12602, N12593);
buf BUF1 (N12603, N12602);
and AND3 (N12604, N12596, N10470, N924);
buf BUF1 (N12605, N12598);
buf BUF1 (N12606, N12591);
or OR4 (N12607, N12599, N3163, N382, N8962);
buf BUF1 (N12608, N12607);
nor NOR3 (N12609, N12597, N4349, N2284);
buf BUF1 (N12610, N12609);
nand NAND4 (N12611, N12594, N9329, N849, N10784);
buf BUF1 (N12612, N12605);
or OR4 (N12613, N12604, N2910, N2574, N455);
nand NAND4 (N12614, N12603, N9758, N10698, N6631);
nand NAND2 (N12615, N12601, N12411);
or OR2 (N12616, N12608, N9828);
nor NOR2 (N12617, N12616, N11242);
xor XOR2 (N12618, N12606, N12344);
and AND3 (N12619, N12614, N7961, N3418);
and AND2 (N12620, N12615, N10956);
and AND3 (N12621, N12613, N7456, N6747);
not NOT1 (N12622, N12619);
nor NOR2 (N12623, N12621, N3804);
and AND3 (N12624, N12573, N7955, N8029);
or OR4 (N12625, N12617, N11185, N1686, N700);
not NOT1 (N12626, N12600);
or OR4 (N12627, N12612, N7952, N11774, N965);
nand NAND4 (N12628, N12626, N4459, N1515, N7486);
and AND2 (N12629, N12625, N11607);
nand NAND2 (N12630, N12623, N2031);
nor NOR4 (N12631, N12630, N8261, N4901, N3350);
not NOT1 (N12632, N12622);
xor XOR2 (N12633, N12610, N2428);
or OR3 (N12634, N12624, N12192, N10873);
xor XOR2 (N12635, N12629, N1209);
not NOT1 (N12636, N12611);
and AND3 (N12637, N12636, N5241, N10206);
not NOT1 (N12638, N12635);
buf BUF1 (N12639, N12632);
nand NAND2 (N12640, N12618, N7359);
buf BUF1 (N12641, N12633);
xor XOR2 (N12642, N12627, N4361);
buf BUF1 (N12643, N12628);
or OR2 (N12644, N12634, N2511);
nand NAND4 (N12645, N12620, N6183, N9447, N8189);
nor NOR4 (N12646, N12644, N6922, N3260, N8975);
nor NOR2 (N12647, N12645, N6614);
not NOT1 (N12648, N12647);
nand NAND2 (N12649, N12643, N8939);
and AND2 (N12650, N12642, N12555);
buf BUF1 (N12651, N12641);
buf BUF1 (N12652, N12638);
not NOT1 (N12653, N12648);
and AND3 (N12654, N12639, N3518, N8915);
nand NAND2 (N12655, N12631, N12622);
nand NAND3 (N12656, N12654, N3694, N2800);
and AND2 (N12657, N12637, N1033);
nand NAND4 (N12658, N12657, N9011, N6551, N10141);
and AND3 (N12659, N12655, N7876, N12430);
buf BUF1 (N12660, N12652);
and AND2 (N12661, N12656, N2450);
or OR2 (N12662, N12651, N2020);
nor NOR4 (N12663, N12653, N1079, N9764, N8128);
and AND2 (N12664, N12659, N2879);
nand NAND4 (N12665, N12658, N5357, N12097, N9026);
not NOT1 (N12666, N12646);
nand NAND3 (N12667, N12664, N8187, N5996);
buf BUF1 (N12668, N12665);
not NOT1 (N12669, N12650);
not NOT1 (N12670, N12668);
and AND2 (N12671, N12667, N11269);
not NOT1 (N12672, N12662);
nor NOR3 (N12673, N12671, N3837, N3091);
buf BUF1 (N12674, N12666);
and AND4 (N12675, N12673, N9882, N12090, N12138);
nand NAND4 (N12676, N12675, N8017, N7728, N11284);
buf BUF1 (N12677, N12661);
xor XOR2 (N12678, N12640, N8668);
nand NAND3 (N12679, N12670, N6298, N10715);
xor XOR2 (N12680, N12678, N10960);
buf BUF1 (N12681, N12677);
and AND3 (N12682, N12681, N1969, N9496);
nand NAND4 (N12683, N12660, N4367, N735, N12289);
nor NOR4 (N12684, N12663, N9710, N10046, N1092);
not NOT1 (N12685, N12682);
nor NOR3 (N12686, N12674, N2358, N11886);
buf BUF1 (N12687, N12685);
or OR4 (N12688, N12676, N9614, N1896, N8386);
not NOT1 (N12689, N12669);
nor NOR2 (N12690, N12687, N6739);
not NOT1 (N12691, N12649);
xor XOR2 (N12692, N12680, N5741);
not NOT1 (N12693, N12684);
nand NAND2 (N12694, N12672, N10765);
and AND2 (N12695, N12679, N554);
buf BUF1 (N12696, N12688);
or OR4 (N12697, N12693, N5085, N9776, N12659);
buf BUF1 (N12698, N12692);
and AND4 (N12699, N12697, N5546, N2473, N7667);
and AND3 (N12700, N12683, N4348, N1599);
buf BUF1 (N12701, N12699);
or OR3 (N12702, N12701, N1015, N9545);
not NOT1 (N12703, N12698);
and AND2 (N12704, N12691, N3659);
nand NAND2 (N12705, N12700, N12685);
nor NOR4 (N12706, N12695, N1158, N9868, N3169);
buf BUF1 (N12707, N12703);
xor XOR2 (N12708, N12707, N130);
and AND2 (N12709, N12708, N6009);
xor XOR2 (N12710, N12689, N8398);
buf BUF1 (N12711, N12710);
nand NAND4 (N12712, N12711, N7624, N5089, N10276);
nor NOR2 (N12713, N12706, N5552);
xor XOR2 (N12714, N12713, N4954);
not NOT1 (N12715, N12714);
or OR3 (N12716, N12712, N8951, N1835);
nor NOR3 (N12717, N12704, N6455, N3736);
or OR2 (N12718, N12709, N3292);
xor XOR2 (N12719, N12686, N11935);
xor XOR2 (N12720, N12718, N7728);
and AND2 (N12721, N12690, N6763);
buf BUF1 (N12722, N12696);
or OR2 (N12723, N12705, N118);
xor XOR2 (N12724, N12717, N9048);
buf BUF1 (N12725, N12702);
or OR2 (N12726, N12720, N12514);
nor NOR3 (N12727, N12724, N4329, N10438);
buf BUF1 (N12728, N12716);
not NOT1 (N12729, N12726);
or OR3 (N12730, N12729, N11779, N3558);
not NOT1 (N12731, N12730);
nand NAND4 (N12732, N12722, N6325, N9194, N289);
not NOT1 (N12733, N12721);
or OR3 (N12734, N12733, N10136, N10279);
nor NOR3 (N12735, N12734, N8658, N5725);
nand NAND3 (N12736, N12715, N10212, N3959);
nor NOR4 (N12737, N12736, N4475, N6999, N11560);
or OR4 (N12738, N12719, N8621, N12640, N12149);
not NOT1 (N12739, N12727);
buf BUF1 (N12740, N12731);
xor XOR2 (N12741, N12723, N11932);
nand NAND3 (N12742, N12725, N884, N11534);
nor NOR2 (N12743, N12739, N406);
and AND4 (N12744, N12728, N9885, N3657, N4039);
and AND3 (N12745, N12694, N629, N5037);
xor XOR2 (N12746, N12740, N10994);
nand NAND3 (N12747, N12742, N826, N10782);
and AND2 (N12748, N12737, N10877);
nand NAND4 (N12749, N12743, N7533, N2901, N12465);
nor NOR2 (N12750, N12749, N6372);
and AND2 (N12751, N12732, N4904);
not NOT1 (N12752, N12741);
or OR4 (N12753, N12746, N4877, N6643, N7762);
or OR2 (N12754, N12747, N6136);
nor NOR2 (N12755, N12738, N2907);
buf BUF1 (N12756, N12751);
xor XOR2 (N12757, N12750, N31);
xor XOR2 (N12758, N12752, N10765);
xor XOR2 (N12759, N12758, N5909);
buf BUF1 (N12760, N12744);
not NOT1 (N12761, N12753);
not NOT1 (N12762, N12748);
buf BUF1 (N12763, N12745);
buf BUF1 (N12764, N12757);
xor XOR2 (N12765, N12759, N5765);
nand NAND4 (N12766, N12763, N7341, N1439, N7322);
not NOT1 (N12767, N12766);
xor XOR2 (N12768, N12760, N7556);
not NOT1 (N12769, N12767);
xor XOR2 (N12770, N12756, N9286);
not NOT1 (N12771, N12735);
not NOT1 (N12772, N12761);
buf BUF1 (N12773, N12770);
nor NOR4 (N12774, N12754, N1035, N10032, N4057);
nor NOR4 (N12775, N12773, N12612, N9863, N10242);
and AND4 (N12776, N12775, N4920, N5583, N11263);
or OR4 (N12777, N12769, N7009, N1483, N1192);
nor NOR2 (N12778, N12774, N10090);
buf BUF1 (N12779, N12776);
and AND3 (N12780, N12768, N1459, N5413);
nor NOR4 (N12781, N12771, N8708, N1413, N11828);
nor NOR2 (N12782, N12778, N1213);
buf BUF1 (N12783, N12765);
buf BUF1 (N12784, N12779);
not NOT1 (N12785, N12782);
xor XOR2 (N12786, N12762, N1229);
or OR2 (N12787, N12780, N3916);
and AND3 (N12788, N12772, N2663, N2441);
not NOT1 (N12789, N12786);
and AND4 (N12790, N12777, N2606, N11674, N10245);
not NOT1 (N12791, N12787);
buf BUF1 (N12792, N12791);
nor NOR4 (N12793, N12783, N10400, N5088, N8304);
nor NOR3 (N12794, N12781, N3418, N9290);
not NOT1 (N12795, N12792);
nand NAND2 (N12796, N12795, N12023);
and AND3 (N12797, N12788, N10161, N7882);
xor XOR2 (N12798, N12796, N1014);
not NOT1 (N12799, N12784);
xor XOR2 (N12800, N12798, N11051);
nand NAND2 (N12801, N12800, N2701);
not NOT1 (N12802, N12790);
xor XOR2 (N12803, N12785, N10137);
not NOT1 (N12804, N12764);
nand NAND3 (N12805, N12804, N9143, N4952);
xor XOR2 (N12806, N12803, N6562);
and AND3 (N12807, N12793, N6087, N4018);
xor XOR2 (N12808, N12806, N5740);
or OR3 (N12809, N12808, N8868, N4782);
nor NOR3 (N12810, N12809, N1809, N7777);
or OR2 (N12811, N12805, N11325);
nand NAND2 (N12812, N12807, N1248);
xor XOR2 (N12813, N12799, N4867);
xor XOR2 (N12814, N12789, N7061);
buf BUF1 (N12815, N12802);
or OR2 (N12816, N12815, N6186);
not NOT1 (N12817, N12816);
xor XOR2 (N12818, N12810, N4617);
buf BUF1 (N12819, N12817);
not NOT1 (N12820, N12801);
buf BUF1 (N12821, N12812);
xor XOR2 (N12822, N12819, N3047);
and AND2 (N12823, N12797, N2224);
and AND2 (N12824, N12823, N2737);
nand NAND3 (N12825, N12813, N10366, N4582);
nor NOR4 (N12826, N12825, N5584, N3656, N8662);
or OR3 (N12827, N12794, N11420, N8091);
xor XOR2 (N12828, N12824, N11219);
not NOT1 (N12829, N12821);
buf BUF1 (N12830, N12814);
nand NAND2 (N12831, N12827, N3462);
not NOT1 (N12832, N12829);
xor XOR2 (N12833, N12830, N468);
not NOT1 (N12834, N12820);
xor XOR2 (N12835, N12826, N8797);
buf BUF1 (N12836, N12818);
nand NAND3 (N12837, N12832, N3734, N6410);
nand NAND4 (N12838, N12833, N820, N1978, N12321);
buf BUF1 (N12839, N12831);
nor NOR4 (N12840, N12839, N12226, N4503, N10004);
not NOT1 (N12841, N12822);
not NOT1 (N12842, N12828);
and AND4 (N12843, N12840, N4093, N271, N5309);
nor NOR2 (N12844, N12838, N521);
not NOT1 (N12845, N12834);
and AND4 (N12846, N12844, N9832, N3974, N7008);
buf BUF1 (N12847, N12755);
or OR2 (N12848, N12811, N11452);
buf BUF1 (N12849, N12841);
not NOT1 (N12850, N12836);
buf BUF1 (N12851, N12835);
nand NAND2 (N12852, N12842, N10213);
xor XOR2 (N12853, N12837, N10502);
and AND3 (N12854, N12853, N10023, N4701);
buf BUF1 (N12855, N12845);
not NOT1 (N12856, N12854);
nor NOR3 (N12857, N12856, N4433, N4473);
buf BUF1 (N12858, N12847);
and AND4 (N12859, N12855, N2260, N8948, N6000);
not NOT1 (N12860, N12850);
not NOT1 (N12861, N12857);
not NOT1 (N12862, N12851);
xor XOR2 (N12863, N12861, N5155);
xor XOR2 (N12864, N12862, N4500);
nand NAND4 (N12865, N12848, N7527, N2652, N3290);
nand NAND4 (N12866, N12843, N9336, N10586, N7692);
and AND4 (N12867, N12860, N6548, N9527, N819);
or OR4 (N12868, N12867, N9512, N11958, N7348);
not NOT1 (N12869, N12852);
xor XOR2 (N12870, N12859, N5539);
xor XOR2 (N12871, N12868, N10513);
not NOT1 (N12872, N12846);
buf BUF1 (N12873, N12870);
nand NAND4 (N12874, N12866, N5245, N4980, N463);
and AND4 (N12875, N12863, N4371, N118, N5811);
xor XOR2 (N12876, N12872, N6636);
or OR4 (N12877, N12858, N2536, N6844, N1970);
or OR4 (N12878, N12874, N1329, N2905, N5292);
buf BUF1 (N12879, N12878);
not NOT1 (N12880, N12871);
nor NOR2 (N12881, N12864, N9335);
not NOT1 (N12882, N12849);
and AND3 (N12883, N12879, N7380, N12250);
not NOT1 (N12884, N12873);
and AND3 (N12885, N12880, N10744, N4274);
and AND3 (N12886, N12884, N12766, N6605);
nor NOR3 (N12887, N12869, N12150, N11627);
or OR2 (N12888, N12865, N1278);
nor NOR3 (N12889, N12887, N3094, N10446);
nor NOR2 (N12890, N12876, N4929);
nand NAND4 (N12891, N12889, N3264, N1646, N12547);
not NOT1 (N12892, N12875);
and AND2 (N12893, N12892, N979);
or OR4 (N12894, N12881, N7656, N11946, N9123);
or OR2 (N12895, N12890, N12701);
nand NAND4 (N12896, N12893, N5262, N7680, N12587);
and AND3 (N12897, N12894, N1551, N12504);
and AND4 (N12898, N12882, N6334, N4559, N5123);
nor NOR2 (N12899, N12888, N4778);
or OR4 (N12900, N12897, N12218, N4454, N5705);
not NOT1 (N12901, N12885);
nor NOR3 (N12902, N12899, N6532, N11337);
not NOT1 (N12903, N12886);
and AND2 (N12904, N12883, N7124);
buf BUF1 (N12905, N12903);
nand NAND2 (N12906, N12891, N6339);
xor XOR2 (N12907, N12877, N10552);
or OR4 (N12908, N12895, N6187, N507, N4416);
nor NOR3 (N12909, N12906, N2240, N6013);
nor NOR3 (N12910, N12908, N4858, N7838);
nand NAND4 (N12911, N12910, N445, N1105, N7313);
and AND4 (N12912, N12901, N11069, N11109, N2289);
and AND2 (N12913, N12907, N4253);
and AND3 (N12914, N12912, N2949, N10827);
or OR2 (N12915, N12898, N8582);
nor NOR2 (N12916, N12896, N3967);
not NOT1 (N12917, N12900);
xor XOR2 (N12918, N12913, N9634);
buf BUF1 (N12919, N12914);
buf BUF1 (N12920, N12911);
and AND2 (N12921, N12917, N8781);
nor NOR4 (N12922, N12921, N614, N2707, N9262);
buf BUF1 (N12923, N12916);
nor NOR2 (N12924, N12909, N3153);
and AND3 (N12925, N12920, N8374, N3737);
not NOT1 (N12926, N12919);
not NOT1 (N12927, N12922);
buf BUF1 (N12928, N12924);
buf BUF1 (N12929, N12902);
xor XOR2 (N12930, N12928, N9172);
not NOT1 (N12931, N12926);
and AND3 (N12932, N12918, N4691, N1191);
xor XOR2 (N12933, N12932, N2806);
xor XOR2 (N12934, N12925, N727);
nor NOR2 (N12935, N12934, N7179);
nand NAND3 (N12936, N12904, N12682, N3741);
buf BUF1 (N12937, N12930);
or OR3 (N12938, N12905, N8505, N3525);
buf BUF1 (N12939, N12938);
nand NAND3 (N12940, N12936, N2778, N7792);
nor NOR4 (N12941, N12927, N1632, N5426, N8464);
nand NAND3 (N12942, N12915, N6980, N2017);
xor XOR2 (N12943, N12940, N9609);
xor XOR2 (N12944, N12923, N9373);
not NOT1 (N12945, N12935);
not NOT1 (N12946, N12943);
buf BUF1 (N12947, N12933);
not NOT1 (N12948, N12942);
xor XOR2 (N12949, N12937, N354);
nor NOR4 (N12950, N12945, N2697, N8931, N2746);
buf BUF1 (N12951, N12947);
nand NAND3 (N12952, N12948, N11789, N7536);
or OR2 (N12953, N12939, N11077);
xor XOR2 (N12954, N12946, N3372);
buf BUF1 (N12955, N12931);
and AND2 (N12956, N12929, N1431);
or OR2 (N12957, N12953, N4055);
or OR4 (N12958, N12954, N1297, N8244, N4395);
not NOT1 (N12959, N12944);
nor NOR4 (N12960, N12959, N11761, N10745, N242);
or OR3 (N12961, N12941, N5246, N3624);
not NOT1 (N12962, N12949);
not NOT1 (N12963, N12957);
nor NOR3 (N12964, N12958, N2283, N10670);
not NOT1 (N12965, N12963);
xor XOR2 (N12966, N12964, N10320);
and AND4 (N12967, N12952, N10832, N6806, N11308);
buf BUF1 (N12968, N12951);
xor XOR2 (N12969, N12968, N11736);
and AND4 (N12970, N12966, N11312, N12931, N10681);
nand NAND4 (N12971, N12969, N12135, N2164, N10914);
not NOT1 (N12972, N12961);
nand NAND3 (N12973, N12962, N3246, N11020);
not NOT1 (N12974, N12970);
buf BUF1 (N12975, N12960);
buf BUF1 (N12976, N12950);
xor XOR2 (N12977, N12971, N9869);
or OR3 (N12978, N12967, N11254, N1065);
nand NAND2 (N12979, N12965, N900);
not NOT1 (N12980, N12974);
nor NOR4 (N12981, N12956, N3405, N3953, N12727);
nand NAND3 (N12982, N12972, N12943, N10822);
nor NOR2 (N12983, N12973, N5077);
nor NOR3 (N12984, N12980, N9195, N1881);
or OR4 (N12985, N12982, N7515, N5923, N1462);
or OR3 (N12986, N12985, N4680, N3478);
nand NAND2 (N12987, N12978, N7783);
xor XOR2 (N12988, N12986, N4470);
not NOT1 (N12989, N12979);
buf BUF1 (N12990, N12988);
nand NAND3 (N12991, N12990, N10574, N9397);
buf BUF1 (N12992, N12987);
nor NOR3 (N12993, N12991, N5302, N11710);
or OR2 (N12994, N12976, N6160);
or OR4 (N12995, N12977, N2644, N1267, N3731);
or OR4 (N12996, N12983, N12910, N8923, N8034);
nor NOR3 (N12997, N12992, N12040, N6013);
nor NOR4 (N12998, N12994, N5066, N10786, N334);
or OR4 (N12999, N12995, N294, N745, N4195);
not NOT1 (N13000, N12981);
not NOT1 (N13001, N12975);
not NOT1 (N13002, N12998);
and AND4 (N13003, N13002, N908, N9883, N9924);
and AND2 (N13004, N12993, N3959);
xor XOR2 (N13005, N12996, N7330);
not NOT1 (N13006, N13000);
nand NAND2 (N13007, N13006, N5661);
and AND3 (N13008, N12997, N4684, N8077);
or OR3 (N13009, N12999, N12598, N7098);
nand NAND2 (N13010, N13004, N9319);
and AND4 (N13011, N13007, N367, N7167, N4028);
xor XOR2 (N13012, N13001, N5518);
and AND4 (N13013, N13010, N968, N3171, N9192);
not NOT1 (N13014, N12984);
buf BUF1 (N13015, N13009);
and AND4 (N13016, N13011, N11016, N8559, N12705);
nand NAND3 (N13017, N13013, N6072, N1346);
and AND4 (N13018, N13017, N11168, N1729, N3323);
not NOT1 (N13019, N13008);
nor NOR2 (N13020, N13014, N5131);
xor XOR2 (N13021, N12989, N3450);
buf BUF1 (N13022, N13005);
or OR3 (N13023, N13020, N8011, N5338);
or OR2 (N13024, N13021, N11740);
not NOT1 (N13025, N13015);
xor XOR2 (N13026, N13025, N11942);
or OR3 (N13027, N12955, N1457, N12602);
not NOT1 (N13028, N13023);
nand NAND4 (N13029, N13012, N4273, N7005, N3319);
and AND3 (N13030, N13026, N7771, N392);
or OR3 (N13031, N13019, N10522, N10015);
not NOT1 (N13032, N13029);
xor XOR2 (N13033, N13003, N1729);
nor NOR2 (N13034, N13024, N8883);
not NOT1 (N13035, N13034);
not NOT1 (N13036, N13018);
xor XOR2 (N13037, N13016, N11863);
buf BUF1 (N13038, N13036);
nor NOR2 (N13039, N13032, N5807);
and AND4 (N13040, N13027, N12441, N5407, N349);
and AND3 (N13041, N13033, N9556, N11791);
buf BUF1 (N13042, N13028);
or OR3 (N13043, N13041, N3371, N5858);
or OR2 (N13044, N13035, N781);
xor XOR2 (N13045, N13022, N6693);
nor NOR2 (N13046, N13045, N336);
and AND2 (N13047, N13040, N4500);
xor XOR2 (N13048, N13038, N4749);
nand NAND2 (N13049, N13043, N334);
buf BUF1 (N13050, N13044);
nor NOR3 (N13051, N13050, N9016, N11966);
not NOT1 (N13052, N13042);
xor XOR2 (N13053, N13051, N11073);
and AND3 (N13054, N13031, N1499, N9197);
buf BUF1 (N13055, N13048);
nor NOR3 (N13056, N13037, N7788, N5287);
nor NOR2 (N13057, N13055, N2205);
or OR4 (N13058, N13049, N9115, N3294, N5564);
and AND2 (N13059, N13056, N691);
nand NAND4 (N13060, N13058, N4113, N5223, N7914);
or OR4 (N13061, N13054, N11458, N7878, N11109);
buf BUF1 (N13062, N13046);
or OR4 (N13063, N13057, N1734, N4388, N6894);
nor NOR3 (N13064, N13053, N9120, N9311);
not NOT1 (N13065, N13063);
and AND2 (N13066, N13059, N3562);
buf BUF1 (N13067, N13047);
nand NAND2 (N13068, N13030, N11755);
not NOT1 (N13069, N13065);
or OR2 (N13070, N13060, N6043);
and AND3 (N13071, N13070, N12169, N8590);
nor NOR3 (N13072, N13064, N1055, N6585);
buf BUF1 (N13073, N13072);
xor XOR2 (N13074, N13069, N3025);
nand NAND4 (N13075, N13067, N10726, N2693, N3826);
nor NOR2 (N13076, N13073, N6128);
or OR3 (N13077, N13076, N1005, N12672);
nand NAND3 (N13078, N13074, N5849, N13032);
nand NAND2 (N13079, N13052, N6866);
nand NAND4 (N13080, N13039, N12885, N7286, N318);
nor NOR2 (N13081, N13075, N12936);
not NOT1 (N13082, N13079);
nor NOR3 (N13083, N13066, N964, N3756);
xor XOR2 (N13084, N13061, N643);
nor NOR4 (N13085, N13083, N6327, N1344, N5006);
xor XOR2 (N13086, N13082, N4901);
and AND3 (N13087, N13071, N9867, N4835);
xor XOR2 (N13088, N13068, N4787);
or OR2 (N13089, N13087, N4327);
not NOT1 (N13090, N13089);
and AND2 (N13091, N13086, N3955);
and AND3 (N13092, N13085, N12915, N7734);
and AND4 (N13093, N13092, N2030, N10056, N744);
nand NAND2 (N13094, N13084, N6162);
nor NOR4 (N13095, N13080, N10521, N2913, N8531);
nand NAND3 (N13096, N13088, N12929, N3563);
and AND2 (N13097, N13091, N1530);
nor NOR2 (N13098, N13096, N3055);
nor NOR4 (N13099, N13095, N2956, N7289, N9617);
xor XOR2 (N13100, N13077, N1551);
or OR4 (N13101, N13093, N2081, N496, N3808);
and AND4 (N13102, N13078, N6942, N12990, N5361);
and AND4 (N13103, N13098, N3745, N10174, N4974);
nand NAND3 (N13104, N13100, N2631, N4681);
buf BUF1 (N13105, N13097);
or OR3 (N13106, N13103, N8977, N6700);
xor XOR2 (N13107, N13099, N7730);
nor NOR2 (N13108, N13090, N5552);
and AND2 (N13109, N13062, N1);
xor XOR2 (N13110, N13108, N11895);
and AND2 (N13111, N13094, N10564);
or OR2 (N13112, N13110, N9232);
xor XOR2 (N13113, N13104, N6509);
xor XOR2 (N13114, N13107, N3780);
nand NAND2 (N13115, N13106, N6270);
not NOT1 (N13116, N13115);
buf BUF1 (N13117, N13081);
and AND3 (N13118, N13105, N1928, N13012);
not NOT1 (N13119, N13114);
not NOT1 (N13120, N13117);
and AND4 (N13121, N13113, N2378, N3244, N2642);
xor XOR2 (N13122, N13101, N6142);
nor NOR2 (N13123, N13109, N8589);
nand NAND2 (N13124, N13121, N3455);
not NOT1 (N13125, N13124);
buf BUF1 (N13126, N13125);
nand NAND4 (N13127, N13112, N9259, N9874, N4639);
or OR4 (N13128, N13120, N5294, N11265, N499);
buf BUF1 (N13129, N13126);
xor XOR2 (N13130, N13116, N9084);
not NOT1 (N13131, N13128);
nor NOR4 (N13132, N13111, N5597, N2339, N1443);
and AND4 (N13133, N13127, N12524, N4787, N8436);
xor XOR2 (N13134, N13131, N10765);
nor NOR2 (N13135, N13118, N7594);
xor XOR2 (N13136, N13133, N2843);
or OR2 (N13137, N13134, N12543);
nand NAND2 (N13138, N13130, N9718);
and AND3 (N13139, N13123, N5752, N4724);
nand NAND3 (N13140, N13139, N8207, N4626);
and AND2 (N13141, N13119, N5754);
and AND2 (N13142, N13138, N6428);
nand NAND3 (N13143, N13135, N8622, N3714);
nand NAND4 (N13144, N13122, N10679, N2270, N3664);
xor XOR2 (N13145, N13143, N6656);
and AND3 (N13146, N13141, N3300, N10701);
nor NOR3 (N13147, N13145, N3752, N9744);
nand NAND4 (N13148, N13142, N11658, N12245, N1615);
xor XOR2 (N13149, N13147, N7951);
and AND2 (N13150, N13146, N7652);
nor NOR2 (N13151, N13140, N9074);
or OR4 (N13152, N13151, N7983, N6293, N3559);
buf BUF1 (N13153, N13129);
not NOT1 (N13154, N13132);
and AND2 (N13155, N13144, N8005);
nand NAND2 (N13156, N13149, N4029);
buf BUF1 (N13157, N13155);
nand NAND3 (N13158, N13157, N737, N5510);
xor XOR2 (N13159, N13137, N714);
not NOT1 (N13160, N13136);
nor NOR2 (N13161, N13156, N8979);
and AND2 (N13162, N13161, N3452);
not NOT1 (N13163, N13160);
and AND3 (N13164, N13153, N10949, N1395);
nor NOR4 (N13165, N13163, N11761, N4926, N11821);
buf BUF1 (N13166, N13159);
or OR4 (N13167, N13166, N5000, N6026, N10454);
or OR3 (N13168, N13148, N3698, N12282);
not NOT1 (N13169, N13162);
or OR2 (N13170, N13150, N9961);
nor NOR4 (N13171, N13164, N7129, N11612, N8781);
nand NAND2 (N13172, N13165, N10719);
or OR3 (N13173, N13167, N5269, N744);
nand NAND3 (N13174, N13173, N4784, N1378);
not NOT1 (N13175, N13152);
nand NAND3 (N13176, N13171, N10975, N12600);
and AND2 (N13177, N13174, N591);
nand NAND4 (N13178, N13154, N2988, N3216, N4855);
and AND4 (N13179, N13172, N7725, N2829, N4818);
or OR2 (N13180, N13178, N1069);
nor NOR3 (N13181, N13168, N8121, N5342);
xor XOR2 (N13182, N13180, N891);
not NOT1 (N13183, N13158);
or OR4 (N13184, N13169, N393, N8406, N611);
and AND3 (N13185, N13170, N4043, N9149);
and AND3 (N13186, N13176, N10758, N306);
not NOT1 (N13187, N13185);
not NOT1 (N13188, N13175);
nor NOR4 (N13189, N13188, N7775, N10897, N492);
nor NOR4 (N13190, N13186, N1143, N13109, N2933);
and AND4 (N13191, N13102, N12357, N10136, N13019);
nor NOR2 (N13192, N13179, N7367);
not NOT1 (N13193, N13187);
and AND3 (N13194, N13177, N3253, N7925);
or OR4 (N13195, N13189, N4715, N11136, N3382);
buf BUF1 (N13196, N13184);
buf BUF1 (N13197, N13191);
nand NAND3 (N13198, N13195, N7436, N10280);
and AND4 (N13199, N13192, N9015, N8023, N573);
nor NOR3 (N13200, N13182, N3101, N10414);
nand NAND3 (N13201, N13193, N3616, N8434);
nor NOR2 (N13202, N13190, N10804);
not NOT1 (N13203, N13202);
nand NAND4 (N13204, N13181, N10936, N916, N7689);
not NOT1 (N13205, N13201);
xor XOR2 (N13206, N13205, N516);
or OR3 (N13207, N13197, N5984, N4550);
or OR2 (N13208, N13203, N345);
nand NAND4 (N13209, N13199, N7759, N3776, N251);
or OR3 (N13210, N13194, N11677, N2706);
nor NOR2 (N13211, N13209, N12584);
buf BUF1 (N13212, N13183);
and AND3 (N13213, N13198, N8423, N12673);
buf BUF1 (N13214, N13200);
not NOT1 (N13215, N13211);
xor XOR2 (N13216, N13208, N3235);
nand NAND4 (N13217, N13196, N2482, N3846, N2254);
xor XOR2 (N13218, N13210, N8503);
xor XOR2 (N13219, N13206, N3526);
nor NOR4 (N13220, N13214, N12734, N2383, N7642);
buf BUF1 (N13221, N13216);
xor XOR2 (N13222, N13217, N1345);
not NOT1 (N13223, N13219);
and AND4 (N13224, N13222, N9551, N679, N13183);
buf BUF1 (N13225, N13212);
xor XOR2 (N13226, N13225, N6668);
buf BUF1 (N13227, N13223);
or OR4 (N13228, N13213, N8234, N5621, N1980);
buf BUF1 (N13229, N13204);
or OR2 (N13230, N13220, N8447);
not NOT1 (N13231, N13227);
or OR2 (N13232, N13218, N2011);
xor XOR2 (N13233, N13231, N260);
nor NOR4 (N13234, N13229, N6564, N12376, N123);
nand NAND3 (N13235, N13221, N11061, N7401);
nor NOR4 (N13236, N13233, N8705, N9142, N9307);
and AND2 (N13237, N13224, N13202);
nor NOR3 (N13238, N13228, N625, N6188);
or OR4 (N13239, N13237, N4512, N8848, N10676);
nand NAND2 (N13240, N13234, N10160);
nand NAND4 (N13241, N13232, N5366, N4994, N12399);
and AND4 (N13242, N13236, N5552, N7065, N8390);
and AND3 (N13243, N13215, N8195, N3608);
xor XOR2 (N13244, N13241, N9154);
nor NOR2 (N13245, N13230, N8456);
nor NOR3 (N13246, N13242, N6593, N10229);
not NOT1 (N13247, N13238);
and AND3 (N13248, N13244, N6991, N6491);
and AND2 (N13249, N13207, N3609);
nand NAND3 (N13250, N13246, N12974, N12381);
nand NAND2 (N13251, N13248, N6132);
and AND3 (N13252, N13247, N12415, N8746);
xor XOR2 (N13253, N13252, N11507);
not NOT1 (N13254, N13235);
nand NAND4 (N13255, N13240, N4031, N74, N3712);
nor NOR2 (N13256, N13249, N12330);
not NOT1 (N13257, N13239);
not NOT1 (N13258, N13257);
nor NOR2 (N13259, N13251, N10381);
and AND4 (N13260, N13256, N8679, N2316, N10081);
nor NOR3 (N13261, N13253, N4145, N3218);
xor XOR2 (N13262, N13258, N12545);
buf BUF1 (N13263, N13261);
buf BUF1 (N13264, N13245);
and AND3 (N13265, N13262, N7958, N12112);
not NOT1 (N13266, N13243);
xor XOR2 (N13267, N13250, N10468);
or OR3 (N13268, N13267, N11885, N1614);
nor NOR4 (N13269, N13259, N10428, N10834, N11990);
nand NAND3 (N13270, N13266, N6818, N3112);
not NOT1 (N13271, N13254);
buf BUF1 (N13272, N13271);
or OR3 (N13273, N13226, N9747, N5729);
buf BUF1 (N13274, N13270);
xor XOR2 (N13275, N13265, N4036);
nor NOR4 (N13276, N13275, N9815, N4179, N208);
and AND2 (N13277, N13269, N3927);
or OR3 (N13278, N13268, N4250, N4891);
xor XOR2 (N13279, N13277, N10479);
xor XOR2 (N13280, N13264, N2502);
or OR3 (N13281, N13260, N4580, N4014);
and AND4 (N13282, N13272, N1224, N7186, N2035);
and AND3 (N13283, N13273, N11970, N5765);
xor XOR2 (N13284, N13282, N7720);
or OR4 (N13285, N13281, N3171, N11275, N7638);
nand NAND2 (N13286, N13255, N7310);
nand NAND4 (N13287, N13274, N1839, N7988, N9490);
xor XOR2 (N13288, N13283, N3485);
buf BUF1 (N13289, N13280);
not NOT1 (N13290, N13278);
not NOT1 (N13291, N13288);
and AND4 (N13292, N13289, N3708, N9913, N10914);
not NOT1 (N13293, N13279);
buf BUF1 (N13294, N13263);
nand NAND4 (N13295, N13293, N5978, N7878, N1935);
or OR2 (N13296, N13286, N862);
or OR3 (N13297, N13291, N7808, N4281);
buf BUF1 (N13298, N13276);
xor XOR2 (N13299, N13298, N9111);
or OR4 (N13300, N13296, N6464, N9706, N9735);
buf BUF1 (N13301, N13284);
not NOT1 (N13302, N13285);
xor XOR2 (N13303, N13292, N3145);
buf BUF1 (N13304, N13302);
and AND3 (N13305, N13294, N247, N10291);
nor NOR2 (N13306, N13287, N4592);
or OR4 (N13307, N13295, N6497, N10763, N10510);
or OR4 (N13308, N13304, N1708, N11963, N1775);
not NOT1 (N13309, N13307);
or OR4 (N13310, N13309, N10102, N6408, N7073);
and AND4 (N13311, N13290, N12996, N8, N12448);
nor NOR4 (N13312, N13299, N8724, N11514, N5706);
not NOT1 (N13313, N13306);
nor NOR3 (N13314, N13297, N12961, N11168);
nand NAND4 (N13315, N13310, N13028, N12625, N12537);
and AND3 (N13316, N13312, N2459, N894);
nor NOR4 (N13317, N13311, N10062, N5645, N4427);
not NOT1 (N13318, N13308);
nor NOR4 (N13319, N13313, N7199, N11491, N1766);
buf BUF1 (N13320, N13305);
xor XOR2 (N13321, N13319, N12752);
nand NAND2 (N13322, N13317, N1683);
or OR2 (N13323, N13303, N13076);
xor XOR2 (N13324, N13318, N8731);
not NOT1 (N13325, N13301);
xor XOR2 (N13326, N13316, N3013);
or OR3 (N13327, N13323, N3678, N5724);
nor NOR4 (N13328, N13325, N8411, N7545, N2959);
not NOT1 (N13329, N13315);
or OR2 (N13330, N13300, N7281);
not NOT1 (N13331, N13321);
or OR3 (N13332, N13324, N5558, N10802);
and AND2 (N13333, N13329, N1092);
or OR2 (N13334, N13328, N7604);
nand NAND4 (N13335, N13332, N818, N6446, N4838);
buf BUF1 (N13336, N13326);
and AND4 (N13337, N13331, N1110, N9743, N8818);
nand NAND4 (N13338, N13334, N10670, N3268, N5810);
or OR4 (N13339, N13330, N11749, N9984, N7349);
or OR4 (N13340, N13333, N2758, N4496, N7960);
xor XOR2 (N13341, N13314, N3567);
not NOT1 (N13342, N13327);
not NOT1 (N13343, N13340);
or OR2 (N13344, N13322, N8161);
buf BUF1 (N13345, N13339);
not NOT1 (N13346, N13343);
or OR4 (N13347, N13336, N7895, N5097, N2776);
not NOT1 (N13348, N13337);
xor XOR2 (N13349, N13345, N2954);
and AND3 (N13350, N13342, N10943, N7153);
nand NAND2 (N13351, N13344, N11991);
not NOT1 (N13352, N13341);
nor NOR4 (N13353, N13350, N8306, N9185, N7736);
nand NAND3 (N13354, N13335, N2302, N8660);
or OR3 (N13355, N13354, N7780, N12283);
xor XOR2 (N13356, N13338, N5655);
and AND3 (N13357, N13349, N7091, N6813);
not NOT1 (N13358, N13355);
nand NAND4 (N13359, N13357, N8905, N5492, N5256);
not NOT1 (N13360, N13358);
buf BUF1 (N13361, N13351);
xor XOR2 (N13362, N13353, N9814);
and AND4 (N13363, N13348, N1594, N11692, N2011);
nand NAND4 (N13364, N13360, N6881, N6381, N12381);
and AND3 (N13365, N13346, N1040, N937);
xor XOR2 (N13366, N13362, N9610);
nor NOR2 (N13367, N13356, N7922);
xor XOR2 (N13368, N13366, N12884);
nand NAND4 (N13369, N13320, N790, N11763, N6000);
buf BUF1 (N13370, N13365);
and AND3 (N13371, N13368, N8890, N12543);
not NOT1 (N13372, N13359);
nor NOR4 (N13373, N13371, N10425, N9573, N9320);
buf BUF1 (N13374, N13363);
xor XOR2 (N13375, N13361, N10910);
nand NAND4 (N13376, N13373, N10447, N792, N4369);
buf BUF1 (N13377, N13367);
xor XOR2 (N13378, N13364, N7352);
not NOT1 (N13379, N13370);
not NOT1 (N13380, N13352);
buf BUF1 (N13381, N13375);
nand NAND3 (N13382, N13376, N1844, N390);
buf BUF1 (N13383, N13374);
buf BUF1 (N13384, N13347);
or OR4 (N13385, N13381, N4736, N3704, N3460);
xor XOR2 (N13386, N13384, N7061);
nor NOR4 (N13387, N13379, N8227, N7416, N6100);
nand NAND3 (N13388, N13377, N8985, N10649);
buf BUF1 (N13389, N13382);
xor XOR2 (N13390, N13369, N10456);
not NOT1 (N13391, N13380);
xor XOR2 (N13392, N13372, N4214);
nor NOR3 (N13393, N13392, N6030, N5055);
and AND2 (N13394, N13389, N11416);
nand NAND3 (N13395, N13394, N3408, N3980);
buf BUF1 (N13396, N13387);
nand NAND3 (N13397, N13390, N7536, N9134);
xor XOR2 (N13398, N13393, N2297);
not NOT1 (N13399, N13395);
or OR3 (N13400, N13383, N9516, N13300);
nand NAND3 (N13401, N13397, N5283, N2242);
nor NOR4 (N13402, N13385, N2717, N12622, N6077);
not NOT1 (N13403, N13391);
nor NOR2 (N13404, N13400, N4937);
nand NAND3 (N13405, N13396, N5438, N7965);
not NOT1 (N13406, N13386);
xor XOR2 (N13407, N13388, N5610);
nand NAND2 (N13408, N13402, N7629);
buf BUF1 (N13409, N13378);
nor NOR2 (N13410, N13408, N6676);
nor NOR3 (N13411, N13399, N717, N355);
not NOT1 (N13412, N13406);
nand NAND2 (N13413, N13403, N9197);
or OR3 (N13414, N13405, N8263, N9082);
or OR3 (N13415, N13404, N7593, N273);
not NOT1 (N13416, N13412);
nor NOR3 (N13417, N13410, N12932, N8266);
not NOT1 (N13418, N13414);
and AND3 (N13419, N13401, N3650, N10646);
not NOT1 (N13420, N13417);
nand NAND2 (N13421, N13413, N1207);
and AND4 (N13422, N13416, N4842, N11232, N577);
xor XOR2 (N13423, N13409, N8112);
nand NAND4 (N13424, N13418, N4574, N9166, N4628);
nor NOR4 (N13425, N13420, N9021, N9209, N10755);
buf BUF1 (N13426, N13411);
nand NAND2 (N13427, N13422, N4618);
not NOT1 (N13428, N13398);
nand NAND3 (N13429, N13426, N2790, N2248);
or OR4 (N13430, N13423, N4057, N11233, N6274);
nand NAND4 (N13431, N13425, N4797, N5450, N10716);
or OR3 (N13432, N13428, N6917, N5507);
nand NAND4 (N13433, N13407, N9582, N38, N4954);
buf BUF1 (N13434, N13424);
nand NAND4 (N13435, N13434, N9413, N6523, N634);
nor NOR3 (N13436, N13421, N13348, N5771);
nor NOR4 (N13437, N13427, N2299, N9874, N2722);
or OR3 (N13438, N13432, N7984, N1029);
xor XOR2 (N13439, N13430, N3591);
buf BUF1 (N13440, N13437);
not NOT1 (N13441, N13415);
or OR3 (N13442, N13441, N5799, N8028);
not NOT1 (N13443, N13433);
nor NOR4 (N13444, N13440, N3849, N7975, N4273);
nor NOR4 (N13445, N13419, N12692, N11707, N6007);
and AND3 (N13446, N13429, N8539, N2979);
nand NAND2 (N13447, N13431, N5399);
and AND3 (N13448, N13435, N2781, N13370);
nand NAND4 (N13449, N13445, N3988, N12694, N5540);
not NOT1 (N13450, N13444);
nor NOR4 (N13451, N13448, N972, N8030, N4001);
buf BUF1 (N13452, N13438);
or OR4 (N13453, N13446, N12265, N5000, N962);
or OR2 (N13454, N13442, N2276);
buf BUF1 (N13455, N13452);
nand NAND2 (N13456, N13454, N10034);
or OR4 (N13457, N13451, N12074, N991, N12723);
nand NAND3 (N13458, N13450, N10315, N5451);
not NOT1 (N13459, N13456);
nor NOR4 (N13460, N13457, N7744, N7278, N3921);
and AND2 (N13461, N13459, N6640);
nor NOR2 (N13462, N13443, N5062);
not NOT1 (N13463, N13460);
buf BUF1 (N13464, N13453);
nand NAND3 (N13465, N13449, N8413, N11930);
nor NOR3 (N13466, N13465, N7688, N2894);
not NOT1 (N13467, N13463);
xor XOR2 (N13468, N13439, N5260);
nor NOR3 (N13469, N13458, N3798, N2306);
xor XOR2 (N13470, N13455, N2547);
and AND2 (N13471, N13447, N7999);
buf BUF1 (N13472, N13471);
buf BUF1 (N13473, N13464);
nor NOR2 (N13474, N13462, N12578);
and AND2 (N13475, N13467, N8272);
not NOT1 (N13476, N13470);
and AND2 (N13477, N13476, N9933);
not NOT1 (N13478, N13473);
nand NAND3 (N13479, N13475, N9578, N8255);
nand NAND2 (N13480, N13479, N7935);
and AND4 (N13481, N13472, N1588, N2967, N9761);
nand NAND3 (N13482, N13480, N5961, N9657);
buf BUF1 (N13483, N13468);
xor XOR2 (N13484, N13482, N10963);
nand NAND2 (N13485, N13484, N9116);
and AND3 (N13486, N13474, N8894, N11679);
nor NOR4 (N13487, N13466, N12636, N2869, N79);
and AND2 (N13488, N13477, N12750);
xor XOR2 (N13489, N13488, N10082);
buf BUF1 (N13490, N13469);
nand NAND4 (N13491, N13461, N9869, N4575, N7418);
xor XOR2 (N13492, N13490, N1604);
not NOT1 (N13493, N13492);
and AND3 (N13494, N13436, N10706, N6432);
buf BUF1 (N13495, N13494);
and AND3 (N13496, N13478, N9839, N3628);
and AND4 (N13497, N13483, N2531, N2765, N10037);
not NOT1 (N13498, N13493);
or OR3 (N13499, N13485, N5886, N5051);
buf BUF1 (N13500, N13499);
not NOT1 (N13501, N13498);
and AND2 (N13502, N13481, N13333);
nand NAND3 (N13503, N13491, N9559, N4849);
or OR2 (N13504, N13497, N7155);
nor NOR2 (N13505, N13504, N9071);
buf BUF1 (N13506, N13505);
and AND2 (N13507, N13495, N7318);
or OR4 (N13508, N13506, N12664, N3813, N11184);
xor XOR2 (N13509, N13496, N2457);
xor XOR2 (N13510, N13502, N12208);
buf BUF1 (N13511, N13507);
xor XOR2 (N13512, N13500, N5435);
buf BUF1 (N13513, N13503);
and AND3 (N13514, N13489, N4686, N10437);
nor NOR4 (N13515, N13509, N8696, N4820, N7580);
not NOT1 (N13516, N13514);
and AND3 (N13517, N13508, N3527, N8759);
nor NOR3 (N13518, N13510, N11615, N13195);
nand NAND2 (N13519, N13487, N2166);
or OR4 (N13520, N13516, N10261, N11562, N4116);
nor NOR3 (N13521, N13501, N6086, N3147);
nand NAND3 (N13522, N13520, N13419, N9795);
buf BUF1 (N13523, N13519);
and AND2 (N13524, N13515, N9591);
nor NOR2 (N13525, N13517, N4927);
nand NAND2 (N13526, N13518, N3121);
nand NAND4 (N13527, N13523, N6550, N8098, N5866);
xor XOR2 (N13528, N13511, N2277);
and AND2 (N13529, N13524, N7012);
buf BUF1 (N13530, N13486);
not NOT1 (N13531, N13529);
or OR2 (N13532, N13531, N3814);
or OR3 (N13533, N13526, N7894, N5020);
nand NAND4 (N13534, N13512, N7308, N11004, N11602);
xor XOR2 (N13535, N13534, N8322);
nor NOR4 (N13536, N13533, N6716, N8264, N7268);
or OR2 (N13537, N13525, N12068);
nand NAND3 (N13538, N13527, N10166, N21);
nand NAND3 (N13539, N13522, N2564, N6936);
nand NAND2 (N13540, N13528, N8590);
buf BUF1 (N13541, N13538);
or OR2 (N13542, N13536, N3183);
and AND2 (N13543, N13513, N8194);
nor NOR4 (N13544, N13535, N13432, N4277, N13035);
buf BUF1 (N13545, N13544);
nand NAND2 (N13546, N13539, N1050);
and AND4 (N13547, N13521, N6509, N3610, N10967);
xor XOR2 (N13548, N13541, N13249);
nor NOR3 (N13549, N13545, N9910, N9667);
or OR2 (N13550, N13548, N7129);
not NOT1 (N13551, N13542);
nor NOR4 (N13552, N13530, N7303, N11124, N2531);
and AND3 (N13553, N13543, N4170, N8489);
buf BUF1 (N13554, N13546);
nor NOR2 (N13555, N13552, N13037);
buf BUF1 (N13556, N13547);
xor XOR2 (N13557, N13549, N2717);
xor XOR2 (N13558, N13555, N2512);
nor NOR2 (N13559, N13554, N2802);
and AND4 (N13560, N13551, N8242, N7958, N4917);
not NOT1 (N13561, N13532);
xor XOR2 (N13562, N13558, N1293);
buf BUF1 (N13563, N13560);
buf BUF1 (N13564, N13563);
xor XOR2 (N13565, N13550, N8206);
not NOT1 (N13566, N13540);
and AND2 (N13567, N13565, N3591);
nor NOR4 (N13568, N13566, N4667, N11229, N9401);
nand NAND2 (N13569, N13553, N10784);
not NOT1 (N13570, N13567);
xor XOR2 (N13571, N13559, N9613);
buf BUF1 (N13572, N13557);
and AND3 (N13573, N13569, N2005, N1736);
buf BUF1 (N13574, N13561);
not NOT1 (N13575, N13564);
nand NAND2 (N13576, N13573, N12955);
or OR3 (N13577, N13562, N4025, N9734);
or OR2 (N13578, N13575, N8297);
not NOT1 (N13579, N13572);
nand NAND3 (N13580, N13577, N6302, N1104);
buf BUF1 (N13581, N13537);
not NOT1 (N13582, N13581);
not NOT1 (N13583, N13582);
xor XOR2 (N13584, N13574, N1253);
or OR4 (N13585, N13579, N4032, N10878, N12006);
buf BUF1 (N13586, N13571);
not NOT1 (N13587, N13585);
and AND4 (N13588, N13570, N2195, N13329, N5198);
not NOT1 (N13589, N13578);
and AND4 (N13590, N13586, N6263, N2566, N3255);
buf BUF1 (N13591, N13568);
or OR3 (N13592, N13591, N3564, N6553);
xor XOR2 (N13593, N13590, N8108);
nor NOR3 (N13594, N13593, N11063, N2541);
xor XOR2 (N13595, N13588, N8087);
and AND4 (N13596, N13594, N1064, N9902, N9880);
buf BUF1 (N13597, N13584);
and AND2 (N13598, N13595, N2799);
buf BUF1 (N13599, N13592);
nor NOR4 (N13600, N13596, N534, N1712, N8428);
nor NOR4 (N13601, N13597, N5849, N8617, N9310);
xor XOR2 (N13602, N13576, N644);
not NOT1 (N13603, N13587);
not NOT1 (N13604, N13602);
or OR3 (N13605, N13599, N5929, N5295);
xor XOR2 (N13606, N13598, N4073);
not NOT1 (N13607, N13603);
and AND4 (N13608, N13604, N1108, N2409, N6263);
not NOT1 (N13609, N13580);
xor XOR2 (N13610, N13600, N4614);
and AND4 (N13611, N13556, N4220, N3138, N6198);
or OR3 (N13612, N13607, N6530, N11649);
xor XOR2 (N13613, N13606, N10226);
or OR2 (N13614, N13589, N6417);
xor XOR2 (N13615, N13614, N1893);
not NOT1 (N13616, N13612);
nand NAND3 (N13617, N13608, N2409, N2674);
not NOT1 (N13618, N13601);
and AND4 (N13619, N13615, N5259, N8054, N9138);
nor NOR2 (N13620, N13610, N6914);
not NOT1 (N13621, N13619);
nand NAND2 (N13622, N13611, N622);
and AND4 (N13623, N13622, N3554, N12744, N12177);
xor XOR2 (N13624, N13617, N1286);
buf BUF1 (N13625, N13613);
and AND2 (N13626, N13624, N11156);
or OR3 (N13627, N13609, N12983, N691);
or OR4 (N13628, N13616, N1852, N10250, N2784);
buf BUF1 (N13629, N13628);
nor NOR4 (N13630, N13629, N4363, N10197, N7198);
nor NOR4 (N13631, N13583, N10657, N10083, N12335);
nand NAND3 (N13632, N13625, N11915, N4549);
nand NAND2 (N13633, N13623, N7509);
nand NAND2 (N13634, N13632, N3244);
not NOT1 (N13635, N13627);
nor NOR4 (N13636, N13631, N13609, N11342, N3227);
and AND4 (N13637, N13626, N3760, N156, N8295);
nor NOR3 (N13638, N13621, N3787, N3696);
not NOT1 (N13639, N13635);
not NOT1 (N13640, N13634);
nand NAND2 (N13641, N13639, N5620);
nor NOR4 (N13642, N13637, N9355, N1594, N8986);
xor XOR2 (N13643, N13605, N4639);
and AND2 (N13644, N13618, N3898);
or OR2 (N13645, N13644, N10667);
buf BUF1 (N13646, N13636);
and AND3 (N13647, N13642, N10683, N9350);
and AND2 (N13648, N13633, N3288);
nand NAND4 (N13649, N13647, N12921, N4771, N12098);
buf BUF1 (N13650, N13640);
nor NOR4 (N13651, N13646, N12051, N537, N4608);
or OR3 (N13652, N13648, N8783, N3246);
not NOT1 (N13653, N13652);
xor XOR2 (N13654, N13638, N11676);
and AND2 (N13655, N13620, N11595);
and AND4 (N13656, N13643, N7867, N13516, N11404);
nor NOR2 (N13657, N13656, N11440);
or OR2 (N13658, N13650, N4970);
nor NOR2 (N13659, N13649, N12383);
not NOT1 (N13660, N13654);
nor NOR4 (N13661, N13658, N9332, N10493, N876);
buf BUF1 (N13662, N13661);
and AND4 (N13663, N13660, N4760, N3761, N8163);
xor XOR2 (N13664, N13663, N10446);
nand NAND2 (N13665, N13664, N8125);
or OR3 (N13666, N13653, N8129, N3763);
not NOT1 (N13667, N13662);
or OR3 (N13668, N13641, N11783, N5660);
nand NAND3 (N13669, N13665, N1369, N2741);
not NOT1 (N13670, N13651);
or OR2 (N13671, N13670, N5196);
xor XOR2 (N13672, N13666, N2863);
buf BUF1 (N13673, N13669);
and AND3 (N13674, N13659, N1666, N7002);
and AND2 (N13675, N13668, N9704);
or OR4 (N13676, N13673, N4736, N11973, N1925);
and AND4 (N13677, N13675, N3888, N7943, N1512);
xor XOR2 (N13678, N13630, N154);
xor XOR2 (N13679, N13655, N6585);
and AND2 (N13680, N13645, N4735);
not NOT1 (N13681, N13667);
xor XOR2 (N13682, N13657, N2850);
and AND4 (N13683, N13681, N10953, N12804, N1573);
nand NAND4 (N13684, N13674, N7792, N2360, N10793);
nor NOR3 (N13685, N13678, N1551, N3880);
or OR4 (N13686, N13684, N7632, N11166, N8800);
buf BUF1 (N13687, N13685);
and AND3 (N13688, N13683, N6910, N3026);
nand NAND3 (N13689, N13682, N7722, N748);
or OR4 (N13690, N13687, N2351, N4824, N5694);
or OR3 (N13691, N13676, N3814, N13111);
xor XOR2 (N13692, N13680, N9647);
not NOT1 (N13693, N13679);
buf BUF1 (N13694, N13693);
xor XOR2 (N13695, N13671, N6849);
or OR3 (N13696, N13686, N10103, N10395);
or OR4 (N13697, N13692, N8912, N1076, N396);
nor NOR4 (N13698, N13672, N13549, N6725, N672);
nor NOR3 (N13699, N13695, N5054, N9831);
nand NAND4 (N13700, N13691, N7563, N12716, N7912);
xor XOR2 (N13701, N13698, N1627);
nand NAND3 (N13702, N13701, N11187, N9027);
or OR4 (N13703, N13700, N1827, N3868, N2740);
nand NAND4 (N13704, N13690, N611, N11201, N3676);
or OR2 (N13705, N13702, N12425);
nand NAND3 (N13706, N13699, N9832, N11599);
or OR4 (N13707, N13706, N12744, N9377, N12811);
buf BUF1 (N13708, N13697);
nor NOR3 (N13709, N13705, N7465, N11025);
nand NAND2 (N13710, N13704, N3481);
nor NOR4 (N13711, N13710, N345, N3057, N10038);
nor NOR3 (N13712, N13708, N12922, N9970);
xor XOR2 (N13713, N13712, N12616);
nor NOR3 (N13714, N13677, N11159, N6650);
nand NAND2 (N13715, N13713, N2169);
xor XOR2 (N13716, N13696, N4177);
or OR3 (N13717, N13716, N8895, N12389);
nor NOR4 (N13718, N13714, N5896, N12716, N2669);
xor XOR2 (N13719, N13689, N3119);
not NOT1 (N13720, N13707);
nand NAND2 (N13721, N13688, N8898);
nor NOR3 (N13722, N13719, N11059, N12094);
xor XOR2 (N13723, N13717, N1742);
or OR3 (N13724, N13721, N12472, N7505);
nor NOR3 (N13725, N13715, N9317, N11187);
not NOT1 (N13726, N13722);
buf BUF1 (N13727, N13718);
or OR2 (N13728, N13726, N4570);
nor NOR4 (N13729, N13694, N11633, N3550, N5206);
or OR2 (N13730, N13703, N8199);
nand NAND2 (N13731, N13709, N10947);
buf BUF1 (N13732, N13711);
and AND3 (N13733, N13729, N11425, N7370);
buf BUF1 (N13734, N13731);
not NOT1 (N13735, N13723);
nor NOR3 (N13736, N13735, N10050, N10498);
nor NOR2 (N13737, N13733, N4758);
xor XOR2 (N13738, N13727, N6034);
xor XOR2 (N13739, N13737, N5791);
and AND2 (N13740, N13739, N2341);
nor NOR4 (N13741, N13724, N8325, N6424, N12878);
or OR2 (N13742, N13740, N4683);
buf BUF1 (N13743, N13734);
buf BUF1 (N13744, N13738);
nand NAND4 (N13745, N13742, N9286, N5551, N7000);
buf BUF1 (N13746, N13732);
nand NAND4 (N13747, N13720, N1506, N9596, N6665);
buf BUF1 (N13748, N13743);
or OR4 (N13749, N13747, N11832, N12277, N1722);
or OR3 (N13750, N13746, N10642, N1419);
nand NAND3 (N13751, N13748, N8402, N9918);
buf BUF1 (N13752, N13745);
not NOT1 (N13753, N13736);
and AND2 (N13754, N13750, N10856);
xor XOR2 (N13755, N13753, N47);
buf BUF1 (N13756, N13755);
or OR3 (N13757, N13725, N2651, N8180);
nand NAND2 (N13758, N13757, N11970);
and AND4 (N13759, N13749, N8606, N716, N6568);
not NOT1 (N13760, N13752);
buf BUF1 (N13761, N13741);
not NOT1 (N13762, N13759);
xor XOR2 (N13763, N13756, N6014);
nor NOR3 (N13764, N13754, N4047, N10747);
not NOT1 (N13765, N13728);
not NOT1 (N13766, N13764);
not NOT1 (N13767, N13765);
not NOT1 (N13768, N13744);
and AND4 (N13769, N13730, N13662, N6195, N2242);
and AND4 (N13770, N13769, N2903, N12488, N6441);
xor XOR2 (N13771, N13758, N12871);
nand NAND3 (N13772, N13767, N4176, N6525);
and AND4 (N13773, N13772, N13220, N12853, N12682);
xor XOR2 (N13774, N13761, N5680);
nand NAND3 (N13775, N13751, N2391, N3302);
not NOT1 (N13776, N13773);
and AND3 (N13777, N13770, N8019, N999);
and AND3 (N13778, N13768, N2874, N426);
or OR3 (N13779, N13776, N11258, N13159);
buf BUF1 (N13780, N13774);
nor NOR2 (N13781, N13762, N8989);
not NOT1 (N13782, N13763);
buf BUF1 (N13783, N13780);
and AND3 (N13784, N13760, N7570, N5728);
nor NOR3 (N13785, N13775, N2170, N13771);
not NOT1 (N13786, N11722);
nor NOR4 (N13787, N13782, N5120, N10575, N5837);
and AND2 (N13788, N13779, N3018);
not NOT1 (N13789, N13766);
buf BUF1 (N13790, N13781);
nor NOR3 (N13791, N13790, N12207, N7549);
buf BUF1 (N13792, N13786);
xor XOR2 (N13793, N13789, N8512);
and AND2 (N13794, N13787, N452);
xor XOR2 (N13795, N13785, N7321);
nand NAND4 (N13796, N13783, N7184, N4651, N9613);
and AND2 (N13797, N13791, N11088);
buf BUF1 (N13798, N13794);
nand NAND4 (N13799, N13798, N6534, N12785, N13629);
buf BUF1 (N13800, N13784);
not NOT1 (N13801, N13799);
buf BUF1 (N13802, N13793);
not NOT1 (N13803, N13792);
nor NOR2 (N13804, N13803, N3759);
xor XOR2 (N13805, N13788, N4639);
nand NAND4 (N13806, N13801, N8562, N7063, N7390);
nor NOR3 (N13807, N13777, N8545, N7939);
and AND2 (N13808, N13800, N5652);
xor XOR2 (N13809, N13808, N13528);
not NOT1 (N13810, N13802);
and AND2 (N13811, N13797, N6335);
xor XOR2 (N13812, N13805, N12184);
and AND4 (N13813, N13796, N904, N10277, N4341);
and AND2 (N13814, N13812, N8867);
buf BUF1 (N13815, N13807);
xor XOR2 (N13816, N13809, N8715);
nor NOR4 (N13817, N13795, N8845, N13020, N9527);
nor NOR3 (N13818, N13817, N269, N570);
buf BUF1 (N13819, N13816);
nand NAND4 (N13820, N13818, N155, N10178, N3382);
xor XOR2 (N13821, N13806, N10516);
buf BUF1 (N13822, N13810);
and AND4 (N13823, N13819, N10009, N9854, N6753);
nor NOR2 (N13824, N13814, N9500);
nand NAND2 (N13825, N13822, N2860);
nand NAND3 (N13826, N13813, N12234, N3390);
or OR3 (N13827, N13811, N4035, N6670);
and AND2 (N13828, N13824, N2170);
or OR3 (N13829, N13826, N8839, N6095);
not NOT1 (N13830, N13827);
nand NAND2 (N13831, N13820, N11749);
nand NAND2 (N13832, N13828, N4209);
buf BUF1 (N13833, N13830);
or OR2 (N13834, N13829, N5071);
not NOT1 (N13835, N13831);
or OR3 (N13836, N13823, N4398, N6473);
nand NAND4 (N13837, N13832, N4130, N8084, N2129);
nand NAND3 (N13838, N13815, N13171, N11033);
or OR2 (N13839, N13821, N3634);
nor NOR2 (N13840, N13778, N9523);
and AND3 (N13841, N13835, N1507, N6715);
not NOT1 (N13842, N13833);
not NOT1 (N13843, N13838);
and AND2 (N13844, N13843, N4251);
nand NAND4 (N13845, N13844, N6059, N8081, N901);
nand NAND3 (N13846, N13840, N11553, N577);
not NOT1 (N13847, N13834);
nand NAND3 (N13848, N13804, N7428, N1297);
buf BUF1 (N13849, N13836);
xor XOR2 (N13850, N13845, N1348);
nor NOR4 (N13851, N13847, N2982, N4102, N4592);
xor XOR2 (N13852, N13849, N1304);
and AND4 (N13853, N13852, N9851, N8790, N8978);
xor XOR2 (N13854, N13853, N6209);
nand NAND2 (N13855, N13846, N11477);
or OR4 (N13856, N13841, N2378, N720, N12121);
not NOT1 (N13857, N13851);
and AND3 (N13858, N13825, N12958, N2516);
xor XOR2 (N13859, N13848, N931);
xor XOR2 (N13860, N13856, N6581);
buf BUF1 (N13861, N13858);
and AND4 (N13862, N13842, N1513, N10159, N4887);
or OR3 (N13863, N13861, N10202, N6941);
nand NAND4 (N13864, N13857, N558, N7017, N441);
nand NAND4 (N13865, N13860, N13075, N11890, N10555);
not NOT1 (N13866, N13859);
and AND3 (N13867, N13854, N12991, N11777);
nor NOR3 (N13868, N13866, N8526, N11005);
and AND2 (N13869, N13863, N11326);
xor XOR2 (N13870, N13855, N5182);
or OR3 (N13871, N13868, N7775, N90);
not NOT1 (N13872, N13869);
or OR4 (N13873, N13839, N4591, N9865, N1709);
xor XOR2 (N13874, N13871, N9918);
or OR2 (N13875, N13872, N12600);
xor XOR2 (N13876, N13874, N11583);
not NOT1 (N13877, N13867);
not NOT1 (N13878, N13864);
xor XOR2 (N13879, N13876, N5949);
or OR3 (N13880, N13875, N2993, N6892);
not NOT1 (N13881, N13865);
buf BUF1 (N13882, N13880);
xor XOR2 (N13883, N13850, N1876);
buf BUF1 (N13884, N13879);
nand NAND2 (N13885, N13870, N4669);
and AND4 (N13886, N13885, N10041, N5815, N12551);
not NOT1 (N13887, N13884);
or OR2 (N13888, N13862, N1269);
not NOT1 (N13889, N13837);
or OR2 (N13890, N13873, N3404);
nand NAND4 (N13891, N13882, N4038, N4999, N1609);
nor NOR2 (N13892, N13890, N3936);
and AND4 (N13893, N13887, N976, N5979, N1106);
and AND3 (N13894, N13888, N8235, N505);
or OR2 (N13895, N13886, N11611);
buf BUF1 (N13896, N13891);
buf BUF1 (N13897, N13894);
or OR3 (N13898, N13896, N2188, N7978);
nand NAND4 (N13899, N13897, N10595, N6316, N11239);
nor NOR3 (N13900, N13877, N7722, N990);
or OR3 (N13901, N13899, N12963, N1328);
xor XOR2 (N13902, N13889, N230);
and AND3 (N13903, N13898, N13900, N11479);
and AND3 (N13904, N11054, N13356, N1464);
and AND4 (N13905, N13892, N12961, N3025, N13358);
buf BUF1 (N13906, N13895);
and AND3 (N13907, N13904, N4979, N12780);
nor NOR3 (N13908, N13893, N5925, N2616);
not NOT1 (N13909, N13881);
buf BUF1 (N13910, N13903);
nand NAND2 (N13911, N13909, N2251);
nand NAND4 (N13912, N13901, N10759, N5807, N6036);
buf BUF1 (N13913, N13907);
xor XOR2 (N13914, N13883, N5166);
and AND3 (N13915, N13912, N4558, N8875);
and AND4 (N13916, N13878, N908, N10813, N1628);
and AND2 (N13917, N13914, N8912);
buf BUF1 (N13918, N13913);
buf BUF1 (N13919, N13905);
nor NOR2 (N13920, N13919, N5099);
buf BUF1 (N13921, N13902);
nor NOR2 (N13922, N13921, N3589);
nand NAND4 (N13923, N13915, N10632, N6998, N5665);
not NOT1 (N13924, N13918);
and AND4 (N13925, N13923, N860, N7700, N9980);
buf BUF1 (N13926, N13906);
not NOT1 (N13927, N13908);
nor NOR3 (N13928, N13926, N7938, N8417);
buf BUF1 (N13929, N13916);
not NOT1 (N13930, N13928);
nand NAND4 (N13931, N13927, N5300, N8752, N4455);
xor XOR2 (N13932, N13931, N6905);
buf BUF1 (N13933, N13925);
and AND3 (N13934, N13922, N9820, N5046);
nor NOR2 (N13935, N13932, N12012);
and AND3 (N13936, N13935, N9264, N7617);
nor NOR3 (N13937, N13929, N933, N3423);
xor XOR2 (N13938, N13910, N6605);
and AND3 (N13939, N13936, N4491, N2433);
buf BUF1 (N13940, N13939);
xor XOR2 (N13941, N13930, N1892);
buf BUF1 (N13942, N13920);
not NOT1 (N13943, N13937);
buf BUF1 (N13944, N13917);
not NOT1 (N13945, N13938);
not NOT1 (N13946, N13941);
not NOT1 (N13947, N13942);
not NOT1 (N13948, N13944);
or OR2 (N13949, N13934, N6738);
or OR2 (N13950, N13945, N1089);
or OR2 (N13951, N13933, N5629);
buf BUF1 (N13952, N13949);
xor XOR2 (N13953, N13950, N12470);
or OR2 (N13954, N13953, N4319);
and AND4 (N13955, N13924, N3444, N7468, N13931);
nand NAND2 (N13956, N13940, N6156);
nand NAND2 (N13957, N13955, N2787);
and AND4 (N13958, N13911, N1200, N7599, N10057);
xor XOR2 (N13959, N13947, N3837);
not NOT1 (N13960, N13946);
nor NOR3 (N13961, N13952, N5856, N7995);
or OR3 (N13962, N13951, N1689, N883);
not NOT1 (N13963, N13956);
nor NOR2 (N13964, N13958, N715);
and AND3 (N13965, N13961, N5187, N6187);
and AND3 (N13966, N13960, N10607, N13736);
not NOT1 (N13967, N13954);
or OR4 (N13968, N13948, N6676, N4008, N6036);
or OR3 (N13969, N13957, N7000, N4306);
nor NOR3 (N13970, N13965, N12804, N256);
nor NOR4 (N13971, N13966, N4922, N7219, N11730);
nor NOR3 (N13972, N13943, N3717, N5642);
xor XOR2 (N13973, N13967, N2644);
or OR2 (N13974, N13971, N10063);
and AND4 (N13975, N13968, N13856, N4621, N12178);
nand NAND4 (N13976, N13959, N11929, N4098, N1079);
nand NAND4 (N13977, N13962, N11530, N3690, N3677);
and AND2 (N13978, N13964, N11479);
xor XOR2 (N13979, N13976, N5258);
nand NAND2 (N13980, N13977, N11379);
and AND4 (N13981, N13974, N2249, N4323, N10210);
or OR4 (N13982, N13980, N9553, N9526, N4135);
nor NOR2 (N13983, N13979, N12112);
nand NAND2 (N13984, N13973, N10706);
buf BUF1 (N13985, N13982);
xor XOR2 (N13986, N13969, N10351);
not NOT1 (N13987, N13981);
xor XOR2 (N13988, N13975, N6917);
xor XOR2 (N13989, N13972, N8103);
nor NOR2 (N13990, N13986, N4102);
nand NAND2 (N13991, N13970, N5051);
or OR4 (N13992, N13963, N3061, N3930, N3167);
or OR3 (N13993, N13990, N8400, N6167);
and AND4 (N13994, N13989, N3464, N12854, N7564);
buf BUF1 (N13995, N13985);
or OR3 (N13996, N13978, N6601, N221);
nor NOR4 (N13997, N13987, N11839, N3755, N11630);
buf BUF1 (N13998, N13993);
and AND4 (N13999, N13998, N2340, N13241, N13011);
or OR4 (N14000, N13997, N3123, N12726, N8638);
xor XOR2 (N14001, N13991, N11082);
buf BUF1 (N14002, N13996);
buf BUF1 (N14003, N13999);
or OR3 (N14004, N13983, N3531, N12635);
or OR4 (N14005, N14000, N9296, N1484, N11936);
not NOT1 (N14006, N14003);
or OR3 (N14007, N13994, N3461, N10312);
and AND4 (N14008, N14006, N4311, N13279, N7862);
and AND4 (N14009, N14008, N11940, N12756, N8736);
nand NAND4 (N14010, N14001, N214, N5212, N3326);
nor NOR2 (N14011, N13995, N9117);
nor NOR3 (N14012, N14010, N1105, N12618);
nor NOR3 (N14013, N13984, N8820, N1741);
and AND4 (N14014, N14013, N8095, N6156, N7397);
or OR4 (N14015, N14007, N3681, N1915, N7483);
or OR4 (N14016, N14014, N98, N11295, N602);
or OR2 (N14017, N13988, N2639);
or OR3 (N14018, N14016, N8736, N2394);
nor NOR4 (N14019, N14009, N11748, N3469, N6930);
or OR3 (N14020, N14005, N2562, N2156);
buf BUF1 (N14021, N14015);
nand NAND3 (N14022, N14017, N5720, N9988);
xor XOR2 (N14023, N14012, N2133);
nor NOR2 (N14024, N14021, N5594);
and AND4 (N14025, N14019, N11366, N10722, N12453);
or OR4 (N14026, N14025, N10781, N9397, N11256);
xor XOR2 (N14027, N14002, N2425);
nor NOR4 (N14028, N14022, N9850, N13308, N10765);
not NOT1 (N14029, N14024);
xor XOR2 (N14030, N14020, N4978);
or OR3 (N14031, N14030, N214, N3216);
buf BUF1 (N14032, N14018);
or OR4 (N14033, N14031, N1316, N1301, N9095);
and AND4 (N14034, N14011, N2807, N7610, N11548);
and AND4 (N14035, N14034, N907, N8298, N8673);
or OR3 (N14036, N14032, N1918, N2609);
and AND2 (N14037, N14029, N12331);
nand NAND4 (N14038, N13992, N4836, N795, N7991);
xor XOR2 (N14039, N14037, N12140);
or OR3 (N14040, N14028, N9468, N12364);
xor XOR2 (N14041, N14038, N6040);
xor XOR2 (N14042, N14033, N850);
or OR4 (N14043, N14026, N4799, N6838, N13874);
and AND3 (N14044, N14035, N4827, N4392);
nand NAND2 (N14045, N14023, N3384);
buf BUF1 (N14046, N14040);
nand NAND4 (N14047, N14043, N11395, N13989, N5362);
xor XOR2 (N14048, N14047, N12679);
or OR4 (N14049, N14045, N1555, N3644, N6834);
not NOT1 (N14050, N14046);
buf BUF1 (N14051, N14048);
buf BUF1 (N14052, N14039);
xor XOR2 (N14053, N14050, N2408);
or OR4 (N14054, N14004, N4907, N13850, N8470);
nor NOR2 (N14055, N14053, N11091);
or OR3 (N14056, N14049, N2496, N12125);
nor NOR4 (N14057, N14036, N2399, N8422, N1476);
xor XOR2 (N14058, N14057, N11212);
nor NOR2 (N14059, N14051, N8538);
or OR2 (N14060, N14054, N9273);
nand NAND2 (N14061, N14044, N634);
buf BUF1 (N14062, N14060);
or OR4 (N14063, N14058, N921, N12967, N5105);
nor NOR3 (N14064, N14042, N10106, N3990);
and AND3 (N14065, N14059, N2571, N8225);
xor XOR2 (N14066, N14061, N11142);
not NOT1 (N14067, N14062);
not NOT1 (N14068, N14065);
not NOT1 (N14069, N14027);
not NOT1 (N14070, N14066);
and AND4 (N14071, N14068, N12266, N13771, N9009);
nand NAND4 (N14072, N14041, N2848, N7651, N7798);
xor XOR2 (N14073, N14056, N6761);
or OR2 (N14074, N14070, N10938);
or OR3 (N14075, N14067, N11209, N6409);
and AND3 (N14076, N14063, N5615, N5068);
not NOT1 (N14077, N14072);
xor XOR2 (N14078, N14075, N11772);
nand NAND3 (N14079, N14078, N6326, N12602);
nand NAND2 (N14080, N14077, N10786);
xor XOR2 (N14081, N14064, N3200);
nand NAND4 (N14082, N14073, N6689, N3833, N564);
buf BUF1 (N14083, N14069);
not NOT1 (N14084, N14083);
not NOT1 (N14085, N14052);
not NOT1 (N14086, N14079);
nand NAND3 (N14087, N14081, N13319, N644);
xor XOR2 (N14088, N14071, N5981);
nor NOR4 (N14089, N14086, N4934, N13701, N12399);
xor XOR2 (N14090, N14084, N7545);
nand NAND3 (N14091, N14074, N249, N4713);
and AND2 (N14092, N14082, N11627);
buf BUF1 (N14093, N14076);
xor XOR2 (N14094, N14088, N863);
or OR4 (N14095, N14087, N940, N8155, N7263);
buf BUF1 (N14096, N14094);
not NOT1 (N14097, N14092);
buf BUF1 (N14098, N14095);
nand NAND4 (N14099, N14093, N13660, N8092, N3647);
not NOT1 (N14100, N14055);
or OR3 (N14101, N14096, N14028, N4838);
buf BUF1 (N14102, N14089);
nor NOR3 (N14103, N14085, N13746, N714);
xor XOR2 (N14104, N14097, N5361);
buf BUF1 (N14105, N14102);
or OR3 (N14106, N14090, N3954, N10691);
not NOT1 (N14107, N14101);
not NOT1 (N14108, N14105);
and AND4 (N14109, N14091, N9190, N9935, N9138);
not NOT1 (N14110, N14103);
and AND3 (N14111, N14080, N7376, N711);
nand NAND4 (N14112, N14100, N534, N2564, N4364);
not NOT1 (N14113, N14109);
xor XOR2 (N14114, N14108, N1231);
not NOT1 (N14115, N14112);
or OR2 (N14116, N14113, N9790);
xor XOR2 (N14117, N14110, N12057);
buf BUF1 (N14118, N14099);
and AND4 (N14119, N14117, N7823, N13560, N7530);
buf BUF1 (N14120, N14114);
nand NAND4 (N14121, N14116, N1849, N5236, N516);
and AND4 (N14122, N14111, N8382, N4415, N9808);
buf BUF1 (N14123, N14119);
not NOT1 (N14124, N14120);
nor NOR2 (N14125, N14123, N1312);
nor NOR3 (N14126, N14118, N12930, N12313);
xor XOR2 (N14127, N14126, N11930);
and AND4 (N14128, N14115, N794, N6324, N11429);
buf BUF1 (N14129, N14098);
buf BUF1 (N14130, N14122);
buf BUF1 (N14131, N14104);
xor XOR2 (N14132, N14127, N1623);
not NOT1 (N14133, N14121);
not NOT1 (N14134, N14125);
and AND3 (N14135, N14134, N11799, N1703);
xor XOR2 (N14136, N14124, N1521);
and AND4 (N14137, N14131, N6442, N5440, N8394);
nand NAND3 (N14138, N14136, N10765, N6810);
nor NOR4 (N14139, N14132, N13971, N9851, N5442);
and AND2 (N14140, N14133, N4946);
buf BUF1 (N14141, N14139);
or OR2 (N14142, N14129, N11537);
xor XOR2 (N14143, N14141, N13393);
xor XOR2 (N14144, N14128, N4694);
buf BUF1 (N14145, N14144);
nor NOR3 (N14146, N14135, N4687, N5107);
buf BUF1 (N14147, N14130);
and AND4 (N14148, N14140, N3860, N8842, N11674);
xor XOR2 (N14149, N14143, N10800);
not NOT1 (N14150, N14107);
not NOT1 (N14151, N14145);
nor NOR2 (N14152, N14106, N13369);
or OR2 (N14153, N14151, N9186);
nand NAND3 (N14154, N14138, N756, N616);
nand NAND2 (N14155, N14137, N616);
and AND3 (N14156, N14146, N8419, N11241);
nand NAND2 (N14157, N14149, N13594);
and AND2 (N14158, N14156, N3313);
not NOT1 (N14159, N14152);
nor NOR3 (N14160, N14147, N4869, N9553);
nand NAND4 (N14161, N14148, N11696, N12904, N7167);
nand NAND2 (N14162, N14157, N9820);
nor NOR2 (N14163, N14161, N13456);
buf BUF1 (N14164, N14142);
nand NAND4 (N14165, N14150, N5687, N10171, N10370);
or OR3 (N14166, N14155, N4459, N8533);
not NOT1 (N14167, N14154);
buf BUF1 (N14168, N14166);
buf BUF1 (N14169, N14168);
xor XOR2 (N14170, N14158, N8178);
and AND2 (N14171, N14167, N11885);
and AND3 (N14172, N14170, N12596, N9647);
buf BUF1 (N14173, N14171);
and AND2 (N14174, N14173, N5005);
nor NOR2 (N14175, N14165, N2870);
or OR3 (N14176, N14162, N6025, N12079);
or OR2 (N14177, N14169, N2190);
not NOT1 (N14178, N14174);
nor NOR4 (N14179, N14153, N14159, N6238, N13978);
nor NOR3 (N14180, N11864, N8601, N207);
nand NAND2 (N14181, N14177, N3164);
nor NOR3 (N14182, N14160, N3959, N2696);
not NOT1 (N14183, N14176);
xor XOR2 (N14184, N14182, N6633);
nand NAND2 (N14185, N14175, N1031);
xor XOR2 (N14186, N14183, N8929);
nand NAND4 (N14187, N14180, N13401, N3210, N10812);
nand NAND4 (N14188, N14172, N12085, N13451, N12073);
not NOT1 (N14189, N14163);
or OR4 (N14190, N14181, N11394, N3063, N4590);
and AND2 (N14191, N14186, N13323);
nor NOR4 (N14192, N14190, N7449, N10794, N2368);
or OR2 (N14193, N14191, N8648);
buf BUF1 (N14194, N14179);
nand NAND2 (N14195, N14192, N6064);
nand NAND4 (N14196, N14193, N5731, N11473, N6973);
not NOT1 (N14197, N14188);
not NOT1 (N14198, N14189);
buf BUF1 (N14199, N14198);
nand NAND3 (N14200, N14184, N731, N13747);
xor XOR2 (N14201, N14197, N2552);
nor NOR3 (N14202, N14196, N11433, N10796);
not NOT1 (N14203, N14199);
not NOT1 (N14204, N14187);
not NOT1 (N14205, N14201);
xor XOR2 (N14206, N14195, N2795);
and AND3 (N14207, N14204, N316, N3825);
buf BUF1 (N14208, N14164);
xor XOR2 (N14209, N14206, N3392);
nor NOR2 (N14210, N14208, N2133);
and AND2 (N14211, N14178, N3195);
xor XOR2 (N14212, N14202, N5715);
xor XOR2 (N14213, N14205, N1919);
nor NOR2 (N14214, N14213, N83);
or OR4 (N14215, N14214, N10825, N10166, N11880);
xor XOR2 (N14216, N14200, N6562);
and AND4 (N14217, N14209, N1969, N4401, N11173);
nor NOR3 (N14218, N14207, N2345, N3134);
xor XOR2 (N14219, N14217, N805);
buf BUF1 (N14220, N14219);
or OR3 (N14221, N14185, N7719, N8238);
or OR3 (N14222, N14211, N14130, N3890);
and AND3 (N14223, N14216, N2240, N2306);
xor XOR2 (N14224, N14215, N9166);
nor NOR4 (N14225, N14203, N1218, N4823, N6223);
nor NOR3 (N14226, N14210, N11192, N2147);
or OR4 (N14227, N14218, N4665, N8948, N11794);
and AND3 (N14228, N14212, N3926, N7734);
and AND3 (N14229, N14225, N11190, N12331);
xor XOR2 (N14230, N14222, N7877);
buf BUF1 (N14231, N14223);
not NOT1 (N14232, N14229);
nand NAND2 (N14233, N14226, N4302);
nor NOR2 (N14234, N14227, N11812);
nor NOR3 (N14235, N14221, N8250, N6600);
nor NOR4 (N14236, N14220, N889, N5855, N3793);
not NOT1 (N14237, N14235);
and AND3 (N14238, N14228, N5715, N420);
and AND2 (N14239, N14236, N11500);
xor XOR2 (N14240, N14234, N3132);
buf BUF1 (N14241, N14238);
nor NOR2 (N14242, N14241, N10130);
and AND3 (N14243, N14231, N5116, N5777);
or OR3 (N14244, N14233, N9618, N2645);
nand NAND3 (N14245, N14242, N6504, N11334);
xor XOR2 (N14246, N14239, N2841);
nand NAND4 (N14247, N14246, N13100, N5703, N1359);
nor NOR3 (N14248, N14244, N13945, N4097);
buf BUF1 (N14249, N14224);
xor XOR2 (N14250, N14230, N6605);
buf BUF1 (N14251, N14237);
and AND4 (N14252, N14249, N3542, N923, N7989);
or OR4 (N14253, N14252, N4057, N13877, N568);
buf BUF1 (N14254, N14248);
not NOT1 (N14255, N14250);
not NOT1 (N14256, N14247);
nor NOR4 (N14257, N14245, N5359, N8376, N11209);
nor NOR3 (N14258, N14243, N4584, N2855);
and AND3 (N14259, N14258, N13267, N9406);
or OR2 (N14260, N14194, N9047);
not NOT1 (N14261, N14253);
or OR4 (N14262, N14240, N1271, N7926, N13977);
or OR2 (N14263, N14256, N9539);
not NOT1 (N14264, N14251);
nand NAND2 (N14265, N14254, N492);
xor XOR2 (N14266, N14232, N4850);
not NOT1 (N14267, N14259);
and AND2 (N14268, N14264, N1478);
nand NAND4 (N14269, N14255, N7500, N7571, N12598);
or OR2 (N14270, N14260, N5021);
nand NAND2 (N14271, N14266, N2326);
or OR4 (N14272, N14271, N12007, N9756, N4229);
buf BUF1 (N14273, N14268);
xor XOR2 (N14274, N14261, N738);
and AND4 (N14275, N14262, N12669, N14150, N13325);
not NOT1 (N14276, N14257);
xor XOR2 (N14277, N14267, N12193);
or OR4 (N14278, N14263, N11386, N10892, N3139);
buf BUF1 (N14279, N14276);
or OR4 (N14280, N14265, N12531, N11086, N5716);
nor NOR4 (N14281, N14275, N12913, N7697, N4674);
not NOT1 (N14282, N14269);
and AND2 (N14283, N14277, N11174);
nand NAND2 (N14284, N14280, N2419);
nand NAND3 (N14285, N14272, N2045, N7705);
nand NAND3 (N14286, N14279, N2718, N6578);
not NOT1 (N14287, N14282);
not NOT1 (N14288, N14274);
and AND2 (N14289, N14281, N4102);
nand NAND2 (N14290, N14270, N1848);
buf BUF1 (N14291, N14286);
xor XOR2 (N14292, N14285, N4122);
nand NAND2 (N14293, N14289, N6612);
nor NOR2 (N14294, N14273, N3110);
nor NOR2 (N14295, N14291, N9136);
nor NOR2 (N14296, N14284, N9927);
xor XOR2 (N14297, N14294, N7812);
nand NAND3 (N14298, N14287, N12696, N9689);
xor XOR2 (N14299, N14292, N10505);
and AND3 (N14300, N14296, N2910, N9763);
nand NAND4 (N14301, N14278, N7880, N5366, N4194);
nand NAND3 (N14302, N14299, N3341, N5584);
xor XOR2 (N14303, N14302, N10744);
buf BUF1 (N14304, N14295);
or OR2 (N14305, N14298, N11220);
and AND4 (N14306, N14293, N1308, N3226, N7644);
and AND2 (N14307, N14283, N9171);
or OR3 (N14308, N14306, N625, N10418);
and AND4 (N14309, N14305, N9977, N1814, N10242);
or OR3 (N14310, N14308, N5024, N7496);
nor NOR2 (N14311, N14301, N11294);
nand NAND3 (N14312, N14300, N8471, N8856);
not NOT1 (N14313, N14288);
buf BUF1 (N14314, N14313);
nand NAND4 (N14315, N14290, N7551, N4637, N6395);
nor NOR4 (N14316, N14311, N6619, N5715, N5374);
xor XOR2 (N14317, N14316, N1403);
not NOT1 (N14318, N14303);
nor NOR4 (N14319, N14318, N5449, N5522, N5710);
nand NAND3 (N14320, N14310, N12299, N8970);
xor XOR2 (N14321, N14304, N7152);
nor NOR2 (N14322, N14319, N13946);
or OR3 (N14323, N14315, N8932, N6411);
and AND2 (N14324, N14297, N11733);
not NOT1 (N14325, N14309);
xor XOR2 (N14326, N14322, N7154);
or OR2 (N14327, N14321, N2655);
xor XOR2 (N14328, N14327, N7806);
or OR4 (N14329, N14323, N7746, N13350, N7717);
not NOT1 (N14330, N14320);
not NOT1 (N14331, N14324);
not NOT1 (N14332, N14331);
or OR3 (N14333, N14312, N4430, N9492);
buf BUF1 (N14334, N14329);
nor NOR2 (N14335, N14326, N5365);
nor NOR4 (N14336, N14335, N6459, N2396, N8644);
or OR3 (N14337, N14333, N7077, N8892);
nand NAND3 (N14338, N14334, N12005, N9515);
xor XOR2 (N14339, N14336, N7519);
nor NOR4 (N14340, N14314, N3066, N10880, N2898);
not NOT1 (N14341, N14332);
not NOT1 (N14342, N14341);
not NOT1 (N14343, N14325);
or OR4 (N14344, N14337, N7950, N827, N2570);
nand NAND3 (N14345, N14338, N11757, N8115);
and AND4 (N14346, N14317, N3379, N13239, N6318);
nor NOR4 (N14347, N14342, N1980, N2157, N10402);
or OR4 (N14348, N14307, N5900, N2680, N3892);
nor NOR2 (N14349, N14340, N13273);
not NOT1 (N14350, N14328);
nand NAND2 (N14351, N14330, N13760);
and AND4 (N14352, N14350, N4559, N9175, N1421);
or OR3 (N14353, N14349, N6904, N460);
nand NAND4 (N14354, N14351, N9031, N7415, N13087);
nor NOR2 (N14355, N14343, N2958);
nor NOR2 (N14356, N14348, N4791);
and AND4 (N14357, N14344, N619, N7047, N12806);
buf BUF1 (N14358, N14339);
buf BUF1 (N14359, N14345);
not NOT1 (N14360, N14355);
and AND4 (N14361, N14356, N11264, N6617, N12434);
and AND2 (N14362, N14360, N13383);
or OR4 (N14363, N14353, N11479, N3324, N9069);
or OR3 (N14364, N14361, N4102, N7599);
xor XOR2 (N14365, N14347, N6725);
not NOT1 (N14366, N14346);
or OR4 (N14367, N14352, N2024, N3143, N6479);
nor NOR3 (N14368, N14359, N6051, N243);
and AND3 (N14369, N14366, N12597, N3936);
not NOT1 (N14370, N14369);
or OR2 (N14371, N14354, N14198);
nor NOR3 (N14372, N14365, N8872, N6109);
or OR4 (N14373, N14372, N13962, N6765, N10945);
not NOT1 (N14374, N14368);
buf BUF1 (N14375, N14358);
and AND4 (N14376, N14373, N7676, N11063, N8784);
nor NOR4 (N14377, N14375, N12949, N11741, N7275);
xor XOR2 (N14378, N14363, N9295);
nor NOR2 (N14379, N14364, N7166);
or OR4 (N14380, N14374, N8236, N13109, N4759);
buf BUF1 (N14381, N14377);
or OR4 (N14382, N14381, N912, N9354, N14045);
not NOT1 (N14383, N14379);
and AND2 (N14384, N14362, N12677);
xor XOR2 (N14385, N14383, N6280);
xor XOR2 (N14386, N14370, N6971);
or OR2 (N14387, N14357, N3204);
nand NAND3 (N14388, N14376, N4167, N4466);
and AND3 (N14389, N14378, N3989, N245);
not NOT1 (N14390, N14385);
or OR3 (N14391, N14389, N2954, N12265);
nand NAND2 (N14392, N14382, N13032);
and AND3 (N14393, N14371, N10340, N7066);
or OR3 (N14394, N14387, N4725, N3452);
nor NOR2 (N14395, N14367, N13778);
and AND4 (N14396, N14380, N3274, N4213, N5749);
nor NOR4 (N14397, N14393, N1833, N4887, N8997);
not NOT1 (N14398, N14391);
nand NAND4 (N14399, N14395, N3542, N6972, N3045);
buf BUF1 (N14400, N14398);
buf BUF1 (N14401, N14390);
buf BUF1 (N14402, N14401);
buf BUF1 (N14403, N14399);
xor XOR2 (N14404, N14392, N8134);
or OR4 (N14405, N14384, N11867, N11219, N996);
nand NAND2 (N14406, N14394, N13602);
and AND2 (N14407, N14388, N4060);
nand NAND4 (N14408, N14402, N3971, N12824, N7798);
or OR4 (N14409, N14403, N10254, N10377, N3737);
xor XOR2 (N14410, N14405, N11761);
or OR3 (N14411, N14396, N9282, N4872);
not NOT1 (N14412, N14386);
or OR4 (N14413, N14411, N5086, N254, N6943);
xor XOR2 (N14414, N14413, N3420);
and AND2 (N14415, N14397, N858);
or OR3 (N14416, N14414, N2986, N1502);
buf BUF1 (N14417, N14406);
buf BUF1 (N14418, N14412);
nor NOR4 (N14419, N14416, N4621, N979, N9412);
or OR4 (N14420, N14407, N1194, N8351, N2930);
nor NOR4 (N14421, N14410, N8027, N14406, N13124);
and AND2 (N14422, N14418, N5451);
buf BUF1 (N14423, N14420);
or OR2 (N14424, N14409, N3125);
and AND4 (N14425, N14400, N9017, N9178, N12244);
or OR2 (N14426, N14419, N8748);
buf BUF1 (N14427, N14417);
buf BUF1 (N14428, N14408);
or OR2 (N14429, N14427, N8639);
xor XOR2 (N14430, N14415, N12434);
xor XOR2 (N14431, N14426, N7938);
buf BUF1 (N14432, N14431);
not NOT1 (N14433, N14423);
xor XOR2 (N14434, N14432, N5286);
xor XOR2 (N14435, N14434, N2604);
buf BUF1 (N14436, N14435);
and AND2 (N14437, N14430, N4724);
xor XOR2 (N14438, N14421, N3436);
and AND3 (N14439, N14429, N11595, N7607);
nor NOR3 (N14440, N14439, N7522, N2297);
or OR3 (N14441, N14425, N5439, N10298);
nand NAND2 (N14442, N14438, N14105);
and AND2 (N14443, N14433, N6875);
nand NAND4 (N14444, N14440, N13362, N9032, N4108);
or OR3 (N14445, N14422, N812, N5937);
or OR3 (N14446, N14437, N10348, N145);
buf BUF1 (N14447, N14441);
and AND2 (N14448, N14442, N7275);
buf BUF1 (N14449, N14444);
nand NAND2 (N14450, N14443, N11775);
not NOT1 (N14451, N14404);
or OR3 (N14452, N14446, N11456, N10456);
nor NOR3 (N14453, N14447, N7294, N7898);
or OR4 (N14454, N14451, N10597, N13329, N2150);
buf BUF1 (N14455, N14453);
and AND3 (N14456, N14454, N299, N10684);
nor NOR4 (N14457, N14448, N175, N3311, N14045);
xor XOR2 (N14458, N14456, N11051);
or OR3 (N14459, N14458, N7970, N5468);
and AND3 (N14460, N14452, N12991, N10747);
not NOT1 (N14461, N14445);
or OR4 (N14462, N14428, N5277, N12462, N8231);
xor XOR2 (N14463, N14450, N14139);
or OR2 (N14464, N14455, N10968);
nand NAND4 (N14465, N14461, N7384, N13485, N13019);
and AND3 (N14466, N14424, N4559, N13833);
xor XOR2 (N14467, N14465, N2618);
xor XOR2 (N14468, N14467, N12421);
or OR3 (N14469, N14464, N4125, N5801);
xor XOR2 (N14470, N14460, N9691);
nor NOR4 (N14471, N14470, N3531, N10796, N11549);
and AND4 (N14472, N14468, N2736, N2881, N8857);
and AND2 (N14473, N14459, N13940);
nor NOR3 (N14474, N14471, N6038, N12752);
and AND2 (N14475, N14472, N7679);
nand NAND2 (N14476, N14463, N13799);
xor XOR2 (N14477, N14457, N10346);
nand NAND2 (N14478, N14462, N553);
buf BUF1 (N14479, N14473);
nand NAND3 (N14480, N14466, N5054, N12629);
buf BUF1 (N14481, N14449);
and AND2 (N14482, N14477, N5526);
xor XOR2 (N14483, N14475, N8467);
nor NOR4 (N14484, N14480, N12880, N5592, N2151);
buf BUF1 (N14485, N14478);
nor NOR2 (N14486, N14436, N12835);
and AND2 (N14487, N14486, N13808);
nand NAND4 (N14488, N14474, N11328, N1005, N425);
nand NAND3 (N14489, N14469, N10535, N2310);
buf BUF1 (N14490, N14483);
and AND4 (N14491, N14479, N11505, N11515, N3355);
nor NOR4 (N14492, N14487, N8516, N10190, N8485);
xor XOR2 (N14493, N14485, N11042);
xor XOR2 (N14494, N14476, N5009);
not NOT1 (N14495, N14482);
and AND4 (N14496, N14490, N10317, N4714, N1848);
or OR4 (N14497, N14488, N9833, N14205, N5776);
not NOT1 (N14498, N14489);
not NOT1 (N14499, N14492);
and AND2 (N14500, N14498, N13320);
buf BUF1 (N14501, N14481);
nor NOR3 (N14502, N14491, N3835, N11446);
not NOT1 (N14503, N14496);
nand NAND4 (N14504, N14501, N3616, N6880, N696);
and AND2 (N14505, N14500, N6536);
nor NOR4 (N14506, N14493, N7297, N10181, N11368);
and AND4 (N14507, N14505, N2084, N6737, N10294);
nor NOR3 (N14508, N14494, N1659, N4155);
not NOT1 (N14509, N14495);
not NOT1 (N14510, N14507);
and AND4 (N14511, N14504, N8948, N8663, N3702);
buf BUF1 (N14512, N14510);
not NOT1 (N14513, N14503);
buf BUF1 (N14514, N14511);
nor NOR3 (N14515, N14502, N50, N13971);
xor XOR2 (N14516, N14514, N6174);
buf BUF1 (N14517, N14497);
buf BUF1 (N14518, N14515);
nand NAND3 (N14519, N14518, N8316, N778);
xor XOR2 (N14520, N14512, N8881);
buf BUF1 (N14521, N14509);
nand NAND2 (N14522, N14516, N173);
or OR2 (N14523, N14519, N14421);
buf BUF1 (N14524, N14508);
nand NAND2 (N14525, N14513, N8052);
and AND3 (N14526, N14522, N3155, N41);
buf BUF1 (N14527, N14506);
and AND3 (N14528, N14527, N6996, N7558);
and AND2 (N14529, N14523, N6824);
xor XOR2 (N14530, N14525, N1373);
nand NAND2 (N14531, N14526, N13220);
nand NAND4 (N14532, N14524, N6050, N11349, N1084);
not NOT1 (N14533, N14528);
or OR4 (N14534, N14499, N11429, N710, N11835);
nor NOR2 (N14535, N14531, N3752);
nor NOR2 (N14536, N14529, N5333);
not NOT1 (N14537, N14484);
or OR4 (N14538, N14536, N2674, N11422, N6094);
buf BUF1 (N14539, N14537);
or OR2 (N14540, N14530, N11725);
nand NAND4 (N14541, N14540, N3033, N10845, N7902);
not NOT1 (N14542, N14533);
nor NOR3 (N14543, N14541, N2878, N8543);
or OR2 (N14544, N14534, N10308);
or OR4 (N14545, N14544, N12050, N6760, N12928);
xor XOR2 (N14546, N14532, N10739);
nand NAND2 (N14547, N14538, N11504);
buf BUF1 (N14548, N14517);
not NOT1 (N14549, N14542);
and AND2 (N14550, N14547, N13456);
or OR4 (N14551, N14543, N5838, N4463, N2459);
or OR2 (N14552, N14548, N13859);
xor XOR2 (N14553, N14546, N6978);
nor NOR2 (N14554, N14550, N7566);
buf BUF1 (N14555, N14553);
not NOT1 (N14556, N14549);
xor XOR2 (N14557, N14521, N3125);
xor XOR2 (N14558, N14552, N13906);
and AND2 (N14559, N14555, N814);
nor NOR3 (N14560, N14539, N6499, N4404);
buf BUF1 (N14561, N14545);
buf BUF1 (N14562, N14557);
nand NAND3 (N14563, N14551, N6339, N8095);
xor XOR2 (N14564, N14563, N8747);
nand NAND4 (N14565, N14562, N10943, N172, N5519);
buf BUF1 (N14566, N14565);
xor XOR2 (N14567, N14561, N7913);
or OR2 (N14568, N14554, N1854);
nand NAND4 (N14569, N14520, N11047, N11377, N13874);
nor NOR4 (N14570, N14568, N6287, N14152, N9120);
and AND3 (N14571, N14569, N11655, N6037);
not NOT1 (N14572, N14558);
and AND2 (N14573, N14572, N12156);
nand NAND3 (N14574, N14571, N4795, N8542);
not NOT1 (N14575, N14559);
or OR3 (N14576, N14556, N10809, N10795);
nor NOR3 (N14577, N14570, N1267, N4430);
nor NOR4 (N14578, N14575, N9872, N12294, N10819);
xor XOR2 (N14579, N14574, N2678);
xor XOR2 (N14580, N14577, N4744);
nand NAND2 (N14581, N14578, N11688);
or OR2 (N14582, N14566, N5305);
buf BUF1 (N14583, N14576);
nand NAND2 (N14584, N14535, N1626);
not NOT1 (N14585, N14580);
nor NOR2 (N14586, N14567, N2241);
not NOT1 (N14587, N14573);
and AND2 (N14588, N14581, N810);
nand NAND2 (N14589, N14587, N9720);
nor NOR2 (N14590, N14560, N10921);
nand NAND3 (N14591, N14582, N5771, N4527);
not NOT1 (N14592, N14579);
nand NAND2 (N14593, N14591, N4024);
buf BUF1 (N14594, N14584);
not NOT1 (N14595, N14590);
buf BUF1 (N14596, N14564);
or OR3 (N14597, N14586, N2219, N8112);
and AND3 (N14598, N14595, N5491, N7887);
nand NAND3 (N14599, N14598, N1128, N9078);
not NOT1 (N14600, N14599);
nand NAND4 (N14601, N14596, N852, N12403, N4796);
or OR2 (N14602, N14588, N13672);
nor NOR3 (N14603, N14602, N7297, N6478);
or OR3 (N14604, N14601, N8798, N8423);
and AND4 (N14605, N14597, N9781, N10440, N4847);
not NOT1 (N14606, N14603);
xor XOR2 (N14607, N14589, N2058);
or OR2 (N14608, N14606, N4278);
not NOT1 (N14609, N14604);
not NOT1 (N14610, N14605);
xor XOR2 (N14611, N14592, N6590);
or OR4 (N14612, N14611, N13975, N12888, N6885);
or OR2 (N14613, N14594, N5905);
nand NAND3 (N14614, N14613, N7786, N10746);
not NOT1 (N14615, N14585);
buf BUF1 (N14616, N14610);
xor XOR2 (N14617, N14609, N13238);
xor XOR2 (N14618, N14600, N10888);
buf BUF1 (N14619, N14607);
nand NAND2 (N14620, N14583, N9423);
and AND3 (N14621, N14618, N14018, N7907);
xor XOR2 (N14622, N14621, N6422);
and AND2 (N14623, N14612, N14525);
and AND3 (N14624, N14614, N732, N3555);
and AND2 (N14625, N14616, N6069);
buf BUF1 (N14626, N14615);
or OR2 (N14627, N14622, N1395);
xor XOR2 (N14628, N14623, N3270);
buf BUF1 (N14629, N14619);
or OR3 (N14630, N14627, N736, N1751);
and AND2 (N14631, N14630, N11631);
not NOT1 (N14632, N14629);
xor XOR2 (N14633, N14631, N5433);
xor XOR2 (N14634, N14628, N5386);
or OR3 (N14635, N14625, N4073, N2531);
and AND2 (N14636, N14632, N7206);
and AND4 (N14637, N14608, N1856, N7578, N8344);
and AND4 (N14638, N14617, N1711, N11952, N11309);
nor NOR3 (N14639, N14593, N2320, N8457);
nor NOR3 (N14640, N14636, N13627, N6585);
or OR2 (N14641, N14633, N2997);
buf BUF1 (N14642, N14624);
nand NAND2 (N14643, N14637, N3184);
xor XOR2 (N14644, N14620, N14186);
nand NAND2 (N14645, N14643, N6327);
not NOT1 (N14646, N14638);
or OR4 (N14647, N14626, N11831, N502, N8258);
xor XOR2 (N14648, N14642, N5311);
buf BUF1 (N14649, N14645);
nand NAND4 (N14650, N14635, N4360, N9190, N13978);
and AND3 (N14651, N14644, N11713, N5630);
nand NAND2 (N14652, N14640, N2580);
and AND4 (N14653, N14634, N7616, N4074, N8858);
nand NAND3 (N14654, N14653, N11350, N13979);
buf BUF1 (N14655, N14649);
and AND2 (N14656, N14646, N5297);
and AND2 (N14657, N14654, N10927);
nor NOR2 (N14658, N14641, N1096);
not NOT1 (N14659, N14656);
not NOT1 (N14660, N14647);
nand NAND3 (N14661, N14659, N1218, N914);
xor XOR2 (N14662, N14655, N6936);
nor NOR4 (N14663, N14661, N1583, N5567, N5353);
nand NAND4 (N14664, N14658, N2143, N356, N9828);
nor NOR4 (N14665, N14639, N1142, N11694, N5066);
nand NAND4 (N14666, N14664, N14013, N9085, N13681);
and AND3 (N14667, N14663, N5796, N1700);
and AND3 (N14668, N14660, N3686, N1652);
nor NOR4 (N14669, N14667, N1404, N11640, N13620);
and AND4 (N14670, N14648, N13114, N5443, N3880);
and AND2 (N14671, N14662, N7136);
not NOT1 (N14672, N14666);
nand NAND3 (N14673, N14670, N5609, N6451);
buf BUF1 (N14674, N14672);
and AND4 (N14675, N14668, N10065, N13705, N722);
nand NAND3 (N14676, N14671, N8900, N7748);
nand NAND4 (N14677, N14675, N4444, N4538, N239);
buf BUF1 (N14678, N14665);
and AND2 (N14679, N14677, N7989);
not NOT1 (N14680, N14679);
nor NOR4 (N14681, N14651, N882, N1128, N13981);
not NOT1 (N14682, N14674);
nor NOR4 (N14683, N14650, N6213, N11150, N1532);
or OR3 (N14684, N14680, N7396, N8912);
nor NOR4 (N14685, N14678, N4400, N4027, N9930);
not NOT1 (N14686, N14682);
nand NAND3 (N14687, N14657, N9295, N10463);
or OR2 (N14688, N14687, N6433);
nor NOR3 (N14689, N14669, N6445, N7554);
xor XOR2 (N14690, N14685, N14460);
xor XOR2 (N14691, N14652, N13333);
and AND2 (N14692, N14673, N11860);
not NOT1 (N14693, N14676);
nor NOR2 (N14694, N14692, N2903);
and AND4 (N14695, N14684, N6939, N12147, N13438);
not NOT1 (N14696, N14693);
nand NAND3 (N14697, N14691, N6018, N5144);
not NOT1 (N14698, N14688);
or OR2 (N14699, N14696, N2287);
not NOT1 (N14700, N14694);
xor XOR2 (N14701, N14698, N8586);
not NOT1 (N14702, N14700);
nor NOR3 (N14703, N14686, N9942, N5184);
buf BUF1 (N14704, N14689);
not NOT1 (N14705, N14695);
or OR4 (N14706, N14683, N6947, N13021, N6952);
nand NAND4 (N14707, N14699, N2241, N12829, N9351);
or OR2 (N14708, N14703, N2228);
xor XOR2 (N14709, N14706, N2608);
xor XOR2 (N14710, N14702, N421);
and AND3 (N14711, N14704, N13547, N3061);
not NOT1 (N14712, N14681);
nor NOR4 (N14713, N14711, N9567, N6253, N7111);
nor NOR2 (N14714, N14701, N14154);
or OR3 (N14715, N14714, N3834, N10456);
or OR4 (N14716, N14713, N8164, N8972, N5057);
nor NOR3 (N14717, N14697, N9357, N1120);
or OR3 (N14718, N14705, N13091, N11895);
not NOT1 (N14719, N14715);
nand NAND2 (N14720, N14690, N8085);
and AND3 (N14721, N14720, N10795, N5355);
not NOT1 (N14722, N14716);
nor NOR4 (N14723, N14709, N10684, N7114, N1028);
or OR3 (N14724, N14721, N1538, N7082);
nand NAND4 (N14725, N14724, N22, N13299, N7046);
xor XOR2 (N14726, N14717, N13517);
nor NOR2 (N14727, N14707, N10142);
not NOT1 (N14728, N14722);
or OR2 (N14729, N14718, N13413);
or OR4 (N14730, N14727, N7962, N9992, N4072);
and AND4 (N14731, N14708, N6860, N2902, N7780);
nor NOR3 (N14732, N14723, N14257, N314);
xor XOR2 (N14733, N14731, N3115);
or OR2 (N14734, N14732, N4686);
not NOT1 (N14735, N14719);
nand NAND3 (N14736, N14735, N10392, N1869);
xor XOR2 (N14737, N14710, N7211);
and AND3 (N14738, N14730, N9025, N214);
not NOT1 (N14739, N14736);
not NOT1 (N14740, N14712);
nor NOR3 (N14741, N14733, N10585, N7086);
not NOT1 (N14742, N14725);
and AND3 (N14743, N14737, N2294, N1857);
xor XOR2 (N14744, N14726, N1241);
not NOT1 (N14745, N14741);
or OR2 (N14746, N14739, N14455);
or OR3 (N14747, N14734, N1757, N13151);
and AND3 (N14748, N14740, N12839, N9859);
nor NOR3 (N14749, N14747, N12849, N150);
not NOT1 (N14750, N14742);
xor XOR2 (N14751, N14728, N8606);
nand NAND2 (N14752, N14729, N4872);
not NOT1 (N14753, N14738);
nor NOR3 (N14754, N14751, N3906, N591);
buf BUF1 (N14755, N14745);
buf BUF1 (N14756, N14754);
nand NAND3 (N14757, N14743, N11527, N6076);
xor XOR2 (N14758, N14755, N3793);
and AND2 (N14759, N14744, N8834);
not NOT1 (N14760, N14756);
or OR4 (N14761, N14746, N13047, N1346, N6979);
nand NAND2 (N14762, N14757, N9362);
or OR4 (N14763, N14758, N13567, N5080, N9455);
nor NOR4 (N14764, N14750, N2372, N1944, N13);
xor XOR2 (N14765, N14759, N11700);
buf BUF1 (N14766, N14764);
nor NOR3 (N14767, N14748, N10599, N3926);
or OR2 (N14768, N14760, N2181);
and AND2 (N14769, N14752, N7064);
or OR4 (N14770, N14765, N2169, N14282, N8373);
nand NAND2 (N14771, N14749, N3296);
not NOT1 (N14772, N14770);
buf BUF1 (N14773, N14768);
xor XOR2 (N14774, N14766, N12439);
not NOT1 (N14775, N14769);
and AND3 (N14776, N14762, N11243, N1469);
or OR4 (N14777, N14772, N12876, N1593, N14322);
xor XOR2 (N14778, N14776, N12249);
nor NOR2 (N14779, N14771, N3376);
and AND3 (N14780, N14778, N11455, N8684);
nand NAND4 (N14781, N14780, N3383, N1958, N7934);
nand NAND2 (N14782, N14774, N13486);
nor NOR2 (N14783, N14779, N6403);
nand NAND2 (N14784, N14775, N7624);
buf BUF1 (N14785, N14783);
or OR3 (N14786, N14782, N4397, N1969);
buf BUF1 (N14787, N14761);
xor XOR2 (N14788, N14763, N4397);
buf BUF1 (N14789, N14785);
and AND2 (N14790, N14777, N8038);
nor NOR3 (N14791, N14784, N4392, N4977);
or OR3 (N14792, N14787, N601, N8531);
nand NAND3 (N14793, N14792, N14317, N14439);
nand NAND4 (N14794, N14790, N13694, N3909, N10058);
not NOT1 (N14795, N14791);
buf BUF1 (N14796, N14781);
or OR3 (N14797, N14753, N11888, N10251);
xor XOR2 (N14798, N14773, N14639);
xor XOR2 (N14799, N14795, N12569);
not NOT1 (N14800, N14796);
xor XOR2 (N14801, N14800, N9307);
nand NAND2 (N14802, N14794, N13530);
and AND4 (N14803, N14797, N14588, N11391, N4709);
buf BUF1 (N14804, N14788);
buf BUF1 (N14805, N14798);
not NOT1 (N14806, N14803);
nand NAND4 (N14807, N14801, N4579, N11371, N3540);
or OR3 (N14808, N14786, N8492, N11907);
nand NAND2 (N14809, N14806, N5276);
nand NAND2 (N14810, N14804, N1002);
or OR4 (N14811, N14807, N2953, N12997, N753);
nor NOR3 (N14812, N14808, N12357, N5053);
xor XOR2 (N14813, N14812, N3554);
and AND3 (N14814, N14799, N2754, N12948);
buf BUF1 (N14815, N14793);
xor XOR2 (N14816, N14767, N14265);
or OR3 (N14817, N14810, N8054, N4952);
buf BUF1 (N14818, N14809);
nor NOR3 (N14819, N14811, N9892, N1467);
and AND4 (N14820, N14815, N8497, N12939, N13893);
and AND4 (N14821, N14817, N14665, N10218, N8111);
buf BUF1 (N14822, N14821);
xor XOR2 (N14823, N14816, N1196);
not NOT1 (N14824, N14822);
or OR4 (N14825, N14820, N11959, N3531, N1696);
and AND4 (N14826, N14818, N10015, N13808, N7506);
nor NOR2 (N14827, N14824, N1018);
nand NAND4 (N14828, N14827, N6691, N4098, N5126);
and AND3 (N14829, N14802, N3793, N12044);
buf BUF1 (N14830, N14829);
nand NAND3 (N14831, N14828, N13160, N12477);
xor XOR2 (N14832, N14823, N4283);
nor NOR2 (N14833, N14813, N14629);
and AND3 (N14834, N14789, N5480, N14529);
and AND2 (N14835, N14814, N871);
nand NAND4 (N14836, N14835, N1980, N4795, N9728);
nand NAND4 (N14837, N14825, N1045, N7468, N6121);
nor NOR4 (N14838, N14836, N9710, N132, N2049);
or OR4 (N14839, N14833, N695, N8106, N470);
nand NAND3 (N14840, N14831, N2847, N865);
xor XOR2 (N14841, N14838, N547);
or OR2 (N14842, N14832, N12703);
or OR2 (N14843, N14830, N2302);
xor XOR2 (N14844, N14826, N9100);
or OR3 (N14845, N14842, N1562, N7859);
and AND4 (N14846, N14844, N14779, N259, N6335);
or OR4 (N14847, N14837, N6116, N8242, N396);
buf BUF1 (N14848, N14845);
not NOT1 (N14849, N14846);
or OR2 (N14850, N14834, N6370);
xor XOR2 (N14851, N14849, N13973);
xor XOR2 (N14852, N14819, N3648);
buf BUF1 (N14853, N14840);
nand NAND2 (N14854, N14847, N3230);
xor XOR2 (N14855, N14853, N7992);
buf BUF1 (N14856, N14854);
or OR4 (N14857, N14850, N14693, N11944, N14089);
nand NAND2 (N14858, N14856, N5855);
or OR2 (N14859, N14843, N6316);
xor XOR2 (N14860, N14848, N12242);
not NOT1 (N14861, N14852);
nor NOR3 (N14862, N14841, N4556, N9740);
or OR2 (N14863, N14859, N8615);
buf BUF1 (N14864, N14862);
buf BUF1 (N14865, N14864);
xor XOR2 (N14866, N14865, N10982);
and AND3 (N14867, N14858, N5646, N6424);
not NOT1 (N14868, N14851);
and AND4 (N14869, N14857, N2342, N11934, N9304);
and AND4 (N14870, N14861, N8145, N9175, N14676);
xor XOR2 (N14871, N14866, N7227);
or OR4 (N14872, N14860, N7393, N10717, N7773);
buf BUF1 (N14873, N14872);
and AND3 (N14874, N14868, N14850, N6986);
xor XOR2 (N14875, N14867, N953);
not NOT1 (N14876, N14870);
buf BUF1 (N14877, N14876);
and AND2 (N14878, N14855, N1268);
nor NOR3 (N14879, N14873, N8166, N585);
xor XOR2 (N14880, N14875, N1);
buf BUF1 (N14881, N14863);
xor XOR2 (N14882, N14869, N1374);
nor NOR4 (N14883, N14877, N4723, N11919, N490);
not NOT1 (N14884, N14839);
and AND4 (N14885, N14880, N2325, N10056, N12513);
and AND4 (N14886, N14884, N5244, N12508, N9308);
nor NOR4 (N14887, N14881, N9711, N6479, N2048);
and AND3 (N14888, N14885, N6631, N179);
or OR4 (N14889, N14805, N5053, N1723, N13723);
or OR2 (N14890, N14886, N9930);
xor XOR2 (N14891, N14883, N8631);
buf BUF1 (N14892, N14874);
not NOT1 (N14893, N14892);
nand NAND3 (N14894, N14888, N6869, N4917);
nand NAND3 (N14895, N14871, N848, N11556);
not NOT1 (N14896, N14879);
not NOT1 (N14897, N14890);
buf BUF1 (N14898, N14895);
and AND4 (N14899, N14897, N1880, N14738, N8738);
xor XOR2 (N14900, N14898, N12661);
or OR4 (N14901, N14882, N5066, N4243, N14755);
xor XOR2 (N14902, N14901, N6222);
or OR2 (N14903, N14893, N1612);
nor NOR3 (N14904, N14903, N3179, N4274);
and AND4 (N14905, N14887, N3976, N10452, N12094);
xor XOR2 (N14906, N14902, N1263);
not NOT1 (N14907, N14900);
nor NOR2 (N14908, N14899, N11458);
nand NAND3 (N14909, N14904, N2466, N13818);
or OR2 (N14910, N14907, N10432);
and AND3 (N14911, N14906, N11435, N10565);
not NOT1 (N14912, N14911);
nor NOR2 (N14913, N14908, N523);
not NOT1 (N14914, N14905);
or OR2 (N14915, N14889, N4549);
nand NAND4 (N14916, N14913, N10728, N982, N14680);
nand NAND3 (N14917, N14910, N4212, N8629);
xor XOR2 (N14918, N14914, N7783);
and AND4 (N14919, N14878, N11282, N12251, N13293);
xor XOR2 (N14920, N14917, N4921);
nand NAND2 (N14921, N14912, N9887);
and AND4 (N14922, N14919, N2098, N9793, N9298);
xor XOR2 (N14923, N14891, N11916);
xor XOR2 (N14924, N14921, N14681);
xor XOR2 (N14925, N14923, N1790);
buf BUF1 (N14926, N14894);
nor NOR4 (N14927, N14909, N11759, N7425, N3823);
and AND3 (N14928, N14926, N59, N4160);
not NOT1 (N14929, N14928);
buf BUF1 (N14930, N14927);
nor NOR2 (N14931, N14929, N5110);
not NOT1 (N14932, N14918);
or OR3 (N14933, N14896, N6891, N12681);
and AND4 (N14934, N14924, N4431, N9484, N6947);
nor NOR3 (N14935, N14931, N6895, N8635);
nor NOR2 (N14936, N14935, N3541);
and AND2 (N14937, N14922, N13555);
nand NAND3 (N14938, N14934, N7893, N4157);
xor XOR2 (N14939, N14930, N9146);
and AND2 (N14940, N14916, N11446);
or OR3 (N14941, N14939, N8954, N3766);
buf BUF1 (N14942, N14936);
and AND4 (N14943, N14920, N8336, N12804, N2376);
nand NAND3 (N14944, N14932, N8031, N10660);
xor XOR2 (N14945, N14938, N579);
or OR2 (N14946, N14915, N7314);
nor NOR2 (N14947, N14944, N2833);
nand NAND2 (N14948, N14946, N5696);
nand NAND3 (N14949, N14943, N494, N713);
nand NAND4 (N14950, N14933, N4018, N4446, N7037);
xor XOR2 (N14951, N14925, N13541);
nor NOR4 (N14952, N14947, N11259, N8029, N12399);
nand NAND2 (N14953, N14940, N7769);
or OR3 (N14954, N14952, N11429, N5195);
or OR4 (N14955, N14954, N8491, N1161, N14044);
xor XOR2 (N14956, N14937, N4762);
not NOT1 (N14957, N14951);
nand NAND4 (N14958, N14941, N1233, N9161, N13431);
not NOT1 (N14959, N14953);
buf BUF1 (N14960, N14949);
and AND2 (N14961, N14942, N8867);
nand NAND4 (N14962, N14945, N464, N6127, N3777);
nand NAND4 (N14963, N14948, N4337, N14547, N1580);
buf BUF1 (N14964, N14955);
buf BUF1 (N14965, N14958);
or OR4 (N14966, N14963, N2367, N8154, N5312);
and AND3 (N14967, N14960, N1499, N2827);
nand NAND3 (N14968, N14962, N12109, N3924);
buf BUF1 (N14969, N14965);
or OR2 (N14970, N14950, N4951);
not NOT1 (N14971, N14966);
nand NAND2 (N14972, N14968, N3329);
nor NOR3 (N14973, N14961, N8265, N6992);
not NOT1 (N14974, N14971);
or OR3 (N14975, N14969, N2724, N10066);
nand NAND2 (N14976, N14973, N14504);
buf BUF1 (N14977, N14959);
buf BUF1 (N14978, N14977);
or OR2 (N14979, N14978, N4166);
xor XOR2 (N14980, N14974, N12202);
not NOT1 (N14981, N14979);
buf BUF1 (N14982, N14964);
xor XOR2 (N14983, N14956, N12838);
xor XOR2 (N14984, N14970, N8180);
and AND2 (N14985, N14980, N9864);
not NOT1 (N14986, N14957);
or OR3 (N14987, N14976, N3983, N7179);
or OR2 (N14988, N14983, N10081);
xor XOR2 (N14989, N14987, N8575);
nor NOR3 (N14990, N14985, N9748, N13977);
not NOT1 (N14991, N14981);
buf BUF1 (N14992, N14989);
not NOT1 (N14993, N14990);
xor XOR2 (N14994, N14993, N10630);
buf BUF1 (N14995, N14982);
or OR4 (N14996, N14995, N5555, N8643, N11564);
nor NOR4 (N14997, N14988, N6616, N4709, N9543);
nand NAND4 (N14998, N14967, N1038, N3536, N774);
buf BUF1 (N14999, N14998);
buf BUF1 (N15000, N14994);
nor NOR4 (N15001, N14992, N12370, N7008, N9240);
or OR3 (N15002, N14999, N10728, N2623);
or OR3 (N15003, N14972, N1063, N6687);
nor NOR4 (N15004, N14996, N14804, N6082, N2621);
xor XOR2 (N15005, N15003, N7753);
not NOT1 (N15006, N14975);
not NOT1 (N15007, N14991);
or OR3 (N15008, N14984, N12917, N10392);
nand NAND2 (N15009, N14986, N5591);
or OR4 (N15010, N15007, N8346, N3428, N8683);
buf BUF1 (N15011, N15004);
xor XOR2 (N15012, N15001, N8188);
buf BUF1 (N15013, N15006);
xor XOR2 (N15014, N15008, N22);
nor NOR2 (N15015, N15014, N12456);
nor NOR2 (N15016, N15009, N8273);
nor NOR3 (N15017, N15015, N4816, N2053);
nand NAND4 (N15018, N15012, N6674, N8605, N14430);
nor NOR4 (N15019, N15013, N7101, N10591, N3585);
nor NOR3 (N15020, N15002, N4456, N7711);
or OR4 (N15021, N15018, N129, N4588, N14056);
nand NAND3 (N15022, N15011, N6319, N5296);
xor XOR2 (N15023, N14997, N43);
xor XOR2 (N15024, N15000, N9826);
buf BUF1 (N15025, N15010);
nor NOR3 (N15026, N15016, N1645, N8608);
and AND4 (N15027, N15005, N14311, N548, N11373);
and AND3 (N15028, N15026, N1124, N14073);
xor XOR2 (N15029, N15019, N13559);
nor NOR2 (N15030, N15021, N10363);
and AND3 (N15031, N15025, N2966, N6902);
or OR3 (N15032, N15028, N1961, N12401);
not NOT1 (N15033, N15022);
and AND4 (N15034, N15020, N9950, N6156, N1546);
and AND4 (N15035, N15032, N5410, N14277, N313);
and AND3 (N15036, N15033, N15029, N10775);
nand NAND4 (N15037, N13310, N4519, N3939, N12152);
buf BUF1 (N15038, N15031);
buf BUF1 (N15039, N15037);
nand NAND2 (N15040, N15027, N3391);
not NOT1 (N15041, N15017);
nor NOR2 (N15042, N15036, N5961);
not NOT1 (N15043, N15041);
or OR3 (N15044, N15023, N7663, N402);
or OR3 (N15045, N15038, N8966, N13478);
buf BUF1 (N15046, N15045);
and AND2 (N15047, N15046, N6252);
and AND2 (N15048, N15035, N7202);
or OR3 (N15049, N15048, N10827, N9504);
nor NOR4 (N15050, N15047, N7960, N10551, N7124);
nand NAND2 (N15051, N15034, N10739);
and AND3 (N15052, N15049, N898, N11943);
or OR2 (N15053, N15050, N11076);
and AND2 (N15054, N15024, N10903);
or OR2 (N15055, N15051, N1670);
not NOT1 (N15056, N15044);
and AND2 (N15057, N15040, N6028);
xor XOR2 (N15058, N15043, N1655);
buf BUF1 (N15059, N15056);
xor XOR2 (N15060, N15042, N12867);
nor NOR2 (N15061, N15057, N8669);
or OR2 (N15062, N15061, N3386);
buf BUF1 (N15063, N15062);
or OR2 (N15064, N15063, N5692);
or OR2 (N15065, N15060, N5773);
xor XOR2 (N15066, N15030, N6911);
nand NAND2 (N15067, N15054, N373);
not NOT1 (N15068, N15059);
and AND4 (N15069, N15064, N8126, N8612, N3688);
or OR2 (N15070, N15052, N827);
nand NAND3 (N15071, N15066, N5379, N3628);
not NOT1 (N15072, N15065);
and AND3 (N15073, N15069, N3219, N11062);
and AND3 (N15074, N15039, N11626, N5131);
buf BUF1 (N15075, N15073);
xor XOR2 (N15076, N15070, N5294);
xor XOR2 (N15077, N15072, N394);
nand NAND3 (N15078, N15075, N3653, N10421);
nor NOR2 (N15079, N15055, N4663);
or OR4 (N15080, N15079, N9601, N966, N3258);
nor NOR2 (N15081, N15076, N806);
nand NAND3 (N15082, N15081, N10177, N9905);
buf BUF1 (N15083, N15077);
xor XOR2 (N15084, N15078, N7772);
nand NAND3 (N15085, N15067, N962, N12027);
not NOT1 (N15086, N15085);
and AND3 (N15087, N15086, N4976, N1270);
nand NAND3 (N15088, N15083, N14207, N3018);
not NOT1 (N15089, N15058);
nor NOR4 (N15090, N15082, N13960, N2166, N2735);
xor XOR2 (N15091, N15053, N7268);
or OR2 (N15092, N15091, N9528);
nor NOR2 (N15093, N15092, N6398);
not NOT1 (N15094, N15087);
not NOT1 (N15095, N15090);
xor XOR2 (N15096, N15095, N3668);
not NOT1 (N15097, N15071);
nor NOR2 (N15098, N15097, N911);
and AND3 (N15099, N15074, N14, N5444);
buf BUF1 (N15100, N15099);
xor XOR2 (N15101, N15094, N10969);
and AND2 (N15102, N15096, N7165);
buf BUF1 (N15103, N15093);
nand NAND2 (N15104, N15102, N6401);
buf BUF1 (N15105, N15103);
and AND3 (N15106, N15104, N3942, N1320);
not NOT1 (N15107, N15088);
nand NAND4 (N15108, N15107, N12312, N14408, N9131);
xor XOR2 (N15109, N15084, N7575);
xor XOR2 (N15110, N15068, N14343);
and AND3 (N15111, N15105, N4779, N2398);
and AND3 (N15112, N15111, N2882, N6124);
buf BUF1 (N15113, N15108);
xor XOR2 (N15114, N15106, N5091);
not NOT1 (N15115, N15109);
not NOT1 (N15116, N15115);
buf BUF1 (N15117, N15101);
nor NOR2 (N15118, N15117, N7251);
nand NAND2 (N15119, N15098, N7384);
xor XOR2 (N15120, N15110, N11420);
nand NAND4 (N15121, N15114, N6491, N13050, N5205);
not NOT1 (N15122, N15113);
nor NOR2 (N15123, N15119, N11649);
buf BUF1 (N15124, N15120);
nand NAND4 (N15125, N15100, N4226, N3617, N14727);
buf BUF1 (N15126, N15080);
not NOT1 (N15127, N15089);
buf BUF1 (N15128, N15127);
or OR2 (N15129, N15118, N5421);
xor XOR2 (N15130, N15125, N6702);
or OR3 (N15131, N15123, N12098, N5937);
not NOT1 (N15132, N15131);
buf BUF1 (N15133, N15126);
nor NOR2 (N15134, N15130, N2844);
xor XOR2 (N15135, N15128, N13303);
nor NOR2 (N15136, N15133, N6224);
nor NOR2 (N15137, N15135, N6117);
not NOT1 (N15138, N15137);
not NOT1 (N15139, N15136);
xor XOR2 (N15140, N15129, N5587);
or OR2 (N15141, N15121, N3152);
nand NAND3 (N15142, N15116, N14870, N7610);
not NOT1 (N15143, N15132);
or OR3 (N15144, N15141, N7798, N6929);
or OR4 (N15145, N15124, N6538, N13640, N8715);
xor XOR2 (N15146, N15140, N12483);
nand NAND3 (N15147, N15138, N719, N6226);
not NOT1 (N15148, N15139);
nor NOR3 (N15149, N15144, N12859, N11742);
nand NAND4 (N15150, N15149, N15108, N944, N2507);
or OR2 (N15151, N15148, N9898);
or OR4 (N15152, N15150, N1746, N8725, N4953);
nor NOR2 (N15153, N15143, N7717);
or OR3 (N15154, N15145, N12681, N5363);
buf BUF1 (N15155, N15153);
and AND2 (N15156, N15122, N3293);
and AND4 (N15157, N15154, N5369, N383, N6796);
xor XOR2 (N15158, N15142, N12182);
and AND4 (N15159, N15152, N3006, N2162, N5978);
xor XOR2 (N15160, N15158, N8603);
and AND3 (N15161, N15155, N8682, N3075);
buf BUF1 (N15162, N15157);
and AND2 (N15163, N15159, N14175);
buf BUF1 (N15164, N15147);
or OR2 (N15165, N15156, N8317);
not NOT1 (N15166, N15146);
not NOT1 (N15167, N15164);
xor XOR2 (N15168, N15161, N8746);
and AND2 (N15169, N15168, N5644);
buf BUF1 (N15170, N15166);
xor XOR2 (N15171, N15160, N13075);
or OR3 (N15172, N15112, N8873, N14961);
buf BUF1 (N15173, N15162);
and AND4 (N15174, N15167, N9356, N13598, N11182);
not NOT1 (N15175, N15151);
or OR4 (N15176, N15170, N1802, N10228, N9954);
xor XOR2 (N15177, N15169, N2597);
and AND4 (N15178, N15163, N9577, N3446, N8787);
xor XOR2 (N15179, N15178, N3194);
nor NOR3 (N15180, N15174, N8881, N14759);
not NOT1 (N15181, N15173);
buf BUF1 (N15182, N15180);
or OR2 (N15183, N15177, N5397);
nor NOR3 (N15184, N15134, N7553, N8338);
nor NOR2 (N15185, N15172, N10708);
or OR3 (N15186, N15171, N9002, N13112);
xor XOR2 (N15187, N15185, N7474);
and AND4 (N15188, N15175, N2612, N12374, N11863);
buf BUF1 (N15189, N15181);
not NOT1 (N15190, N15182);
buf BUF1 (N15191, N15184);
xor XOR2 (N15192, N15183, N13482);
nand NAND4 (N15193, N15186, N7357, N12293, N2035);
buf BUF1 (N15194, N15187);
and AND2 (N15195, N15192, N14691);
xor XOR2 (N15196, N15165, N13939);
buf BUF1 (N15197, N15189);
or OR2 (N15198, N15193, N13754);
not NOT1 (N15199, N15191);
buf BUF1 (N15200, N15196);
and AND3 (N15201, N15197, N2813, N5009);
and AND3 (N15202, N15176, N7257, N14464);
nor NOR4 (N15203, N15201, N11952, N7345, N6933);
or OR2 (N15204, N15202, N2677);
and AND2 (N15205, N15195, N2663);
nand NAND4 (N15206, N15194, N2897, N10340, N15179);
xor XOR2 (N15207, N11260, N13551);
or OR3 (N15208, N15205, N2722, N7124);
nand NAND4 (N15209, N15200, N104, N8028, N13612);
not NOT1 (N15210, N15198);
nor NOR4 (N15211, N15209, N5112, N14244, N2256);
or OR4 (N15212, N15211, N10710, N12921, N12518);
nor NOR4 (N15213, N15212, N12742, N5361, N10847);
nand NAND2 (N15214, N15206, N2437);
xor XOR2 (N15215, N15208, N9965);
not NOT1 (N15216, N15190);
xor XOR2 (N15217, N15215, N3077);
xor XOR2 (N15218, N15213, N12028);
xor XOR2 (N15219, N15216, N7603);
or OR4 (N15220, N15217, N9176, N11878, N5064);
nand NAND4 (N15221, N15203, N9882, N6428, N14453);
buf BUF1 (N15222, N15220);
nor NOR3 (N15223, N15188, N6237, N5855);
buf BUF1 (N15224, N15204);
or OR4 (N15225, N15221, N3589, N4797, N9289);
nand NAND3 (N15226, N15199, N6059, N13133);
xor XOR2 (N15227, N15207, N3755);
xor XOR2 (N15228, N15223, N2972);
and AND3 (N15229, N15210, N7774, N14960);
nor NOR3 (N15230, N15218, N9904, N7375);
xor XOR2 (N15231, N15225, N12278);
and AND4 (N15232, N15226, N4425, N2336, N11755);
nor NOR4 (N15233, N15229, N12256, N14590, N10420);
buf BUF1 (N15234, N15233);
xor XOR2 (N15235, N15230, N4961);
nor NOR2 (N15236, N15227, N3805);
and AND3 (N15237, N15234, N14429, N14392);
nor NOR2 (N15238, N15237, N5884);
buf BUF1 (N15239, N15228);
nor NOR2 (N15240, N15239, N9786);
and AND3 (N15241, N15214, N1259, N7440);
xor XOR2 (N15242, N15219, N13763);
nor NOR4 (N15243, N15238, N5807, N3463, N11321);
or OR2 (N15244, N15236, N1490);
not NOT1 (N15245, N15222);
xor XOR2 (N15246, N15241, N2363);
and AND2 (N15247, N15244, N1095);
or OR2 (N15248, N15245, N8525);
xor XOR2 (N15249, N15246, N69);
not NOT1 (N15250, N15231);
or OR4 (N15251, N15247, N928, N4951, N11292);
or OR3 (N15252, N15248, N1390, N11992);
not NOT1 (N15253, N15240);
and AND4 (N15254, N15253, N13129, N10951, N11108);
buf BUF1 (N15255, N15242);
or OR3 (N15256, N15250, N10597, N8767);
nor NOR4 (N15257, N15224, N15215, N2138, N1560);
and AND3 (N15258, N15251, N974, N10215);
buf BUF1 (N15259, N15255);
or OR3 (N15260, N15256, N233, N4151);
and AND4 (N15261, N15249, N10228, N11359, N2848);
nor NOR3 (N15262, N15260, N13938, N4626);
not NOT1 (N15263, N15232);
not NOT1 (N15264, N15243);
or OR4 (N15265, N15264, N5442, N5092, N190);
not NOT1 (N15266, N15252);
buf BUF1 (N15267, N15259);
not NOT1 (N15268, N15262);
or OR4 (N15269, N15235, N11307, N13318, N15080);
nand NAND3 (N15270, N15269, N5319, N11476);
buf BUF1 (N15271, N15254);
nand NAND2 (N15272, N15266, N10621);
and AND3 (N15273, N15257, N7624, N2200);
nor NOR4 (N15274, N15261, N13302, N13133, N5069);
xor XOR2 (N15275, N15267, N1178);
or OR2 (N15276, N15268, N3664);
nand NAND4 (N15277, N15276, N9154, N888, N3777);
buf BUF1 (N15278, N15272);
not NOT1 (N15279, N15263);
xor XOR2 (N15280, N15270, N5679);
and AND2 (N15281, N15280, N4616);
or OR2 (N15282, N15275, N5994);
xor XOR2 (N15283, N15273, N11181);
not NOT1 (N15284, N15282);
nor NOR3 (N15285, N15283, N518, N4393);
nand NAND4 (N15286, N15278, N66, N8498, N2414);
xor XOR2 (N15287, N15271, N6326);
nor NOR3 (N15288, N15281, N10529, N7936);
nand NAND2 (N15289, N15284, N14515);
and AND2 (N15290, N15265, N6335);
not NOT1 (N15291, N15289);
not NOT1 (N15292, N15277);
xor XOR2 (N15293, N15288, N11503);
nand NAND3 (N15294, N15279, N11462, N3149);
nand NAND3 (N15295, N15286, N9679, N5863);
or OR3 (N15296, N15285, N12215, N10380);
and AND2 (N15297, N15292, N15189);
not NOT1 (N15298, N15297);
nand NAND4 (N15299, N15298, N6924, N12089, N3069);
and AND2 (N15300, N15291, N8163);
or OR3 (N15301, N15294, N12934, N4860);
or OR2 (N15302, N15296, N12951);
nand NAND2 (N15303, N15301, N714);
nand NAND4 (N15304, N15293, N11493, N11126, N2410);
not NOT1 (N15305, N15295);
nor NOR3 (N15306, N15303, N8746, N3228);
xor XOR2 (N15307, N15304, N8575);
and AND3 (N15308, N15302, N12534, N1409);
buf BUF1 (N15309, N15258);
nand NAND4 (N15310, N15308, N8374, N7611, N3007);
and AND4 (N15311, N15274, N5579, N6016, N6366);
xor XOR2 (N15312, N15307, N2335);
nand NAND3 (N15313, N15290, N9419, N14891);
not NOT1 (N15314, N15299);
and AND3 (N15315, N15312, N13479, N5927);
buf BUF1 (N15316, N15309);
buf BUF1 (N15317, N15315);
or OR3 (N15318, N15305, N11486, N11587);
nor NOR4 (N15319, N15316, N11764, N14943, N6045);
not NOT1 (N15320, N15314);
xor XOR2 (N15321, N15311, N2221);
xor XOR2 (N15322, N15318, N1923);
buf BUF1 (N15323, N15313);
xor XOR2 (N15324, N15287, N8602);
buf BUF1 (N15325, N15323);
buf BUF1 (N15326, N15317);
not NOT1 (N15327, N15322);
or OR3 (N15328, N15306, N14859, N5577);
xor XOR2 (N15329, N15327, N14269);
and AND4 (N15330, N15319, N11615, N10280, N9154);
not NOT1 (N15331, N15325);
buf BUF1 (N15332, N15326);
and AND4 (N15333, N15321, N10395, N6648, N7209);
and AND3 (N15334, N15333, N10089, N13855);
not NOT1 (N15335, N15300);
nand NAND4 (N15336, N15335, N2572, N11035, N6408);
xor XOR2 (N15337, N15334, N3068);
xor XOR2 (N15338, N15328, N2445);
buf BUF1 (N15339, N15337);
not NOT1 (N15340, N15310);
not NOT1 (N15341, N15338);
or OR2 (N15342, N15330, N12619);
buf BUF1 (N15343, N15332);
nand NAND3 (N15344, N15342, N8032, N424);
not NOT1 (N15345, N15324);
and AND2 (N15346, N15341, N10879);
or OR4 (N15347, N15331, N5177, N13091, N8450);
nand NAND4 (N15348, N15336, N10301, N7879, N12027);
nand NAND2 (N15349, N15348, N9277);
nor NOR4 (N15350, N15346, N135, N3626, N12562);
xor XOR2 (N15351, N15349, N3937);
buf BUF1 (N15352, N15351);
or OR4 (N15353, N15344, N303, N14074, N9629);
not NOT1 (N15354, N15352);
or OR3 (N15355, N15353, N12324, N4019);
buf BUF1 (N15356, N15355);
or OR4 (N15357, N15340, N3538, N5195, N3576);
and AND4 (N15358, N15343, N1718, N2474, N11654);
nor NOR2 (N15359, N15357, N9132);
nand NAND3 (N15360, N15345, N8596, N219);
nand NAND2 (N15361, N15347, N5942);
or OR4 (N15362, N15320, N9913, N12439, N13180);
xor XOR2 (N15363, N15339, N13936);
or OR3 (N15364, N15361, N13202, N6635);
or OR2 (N15365, N15358, N10147);
not NOT1 (N15366, N15360);
buf BUF1 (N15367, N15329);
or OR3 (N15368, N15362, N11553, N114);
and AND4 (N15369, N15366, N11882, N3082, N8053);
not NOT1 (N15370, N15364);
and AND2 (N15371, N15356, N3786);
xor XOR2 (N15372, N15369, N4652);
not NOT1 (N15373, N15372);
or OR3 (N15374, N15367, N1287, N4091);
or OR3 (N15375, N15359, N9623, N11349);
nand NAND2 (N15376, N15373, N7149);
nand NAND2 (N15377, N15365, N12794);
nand NAND4 (N15378, N15375, N14742, N5918, N2488);
and AND4 (N15379, N15370, N1452, N2804, N6636);
not NOT1 (N15380, N15363);
buf BUF1 (N15381, N15374);
nand NAND3 (N15382, N15371, N8346, N6526);
nand NAND3 (N15383, N15368, N12523, N15068);
buf BUF1 (N15384, N15380);
nand NAND3 (N15385, N15350, N9933, N2157);
nand NAND4 (N15386, N15383, N13561, N5845, N1268);
xor XOR2 (N15387, N15377, N3426);
nor NOR2 (N15388, N15381, N455);
nor NOR4 (N15389, N15379, N10105, N12793, N9527);
or OR2 (N15390, N15386, N6940);
buf BUF1 (N15391, N15388);
nand NAND2 (N15392, N15385, N9438);
not NOT1 (N15393, N15378);
nor NOR2 (N15394, N15389, N12180);
xor XOR2 (N15395, N15392, N14943);
nor NOR4 (N15396, N15354, N3306, N12992, N13181);
and AND4 (N15397, N15396, N7029, N12903, N4640);
xor XOR2 (N15398, N15395, N8460);
not NOT1 (N15399, N15376);
buf BUF1 (N15400, N15394);
or OR4 (N15401, N15400, N7238, N3781, N9800);
xor XOR2 (N15402, N15397, N534);
nand NAND3 (N15403, N15399, N8856, N4330);
buf BUF1 (N15404, N15403);
nand NAND4 (N15405, N15391, N11155, N8879, N535);
nor NOR4 (N15406, N15387, N7499, N1560, N9162);
or OR2 (N15407, N15393, N882);
buf BUF1 (N15408, N15402);
or OR3 (N15409, N15407, N13934, N3538);
nand NAND2 (N15410, N15384, N14041);
nor NOR3 (N15411, N15382, N11143, N2957);
or OR3 (N15412, N15398, N2570, N6599);
nand NAND4 (N15413, N15411, N2885, N12650, N4788);
not NOT1 (N15414, N15404);
nor NOR3 (N15415, N15413, N1776, N279);
nor NOR2 (N15416, N15415, N11707);
not NOT1 (N15417, N15409);
nor NOR4 (N15418, N15412, N3612, N7035, N11669);
nand NAND4 (N15419, N15417, N12958, N9511, N13132);
and AND2 (N15420, N15416, N9439);
nor NOR4 (N15421, N15406, N944, N3026, N4895);
or OR4 (N15422, N15414, N9046, N12420, N3401);
and AND4 (N15423, N15420, N8838, N175, N2214);
and AND2 (N15424, N15421, N4474);
nor NOR4 (N15425, N15422, N12203, N14083, N4197);
xor XOR2 (N15426, N15410, N14346);
not NOT1 (N15427, N15401);
or OR3 (N15428, N15418, N427, N10261);
nor NOR3 (N15429, N15419, N4001, N10033);
and AND2 (N15430, N15428, N14262);
not NOT1 (N15431, N15405);
xor XOR2 (N15432, N15424, N10534);
nand NAND3 (N15433, N15425, N11378, N13201);
and AND3 (N15434, N15426, N311, N10047);
nand NAND3 (N15435, N15433, N4757, N4205);
nor NOR3 (N15436, N15423, N4052, N12497);
xor XOR2 (N15437, N15408, N1491);
nor NOR4 (N15438, N15437, N8793, N5299, N12252);
nor NOR3 (N15439, N15430, N1152, N9992);
or OR4 (N15440, N15436, N13590, N9130, N2340);
xor XOR2 (N15441, N15435, N6613);
not NOT1 (N15442, N15390);
nor NOR4 (N15443, N15429, N9485, N13174, N14535);
not NOT1 (N15444, N15432);
or OR3 (N15445, N15434, N4418, N7876);
or OR4 (N15446, N15440, N4378, N13085, N13975);
and AND2 (N15447, N15442, N15116);
nor NOR2 (N15448, N15441, N12468);
buf BUF1 (N15449, N15445);
buf BUF1 (N15450, N15448);
buf BUF1 (N15451, N15427);
buf BUF1 (N15452, N15438);
nor NOR3 (N15453, N15443, N2916, N15036);
nor NOR2 (N15454, N15450, N1114);
nor NOR3 (N15455, N15439, N7949, N446);
buf BUF1 (N15456, N15444);
not NOT1 (N15457, N15451);
buf BUF1 (N15458, N15457);
buf BUF1 (N15459, N15453);
not NOT1 (N15460, N15447);
nand NAND3 (N15461, N15431, N8741, N6867);
nand NAND2 (N15462, N15456, N4515);
and AND2 (N15463, N15446, N3636);
xor XOR2 (N15464, N15463, N13021);
nand NAND2 (N15465, N15462, N6565);
and AND3 (N15466, N15464, N3589, N9167);
not NOT1 (N15467, N15454);
buf BUF1 (N15468, N15466);
xor XOR2 (N15469, N15461, N12915);
nand NAND3 (N15470, N15469, N3909, N6984);
or OR2 (N15471, N15465, N10172);
xor XOR2 (N15472, N15470, N9622);
nor NOR2 (N15473, N15459, N12768);
xor XOR2 (N15474, N15473, N13795);
not NOT1 (N15475, N15460);
and AND4 (N15476, N15475, N13795, N5038, N9739);
and AND4 (N15477, N15472, N10397, N14771, N11198);
nand NAND4 (N15478, N15449, N15231, N11488, N12340);
nand NAND4 (N15479, N15478, N11898, N11994, N2169);
nor NOR3 (N15480, N15476, N8715, N4044);
nor NOR2 (N15481, N15479, N1250);
nor NOR2 (N15482, N15458, N8168);
xor XOR2 (N15483, N15471, N11240);
or OR4 (N15484, N15482, N13231, N1994, N5156);
not NOT1 (N15485, N15481);
nor NOR2 (N15486, N15480, N14471);
nand NAND3 (N15487, N15477, N11516, N4798);
nand NAND2 (N15488, N15485, N337);
and AND3 (N15489, N15455, N9403, N8951);
or OR2 (N15490, N15488, N10453);
buf BUF1 (N15491, N15474);
xor XOR2 (N15492, N15490, N12356);
buf BUF1 (N15493, N15489);
xor XOR2 (N15494, N15493, N5366);
nand NAND2 (N15495, N15468, N2619);
or OR2 (N15496, N15491, N6684);
nor NOR2 (N15497, N15452, N14788);
xor XOR2 (N15498, N15496, N5573);
nor NOR4 (N15499, N15492, N4944, N9272, N14501);
xor XOR2 (N15500, N15498, N5169);
and AND2 (N15501, N15467, N3371);
and AND2 (N15502, N15483, N3847);
not NOT1 (N15503, N15484);
and AND4 (N15504, N15501, N5863, N1619, N14324);
buf BUF1 (N15505, N15503);
and AND3 (N15506, N15502, N15021, N2736);
nor NOR4 (N15507, N15505, N14031, N14715, N1925);
buf BUF1 (N15508, N15506);
not NOT1 (N15509, N15499);
xor XOR2 (N15510, N15487, N13127);
or OR4 (N15511, N15510, N9515, N5765, N14136);
nor NOR2 (N15512, N15511, N225);
nor NOR3 (N15513, N15494, N1789, N12082);
buf BUF1 (N15514, N15512);
buf BUF1 (N15515, N15500);
or OR2 (N15516, N15513, N372);
nand NAND2 (N15517, N15495, N4431);
nand NAND2 (N15518, N15514, N1342);
nor NOR3 (N15519, N15516, N603, N10477);
xor XOR2 (N15520, N15508, N1259);
xor XOR2 (N15521, N15497, N5675);
xor XOR2 (N15522, N15509, N15106);
nand NAND3 (N15523, N15522, N7157, N12251);
xor XOR2 (N15524, N15523, N8821);
nor NOR3 (N15525, N15518, N98, N5292);
or OR3 (N15526, N15519, N7353, N8997);
xor XOR2 (N15527, N15524, N15508);
nand NAND3 (N15528, N15520, N11442, N7798);
nor NOR2 (N15529, N15515, N2726);
and AND4 (N15530, N15529, N1862, N12412, N3751);
not NOT1 (N15531, N15504);
buf BUF1 (N15532, N15525);
buf BUF1 (N15533, N15517);
or OR2 (N15534, N15530, N1480);
buf BUF1 (N15535, N15533);
or OR3 (N15536, N15526, N11216, N8477);
or OR2 (N15537, N15528, N3452);
nand NAND3 (N15538, N15521, N14094, N6844);
not NOT1 (N15539, N15536);
nand NAND2 (N15540, N15486, N4712);
and AND3 (N15541, N15531, N11693, N2330);
nand NAND4 (N15542, N15540, N14387, N3559, N5457);
xor XOR2 (N15543, N15537, N11295);
nand NAND3 (N15544, N15541, N8874, N11923);
nand NAND2 (N15545, N15535, N10798);
buf BUF1 (N15546, N15545);
xor XOR2 (N15547, N15538, N1999);
or OR2 (N15548, N15544, N4885);
nor NOR3 (N15549, N15547, N8539, N4550);
buf BUF1 (N15550, N15546);
or OR3 (N15551, N15534, N8259, N10598);
nand NAND2 (N15552, N15543, N6249);
buf BUF1 (N15553, N15548);
buf BUF1 (N15554, N15527);
xor XOR2 (N15555, N15539, N12375);
buf BUF1 (N15556, N15555);
not NOT1 (N15557, N15551);
xor XOR2 (N15558, N15557, N3399);
or OR3 (N15559, N15552, N12493, N1143);
not NOT1 (N15560, N15559);
nand NAND2 (N15561, N15560, N6491);
nor NOR2 (N15562, N15561, N14390);
and AND2 (N15563, N15542, N4099);
not NOT1 (N15564, N15563);
nand NAND3 (N15565, N15550, N14940, N2139);
xor XOR2 (N15566, N15565, N6187);
not NOT1 (N15567, N15532);
buf BUF1 (N15568, N15549);
not NOT1 (N15569, N15566);
xor XOR2 (N15570, N15554, N8591);
xor XOR2 (N15571, N15567, N14772);
nand NAND2 (N15572, N15562, N14613);
xor XOR2 (N15573, N15572, N14164);
and AND4 (N15574, N15573, N7587, N6493, N4213);
not NOT1 (N15575, N15568);
or OR3 (N15576, N15569, N10401, N9833);
nor NOR3 (N15577, N15570, N10580, N3835);
xor XOR2 (N15578, N15558, N8291);
not NOT1 (N15579, N15574);
or OR4 (N15580, N15577, N11343, N14165, N2430);
nand NAND2 (N15581, N15575, N7801);
not NOT1 (N15582, N15579);
buf BUF1 (N15583, N15581);
not NOT1 (N15584, N15507);
buf BUF1 (N15585, N15564);
buf BUF1 (N15586, N15571);
or OR3 (N15587, N15556, N15397, N12570);
and AND4 (N15588, N15586, N9819, N14878, N1039);
xor XOR2 (N15589, N15583, N10657);
nand NAND2 (N15590, N15578, N6624);
xor XOR2 (N15591, N15589, N12830);
and AND2 (N15592, N15582, N9331);
not NOT1 (N15593, N15591);
or OR2 (N15594, N15588, N7477);
or OR2 (N15595, N15553, N11172);
nand NAND4 (N15596, N15595, N8919, N797, N1349);
and AND3 (N15597, N15596, N7646, N11707);
or OR3 (N15598, N15584, N2486, N9511);
or OR3 (N15599, N15576, N14094, N2620);
nor NOR2 (N15600, N15580, N9575);
not NOT1 (N15601, N15599);
xor XOR2 (N15602, N15597, N8595);
buf BUF1 (N15603, N15592);
nand NAND4 (N15604, N15601, N6349, N3421, N12217);
not NOT1 (N15605, N15604);
and AND3 (N15606, N15590, N9029, N8964);
nor NOR4 (N15607, N15593, N103, N6188, N4857);
xor XOR2 (N15608, N15603, N11034);
nand NAND4 (N15609, N15602, N8296, N12015, N6069);
not NOT1 (N15610, N15608);
nand NAND3 (N15611, N15606, N9542, N2419);
or OR2 (N15612, N15605, N6692);
nor NOR3 (N15613, N15610, N12221, N4043);
nand NAND3 (N15614, N15598, N1682, N9447);
or OR3 (N15615, N15587, N11839, N11357);
xor XOR2 (N15616, N15612, N13664);
not NOT1 (N15617, N15614);
buf BUF1 (N15618, N15617);
nor NOR4 (N15619, N15616, N12740, N3185, N1462);
and AND3 (N15620, N15618, N5209, N6287);
nand NAND3 (N15621, N15594, N11084, N10619);
nor NOR2 (N15622, N15619, N15465);
and AND2 (N15623, N15609, N868);
xor XOR2 (N15624, N15620, N7051);
nor NOR4 (N15625, N15622, N2209, N11697, N6912);
buf BUF1 (N15626, N15607);
not NOT1 (N15627, N15600);
not NOT1 (N15628, N15625);
and AND4 (N15629, N15624, N10405, N14916, N12267);
not NOT1 (N15630, N15626);
buf BUF1 (N15631, N15629);
not NOT1 (N15632, N15615);
and AND2 (N15633, N15632, N657);
and AND2 (N15634, N15623, N281);
nand NAND3 (N15635, N15630, N5660, N5516);
not NOT1 (N15636, N15631);
not NOT1 (N15637, N15634);
or OR4 (N15638, N15635, N7856, N7967, N4567);
or OR2 (N15639, N15638, N4914);
nor NOR4 (N15640, N15636, N6802, N5705, N1934);
and AND2 (N15641, N15639, N5745);
not NOT1 (N15642, N15640);
buf BUF1 (N15643, N15641);
or OR3 (N15644, N15627, N7994, N10464);
not NOT1 (N15645, N15642);
buf BUF1 (N15646, N15645);
nand NAND2 (N15647, N15646, N2109);
not NOT1 (N15648, N15585);
xor XOR2 (N15649, N15633, N13494);
nor NOR3 (N15650, N15621, N7693, N4223);
buf BUF1 (N15651, N15637);
xor XOR2 (N15652, N15628, N3778);
nand NAND3 (N15653, N15650, N6174, N13935);
not NOT1 (N15654, N15611);
or OR4 (N15655, N15613, N4442, N7857, N2521);
buf BUF1 (N15656, N15649);
xor XOR2 (N15657, N15653, N10695);
not NOT1 (N15658, N15656);
nand NAND2 (N15659, N15644, N9986);
xor XOR2 (N15660, N15659, N8410);
not NOT1 (N15661, N15658);
not NOT1 (N15662, N15660);
or OR3 (N15663, N15655, N11830, N6045);
nand NAND4 (N15664, N15661, N10051, N4527, N11694);
buf BUF1 (N15665, N15651);
or OR2 (N15666, N15652, N829);
nor NOR4 (N15667, N15643, N8410, N12306, N5424);
or OR4 (N15668, N15664, N8987, N10208, N14886);
buf BUF1 (N15669, N15663);
not NOT1 (N15670, N15654);
nand NAND3 (N15671, N15670, N7647, N11456);
and AND2 (N15672, N15668, N4603);
nand NAND3 (N15673, N15662, N12869, N2739);
nand NAND2 (N15674, N15672, N12187);
or OR2 (N15675, N15674, N10988);
not NOT1 (N15676, N15665);
nand NAND3 (N15677, N15669, N10830, N8991);
or OR3 (N15678, N15671, N284, N15523);
buf BUF1 (N15679, N15648);
nand NAND2 (N15680, N15678, N14254);
or OR4 (N15681, N15673, N7905, N9984, N12904);
nand NAND2 (N15682, N15681, N1452);
nand NAND3 (N15683, N15667, N6160, N8275);
buf BUF1 (N15684, N15657);
or OR4 (N15685, N15675, N8952, N9544, N10219);
or OR4 (N15686, N15685, N12713, N7539, N13152);
xor XOR2 (N15687, N15647, N11450);
not NOT1 (N15688, N15677);
buf BUF1 (N15689, N15684);
nand NAND3 (N15690, N15686, N9146, N2113);
nor NOR4 (N15691, N15679, N8926, N10016, N8174);
nor NOR2 (N15692, N15687, N4034);
nor NOR3 (N15693, N15682, N11545, N8683);
not NOT1 (N15694, N15683);
buf BUF1 (N15695, N15690);
buf BUF1 (N15696, N15695);
not NOT1 (N15697, N15666);
not NOT1 (N15698, N15692);
not NOT1 (N15699, N15697);
xor XOR2 (N15700, N15699, N3446);
nand NAND2 (N15701, N15694, N5843);
or OR2 (N15702, N15693, N5786);
nor NOR2 (N15703, N15676, N812);
and AND2 (N15704, N15701, N15558);
nand NAND4 (N15705, N15702, N6774, N12890, N9780);
xor XOR2 (N15706, N15705, N3058);
or OR2 (N15707, N15691, N14531);
and AND2 (N15708, N15704, N12913);
or OR2 (N15709, N15688, N7079);
nand NAND3 (N15710, N15708, N11791, N10124);
and AND3 (N15711, N15709, N1968, N1065);
buf BUF1 (N15712, N15710);
or OR2 (N15713, N15698, N4288);
and AND3 (N15714, N15703, N295, N8116);
not NOT1 (N15715, N15712);
or OR4 (N15716, N15713, N1481, N4243, N8106);
nor NOR3 (N15717, N15706, N14742, N96);
and AND4 (N15718, N15711, N3880, N12527, N11494);
nand NAND2 (N15719, N15696, N10465);
or OR2 (N15720, N15719, N6171);
xor XOR2 (N15721, N15680, N13686);
not NOT1 (N15722, N15714);
and AND2 (N15723, N15717, N14464);
buf BUF1 (N15724, N15723);
not NOT1 (N15725, N15718);
nor NOR4 (N15726, N15721, N5092, N4077, N15386);
xor XOR2 (N15727, N15716, N990);
xor XOR2 (N15728, N15715, N10916);
nor NOR4 (N15729, N15725, N6320, N174, N421);
nand NAND4 (N15730, N15728, N1159, N415, N13621);
not NOT1 (N15731, N15707);
or OR2 (N15732, N15722, N8795);
or OR2 (N15733, N15720, N3384);
buf BUF1 (N15734, N15733);
xor XOR2 (N15735, N15724, N391);
or OR3 (N15736, N15735, N14959, N3753);
not NOT1 (N15737, N15734);
xor XOR2 (N15738, N15732, N10740);
buf BUF1 (N15739, N15730);
or OR3 (N15740, N15727, N12426, N7027);
not NOT1 (N15741, N15738);
or OR4 (N15742, N15700, N2108, N304, N3077);
xor XOR2 (N15743, N15739, N13942);
nor NOR4 (N15744, N15743, N1964, N5061, N1220);
not NOT1 (N15745, N15729);
not NOT1 (N15746, N15726);
not NOT1 (N15747, N15731);
nand NAND3 (N15748, N15740, N10056, N909);
not NOT1 (N15749, N15744);
not NOT1 (N15750, N15736);
buf BUF1 (N15751, N15741);
buf BUF1 (N15752, N15745);
and AND2 (N15753, N15746, N15419);
xor XOR2 (N15754, N15751, N1164);
buf BUF1 (N15755, N15689);
buf BUF1 (N15756, N15755);
and AND3 (N15757, N15756, N6057, N573);
not NOT1 (N15758, N15749);
nor NOR3 (N15759, N15757, N15438, N14065);
xor XOR2 (N15760, N15752, N12677);
and AND4 (N15761, N15747, N7534, N6960, N13561);
or OR3 (N15762, N15748, N2934, N13201);
and AND3 (N15763, N15754, N4588, N2244);
not NOT1 (N15764, N15763);
not NOT1 (N15765, N15761);
nand NAND4 (N15766, N15737, N15745, N12620, N11206);
or OR2 (N15767, N15764, N10299);
not NOT1 (N15768, N15760);
xor XOR2 (N15769, N15766, N15229);
nor NOR2 (N15770, N15750, N7415);
nor NOR2 (N15771, N15765, N5065);
xor XOR2 (N15772, N15769, N9026);
or OR3 (N15773, N15762, N1634, N8303);
buf BUF1 (N15774, N15759);
nand NAND3 (N15775, N15753, N13404, N8298);
nand NAND2 (N15776, N15770, N9893);
xor XOR2 (N15777, N15767, N2084);
nor NOR3 (N15778, N15771, N686, N2526);
not NOT1 (N15779, N15758);
or OR4 (N15780, N15768, N2146, N4194, N1041);
and AND3 (N15781, N15777, N11733, N3636);
nand NAND2 (N15782, N15779, N4169);
nand NAND4 (N15783, N15782, N7049, N2028, N2750);
buf BUF1 (N15784, N15772);
not NOT1 (N15785, N15778);
not NOT1 (N15786, N15774);
and AND4 (N15787, N15781, N14332, N13621, N365);
and AND2 (N15788, N15784, N15186);
not NOT1 (N15789, N15776);
nor NOR3 (N15790, N15789, N8091, N756);
xor XOR2 (N15791, N15773, N8342);
buf BUF1 (N15792, N15790);
buf BUF1 (N15793, N15783);
nand NAND2 (N15794, N15793, N15273);
not NOT1 (N15795, N15794);
not NOT1 (N15796, N15742);
or OR2 (N15797, N15786, N10417);
nand NAND3 (N15798, N15792, N13292, N2234);
and AND3 (N15799, N15780, N8626, N6094);
nand NAND4 (N15800, N15795, N7554, N10152, N11413);
not NOT1 (N15801, N15791);
xor XOR2 (N15802, N15800, N10765);
or OR2 (N15803, N15798, N15423);
and AND2 (N15804, N15803, N9765);
and AND2 (N15805, N15802, N4699);
xor XOR2 (N15806, N15805, N8542);
xor XOR2 (N15807, N15804, N4036);
xor XOR2 (N15808, N15801, N8257);
nand NAND4 (N15809, N15775, N626, N598, N10061);
and AND3 (N15810, N15797, N2908, N9036);
nand NAND2 (N15811, N15806, N8807);
and AND4 (N15812, N15799, N14835, N7013, N5516);
nand NAND4 (N15813, N15809, N5081, N11396, N6973);
and AND4 (N15814, N15808, N7451, N8517, N6762);
and AND2 (N15815, N15812, N13603);
not NOT1 (N15816, N15815);
xor XOR2 (N15817, N15816, N11580);
xor XOR2 (N15818, N15788, N10211);
not NOT1 (N15819, N15818);
or OR3 (N15820, N15813, N3774, N6475);
nor NOR3 (N15821, N15787, N11623, N2635);
buf BUF1 (N15822, N15807);
not NOT1 (N15823, N15821);
or OR2 (N15824, N15814, N4780);
buf BUF1 (N15825, N15822);
nor NOR4 (N15826, N15785, N7773, N2556, N5337);
or OR4 (N15827, N15824, N5121, N7773, N11788);
xor XOR2 (N15828, N15810, N9510);
buf BUF1 (N15829, N15796);
or OR3 (N15830, N15827, N8105, N8920);
buf BUF1 (N15831, N15811);
or OR2 (N15832, N15831, N1002);
buf BUF1 (N15833, N15829);
nor NOR2 (N15834, N15826, N14461);
nand NAND4 (N15835, N15823, N7237, N4928, N10110);
buf BUF1 (N15836, N15828);
buf BUF1 (N15837, N15830);
buf BUF1 (N15838, N15825);
or OR4 (N15839, N15817, N5248, N9666, N9540);
not NOT1 (N15840, N15839);
or OR2 (N15841, N15840, N2422);
nand NAND3 (N15842, N15819, N15730, N9224);
and AND2 (N15843, N15841, N326);
nor NOR2 (N15844, N15843, N6824);
nor NOR2 (N15845, N15836, N5438);
nor NOR2 (N15846, N15845, N2207);
buf BUF1 (N15847, N15832);
or OR3 (N15848, N15847, N8694, N2867);
not NOT1 (N15849, N15834);
or OR3 (N15850, N15846, N4012, N1346);
not NOT1 (N15851, N15849);
nor NOR2 (N15852, N15838, N14744);
xor XOR2 (N15853, N15848, N4511);
nor NOR3 (N15854, N15820, N15452, N15468);
xor XOR2 (N15855, N15854, N5208);
not NOT1 (N15856, N15852);
buf BUF1 (N15857, N15856);
or OR2 (N15858, N15851, N11405);
buf BUF1 (N15859, N15835);
or OR2 (N15860, N15837, N6717);
or OR2 (N15861, N15860, N12648);
buf BUF1 (N15862, N15859);
buf BUF1 (N15863, N15853);
buf BUF1 (N15864, N15862);
or OR3 (N15865, N15858, N1959, N5919);
not NOT1 (N15866, N15833);
not NOT1 (N15867, N15855);
or OR2 (N15868, N15844, N13282);
or OR3 (N15869, N15864, N182, N5893);
buf BUF1 (N15870, N15868);
nor NOR3 (N15871, N15850, N2881, N9536);
nor NOR3 (N15872, N15857, N5754, N1686);
buf BUF1 (N15873, N15869);
nand NAND4 (N15874, N15867, N13828, N14230, N15167);
and AND3 (N15875, N15863, N14702, N10501);
buf BUF1 (N15876, N15874);
nand NAND2 (N15877, N15865, N14303);
and AND2 (N15878, N15872, N11089);
buf BUF1 (N15879, N15873);
or OR4 (N15880, N15875, N5567, N7149, N2302);
not NOT1 (N15881, N15876);
nor NOR4 (N15882, N15870, N6639, N15093, N6780);
buf BUF1 (N15883, N15866);
or OR4 (N15884, N15871, N13078, N9496, N10758);
xor XOR2 (N15885, N15881, N12363);
or OR4 (N15886, N15883, N7240, N11207, N1224);
or OR2 (N15887, N15880, N8562);
buf BUF1 (N15888, N15886);
nor NOR4 (N15889, N15887, N7564, N592, N6125);
and AND2 (N15890, N15884, N9195);
xor XOR2 (N15891, N15877, N13251);
or OR3 (N15892, N15878, N9860, N1393);
not NOT1 (N15893, N15890);
not NOT1 (N15894, N15885);
buf BUF1 (N15895, N15891);
or OR3 (N15896, N15888, N12144, N3028);
or OR2 (N15897, N15894, N5007);
nand NAND2 (N15898, N15892, N8725);
xor XOR2 (N15899, N15879, N11238);
buf BUF1 (N15900, N15897);
nor NOR4 (N15901, N15896, N15473, N13884, N13189);
nor NOR2 (N15902, N15893, N1522);
nor NOR3 (N15903, N15899, N4019, N4485);
nor NOR4 (N15904, N15895, N11938, N5934, N7054);
and AND3 (N15905, N15904, N13796, N3308);
nand NAND2 (N15906, N15902, N11069);
or OR4 (N15907, N15898, N12417, N13822, N9886);
xor XOR2 (N15908, N15861, N1136);
and AND2 (N15909, N15903, N1863);
and AND3 (N15910, N15901, N9594, N2340);
or OR2 (N15911, N15905, N13576);
not NOT1 (N15912, N15906);
and AND3 (N15913, N15910, N12725, N7306);
and AND3 (N15914, N15908, N10, N6700);
nand NAND2 (N15915, N15882, N5150);
nand NAND2 (N15916, N15889, N3355);
and AND4 (N15917, N15912, N8286, N2038, N11715);
and AND4 (N15918, N15911, N1530, N14798, N4174);
nor NOR2 (N15919, N15913, N13719);
nand NAND2 (N15920, N15914, N12448);
xor XOR2 (N15921, N15918, N6727);
buf BUF1 (N15922, N15916);
and AND4 (N15923, N15909, N2954, N3297, N15398);
xor XOR2 (N15924, N15917, N13955);
xor XOR2 (N15925, N15921, N4872);
and AND2 (N15926, N15924, N5101);
and AND4 (N15927, N15842, N13543, N10808, N15790);
not NOT1 (N15928, N15926);
nand NAND2 (N15929, N15922, N12547);
not NOT1 (N15930, N15927);
buf BUF1 (N15931, N15920);
not NOT1 (N15932, N15900);
or OR3 (N15933, N15923, N9281, N3762);
and AND3 (N15934, N15929, N15399, N1404);
buf BUF1 (N15935, N15925);
nor NOR2 (N15936, N15928, N14877);
nand NAND3 (N15937, N15933, N7439, N4652);
and AND4 (N15938, N15915, N3873, N11411, N13394);
or OR2 (N15939, N15935, N1304);
buf BUF1 (N15940, N15930);
nor NOR4 (N15941, N15936, N6145, N2792, N14754);
buf BUF1 (N15942, N15932);
not NOT1 (N15943, N15940);
xor XOR2 (N15944, N15938, N7622);
nand NAND4 (N15945, N15934, N1516, N3962, N4922);
nand NAND3 (N15946, N15945, N13783, N7425);
or OR2 (N15947, N15919, N2693);
xor XOR2 (N15948, N15931, N3128);
nand NAND4 (N15949, N15942, N11701, N12174, N13309);
not NOT1 (N15950, N15944);
buf BUF1 (N15951, N15939);
not NOT1 (N15952, N15943);
buf BUF1 (N15953, N15907);
or OR2 (N15954, N15946, N9186);
nand NAND2 (N15955, N15948, N2127);
or OR4 (N15956, N15941, N12227, N10633, N2845);
not NOT1 (N15957, N15954);
not NOT1 (N15958, N15953);
or OR2 (N15959, N15951, N13566);
nor NOR3 (N15960, N15958, N8492, N8846);
xor XOR2 (N15961, N15952, N3260);
and AND3 (N15962, N15950, N2998, N7778);
and AND2 (N15963, N15959, N631);
nand NAND2 (N15964, N15960, N9919);
nor NOR2 (N15965, N15963, N12684);
not NOT1 (N15966, N15949);
or OR4 (N15967, N15955, N14989, N4500, N12312);
not NOT1 (N15968, N15961);
not NOT1 (N15969, N15965);
not NOT1 (N15970, N15964);
nor NOR3 (N15971, N15957, N14842, N13171);
xor XOR2 (N15972, N15968, N151);
or OR2 (N15973, N15937, N11519);
nor NOR3 (N15974, N15966, N15833, N4227);
and AND3 (N15975, N15947, N5429, N227);
xor XOR2 (N15976, N15972, N7206);
xor XOR2 (N15977, N15973, N15907);
and AND4 (N15978, N15970, N11325, N1867, N6867);
not NOT1 (N15979, N15974);
nor NOR2 (N15980, N15962, N13529);
not NOT1 (N15981, N15980);
and AND2 (N15982, N15981, N2310);
or OR3 (N15983, N15971, N9225, N10593);
or OR4 (N15984, N15982, N8210, N7388, N8642);
or OR3 (N15985, N15976, N2757, N14102);
buf BUF1 (N15986, N15985);
not NOT1 (N15987, N15967);
buf BUF1 (N15988, N15977);
nand NAND4 (N15989, N15986, N15494, N11027, N15380);
not NOT1 (N15990, N15988);
or OR2 (N15991, N15969, N5570);
and AND2 (N15992, N15990, N9884);
xor XOR2 (N15993, N15984, N1491);
or OR2 (N15994, N15987, N10972);
not NOT1 (N15995, N15978);
and AND2 (N15996, N15992, N7867);
not NOT1 (N15997, N15991);
nor NOR4 (N15998, N15997, N2861, N7123, N12220);
or OR2 (N15999, N15996, N956);
xor XOR2 (N16000, N15975, N10273);
nand NAND3 (N16001, N15956, N7417, N5469);
nor NOR4 (N16002, N15993, N15698, N5342, N7560);
nand NAND4 (N16003, N16002, N4173, N5797, N11305);
not NOT1 (N16004, N16000);
buf BUF1 (N16005, N16004);
and AND2 (N16006, N15979, N13315);
not NOT1 (N16007, N16006);
nand NAND4 (N16008, N15998, N13936, N7139, N1303);
not NOT1 (N16009, N16007);
nand NAND2 (N16010, N15983, N2266);
nor NOR3 (N16011, N15989, N4068, N11169);
or OR4 (N16012, N16011, N829, N10480, N10136);
endmodule