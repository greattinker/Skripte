// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23;

output N911,N919,N904,N922,N921,N918,N897,N917,N913,N923;

or OR3 (N24, N12, N15, N15);
buf BUF1 (N25, N15);
xor XOR2 (N26, N7, N22);
and AND2 (N27, N10, N22);
not NOT1 (N28, N21);
nor NOR3 (N29, N10, N4, N21);
or OR2 (N30, N3, N3);
and AND3 (N31, N22, N5, N24);
buf BUF1 (N32, N25);
nor NOR4 (N33, N25, N11, N21, N24);
not NOT1 (N34, N17);
buf BUF1 (N35, N29);
nor NOR3 (N36, N19, N21, N2);
or OR4 (N37, N28, N11, N14, N18);
nor NOR3 (N38, N33, N24, N14);
nand NAND2 (N39, N35, N3);
xor XOR2 (N40, N37, N7);
or OR4 (N41, N40, N34, N29, N23);
buf BUF1 (N42, N22);
nor NOR3 (N43, N41, N14, N37);
xor XOR2 (N44, N43, N9);
nor NOR3 (N45, N44, N43, N18);
buf BUF1 (N46, N32);
not NOT1 (N47, N39);
or OR2 (N48, N26, N21);
nor NOR2 (N49, N48, N28);
nand NAND2 (N50, N30, N4);
xor XOR2 (N51, N27, N6);
or OR2 (N52, N46, N45);
nand NAND3 (N53, N44, N10, N10);
and AND3 (N54, N53, N31, N4);
nand NAND3 (N55, N52, N40, N4);
nor NOR2 (N56, N4, N20);
nor NOR4 (N57, N42, N38, N6, N33);
xor XOR2 (N58, N15, N22);
or OR3 (N59, N36, N7, N21);
xor XOR2 (N60, N55, N52);
and AND3 (N61, N59, N15, N34);
buf BUF1 (N62, N51);
xor XOR2 (N63, N57, N39);
and AND2 (N64, N54, N34);
nor NOR4 (N65, N60, N37, N15, N18);
and AND2 (N66, N61, N35);
and AND4 (N67, N66, N49, N25, N58);
buf BUF1 (N68, N65);
xor XOR2 (N69, N9, N7);
not NOT1 (N70, N31);
xor XOR2 (N71, N47, N19);
nor NOR3 (N72, N64, N40, N47);
nand NAND2 (N73, N69, N33);
buf BUF1 (N74, N50);
or OR3 (N75, N67, N30, N18);
buf BUF1 (N76, N68);
xor XOR2 (N77, N71, N21);
nor NOR2 (N78, N74, N36);
buf BUF1 (N79, N70);
nor NOR2 (N80, N79, N59);
not NOT1 (N81, N80);
xor XOR2 (N82, N75, N55);
xor XOR2 (N83, N63, N55);
nor NOR2 (N84, N73, N65);
nand NAND3 (N85, N77, N26, N22);
nand NAND3 (N86, N76, N15, N63);
not NOT1 (N87, N85);
not NOT1 (N88, N82);
and AND2 (N89, N86, N73);
nand NAND3 (N90, N56, N3, N87);
or OR2 (N91, N23, N74);
and AND2 (N92, N91, N48);
nand NAND3 (N93, N90, N54, N35);
nand NAND3 (N94, N72, N63, N8);
xor XOR2 (N95, N83, N30);
nor NOR2 (N96, N62, N71);
and AND4 (N97, N96, N46, N12, N80);
not NOT1 (N98, N78);
buf BUF1 (N99, N81);
nor NOR3 (N100, N93, N82, N17);
or OR4 (N101, N88, N48, N4, N72);
xor XOR2 (N102, N98, N58);
xor XOR2 (N103, N95, N84);
xor XOR2 (N104, N90, N34);
buf BUF1 (N105, N101);
nand NAND3 (N106, N94, N22, N14);
not NOT1 (N107, N103);
xor XOR2 (N108, N100, N36);
nor NOR2 (N109, N108, N23);
and AND3 (N110, N89, N61, N11);
nor NOR3 (N111, N97, N19, N42);
and AND3 (N112, N109, N60, N15);
nand NAND3 (N113, N110, N13, N40);
nand NAND4 (N114, N106, N19, N86, N47);
nand NAND2 (N115, N107, N113);
nor NOR4 (N116, N113, N35, N108, N48);
not NOT1 (N117, N102);
nand NAND2 (N118, N117, N88);
xor XOR2 (N119, N116, N64);
xor XOR2 (N120, N92, N88);
nor NOR4 (N121, N114, N109, N64, N75);
or OR3 (N122, N121, N65, N103);
not NOT1 (N123, N104);
nand NAND3 (N124, N119, N9, N123);
nand NAND2 (N125, N57, N48);
or OR3 (N126, N125, N30, N111);
nor NOR2 (N127, N56, N7);
nor NOR2 (N128, N105, N2);
xor XOR2 (N129, N127, N74);
or OR3 (N130, N128, N91, N30);
or OR2 (N131, N118, N49);
nor NOR4 (N132, N122, N87, N39, N79);
nor NOR3 (N133, N132, N75, N63);
buf BUF1 (N134, N99);
xor XOR2 (N135, N129, N114);
and AND2 (N136, N135, N131);
or OR4 (N137, N14, N11, N62, N76);
nor NOR4 (N138, N137, N91, N77, N119);
nand NAND2 (N139, N126, N97);
or OR3 (N140, N138, N55, N120);
nand NAND2 (N141, N101, N55);
xor XOR2 (N142, N130, N86);
buf BUF1 (N143, N142);
not NOT1 (N144, N124);
xor XOR2 (N145, N140, N82);
and AND4 (N146, N141, N85, N54, N61);
nand NAND2 (N147, N115, N17);
or OR3 (N148, N144, N117, N81);
nor NOR4 (N149, N148, N45, N35, N146);
not NOT1 (N150, N76);
xor XOR2 (N151, N134, N130);
not NOT1 (N152, N136);
nand NAND3 (N153, N147, N113, N21);
nor NOR2 (N154, N139, N16);
xor XOR2 (N155, N149, N112);
xor XOR2 (N156, N4, N32);
buf BUF1 (N157, N143);
xor XOR2 (N158, N154, N14);
buf BUF1 (N159, N151);
buf BUF1 (N160, N157);
xor XOR2 (N161, N152, N15);
nand NAND3 (N162, N155, N16, N68);
not NOT1 (N163, N160);
nand NAND2 (N164, N161, N96);
not NOT1 (N165, N159);
buf BUF1 (N166, N153);
and AND4 (N167, N165, N83, N40, N40);
nor NOR2 (N168, N150, N167);
not NOT1 (N169, N71);
not NOT1 (N170, N169);
not NOT1 (N171, N158);
and AND4 (N172, N168, N65, N50, N166);
not NOT1 (N173, N82);
nand NAND2 (N174, N172, N14);
and AND3 (N175, N171, N4, N27);
nor NOR3 (N176, N156, N132, N114);
and AND4 (N177, N173, N89, N83, N149);
nor NOR3 (N178, N170, N172, N135);
and AND4 (N179, N175, N49, N150, N165);
nor NOR3 (N180, N176, N5, N96);
or OR3 (N181, N174, N173, N88);
nor NOR2 (N182, N162, N108);
nand NAND3 (N183, N180, N136, N20);
buf BUF1 (N184, N183);
xor XOR2 (N185, N163, N85);
xor XOR2 (N186, N185, N42);
or OR4 (N187, N178, N51, N101, N168);
and AND3 (N188, N133, N85, N186);
buf BUF1 (N189, N1);
nand NAND2 (N190, N182, N36);
xor XOR2 (N191, N181, N168);
buf BUF1 (N192, N187);
or OR3 (N193, N177, N171, N95);
buf BUF1 (N194, N184);
xor XOR2 (N195, N164, N152);
nor NOR2 (N196, N188, N145);
and AND4 (N197, N139, N190, N98, N107);
nor NOR2 (N198, N18, N47);
buf BUF1 (N199, N189);
buf BUF1 (N200, N179);
nand NAND2 (N201, N198, N162);
or OR4 (N202, N201, N32, N43, N179);
nor NOR2 (N203, N192, N1);
and AND4 (N204, N193, N124, N203, N29);
or OR3 (N205, N98, N95, N3);
buf BUF1 (N206, N191);
xor XOR2 (N207, N197, N33);
nand NAND4 (N208, N202, N72, N187, N127);
not NOT1 (N209, N208);
or OR2 (N210, N206, N84);
nand NAND4 (N211, N195, N70, N71, N38);
and AND3 (N212, N205, N123, N197);
nand NAND3 (N213, N210, N64, N62);
buf BUF1 (N214, N199);
buf BUF1 (N215, N200);
nand NAND3 (N216, N215, N179, N98);
xor XOR2 (N217, N194, N96);
xor XOR2 (N218, N207, N36);
buf BUF1 (N219, N209);
and AND3 (N220, N212, N106, N110);
buf BUF1 (N221, N214);
xor XOR2 (N222, N196, N47);
or OR2 (N223, N216, N204);
nor NOR3 (N224, N144, N143, N16);
and AND4 (N225, N218, N3, N11, N115);
or OR3 (N226, N211, N200, N140);
not NOT1 (N227, N219);
nor NOR4 (N228, N227, N88, N152, N12);
nand NAND4 (N229, N223, N53, N66, N41);
nor NOR3 (N230, N229, N1, N165);
not NOT1 (N231, N224);
or OR2 (N232, N230, N57);
nand NAND2 (N233, N228, N167);
not NOT1 (N234, N231);
and AND4 (N235, N225, N181, N70, N25);
and AND3 (N236, N217, N69, N186);
xor XOR2 (N237, N220, N15);
xor XOR2 (N238, N236, N117);
not NOT1 (N239, N238);
nand NAND4 (N240, N234, N35, N95, N189);
nor NOR3 (N241, N232, N57, N175);
or OR3 (N242, N213, N219, N221);
nor NOR4 (N243, N190, N46, N24, N139);
and AND3 (N244, N241, N92, N175);
nor NOR4 (N245, N235, N217, N71, N51);
and AND3 (N246, N240, N175, N165);
nand NAND4 (N247, N222, N242, N63, N156);
not NOT1 (N248, N196);
or OR3 (N249, N244, N207, N165);
and AND3 (N250, N226, N76, N191);
nand NAND3 (N251, N233, N140, N9);
nor NOR4 (N252, N249, N51, N67, N35);
nor NOR4 (N253, N248, N245, N48, N199);
nor NOR4 (N254, N202, N71, N148, N15);
nor NOR4 (N255, N237, N24, N8, N131);
not NOT1 (N256, N250);
nor NOR4 (N257, N246, N216, N123, N41);
xor XOR2 (N258, N247, N159);
nand NAND4 (N259, N239, N92, N139, N17);
nor NOR4 (N260, N251, N36, N163, N99);
nand NAND4 (N261, N243, N11, N16, N104);
nand NAND3 (N262, N259, N40, N54);
and AND4 (N263, N254, N10, N201, N160);
nor NOR3 (N264, N260, N47, N43);
nor NOR2 (N265, N264, N263);
nor NOR4 (N266, N55, N14, N29, N211);
nand NAND4 (N267, N252, N90, N200, N246);
xor XOR2 (N268, N265, N178);
and AND3 (N269, N256, N48, N33);
and AND2 (N270, N257, N30);
not NOT1 (N271, N253);
and AND3 (N272, N262, N130, N118);
and AND2 (N273, N258, N150);
buf BUF1 (N274, N255);
and AND3 (N275, N273, N262, N165);
xor XOR2 (N276, N270, N261);
buf BUF1 (N277, N176);
nand NAND3 (N278, N266, N258, N96);
or OR3 (N279, N274, N51, N227);
or OR2 (N280, N272, N97);
not NOT1 (N281, N277);
nor NOR2 (N282, N269, N276);
not NOT1 (N283, N168);
nor NOR2 (N284, N267, N277);
nor NOR3 (N285, N284, N19, N23);
and AND3 (N286, N271, N151, N278);
nor NOR3 (N287, N168, N77, N179);
xor XOR2 (N288, N286, N283);
buf BUF1 (N289, N191);
nand NAND4 (N290, N281, N20, N176, N278);
and AND4 (N291, N280, N172, N276, N263);
nand NAND4 (N292, N288, N78, N108, N245);
buf BUF1 (N293, N268);
xor XOR2 (N294, N282, N168);
nand NAND2 (N295, N285, N201);
or OR4 (N296, N275, N90, N247, N54);
or OR3 (N297, N295, N237, N87);
not NOT1 (N298, N296);
nor NOR2 (N299, N290, N57);
and AND4 (N300, N299, N73, N155, N297);
nor NOR3 (N301, N219, N270, N243);
xor XOR2 (N302, N293, N124);
xor XOR2 (N303, N298, N189);
not NOT1 (N304, N291);
not NOT1 (N305, N287);
not NOT1 (N306, N305);
buf BUF1 (N307, N300);
or OR3 (N308, N307, N167, N126);
buf BUF1 (N309, N301);
nor NOR3 (N310, N289, N271, N252);
and AND4 (N311, N302, N135, N193, N45);
not NOT1 (N312, N294);
not NOT1 (N313, N303);
and AND3 (N314, N312, N25, N278);
not NOT1 (N315, N292);
buf BUF1 (N316, N309);
not NOT1 (N317, N310);
or OR3 (N318, N304, N63, N95);
and AND4 (N319, N318, N244, N152, N236);
nand NAND3 (N320, N315, N270, N97);
nand NAND4 (N321, N279, N213, N64, N45);
nor NOR3 (N322, N311, N305, N127);
nand NAND2 (N323, N306, N135);
or OR2 (N324, N308, N251);
xor XOR2 (N325, N323, N276);
xor XOR2 (N326, N313, N246);
xor XOR2 (N327, N322, N239);
or OR3 (N328, N321, N153, N266);
nor NOR2 (N329, N328, N126);
or OR3 (N330, N329, N176, N275);
nor NOR3 (N331, N314, N29, N38);
buf BUF1 (N332, N330);
or OR2 (N333, N316, N1);
and AND2 (N334, N319, N42);
not NOT1 (N335, N317);
nand NAND4 (N336, N334, N203, N187, N138);
and AND4 (N337, N336, N96, N170, N171);
not NOT1 (N338, N327);
or OR3 (N339, N320, N141, N54);
not NOT1 (N340, N339);
and AND2 (N341, N325, N152);
xor XOR2 (N342, N340, N267);
nor NOR3 (N343, N333, N290, N148);
buf BUF1 (N344, N326);
not NOT1 (N345, N344);
not NOT1 (N346, N343);
or OR4 (N347, N346, N42, N149, N297);
xor XOR2 (N348, N335, N60);
buf BUF1 (N349, N341);
xor XOR2 (N350, N324, N216);
nand NAND3 (N351, N350, N42, N338);
not NOT1 (N352, N257);
and AND2 (N353, N351, N86);
nor NOR2 (N354, N342, N269);
or OR2 (N355, N352, N351);
or OR3 (N356, N347, N19, N127);
or OR4 (N357, N353, N335, N340, N28);
not NOT1 (N358, N345);
xor XOR2 (N359, N358, N134);
nand NAND2 (N360, N355, N113);
or OR2 (N361, N337, N273);
buf BUF1 (N362, N360);
nand NAND2 (N363, N348, N100);
nand NAND3 (N364, N349, N198, N332);
buf BUF1 (N365, N44);
not NOT1 (N366, N362);
nand NAND2 (N367, N364, N37);
buf BUF1 (N368, N359);
nand NAND2 (N369, N365, N136);
buf BUF1 (N370, N361);
or OR3 (N371, N331, N319, N316);
nand NAND2 (N372, N357, N24);
buf BUF1 (N373, N356);
or OR4 (N374, N370, N342, N196, N101);
xor XOR2 (N375, N374, N170);
and AND2 (N376, N368, N204);
xor XOR2 (N377, N371, N16);
or OR3 (N378, N372, N171, N330);
not NOT1 (N379, N354);
nand NAND3 (N380, N376, N334, N9);
nor NOR3 (N381, N378, N100, N14);
nor NOR2 (N382, N363, N200);
and AND4 (N383, N382, N165, N219, N60);
and AND3 (N384, N379, N215, N55);
xor XOR2 (N385, N366, N188);
nand NAND3 (N386, N377, N298, N303);
buf BUF1 (N387, N375);
nor NOR4 (N388, N369, N77, N313, N172);
not NOT1 (N389, N384);
nor NOR3 (N390, N389, N352, N234);
or OR2 (N391, N381, N150);
or OR3 (N392, N391, N379, N334);
xor XOR2 (N393, N386, N358);
nand NAND4 (N394, N385, N71, N249, N63);
xor XOR2 (N395, N394, N203);
xor XOR2 (N396, N395, N291);
not NOT1 (N397, N383);
not NOT1 (N398, N380);
nor NOR3 (N399, N392, N398, N301);
xor XOR2 (N400, N212, N115);
xor XOR2 (N401, N400, N187);
and AND2 (N402, N399, N36);
nand NAND4 (N403, N367, N191, N101, N339);
nor NOR4 (N404, N390, N236, N248, N397);
or OR2 (N405, N193, N151);
and AND2 (N406, N404, N305);
not NOT1 (N407, N393);
not NOT1 (N408, N403);
and AND3 (N409, N406, N208, N110);
xor XOR2 (N410, N409, N393);
xor XOR2 (N411, N387, N354);
not NOT1 (N412, N373);
nor NOR2 (N413, N402, N102);
xor XOR2 (N414, N401, N82);
nor NOR4 (N415, N410, N237, N171, N142);
and AND4 (N416, N408, N382, N177, N231);
nand NAND4 (N417, N413, N273, N130, N359);
xor XOR2 (N418, N417, N247);
buf BUF1 (N419, N412);
xor XOR2 (N420, N396, N64);
and AND3 (N421, N419, N237, N275);
nor NOR3 (N422, N420, N358, N162);
xor XOR2 (N423, N421, N139);
xor XOR2 (N424, N411, N389);
not NOT1 (N425, N388);
or OR4 (N426, N423, N402, N50, N339);
nand NAND2 (N427, N415, N386);
nor NOR4 (N428, N416, N283, N17, N396);
nor NOR2 (N429, N405, N426);
nor NOR2 (N430, N254, N279);
or OR2 (N431, N427, N312);
xor XOR2 (N432, N414, N341);
not NOT1 (N433, N430);
or OR4 (N434, N407, N153, N20, N355);
buf BUF1 (N435, N422);
nor NOR4 (N436, N434, N287, N228, N25);
xor XOR2 (N437, N429, N179);
and AND4 (N438, N424, N409, N141, N95);
nand NAND3 (N439, N428, N178, N154);
and AND4 (N440, N433, N74, N407, N259);
or OR3 (N441, N432, N114, N229);
or OR3 (N442, N441, N421, N190);
nand NAND3 (N443, N438, N194, N185);
nor NOR3 (N444, N437, N439, N228);
xor XOR2 (N445, N280, N159);
buf BUF1 (N446, N431);
buf BUF1 (N447, N443);
not NOT1 (N448, N440);
not NOT1 (N449, N442);
nand NAND3 (N450, N444, N437, N300);
nand NAND2 (N451, N446, N449);
nand NAND3 (N452, N338, N149, N276);
or OR2 (N453, N445, N15);
or OR4 (N454, N418, N299, N331, N328);
or OR4 (N455, N452, N175, N224, N436);
or OR3 (N456, N81, N160, N407);
xor XOR2 (N457, N451, N98);
xor XOR2 (N458, N457, N78);
nand NAND2 (N459, N448, N18);
xor XOR2 (N460, N455, N34);
not NOT1 (N461, N456);
xor XOR2 (N462, N460, N393);
nor NOR3 (N463, N425, N379, N89);
nor NOR3 (N464, N454, N10, N395);
nor NOR2 (N465, N435, N315);
nand NAND4 (N466, N463, N373, N52, N114);
not NOT1 (N467, N459);
not NOT1 (N468, N464);
nor NOR4 (N469, N458, N216, N128, N420);
and AND4 (N470, N467, N422, N125, N86);
not NOT1 (N471, N470);
buf BUF1 (N472, N471);
xor XOR2 (N473, N469, N155);
nor NOR2 (N474, N453, N369);
or OR3 (N475, N473, N345, N323);
nand NAND2 (N476, N447, N244);
or OR3 (N477, N474, N357, N468);
or OR3 (N478, N459, N114, N305);
not NOT1 (N479, N478);
buf BUF1 (N480, N466);
or OR4 (N481, N472, N38, N454, N73);
or OR3 (N482, N475, N14, N68);
buf BUF1 (N483, N482);
nand NAND3 (N484, N476, N118, N142);
buf BUF1 (N485, N450);
not NOT1 (N486, N481);
xor XOR2 (N487, N461, N228);
and AND3 (N488, N477, N340, N374);
nand NAND3 (N489, N486, N261, N123);
or OR3 (N490, N485, N165, N145);
xor XOR2 (N491, N480, N420);
buf BUF1 (N492, N483);
nor NOR3 (N493, N487, N209, N292);
not NOT1 (N494, N492);
buf BUF1 (N495, N488);
buf BUF1 (N496, N465);
or OR3 (N497, N489, N8, N160);
and AND2 (N498, N462, N493);
xor XOR2 (N499, N309, N125);
xor XOR2 (N500, N496, N81);
nand NAND4 (N501, N497, N391, N284, N271);
or OR4 (N502, N498, N5, N113, N141);
nor NOR4 (N503, N499, N206, N60, N301);
buf BUF1 (N504, N501);
not NOT1 (N505, N503);
nor NOR4 (N506, N504, N453, N394, N382);
xor XOR2 (N507, N490, N494);
and AND2 (N508, N233, N74);
buf BUF1 (N509, N505);
or OR3 (N510, N502, N183, N372);
nor NOR4 (N511, N500, N301, N408, N127);
and AND3 (N512, N484, N263, N315);
or OR3 (N513, N512, N161, N246);
buf BUF1 (N514, N491);
nor NOR2 (N515, N508, N5);
not NOT1 (N516, N507);
or OR3 (N517, N506, N33, N461);
xor XOR2 (N518, N479, N392);
or OR3 (N519, N510, N325, N69);
or OR3 (N520, N519, N47, N378);
nand NAND2 (N521, N518, N408);
buf BUF1 (N522, N514);
nor NOR2 (N523, N522, N328);
nand NAND2 (N524, N516, N91);
not NOT1 (N525, N524);
or OR3 (N526, N515, N305, N208);
or OR2 (N527, N525, N156);
not NOT1 (N528, N495);
buf BUF1 (N529, N523);
or OR2 (N530, N520, N134);
xor XOR2 (N531, N517, N487);
buf BUF1 (N532, N521);
not NOT1 (N533, N513);
buf BUF1 (N534, N509);
nor NOR3 (N535, N534, N348, N187);
or OR4 (N536, N535, N187, N179, N11);
xor XOR2 (N537, N530, N196);
xor XOR2 (N538, N527, N47);
and AND4 (N539, N532, N332, N425, N356);
and AND3 (N540, N529, N522, N429);
and AND3 (N541, N537, N367, N146);
not NOT1 (N542, N511);
nand NAND3 (N543, N540, N273, N131);
nor NOR3 (N544, N542, N85, N187);
not NOT1 (N545, N541);
nor NOR2 (N546, N543, N177);
xor XOR2 (N547, N536, N59);
or OR3 (N548, N533, N98, N106);
or OR3 (N549, N531, N419, N472);
buf BUF1 (N550, N539);
nand NAND4 (N551, N546, N256, N411, N215);
or OR3 (N552, N538, N271, N465);
nor NOR4 (N553, N548, N383, N511, N462);
nor NOR3 (N554, N552, N460, N516);
and AND4 (N555, N547, N447, N443, N110);
xor XOR2 (N556, N528, N110);
and AND3 (N557, N553, N524, N37);
and AND2 (N558, N544, N388);
xor XOR2 (N559, N550, N474);
nand NAND3 (N560, N545, N512, N188);
nand NAND3 (N561, N526, N112, N114);
buf BUF1 (N562, N557);
buf BUF1 (N563, N555);
nor NOR3 (N564, N549, N236, N268);
buf BUF1 (N565, N564);
nor NOR2 (N566, N551, N358);
nor NOR3 (N567, N561, N559, N425);
xor XOR2 (N568, N181, N188);
xor XOR2 (N569, N556, N401);
or OR4 (N570, N569, N308, N187, N280);
buf BUF1 (N571, N570);
nor NOR3 (N572, N554, N260, N282);
nand NAND3 (N573, N566, N8, N359);
and AND3 (N574, N563, N419, N286);
xor XOR2 (N575, N562, N237);
not NOT1 (N576, N573);
and AND3 (N577, N558, N347, N293);
buf BUF1 (N578, N567);
nand NAND3 (N579, N575, N200, N530);
nor NOR3 (N580, N576, N457, N341);
not NOT1 (N581, N578);
nand NAND2 (N582, N579, N125);
xor XOR2 (N583, N568, N195);
buf BUF1 (N584, N560);
or OR2 (N585, N565, N419);
buf BUF1 (N586, N582);
nand NAND3 (N587, N572, N404, N389);
nor NOR3 (N588, N584, N240, N304);
nand NAND2 (N589, N580, N74);
not NOT1 (N590, N585);
or OR4 (N591, N590, N425, N246, N270);
or OR3 (N592, N574, N301, N478);
xor XOR2 (N593, N591, N223);
and AND3 (N594, N577, N452, N404);
and AND2 (N595, N583, N95);
xor XOR2 (N596, N586, N203);
buf BUF1 (N597, N595);
nand NAND4 (N598, N596, N262, N266, N355);
and AND3 (N599, N594, N589, N401);
not NOT1 (N600, N96);
buf BUF1 (N601, N600);
buf BUF1 (N602, N592);
and AND3 (N603, N588, N220, N518);
or OR2 (N604, N602, N37);
and AND3 (N605, N598, N217, N184);
not NOT1 (N606, N571);
not NOT1 (N607, N601);
nand NAND3 (N608, N606, N479, N388);
or OR3 (N609, N587, N252, N443);
nor NOR2 (N610, N608, N432);
or OR2 (N611, N593, N127);
and AND3 (N612, N611, N45, N321);
nor NOR3 (N613, N610, N292, N559);
xor XOR2 (N614, N599, N334);
xor XOR2 (N615, N603, N425);
buf BUF1 (N616, N581);
not NOT1 (N617, N613);
xor XOR2 (N618, N615, N183);
not NOT1 (N619, N617);
not NOT1 (N620, N607);
nor NOR3 (N621, N605, N106, N146);
buf BUF1 (N622, N597);
or OR3 (N623, N620, N430, N537);
nor NOR2 (N624, N623, N278);
and AND3 (N625, N616, N448, N85);
or OR3 (N626, N625, N445, N362);
or OR2 (N627, N609, N601);
and AND4 (N628, N627, N250, N140, N243);
xor XOR2 (N629, N618, N461);
buf BUF1 (N630, N619);
nor NOR2 (N631, N612, N114);
and AND2 (N632, N628, N283);
not NOT1 (N633, N621);
not NOT1 (N634, N630);
and AND3 (N635, N622, N476, N130);
and AND4 (N636, N629, N75, N172, N361);
xor XOR2 (N637, N633, N303);
not NOT1 (N638, N614);
not NOT1 (N639, N632);
xor XOR2 (N640, N638, N531);
and AND2 (N641, N635, N473);
or OR3 (N642, N639, N59, N494);
nand NAND3 (N643, N624, N174, N574);
xor XOR2 (N644, N636, N169);
and AND3 (N645, N641, N518, N623);
and AND4 (N646, N644, N221, N374, N61);
and AND3 (N647, N634, N91, N599);
or OR3 (N648, N626, N242, N424);
and AND2 (N649, N643, N502);
not NOT1 (N650, N631);
not NOT1 (N651, N649);
buf BUF1 (N652, N640);
xor XOR2 (N653, N650, N79);
nand NAND3 (N654, N642, N611, N652);
buf BUF1 (N655, N382);
nand NAND3 (N656, N653, N578, N339);
nor NOR4 (N657, N647, N277, N476, N462);
nor NOR2 (N658, N651, N325);
nor NOR3 (N659, N655, N500, N104);
not NOT1 (N660, N645);
or OR2 (N661, N654, N405);
or OR3 (N662, N658, N628, N628);
and AND4 (N663, N660, N21, N513, N362);
buf BUF1 (N664, N648);
xor XOR2 (N665, N646, N252);
buf BUF1 (N666, N637);
nor NOR4 (N667, N656, N554, N300, N76);
and AND3 (N668, N661, N226, N615);
and AND3 (N669, N668, N430, N222);
nor NOR3 (N670, N666, N34, N241);
buf BUF1 (N671, N657);
nor NOR4 (N672, N604, N494, N141, N296);
not NOT1 (N673, N672);
or OR3 (N674, N663, N254, N244);
nand NAND4 (N675, N673, N230, N299, N53);
and AND4 (N676, N669, N638, N372, N488);
not NOT1 (N677, N665);
xor XOR2 (N678, N676, N413);
nand NAND4 (N679, N671, N543, N177, N38);
nor NOR4 (N680, N667, N494, N230, N544);
xor XOR2 (N681, N664, N94);
buf BUF1 (N682, N677);
nand NAND4 (N683, N679, N232, N170, N100);
buf BUF1 (N684, N659);
xor XOR2 (N685, N678, N211);
and AND2 (N686, N684, N232);
and AND2 (N687, N675, N431);
nor NOR2 (N688, N680, N415);
not NOT1 (N689, N670);
or OR3 (N690, N689, N139, N562);
and AND2 (N691, N682, N525);
nor NOR2 (N692, N674, N564);
not NOT1 (N693, N690);
or OR4 (N694, N687, N504, N128, N189);
and AND2 (N695, N688, N303);
not NOT1 (N696, N692);
xor XOR2 (N697, N691, N441);
buf BUF1 (N698, N683);
xor XOR2 (N699, N698, N449);
buf BUF1 (N700, N685);
nand NAND2 (N701, N696, N143);
or OR3 (N702, N700, N219, N445);
and AND4 (N703, N681, N357, N395, N83);
nor NOR3 (N704, N695, N291, N529);
or OR3 (N705, N662, N1, N569);
not NOT1 (N706, N693);
nand NAND4 (N707, N702, N172, N253, N559);
nor NOR2 (N708, N697, N408);
nand NAND4 (N709, N686, N35, N552, N692);
and AND4 (N710, N699, N310, N32, N514);
or OR2 (N711, N703, N95);
nand NAND4 (N712, N710, N561, N350, N332);
and AND4 (N713, N705, N153, N424, N82);
xor XOR2 (N714, N709, N258);
or OR2 (N715, N711, N385);
nor NOR4 (N716, N708, N627, N508, N627);
xor XOR2 (N717, N707, N693);
buf BUF1 (N718, N712);
nor NOR3 (N719, N717, N415, N293);
buf BUF1 (N720, N719);
xor XOR2 (N721, N716, N575);
or OR3 (N722, N694, N32, N569);
nor NOR2 (N723, N714, N305);
nor NOR3 (N724, N723, N2, N64);
or OR2 (N725, N720, N511);
nor NOR2 (N726, N706, N205);
nand NAND4 (N727, N715, N385, N337, N484);
or OR3 (N728, N725, N292, N252);
buf BUF1 (N729, N718);
and AND2 (N730, N727, N342);
xor XOR2 (N731, N730, N593);
not NOT1 (N732, N722);
nand NAND4 (N733, N713, N102, N552, N728);
buf BUF1 (N734, N579);
not NOT1 (N735, N724);
not NOT1 (N736, N726);
not NOT1 (N737, N704);
nand NAND3 (N738, N733, N524, N491);
and AND4 (N739, N736, N538, N715, N496);
and AND2 (N740, N729, N56);
nor NOR2 (N741, N739, N350);
and AND2 (N742, N701, N276);
nand NAND4 (N743, N740, N463, N419, N370);
nor NOR4 (N744, N742, N528, N34, N447);
or OR2 (N745, N734, N551);
nor NOR3 (N746, N745, N386, N297);
buf BUF1 (N747, N721);
nor NOR3 (N748, N732, N542, N546);
nor NOR3 (N749, N744, N514, N646);
buf BUF1 (N750, N743);
xor XOR2 (N751, N737, N237);
nor NOR3 (N752, N748, N500, N561);
xor XOR2 (N753, N749, N644);
or OR2 (N754, N751, N491);
not NOT1 (N755, N752);
buf BUF1 (N756, N755);
nand NAND4 (N757, N731, N707, N365, N697);
nand NAND3 (N758, N750, N605, N533);
nor NOR4 (N759, N757, N21, N259, N72);
nor NOR2 (N760, N753, N406);
nor NOR4 (N761, N754, N390, N506, N416);
xor XOR2 (N762, N759, N700);
not NOT1 (N763, N741);
xor XOR2 (N764, N756, N454);
nor NOR2 (N765, N760, N315);
and AND4 (N766, N762, N12, N193, N203);
nor NOR4 (N767, N747, N313, N468, N144);
and AND2 (N768, N765, N63);
nand NAND3 (N769, N767, N623, N224);
buf BUF1 (N770, N758);
nor NOR3 (N771, N769, N106, N149);
buf BUF1 (N772, N764);
nor NOR3 (N773, N772, N389, N422);
buf BUF1 (N774, N770);
and AND4 (N775, N738, N142, N611, N267);
and AND4 (N776, N773, N544, N661, N510);
or OR2 (N777, N735, N687);
buf BUF1 (N778, N775);
or OR3 (N779, N761, N767, N716);
not NOT1 (N780, N776);
or OR2 (N781, N771, N761);
buf BUF1 (N782, N777);
nand NAND4 (N783, N779, N137, N50, N54);
nand NAND4 (N784, N782, N118, N559, N575);
and AND4 (N785, N780, N424, N450, N605);
or OR4 (N786, N778, N663, N141, N203);
or OR3 (N787, N763, N570, N79);
not NOT1 (N788, N784);
not NOT1 (N789, N768);
xor XOR2 (N790, N781, N235);
or OR4 (N791, N746, N187, N757, N623);
nand NAND4 (N792, N774, N719, N186, N514);
or OR4 (N793, N786, N500, N248, N506);
nor NOR4 (N794, N791, N305, N344, N114);
nor NOR4 (N795, N792, N313, N650, N125);
buf BUF1 (N796, N794);
nor NOR3 (N797, N783, N229, N362);
and AND4 (N798, N790, N646, N222, N177);
and AND3 (N799, N797, N48, N458);
or OR3 (N800, N788, N516, N386);
nand NAND3 (N801, N795, N117, N260);
or OR2 (N802, N766, N206);
and AND3 (N803, N802, N587, N784);
nand NAND2 (N804, N785, N600);
buf BUF1 (N805, N801);
xor XOR2 (N806, N799, N498);
nand NAND4 (N807, N796, N478, N12, N790);
buf BUF1 (N808, N800);
not NOT1 (N809, N808);
or OR3 (N810, N793, N607, N787);
nor NOR2 (N811, N293, N410);
not NOT1 (N812, N810);
buf BUF1 (N813, N798);
not NOT1 (N814, N789);
nor NOR3 (N815, N811, N760, N396);
or OR3 (N816, N809, N252, N374);
and AND2 (N817, N814, N89);
nand NAND2 (N818, N817, N191);
nand NAND4 (N819, N806, N371, N567, N606);
nor NOR3 (N820, N812, N89, N207);
not NOT1 (N821, N807);
buf BUF1 (N822, N805);
not NOT1 (N823, N822);
xor XOR2 (N824, N819, N371);
or OR3 (N825, N813, N673, N4);
nand NAND2 (N826, N803, N615);
nor NOR3 (N827, N825, N520, N23);
nand NAND3 (N828, N815, N353, N605);
nand NAND3 (N829, N804, N618, N226);
buf BUF1 (N830, N816);
not NOT1 (N831, N818);
or OR3 (N832, N829, N631, N268);
not NOT1 (N833, N830);
not NOT1 (N834, N832);
or OR2 (N835, N827, N380);
xor XOR2 (N836, N821, N84);
or OR3 (N837, N828, N143, N102);
nand NAND4 (N838, N823, N64, N803, N364);
nand NAND4 (N839, N833, N209, N285, N196);
or OR2 (N840, N839, N789);
xor XOR2 (N841, N831, N341);
nand NAND3 (N842, N837, N403, N202);
and AND4 (N843, N826, N813, N523, N493);
not NOT1 (N844, N842);
nor NOR2 (N845, N844, N82);
xor XOR2 (N846, N845, N637);
not NOT1 (N847, N841);
nor NOR3 (N848, N838, N660, N718);
nor NOR4 (N849, N848, N280, N455, N802);
and AND4 (N850, N846, N546, N769, N500);
or OR4 (N851, N835, N264, N85, N555);
xor XOR2 (N852, N849, N107);
xor XOR2 (N853, N834, N380);
nand NAND3 (N854, N850, N411, N541);
xor XOR2 (N855, N840, N819);
xor XOR2 (N856, N824, N426);
or OR3 (N857, N843, N250, N458);
or OR2 (N858, N854, N270);
not NOT1 (N859, N853);
or OR2 (N860, N820, N47);
or OR2 (N861, N857, N795);
and AND4 (N862, N858, N590, N194, N235);
or OR2 (N863, N859, N68);
nor NOR3 (N864, N855, N310, N489);
nand NAND4 (N865, N864, N227, N780, N547);
not NOT1 (N866, N862);
nor NOR2 (N867, N836, N807);
nor NOR2 (N868, N847, N78);
nand NAND3 (N869, N856, N438, N172);
nand NAND4 (N870, N852, N245, N43, N89);
nand NAND3 (N871, N870, N187, N755);
nand NAND4 (N872, N865, N735, N412, N543);
and AND4 (N873, N866, N345, N466, N862);
nor NOR4 (N874, N871, N790, N370, N475);
buf BUF1 (N875, N872);
xor XOR2 (N876, N875, N511);
not NOT1 (N877, N851);
nor NOR2 (N878, N868, N440);
nand NAND4 (N879, N863, N654, N645, N620);
nor NOR2 (N880, N867, N262);
or OR3 (N881, N874, N372, N107);
nand NAND3 (N882, N873, N529, N569);
or OR3 (N883, N869, N776, N447);
or OR2 (N884, N881, N135);
nor NOR2 (N885, N883, N698);
and AND3 (N886, N876, N7, N813);
not NOT1 (N887, N884);
or OR2 (N888, N885, N495);
xor XOR2 (N889, N878, N27);
xor XOR2 (N890, N877, N594);
nor NOR3 (N891, N890, N239, N169);
not NOT1 (N892, N861);
nor NOR3 (N893, N879, N328, N854);
nand NAND4 (N894, N888, N531, N715, N174);
not NOT1 (N895, N882);
nand NAND3 (N896, N886, N406, N22);
or OR2 (N897, N894, N699);
buf BUF1 (N898, N860);
or OR2 (N899, N898, N310);
buf BUF1 (N900, N887);
nand NAND2 (N901, N899, N694);
nor NOR4 (N902, N896, N45, N295, N396);
or OR2 (N903, N880, N389);
xor XOR2 (N904, N902, N752);
nor NOR3 (N905, N889, N671, N231);
and AND4 (N906, N901, N483, N53, N848);
not NOT1 (N907, N903);
buf BUF1 (N908, N892);
and AND3 (N909, N908, N236, N796);
or OR2 (N910, N907, N131);
not NOT1 (N911, N900);
nand NAND4 (N912, N893, N779, N896, N825);
buf BUF1 (N913, N909);
xor XOR2 (N914, N895, N507);
not NOT1 (N915, N914);
not NOT1 (N916, N891);
and AND4 (N917, N915, N806, N536, N896);
nor NOR2 (N918, N910, N613);
buf BUF1 (N919, N906);
not NOT1 (N920, N916);
and AND4 (N921, N905, N19, N891, N896);
nand NAND4 (N922, N920, N526, N442, N190);
and AND3 (N923, N912, N909, N148);
endmodule