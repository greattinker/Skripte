// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12;

output N1511,N1504,N1505,N1491,N1508,N1484,N1486,N1502,N1510,N1512;

nand NAND3 (N13, N1, N9, N7);
not NOT1 (N14, N7);
nor NOR3 (N15, N5, N14, N2);
buf BUF1 (N16, N14);
and AND4 (N17, N14, N2, N4, N8);
nor NOR3 (N18, N15, N9, N7);
not NOT1 (N19, N2);
not NOT1 (N20, N7);
nor NOR4 (N21, N15, N13, N1, N1);
and AND4 (N22, N16, N7, N4, N9);
nand NAND2 (N23, N21, N14);
xor XOR2 (N24, N20, N9);
not NOT1 (N25, N14);
not NOT1 (N26, N25);
xor XOR2 (N27, N21, N10);
and AND2 (N28, N6, N15);
and AND4 (N29, N27, N21, N23, N26);
nand NAND3 (N30, N6, N25, N25);
not NOT1 (N31, N22);
buf BUF1 (N32, N17);
not NOT1 (N33, N21);
or OR4 (N34, N4, N1, N10, N14);
not NOT1 (N35, N24);
and AND4 (N36, N32, N34, N10, N24);
or OR3 (N37, N26, N22, N17);
or OR4 (N38, N18, N18, N22, N18);
not NOT1 (N39, N35);
and AND4 (N40, N28, N30, N28, N2);
nor NOR3 (N41, N14, N35, N34);
nand NAND4 (N42, N19, N19, N41, N16);
buf BUF1 (N43, N39);
not NOT1 (N44, N43);
not NOT1 (N45, N9);
xor XOR2 (N46, N31, N12);
and AND2 (N47, N36, N2);
not NOT1 (N48, N38);
buf BUF1 (N49, N33);
not NOT1 (N50, N44);
nor NOR3 (N51, N46, N46, N20);
not NOT1 (N52, N48);
xor XOR2 (N53, N45, N13);
and AND3 (N54, N49, N38, N32);
nand NAND3 (N55, N40, N32, N39);
buf BUF1 (N56, N29);
xor XOR2 (N57, N54, N52);
nand NAND4 (N58, N33, N4, N9, N35);
or OR3 (N59, N42, N29, N52);
not NOT1 (N60, N51);
nor NOR2 (N61, N53, N35);
buf BUF1 (N62, N56);
or OR2 (N63, N50, N33);
not NOT1 (N64, N55);
xor XOR2 (N65, N60, N6);
and AND4 (N66, N58, N23, N47, N52);
buf BUF1 (N67, N36);
or OR4 (N68, N57, N12, N17, N26);
nand NAND3 (N69, N62, N50, N23);
buf BUF1 (N70, N64);
xor XOR2 (N71, N69, N46);
buf BUF1 (N72, N63);
not NOT1 (N73, N70);
or OR3 (N74, N65, N11, N35);
or OR4 (N75, N59, N26, N6, N55);
nand NAND2 (N76, N61, N22);
or OR4 (N77, N37, N30, N69, N28);
nand NAND3 (N78, N74, N76, N32);
and AND2 (N79, N37, N5);
nor NOR2 (N80, N67, N37);
buf BUF1 (N81, N66);
or OR2 (N82, N73, N70);
and AND4 (N83, N77, N63, N64, N58);
nand NAND4 (N84, N79, N55, N83, N18);
nand NAND4 (N85, N14, N41, N52, N59);
and AND4 (N86, N75, N62, N31, N26);
buf BUF1 (N87, N85);
or OR2 (N88, N72, N42);
not NOT1 (N89, N78);
buf BUF1 (N90, N68);
and AND2 (N91, N84, N20);
buf BUF1 (N92, N71);
xor XOR2 (N93, N89, N38);
xor XOR2 (N94, N86, N31);
and AND4 (N95, N92, N29, N27, N4);
nand NAND3 (N96, N91, N51, N74);
not NOT1 (N97, N82);
and AND4 (N98, N97, N63, N27, N75);
xor XOR2 (N99, N93, N96);
buf BUF1 (N100, N48);
buf BUF1 (N101, N99);
buf BUF1 (N102, N90);
nor NOR2 (N103, N100, N48);
nand NAND3 (N104, N95, N90, N55);
buf BUF1 (N105, N102);
nand NAND2 (N106, N105, N59);
nand NAND4 (N107, N88, N51, N91, N81);
nand NAND2 (N108, N38, N81);
or OR2 (N109, N104, N29);
or OR2 (N110, N101, N31);
nand NAND2 (N111, N109, N94);
and AND3 (N112, N108, N35, N34);
buf BUF1 (N113, N20);
nand NAND3 (N114, N106, N70, N13);
or OR4 (N115, N110, N69, N8, N57);
xor XOR2 (N116, N80, N27);
not NOT1 (N117, N107);
not NOT1 (N118, N114);
buf BUF1 (N119, N116);
or OR2 (N120, N119, N47);
and AND3 (N121, N111, N4, N30);
nor NOR4 (N122, N120, N50, N21, N112);
buf BUF1 (N123, N45);
xor XOR2 (N124, N121, N68);
buf BUF1 (N125, N103);
nor NOR4 (N126, N113, N79, N32, N50);
not NOT1 (N127, N98);
not NOT1 (N128, N125);
and AND2 (N129, N117, N124);
or OR4 (N130, N119, N122, N40, N24);
not NOT1 (N131, N36);
nand NAND4 (N132, N126, N99, N48, N79);
and AND4 (N133, N87, N24, N71, N112);
not NOT1 (N134, N128);
or OR2 (N135, N131, N72);
xor XOR2 (N136, N129, N117);
nand NAND3 (N137, N130, N82, N127);
xor XOR2 (N138, N117, N66);
buf BUF1 (N139, N138);
or OR4 (N140, N139, N11, N98, N21);
not NOT1 (N141, N132);
and AND4 (N142, N115, N88, N6, N37);
or OR4 (N143, N140, N3, N38, N97);
and AND4 (N144, N118, N141, N83, N32);
not NOT1 (N145, N52);
nor NOR3 (N146, N136, N50, N138);
nand NAND3 (N147, N133, N10, N75);
and AND2 (N148, N147, N41);
xor XOR2 (N149, N142, N119);
nor NOR2 (N150, N137, N1);
or OR3 (N151, N135, N133, N65);
nand NAND2 (N152, N148, N34);
xor XOR2 (N153, N151, N23);
and AND3 (N154, N152, N88, N68);
not NOT1 (N155, N123);
buf BUF1 (N156, N154);
and AND2 (N157, N149, N87);
or OR2 (N158, N134, N45);
nor NOR4 (N159, N153, N126, N28, N102);
nor NOR3 (N160, N146, N89, N102);
nor NOR4 (N161, N156, N46, N157, N156);
nand NAND3 (N162, N56, N141, N79);
not NOT1 (N163, N143);
xor XOR2 (N164, N155, N12);
nor NOR4 (N165, N160, N144, N69, N134);
or OR3 (N166, N91, N8, N46);
xor XOR2 (N167, N162, N59);
buf BUF1 (N168, N159);
and AND2 (N169, N158, N129);
not NOT1 (N170, N165);
or OR2 (N171, N145, N26);
and AND2 (N172, N171, N97);
buf BUF1 (N173, N167);
buf BUF1 (N174, N164);
nand NAND2 (N175, N170, N22);
not NOT1 (N176, N161);
nand NAND2 (N177, N174, N106);
or OR3 (N178, N150, N151, N132);
xor XOR2 (N179, N172, N74);
nor NOR4 (N180, N168, N15, N153, N131);
or OR4 (N181, N179, N61, N75, N100);
buf BUF1 (N182, N178);
not NOT1 (N183, N173);
nor NOR2 (N184, N181, N87);
buf BUF1 (N185, N184);
or OR4 (N186, N163, N51, N16, N145);
nand NAND4 (N187, N186, N118, N98, N138);
nand NAND3 (N188, N182, N34, N35);
not NOT1 (N189, N187);
buf BUF1 (N190, N169);
buf BUF1 (N191, N180);
or OR3 (N192, N190, N151, N43);
buf BUF1 (N193, N166);
not NOT1 (N194, N183);
or OR3 (N195, N176, N48, N171);
xor XOR2 (N196, N193, N19);
and AND3 (N197, N185, N67, N72);
or OR3 (N198, N196, N146, N136);
or OR4 (N199, N175, N9, N177, N143);
xor XOR2 (N200, N146, N109);
nor NOR4 (N201, N200, N47, N155, N187);
or OR3 (N202, N191, N48, N135);
or OR2 (N203, N198, N11);
or OR3 (N204, N201, N200, N9);
nand NAND3 (N205, N203, N101, N160);
and AND3 (N206, N205, N105, N153);
or OR2 (N207, N188, N177);
xor XOR2 (N208, N195, N52);
or OR2 (N209, N208, N167);
xor XOR2 (N210, N204, N88);
nand NAND4 (N211, N194, N83, N176, N181);
xor XOR2 (N212, N207, N70);
not NOT1 (N213, N202);
nand NAND3 (N214, N192, N177, N191);
or OR3 (N215, N209, N128, N196);
or OR3 (N216, N199, N154, N23);
buf BUF1 (N217, N213);
not NOT1 (N218, N189);
and AND2 (N219, N215, N20);
and AND4 (N220, N197, N180, N30, N26);
or OR4 (N221, N218, N136, N53, N39);
buf BUF1 (N222, N211);
and AND3 (N223, N206, N176, N99);
nand NAND3 (N224, N216, N202, N190);
or OR2 (N225, N220, N148);
and AND2 (N226, N210, N212);
or OR2 (N227, N52, N132);
nor NOR2 (N228, N226, N89);
nor NOR3 (N229, N225, N147, N70);
buf BUF1 (N230, N214);
nor NOR3 (N231, N224, N44, N170);
and AND2 (N232, N231, N125);
not NOT1 (N233, N228);
nand NAND4 (N234, N222, N221, N220, N97);
nor NOR2 (N235, N19, N28);
nor NOR2 (N236, N227, N172);
or OR3 (N237, N235, N58, N229);
not NOT1 (N238, N231);
nand NAND2 (N239, N238, N59);
and AND3 (N240, N219, N87, N19);
buf BUF1 (N241, N232);
or OR2 (N242, N234, N241);
or OR3 (N243, N238, N90, N82);
xor XOR2 (N244, N239, N8);
nor NOR3 (N245, N242, N214, N211);
and AND4 (N246, N240, N31, N90, N164);
nor NOR3 (N247, N217, N108, N26);
buf BUF1 (N248, N230);
buf BUF1 (N249, N237);
or OR2 (N250, N247, N145);
nor NOR3 (N251, N233, N210, N150);
buf BUF1 (N252, N249);
nor NOR3 (N253, N245, N29, N54);
not NOT1 (N254, N252);
not NOT1 (N255, N254);
nand NAND2 (N256, N223, N197);
not NOT1 (N257, N251);
buf BUF1 (N258, N248);
nand NAND4 (N259, N246, N204, N164, N196);
or OR4 (N260, N257, N132, N114, N146);
and AND4 (N261, N260, N241, N137, N215);
or OR3 (N262, N256, N182, N226);
xor XOR2 (N263, N236, N122);
xor XOR2 (N264, N261, N146);
nand NAND2 (N265, N255, N25);
not NOT1 (N266, N263);
not NOT1 (N267, N244);
xor XOR2 (N268, N266, N174);
not NOT1 (N269, N259);
buf BUF1 (N270, N264);
not NOT1 (N271, N265);
and AND3 (N272, N267, N98, N182);
nor NOR4 (N273, N268, N150, N63, N125);
nand NAND2 (N274, N253, N86);
nor NOR3 (N275, N269, N5, N270);
buf BUF1 (N276, N157);
not NOT1 (N277, N271);
or OR3 (N278, N273, N176, N151);
and AND3 (N279, N277, N198, N278);
nand NAND2 (N280, N234, N17);
buf BUF1 (N281, N250);
and AND2 (N282, N262, N195);
xor XOR2 (N283, N274, N32);
nand NAND3 (N284, N258, N21, N75);
or OR2 (N285, N276, N57);
nand NAND3 (N286, N283, N190, N199);
or OR3 (N287, N243, N32, N204);
buf BUF1 (N288, N284);
xor XOR2 (N289, N279, N251);
xor XOR2 (N290, N282, N213);
and AND4 (N291, N272, N246, N57, N59);
nor NOR2 (N292, N290, N144);
not NOT1 (N293, N286);
nand NAND4 (N294, N280, N26, N189, N168);
nor NOR2 (N295, N292, N167);
not NOT1 (N296, N288);
xor XOR2 (N297, N287, N31);
not NOT1 (N298, N289);
and AND2 (N299, N281, N46);
not NOT1 (N300, N299);
buf BUF1 (N301, N295);
xor XOR2 (N302, N294, N43);
not NOT1 (N303, N296);
buf BUF1 (N304, N275);
or OR4 (N305, N298, N152, N201, N14);
buf BUF1 (N306, N300);
nand NAND2 (N307, N306, N43);
xor XOR2 (N308, N291, N275);
not NOT1 (N309, N304);
nand NAND2 (N310, N301, N28);
buf BUF1 (N311, N303);
buf BUF1 (N312, N285);
buf BUF1 (N313, N297);
not NOT1 (N314, N293);
buf BUF1 (N315, N305);
not NOT1 (N316, N315);
buf BUF1 (N317, N313);
not NOT1 (N318, N311);
not NOT1 (N319, N308);
xor XOR2 (N320, N314, N233);
and AND3 (N321, N312, N276, N151);
nand NAND3 (N322, N309, N308, N6);
not NOT1 (N323, N302);
not NOT1 (N324, N319);
and AND2 (N325, N318, N242);
not NOT1 (N326, N317);
nor NOR4 (N327, N321, N107, N307, N168);
not NOT1 (N328, N41);
and AND3 (N329, N324, N206, N119);
or OR4 (N330, N310, N304, N12, N55);
nand NAND2 (N331, N322, N191);
nand NAND3 (N332, N323, N94, N162);
nor NOR3 (N333, N325, N196, N264);
not NOT1 (N334, N316);
buf BUF1 (N335, N330);
buf BUF1 (N336, N329);
nor NOR3 (N337, N335, N223, N138);
or OR2 (N338, N332, N240);
nor NOR4 (N339, N320, N95, N315, N130);
and AND2 (N340, N328, N141);
nor NOR4 (N341, N331, N46, N262, N149);
not NOT1 (N342, N340);
or OR4 (N343, N336, N208, N103, N274);
or OR3 (N344, N334, N184, N338);
buf BUF1 (N345, N311);
and AND3 (N346, N327, N134, N2);
nor NOR2 (N347, N346, N94);
or OR3 (N348, N343, N64, N315);
xor XOR2 (N349, N347, N99);
not NOT1 (N350, N342);
not NOT1 (N351, N337);
xor XOR2 (N352, N341, N12);
buf BUF1 (N353, N349);
not NOT1 (N354, N351);
buf BUF1 (N355, N352);
xor XOR2 (N356, N339, N109);
not NOT1 (N357, N356);
or OR2 (N358, N326, N168);
xor XOR2 (N359, N358, N122);
nand NAND2 (N360, N344, N107);
or OR4 (N361, N345, N218, N247, N235);
and AND4 (N362, N353, N31, N143, N268);
nand NAND4 (N363, N362, N180, N176, N179);
and AND3 (N364, N361, N52, N276);
xor XOR2 (N365, N363, N292);
buf BUF1 (N366, N350);
xor XOR2 (N367, N348, N351);
nand NAND4 (N368, N333, N278, N357, N127);
or OR4 (N369, N127, N96, N278, N248);
xor XOR2 (N370, N359, N364);
nand NAND2 (N371, N178, N68);
or OR4 (N372, N369, N250, N260, N131);
nand NAND4 (N373, N372, N80, N228, N123);
and AND2 (N374, N373, N269);
not NOT1 (N375, N368);
buf BUF1 (N376, N375);
and AND2 (N377, N365, N1);
and AND2 (N378, N371, N31);
not NOT1 (N379, N360);
nor NOR2 (N380, N374, N42);
and AND3 (N381, N380, N104, N114);
xor XOR2 (N382, N376, N34);
and AND3 (N383, N377, N171, N194);
or OR4 (N384, N355, N311, N356, N154);
or OR2 (N385, N383, N120);
nand NAND2 (N386, N382, N380);
not NOT1 (N387, N367);
and AND4 (N388, N366, N88, N105, N287);
not NOT1 (N389, N388);
nor NOR2 (N390, N354, N211);
and AND3 (N391, N389, N18, N222);
or OR4 (N392, N370, N334, N187, N120);
or OR3 (N393, N386, N350, N112);
xor XOR2 (N394, N379, N356);
nor NOR4 (N395, N381, N360, N9, N205);
and AND4 (N396, N390, N166, N101, N157);
not NOT1 (N397, N384);
or OR3 (N398, N378, N343, N134);
buf BUF1 (N399, N395);
nor NOR3 (N400, N391, N288, N28);
xor XOR2 (N401, N393, N7);
nand NAND3 (N402, N387, N82, N129);
buf BUF1 (N403, N385);
buf BUF1 (N404, N401);
or OR2 (N405, N403, N370);
nor NOR4 (N406, N405, N330, N372, N292);
buf BUF1 (N407, N399);
nand NAND2 (N408, N398, N342);
buf BUF1 (N409, N406);
and AND2 (N410, N394, N10);
nor NOR2 (N411, N402, N40);
or OR2 (N412, N407, N301);
or OR3 (N413, N392, N340, N186);
nand NAND3 (N414, N396, N354, N121);
buf BUF1 (N415, N410);
or OR2 (N416, N400, N279);
xor XOR2 (N417, N411, N360);
buf BUF1 (N418, N417);
xor XOR2 (N419, N408, N149);
not NOT1 (N420, N418);
not NOT1 (N421, N412);
buf BUF1 (N422, N414);
nor NOR3 (N423, N413, N243, N75);
nor NOR3 (N424, N415, N60, N379);
xor XOR2 (N425, N397, N348);
or OR3 (N426, N423, N362, N250);
nand NAND3 (N427, N420, N277, N37);
nand NAND4 (N428, N404, N427, N90, N268);
buf BUF1 (N429, N352);
not NOT1 (N430, N419);
and AND3 (N431, N425, N362, N312);
xor XOR2 (N432, N426, N170);
and AND3 (N433, N430, N253, N319);
nor NOR3 (N434, N424, N196, N207);
xor XOR2 (N435, N421, N398);
not NOT1 (N436, N429);
buf BUF1 (N437, N435);
nor NOR2 (N438, N436, N415);
buf BUF1 (N439, N431);
xor XOR2 (N440, N434, N326);
and AND3 (N441, N438, N417, N8);
nor NOR3 (N442, N409, N240, N37);
buf BUF1 (N443, N441);
not NOT1 (N444, N428);
or OR4 (N445, N416, N221, N210, N126);
buf BUF1 (N446, N443);
and AND4 (N447, N432, N341, N79, N186);
not NOT1 (N448, N433);
nand NAND3 (N449, N422, N298, N422);
or OR2 (N450, N448, N286);
nor NOR2 (N451, N447, N376);
buf BUF1 (N452, N444);
nor NOR3 (N453, N439, N219, N297);
nor NOR2 (N454, N453, N374);
or OR2 (N455, N451, N143);
xor XOR2 (N456, N442, N39);
not NOT1 (N457, N440);
not NOT1 (N458, N457);
buf BUF1 (N459, N455);
nor NOR4 (N460, N452, N438, N124, N396);
or OR4 (N461, N454, N211, N388, N72);
and AND3 (N462, N445, N5, N244);
buf BUF1 (N463, N450);
nor NOR3 (N464, N463, N341, N58);
or OR2 (N465, N459, N133);
and AND3 (N466, N461, N219, N171);
and AND4 (N467, N466, N422, N388, N375);
buf BUF1 (N468, N465);
nor NOR4 (N469, N467, N122, N116, N194);
nor NOR3 (N470, N460, N137, N161);
xor XOR2 (N471, N468, N201);
xor XOR2 (N472, N462, N80);
not NOT1 (N473, N471);
nand NAND4 (N474, N464, N296, N90, N72);
not NOT1 (N475, N446);
nor NOR2 (N476, N458, N271);
xor XOR2 (N477, N476, N239);
or OR2 (N478, N469, N189);
and AND3 (N479, N472, N432, N97);
not NOT1 (N480, N449);
xor XOR2 (N481, N480, N376);
and AND4 (N482, N474, N88, N195, N27);
and AND4 (N483, N470, N280, N176, N250);
nor NOR3 (N484, N479, N159, N419);
and AND2 (N485, N484, N301);
not NOT1 (N486, N477);
or OR2 (N487, N483, N472);
and AND2 (N488, N473, N438);
and AND3 (N489, N456, N416, N13);
and AND2 (N490, N486, N142);
nor NOR3 (N491, N478, N485, N32);
or OR3 (N492, N408, N62, N477);
nor NOR4 (N493, N492, N400, N256, N394);
nor NOR2 (N494, N487, N41);
xor XOR2 (N495, N493, N141);
nand NAND4 (N496, N475, N122, N480, N301);
nor NOR2 (N497, N482, N325);
xor XOR2 (N498, N495, N130);
and AND3 (N499, N481, N79, N192);
and AND3 (N500, N494, N357, N134);
or OR4 (N501, N489, N292, N76, N3);
nor NOR4 (N502, N500, N117, N257, N469);
xor XOR2 (N503, N491, N346);
not NOT1 (N504, N488);
buf BUF1 (N505, N502);
xor XOR2 (N506, N499, N15);
nor NOR4 (N507, N490, N151, N195, N278);
nor NOR2 (N508, N496, N237);
nand NAND2 (N509, N506, N40);
nand NAND3 (N510, N508, N332, N395);
and AND3 (N511, N505, N339, N389);
and AND2 (N512, N509, N139);
nand NAND2 (N513, N510, N241);
nand NAND4 (N514, N498, N399, N161, N148);
nand NAND2 (N515, N512, N431);
nand NAND2 (N516, N511, N330);
nand NAND2 (N517, N504, N339);
or OR2 (N518, N497, N265);
not NOT1 (N519, N513);
or OR4 (N520, N515, N48, N253, N430);
buf BUF1 (N521, N519);
or OR2 (N522, N501, N176);
xor XOR2 (N523, N522, N152);
and AND3 (N524, N437, N245, N331);
nand NAND4 (N525, N507, N250, N85, N259);
xor XOR2 (N526, N521, N490);
xor XOR2 (N527, N523, N20);
or OR4 (N528, N527, N67, N510, N161);
not NOT1 (N529, N516);
buf BUF1 (N530, N518);
or OR2 (N531, N520, N382);
nand NAND3 (N532, N524, N123, N374);
buf BUF1 (N533, N514);
nor NOR3 (N534, N525, N132, N488);
buf BUF1 (N535, N526);
nor NOR4 (N536, N517, N412, N71, N426);
not NOT1 (N537, N534);
buf BUF1 (N538, N531);
xor XOR2 (N539, N537, N72);
nand NAND3 (N540, N528, N352, N533);
nor NOR2 (N541, N384, N69);
buf BUF1 (N542, N536);
buf BUF1 (N543, N535);
xor XOR2 (N544, N543, N11);
buf BUF1 (N545, N542);
nand NAND2 (N546, N540, N41);
not NOT1 (N547, N539);
buf BUF1 (N548, N546);
buf BUF1 (N549, N530);
and AND2 (N550, N532, N48);
nor NOR2 (N551, N545, N544);
xor XOR2 (N552, N5, N278);
xor XOR2 (N553, N550, N304);
nand NAND2 (N554, N553, N177);
nor NOR2 (N555, N554, N171);
and AND4 (N556, N538, N70, N230, N262);
and AND3 (N557, N541, N469, N236);
or OR2 (N558, N552, N319);
xor XOR2 (N559, N529, N536);
not NOT1 (N560, N551);
or OR3 (N561, N549, N284, N417);
nor NOR3 (N562, N548, N498, N133);
not NOT1 (N563, N555);
buf BUF1 (N564, N503);
not NOT1 (N565, N556);
and AND2 (N566, N557, N68);
nand NAND2 (N567, N563, N563);
not NOT1 (N568, N566);
not NOT1 (N569, N562);
and AND2 (N570, N568, N171);
nand NAND4 (N571, N558, N385, N472, N206);
xor XOR2 (N572, N571, N309);
xor XOR2 (N573, N572, N507);
and AND4 (N574, N569, N270, N287, N522);
or OR2 (N575, N559, N156);
buf BUF1 (N576, N565);
nor NOR2 (N577, N575, N264);
nand NAND2 (N578, N574, N142);
or OR3 (N579, N547, N275, N249);
and AND2 (N580, N564, N266);
nor NOR4 (N581, N561, N162, N399, N424);
nand NAND4 (N582, N570, N499, N228, N51);
or OR4 (N583, N567, N578, N370, N57);
nor NOR4 (N584, N446, N348, N542, N109);
not NOT1 (N585, N573);
nand NAND3 (N586, N579, N63, N333);
xor XOR2 (N587, N585, N507);
nor NOR2 (N588, N584, N224);
or OR2 (N589, N560, N166);
not NOT1 (N590, N586);
not NOT1 (N591, N582);
nand NAND4 (N592, N591, N47, N335, N187);
nor NOR4 (N593, N576, N467, N490, N124);
nand NAND4 (N594, N587, N121, N541, N67);
xor XOR2 (N595, N589, N252);
xor XOR2 (N596, N592, N490);
or OR2 (N597, N590, N437);
buf BUF1 (N598, N580);
or OR2 (N599, N588, N273);
xor XOR2 (N600, N597, N538);
or OR2 (N601, N577, N551);
not NOT1 (N602, N595);
xor XOR2 (N603, N594, N565);
nand NAND2 (N604, N598, N488);
xor XOR2 (N605, N600, N550);
and AND3 (N606, N596, N475, N464);
nand NAND3 (N607, N606, N495, N343);
and AND2 (N608, N607, N356);
nor NOR2 (N609, N599, N81);
nor NOR3 (N610, N604, N98, N504);
nor NOR3 (N611, N610, N208, N274);
not NOT1 (N612, N593);
not NOT1 (N613, N583);
buf BUF1 (N614, N603);
buf BUF1 (N615, N612);
or OR3 (N616, N614, N119, N527);
nor NOR4 (N617, N601, N450, N51, N394);
and AND4 (N618, N581, N437, N402, N569);
nand NAND2 (N619, N616, N172);
nor NOR3 (N620, N602, N363, N389);
not NOT1 (N621, N615);
xor XOR2 (N622, N618, N526);
and AND3 (N623, N609, N569, N381);
and AND3 (N624, N617, N383, N269);
or OR2 (N625, N613, N231);
xor XOR2 (N626, N611, N255);
xor XOR2 (N627, N626, N382);
not NOT1 (N628, N608);
xor XOR2 (N629, N625, N179);
nor NOR4 (N630, N622, N484, N297, N300);
nand NAND4 (N631, N627, N61, N213, N336);
nand NAND2 (N632, N631, N552);
and AND2 (N633, N629, N103);
or OR2 (N634, N619, N318);
xor XOR2 (N635, N633, N143);
buf BUF1 (N636, N605);
xor XOR2 (N637, N623, N46);
not NOT1 (N638, N632);
xor XOR2 (N639, N637, N403);
xor XOR2 (N640, N624, N452);
buf BUF1 (N641, N640);
buf BUF1 (N642, N636);
xor XOR2 (N643, N642, N448);
nor NOR2 (N644, N638, N592);
and AND3 (N645, N630, N341, N213);
nand NAND4 (N646, N645, N619, N629, N438);
buf BUF1 (N647, N639);
or OR3 (N648, N644, N197, N153);
xor XOR2 (N649, N620, N384);
nand NAND4 (N650, N647, N498, N222, N170);
and AND4 (N651, N650, N544, N329, N317);
or OR4 (N652, N634, N301, N525, N573);
nand NAND2 (N653, N651, N326);
xor XOR2 (N654, N648, N177);
not NOT1 (N655, N643);
nand NAND4 (N656, N649, N654, N393, N381);
and AND4 (N657, N344, N109, N530, N421);
and AND2 (N658, N653, N232);
buf BUF1 (N659, N655);
nand NAND3 (N660, N656, N554, N58);
nand NAND2 (N661, N652, N47);
and AND2 (N662, N646, N463);
nand NAND4 (N663, N621, N361, N80, N519);
nor NOR2 (N664, N658, N98);
not NOT1 (N665, N641);
not NOT1 (N666, N628);
nor NOR3 (N667, N662, N476, N13);
or OR3 (N668, N661, N649, N614);
nor NOR4 (N669, N667, N475, N336, N262);
nand NAND3 (N670, N663, N371, N440);
nand NAND3 (N671, N668, N422, N275);
buf BUF1 (N672, N659);
nand NAND2 (N673, N671, N321);
and AND4 (N674, N670, N319, N379, N598);
and AND2 (N675, N635, N107);
nand NAND3 (N676, N672, N288, N508);
xor XOR2 (N677, N660, N542);
not NOT1 (N678, N675);
xor XOR2 (N679, N665, N186);
or OR2 (N680, N678, N155);
or OR2 (N681, N666, N452);
not NOT1 (N682, N680);
nor NOR4 (N683, N674, N119, N665, N632);
not NOT1 (N684, N683);
buf BUF1 (N685, N676);
xor XOR2 (N686, N664, N15);
or OR3 (N687, N669, N511, N637);
buf BUF1 (N688, N681);
buf BUF1 (N689, N688);
buf BUF1 (N690, N673);
buf BUF1 (N691, N684);
nor NOR3 (N692, N686, N291, N654);
buf BUF1 (N693, N682);
nand NAND2 (N694, N690, N267);
or OR2 (N695, N694, N390);
nand NAND3 (N696, N695, N670, N215);
not NOT1 (N697, N696);
nor NOR2 (N698, N697, N583);
xor XOR2 (N699, N685, N469);
xor XOR2 (N700, N691, N500);
xor XOR2 (N701, N677, N108);
nand NAND4 (N702, N698, N474, N281, N94);
buf BUF1 (N703, N687);
and AND2 (N704, N679, N655);
nor NOR3 (N705, N701, N73, N616);
buf BUF1 (N706, N699);
or OR4 (N707, N702, N566, N295, N318);
xor XOR2 (N708, N657, N320);
nor NOR3 (N709, N707, N123, N254);
buf BUF1 (N710, N692);
xor XOR2 (N711, N705, N51);
or OR4 (N712, N708, N58, N401, N275);
xor XOR2 (N713, N703, N643);
nand NAND2 (N714, N712, N492);
xor XOR2 (N715, N709, N565);
xor XOR2 (N716, N689, N245);
nor NOR3 (N717, N715, N60, N696);
not NOT1 (N718, N704);
nand NAND4 (N719, N693, N22, N37, N674);
xor XOR2 (N720, N713, N693);
nor NOR4 (N721, N700, N408, N161, N635);
nand NAND2 (N722, N706, N59);
and AND3 (N723, N714, N679, N73);
or OR3 (N724, N718, N375, N81);
or OR2 (N725, N717, N685);
nor NOR4 (N726, N710, N1, N521, N413);
nor NOR3 (N727, N725, N323, N401);
nand NAND2 (N728, N720, N64);
not NOT1 (N729, N727);
nand NAND4 (N730, N716, N493, N686, N345);
buf BUF1 (N731, N721);
xor XOR2 (N732, N729, N269);
buf BUF1 (N733, N723);
and AND3 (N734, N728, N351, N432);
not NOT1 (N735, N733);
and AND2 (N736, N711, N100);
or OR2 (N737, N724, N500);
nand NAND2 (N738, N730, N709);
nor NOR3 (N739, N735, N392, N665);
xor XOR2 (N740, N736, N284);
xor XOR2 (N741, N738, N469);
not NOT1 (N742, N734);
buf BUF1 (N743, N737);
xor XOR2 (N744, N743, N14);
nor NOR3 (N745, N731, N559, N167);
nor NOR2 (N746, N742, N160);
buf BUF1 (N747, N719);
nor NOR4 (N748, N745, N306, N450, N382);
xor XOR2 (N749, N741, N271);
buf BUF1 (N750, N726);
nand NAND2 (N751, N746, N33);
and AND3 (N752, N732, N166, N568);
nand NAND4 (N753, N750, N504, N658, N475);
nand NAND3 (N754, N753, N383, N172);
nand NAND2 (N755, N739, N316);
xor XOR2 (N756, N722, N272);
nor NOR2 (N757, N747, N737);
and AND4 (N758, N744, N164, N158, N118);
nand NAND4 (N759, N752, N457, N302, N521);
xor XOR2 (N760, N756, N266);
buf BUF1 (N761, N760);
buf BUF1 (N762, N740);
and AND2 (N763, N762, N88);
buf BUF1 (N764, N749);
nor NOR2 (N765, N755, N699);
nor NOR2 (N766, N751, N681);
or OR2 (N767, N763, N413);
buf BUF1 (N768, N758);
xor XOR2 (N769, N765, N179);
nor NOR2 (N770, N754, N74);
buf BUF1 (N771, N757);
not NOT1 (N772, N766);
xor XOR2 (N773, N764, N445);
nand NAND3 (N774, N772, N459, N203);
and AND2 (N775, N748, N171);
not NOT1 (N776, N774);
nand NAND2 (N777, N767, N543);
buf BUF1 (N778, N776);
or OR4 (N779, N778, N61, N671, N117);
nand NAND3 (N780, N777, N330, N370);
buf BUF1 (N781, N780);
or OR3 (N782, N775, N213, N480);
or OR4 (N783, N770, N610, N540, N251);
or OR2 (N784, N771, N427);
and AND4 (N785, N769, N734, N141, N661);
xor XOR2 (N786, N773, N570);
and AND2 (N787, N779, N332);
and AND2 (N788, N783, N673);
nor NOR3 (N789, N784, N560, N345);
not NOT1 (N790, N789);
not NOT1 (N791, N759);
buf BUF1 (N792, N786);
or OR3 (N793, N761, N229, N229);
and AND3 (N794, N785, N439, N591);
or OR4 (N795, N788, N442, N229, N781);
nor NOR2 (N796, N197, N653);
xor XOR2 (N797, N793, N153);
buf BUF1 (N798, N782);
nor NOR2 (N799, N798, N599);
nor NOR2 (N800, N792, N449);
xor XOR2 (N801, N797, N9);
and AND4 (N802, N795, N35, N449, N628);
xor XOR2 (N803, N794, N266);
xor XOR2 (N804, N790, N661);
nand NAND3 (N805, N804, N460, N570);
nand NAND2 (N806, N791, N585);
xor XOR2 (N807, N802, N793);
not NOT1 (N808, N801);
and AND3 (N809, N807, N54, N316);
buf BUF1 (N810, N796);
buf BUF1 (N811, N803);
and AND4 (N812, N805, N690, N471, N485);
or OR3 (N813, N812, N120, N82);
not NOT1 (N814, N813);
not NOT1 (N815, N768);
not NOT1 (N816, N806);
or OR2 (N817, N815, N170);
not NOT1 (N818, N811);
buf BUF1 (N819, N810);
nor NOR3 (N820, N814, N769, N113);
nand NAND2 (N821, N799, N625);
xor XOR2 (N822, N820, N620);
not NOT1 (N823, N808);
nand NAND4 (N824, N819, N5, N415, N87);
and AND4 (N825, N824, N354, N470, N490);
buf BUF1 (N826, N816);
buf BUF1 (N827, N825);
or OR4 (N828, N787, N275, N532, N118);
xor XOR2 (N829, N800, N151);
and AND3 (N830, N826, N599, N148);
nand NAND4 (N831, N818, N551, N656, N31);
nor NOR4 (N832, N822, N242, N19, N532);
not NOT1 (N833, N830);
xor XOR2 (N834, N833, N494);
and AND3 (N835, N832, N301, N216);
nand NAND4 (N836, N828, N749, N100, N470);
and AND3 (N837, N821, N489, N167);
and AND2 (N838, N827, N105);
nand NAND2 (N839, N835, N790);
xor XOR2 (N840, N817, N202);
nor NOR3 (N841, N831, N770, N722);
not NOT1 (N842, N839);
not NOT1 (N843, N809);
not NOT1 (N844, N837);
nand NAND4 (N845, N834, N835, N227, N786);
nand NAND3 (N846, N844, N612, N841);
nand NAND3 (N847, N174, N129, N104);
and AND2 (N848, N838, N385);
xor XOR2 (N849, N823, N443);
and AND2 (N850, N845, N383);
nand NAND4 (N851, N840, N393, N727, N486);
and AND2 (N852, N851, N528);
nor NOR3 (N853, N843, N429, N424);
nand NAND3 (N854, N848, N302, N508);
and AND3 (N855, N847, N183, N385);
nor NOR3 (N856, N829, N115, N609);
or OR3 (N857, N853, N446, N550);
not NOT1 (N858, N846);
nor NOR2 (N859, N854, N16);
or OR4 (N860, N836, N543, N549, N95);
buf BUF1 (N861, N842);
nand NAND2 (N862, N859, N787);
not NOT1 (N863, N850);
xor XOR2 (N864, N856, N148);
or OR3 (N865, N852, N292, N309);
not NOT1 (N866, N849);
nor NOR2 (N867, N861, N128);
buf BUF1 (N868, N863);
and AND4 (N869, N855, N467, N467, N773);
nor NOR3 (N870, N867, N325, N514);
nor NOR3 (N871, N864, N434, N657);
xor XOR2 (N872, N870, N337);
not NOT1 (N873, N868);
buf BUF1 (N874, N865);
nand NAND2 (N875, N857, N376);
xor XOR2 (N876, N862, N298);
nor NOR3 (N877, N858, N519, N271);
buf BUF1 (N878, N872);
nor NOR2 (N879, N871, N590);
and AND3 (N880, N874, N329, N817);
buf BUF1 (N881, N866);
or OR4 (N882, N875, N825, N702, N510);
or OR3 (N883, N876, N72, N223);
or OR4 (N884, N873, N721, N104, N157);
or OR3 (N885, N877, N615, N664);
not NOT1 (N886, N885);
buf BUF1 (N887, N860);
buf BUF1 (N888, N887);
not NOT1 (N889, N880);
nor NOR4 (N890, N869, N80, N508, N799);
xor XOR2 (N891, N879, N298);
buf BUF1 (N892, N890);
or OR3 (N893, N888, N651, N489);
not NOT1 (N894, N891);
or OR3 (N895, N882, N81, N425);
nand NAND4 (N896, N884, N232, N198, N41);
xor XOR2 (N897, N886, N532);
or OR4 (N898, N894, N457, N657, N534);
nand NAND2 (N899, N881, N816);
not NOT1 (N900, N899);
or OR2 (N901, N889, N893);
or OR4 (N902, N754, N851, N386, N761);
and AND4 (N903, N883, N614, N552, N848);
nand NAND4 (N904, N901, N454, N290, N30);
nor NOR3 (N905, N878, N716, N123);
nand NAND2 (N906, N895, N208);
and AND2 (N907, N906, N10);
not NOT1 (N908, N896);
xor XOR2 (N909, N902, N596);
nand NAND2 (N910, N903, N597);
nand NAND2 (N911, N900, N64);
xor XOR2 (N912, N909, N46);
xor XOR2 (N913, N897, N436);
not NOT1 (N914, N905);
nand NAND2 (N915, N910, N422);
and AND2 (N916, N904, N906);
nand NAND2 (N917, N907, N742);
nand NAND3 (N918, N915, N427, N912);
nor NOR2 (N919, N798, N220);
nor NOR4 (N920, N918, N74, N483, N650);
xor XOR2 (N921, N917, N646);
buf BUF1 (N922, N911);
or OR4 (N923, N908, N689, N697, N238);
buf BUF1 (N924, N892);
not NOT1 (N925, N923);
nor NOR2 (N926, N921, N368);
and AND4 (N927, N924, N135, N357, N17);
nand NAND3 (N928, N919, N5, N844);
not NOT1 (N929, N914);
nor NOR2 (N930, N922, N782);
or OR3 (N931, N926, N640, N113);
or OR3 (N932, N920, N803, N805);
nor NOR3 (N933, N932, N249, N181);
or OR3 (N934, N929, N652, N585);
nor NOR4 (N935, N898, N917, N325, N383);
nor NOR2 (N936, N931, N667);
or OR3 (N937, N936, N54, N696);
nor NOR2 (N938, N934, N623);
or OR4 (N939, N916, N400, N60, N643);
not NOT1 (N940, N927);
not NOT1 (N941, N925);
not NOT1 (N942, N939);
not NOT1 (N943, N933);
nor NOR4 (N944, N943, N756, N627, N101);
xor XOR2 (N945, N940, N128);
or OR3 (N946, N913, N319, N87);
nand NAND2 (N947, N942, N547);
buf BUF1 (N948, N938);
or OR4 (N949, N948, N282, N318, N604);
nand NAND3 (N950, N941, N540, N866);
nand NAND4 (N951, N950, N679, N594, N812);
not NOT1 (N952, N946);
xor XOR2 (N953, N949, N173);
nor NOR2 (N954, N944, N177);
or OR3 (N955, N930, N872, N308);
or OR3 (N956, N952, N186, N48);
buf BUF1 (N957, N951);
or OR4 (N958, N955, N909, N412, N463);
buf BUF1 (N959, N953);
not NOT1 (N960, N937);
nand NAND3 (N961, N958, N544, N856);
and AND2 (N962, N947, N557);
not NOT1 (N963, N954);
nand NAND2 (N964, N959, N268);
nand NAND4 (N965, N957, N155, N316, N776);
nand NAND3 (N966, N928, N529, N338);
nor NOR4 (N967, N945, N410, N910, N302);
nor NOR2 (N968, N961, N8);
or OR4 (N969, N968, N728, N460, N25);
or OR2 (N970, N969, N537);
buf BUF1 (N971, N965);
xor XOR2 (N972, N963, N58);
not NOT1 (N973, N964);
and AND4 (N974, N960, N446, N429, N484);
nand NAND3 (N975, N966, N718, N208);
nand NAND4 (N976, N973, N841, N479, N643);
nand NAND4 (N977, N975, N880, N970, N698);
or OR2 (N978, N375, N243);
nor NOR4 (N979, N977, N62, N592, N588);
not NOT1 (N980, N978);
or OR2 (N981, N980, N739);
buf BUF1 (N982, N962);
and AND2 (N983, N956, N765);
not NOT1 (N984, N972);
or OR3 (N985, N935, N547, N829);
nor NOR3 (N986, N983, N154, N533);
xor XOR2 (N987, N984, N349);
or OR2 (N988, N986, N644);
or OR2 (N989, N979, N244);
or OR3 (N990, N976, N863, N651);
not NOT1 (N991, N990);
nor NOR3 (N992, N981, N103, N914);
and AND2 (N993, N974, N383);
and AND2 (N994, N988, N568);
xor XOR2 (N995, N989, N503);
nor NOR3 (N996, N967, N146, N989);
or OR3 (N997, N985, N4, N502);
and AND4 (N998, N993, N216, N832, N834);
not NOT1 (N999, N971);
nand NAND3 (N1000, N999, N312, N516);
buf BUF1 (N1001, N994);
and AND4 (N1002, N982, N230, N73, N794);
nor NOR3 (N1003, N998, N971, N489);
and AND4 (N1004, N992, N860, N189, N974);
not NOT1 (N1005, N1003);
not NOT1 (N1006, N1004);
nand NAND2 (N1007, N1000, N457);
buf BUF1 (N1008, N1002);
and AND3 (N1009, N1006, N525, N417);
buf BUF1 (N1010, N997);
nor NOR2 (N1011, N995, N736);
and AND3 (N1012, N1001, N505, N972);
or OR4 (N1013, N1010, N673, N777, N772);
or OR2 (N1014, N1007, N714);
nor NOR4 (N1015, N1013, N180, N551, N345);
xor XOR2 (N1016, N1005, N178);
nor NOR4 (N1017, N1009, N521, N783, N348);
buf BUF1 (N1018, N991);
not NOT1 (N1019, N1008);
nand NAND2 (N1020, N1014, N178);
or OR2 (N1021, N1017, N388);
not NOT1 (N1022, N1016);
buf BUF1 (N1023, N1020);
nor NOR3 (N1024, N1015, N748, N91);
xor XOR2 (N1025, N1018, N540);
xor XOR2 (N1026, N1023, N533);
and AND3 (N1027, N1011, N555, N211);
not NOT1 (N1028, N1024);
and AND2 (N1029, N1012, N563);
nand NAND3 (N1030, N987, N391, N347);
xor XOR2 (N1031, N996, N901);
not NOT1 (N1032, N1030);
not NOT1 (N1033, N1032);
xor XOR2 (N1034, N1021, N865);
xor XOR2 (N1035, N1026, N258);
nand NAND3 (N1036, N1022, N146, N757);
nor NOR2 (N1037, N1031, N919);
or OR3 (N1038, N1037, N711, N471);
or OR2 (N1039, N1033, N609);
xor XOR2 (N1040, N1039, N776);
and AND2 (N1041, N1028, N815);
buf BUF1 (N1042, N1019);
nand NAND4 (N1043, N1025, N384, N251, N897);
or OR4 (N1044, N1034, N707, N1014, N34);
and AND2 (N1045, N1038, N842);
nand NAND3 (N1046, N1044, N979, N909);
nor NOR4 (N1047, N1035, N53, N52, N1044);
or OR3 (N1048, N1043, N588, N870);
not NOT1 (N1049, N1042);
and AND4 (N1050, N1029, N243, N994, N5);
xor XOR2 (N1051, N1050, N581);
nor NOR2 (N1052, N1049, N467);
and AND3 (N1053, N1036, N281, N1047);
and AND3 (N1054, N187, N405, N938);
not NOT1 (N1055, N1052);
nor NOR2 (N1056, N1048, N510);
or OR4 (N1057, N1053, N969, N655, N406);
and AND2 (N1058, N1057, N809);
xor XOR2 (N1059, N1056, N715);
not NOT1 (N1060, N1041);
xor XOR2 (N1061, N1045, N466);
or OR3 (N1062, N1061, N813, N782);
buf BUF1 (N1063, N1055);
or OR4 (N1064, N1051, N555, N609, N821);
buf BUF1 (N1065, N1058);
not NOT1 (N1066, N1065);
buf BUF1 (N1067, N1040);
and AND2 (N1068, N1066, N975);
or OR2 (N1069, N1027, N709);
nor NOR2 (N1070, N1068, N1029);
buf BUF1 (N1071, N1069);
or OR4 (N1072, N1070, N268, N1028, N241);
buf BUF1 (N1073, N1060);
xor XOR2 (N1074, N1064, N193);
nor NOR3 (N1075, N1046, N406, N291);
or OR2 (N1076, N1063, N98);
and AND3 (N1077, N1071, N8, N837);
nand NAND4 (N1078, N1067, N435, N113, N630);
nor NOR2 (N1079, N1054, N412);
buf BUF1 (N1080, N1059);
nand NAND3 (N1081, N1076, N736, N466);
nor NOR2 (N1082, N1081, N229);
or OR4 (N1083, N1080, N483, N41, N417);
or OR2 (N1084, N1073, N550);
xor XOR2 (N1085, N1078, N747);
nand NAND3 (N1086, N1074, N4, N431);
buf BUF1 (N1087, N1079);
nand NAND3 (N1088, N1084, N837, N118);
or OR2 (N1089, N1088, N344);
xor XOR2 (N1090, N1085, N940);
nor NOR3 (N1091, N1087, N287, N688);
not NOT1 (N1092, N1077);
and AND2 (N1093, N1091, N510);
nand NAND3 (N1094, N1089, N726, N340);
not NOT1 (N1095, N1094);
and AND4 (N1096, N1086, N763, N1053, N2);
nand NAND3 (N1097, N1090, N577, N1069);
nor NOR3 (N1098, N1092, N16, N382);
nand NAND4 (N1099, N1093, N478, N670, N508);
xor XOR2 (N1100, N1062, N841);
buf BUF1 (N1101, N1100);
not NOT1 (N1102, N1095);
or OR4 (N1103, N1083, N935, N602, N133);
xor XOR2 (N1104, N1097, N588);
nand NAND4 (N1105, N1082, N288, N712, N239);
or OR2 (N1106, N1099, N406);
not NOT1 (N1107, N1106);
xor XOR2 (N1108, N1072, N804);
xor XOR2 (N1109, N1075, N867);
not NOT1 (N1110, N1096);
not NOT1 (N1111, N1101);
and AND2 (N1112, N1110, N117);
and AND4 (N1113, N1105, N687, N1086, N588);
xor XOR2 (N1114, N1103, N335);
nand NAND4 (N1115, N1112, N457, N652, N969);
and AND4 (N1116, N1113, N950, N341, N434);
and AND4 (N1117, N1102, N415, N984, N462);
xor XOR2 (N1118, N1115, N275);
not NOT1 (N1119, N1109);
or OR2 (N1120, N1107, N57);
buf BUF1 (N1121, N1118);
and AND3 (N1122, N1111, N450, N758);
buf BUF1 (N1123, N1117);
and AND3 (N1124, N1121, N752, N1061);
nor NOR2 (N1125, N1122, N791);
nand NAND3 (N1126, N1120, N1043, N699);
not NOT1 (N1127, N1124);
nor NOR3 (N1128, N1125, N378, N145);
and AND4 (N1129, N1123, N798, N753, N1088);
nand NAND3 (N1130, N1114, N587, N1025);
or OR3 (N1131, N1119, N305, N435);
or OR3 (N1132, N1126, N310, N870);
nand NAND3 (N1133, N1127, N842, N704);
buf BUF1 (N1134, N1130);
or OR2 (N1135, N1116, N626);
nor NOR4 (N1136, N1135, N213, N221, N412);
nand NAND3 (N1137, N1136, N1111, N552);
nand NAND2 (N1138, N1134, N1125);
xor XOR2 (N1139, N1131, N500);
xor XOR2 (N1140, N1108, N1032);
buf BUF1 (N1141, N1140);
nor NOR4 (N1142, N1141, N550, N43, N283);
nand NAND3 (N1143, N1139, N621, N91);
or OR4 (N1144, N1104, N20, N191, N212);
nand NAND2 (N1145, N1144, N1092);
xor XOR2 (N1146, N1128, N595);
buf BUF1 (N1147, N1146);
not NOT1 (N1148, N1145);
buf BUF1 (N1149, N1098);
not NOT1 (N1150, N1149);
not NOT1 (N1151, N1138);
buf BUF1 (N1152, N1129);
not NOT1 (N1153, N1132);
not NOT1 (N1154, N1142);
and AND2 (N1155, N1148, N1036);
not NOT1 (N1156, N1155);
xor XOR2 (N1157, N1137, N385);
and AND4 (N1158, N1152, N586, N661, N636);
nor NOR3 (N1159, N1154, N37, N247);
xor XOR2 (N1160, N1158, N364);
nor NOR4 (N1161, N1151, N16, N551, N327);
or OR4 (N1162, N1159, N911, N205, N25);
or OR2 (N1163, N1157, N522);
nand NAND4 (N1164, N1133, N1158, N1145, N761);
not NOT1 (N1165, N1162);
not NOT1 (N1166, N1164);
or OR4 (N1167, N1166, N332, N28, N503);
and AND4 (N1168, N1163, N1073, N853, N39);
or OR3 (N1169, N1168, N631, N294);
nor NOR3 (N1170, N1165, N217, N539);
not NOT1 (N1171, N1143);
or OR3 (N1172, N1147, N33, N485);
nor NOR4 (N1173, N1172, N130, N812, N150);
and AND3 (N1174, N1170, N827, N214);
or OR2 (N1175, N1174, N342);
nand NAND2 (N1176, N1173, N1144);
nor NOR3 (N1177, N1167, N229, N238);
xor XOR2 (N1178, N1169, N11);
not NOT1 (N1179, N1156);
nor NOR2 (N1180, N1171, N1080);
buf BUF1 (N1181, N1180);
buf BUF1 (N1182, N1161);
xor XOR2 (N1183, N1176, N168);
not NOT1 (N1184, N1177);
or OR4 (N1185, N1179, N957, N416, N449);
or OR4 (N1186, N1183, N743, N817, N280);
xor XOR2 (N1187, N1178, N325);
xor XOR2 (N1188, N1150, N963);
xor XOR2 (N1189, N1184, N762);
nand NAND2 (N1190, N1187, N615);
nand NAND4 (N1191, N1175, N204, N906, N1072);
and AND3 (N1192, N1181, N660, N322);
nand NAND3 (N1193, N1188, N1075, N24);
not NOT1 (N1194, N1185);
nor NOR3 (N1195, N1189, N130, N1041);
and AND4 (N1196, N1191, N211, N229, N313);
xor XOR2 (N1197, N1153, N872);
nor NOR4 (N1198, N1193, N1100, N995, N576);
or OR2 (N1199, N1194, N300);
nand NAND4 (N1200, N1182, N631, N288, N1164);
not NOT1 (N1201, N1190);
buf BUF1 (N1202, N1201);
and AND2 (N1203, N1202, N1123);
and AND2 (N1204, N1186, N713);
nand NAND4 (N1205, N1195, N788, N725, N400);
not NOT1 (N1206, N1200);
buf BUF1 (N1207, N1196);
nand NAND4 (N1208, N1207, N1141, N1141, N76);
xor XOR2 (N1209, N1208, N924);
and AND2 (N1210, N1205, N36);
buf BUF1 (N1211, N1192);
and AND4 (N1212, N1206, N783, N610, N1074);
buf BUF1 (N1213, N1204);
buf BUF1 (N1214, N1210);
buf BUF1 (N1215, N1211);
and AND2 (N1216, N1215, N15);
or OR2 (N1217, N1209, N18);
and AND2 (N1218, N1216, N534);
or OR4 (N1219, N1160, N1008, N1023, N1136);
and AND2 (N1220, N1213, N294);
and AND4 (N1221, N1197, N358, N487, N1138);
nor NOR4 (N1222, N1217, N749, N16, N239);
and AND2 (N1223, N1198, N469);
nor NOR3 (N1224, N1222, N553, N924);
not NOT1 (N1225, N1214);
or OR3 (N1226, N1218, N1032, N930);
not NOT1 (N1227, N1226);
nor NOR3 (N1228, N1224, N183, N572);
xor XOR2 (N1229, N1221, N707);
nand NAND2 (N1230, N1225, N1098);
and AND2 (N1231, N1212, N241);
or OR2 (N1232, N1199, N1003);
nand NAND3 (N1233, N1232, N606, N752);
or OR2 (N1234, N1229, N262);
nor NOR3 (N1235, N1203, N994, N1146);
not NOT1 (N1236, N1234);
not NOT1 (N1237, N1223);
nor NOR2 (N1238, N1233, N252);
buf BUF1 (N1239, N1235);
buf BUF1 (N1240, N1230);
buf BUF1 (N1241, N1238);
nor NOR2 (N1242, N1240, N172);
nand NAND4 (N1243, N1242, N408, N169, N835);
or OR3 (N1244, N1219, N29, N476);
buf BUF1 (N1245, N1241);
nor NOR3 (N1246, N1237, N700, N75);
nor NOR2 (N1247, N1227, N272);
not NOT1 (N1248, N1245);
nor NOR3 (N1249, N1220, N111, N837);
not NOT1 (N1250, N1247);
buf BUF1 (N1251, N1243);
nand NAND4 (N1252, N1246, N437, N138, N935);
or OR2 (N1253, N1244, N604);
or OR3 (N1254, N1231, N896, N132);
not NOT1 (N1255, N1236);
not NOT1 (N1256, N1253);
or OR2 (N1257, N1250, N34);
and AND4 (N1258, N1256, N1238, N1187, N1172);
not NOT1 (N1259, N1252);
buf BUF1 (N1260, N1258);
or OR4 (N1261, N1239, N891, N18, N1185);
and AND4 (N1262, N1261, N760, N557, N187);
nand NAND2 (N1263, N1255, N1036);
or OR2 (N1264, N1263, N980);
or OR2 (N1265, N1254, N494);
nor NOR4 (N1266, N1248, N167, N110, N455);
or OR2 (N1267, N1251, N427);
not NOT1 (N1268, N1257);
not NOT1 (N1269, N1264);
xor XOR2 (N1270, N1259, N117);
nand NAND4 (N1271, N1249, N1131, N1259, N202);
xor XOR2 (N1272, N1228, N99);
not NOT1 (N1273, N1262);
not NOT1 (N1274, N1273);
or OR3 (N1275, N1271, N901, N666);
and AND3 (N1276, N1275, N437, N230);
xor XOR2 (N1277, N1267, N112);
nor NOR2 (N1278, N1266, N955);
buf BUF1 (N1279, N1274);
nand NAND4 (N1280, N1277, N1129, N532, N1203);
and AND2 (N1281, N1265, N43);
nor NOR4 (N1282, N1281, N1023, N569, N25);
and AND4 (N1283, N1282, N478, N102, N1024);
buf BUF1 (N1284, N1278);
and AND2 (N1285, N1269, N1245);
or OR4 (N1286, N1279, N864, N984, N193);
or OR2 (N1287, N1276, N1268);
xor XOR2 (N1288, N603, N297);
xor XOR2 (N1289, N1272, N587);
or OR3 (N1290, N1289, N336, N1246);
or OR4 (N1291, N1260, N402, N283, N355);
xor XOR2 (N1292, N1283, N28);
nand NAND4 (N1293, N1287, N950, N591, N886);
or OR2 (N1294, N1288, N75);
buf BUF1 (N1295, N1284);
and AND2 (N1296, N1295, N987);
or OR4 (N1297, N1292, N1224, N363, N1162);
buf BUF1 (N1298, N1297);
buf BUF1 (N1299, N1298);
not NOT1 (N1300, N1296);
nand NAND4 (N1301, N1294, N757, N133, N88);
and AND2 (N1302, N1300, N673);
buf BUF1 (N1303, N1285);
or OR3 (N1304, N1299, N400, N887);
and AND4 (N1305, N1302, N959, N1144, N588);
and AND3 (N1306, N1303, N435, N959);
nand NAND2 (N1307, N1286, N1280);
nor NOR4 (N1308, N1180, N64, N589, N313);
buf BUF1 (N1309, N1304);
xor XOR2 (N1310, N1308, N1268);
xor XOR2 (N1311, N1270, N990);
not NOT1 (N1312, N1306);
nor NOR4 (N1313, N1305, N460, N250, N927);
nand NAND3 (N1314, N1312, N560, N716);
nor NOR4 (N1315, N1311, N911, N176, N383);
or OR3 (N1316, N1301, N1214, N694);
buf BUF1 (N1317, N1307);
nand NAND4 (N1318, N1291, N736, N188, N178);
xor XOR2 (N1319, N1309, N1105);
not NOT1 (N1320, N1316);
not NOT1 (N1321, N1319);
buf BUF1 (N1322, N1321);
nand NAND3 (N1323, N1320, N911, N694);
nor NOR3 (N1324, N1315, N1010, N256);
not NOT1 (N1325, N1290);
buf BUF1 (N1326, N1324);
xor XOR2 (N1327, N1326, N675);
nor NOR3 (N1328, N1325, N378, N187);
or OR4 (N1329, N1314, N55, N91, N74);
or OR2 (N1330, N1327, N319);
buf BUF1 (N1331, N1329);
buf BUF1 (N1332, N1313);
not NOT1 (N1333, N1310);
buf BUF1 (N1334, N1317);
nor NOR3 (N1335, N1323, N293, N1058);
and AND3 (N1336, N1293, N815, N1193);
not NOT1 (N1337, N1336);
and AND3 (N1338, N1334, N1143, N1302);
and AND3 (N1339, N1322, N919, N92);
nand NAND4 (N1340, N1339, N1018, N552, N238);
or OR4 (N1341, N1335, N823, N511, N777);
or OR4 (N1342, N1332, N1118, N197, N836);
or OR3 (N1343, N1331, N509, N1299);
or OR3 (N1344, N1330, N604, N165);
xor XOR2 (N1345, N1333, N888);
or OR4 (N1346, N1341, N798, N1227, N900);
or OR2 (N1347, N1343, N190);
or OR4 (N1348, N1337, N671, N485, N50);
nor NOR2 (N1349, N1348, N1269);
buf BUF1 (N1350, N1349);
nand NAND2 (N1351, N1347, N954);
nor NOR4 (N1352, N1344, N1097, N663, N240);
xor XOR2 (N1353, N1338, N409);
not NOT1 (N1354, N1328);
and AND2 (N1355, N1350, N348);
not NOT1 (N1356, N1340);
nor NOR2 (N1357, N1346, N1223);
nor NOR4 (N1358, N1318, N257, N745, N47);
nor NOR2 (N1359, N1353, N256);
xor XOR2 (N1360, N1359, N458);
nand NAND2 (N1361, N1360, N38);
or OR4 (N1362, N1357, N78, N1276, N1109);
or OR3 (N1363, N1345, N845, N466);
and AND3 (N1364, N1342, N321, N372);
and AND2 (N1365, N1361, N285);
nand NAND3 (N1366, N1363, N1258, N798);
or OR2 (N1367, N1355, N768);
and AND4 (N1368, N1365, N1126, N90, N480);
xor XOR2 (N1369, N1354, N795);
buf BUF1 (N1370, N1358);
nor NOR4 (N1371, N1362, N509, N787, N151);
or OR2 (N1372, N1356, N1085);
nor NOR4 (N1373, N1370, N692, N710, N478);
nor NOR3 (N1374, N1369, N979, N601);
not NOT1 (N1375, N1372);
nand NAND3 (N1376, N1375, N790, N73);
not NOT1 (N1377, N1352);
nor NOR3 (N1378, N1367, N1264, N706);
nand NAND4 (N1379, N1374, N851, N51, N39);
nand NAND2 (N1380, N1351, N772);
not NOT1 (N1381, N1366);
nor NOR4 (N1382, N1380, N83, N336, N851);
or OR2 (N1383, N1376, N40);
and AND3 (N1384, N1364, N532, N1097);
xor XOR2 (N1385, N1379, N91);
or OR3 (N1386, N1382, N64, N622);
buf BUF1 (N1387, N1371);
or OR3 (N1388, N1385, N235, N1382);
not NOT1 (N1389, N1387);
nand NAND3 (N1390, N1389, N814, N245);
buf BUF1 (N1391, N1377);
buf BUF1 (N1392, N1368);
nand NAND4 (N1393, N1384, N624, N631, N836);
and AND2 (N1394, N1386, N699);
buf BUF1 (N1395, N1381);
or OR4 (N1396, N1391, N899, N100, N1180);
and AND2 (N1397, N1394, N496);
and AND4 (N1398, N1383, N714, N383, N170);
or OR3 (N1399, N1388, N1077, N629);
nor NOR3 (N1400, N1393, N623, N1244);
xor XOR2 (N1401, N1396, N189);
and AND3 (N1402, N1400, N1234, N330);
or OR2 (N1403, N1397, N590);
and AND3 (N1404, N1378, N511, N1314);
xor XOR2 (N1405, N1395, N204);
or OR4 (N1406, N1404, N1080, N945, N1014);
xor XOR2 (N1407, N1406, N90);
and AND4 (N1408, N1399, N1057, N1280, N1331);
nor NOR4 (N1409, N1401, N491, N170, N1097);
xor XOR2 (N1410, N1409, N569);
nand NAND3 (N1411, N1402, N477, N1344);
xor XOR2 (N1412, N1411, N168);
not NOT1 (N1413, N1410);
xor XOR2 (N1414, N1403, N137);
buf BUF1 (N1415, N1407);
and AND2 (N1416, N1392, N138);
nand NAND3 (N1417, N1416, N775, N910);
nor NOR2 (N1418, N1373, N432);
or OR2 (N1419, N1405, N30);
nor NOR2 (N1420, N1414, N511);
buf BUF1 (N1421, N1413);
xor XOR2 (N1422, N1421, N597);
not NOT1 (N1423, N1398);
not NOT1 (N1424, N1412);
nor NOR2 (N1425, N1422, N491);
not NOT1 (N1426, N1423);
xor XOR2 (N1427, N1424, N970);
and AND4 (N1428, N1427, N107, N1182, N919);
and AND4 (N1429, N1419, N562, N1041, N639);
and AND3 (N1430, N1417, N1110, N366);
not NOT1 (N1431, N1408);
and AND2 (N1432, N1430, N352);
nand NAND3 (N1433, N1418, N1085, N791);
and AND3 (N1434, N1432, N1117, N1222);
and AND2 (N1435, N1433, N412);
or OR4 (N1436, N1429, N760, N872, N93);
or OR4 (N1437, N1420, N884, N872, N364);
xor XOR2 (N1438, N1415, N523);
or OR4 (N1439, N1425, N1318, N68, N1366);
and AND2 (N1440, N1428, N68);
xor XOR2 (N1441, N1439, N127);
and AND2 (N1442, N1435, N1359);
not NOT1 (N1443, N1434);
xor XOR2 (N1444, N1431, N842);
or OR2 (N1445, N1440, N152);
buf BUF1 (N1446, N1437);
buf BUF1 (N1447, N1442);
xor XOR2 (N1448, N1436, N203);
nand NAND2 (N1449, N1390, N904);
or OR2 (N1450, N1444, N855);
nor NOR3 (N1451, N1445, N945, N175);
nand NAND4 (N1452, N1438, N455, N652, N1033);
buf BUF1 (N1453, N1443);
and AND2 (N1454, N1450, N206);
buf BUF1 (N1455, N1449);
and AND3 (N1456, N1453, N1331, N372);
not NOT1 (N1457, N1454);
nor NOR2 (N1458, N1457, N112);
nor NOR3 (N1459, N1455, N928, N143);
buf BUF1 (N1460, N1426);
xor XOR2 (N1461, N1456, N776);
nor NOR4 (N1462, N1460, N468, N851, N660);
nand NAND2 (N1463, N1441, N474);
and AND4 (N1464, N1451, N342, N716, N269);
not NOT1 (N1465, N1446);
and AND2 (N1466, N1452, N236);
nor NOR4 (N1467, N1448, N1214, N714, N708);
xor XOR2 (N1468, N1459, N1185);
xor XOR2 (N1469, N1465, N298);
buf BUF1 (N1470, N1461);
not NOT1 (N1471, N1463);
buf BUF1 (N1472, N1447);
or OR4 (N1473, N1470, N935, N797, N491);
buf BUF1 (N1474, N1462);
xor XOR2 (N1475, N1458, N221);
nand NAND2 (N1476, N1471, N428);
nand NAND2 (N1477, N1468, N172);
not NOT1 (N1478, N1466);
xor XOR2 (N1479, N1474, N1444);
xor XOR2 (N1480, N1467, N1333);
not NOT1 (N1481, N1473);
not NOT1 (N1482, N1472);
buf BUF1 (N1483, N1475);
not NOT1 (N1484, N1476);
nand NAND4 (N1485, N1477, N185, N245, N551);
xor XOR2 (N1486, N1481, N328);
or OR3 (N1487, N1480, N476, N1443);
xor XOR2 (N1488, N1469, N916);
buf BUF1 (N1489, N1482);
nor NOR3 (N1490, N1479, N755, N1375);
nor NOR3 (N1491, N1490, N7, N1013);
buf BUF1 (N1492, N1483);
xor XOR2 (N1493, N1464, N714);
or OR4 (N1494, N1488, N838, N964, N285);
xor XOR2 (N1495, N1478, N32);
xor XOR2 (N1496, N1487, N26);
buf BUF1 (N1497, N1494);
buf BUF1 (N1498, N1495);
and AND3 (N1499, N1496, N951, N312);
nand NAND3 (N1500, N1498, N257, N62);
xor XOR2 (N1501, N1493, N499);
and AND4 (N1502, N1500, N61, N707, N1185);
not NOT1 (N1503, N1501);
or OR3 (N1504, N1497, N190, N1346);
or OR2 (N1505, N1485, N690);
or OR4 (N1506, N1503, N339, N1204, N1094);
not NOT1 (N1507, N1506);
or OR3 (N1508, N1492, N159, N825);
buf BUF1 (N1509, N1489);
nor NOR3 (N1510, N1499, N194, N269);
xor XOR2 (N1511, N1507, N254);
xor XOR2 (N1512, N1509, N1117);
endmodule