// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13;

output N808,N802,N810,N807,N792,N796,N809,N799,N812,N813;

buf BUF1 (N14, N3);
not NOT1 (N15, N10);
xor XOR2 (N16, N7, N15);
not NOT1 (N17, N10);
not NOT1 (N18, N3);
not NOT1 (N19, N6);
not NOT1 (N20, N3);
xor XOR2 (N21, N6, N1);
nand NAND3 (N22, N3, N17, N8);
and AND4 (N23, N10, N1, N10, N14);
or OR3 (N24, N6, N17, N3);
nor NOR3 (N25, N2, N8, N14);
nor NOR4 (N26, N16, N5, N6, N12);
nor NOR4 (N27, N20, N16, N24, N6);
and AND4 (N28, N10, N15, N22, N20);
nand NAND2 (N29, N13, N25);
xor XOR2 (N30, N10, N22);
xor XOR2 (N31, N15, N19);
xor XOR2 (N32, N18, N24);
buf BUF1 (N33, N11);
nand NAND2 (N34, N28, N31);
xor XOR2 (N35, N22, N8);
buf BUF1 (N36, N23);
or OR3 (N37, N33, N17, N35);
xor XOR2 (N38, N22, N35);
xor XOR2 (N39, N32, N6);
or OR2 (N40, N37, N6);
or OR2 (N41, N40, N3);
and AND3 (N42, N39, N9, N25);
buf BUF1 (N43, N38);
and AND2 (N44, N36, N13);
nor NOR3 (N45, N30, N34, N24);
buf BUF1 (N46, N21);
or OR4 (N47, N7, N23, N5, N15);
and AND2 (N48, N46, N18);
buf BUF1 (N49, N41);
buf BUF1 (N50, N48);
and AND3 (N51, N45, N5, N46);
xor XOR2 (N52, N47, N28);
or OR2 (N53, N42, N32);
xor XOR2 (N54, N50, N32);
or OR2 (N55, N44, N45);
buf BUF1 (N56, N55);
nand NAND4 (N57, N27, N4, N16, N33);
nor NOR2 (N58, N53, N25);
nor NOR3 (N59, N43, N6, N33);
nand NAND4 (N60, N57, N21, N49, N8);
xor XOR2 (N61, N4, N13);
and AND2 (N62, N60, N13);
or OR4 (N63, N29, N1, N60, N5);
buf BUF1 (N64, N56);
buf BUF1 (N65, N59);
xor XOR2 (N66, N51, N19);
and AND3 (N67, N65, N33, N7);
xor XOR2 (N68, N67, N30);
not NOT1 (N69, N26);
nand NAND3 (N70, N61, N43, N17);
buf BUF1 (N71, N54);
xor XOR2 (N72, N66, N71);
and AND3 (N73, N22, N63, N65);
not NOT1 (N74, N73);
not NOT1 (N75, N55);
xor XOR2 (N76, N62, N1);
and AND3 (N77, N70, N35, N46);
xor XOR2 (N78, N74, N58);
and AND2 (N79, N10, N8);
not NOT1 (N80, N79);
xor XOR2 (N81, N76, N11);
buf BUF1 (N82, N52);
not NOT1 (N83, N64);
xor XOR2 (N84, N72, N49);
and AND3 (N85, N84, N29, N23);
not NOT1 (N86, N80);
not NOT1 (N87, N68);
buf BUF1 (N88, N83);
buf BUF1 (N89, N69);
or OR2 (N90, N87, N53);
nand NAND3 (N91, N82, N38, N48);
and AND4 (N92, N89, N76, N69, N14);
nand NAND3 (N93, N91, N27, N25);
xor XOR2 (N94, N75, N60);
xor XOR2 (N95, N90, N14);
nor NOR2 (N96, N93, N71);
buf BUF1 (N97, N85);
not NOT1 (N98, N96);
xor XOR2 (N99, N97, N96);
buf BUF1 (N100, N81);
and AND3 (N101, N88, N57, N17);
buf BUF1 (N102, N99);
buf BUF1 (N103, N86);
buf BUF1 (N104, N94);
nor NOR2 (N105, N92, N14);
not NOT1 (N106, N95);
nand NAND4 (N107, N100, N30, N60, N85);
xor XOR2 (N108, N105, N88);
and AND2 (N109, N107, N105);
nor NOR2 (N110, N101, N51);
not NOT1 (N111, N108);
nor NOR4 (N112, N106, N31, N53, N31);
or OR4 (N113, N78, N65, N18, N60);
and AND2 (N114, N110, N102);
xor XOR2 (N115, N31, N65);
xor XOR2 (N116, N109, N26);
and AND3 (N117, N114, N30, N77);
nand NAND3 (N118, N52, N65, N30);
and AND3 (N119, N104, N56, N54);
nor NOR4 (N120, N112, N62, N89, N63);
nor NOR4 (N121, N98, N77, N68, N58);
buf BUF1 (N122, N116);
not NOT1 (N123, N111);
buf BUF1 (N124, N113);
xor XOR2 (N125, N121, N79);
buf BUF1 (N126, N117);
buf BUF1 (N127, N103);
nand NAND2 (N128, N123, N38);
and AND4 (N129, N119, N38, N10, N112);
nor NOR2 (N130, N126, N85);
or OR2 (N131, N125, N67);
and AND2 (N132, N118, N35);
xor XOR2 (N133, N122, N39);
buf BUF1 (N134, N129);
nor NOR4 (N135, N133, N107, N52, N11);
nand NAND2 (N136, N115, N24);
nand NAND4 (N137, N134, N103, N127, N6);
nand NAND2 (N138, N91, N77);
nor NOR3 (N139, N128, N77, N16);
or OR4 (N140, N131, N28, N95, N94);
or OR4 (N141, N130, N29, N79, N89);
not NOT1 (N142, N135);
nor NOR4 (N143, N132, N63, N40, N133);
not NOT1 (N144, N142);
and AND2 (N145, N143, N66);
not NOT1 (N146, N140);
not NOT1 (N147, N120);
buf BUF1 (N148, N136);
nor NOR2 (N149, N138, N28);
or OR3 (N150, N141, N15, N104);
or OR3 (N151, N147, N87, N33);
nand NAND2 (N152, N145, N73);
and AND3 (N153, N137, N6, N146);
xor XOR2 (N154, N136, N127);
nor NOR3 (N155, N139, N112, N59);
buf BUF1 (N156, N155);
buf BUF1 (N157, N149);
nand NAND4 (N158, N144, N107, N139, N115);
and AND2 (N159, N156, N45);
or OR3 (N160, N124, N94, N19);
nand NAND2 (N161, N153, N71);
buf BUF1 (N162, N160);
buf BUF1 (N163, N157);
nand NAND4 (N164, N154, N136, N32, N111);
not NOT1 (N165, N162);
nor NOR4 (N166, N151, N125, N108, N139);
and AND3 (N167, N166, N50, N156);
or OR3 (N168, N159, N123, N124);
xor XOR2 (N169, N163, N125);
xor XOR2 (N170, N158, N125);
nand NAND2 (N171, N152, N102);
buf BUF1 (N172, N167);
xor XOR2 (N173, N165, N36);
nand NAND2 (N174, N172, N54);
and AND4 (N175, N164, N135, N34, N101);
or OR2 (N176, N170, N106);
not NOT1 (N177, N148);
buf BUF1 (N178, N168);
nor NOR4 (N179, N175, N158, N166, N102);
not NOT1 (N180, N161);
buf BUF1 (N181, N150);
buf BUF1 (N182, N171);
xor XOR2 (N183, N178, N155);
buf BUF1 (N184, N174);
not NOT1 (N185, N183);
not NOT1 (N186, N179);
and AND4 (N187, N176, N11, N72, N119);
nor NOR4 (N188, N187, N48, N88, N81);
nand NAND2 (N189, N181, N174);
not NOT1 (N190, N186);
xor XOR2 (N191, N182, N144);
nand NAND4 (N192, N191, N151, N5, N124);
and AND3 (N193, N188, N86, N76);
and AND3 (N194, N177, N184, N152);
and AND3 (N195, N73, N96, N120);
and AND2 (N196, N195, N45);
or OR3 (N197, N169, N148, N118);
buf BUF1 (N198, N185);
nand NAND2 (N199, N190, N44);
nor NOR4 (N200, N199, N130, N99, N75);
xor XOR2 (N201, N198, N160);
or OR4 (N202, N180, N102, N75, N145);
not NOT1 (N203, N189);
nand NAND2 (N204, N196, N57);
nor NOR4 (N205, N201, N25, N53, N113);
not NOT1 (N206, N197);
or OR4 (N207, N204, N101, N80, N194);
and AND4 (N208, N106, N171, N52, N150);
nand NAND2 (N209, N202, N41);
nand NAND3 (N210, N200, N36, N141);
nor NOR3 (N211, N193, N85, N49);
or OR2 (N212, N210, N62);
not NOT1 (N213, N192);
buf BUF1 (N214, N209);
nor NOR4 (N215, N212, N174, N100, N56);
or OR3 (N216, N215, N163, N186);
nand NAND2 (N217, N205, N5);
and AND2 (N218, N213, N77);
and AND2 (N219, N214, N129);
buf BUF1 (N220, N206);
nor NOR3 (N221, N218, N205, N189);
buf BUF1 (N222, N217);
not NOT1 (N223, N211);
or OR4 (N224, N203, N156, N111, N158);
buf BUF1 (N225, N221);
not NOT1 (N226, N207);
not NOT1 (N227, N173);
not NOT1 (N228, N225);
and AND3 (N229, N222, N28, N189);
xor XOR2 (N230, N219, N69);
or OR4 (N231, N216, N78, N137, N204);
buf BUF1 (N232, N228);
xor XOR2 (N233, N231, N15);
nor NOR4 (N234, N220, N104, N168, N182);
nand NAND3 (N235, N227, N42, N73);
nand NAND2 (N236, N224, N167);
nor NOR3 (N237, N208, N104, N133);
buf BUF1 (N238, N232);
xor XOR2 (N239, N235, N101);
buf BUF1 (N240, N238);
not NOT1 (N241, N240);
not NOT1 (N242, N229);
nor NOR3 (N243, N241, N54, N16);
and AND2 (N244, N230, N5);
not NOT1 (N245, N233);
not NOT1 (N246, N236);
buf BUF1 (N247, N239);
nor NOR3 (N248, N226, N186, N124);
nor NOR3 (N249, N243, N97, N187);
buf BUF1 (N250, N237);
nand NAND4 (N251, N247, N9, N160, N190);
nand NAND4 (N252, N244, N85, N152, N5);
nand NAND4 (N253, N250, N152, N239, N29);
not NOT1 (N254, N245);
or OR2 (N255, N252, N74);
or OR3 (N256, N255, N16, N23);
not NOT1 (N257, N242);
and AND3 (N258, N249, N40, N31);
not NOT1 (N259, N258);
not NOT1 (N260, N223);
not NOT1 (N261, N253);
xor XOR2 (N262, N257, N258);
or OR3 (N263, N246, N4, N179);
or OR4 (N264, N254, N33, N137, N164);
nand NAND3 (N265, N248, N11, N179);
not NOT1 (N266, N261);
nor NOR3 (N267, N263, N139, N219);
and AND3 (N268, N264, N197, N256);
xor XOR2 (N269, N244, N75);
nand NAND2 (N270, N269, N218);
nand NAND3 (N271, N265, N237, N21);
and AND2 (N272, N260, N137);
or OR3 (N273, N268, N182, N127);
nor NOR4 (N274, N234, N143, N36, N267);
nand NAND4 (N275, N195, N123, N124, N143);
or OR3 (N276, N273, N154, N27);
nor NOR3 (N277, N262, N37, N250);
nor NOR4 (N278, N275, N34, N195, N38);
nor NOR4 (N279, N278, N138, N228, N45);
and AND4 (N280, N266, N209, N236, N152);
nand NAND3 (N281, N276, N111, N261);
not NOT1 (N282, N259);
xor XOR2 (N283, N280, N163);
not NOT1 (N284, N277);
xor XOR2 (N285, N270, N270);
buf BUF1 (N286, N283);
and AND2 (N287, N251, N178);
buf BUF1 (N288, N281);
not NOT1 (N289, N271);
or OR2 (N290, N284, N105);
xor XOR2 (N291, N274, N157);
and AND3 (N292, N291, N100, N182);
or OR4 (N293, N290, N122, N36, N6);
and AND4 (N294, N292, N34, N108, N278);
buf BUF1 (N295, N294);
nand NAND2 (N296, N288, N19);
nand NAND3 (N297, N287, N139, N286);
and AND3 (N298, N217, N117, N189);
nor NOR2 (N299, N279, N92);
nand NAND2 (N300, N298, N255);
nand NAND4 (N301, N300, N239, N56, N196);
nand NAND3 (N302, N293, N285, N260);
not NOT1 (N303, N242);
not NOT1 (N304, N295);
buf BUF1 (N305, N303);
nand NAND4 (N306, N305, N160, N260, N276);
and AND2 (N307, N296, N133);
and AND2 (N308, N306, N84);
not NOT1 (N309, N299);
xor XOR2 (N310, N301, N254);
nor NOR4 (N311, N309, N130, N110, N55);
buf BUF1 (N312, N282);
buf BUF1 (N313, N289);
nor NOR3 (N314, N302, N91, N58);
nor NOR4 (N315, N312, N279, N133, N283);
or OR3 (N316, N310, N42, N20);
nor NOR3 (N317, N311, N186, N188);
xor XOR2 (N318, N304, N55);
and AND2 (N319, N317, N197);
not NOT1 (N320, N314);
nor NOR2 (N321, N318, N254);
or OR2 (N322, N307, N101);
buf BUF1 (N323, N313);
nand NAND3 (N324, N322, N19, N316);
xor XOR2 (N325, N136, N203);
nor NOR2 (N326, N315, N263);
and AND2 (N327, N324, N270);
buf BUF1 (N328, N297);
not NOT1 (N329, N325);
buf BUF1 (N330, N272);
nand NAND4 (N331, N327, N282, N12, N12);
not NOT1 (N332, N308);
and AND4 (N333, N319, N152, N50, N110);
not NOT1 (N334, N333);
or OR2 (N335, N329, N151);
nand NAND4 (N336, N330, N41, N218, N7);
buf BUF1 (N337, N331);
or OR2 (N338, N332, N123);
or OR3 (N339, N320, N13, N334);
nand NAND4 (N340, N30, N169, N271, N112);
buf BUF1 (N341, N323);
nor NOR3 (N342, N321, N338, N43);
nor NOR2 (N343, N341, N129);
not NOT1 (N344, N248);
nand NAND2 (N345, N326, N74);
and AND3 (N346, N335, N96, N25);
nand NAND2 (N347, N342, N221);
nor NOR2 (N348, N339, N250);
or OR4 (N349, N337, N322, N283, N97);
nand NAND3 (N350, N347, N308, N116);
and AND4 (N351, N343, N21, N127, N40);
nand NAND4 (N352, N336, N260, N58, N169);
buf BUF1 (N353, N345);
nand NAND2 (N354, N350, N41);
nand NAND4 (N355, N354, N340, N193, N163);
xor XOR2 (N356, N239, N72);
nand NAND3 (N357, N352, N302, N356);
nand NAND3 (N358, N11, N22, N340);
nor NOR3 (N359, N357, N78, N166);
nor NOR3 (N360, N328, N27, N269);
not NOT1 (N361, N346);
not NOT1 (N362, N344);
and AND2 (N363, N353, N19);
and AND4 (N364, N361, N58, N338, N351);
buf BUF1 (N365, N3);
or OR3 (N366, N348, N275, N221);
and AND2 (N367, N349, N310);
or OR4 (N368, N366, N11, N334, N62);
xor XOR2 (N369, N358, N20);
or OR3 (N370, N360, N178, N320);
buf BUF1 (N371, N364);
not NOT1 (N372, N370);
nor NOR2 (N373, N368, N355);
buf BUF1 (N374, N150);
xor XOR2 (N375, N367, N8);
nand NAND3 (N376, N373, N189, N330);
xor XOR2 (N377, N365, N267);
buf BUF1 (N378, N371);
buf BUF1 (N379, N362);
or OR3 (N380, N363, N191, N97);
nor NOR3 (N381, N380, N185, N219);
nand NAND2 (N382, N359, N48);
and AND3 (N383, N369, N150, N203);
and AND3 (N384, N372, N366, N354);
or OR4 (N385, N379, N162, N241, N341);
nor NOR4 (N386, N384, N35, N122, N266);
not NOT1 (N387, N378);
not NOT1 (N388, N381);
xor XOR2 (N389, N376, N178);
nor NOR2 (N390, N386, N235);
not NOT1 (N391, N390);
and AND2 (N392, N385, N81);
nor NOR2 (N393, N382, N384);
nor NOR2 (N394, N388, N229);
buf BUF1 (N395, N389);
or OR4 (N396, N387, N161, N78, N285);
buf BUF1 (N397, N383);
nor NOR3 (N398, N395, N334, N124);
nand NAND2 (N399, N393, N331);
or OR4 (N400, N397, N191, N212, N9);
nor NOR3 (N401, N400, N84, N102);
buf BUF1 (N402, N375);
xor XOR2 (N403, N399, N108);
buf BUF1 (N404, N394);
nor NOR4 (N405, N404, N64, N241, N151);
nand NAND2 (N406, N391, N397);
buf BUF1 (N407, N403);
nand NAND3 (N408, N374, N167, N218);
nand NAND3 (N409, N401, N174, N122);
xor XOR2 (N410, N392, N234);
xor XOR2 (N411, N402, N106);
buf BUF1 (N412, N409);
nor NOR4 (N413, N406, N234, N296, N337);
xor XOR2 (N414, N408, N381);
and AND3 (N415, N412, N220, N332);
not NOT1 (N416, N405);
and AND2 (N417, N398, N333);
nand NAND3 (N418, N416, N249, N401);
not NOT1 (N419, N377);
xor XOR2 (N420, N414, N62);
buf BUF1 (N421, N407);
nand NAND3 (N422, N418, N263, N96);
buf BUF1 (N423, N421);
or OR2 (N424, N415, N110);
or OR3 (N425, N422, N109, N137);
buf BUF1 (N426, N425);
or OR4 (N427, N419, N176, N129, N19);
nand NAND4 (N428, N424, N83, N54, N94);
xor XOR2 (N429, N413, N423);
not NOT1 (N430, N210);
nor NOR3 (N431, N410, N403, N337);
and AND4 (N432, N429, N302, N3, N363);
xor XOR2 (N433, N427, N327);
nor NOR2 (N434, N433, N354);
xor XOR2 (N435, N396, N412);
nand NAND3 (N436, N411, N107, N195);
nor NOR4 (N437, N436, N38, N292, N303);
nand NAND3 (N438, N420, N392, N231);
buf BUF1 (N439, N428);
nor NOR4 (N440, N434, N6, N311, N175);
and AND2 (N441, N437, N17);
not NOT1 (N442, N426);
or OR3 (N443, N430, N96, N279);
nor NOR2 (N444, N435, N430);
or OR4 (N445, N432, N386, N430, N427);
not NOT1 (N446, N443);
nand NAND2 (N447, N441, N394);
and AND3 (N448, N438, N132, N349);
not NOT1 (N449, N446);
nor NOR4 (N450, N431, N414, N25, N11);
xor XOR2 (N451, N417, N316);
xor XOR2 (N452, N445, N407);
nor NOR2 (N453, N449, N439);
xor XOR2 (N454, N234, N134);
nor NOR4 (N455, N440, N404, N6, N445);
and AND4 (N456, N448, N308, N34, N331);
and AND3 (N457, N442, N146, N287);
buf BUF1 (N458, N456);
nand NAND3 (N459, N447, N169, N56);
xor XOR2 (N460, N459, N73);
or OR3 (N461, N451, N242, N377);
not NOT1 (N462, N454);
xor XOR2 (N463, N457, N48);
and AND4 (N464, N458, N186, N321, N348);
not NOT1 (N465, N460);
xor XOR2 (N466, N453, N29);
nor NOR4 (N467, N461, N434, N233, N444);
xor XOR2 (N468, N126, N412);
nand NAND4 (N469, N452, N146, N375, N245);
xor XOR2 (N470, N464, N192);
nand NAND3 (N471, N466, N352, N49);
or OR3 (N472, N467, N431, N35);
nor NOR4 (N473, N471, N174, N469, N328);
not NOT1 (N474, N221);
xor XOR2 (N475, N474, N139);
not NOT1 (N476, N470);
nor NOR3 (N477, N450, N224, N440);
not NOT1 (N478, N473);
not NOT1 (N479, N468);
or OR2 (N480, N465, N454);
and AND2 (N481, N472, N207);
xor XOR2 (N482, N463, N60);
buf BUF1 (N483, N475);
not NOT1 (N484, N455);
nor NOR2 (N485, N478, N477);
nand NAND3 (N486, N310, N141, N378);
nor NOR4 (N487, N479, N324, N424, N428);
and AND2 (N488, N483, N429);
nor NOR2 (N489, N481, N208);
buf BUF1 (N490, N482);
buf BUF1 (N491, N490);
nor NOR4 (N492, N488, N115, N89, N419);
xor XOR2 (N493, N476, N356);
xor XOR2 (N494, N484, N434);
and AND4 (N495, N485, N417, N101, N82);
not NOT1 (N496, N491);
nor NOR4 (N497, N496, N433, N425, N50);
xor XOR2 (N498, N489, N264);
or OR4 (N499, N462, N268, N369, N319);
not NOT1 (N500, N499);
and AND2 (N501, N495, N107);
nand NAND3 (N502, N480, N186, N34);
and AND4 (N503, N502, N36, N255, N79);
not NOT1 (N504, N486);
buf BUF1 (N505, N500);
buf BUF1 (N506, N492);
nor NOR2 (N507, N487, N463);
not NOT1 (N508, N498);
nor NOR4 (N509, N508, N408, N346, N307);
xor XOR2 (N510, N509, N246);
nor NOR4 (N511, N507, N427, N243, N484);
and AND2 (N512, N511, N97);
and AND4 (N513, N501, N270, N111, N314);
and AND2 (N514, N504, N398);
nor NOR3 (N515, N506, N354, N80);
or OR2 (N516, N505, N45);
and AND4 (N517, N494, N372, N267, N269);
nand NAND2 (N518, N503, N206);
buf BUF1 (N519, N518);
nor NOR4 (N520, N512, N214, N31, N261);
nor NOR4 (N521, N514, N138, N347, N430);
or OR4 (N522, N510, N377, N424, N167);
and AND2 (N523, N519, N347);
and AND4 (N524, N515, N136, N126, N98);
buf BUF1 (N525, N497);
nor NOR2 (N526, N520, N448);
nand NAND4 (N527, N526, N450, N469, N430);
nand NAND2 (N528, N523, N22);
xor XOR2 (N529, N527, N372);
xor XOR2 (N530, N516, N383);
xor XOR2 (N531, N530, N207);
nor NOR4 (N532, N528, N349, N107, N198);
nand NAND2 (N533, N525, N104);
and AND4 (N534, N513, N350, N158, N143);
nand NAND2 (N535, N532, N408);
or OR4 (N536, N521, N8, N506, N181);
or OR4 (N537, N535, N512, N283, N511);
or OR2 (N538, N493, N279);
or OR3 (N539, N524, N47, N405);
not NOT1 (N540, N537);
nand NAND2 (N541, N533, N121);
nand NAND4 (N542, N517, N341, N262, N129);
nand NAND2 (N543, N536, N374);
not NOT1 (N544, N522);
nor NOR2 (N545, N542, N333);
nor NOR3 (N546, N544, N487, N177);
not NOT1 (N547, N545);
xor XOR2 (N548, N543, N16);
nor NOR3 (N549, N539, N52, N103);
nand NAND2 (N550, N547, N6);
xor XOR2 (N551, N534, N523);
buf BUF1 (N552, N548);
or OR3 (N553, N529, N104, N315);
nor NOR2 (N554, N531, N128);
nand NAND2 (N555, N550, N224);
and AND2 (N556, N541, N341);
buf BUF1 (N557, N540);
and AND2 (N558, N538, N482);
or OR3 (N559, N558, N40, N162);
buf BUF1 (N560, N555);
or OR2 (N561, N551, N138);
xor XOR2 (N562, N561, N409);
xor XOR2 (N563, N560, N224);
and AND4 (N564, N554, N275, N560, N87);
not NOT1 (N565, N552);
xor XOR2 (N566, N549, N37);
xor XOR2 (N567, N553, N111);
not NOT1 (N568, N567);
xor XOR2 (N569, N557, N545);
xor XOR2 (N570, N569, N423);
nand NAND3 (N571, N559, N519, N291);
or OR3 (N572, N568, N399, N235);
buf BUF1 (N573, N556);
or OR3 (N574, N564, N238, N152);
and AND3 (N575, N572, N390, N37);
xor XOR2 (N576, N563, N431);
xor XOR2 (N577, N546, N569);
xor XOR2 (N578, N577, N256);
not NOT1 (N579, N566);
and AND4 (N580, N570, N531, N359, N361);
nand NAND3 (N581, N574, N172, N507);
and AND3 (N582, N576, N127, N494);
buf BUF1 (N583, N575);
and AND3 (N584, N581, N221, N214);
not NOT1 (N585, N571);
not NOT1 (N586, N580);
and AND4 (N587, N578, N125, N552, N87);
xor XOR2 (N588, N586, N432);
or OR2 (N589, N579, N319);
xor XOR2 (N590, N589, N109);
and AND3 (N591, N584, N194, N122);
buf BUF1 (N592, N573);
xor XOR2 (N593, N590, N235);
nand NAND3 (N594, N583, N229, N106);
xor XOR2 (N595, N562, N584);
or OR2 (N596, N565, N139);
xor XOR2 (N597, N587, N345);
buf BUF1 (N598, N592);
nand NAND4 (N599, N596, N471, N541, N4);
buf BUF1 (N600, N588);
not NOT1 (N601, N585);
nor NOR4 (N602, N598, N71, N431, N496);
and AND3 (N603, N599, N2, N132);
not NOT1 (N604, N602);
and AND3 (N605, N604, N49, N132);
xor XOR2 (N606, N595, N203);
and AND4 (N607, N593, N379, N64, N61);
and AND2 (N608, N607, N115);
nand NAND4 (N609, N600, N581, N323, N280);
xor XOR2 (N610, N601, N418);
and AND4 (N611, N591, N215, N56, N117);
and AND2 (N612, N609, N142);
xor XOR2 (N613, N606, N336);
nor NOR3 (N614, N612, N188, N563);
or OR3 (N615, N603, N422, N570);
or OR2 (N616, N614, N533);
and AND3 (N617, N605, N441, N137);
nand NAND2 (N618, N616, N374);
nand NAND3 (N619, N594, N22, N431);
buf BUF1 (N620, N618);
buf BUF1 (N621, N620);
nand NAND4 (N622, N621, N544, N361, N562);
not NOT1 (N623, N615);
nand NAND3 (N624, N622, N340, N576);
or OR4 (N625, N597, N609, N253, N530);
xor XOR2 (N626, N617, N332);
buf BUF1 (N627, N613);
and AND2 (N628, N619, N528);
xor XOR2 (N629, N624, N467);
nor NOR4 (N630, N628, N152, N39, N189);
or OR3 (N631, N608, N498, N245);
nor NOR4 (N632, N623, N227, N557, N89);
nand NAND3 (N633, N629, N501, N261);
or OR3 (N634, N625, N121, N64);
nand NAND4 (N635, N633, N523, N215, N17);
not NOT1 (N636, N632);
nand NAND4 (N637, N627, N402, N135, N380);
nand NAND3 (N638, N582, N357, N621);
xor XOR2 (N639, N636, N585);
nand NAND2 (N640, N637, N194);
not NOT1 (N641, N630);
not NOT1 (N642, N634);
nand NAND3 (N643, N631, N216, N24);
or OR4 (N644, N611, N18, N48, N181);
or OR4 (N645, N635, N475, N555, N204);
nand NAND3 (N646, N642, N490, N443);
and AND3 (N647, N640, N308, N507);
not NOT1 (N648, N639);
nand NAND4 (N649, N626, N49, N367, N584);
nor NOR3 (N650, N649, N363, N566);
nor NOR2 (N651, N647, N564);
nand NAND4 (N652, N644, N338, N522, N505);
buf BUF1 (N653, N641);
nor NOR2 (N654, N643, N190);
nor NOR4 (N655, N648, N28, N98, N142);
buf BUF1 (N656, N610);
xor XOR2 (N657, N650, N122);
or OR2 (N658, N655, N432);
buf BUF1 (N659, N638);
not NOT1 (N660, N654);
not NOT1 (N661, N645);
nand NAND4 (N662, N660, N352, N257, N146);
not NOT1 (N663, N656);
nor NOR3 (N664, N659, N513, N377);
xor XOR2 (N665, N663, N108);
or OR3 (N666, N658, N632, N605);
nor NOR2 (N667, N662, N625);
nor NOR3 (N668, N651, N61, N620);
buf BUF1 (N669, N653);
xor XOR2 (N670, N667, N28);
or OR4 (N671, N666, N254, N581, N24);
nor NOR4 (N672, N669, N405, N630, N306);
not NOT1 (N673, N664);
not NOT1 (N674, N671);
or OR4 (N675, N670, N129, N541, N197);
xor XOR2 (N676, N668, N414);
nand NAND3 (N677, N661, N585, N199);
buf BUF1 (N678, N674);
xor XOR2 (N679, N652, N276);
not NOT1 (N680, N679);
and AND4 (N681, N678, N634, N584, N338);
nor NOR4 (N682, N665, N105, N399, N332);
or OR2 (N683, N682, N273);
buf BUF1 (N684, N681);
xor XOR2 (N685, N672, N282);
and AND3 (N686, N675, N337, N77);
xor XOR2 (N687, N680, N81);
nand NAND3 (N688, N676, N305, N485);
not NOT1 (N689, N688);
buf BUF1 (N690, N646);
nand NAND4 (N691, N686, N645, N334, N154);
nor NOR3 (N692, N657, N471, N243);
not NOT1 (N693, N687);
buf BUF1 (N694, N673);
not NOT1 (N695, N677);
buf BUF1 (N696, N684);
or OR4 (N697, N693, N199, N390, N120);
buf BUF1 (N698, N685);
or OR2 (N699, N695, N689);
or OR4 (N700, N41, N629, N108, N692);
xor XOR2 (N701, N427, N82);
and AND2 (N702, N683, N591);
or OR3 (N703, N691, N154, N490);
and AND2 (N704, N703, N432);
not NOT1 (N705, N696);
and AND2 (N706, N705, N214);
and AND3 (N707, N706, N259, N225);
buf BUF1 (N708, N698);
not NOT1 (N709, N700);
and AND3 (N710, N707, N471, N133);
xor XOR2 (N711, N699, N685);
or OR4 (N712, N704, N381, N276, N424);
nor NOR2 (N713, N701, N344);
nor NOR2 (N714, N708, N675);
nand NAND4 (N715, N709, N366, N233, N292);
xor XOR2 (N716, N690, N516);
nand NAND3 (N717, N697, N58, N298);
or OR3 (N718, N714, N370, N436);
nor NOR4 (N719, N702, N127, N411, N167);
nand NAND3 (N720, N712, N445, N405);
nand NAND2 (N721, N710, N600);
nor NOR3 (N722, N694, N234, N695);
not NOT1 (N723, N722);
or OR4 (N724, N711, N397, N117, N449);
and AND3 (N725, N716, N195, N204);
and AND4 (N726, N717, N333, N80, N242);
xor XOR2 (N727, N720, N594);
not NOT1 (N728, N719);
nor NOR3 (N729, N723, N342, N461);
not NOT1 (N730, N727);
or OR2 (N731, N728, N572);
not NOT1 (N732, N721);
nor NOR2 (N733, N726, N365);
or OR2 (N734, N733, N421);
nand NAND2 (N735, N734, N154);
not NOT1 (N736, N735);
nand NAND3 (N737, N718, N726, N369);
or OR4 (N738, N729, N75, N369, N234);
nand NAND4 (N739, N732, N42, N208, N39);
and AND4 (N740, N725, N442, N369, N581);
nand NAND3 (N741, N724, N172, N624);
or OR2 (N742, N731, N25);
xor XOR2 (N743, N738, N728);
nor NOR3 (N744, N743, N582, N485);
or OR2 (N745, N730, N719);
buf BUF1 (N746, N740);
and AND4 (N747, N713, N138, N614, N548);
xor XOR2 (N748, N744, N194);
nand NAND2 (N749, N736, N177);
or OR2 (N750, N741, N436);
not NOT1 (N751, N745);
buf BUF1 (N752, N751);
not NOT1 (N753, N749);
not NOT1 (N754, N715);
buf BUF1 (N755, N748);
or OR4 (N756, N739, N55, N485, N287);
not NOT1 (N757, N747);
buf BUF1 (N758, N753);
nor NOR4 (N759, N750, N382, N130, N206);
or OR4 (N760, N758, N158, N687, N364);
buf BUF1 (N761, N757);
nor NOR2 (N762, N742, N218);
not NOT1 (N763, N746);
xor XOR2 (N764, N763, N651);
nor NOR3 (N765, N752, N405, N445);
or OR4 (N766, N762, N429, N595, N34);
nor NOR4 (N767, N756, N720, N97, N618);
nand NAND4 (N768, N766, N315, N767, N142);
or OR2 (N769, N649, N320);
nand NAND3 (N770, N760, N438, N268);
nand NAND2 (N771, N759, N622);
nor NOR4 (N772, N768, N284, N766, N565);
or OR3 (N773, N755, N529, N45);
nand NAND4 (N774, N765, N441, N513, N80);
buf BUF1 (N775, N769);
buf BUF1 (N776, N772);
xor XOR2 (N777, N771, N482);
xor XOR2 (N778, N754, N515);
xor XOR2 (N779, N761, N543);
nand NAND4 (N780, N775, N113, N243, N639);
buf BUF1 (N781, N764);
nand NAND4 (N782, N774, N465, N391, N657);
buf BUF1 (N783, N773);
nor NOR3 (N784, N782, N617, N363);
nor NOR3 (N785, N779, N742, N233);
nand NAND2 (N786, N783, N386);
xor XOR2 (N787, N786, N784);
buf BUF1 (N788, N59);
nand NAND2 (N789, N787, N645);
nand NAND3 (N790, N781, N691, N484);
or OR4 (N791, N776, N750, N517, N422);
not NOT1 (N792, N789);
nand NAND2 (N793, N791, N428);
xor XOR2 (N794, N785, N641);
xor XOR2 (N795, N778, N78);
xor XOR2 (N796, N780, N340);
nand NAND4 (N797, N737, N245, N262, N438);
not NOT1 (N798, N770);
and AND3 (N799, N793, N176, N584);
not NOT1 (N800, N797);
nand NAND2 (N801, N794, N236);
nor NOR4 (N802, N795, N235, N223, N253);
and AND4 (N803, N800, N46, N682, N527);
nand NAND2 (N804, N788, N125);
or OR4 (N805, N803, N611, N327, N482);
nand NAND2 (N806, N777, N95);
xor XOR2 (N807, N790, N206);
xor XOR2 (N808, N805, N322);
not NOT1 (N809, N801);
xor XOR2 (N810, N798, N765);
or OR2 (N811, N804, N672);
nor NOR3 (N812, N806, N589, N811);
buf BUF1 (N813, N676);
endmodule