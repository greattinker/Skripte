// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13;

output N611,N609,N610,N600,N597,N612,N588,N603,N602,N613;

nand NAND4 (N14, N11, N1, N12, N8);
nor NOR2 (N15, N9, N12);
not NOT1 (N16, N7);
and AND2 (N17, N10, N3);
xor XOR2 (N18, N5, N7);
buf BUF1 (N19, N12);
nand NAND4 (N20, N1, N9, N6, N13);
xor XOR2 (N21, N15, N16);
nor NOR3 (N22, N11, N16, N11);
buf BUF1 (N23, N16);
and AND4 (N24, N15, N16, N6, N19);
and AND2 (N25, N20, N19);
or OR2 (N26, N7, N24);
xor XOR2 (N27, N19, N18);
nand NAND2 (N28, N5, N15);
not NOT1 (N29, N7);
or OR3 (N30, N22, N3, N18);
or OR2 (N31, N25, N22);
buf BUF1 (N32, N26);
nor NOR4 (N33, N14, N21, N7, N27);
not NOT1 (N34, N5);
and AND3 (N35, N5, N27, N21);
xor XOR2 (N36, N29, N32);
buf BUF1 (N37, N18);
not NOT1 (N38, N31);
not NOT1 (N39, N23);
nand NAND2 (N40, N28, N14);
buf BUF1 (N41, N34);
or OR2 (N42, N38, N37);
nand NAND2 (N43, N9, N9);
or OR2 (N44, N36, N22);
not NOT1 (N45, N44);
nor NOR3 (N46, N41, N2, N39);
nor NOR4 (N47, N40, N44, N6, N44);
buf BUF1 (N48, N20);
and AND3 (N49, N47, N17, N35);
nor NOR3 (N50, N45, N16, N46);
nand NAND3 (N51, N18, N7, N24);
nand NAND3 (N52, N4, N21, N25);
not NOT1 (N53, N3);
not NOT1 (N54, N53);
and AND3 (N55, N48, N25, N3);
xor XOR2 (N56, N51, N32);
or OR4 (N57, N49, N3, N17, N24);
buf BUF1 (N58, N30);
xor XOR2 (N59, N57, N5);
xor XOR2 (N60, N58, N35);
and AND3 (N61, N33, N60, N60);
not NOT1 (N62, N11);
and AND3 (N63, N54, N16, N37);
nor NOR4 (N64, N43, N9, N46, N58);
nor NOR4 (N65, N52, N30, N62, N27);
buf BUF1 (N66, N10);
nor NOR2 (N67, N59, N45);
or OR3 (N68, N66, N2, N2);
or OR2 (N69, N50, N7);
nor NOR3 (N70, N42, N35, N45);
xor XOR2 (N71, N68, N23);
or OR2 (N72, N65, N23);
and AND4 (N73, N67, N49, N46, N21);
xor XOR2 (N74, N64, N29);
nor NOR2 (N75, N73, N42);
not NOT1 (N76, N69);
nor NOR2 (N77, N71, N63);
nand NAND3 (N78, N50, N22, N24);
and AND2 (N79, N55, N64);
and AND4 (N80, N61, N42, N79, N20);
xor XOR2 (N81, N53, N77);
buf BUF1 (N82, N79);
or OR4 (N83, N81, N61, N43, N14);
nor NOR4 (N84, N74, N70, N20, N53);
not NOT1 (N85, N38);
and AND4 (N86, N84, N69, N28, N85);
nand NAND4 (N87, N23, N44, N33, N65);
buf BUF1 (N88, N78);
nand NAND3 (N89, N80, N78, N72);
nand NAND3 (N90, N47, N27, N79);
and AND4 (N91, N87, N59, N75, N37);
or OR2 (N92, N70, N80);
nand NAND3 (N93, N88, N85, N82);
xor XOR2 (N94, N38, N76);
and AND3 (N95, N3, N13, N85);
nand NAND4 (N96, N89, N20, N25, N7);
nand NAND3 (N97, N95, N4, N51);
nand NAND4 (N98, N96, N21, N5, N4);
or OR3 (N99, N92, N90, N60);
xor XOR2 (N100, N50, N54);
nor NOR4 (N101, N91, N7, N27, N94);
nor NOR4 (N102, N12, N89, N67, N53);
and AND4 (N103, N100, N11, N76, N97);
buf BUF1 (N104, N26);
nand NAND2 (N105, N102, N70);
or OR2 (N106, N101, N86);
not NOT1 (N107, N18);
not NOT1 (N108, N99);
or OR2 (N109, N104, N62);
xor XOR2 (N110, N107, N12);
and AND3 (N111, N93, N61, N81);
not NOT1 (N112, N83);
nor NOR4 (N113, N105, N60, N29, N2);
xor XOR2 (N114, N113, N42);
and AND2 (N115, N103, N7);
nand NAND2 (N116, N98, N78);
and AND2 (N117, N111, N4);
xor XOR2 (N118, N116, N34);
or OR4 (N119, N117, N75, N70, N108);
xor XOR2 (N120, N59, N38);
buf BUF1 (N121, N110);
xor XOR2 (N122, N120, N111);
not NOT1 (N123, N112);
buf BUF1 (N124, N106);
nor NOR3 (N125, N119, N64, N85);
not NOT1 (N126, N122);
xor XOR2 (N127, N126, N39);
xor XOR2 (N128, N115, N85);
buf BUF1 (N129, N109);
nand NAND4 (N130, N114, N38, N35, N18);
or OR3 (N131, N125, N13, N118);
and AND3 (N132, N20, N103, N110);
not NOT1 (N133, N127);
buf BUF1 (N134, N123);
not NOT1 (N135, N131);
or OR2 (N136, N135, N36);
not NOT1 (N137, N136);
nor NOR4 (N138, N56, N123, N25, N80);
nand NAND2 (N139, N134, N38);
nand NAND3 (N140, N130, N19, N9);
buf BUF1 (N141, N124);
or OR2 (N142, N132, N67);
not NOT1 (N143, N142);
xor XOR2 (N144, N143, N46);
xor XOR2 (N145, N144, N99);
and AND3 (N146, N128, N71, N117);
or OR3 (N147, N140, N85, N127);
nand NAND3 (N148, N137, N76, N7);
and AND3 (N149, N141, N1, N90);
xor XOR2 (N150, N121, N39);
xor XOR2 (N151, N138, N85);
not NOT1 (N152, N147);
or OR4 (N153, N150, N127, N18, N135);
and AND3 (N154, N149, N83, N30);
nand NAND4 (N155, N146, N34, N44, N68);
xor XOR2 (N156, N153, N83);
and AND2 (N157, N151, N147);
or OR2 (N158, N133, N43);
or OR2 (N159, N152, N135);
nor NOR4 (N160, N157, N59, N85, N89);
xor XOR2 (N161, N158, N137);
and AND4 (N162, N139, N99, N23, N52);
and AND2 (N163, N154, N78);
nand NAND3 (N164, N160, N59, N59);
nand NAND4 (N165, N162, N29, N76, N40);
not NOT1 (N166, N156);
nor NOR4 (N167, N163, N133, N59, N88);
buf BUF1 (N168, N148);
nor NOR3 (N169, N129, N124, N16);
xor XOR2 (N170, N159, N167);
or OR2 (N171, N12, N77);
xor XOR2 (N172, N164, N153);
buf BUF1 (N173, N166);
nand NAND4 (N174, N169, N90, N94, N47);
buf BUF1 (N175, N161);
or OR2 (N176, N174, N111);
nor NOR2 (N177, N171, N40);
buf BUF1 (N178, N176);
xor XOR2 (N179, N168, N71);
nor NOR2 (N180, N173, N76);
buf BUF1 (N181, N177);
and AND2 (N182, N179, N94);
not NOT1 (N183, N178);
xor XOR2 (N184, N165, N143);
xor XOR2 (N185, N175, N112);
nand NAND3 (N186, N184, N53, N75);
nor NOR2 (N187, N145, N34);
or OR2 (N188, N186, N101);
nor NOR2 (N189, N188, N2);
or OR4 (N190, N189, N169, N103, N80);
or OR2 (N191, N170, N144);
nor NOR4 (N192, N183, N187, N180, N174);
buf BUF1 (N193, N15);
nor NOR2 (N194, N83, N171);
and AND3 (N195, N191, N127, N27);
nand NAND3 (N196, N193, N194, N149);
nor NOR3 (N197, N81, N76, N185);
buf BUF1 (N198, N101);
not NOT1 (N199, N181);
buf BUF1 (N200, N172);
nand NAND2 (N201, N197, N63);
and AND4 (N202, N190, N89, N151, N183);
not NOT1 (N203, N155);
not NOT1 (N204, N198);
nor NOR2 (N205, N199, N144);
nor NOR3 (N206, N200, N152, N28);
xor XOR2 (N207, N204, N47);
nand NAND4 (N208, N205, N60, N69, N31);
buf BUF1 (N209, N196);
nor NOR4 (N210, N209, N166, N110, N83);
not NOT1 (N211, N208);
and AND2 (N212, N195, N159);
xor XOR2 (N213, N206, N165);
buf BUF1 (N214, N213);
or OR4 (N215, N202, N60, N202, N205);
and AND3 (N216, N211, N107, N125);
nand NAND3 (N217, N210, N60, N92);
and AND4 (N218, N201, N39, N86, N213);
and AND4 (N219, N203, N138, N175, N150);
xor XOR2 (N220, N219, N146);
xor XOR2 (N221, N218, N182);
not NOT1 (N222, N104);
or OR3 (N223, N207, N121, N95);
not NOT1 (N224, N214);
xor XOR2 (N225, N221, N143);
buf BUF1 (N226, N212);
nand NAND4 (N227, N222, N117, N129, N53);
or OR2 (N228, N220, N207);
not NOT1 (N229, N217);
or OR2 (N230, N223, N229);
and AND2 (N231, N229, N108);
xor XOR2 (N232, N228, N147);
and AND3 (N233, N225, N218, N223);
xor XOR2 (N234, N216, N157);
buf BUF1 (N235, N230);
and AND2 (N236, N233, N20);
and AND4 (N237, N192, N234, N179, N1);
xor XOR2 (N238, N186, N218);
or OR3 (N239, N235, N140, N165);
or OR4 (N240, N215, N111, N213, N198);
xor XOR2 (N241, N227, N70);
buf BUF1 (N242, N224);
and AND2 (N243, N231, N82);
nand NAND4 (N244, N238, N186, N103, N31);
nor NOR3 (N245, N237, N169, N182);
or OR4 (N246, N245, N205, N146, N44);
not NOT1 (N247, N236);
xor XOR2 (N248, N226, N48);
or OR4 (N249, N244, N31, N194, N175);
nand NAND3 (N250, N232, N20, N128);
and AND4 (N251, N241, N19, N46, N84);
or OR3 (N252, N249, N195, N182);
or OR3 (N253, N250, N117, N87);
nand NAND2 (N254, N253, N195);
xor XOR2 (N255, N251, N218);
nand NAND2 (N256, N239, N109);
buf BUF1 (N257, N243);
and AND2 (N258, N254, N235);
xor XOR2 (N259, N257, N7);
nor NOR3 (N260, N256, N204, N199);
nor NOR2 (N261, N255, N82);
nor NOR3 (N262, N247, N66, N139);
nand NAND2 (N263, N246, N133);
xor XOR2 (N264, N248, N143);
nor NOR3 (N265, N260, N115, N169);
nor NOR2 (N266, N265, N25);
and AND3 (N267, N266, N266, N113);
nor NOR4 (N268, N263, N147, N211, N135);
not NOT1 (N269, N264);
xor XOR2 (N270, N262, N138);
nor NOR4 (N271, N269, N173, N173, N108);
and AND2 (N272, N271, N226);
and AND3 (N273, N272, N151, N226);
nor NOR3 (N274, N242, N97, N102);
or OR3 (N275, N258, N43, N191);
nand NAND3 (N276, N259, N114, N57);
nor NOR4 (N277, N268, N64, N130, N165);
and AND3 (N278, N277, N161, N82);
xor XOR2 (N279, N276, N145);
nand NAND2 (N280, N279, N185);
nor NOR3 (N281, N240, N147, N43);
xor XOR2 (N282, N275, N41);
buf BUF1 (N283, N280);
not NOT1 (N284, N267);
xor XOR2 (N285, N270, N87);
xor XOR2 (N286, N283, N155);
nand NAND4 (N287, N285, N209, N26, N234);
or OR4 (N288, N284, N140, N153, N264);
or OR2 (N289, N287, N7);
and AND3 (N290, N274, N286, N192);
not NOT1 (N291, N60);
nor NOR2 (N292, N290, N8);
nand NAND3 (N293, N252, N193, N52);
and AND4 (N294, N289, N289, N109, N254);
nor NOR2 (N295, N292, N124);
and AND3 (N296, N291, N229, N13);
or OR2 (N297, N296, N100);
not NOT1 (N298, N278);
nor NOR2 (N299, N282, N37);
and AND2 (N300, N294, N214);
not NOT1 (N301, N298);
or OR3 (N302, N288, N53, N244);
and AND4 (N303, N300, N85, N90, N35);
nor NOR4 (N304, N303, N157, N102, N149);
nor NOR2 (N305, N273, N27);
or OR3 (N306, N302, N221, N91);
and AND3 (N307, N261, N142, N170);
buf BUF1 (N308, N306);
nor NOR4 (N309, N281, N68, N128, N218);
or OR4 (N310, N305, N63, N95, N22);
buf BUF1 (N311, N310);
and AND2 (N312, N304, N188);
buf BUF1 (N313, N295);
nand NAND2 (N314, N293, N124);
and AND2 (N315, N313, N308);
and AND2 (N316, N73, N45);
not NOT1 (N317, N316);
nor NOR2 (N318, N317, N23);
buf BUF1 (N319, N301);
or OR4 (N320, N319, N203, N125, N50);
nor NOR2 (N321, N309, N15);
xor XOR2 (N322, N307, N154);
nor NOR3 (N323, N318, N306, N289);
or OR2 (N324, N314, N41);
nand NAND3 (N325, N311, N92, N290);
nand NAND3 (N326, N321, N267, N91);
nor NOR4 (N327, N299, N157, N193, N203);
nand NAND2 (N328, N323, N54);
nand NAND2 (N329, N328, N107);
not NOT1 (N330, N326);
nor NOR3 (N331, N322, N157, N298);
buf BUF1 (N332, N320);
or OR4 (N333, N327, N64, N192, N219);
buf BUF1 (N334, N332);
nand NAND2 (N335, N333, N30);
xor XOR2 (N336, N315, N12);
xor XOR2 (N337, N330, N291);
nand NAND2 (N338, N336, N184);
and AND4 (N339, N337, N141, N4, N165);
or OR2 (N340, N331, N151);
xor XOR2 (N341, N338, N212);
or OR4 (N342, N324, N215, N241, N162);
not NOT1 (N343, N334);
nor NOR3 (N344, N341, N288, N201);
nor NOR3 (N345, N312, N313, N167);
buf BUF1 (N346, N345);
not NOT1 (N347, N325);
not NOT1 (N348, N343);
or OR2 (N349, N342, N210);
or OR3 (N350, N329, N292, N328);
and AND4 (N351, N340, N129, N157, N25);
nand NAND3 (N352, N339, N274, N148);
buf BUF1 (N353, N335);
or OR3 (N354, N346, N10, N215);
or OR3 (N355, N348, N150, N64);
and AND3 (N356, N354, N34, N125);
not NOT1 (N357, N350);
nor NOR4 (N358, N356, N289, N171, N6);
buf BUF1 (N359, N352);
buf BUF1 (N360, N344);
nor NOR2 (N361, N351, N104);
buf BUF1 (N362, N357);
nor NOR4 (N363, N347, N78, N2, N127);
xor XOR2 (N364, N297, N307);
buf BUF1 (N365, N355);
nand NAND3 (N366, N361, N283, N68);
not NOT1 (N367, N353);
buf BUF1 (N368, N360);
nor NOR2 (N369, N363, N263);
buf BUF1 (N370, N358);
xor XOR2 (N371, N365, N273);
or OR3 (N372, N371, N85, N362);
and AND3 (N373, N149, N33, N372);
nand NAND4 (N374, N35, N108, N267, N315);
buf BUF1 (N375, N364);
xor XOR2 (N376, N359, N32);
and AND3 (N377, N366, N113, N296);
nand NAND3 (N378, N375, N314, N39);
nor NOR4 (N379, N367, N349, N185, N148);
and AND3 (N380, N86, N365, N74);
or OR4 (N381, N373, N262, N127, N378);
xor XOR2 (N382, N32, N362);
not NOT1 (N383, N369);
xor XOR2 (N384, N377, N324);
xor XOR2 (N385, N368, N252);
xor XOR2 (N386, N374, N268);
nand NAND3 (N387, N379, N113, N198);
and AND4 (N388, N381, N306, N184, N313);
xor XOR2 (N389, N380, N265);
buf BUF1 (N390, N370);
nand NAND3 (N391, N387, N63, N86);
nor NOR2 (N392, N384, N379);
nand NAND2 (N393, N392, N70);
nor NOR3 (N394, N388, N6, N255);
nand NAND4 (N395, N390, N27, N290, N369);
nor NOR3 (N396, N386, N135, N276);
not NOT1 (N397, N389);
not NOT1 (N398, N382);
buf BUF1 (N399, N393);
not NOT1 (N400, N398);
buf BUF1 (N401, N391);
buf BUF1 (N402, N376);
not NOT1 (N403, N401);
buf BUF1 (N404, N394);
and AND2 (N405, N397, N400);
nand NAND2 (N406, N313, N378);
xor XOR2 (N407, N396, N84);
not NOT1 (N408, N402);
or OR3 (N409, N385, N245, N2);
nand NAND3 (N410, N409, N334, N364);
not NOT1 (N411, N395);
and AND4 (N412, N407, N242, N288, N268);
or OR4 (N413, N404, N84, N53, N41);
not NOT1 (N414, N406);
or OR3 (N415, N403, N193, N303);
and AND3 (N416, N414, N179, N169);
nor NOR3 (N417, N415, N411, N200);
and AND3 (N418, N1, N55, N112);
xor XOR2 (N419, N416, N179);
or OR4 (N420, N405, N25, N240, N361);
xor XOR2 (N421, N408, N89);
and AND2 (N422, N410, N254);
buf BUF1 (N423, N418);
and AND2 (N424, N421, N130);
nand NAND2 (N425, N423, N290);
buf BUF1 (N426, N417);
nor NOR3 (N427, N420, N393, N394);
buf BUF1 (N428, N425);
not NOT1 (N429, N424);
or OR3 (N430, N419, N235, N376);
or OR2 (N431, N428, N254);
xor XOR2 (N432, N429, N391);
xor XOR2 (N433, N426, N156);
or OR4 (N434, N427, N59, N360, N252);
nand NAND3 (N435, N413, N269, N95);
nand NAND3 (N436, N422, N247, N72);
buf BUF1 (N437, N433);
buf BUF1 (N438, N436);
xor XOR2 (N439, N434, N273);
nand NAND2 (N440, N412, N337);
xor XOR2 (N441, N435, N220);
and AND2 (N442, N439, N101);
xor XOR2 (N443, N437, N258);
and AND2 (N444, N399, N274);
nand NAND2 (N445, N431, N55);
xor XOR2 (N446, N442, N9);
nor NOR4 (N447, N445, N24, N9, N410);
xor XOR2 (N448, N443, N294);
and AND4 (N449, N441, N34, N351, N86);
and AND2 (N450, N383, N157);
xor XOR2 (N451, N450, N130);
and AND4 (N452, N449, N356, N400, N443);
nand NAND2 (N453, N440, N305);
and AND2 (N454, N430, N42);
xor XOR2 (N455, N444, N247);
xor XOR2 (N456, N454, N173);
nand NAND3 (N457, N447, N71, N394);
not NOT1 (N458, N432);
or OR2 (N459, N438, N24);
and AND3 (N460, N453, N101, N7);
xor XOR2 (N461, N456, N401);
not NOT1 (N462, N452);
xor XOR2 (N463, N458, N347);
nand NAND2 (N464, N451, N382);
not NOT1 (N465, N457);
nor NOR2 (N466, N448, N187);
or OR4 (N467, N462, N92, N126, N420);
and AND3 (N468, N464, N219, N211);
and AND2 (N469, N446, N202);
not NOT1 (N470, N461);
nand NAND4 (N471, N459, N118, N288, N200);
not NOT1 (N472, N455);
xor XOR2 (N473, N469, N106);
nor NOR3 (N474, N463, N143, N106);
or OR3 (N475, N474, N233, N32);
and AND2 (N476, N473, N199);
not NOT1 (N477, N460);
nand NAND4 (N478, N468, N305, N340, N322);
and AND2 (N479, N472, N211);
xor XOR2 (N480, N470, N346);
or OR2 (N481, N478, N115);
or OR2 (N482, N479, N154);
nand NAND3 (N483, N475, N189, N478);
not NOT1 (N484, N471);
buf BUF1 (N485, N467);
not NOT1 (N486, N485);
xor XOR2 (N487, N484, N182);
nor NOR3 (N488, N487, N208, N75);
xor XOR2 (N489, N482, N19);
nor NOR4 (N490, N483, N319, N70, N26);
not NOT1 (N491, N466);
not NOT1 (N492, N490);
buf BUF1 (N493, N476);
or OR2 (N494, N477, N31);
and AND3 (N495, N489, N303, N366);
or OR4 (N496, N492, N465, N294, N263);
or OR4 (N497, N462, N312, N90, N128);
buf BUF1 (N498, N481);
nor NOR4 (N499, N496, N371, N354, N62);
nor NOR2 (N500, N495, N49);
buf BUF1 (N501, N493);
nand NAND2 (N502, N499, N335);
and AND3 (N503, N480, N49, N433);
or OR2 (N504, N500, N224);
or OR3 (N505, N498, N392, N324);
nand NAND3 (N506, N505, N49, N307);
nand NAND4 (N507, N504, N502, N474, N434);
not NOT1 (N508, N284);
not NOT1 (N509, N497);
xor XOR2 (N510, N503, N316);
buf BUF1 (N511, N510);
nor NOR3 (N512, N494, N307, N239);
not NOT1 (N513, N508);
not NOT1 (N514, N507);
or OR2 (N515, N506, N416);
nand NAND3 (N516, N488, N479, N322);
nand NAND2 (N517, N515, N397);
and AND2 (N518, N491, N36);
and AND3 (N519, N501, N4, N365);
not NOT1 (N520, N517);
nand NAND2 (N521, N512, N504);
nor NOR4 (N522, N520, N481, N484, N165);
nor NOR3 (N523, N514, N518, N160);
xor XOR2 (N524, N410, N181);
nor NOR4 (N525, N511, N67, N153, N335);
buf BUF1 (N526, N523);
buf BUF1 (N527, N524);
buf BUF1 (N528, N513);
nor NOR2 (N529, N486, N113);
and AND2 (N530, N528, N237);
xor XOR2 (N531, N521, N74);
xor XOR2 (N532, N526, N239);
nand NAND2 (N533, N530, N211);
nand NAND2 (N534, N529, N279);
xor XOR2 (N535, N534, N162);
nand NAND3 (N536, N531, N148, N124);
not NOT1 (N537, N516);
buf BUF1 (N538, N525);
nor NOR4 (N539, N535, N298, N29, N273);
nor NOR2 (N540, N538, N303);
or OR2 (N541, N536, N151);
nor NOR2 (N542, N522, N536);
xor XOR2 (N543, N533, N28);
xor XOR2 (N544, N532, N209);
xor XOR2 (N545, N509, N306);
nor NOR2 (N546, N540, N510);
nor NOR4 (N547, N545, N285, N9, N28);
nor NOR3 (N548, N547, N144, N272);
nand NAND2 (N549, N543, N233);
not NOT1 (N550, N537);
nand NAND3 (N551, N519, N239, N105);
buf BUF1 (N552, N544);
not NOT1 (N553, N542);
nand NAND3 (N554, N550, N462, N411);
and AND2 (N555, N551, N178);
or OR4 (N556, N549, N380, N61, N408);
not NOT1 (N557, N554);
nor NOR3 (N558, N539, N112, N454);
and AND3 (N559, N557, N378, N61);
nor NOR4 (N560, N556, N226, N55, N343);
buf BUF1 (N561, N546);
nand NAND2 (N562, N527, N6);
nand NAND4 (N563, N548, N139, N165, N49);
not NOT1 (N564, N563);
nor NOR2 (N565, N541, N183);
and AND4 (N566, N561, N524, N466, N559);
not NOT1 (N567, N290);
and AND3 (N568, N567, N493, N402);
nand NAND4 (N569, N568, N165, N135, N12);
buf BUF1 (N570, N569);
nand NAND4 (N571, N566, N285, N385, N130);
nand NAND4 (N572, N553, N165, N264, N530);
nand NAND4 (N573, N560, N546, N515, N54);
or OR4 (N574, N565, N314, N186, N173);
and AND3 (N575, N571, N114, N80);
nand NAND2 (N576, N575, N153);
or OR4 (N577, N570, N92, N384, N371);
nand NAND2 (N578, N576, N306);
buf BUF1 (N579, N574);
xor XOR2 (N580, N577, N248);
xor XOR2 (N581, N580, N559);
nand NAND2 (N582, N573, N442);
nor NOR4 (N583, N572, N578, N124, N287);
nand NAND2 (N584, N42, N217);
or OR3 (N585, N552, N50, N282);
buf BUF1 (N586, N562);
not NOT1 (N587, N586);
or OR3 (N588, N558, N365, N443);
xor XOR2 (N589, N582, N277);
nor NOR2 (N590, N581, N49);
not NOT1 (N591, N564);
or OR2 (N592, N589, N54);
nor NOR3 (N593, N579, N298, N589);
buf BUF1 (N594, N591);
buf BUF1 (N595, N583);
or OR3 (N596, N593, N159, N382);
or OR3 (N597, N595, N309, N508);
buf BUF1 (N598, N585);
nor NOR3 (N599, N590, N139, N337);
or OR3 (N600, N555, N382, N591);
nand NAND3 (N601, N587, N154, N397);
nand NAND4 (N602, N601, N502, N64, N37);
or OR4 (N603, N596, N174, N601, N226);
xor XOR2 (N604, N592, N82);
buf BUF1 (N605, N584);
or OR3 (N606, N598, N401, N312);
xor XOR2 (N607, N605, N574);
nand NAND4 (N608, N604, N587, N34, N531);
xor XOR2 (N609, N594, N420);
nor NOR2 (N610, N599, N496);
or OR3 (N611, N608, N535, N171);
not NOT1 (N612, N607);
or OR4 (N613, N606, N534, N103, N438);
endmodule