// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19;

output N1515,N1517,N1505,N1512,N1500,N1486,N1516,N1506,N1514,N1519;

nor NOR4 (N20, N7, N7, N1, N16);
and AND2 (N21, N7, N7);
not NOT1 (N22, N8);
nand NAND3 (N23, N1, N1, N1);
xor XOR2 (N24, N15, N23);
or OR4 (N25, N24, N19, N11, N13);
buf BUF1 (N26, N8);
and AND3 (N27, N24, N21, N10);
nor NOR2 (N28, N1, N18);
xor XOR2 (N29, N28, N2);
or OR4 (N30, N1, N2, N21, N3);
nand NAND2 (N31, N12, N12);
xor XOR2 (N32, N30, N13);
nor NOR4 (N33, N5, N9, N30, N16);
not NOT1 (N34, N20);
nand NAND3 (N35, N5, N31, N5);
xor XOR2 (N36, N34, N24);
xor XOR2 (N37, N25, N35);
buf BUF1 (N38, N29);
nand NAND3 (N39, N29, N7, N34);
or OR3 (N40, N18, N21, N7);
not NOT1 (N41, N40);
nand NAND4 (N42, N26, N21, N15, N14);
not NOT1 (N43, N41);
not NOT1 (N44, N36);
nand NAND4 (N45, N44, N40, N15, N11);
buf BUF1 (N46, N22);
nand NAND4 (N47, N43, N19, N1, N35);
xor XOR2 (N48, N42, N17);
and AND2 (N49, N33, N1);
or OR4 (N50, N49, N34, N40, N6);
and AND4 (N51, N39, N42, N4, N11);
or OR4 (N52, N32, N36, N15, N39);
nor NOR2 (N53, N50, N45);
buf BUF1 (N54, N42);
or OR2 (N55, N52, N44);
nand NAND2 (N56, N55, N20);
nor NOR3 (N57, N47, N2, N47);
and AND2 (N58, N56, N9);
buf BUF1 (N59, N37);
nand NAND4 (N60, N27, N5, N17, N45);
buf BUF1 (N61, N48);
nor NOR2 (N62, N57, N23);
nor NOR3 (N63, N54, N44, N62);
nor NOR2 (N64, N20, N21);
nor NOR4 (N65, N64, N47, N55, N18);
nand NAND3 (N66, N53, N34, N27);
nor NOR3 (N67, N51, N38, N56);
nor NOR2 (N68, N54, N11);
xor XOR2 (N69, N46, N55);
not NOT1 (N70, N63);
xor XOR2 (N71, N70, N66);
or OR2 (N72, N32, N44);
and AND4 (N73, N65, N57, N32, N22);
and AND4 (N74, N69, N22, N3, N33);
and AND4 (N75, N71, N3, N15, N1);
nor NOR3 (N76, N60, N41, N51);
nand NAND2 (N77, N75, N46);
xor XOR2 (N78, N58, N52);
or OR4 (N79, N76, N12, N75, N28);
xor XOR2 (N80, N72, N4);
and AND4 (N81, N80, N4, N8, N45);
not NOT1 (N82, N68);
nor NOR4 (N83, N59, N44, N14, N65);
nor NOR3 (N84, N73, N33, N26);
not NOT1 (N85, N82);
buf BUF1 (N86, N67);
or OR3 (N87, N78, N54, N79);
and AND3 (N88, N69, N45, N19);
nor NOR4 (N89, N61, N35, N57, N25);
and AND4 (N90, N88, N1, N53, N54);
xor XOR2 (N91, N74, N27);
nor NOR4 (N92, N90, N4, N55, N13);
and AND4 (N93, N89, N9, N79, N18);
buf BUF1 (N94, N84);
buf BUF1 (N95, N92);
or OR3 (N96, N85, N14, N11);
xor XOR2 (N97, N81, N83);
buf BUF1 (N98, N41);
nor NOR3 (N99, N97, N31, N45);
buf BUF1 (N100, N93);
nand NAND3 (N101, N95, N88, N43);
nand NAND2 (N102, N99, N75);
or OR3 (N103, N91, N25, N77);
nor NOR4 (N104, N65, N35, N15, N35);
and AND3 (N105, N101, N79, N24);
or OR4 (N106, N100, N47, N20, N57);
and AND3 (N107, N87, N17, N55);
nand NAND3 (N108, N86, N38, N75);
nand NAND3 (N109, N105, N30, N83);
xor XOR2 (N110, N102, N16);
nor NOR3 (N111, N110, N36, N17);
nor NOR4 (N112, N96, N23, N67, N91);
nor NOR3 (N113, N103, N21, N70);
xor XOR2 (N114, N112, N49);
nand NAND2 (N115, N106, N103);
not NOT1 (N116, N109);
buf BUF1 (N117, N116);
nor NOR4 (N118, N94, N24, N22, N80);
not NOT1 (N119, N98);
not NOT1 (N120, N108);
and AND4 (N121, N107, N108, N41, N14);
nand NAND4 (N122, N115, N52, N70, N66);
xor XOR2 (N123, N119, N41);
nand NAND4 (N124, N121, N12, N34, N38);
nand NAND2 (N125, N111, N103);
xor XOR2 (N126, N114, N43);
nand NAND3 (N127, N125, N75, N41);
not NOT1 (N128, N118);
nor NOR2 (N129, N122, N104);
nor NOR4 (N130, N47, N42, N58, N52);
nand NAND4 (N131, N113, N48, N93, N122);
xor XOR2 (N132, N124, N28);
nand NAND3 (N133, N132, N40, N61);
and AND3 (N134, N133, N11, N25);
buf BUF1 (N135, N134);
or OR3 (N136, N117, N108, N50);
or OR2 (N137, N128, N2);
nand NAND3 (N138, N130, N86, N45);
and AND4 (N139, N129, N65, N116, N124);
buf BUF1 (N140, N126);
and AND3 (N141, N136, N122, N114);
nor NOR4 (N142, N127, N24, N109, N26);
and AND3 (N143, N138, N35, N17);
or OR4 (N144, N137, N8, N83, N33);
and AND4 (N145, N144, N46, N41, N30);
buf BUF1 (N146, N139);
nand NAND4 (N147, N145, N137, N63, N36);
nand NAND3 (N148, N143, N9, N123);
xor XOR2 (N149, N143, N29);
not NOT1 (N150, N141);
nor NOR3 (N151, N150, N105, N23);
nor NOR4 (N152, N151, N130, N107, N45);
nor NOR2 (N153, N146, N87);
or OR3 (N154, N152, N19, N74);
nand NAND2 (N155, N147, N34);
nor NOR2 (N156, N155, N145);
nand NAND4 (N157, N142, N117, N64, N81);
and AND2 (N158, N131, N112);
nor NOR3 (N159, N154, N18, N7);
nand NAND2 (N160, N120, N4);
or OR4 (N161, N157, N43, N120, N55);
not NOT1 (N162, N160);
not NOT1 (N163, N162);
nand NAND4 (N164, N159, N82, N128, N47);
xor XOR2 (N165, N164, N147);
nand NAND4 (N166, N149, N94, N102, N3);
buf BUF1 (N167, N158);
nand NAND3 (N168, N167, N129, N44);
not NOT1 (N169, N168);
buf BUF1 (N170, N166);
and AND4 (N171, N169, N105, N46, N37);
nand NAND3 (N172, N163, N49, N70);
xor XOR2 (N173, N135, N90);
and AND2 (N174, N140, N142);
or OR3 (N175, N171, N153, N48);
or OR3 (N176, N29, N155, N135);
not NOT1 (N177, N172);
not NOT1 (N178, N173);
xor XOR2 (N179, N174, N141);
and AND2 (N180, N170, N149);
xor XOR2 (N181, N176, N174);
nand NAND2 (N182, N180, N39);
and AND4 (N183, N178, N38, N119, N23);
or OR3 (N184, N148, N183, N182);
nand NAND3 (N185, N101, N100, N74);
nor NOR3 (N186, N84, N17, N48);
nand NAND3 (N187, N185, N57, N19);
nand NAND3 (N188, N177, N67, N166);
buf BUF1 (N189, N179);
not NOT1 (N190, N156);
nand NAND2 (N191, N190, N104);
not NOT1 (N192, N184);
nor NOR4 (N193, N191, N28, N121, N14);
buf BUF1 (N194, N193);
or OR4 (N195, N189, N99, N12, N36);
or OR2 (N196, N161, N33);
or OR2 (N197, N186, N101);
and AND2 (N198, N181, N13);
not NOT1 (N199, N188);
and AND2 (N200, N175, N42);
and AND3 (N201, N165, N165, N156);
nand NAND3 (N202, N187, N8, N75);
not NOT1 (N203, N199);
or OR3 (N204, N201, N15, N195);
xor XOR2 (N205, N77, N162);
xor XOR2 (N206, N204, N63);
or OR3 (N207, N203, N28, N172);
xor XOR2 (N208, N207, N17);
xor XOR2 (N209, N194, N125);
or OR2 (N210, N206, N9);
xor XOR2 (N211, N205, N194);
nor NOR2 (N212, N192, N113);
not NOT1 (N213, N208);
and AND2 (N214, N198, N108);
not NOT1 (N215, N214);
or OR4 (N216, N213, N181, N208, N32);
or OR2 (N217, N209, N96);
not NOT1 (N218, N217);
and AND2 (N219, N210, N78);
nand NAND4 (N220, N215, N111, N159, N113);
or OR2 (N221, N218, N202);
and AND2 (N222, N33, N154);
xor XOR2 (N223, N197, N189);
or OR2 (N224, N220, N99);
and AND4 (N225, N224, N151, N6, N176);
and AND4 (N226, N212, N44, N102, N148);
buf BUF1 (N227, N225);
not NOT1 (N228, N221);
nor NOR4 (N229, N219, N183, N21, N74);
or OR3 (N230, N196, N225, N42);
and AND4 (N231, N228, N175, N195, N32);
xor XOR2 (N232, N226, N159);
nand NAND3 (N233, N231, N21, N229);
buf BUF1 (N234, N93);
or OR2 (N235, N230, N154);
and AND2 (N236, N223, N42);
nand NAND4 (N237, N222, N211, N165, N175);
xor XOR2 (N238, N140, N224);
xor XOR2 (N239, N232, N106);
nor NOR4 (N240, N239, N21, N59, N9);
nand NAND3 (N241, N216, N121, N105);
xor XOR2 (N242, N234, N49);
buf BUF1 (N243, N242);
buf BUF1 (N244, N233);
and AND2 (N245, N241, N150);
nor NOR3 (N246, N200, N70, N155);
xor XOR2 (N247, N246, N72);
nand NAND4 (N248, N237, N198, N91, N180);
xor XOR2 (N249, N240, N77);
nand NAND4 (N250, N245, N49, N184, N13);
or OR4 (N251, N227, N40, N70, N4);
not NOT1 (N252, N251);
xor XOR2 (N253, N248, N13);
or OR3 (N254, N238, N83, N173);
or OR3 (N255, N235, N183, N142);
nand NAND2 (N256, N255, N108);
not NOT1 (N257, N252);
xor XOR2 (N258, N243, N151);
and AND2 (N259, N253, N89);
nand NAND3 (N260, N256, N148, N50);
not NOT1 (N261, N259);
xor XOR2 (N262, N244, N26);
not NOT1 (N263, N261);
not NOT1 (N264, N247);
not NOT1 (N265, N264);
not NOT1 (N266, N262);
buf BUF1 (N267, N258);
or OR2 (N268, N266, N151);
xor XOR2 (N269, N268, N124);
nand NAND4 (N270, N250, N158, N158, N71);
xor XOR2 (N271, N269, N30);
buf BUF1 (N272, N263);
not NOT1 (N273, N257);
and AND2 (N274, N249, N255);
buf BUF1 (N275, N274);
or OR4 (N276, N236, N257, N158, N44);
and AND2 (N277, N270, N218);
and AND3 (N278, N254, N50, N170);
or OR3 (N279, N271, N147, N66);
nor NOR3 (N280, N260, N10, N234);
and AND4 (N281, N278, N174, N51, N164);
not NOT1 (N282, N273);
and AND3 (N283, N280, N153, N228);
buf BUF1 (N284, N281);
not NOT1 (N285, N284);
or OR3 (N286, N267, N19, N37);
xor XOR2 (N287, N285, N251);
xor XOR2 (N288, N277, N3);
nor NOR4 (N289, N276, N273, N139, N176);
or OR4 (N290, N282, N19, N31, N26);
buf BUF1 (N291, N279);
not NOT1 (N292, N275);
nor NOR2 (N293, N292, N7);
buf BUF1 (N294, N290);
or OR4 (N295, N287, N132, N289, N174);
xor XOR2 (N296, N233, N291);
buf BUF1 (N297, N162);
xor XOR2 (N298, N295, N236);
and AND4 (N299, N297, N135, N71, N165);
nor NOR2 (N300, N288, N248);
buf BUF1 (N301, N299);
nand NAND3 (N302, N294, N148, N44);
nand NAND3 (N303, N293, N192, N98);
nand NAND2 (N304, N303, N129);
xor XOR2 (N305, N296, N75);
nor NOR4 (N306, N300, N3, N131, N109);
xor XOR2 (N307, N265, N86);
xor XOR2 (N308, N305, N149);
or OR2 (N309, N307, N280);
nand NAND3 (N310, N308, N155, N258);
nor NOR4 (N311, N301, N106, N186, N214);
nand NAND2 (N312, N298, N228);
and AND2 (N313, N310, N4);
xor XOR2 (N314, N311, N268);
nor NOR4 (N315, N309, N56, N93, N299);
not NOT1 (N316, N272);
or OR2 (N317, N313, N231);
and AND3 (N318, N286, N160, N199);
not NOT1 (N319, N316);
not NOT1 (N320, N317);
buf BUF1 (N321, N302);
buf BUF1 (N322, N315);
or OR2 (N323, N318, N44);
nor NOR3 (N324, N322, N151, N71);
xor XOR2 (N325, N323, N34);
nor NOR2 (N326, N320, N232);
and AND3 (N327, N325, N304, N106);
xor XOR2 (N328, N313, N282);
xor XOR2 (N329, N319, N290);
buf BUF1 (N330, N327);
or OR3 (N331, N330, N318, N37);
or OR2 (N332, N328, N107);
or OR2 (N333, N283, N145);
not NOT1 (N334, N331);
xor XOR2 (N335, N329, N72);
and AND4 (N336, N321, N3, N202, N160);
nor NOR3 (N337, N326, N143, N323);
nor NOR4 (N338, N312, N26, N220, N133);
nor NOR2 (N339, N334, N18);
buf BUF1 (N340, N324);
nor NOR3 (N341, N339, N263, N76);
xor XOR2 (N342, N340, N225);
not NOT1 (N343, N342);
xor XOR2 (N344, N314, N158);
buf BUF1 (N345, N341);
and AND4 (N346, N332, N15, N243, N60);
buf BUF1 (N347, N338);
not NOT1 (N348, N347);
nand NAND4 (N349, N336, N323, N348, N65);
xor XOR2 (N350, N295, N232);
nand NAND4 (N351, N306, N189, N115, N89);
or OR3 (N352, N345, N257, N326);
not NOT1 (N353, N351);
xor XOR2 (N354, N350, N295);
not NOT1 (N355, N349);
buf BUF1 (N356, N353);
and AND3 (N357, N335, N167, N288);
nand NAND3 (N358, N352, N285, N18);
xor XOR2 (N359, N356, N22);
buf BUF1 (N360, N337);
and AND4 (N361, N343, N175, N79, N123);
buf BUF1 (N362, N355);
and AND3 (N363, N359, N207, N275);
buf BUF1 (N364, N362);
not NOT1 (N365, N357);
or OR4 (N366, N358, N213, N358, N43);
buf BUF1 (N367, N333);
and AND4 (N368, N366, N151, N261, N202);
not NOT1 (N369, N360);
or OR2 (N370, N354, N214);
nor NOR3 (N371, N370, N256, N261);
nor NOR2 (N372, N365, N74);
buf BUF1 (N373, N372);
buf BUF1 (N374, N361);
not NOT1 (N375, N344);
nand NAND4 (N376, N367, N301, N297, N145);
not NOT1 (N377, N374);
nand NAND4 (N378, N377, N226, N62, N247);
nand NAND2 (N379, N368, N358);
nand NAND2 (N380, N371, N258);
not NOT1 (N381, N375);
nor NOR2 (N382, N373, N112);
not NOT1 (N383, N380);
xor XOR2 (N384, N383, N25);
nand NAND4 (N385, N376, N378, N282, N72);
nor NOR3 (N386, N294, N75, N210);
or OR4 (N387, N364, N11, N352, N356);
nor NOR3 (N388, N346, N76, N122);
and AND3 (N389, N386, N388, N378);
xor XOR2 (N390, N242, N346);
xor XOR2 (N391, N389, N217);
not NOT1 (N392, N384);
or OR2 (N393, N391, N215);
not NOT1 (N394, N382);
nand NAND3 (N395, N394, N25, N129);
or OR3 (N396, N369, N364, N109);
xor XOR2 (N397, N390, N188);
nand NAND4 (N398, N397, N336, N142, N119);
nand NAND3 (N399, N363, N311, N359);
and AND4 (N400, N393, N241, N187, N26);
xor XOR2 (N401, N396, N368);
or OR4 (N402, N401, N107, N395, N354);
buf BUF1 (N403, N269);
not NOT1 (N404, N398);
or OR2 (N405, N399, N146);
nor NOR3 (N406, N381, N39, N113);
nand NAND3 (N407, N392, N139, N89);
nand NAND4 (N408, N403, N270, N306, N241);
nand NAND2 (N409, N408, N132);
or OR3 (N410, N387, N13, N282);
buf BUF1 (N411, N409);
nand NAND2 (N412, N406, N107);
nor NOR2 (N413, N379, N19);
xor XOR2 (N414, N405, N216);
xor XOR2 (N415, N400, N71);
buf BUF1 (N416, N410);
buf BUF1 (N417, N415);
nor NOR4 (N418, N411, N239, N259, N292);
nor NOR3 (N419, N418, N349, N115);
not NOT1 (N420, N417);
nor NOR4 (N421, N407, N367, N48, N81);
not NOT1 (N422, N413);
nor NOR4 (N423, N421, N265, N323, N134);
nand NAND4 (N424, N420, N87, N216, N130);
nor NOR3 (N425, N423, N95, N305);
nand NAND3 (N426, N425, N274, N207);
not NOT1 (N427, N419);
nand NAND3 (N428, N427, N116, N69);
not NOT1 (N429, N385);
or OR4 (N430, N414, N99, N188, N318);
nand NAND3 (N431, N416, N232, N146);
buf BUF1 (N432, N404);
xor XOR2 (N433, N428, N67);
nor NOR2 (N434, N432, N381);
nor NOR2 (N435, N434, N49);
not NOT1 (N436, N435);
not NOT1 (N437, N402);
and AND4 (N438, N433, N437, N121, N12);
xor XOR2 (N439, N42, N259);
nor NOR3 (N440, N430, N330, N427);
not NOT1 (N441, N429);
nor NOR3 (N442, N422, N170, N146);
nand NAND2 (N443, N440, N67);
buf BUF1 (N444, N442);
xor XOR2 (N445, N441, N217);
xor XOR2 (N446, N436, N2);
nand NAND4 (N447, N426, N186, N210, N110);
not NOT1 (N448, N439);
nand NAND2 (N449, N445, N109);
xor XOR2 (N450, N449, N226);
nand NAND4 (N451, N446, N159, N144, N99);
and AND4 (N452, N424, N296, N420, N263);
or OR3 (N453, N412, N262, N324);
xor XOR2 (N454, N431, N82);
buf BUF1 (N455, N438);
buf BUF1 (N456, N454);
and AND2 (N457, N444, N388);
xor XOR2 (N458, N456, N130);
or OR3 (N459, N443, N425, N216);
xor XOR2 (N460, N451, N227);
not NOT1 (N461, N453);
not NOT1 (N462, N452);
buf BUF1 (N463, N461);
buf BUF1 (N464, N460);
buf BUF1 (N465, N457);
and AND4 (N466, N448, N107, N163, N456);
nand NAND2 (N467, N465, N450);
or OR3 (N468, N250, N448, N22);
nand NAND2 (N469, N467, N142);
buf BUF1 (N470, N468);
not NOT1 (N471, N458);
buf BUF1 (N472, N469);
nand NAND2 (N473, N447, N443);
or OR3 (N474, N459, N21, N211);
or OR4 (N475, N463, N391, N287, N256);
and AND3 (N476, N462, N360, N9);
nor NOR4 (N477, N476, N277, N188, N179);
not NOT1 (N478, N473);
or OR3 (N479, N455, N256, N132);
buf BUF1 (N480, N472);
nor NOR4 (N481, N480, N142, N251, N279);
nor NOR2 (N482, N464, N150);
or OR3 (N483, N470, N341, N241);
nand NAND3 (N484, N475, N267, N347);
buf BUF1 (N485, N474);
nand NAND2 (N486, N477, N268);
buf BUF1 (N487, N479);
nor NOR4 (N488, N486, N108, N473, N294);
and AND4 (N489, N488, N282, N458, N172);
xor XOR2 (N490, N483, N118);
buf BUF1 (N491, N481);
and AND2 (N492, N484, N456);
xor XOR2 (N493, N489, N474);
buf BUF1 (N494, N493);
nand NAND4 (N495, N482, N455, N375, N285);
or OR4 (N496, N471, N437, N116, N236);
nand NAND4 (N497, N490, N63, N402, N64);
nand NAND3 (N498, N496, N479, N319);
not NOT1 (N499, N498);
and AND3 (N500, N478, N331, N14);
nand NAND3 (N501, N492, N36, N257);
not NOT1 (N502, N491);
or OR2 (N503, N487, N161);
xor XOR2 (N504, N497, N205);
nand NAND4 (N505, N501, N361, N256, N59);
or OR2 (N506, N502, N328);
buf BUF1 (N507, N506);
nand NAND2 (N508, N507, N406);
xor XOR2 (N509, N508, N1);
nor NOR2 (N510, N494, N354);
and AND4 (N511, N466, N365, N382, N103);
buf BUF1 (N512, N505);
xor XOR2 (N513, N500, N381);
and AND2 (N514, N485, N100);
not NOT1 (N515, N509);
not NOT1 (N516, N495);
xor XOR2 (N517, N504, N255);
nor NOR3 (N518, N516, N136, N323);
or OR3 (N519, N503, N454, N381);
or OR2 (N520, N519, N202);
nor NOR4 (N521, N512, N115, N77, N220);
not NOT1 (N522, N518);
not NOT1 (N523, N521);
not NOT1 (N524, N514);
nor NOR4 (N525, N499, N211, N288, N516);
and AND4 (N526, N524, N132, N437, N322);
xor XOR2 (N527, N513, N301);
nand NAND3 (N528, N515, N60, N336);
or OR3 (N529, N523, N155, N273);
nand NAND4 (N530, N511, N92, N69, N273);
buf BUF1 (N531, N530);
buf BUF1 (N532, N526);
nand NAND2 (N533, N528, N387);
not NOT1 (N534, N525);
xor XOR2 (N535, N531, N153);
and AND4 (N536, N532, N84, N11, N339);
and AND2 (N537, N522, N46);
or OR2 (N538, N537, N4);
buf BUF1 (N539, N538);
or OR2 (N540, N520, N198);
not NOT1 (N541, N533);
and AND2 (N542, N536, N55);
nand NAND3 (N543, N539, N424, N46);
xor XOR2 (N544, N542, N219);
buf BUF1 (N545, N534);
or OR3 (N546, N544, N489, N135);
or OR3 (N547, N546, N229, N218);
buf BUF1 (N548, N535);
buf BUF1 (N549, N541);
and AND4 (N550, N529, N298, N246, N96);
or OR4 (N551, N550, N125, N544, N100);
buf BUF1 (N552, N551);
nor NOR2 (N553, N549, N406);
xor XOR2 (N554, N527, N446);
not NOT1 (N555, N548);
or OR3 (N556, N543, N214, N320);
and AND4 (N557, N545, N32, N463, N396);
not NOT1 (N558, N540);
xor XOR2 (N559, N557, N16);
or OR3 (N560, N517, N509, N435);
or OR3 (N561, N560, N359, N18);
nand NAND4 (N562, N559, N393, N152, N506);
xor XOR2 (N563, N552, N500);
or OR3 (N564, N555, N270, N29);
nor NOR2 (N565, N553, N301);
nor NOR3 (N566, N564, N109, N412);
xor XOR2 (N567, N563, N456);
buf BUF1 (N568, N554);
not NOT1 (N569, N561);
nand NAND2 (N570, N556, N240);
buf BUF1 (N571, N567);
and AND2 (N572, N568, N428);
and AND3 (N573, N558, N291, N279);
nor NOR3 (N574, N566, N223, N52);
nor NOR3 (N575, N573, N203, N268);
nor NOR4 (N576, N572, N85, N238, N202);
not NOT1 (N577, N571);
nor NOR4 (N578, N575, N461, N456, N283);
nor NOR3 (N579, N577, N495, N303);
buf BUF1 (N580, N570);
xor XOR2 (N581, N562, N88);
nand NAND3 (N582, N574, N440, N172);
buf BUF1 (N583, N510);
nor NOR4 (N584, N579, N238, N76, N376);
nor NOR4 (N585, N582, N400, N46, N174);
buf BUF1 (N586, N547);
or OR3 (N587, N581, N189, N551);
nor NOR2 (N588, N583, N161);
or OR3 (N589, N578, N529, N135);
buf BUF1 (N590, N585);
xor XOR2 (N591, N586, N532);
not NOT1 (N592, N584);
or OR4 (N593, N590, N374, N274, N366);
nor NOR3 (N594, N576, N284, N250);
buf BUF1 (N595, N589);
buf BUF1 (N596, N588);
nor NOR2 (N597, N565, N448);
not NOT1 (N598, N596);
buf BUF1 (N599, N569);
buf BUF1 (N600, N587);
and AND3 (N601, N593, N39, N434);
nor NOR3 (N602, N601, N267, N571);
and AND3 (N603, N597, N120, N430);
xor XOR2 (N604, N595, N537);
and AND2 (N605, N603, N470);
nor NOR4 (N606, N605, N233, N241, N124);
and AND2 (N607, N592, N462);
and AND3 (N608, N591, N438, N5);
or OR3 (N609, N598, N468, N574);
or OR4 (N610, N599, N188, N352, N356);
and AND3 (N611, N594, N306, N396);
not NOT1 (N612, N608);
not NOT1 (N613, N607);
and AND4 (N614, N604, N261, N16, N246);
xor XOR2 (N615, N602, N138);
buf BUF1 (N616, N615);
buf BUF1 (N617, N614);
nand NAND4 (N618, N610, N400, N279, N198);
xor XOR2 (N619, N616, N462);
buf BUF1 (N620, N600);
xor XOR2 (N621, N609, N533);
not NOT1 (N622, N621);
buf BUF1 (N623, N613);
buf BUF1 (N624, N606);
nor NOR4 (N625, N622, N52, N369, N213);
buf BUF1 (N626, N624);
not NOT1 (N627, N612);
xor XOR2 (N628, N611, N226);
or OR2 (N629, N623, N15);
buf BUF1 (N630, N626);
nor NOR2 (N631, N620, N411);
nand NAND4 (N632, N627, N28, N495, N103);
nand NAND2 (N633, N629, N371);
nand NAND3 (N634, N628, N36, N623);
nor NOR3 (N635, N618, N204, N218);
or OR2 (N636, N633, N422);
nor NOR3 (N637, N631, N240, N482);
xor XOR2 (N638, N625, N302);
and AND4 (N639, N619, N556, N10, N584);
buf BUF1 (N640, N630);
xor XOR2 (N641, N636, N271);
nand NAND3 (N642, N638, N365, N623);
and AND2 (N643, N639, N244);
buf BUF1 (N644, N632);
nor NOR2 (N645, N580, N511);
nand NAND2 (N646, N641, N287);
xor XOR2 (N647, N646, N600);
or OR3 (N648, N647, N632, N179);
buf BUF1 (N649, N648);
nor NOR3 (N650, N637, N312, N524);
nand NAND3 (N651, N650, N535, N149);
not NOT1 (N652, N617);
not NOT1 (N653, N649);
nor NOR3 (N654, N651, N181, N526);
xor XOR2 (N655, N642, N419);
not NOT1 (N656, N645);
buf BUF1 (N657, N656);
xor XOR2 (N658, N643, N207);
and AND2 (N659, N634, N93);
nor NOR4 (N660, N652, N405, N28, N331);
xor XOR2 (N661, N640, N653);
nand NAND3 (N662, N246, N154, N527);
nand NAND2 (N663, N658, N486);
and AND4 (N664, N654, N245, N318, N89);
xor XOR2 (N665, N664, N196);
or OR3 (N666, N661, N34, N347);
not NOT1 (N667, N662);
nand NAND3 (N668, N660, N161, N303);
and AND4 (N669, N644, N458, N585, N370);
not NOT1 (N670, N665);
and AND4 (N671, N663, N597, N36, N667);
and AND2 (N672, N26, N91);
not NOT1 (N673, N635);
xor XOR2 (N674, N657, N103);
xor XOR2 (N675, N669, N587);
and AND3 (N676, N675, N335, N664);
and AND4 (N677, N659, N324, N444, N50);
buf BUF1 (N678, N674);
xor XOR2 (N679, N676, N77);
buf BUF1 (N680, N673);
buf BUF1 (N681, N655);
or OR4 (N682, N670, N254, N380, N228);
or OR4 (N683, N682, N213, N527, N381);
xor XOR2 (N684, N677, N578);
not NOT1 (N685, N666);
buf BUF1 (N686, N685);
buf BUF1 (N687, N679);
or OR2 (N688, N671, N567);
nand NAND4 (N689, N687, N295, N45, N256);
nand NAND4 (N690, N672, N254, N163, N371);
buf BUF1 (N691, N681);
nand NAND2 (N692, N683, N333);
and AND4 (N693, N680, N400, N585, N541);
and AND2 (N694, N668, N439);
buf BUF1 (N695, N678);
not NOT1 (N696, N690);
buf BUF1 (N697, N691);
nor NOR2 (N698, N697, N691);
nand NAND2 (N699, N688, N642);
nor NOR4 (N700, N686, N459, N299, N104);
not NOT1 (N701, N696);
nor NOR3 (N702, N694, N676, N600);
nor NOR3 (N703, N695, N414, N632);
not NOT1 (N704, N693);
not NOT1 (N705, N698);
not NOT1 (N706, N703);
buf BUF1 (N707, N700);
and AND4 (N708, N692, N634, N405, N466);
xor XOR2 (N709, N699, N121);
nand NAND3 (N710, N708, N673, N466);
not NOT1 (N711, N704);
nor NOR4 (N712, N707, N186, N376, N630);
nor NOR2 (N713, N702, N231);
xor XOR2 (N714, N709, N165);
xor XOR2 (N715, N713, N519);
or OR2 (N716, N684, N563);
or OR4 (N717, N701, N226, N494, N708);
or OR2 (N718, N710, N184);
buf BUF1 (N719, N716);
nand NAND4 (N720, N714, N80, N619, N396);
and AND3 (N721, N719, N672, N466);
not NOT1 (N722, N689);
xor XOR2 (N723, N711, N570);
and AND2 (N724, N723, N514);
not NOT1 (N725, N721);
xor XOR2 (N726, N706, N259);
xor XOR2 (N727, N718, N43);
or OR4 (N728, N725, N418, N572, N589);
not NOT1 (N729, N726);
nand NAND4 (N730, N717, N460, N445, N439);
nand NAND2 (N731, N729, N557);
not NOT1 (N732, N712);
xor XOR2 (N733, N730, N463);
and AND3 (N734, N715, N439, N572);
buf BUF1 (N735, N720);
xor XOR2 (N736, N722, N684);
not NOT1 (N737, N727);
nor NOR3 (N738, N724, N257, N277);
nor NOR4 (N739, N737, N327, N50, N505);
nor NOR2 (N740, N738, N405);
and AND4 (N741, N728, N484, N353, N267);
nand NAND3 (N742, N734, N69, N517);
buf BUF1 (N743, N739);
or OR3 (N744, N736, N362, N632);
and AND3 (N745, N740, N19, N511);
xor XOR2 (N746, N741, N378);
or OR2 (N747, N705, N426);
buf BUF1 (N748, N744);
buf BUF1 (N749, N732);
nor NOR4 (N750, N747, N17, N704, N94);
nor NOR4 (N751, N749, N131, N428, N445);
not NOT1 (N752, N746);
buf BUF1 (N753, N748);
xor XOR2 (N754, N731, N313);
and AND4 (N755, N754, N132, N739, N233);
xor XOR2 (N756, N750, N578);
xor XOR2 (N757, N751, N13);
not NOT1 (N758, N755);
or OR3 (N759, N757, N173, N159);
and AND2 (N760, N745, N115);
or OR3 (N761, N743, N177, N490);
nand NAND3 (N762, N733, N697, N457);
or OR4 (N763, N760, N480, N411, N513);
buf BUF1 (N764, N763);
xor XOR2 (N765, N759, N521);
nand NAND2 (N766, N764, N154);
and AND4 (N767, N766, N147, N666, N252);
and AND3 (N768, N735, N80, N546);
or OR2 (N769, N762, N27);
not NOT1 (N770, N752);
xor XOR2 (N771, N768, N206);
or OR2 (N772, N767, N399);
nor NOR2 (N773, N756, N223);
nand NAND2 (N774, N758, N449);
nand NAND4 (N775, N771, N293, N552, N255);
and AND4 (N776, N773, N580, N438, N167);
nor NOR2 (N777, N753, N299);
not NOT1 (N778, N770);
or OR3 (N779, N742, N606, N349);
xor XOR2 (N780, N774, N176);
or OR2 (N781, N776, N528);
xor XOR2 (N782, N777, N39);
and AND4 (N783, N765, N213, N474, N31);
nand NAND4 (N784, N778, N606, N363, N617);
not NOT1 (N785, N761);
nor NOR3 (N786, N783, N625, N521);
nand NAND4 (N787, N779, N109, N740, N759);
and AND2 (N788, N780, N556);
and AND3 (N789, N772, N249, N232);
buf BUF1 (N790, N789);
xor XOR2 (N791, N788, N751);
buf BUF1 (N792, N781);
xor XOR2 (N793, N792, N239);
xor XOR2 (N794, N790, N549);
not NOT1 (N795, N787);
nand NAND3 (N796, N786, N398, N156);
and AND4 (N797, N796, N300, N486, N641);
buf BUF1 (N798, N793);
xor XOR2 (N799, N791, N706);
and AND3 (N800, N795, N164, N526);
nor NOR2 (N801, N769, N31);
nor NOR2 (N802, N794, N325);
buf BUF1 (N803, N802);
or OR3 (N804, N798, N356, N599);
nor NOR3 (N805, N785, N256, N383);
nor NOR3 (N806, N801, N740, N663);
xor XOR2 (N807, N775, N209);
buf BUF1 (N808, N799);
xor XOR2 (N809, N782, N389);
xor XOR2 (N810, N806, N241);
not NOT1 (N811, N803);
and AND3 (N812, N797, N543, N362);
nand NAND2 (N813, N811, N311);
not NOT1 (N814, N800);
buf BUF1 (N815, N810);
and AND2 (N816, N812, N20);
or OR2 (N817, N809, N705);
or OR3 (N818, N816, N733, N632);
xor XOR2 (N819, N814, N94);
buf BUF1 (N820, N817);
xor XOR2 (N821, N807, N329);
not NOT1 (N822, N784);
xor XOR2 (N823, N815, N640);
not NOT1 (N824, N821);
nand NAND2 (N825, N824, N317);
not NOT1 (N826, N819);
and AND2 (N827, N820, N466);
or OR3 (N828, N822, N280, N536);
nor NOR3 (N829, N823, N44, N94);
and AND2 (N830, N805, N594);
not NOT1 (N831, N808);
buf BUF1 (N832, N818);
or OR2 (N833, N827, N325);
nand NAND4 (N834, N826, N748, N611, N705);
nor NOR3 (N835, N831, N136, N229);
nor NOR2 (N836, N830, N792);
xor XOR2 (N837, N835, N474);
nor NOR4 (N838, N829, N280, N832, N835);
or OR3 (N839, N357, N690, N240);
nor NOR3 (N840, N834, N495, N540);
buf BUF1 (N841, N833);
buf BUF1 (N842, N836);
and AND3 (N843, N837, N313, N814);
buf BUF1 (N844, N825);
nor NOR2 (N845, N838, N281);
xor XOR2 (N846, N844, N26);
nor NOR2 (N847, N813, N171);
nand NAND4 (N848, N839, N794, N647, N165);
nor NOR2 (N849, N828, N151);
not NOT1 (N850, N846);
xor XOR2 (N851, N804, N779);
not NOT1 (N852, N843);
buf BUF1 (N853, N840);
or OR3 (N854, N853, N702, N114);
nor NOR3 (N855, N847, N36, N633);
nor NOR4 (N856, N852, N759, N499, N450);
buf BUF1 (N857, N842);
nor NOR2 (N858, N851, N539);
not NOT1 (N859, N857);
buf BUF1 (N860, N849);
buf BUF1 (N861, N854);
and AND4 (N862, N860, N406, N697, N498);
nand NAND3 (N863, N845, N120, N589);
nor NOR4 (N864, N856, N626, N603, N281);
and AND2 (N865, N861, N67);
or OR4 (N866, N855, N731, N304, N56);
nor NOR4 (N867, N865, N415, N596, N531);
not NOT1 (N868, N864);
not NOT1 (N869, N841);
nand NAND3 (N870, N850, N307, N65);
nand NAND2 (N871, N862, N163);
nor NOR4 (N872, N848, N628, N589, N184);
nor NOR3 (N873, N859, N68, N781);
and AND3 (N874, N866, N348, N113);
xor XOR2 (N875, N868, N241);
not NOT1 (N876, N869);
not NOT1 (N877, N875);
nand NAND3 (N878, N870, N129, N133);
or OR3 (N879, N873, N541, N571);
buf BUF1 (N880, N872);
xor XOR2 (N881, N871, N674);
nand NAND2 (N882, N858, N358);
nand NAND2 (N883, N878, N64);
not NOT1 (N884, N882);
buf BUF1 (N885, N863);
nand NAND4 (N886, N880, N130, N146, N635);
buf BUF1 (N887, N876);
and AND3 (N888, N874, N8, N252);
not NOT1 (N889, N884);
not NOT1 (N890, N888);
buf BUF1 (N891, N887);
nor NOR4 (N892, N877, N105, N43, N559);
buf BUF1 (N893, N867);
xor XOR2 (N894, N892, N597);
nor NOR2 (N895, N889, N6);
or OR2 (N896, N881, N643);
nor NOR3 (N897, N885, N632, N500);
xor XOR2 (N898, N883, N384);
xor XOR2 (N899, N891, N271);
not NOT1 (N900, N893);
nor NOR4 (N901, N899, N568, N797, N244);
and AND3 (N902, N886, N803, N469);
nor NOR3 (N903, N879, N401, N424);
nor NOR4 (N904, N895, N222, N133, N152);
xor XOR2 (N905, N900, N344);
xor XOR2 (N906, N901, N530);
nand NAND2 (N907, N905, N138);
xor XOR2 (N908, N903, N677);
and AND3 (N909, N904, N540, N71);
nor NOR2 (N910, N909, N339);
not NOT1 (N911, N908);
not NOT1 (N912, N906);
nor NOR2 (N913, N912, N879);
nor NOR3 (N914, N913, N683, N75);
nor NOR4 (N915, N914, N404, N2, N343);
xor XOR2 (N916, N907, N420);
buf BUF1 (N917, N902);
not NOT1 (N918, N896);
not NOT1 (N919, N897);
and AND3 (N920, N898, N256, N582);
xor XOR2 (N921, N910, N361);
not NOT1 (N922, N918);
not NOT1 (N923, N915);
nor NOR2 (N924, N916, N842);
nand NAND2 (N925, N919, N268);
nor NOR4 (N926, N920, N214, N75, N342);
nor NOR3 (N927, N925, N41, N854);
nor NOR4 (N928, N927, N717, N863, N398);
xor XOR2 (N929, N922, N819);
not NOT1 (N930, N928);
xor XOR2 (N931, N890, N60);
nand NAND4 (N932, N921, N649, N349, N3);
not NOT1 (N933, N917);
nor NOR2 (N934, N931, N372);
nand NAND4 (N935, N926, N925, N54, N325);
buf BUF1 (N936, N929);
or OR4 (N937, N930, N590, N726, N765);
not NOT1 (N938, N924);
or OR3 (N939, N933, N679, N9);
buf BUF1 (N940, N939);
or OR2 (N941, N937, N901);
buf BUF1 (N942, N936);
not NOT1 (N943, N938);
nor NOR2 (N944, N943, N647);
buf BUF1 (N945, N911);
or OR3 (N946, N935, N23, N656);
buf BUF1 (N947, N945);
nor NOR3 (N948, N942, N317, N442);
and AND4 (N949, N934, N743, N424, N217);
nor NOR2 (N950, N932, N542);
buf BUF1 (N951, N944);
and AND2 (N952, N951, N717);
buf BUF1 (N953, N940);
and AND3 (N954, N953, N491, N656);
buf BUF1 (N955, N949);
and AND3 (N956, N950, N899, N448);
and AND4 (N957, N894, N674, N768, N35);
not NOT1 (N958, N941);
buf BUF1 (N959, N948);
nor NOR2 (N960, N954, N296);
nand NAND4 (N961, N958, N542, N333, N833);
xor XOR2 (N962, N957, N418);
nand NAND2 (N963, N956, N702);
nand NAND3 (N964, N923, N708, N172);
or OR4 (N965, N962, N320, N144, N423);
nand NAND4 (N966, N965, N556, N775, N608);
and AND2 (N967, N966, N440);
not NOT1 (N968, N961);
nor NOR3 (N969, N955, N118, N428);
buf BUF1 (N970, N946);
not NOT1 (N971, N947);
nor NOR2 (N972, N971, N146);
not NOT1 (N973, N967);
not NOT1 (N974, N969);
xor XOR2 (N975, N970, N78);
and AND2 (N976, N963, N72);
or OR2 (N977, N976, N131);
or OR4 (N978, N972, N960, N235, N946);
and AND2 (N979, N836, N98);
and AND2 (N980, N973, N214);
and AND4 (N981, N980, N277, N97, N57);
buf BUF1 (N982, N978);
nand NAND3 (N983, N975, N453, N264);
xor XOR2 (N984, N979, N96);
and AND2 (N985, N964, N417);
buf BUF1 (N986, N983);
xor XOR2 (N987, N974, N100);
and AND4 (N988, N984, N660, N895, N847);
not NOT1 (N989, N977);
nand NAND3 (N990, N968, N763, N123);
nand NAND4 (N991, N982, N60, N231, N467);
not NOT1 (N992, N985);
xor XOR2 (N993, N990, N603);
or OR2 (N994, N981, N127);
nor NOR2 (N995, N992, N522);
and AND2 (N996, N987, N274);
buf BUF1 (N997, N952);
xor XOR2 (N998, N997, N915);
and AND4 (N999, N989, N336, N900, N250);
buf BUF1 (N1000, N991);
nor NOR4 (N1001, N986, N907, N897, N884);
nor NOR2 (N1002, N999, N960);
or OR2 (N1003, N959, N962);
buf BUF1 (N1004, N996);
nand NAND3 (N1005, N998, N912, N426);
nor NOR2 (N1006, N1001, N63);
or OR4 (N1007, N1004, N155, N612, N145);
or OR3 (N1008, N994, N604, N963);
buf BUF1 (N1009, N1005);
and AND4 (N1010, N1006, N159, N191, N698);
nor NOR4 (N1011, N1010, N785, N964, N438);
or OR2 (N1012, N1000, N498);
xor XOR2 (N1013, N988, N162);
or OR4 (N1014, N1008, N699, N718, N576);
or OR3 (N1015, N1002, N554, N714);
nor NOR3 (N1016, N995, N760, N148);
xor XOR2 (N1017, N1007, N346);
not NOT1 (N1018, N1003);
xor XOR2 (N1019, N1012, N511);
or OR2 (N1020, N1016, N35);
nor NOR4 (N1021, N1020, N121, N119, N805);
xor XOR2 (N1022, N1015, N845);
buf BUF1 (N1023, N1017);
and AND4 (N1024, N1021, N285, N132, N248);
not NOT1 (N1025, N1011);
buf BUF1 (N1026, N1019);
nor NOR2 (N1027, N1014, N257);
xor XOR2 (N1028, N1022, N50);
xor XOR2 (N1029, N1027, N980);
or OR3 (N1030, N1028, N683, N583);
and AND4 (N1031, N1013, N665, N79, N438);
not NOT1 (N1032, N1031);
buf BUF1 (N1033, N1030);
xor XOR2 (N1034, N1023, N537);
and AND4 (N1035, N1029, N563, N690, N76);
nor NOR4 (N1036, N1032, N849, N1004, N870);
buf BUF1 (N1037, N1009);
not NOT1 (N1038, N1026);
or OR4 (N1039, N993, N949, N354, N400);
or OR3 (N1040, N1035, N644, N308);
not NOT1 (N1041, N1037);
not NOT1 (N1042, N1041);
xor XOR2 (N1043, N1033, N1005);
and AND4 (N1044, N1018, N884, N437, N498);
buf BUF1 (N1045, N1039);
or OR2 (N1046, N1043, N469);
or OR4 (N1047, N1045, N330, N456, N39);
nand NAND4 (N1048, N1034, N601, N284, N713);
xor XOR2 (N1049, N1048, N347);
xor XOR2 (N1050, N1038, N499);
not NOT1 (N1051, N1050);
nor NOR3 (N1052, N1025, N264, N932);
or OR3 (N1053, N1046, N569, N579);
or OR4 (N1054, N1040, N123, N510, N602);
or OR3 (N1055, N1053, N511, N680);
not NOT1 (N1056, N1049);
nand NAND2 (N1057, N1044, N567);
xor XOR2 (N1058, N1057, N1020);
and AND3 (N1059, N1036, N347, N834);
nor NOR4 (N1060, N1055, N13, N703, N199);
xor XOR2 (N1061, N1052, N779);
buf BUF1 (N1062, N1060);
xor XOR2 (N1063, N1058, N337);
xor XOR2 (N1064, N1047, N737);
not NOT1 (N1065, N1064);
xor XOR2 (N1066, N1059, N256);
nand NAND2 (N1067, N1063, N138);
buf BUF1 (N1068, N1054);
nor NOR2 (N1069, N1056, N380);
xor XOR2 (N1070, N1061, N814);
and AND4 (N1071, N1051, N334, N951, N122);
nand NAND4 (N1072, N1068, N443, N144, N214);
buf BUF1 (N1073, N1072);
nand NAND3 (N1074, N1067, N666, N646);
not NOT1 (N1075, N1024);
xor XOR2 (N1076, N1042, N853);
nor NOR3 (N1077, N1074, N950, N796);
and AND3 (N1078, N1076, N684, N492);
nand NAND2 (N1079, N1066, N405);
not NOT1 (N1080, N1078);
and AND2 (N1081, N1079, N43);
or OR3 (N1082, N1070, N1029, N1013);
xor XOR2 (N1083, N1069, N480);
not NOT1 (N1084, N1077);
xor XOR2 (N1085, N1071, N924);
buf BUF1 (N1086, N1062);
buf BUF1 (N1087, N1075);
not NOT1 (N1088, N1081);
not NOT1 (N1089, N1073);
not NOT1 (N1090, N1080);
nand NAND2 (N1091, N1084, N759);
nor NOR4 (N1092, N1087, N642, N746, N1003);
buf BUF1 (N1093, N1083);
not NOT1 (N1094, N1082);
buf BUF1 (N1095, N1065);
buf BUF1 (N1096, N1094);
or OR3 (N1097, N1088, N593, N303);
and AND2 (N1098, N1092, N108);
nand NAND4 (N1099, N1090, N826, N327, N1095);
or OR3 (N1100, N1032, N52, N1034);
nand NAND3 (N1101, N1097, N583, N26);
buf BUF1 (N1102, N1096);
xor XOR2 (N1103, N1101, N714);
nor NOR3 (N1104, N1086, N39, N1081);
buf BUF1 (N1105, N1103);
not NOT1 (N1106, N1089);
not NOT1 (N1107, N1093);
xor XOR2 (N1108, N1098, N521);
not NOT1 (N1109, N1085);
nor NOR2 (N1110, N1099, N674);
nor NOR2 (N1111, N1105, N862);
or OR3 (N1112, N1107, N769, N205);
buf BUF1 (N1113, N1108);
or OR3 (N1114, N1110, N695, N688);
or OR4 (N1115, N1113, N173, N910, N839);
and AND4 (N1116, N1104, N669, N165, N221);
nand NAND2 (N1117, N1106, N531);
nand NAND3 (N1118, N1091, N491, N1017);
xor XOR2 (N1119, N1118, N236);
or OR2 (N1120, N1114, N652);
or OR2 (N1121, N1117, N874);
nand NAND3 (N1122, N1116, N440, N700);
and AND4 (N1123, N1120, N128, N278, N736);
nor NOR4 (N1124, N1123, N656, N613, N1053);
nand NAND4 (N1125, N1112, N1051, N451, N491);
or OR3 (N1126, N1121, N1111, N1004);
or OR4 (N1127, N1092, N21, N565, N371);
nor NOR4 (N1128, N1127, N922, N792, N1032);
and AND2 (N1129, N1119, N394);
and AND3 (N1130, N1128, N504, N563);
nand NAND3 (N1131, N1122, N658, N100);
not NOT1 (N1132, N1131);
not NOT1 (N1133, N1100);
not NOT1 (N1134, N1125);
nor NOR2 (N1135, N1102, N287);
buf BUF1 (N1136, N1133);
or OR4 (N1137, N1109, N475, N517, N96);
nand NAND4 (N1138, N1115, N613, N1112, N68);
or OR4 (N1139, N1135, N964, N276, N1032);
nor NOR3 (N1140, N1139, N786, N710);
not NOT1 (N1141, N1129);
and AND4 (N1142, N1130, N456, N819, N935);
xor XOR2 (N1143, N1140, N382);
or OR2 (N1144, N1143, N547);
nor NOR3 (N1145, N1134, N672, N609);
buf BUF1 (N1146, N1142);
buf BUF1 (N1147, N1137);
not NOT1 (N1148, N1141);
or OR2 (N1149, N1145, N183);
buf BUF1 (N1150, N1146);
nand NAND2 (N1151, N1126, N347);
nor NOR4 (N1152, N1132, N306, N237, N1114);
nand NAND3 (N1153, N1136, N662, N84);
buf BUF1 (N1154, N1148);
or OR4 (N1155, N1151, N154, N228, N109);
or OR2 (N1156, N1138, N84);
buf BUF1 (N1157, N1155);
xor XOR2 (N1158, N1124, N123);
or OR3 (N1159, N1158, N1018, N357);
nor NOR3 (N1160, N1156, N81, N205);
nand NAND3 (N1161, N1147, N704, N213);
and AND4 (N1162, N1149, N495, N317, N675);
not NOT1 (N1163, N1153);
not NOT1 (N1164, N1144);
nor NOR3 (N1165, N1164, N710, N316);
xor XOR2 (N1166, N1162, N138);
xor XOR2 (N1167, N1159, N832);
xor XOR2 (N1168, N1160, N535);
and AND3 (N1169, N1152, N624, N640);
or OR3 (N1170, N1163, N586, N796);
or OR3 (N1171, N1166, N726, N1143);
and AND2 (N1172, N1170, N137);
and AND2 (N1173, N1169, N749);
nor NOR3 (N1174, N1167, N1023, N708);
and AND2 (N1175, N1150, N584);
nor NOR2 (N1176, N1173, N370);
xor XOR2 (N1177, N1154, N491);
or OR3 (N1178, N1175, N282, N350);
nor NOR3 (N1179, N1174, N112, N665);
buf BUF1 (N1180, N1172);
not NOT1 (N1181, N1157);
buf BUF1 (N1182, N1165);
not NOT1 (N1183, N1161);
buf BUF1 (N1184, N1180);
nor NOR3 (N1185, N1168, N449, N23);
buf BUF1 (N1186, N1183);
or OR2 (N1187, N1176, N541);
and AND2 (N1188, N1181, N628);
nor NOR3 (N1189, N1179, N510, N1112);
buf BUF1 (N1190, N1184);
not NOT1 (N1191, N1187);
xor XOR2 (N1192, N1190, N843);
nand NAND3 (N1193, N1192, N198, N575);
nand NAND4 (N1194, N1177, N249, N1126, N335);
and AND2 (N1195, N1191, N267);
xor XOR2 (N1196, N1178, N604);
or OR4 (N1197, N1171, N1111, N579, N499);
and AND3 (N1198, N1193, N277, N1147);
not NOT1 (N1199, N1182);
nand NAND2 (N1200, N1198, N426);
not NOT1 (N1201, N1186);
buf BUF1 (N1202, N1197);
not NOT1 (N1203, N1185);
nor NOR4 (N1204, N1195, N528, N966, N265);
not NOT1 (N1205, N1194);
and AND3 (N1206, N1202, N119, N358);
and AND2 (N1207, N1188, N446);
not NOT1 (N1208, N1206);
nor NOR4 (N1209, N1207, N563, N421, N749);
nand NAND3 (N1210, N1208, N437, N475);
nor NOR4 (N1211, N1200, N331, N51, N530);
and AND3 (N1212, N1211, N625, N1024);
buf BUF1 (N1213, N1204);
xor XOR2 (N1214, N1201, N1168);
not NOT1 (N1215, N1209);
xor XOR2 (N1216, N1203, N360);
and AND3 (N1217, N1205, N95, N1134);
nand NAND4 (N1218, N1210, N1094, N411, N1034);
nor NOR3 (N1219, N1215, N672, N1066);
xor XOR2 (N1220, N1218, N544);
not NOT1 (N1221, N1199);
xor XOR2 (N1222, N1196, N422);
not NOT1 (N1223, N1217);
buf BUF1 (N1224, N1216);
not NOT1 (N1225, N1221);
not NOT1 (N1226, N1222);
not NOT1 (N1227, N1214);
buf BUF1 (N1228, N1227);
not NOT1 (N1229, N1213);
or OR3 (N1230, N1228, N996, N826);
or OR3 (N1231, N1223, N571, N1181);
and AND2 (N1232, N1224, N419);
not NOT1 (N1233, N1189);
nor NOR3 (N1234, N1225, N948, N394);
not NOT1 (N1235, N1229);
not NOT1 (N1236, N1232);
nand NAND2 (N1237, N1220, N329);
not NOT1 (N1238, N1233);
nand NAND2 (N1239, N1236, N561);
and AND3 (N1240, N1237, N57, N10);
nor NOR2 (N1241, N1231, N1060);
or OR4 (N1242, N1235, N545, N949, N619);
not NOT1 (N1243, N1212);
and AND2 (N1244, N1234, N1046);
nand NAND4 (N1245, N1230, N904, N663, N939);
nand NAND4 (N1246, N1239, N470, N659, N583);
nand NAND3 (N1247, N1246, N1066, N1219);
buf BUF1 (N1248, N339);
nor NOR3 (N1249, N1226, N35, N12);
nand NAND4 (N1250, N1247, N831, N312, N294);
buf BUF1 (N1251, N1248);
nand NAND4 (N1252, N1240, N1220, N1032, N124);
or OR4 (N1253, N1251, N321, N353, N348);
or OR3 (N1254, N1238, N692, N972);
xor XOR2 (N1255, N1254, N1088);
nor NOR3 (N1256, N1250, N247, N263);
buf BUF1 (N1257, N1241);
buf BUF1 (N1258, N1242);
xor XOR2 (N1259, N1255, N151);
buf BUF1 (N1260, N1259);
and AND2 (N1261, N1244, N852);
not NOT1 (N1262, N1243);
xor XOR2 (N1263, N1260, N214);
or OR4 (N1264, N1258, N522, N514, N556);
xor XOR2 (N1265, N1253, N639);
nor NOR4 (N1266, N1257, N984, N1169, N412);
and AND4 (N1267, N1264, N1151, N820, N1149);
nor NOR4 (N1268, N1261, N1096, N758, N704);
buf BUF1 (N1269, N1252);
and AND4 (N1270, N1263, N790, N797, N455);
buf BUF1 (N1271, N1245);
not NOT1 (N1272, N1266);
not NOT1 (N1273, N1272);
or OR2 (N1274, N1265, N493);
nand NAND2 (N1275, N1249, N212);
nand NAND3 (N1276, N1274, N779, N781);
nor NOR4 (N1277, N1269, N1126, N1159, N436);
nor NOR2 (N1278, N1271, N79);
nand NAND2 (N1279, N1270, N174);
not NOT1 (N1280, N1279);
nand NAND3 (N1281, N1256, N353, N224);
xor XOR2 (N1282, N1280, N384);
nand NAND4 (N1283, N1282, N605, N185, N309);
or OR4 (N1284, N1275, N112, N132, N821);
or OR4 (N1285, N1278, N837, N1011, N215);
nor NOR4 (N1286, N1285, N608, N767, N746);
nor NOR2 (N1287, N1267, N283);
and AND3 (N1288, N1276, N96, N586);
buf BUF1 (N1289, N1281);
not NOT1 (N1290, N1289);
nand NAND2 (N1291, N1288, N1182);
or OR4 (N1292, N1287, N932, N277, N895);
or OR3 (N1293, N1284, N631, N856);
xor XOR2 (N1294, N1262, N439);
and AND3 (N1295, N1291, N55, N1105);
nor NOR4 (N1296, N1277, N1053, N1006, N1147);
or OR3 (N1297, N1294, N310, N1060);
or OR2 (N1298, N1296, N49);
nand NAND4 (N1299, N1283, N72, N730, N1165);
nand NAND2 (N1300, N1293, N102);
or OR4 (N1301, N1286, N621, N294, N249);
nor NOR4 (N1302, N1295, N523, N219, N498);
buf BUF1 (N1303, N1297);
nand NAND2 (N1304, N1302, N1027);
buf BUF1 (N1305, N1301);
nor NOR4 (N1306, N1305, N1067, N921, N922);
or OR3 (N1307, N1306, N196, N360);
nor NOR4 (N1308, N1290, N409, N1076, N1254);
nand NAND3 (N1309, N1304, N1307, N1131);
and AND2 (N1310, N984, N927);
not NOT1 (N1311, N1303);
nand NAND2 (N1312, N1273, N556);
nor NOR2 (N1313, N1268, N917);
and AND2 (N1314, N1309, N768);
and AND4 (N1315, N1308, N668, N319, N682);
buf BUF1 (N1316, N1310);
nor NOR4 (N1317, N1299, N522, N539, N835);
or OR3 (N1318, N1317, N1260, N380);
and AND3 (N1319, N1315, N767, N174);
not NOT1 (N1320, N1313);
buf BUF1 (N1321, N1318);
buf BUF1 (N1322, N1316);
not NOT1 (N1323, N1311);
not NOT1 (N1324, N1298);
nor NOR2 (N1325, N1314, N872);
nor NOR4 (N1326, N1324, N482, N121, N971);
nor NOR3 (N1327, N1325, N1008, N1287);
buf BUF1 (N1328, N1327);
xor XOR2 (N1329, N1322, N687);
not NOT1 (N1330, N1300);
nand NAND4 (N1331, N1323, N291, N432, N232);
xor XOR2 (N1332, N1329, N590);
xor XOR2 (N1333, N1321, N818);
buf BUF1 (N1334, N1331);
and AND3 (N1335, N1332, N934, N460);
xor XOR2 (N1336, N1335, N596);
not NOT1 (N1337, N1320);
xor XOR2 (N1338, N1333, N513);
buf BUF1 (N1339, N1334);
buf BUF1 (N1340, N1312);
xor XOR2 (N1341, N1336, N523);
and AND2 (N1342, N1341, N558);
nand NAND3 (N1343, N1292, N1215, N105);
nand NAND4 (N1344, N1339, N430, N482, N98);
not NOT1 (N1345, N1330);
or OR4 (N1346, N1328, N511, N1185, N1272);
xor XOR2 (N1347, N1345, N356);
buf BUF1 (N1348, N1326);
not NOT1 (N1349, N1348);
buf BUF1 (N1350, N1342);
or OR3 (N1351, N1350, N1039, N1006);
or OR4 (N1352, N1337, N300, N1093, N1262);
not NOT1 (N1353, N1351);
xor XOR2 (N1354, N1353, N57);
nand NAND4 (N1355, N1347, N936, N744, N512);
nor NOR2 (N1356, N1343, N765);
and AND3 (N1357, N1349, N482, N944);
nor NOR4 (N1358, N1346, N77, N922, N957);
or OR2 (N1359, N1340, N930);
not NOT1 (N1360, N1344);
not NOT1 (N1361, N1355);
buf BUF1 (N1362, N1356);
and AND2 (N1363, N1362, N1128);
buf BUF1 (N1364, N1360);
nor NOR4 (N1365, N1354, N1335, N910, N80);
xor XOR2 (N1366, N1352, N360);
not NOT1 (N1367, N1363);
or OR2 (N1368, N1365, N1188);
and AND2 (N1369, N1366, N704);
xor XOR2 (N1370, N1358, N735);
buf BUF1 (N1371, N1319);
nand NAND3 (N1372, N1338, N1214, N485);
xor XOR2 (N1373, N1367, N682);
and AND2 (N1374, N1371, N366);
or OR4 (N1375, N1370, N1248, N99, N424);
nor NOR4 (N1376, N1364, N899, N553, N816);
not NOT1 (N1377, N1361);
buf BUF1 (N1378, N1372);
xor XOR2 (N1379, N1377, N531);
xor XOR2 (N1380, N1374, N626);
or OR3 (N1381, N1357, N412, N794);
buf BUF1 (N1382, N1381);
buf BUF1 (N1383, N1373);
nand NAND3 (N1384, N1359, N673, N143);
not NOT1 (N1385, N1368);
not NOT1 (N1386, N1383);
and AND4 (N1387, N1379, N1226, N1155, N1090);
nand NAND4 (N1388, N1387, N790, N585, N103);
not NOT1 (N1389, N1384);
not NOT1 (N1390, N1382);
nor NOR4 (N1391, N1386, N1218, N529, N162);
xor XOR2 (N1392, N1391, N1290);
nand NAND2 (N1393, N1369, N574);
buf BUF1 (N1394, N1380);
buf BUF1 (N1395, N1389);
not NOT1 (N1396, N1394);
xor XOR2 (N1397, N1378, N652);
not NOT1 (N1398, N1393);
nor NOR3 (N1399, N1376, N104, N952);
xor XOR2 (N1400, N1385, N1095);
or OR3 (N1401, N1397, N35, N1061);
and AND2 (N1402, N1401, N1324);
xor XOR2 (N1403, N1390, N1327);
nand NAND4 (N1404, N1388, N413, N3, N482);
and AND2 (N1405, N1404, N1241);
not NOT1 (N1406, N1375);
nor NOR2 (N1407, N1399, N516);
buf BUF1 (N1408, N1400);
xor XOR2 (N1409, N1406, N119);
or OR2 (N1410, N1395, N607);
buf BUF1 (N1411, N1402);
buf BUF1 (N1412, N1405);
nand NAND2 (N1413, N1396, N73);
not NOT1 (N1414, N1413);
or OR4 (N1415, N1407, N999, N138, N646);
nor NOR4 (N1416, N1392, N735, N79, N385);
buf BUF1 (N1417, N1416);
not NOT1 (N1418, N1412);
or OR2 (N1419, N1415, N114);
nand NAND3 (N1420, N1408, N381, N445);
buf BUF1 (N1421, N1403);
and AND2 (N1422, N1410, N301);
xor XOR2 (N1423, N1421, N351);
or OR3 (N1424, N1398, N268, N781);
or OR4 (N1425, N1419, N337, N1329, N219);
xor XOR2 (N1426, N1417, N429);
xor XOR2 (N1427, N1425, N293);
nand NAND2 (N1428, N1422, N505);
xor XOR2 (N1429, N1423, N574);
buf BUF1 (N1430, N1420);
nor NOR3 (N1431, N1430, N306, N75);
and AND2 (N1432, N1409, N337);
not NOT1 (N1433, N1424);
xor XOR2 (N1434, N1426, N105);
not NOT1 (N1435, N1411);
buf BUF1 (N1436, N1429);
not NOT1 (N1437, N1433);
or OR3 (N1438, N1434, N1057, N423);
or OR2 (N1439, N1431, N1421);
or OR3 (N1440, N1418, N291, N139);
nand NAND4 (N1441, N1414, N1016, N1030, N1102);
not NOT1 (N1442, N1427);
buf BUF1 (N1443, N1438);
nand NAND4 (N1444, N1432, N1330, N835, N760);
xor XOR2 (N1445, N1437, N88);
xor XOR2 (N1446, N1444, N61);
or OR2 (N1447, N1443, N1354);
buf BUF1 (N1448, N1446);
and AND4 (N1449, N1442, N201, N1311, N1391);
and AND2 (N1450, N1447, N679);
not NOT1 (N1451, N1428);
nand NAND4 (N1452, N1449, N29, N209, N326);
xor XOR2 (N1453, N1448, N1387);
and AND3 (N1454, N1450, N574, N1374);
nand NAND2 (N1455, N1436, N1205);
nand NAND4 (N1456, N1453, N1094, N91, N805);
xor XOR2 (N1457, N1456, N1323);
not NOT1 (N1458, N1451);
or OR4 (N1459, N1458, N720, N20, N1313);
and AND3 (N1460, N1440, N199, N236);
nand NAND4 (N1461, N1452, N768, N403, N888);
buf BUF1 (N1462, N1459);
xor XOR2 (N1463, N1457, N281);
or OR2 (N1464, N1462, N797);
nand NAND2 (N1465, N1460, N1429);
and AND3 (N1466, N1463, N260, N37);
and AND4 (N1467, N1435, N1296, N667, N1450);
not NOT1 (N1468, N1441);
or OR3 (N1469, N1461, N650, N815);
xor XOR2 (N1470, N1465, N1373);
and AND2 (N1471, N1454, N1168);
xor XOR2 (N1472, N1464, N667);
nor NOR3 (N1473, N1455, N424, N1065);
xor XOR2 (N1474, N1471, N147);
nor NOR4 (N1475, N1445, N1377, N268, N29);
and AND2 (N1476, N1439, N90);
and AND2 (N1477, N1473, N228);
nand NAND3 (N1478, N1475, N1384, N1377);
not NOT1 (N1479, N1468);
and AND2 (N1480, N1477, N236);
and AND3 (N1481, N1469, N967, N157);
xor XOR2 (N1482, N1481, N1334);
xor XOR2 (N1483, N1467, N304);
nor NOR3 (N1484, N1480, N858, N732);
nand NAND2 (N1485, N1476, N149);
nor NOR4 (N1486, N1483, N225, N1126, N245);
nand NAND3 (N1487, N1479, N955, N1245);
nand NAND4 (N1488, N1472, N337, N909, N1279);
nor NOR2 (N1489, N1487, N921);
xor XOR2 (N1490, N1489, N1087);
nor NOR4 (N1491, N1466, N933, N856, N665);
not NOT1 (N1492, N1491);
buf BUF1 (N1493, N1484);
not NOT1 (N1494, N1493);
not NOT1 (N1495, N1478);
not NOT1 (N1496, N1495);
and AND3 (N1497, N1490, N902, N1372);
or OR3 (N1498, N1496, N407, N408);
xor XOR2 (N1499, N1470, N1147);
buf BUF1 (N1500, N1499);
xor XOR2 (N1501, N1474, N1293);
buf BUF1 (N1502, N1488);
nor NOR3 (N1503, N1482, N521, N701);
not NOT1 (N1504, N1501);
nand NAND2 (N1505, N1494, N560);
xor XOR2 (N1506, N1485, N1109);
or OR3 (N1507, N1498, N1257, N541);
nand NAND4 (N1508, N1497, N1333, N30, N581);
nand NAND3 (N1509, N1492, N1159, N744);
xor XOR2 (N1510, N1503, N183);
or OR4 (N1511, N1510, N596, N544, N44);
nand NAND4 (N1512, N1511, N365, N407, N594);
buf BUF1 (N1513, N1509);
buf BUF1 (N1514, N1513);
nand NAND4 (N1515, N1507, N45, N1279, N621);
or OR4 (N1516, N1502, N870, N180, N1306);
xor XOR2 (N1517, N1504, N33);
xor XOR2 (N1518, N1508, N739);
nand NAND3 (N1519, N1518, N323, N94);
endmodule