// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16;

output N1603,N1599,N1611,N1613,N1597,N1581,N1615,N1610,N1609,N1616;

nor NOR2 (N17, N15, N15);
nor NOR3 (N18, N12, N3, N5);
and AND3 (N19, N17, N18, N9);
buf BUF1 (N20, N17);
nor NOR4 (N21, N14, N5, N1, N2);
buf BUF1 (N22, N20);
nand NAND4 (N23, N11, N7, N9, N11);
buf BUF1 (N24, N16);
nor NOR4 (N25, N18, N6, N4, N7);
buf BUF1 (N26, N16);
or OR2 (N27, N15, N4);
buf BUF1 (N28, N5);
and AND3 (N29, N17, N6, N4);
nand NAND2 (N30, N28, N1);
and AND3 (N31, N30, N28, N22);
and AND3 (N32, N12, N6, N11);
or OR3 (N33, N23, N3, N23);
and AND2 (N34, N25, N1);
or OR2 (N35, N32, N31);
not NOT1 (N36, N7);
nor NOR2 (N37, N29, N14);
buf BUF1 (N38, N27);
and AND4 (N39, N37, N13, N32, N29);
buf BUF1 (N40, N33);
and AND4 (N41, N19, N29, N36, N6);
not NOT1 (N42, N41);
nor NOR4 (N43, N10, N8, N20, N30);
nor NOR3 (N44, N24, N22, N8);
xor XOR2 (N45, N44, N30);
not NOT1 (N46, N43);
nand NAND3 (N47, N46, N17, N28);
nor NOR4 (N48, N47, N31, N47, N28);
buf BUF1 (N49, N34);
not NOT1 (N50, N45);
or OR4 (N51, N35, N46, N2, N49);
not NOT1 (N52, N11);
nand NAND4 (N53, N50, N32, N32, N31);
nand NAND4 (N54, N38, N15, N48, N45);
or OR2 (N55, N41, N32);
buf BUF1 (N56, N54);
buf BUF1 (N57, N26);
buf BUF1 (N58, N57);
not NOT1 (N59, N21);
buf BUF1 (N60, N58);
nand NAND3 (N61, N56, N4, N49);
nand NAND4 (N62, N39, N37, N42, N36);
not NOT1 (N63, N47);
or OR4 (N64, N59, N11, N33, N46);
nand NAND2 (N65, N53, N2);
and AND3 (N66, N65, N2, N59);
or OR2 (N67, N60, N31);
xor XOR2 (N68, N67, N4);
nor NOR3 (N69, N63, N14, N60);
nor NOR3 (N70, N69, N48, N36);
nand NAND4 (N71, N51, N23, N36, N38);
or OR4 (N72, N70, N37, N32, N63);
not NOT1 (N73, N52);
or OR3 (N74, N61, N61, N6);
not NOT1 (N75, N64);
or OR4 (N76, N75, N14, N54, N70);
or OR4 (N77, N72, N70, N53, N43);
nand NAND3 (N78, N62, N74, N51);
not NOT1 (N79, N15);
or OR3 (N80, N79, N43, N75);
not NOT1 (N81, N68);
buf BUF1 (N82, N55);
nor NOR2 (N83, N80, N54);
not NOT1 (N84, N40);
buf BUF1 (N85, N78);
xor XOR2 (N86, N66, N22);
buf BUF1 (N87, N73);
not NOT1 (N88, N87);
buf BUF1 (N89, N84);
or OR2 (N90, N81, N68);
nor NOR2 (N91, N76, N13);
and AND3 (N92, N86, N66, N57);
nor NOR4 (N93, N92, N83, N38, N69);
or OR2 (N94, N91, N8);
xor XOR2 (N95, N47, N11);
nor NOR3 (N96, N77, N80, N30);
and AND2 (N97, N96, N96);
and AND4 (N98, N82, N6, N35, N38);
xor XOR2 (N99, N88, N51);
nor NOR2 (N100, N98, N35);
nand NAND4 (N101, N100, N11, N49, N13);
not NOT1 (N102, N93);
xor XOR2 (N103, N94, N25);
not NOT1 (N104, N99);
not NOT1 (N105, N85);
not NOT1 (N106, N105);
buf BUF1 (N107, N101);
xor XOR2 (N108, N107, N30);
nor NOR4 (N109, N95, N89, N100, N51);
and AND4 (N110, N12, N19, N13, N62);
nor NOR4 (N111, N106, N1, N82, N23);
or OR2 (N112, N90, N106);
nand NAND2 (N113, N108, N92);
not NOT1 (N114, N103);
and AND2 (N115, N97, N102);
nand NAND4 (N116, N103, N113, N36, N88);
buf BUF1 (N117, N74);
nor NOR2 (N118, N112, N88);
or OR2 (N119, N104, N54);
nor NOR3 (N120, N117, N43, N38);
xor XOR2 (N121, N71, N45);
nor NOR3 (N122, N114, N4, N87);
nor NOR2 (N123, N121, N92);
or OR4 (N124, N115, N121, N106, N122);
buf BUF1 (N125, N121);
xor XOR2 (N126, N109, N24);
or OR4 (N127, N126, N50, N87, N114);
not NOT1 (N128, N116);
not NOT1 (N129, N125);
and AND2 (N130, N120, N113);
nor NOR4 (N131, N127, N103, N41, N130);
and AND2 (N132, N6, N78);
or OR2 (N133, N111, N44);
nor NOR2 (N134, N124, N52);
nor NOR4 (N135, N118, N51, N13, N42);
not NOT1 (N136, N119);
xor XOR2 (N137, N135, N1);
or OR4 (N138, N123, N50, N71, N112);
xor XOR2 (N139, N138, N72);
xor XOR2 (N140, N139, N77);
not NOT1 (N141, N129);
not NOT1 (N142, N128);
xor XOR2 (N143, N110, N123);
nand NAND4 (N144, N137, N80, N62, N66);
or OR2 (N145, N143, N103);
not NOT1 (N146, N145);
buf BUF1 (N147, N132);
buf BUF1 (N148, N146);
nor NOR3 (N149, N144, N99, N64);
buf BUF1 (N150, N134);
or OR2 (N151, N141, N145);
nand NAND4 (N152, N136, N142, N119, N44);
nand NAND3 (N153, N131, N54, N143);
buf BUF1 (N154, N32);
buf BUF1 (N155, N133);
or OR3 (N156, N140, N91, N61);
nor NOR3 (N157, N156, N71, N34);
xor XOR2 (N158, N153, N107);
and AND3 (N159, N151, N27, N78);
or OR2 (N160, N155, N157);
not NOT1 (N161, N111);
not NOT1 (N162, N160);
buf BUF1 (N163, N161);
not NOT1 (N164, N158);
xor XOR2 (N165, N149, N142);
buf BUF1 (N166, N163);
and AND4 (N167, N148, N111, N137, N6);
xor XOR2 (N168, N150, N80);
buf BUF1 (N169, N159);
nand NAND3 (N170, N165, N19, N13);
and AND2 (N171, N166, N134);
buf BUF1 (N172, N168);
nor NOR4 (N173, N147, N72, N78, N109);
or OR4 (N174, N171, N71, N123, N165);
not NOT1 (N175, N173);
not NOT1 (N176, N162);
or OR2 (N177, N175, N7);
and AND4 (N178, N176, N31, N157, N117);
nand NAND2 (N179, N164, N86);
not NOT1 (N180, N152);
or OR4 (N181, N167, N171, N50, N107);
and AND2 (N182, N169, N46);
xor XOR2 (N183, N181, N9);
xor XOR2 (N184, N178, N155);
not NOT1 (N185, N180);
or OR4 (N186, N182, N31, N75, N2);
not NOT1 (N187, N179);
buf BUF1 (N188, N174);
nand NAND4 (N189, N184, N155, N1, N29);
or OR3 (N190, N185, N90, N142);
nor NOR3 (N191, N188, N39, N45);
buf BUF1 (N192, N177);
nor NOR2 (N193, N186, N31);
buf BUF1 (N194, N183);
nor NOR3 (N195, N170, N124, N144);
nand NAND4 (N196, N191, N26, N27, N95);
not NOT1 (N197, N189);
and AND3 (N198, N196, N170, N66);
nand NAND2 (N199, N154, N116);
nor NOR2 (N200, N198, N84);
xor XOR2 (N201, N190, N189);
or OR3 (N202, N193, N73, N171);
buf BUF1 (N203, N202);
and AND2 (N204, N194, N52);
nor NOR4 (N205, N200, N60, N19, N36);
xor XOR2 (N206, N187, N184);
nor NOR4 (N207, N172, N145, N59, N159);
or OR4 (N208, N201, N134, N140, N113);
not NOT1 (N209, N192);
not NOT1 (N210, N195);
buf BUF1 (N211, N204);
and AND2 (N212, N206, N147);
xor XOR2 (N213, N209, N201);
not NOT1 (N214, N211);
buf BUF1 (N215, N213);
nor NOR3 (N216, N197, N9, N80);
nor NOR4 (N217, N210, N84, N82, N111);
and AND2 (N218, N207, N91);
nor NOR4 (N219, N203, N18, N86, N208);
not NOT1 (N220, N46);
buf BUF1 (N221, N212);
or OR2 (N222, N217, N41);
and AND3 (N223, N199, N147, N38);
and AND3 (N224, N215, N33, N37);
buf BUF1 (N225, N223);
xor XOR2 (N226, N218, N73);
nor NOR3 (N227, N221, N87, N33);
nand NAND2 (N228, N216, N160);
nand NAND2 (N229, N214, N214);
buf BUF1 (N230, N224);
buf BUF1 (N231, N219);
xor XOR2 (N232, N229, N75);
and AND3 (N233, N231, N197, N171);
xor XOR2 (N234, N220, N198);
buf BUF1 (N235, N234);
nand NAND4 (N236, N228, N212, N85, N46);
xor XOR2 (N237, N225, N151);
xor XOR2 (N238, N236, N58);
and AND2 (N239, N238, N32);
or OR4 (N240, N222, N43, N171, N141);
and AND2 (N241, N205, N142);
not NOT1 (N242, N237);
nor NOR2 (N243, N233, N41);
or OR2 (N244, N239, N180);
nand NAND2 (N245, N242, N169);
nand NAND3 (N246, N230, N125, N148);
or OR4 (N247, N244, N152, N215, N55);
buf BUF1 (N248, N247);
not NOT1 (N249, N246);
or OR2 (N250, N245, N45);
nor NOR2 (N251, N232, N27);
buf BUF1 (N252, N249);
or OR3 (N253, N240, N75, N232);
not NOT1 (N254, N226);
buf BUF1 (N255, N241);
nand NAND4 (N256, N253, N24, N57, N229);
xor XOR2 (N257, N252, N104);
or OR2 (N258, N227, N209);
nor NOR4 (N259, N235, N145, N4, N108);
nand NAND2 (N260, N243, N83);
nand NAND2 (N261, N259, N68);
nand NAND3 (N262, N260, N219, N150);
xor XOR2 (N263, N262, N173);
nor NOR3 (N264, N251, N152, N127);
not NOT1 (N265, N250);
buf BUF1 (N266, N264);
and AND4 (N267, N256, N139, N207, N63);
and AND4 (N268, N257, N99, N144, N45);
not NOT1 (N269, N254);
and AND4 (N270, N265, N249, N181, N252);
and AND2 (N271, N258, N150);
nor NOR2 (N272, N266, N99);
buf BUF1 (N273, N272);
nand NAND3 (N274, N269, N201, N83);
and AND2 (N275, N274, N163);
xor XOR2 (N276, N275, N259);
or OR3 (N277, N267, N106, N103);
nor NOR4 (N278, N261, N222, N192, N155);
buf BUF1 (N279, N268);
nor NOR4 (N280, N273, N107, N263, N265);
not NOT1 (N281, N156);
or OR4 (N282, N276, N3, N143, N50);
nand NAND3 (N283, N280, N98, N153);
or OR2 (N284, N282, N226);
nor NOR4 (N285, N271, N179, N259, N68);
buf BUF1 (N286, N270);
or OR4 (N287, N281, N165, N274, N48);
nor NOR3 (N288, N287, N212, N278);
buf BUF1 (N289, N15);
buf BUF1 (N290, N279);
not NOT1 (N291, N286);
xor XOR2 (N292, N255, N153);
or OR4 (N293, N289, N261, N110, N209);
and AND3 (N294, N291, N179, N110);
xor XOR2 (N295, N285, N153);
xor XOR2 (N296, N288, N133);
or OR4 (N297, N295, N41, N28, N74);
xor XOR2 (N298, N296, N169);
nor NOR3 (N299, N294, N92, N242);
not NOT1 (N300, N293);
or OR2 (N301, N284, N213);
nor NOR3 (N302, N301, N260, N198);
nor NOR2 (N303, N292, N139);
buf BUF1 (N304, N277);
buf BUF1 (N305, N303);
nor NOR4 (N306, N297, N211, N72, N270);
xor XOR2 (N307, N298, N31);
not NOT1 (N308, N306);
and AND3 (N309, N299, N44, N34);
nor NOR4 (N310, N283, N13, N274, N242);
not NOT1 (N311, N305);
xor XOR2 (N312, N309, N137);
nand NAND3 (N313, N300, N223, N213);
and AND3 (N314, N313, N264, N153);
or OR2 (N315, N290, N66);
and AND4 (N316, N314, N142, N207, N249);
nand NAND2 (N317, N302, N123);
nand NAND2 (N318, N310, N180);
nand NAND3 (N319, N317, N163, N222);
and AND4 (N320, N248, N81, N40, N133);
nor NOR3 (N321, N318, N165, N246);
nand NAND4 (N322, N307, N153, N294, N46);
and AND2 (N323, N321, N238);
and AND2 (N324, N320, N45);
nor NOR4 (N325, N304, N50, N112, N75);
or OR2 (N326, N315, N184);
buf BUF1 (N327, N326);
not NOT1 (N328, N308);
and AND2 (N329, N328, N261);
and AND2 (N330, N324, N31);
and AND2 (N331, N322, N58);
buf BUF1 (N332, N316);
buf BUF1 (N333, N312);
buf BUF1 (N334, N319);
not NOT1 (N335, N311);
xor XOR2 (N336, N333, N332);
xor XOR2 (N337, N59, N186);
nor NOR3 (N338, N329, N319, N44);
not NOT1 (N339, N325);
and AND4 (N340, N337, N38, N239, N100);
and AND3 (N341, N339, N188, N250);
buf BUF1 (N342, N341);
and AND4 (N343, N335, N157, N235, N185);
nor NOR4 (N344, N343, N165, N303, N284);
xor XOR2 (N345, N340, N243);
not NOT1 (N346, N331);
and AND4 (N347, N327, N169, N296, N123);
and AND4 (N348, N345, N284, N96, N40);
buf BUF1 (N349, N323);
nand NAND3 (N350, N338, N208, N312);
nor NOR2 (N351, N330, N225);
buf BUF1 (N352, N349);
buf BUF1 (N353, N342);
buf BUF1 (N354, N344);
nor NOR3 (N355, N350, N227, N177);
nor NOR3 (N356, N347, N198, N105);
xor XOR2 (N357, N334, N26);
not NOT1 (N358, N354);
nor NOR3 (N359, N336, N306, N119);
buf BUF1 (N360, N352);
nor NOR2 (N361, N355, N219);
nor NOR2 (N362, N348, N225);
and AND4 (N363, N358, N65, N295, N349);
buf BUF1 (N364, N351);
xor XOR2 (N365, N359, N243);
buf BUF1 (N366, N346);
buf BUF1 (N367, N356);
not NOT1 (N368, N363);
and AND4 (N369, N360, N9, N214, N64);
not NOT1 (N370, N357);
or OR2 (N371, N370, N368);
xor XOR2 (N372, N137, N116);
or OR2 (N373, N367, N246);
and AND4 (N374, N372, N70, N5, N17);
nand NAND4 (N375, N366, N167, N288, N74);
or OR3 (N376, N369, N215, N357);
and AND2 (N377, N361, N178);
xor XOR2 (N378, N374, N82);
and AND4 (N379, N364, N264, N270, N335);
nor NOR3 (N380, N365, N41, N46);
xor XOR2 (N381, N380, N55);
not NOT1 (N382, N373);
xor XOR2 (N383, N377, N51);
not NOT1 (N384, N378);
or OR4 (N385, N383, N113, N334, N235);
not NOT1 (N386, N382);
nand NAND4 (N387, N379, N79, N171, N253);
and AND3 (N388, N384, N243, N7);
and AND3 (N389, N376, N173, N128);
or OR4 (N390, N375, N263, N15, N256);
nor NOR4 (N391, N362, N159, N166, N240);
or OR2 (N392, N381, N319);
nor NOR2 (N393, N389, N250);
and AND2 (N394, N386, N360);
and AND4 (N395, N391, N200, N260, N29);
not NOT1 (N396, N371);
nor NOR2 (N397, N396, N143);
or OR4 (N398, N388, N151, N13, N46);
buf BUF1 (N399, N385);
and AND3 (N400, N395, N314, N52);
xor XOR2 (N401, N387, N267);
buf BUF1 (N402, N400);
buf BUF1 (N403, N393);
and AND3 (N404, N397, N332, N322);
xor XOR2 (N405, N402, N47);
nor NOR4 (N406, N398, N16, N383, N302);
buf BUF1 (N407, N406);
or OR4 (N408, N404, N344, N308, N245);
buf BUF1 (N409, N401);
or OR3 (N410, N390, N245, N202);
not NOT1 (N411, N403);
or OR4 (N412, N399, N238, N389, N3);
or OR2 (N413, N392, N268);
nor NOR3 (N414, N410, N411, N406);
or OR2 (N415, N374, N161);
nand NAND4 (N416, N394, N377, N169, N289);
xor XOR2 (N417, N408, N119);
nor NOR4 (N418, N414, N150, N370, N29);
not NOT1 (N419, N409);
buf BUF1 (N420, N353);
xor XOR2 (N421, N420, N359);
or OR3 (N422, N405, N102, N275);
or OR3 (N423, N421, N58, N70);
xor XOR2 (N424, N417, N289);
nor NOR4 (N425, N423, N345, N196, N250);
nor NOR4 (N426, N416, N313, N305, N69);
nand NAND2 (N427, N426, N106);
nor NOR3 (N428, N422, N50, N425);
or OR2 (N429, N65, N329);
and AND4 (N430, N413, N118, N98, N329);
and AND3 (N431, N429, N162, N224);
not NOT1 (N432, N415);
not NOT1 (N433, N430);
and AND4 (N434, N432, N338, N136, N202);
and AND2 (N435, N407, N417);
nor NOR3 (N436, N418, N87, N127);
nand NAND2 (N437, N431, N196);
not NOT1 (N438, N428);
xor XOR2 (N439, N412, N14);
xor XOR2 (N440, N434, N227);
buf BUF1 (N441, N427);
xor XOR2 (N442, N435, N181);
nand NAND4 (N443, N436, N256, N136, N94);
nand NAND2 (N444, N442, N398);
nand NAND4 (N445, N438, N146, N177, N375);
nor NOR2 (N446, N440, N367);
nand NAND2 (N447, N433, N419);
xor XOR2 (N448, N311, N84);
xor XOR2 (N449, N445, N442);
nand NAND2 (N450, N437, N391);
and AND4 (N451, N441, N217, N427, N29);
nand NAND4 (N452, N449, N191, N63, N391);
xor XOR2 (N453, N452, N451);
nand NAND2 (N454, N31, N311);
xor XOR2 (N455, N447, N271);
or OR2 (N456, N455, N115);
and AND4 (N457, N444, N5, N298, N413);
not NOT1 (N458, N456);
not NOT1 (N459, N454);
and AND4 (N460, N457, N46, N113, N95);
nand NAND4 (N461, N424, N155, N285, N180);
not NOT1 (N462, N439);
xor XOR2 (N463, N458, N137);
buf BUF1 (N464, N460);
buf BUF1 (N465, N464);
xor XOR2 (N466, N448, N289);
xor XOR2 (N467, N450, N356);
xor XOR2 (N468, N461, N9);
and AND2 (N469, N465, N130);
buf BUF1 (N470, N462);
nor NOR2 (N471, N453, N124);
and AND4 (N472, N443, N118, N112, N39);
and AND2 (N473, N446, N311);
nor NOR2 (N474, N473, N81);
nor NOR2 (N475, N474, N35);
not NOT1 (N476, N459);
nand NAND2 (N477, N468, N385);
and AND4 (N478, N469, N23, N405, N340);
or OR3 (N479, N476, N78, N285);
or OR4 (N480, N467, N446, N473, N101);
or OR3 (N481, N480, N355, N302);
nor NOR3 (N482, N477, N257, N442);
not NOT1 (N483, N466);
buf BUF1 (N484, N479);
or OR2 (N485, N482, N410);
and AND3 (N486, N478, N8, N80);
and AND4 (N487, N483, N100, N114, N56);
not NOT1 (N488, N481);
and AND4 (N489, N470, N320, N86, N8);
nor NOR2 (N490, N489, N363);
buf BUF1 (N491, N472);
or OR3 (N492, N471, N2, N150);
nand NAND2 (N493, N463, N36);
xor XOR2 (N494, N490, N116);
nor NOR2 (N495, N484, N112);
buf BUF1 (N496, N492);
or OR4 (N497, N475, N285, N451, N287);
nor NOR4 (N498, N497, N87, N391, N212);
not NOT1 (N499, N485);
and AND3 (N500, N486, N307, N188);
nand NAND4 (N501, N493, N237, N372, N223);
xor XOR2 (N502, N498, N300);
buf BUF1 (N503, N502);
or OR2 (N504, N501, N468);
or OR3 (N505, N494, N148, N315);
or OR2 (N506, N504, N108);
nor NOR3 (N507, N499, N155, N463);
nand NAND2 (N508, N496, N116);
and AND3 (N509, N491, N362, N20);
nor NOR2 (N510, N508, N129);
xor XOR2 (N511, N500, N483);
xor XOR2 (N512, N510, N9);
nand NAND3 (N513, N503, N213, N274);
not NOT1 (N514, N506);
and AND2 (N515, N507, N335);
nor NOR2 (N516, N514, N437);
buf BUF1 (N517, N509);
and AND4 (N518, N488, N241, N43, N322);
nor NOR4 (N519, N511, N88, N468, N110);
nor NOR3 (N520, N487, N119, N115);
nand NAND4 (N521, N505, N278, N485, N484);
or OR4 (N522, N519, N478, N26, N345);
xor XOR2 (N523, N512, N101);
not NOT1 (N524, N518);
not NOT1 (N525, N520);
or OR3 (N526, N525, N14, N343);
nor NOR3 (N527, N516, N305, N468);
buf BUF1 (N528, N495);
and AND3 (N529, N527, N394, N287);
or OR4 (N530, N524, N427, N416, N93);
buf BUF1 (N531, N522);
or OR4 (N532, N521, N309, N394, N72);
xor XOR2 (N533, N523, N14);
xor XOR2 (N534, N513, N224);
nand NAND3 (N535, N528, N203, N484);
or OR4 (N536, N531, N498, N230, N254);
and AND3 (N537, N530, N67, N75);
nand NAND3 (N538, N517, N256, N465);
not NOT1 (N539, N537);
or OR3 (N540, N529, N405, N349);
and AND4 (N541, N536, N476, N142, N274);
xor XOR2 (N542, N539, N160);
nor NOR4 (N543, N538, N536, N2, N71);
nand NAND4 (N544, N532, N102, N337, N106);
nand NAND2 (N545, N544, N401);
nand NAND2 (N546, N533, N474);
nand NAND3 (N547, N543, N141, N125);
and AND2 (N548, N526, N271);
xor XOR2 (N549, N546, N487);
nand NAND4 (N550, N549, N385, N108, N74);
nand NAND3 (N551, N515, N209, N493);
nand NAND2 (N552, N534, N15);
nand NAND3 (N553, N547, N235, N130);
not NOT1 (N554, N548);
nand NAND2 (N555, N553, N52);
or OR2 (N556, N554, N144);
xor XOR2 (N557, N541, N469);
buf BUF1 (N558, N551);
nand NAND4 (N559, N555, N5, N433, N470);
nor NOR3 (N560, N559, N530, N226);
nor NOR3 (N561, N542, N258, N255);
not NOT1 (N562, N535);
buf BUF1 (N563, N560);
or OR2 (N564, N563, N125);
nor NOR4 (N565, N545, N101, N102, N39);
or OR4 (N566, N562, N370, N70, N433);
nand NAND2 (N567, N557, N327);
nand NAND3 (N568, N550, N307, N434);
xor XOR2 (N569, N558, N426);
nor NOR2 (N570, N564, N338);
buf BUF1 (N571, N566);
and AND4 (N572, N556, N21, N312, N49);
nor NOR2 (N573, N570, N320);
not NOT1 (N574, N552);
not NOT1 (N575, N540);
and AND4 (N576, N571, N392, N54, N526);
nand NAND4 (N577, N567, N222, N550, N327);
nor NOR4 (N578, N576, N551, N234, N279);
nand NAND3 (N579, N568, N109, N49);
xor XOR2 (N580, N579, N535);
buf BUF1 (N581, N561);
not NOT1 (N582, N581);
and AND3 (N583, N582, N178, N338);
buf BUF1 (N584, N572);
nor NOR4 (N585, N573, N47, N505, N501);
nor NOR2 (N586, N578, N186);
not NOT1 (N587, N580);
nor NOR3 (N588, N587, N63, N343);
buf BUF1 (N589, N575);
buf BUF1 (N590, N589);
or OR2 (N591, N577, N316);
or OR3 (N592, N565, N226, N337);
and AND2 (N593, N588, N506);
nand NAND3 (N594, N591, N402, N357);
xor XOR2 (N595, N590, N208);
or OR4 (N596, N586, N345, N415, N42);
buf BUF1 (N597, N584);
xor XOR2 (N598, N583, N391);
buf BUF1 (N599, N595);
nor NOR3 (N600, N593, N396, N33);
nor NOR4 (N601, N569, N573, N91, N290);
nand NAND3 (N602, N585, N340, N105);
and AND4 (N603, N592, N263, N374, N428);
and AND2 (N604, N603, N479);
not NOT1 (N605, N574);
xor XOR2 (N606, N596, N535);
xor XOR2 (N607, N601, N510);
not NOT1 (N608, N602);
and AND3 (N609, N599, N140, N2);
not NOT1 (N610, N609);
and AND3 (N611, N608, N475, N305);
xor XOR2 (N612, N606, N424);
nand NAND2 (N613, N607, N457);
and AND3 (N614, N610, N571, N141);
or OR4 (N615, N611, N300, N54, N233);
buf BUF1 (N616, N604);
and AND2 (N617, N615, N229);
and AND3 (N618, N614, N596, N436);
and AND2 (N619, N618, N541);
and AND3 (N620, N616, N335, N125);
xor XOR2 (N621, N612, N482);
buf BUF1 (N622, N613);
and AND4 (N623, N622, N186, N290, N293);
or OR2 (N624, N617, N210);
or OR3 (N625, N619, N130, N434);
nand NAND3 (N626, N624, N586, N363);
buf BUF1 (N627, N621);
nand NAND4 (N628, N623, N67, N481, N461);
xor XOR2 (N629, N597, N368);
xor XOR2 (N630, N620, N582);
or OR2 (N631, N626, N322);
and AND4 (N632, N627, N426, N346, N347);
nand NAND2 (N633, N600, N592);
and AND4 (N634, N630, N231, N452, N477);
nor NOR3 (N635, N633, N253, N620);
xor XOR2 (N636, N631, N111);
and AND2 (N637, N635, N626);
xor XOR2 (N638, N594, N151);
or OR4 (N639, N637, N355, N90, N256);
nand NAND4 (N640, N598, N176, N212, N577);
and AND2 (N641, N605, N376);
or OR2 (N642, N636, N4);
not NOT1 (N643, N628);
or OR4 (N644, N642, N485, N260, N308);
or OR2 (N645, N625, N594);
nor NOR3 (N646, N643, N367, N188);
not NOT1 (N647, N632);
xor XOR2 (N648, N638, N439);
buf BUF1 (N649, N645);
nand NAND2 (N650, N629, N522);
and AND3 (N651, N647, N530, N539);
buf BUF1 (N652, N651);
xor XOR2 (N653, N652, N478);
and AND4 (N654, N650, N608, N316, N114);
xor XOR2 (N655, N641, N343);
or OR4 (N656, N654, N567, N602, N458);
not NOT1 (N657, N634);
nand NAND2 (N658, N640, N341);
or OR4 (N659, N653, N346, N600, N70);
not NOT1 (N660, N655);
or OR2 (N661, N658, N314);
nand NAND3 (N662, N656, N554, N286);
xor XOR2 (N663, N648, N464);
nor NOR3 (N664, N661, N446, N362);
buf BUF1 (N665, N660);
or OR3 (N666, N664, N211, N375);
nand NAND4 (N667, N659, N302, N122, N385);
and AND3 (N668, N649, N479, N428);
xor XOR2 (N669, N667, N447);
and AND2 (N670, N644, N578);
nand NAND2 (N671, N666, N237);
not NOT1 (N672, N657);
not NOT1 (N673, N663);
nand NAND2 (N674, N665, N192);
or OR3 (N675, N670, N412, N405);
and AND3 (N676, N668, N242, N433);
buf BUF1 (N677, N662);
and AND2 (N678, N673, N604);
and AND4 (N679, N672, N452, N17, N654);
nor NOR2 (N680, N639, N12);
not NOT1 (N681, N677);
xor XOR2 (N682, N680, N31);
nor NOR3 (N683, N682, N360, N288);
and AND4 (N684, N683, N168, N412, N8);
or OR3 (N685, N681, N278, N318);
nand NAND3 (N686, N685, N648, N374);
nand NAND3 (N687, N676, N647, N162);
buf BUF1 (N688, N646);
nor NOR3 (N689, N669, N384, N648);
xor XOR2 (N690, N687, N151);
and AND4 (N691, N688, N620, N587, N60);
nand NAND4 (N692, N691, N500, N486, N228);
xor XOR2 (N693, N678, N243);
or OR3 (N694, N690, N163, N561);
xor XOR2 (N695, N692, N33);
nor NOR2 (N696, N689, N557);
nand NAND3 (N697, N675, N317, N204);
buf BUF1 (N698, N695);
buf BUF1 (N699, N671);
not NOT1 (N700, N694);
not NOT1 (N701, N699);
xor XOR2 (N702, N679, N229);
and AND3 (N703, N686, N210, N177);
buf BUF1 (N704, N696);
nand NAND2 (N705, N700, N683);
or OR2 (N706, N693, N540);
xor XOR2 (N707, N702, N302);
not NOT1 (N708, N704);
nand NAND4 (N709, N707, N677, N37, N555);
xor XOR2 (N710, N703, N289);
buf BUF1 (N711, N708);
nor NOR2 (N712, N706, N471);
nor NOR3 (N713, N698, N68, N387);
buf BUF1 (N714, N674);
xor XOR2 (N715, N709, N88);
nand NAND4 (N716, N713, N15, N171, N565);
xor XOR2 (N717, N684, N219);
xor XOR2 (N718, N716, N319);
and AND2 (N719, N711, N500);
nand NAND4 (N720, N718, N111, N718, N328);
and AND2 (N721, N705, N525);
not NOT1 (N722, N721);
not NOT1 (N723, N710);
nor NOR2 (N724, N720, N101);
xor XOR2 (N725, N714, N682);
not NOT1 (N726, N724);
nand NAND4 (N727, N717, N668, N220, N220);
xor XOR2 (N728, N725, N503);
nand NAND2 (N729, N728, N657);
not NOT1 (N730, N719);
and AND3 (N731, N727, N44, N362);
not NOT1 (N732, N726);
nor NOR3 (N733, N697, N701, N420);
or OR2 (N734, N688, N612);
xor XOR2 (N735, N732, N720);
or OR3 (N736, N723, N639, N680);
nand NAND4 (N737, N722, N134, N561, N8);
buf BUF1 (N738, N733);
xor XOR2 (N739, N712, N542);
buf BUF1 (N740, N739);
xor XOR2 (N741, N734, N103);
nor NOR2 (N742, N740, N310);
and AND2 (N743, N737, N261);
or OR4 (N744, N742, N265, N658, N29);
xor XOR2 (N745, N741, N656);
xor XOR2 (N746, N736, N10);
xor XOR2 (N747, N745, N451);
buf BUF1 (N748, N715);
nor NOR4 (N749, N729, N38, N724, N498);
or OR3 (N750, N749, N415, N620);
and AND2 (N751, N747, N545);
nand NAND2 (N752, N730, N611);
not NOT1 (N753, N746);
buf BUF1 (N754, N750);
buf BUF1 (N755, N731);
nand NAND3 (N756, N753, N223, N394);
nor NOR4 (N757, N743, N60, N407, N258);
and AND3 (N758, N752, N588, N8);
or OR2 (N759, N748, N265);
not NOT1 (N760, N751);
nor NOR4 (N761, N755, N389, N326, N247);
not NOT1 (N762, N744);
nand NAND4 (N763, N759, N462, N693, N700);
xor XOR2 (N764, N757, N676);
or OR2 (N765, N763, N164);
buf BUF1 (N766, N765);
xor XOR2 (N767, N738, N207);
buf BUF1 (N768, N761);
and AND3 (N769, N766, N585, N69);
and AND3 (N770, N769, N740, N222);
and AND2 (N771, N760, N231);
and AND4 (N772, N767, N505, N84, N509);
and AND4 (N773, N771, N185, N192, N289);
nand NAND4 (N774, N770, N64, N573, N187);
and AND4 (N775, N774, N560, N426, N78);
xor XOR2 (N776, N754, N98);
nor NOR2 (N777, N758, N51);
buf BUF1 (N778, N756);
not NOT1 (N779, N762);
nand NAND2 (N780, N768, N766);
not NOT1 (N781, N777);
xor XOR2 (N782, N772, N114);
or OR3 (N783, N764, N517, N391);
or OR4 (N784, N779, N590, N564, N547);
buf BUF1 (N785, N783);
not NOT1 (N786, N785);
xor XOR2 (N787, N780, N110);
nand NAND2 (N788, N778, N295);
or OR4 (N789, N775, N741, N353, N179);
nand NAND4 (N790, N788, N343, N520, N560);
not NOT1 (N791, N773);
and AND4 (N792, N790, N403, N447, N597);
and AND4 (N793, N791, N16, N217, N71);
buf BUF1 (N794, N787);
nor NOR3 (N795, N792, N570, N7);
and AND4 (N796, N781, N368, N45, N751);
nor NOR4 (N797, N795, N122, N784, N536);
not NOT1 (N798, N192);
xor XOR2 (N799, N797, N260);
or OR3 (N800, N796, N748, N157);
xor XOR2 (N801, N793, N90);
xor XOR2 (N802, N735, N59);
buf BUF1 (N803, N801);
nand NAND2 (N804, N794, N170);
or OR2 (N805, N786, N67);
nor NOR4 (N806, N789, N697, N804, N666);
nand NAND4 (N807, N47, N504, N576, N337);
xor XOR2 (N808, N806, N261);
buf BUF1 (N809, N799);
buf BUF1 (N810, N807);
nand NAND4 (N811, N810, N105, N296, N625);
xor XOR2 (N812, N800, N612);
xor XOR2 (N813, N802, N141);
nand NAND4 (N814, N803, N291, N639, N191);
not NOT1 (N815, N798);
not NOT1 (N816, N782);
and AND4 (N817, N776, N483, N738, N758);
or OR2 (N818, N812, N678);
xor XOR2 (N819, N813, N142);
buf BUF1 (N820, N819);
or OR3 (N821, N808, N775, N648);
buf BUF1 (N822, N817);
buf BUF1 (N823, N818);
or OR3 (N824, N820, N796, N648);
not NOT1 (N825, N809);
or OR4 (N826, N811, N528, N789, N648);
buf BUF1 (N827, N824);
nor NOR3 (N828, N814, N8, N63);
nor NOR4 (N829, N827, N812, N41, N346);
or OR2 (N830, N823, N721);
nand NAND2 (N831, N822, N62);
nor NOR4 (N832, N830, N277, N656, N48);
and AND3 (N833, N829, N694, N359);
buf BUF1 (N834, N825);
buf BUF1 (N835, N833);
and AND2 (N836, N828, N57);
xor XOR2 (N837, N836, N755);
and AND4 (N838, N832, N147, N274, N133);
xor XOR2 (N839, N821, N575);
not NOT1 (N840, N816);
nand NAND4 (N841, N837, N69, N251, N825);
nand NAND3 (N842, N835, N834, N495);
buf BUF1 (N843, N318);
not NOT1 (N844, N826);
buf BUF1 (N845, N842);
and AND2 (N846, N841, N495);
nor NOR3 (N847, N839, N213, N281);
xor XOR2 (N848, N840, N645);
xor XOR2 (N849, N843, N342);
xor XOR2 (N850, N831, N375);
nand NAND4 (N851, N848, N603, N442, N770);
or OR4 (N852, N847, N791, N387, N391);
not NOT1 (N853, N805);
nor NOR4 (N854, N850, N747, N194, N797);
buf BUF1 (N855, N838);
and AND2 (N856, N854, N717);
or OR2 (N857, N853, N502);
or OR3 (N858, N857, N382, N298);
not NOT1 (N859, N846);
buf BUF1 (N860, N856);
buf BUF1 (N861, N851);
buf BUF1 (N862, N844);
not NOT1 (N863, N858);
nand NAND2 (N864, N849, N94);
not NOT1 (N865, N859);
and AND3 (N866, N864, N375, N699);
buf BUF1 (N867, N863);
not NOT1 (N868, N865);
and AND4 (N869, N861, N503, N428, N639);
or OR3 (N870, N868, N849, N783);
nand NAND3 (N871, N869, N671, N657);
nor NOR2 (N872, N860, N105);
xor XOR2 (N873, N862, N300);
and AND2 (N874, N871, N218);
nand NAND2 (N875, N855, N19);
xor XOR2 (N876, N870, N76);
nand NAND2 (N877, N872, N663);
xor XOR2 (N878, N875, N605);
or OR4 (N879, N874, N779, N157, N547);
not NOT1 (N880, N866);
nor NOR3 (N881, N845, N133, N362);
or OR2 (N882, N878, N50);
not NOT1 (N883, N852);
xor XOR2 (N884, N877, N683);
not NOT1 (N885, N882);
or OR2 (N886, N879, N837);
nor NOR3 (N887, N873, N755, N437);
buf BUF1 (N888, N815);
and AND3 (N889, N881, N393, N547);
or OR4 (N890, N880, N370, N57, N107);
nand NAND3 (N891, N888, N329, N218);
nand NAND3 (N892, N889, N649, N492);
not NOT1 (N893, N883);
xor XOR2 (N894, N867, N822);
or OR3 (N895, N885, N308, N268);
and AND2 (N896, N894, N278);
xor XOR2 (N897, N890, N393);
not NOT1 (N898, N895);
xor XOR2 (N899, N884, N450);
not NOT1 (N900, N899);
nor NOR4 (N901, N897, N152, N495, N703);
and AND4 (N902, N900, N534, N850, N4);
nor NOR3 (N903, N893, N799, N198);
xor XOR2 (N904, N892, N2);
nand NAND4 (N905, N901, N184, N152, N751);
nor NOR4 (N906, N902, N818, N21, N857);
not NOT1 (N907, N876);
not NOT1 (N908, N891);
xor XOR2 (N909, N898, N463);
xor XOR2 (N910, N909, N801);
or OR3 (N911, N907, N312, N285);
nor NOR4 (N912, N896, N566, N676, N481);
not NOT1 (N913, N905);
and AND2 (N914, N910, N384);
nand NAND2 (N915, N904, N885);
buf BUF1 (N916, N912);
nor NOR4 (N917, N908, N198, N513, N559);
nand NAND3 (N918, N916, N864, N663);
nor NOR2 (N919, N914, N652);
or OR4 (N920, N903, N774, N489, N206);
not NOT1 (N921, N911);
nand NAND3 (N922, N886, N473, N302);
not NOT1 (N923, N922);
and AND3 (N924, N919, N592, N831);
buf BUF1 (N925, N913);
nor NOR4 (N926, N923, N211, N646, N336);
and AND2 (N927, N887, N638);
xor XOR2 (N928, N915, N407);
nand NAND3 (N929, N927, N173, N861);
and AND4 (N930, N920, N701, N815, N598);
nand NAND2 (N931, N921, N891);
nand NAND3 (N932, N906, N529, N96);
nor NOR3 (N933, N932, N188, N402);
nor NOR2 (N934, N928, N756);
nor NOR4 (N935, N924, N295, N336, N251);
not NOT1 (N936, N931);
nor NOR2 (N937, N918, N284);
xor XOR2 (N938, N933, N224);
not NOT1 (N939, N917);
and AND3 (N940, N936, N481, N907);
nor NOR2 (N941, N926, N290);
and AND3 (N942, N939, N342, N768);
xor XOR2 (N943, N934, N883);
and AND3 (N944, N940, N11, N494);
not NOT1 (N945, N943);
buf BUF1 (N946, N938);
nand NAND4 (N947, N930, N803, N876, N109);
and AND4 (N948, N942, N702, N907, N259);
and AND4 (N949, N948, N590, N705, N585);
buf BUF1 (N950, N946);
nand NAND2 (N951, N929, N916);
or OR4 (N952, N935, N741, N560, N753);
and AND4 (N953, N945, N478, N314, N492);
nand NAND4 (N954, N952, N316, N695, N494);
xor XOR2 (N955, N953, N944);
nor NOR3 (N956, N501, N593, N548);
and AND4 (N957, N956, N20, N882, N874);
buf BUF1 (N958, N950);
not NOT1 (N959, N955);
and AND4 (N960, N949, N604, N369, N217);
nor NOR4 (N961, N947, N550, N882, N619);
or OR3 (N962, N957, N383, N781);
or OR2 (N963, N961, N955);
and AND3 (N964, N962, N297, N28);
and AND4 (N965, N954, N901, N235, N902);
not NOT1 (N966, N963);
xor XOR2 (N967, N958, N836);
nand NAND4 (N968, N965, N803, N5, N146);
xor XOR2 (N969, N966, N651);
and AND4 (N970, N941, N705, N144, N843);
nand NAND4 (N971, N968, N397, N642, N273);
buf BUF1 (N972, N959);
xor XOR2 (N973, N937, N322);
not NOT1 (N974, N973);
and AND4 (N975, N951, N712, N939, N215);
or OR3 (N976, N972, N93, N787);
buf BUF1 (N977, N974);
not NOT1 (N978, N971);
xor XOR2 (N979, N964, N14);
and AND4 (N980, N976, N400, N204, N779);
buf BUF1 (N981, N980);
and AND4 (N982, N970, N980, N652, N1);
or OR2 (N983, N982, N188);
xor XOR2 (N984, N981, N627);
and AND2 (N985, N975, N150);
and AND3 (N986, N969, N229, N411);
and AND4 (N987, N979, N435, N952, N156);
buf BUF1 (N988, N967);
xor XOR2 (N989, N978, N548);
not NOT1 (N990, N977);
and AND3 (N991, N986, N121, N246);
nor NOR3 (N992, N983, N256, N285);
nand NAND2 (N993, N925, N336);
nand NAND3 (N994, N991, N953, N676);
not NOT1 (N995, N993);
or OR2 (N996, N988, N305);
buf BUF1 (N997, N987);
or OR4 (N998, N960, N862, N644, N453);
and AND4 (N999, N984, N140, N856, N183);
buf BUF1 (N1000, N997);
or OR3 (N1001, N994, N787, N387);
or OR4 (N1002, N999, N987, N85, N341);
xor XOR2 (N1003, N989, N885);
not NOT1 (N1004, N992);
and AND2 (N1005, N998, N113);
not NOT1 (N1006, N1002);
xor XOR2 (N1007, N985, N929);
and AND4 (N1008, N1005, N188, N364, N212);
nand NAND4 (N1009, N995, N737, N742, N910);
nor NOR3 (N1010, N1000, N201, N661);
buf BUF1 (N1011, N1004);
nand NAND2 (N1012, N1008, N38);
or OR2 (N1013, N990, N788);
xor XOR2 (N1014, N1009, N485);
nand NAND3 (N1015, N1003, N845, N881);
nor NOR2 (N1016, N1001, N474);
and AND3 (N1017, N1013, N290, N600);
nand NAND3 (N1018, N1007, N394, N298);
buf BUF1 (N1019, N1006);
nor NOR4 (N1020, N1015, N644, N132, N385);
buf BUF1 (N1021, N1014);
buf BUF1 (N1022, N1012);
or OR2 (N1023, N1010, N504);
nand NAND3 (N1024, N1023, N304, N586);
and AND3 (N1025, N1021, N481, N855);
or OR2 (N1026, N1024, N212);
xor XOR2 (N1027, N1025, N313);
xor XOR2 (N1028, N1022, N140);
and AND3 (N1029, N996, N522, N511);
nor NOR3 (N1030, N1029, N714, N909);
buf BUF1 (N1031, N1016);
nand NAND3 (N1032, N1011, N871, N570);
buf BUF1 (N1033, N1017);
nor NOR3 (N1034, N1030, N848, N683);
and AND3 (N1035, N1034, N9, N826);
nor NOR4 (N1036, N1032, N858, N910, N457);
xor XOR2 (N1037, N1019, N833);
buf BUF1 (N1038, N1018);
nor NOR4 (N1039, N1037, N625, N198, N452);
xor XOR2 (N1040, N1035, N532);
nor NOR3 (N1041, N1038, N1017, N796);
buf BUF1 (N1042, N1031);
and AND3 (N1043, N1027, N419, N600);
nand NAND3 (N1044, N1041, N59, N834);
nor NOR3 (N1045, N1036, N315, N338);
nor NOR4 (N1046, N1033, N521, N280, N95);
or OR2 (N1047, N1020, N629);
or OR4 (N1048, N1039, N450, N642, N1015);
or OR3 (N1049, N1026, N399, N1042);
and AND2 (N1050, N268, N156);
nand NAND2 (N1051, N1047, N857);
or OR2 (N1052, N1050, N130);
nand NAND4 (N1053, N1046, N849, N346, N395);
and AND3 (N1054, N1053, N125, N885);
not NOT1 (N1055, N1051);
nand NAND3 (N1056, N1044, N409, N710);
and AND2 (N1057, N1056, N622);
or OR2 (N1058, N1040, N273);
buf BUF1 (N1059, N1058);
xor XOR2 (N1060, N1054, N550);
buf BUF1 (N1061, N1052);
xor XOR2 (N1062, N1061, N751);
or OR4 (N1063, N1059, N224, N890, N282);
or OR3 (N1064, N1057, N675, N853);
nand NAND4 (N1065, N1062, N797, N657, N632);
nand NAND4 (N1066, N1065, N398, N521, N888);
nor NOR4 (N1067, N1055, N1044, N50, N223);
nor NOR4 (N1068, N1066, N234, N656, N271);
and AND3 (N1069, N1049, N771, N271);
nand NAND3 (N1070, N1048, N672, N679);
not NOT1 (N1071, N1069);
nand NAND2 (N1072, N1071, N890);
nor NOR4 (N1073, N1064, N629, N717, N92);
not NOT1 (N1074, N1067);
or OR2 (N1075, N1070, N656);
xor XOR2 (N1076, N1043, N770);
or OR3 (N1077, N1075, N1056, N129);
nand NAND2 (N1078, N1063, N932);
nor NOR3 (N1079, N1045, N961, N566);
xor XOR2 (N1080, N1073, N1044);
buf BUF1 (N1081, N1076);
or OR4 (N1082, N1081, N1050, N740, N438);
or OR3 (N1083, N1068, N381, N897);
not NOT1 (N1084, N1079);
and AND3 (N1085, N1074, N702, N488);
nor NOR3 (N1086, N1060, N447, N224);
buf BUF1 (N1087, N1077);
and AND3 (N1088, N1085, N622, N847);
or OR3 (N1089, N1082, N528, N481);
not NOT1 (N1090, N1089);
and AND4 (N1091, N1083, N224, N563, N957);
nand NAND4 (N1092, N1088, N961, N563, N764);
nor NOR3 (N1093, N1080, N273, N824);
or OR4 (N1094, N1093, N617, N979, N428);
buf BUF1 (N1095, N1078);
xor XOR2 (N1096, N1095, N940);
buf BUF1 (N1097, N1094);
not NOT1 (N1098, N1087);
or OR3 (N1099, N1092, N1083, N563);
nand NAND2 (N1100, N1097, N1080);
buf BUF1 (N1101, N1099);
not NOT1 (N1102, N1072);
or OR2 (N1103, N1102, N433);
not NOT1 (N1104, N1090);
buf BUF1 (N1105, N1103);
nand NAND4 (N1106, N1091, N883, N586, N873);
or OR3 (N1107, N1100, N831, N124);
or OR4 (N1108, N1104, N1044, N805, N839);
and AND3 (N1109, N1096, N86, N788);
or OR3 (N1110, N1084, N326, N357);
not NOT1 (N1111, N1098);
or OR3 (N1112, N1111, N632, N1000);
buf BUF1 (N1113, N1112);
nor NOR3 (N1114, N1108, N662, N700);
nor NOR2 (N1115, N1105, N334);
not NOT1 (N1116, N1028);
nand NAND2 (N1117, N1115, N1041);
buf BUF1 (N1118, N1113);
not NOT1 (N1119, N1116);
or OR3 (N1120, N1101, N44, N393);
nand NAND2 (N1121, N1109, N516);
nor NOR4 (N1122, N1119, N180, N1030, N378);
and AND3 (N1123, N1107, N1100, N40);
not NOT1 (N1124, N1086);
buf BUF1 (N1125, N1122);
not NOT1 (N1126, N1121);
nor NOR3 (N1127, N1120, N558, N87);
or OR2 (N1128, N1126, N905);
not NOT1 (N1129, N1118);
or OR2 (N1130, N1124, N498);
or OR4 (N1131, N1123, N795, N775, N958);
xor XOR2 (N1132, N1125, N992);
or OR3 (N1133, N1114, N599, N894);
not NOT1 (N1134, N1127);
or OR3 (N1135, N1110, N146, N332);
not NOT1 (N1136, N1132);
nand NAND4 (N1137, N1135, N867, N7, N254);
and AND3 (N1138, N1129, N856, N1079);
buf BUF1 (N1139, N1136);
buf BUF1 (N1140, N1117);
nand NAND4 (N1141, N1128, N389, N783, N88);
or OR3 (N1142, N1139, N103, N119);
or OR2 (N1143, N1131, N127);
buf BUF1 (N1144, N1141);
or OR2 (N1145, N1142, N281);
nand NAND3 (N1146, N1130, N848, N903);
nand NAND3 (N1147, N1146, N485, N353);
or OR2 (N1148, N1144, N1103);
buf BUF1 (N1149, N1143);
buf BUF1 (N1150, N1137);
nor NOR2 (N1151, N1149, N1110);
nand NAND4 (N1152, N1147, N11, N1119, N961);
or OR4 (N1153, N1152, N79, N161, N1111);
xor XOR2 (N1154, N1133, N666);
and AND2 (N1155, N1150, N489);
nand NAND2 (N1156, N1138, N1101);
or OR3 (N1157, N1134, N895, N70);
and AND3 (N1158, N1145, N1045, N887);
and AND4 (N1159, N1154, N886, N865, N845);
nor NOR2 (N1160, N1153, N521);
nand NAND3 (N1161, N1148, N579, N112);
and AND4 (N1162, N1159, N589, N382, N134);
nand NAND4 (N1163, N1158, N961, N523, N793);
nand NAND4 (N1164, N1160, N883, N584, N776);
or OR3 (N1165, N1155, N77, N602);
or OR4 (N1166, N1106, N772, N559, N316);
and AND4 (N1167, N1157, N201, N1134, N58);
xor XOR2 (N1168, N1151, N406);
and AND4 (N1169, N1168, N44, N366, N534);
not NOT1 (N1170, N1167);
and AND2 (N1171, N1166, N819);
not NOT1 (N1172, N1156);
buf BUF1 (N1173, N1165);
or OR2 (N1174, N1163, N497);
xor XOR2 (N1175, N1169, N723);
and AND2 (N1176, N1174, N125);
nor NOR3 (N1177, N1164, N153, N489);
not NOT1 (N1178, N1161);
nor NOR4 (N1179, N1175, N193, N136, N422);
or OR3 (N1180, N1178, N652, N4);
or OR3 (N1181, N1170, N738, N816);
nand NAND3 (N1182, N1162, N554, N311);
buf BUF1 (N1183, N1182);
nand NAND3 (N1184, N1181, N1107, N1055);
buf BUF1 (N1185, N1183);
or OR4 (N1186, N1172, N1086, N1034, N884);
and AND4 (N1187, N1176, N875, N77, N28);
not NOT1 (N1188, N1180);
not NOT1 (N1189, N1179);
not NOT1 (N1190, N1177);
nand NAND2 (N1191, N1171, N960);
not NOT1 (N1192, N1190);
buf BUF1 (N1193, N1186);
buf BUF1 (N1194, N1140);
xor XOR2 (N1195, N1194, N135);
and AND2 (N1196, N1187, N86);
or OR3 (N1197, N1185, N729, N458);
xor XOR2 (N1198, N1173, N446);
buf BUF1 (N1199, N1193);
or OR4 (N1200, N1195, N493, N602, N255);
nor NOR2 (N1201, N1198, N774);
nand NAND4 (N1202, N1201, N693, N767, N246);
or OR4 (N1203, N1197, N847, N991, N856);
nor NOR2 (N1204, N1199, N684);
or OR2 (N1205, N1191, N57);
buf BUF1 (N1206, N1200);
xor XOR2 (N1207, N1202, N162);
or OR2 (N1208, N1189, N683);
buf BUF1 (N1209, N1207);
nand NAND3 (N1210, N1208, N133, N1142);
or OR3 (N1211, N1196, N1152, N1149);
xor XOR2 (N1212, N1211, N370);
nand NAND4 (N1213, N1205, N384, N27, N1092);
and AND4 (N1214, N1204, N181, N284, N402);
nand NAND4 (N1215, N1184, N938, N376, N687);
or OR4 (N1216, N1188, N111, N983, N613);
or OR3 (N1217, N1203, N592, N75);
not NOT1 (N1218, N1214);
not NOT1 (N1219, N1206);
xor XOR2 (N1220, N1213, N962);
and AND2 (N1221, N1210, N132);
nor NOR2 (N1222, N1217, N916);
buf BUF1 (N1223, N1221);
xor XOR2 (N1224, N1212, N860);
buf BUF1 (N1225, N1215);
nor NOR3 (N1226, N1222, N775, N808);
or OR4 (N1227, N1225, N143, N271, N709);
xor XOR2 (N1228, N1220, N898);
or OR2 (N1229, N1226, N511);
or OR4 (N1230, N1224, N1144, N21, N102);
and AND4 (N1231, N1209, N1058, N767, N68);
buf BUF1 (N1232, N1216);
buf BUF1 (N1233, N1219);
buf BUF1 (N1234, N1218);
xor XOR2 (N1235, N1223, N243);
buf BUF1 (N1236, N1227);
and AND4 (N1237, N1231, N301, N1085, N974);
and AND2 (N1238, N1237, N759);
or OR4 (N1239, N1235, N1103, N51, N1177);
and AND4 (N1240, N1234, N882, N41, N572);
or OR3 (N1241, N1236, N894, N318);
buf BUF1 (N1242, N1232);
and AND2 (N1243, N1228, N144);
nand NAND2 (N1244, N1243, N292);
or OR4 (N1245, N1241, N420, N1062, N720);
or OR2 (N1246, N1242, N528);
buf BUF1 (N1247, N1229);
xor XOR2 (N1248, N1240, N866);
nor NOR3 (N1249, N1244, N97, N485);
nand NAND4 (N1250, N1246, N608, N105, N587);
nand NAND3 (N1251, N1230, N789, N152);
xor XOR2 (N1252, N1248, N430);
nor NOR4 (N1253, N1252, N767, N886, N14);
and AND3 (N1254, N1245, N200, N629);
and AND2 (N1255, N1251, N364);
buf BUF1 (N1256, N1192);
not NOT1 (N1257, N1253);
or OR4 (N1258, N1238, N630, N462, N521);
buf BUF1 (N1259, N1249);
xor XOR2 (N1260, N1257, N49);
buf BUF1 (N1261, N1239);
nand NAND2 (N1262, N1233, N1194);
and AND4 (N1263, N1262, N268, N210, N541);
or OR3 (N1264, N1259, N1016, N1106);
and AND4 (N1265, N1258, N1059, N908, N797);
nor NOR3 (N1266, N1263, N986, N561);
buf BUF1 (N1267, N1250);
and AND4 (N1268, N1261, N1148, N151, N469);
nor NOR4 (N1269, N1260, N918, N976, N337);
or OR3 (N1270, N1256, N334, N1024);
not NOT1 (N1271, N1254);
not NOT1 (N1272, N1271);
or OR4 (N1273, N1266, N180, N113, N115);
xor XOR2 (N1274, N1272, N862);
nand NAND4 (N1275, N1274, N111, N71, N375);
and AND2 (N1276, N1268, N942);
not NOT1 (N1277, N1270);
xor XOR2 (N1278, N1275, N922);
and AND4 (N1279, N1255, N286, N189, N607);
not NOT1 (N1280, N1264);
nor NOR2 (N1281, N1273, N363);
nor NOR4 (N1282, N1267, N484, N474, N99);
buf BUF1 (N1283, N1277);
nor NOR4 (N1284, N1279, N848, N515, N925);
nor NOR3 (N1285, N1276, N740, N904);
buf BUF1 (N1286, N1283);
and AND3 (N1287, N1280, N258, N482);
xor XOR2 (N1288, N1281, N1282);
xor XOR2 (N1289, N664, N700);
buf BUF1 (N1290, N1288);
and AND2 (N1291, N1269, N408);
not NOT1 (N1292, N1278);
not NOT1 (N1293, N1286);
and AND3 (N1294, N1293, N632, N755);
nand NAND3 (N1295, N1294, N89, N1240);
buf BUF1 (N1296, N1292);
xor XOR2 (N1297, N1290, N901);
nor NOR2 (N1298, N1287, N110);
xor XOR2 (N1299, N1289, N226);
buf BUF1 (N1300, N1297);
nor NOR2 (N1301, N1265, N439);
and AND2 (N1302, N1291, N47);
or OR2 (N1303, N1302, N376);
and AND4 (N1304, N1298, N1219, N878, N1102);
nor NOR2 (N1305, N1284, N1161);
nand NAND2 (N1306, N1304, N714);
xor XOR2 (N1307, N1247, N381);
xor XOR2 (N1308, N1299, N95);
nand NAND2 (N1309, N1308, N1125);
not NOT1 (N1310, N1285);
not NOT1 (N1311, N1301);
or OR3 (N1312, N1307, N239, N154);
xor XOR2 (N1313, N1309, N47);
buf BUF1 (N1314, N1312);
and AND4 (N1315, N1314, N482, N772, N437);
not NOT1 (N1316, N1311);
xor XOR2 (N1317, N1296, N974);
buf BUF1 (N1318, N1310);
and AND3 (N1319, N1318, N635, N616);
nand NAND3 (N1320, N1295, N511, N532);
and AND4 (N1321, N1300, N781, N21, N142);
and AND3 (N1322, N1315, N362, N199);
nand NAND2 (N1323, N1320, N368);
not NOT1 (N1324, N1321);
buf BUF1 (N1325, N1323);
or OR3 (N1326, N1306, N346, N114);
buf BUF1 (N1327, N1313);
buf BUF1 (N1328, N1326);
or OR3 (N1329, N1316, N378, N497);
nor NOR4 (N1330, N1329, N1216, N941, N681);
or OR2 (N1331, N1325, N381);
not NOT1 (N1332, N1331);
and AND4 (N1333, N1324, N704, N1085, N1126);
not NOT1 (N1334, N1333);
or OR2 (N1335, N1317, N556);
nor NOR2 (N1336, N1330, N715);
nand NAND2 (N1337, N1327, N977);
nor NOR3 (N1338, N1337, N1249, N694);
buf BUF1 (N1339, N1328);
and AND2 (N1340, N1336, N911);
and AND2 (N1341, N1338, N385);
not NOT1 (N1342, N1335);
not NOT1 (N1343, N1341);
buf BUF1 (N1344, N1322);
nand NAND2 (N1345, N1342, N1293);
and AND3 (N1346, N1303, N637, N671);
buf BUF1 (N1347, N1334);
nor NOR3 (N1348, N1319, N132, N480);
xor XOR2 (N1349, N1343, N777);
not NOT1 (N1350, N1340);
nor NOR4 (N1351, N1332, N422, N342, N551);
nand NAND4 (N1352, N1345, N618, N1191, N844);
and AND3 (N1353, N1351, N1186, N499);
nand NAND4 (N1354, N1347, N981, N496, N218);
nor NOR4 (N1355, N1354, N1055, N71, N902);
nand NAND2 (N1356, N1355, N1059);
nor NOR2 (N1357, N1349, N623);
or OR2 (N1358, N1344, N361);
nand NAND4 (N1359, N1339, N973, N1173, N402);
or OR3 (N1360, N1350, N784, N181);
nand NAND4 (N1361, N1352, N1167, N426, N327);
and AND2 (N1362, N1360, N1234);
and AND3 (N1363, N1357, N124, N814);
and AND4 (N1364, N1358, N807, N363, N1280);
nand NAND3 (N1365, N1353, N931, N967);
not NOT1 (N1366, N1362);
xor XOR2 (N1367, N1346, N19);
nand NAND3 (N1368, N1364, N11, N352);
nand NAND3 (N1369, N1348, N1226, N385);
buf BUF1 (N1370, N1356);
and AND4 (N1371, N1305, N515, N154, N831);
xor XOR2 (N1372, N1365, N402);
and AND3 (N1373, N1371, N555, N835);
or OR4 (N1374, N1359, N928, N1258, N664);
not NOT1 (N1375, N1366);
nor NOR3 (N1376, N1369, N918, N233);
not NOT1 (N1377, N1368);
or OR4 (N1378, N1377, N444, N713, N2);
nand NAND4 (N1379, N1367, N1016, N844, N1197);
nor NOR3 (N1380, N1373, N874, N337);
xor XOR2 (N1381, N1376, N361);
xor XOR2 (N1382, N1375, N1206);
and AND4 (N1383, N1372, N1128, N1018, N857);
nand NAND3 (N1384, N1378, N406, N912);
xor XOR2 (N1385, N1382, N125);
or OR2 (N1386, N1370, N1012);
nand NAND2 (N1387, N1361, N630);
nor NOR2 (N1388, N1385, N1361);
and AND2 (N1389, N1388, N339);
nand NAND4 (N1390, N1389, N951, N716, N270);
and AND3 (N1391, N1384, N460, N647);
buf BUF1 (N1392, N1380);
and AND2 (N1393, N1386, N237);
buf BUF1 (N1394, N1393);
nor NOR2 (N1395, N1392, N117);
or OR2 (N1396, N1381, N419);
nand NAND2 (N1397, N1390, N735);
not NOT1 (N1398, N1396);
not NOT1 (N1399, N1391);
or OR3 (N1400, N1395, N624, N1025);
nor NOR4 (N1401, N1374, N1144, N620, N4);
xor XOR2 (N1402, N1394, N766);
buf BUF1 (N1403, N1397);
and AND3 (N1404, N1387, N1029, N1171);
xor XOR2 (N1405, N1401, N925);
buf BUF1 (N1406, N1404);
xor XOR2 (N1407, N1399, N366);
xor XOR2 (N1408, N1405, N382);
or OR2 (N1409, N1408, N1262);
and AND2 (N1410, N1383, N1180);
or OR4 (N1411, N1400, N651, N441, N1127);
buf BUF1 (N1412, N1407);
not NOT1 (N1413, N1403);
not NOT1 (N1414, N1363);
or OR2 (N1415, N1414, N446);
or OR2 (N1416, N1415, N962);
or OR3 (N1417, N1379, N203, N458);
or OR3 (N1418, N1409, N970, N409);
and AND3 (N1419, N1416, N808, N1321);
nor NOR4 (N1420, N1418, N382, N652, N847);
or OR3 (N1421, N1419, N861, N1381);
buf BUF1 (N1422, N1417);
nor NOR3 (N1423, N1398, N962, N694);
not NOT1 (N1424, N1421);
not NOT1 (N1425, N1423);
nand NAND3 (N1426, N1411, N1185, N356);
not NOT1 (N1427, N1406);
nand NAND2 (N1428, N1412, N1226);
not NOT1 (N1429, N1410);
nor NOR2 (N1430, N1424, N939);
nand NAND4 (N1431, N1427, N1001, N1182, N182);
xor XOR2 (N1432, N1430, N1327);
nor NOR4 (N1433, N1422, N928, N1281, N1178);
and AND4 (N1434, N1433, N1222, N739, N613);
nor NOR3 (N1435, N1420, N1214, N1075);
xor XOR2 (N1436, N1413, N211);
nand NAND2 (N1437, N1426, N169);
or OR3 (N1438, N1432, N939, N1257);
buf BUF1 (N1439, N1425);
or OR4 (N1440, N1434, N1268, N11, N300);
buf BUF1 (N1441, N1439);
nand NAND2 (N1442, N1402, N1405);
xor XOR2 (N1443, N1428, N488);
and AND3 (N1444, N1436, N1252, N1132);
nor NOR3 (N1445, N1442, N1361, N186);
buf BUF1 (N1446, N1438);
and AND3 (N1447, N1446, N829, N436);
buf BUF1 (N1448, N1441);
or OR4 (N1449, N1437, N481, N1420, N975);
xor XOR2 (N1450, N1443, N856);
not NOT1 (N1451, N1449);
not NOT1 (N1452, N1447);
and AND4 (N1453, N1429, N1400, N134, N1300);
nor NOR3 (N1454, N1451, N739, N790);
nor NOR2 (N1455, N1431, N324);
nor NOR4 (N1456, N1440, N365, N1437, N391);
or OR3 (N1457, N1455, N514, N1043);
xor XOR2 (N1458, N1453, N634);
xor XOR2 (N1459, N1456, N754);
and AND3 (N1460, N1457, N530, N921);
and AND2 (N1461, N1454, N18);
and AND4 (N1462, N1452, N94, N1368, N500);
buf BUF1 (N1463, N1448);
or OR4 (N1464, N1462, N1095, N472, N622);
nor NOR2 (N1465, N1435, N516);
and AND2 (N1466, N1464, N1411);
nor NOR3 (N1467, N1461, N794, N572);
buf BUF1 (N1468, N1460);
or OR4 (N1469, N1463, N897, N320, N357);
nand NAND3 (N1470, N1465, N521, N97);
buf BUF1 (N1471, N1467);
nand NAND2 (N1472, N1458, N1245);
xor XOR2 (N1473, N1472, N478);
and AND2 (N1474, N1469, N633);
buf BUF1 (N1475, N1471);
and AND2 (N1476, N1470, N595);
or OR2 (N1477, N1459, N164);
buf BUF1 (N1478, N1473);
xor XOR2 (N1479, N1476, N1433);
or OR3 (N1480, N1444, N817, N400);
xor XOR2 (N1481, N1474, N1350);
buf BUF1 (N1482, N1478);
xor XOR2 (N1483, N1477, N1430);
xor XOR2 (N1484, N1479, N434);
nand NAND3 (N1485, N1483, N188, N342);
nand NAND2 (N1486, N1475, N700);
buf BUF1 (N1487, N1445);
nand NAND4 (N1488, N1484, N1482, N1072, N287);
nand NAND4 (N1489, N720, N1204, N425, N1165);
and AND2 (N1490, N1481, N597);
and AND2 (N1491, N1490, N340);
nand NAND3 (N1492, N1450, N1169, N180);
nand NAND4 (N1493, N1468, N806, N268, N1458);
nand NAND2 (N1494, N1485, N403);
nand NAND2 (N1495, N1489, N384);
buf BUF1 (N1496, N1486);
nand NAND3 (N1497, N1493, N1173, N64);
not NOT1 (N1498, N1494);
nand NAND4 (N1499, N1480, N1061, N1273, N868);
buf BUF1 (N1500, N1499);
or OR3 (N1501, N1498, N1199, N495);
nand NAND4 (N1502, N1501, N685, N634, N1292);
or OR4 (N1503, N1495, N1347, N775, N1137);
or OR3 (N1504, N1503, N790, N162);
or OR4 (N1505, N1487, N1481, N993, N896);
and AND4 (N1506, N1488, N554, N844, N652);
not NOT1 (N1507, N1505);
nand NAND2 (N1508, N1491, N628);
or OR4 (N1509, N1500, N814, N171, N105);
nand NAND2 (N1510, N1509, N66);
nor NOR4 (N1511, N1506, N160, N120, N249);
or OR4 (N1512, N1507, N85, N1373, N60);
or OR3 (N1513, N1497, N761, N368);
buf BUF1 (N1514, N1508);
nand NAND2 (N1515, N1492, N54);
not NOT1 (N1516, N1513);
nor NOR2 (N1517, N1511, N374);
buf BUF1 (N1518, N1466);
or OR2 (N1519, N1516, N661);
xor XOR2 (N1520, N1512, N795);
xor XOR2 (N1521, N1510, N193);
nand NAND4 (N1522, N1521, N313, N435, N316);
xor XOR2 (N1523, N1518, N84);
buf BUF1 (N1524, N1514);
nand NAND2 (N1525, N1524, N480);
not NOT1 (N1526, N1519);
xor XOR2 (N1527, N1502, N863);
not NOT1 (N1528, N1496);
buf BUF1 (N1529, N1515);
or OR4 (N1530, N1517, N349, N1024, N459);
and AND4 (N1531, N1525, N826, N2, N57);
buf BUF1 (N1532, N1527);
buf BUF1 (N1533, N1526);
buf BUF1 (N1534, N1528);
buf BUF1 (N1535, N1523);
nand NAND3 (N1536, N1504, N1040, N1036);
buf BUF1 (N1537, N1520);
nand NAND3 (N1538, N1534, N1180, N1043);
nand NAND2 (N1539, N1522, N1334);
xor XOR2 (N1540, N1536, N434);
nand NAND2 (N1541, N1531, N1077);
or OR4 (N1542, N1540, N1173, N558, N649);
nor NOR4 (N1543, N1537, N219, N1401, N946);
nor NOR4 (N1544, N1542, N1486, N28, N914);
xor XOR2 (N1545, N1535, N481);
nand NAND3 (N1546, N1543, N1515, N850);
buf BUF1 (N1547, N1539);
not NOT1 (N1548, N1541);
and AND4 (N1549, N1530, N709, N612, N477);
or OR3 (N1550, N1538, N841, N831);
not NOT1 (N1551, N1533);
nand NAND3 (N1552, N1549, N1044, N363);
xor XOR2 (N1553, N1529, N718);
buf BUF1 (N1554, N1551);
not NOT1 (N1555, N1553);
nor NOR2 (N1556, N1550, N1438);
nor NOR2 (N1557, N1547, N1332);
nor NOR4 (N1558, N1548, N649, N1157, N686);
nor NOR4 (N1559, N1532, N326, N1118, N791);
nor NOR4 (N1560, N1552, N904, N1519, N1477);
or OR4 (N1561, N1558, N759, N1333, N1295);
nand NAND4 (N1562, N1561, N195, N248, N682);
xor XOR2 (N1563, N1557, N110);
buf BUF1 (N1564, N1554);
and AND2 (N1565, N1560, N161);
or OR2 (N1566, N1555, N1535);
or OR2 (N1567, N1556, N220);
and AND2 (N1568, N1566, N454);
nand NAND3 (N1569, N1559, N758, N346);
nand NAND4 (N1570, N1565, N291, N1185, N449);
buf BUF1 (N1571, N1545);
nor NOR4 (N1572, N1569, N252, N71, N1191);
nor NOR2 (N1573, N1544, N300);
nor NOR2 (N1574, N1568, N1435);
and AND3 (N1575, N1571, N434, N1311);
xor XOR2 (N1576, N1572, N745);
or OR3 (N1577, N1564, N1427, N936);
not NOT1 (N1578, N1570);
not NOT1 (N1579, N1573);
nand NAND3 (N1580, N1579, N1169, N1546);
xor XOR2 (N1581, N1335, N1510);
nand NAND3 (N1582, N1563, N1462, N1509);
nor NOR4 (N1583, N1567, N643, N1270, N960);
buf BUF1 (N1584, N1577);
nand NAND3 (N1585, N1574, N965, N1571);
xor XOR2 (N1586, N1578, N715);
buf BUF1 (N1587, N1562);
or OR3 (N1588, N1587, N486, N1055);
and AND3 (N1589, N1588, N1261, N468);
xor XOR2 (N1590, N1584, N300);
xor XOR2 (N1591, N1589, N670);
or OR4 (N1592, N1583, N272, N1264, N480);
and AND2 (N1593, N1592, N27);
or OR3 (N1594, N1575, N964, N908);
nor NOR2 (N1595, N1582, N1490);
nor NOR2 (N1596, N1585, N646);
xor XOR2 (N1597, N1593, N1090);
nor NOR2 (N1598, N1591, N1027);
not NOT1 (N1599, N1580);
xor XOR2 (N1600, N1590, N472);
buf BUF1 (N1601, N1598);
and AND2 (N1602, N1595, N347);
not NOT1 (N1603, N1601);
nand NAND4 (N1604, N1586, N1340, N218, N1396);
nand NAND2 (N1605, N1604, N1087);
and AND4 (N1606, N1605, N874, N1004, N1095);
nor NOR2 (N1607, N1576, N433);
nor NOR3 (N1608, N1594, N300, N366);
or OR2 (N1609, N1606, N1233);
buf BUF1 (N1610, N1600);
nor NOR2 (N1611, N1596, N379);
buf BUF1 (N1612, N1608);
nor NOR2 (N1613, N1607, N1297);
not NOT1 (N1614, N1602);
nor NOR4 (N1615, N1612, N380, N1166, N1113);
or OR3 (N1616, N1614, N353, N238);
endmodule