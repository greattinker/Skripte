// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22;

output N203,N210,N209,N221,N215,N216,N207,N214,N220,N222;

nand NAND4 (N23, N3, N19, N20, N17);
nand NAND4 (N24, N20, N2, N8, N21);
xor XOR2 (N25, N4, N13);
and AND4 (N26, N12, N7, N21, N20);
buf BUF1 (N27, N16);
not NOT1 (N28, N22);
nor NOR4 (N29, N20, N10, N21, N18);
nand NAND4 (N30, N21, N7, N24, N6);
nand NAND4 (N31, N13, N16, N15, N25);
or OR3 (N32, N16, N29, N23);
buf BUF1 (N33, N12);
xor XOR2 (N34, N19, N19);
or OR3 (N35, N21, N13, N14);
not NOT1 (N36, N6);
or OR3 (N37, N34, N35, N26);
and AND2 (N38, N2, N6);
xor XOR2 (N39, N29, N31);
buf BUF1 (N40, N2);
buf BUF1 (N41, N39);
nand NAND3 (N42, N33, N29, N5);
and AND4 (N43, N30, N11, N3, N19);
and AND3 (N44, N42, N3, N27);
xor XOR2 (N45, N11, N15);
xor XOR2 (N46, N41, N45);
nand NAND2 (N47, N43, N34);
buf BUF1 (N48, N8);
buf BUF1 (N49, N48);
and AND3 (N50, N46, N45, N28);
nor NOR4 (N51, N4, N11, N26, N36);
and AND2 (N52, N50, N4);
nor NOR3 (N53, N20, N11, N49);
xor XOR2 (N54, N37, N51);
xor XOR2 (N55, N31, N39);
buf BUF1 (N56, N22);
xor XOR2 (N57, N55, N19);
nor NOR3 (N58, N47, N46, N29);
xor XOR2 (N59, N52, N24);
nor NOR3 (N60, N59, N18, N4);
and AND2 (N61, N40, N14);
and AND3 (N62, N60, N33, N40);
buf BUF1 (N63, N62);
and AND2 (N64, N57, N11);
and AND3 (N65, N54, N45, N32);
or OR2 (N66, N7, N34);
not NOT1 (N67, N44);
or OR4 (N68, N53, N25, N11, N38);
xor XOR2 (N69, N25, N58);
nand NAND3 (N70, N19, N16, N6);
nand NAND2 (N71, N66, N57);
nor NOR2 (N72, N61, N7);
or OR2 (N73, N68, N56);
nor NOR4 (N74, N30, N47, N44, N64);
nand NAND3 (N75, N40, N1, N30);
not NOT1 (N76, N74);
not NOT1 (N77, N75);
buf BUF1 (N78, N72);
not NOT1 (N79, N65);
and AND3 (N80, N70, N16, N55);
not NOT1 (N81, N67);
nor NOR2 (N82, N81, N29);
not NOT1 (N83, N76);
nand NAND4 (N84, N77, N30, N29, N10);
nand NAND4 (N85, N82, N29, N74, N79);
buf BUF1 (N86, N27);
nand NAND4 (N87, N78, N77, N45, N39);
not NOT1 (N88, N85);
nor NOR4 (N89, N87, N6, N58, N29);
xor XOR2 (N90, N89, N71);
xor XOR2 (N91, N16, N11);
not NOT1 (N92, N88);
not NOT1 (N93, N69);
not NOT1 (N94, N80);
or OR3 (N95, N92, N57, N6);
nand NAND2 (N96, N84, N75);
and AND2 (N97, N91, N34);
buf BUF1 (N98, N90);
xor XOR2 (N99, N97, N52);
not NOT1 (N100, N93);
nand NAND2 (N101, N83, N20);
xor XOR2 (N102, N96, N95);
or OR4 (N103, N55, N102, N84, N60);
not NOT1 (N104, N79);
and AND4 (N105, N73, N44, N54, N40);
nor NOR3 (N106, N103, N74, N44);
buf BUF1 (N107, N101);
xor XOR2 (N108, N100, N78);
buf BUF1 (N109, N98);
xor XOR2 (N110, N106, N54);
and AND4 (N111, N104, N98, N29, N99);
xor XOR2 (N112, N3, N106);
nor NOR3 (N113, N94, N54, N111);
nor NOR2 (N114, N47, N75);
buf BUF1 (N115, N86);
or OR2 (N116, N108, N42);
and AND2 (N117, N113, N75);
or OR3 (N118, N63, N25, N30);
not NOT1 (N119, N109);
or OR2 (N120, N105, N98);
nand NAND4 (N121, N115, N48, N6, N73);
and AND2 (N122, N117, N16);
buf BUF1 (N123, N120);
xor XOR2 (N124, N121, N64);
nand NAND4 (N125, N119, N70, N100, N73);
nor NOR3 (N126, N116, N54, N2);
nand NAND3 (N127, N123, N62, N35);
or OR2 (N128, N112, N64);
and AND2 (N129, N124, N63);
and AND2 (N130, N114, N81);
nand NAND3 (N131, N127, N99, N51);
buf BUF1 (N132, N107);
buf BUF1 (N133, N129);
buf BUF1 (N134, N110);
nor NOR4 (N135, N126, N63, N40, N107);
and AND3 (N136, N132, N135, N32);
nand NAND3 (N137, N124, N58, N18);
not NOT1 (N138, N130);
not NOT1 (N139, N125);
nor NOR3 (N140, N138, N72, N107);
nor NOR3 (N141, N139, N55, N22);
nand NAND3 (N142, N133, N130, N93);
xor XOR2 (N143, N128, N37);
not NOT1 (N144, N122);
or OR3 (N145, N136, N129, N37);
and AND2 (N146, N142, N80);
nor NOR4 (N147, N137, N131, N117, N65);
buf BUF1 (N148, N77);
buf BUF1 (N149, N141);
xor XOR2 (N150, N148, N61);
and AND2 (N151, N118, N17);
not NOT1 (N152, N151);
nand NAND2 (N153, N145, N45);
nor NOR4 (N154, N153, N44, N141, N93);
xor XOR2 (N155, N143, N121);
and AND4 (N156, N149, N136, N32, N2);
or OR3 (N157, N140, N37, N146);
nor NOR2 (N158, N62, N12);
nand NAND3 (N159, N134, N50, N135);
xor XOR2 (N160, N157, N118);
and AND3 (N161, N144, N105, N47);
nand NAND4 (N162, N161, N101, N132, N43);
nand NAND3 (N163, N162, N47, N66);
nor NOR3 (N164, N159, N52, N31);
or OR4 (N165, N160, N9, N61, N47);
xor XOR2 (N166, N152, N118);
buf BUF1 (N167, N154);
nand NAND2 (N168, N158, N124);
buf BUF1 (N169, N163);
buf BUF1 (N170, N166);
or OR4 (N171, N164, N139, N168, N2);
not NOT1 (N172, N89);
buf BUF1 (N173, N155);
and AND2 (N174, N172, N149);
buf BUF1 (N175, N174);
buf BUF1 (N176, N165);
nand NAND3 (N177, N171, N53, N160);
and AND2 (N178, N169, N170);
not NOT1 (N179, N137);
buf BUF1 (N180, N156);
or OR2 (N181, N147, N176);
or OR3 (N182, N55, N30, N152);
or OR2 (N183, N178, N100);
and AND4 (N184, N181, N56, N65, N103);
nand NAND4 (N185, N167, N7, N22, N159);
xor XOR2 (N186, N175, N37);
nand NAND2 (N187, N184, N136);
xor XOR2 (N188, N185, N173);
or OR3 (N189, N121, N93, N30);
xor XOR2 (N190, N187, N150);
or OR3 (N191, N81, N57, N104);
nor NOR3 (N192, N191, N166, N72);
nor NOR2 (N193, N189, N58);
or OR3 (N194, N190, N31, N3);
not NOT1 (N195, N177);
buf BUF1 (N196, N183);
not NOT1 (N197, N192);
or OR4 (N198, N182, N173, N180, N159);
xor XOR2 (N199, N106, N91);
buf BUF1 (N200, N186);
not NOT1 (N201, N200);
not NOT1 (N202, N195);
or OR3 (N203, N201, N121, N162);
xor XOR2 (N204, N194, N49);
xor XOR2 (N205, N204, N99);
or OR3 (N206, N205, N199, N205);
buf BUF1 (N207, N161);
not NOT1 (N208, N202);
xor XOR2 (N209, N208, N50);
and AND3 (N210, N188, N65, N101);
not NOT1 (N211, N206);
nand NAND2 (N212, N197, N47);
buf BUF1 (N213, N193);
and AND3 (N214, N212, N120, N134);
xor XOR2 (N215, N198, N131);
nand NAND2 (N216, N179, N180);
and AND2 (N217, N211, N173);
nor NOR3 (N218, N217, N135, N205);
not NOT1 (N219, N213);
xor XOR2 (N220, N218, N174);
nor NOR4 (N221, N219, N37, N5, N176);
or OR4 (N222, N196, N126, N99, N160);
endmodule