// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20;

output N8012,N8005,N7984,N8017,N8018,N8010,N8011,N8019,N7981,N8020;

nor NOR2 (N21, N8, N16);
not NOT1 (N22, N20);
and AND4 (N23, N14, N18, N13, N7);
not NOT1 (N24, N2);
xor XOR2 (N25, N22, N19);
nor NOR4 (N26, N21, N16, N21, N14);
xor XOR2 (N27, N8, N12);
nand NAND2 (N28, N14, N9);
or OR2 (N29, N25, N4);
nor NOR4 (N30, N4, N24, N5, N10);
nand NAND3 (N31, N17, N11, N17);
buf BUF1 (N32, N31);
not NOT1 (N33, N31);
or OR2 (N34, N8, N26);
nor NOR3 (N35, N26, N17, N18);
nor NOR2 (N36, N12, N21);
nor NOR3 (N37, N32, N17, N23);
or OR3 (N38, N27, N15, N15);
xor XOR2 (N39, N2, N23);
or OR4 (N40, N36, N16, N26, N10);
and AND4 (N41, N38, N22, N38, N37);
or OR3 (N42, N15, N5, N6);
nand NAND4 (N43, N33, N41, N19, N34);
xor XOR2 (N44, N22, N26);
not NOT1 (N45, N23);
nand NAND4 (N46, N30, N37, N33, N22);
xor XOR2 (N47, N42, N20);
xor XOR2 (N48, N44, N10);
nor NOR4 (N49, N28, N37, N20, N15);
buf BUF1 (N50, N49);
nor NOR3 (N51, N29, N35, N23);
nor NOR2 (N52, N45, N7);
not NOT1 (N53, N16);
nor NOR3 (N54, N40, N49, N47);
nor NOR2 (N55, N19, N38);
or OR2 (N56, N50, N12);
and AND2 (N57, N52, N23);
nor NOR3 (N58, N53, N17, N47);
xor XOR2 (N59, N46, N41);
not NOT1 (N60, N54);
xor XOR2 (N61, N43, N22);
nand NAND4 (N62, N48, N29, N20, N19);
not NOT1 (N63, N59);
buf BUF1 (N64, N60);
xor XOR2 (N65, N39, N16);
xor XOR2 (N66, N57, N45);
xor XOR2 (N67, N51, N11);
not NOT1 (N68, N55);
and AND2 (N69, N64, N16);
or OR4 (N70, N65, N58, N64, N16);
and AND3 (N71, N52, N58, N55);
not NOT1 (N72, N70);
not NOT1 (N73, N67);
nand NAND3 (N74, N73, N28, N40);
nor NOR3 (N75, N68, N47, N36);
and AND2 (N76, N71, N32);
buf BUF1 (N77, N63);
buf BUF1 (N78, N77);
nor NOR4 (N79, N72, N48, N10, N39);
or OR2 (N80, N74, N45);
buf BUF1 (N81, N56);
nand NAND3 (N82, N75, N7, N56);
not NOT1 (N83, N78);
xor XOR2 (N84, N83, N16);
or OR4 (N85, N84, N11, N31, N3);
or OR2 (N86, N62, N77);
nor NOR4 (N87, N82, N79, N35, N3);
or OR4 (N88, N2, N23, N74, N47);
nand NAND4 (N89, N81, N61, N86, N51);
nand NAND3 (N90, N50, N1, N37);
nand NAND4 (N91, N90, N33, N8, N38);
or OR2 (N92, N3, N31);
or OR3 (N93, N92, N59, N80);
not NOT1 (N94, N28);
buf BUF1 (N95, N91);
buf BUF1 (N96, N85);
buf BUF1 (N97, N93);
xor XOR2 (N98, N66, N49);
and AND4 (N99, N69, N43, N35, N57);
xor XOR2 (N100, N76, N35);
xor XOR2 (N101, N94, N33);
not NOT1 (N102, N97);
buf BUF1 (N103, N89);
nor NOR2 (N104, N98, N50);
nor NOR3 (N105, N102, N64, N80);
not NOT1 (N106, N88);
xor XOR2 (N107, N100, N14);
buf BUF1 (N108, N99);
and AND3 (N109, N87, N82, N71);
not NOT1 (N110, N109);
and AND3 (N111, N103, N31, N79);
buf BUF1 (N112, N95);
not NOT1 (N113, N101);
nor NOR4 (N114, N110, N26, N26, N25);
xor XOR2 (N115, N113, N70);
not NOT1 (N116, N115);
xor XOR2 (N117, N112, N7);
buf BUF1 (N118, N107);
nor NOR2 (N119, N116, N90);
xor XOR2 (N120, N111, N21);
buf BUF1 (N121, N117);
nor NOR3 (N122, N119, N113, N40);
xor XOR2 (N123, N118, N41);
buf BUF1 (N124, N114);
and AND4 (N125, N121, N118, N95, N67);
buf BUF1 (N126, N122);
nor NOR2 (N127, N120, N5);
nor NOR3 (N128, N125, N46, N73);
not NOT1 (N129, N124);
buf BUF1 (N130, N104);
and AND4 (N131, N106, N42, N58, N78);
nor NOR4 (N132, N105, N129, N41, N13);
and AND3 (N133, N16, N106, N60);
buf BUF1 (N134, N96);
not NOT1 (N135, N108);
or OR3 (N136, N132, N118, N31);
nor NOR2 (N137, N128, N42);
not NOT1 (N138, N136);
not NOT1 (N139, N135);
xor XOR2 (N140, N123, N96);
xor XOR2 (N141, N131, N59);
and AND2 (N142, N127, N72);
not NOT1 (N143, N139);
not NOT1 (N144, N137);
buf BUF1 (N145, N126);
xor XOR2 (N146, N144, N19);
or OR2 (N147, N143, N83);
xor XOR2 (N148, N142, N97);
nor NOR4 (N149, N146, N51, N9, N90);
and AND4 (N150, N145, N3, N87, N105);
nand NAND2 (N151, N149, N74);
or OR4 (N152, N130, N67, N115, N142);
and AND3 (N153, N133, N66, N66);
or OR2 (N154, N150, N115);
not NOT1 (N155, N138);
nor NOR3 (N156, N152, N54, N155);
or OR2 (N157, N136, N109);
not NOT1 (N158, N140);
xor XOR2 (N159, N156, N12);
or OR3 (N160, N153, N9, N26);
or OR3 (N161, N134, N90, N127);
or OR4 (N162, N141, N111, N71, N156);
and AND4 (N163, N160, N90, N10, N36);
nand NAND3 (N164, N162, N87, N104);
or OR2 (N165, N147, N156);
not NOT1 (N166, N157);
nand NAND3 (N167, N166, N33, N157);
and AND3 (N168, N158, N48, N22);
buf BUF1 (N169, N167);
buf BUF1 (N170, N168);
buf BUF1 (N171, N154);
and AND3 (N172, N151, N13, N117);
not NOT1 (N173, N159);
nand NAND3 (N174, N172, N61, N134);
or OR4 (N175, N174, N99, N48, N86);
nor NOR4 (N176, N173, N46, N116, N14);
and AND2 (N177, N170, N11);
buf BUF1 (N178, N148);
xor XOR2 (N179, N175, N153);
nand NAND2 (N180, N177, N165);
xor XOR2 (N181, N114, N119);
and AND4 (N182, N179, N142, N158, N93);
or OR4 (N183, N182, N127, N32, N87);
buf BUF1 (N184, N164);
not NOT1 (N185, N183);
buf BUF1 (N186, N178);
or OR2 (N187, N181, N39);
not NOT1 (N188, N180);
and AND3 (N189, N176, N5, N59);
buf BUF1 (N190, N169);
and AND4 (N191, N163, N90, N150, N118);
xor XOR2 (N192, N186, N47);
nand NAND4 (N193, N187, N137, N7, N123);
xor XOR2 (N194, N192, N190);
xor XOR2 (N195, N124, N188);
nand NAND3 (N196, N98, N101, N118);
and AND4 (N197, N193, N193, N136, N17);
nor NOR2 (N198, N195, N196);
nor NOR2 (N199, N125, N185);
xor XOR2 (N200, N71, N165);
or OR4 (N201, N194, N41, N102, N37);
buf BUF1 (N202, N199);
buf BUF1 (N203, N202);
nor NOR2 (N204, N184, N139);
nand NAND2 (N205, N191, N95);
buf BUF1 (N206, N161);
buf BUF1 (N207, N205);
and AND4 (N208, N200, N182, N120, N11);
not NOT1 (N209, N207);
nor NOR3 (N210, N204, N162, N191);
xor XOR2 (N211, N189, N56);
not NOT1 (N212, N206);
xor XOR2 (N213, N208, N174);
nand NAND4 (N214, N197, N67, N32, N68);
buf BUF1 (N215, N209);
buf BUF1 (N216, N198);
or OR3 (N217, N211, N101, N137);
nand NAND2 (N218, N212, N69);
nand NAND2 (N219, N201, N151);
or OR4 (N220, N217, N71, N63, N96);
xor XOR2 (N221, N215, N14);
and AND3 (N222, N203, N4, N98);
xor XOR2 (N223, N216, N98);
nand NAND4 (N224, N218, N176, N30, N68);
or OR2 (N225, N213, N140);
buf BUF1 (N226, N220);
and AND4 (N227, N224, N221, N62, N177);
buf BUF1 (N228, N56);
buf BUF1 (N229, N214);
nand NAND4 (N230, N226, N160, N223, N152);
and AND4 (N231, N230, N209, N229, N109);
or OR3 (N232, N86, N208, N154);
nand NAND3 (N233, N104, N78, N76);
xor XOR2 (N234, N231, N94);
not NOT1 (N235, N227);
or OR3 (N236, N219, N38, N230);
not NOT1 (N237, N222);
not NOT1 (N238, N235);
and AND3 (N239, N238, N226, N186);
or OR2 (N240, N236, N140);
and AND4 (N241, N233, N179, N207, N200);
nor NOR3 (N242, N171, N76, N55);
or OR2 (N243, N240, N182);
buf BUF1 (N244, N234);
or OR4 (N245, N237, N106, N189, N45);
and AND3 (N246, N241, N87, N13);
not NOT1 (N247, N225);
not NOT1 (N248, N239);
xor XOR2 (N249, N243, N205);
not NOT1 (N250, N248);
buf BUF1 (N251, N250);
buf BUF1 (N252, N232);
nor NOR4 (N253, N251, N27, N130, N46);
nor NOR3 (N254, N249, N43, N246);
nand NAND2 (N255, N118, N98);
nor NOR2 (N256, N228, N181);
not NOT1 (N257, N256);
nor NOR3 (N258, N245, N184, N161);
and AND4 (N259, N254, N33, N209, N141);
nand NAND2 (N260, N210, N160);
xor XOR2 (N261, N259, N164);
xor XOR2 (N262, N260, N167);
buf BUF1 (N263, N258);
buf BUF1 (N264, N257);
and AND4 (N265, N242, N151, N175, N215);
nor NOR2 (N266, N265, N72);
or OR3 (N267, N261, N169, N251);
buf BUF1 (N268, N262);
nand NAND3 (N269, N253, N9, N58);
xor XOR2 (N270, N266, N206);
and AND2 (N271, N247, N198);
buf BUF1 (N272, N263);
nor NOR4 (N273, N267, N26, N269, N36);
buf BUF1 (N274, N3);
and AND4 (N275, N268, N201, N174, N99);
and AND2 (N276, N244, N50);
and AND3 (N277, N276, N61, N32);
or OR4 (N278, N271, N46, N185, N219);
not NOT1 (N279, N273);
and AND4 (N280, N264, N196, N12, N162);
buf BUF1 (N281, N280);
not NOT1 (N282, N278);
not NOT1 (N283, N255);
xor XOR2 (N284, N277, N5);
and AND3 (N285, N283, N113, N205);
xor XOR2 (N286, N275, N218);
xor XOR2 (N287, N281, N80);
and AND3 (N288, N272, N249, N162);
xor XOR2 (N289, N288, N187);
buf BUF1 (N290, N285);
nor NOR2 (N291, N270, N180);
nor NOR4 (N292, N289, N44, N48, N243);
xor XOR2 (N293, N290, N165);
or OR4 (N294, N274, N162, N31, N243);
nor NOR4 (N295, N282, N5, N160, N106);
nor NOR3 (N296, N284, N252, N126);
nor NOR2 (N297, N187, N225);
not NOT1 (N298, N286);
xor XOR2 (N299, N295, N123);
buf BUF1 (N300, N299);
nand NAND3 (N301, N298, N227, N179);
buf BUF1 (N302, N291);
buf BUF1 (N303, N292);
not NOT1 (N304, N297);
nand NAND3 (N305, N300, N123, N198);
xor XOR2 (N306, N293, N63);
nand NAND4 (N307, N304, N158, N230, N11);
buf BUF1 (N308, N302);
nor NOR3 (N309, N303, N14, N215);
nand NAND3 (N310, N287, N198, N279);
nand NAND2 (N311, N299, N267);
nand NAND4 (N312, N305, N240, N143, N184);
or OR2 (N313, N307, N40);
xor XOR2 (N314, N301, N313);
and AND2 (N315, N225, N254);
xor XOR2 (N316, N296, N95);
or OR3 (N317, N310, N50, N34);
not NOT1 (N318, N316);
nand NAND3 (N319, N308, N117, N63);
or OR3 (N320, N294, N129, N66);
nor NOR3 (N321, N311, N291, N54);
xor XOR2 (N322, N317, N313);
not NOT1 (N323, N314);
nand NAND2 (N324, N306, N154);
nand NAND3 (N325, N322, N169, N179);
buf BUF1 (N326, N312);
not NOT1 (N327, N325);
nor NOR2 (N328, N326, N189);
nand NAND2 (N329, N328, N71);
buf BUF1 (N330, N309);
nand NAND3 (N331, N319, N51, N122);
xor XOR2 (N332, N331, N121);
or OR2 (N333, N329, N196);
buf BUF1 (N334, N320);
and AND2 (N335, N334, N118);
nand NAND4 (N336, N333, N146, N120, N271);
nand NAND4 (N337, N318, N54, N44, N39);
not NOT1 (N338, N315);
nand NAND4 (N339, N336, N70, N172, N300);
and AND2 (N340, N323, N99);
and AND3 (N341, N340, N272, N57);
xor XOR2 (N342, N338, N198);
nand NAND4 (N343, N341, N93, N307, N325);
xor XOR2 (N344, N343, N309);
buf BUF1 (N345, N337);
xor XOR2 (N346, N342, N28);
buf BUF1 (N347, N330);
not NOT1 (N348, N324);
xor XOR2 (N349, N321, N98);
or OR2 (N350, N335, N22);
nand NAND3 (N351, N347, N296, N256);
or OR4 (N352, N344, N338, N11, N296);
buf BUF1 (N353, N327);
nand NAND3 (N354, N350, N238, N346);
and AND3 (N355, N153, N115, N214);
not NOT1 (N356, N354);
not NOT1 (N357, N339);
or OR2 (N358, N356, N330);
xor XOR2 (N359, N351, N268);
or OR2 (N360, N349, N85);
nor NOR2 (N361, N355, N10);
nand NAND4 (N362, N353, N278, N140, N94);
xor XOR2 (N363, N332, N338);
xor XOR2 (N364, N345, N102);
buf BUF1 (N365, N348);
buf BUF1 (N366, N357);
buf BUF1 (N367, N361);
nor NOR2 (N368, N365, N314);
nand NAND2 (N369, N352, N109);
or OR3 (N370, N366, N255, N311);
buf BUF1 (N371, N364);
or OR2 (N372, N369, N306);
nor NOR3 (N373, N363, N118, N91);
not NOT1 (N374, N358);
xor XOR2 (N375, N372, N234);
nor NOR2 (N376, N374, N290);
buf BUF1 (N377, N360);
nor NOR4 (N378, N373, N366, N309, N318);
buf BUF1 (N379, N375);
not NOT1 (N380, N368);
xor XOR2 (N381, N362, N350);
xor XOR2 (N382, N379, N326);
nor NOR4 (N383, N382, N279, N209, N3);
not NOT1 (N384, N380);
and AND4 (N385, N384, N220, N318, N185);
buf BUF1 (N386, N385);
nor NOR2 (N387, N386, N86);
nor NOR3 (N388, N370, N196, N231);
and AND2 (N389, N378, N243);
or OR4 (N390, N388, N377, N129, N245);
nand NAND2 (N391, N255, N58);
not NOT1 (N392, N371);
nor NOR3 (N393, N381, N57, N371);
nand NAND4 (N394, N383, N267, N47, N192);
and AND4 (N395, N391, N145, N393, N392);
not NOT1 (N396, N141);
not NOT1 (N397, N11);
xor XOR2 (N398, N387, N73);
and AND2 (N399, N376, N118);
xor XOR2 (N400, N399, N224);
and AND4 (N401, N396, N258, N222, N208);
and AND3 (N402, N359, N15, N329);
nand NAND2 (N403, N395, N233);
nor NOR2 (N404, N403, N270);
nand NAND3 (N405, N390, N216, N245);
nor NOR4 (N406, N400, N113, N17, N87);
not NOT1 (N407, N405);
nand NAND4 (N408, N367, N139, N373, N350);
nand NAND4 (N409, N401, N4, N103, N238);
xor XOR2 (N410, N394, N120);
not NOT1 (N411, N406);
xor XOR2 (N412, N398, N164);
not NOT1 (N413, N389);
not NOT1 (N414, N407);
buf BUF1 (N415, N404);
xor XOR2 (N416, N411, N329);
xor XOR2 (N417, N412, N125);
and AND3 (N418, N397, N175, N115);
xor XOR2 (N419, N417, N382);
nor NOR3 (N420, N414, N210, N355);
and AND3 (N421, N413, N109, N82);
buf BUF1 (N422, N419);
xor XOR2 (N423, N422, N285);
buf BUF1 (N424, N418);
nand NAND2 (N425, N424, N387);
and AND2 (N426, N423, N38);
and AND2 (N427, N415, N5);
nor NOR2 (N428, N421, N166);
and AND2 (N429, N410, N81);
nor NOR2 (N430, N427, N66);
not NOT1 (N431, N420);
nor NOR4 (N432, N409, N197, N43, N424);
nor NOR3 (N433, N402, N31, N176);
xor XOR2 (N434, N408, N285);
not NOT1 (N435, N430);
nor NOR4 (N436, N429, N304, N169, N53);
nor NOR3 (N437, N416, N424, N371);
nor NOR4 (N438, N425, N121, N270, N173);
nand NAND4 (N439, N426, N276, N47, N367);
xor XOR2 (N440, N431, N12);
buf BUF1 (N441, N435);
not NOT1 (N442, N433);
or OR3 (N443, N428, N207, N128);
nand NAND2 (N444, N442, N119);
buf BUF1 (N445, N439);
and AND2 (N446, N438, N135);
not NOT1 (N447, N446);
nand NAND3 (N448, N440, N88, N443);
and AND3 (N449, N142, N415, N8);
not NOT1 (N450, N436);
or OR3 (N451, N437, N153, N207);
and AND3 (N452, N445, N303, N274);
nand NAND2 (N453, N432, N375);
nand NAND2 (N454, N452, N407);
not NOT1 (N455, N448);
or OR3 (N456, N449, N238, N47);
xor XOR2 (N457, N453, N368);
not NOT1 (N458, N457);
xor XOR2 (N459, N444, N267);
and AND2 (N460, N455, N4);
or OR4 (N461, N450, N113, N310, N252);
nor NOR3 (N462, N458, N123, N286);
nand NAND2 (N463, N456, N300);
buf BUF1 (N464, N441);
nand NAND4 (N465, N447, N86, N13, N59);
buf BUF1 (N466, N460);
or OR2 (N467, N465, N262);
or OR4 (N468, N462, N120, N136, N165);
xor XOR2 (N469, N464, N378);
not NOT1 (N470, N451);
not NOT1 (N471, N466);
not NOT1 (N472, N434);
and AND2 (N473, N467, N346);
nor NOR4 (N474, N473, N422, N439, N22);
and AND4 (N475, N468, N133, N157, N450);
nor NOR2 (N476, N454, N233);
nor NOR3 (N477, N471, N69, N174);
and AND2 (N478, N474, N87);
buf BUF1 (N479, N469);
not NOT1 (N480, N470);
nor NOR4 (N481, N476, N65, N321, N213);
xor XOR2 (N482, N472, N107);
xor XOR2 (N483, N463, N155);
or OR3 (N484, N461, N421, N443);
buf BUF1 (N485, N484);
nand NAND4 (N486, N477, N89, N288, N117);
nand NAND3 (N487, N485, N186, N85);
and AND2 (N488, N486, N85);
nor NOR4 (N489, N478, N442, N386, N417);
or OR2 (N490, N482, N309);
and AND2 (N491, N488, N449);
and AND3 (N492, N480, N270, N222);
not NOT1 (N493, N459);
not NOT1 (N494, N487);
or OR3 (N495, N483, N491, N158);
xor XOR2 (N496, N465, N213);
or OR3 (N497, N490, N491, N434);
buf BUF1 (N498, N481);
or OR3 (N499, N497, N208, N487);
nor NOR2 (N500, N499, N240);
and AND3 (N501, N496, N461, N389);
not NOT1 (N502, N494);
xor XOR2 (N503, N475, N323);
nor NOR4 (N504, N502, N225, N470, N131);
nor NOR2 (N505, N489, N343);
and AND3 (N506, N501, N243, N186);
nor NOR3 (N507, N479, N108, N335);
nand NAND3 (N508, N498, N269, N21);
nand NAND4 (N509, N506, N184, N235, N12);
buf BUF1 (N510, N493);
and AND3 (N511, N503, N189, N388);
or OR4 (N512, N511, N363, N257, N359);
xor XOR2 (N513, N510, N282);
or OR3 (N514, N513, N455, N116);
or OR3 (N515, N514, N59, N254);
nor NOR4 (N516, N509, N205, N157, N420);
buf BUF1 (N517, N507);
nand NAND2 (N518, N492, N6);
or OR4 (N519, N518, N68, N223, N286);
or OR2 (N520, N508, N109);
nand NAND4 (N521, N520, N144, N83, N361);
not NOT1 (N522, N504);
nand NAND4 (N523, N519, N46, N507, N171);
xor XOR2 (N524, N523, N296);
and AND3 (N525, N500, N209, N447);
and AND2 (N526, N521, N154);
buf BUF1 (N527, N525);
xor XOR2 (N528, N517, N144);
not NOT1 (N529, N512);
nand NAND3 (N530, N515, N457, N377);
xor XOR2 (N531, N528, N75);
nand NAND2 (N532, N505, N515);
buf BUF1 (N533, N529);
nor NOR4 (N534, N524, N159, N371, N394);
not NOT1 (N535, N516);
xor XOR2 (N536, N530, N138);
and AND3 (N537, N522, N334, N342);
nor NOR4 (N538, N532, N452, N348, N180);
and AND3 (N539, N527, N356, N251);
xor XOR2 (N540, N536, N50);
not NOT1 (N541, N526);
nand NAND4 (N542, N538, N212, N501, N340);
nor NOR3 (N543, N542, N379, N326);
buf BUF1 (N544, N533);
nand NAND2 (N545, N531, N407);
buf BUF1 (N546, N534);
buf BUF1 (N547, N543);
nand NAND4 (N548, N544, N437, N11, N252);
xor XOR2 (N549, N548, N536);
xor XOR2 (N550, N547, N328);
xor XOR2 (N551, N550, N458);
nor NOR2 (N552, N541, N406);
and AND2 (N553, N539, N229);
or OR3 (N554, N551, N97, N28);
xor XOR2 (N555, N554, N402);
buf BUF1 (N556, N555);
and AND4 (N557, N540, N262, N329, N540);
xor XOR2 (N558, N537, N458);
and AND4 (N559, N557, N187, N381, N112);
nand NAND2 (N560, N552, N156);
and AND2 (N561, N556, N405);
not NOT1 (N562, N549);
not NOT1 (N563, N545);
xor XOR2 (N564, N546, N523);
and AND4 (N565, N495, N550, N172, N166);
xor XOR2 (N566, N563, N37);
buf BUF1 (N567, N558);
nor NOR2 (N568, N553, N156);
nand NAND3 (N569, N564, N20, N73);
or OR2 (N570, N561, N148);
nor NOR2 (N571, N568, N346);
not NOT1 (N572, N571);
not NOT1 (N573, N569);
xor XOR2 (N574, N559, N336);
nor NOR4 (N575, N560, N350, N185, N510);
and AND4 (N576, N573, N343, N354, N285);
not NOT1 (N577, N565);
xor XOR2 (N578, N576, N352);
nor NOR4 (N579, N567, N522, N468, N267);
nor NOR4 (N580, N566, N14, N238, N527);
and AND3 (N581, N578, N133, N317);
or OR3 (N582, N580, N445, N407);
buf BUF1 (N583, N574);
and AND2 (N584, N577, N6);
xor XOR2 (N585, N575, N139);
xor XOR2 (N586, N579, N325);
not NOT1 (N587, N586);
nand NAND4 (N588, N570, N482, N308, N409);
xor XOR2 (N589, N582, N537);
nor NOR2 (N590, N587, N92);
nor NOR3 (N591, N581, N576, N224);
not NOT1 (N592, N584);
nand NAND4 (N593, N572, N49, N443, N541);
xor XOR2 (N594, N592, N314);
not NOT1 (N595, N594);
not NOT1 (N596, N562);
or OR3 (N597, N589, N181, N23);
nand NAND4 (N598, N583, N111, N204, N61);
nand NAND4 (N599, N591, N350, N494, N156);
or OR2 (N600, N590, N502);
xor XOR2 (N601, N599, N167);
nor NOR3 (N602, N600, N582, N80);
nor NOR2 (N603, N602, N403);
nand NAND2 (N604, N585, N217);
nand NAND3 (N605, N595, N563, N49);
buf BUF1 (N606, N593);
not NOT1 (N607, N535);
or OR2 (N608, N596, N380);
or OR3 (N609, N607, N556, N172);
xor XOR2 (N610, N598, N212);
xor XOR2 (N611, N610, N17);
and AND3 (N612, N604, N556, N202);
and AND4 (N613, N606, N353, N266, N564);
nor NOR2 (N614, N601, N545);
buf BUF1 (N615, N609);
nand NAND3 (N616, N611, N77, N250);
xor XOR2 (N617, N615, N240);
buf BUF1 (N618, N614);
not NOT1 (N619, N618);
buf BUF1 (N620, N588);
or OR3 (N621, N619, N298, N424);
nor NOR2 (N622, N597, N394);
xor XOR2 (N623, N622, N489);
nand NAND2 (N624, N617, N18);
or OR4 (N625, N612, N522, N193, N195);
nor NOR4 (N626, N624, N44, N409, N154);
buf BUF1 (N627, N616);
not NOT1 (N628, N621);
nor NOR3 (N629, N626, N146, N291);
and AND2 (N630, N608, N551);
or OR2 (N631, N630, N164);
nand NAND4 (N632, N613, N434, N396, N255);
and AND2 (N633, N629, N593);
xor XOR2 (N634, N628, N474);
xor XOR2 (N635, N633, N399);
nand NAND4 (N636, N623, N53, N246, N28);
xor XOR2 (N637, N632, N101);
or OR4 (N638, N637, N350, N335, N124);
nand NAND3 (N639, N620, N543, N306);
buf BUF1 (N640, N634);
buf BUF1 (N641, N603);
xor XOR2 (N642, N641, N166);
not NOT1 (N643, N635);
xor XOR2 (N644, N639, N439);
not NOT1 (N645, N636);
not NOT1 (N646, N640);
buf BUF1 (N647, N646);
not NOT1 (N648, N605);
nand NAND4 (N649, N625, N517, N470, N169);
nor NOR2 (N650, N647, N141);
nor NOR4 (N651, N642, N222, N545, N147);
nand NAND2 (N652, N650, N31);
buf BUF1 (N653, N651);
not NOT1 (N654, N648);
and AND2 (N655, N627, N585);
or OR4 (N656, N631, N36, N224, N412);
buf BUF1 (N657, N652);
xor XOR2 (N658, N644, N546);
xor XOR2 (N659, N653, N1);
not NOT1 (N660, N638);
buf BUF1 (N661, N660);
or OR2 (N662, N645, N413);
or OR3 (N663, N658, N217, N523);
or OR4 (N664, N661, N294, N211, N386);
and AND2 (N665, N655, N589);
nor NOR3 (N666, N663, N355, N456);
or OR2 (N667, N665, N1);
nor NOR4 (N668, N657, N552, N512, N348);
nand NAND4 (N669, N656, N282, N7, N571);
and AND3 (N670, N654, N343, N658);
not NOT1 (N671, N670);
or OR4 (N672, N659, N506, N190, N44);
nor NOR3 (N673, N666, N64, N501);
buf BUF1 (N674, N668);
nand NAND2 (N675, N674, N304);
nor NOR3 (N676, N643, N134, N445);
and AND2 (N677, N649, N17);
not NOT1 (N678, N669);
or OR3 (N679, N678, N428, N353);
nor NOR3 (N680, N677, N117, N559);
nand NAND2 (N681, N680, N415);
buf BUF1 (N682, N667);
nor NOR2 (N683, N675, N51);
buf BUF1 (N684, N673);
nor NOR3 (N685, N683, N440, N404);
nor NOR4 (N686, N662, N234, N419, N565);
or OR4 (N687, N671, N563, N160, N393);
xor XOR2 (N688, N679, N102);
buf BUF1 (N689, N688);
xor XOR2 (N690, N689, N469);
and AND3 (N691, N687, N205, N659);
nor NOR3 (N692, N681, N202, N443);
or OR3 (N693, N664, N3, N401);
nand NAND3 (N694, N672, N364, N258);
and AND2 (N695, N691, N476);
nand NAND3 (N696, N685, N79, N522);
nor NOR2 (N697, N692, N542);
and AND4 (N698, N684, N593, N195, N601);
and AND3 (N699, N690, N471, N220);
or OR3 (N700, N696, N569, N430);
and AND2 (N701, N686, N202);
xor XOR2 (N702, N698, N678);
or OR4 (N703, N702, N14, N177, N449);
buf BUF1 (N704, N695);
and AND4 (N705, N697, N260, N32, N451);
or OR4 (N706, N676, N314, N275, N239);
nor NOR4 (N707, N699, N389, N627, N8);
and AND3 (N708, N707, N454, N227);
or OR2 (N709, N704, N206);
nand NAND2 (N710, N705, N493);
buf BUF1 (N711, N700);
nor NOR4 (N712, N709, N629, N485, N404);
buf BUF1 (N713, N682);
nor NOR3 (N714, N703, N230, N222);
not NOT1 (N715, N694);
xor XOR2 (N716, N710, N506);
buf BUF1 (N717, N714);
buf BUF1 (N718, N717);
and AND2 (N719, N708, N201);
or OR3 (N720, N693, N632, N314);
not NOT1 (N721, N713);
buf BUF1 (N722, N715);
nor NOR3 (N723, N718, N635, N597);
buf BUF1 (N724, N711);
nor NOR3 (N725, N723, N555, N601);
xor XOR2 (N726, N722, N706);
or OR3 (N727, N594, N285, N504);
not NOT1 (N728, N724);
xor XOR2 (N729, N720, N216);
or OR2 (N730, N725, N725);
not NOT1 (N731, N730);
nand NAND2 (N732, N729, N580);
xor XOR2 (N733, N721, N427);
and AND2 (N734, N731, N133);
or OR3 (N735, N728, N618, N190);
nand NAND3 (N736, N716, N98, N701);
and AND4 (N737, N736, N712, N6, N121);
nand NAND4 (N738, N137, N522, N21, N569);
xor XOR2 (N739, N277, N464);
not NOT1 (N740, N737);
and AND3 (N741, N734, N299, N55);
buf BUF1 (N742, N732);
not NOT1 (N743, N735);
buf BUF1 (N744, N727);
nor NOR4 (N745, N741, N387, N422, N115);
and AND3 (N746, N744, N526, N502);
nand NAND2 (N747, N738, N96);
nand NAND2 (N748, N747, N145);
or OR3 (N749, N745, N51, N735);
and AND3 (N750, N719, N91, N326);
and AND4 (N751, N739, N713, N27, N296);
not NOT1 (N752, N746);
buf BUF1 (N753, N749);
or OR4 (N754, N743, N675, N225, N136);
nand NAND4 (N755, N754, N319, N89, N57);
not NOT1 (N756, N726);
or OR2 (N757, N742, N741);
buf BUF1 (N758, N751);
or OR2 (N759, N748, N56);
nand NAND4 (N760, N753, N440, N266, N300);
nand NAND3 (N761, N740, N543, N227);
nand NAND2 (N762, N757, N464);
or OR3 (N763, N755, N486, N616);
nand NAND4 (N764, N762, N190, N111, N347);
not NOT1 (N765, N756);
xor XOR2 (N766, N750, N288);
nand NAND2 (N767, N758, N196);
nor NOR2 (N768, N765, N2);
xor XOR2 (N769, N763, N165);
buf BUF1 (N770, N767);
nand NAND2 (N771, N770, N118);
nand NAND4 (N772, N766, N290, N707, N512);
nand NAND3 (N773, N768, N677, N653);
xor XOR2 (N774, N759, N629);
nor NOR3 (N775, N760, N668, N699);
not NOT1 (N776, N752);
and AND2 (N777, N776, N318);
buf BUF1 (N778, N773);
xor XOR2 (N779, N775, N427);
nor NOR3 (N780, N733, N280, N697);
and AND3 (N781, N778, N42, N227);
nor NOR3 (N782, N764, N636, N375);
xor XOR2 (N783, N774, N273);
xor XOR2 (N784, N769, N21);
not NOT1 (N785, N784);
buf BUF1 (N786, N781);
and AND4 (N787, N786, N169, N228, N307);
and AND4 (N788, N785, N638, N669, N444);
or OR4 (N789, N779, N732, N530, N523);
or OR4 (N790, N783, N280, N637, N411);
and AND2 (N791, N782, N735);
and AND2 (N792, N777, N47);
not NOT1 (N793, N792);
and AND2 (N794, N771, N139);
and AND3 (N795, N761, N66, N601);
not NOT1 (N796, N789);
or OR2 (N797, N790, N229);
buf BUF1 (N798, N791);
buf BUF1 (N799, N772);
not NOT1 (N800, N798);
not NOT1 (N801, N799);
nand NAND3 (N802, N800, N108, N159);
and AND4 (N803, N802, N742, N589, N668);
nor NOR4 (N804, N788, N37, N37, N218);
and AND3 (N805, N803, N362, N613);
or OR3 (N806, N796, N80, N172);
xor XOR2 (N807, N797, N146);
not NOT1 (N808, N794);
nor NOR3 (N809, N808, N303, N116);
nand NAND2 (N810, N801, N518);
or OR4 (N811, N804, N142, N218, N79);
buf BUF1 (N812, N806);
buf BUF1 (N813, N810);
buf BUF1 (N814, N780);
nand NAND2 (N815, N814, N705);
buf BUF1 (N816, N793);
buf BUF1 (N817, N787);
nand NAND3 (N818, N811, N698, N86);
not NOT1 (N819, N818);
xor XOR2 (N820, N807, N763);
not NOT1 (N821, N815);
nor NOR3 (N822, N821, N555, N305);
or OR3 (N823, N820, N466, N456);
or OR4 (N824, N819, N495, N190, N182);
not NOT1 (N825, N816);
nand NAND4 (N826, N805, N368, N173, N38);
and AND3 (N827, N809, N333, N85);
and AND4 (N828, N813, N620, N546, N706);
nand NAND4 (N829, N823, N166, N324, N44);
not NOT1 (N830, N824);
buf BUF1 (N831, N828);
not NOT1 (N832, N829);
xor XOR2 (N833, N812, N616);
or OR2 (N834, N825, N762);
nand NAND3 (N835, N832, N685, N528);
buf BUF1 (N836, N817);
nand NAND4 (N837, N795, N604, N339, N86);
nor NOR4 (N838, N835, N179, N336, N477);
nand NAND3 (N839, N830, N79, N12);
nand NAND3 (N840, N837, N117, N724);
nand NAND3 (N841, N822, N320, N800);
nand NAND3 (N842, N833, N494, N489);
nor NOR3 (N843, N836, N698, N145);
and AND2 (N844, N831, N378);
not NOT1 (N845, N838);
not NOT1 (N846, N834);
nor NOR4 (N847, N840, N816, N389, N248);
buf BUF1 (N848, N847);
or OR4 (N849, N844, N65, N760, N74);
buf BUF1 (N850, N826);
xor XOR2 (N851, N842, N67);
buf BUF1 (N852, N850);
not NOT1 (N853, N845);
xor XOR2 (N854, N851, N163);
xor XOR2 (N855, N843, N58);
buf BUF1 (N856, N848);
buf BUF1 (N857, N855);
nand NAND3 (N858, N854, N51, N628);
and AND2 (N859, N853, N384);
nand NAND2 (N860, N858, N795);
xor XOR2 (N861, N857, N724);
nand NAND4 (N862, N839, N168, N733, N49);
or OR2 (N863, N862, N85);
nand NAND4 (N864, N859, N845, N340, N522);
buf BUF1 (N865, N863);
xor XOR2 (N866, N856, N279);
buf BUF1 (N867, N864);
nor NOR4 (N868, N861, N33, N505, N252);
not NOT1 (N869, N852);
buf BUF1 (N870, N841);
xor XOR2 (N871, N860, N417);
xor XOR2 (N872, N865, N445);
not NOT1 (N873, N868);
or OR4 (N874, N869, N230, N432, N753);
not NOT1 (N875, N866);
nand NAND2 (N876, N846, N650);
or OR2 (N877, N872, N102);
or OR4 (N878, N874, N786, N297, N638);
nand NAND3 (N879, N876, N207, N404);
nor NOR2 (N880, N877, N30);
nor NOR2 (N881, N870, N247);
not NOT1 (N882, N827);
nor NOR2 (N883, N867, N717);
nand NAND3 (N884, N881, N157, N399);
nor NOR2 (N885, N883, N847);
buf BUF1 (N886, N879);
nand NAND2 (N887, N871, N531);
not NOT1 (N888, N880);
and AND3 (N889, N888, N385, N693);
not NOT1 (N890, N885);
or OR4 (N891, N886, N413, N549, N416);
and AND3 (N892, N889, N465, N682);
and AND4 (N893, N892, N137, N243, N176);
and AND2 (N894, N882, N845);
nor NOR4 (N895, N873, N522, N769, N628);
xor XOR2 (N896, N884, N578);
buf BUF1 (N897, N887);
xor XOR2 (N898, N893, N225);
nor NOR2 (N899, N890, N651);
not NOT1 (N900, N891);
xor XOR2 (N901, N875, N5);
or OR4 (N902, N896, N586, N265, N549);
nand NAND2 (N903, N895, N127);
buf BUF1 (N904, N903);
nand NAND3 (N905, N878, N767, N139);
or OR2 (N906, N902, N101);
buf BUF1 (N907, N904);
not NOT1 (N908, N894);
buf BUF1 (N909, N897);
or OR2 (N910, N909, N292);
not NOT1 (N911, N907);
xor XOR2 (N912, N898, N811);
or OR2 (N913, N910, N799);
nor NOR4 (N914, N911, N111, N332, N477);
or OR3 (N915, N899, N130, N909);
not NOT1 (N916, N915);
xor XOR2 (N917, N912, N249);
buf BUF1 (N918, N908);
buf BUF1 (N919, N916);
or OR3 (N920, N849, N915, N912);
buf BUF1 (N921, N900);
and AND3 (N922, N918, N55, N631);
nand NAND2 (N923, N914, N527);
not NOT1 (N924, N919);
or OR3 (N925, N924, N614, N534);
or OR2 (N926, N906, N132);
and AND4 (N927, N905, N175, N381, N639);
or OR4 (N928, N926, N594, N306, N854);
nand NAND4 (N929, N920, N585, N798, N291);
nand NAND3 (N930, N929, N331, N426);
or OR4 (N931, N901, N748, N326, N525);
xor XOR2 (N932, N923, N350);
buf BUF1 (N933, N925);
xor XOR2 (N934, N933, N815);
and AND3 (N935, N930, N119, N703);
and AND4 (N936, N931, N84, N290, N691);
xor XOR2 (N937, N936, N811);
nand NAND2 (N938, N935, N873);
xor XOR2 (N939, N917, N726);
nor NOR4 (N940, N921, N515, N482, N124);
nor NOR3 (N941, N934, N907, N652);
buf BUF1 (N942, N932);
and AND4 (N943, N928, N195, N715, N767);
nor NOR4 (N944, N940, N333, N570, N805);
nand NAND3 (N945, N943, N102, N560);
not NOT1 (N946, N941);
not NOT1 (N947, N944);
and AND4 (N948, N947, N502, N48, N836);
not NOT1 (N949, N913);
or OR2 (N950, N946, N872);
not NOT1 (N951, N939);
buf BUF1 (N952, N937);
nand NAND4 (N953, N948, N720, N382, N49);
xor XOR2 (N954, N951, N410);
not NOT1 (N955, N949);
or OR3 (N956, N927, N229, N866);
nand NAND2 (N957, N953, N783);
buf BUF1 (N958, N956);
nor NOR2 (N959, N955, N357);
nor NOR3 (N960, N950, N120, N828);
not NOT1 (N961, N942);
buf BUF1 (N962, N958);
or OR3 (N963, N945, N581, N693);
nand NAND2 (N964, N938, N183);
or OR4 (N965, N964, N350, N270, N837);
buf BUF1 (N966, N954);
xor XOR2 (N967, N922, N369);
nand NAND3 (N968, N963, N582, N484);
xor XOR2 (N969, N962, N275);
not NOT1 (N970, N960);
nand NAND4 (N971, N965, N340, N729, N963);
not NOT1 (N972, N970);
nand NAND2 (N973, N967, N793);
or OR2 (N974, N971, N483);
and AND2 (N975, N959, N56);
xor XOR2 (N976, N975, N498);
xor XOR2 (N977, N976, N80);
nor NOR3 (N978, N969, N547, N59);
xor XOR2 (N979, N973, N725);
or OR4 (N980, N961, N698, N533, N336);
not NOT1 (N981, N978);
xor XOR2 (N982, N974, N503);
or OR3 (N983, N981, N282, N111);
nand NAND3 (N984, N957, N686, N749);
nand NAND3 (N985, N952, N154, N766);
nor NOR4 (N986, N980, N338, N444, N14);
and AND2 (N987, N968, N725);
or OR2 (N988, N984, N369);
or OR3 (N989, N977, N599, N432);
buf BUF1 (N990, N985);
buf BUF1 (N991, N966);
buf BUF1 (N992, N983);
and AND4 (N993, N992, N922, N857, N347);
xor XOR2 (N994, N979, N86);
nor NOR4 (N995, N986, N762, N758, N71);
not NOT1 (N996, N987);
xor XOR2 (N997, N993, N642);
xor XOR2 (N998, N991, N14);
xor XOR2 (N999, N988, N755);
or OR4 (N1000, N990, N257, N816, N311);
not NOT1 (N1001, N972);
nor NOR4 (N1002, N989, N354, N36, N862);
or OR4 (N1003, N998, N643, N377, N974);
buf BUF1 (N1004, N1003);
or OR3 (N1005, N1002, N832, N666);
or OR3 (N1006, N994, N389, N327);
xor XOR2 (N1007, N1006, N941);
not NOT1 (N1008, N997);
or OR2 (N1009, N996, N593);
buf BUF1 (N1010, N1004);
buf BUF1 (N1011, N995);
xor XOR2 (N1012, N1010, N391);
buf BUF1 (N1013, N1012);
buf BUF1 (N1014, N1011);
nand NAND3 (N1015, N1014, N795, N43);
xor XOR2 (N1016, N999, N928);
nand NAND2 (N1017, N1005, N724);
not NOT1 (N1018, N1017);
nand NAND4 (N1019, N1015, N871, N809, N413);
and AND2 (N1020, N1001, N234);
not NOT1 (N1021, N1020);
not NOT1 (N1022, N1019);
and AND3 (N1023, N1021, N773, N875);
not NOT1 (N1024, N1013);
nor NOR3 (N1025, N1000, N541, N599);
nor NOR2 (N1026, N1023, N770);
or OR3 (N1027, N1026, N173, N964);
xor XOR2 (N1028, N1027, N702);
or OR3 (N1029, N1007, N620, N951);
nor NOR3 (N1030, N1008, N255, N380);
nand NAND4 (N1031, N1024, N860, N679, N772);
buf BUF1 (N1032, N1031);
nand NAND3 (N1033, N1009, N511, N391);
or OR3 (N1034, N1033, N241, N787);
buf BUF1 (N1035, N1022);
nand NAND2 (N1036, N1016, N767);
not NOT1 (N1037, N1029);
and AND3 (N1038, N1034, N277, N228);
not NOT1 (N1039, N1032);
nand NAND4 (N1040, N1028, N723, N961, N284);
or OR4 (N1041, N1030, N2, N103, N64);
buf BUF1 (N1042, N1039);
and AND3 (N1043, N1035, N399, N503);
and AND3 (N1044, N1037, N340, N112);
xor XOR2 (N1045, N1040, N256);
not NOT1 (N1046, N1038);
nand NAND4 (N1047, N1043, N641, N303, N601);
nand NAND3 (N1048, N1045, N912, N756);
xor XOR2 (N1049, N1047, N326);
not NOT1 (N1050, N982);
buf BUF1 (N1051, N1044);
nand NAND3 (N1052, N1050, N195, N522);
nand NAND2 (N1053, N1041, N724);
and AND3 (N1054, N1048, N848, N28);
not NOT1 (N1055, N1054);
nand NAND3 (N1056, N1051, N457, N265);
xor XOR2 (N1057, N1025, N298);
or OR4 (N1058, N1055, N189, N557, N284);
xor XOR2 (N1059, N1042, N196);
and AND3 (N1060, N1056, N12, N763);
buf BUF1 (N1061, N1053);
and AND4 (N1062, N1046, N7, N136, N393);
xor XOR2 (N1063, N1049, N992);
nor NOR4 (N1064, N1057, N545, N294, N575);
nand NAND2 (N1065, N1062, N271);
not NOT1 (N1066, N1052);
or OR3 (N1067, N1064, N409, N683);
buf BUF1 (N1068, N1067);
nor NOR2 (N1069, N1036, N318);
nor NOR3 (N1070, N1059, N313, N9);
not NOT1 (N1071, N1058);
xor XOR2 (N1072, N1066, N757);
nand NAND2 (N1073, N1061, N157);
buf BUF1 (N1074, N1068);
buf BUF1 (N1075, N1073);
or OR4 (N1076, N1069, N462, N805, N660);
buf BUF1 (N1077, N1072);
nor NOR2 (N1078, N1070, N314);
or OR4 (N1079, N1077, N564, N796, N771);
buf BUF1 (N1080, N1078);
xor XOR2 (N1081, N1065, N884);
xor XOR2 (N1082, N1079, N850);
or OR3 (N1083, N1081, N580, N997);
not NOT1 (N1084, N1082);
not NOT1 (N1085, N1071);
buf BUF1 (N1086, N1060);
nor NOR2 (N1087, N1063, N272);
xor XOR2 (N1088, N1074, N361);
not NOT1 (N1089, N1085);
and AND4 (N1090, N1075, N891, N333, N1036);
nor NOR4 (N1091, N1090, N474, N1080, N617);
not NOT1 (N1092, N790);
nand NAND4 (N1093, N1089, N747, N362, N29);
and AND2 (N1094, N1091, N157);
nor NOR3 (N1095, N1018, N717, N386);
or OR2 (N1096, N1087, N27);
and AND2 (N1097, N1088, N200);
and AND4 (N1098, N1096, N1016, N1086, N758);
and AND4 (N1099, N743, N487, N992, N384);
or OR4 (N1100, N1094, N58, N756, N352);
xor XOR2 (N1101, N1076, N1081);
nand NAND2 (N1102, N1100, N975);
buf BUF1 (N1103, N1101);
and AND3 (N1104, N1099, N516, N68);
xor XOR2 (N1105, N1093, N270);
buf BUF1 (N1106, N1102);
nand NAND2 (N1107, N1097, N784);
buf BUF1 (N1108, N1092);
xor XOR2 (N1109, N1083, N610);
nor NOR4 (N1110, N1108, N796, N330, N758);
buf BUF1 (N1111, N1110);
and AND2 (N1112, N1106, N983);
buf BUF1 (N1113, N1098);
xor XOR2 (N1114, N1084, N230);
and AND4 (N1115, N1111, N1043, N986, N1059);
and AND4 (N1116, N1107, N267, N970, N696);
nor NOR3 (N1117, N1116, N114, N232);
nor NOR3 (N1118, N1105, N826, N366);
not NOT1 (N1119, N1118);
and AND3 (N1120, N1103, N479, N454);
nor NOR2 (N1121, N1095, N149);
and AND4 (N1122, N1114, N469, N41, N930);
not NOT1 (N1123, N1121);
nor NOR2 (N1124, N1122, N601);
buf BUF1 (N1125, N1119);
nor NOR4 (N1126, N1120, N701, N939, N661);
not NOT1 (N1127, N1125);
not NOT1 (N1128, N1104);
and AND3 (N1129, N1127, N674, N639);
not NOT1 (N1130, N1117);
nor NOR2 (N1131, N1112, N643);
nor NOR2 (N1132, N1115, N335);
or OR2 (N1133, N1132, N935);
and AND4 (N1134, N1109, N1123, N273, N457);
xor XOR2 (N1135, N797, N300);
or OR2 (N1136, N1113, N1126);
or OR3 (N1137, N1060, N388, N369);
or OR4 (N1138, N1124, N103, N119, N417);
buf BUF1 (N1139, N1128);
nand NAND3 (N1140, N1136, N375, N34);
and AND4 (N1141, N1129, N78, N21, N340);
nor NOR4 (N1142, N1140, N593, N1120, N415);
and AND2 (N1143, N1133, N925);
or OR2 (N1144, N1141, N878);
xor XOR2 (N1145, N1130, N123);
buf BUF1 (N1146, N1131);
nor NOR2 (N1147, N1143, N93);
buf BUF1 (N1148, N1135);
nor NOR4 (N1149, N1144, N1037, N1009, N668);
nand NAND4 (N1150, N1139, N501, N788, N1001);
or OR2 (N1151, N1149, N808);
or OR3 (N1152, N1142, N1104, N745);
buf BUF1 (N1153, N1138);
xor XOR2 (N1154, N1147, N422);
or OR2 (N1155, N1145, N189);
not NOT1 (N1156, N1146);
not NOT1 (N1157, N1152);
nor NOR4 (N1158, N1157, N1106, N848, N135);
buf BUF1 (N1159, N1153);
nor NOR2 (N1160, N1134, N344);
buf BUF1 (N1161, N1155);
nor NOR4 (N1162, N1161, N734, N55, N591);
or OR3 (N1163, N1150, N659, N21);
not NOT1 (N1164, N1151);
not NOT1 (N1165, N1148);
nand NAND4 (N1166, N1162, N1023, N1, N337);
nor NOR4 (N1167, N1137, N1153, N592, N425);
xor XOR2 (N1168, N1164, N105);
or OR3 (N1169, N1156, N1043, N121);
nand NAND4 (N1170, N1158, N1125, N87, N1004);
nand NAND2 (N1171, N1170, N991);
not NOT1 (N1172, N1171);
xor XOR2 (N1173, N1159, N39);
not NOT1 (N1174, N1168);
or OR2 (N1175, N1166, N406);
and AND2 (N1176, N1163, N541);
and AND4 (N1177, N1160, N88, N398, N212);
and AND4 (N1178, N1172, N813, N762, N606);
not NOT1 (N1179, N1176);
xor XOR2 (N1180, N1177, N1093);
buf BUF1 (N1181, N1179);
not NOT1 (N1182, N1173);
nand NAND3 (N1183, N1174, N816, N556);
nand NAND3 (N1184, N1154, N1147, N98);
buf BUF1 (N1185, N1184);
xor XOR2 (N1186, N1167, N495);
not NOT1 (N1187, N1180);
or OR4 (N1188, N1181, N87, N270, N862);
nand NAND3 (N1189, N1165, N1141, N733);
or OR3 (N1190, N1189, N310, N948);
xor XOR2 (N1191, N1175, N104);
not NOT1 (N1192, N1191);
and AND4 (N1193, N1186, N559, N640, N981);
buf BUF1 (N1194, N1190);
nand NAND3 (N1195, N1185, N260, N189);
not NOT1 (N1196, N1193);
and AND2 (N1197, N1178, N249);
or OR4 (N1198, N1182, N966, N943, N402);
nor NOR4 (N1199, N1197, N622, N363, N697);
and AND4 (N1200, N1188, N131, N396, N867);
nand NAND2 (N1201, N1194, N1186);
or OR2 (N1202, N1200, N941);
not NOT1 (N1203, N1183);
nand NAND3 (N1204, N1201, N39, N258);
nand NAND2 (N1205, N1202, N29);
and AND2 (N1206, N1196, N56);
not NOT1 (N1207, N1203);
buf BUF1 (N1208, N1198);
buf BUF1 (N1209, N1207);
not NOT1 (N1210, N1208);
and AND4 (N1211, N1204, N675, N942, N955);
and AND2 (N1212, N1206, N1143);
buf BUF1 (N1213, N1211);
and AND2 (N1214, N1210, N883);
or OR4 (N1215, N1214, N571, N910, N540);
nor NOR2 (N1216, N1169, N1179);
or OR4 (N1217, N1213, N213, N508, N378);
not NOT1 (N1218, N1199);
xor XOR2 (N1219, N1218, N539);
nand NAND4 (N1220, N1212, N470, N941, N1047);
nor NOR4 (N1221, N1217, N208, N872, N849);
not NOT1 (N1222, N1215);
nor NOR2 (N1223, N1222, N130);
nand NAND3 (N1224, N1220, N639, N36);
xor XOR2 (N1225, N1195, N875);
buf BUF1 (N1226, N1209);
or OR4 (N1227, N1226, N468, N509, N156);
xor XOR2 (N1228, N1187, N1160);
nand NAND3 (N1229, N1219, N102, N825);
nand NAND4 (N1230, N1225, N366, N514, N714);
buf BUF1 (N1231, N1227);
or OR4 (N1232, N1224, N1176, N750, N809);
nand NAND2 (N1233, N1221, N1128);
xor XOR2 (N1234, N1192, N815);
nor NOR4 (N1235, N1228, N536, N152, N1069);
nand NAND4 (N1236, N1230, N561, N1024, N135);
or OR2 (N1237, N1229, N342);
nand NAND4 (N1238, N1232, N878, N27, N578);
not NOT1 (N1239, N1236);
and AND4 (N1240, N1223, N850, N529, N250);
not NOT1 (N1241, N1216);
xor XOR2 (N1242, N1241, N349);
not NOT1 (N1243, N1205);
not NOT1 (N1244, N1240);
xor XOR2 (N1245, N1239, N313);
xor XOR2 (N1246, N1235, N669);
or OR2 (N1247, N1238, N189);
nor NOR2 (N1248, N1237, N1035);
nand NAND2 (N1249, N1245, N777);
or OR3 (N1250, N1231, N1239, N184);
and AND4 (N1251, N1249, N805, N888, N56);
nand NAND2 (N1252, N1234, N1011);
and AND3 (N1253, N1242, N939, N920);
nor NOR2 (N1254, N1248, N32);
nand NAND3 (N1255, N1247, N37, N868);
nand NAND4 (N1256, N1253, N239, N726, N767);
nor NOR4 (N1257, N1233, N139, N896, N601);
and AND3 (N1258, N1254, N1083, N920);
nor NOR3 (N1259, N1256, N466, N505);
and AND3 (N1260, N1257, N93, N807);
xor XOR2 (N1261, N1244, N63);
not NOT1 (N1262, N1246);
nor NOR2 (N1263, N1259, N1066);
nand NAND2 (N1264, N1260, N910);
not NOT1 (N1265, N1252);
nor NOR2 (N1266, N1255, N185);
xor XOR2 (N1267, N1251, N228);
nand NAND4 (N1268, N1262, N1241, N1214, N1231);
nand NAND3 (N1269, N1265, N316, N231);
or OR3 (N1270, N1261, N268, N1043);
buf BUF1 (N1271, N1266);
or OR4 (N1272, N1271, N1197, N826, N1073);
and AND3 (N1273, N1263, N373, N784);
not NOT1 (N1274, N1264);
and AND3 (N1275, N1258, N623, N496);
and AND2 (N1276, N1269, N558);
or OR2 (N1277, N1272, N970);
and AND3 (N1278, N1250, N550, N1037);
and AND2 (N1279, N1270, N1069);
nand NAND4 (N1280, N1276, N417, N402, N521);
and AND3 (N1281, N1275, N812, N1166);
xor XOR2 (N1282, N1243, N1059);
nor NOR2 (N1283, N1281, N180);
not NOT1 (N1284, N1274);
buf BUF1 (N1285, N1282);
and AND4 (N1286, N1277, N320, N1122, N434);
nor NOR2 (N1287, N1278, N942);
or OR4 (N1288, N1268, N1153, N903, N226);
or OR2 (N1289, N1288, N214);
not NOT1 (N1290, N1289);
or OR2 (N1291, N1284, N1073);
nand NAND2 (N1292, N1273, N540);
or OR3 (N1293, N1267, N1244, N413);
xor XOR2 (N1294, N1290, N722);
not NOT1 (N1295, N1291);
nand NAND2 (N1296, N1285, N579);
or OR2 (N1297, N1286, N876);
buf BUF1 (N1298, N1296);
nor NOR4 (N1299, N1295, N924, N433, N469);
or OR4 (N1300, N1298, N727, N172, N252);
buf BUF1 (N1301, N1294);
nor NOR3 (N1302, N1287, N967, N917);
nor NOR2 (N1303, N1300, N141);
and AND2 (N1304, N1280, N123);
buf BUF1 (N1305, N1283);
xor XOR2 (N1306, N1302, N1087);
and AND4 (N1307, N1306, N558, N557, N30);
buf BUF1 (N1308, N1297);
nand NAND3 (N1309, N1307, N113, N992);
and AND3 (N1310, N1279, N402, N1217);
buf BUF1 (N1311, N1308);
not NOT1 (N1312, N1293);
and AND4 (N1313, N1305, N613, N307, N886);
nor NOR4 (N1314, N1310, N738, N39, N936);
not NOT1 (N1315, N1312);
or OR2 (N1316, N1303, N775);
xor XOR2 (N1317, N1309, N475);
buf BUF1 (N1318, N1304);
xor XOR2 (N1319, N1318, N1173);
or OR2 (N1320, N1313, N419);
or OR2 (N1321, N1314, N487);
xor XOR2 (N1322, N1315, N579);
not NOT1 (N1323, N1292);
or OR3 (N1324, N1322, N1259, N867);
and AND4 (N1325, N1320, N258, N1274, N50);
or OR4 (N1326, N1316, N1009, N1183, N772);
nor NOR3 (N1327, N1324, N1014, N528);
buf BUF1 (N1328, N1323);
not NOT1 (N1329, N1325);
nor NOR3 (N1330, N1326, N1176, N678);
and AND4 (N1331, N1327, N673, N483, N26);
nand NAND4 (N1332, N1328, N195, N377, N478);
not NOT1 (N1333, N1332);
or OR2 (N1334, N1331, N708);
not NOT1 (N1335, N1317);
buf BUF1 (N1336, N1334);
or OR2 (N1337, N1319, N1109);
nand NAND3 (N1338, N1321, N830, N183);
xor XOR2 (N1339, N1330, N600);
nand NAND4 (N1340, N1311, N485, N1041, N1137);
buf BUF1 (N1341, N1338);
buf BUF1 (N1342, N1341);
xor XOR2 (N1343, N1339, N792);
or OR3 (N1344, N1301, N962, N1159);
nor NOR2 (N1345, N1343, N215);
xor XOR2 (N1346, N1333, N90);
or OR4 (N1347, N1299, N359, N586, N189);
nor NOR3 (N1348, N1337, N1194, N1064);
nor NOR4 (N1349, N1340, N675, N963, N120);
nor NOR3 (N1350, N1347, N745, N1246);
nand NAND4 (N1351, N1342, N1284, N81, N75);
nand NAND4 (N1352, N1348, N783, N227, N1318);
and AND2 (N1353, N1349, N942);
not NOT1 (N1354, N1353);
or OR2 (N1355, N1335, N283);
or OR3 (N1356, N1355, N90, N606);
not NOT1 (N1357, N1345);
nor NOR3 (N1358, N1357, N812, N43);
buf BUF1 (N1359, N1352);
nand NAND4 (N1360, N1346, N706, N1081, N801);
and AND4 (N1361, N1329, N520, N1287, N748);
or OR3 (N1362, N1354, N1209, N1027);
not NOT1 (N1363, N1358);
and AND2 (N1364, N1359, N1018);
xor XOR2 (N1365, N1344, N259);
nor NOR4 (N1366, N1356, N679, N691, N538);
not NOT1 (N1367, N1363);
not NOT1 (N1368, N1350);
not NOT1 (N1369, N1351);
not NOT1 (N1370, N1336);
xor XOR2 (N1371, N1364, N408);
xor XOR2 (N1372, N1365, N566);
and AND3 (N1373, N1368, N416, N801);
nand NAND2 (N1374, N1366, N1092);
xor XOR2 (N1375, N1372, N51);
nor NOR2 (N1376, N1369, N410);
nand NAND2 (N1377, N1371, N391);
or OR2 (N1378, N1375, N686);
xor XOR2 (N1379, N1360, N1352);
not NOT1 (N1380, N1361);
nand NAND4 (N1381, N1374, N303, N1133, N1232);
not NOT1 (N1382, N1381);
xor XOR2 (N1383, N1362, N1211);
xor XOR2 (N1384, N1378, N1150);
nor NOR3 (N1385, N1373, N1345, N833);
nand NAND2 (N1386, N1376, N1342);
or OR2 (N1387, N1367, N116);
not NOT1 (N1388, N1386);
buf BUF1 (N1389, N1384);
xor XOR2 (N1390, N1370, N729);
buf BUF1 (N1391, N1388);
or OR3 (N1392, N1385, N717, N411);
nor NOR3 (N1393, N1387, N23, N744);
buf BUF1 (N1394, N1383);
buf BUF1 (N1395, N1382);
nor NOR2 (N1396, N1391, N801);
nor NOR4 (N1397, N1377, N750, N1289, N537);
xor XOR2 (N1398, N1393, N708);
nor NOR4 (N1399, N1394, N211, N1337, N1336);
nor NOR4 (N1400, N1390, N306, N682, N232);
buf BUF1 (N1401, N1397);
not NOT1 (N1402, N1400);
not NOT1 (N1403, N1379);
nor NOR3 (N1404, N1399, N405, N658);
or OR4 (N1405, N1392, N889, N1334, N689);
and AND2 (N1406, N1380, N223);
nand NAND3 (N1407, N1406, N835, N1124);
nand NAND2 (N1408, N1395, N534);
and AND2 (N1409, N1396, N1094);
nor NOR2 (N1410, N1402, N220);
and AND3 (N1411, N1398, N462, N1187);
nor NOR4 (N1412, N1403, N1226, N1108, N1296);
not NOT1 (N1413, N1407);
or OR4 (N1414, N1411, N468, N338, N702);
or OR3 (N1415, N1404, N921, N971);
and AND3 (N1416, N1414, N278, N550);
nand NAND3 (N1417, N1389, N858, N805);
xor XOR2 (N1418, N1415, N36);
not NOT1 (N1419, N1418);
xor XOR2 (N1420, N1413, N906);
and AND4 (N1421, N1412, N354, N1007, N547);
and AND2 (N1422, N1410, N1286);
not NOT1 (N1423, N1419);
and AND3 (N1424, N1417, N1340, N144);
nor NOR2 (N1425, N1401, N171);
or OR3 (N1426, N1424, N200, N1095);
xor XOR2 (N1427, N1421, N1068);
xor XOR2 (N1428, N1409, N560);
buf BUF1 (N1429, N1416);
not NOT1 (N1430, N1423);
not NOT1 (N1431, N1427);
xor XOR2 (N1432, N1426, N1421);
and AND4 (N1433, N1432, N921, N778, N1270);
not NOT1 (N1434, N1433);
not NOT1 (N1435, N1405);
not NOT1 (N1436, N1429);
and AND2 (N1437, N1422, N614);
and AND4 (N1438, N1420, N577, N1127, N867);
or OR2 (N1439, N1431, N445);
nand NAND4 (N1440, N1435, N398, N554, N720);
xor XOR2 (N1441, N1430, N749);
nor NOR2 (N1442, N1425, N924);
buf BUF1 (N1443, N1437);
and AND3 (N1444, N1439, N283, N1072);
not NOT1 (N1445, N1438);
xor XOR2 (N1446, N1440, N860);
nor NOR2 (N1447, N1441, N707);
nor NOR4 (N1448, N1444, N83, N127, N1045);
or OR3 (N1449, N1445, N133, N682);
xor XOR2 (N1450, N1447, N273);
xor XOR2 (N1451, N1448, N206);
buf BUF1 (N1452, N1442);
nand NAND4 (N1453, N1452, N989, N859, N1148);
buf BUF1 (N1454, N1428);
nor NOR4 (N1455, N1449, N54, N94, N444);
not NOT1 (N1456, N1454);
xor XOR2 (N1457, N1451, N1244);
buf BUF1 (N1458, N1455);
not NOT1 (N1459, N1408);
xor XOR2 (N1460, N1443, N1138);
nor NOR2 (N1461, N1459, N54);
or OR4 (N1462, N1450, N338, N955, N420);
nand NAND4 (N1463, N1458, N920, N489, N1107);
nor NOR3 (N1464, N1461, N989, N623);
and AND3 (N1465, N1434, N1105, N838);
xor XOR2 (N1466, N1464, N905);
nand NAND2 (N1467, N1436, N1383);
nand NAND2 (N1468, N1446, N436);
nor NOR3 (N1469, N1462, N1253, N1265);
nand NAND3 (N1470, N1463, N865, N1376);
and AND4 (N1471, N1460, N1132, N733, N35);
xor XOR2 (N1472, N1465, N1256);
not NOT1 (N1473, N1469);
nand NAND2 (N1474, N1470, N244);
or OR4 (N1475, N1474, N211, N1055, N1379);
and AND2 (N1476, N1457, N1009);
xor XOR2 (N1477, N1467, N711);
xor XOR2 (N1478, N1472, N690);
xor XOR2 (N1479, N1466, N1112);
buf BUF1 (N1480, N1453);
and AND3 (N1481, N1479, N786, N771);
xor XOR2 (N1482, N1456, N29);
buf BUF1 (N1483, N1468);
not NOT1 (N1484, N1473);
nor NOR4 (N1485, N1475, N505, N520, N461);
and AND3 (N1486, N1477, N293, N702);
and AND4 (N1487, N1481, N1077, N257, N463);
not NOT1 (N1488, N1482);
buf BUF1 (N1489, N1485);
buf BUF1 (N1490, N1489);
xor XOR2 (N1491, N1480, N1206);
or OR2 (N1492, N1483, N105);
buf BUF1 (N1493, N1478);
buf BUF1 (N1494, N1493);
and AND4 (N1495, N1494, N1065, N1042, N1326);
or OR3 (N1496, N1488, N185, N468);
or OR2 (N1497, N1476, N885);
not NOT1 (N1498, N1471);
and AND4 (N1499, N1495, N260, N1007, N758);
xor XOR2 (N1500, N1490, N366);
xor XOR2 (N1501, N1486, N899);
or OR4 (N1502, N1484, N146, N1478, N414);
and AND3 (N1503, N1491, N483, N922);
xor XOR2 (N1504, N1500, N720);
and AND3 (N1505, N1502, N7, N390);
nor NOR3 (N1506, N1487, N445, N1269);
or OR2 (N1507, N1499, N605);
buf BUF1 (N1508, N1501);
buf BUF1 (N1509, N1496);
xor XOR2 (N1510, N1503, N280);
xor XOR2 (N1511, N1510, N1046);
xor XOR2 (N1512, N1507, N1340);
or OR4 (N1513, N1505, N774, N1315, N1285);
not NOT1 (N1514, N1506);
or OR2 (N1515, N1509, N429);
and AND2 (N1516, N1514, N1040);
and AND2 (N1517, N1497, N93);
xor XOR2 (N1518, N1504, N1380);
xor XOR2 (N1519, N1518, N764);
nand NAND3 (N1520, N1508, N1172, N573);
and AND2 (N1521, N1492, N784);
buf BUF1 (N1522, N1515);
xor XOR2 (N1523, N1522, N1062);
xor XOR2 (N1524, N1512, N347);
xor XOR2 (N1525, N1524, N1204);
not NOT1 (N1526, N1511);
and AND3 (N1527, N1519, N1515, N853);
not NOT1 (N1528, N1498);
nor NOR3 (N1529, N1516, N10, N1449);
nor NOR2 (N1530, N1521, N155);
buf BUF1 (N1531, N1529);
nor NOR3 (N1532, N1531, N466, N1463);
nand NAND2 (N1533, N1528, N1122);
nor NOR2 (N1534, N1526, N981);
or OR3 (N1535, N1532, N1295, N1369);
and AND4 (N1536, N1530, N1303, N1408, N1449);
xor XOR2 (N1537, N1535, N946);
not NOT1 (N1538, N1520);
or OR3 (N1539, N1534, N97, N360);
nand NAND2 (N1540, N1517, N164);
or OR3 (N1541, N1538, N904, N436);
not NOT1 (N1542, N1523);
not NOT1 (N1543, N1540);
or OR3 (N1544, N1542, N746, N889);
xor XOR2 (N1545, N1537, N1194);
and AND3 (N1546, N1525, N743, N1286);
or OR3 (N1547, N1546, N1486, N1015);
or OR4 (N1548, N1536, N1419, N844, N1358);
buf BUF1 (N1549, N1543);
and AND3 (N1550, N1541, N1141, N1173);
not NOT1 (N1551, N1549);
not NOT1 (N1552, N1545);
not NOT1 (N1553, N1547);
nand NAND2 (N1554, N1533, N553);
nand NAND3 (N1555, N1539, N918, N162);
or OR4 (N1556, N1550, N794, N1184, N190);
and AND3 (N1557, N1555, N924, N383);
or OR3 (N1558, N1553, N1204, N235);
not NOT1 (N1559, N1554);
nand NAND3 (N1560, N1559, N757, N1395);
nor NOR2 (N1561, N1513, N804);
nand NAND4 (N1562, N1556, N648, N496, N841);
xor XOR2 (N1563, N1562, N1202);
and AND4 (N1564, N1558, N1427, N1436, N1015);
buf BUF1 (N1565, N1561);
not NOT1 (N1566, N1563);
buf BUF1 (N1567, N1564);
buf BUF1 (N1568, N1544);
or OR3 (N1569, N1527, N59, N742);
nor NOR2 (N1570, N1568, N141);
and AND3 (N1571, N1548, N546, N212);
nor NOR4 (N1572, N1565, N1239, N1371, N1569);
not NOT1 (N1573, N1046);
and AND4 (N1574, N1557, N27, N318, N1322);
buf BUF1 (N1575, N1570);
or OR2 (N1576, N1560, N867);
buf BUF1 (N1577, N1575);
nand NAND4 (N1578, N1566, N1359, N318, N762);
buf BUF1 (N1579, N1578);
nor NOR3 (N1580, N1576, N766, N771);
nand NAND3 (N1581, N1579, N629, N611);
and AND3 (N1582, N1580, N590, N310);
or OR3 (N1583, N1574, N1492, N767);
buf BUF1 (N1584, N1551);
not NOT1 (N1585, N1572);
buf BUF1 (N1586, N1573);
nand NAND3 (N1587, N1581, N521, N801);
not NOT1 (N1588, N1577);
xor XOR2 (N1589, N1588, N839);
and AND4 (N1590, N1584, N520, N924, N1217);
nand NAND4 (N1591, N1552, N1344, N1010, N388);
xor XOR2 (N1592, N1590, N330);
nor NOR4 (N1593, N1571, N457, N180, N434);
nor NOR3 (N1594, N1592, N199, N730);
nor NOR2 (N1595, N1594, N350);
not NOT1 (N1596, N1582);
nand NAND4 (N1597, N1596, N181, N1505, N702);
or OR2 (N1598, N1585, N371);
and AND3 (N1599, N1586, N1053, N214);
or OR2 (N1600, N1598, N1567);
and AND2 (N1601, N773, N790);
buf BUF1 (N1602, N1593);
and AND3 (N1603, N1602, N654, N1377);
buf BUF1 (N1604, N1591);
not NOT1 (N1605, N1601);
not NOT1 (N1606, N1589);
or OR3 (N1607, N1603, N306, N262);
and AND4 (N1608, N1606, N1567, N670, N760);
not NOT1 (N1609, N1604);
xor XOR2 (N1610, N1605, N852);
or OR2 (N1611, N1583, N878);
buf BUF1 (N1612, N1609);
nand NAND2 (N1613, N1611, N629);
and AND2 (N1614, N1595, N1333);
and AND4 (N1615, N1608, N499, N194, N981);
nor NOR2 (N1616, N1615, N92);
nor NOR3 (N1617, N1612, N482, N325);
nand NAND2 (N1618, N1613, N823);
buf BUF1 (N1619, N1599);
xor XOR2 (N1620, N1617, N887);
buf BUF1 (N1621, N1619);
and AND4 (N1622, N1600, N1135, N425, N1609);
not NOT1 (N1623, N1620);
and AND2 (N1624, N1621, N1469);
buf BUF1 (N1625, N1623);
not NOT1 (N1626, N1616);
xor XOR2 (N1627, N1625, N491);
nor NOR4 (N1628, N1587, N1550, N764, N1406);
xor XOR2 (N1629, N1628, N910);
xor XOR2 (N1630, N1607, N899);
and AND4 (N1631, N1624, N1462, N436, N43);
xor XOR2 (N1632, N1614, N465);
xor XOR2 (N1633, N1597, N1120);
buf BUF1 (N1634, N1630);
and AND3 (N1635, N1627, N1393, N996);
and AND4 (N1636, N1629, N1400, N419, N969);
xor XOR2 (N1637, N1633, N1530);
buf BUF1 (N1638, N1632);
xor XOR2 (N1639, N1638, N612);
xor XOR2 (N1640, N1622, N186);
not NOT1 (N1641, N1640);
nand NAND4 (N1642, N1610, N21, N876, N542);
xor XOR2 (N1643, N1626, N30);
and AND4 (N1644, N1618, N1453, N486, N326);
not NOT1 (N1645, N1636);
nor NOR4 (N1646, N1639, N609, N1154, N670);
nand NAND2 (N1647, N1646, N707);
or OR4 (N1648, N1643, N1156, N981, N1389);
not NOT1 (N1649, N1631);
nand NAND3 (N1650, N1645, N90, N1513);
not NOT1 (N1651, N1649);
and AND3 (N1652, N1651, N587, N356);
nand NAND2 (N1653, N1635, N1391);
and AND4 (N1654, N1653, N1400, N317, N1089);
buf BUF1 (N1655, N1634);
nor NOR4 (N1656, N1654, N658, N3, N242);
nand NAND3 (N1657, N1648, N1346, N293);
or OR2 (N1658, N1657, N80);
xor XOR2 (N1659, N1652, N93);
not NOT1 (N1660, N1637);
not NOT1 (N1661, N1656);
xor XOR2 (N1662, N1641, N1164);
buf BUF1 (N1663, N1662);
and AND2 (N1664, N1660, N68);
nand NAND4 (N1665, N1664, N220, N1656, N732);
nand NAND3 (N1666, N1659, N864, N713);
and AND2 (N1667, N1647, N186);
nor NOR4 (N1668, N1644, N499, N579, N1146);
nand NAND4 (N1669, N1661, N465, N537, N1509);
buf BUF1 (N1670, N1642);
nor NOR2 (N1671, N1665, N472);
buf BUF1 (N1672, N1671);
xor XOR2 (N1673, N1663, N362);
not NOT1 (N1674, N1670);
nor NOR2 (N1675, N1667, N1565);
xor XOR2 (N1676, N1673, N71);
and AND3 (N1677, N1666, N1228, N162);
not NOT1 (N1678, N1676);
nand NAND2 (N1679, N1674, N900);
xor XOR2 (N1680, N1668, N355);
nand NAND3 (N1681, N1669, N381, N1116);
nor NOR2 (N1682, N1678, N778);
xor XOR2 (N1683, N1681, N282);
not NOT1 (N1684, N1672);
xor XOR2 (N1685, N1675, N672);
nor NOR2 (N1686, N1682, N1543);
not NOT1 (N1687, N1686);
and AND2 (N1688, N1687, N1252);
and AND3 (N1689, N1679, N610, N425);
nor NOR2 (N1690, N1689, N1087);
nor NOR2 (N1691, N1677, N1682);
xor XOR2 (N1692, N1683, N360);
buf BUF1 (N1693, N1650);
buf BUF1 (N1694, N1690);
buf BUF1 (N1695, N1684);
nor NOR2 (N1696, N1658, N851);
buf BUF1 (N1697, N1691);
or OR3 (N1698, N1694, N1511, N1139);
or OR3 (N1699, N1698, N1230, N235);
buf BUF1 (N1700, N1699);
buf BUF1 (N1701, N1685);
or OR3 (N1702, N1680, N1377, N1406);
buf BUF1 (N1703, N1688);
not NOT1 (N1704, N1693);
buf BUF1 (N1705, N1692);
nor NOR3 (N1706, N1696, N540, N537);
xor XOR2 (N1707, N1655, N1588);
nand NAND2 (N1708, N1704, N223);
xor XOR2 (N1709, N1703, N1388);
buf BUF1 (N1710, N1707);
not NOT1 (N1711, N1710);
buf BUF1 (N1712, N1705);
nor NOR4 (N1713, N1701, N1360, N320, N472);
xor XOR2 (N1714, N1708, N460);
xor XOR2 (N1715, N1702, N1146);
xor XOR2 (N1716, N1711, N535);
nor NOR4 (N1717, N1700, N901, N302, N993);
nor NOR2 (N1718, N1697, N338);
buf BUF1 (N1719, N1706);
not NOT1 (N1720, N1715);
and AND2 (N1721, N1714, N1458);
not NOT1 (N1722, N1719);
buf BUF1 (N1723, N1717);
and AND3 (N1724, N1722, N215, N1445);
nand NAND4 (N1725, N1721, N578, N1335, N970);
buf BUF1 (N1726, N1712);
buf BUF1 (N1727, N1716);
and AND3 (N1728, N1724, N1601, N1592);
nand NAND4 (N1729, N1728, N650, N1540, N108);
xor XOR2 (N1730, N1729, N166);
and AND2 (N1731, N1727, N1255);
not NOT1 (N1732, N1730);
or OR3 (N1733, N1731, N643, N727);
xor XOR2 (N1734, N1723, N219);
and AND4 (N1735, N1713, N1043, N810, N719);
and AND2 (N1736, N1695, N597);
nand NAND4 (N1737, N1709, N182, N16, N54);
nand NAND2 (N1738, N1735, N1092);
xor XOR2 (N1739, N1726, N891);
nor NOR2 (N1740, N1738, N423);
nor NOR4 (N1741, N1737, N44, N1382, N1140);
xor XOR2 (N1742, N1720, N1384);
nor NOR3 (N1743, N1736, N1669, N1555);
xor XOR2 (N1744, N1725, N1235);
nand NAND2 (N1745, N1744, N473);
nor NOR3 (N1746, N1739, N427, N987);
nor NOR3 (N1747, N1743, N1079, N1537);
or OR3 (N1748, N1741, N474, N935);
buf BUF1 (N1749, N1746);
nor NOR4 (N1750, N1740, N622, N338, N1273);
or OR2 (N1751, N1749, N1579);
and AND2 (N1752, N1750, N1243);
nor NOR3 (N1753, N1742, N709, N1132);
xor XOR2 (N1754, N1745, N187);
nand NAND3 (N1755, N1718, N1746, N577);
and AND4 (N1756, N1747, N939, N500, N178);
or OR4 (N1757, N1751, N644, N626, N417);
buf BUF1 (N1758, N1756);
and AND3 (N1759, N1734, N638, N758);
not NOT1 (N1760, N1732);
not NOT1 (N1761, N1733);
not NOT1 (N1762, N1755);
or OR3 (N1763, N1754, N1111, N682);
nand NAND4 (N1764, N1759, N286, N679, N770);
nand NAND3 (N1765, N1753, N722, N1333);
nor NOR4 (N1766, N1757, N773, N520, N1319);
not NOT1 (N1767, N1766);
or OR4 (N1768, N1765, N950, N1291, N1340);
buf BUF1 (N1769, N1768);
and AND3 (N1770, N1763, N1009, N894);
not NOT1 (N1771, N1770);
and AND3 (N1772, N1760, N389, N1282);
nor NOR2 (N1773, N1748, N741);
and AND4 (N1774, N1769, N48, N1729, N1359);
nand NAND2 (N1775, N1772, N1171);
xor XOR2 (N1776, N1767, N1344);
nand NAND4 (N1777, N1758, N513, N938, N1182);
nand NAND2 (N1778, N1762, N1517);
nor NOR4 (N1779, N1773, N1731, N80, N1155);
not NOT1 (N1780, N1776);
or OR4 (N1781, N1775, N500, N103, N712);
nor NOR3 (N1782, N1764, N1223, N685);
xor XOR2 (N1783, N1779, N441);
not NOT1 (N1784, N1774);
and AND3 (N1785, N1778, N1760, N1382);
not NOT1 (N1786, N1781);
nand NAND4 (N1787, N1752, N1243, N1265, N887);
or OR2 (N1788, N1783, N836);
xor XOR2 (N1789, N1777, N461);
buf BUF1 (N1790, N1784);
nor NOR3 (N1791, N1787, N1313, N754);
xor XOR2 (N1792, N1782, N1280);
xor XOR2 (N1793, N1785, N369);
not NOT1 (N1794, N1793);
buf BUF1 (N1795, N1786);
nor NOR2 (N1796, N1761, N1060);
not NOT1 (N1797, N1790);
xor XOR2 (N1798, N1780, N1535);
nand NAND4 (N1799, N1791, N397, N1507, N184);
xor XOR2 (N1800, N1797, N280);
or OR4 (N1801, N1789, N1755, N1136, N1440);
buf BUF1 (N1802, N1788);
xor XOR2 (N1803, N1798, N1207);
xor XOR2 (N1804, N1796, N728);
nor NOR2 (N1805, N1799, N884);
not NOT1 (N1806, N1800);
not NOT1 (N1807, N1794);
nand NAND3 (N1808, N1806, N1250, N860);
not NOT1 (N1809, N1792);
xor XOR2 (N1810, N1809, N160);
and AND2 (N1811, N1771, N575);
buf BUF1 (N1812, N1802);
xor XOR2 (N1813, N1807, N236);
nand NAND3 (N1814, N1805, N1410, N1069);
buf BUF1 (N1815, N1814);
nor NOR3 (N1816, N1795, N1529, N1695);
not NOT1 (N1817, N1813);
nand NAND2 (N1818, N1810, N821);
nand NAND3 (N1819, N1815, N319, N182);
xor XOR2 (N1820, N1804, N651);
not NOT1 (N1821, N1812);
xor XOR2 (N1822, N1817, N1432);
xor XOR2 (N1823, N1811, N928);
xor XOR2 (N1824, N1823, N870);
nand NAND3 (N1825, N1819, N411, N771);
nand NAND2 (N1826, N1803, N1174);
nor NOR2 (N1827, N1808, N1222);
xor XOR2 (N1828, N1818, N1095);
nor NOR4 (N1829, N1816, N1602, N1485, N1627);
not NOT1 (N1830, N1828);
xor XOR2 (N1831, N1825, N1517);
or OR2 (N1832, N1821, N920);
xor XOR2 (N1833, N1820, N740);
nand NAND2 (N1834, N1832, N43);
nor NOR3 (N1835, N1822, N1550, N518);
nand NAND2 (N1836, N1831, N492);
not NOT1 (N1837, N1801);
nor NOR2 (N1838, N1829, N884);
not NOT1 (N1839, N1824);
xor XOR2 (N1840, N1837, N498);
not NOT1 (N1841, N1833);
not NOT1 (N1842, N1840);
not NOT1 (N1843, N1827);
and AND4 (N1844, N1842, N879, N247, N1585);
xor XOR2 (N1845, N1843, N306);
and AND3 (N1846, N1835, N1229, N600);
nor NOR4 (N1847, N1830, N939, N1051, N1390);
xor XOR2 (N1848, N1844, N266);
and AND3 (N1849, N1847, N881, N1546);
nor NOR2 (N1850, N1826, N1034);
nand NAND4 (N1851, N1836, N1576, N1453, N891);
nand NAND4 (N1852, N1851, N259, N1676, N883);
buf BUF1 (N1853, N1848);
or OR3 (N1854, N1853, N1826, N878);
buf BUF1 (N1855, N1849);
or OR4 (N1856, N1850, N1030, N1297, N662);
or OR2 (N1857, N1856, N1136);
or OR4 (N1858, N1839, N245, N1535, N12);
nor NOR4 (N1859, N1854, N1450, N977, N80);
xor XOR2 (N1860, N1841, N1408);
nand NAND2 (N1861, N1838, N1428);
buf BUF1 (N1862, N1858);
or OR2 (N1863, N1834, N259);
xor XOR2 (N1864, N1862, N891);
and AND4 (N1865, N1855, N267, N48, N700);
xor XOR2 (N1866, N1864, N138);
nor NOR3 (N1867, N1860, N447, N939);
xor XOR2 (N1868, N1846, N1048);
nor NOR3 (N1869, N1867, N965, N20);
xor XOR2 (N1870, N1868, N1094);
buf BUF1 (N1871, N1866);
or OR4 (N1872, N1857, N993, N113, N919);
not NOT1 (N1873, N1871);
nor NOR2 (N1874, N1865, N1790);
or OR4 (N1875, N1861, N1020, N256, N1586);
and AND4 (N1876, N1869, N607, N1035, N860);
not NOT1 (N1877, N1875);
nand NAND4 (N1878, N1872, N1869, N976, N1333);
buf BUF1 (N1879, N1873);
xor XOR2 (N1880, N1852, N948);
nor NOR4 (N1881, N1879, N748, N1195, N1163);
or OR3 (N1882, N1877, N1005, N1660);
nand NAND4 (N1883, N1845, N1758, N247, N1588);
or OR4 (N1884, N1874, N1874, N1, N1116);
or OR4 (N1885, N1878, N460, N15, N1539);
nor NOR2 (N1886, N1876, N433);
not NOT1 (N1887, N1881);
xor XOR2 (N1888, N1885, N1023);
xor XOR2 (N1889, N1870, N1037);
nor NOR2 (N1890, N1886, N1685);
or OR3 (N1891, N1882, N88, N1253);
and AND3 (N1892, N1888, N768, N1301);
and AND4 (N1893, N1891, N963, N1276, N760);
and AND2 (N1894, N1889, N1049);
buf BUF1 (N1895, N1859);
and AND3 (N1896, N1890, N1759, N1867);
buf BUF1 (N1897, N1884);
nand NAND3 (N1898, N1883, N1774, N1368);
or OR3 (N1899, N1898, N478, N889);
and AND4 (N1900, N1893, N990, N1764, N371);
and AND2 (N1901, N1896, N535);
not NOT1 (N1902, N1900);
or OR2 (N1903, N1894, N1532);
not NOT1 (N1904, N1897);
xor XOR2 (N1905, N1895, N771);
nor NOR3 (N1906, N1903, N711, N1883);
nor NOR2 (N1907, N1902, N1800);
and AND3 (N1908, N1904, N1172, N841);
and AND4 (N1909, N1901, N1617, N580, N1321);
or OR4 (N1910, N1863, N929, N857, N1552);
not NOT1 (N1911, N1892);
buf BUF1 (N1912, N1906);
nor NOR2 (N1913, N1899, N1061);
buf BUF1 (N1914, N1911);
not NOT1 (N1915, N1907);
nand NAND2 (N1916, N1914, N1533);
nor NOR2 (N1917, N1912, N1101);
not NOT1 (N1918, N1915);
not NOT1 (N1919, N1916);
not NOT1 (N1920, N1887);
xor XOR2 (N1921, N1905, N1787);
buf BUF1 (N1922, N1909);
not NOT1 (N1923, N1910);
or OR4 (N1924, N1918, N1326, N1843, N604);
xor XOR2 (N1925, N1924, N4);
and AND2 (N1926, N1908, N1499);
buf BUF1 (N1927, N1926);
nand NAND3 (N1928, N1927, N1205, N1305);
nand NAND4 (N1929, N1919, N1131, N1758, N1654);
and AND4 (N1930, N1920, N1843, N978, N577);
nand NAND3 (N1931, N1928, N1742, N75);
not NOT1 (N1932, N1922);
or OR3 (N1933, N1930, N1338, N1529);
not NOT1 (N1934, N1913);
or OR2 (N1935, N1925, N791);
xor XOR2 (N1936, N1932, N539);
not NOT1 (N1937, N1880);
buf BUF1 (N1938, N1936);
nor NOR4 (N1939, N1934, N1850, N1114, N61);
xor XOR2 (N1940, N1929, N466);
and AND2 (N1941, N1937, N1054);
nand NAND4 (N1942, N1938, N951, N1095, N466);
and AND4 (N1943, N1923, N549, N106, N1625);
nand NAND2 (N1944, N1940, N281);
nand NAND3 (N1945, N1939, N402, N1893);
buf BUF1 (N1946, N1945);
and AND2 (N1947, N1917, N413);
and AND2 (N1948, N1942, N921);
buf BUF1 (N1949, N1935);
nor NOR2 (N1950, N1931, N184);
or OR4 (N1951, N1943, N377, N857, N116);
nand NAND2 (N1952, N1946, N227);
nand NAND3 (N1953, N1947, N1533, N558);
not NOT1 (N1954, N1948);
or OR2 (N1955, N1954, N1493);
and AND2 (N1956, N1933, N1467);
and AND4 (N1957, N1950, N456, N216, N338);
and AND2 (N1958, N1957, N820);
and AND3 (N1959, N1952, N1796, N277);
nand NAND3 (N1960, N1951, N1406, N386);
xor XOR2 (N1961, N1960, N1081);
nor NOR4 (N1962, N1949, N133, N116, N1460);
and AND3 (N1963, N1953, N184, N887);
not NOT1 (N1964, N1956);
and AND4 (N1965, N1944, N1518, N1110, N1720);
not NOT1 (N1966, N1965);
or OR4 (N1967, N1963, N619, N1185, N909);
nand NAND4 (N1968, N1961, N1784, N1214, N1723);
nand NAND4 (N1969, N1964, N1761, N392, N104);
and AND4 (N1970, N1968, N489, N278, N1727);
and AND3 (N1971, N1959, N306, N1724);
nand NAND2 (N1972, N1941, N34);
or OR2 (N1973, N1970, N1385);
nor NOR2 (N1974, N1971, N566);
and AND4 (N1975, N1969, N1429, N912, N820);
xor XOR2 (N1976, N1973, N716);
nand NAND2 (N1977, N1966, N906);
or OR3 (N1978, N1977, N359, N1676);
xor XOR2 (N1979, N1978, N348);
xor XOR2 (N1980, N1974, N159);
buf BUF1 (N1981, N1955);
or OR4 (N1982, N1962, N892, N1242, N1827);
buf BUF1 (N1983, N1980);
buf BUF1 (N1984, N1982);
buf BUF1 (N1985, N1981);
or OR4 (N1986, N1985, N1523, N833, N515);
xor XOR2 (N1987, N1983, N1421);
nand NAND3 (N1988, N1984, N792, N657);
nand NAND3 (N1989, N1976, N1579, N581);
or OR2 (N1990, N1989, N803);
nor NOR4 (N1991, N1990, N916, N308, N1162);
nand NAND3 (N1992, N1921, N1863, N401);
nor NOR3 (N1993, N1992, N1919, N728);
nor NOR4 (N1994, N1979, N1364, N1406, N705);
buf BUF1 (N1995, N1967);
or OR3 (N1996, N1972, N1540, N1027);
xor XOR2 (N1997, N1975, N914);
not NOT1 (N1998, N1987);
xor XOR2 (N1999, N1994, N974);
and AND3 (N2000, N1997, N860, N1867);
nor NOR4 (N2001, N1988, N966, N1715, N715);
nand NAND4 (N2002, N1991, N1853, N306, N705);
xor XOR2 (N2003, N1999, N432);
buf BUF1 (N2004, N1995);
and AND2 (N2005, N2004, N1100);
nand NAND4 (N2006, N1996, N834, N1043, N1641);
not NOT1 (N2007, N2000);
nand NAND3 (N2008, N1998, N205, N1826);
buf BUF1 (N2009, N1993);
nor NOR4 (N2010, N2006, N131, N1865, N9);
not NOT1 (N2011, N2001);
and AND2 (N2012, N1986, N1676);
nand NAND3 (N2013, N2005, N1224, N1388);
not NOT1 (N2014, N2003);
nor NOR4 (N2015, N2014, N1485, N586, N373);
or OR3 (N2016, N1958, N1016, N376);
buf BUF1 (N2017, N2002);
nand NAND2 (N2018, N2016, N885);
not NOT1 (N2019, N2009);
and AND4 (N2020, N2015, N1849, N1786, N1338);
buf BUF1 (N2021, N2007);
buf BUF1 (N2022, N2021);
xor XOR2 (N2023, N2013, N1087);
nor NOR4 (N2024, N2022, N595, N47, N1429);
buf BUF1 (N2025, N2020);
not NOT1 (N2026, N2019);
or OR4 (N2027, N2018, N1819, N738, N157);
or OR3 (N2028, N2024, N1291, N1632);
not NOT1 (N2029, N2023);
xor XOR2 (N2030, N2027, N1085);
not NOT1 (N2031, N2017);
and AND4 (N2032, N2031, N1064, N1307, N604);
buf BUF1 (N2033, N2012);
or OR4 (N2034, N2030, N259, N357, N1926);
or OR4 (N2035, N2011, N1803, N471, N605);
xor XOR2 (N2036, N2033, N1807);
or OR2 (N2037, N2008, N1440);
buf BUF1 (N2038, N2034);
not NOT1 (N2039, N2036);
or OR3 (N2040, N2037, N466, N4);
nand NAND2 (N2041, N2038, N1620);
nor NOR4 (N2042, N2025, N1256, N1733, N65);
not NOT1 (N2043, N2028);
nand NAND3 (N2044, N2043, N1537, N798);
nand NAND4 (N2045, N2042, N555, N1306, N937);
and AND3 (N2046, N2029, N874, N457);
nor NOR2 (N2047, N2026, N1971);
xor XOR2 (N2048, N2041, N897);
nand NAND2 (N2049, N2045, N1762);
xor XOR2 (N2050, N2048, N1260);
not NOT1 (N2051, N2050);
not NOT1 (N2052, N2051);
nand NAND3 (N2053, N2035, N15, N1023);
and AND2 (N2054, N2044, N1255);
nand NAND3 (N2055, N2040, N950, N935);
nor NOR3 (N2056, N2053, N967, N305);
buf BUF1 (N2057, N2046);
buf BUF1 (N2058, N2055);
xor XOR2 (N2059, N2049, N1157);
nand NAND3 (N2060, N2059, N1468, N1167);
or OR3 (N2061, N2058, N696, N1351);
and AND4 (N2062, N2047, N243, N312, N743);
or OR3 (N2063, N2054, N1028, N1848);
nor NOR4 (N2064, N2052, N659, N843, N380);
xor XOR2 (N2065, N2039, N573);
xor XOR2 (N2066, N2063, N821);
and AND3 (N2067, N2032, N362, N584);
buf BUF1 (N2068, N2065);
buf BUF1 (N2069, N2068);
not NOT1 (N2070, N2061);
xor XOR2 (N2071, N2066, N1152);
nor NOR3 (N2072, N2056, N340, N348);
nand NAND2 (N2073, N2010, N925);
buf BUF1 (N2074, N2071);
or OR2 (N2075, N2060, N333);
nand NAND3 (N2076, N2062, N1003, N414);
and AND4 (N2077, N2073, N158, N260, N1183);
nand NAND2 (N2078, N2057, N1581);
not NOT1 (N2079, N2078);
and AND4 (N2080, N2077, N1060, N888, N875);
and AND2 (N2081, N2075, N478);
nor NOR4 (N2082, N2076, N1581, N915, N758);
nand NAND2 (N2083, N2074, N1792);
or OR4 (N2084, N2082, N2028, N243, N590);
nor NOR4 (N2085, N2069, N1897, N1147, N1284);
not NOT1 (N2086, N2064);
nor NOR4 (N2087, N2079, N520, N855, N1439);
and AND4 (N2088, N2083, N1891, N1024, N1408);
and AND3 (N2089, N2085, N242, N461);
and AND2 (N2090, N2080, N1796);
not NOT1 (N2091, N2090);
buf BUF1 (N2092, N2088);
xor XOR2 (N2093, N2067, N1519);
and AND3 (N2094, N2087, N302, N208);
and AND4 (N2095, N2084, N723, N1990, N1979);
nor NOR4 (N2096, N2091, N151, N1316, N59);
xor XOR2 (N2097, N2081, N1434);
nand NAND3 (N2098, N2086, N1935, N1699);
nand NAND3 (N2099, N2070, N1358, N1498);
and AND4 (N2100, N2098, N650, N1718, N180);
nor NOR4 (N2101, N2100, N1810, N1373, N538);
or OR4 (N2102, N2099, N1116, N445, N1753);
and AND3 (N2103, N2093, N1304, N1753);
nor NOR2 (N2104, N2095, N197);
not NOT1 (N2105, N2089);
not NOT1 (N2106, N2104);
or OR4 (N2107, N2102, N377, N1848, N1630);
not NOT1 (N2108, N2103);
nand NAND2 (N2109, N2094, N536);
or OR2 (N2110, N2105, N19);
nand NAND3 (N2111, N2106, N366, N687);
nor NOR3 (N2112, N2096, N868, N1648);
nand NAND4 (N2113, N2109, N982, N1721, N526);
not NOT1 (N2114, N2108);
or OR4 (N2115, N2101, N2083, N28, N66);
and AND4 (N2116, N2115, N753, N1129, N1283);
or OR2 (N2117, N2092, N1704);
xor XOR2 (N2118, N2107, N1746);
xor XOR2 (N2119, N2072, N1693);
nor NOR4 (N2120, N2111, N1406, N451, N1871);
xor XOR2 (N2121, N2097, N1343);
nor NOR4 (N2122, N2114, N1584, N377, N820);
nand NAND4 (N2123, N2116, N887, N1121, N2017);
and AND2 (N2124, N2110, N1811);
nand NAND4 (N2125, N2117, N882, N107, N1546);
or OR2 (N2126, N2123, N2074);
or OR3 (N2127, N2118, N1104, N1885);
nor NOR4 (N2128, N2121, N660, N2092, N1329);
nand NAND4 (N2129, N2124, N1431, N853, N581);
nor NOR4 (N2130, N2129, N1803, N1794, N633);
not NOT1 (N2131, N2119);
not NOT1 (N2132, N2128);
not NOT1 (N2133, N2122);
and AND3 (N2134, N2125, N74, N2101);
xor XOR2 (N2135, N2112, N67);
nor NOR2 (N2136, N2113, N1327);
nor NOR4 (N2137, N2126, N457, N184, N702);
and AND4 (N2138, N2137, N169, N205, N480);
xor XOR2 (N2139, N2135, N1185);
buf BUF1 (N2140, N2132);
nand NAND4 (N2141, N2131, N320, N1694, N1079);
not NOT1 (N2142, N2130);
buf BUF1 (N2143, N2138);
nor NOR3 (N2144, N2134, N1283, N1052);
xor XOR2 (N2145, N2143, N112);
or OR4 (N2146, N2144, N304, N1302, N1177);
xor XOR2 (N2147, N2141, N2140);
buf BUF1 (N2148, N660);
xor XOR2 (N2149, N2147, N749);
nor NOR4 (N2150, N2127, N1624, N2096, N1188);
or OR3 (N2151, N2133, N1719, N1945);
xor XOR2 (N2152, N2120, N343);
buf BUF1 (N2153, N2150);
and AND4 (N2154, N2153, N1970, N1524, N169);
nor NOR4 (N2155, N2154, N1419, N940, N647);
not NOT1 (N2156, N2149);
nor NOR2 (N2157, N2155, N1297);
buf BUF1 (N2158, N2142);
or OR2 (N2159, N2151, N1359);
not NOT1 (N2160, N2136);
and AND2 (N2161, N2159, N358);
not NOT1 (N2162, N2139);
nand NAND2 (N2163, N2160, N242);
buf BUF1 (N2164, N2152);
xor XOR2 (N2165, N2148, N259);
xor XOR2 (N2166, N2162, N434);
xor XOR2 (N2167, N2145, N768);
buf BUF1 (N2168, N2161);
xor XOR2 (N2169, N2168, N1418);
nor NOR4 (N2170, N2163, N188, N842, N1530);
or OR2 (N2171, N2158, N331);
nor NOR2 (N2172, N2169, N11);
nand NAND2 (N2173, N2164, N921);
nand NAND3 (N2174, N2157, N945, N2121);
nor NOR3 (N2175, N2173, N1161, N931);
not NOT1 (N2176, N2156);
xor XOR2 (N2177, N2175, N1622);
and AND4 (N2178, N2167, N284, N1505, N588);
buf BUF1 (N2179, N2176);
and AND2 (N2180, N2172, N539);
and AND2 (N2181, N2171, N2028);
or OR4 (N2182, N2181, N2010, N2135, N1863);
nand NAND3 (N2183, N2170, N1284, N173);
or OR4 (N2184, N2183, N1617, N27, N1740);
nand NAND3 (N2185, N2179, N1614, N2041);
buf BUF1 (N2186, N2177);
or OR4 (N2187, N2165, N732, N1597, N1549);
nand NAND4 (N2188, N2166, N1913, N2098, N2150);
nor NOR2 (N2189, N2188, N757);
and AND2 (N2190, N2186, N1567);
nor NOR2 (N2191, N2180, N1639);
xor XOR2 (N2192, N2185, N953);
not NOT1 (N2193, N2184);
and AND4 (N2194, N2187, N1881, N903, N388);
or OR4 (N2195, N2191, N153, N1000, N42);
and AND3 (N2196, N2193, N1920, N2005);
or OR2 (N2197, N2146, N948);
nor NOR2 (N2198, N2190, N2064);
xor XOR2 (N2199, N2197, N922);
nor NOR2 (N2200, N2189, N582);
nand NAND2 (N2201, N2192, N1617);
and AND4 (N2202, N2198, N1352, N863, N1687);
nand NAND4 (N2203, N2200, N1806, N20, N2172);
buf BUF1 (N2204, N2203);
buf BUF1 (N2205, N2182);
xor XOR2 (N2206, N2195, N616);
and AND2 (N2207, N2199, N290);
or OR3 (N2208, N2205, N577, N186);
or OR2 (N2209, N2201, N1533);
nand NAND2 (N2210, N2194, N1501);
nor NOR3 (N2211, N2174, N1562, N986);
and AND3 (N2212, N2206, N673, N876);
and AND4 (N2213, N2211, N1812, N324, N1346);
xor XOR2 (N2214, N2204, N320);
xor XOR2 (N2215, N2212, N352);
and AND4 (N2216, N2196, N2043, N490, N30);
or OR4 (N2217, N2210, N1000, N1360, N356);
buf BUF1 (N2218, N2213);
or OR3 (N2219, N2214, N1880, N1040);
xor XOR2 (N2220, N2207, N1780);
not NOT1 (N2221, N2217);
not NOT1 (N2222, N2219);
xor XOR2 (N2223, N2208, N1484);
and AND2 (N2224, N2221, N606);
buf BUF1 (N2225, N2224);
xor XOR2 (N2226, N2202, N1449);
or OR2 (N2227, N2178, N2006);
buf BUF1 (N2228, N2215);
nor NOR2 (N2229, N2226, N1146);
or OR3 (N2230, N2223, N277, N1170);
xor XOR2 (N2231, N2218, N1597);
nor NOR4 (N2232, N2225, N1790, N1968, N1396);
nand NAND2 (N2233, N2222, N965);
nand NAND3 (N2234, N2228, N2185, N408);
or OR2 (N2235, N2234, N1331);
and AND2 (N2236, N2229, N2033);
not NOT1 (N2237, N2230);
not NOT1 (N2238, N2235);
nand NAND4 (N2239, N2236, N1974, N1011, N1635);
not NOT1 (N2240, N2232);
buf BUF1 (N2241, N2220);
nor NOR2 (N2242, N2233, N2083);
not NOT1 (N2243, N2227);
xor XOR2 (N2244, N2209, N401);
not NOT1 (N2245, N2238);
nor NOR4 (N2246, N2237, N385, N2141, N201);
or OR3 (N2247, N2240, N845, N2184);
nor NOR3 (N2248, N2245, N2168, N93);
xor XOR2 (N2249, N2231, N577);
or OR2 (N2250, N2242, N1883);
nand NAND2 (N2251, N2216, N360);
not NOT1 (N2252, N2248);
buf BUF1 (N2253, N2243);
nand NAND2 (N2254, N2250, N956);
and AND2 (N2255, N2241, N1214);
nor NOR4 (N2256, N2246, N1917, N253, N322);
xor XOR2 (N2257, N2251, N1742);
xor XOR2 (N2258, N2252, N2051);
buf BUF1 (N2259, N2247);
xor XOR2 (N2260, N2256, N2030);
not NOT1 (N2261, N2254);
nor NOR2 (N2262, N2261, N1911);
xor XOR2 (N2263, N2262, N1155);
or OR3 (N2264, N2259, N1297, N1665);
and AND4 (N2265, N2263, N540, N403, N1497);
not NOT1 (N2266, N2260);
and AND3 (N2267, N2258, N274, N84);
buf BUF1 (N2268, N2266);
buf BUF1 (N2269, N2268);
and AND3 (N2270, N2265, N1661, N1181);
and AND3 (N2271, N2253, N191, N328);
and AND3 (N2272, N2271, N142, N2202);
xor XOR2 (N2273, N2255, N1239);
nand NAND4 (N2274, N2269, N2150, N979, N753);
nor NOR4 (N2275, N2272, N1559, N600, N2264);
and AND4 (N2276, N681, N539, N1008, N1034);
xor XOR2 (N2277, N2239, N974);
xor XOR2 (N2278, N2270, N1651);
buf BUF1 (N2279, N2257);
nand NAND4 (N2280, N2278, N88, N819, N1683);
buf BUF1 (N2281, N2274);
xor XOR2 (N2282, N2277, N661);
buf BUF1 (N2283, N2282);
buf BUF1 (N2284, N2281);
buf BUF1 (N2285, N2273);
and AND4 (N2286, N2280, N537, N350, N313);
or OR2 (N2287, N2249, N100);
nor NOR4 (N2288, N2283, N59, N1487, N2036);
nor NOR4 (N2289, N2275, N2083, N119, N29);
xor XOR2 (N2290, N2279, N2051);
and AND4 (N2291, N2289, N916, N1417, N161);
or OR4 (N2292, N2288, N1390, N1863, N257);
or OR4 (N2293, N2285, N370, N1298, N1872);
nand NAND3 (N2294, N2267, N1029, N1227);
buf BUF1 (N2295, N2286);
nand NAND3 (N2296, N2292, N869, N757);
or OR2 (N2297, N2295, N1377);
nor NOR4 (N2298, N2290, N808, N445, N685);
xor XOR2 (N2299, N2284, N1125);
and AND4 (N2300, N2244, N567, N319, N1979);
xor XOR2 (N2301, N2297, N1679);
or OR4 (N2302, N2296, N1429, N1557, N1461);
not NOT1 (N2303, N2276);
xor XOR2 (N2304, N2302, N2026);
and AND2 (N2305, N2298, N1124);
nor NOR2 (N2306, N2299, N494);
not NOT1 (N2307, N2304);
nor NOR3 (N2308, N2294, N992, N690);
nor NOR4 (N2309, N2301, N2127, N2179, N1255);
and AND3 (N2310, N2291, N697, N604);
buf BUF1 (N2311, N2287);
nand NAND2 (N2312, N2303, N388);
nand NAND2 (N2313, N2307, N1694);
nand NAND2 (N2314, N2312, N1904);
nor NOR4 (N2315, N2308, N1390, N2002, N311);
or OR2 (N2316, N2313, N961);
nor NOR2 (N2317, N2305, N437);
and AND3 (N2318, N2310, N1685, N729);
or OR2 (N2319, N2311, N1835);
xor XOR2 (N2320, N2306, N149);
and AND3 (N2321, N2320, N1232, N1884);
or OR4 (N2322, N2309, N1324, N428, N734);
and AND4 (N2323, N2314, N1473, N1271, N292);
not NOT1 (N2324, N2300);
nor NOR2 (N2325, N2315, N669);
and AND3 (N2326, N2317, N545, N1129);
buf BUF1 (N2327, N2319);
xor XOR2 (N2328, N2316, N392);
xor XOR2 (N2329, N2328, N1486);
nor NOR3 (N2330, N2321, N1508, N571);
or OR4 (N2331, N2327, N331, N1388, N2287);
buf BUF1 (N2332, N2325);
and AND2 (N2333, N2330, N1865);
xor XOR2 (N2334, N2326, N472);
nand NAND3 (N2335, N2331, N2269, N598);
nor NOR4 (N2336, N2334, N378, N1898, N997);
and AND4 (N2337, N2332, N95, N681, N2062);
nor NOR2 (N2338, N2324, N719);
not NOT1 (N2339, N2293);
xor XOR2 (N2340, N2333, N2339);
or OR2 (N2341, N517, N1767);
xor XOR2 (N2342, N2318, N1113);
and AND2 (N2343, N2323, N988);
buf BUF1 (N2344, N2337);
nor NOR3 (N2345, N2344, N339, N515);
nand NAND2 (N2346, N2329, N442);
xor XOR2 (N2347, N2336, N1253);
nand NAND3 (N2348, N2341, N270, N888);
xor XOR2 (N2349, N2343, N484);
nand NAND4 (N2350, N2348, N2178, N1284, N405);
nor NOR2 (N2351, N2349, N373);
xor XOR2 (N2352, N2342, N2217);
nor NOR3 (N2353, N2351, N1691, N2038);
or OR3 (N2354, N2340, N1140, N1051);
not NOT1 (N2355, N2353);
not NOT1 (N2356, N2335);
and AND3 (N2357, N2354, N1900, N715);
buf BUF1 (N2358, N2338);
or OR4 (N2359, N2352, N1292, N200, N1448);
and AND4 (N2360, N2345, N1357, N710, N1557);
and AND3 (N2361, N2355, N1905, N1975);
buf BUF1 (N2362, N2357);
or OR3 (N2363, N2347, N2082, N2161);
and AND2 (N2364, N2350, N1762);
buf BUF1 (N2365, N2364);
nand NAND2 (N2366, N2365, N1547);
buf BUF1 (N2367, N2359);
buf BUF1 (N2368, N2322);
buf BUF1 (N2369, N2360);
or OR2 (N2370, N2366, N1374);
buf BUF1 (N2371, N2370);
buf BUF1 (N2372, N2367);
not NOT1 (N2373, N2358);
nor NOR2 (N2374, N2361, N766);
nor NOR2 (N2375, N2372, N2033);
nor NOR2 (N2376, N2375, N1204);
nor NOR3 (N2377, N2346, N1337, N1520);
nand NAND2 (N2378, N2369, N1864);
not NOT1 (N2379, N2371);
not NOT1 (N2380, N2374);
buf BUF1 (N2381, N2379);
xor XOR2 (N2382, N2373, N1549);
nor NOR2 (N2383, N2377, N644);
and AND3 (N2384, N2376, N1588, N1877);
xor XOR2 (N2385, N2363, N1544);
nand NAND4 (N2386, N2384, N183, N1874, N1002);
or OR4 (N2387, N2381, N1887, N593, N468);
nor NOR4 (N2388, N2382, N38, N2133, N2322);
not NOT1 (N2389, N2368);
or OR2 (N2390, N2385, N714);
nand NAND4 (N2391, N2387, N1518, N2278, N2290);
nand NAND2 (N2392, N2386, N1092);
not NOT1 (N2393, N2383);
xor XOR2 (N2394, N2389, N761);
or OR2 (N2395, N2378, N895);
and AND2 (N2396, N2394, N2308);
or OR3 (N2397, N2391, N1741, N355);
or OR2 (N2398, N2396, N547);
buf BUF1 (N2399, N2395);
or OR3 (N2400, N2356, N1063, N728);
nand NAND4 (N2401, N2390, N2397, N1776, N1266);
xor XOR2 (N2402, N1163, N1423);
buf BUF1 (N2403, N2362);
xor XOR2 (N2404, N2399, N2104);
xor XOR2 (N2405, N2392, N39);
xor XOR2 (N2406, N2393, N1289);
nand NAND3 (N2407, N2380, N1520, N724);
and AND2 (N2408, N2388, N1079);
xor XOR2 (N2409, N2406, N101);
buf BUF1 (N2410, N2401);
not NOT1 (N2411, N2402);
or OR2 (N2412, N2407, N2115);
nor NOR3 (N2413, N2405, N1911, N1227);
xor XOR2 (N2414, N2409, N773);
nor NOR3 (N2415, N2400, N2132, N1457);
and AND4 (N2416, N2408, N1488, N72, N1361);
nor NOR4 (N2417, N2403, N362, N1870, N1628);
nand NAND4 (N2418, N2415, N1783, N229, N578);
xor XOR2 (N2419, N2417, N2223);
buf BUF1 (N2420, N2413);
nor NOR2 (N2421, N2404, N365);
and AND3 (N2422, N2420, N1492, N1432);
not NOT1 (N2423, N2418);
xor XOR2 (N2424, N2414, N1798);
or OR4 (N2425, N2422, N1521, N2194, N1719);
buf BUF1 (N2426, N2424);
nand NAND3 (N2427, N2423, N2231, N2349);
xor XOR2 (N2428, N2421, N47);
and AND2 (N2429, N2425, N771);
buf BUF1 (N2430, N2419);
nor NOR2 (N2431, N2416, N2240);
or OR2 (N2432, N2430, N1658);
not NOT1 (N2433, N2431);
nor NOR3 (N2434, N2432, N1409, N235);
nor NOR2 (N2435, N2427, N1930);
not NOT1 (N2436, N2429);
and AND2 (N2437, N2436, N552);
not NOT1 (N2438, N2435);
xor XOR2 (N2439, N2438, N2346);
nand NAND4 (N2440, N2410, N1280, N581, N836);
xor XOR2 (N2441, N2412, N195);
nor NOR2 (N2442, N2434, N1258);
nor NOR3 (N2443, N2437, N388, N44);
nand NAND4 (N2444, N2426, N661, N1551, N294);
and AND4 (N2445, N2411, N2336, N1899, N1274);
not NOT1 (N2446, N2444);
not NOT1 (N2447, N2439);
and AND2 (N2448, N2447, N1348);
xor XOR2 (N2449, N2398, N2435);
nor NOR4 (N2450, N2445, N1593, N1186, N1267);
not NOT1 (N2451, N2428);
or OR4 (N2452, N2441, N1504, N2065, N387);
and AND2 (N2453, N2450, N1745);
buf BUF1 (N2454, N2452);
nand NAND2 (N2455, N2433, N724);
nor NOR2 (N2456, N2446, N1638);
and AND3 (N2457, N2440, N594, N428);
and AND3 (N2458, N2442, N1301, N880);
not NOT1 (N2459, N2451);
or OR2 (N2460, N2458, N1318);
or OR3 (N2461, N2449, N772, N1174);
nand NAND2 (N2462, N2461, N218);
buf BUF1 (N2463, N2455);
xor XOR2 (N2464, N2454, N1426);
xor XOR2 (N2465, N2464, N1943);
nand NAND3 (N2466, N2463, N2321, N1488);
not NOT1 (N2467, N2448);
nand NAND3 (N2468, N2462, N1252, N312);
nand NAND4 (N2469, N2468, N451, N226, N1933);
xor XOR2 (N2470, N2467, N877);
not NOT1 (N2471, N2460);
xor XOR2 (N2472, N2459, N1751);
buf BUF1 (N2473, N2453);
and AND4 (N2474, N2472, N1694, N852, N1511);
and AND2 (N2475, N2471, N481);
or OR4 (N2476, N2473, N1768, N407, N737);
nor NOR3 (N2477, N2443, N2368, N1021);
and AND3 (N2478, N2474, N1365, N1321);
nand NAND4 (N2479, N2478, N890, N557, N898);
buf BUF1 (N2480, N2466);
xor XOR2 (N2481, N2456, N342);
xor XOR2 (N2482, N2465, N418);
and AND4 (N2483, N2479, N1012, N1493, N1558);
nor NOR2 (N2484, N2483, N1916);
not NOT1 (N2485, N2469);
or OR3 (N2486, N2480, N442, N255);
buf BUF1 (N2487, N2457);
xor XOR2 (N2488, N2487, N1690);
or OR3 (N2489, N2475, N985, N172);
buf BUF1 (N2490, N2470);
buf BUF1 (N2491, N2489);
or OR3 (N2492, N2477, N1935, N410);
xor XOR2 (N2493, N2486, N413);
xor XOR2 (N2494, N2488, N104);
xor XOR2 (N2495, N2484, N1569);
buf BUF1 (N2496, N2491);
not NOT1 (N2497, N2476);
xor XOR2 (N2498, N2493, N1307);
buf BUF1 (N2499, N2481);
not NOT1 (N2500, N2496);
nand NAND4 (N2501, N2494, N338, N1170, N1273);
not NOT1 (N2502, N2500);
and AND3 (N2503, N2499, N847, N1175);
not NOT1 (N2504, N2502);
or OR4 (N2505, N2504, N1169, N1163, N824);
and AND2 (N2506, N2505, N2423);
or OR4 (N2507, N2490, N2250, N2389, N301);
xor XOR2 (N2508, N2497, N1631);
nor NOR4 (N2509, N2501, N203, N946, N1882);
or OR3 (N2510, N2507, N566, N2113);
not NOT1 (N2511, N2482);
buf BUF1 (N2512, N2506);
nand NAND3 (N2513, N2508, N517, N1058);
nand NAND4 (N2514, N2510, N96, N779, N1794);
nor NOR4 (N2515, N2498, N1839, N356, N1144);
nor NOR3 (N2516, N2503, N576, N17);
and AND3 (N2517, N2514, N1435, N1416);
and AND4 (N2518, N2517, N2271, N612, N1899);
or OR3 (N2519, N2513, N1093, N2265);
nor NOR2 (N2520, N2492, N1755);
and AND4 (N2521, N2520, N1304, N701, N1752);
nor NOR4 (N2522, N2516, N1132, N1727, N1913);
not NOT1 (N2523, N2519);
not NOT1 (N2524, N2522);
buf BUF1 (N2525, N2518);
xor XOR2 (N2526, N2511, N2114);
and AND2 (N2527, N2512, N860);
nand NAND3 (N2528, N2525, N2259, N21);
not NOT1 (N2529, N2526);
or OR4 (N2530, N2485, N1674, N772, N1638);
not NOT1 (N2531, N2515);
xor XOR2 (N2532, N2524, N2330);
or OR4 (N2533, N2521, N2042, N601, N894);
and AND3 (N2534, N2527, N1860, N345);
xor XOR2 (N2535, N2530, N2066);
buf BUF1 (N2536, N2535);
xor XOR2 (N2537, N2536, N1566);
and AND4 (N2538, N2528, N143, N1910, N561);
buf BUF1 (N2539, N2532);
not NOT1 (N2540, N2533);
nand NAND4 (N2541, N2538, N2464, N1094, N909);
or OR2 (N2542, N2495, N43);
and AND4 (N2543, N2539, N1384, N172, N2326);
and AND3 (N2544, N2543, N206, N57);
nand NAND2 (N2545, N2540, N195);
nand NAND2 (N2546, N2509, N1568);
nand NAND3 (N2547, N2542, N395, N385);
nand NAND3 (N2548, N2546, N1515, N1256);
and AND4 (N2549, N2534, N1125, N384, N2294);
or OR3 (N2550, N2544, N1139, N577);
nand NAND3 (N2551, N2545, N117, N56);
and AND2 (N2552, N2547, N967);
and AND3 (N2553, N2552, N617, N1061);
buf BUF1 (N2554, N2523);
xor XOR2 (N2555, N2550, N1974);
nor NOR3 (N2556, N2531, N1787, N2352);
and AND3 (N2557, N2554, N1276, N1687);
xor XOR2 (N2558, N2541, N2258);
buf BUF1 (N2559, N2549);
nor NOR2 (N2560, N2559, N1559);
buf BUF1 (N2561, N2560);
and AND3 (N2562, N2529, N2348, N2360);
and AND3 (N2563, N2553, N578, N382);
and AND4 (N2564, N2558, N963, N874, N1982);
nor NOR2 (N2565, N2551, N790);
buf BUF1 (N2566, N2557);
not NOT1 (N2567, N2537);
not NOT1 (N2568, N2562);
and AND2 (N2569, N2561, N1151);
xor XOR2 (N2570, N2556, N983);
and AND3 (N2571, N2566, N2165, N2274);
buf BUF1 (N2572, N2548);
and AND2 (N2573, N2564, N389);
nor NOR2 (N2574, N2567, N2123);
nor NOR3 (N2575, N2570, N1602, N1656);
not NOT1 (N2576, N2565);
nand NAND3 (N2577, N2569, N1271, N1956);
not NOT1 (N2578, N2563);
xor XOR2 (N2579, N2571, N2287);
or OR2 (N2580, N2568, N1112);
and AND4 (N2581, N2577, N1295, N943, N2107);
or OR4 (N2582, N2580, N2202, N1136, N74);
or OR2 (N2583, N2579, N418);
buf BUF1 (N2584, N2574);
or OR4 (N2585, N2578, N1129, N2004, N1584);
nor NOR3 (N2586, N2582, N2211, N260);
nand NAND4 (N2587, N2586, N239, N1785, N1962);
not NOT1 (N2588, N2587);
buf BUF1 (N2589, N2584);
and AND3 (N2590, N2575, N1732, N2162);
or OR2 (N2591, N2581, N222);
or OR2 (N2592, N2590, N2170);
buf BUF1 (N2593, N2573);
or OR3 (N2594, N2576, N90, N417);
not NOT1 (N2595, N2583);
nor NOR4 (N2596, N2589, N1537, N160, N2249);
nor NOR3 (N2597, N2588, N1653, N1442);
not NOT1 (N2598, N2585);
nor NOR4 (N2599, N2596, N51, N340, N57);
nand NAND4 (N2600, N2597, N306, N1980, N1117);
and AND2 (N2601, N2593, N2149);
nand NAND3 (N2602, N2601, N1444, N489);
nand NAND2 (N2603, N2595, N363);
and AND4 (N2604, N2592, N750, N703, N927);
and AND3 (N2605, N2604, N2377, N189);
buf BUF1 (N2606, N2600);
and AND4 (N2607, N2605, N1666, N384, N619);
and AND2 (N2608, N2603, N1643);
xor XOR2 (N2609, N2591, N1007);
or OR2 (N2610, N2602, N141);
nand NAND2 (N2611, N2555, N2214);
not NOT1 (N2612, N2572);
nand NAND2 (N2613, N2610, N1636);
nand NAND3 (N2614, N2606, N751, N555);
nand NAND3 (N2615, N2611, N1135, N387);
nand NAND3 (N2616, N2598, N2116, N831);
nand NAND3 (N2617, N2616, N1936, N427);
buf BUF1 (N2618, N2594);
not NOT1 (N2619, N2617);
not NOT1 (N2620, N2618);
nor NOR2 (N2621, N2615, N1541);
buf BUF1 (N2622, N2614);
xor XOR2 (N2623, N2609, N2345);
nand NAND3 (N2624, N2623, N69, N1770);
buf BUF1 (N2625, N2622);
not NOT1 (N2626, N2621);
xor XOR2 (N2627, N2608, N291);
buf BUF1 (N2628, N2599);
not NOT1 (N2629, N2619);
buf BUF1 (N2630, N2607);
not NOT1 (N2631, N2626);
nand NAND4 (N2632, N2627, N571, N175, N391);
nor NOR4 (N2633, N2630, N644, N1624, N1949);
nand NAND4 (N2634, N2620, N1511, N871, N1083);
xor XOR2 (N2635, N2634, N2071);
nor NOR4 (N2636, N2624, N544, N1011, N643);
nor NOR4 (N2637, N2628, N1995, N555, N2143);
nor NOR4 (N2638, N2631, N1197, N2240, N1304);
buf BUF1 (N2639, N2613);
xor XOR2 (N2640, N2625, N2126);
and AND4 (N2641, N2633, N1665, N1677, N755);
and AND4 (N2642, N2638, N483, N548, N190);
buf BUF1 (N2643, N2635);
and AND2 (N2644, N2632, N2012);
and AND2 (N2645, N2629, N2471);
or OR3 (N2646, N2645, N871, N677);
and AND4 (N2647, N2641, N705, N2304, N1296);
buf BUF1 (N2648, N2640);
xor XOR2 (N2649, N2639, N793);
xor XOR2 (N2650, N2644, N681);
xor XOR2 (N2651, N2643, N634);
xor XOR2 (N2652, N2646, N2207);
nor NOR4 (N2653, N2650, N1532, N722, N1561);
buf BUF1 (N2654, N2647);
nor NOR2 (N2655, N2653, N247);
nor NOR3 (N2656, N2612, N2557, N307);
and AND4 (N2657, N2656, N2138, N1368, N1031);
nand NAND3 (N2658, N2657, N159, N2121);
or OR2 (N2659, N2648, N686);
and AND4 (N2660, N2637, N2456, N413, N1268);
or OR4 (N2661, N2636, N292, N915, N802);
buf BUF1 (N2662, N2659);
or OR3 (N2663, N2652, N1799, N2468);
xor XOR2 (N2664, N2642, N1553);
nor NOR4 (N2665, N2660, N150, N62, N647);
xor XOR2 (N2666, N2662, N2636);
nand NAND4 (N2667, N2661, N1921, N1649, N1323);
or OR4 (N2668, N2665, N2379, N9, N2587);
nand NAND4 (N2669, N2668, N1695, N1562, N762);
nor NOR3 (N2670, N2669, N177, N1963);
buf BUF1 (N2671, N2655);
and AND3 (N2672, N2664, N2374, N2520);
and AND3 (N2673, N2663, N1331, N848);
nor NOR4 (N2674, N2649, N59, N1439, N1986);
or OR3 (N2675, N2658, N2526, N234);
and AND3 (N2676, N2667, N819, N404);
nor NOR3 (N2677, N2672, N1200, N2636);
or OR3 (N2678, N2677, N1838, N1349);
nand NAND2 (N2679, N2671, N983);
buf BUF1 (N2680, N2654);
nor NOR2 (N2681, N2680, N1240);
nor NOR2 (N2682, N2678, N2354);
nand NAND3 (N2683, N2674, N702, N1218);
not NOT1 (N2684, N2666);
nand NAND3 (N2685, N2684, N1304, N2150);
nor NOR4 (N2686, N2679, N213, N911, N1007);
buf BUF1 (N2687, N2673);
xor XOR2 (N2688, N2681, N2437);
nand NAND3 (N2689, N2675, N382, N457);
and AND4 (N2690, N2682, N1481, N2307, N1864);
nand NAND2 (N2691, N2687, N646);
and AND3 (N2692, N2688, N2366, N1039);
or OR2 (N2693, N2689, N628);
nand NAND3 (N2694, N2686, N146, N1761);
not NOT1 (N2695, N2651);
xor XOR2 (N2696, N2695, N1992);
and AND3 (N2697, N2670, N2179, N1954);
xor XOR2 (N2698, N2696, N770);
not NOT1 (N2699, N2698);
nand NAND2 (N2700, N2691, N1820);
not NOT1 (N2701, N2685);
and AND2 (N2702, N2701, N2124);
or OR3 (N2703, N2683, N1935, N144);
or OR2 (N2704, N2700, N274);
buf BUF1 (N2705, N2693);
nor NOR3 (N2706, N2694, N1048, N381);
xor XOR2 (N2707, N2706, N1517);
nand NAND4 (N2708, N2692, N1754, N397, N1758);
buf BUF1 (N2709, N2707);
and AND2 (N2710, N2697, N955);
nor NOR4 (N2711, N2676, N2496, N529, N447);
xor XOR2 (N2712, N2704, N2708);
nand NAND3 (N2713, N2080, N2299, N1014);
xor XOR2 (N2714, N2711, N1602);
nand NAND3 (N2715, N2699, N1184, N1741);
and AND2 (N2716, N2703, N1439);
and AND2 (N2717, N2716, N36);
nor NOR3 (N2718, N2710, N2693, N2270);
and AND2 (N2719, N2718, N129);
xor XOR2 (N2720, N2713, N782);
buf BUF1 (N2721, N2720);
and AND2 (N2722, N2714, N1243);
xor XOR2 (N2723, N2722, N953);
and AND2 (N2724, N2709, N2504);
nand NAND3 (N2725, N2717, N1040, N2623);
nor NOR3 (N2726, N2702, N1374, N901);
buf BUF1 (N2727, N2726);
or OR3 (N2728, N2705, N2573, N784);
nand NAND2 (N2729, N2719, N196);
and AND4 (N2730, N2723, N1113, N2603, N375);
not NOT1 (N2731, N2730);
nand NAND4 (N2732, N2715, N745, N1581, N543);
not NOT1 (N2733, N2725);
or OR2 (N2734, N2724, N2653);
nand NAND4 (N2735, N2690, N889, N1446, N1363);
nor NOR4 (N2736, N2721, N2321, N474, N1407);
xor XOR2 (N2737, N2712, N1531);
or OR4 (N2738, N2729, N547, N1966, N1485);
not NOT1 (N2739, N2733);
or OR3 (N2740, N2735, N1611, N2144);
or OR2 (N2741, N2734, N1465);
xor XOR2 (N2742, N2732, N2410);
and AND3 (N2743, N2739, N1652, N158);
or OR4 (N2744, N2740, N2423, N1158, N647);
or OR3 (N2745, N2738, N344, N2355);
buf BUF1 (N2746, N2741);
and AND2 (N2747, N2737, N859);
and AND2 (N2748, N2742, N1218);
or OR2 (N2749, N2727, N2028);
xor XOR2 (N2750, N2744, N2125);
not NOT1 (N2751, N2745);
xor XOR2 (N2752, N2751, N1294);
or OR4 (N2753, N2743, N1462, N2580, N2703);
xor XOR2 (N2754, N2747, N186);
xor XOR2 (N2755, N2753, N776);
nand NAND4 (N2756, N2731, N2059, N1164, N2272);
not NOT1 (N2757, N2748);
xor XOR2 (N2758, N2750, N184);
buf BUF1 (N2759, N2755);
nor NOR3 (N2760, N2758, N2092, N1162);
xor XOR2 (N2761, N2736, N47);
or OR3 (N2762, N2757, N2148, N1477);
not NOT1 (N2763, N2759);
or OR4 (N2764, N2752, N1230, N169, N655);
nand NAND4 (N2765, N2749, N1771, N1112, N2091);
xor XOR2 (N2766, N2746, N1335);
xor XOR2 (N2767, N2766, N1066);
buf BUF1 (N2768, N2765);
nor NOR4 (N2769, N2756, N646, N2124, N724);
buf BUF1 (N2770, N2769);
buf BUF1 (N2771, N2764);
not NOT1 (N2772, N2760);
or OR3 (N2773, N2771, N262, N2710);
or OR2 (N2774, N2763, N1608);
xor XOR2 (N2775, N2772, N612);
buf BUF1 (N2776, N2768);
not NOT1 (N2777, N2775);
not NOT1 (N2778, N2776);
and AND3 (N2779, N2767, N1223, N1506);
or OR2 (N2780, N2773, N2669);
nand NAND4 (N2781, N2774, N1342, N1176, N159);
nand NAND2 (N2782, N2728, N657);
nand NAND3 (N2783, N2779, N2182, N194);
or OR3 (N2784, N2778, N288, N158);
nand NAND4 (N2785, N2761, N1090, N2113, N1759);
xor XOR2 (N2786, N2762, N249);
nor NOR3 (N2787, N2785, N2175, N2215);
or OR2 (N2788, N2770, N2215);
buf BUF1 (N2789, N2787);
not NOT1 (N2790, N2754);
buf BUF1 (N2791, N2789);
xor XOR2 (N2792, N2788, N327);
nor NOR3 (N2793, N2783, N230, N699);
and AND2 (N2794, N2777, N1592);
and AND4 (N2795, N2786, N2436, N1236, N1303);
not NOT1 (N2796, N2780);
buf BUF1 (N2797, N2794);
nor NOR3 (N2798, N2793, N1269, N701);
buf BUF1 (N2799, N2782);
xor XOR2 (N2800, N2799, N1366);
xor XOR2 (N2801, N2791, N19);
or OR4 (N2802, N2781, N953, N2491, N2222);
or OR4 (N2803, N2801, N2133, N2631, N2721);
nor NOR3 (N2804, N2795, N20, N388);
buf BUF1 (N2805, N2798);
nor NOR4 (N2806, N2805, N2610, N207, N676);
not NOT1 (N2807, N2784);
buf BUF1 (N2808, N2797);
nand NAND4 (N2809, N2790, N327, N1626, N2045);
nor NOR2 (N2810, N2808, N157);
nand NAND2 (N2811, N2803, N2347);
nor NOR3 (N2812, N2802, N387, N2668);
or OR4 (N2813, N2812, N757, N50, N1304);
and AND2 (N2814, N2811, N1000);
nand NAND3 (N2815, N2814, N2482, N1108);
or OR2 (N2816, N2813, N594);
nand NAND2 (N2817, N2809, N1747);
and AND4 (N2818, N2815, N823, N2574, N692);
nand NAND4 (N2819, N2816, N2587, N2589, N166);
buf BUF1 (N2820, N2796);
or OR2 (N2821, N2792, N2340);
buf BUF1 (N2822, N2807);
or OR3 (N2823, N2804, N2034, N1984);
not NOT1 (N2824, N2817);
buf BUF1 (N2825, N2819);
nor NOR3 (N2826, N2825, N1239, N50);
and AND2 (N2827, N2823, N636);
xor XOR2 (N2828, N2800, N1823);
and AND2 (N2829, N2827, N2824);
or OR2 (N2830, N975, N2028);
or OR3 (N2831, N2820, N1064, N1793);
xor XOR2 (N2832, N2830, N690);
or OR2 (N2833, N2821, N2176);
nor NOR2 (N2834, N2829, N1348);
buf BUF1 (N2835, N2834);
nand NAND4 (N2836, N2826, N2431, N2471, N694);
buf BUF1 (N2837, N2818);
nand NAND2 (N2838, N2822, N2308);
buf BUF1 (N2839, N2836);
or OR2 (N2840, N2828, N1113);
nor NOR4 (N2841, N2840, N1085, N2056, N185);
buf BUF1 (N2842, N2833);
nand NAND4 (N2843, N2832, N2662, N2135, N2708);
not NOT1 (N2844, N2810);
and AND3 (N2845, N2841, N876, N813);
and AND2 (N2846, N2839, N797);
not NOT1 (N2847, N2806);
or OR4 (N2848, N2845, N103, N2280, N295);
and AND4 (N2849, N2838, N1159, N2106, N2270);
nand NAND3 (N2850, N2831, N919, N285);
nand NAND3 (N2851, N2850, N1943, N2701);
and AND2 (N2852, N2844, N820);
xor XOR2 (N2853, N2849, N1305);
buf BUF1 (N2854, N2837);
nor NOR3 (N2855, N2842, N2792, N2130);
not NOT1 (N2856, N2843);
buf BUF1 (N2857, N2846);
not NOT1 (N2858, N2855);
xor XOR2 (N2859, N2851, N1429);
nor NOR2 (N2860, N2852, N2788);
not NOT1 (N2861, N2857);
and AND2 (N2862, N2853, N2168);
or OR2 (N2863, N2861, N1356);
nor NOR4 (N2864, N2856, N1483, N2107, N699);
xor XOR2 (N2865, N2862, N1816);
not NOT1 (N2866, N2864);
or OR2 (N2867, N2835, N1291);
or OR2 (N2868, N2865, N1915);
not NOT1 (N2869, N2866);
nand NAND2 (N2870, N2858, N1505);
buf BUF1 (N2871, N2867);
not NOT1 (N2872, N2871);
buf BUF1 (N2873, N2847);
not NOT1 (N2874, N2860);
nand NAND4 (N2875, N2863, N1738, N786, N2780);
nand NAND4 (N2876, N2875, N2188, N1567, N936);
buf BUF1 (N2877, N2874);
or OR2 (N2878, N2873, N1621);
nor NOR3 (N2879, N2868, N2861, N1277);
not NOT1 (N2880, N2879);
and AND4 (N2881, N2870, N1850, N71, N840);
not NOT1 (N2882, N2878);
and AND4 (N2883, N2877, N1549, N2313, N2127);
nor NOR2 (N2884, N2859, N1995);
nand NAND4 (N2885, N2876, N857, N1544, N2642);
buf BUF1 (N2886, N2848);
buf BUF1 (N2887, N2872);
xor XOR2 (N2888, N2880, N240);
and AND3 (N2889, N2885, N1052, N254);
or OR4 (N2890, N2889, N1860, N355, N2485);
buf BUF1 (N2891, N2886);
or OR3 (N2892, N2890, N2001, N2239);
not NOT1 (N2893, N2854);
nor NOR2 (N2894, N2882, N2373);
nand NAND4 (N2895, N2883, N1605, N1329, N970);
or OR3 (N2896, N2892, N393, N1011);
nor NOR2 (N2897, N2895, N1634);
or OR2 (N2898, N2869, N2474);
and AND3 (N2899, N2893, N248, N438);
nor NOR3 (N2900, N2899, N1089, N1496);
and AND3 (N2901, N2884, N1450, N1409);
nand NAND3 (N2902, N2891, N1786, N1151);
and AND2 (N2903, N2894, N2266);
buf BUF1 (N2904, N2902);
nor NOR3 (N2905, N2897, N2404, N1172);
buf BUF1 (N2906, N2901);
buf BUF1 (N2907, N2881);
or OR4 (N2908, N2887, N405, N284, N549);
nand NAND2 (N2909, N2898, N312);
nand NAND3 (N2910, N2909, N2824, N319);
and AND2 (N2911, N2908, N1134);
or OR4 (N2912, N2904, N1911, N1438, N2035);
nand NAND2 (N2913, N2900, N1410);
nand NAND4 (N2914, N2907, N2585, N1885, N2225);
xor XOR2 (N2915, N2913, N1533);
xor XOR2 (N2916, N2906, N2423);
buf BUF1 (N2917, N2914);
xor XOR2 (N2918, N2917, N2509);
and AND3 (N2919, N2912, N2105, N608);
nor NOR4 (N2920, N2918, N908, N430, N2316);
not NOT1 (N2921, N2888);
xor XOR2 (N2922, N2919, N1668);
buf BUF1 (N2923, N2905);
nand NAND3 (N2924, N2916, N302, N376);
nand NAND4 (N2925, N2911, N1023, N2563, N545);
buf BUF1 (N2926, N2921);
nand NAND3 (N2927, N2923, N1351, N1666);
or OR4 (N2928, N2903, N851, N1286, N1504);
nand NAND4 (N2929, N2915, N1951, N2602, N1621);
nand NAND2 (N2930, N2926, N1201);
not NOT1 (N2931, N2929);
and AND2 (N2932, N2928, N167);
nand NAND2 (N2933, N2925, N1649);
nand NAND3 (N2934, N2931, N2605, N2237);
nor NOR3 (N2935, N2922, N421, N1705);
not NOT1 (N2936, N2910);
or OR3 (N2937, N2930, N2320, N1025);
nor NOR4 (N2938, N2927, N1726, N2607, N1963);
and AND2 (N2939, N2938, N633);
not NOT1 (N2940, N2935);
nor NOR2 (N2941, N2934, N1879);
not NOT1 (N2942, N2937);
nor NOR4 (N2943, N2942, N920, N2448, N962);
xor XOR2 (N2944, N2943, N431);
buf BUF1 (N2945, N2896);
xor XOR2 (N2946, N2941, N2856);
or OR3 (N2947, N2939, N2661, N512);
and AND3 (N2948, N2924, N1716, N658);
not NOT1 (N2949, N2945);
and AND4 (N2950, N2948, N2314, N1625, N320);
buf BUF1 (N2951, N2944);
buf BUF1 (N2952, N2946);
or OR3 (N2953, N2940, N2472, N2470);
or OR2 (N2954, N2952, N2210);
and AND3 (N2955, N2950, N2322, N2537);
xor XOR2 (N2956, N2933, N276);
nor NOR4 (N2957, N2932, N1986, N43, N2788);
and AND4 (N2958, N2956, N177, N409, N2386);
buf BUF1 (N2959, N2949);
or OR2 (N2960, N2954, N2128);
and AND4 (N2961, N2958, N2011, N1037, N1590);
and AND3 (N2962, N2957, N1420, N138);
nor NOR4 (N2963, N2960, N1793, N1052, N1671);
buf BUF1 (N2964, N2953);
nand NAND3 (N2965, N2962, N1154, N633);
or OR2 (N2966, N2963, N1120);
or OR4 (N2967, N2961, N2748, N1995, N1894);
xor XOR2 (N2968, N2965, N1011);
nor NOR2 (N2969, N2959, N860);
not NOT1 (N2970, N2951);
nand NAND4 (N2971, N2947, N645, N928, N493);
not NOT1 (N2972, N2920);
nor NOR2 (N2973, N2969, N959);
or OR2 (N2974, N2972, N1650);
buf BUF1 (N2975, N2971);
buf BUF1 (N2976, N2974);
buf BUF1 (N2977, N2976);
or OR4 (N2978, N2936, N918, N171, N854);
xor XOR2 (N2979, N2978, N2141);
xor XOR2 (N2980, N2970, N715);
buf BUF1 (N2981, N2967);
xor XOR2 (N2982, N2981, N2478);
nand NAND2 (N2983, N2966, N510);
xor XOR2 (N2984, N2968, N2764);
nor NOR4 (N2985, N2982, N102, N997, N1793);
buf BUF1 (N2986, N2984);
buf BUF1 (N2987, N2964);
buf BUF1 (N2988, N2979);
and AND2 (N2989, N2975, N1313);
not NOT1 (N2990, N2985);
xor XOR2 (N2991, N2955, N1120);
and AND2 (N2992, N2990, N491);
or OR4 (N2993, N2977, N710, N2116, N2757);
buf BUF1 (N2994, N2986);
not NOT1 (N2995, N2993);
or OR2 (N2996, N2983, N632);
xor XOR2 (N2997, N2996, N1075);
not NOT1 (N2998, N2987);
nor NOR3 (N2999, N2997, N2128, N944);
buf BUF1 (N3000, N2989);
and AND3 (N3001, N2999, N1145, N1995);
xor XOR2 (N3002, N3000, N968);
buf BUF1 (N3003, N3001);
buf BUF1 (N3004, N2991);
buf BUF1 (N3005, N3003);
not NOT1 (N3006, N3002);
nand NAND3 (N3007, N2995, N2958, N1271);
buf BUF1 (N3008, N2994);
and AND3 (N3009, N2973, N1609, N1089);
nor NOR2 (N3010, N3005, N672);
xor XOR2 (N3011, N2988, N787);
not NOT1 (N3012, N3006);
buf BUF1 (N3013, N3012);
xor XOR2 (N3014, N3013, N1737);
and AND3 (N3015, N3008, N1289, N2645);
or OR2 (N3016, N2980, N2352);
buf BUF1 (N3017, N3010);
xor XOR2 (N3018, N3007, N352);
and AND3 (N3019, N3004, N477, N1512);
and AND3 (N3020, N2992, N1521, N1765);
buf BUF1 (N3021, N2998);
xor XOR2 (N3022, N3018, N1208);
or OR4 (N3023, N3016, N337, N2383, N2295);
nand NAND4 (N3024, N3017, N2421, N1838, N2823);
buf BUF1 (N3025, N3021);
buf BUF1 (N3026, N3023);
or OR3 (N3027, N3009, N596, N2272);
and AND3 (N3028, N3020, N1173, N980);
or OR2 (N3029, N3019, N1171);
and AND3 (N3030, N3026, N1289, N440);
buf BUF1 (N3031, N3014);
not NOT1 (N3032, N3024);
nand NAND2 (N3033, N3015, N2878);
nand NAND4 (N3034, N3029, N195, N2442, N2114);
or OR3 (N3035, N3032, N1414, N1759);
or OR2 (N3036, N3027, N2879);
or OR4 (N3037, N3035, N2786, N1387, N421);
buf BUF1 (N3038, N3034);
not NOT1 (N3039, N3037);
and AND3 (N3040, N3011, N1307, N2219);
not NOT1 (N3041, N3028);
xor XOR2 (N3042, N3025, N1482);
buf BUF1 (N3043, N3039);
nand NAND3 (N3044, N3022, N2539, N518);
not NOT1 (N3045, N3043);
or OR4 (N3046, N3042, N376, N2115, N2017);
xor XOR2 (N3047, N3044, N532);
xor XOR2 (N3048, N3033, N1257);
buf BUF1 (N3049, N3038);
nand NAND4 (N3050, N3045, N758, N2500, N195);
and AND3 (N3051, N3031, N1221, N2995);
buf BUF1 (N3052, N3030);
or OR2 (N3053, N3049, N2158);
buf BUF1 (N3054, N3051);
nand NAND2 (N3055, N3040, N475);
nand NAND4 (N3056, N3036, N826, N994, N2581);
buf BUF1 (N3057, N3052);
xor XOR2 (N3058, N3047, N372);
buf BUF1 (N3059, N3055);
nand NAND2 (N3060, N3046, N863);
not NOT1 (N3061, N3041);
buf BUF1 (N3062, N3060);
or OR3 (N3063, N3048, N1360, N429);
and AND3 (N3064, N3058, N954, N469);
buf BUF1 (N3065, N3063);
not NOT1 (N3066, N3065);
not NOT1 (N3067, N3056);
or OR2 (N3068, N3066, N2025);
buf BUF1 (N3069, N3053);
buf BUF1 (N3070, N3064);
or OR4 (N3071, N3068, N1206, N1496, N1871);
nand NAND2 (N3072, N3071, N2845);
nor NOR2 (N3073, N3061, N906);
nor NOR2 (N3074, N3057, N862);
buf BUF1 (N3075, N3059);
nor NOR4 (N3076, N3074, N2046, N931, N294);
not NOT1 (N3077, N3075);
not NOT1 (N3078, N3072);
nor NOR3 (N3079, N3073, N1355, N490);
xor XOR2 (N3080, N3067, N2500);
nor NOR3 (N3081, N3078, N1194, N2831);
not NOT1 (N3082, N3054);
buf BUF1 (N3083, N3080);
not NOT1 (N3084, N3076);
not NOT1 (N3085, N3050);
xor XOR2 (N3086, N3082, N557);
buf BUF1 (N3087, N3086);
xor XOR2 (N3088, N3062, N579);
nand NAND2 (N3089, N3069, N65);
and AND4 (N3090, N3070, N914, N1806, N249);
nand NAND4 (N3091, N3090, N1726, N898, N275);
nor NOR2 (N3092, N3087, N1410);
xor XOR2 (N3093, N3089, N556);
buf BUF1 (N3094, N3083);
buf BUF1 (N3095, N3092);
xor XOR2 (N3096, N3077, N674);
buf BUF1 (N3097, N3093);
and AND3 (N3098, N3096, N2912, N1771);
and AND3 (N3099, N3097, N1703, N1025);
or OR2 (N3100, N3095, N2959);
or OR3 (N3101, N3085, N2130, N1998);
and AND2 (N3102, N3100, N889);
nor NOR3 (N3103, N3099, N245, N1651);
and AND2 (N3104, N3101, N705);
xor XOR2 (N3105, N3102, N317);
or OR4 (N3106, N3103, N1396, N809, N1889);
nor NOR4 (N3107, N3098, N215, N2738, N1345);
buf BUF1 (N3108, N3084);
nand NAND4 (N3109, N3108, N2964, N494, N302);
nor NOR3 (N3110, N3104, N2874, N570);
not NOT1 (N3111, N3105);
xor XOR2 (N3112, N3088, N1135);
or OR3 (N3113, N3109, N626, N1002);
buf BUF1 (N3114, N3094);
and AND3 (N3115, N3091, N1015, N983);
xor XOR2 (N3116, N3115, N2583);
nand NAND2 (N3117, N3114, N1194);
nor NOR4 (N3118, N3117, N526, N1676, N2760);
or OR2 (N3119, N3110, N25);
xor XOR2 (N3120, N3079, N1176);
and AND4 (N3121, N3081, N2944, N2535, N185);
nor NOR3 (N3122, N3111, N567, N1913);
or OR4 (N3123, N3118, N2246, N2706, N2303);
nand NAND4 (N3124, N3106, N2549, N2980, N2746);
or OR4 (N3125, N3112, N176, N582, N1575);
nand NAND4 (N3126, N3123, N3055, N2868, N3097);
xor XOR2 (N3127, N3124, N2533);
or OR3 (N3128, N3119, N1477, N661);
nor NOR2 (N3129, N3113, N306);
buf BUF1 (N3130, N3126);
nor NOR3 (N3131, N3128, N1149, N828);
or OR3 (N3132, N3122, N1771, N2164);
or OR2 (N3133, N3129, N190);
nor NOR4 (N3134, N3132, N1849, N2584, N1050);
xor XOR2 (N3135, N3107, N22);
nor NOR2 (N3136, N3133, N99);
and AND3 (N3137, N3134, N1916, N2110);
xor XOR2 (N3138, N3137, N1038);
xor XOR2 (N3139, N3138, N2164);
xor XOR2 (N3140, N3127, N3022);
nor NOR3 (N3141, N3121, N1412, N308);
and AND4 (N3142, N3131, N2579, N1788, N1821);
nand NAND3 (N3143, N3136, N967, N2080);
and AND4 (N3144, N3120, N775, N2609, N551);
and AND4 (N3145, N3139, N2649, N2272, N492);
not NOT1 (N3146, N3130);
buf BUF1 (N3147, N3141);
nor NOR2 (N3148, N3145, N1815);
not NOT1 (N3149, N3125);
or OR4 (N3150, N3142, N80, N1323, N600);
xor XOR2 (N3151, N3147, N2016);
nor NOR3 (N3152, N3140, N164, N590);
and AND2 (N3153, N3149, N2835);
or OR4 (N3154, N3143, N37, N954, N2996);
and AND2 (N3155, N3153, N1655);
and AND4 (N3156, N3146, N1449, N265, N1773);
buf BUF1 (N3157, N3148);
or OR2 (N3158, N3150, N606);
nand NAND3 (N3159, N3116, N1871, N2425);
nor NOR4 (N3160, N3158, N2396, N2050, N1270);
or OR3 (N3161, N3160, N2613, N1266);
nand NAND2 (N3162, N3155, N1959);
xor XOR2 (N3163, N3156, N397);
nor NOR3 (N3164, N3144, N310, N153);
nand NAND3 (N3165, N3151, N1997, N1901);
buf BUF1 (N3166, N3152);
xor XOR2 (N3167, N3161, N2978);
nand NAND3 (N3168, N3166, N2292, N2563);
and AND2 (N3169, N3165, N2139);
nand NAND2 (N3170, N3167, N2177);
buf BUF1 (N3171, N3168);
buf BUF1 (N3172, N3154);
xor XOR2 (N3173, N3164, N407);
xor XOR2 (N3174, N3157, N2531);
nand NAND2 (N3175, N3135, N555);
xor XOR2 (N3176, N3169, N2683);
nor NOR2 (N3177, N3163, N114);
nor NOR3 (N3178, N3173, N1278, N1715);
nor NOR3 (N3179, N3174, N2141, N2009);
nor NOR2 (N3180, N3176, N3051);
or OR2 (N3181, N3179, N1373);
xor XOR2 (N3182, N3175, N1502);
nand NAND3 (N3183, N3162, N1468, N1203);
or OR2 (N3184, N3159, N702);
and AND3 (N3185, N3182, N628, N2097);
and AND2 (N3186, N3178, N1824);
not NOT1 (N3187, N3170);
buf BUF1 (N3188, N3186);
not NOT1 (N3189, N3177);
buf BUF1 (N3190, N3184);
nand NAND4 (N3191, N3188, N400, N1586, N58);
nand NAND4 (N3192, N3185, N2703, N937, N317);
xor XOR2 (N3193, N3190, N1634);
nor NOR4 (N3194, N3191, N552, N2052, N1989);
and AND2 (N3195, N3187, N204);
nor NOR3 (N3196, N3183, N1140, N2344);
nand NAND2 (N3197, N3181, N1861);
and AND2 (N3198, N3172, N1925);
nand NAND3 (N3199, N3196, N2214, N2517);
buf BUF1 (N3200, N3199);
nor NOR2 (N3201, N3171, N1489);
or OR4 (N3202, N3189, N2541, N2997, N1614);
and AND2 (N3203, N3201, N3174);
or OR3 (N3204, N3200, N2519, N1856);
nand NAND2 (N3205, N3192, N2902);
nand NAND4 (N3206, N3195, N372, N994, N458);
xor XOR2 (N3207, N3180, N213);
not NOT1 (N3208, N3204);
and AND3 (N3209, N3205, N1976, N1843);
or OR3 (N3210, N3206, N2880, N1621);
xor XOR2 (N3211, N3207, N87);
xor XOR2 (N3212, N3209, N3076);
xor XOR2 (N3213, N3208, N567);
or OR4 (N3214, N3211, N2284, N51, N1313);
nor NOR2 (N3215, N3214, N759);
or OR4 (N3216, N3213, N2760, N2075, N3117);
xor XOR2 (N3217, N3216, N1835);
nand NAND2 (N3218, N3197, N315);
buf BUF1 (N3219, N3215);
nor NOR3 (N3220, N3210, N2653, N2907);
nand NAND4 (N3221, N3212, N1597, N2697, N2915);
buf BUF1 (N3222, N3203);
xor XOR2 (N3223, N3220, N505);
and AND3 (N3224, N3218, N2436, N1937);
not NOT1 (N3225, N3193);
or OR3 (N3226, N3194, N2501, N2812);
and AND3 (N3227, N3198, N1840, N2083);
or OR4 (N3228, N3222, N652, N529, N25);
xor XOR2 (N3229, N3228, N2844);
and AND4 (N3230, N3217, N1039, N1456, N82);
buf BUF1 (N3231, N3226);
or OR2 (N3232, N3219, N3195);
not NOT1 (N3233, N3227);
nand NAND3 (N3234, N3231, N1357, N806);
or OR3 (N3235, N3225, N1567, N863);
not NOT1 (N3236, N3224);
nor NOR3 (N3237, N3229, N84, N2446);
nand NAND4 (N3238, N3233, N1293, N1684, N644);
not NOT1 (N3239, N3235);
and AND4 (N3240, N3238, N1259, N555, N3204);
xor XOR2 (N3241, N3232, N1258);
nor NOR2 (N3242, N3239, N1250);
xor XOR2 (N3243, N3221, N574);
nand NAND4 (N3244, N3242, N1629, N1604, N1158);
or OR2 (N3245, N3243, N2203);
xor XOR2 (N3246, N3234, N632);
not NOT1 (N3247, N3244);
nand NAND3 (N3248, N3247, N1946, N304);
buf BUF1 (N3249, N3237);
or OR4 (N3250, N3230, N3146, N3024, N1375);
or OR4 (N3251, N3248, N1184, N651, N1871);
buf BUF1 (N3252, N3250);
nor NOR2 (N3253, N3245, N3244);
nor NOR3 (N3254, N3249, N673, N506);
and AND2 (N3255, N3202, N2047);
nor NOR4 (N3256, N3255, N2107, N296, N1161);
buf BUF1 (N3257, N3253);
nor NOR4 (N3258, N3256, N1902, N1165, N999);
and AND3 (N3259, N3251, N2963, N3131);
nand NAND3 (N3260, N3252, N809, N1710);
or OR3 (N3261, N3260, N2906, N1196);
nand NAND3 (N3262, N3240, N1295, N37);
nand NAND4 (N3263, N3246, N1008, N2141, N717);
or OR3 (N3264, N3254, N2400, N2031);
buf BUF1 (N3265, N3236);
buf BUF1 (N3266, N3257);
or OR2 (N3267, N3259, N3115);
xor XOR2 (N3268, N3264, N2821);
nor NOR3 (N3269, N3241, N3156, N2728);
nor NOR2 (N3270, N3266, N1995);
buf BUF1 (N3271, N3258);
buf BUF1 (N3272, N3263);
not NOT1 (N3273, N3270);
not NOT1 (N3274, N3223);
xor XOR2 (N3275, N3268, N268);
buf BUF1 (N3276, N3272);
and AND2 (N3277, N3269, N3137);
nor NOR3 (N3278, N3275, N2135, N2428);
xor XOR2 (N3279, N3265, N1593);
or OR4 (N3280, N3271, N2070, N1278, N175);
nor NOR2 (N3281, N3278, N2842);
nor NOR2 (N3282, N3274, N1505);
buf BUF1 (N3283, N3276);
and AND2 (N3284, N3283, N2820);
not NOT1 (N3285, N3273);
or OR2 (N3286, N3262, N1688);
buf BUF1 (N3287, N3279);
and AND4 (N3288, N3277, N721, N748, N813);
and AND2 (N3289, N3286, N1462);
buf BUF1 (N3290, N3267);
not NOT1 (N3291, N3282);
buf BUF1 (N3292, N3289);
or OR2 (N3293, N3292, N84);
xor XOR2 (N3294, N3281, N370);
or OR3 (N3295, N3293, N745, N1737);
buf BUF1 (N3296, N3290);
nand NAND4 (N3297, N3284, N2732, N2083, N1091);
and AND2 (N3298, N3297, N630);
not NOT1 (N3299, N3295);
buf BUF1 (N3300, N3291);
and AND4 (N3301, N3294, N1141, N3001, N1753);
xor XOR2 (N3302, N3287, N1671);
and AND4 (N3303, N3261, N1036, N3171, N2961);
or OR2 (N3304, N3303, N181);
nor NOR4 (N3305, N3302, N189, N9, N132);
and AND4 (N3306, N3299, N2778, N1599, N482);
nand NAND2 (N3307, N3306, N639);
nand NAND2 (N3308, N3301, N362);
xor XOR2 (N3309, N3307, N2870);
or OR3 (N3310, N3305, N2306, N445);
nand NAND4 (N3311, N3298, N795, N1382, N759);
xor XOR2 (N3312, N3288, N2687);
or OR3 (N3313, N3280, N1129, N3059);
not NOT1 (N3314, N3310);
or OR4 (N3315, N3311, N454, N1451, N294);
nand NAND3 (N3316, N3308, N3107, N1070);
and AND4 (N3317, N3312, N608, N1400, N178);
or OR3 (N3318, N3304, N9, N2548);
not NOT1 (N3319, N3309);
or OR4 (N3320, N3315, N2597, N2906, N2011);
and AND3 (N3321, N3300, N2938, N453);
xor XOR2 (N3322, N3319, N3086);
nand NAND4 (N3323, N3317, N943, N1158, N2853);
buf BUF1 (N3324, N3316);
buf BUF1 (N3325, N3318);
xor XOR2 (N3326, N3323, N2523);
not NOT1 (N3327, N3322);
not NOT1 (N3328, N3314);
or OR3 (N3329, N3285, N2049, N2560);
or OR3 (N3330, N3320, N1468, N993);
nand NAND2 (N3331, N3296, N2439);
nand NAND3 (N3332, N3324, N2174, N3071);
not NOT1 (N3333, N3329);
not NOT1 (N3334, N3327);
buf BUF1 (N3335, N3330);
and AND2 (N3336, N3331, N169);
nor NOR2 (N3337, N3321, N699);
nand NAND3 (N3338, N3334, N2785, N1264);
xor XOR2 (N3339, N3325, N1543);
or OR3 (N3340, N3335, N1279, N1341);
not NOT1 (N3341, N3337);
or OR3 (N3342, N3341, N1487, N2753);
or OR3 (N3343, N3313, N3258, N1437);
nor NOR2 (N3344, N3336, N2170);
nand NAND3 (N3345, N3332, N1642, N391);
nor NOR2 (N3346, N3328, N2070);
buf BUF1 (N3347, N3339);
and AND2 (N3348, N3346, N1227);
xor XOR2 (N3349, N3347, N1589);
xor XOR2 (N3350, N3333, N3142);
and AND2 (N3351, N3350, N593);
nand NAND4 (N3352, N3340, N1684, N114, N3000);
nand NAND2 (N3353, N3352, N605);
buf BUF1 (N3354, N3342);
not NOT1 (N3355, N3343);
and AND3 (N3356, N3326, N2993, N209);
buf BUF1 (N3357, N3338);
buf BUF1 (N3358, N3344);
buf BUF1 (N3359, N3345);
and AND4 (N3360, N3351, N1161, N2625, N1370);
not NOT1 (N3361, N3357);
xor XOR2 (N3362, N3354, N988);
xor XOR2 (N3363, N3359, N2952);
nand NAND4 (N3364, N3362, N313, N601, N2646);
buf BUF1 (N3365, N3364);
buf BUF1 (N3366, N3358);
nand NAND2 (N3367, N3363, N1080);
not NOT1 (N3368, N3349);
not NOT1 (N3369, N3361);
and AND2 (N3370, N3348, N2324);
nand NAND3 (N3371, N3356, N2008, N2417);
buf BUF1 (N3372, N3353);
buf BUF1 (N3373, N3369);
nor NOR3 (N3374, N3372, N1127, N1167);
not NOT1 (N3375, N3370);
or OR4 (N3376, N3366, N2569, N3003, N685);
nor NOR3 (N3377, N3371, N1353, N3023);
and AND2 (N3378, N3355, N206);
not NOT1 (N3379, N3365);
nor NOR4 (N3380, N3375, N701, N2243, N1308);
nor NOR4 (N3381, N3367, N2155, N1876, N257);
xor XOR2 (N3382, N3368, N196);
buf BUF1 (N3383, N3373);
buf BUF1 (N3384, N3379);
buf BUF1 (N3385, N3383);
not NOT1 (N3386, N3374);
not NOT1 (N3387, N3385);
nor NOR4 (N3388, N3376, N2177, N2556, N1711);
xor XOR2 (N3389, N3384, N2588);
or OR2 (N3390, N3378, N1346);
xor XOR2 (N3391, N3386, N1588);
nor NOR4 (N3392, N3360, N600, N1472, N1913);
nor NOR2 (N3393, N3388, N924);
xor XOR2 (N3394, N3390, N2926);
xor XOR2 (N3395, N3391, N35);
nor NOR3 (N3396, N3394, N965, N3014);
nor NOR2 (N3397, N3380, N2066);
and AND4 (N3398, N3392, N1555, N371, N1589);
not NOT1 (N3399, N3393);
and AND2 (N3400, N3381, N2378);
and AND4 (N3401, N3399, N1260, N2717, N1574);
xor XOR2 (N3402, N3397, N1011);
nor NOR3 (N3403, N3389, N2805, N2052);
and AND2 (N3404, N3400, N1598);
or OR3 (N3405, N3387, N1084, N1587);
buf BUF1 (N3406, N3403);
nand NAND4 (N3407, N3402, N996, N624, N2267);
and AND4 (N3408, N3405, N1828, N2898, N693);
buf BUF1 (N3409, N3408);
and AND4 (N3410, N3382, N3244, N1816, N1040);
nand NAND4 (N3411, N3377, N563, N1168, N1808);
buf BUF1 (N3412, N3409);
not NOT1 (N3413, N3407);
nand NAND2 (N3414, N3401, N610);
nor NOR3 (N3415, N3395, N979, N1579);
and AND4 (N3416, N3406, N3079, N230, N3315);
buf BUF1 (N3417, N3396);
or OR2 (N3418, N3415, N2278);
or OR4 (N3419, N3411, N2503, N940, N1268);
and AND3 (N3420, N3410, N2101, N2200);
or OR4 (N3421, N3417, N1378, N3350, N1731);
nor NOR4 (N3422, N3420, N1410, N1055, N1976);
and AND2 (N3423, N3404, N344);
or OR2 (N3424, N3419, N1508);
nor NOR2 (N3425, N3398, N1501);
xor XOR2 (N3426, N3423, N2764);
nand NAND3 (N3427, N3416, N1505, N389);
nor NOR2 (N3428, N3425, N1091);
buf BUF1 (N3429, N3422);
and AND3 (N3430, N3413, N3214, N1483);
xor XOR2 (N3431, N3424, N3385);
not NOT1 (N3432, N3412);
buf BUF1 (N3433, N3430);
nor NOR2 (N3434, N3432, N2807);
or OR2 (N3435, N3426, N1618);
nand NAND3 (N3436, N3431, N536, N177);
and AND4 (N3437, N3435, N3059, N24, N2193);
not NOT1 (N3438, N3427);
xor XOR2 (N3439, N3436, N2738);
not NOT1 (N3440, N3429);
or OR3 (N3441, N3434, N1677, N2740);
not NOT1 (N3442, N3439);
buf BUF1 (N3443, N3418);
buf BUF1 (N3444, N3414);
not NOT1 (N3445, N3442);
xor XOR2 (N3446, N3433, N1770);
or OR4 (N3447, N3440, N235, N2515, N2782);
nor NOR4 (N3448, N3447, N14, N1572, N2204);
nand NAND4 (N3449, N3428, N2343, N3350, N540);
or OR4 (N3450, N3449, N1492, N2964, N2797);
nand NAND2 (N3451, N3441, N364);
not NOT1 (N3452, N3438);
buf BUF1 (N3453, N3437);
or OR4 (N3454, N3452, N3115, N827, N1395);
and AND4 (N3455, N3445, N1507, N2725, N2404);
or OR4 (N3456, N3444, N2741, N771, N2367);
buf BUF1 (N3457, N3451);
and AND4 (N3458, N3450, N121, N1046, N2442);
or OR4 (N3459, N3453, N2106, N2353, N299);
not NOT1 (N3460, N3458);
xor XOR2 (N3461, N3460, N2878);
nor NOR4 (N3462, N3455, N3330, N895, N673);
or OR4 (N3463, N3461, N785, N1125, N809);
and AND2 (N3464, N3462, N2800);
xor XOR2 (N3465, N3464, N991);
xor XOR2 (N3466, N3443, N207);
and AND2 (N3467, N3454, N1695);
and AND3 (N3468, N3465, N1924, N735);
xor XOR2 (N3469, N3466, N2963);
buf BUF1 (N3470, N3469);
nand NAND2 (N3471, N3468, N153);
xor XOR2 (N3472, N3421, N1178);
buf BUF1 (N3473, N3471);
xor XOR2 (N3474, N3463, N2070);
nand NAND4 (N3475, N3456, N1118, N2018, N2456);
nor NOR4 (N3476, N3459, N602, N623, N2541);
or OR3 (N3477, N3475, N2227, N94);
xor XOR2 (N3478, N3467, N3115);
nand NAND4 (N3479, N3474, N3255, N2387, N760);
or OR3 (N3480, N3476, N556, N112);
and AND4 (N3481, N3457, N2534, N3149, N1176);
xor XOR2 (N3482, N3470, N284);
buf BUF1 (N3483, N3482);
not NOT1 (N3484, N3483);
not NOT1 (N3485, N3448);
xor XOR2 (N3486, N3480, N173);
nor NOR3 (N3487, N3484, N2480, N51);
and AND3 (N3488, N3481, N247, N507);
buf BUF1 (N3489, N3486);
or OR2 (N3490, N3473, N2326);
not NOT1 (N3491, N3478);
nand NAND2 (N3492, N3485, N2496);
and AND3 (N3493, N3491, N1258, N1990);
or OR2 (N3494, N3488, N1699);
nand NAND4 (N3495, N3492, N3389, N2378, N1945);
not NOT1 (N3496, N3446);
buf BUF1 (N3497, N3496);
or OR3 (N3498, N3493, N1245, N1429);
not NOT1 (N3499, N3489);
nor NOR2 (N3500, N3472, N1571);
not NOT1 (N3501, N3479);
or OR3 (N3502, N3501, N714, N885);
xor XOR2 (N3503, N3500, N424);
nor NOR4 (N3504, N3487, N2647, N3076, N2464);
not NOT1 (N3505, N3499);
not NOT1 (N3506, N3505);
and AND2 (N3507, N3490, N81);
xor XOR2 (N3508, N3498, N3215);
not NOT1 (N3509, N3494);
xor XOR2 (N3510, N3495, N755);
nor NOR2 (N3511, N3503, N14);
or OR3 (N3512, N3509, N1413, N2816);
nand NAND2 (N3513, N3508, N2003);
buf BUF1 (N3514, N3502);
or OR2 (N3515, N3511, N1742);
nor NOR2 (N3516, N3477, N2530);
and AND4 (N3517, N3507, N1869, N3256, N1171);
xor XOR2 (N3518, N3514, N2389);
xor XOR2 (N3519, N3516, N3442);
and AND4 (N3520, N3515, N2518, N354, N1765);
not NOT1 (N3521, N3497);
xor XOR2 (N3522, N3512, N822);
nor NOR2 (N3523, N3504, N2191);
nand NAND3 (N3524, N3510, N2287, N772);
buf BUF1 (N3525, N3520);
or OR2 (N3526, N3517, N2295);
not NOT1 (N3527, N3506);
or OR3 (N3528, N3518, N650, N266);
nor NOR3 (N3529, N3519, N368, N1635);
xor XOR2 (N3530, N3523, N506);
and AND4 (N3531, N3528, N1271, N952, N1776);
or OR4 (N3532, N3526, N1087, N3098, N1510);
or OR3 (N3533, N3532, N3027, N2216);
buf BUF1 (N3534, N3529);
or OR2 (N3535, N3522, N1166);
nand NAND3 (N3536, N3527, N2217, N1817);
nor NOR4 (N3537, N3531, N1041, N2333, N3382);
nor NOR3 (N3538, N3536, N1647, N2241);
or OR3 (N3539, N3524, N663, N1517);
xor XOR2 (N3540, N3521, N517);
nor NOR4 (N3541, N3535, N3234, N385, N969);
nand NAND2 (N3542, N3537, N888);
nor NOR3 (N3543, N3541, N17, N953);
xor XOR2 (N3544, N3543, N39);
nand NAND2 (N3545, N3538, N425);
and AND2 (N3546, N3544, N1962);
nor NOR2 (N3547, N3545, N3004);
nor NOR3 (N3548, N3539, N735, N1499);
nand NAND4 (N3549, N3525, N2776, N2947, N3303);
xor XOR2 (N3550, N3549, N84);
buf BUF1 (N3551, N3542);
xor XOR2 (N3552, N3550, N3024);
not NOT1 (N3553, N3552);
nand NAND2 (N3554, N3546, N2444);
or OR2 (N3555, N3540, N1408);
and AND3 (N3556, N3551, N1562, N48);
not NOT1 (N3557, N3533);
buf BUF1 (N3558, N3534);
buf BUF1 (N3559, N3548);
xor XOR2 (N3560, N3555, N1990);
nand NAND2 (N3561, N3513, N3514);
or OR4 (N3562, N3554, N1106, N3502, N2191);
nand NAND4 (N3563, N3553, N3459, N2457, N1482);
not NOT1 (N3564, N3557);
buf BUF1 (N3565, N3547);
nand NAND4 (N3566, N3561, N205, N2697, N2897);
not NOT1 (N3567, N3530);
nor NOR2 (N3568, N3563, N2624);
nor NOR2 (N3569, N3564, N2354);
nand NAND3 (N3570, N3562, N1903, N1541);
or OR3 (N3571, N3567, N2262, N1223);
not NOT1 (N3572, N3565);
and AND4 (N3573, N3571, N1485, N2252, N2897);
nor NOR3 (N3574, N3560, N1755, N726);
nand NAND3 (N3575, N3558, N1128, N716);
not NOT1 (N3576, N3572);
not NOT1 (N3577, N3574);
nand NAND3 (N3578, N3575, N508, N1610);
nand NAND2 (N3579, N3578, N239);
and AND3 (N3580, N3568, N2792, N2630);
buf BUF1 (N3581, N3569);
and AND4 (N3582, N3556, N735, N275, N496);
buf BUF1 (N3583, N3580);
buf BUF1 (N3584, N3579);
and AND3 (N3585, N3559, N1431, N3326);
and AND2 (N3586, N3584, N2249);
not NOT1 (N3587, N3581);
nand NAND3 (N3588, N3577, N2985, N1552);
xor XOR2 (N3589, N3586, N2438);
or OR4 (N3590, N3588, N3207, N3138, N299);
xor XOR2 (N3591, N3590, N2941);
or OR3 (N3592, N3591, N605, N2062);
or OR4 (N3593, N3585, N1081, N2549, N1418);
buf BUF1 (N3594, N3592);
nor NOR2 (N3595, N3583, N990);
or OR3 (N3596, N3589, N1797, N1032);
nor NOR3 (N3597, N3570, N1759, N556);
xor XOR2 (N3598, N3573, N351);
nand NAND4 (N3599, N3596, N376, N2546, N2376);
nor NOR4 (N3600, N3576, N1943, N3152, N2879);
buf BUF1 (N3601, N3587);
nand NAND4 (N3602, N3595, N442, N2230, N3043);
xor XOR2 (N3603, N3602, N1821);
nor NOR4 (N3604, N3599, N37, N406, N1171);
or OR4 (N3605, N3594, N2454, N2859, N3527);
buf BUF1 (N3606, N3566);
buf BUF1 (N3607, N3593);
buf BUF1 (N3608, N3598);
nand NAND3 (N3609, N3608, N3175, N2307);
or OR4 (N3610, N3607, N870, N3538, N3104);
buf BUF1 (N3611, N3582);
buf BUF1 (N3612, N3600);
or OR3 (N3613, N3601, N3591, N1646);
buf BUF1 (N3614, N3605);
or OR2 (N3615, N3611, N3109);
or OR3 (N3616, N3609, N3449, N2515);
xor XOR2 (N3617, N3613, N1295);
nand NAND4 (N3618, N3610, N2058, N3056, N2272);
nor NOR4 (N3619, N3612, N2230, N3207, N2797);
or OR2 (N3620, N3606, N2573);
xor XOR2 (N3621, N3617, N1557);
buf BUF1 (N3622, N3616);
buf BUF1 (N3623, N3615);
not NOT1 (N3624, N3618);
or OR3 (N3625, N3597, N3407, N1161);
nor NOR2 (N3626, N3619, N2826);
nor NOR3 (N3627, N3620, N203, N1074);
and AND3 (N3628, N3614, N3579, N2825);
or OR4 (N3629, N3621, N638, N285, N2067);
not NOT1 (N3630, N3629);
nor NOR2 (N3631, N3604, N2998);
nand NAND4 (N3632, N3622, N802, N3419, N1097);
not NOT1 (N3633, N3631);
buf BUF1 (N3634, N3632);
nor NOR2 (N3635, N3624, N3623);
not NOT1 (N3636, N846);
and AND3 (N3637, N3630, N312, N2413);
nor NOR3 (N3638, N3626, N2787, N2267);
nand NAND4 (N3639, N3636, N3531, N1519, N3390);
xor XOR2 (N3640, N3639, N1292);
xor XOR2 (N3641, N3638, N3079);
not NOT1 (N3642, N3640);
and AND4 (N3643, N3603, N2266, N2516, N2543);
and AND3 (N3644, N3635, N240, N1262);
or OR3 (N3645, N3628, N3623, N129);
nor NOR4 (N3646, N3645, N1084, N3491, N189);
xor XOR2 (N3647, N3633, N1202);
xor XOR2 (N3648, N3625, N2211);
not NOT1 (N3649, N3647);
or OR2 (N3650, N3646, N2081);
buf BUF1 (N3651, N3650);
nor NOR2 (N3652, N3634, N2824);
and AND4 (N3653, N3643, N1118, N1094, N469);
or OR2 (N3654, N3653, N2195);
xor XOR2 (N3655, N3644, N2274);
and AND2 (N3656, N3642, N3219);
nand NAND3 (N3657, N3654, N2361, N2153);
or OR2 (N3658, N3648, N2739);
nand NAND4 (N3659, N3649, N2396, N1335, N1428);
nor NOR4 (N3660, N3637, N480, N3404, N3159);
xor XOR2 (N3661, N3651, N1879);
and AND3 (N3662, N3641, N3327, N1817);
nor NOR3 (N3663, N3657, N2077, N1924);
buf BUF1 (N3664, N3652);
nor NOR3 (N3665, N3664, N2524, N600);
not NOT1 (N3666, N3663);
and AND4 (N3667, N3660, N990, N627, N3207);
not NOT1 (N3668, N3667);
not NOT1 (N3669, N3666);
not NOT1 (N3670, N3656);
or OR3 (N3671, N3669, N2415, N2577);
nor NOR3 (N3672, N3662, N871, N3099);
nor NOR2 (N3673, N3670, N2958);
not NOT1 (N3674, N3671);
not NOT1 (N3675, N3665);
buf BUF1 (N3676, N3675);
not NOT1 (N3677, N3672);
nor NOR4 (N3678, N3658, N199, N2529, N3375);
and AND2 (N3679, N3676, N3146);
or OR2 (N3680, N3668, N2876);
not NOT1 (N3681, N3655);
and AND2 (N3682, N3677, N2480);
and AND3 (N3683, N3661, N3394, N2979);
or OR2 (N3684, N3673, N97);
nand NAND2 (N3685, N3680, N3061);
or OR4 (N3686, N3681, N1, N2206, N1645);
buf BUF1 (N3687, N3685);
buf BUF1 (N3688, N3627);
or OR4 (N3689, N3686, N329, N1613, N883);
nor NOR3 (N3690, N3687, N3430, N2882);
xor XOR2 (N3691, N3690, N1237);
buf BUF1 (N3692, N3691);
buf BUF1 (N3693, N3682);
nand NAND4 (N3694, N3679, N136, N1448, N1630);
and AND3 (N3695, N3674, N1781, N3646);
buf BUF1 (N3696, N3678);
not NOT1 (N3697, N3693);
xor XOR2 (N3698, N3694, N377);
nor NOR2 (N3699, N3684, N1210);
buf BUF1 (N3700, N3696);
xor XOR2 (N3701, N3683, N610);
and AND2 (N3702, N3700, N953);
nand NAND2 (N3703, N3659, N1042);
buf BUF1 (N3704, N3689);
nor NOR2 (N3705, N3688, N2835);
not NOT1 (N3706, N3695);
xor XOR2 (N3707, N3697, N401);
not NOT1 (N3708, N3704);
and AND2 (N3709, N3702, N69);
and AND2 (N3710, N3703, N2141);
and AND2 (N3711, N3692, N3541);
or OR2 (N3712, N3706, N369);
or OR2 (N3713, N3699, N2433);
buf BUF1 (N3714, N3708);
or OR2 (N3715, N3712, N76);
nand NAND3 (N3716, N3709, N485, N641);
or OR3 (N3717, N3710, N3384, N23);
or OR3 (N3718, N3701, N774, N1319);
buf BUF1 (N3719, N3717);
xor XOR2 (N3720, N3714, N2920);
nor NOR3 (N3721, N3718, N1789, N2844);
nor NOR2 (N3722, N3715, N271);
and AND2 (N3723, N3716, N1436);
buf BUF1 (N3724, N3720);
and AND3 (N3725, N3707, N1685, N2784);
and AND3 (N3726, N3721, N265, N342);
buf BUF1 (N3727, N3698);
not NOT1 (N3728, N3713);
buf BUF1 (N3729, N3727);
buf BUF1 (N3730, N3729);
nor NOR3 (N3731, N3722, N3104, N1141);
not NOT1 (N3732, N3731);
xor XOR2 (N3733, N3723, N3722);
or OR4 (N3734, N3724, N2520, N3047, N3211);
buf BUF1 (N3735, N3725);
not NOT1 (N3736, N3705);
and AND4 (N3737, N3735, N1713, N7, N1956);
buf BUF1 (N3738, N3728);
nand NAND2 (N3739, N3711, N1270);
not NOT1 (N3740, N3726);
buf BUF1 (N3741, N3736);
xor XOR2 (N3742, N3741, N3168);
nor NOR4 (N3743, N3738, N3458, N3247, N47);
xor XOR2 (N3744, N3743, N2459);
nand NAND3 (N3745, N3737, N1588, N1377);
xor XOR2 (N3746, N3739, N999);
nand NAND4 (N3747, N3732, N689, N648, N2010);
nand NAND2 (N3748, N3733, N3648);
nand NAND3 (N3749, N3748, N3077, N887);
buf BUF1 (N3750, N3745);
and AND2 (N3751, N3734, N808);
xor XOR2 (N3752, N3751, N102);
not NOT1 (N3753, N3730);
xor XOR2 (N3754, N3742, N3649);
not NOT1 (N3755, N3740);
or OR2 (N3756, N3719, N548);
and AND3 (N3757, N3744, N456, N3429);
or OR2 (N3758, N3747, N3641);
or OR4 (N3759, N3749, N3305, N262, N2952);
not NOT1 (N3760, N3754);
nor NOR4 (N3761, N3753, N2718, N3528, N1092);
nand NAND4 (N3762, N3755, N2304, N231, N2913);
nand NAND3 (N3763, N3762, N1926, N1782);
nor NOR2 (N3764, N3759, N193);
nand NAND2 (N3765, N3750, N2511);
not NOT1 (N3766, N3746);
buf BUF1 (N3767, N3764);
xor XOR2 (N3768, N3752, N1072);
nand NAND2 (N3769, N3761, N645);
and AND3 (N3770, N3769, N784, N2205);
not NOT1 (N3771, N3760);
nand NAND4 (N3772, N3757, N1833, N1825, N195);
nor NOR3 (N3773, N3763, N2490, N1259);
nor NOR3 (N3774, N3771, N441, N1387);
not NOT1 (N3775, N3768);
or OR3 (N3776, N3758, N270, N3265);
and AND3 (N3777, N3775, N565, N1167);
not NOT1 (N3778, N3765);
nand NAND2 (N3779, N3756, N800);
nor NOR3 (N3780, N3766, N2575, N1527);
xor XOR2 (N3781, N3773, N2369);
xor XOR2 (N3782, N3772, N534);
nor NOR4 (N3783, N3779, N1812, N1086, N1125);
xor XOR2 (N3784, N3776, N1685);
or OR2 (N3785, N3783, N3032);
not NOT1 (N3786, N3781);
or OR3 (N3787, N3785, N2493, N2493);
buf BUF1 (N3788, N3770);
or OR4 (N3789, N3782, N224, N2213, N3279);
or OR4 (N3790, N3777, N4, N3500, N619);
and AND4 (N3791, N3778, N3372, N337, N163);
xor XOR2 (N3792, N3790, N461);
xor XOR2 (N3793, N3792, N3183);
or OR4 (N3794, N3788, N1972, N2139, N3484);
buf BUF1 (N3795, N3787);
nand NAND3 (N3796, N3780, N349, N1856);
nor NOR4 (N3797, N3793, N1064, N1989, N3735);
and AND4 (N3798, N3767, N3132, N2009, N2149);
nor NOR4 (N3799, N3786, N2386, N215, N1221);
not NOT1 (N3800, N3784);
or OR4 (N3801, N3789, N847, N2782, N3347);
or OR2 (N3802, N3799, N810);
or OR3 (N3803, N3795, N3523, N2563);
or OR4 (N3804, N3794, N1639, N1934, N3403);
and AND4 (N3805, N3802, N1153, N2330, N1487);
and AND3 (N3806, N3796, N1160, N3017);
buf BUF1 (N3807, N3791);
and AND4 (N3808, N3805, N581, N1406, N613);
or OR4 (N3809, N3806, N2484, N2405, N1435);
not NOT1 (N3810, N3800);
xor XOR2 (N3811, N3774, N1907);
buf BUF1 (N3812, N3809);
nand NAND4 (N3813, N3810, N2427, N2617, N1567);
or OR2 (N3814, N3803, N1482);
and AND3 (N3815, N3801, N495, N2623);
buf BUF1 (N3816, N3815);
not NOT1 (N3817, N3816);
buf BUF1 (N3818, N3817);
and AND3 (N3819, N3811, N2537, N679);
nor NOR3 (N3820, N3819, N2876, N2675);
xor XOR2 (N3821, N3804, N2000);
not NOT1 (N3822, N3812);
nand NAND3 (N3823, N3814, N1367, N639);
and AND2 (N3824, N3807, N3280);
or OR2 (N3825, N3798, N2371);
buf BUF1 (N3826, N3824);
nor NOR2 (N3827, N3826, N3537);
and AND4 (N3828, N3813, N1870, N1092, N202);
nor NOR3 (N3829, N3818, N598, N501);
xor XOR2 (N3830, N3825, N780);
not NOT1 (N3831, N3827);
or OR2 (N3832, N3821, N1445);
or OR3 (N3833, N3830, N2803, N267);
not NOT1 (N3834, N3828);
nor NOR3 (N3835, N3833, N2198, N3634);
and AND3 (N3836, N3823, N719, N2014);
buf BUF1 (N3837, N3808);
or OR4 (N3838, N3822, N1872, N373, N3801);
nand NAND2 (N3839, N3832, N3458);
and AND2 (N3840, N3836, N2824);
buf BUF1 (N3841, N3839);
not NOT1 (N3842, N3838);
and AND2 (N3843, N3835, N1726);
xor XOR2 (N3844, N3829, N2597);
nor NOR3 (N3845, N3841, N3272, N2201);
and AND2 (N3846, N3843, N502);
xor XOR2 (N3847, N3797, N723);
and AND2 (N3848, N3844, N2562);
xor XOR2 (N3849, N3820, N1026);
xor XOR2 (N3850, N3831, N3317);
nand NAND2 (N3851, N3834, N1373);
and AND4 (N3852, N3849, N893, N3385, N74);
not NOT1 (N3853, N3837);
not NOT1 (N3854, N3852);
not NOT1 (N3855, N3854);
nor NOR4 (N3856, N3846, N2883, N1233, N3084);
nand NAND3 (N3857, N3851, N2776, N242);
nor NOR4 (N3858, N3855, N738, N3206, N3684);
not NOT1 (N3859, N3858);
buf BUF1 (N3860, N3853);
or OR2 (N3861, N3845, N500);
nor NOR3 (N3862, N3856, N1087, N390);
and AND2 (N3863, N3842, N2747);
buf BUF1 (N3864, N3863);
nor NOR2 (N3865, N3861, N1971);
or OR3 (N3866, N3860, N3618, N1970);
buf BUF1 (N3867, N3866);
nand NAND2 (N3868, N3848, N202);
not NOT1 (N3869, N3840);
buf BUF1 (N3870, N3865);
xor XOR2 (N3871, N3862, N1681);
buf BUF1 (N3872, N3867);
nand NAND4 (N3873, N3847, N1645, N2498, N3721);
xor XOR2 (N3874, N3850, N1232);
xor XOR2 (N3875, N3864, N1597);
and AND4 (N3876, N3869, N398, N3485, N748);
xor XOR2 (N3877, N3868, N2023);
nor NOR3 (N3878, N3857, N2417, N2248);
buf BUF1 (N3879, N3872);
or OR2 (N3880, N3870, N265);
and AND2 (N3881, N3871, N3462);
or OR2 (N3882, N3875, N796);
nand NAND4 (N3883, N3859, N491, N2025, N545);
buf BUF1 (N3884, N3882);
or OR4 (N3885, N3878, N3624, N2268, N962);
or OR4 (N3886, N3884, N1488, N3568, N2384);
buf BUF1 (N3887, N3876);
or OR2 (N3888, N3886, N2289);
nor NOR2 (N3889, N3880, N676);
or OR4 (N3890, N3885, N3399, N1099, N3466);
or OR3 (N3891, N3881, N2314, N3089);
buf BUF1 (N3892, N3888);
nor NOR3 (N3893, N3879, N2030, N3741);
nor NOR3 (N3894, N3883, N3356, N476);
nor NOR3 (N3895, N3891, N3875, N1832);
not NOT1 (N3896, N3873);
xor XOR2 (N3897, N3896, N1177);
nand NAND2 (N3898, N3890, N374);
nand NAND3 (N3899, N3895, N821, N3790);
buf BUF1 (N3900, N3897);
and AND4 (N3901, N3894, N259, N2034, N1870);
buf BUF1 (N3902, N3898);
xor XOR2 (N3903, N3901, N1071);
nand NAND3 (N3904, N3893, N2093, N3534);
xor XOR2 (N3905, N3903, N146);
nand NAND4 (N3906, N3874, N1704, N3261, N738);
xor XOR2 (N3907, N3899, N1229);
and AND4 (N3908, N3905, N1485, N2777, N2176);
or OR2 (N3909, N3900, N428);
buf BUF1 (N3910, N3892);
xor XOR2 (N3911, N3907, N498);
and AND4 (N3912, N3908, N1213, N3414, N1273);
xor XOR2 (N3913, N3906, N1720);
not NOT1 (N3914, N3912);
and AND4 (N3915, N3902, N207, N2159, N1140);
nor NOR2 (N3916, N3911, N737);
xor XOR2 (N3917, N3877, N2939);
nor NOR3 (N3918, N3889, N235, N2279);
xor XOR2 (N3919, N3914, N2013);
and AND2 (N3920, N3910, N1407);
buf BUF1 (N3921, N3917);
nand NAND4 (N3922, N3919, N1269, N90, N1815);
nand NAND2 (N3923, N3918, N695);
nor NOR4 (N3924, N3923, N674, N1142, N199);
xor XOR2 (N3925, N3921, N2052);
xor XOR2 (N3926, N3887, N484);
nand NAND3 (N3927, N3926, N1005, N651);
xor XOR2 (N3928, N3924, N683);
buf BUF1 (N3929, N3916);
or OR4 (N3930, N3925, N37, N2933, N2235);
and AND2 (N3931, N3920, N1904);
nand NAND2 (N3932, N3928, N482);
xor XOR2 (N3933, N3909, N3272);
xor XOR2 (N3934, N3929, N3561);
and AND4 (N3935, N3930, N51, N1181, N881);
not NOT1 (N3936, N3922);
xor XOR2 (N3937, N3913, N3560);
and AND2 (N3938, N3931, N730);
nand NAND2 (N3939, N3934, N2005);
nor NOR3 (N3940, N3938, N3535, N2774);
xor XOR2 (N3941, N3927, N480);
not NOT1 (N3942, N3904);
xor XOR2 (N3943, N3942, N3890);
and AND3 (N3944, N3937, N2379, N2628);
xor XOR2 (N3945, N3932, N3639);
or OR3 (N3946, N3941, N2273, N3289);
buf BUF1 (N3947, N3915);
nor NOR3 (N3948, N3945, N1011, N2536);
nor NOR4 (N3949, N3947, N993, N587, N3415);
nand NAND2 (N3950, N3948, N3819);
not NOT1 (N3951, N3943);
nand NAND4 (N3952, N3951, N457, N3169, N2234);
buf BUF1 (N3953, N3940);
xor XOR2 (N3954, N3949, N2956);
not NOT1 (N3955, N3944);
xor XOR2 (N3956, N3952, N2075);
xor XOR2 (N3957, N3954, N3918);
buf BUF1 (N3958, N3950);
not NOT1 (N3959, N3958);
xor XOR2 (N3960, N3953, N849);
xor XOR2 (N3961, N3935, N1115);
buf BUF1 (N3962, N3957);
nand NAND2 (N3963, N3961, N1661);
or OR4 (N3964, N3955, N2929, N1219, N1886);
nor NOR3 (N3965, N3964, N670, N784);
nor NOR3 (N3966, N3946, N2591, N1430);
buf BUF1 (N3967, N3966);
and AND2 (N3968, N3960, N1348);
nand NAND2 (N3969, N3936, N1551);
nand NAND2 (N3970, N3956, N571);
or OR4 (N3971, N3970, N3748, N1067, N3663);
and AND2 (N3972, N3969, N3890);
nor NOR3 (N3973, N3939, N3844, N64);
buf BUF1 (N3974, N3972);
nor NOR4 (N3975, N3973, N2983, N1751, N3582);
nor NOR4 (N3976, N3974, N2395, N1282, N629);
nand NAND2 (N3977, N3959, N311);
xor XOR2 (N3978, N3963, N1414);
buf BUF1 (N3979, N3976);
nand NAND3 (N3980, N3977, N927, N1002);
buf BUF1 (N3981, N3967);
not NOT1 (N3982, N3975);
nor NOR2 (N3983, N3979, N1322);
not NOT1 (N3984, N3968);
not NOT1 (N3985, N3984);
not NOT1 (N3986, N3980);
and AND3 (N3987, N3933, N1181, N2160);
and AND3 (N3988, N3985, N2020, N3567);
xor XOR2 (N3989, N3983, N1578);
buf BUF1 (N3990, N3988);
and AND2 (N3991, N3989, N2730);
or OR2 (N3992, N3978, N1546);
not NOT1 (N3993, N3971);
nand NAND4 (N3994, N3962, N2398, N2414, N3528);
buf BUF1 (N3995, N3994);
nand NAND3 (N3996, N3986, N3782, N2016);
nand NAND4 (N3997, N3981, N312, N3015, N1627);
buf BUF1 (N3998, N3965);
and AND3 (N3999, N3990, N1430, N2924);
nor NOR2 (N4000, N3997, N3462);
buf BUF1 (N4001, N3999);
and AND3 (N4002, N3982, N1803, N1277);
buf BUF1 (N4003, N3995);
nand NAND3 (N4004, N3996, N2170, N2419);
or OR2 (N4005, N3987, N2072);
not NOT1 (N4006, N4003);
xor XOR2 (N4007, N4002, N3032);
and AND3 (N4008, N3993, N3593, N443);
or OR2 (N4009, N4006, N1727);
or OR4 (N4010, N4005, N1926, N2939, N2974);
nor NOR3 (N4011, N4009, N1377, N3402);
and AND3 (N4012, N4007, N1132, N2790);
not NOT1 (N4013, N4012);
buf BUF1 (N4014, N4011);
not NOT1 (N4015, N4014);
nand NAND2 (N4016, N4000, N616);
not NOT1 (N4017, N4016);
buf BUF1 (N4018, N4013);
xor XOR2 (N4019, N4018, N800);
buf BUF1 (N4020, N4017);
xor XOR2 (N4021, N4020, N1606);
and AND4 (N4022, N4015, N2600, N2042, N3246);
nand NAND4 (N4023, N3991, N1300, N1839, N3719);
buf BUF1 (N4024, N3998);
buf BUF1 (N4025, N3992);
nor NOR4 (N4026, N4008, N1287, N1102, N3586);
nand NAND2 (N4027, N4022, N2968);
or OR2 (N4028, N4001, N3091);
and AND3 (N4029, N4024, N1039, N336);
buf BUF1 (N4030, N4023);
nand NAND4 (N4031, N4025, N3212, N1558, N3244);
buf BUF1 (N4032, N4029);
and AND2 (N4033, N4010, N375);
and AND3 (N4034, N4032, N3440, N3785);
nand NAND3 (N4035, N4028, N3287, N2959);
nand NAND4 (N4036, N4031, N2525, N1457, N1618);
nor NOR3 (N4037, N4035, N1680, N1228);
xor XOR2 (N4038, N4036, N3087);
or OR4 (N4039, N4030, N337, N659, N793);
nand NAND2 (N4040, N4037, N3463);
not NOT1 (N4041, N4019);
not NOT1 (N4042, N4039);
or OR3 (N4043, N4033, N497, N510);
or OR3 (N4044, N4041, N3584, N1679);
nor NOR2 (N4045, N4040, N2930);
nand NAND4 (N4046, N4043, N1970, N2279, N581);
not NOT1 (N4047, N4046);
xor XOR2 (N4048, N4034, N2473);
nand NAND3 (N4049, N4021, N2612, N536);
buf BUF1 (N4050, N4042);
or OR4 (N4051, N4048, N1900, N2163, N1949);
buf BUF1 (N4052, N4044);
buf BUF1 (N4053, N4049);
buf BUF1 (N4054, N4045);
not NOT1 (N4055, N4051);
nand NAND3 (N4056, N4004, N3266, N3369);
nor NOR3 (N4057, N4047, N3269, N327);
buf BUF1 (N4058, N4027);
buf BUF1 (N4059, N4055);
and AND2 (N4060, N4026, N3037);
not NOT1 (N4061, N4056);
or OR3 (N4062, N4058, N1642, N3436);
or OR2 (N4063, N4054, N1060);
nand NAND3 (N4064, N4052, N3576, N1176);
or OR4 (N4065, N4057, N1081, N1814, N3632);
nand NAND3 (N4066, N4065, N1090, N2744);
nor NOR3 (N4067, N4050, N2816, N82);
nor NOR3 (N4068, N4038, N1643, N2838);
and AND2 (N4069, N4067, N3984);
and AND2 (N4070, N4059, N328);
buf BUF1 (N4071, N4063);
nor NOR4 (N4072, N4066, N2073, N1533, N1096);
or OR3 (N4073, N4072, N2288, N1740);
xor XOR2 (N4074, N4073, N356);
buf BUF1 (N4075, N4070);
nand NAND2 (N4076, N4060, N1590);
or OR2 (N4077, N4062, N1867);
buf BUF1 (N4078, N4064);
buf BUF1 (N4079, N4071);
nand NAND4 (N4080, N4078, N2377, N3459, N1276);
nor NOR2 (N4081, N4069, N81);
buf BUF1 (N4082, N4081);
xor XOR2 (N4083, N4077, N1591);
and AND4 (N4084, N4075, N2104, N303, N3489);
nor NOR2 (N4085, N4074, N1078);
nor NOR3 (N4086, N4082, N1540, N2174);
nand NAND2 (N4087, N4086, N2983);
xor XOR2 (N4088, N4087, N3781);
xor XOR2 (N4089, N4084, N1432);
and AND2 (N4090, N4079, N607);
or OR2 (N4091, N4053, N1839);
nor NOR2 (N4092, N4068, N382);
and AND4 (N4093, N4076, N3653, N3616, N3805);
nand NAND3 (N4094, N4093, N3902, N2658);
and AND2 (N4095, N4085, N3150);
not NOT1 (N4096, N4090);
nand NAND2 (N4097, N4083, N3561);
nor NOR2 (N4098, N4094, N625);
not NOT1 (N4099, N4098);
nor NOR2 (N4100, N4095, N1218);
nor NOR2 (N4101, N4100, N1753);
xor XOR2 (N4102, N4092, N1967);
xor XOR2 (N4103, N4096, N2038);
or OR2 (N4104, N4099, N516);
xor XOR2 (N4105, N4103, N3847);
buf BUF1 (N4106, N4101);
nor NOR2 (N4107, N4091, N1075);
and AND4 (N4108, N4102, N552, N3251, N2263);
nor NOR4 (N4109, N4080, N2606, N3801, N764);
nor NOR4 (N4110, N4061, N2132, N1186, N2361);
not NOT1 (N4111, N4110);
xor XOR2 (N4112, N4097, N1691);
or OR3 (N4113, N4107, N234, N342);
not NOT1 (N4114, N4109);
xor XOR2 (N4115, N4106, N2918);
not NOT1 (N4116, N4113);
xor XOR2 (N4117, N4116, N661);
nand NAND4 (N4118, N4111, N2218, N1045, N2537);
nor NOR4 (N4119, N4112, N3135, N2408, N4003);
xor XOR2 (N4120, N4108, N3915);
nand NAND2 (N4121, N4114, N2998);
nor NOR3 (N4122, N4088, N1878, N1170);
and AND2 (N4123, N4115, N2147);
nor NOR3 (N4124, N4117, N3205, N629);
not NOT1 (N4125, N4123);
nor NOR3 (N4126, N4124, N971, N2901);
buf BUF1 (N4127, N4126);
and AND2 (N4128, N4104, N2901);
xor XOR2 (N4129, N4105, N671);
or OR2 (N4130, N4127, N2323);
nand NAND4 (N4131, N4120, N2933, N1530, N2582);
nor NOR4 (N4132, N4129, N2926, N3052, N2745);
nor NOR3 (N4133, N4119, N452, N545);
not NOT1 (N4134, N4121);
nor NOR2 (N4135, N4132, N1592);
and AND4 (N4136, N4128, N1276, N2957, N1979);
and AND2 (N4137, N4130, N4102);
or OR4 (N4138, N4133, N1754, N2860, N2117);
buf BUF1 (N4139, N4138);
xor XOR2 (N4140, N4131, N3643);
or OR4 (N4141, N4125, N102, N2129, N1490);
not NOT1 (N4142, N4137);
or OR3 (N4143, N4141, N3733, N2310);
and AND3 (N4144, N4140, N4074, N108);
nand NAND2 (N4145, N4089, N1944);
nand NAND2 (N4146, N4143, N2079);
and AND4 (N4147, N4139, N2016, N516, N2325);
xor XOR2 (N4148, N4134, N48);
nor NOR3 (N4149, N4144, N237, N3318);
and AND4 (N4150, N4118, N560, N2601, N2112);
nor NOR3 (N4151, N4147, N4143, N267);
xor XOR2 (N4152, N4142, N781);
or OR4 (N4153, N4145, N217, N5, N661);
xor XOR2 (N4154, N4146, N1383);
xor XOR2 (N4155, N4135, N2115);
xor XOR2 (N4156, N4152, N972);
buf BUF1 (N4157, N4155);
nor NOR4 (N4158, N4151, N635, N4143, N590);
nor NOR4 (N4159, N4149, N3296, N31, N3487);
xor XOR2 (N4160, N4157, N3907);
not NOT1 (N4161, N4160);
and AND4 (N4162, N4154, N1381, N1376, N4119);
xor XOR2 (N4163, N4158, N1080);
not NOT1 (N4164, N4161);
xor XOR2 (N4165, N4162, N3107);
and AND3 (N4166, N4153, N3813, N1338);
buf BUF1 (N4167, N4156);
not NOT1 (N4168, N4148);
nor NOR2 (N4169, N4166, N3449);
not NOT1 (N4170, N4164);
nor NOR2 (N4171, N4159, N74);
not NOT1 (N4172, N4169);
xor XOR2 (N4173, N4168, N859);
nand NAND2 (N4174, N4171, N2292);
or OR3 (N4175, N4174, N1039, N689);
nor NOR2 (N4176, N4165, N78);
xor XOR2 (N4177, N4176, N3911);
nand NAND2 (N4178, N4163, N1040);
not NOT1 (N4179, N4150);
and AND4 (N4180, N4136, N3769, N3518, N724);
not NOT1 (N4181, N4179);
not NOT1 (N4182, N4170);
nor NOR4 (N4183, N4167, N3778, N1364, N854);
or OR2 (N4184, N4181, N3316);
not NOT1 (N4185, N4175);
nand NAND2 (N4186, N4122, N227);
xor XOR2 (N4187, N4182, N3298);
nand NAND3 (N4188, N4185, N3162, N3472);
xor XOR2 (N4189, N4183, N2777);
not NOT1 (N4190, N4172);
nor NOR3 (N4191, N4190, N478, N1149);
buf BUF1 (N4192, N4189);
buf BUF1 (N4193, N4191);
nand NAND4 (N4194, N4187, N1247, N952, N1435);
and AND2 (N4195, N4184, N2431);
not NOT1 (N4196, N4186);
and AND4 (N4197, N4178, N2578, N1153, N1782);
buf BUF1 (N4198, N4197);
and AND4 (N4199, N4193, N3462, N3413, N3583);
xor XOR2 (N4200, N4177, N4152);
xor XOR2 (N4201, N4200, N910);
not NOT1 (N4202, N4173);
or OR3 (N4203, N4180, N3865, N4052);
and AND2 (N4204, N4195, N1371);
not NOT1 (N4205, N4201);
buf BUF1 (N4206, N4198);
xor XOR2 (N4207, N4204, N2113);
nor NOR4 (N4208, N4207, N1775, N1850, N549);
nand NAND2 (N4209, N4205, N1862);
and AND2 (N4210, N4209, N2801);
xor XOR2 (N4211, N4208, N790);
not NOT1 (N4212, N4192);
or OR4 (N4213, N4196, N1901, N3796, N656);
or OR4 (N4214, N4188, N3544, N2682, N2257);
and AND3 (N4215, N4194, N3658, N2791);
buf BUF1 (N4216, N4210);
or OR4 (N4217, N4202, N1397, N3709, N3499);
xor XOR2 (N4218, N4217, N820);
not NOT1 (N4219, N4203);
and AND2 (N4220, N4214, N3745);
and AND3 (N4221, N4212, N3775, N1359);
nor NOR3 (N4222, N4206, N1923, N3310);
and AND3 (N4223, N4213, N509, N3328);
and AND2 (N4224, N4216, N1077);
or OR2 (N4225, N4222, N3300);
nor NOR3 (N4226, N4223, N1832, N274);
nor NOR4 (N4227, N4224, N1731, N1526, N4005);
buf BUF1 (N4228, N4211);
nand NAND2 (N4229, N4226, N1243);
nand NAND2 (N4230, N4215, N3053);
buf BUF1 (N4231, N4229);
and AND4 (N4232, N4221, N567, N3864, N772);
and AND3 (N4233, N4219, N2459, N3484);
buf BUF1 (N4234, N4199);
not NOT1 (N4235, N4218);
nor NOR3 (N4236, N4235, N1656, N3788);
not NOT1 (N4237, N4234);
nor NOR4 (N4238, N4231, N824, N203, N2760);
nand NAND2 (N4239, N4232, N3893);
and AND2 (N4240, N4236, N2882);
or OR2 (N4241, N4233, N2751);
nand NAND2 (N4242, N4228, N1490);
xor XOR2 (N4243, N4227, N4);
not NOT1 (N4244, N4241);
xor XOR2 (N4245, N4225, N1444);
nor NOR4 (N4246, N4237, N2387, N887, N2120);
xor XOR2 (N4247, N4240, N1275);
nand NAND2 (N4248, N4247, N3709);
nor NOR3 (N4249, N4248, N1686, N2097);
buf BUF1 (N4250, N4245);
xor XOR2 (N4251, N4242, N455);
nand NAND3 (N4252, N4244, N3491, N3519);
xor XOR2 (N4253, N4243, N1186);
nand NAND3 (N4254, N4238, N412, N2839);
nor NOR2 (N4255, N4220, N370);
buf BUF1 (N4256, N4253);
nand NAND2 (N4257, N4230, N2482);
nand NAND2 (N4258, N4250, N332);
buf BUF1 (N4259, N4251);
and AND2 (N4260, N4256, N604);
or OR2 (N4261, N4258, N835);
or OR4 (N4262, N4239, N3327, N2452, N3969);
and AND3 (N4263, N4254, N924, N1492);
not NOT1 (N4264, N4249);
or OR2 (N4265, N4246, N667);
buf BUF1 (N4266, N4264);
not NOT1 (N4267, N4257);
not NOT1 (N4268, N4266);
not NOT1 (N4269, N4262);
or OR3 (N4270, N4268, N2646, N2137);
or OR2 (N4271, N4259, N2007);
nor NOR3 (N4272, N4255, N2526, N435);
xor XOR2 (N4273, N4261, N2046);
xor XOR2 (N4274, N4267, N3889);
not NOT1 (N4275, N4252);
buf BUF1 (N4276, N4270);
buf BUF1 (N4277, N4273);
not NOT1 (N4278, N4263);
and AND3 (N4279, N4276, N1310, N2852);
xor XOR2 (N4280, N4260, N651);
buf BUF1 (N4281, N4272);
xor XOR2 (N4282, N4269, N3325);
xor XOR2 (N4283, N4274, N1185);
or OR3 (N4284, N4281, N4030, N3982);
and AND3 (N4285, N4284, N1572, N2854);
and AND3 (N4286, N4285, N850, N1869);
not NOT1 (N4287, N4275);
nand NAND2 (N4288, N4287, N3626);
nand NAND3 (N4289, N4278, N3877, N2255);
not NOT1 (N4290, N4280);
buf BUF1 (N4291, N4289);
nand NAND4 (N4292, N4271, N1150, N539, N2110);
nor NOR3 (N4293, N4277, N1095, N2738);
nor NOR2 (N4294, N4282, N1001);
nand NAND3 (N4295, N4286, N670, N1830);
nand NAND4 (N4296, N4295, N3129, N2407, N4086);
or OR2 (N4297, N4288, N3044);
not NOT1 (N4298, N4292);
nand NAND3 (N4299, N4293, N2133, N3996);
nor NOR4 (N4300, N4291, N3231, N341, N3374);
xor XOR2 (N4301, N4298, N3052);
not NOT1 (N4302, N4296);
and AND4 (N4303, N4300, N1028, N3147, N2481);
or OR2 (N4304, N4294, N2635);
nor NOR4 (N4305, N4279, N807, N1538, N2356);
or OR3 (N4306, N4290, N1180, N2256);
xor XOR2 (N4307, N4303, N1585);
and AND2 (N4308, N4297, N1495);
or OR4 (N4309, N4308, N4174, N1283, N655);
or OR4 (N4310, N4302, N342, N4117, N3072);
not NOT1 (N4311, N4283);
nand NAND3 (N4312, N4265, N4127, N1357);
nor NOR2 (N4313, N4306, N1892);
nand NAND3 (N4314, N4309, N525, N2349);
nand NAND3 (N4315, N4310, N1090, N3832);
xor XOR2 (N4316, N4299, N2360);
xor XOR2 (N4317, N4305, N2577);
or OR4 (N4318, N4301, N3305, N1151, N2127);
nor NOR4 (N4319, N4311, N2204, N3348, N1484);
nor NOR3 (N4320, N4314, N1266, N1875);
or OR4 (N4321, N4318, N3192, N1244, N3763);
buf BUF1 (N4322, N4317);
and AND4 (N4323, N4312, N459, N2909, N946);
not NOT1 (N4324, N4304);
and AND2 (N4325, N4321, N1722);
not NOT1 (N4326, N4313);
not NOT1 (N4327, N4315);
or OR4 (N4328, N4325, N3056, N1977, N3456);
nor NOR3 (N4329, N4319, N2205, N2263);
nor NOR3 (N4330, N4329, N2382, N3200);
buf BUF1 (N4331, N4326);
and AND4 (N4332, N4323, N3516, N2439, N4043);
buf BUF1 (N4333, N4322);
and AND3 (N4334, N4328, N272, N2208);
buf BUF1 (N4335, N4331);
xor XOR2 (N4336, N4320, N1510);
or OR2 (N4337, N4332, N2513);
nand NAND4 (N4338, N4336, N3869, N428, N3826);
buf BUF1 (N4339, N4335);
not NOT1 (N4340, N4339);
nand NAND4 (N4341, N4327, N1555, N3512, N3604);
xor XOR2 (N4342, N4334, N911);
and AND4 (N4343, N4340, N1418, N2898, N1917);
buf BUF1 (N4344, N4330);
not NOT1 (N4345, N4342);
nand NAND3 (N4346, N4307, N3334, N654);
or OR4 (N4347, N4346, N3045, N617, N3874);
and AND2 (N4348, N4344, N3603);
not NOT1 (N4349, N4348);
not NOT1 (N4350, N4337);
or OR2 (N4351, N4341, N3678);
xor XOR2 (N4352, N4350, N382);
xor XOR2 (N4353, N4324, N2463);
or OR3 (N4354, N4333, N3322, N2930);
nor NOR3 (N4355, N4338, N4083, N1149);
buf BUF1 (N4356, N4353);
or OR4 (N4357, N4351, N873, N3252, N2986);
not NOT1 (N4358, N4347);
and AND3 (N4359, N4354, N2502, N903);
nor NOR2 (N4360, N4356, N1557);
not NOT1 (N4361, N4358);
nand NAND4 (N4362, N4361, N1408, N4300, N3319);
or OR3 (N4363, N4316, N700, N3995);
nand NAND3 (N4364, N4357, N4181, N1460);
nor NOR3 (N4365, N4355, N3952, N201);
nor NOR4 (N4366, N4349, N41, N2184, N1781);
nor NOR2 (N4367, N4352, N1148);
nor NOR3 (N4368, N4364, N1264, N565);
and AND2 (N4369, N4359, N3215);
not NOT1 (N4370, N4368);
nand NAND4 (N4371, N4370, N4319, N3236, N794);
nor NOR4 (N4372, N4343, N1467, N3077, N3896);
nor NOR2 (N4373, N4367, N1481);
nor NOR2 (N4374, N4363, N3679);
or OR3 (N4375, N4366, N389, N4122);
nor NOR2 (N4376, N4373, N1669);
nand NAND2 (N4377, N4374, N4111);
xor XOR2 (N4378, N4362, N2859);
nor NOR4 (N4379, N4376, N1593, N2559, N2807);
nor NOR4 (N4380, N4377, N690, N2250, N3391);
xor XOR2 (N4381, N4378, N3953);
buf BUF1 (N4382, N4365);
nand NAND3 (N4383, N4371, N2500, N877);
and AND4 (N4384, N4345, N789, N1516, N3691);
buf BUF1 (N4385, N4382);
xor XOR2 (N4386, N4369, N4192);
not NOT1 (N4387, N4383);
and AND2 (N4388, N4381, N1035);
xor XOR2 (N4389, N4379, N1536);
xor XOR2 (N4390, N4375, N1507);
and AND3 (N4391, N4385, N292, N3516);
nor NOR2 (N4392, N4360, N1301);
nand NAND2 (N4393, N4388, N2628);
nand NAND2 (N4394, N4380, N1890);
or OR2 (N4395, N4387, N450);
nand NAND4 (N4396, N4372, N3064, N1581, N1319);
not NOT1 (N4397, N4389);
nand NAND2 (N4398, N4391, N3091);
nor NOR2 (N4399, N4395, N4273);
buf BUF1 (N4400, N4396);
and AND3 (N4401, N4394, N4356, N2281);
nor NOR4 (N4402, N4390, N1341, N2050, N4111);
buf BUF1 (N4403, N4400);
buf BUF1 (N4404, N4384);
buf BUF1 (N4405, N4402);
nor NOR2 (N4406, N4405, N2535);
nand NAND4 (N4407, N4399, N770, N3360, N3156);
xor XOR2 (N4408, N4393, N2673);
nor NOR4 (N4409, N4404, N866, N1234, N1679);
xor XOR2 (N4410, N4409, N3665);
nand NAND2 (N4411, N4386, N2243);
or OR4 (N4412, N4410, N3565, N2363, N556);
nand NAND4 (N4413, N4398, N3609, N3936, N3631);
and AND3 (N4414, N4411, N2595, N1683);
xor XOR2 (N4415, N4392, N2339);
nand NAND4 (N4416, N4407, N3908, N235, N1678);
nand NAND3 (N4417, N4397, N899, N3048);
nand NAND3 (N4418, N4403, N274, N4346);
not NOT1 (N4419, N4414);
nand NAND2 (N4420, N4408, N1316);
buf BUF1 (N4421, N4420);
nand NAND3 (N4422, N4415, N1862, N29);
or OR3 (N4423, N4417, N3198, N1892);
or OR3 (N4424, N4413, N4254, N1356);
buf BUF1 (N4425, N4416);
nor NOR4 (N4426, N4406, N421, N4323, N698);
or OR4 (N4427, N4418, N2702, N356, N1823);
xor XOR2 (N4428, N4419, N1279);
not NOT1 (N4429, N4427);
buf BUF1 (N4430, N4423);
not NOT1 (N4431, N4421);
xor XOR2 (N4432, N4422, N508);
nor NOR2 (N4433, N4431, N3222);
nand NAND4 (N4434, N4412, N3165, N826, N1073);
xor XOR2 (N4435, N4425, N2955);
buf BUF1 (N4436, N4429);
not NOT1 (N4437, N4428);
and AND2 (N4438, N4424, N3179);
and AND3 (N4439, N4433, N2721, N472);
nand NAND2 (N4440, N4430, N794);
and AND2 (N4441, N4434, N3726);
nand NAND2 (N4442, N4435, N1499);
nand NAND3 (N4443, N4436, N2736, N3189);
nand NAND4 (N4444, N4437, N4213, N530, N1068);
or OR4 (N4445, N4426, N4377, N3189, N3081);
buf BUF1 (N4446, N4444);
nand NAND4 (N4447, N4439, N75, N2237, N3977);
or OR4 (N4448, N4441, N2436, N2465, N2011);
nor NOR3 (N4449, N4432, N1046, N3390);
nand NAND3 (N4450, N4442, N2963, N1974);
not NOT1 (N4451, N4446);
or OR4 (N4452, N4445, N44, N1148, N1354);
nor NOR3 (N4453, N4447, N2654, N2863);
not NOT1 (N4454, N4401);
and AND3 (N4455, N4449, N1207, N523);
not NOT1 (N4456, N4455);
not NOT1 (N4457, N4450);
not NOT1 (N4458, N4452);
not NOT1 (N4459, N4451);
and AND4 (N4460, N4454, N2587, N1181, N3851);
nand NAND2 (N4461, N4438, N998);
xor XOR2 (N4462, N4458, N4139);
and AND4 (N4463, N4456, N2266, N4064, N4422);
xor XOR2 (N4464, N4462, N1347);
nor NOR3 (N4465, N4453, N1230, N3373);
nor NOR4 (N4466, N4457, N2415, N2375, N2967);
xor XOR2 (N4467, N4448, N536);
and AND2 (N4468, N4443, N1943);
nor NOR4 (N4469, N4468, N6, N164, N3757);
not NOT1 (N4470, N4467);
nor NOR4 (N4471, N4466, N300, N341, N2481);
and AND3 (N4472, N4470, N955, N985);
nor NOR4 (N4473, N4472, N2427, N1641, N2207);
xor XOR2 (N4474, N4471, N1370);
nand NAND2 (N4475, N4473, N2499);
and AND3 (N4476, N4464, N2590, N3226);
buf BUF1 (N4477, N4465);
nand NAND2 (N4478, N4469, N106);
and AND2 (N4479, N4476, N2203);
not NOT1 (N4480, N4478);
not NOT1 (N4481, N4480);
xor XOR2 (N4482, N4477, N3117);
buf BUF1 (N4483, N4474);
xor XOR2 (N4484, N4460, N1728);
not NOT1 (N4485, N4459);
nor NOR4 (N4486, N4485, N157, N229, N1448);
buf BUF1 (N4487, N4461);
nand NAND3 (N4488, N4484, N4472, N1916);
nand NAND4 (N4489, N4440, N2264, N1306, N3492);
and AND4 (N4490, N4489, N2304, N3881, N1099);
buf BUF1 (N4491, N4486);
nand NAND2 (N4492, N4475, N1060);
or OR4 (N4493, N4483, N2678, N1464, N3787);
xor XOR2 (N4494, N4481, N3894);
buf BUF1 (N4495, N4490);
xor XOR2 (N4496, N4495, N3031);
or OR4 (N4497, N4482, N4265, N2313, N67);
and AND2 (N4498, N4488, N200);
or OR2 (N4499, N4497, N3184);
nand NAND4 (N4500, N4491, N1792, N3694, N3962);
not NOT1 (N4501, N4479);
buf BUF1 (N4502, N4492);
or OR2 (N4503, N4500, N1217);
and AND3 (N4504, N4499, N929, N2952);
nor NOR3 (N4505, N4493, N3911, N749);
or OR3 (N4506, N4503, N2396, N3069);
and AND3 (N4507, N4504, N3751, N867);
nor NOR3 (N4508, N4507, N1683, N4247);
and AND2 (N4509, N4508, N758);
nor NOR2 (N4510, N4496, N3683);
or OR4 (N4511, N4505, N1773, N2283, N1604);
or OR2 (N4512, N4506, N4433);
and AND4 (N4513, N4498, N2931, N2060, N1164);
nand NAND4 (N4514, N4463, N1455, N4449, N3404);
xor XOR2 (N4515, N4494, N3399);
or OR2 (N4516, N4511, N3961);
nor NOR4 (N4517, N4512, N111, N1306, N1132);
nand NAND3 (N4518, N4514, N4045, N3780);
nor NOR3 (N4519, N4516, N2608, N1590);
buf BUF1 (N4520, N4502);
not NOT1 (N4521, N4487);
xor XOR2 (N4522, N4521, N1577);
buf BUF1 (N4523, N4517);
nor NOR2 (N4524, N4510, N2054);
nor NOR4 (N4525, N4523, N3793, N739, N4375);
buf BUF1 (N4526, N4518);
or OR3 (N4527, N4526, N1169, N1792);
nor NOR4 (N4528, N4522, N1431, N3981, N4492);
nor NOR4 (N4529, N4515, N2018, N1261, N1338);
nor NOR2 (N4530, N4525, N1612);
buf BUF1 (N4531, N4513);
and AND3 (N4532, N4530, N2003, N982);
not NOT1 (N4533, N4520);
xor XOR2 (N4534, N4501, N3500);
nand NAND2 (N4535, N4534, N763);
nand NAND2 (N4536, N4529, N1462);
nand NAND2 (N4537, N4532, N1847);
buf BUF1 (N4538, N4519);
nor NOR2 (N4539, N4527, N1242);
nor NOR2 (N4540, N4509, N2306);
and AND3 (N4541, N4536, N3693, N2294);
buf BUF1 (N4542, N4541);
buf BUF1 (N4543, N4539);
and AND3 (N4544, N4538, N441, N4380);
or OR2 (N4545, N4533, N2505);
or OR2 (N4546, N4540, N4447);
xor XOR2 (N4547, N4528, N2634);
buf BUF1 (N4548, N4531);
nor NOR2 (N4549, N4524, N2296);
and AND3 (N4550, N4546, N479, N613);
nor NOR4 (N4551, N4537, N1206, N680, N811);
and AND3 (N4552, N4551, N2655, N3247);
not NOT1 (N4553, N4545);
or OR4 (N4554, N4544, N3316, N966, N2196);
buf BUF1 (N4555, N4548);
xor XOR2 (N4556, N4542, N3004);
nor NOR4 (N4557, N4535, N365, N1458, N4425);
not NOT1 (N4558, N4552);
xor XOR2 (N4559, N4543, N2826);
not NOT1 (N4560, N4554);
or OR2 (N4561, N4547, N3432);
buf BUF1 (N4562, N4550);
xor XOR2 (N4563, N4562, N307);
xor XOR2 (N4564, N4559, N35);
nand NAND3 (N4565, N4556, N1046, N3436);
buf BUF1 (N4566, N4560);
nand NAND2 (N4567, N4563, N3118);
not NOT1 (N4568, N4564);
or OR3 (N4569, N4567, N2239, N4519);
xor XOR2 (N4570, N4557, N1863);
or OR2 (N4571, N4568, N1550);
nor NOR2 (N4572, N4571, N598);
or OR4 (N4573, N4569, N3236, N357, N2699);
nor NOR2 (N4574, N4570, N1673);
xor XOR2 (N4575, N4565, N2943);
xor XOR2 (N4576, N4558, N803);
and AND2 (N4577, N4573, N1651);
or OR3 (N4578, N4572, N4424, N1537);
buf BUF1 (N4579, N4553);
and AND4 (N4580, N4579, N4455, N520, N440);
not NOT1 (N4581, N4576);
nand NAND3 (N4582, N4577, N4417, N1059);
and AND4 (N4583, N4582, N565, N3066, N2158);
or OR4 (N4584, N4561, N3654, N3518, N3944);
nand NAND3 (N4585, N4555, N999, N801);
or OR4 (N4586, N4574, N1529, N644, N1663);
nand NAND2 (N4587, N4580, N517);
not NOT1 (N4588, N4586);
nor NOR4 (N4589, N4585, N2745, N1959, N2350);
or OR3 (N4590, N4575, N1727, N4027);
and AND4 (N4591, N4587, N3871, N2898, N3129);
nor NOR2 (N4592, N4578, N2788);
xor XOR2 (N4593, N4584, N1075);
buf BUF1 (N4594, N4591);
buf BUF1 (N4595, N4593);
xor XOR2 (N4596, N4581, N3697);
and AND3 (N4597, N4588, N4548, N3311);
xor XOR2 (N4598, N4594, N1532);
not NOT1 (N4599, N4589);
nor NOR3 (N4600, N4595, N3617, N3564);
xor XOR2 (N4601, N4597, N1339);
nor NOR4 (N4602, N4549, N2456, N1385, N1408);
xor XOR2 (N4603, N4602, N4090);
and AND3 (N4604, N4566, N1401, N4138);
not NOT1 (N4605, N4601);
nor NOR2 (N4606, N4605, N1818);
buf BUF1 (N4607, N4583);
not NOT1 (N4608, N4603);
and AND2 (N4609, N4600, N866);
and AND2 (N4610, N4607, N1917);
xor XOR2 (N4611, N4599, N1006);
or OR3 (N4612, N4610, N1885, N719);
buf BUF1 (N4613, N4598);
xor XOR2 (N4614, N4611, N1277);
xor XOR2 (N4615, N4606, N249);
nand NAND3 (N4616, N4615, N4524, N4003);
buf BUF1 (N4617, N4613);
not NOT1 (N4618, N4617);
buf BUF1 (N4619, N4608);
and AND2 (N4620, N4618, N4289);
nand NAND3 (N4621, N4604, N4051, N748);
nand NAND2 (N4622, N4596, N2988);
buf BUF1 (N4623, N4621);
nand NAND2 (N4624, N4620, N1083);
and AND3 (N4625, N4614, N609, N2426);
or OR2 (N4626, N4624, N2325);
buf BUF1 (N4627, N4623);
not NOT1 (N4628, N4592);
nand NAND2 (N4629, N4626, N2640);
buf BUF1 (N4630, N4622);
and AND2 (N4631, N4628, N2572);
and AND4 (N4632, N4612, N605, N882, N3474);
not NOT1 (N4633, N4619);
buf BUF1 (N4634, N4632);
not NOT1 (N4635, N4633);
or OR3 (N4636, N4627, N4469, N784);
xor XOR2 (N4637, N4634, N2042);
nor NOR4 (N4638, N4636, N4500, N3024, N1400);
nor NOR2 (N4639, N4638, N1808);
and AND3 (N4640, N4629, N3216, N4462);
buf BUF1 (N4641, N4609);
xor XOR2 (N4642, N4630, N2111);
nor NOR2 (N4643, N4590, N2325);
buf BUF1 (N4644, N4637);
xor XOR2 (N4645, N4625, N978);
buf BUF1 (N4646, N4631);
buf BUF1 (N4647, N4616);
nand NAND4 (N4648, N4646, N2392, N3024, N881);
not NOT1 (N4649, N4641);
or OR4 (N4650, N4644, N2490, N1050, N3500);
or OR2 (N4651, N4643, N2751);
or OR2 (N4652, N4651, N1783);
or OR2 (N4653, N4649, N4163);
buf BUF1 (N4654, N4653);
xor XOR2 (N4655, N4647, N3796);
buf BUF1 (N4656, N4645);
or OR4 (N4657, N4656, N1575, N3389, N2463);
or OR4 (N4658, N4639, N3519, N3596, N2928);
nand NAND3 (N4659, N4648, N4420, N4030);
or OR3 (N4660, N4657, N1766, N347);
not NOT1 (N4661, N4650);
or OR2 (N4662, N4640, N3271);
nand NAND4 (N4663, N4652, N2254, N528, N1907);
or OR3 (N4664, N4659, N3292, N1276);
buf BUF1 (N4665, N4658);
or OR3 (N4666, N4642, N3359, N2726);
nand NAND2 (N4667, N4655, N3);
nand NAND2 (N4668, N4663, N392);
nor NOR4 (N4669, N4660, N4396, N97, N718);
nor NOR3 (N4670, N4665, N2909, N1284);
or OR2 (N4671, N4664, N1841);
xor XOR2 (N4672, N4669, N1244);
nor NOR4 (N4673, N4670, N2285, N1602, N1677);
buf BUF1 (N4674, N4635);
nor NOR2 (N4675, N4671, N4417);
nor NOR3 (N4676, N4661, N1423, N3553);
nand NAND4 (N4677, N4666, N4182, N1338, N4634);
xor XOR2 (N4678, N4674, N1317);
and AND4 (N4679, N4678, N358, N936, N522);
xor XOR2 (N4680, N4679, N1099);
or OR4 (N4681, N4676, N3862, N320, N2782);
and AND3 (N4682, N4675, N3541, N2790);
nor NOR3 (N4683, N4668, N673, N70);
and AND3 (N4684, N4654, N4127, N4645);
or OR2 (N4685, N4681, N370);
xor XOR2 (N4686, N4685, N1464);
xor XOR2 (N4687, N4672, N1971);
or OR4 (N4688, N4680, N4273, N2582, N1965);
buf BUF1 (N4689, N4667);
and AND3 (N4690, N4686, N1163, N2352);
not NOT1 (N4691, N4677);
xor XOR2 (N4692, N4689, N1499);
xor XOR2 (N4693, N4687, N3852);
nand NAND3 (N4694, N4693, N1910, N3281);
buf BUF1 (N4695, N4692);
not NOT1 (N4696, N4683);
nor NOR2 (N4697, N4684, N257);
or OR3 (N4698, N4695, N3545, N3359);
buf BUF1 (N4699, N4662);
buf BUF1 (N4700, N4673);
nand NAND3 (N4701, N4699, N840, N60);
nor NOR2 (N4702, N4688, N621);
or OR2 (N4703, N4700, N23);
not NOT1 (N4704, N4694);
and AND2 (N4705, N4697, N49);
and AND3 (N4706, N4702, N3234, N1656);
nand NAND2 (N4707, N4706, N1839);
nand NAND3 (N4708, N4691, N4462, N3105);
xor XOR2 (N4709, N4698, N4688);
nor NOR4 (N4710, N4707, N1786, N2174, N3219);
buf BUF1 (N4711, N4708);
nor NOR3 (N4712, N4703, N4152, N1442);
and AND3 (N4713, N4690, N771, N3151);
nand NAND4 (N4714, N4701, N500, N4217, N25);
buf BUF1 (N4715, N4696);
nand NAND4 (N4716, N4704, N2743, N4496, N4673);
buf BUF1 (N4717, N4711);
and AND3 (N4718, N4714, N393, N3802);
xor XOR2 (N4719, N4717, N963);
nand NAND2 (N4720, N4705, N689);
or OR3 (N4721, N4718, N831, N1591);
or OR4 (N4722, N4720, N1522, N1782, N1418);
not NOT1 (N4723, N4721);
nand NAND3 (N4724, N4719, N1476, N309);
nand NAND2 (N4725, N4722, N2327);
or OR4 (N4726, N4682, N2420, N3174, N2282);
xor XOR2 (N4727, N4712, N1008);
buf BUF1 (N4728, N4724);
or OR4 (N4729, N4710, N236, N1499, N1887);
or OR3 (N4730, N4726, N579, N4680);
not NOT1 (N4731, N4729);
buf BUF1 (N4732, N4709);
nand NAND3 (N4733, N4728, N2261, N4084);
nand NAND4 (N4734, N4715, N3560, N400, N2802);
and AND2 (N4735, N4732, N3557);
buf BUF1 (N4736, N4735);
buf BUF1 (N4737, N4716);
or OR3 (N4738, N4730, N1124, N1682);
nor NOR3 (N4739, N4723, N2082, N466);
not NOT1 (N4740, N4739);
xor XOR2 (N4741, N4713, N1037);
or OR3 (N4742, N4737, N3359, N4094);
nor NOR2 (N4743, N4733, N827);
xor XOR2 (N4744, N4734, N826);
nor NOR4 (N4745, N4744, N2934, N3211, N2090);
buf BUF1 (N4746, N4738);
xor XOR2 (N4747, N4743, N1743);
nor NOR3 (N4748, N4731, N1915, N1453);
nor NOR4 (N4749, N4740, N2724, N3073, N3476);
nand NAND4 (N4750, N4727, N211, N3556, N1172);
or OR2 (N4751, N4749, N552);
and AND4 (N4752, N4747, N18, N2401, N4729);
nand NAND4 (N4753, N4741, N271, N834, N144);
nor NOR4 (N4754, N4725, N852, N441, N2456);
and AND2 (N4755, N4750, N4748);
nor NOR2 (N4756, N3694, N2253);
or OR2 (N4757, N4736, N3562);
not NOT1 (N4758, N4752);
nor NOR4 (N4759, N4755, N2552, N3317, N3094);
nor NOR4 (N4760, N4754, N764, N3510, N3667);
buf BUF1 (N4761, N4746);
and AND3 (N4762, N4756, N843, N1432);
nand NAND2 (N4763, N4742, N4661);
and AND2 (N4764, N4758, N1425);
buf BUF1 (N4765, N4753);
or OR3 (N4766, N4757, N4507, N4334);
buf BUF1 (N4767, N4759);
xor XOR2 (N4768, N4751, N4718);
or OR3 (N4769, N4768, N3644, N1509);
or OR4 (N4770, N4762, N4650, N1029, N342);
not NOT1 (N4771, N4766);
buf BUF1 (N4772, N4770);
buf BUF1 (N4773, N4765);
nand NAND4 (N4774, N4773, N3709, N1059, N2704);
or OR2 (N4775, N4774, N277);
and AND3 (N4776, N4771, N2020, N477);
not NOT1 (N4777, N4776);
buf BUF1 (N4778, N4777);
nor NOR4 (N4779, N4775, N236, N3570, N886);
nor NOR4 (N4780, N4767, N4108, N1701, N4337);
nand NAND3 (N4781, N4778, N2409, N3339);
or OR3 (N4782, N4745, N4530, N2888);
buf BUF1 (N4783, N4780);
nor NOR4 (N4784, N4781, N2687, N4728, N39);
xor XOR2 (N4785, N4772, N2515);
not NOT1 (N4786, N4760);
or OR4 (N4787, N4769, N3664, N934, N1598);
or OR3 (N4788, N4786, N2983, N4479);
and AND4 (N4789, N4783, N752, N409, N4035);
buf BUF1 (N4790, N4763);
nand NAND3 (N4791, N4785, N878, N3057);
xor XOR2 (N4792, N4782, N2372);
nand NAND2 (N4793, N4784, N2725);
nand NAND4 (N4794, N4761, N1544, N2462, N2876);
nand NAND2 (N4795, N4794, N2493);
not NOT1 (N4796, N4788);
xor XOR2 (N4797, N4792, N1);
buf BUF1 (N4798, N4791);
nand NAND2 (N4799, N4795, N3295);
xor XOR2 (N4800, N4790, N4740);
xor XOR2 (N4801, N4798, N4754);
nor NOR2 (N4802, N4800, N3050);
nand NAND4 (N4803, N4789, N2831, N2836, N1842);
not NOT1 (N4804, N4801);
and AND3 (N4805, N4803, N3347, N4551);
xor XOR2 (N4806, N4799, N3567);
xor XOR2 (N4807, N4793, N3910);
buf BUF1 (N4808, N4796);
nor NOR3 (N4809, N4808, N2955, N2079);
or OR4 (N4810, N4764, N440, N2420, N1000);
nand NAND2 (N4811, N4805, N1209);
and AND4 (N4812, N4806, N3639, N1617, N2637);
nand NAND3 (N4813, N4797, N3396, N4076);
nand NAND3 (N4814, N4804, N917, N4709);
nand NAND2 (N4815, N4813, N331);
nand NAND3 (N4816, N4814, N938, N3756);
buf BUF1 (N4817, N4811);
nand NAND4 (N4818, N4812, N2081, N448, N2546);
not NOT1 (N4819, N4802);
nor NOR3 (N4820, N4807, N3456, N109);
or OR2 (N4821, N4818, N3285);
xor XOR2 (N4822, N4810, N364);
xor XOR2 (N4823, N4787, N1481);
buf BUF1 (N4824, N4779);
or OR3 (N4825, N4822, N1753, N3522);
xor XOR2 (N4826, N4815, N958);
or OR2 (N4827, N4817, N2681);
nand NAND4 (N4828, N4824, N1869, N1633, N2522);
or OR3 (N4829, N4826, N3021, N4622);
and AND2 (N4830, N4825, N1968);
and AND3 (N4831, N4816, N4152, N1085);
and AND2 (N4832, N4827, N1220);
not NOT1 (N4833, N4809);
and AND4 (N4834, N4829, N3123, N2700, N3826);
xor XOR2 (N4835, N4820, N3040);
buf BUF1 (N4836, N4835);
nor NOR4 (N4837, N4828, N1016, N3171, N3691);
buf BUF1 (N4838, N4834);
xor XOR2 (N4839, N4823, N4818);
not NOT1 (N4840, N4833);
or OR2 (N4841, N4831, N2853);
xor XOR2 (N4842, N4839, N3512);
xor XOR2 (N4843, N4841, N2008);
buf BUF1 (N4844, N4837);
buf BUF1 (N4845, N4819);
xor XOR2 (N4846, N4842, N2842);
nor NOR2 (N4847, N4838, N704);
buf BUF1 (N4848, N4844);
and AND4 (N4849, N4843, N1806, N813, N2941);
not NOT1 (N4850, N4849);
nor NOR2 (N4851, N4845, N4039);
buf BUF1 (N4852, N4840);
xor XOR2 (N4853, N4852, N4374);
buf BUF1 (N4854, N4830);
not NOT1 (N4855, N4853);
buf BUF1 (N4856, N4854);
nor NOR2 (N4857, N4848, N3221);
and AND2 (N4858, N4851, N2484);
nand NAND2 (N4859, N4836, N1150);
or OR3 (N4860, N4856, N2935, N4431);
nor NOR4 (N4861, N4859, N1603, N2833, N2782);
not NOT1 (N4862, N4855);
not NOT1 (N4863, N4857);
buf BUF1 (N4864, N4821);
not NOT1 (N4865, N4832);
xor XOR2 (N4866, N4858, N3902);
not NOT1 (N4867, N4862);
xor XOR2 (N4868, N4866, N3271);
and AND2 (N4869, N4867, N4271);
not NOT1 (N4870, N4860);
or OR4 (N4871, N4863, N4036, N3119, N1577);
buf BUF1 (N4872, N4870);
nand NAND4 (N4873, N4846, N303, N4483, N629);
xor XOR2 (N4874, N4868, N163);
xor XOR2 (N4875, N4847, N2548);
buf BUF1 (N4876, N4869);
or OR3 (N4877, N4873, N4320, N2081);
nand NAND2 (N4878, N4865, N4009);
and AND3 (N4879, N4861, N3509, N60);
nor NOR4 (N4880, N4876, N3726, N529, N1445);
not NOT1 (N4881, N4879);
nor NOR2 (N4882, N4875, N1257);
nor NOR4 (N4883, N4878, N1706, N460, N2518);
nand NAND3 (N4884, N4881, N376, N2047);
not NOT1 (N4885, N4871);
and AND2 (N4886, N4864, N3651);
nand NAND4 (N4887, N4880, N3637, N474, N484);
buf BUF1 (N4888, N4885);
not NOT1 (N4889, N4884);
xor XOR2 (N4890, N4850, N3731);
not NOT1 (N4891, N4886);
buf BUF1 (N4892, N4889);
or OR2 (N4893, N4887, N2421);
xor XOR2 (N4894, N4890, N2068);
nand NAND2 (N4895, N4892, N2675);
not NOT1 (N4896, N4895);
not NOT1 (N4897, N4891);
nor NOR4 (N4898, N4896, N4034, N3234, N2973);
nand NAND2 (N4899, N4894, N1232);
or OR3 (N4900, N4893, N1297, N236);
buf BUF1 (N4901, N4899);
or OR3 (N4902, N4882, N1227, N1632);
or OR3 (N4903, N4900, N4261, N4087);
or OR3 (N4904, N4903, N2430, N3948);
not NOT1 (N4905, N4898);
nand NAND2 (N4906, N4888, N2504);
nand NAND4 (N4907, N4877, N3060, N4190, N888);
nand NAND2 (N4908, N4902, N4799);
buf BUF1 (N4909, N4908);
and AND3 (N4910, N4909, N4630, N4520);
and AND3 (N4911, N4897, N1796, N485);
or OR2 (N4912, N4906, N3875);
xor XOR2 (N4913, N4883, N832);
and AND3 (N4914, N4913, N1312, N472);
nor NOR4 (N4915, N4901, N1829, N1820, N2404);
buf BUF1 (N4916, N4912);
nor NOR2 (N4917, N4916, N2988);
nor NOR4 (N4918, N4917, N4098, N434, N1988);
nor NOR4 (N4919, N4905, N1013, N651, N4224);
or OR4 (N4920, N4904, N2060, N993, N4876);
buf BUF1 (N4921, N4910);
nor NOR2 (N4922, N4920, N3212);
and AND4 (N4923, N4915, N4003, N1347, N4484);
buf BUF1 (N4924, N4921);
xor XOR2 (N4925, N4911, N1783);
or OR2 (N4926, N4922, N252);
xor XOR2 (N4927, N4919, N2291);
xor XOR2 (N4928, N4874, N986);
not NOT1 (N4929, N4924);
or OR3 (N4930, N4914, N3589, N4016);
or OR4 (N4931, N4925, N1157, N4605, N3752);
not NOT1 (N4932, N4928);
xor XOR2 (N4933, N4931, N85);
xor XOR2 (N4934, N4926, N4603);
or OR2 (N4935, N4872, N2576);
nand NAND4 (N4936, N4930, N2131, N4530, N2847);
buf BUF1 (N4937, N4932);
nor NOR2 (N4938, N4907, N4177);
not NOT1 (N4939, N4933);
and AND4 (N4940, N4918, N1729, N3543, N2548);
nor NOR2 (N4941, N4937, N4659);
or OR4 (N4942, N4934, N2629, N3985, N4565);
buf BUF1 (N4943, N4942);
not NOT1 (N4944, N4940);
or OR3 (N4945, N4927, N4029, N4103);
buf BUF1 (N4946, N4929);
or OR3 (N4947, N4938, N2253, N4886);
not NOT1 (N4948, N4935);
xor XOR2 (N4949, N4946, N1930);
nand NAND3 (N4950, N4948, N3374, N4033);
xor XOR2 (N4951, N4943, N2500);
and AND2 (N4952, N4947, N3494);
nand NAND2 (N4953, N4936, N4738);
buf BUF1 (N4954, N4953);
or OR3 (N4955, N4951, N4209, N317);
and AND2 (N4956, N4923, N4313);
or OR2 (N4957, N4941, N1385);
nor NOR3 (N4958, N4955, N4644, N1416);
not NOT1 (N4959, N4952);
buf BUF1 (N4960, N4950);
xor XOR2 (N4961, N4957, N3228);
or OR2 (N4962, N4945, N2440);
not NOT1 (N4963, N4949);
or OR4 (N4964, N4939, N258, N2928, N608);
or OR2 (N4965, N4962, N3037);
buf BUF1 (N4966, N4954);
buf BUF1 (N4967, N4963);
buf BUF1 (N4968, N4965);
nand NAND2 (N4969, N4959, N3164);
nor NOR2 (N4970, N4958, N3250);
or OR3 (N4971, N4961, N3654, N65);
nor NOR4 (N4972, N4971, N269, N4040, N2118);
nand NAND2 (N4973, N4960, N2499);
nor NOR3 (N4974, N4972, N302, N4271);
or OR3 (N4975, N4969, N945, N1470);
or OR4 (N4976, N4956, N2205, N3427, N200);
nor NOR2 (N4977, N4944, N2018);
not NOT1 (N4978, N4967);
or OR2 (N4979, N4976, N617);
nor NOR4 (N4980, N4966, N903, N3426, N1990);
buf BUF1 (N4981, N4970);
nor NOR3 (N4982, N4975, N576, N355);
and AND2 (N4983, N4980, N3563);
nor NOR3 (N4984, N4983, N788, N3447);
nand NAND4 (N4985, N4964, N696, N4353, N925);
not NOT1 (N4986, N4968);
or OR2 (N4987, N4979, N2293);
nand NAND2 (N4988, N4978, N2595);
nor NOR2 (N4989, N4977, N3833);
nor NOR3 (N4990, N4987, N1281, N1443);
xor XOR2 (N4991, N4986, N185);
and AND2 (N4992, N4973, N804);
not NOT1 (N4993, N4984);
not NOT1 (N4994, N4982);
nor NOR4 (N4995, N4992, N1420, N2867, N4576);
or OR2 (N4996, N4993, N3945);
xor XOR2 (N4997, N4988, N3245);
or OR3 (N4998, N4997, N1487, N1071);
not NOT1 (N4999, N4989);
not NOT1 (N5000, N4981);
not NOT1 (N5001, N4990);
and AND4 (N5002, N4998, N1056, N4572, N778);
buf BUF1 (N5003, N4994);
buf BUF1 (N5004, N5000);
nand NAND4 (N5005, N4985, N3361, N3678, N4536);
buf BUF1 (N5006, N4974);
and AND3 (N5007, N5006, N4316, N3797);
or OR2 (N5008, N4999, N4084);
nand NAND4 (N5009, N5001, N2025, N4735, N1299);
xor XOR2 (N5010, N5005, N2266);
nand NAND4 (N5011, N5007, N1849, N525, N4952);
and AND4 (N5012, N5008, N633, N749, N1929);
not NOT1 (N5013, N4995);
xor XOR2 (N5014, N5010, N4476);
and AND2 (N5015, N5002, N588);
nand NAND2 (N5016, N4996, N740);
nor NOR4 (N5017, N5004, N969, N158, N773);
buf BUF1 (N5018, N5009);
not NOT1 (N5019, N5013);
buf BUF1 (N5020, N5016);
nor NOR2 (N5021, N5015, N3489);
or OR2 (N5022, N5011, N3572);
and AND3 (N5023, N5012, N1431, N1141);
not NOT1 (N5024, N5019);
and AND3 (N5025, N5021, N1156, N2967);
or OR2 (N5026, N5020, N825);
and AND2 (N5027, N5014, N4790);
or OR3 (N5028, N5027, N2974, N4839);
not NOT1 (N5029, N5003);
nor NOR4 (N5030, N5018, N4056, N1531, N544);
and AND4 (N5031, N5023, N273, N656, N1567);
xor XOR2 (N5032, N5028, N4084);
or OR4 (N5033, N5032, N89, N3317, N4066);
nand NAND3 (N5034, N5031, N986, N2727);
xor XOR2 (N5035, N5022, N77);
nor NOR3 (N5036, N5034, N1901, N785);
not NOT1 (N5037, N5030);
xor XOR2 (N5038, N5035, N2212);
nand NAND3 (N5039, N5036, N2111, N4911);
and AND4 (N5040, N5039, N1606, N225, N723);
nand NAND2 (N5041, N5025, N822);
or OR3 (N5042, N5041, N2140, N3166);
and AND4 (N5043, N4991, N2352, N846, N3253);
and AND2 (N5044, N5038, N3683);
and AND4 (N5045, N5017, N475, N1815, N705);
and AND3 (N5046, N5044, N386, N1212);
not NOT1 (N5047, N5026);
nor NOR2 (N5048, N5033, N3828);
not NOT1 (N5049, N5048);
nor NOR3 (N5050, N5046, N4860, N1209);
and AND3 (N5051, N5042, N3204, N1355);
nor NOR4 (N5052, N5040, N3531, N4313, N3629);
or OR4 (N5053, N5029, N3261, N3799, N2380);
nand NAND4 (N5054, N5052, N2315, N505, N1743);
and AND4 (N5055, N5024, N2598, N3062, N5014);
not NOT1 (N5056, N5045);
nand NAND2 (N5057, N5053, N3163);
nand NAND3 (N5058, N5056, N1032, N3916);
not NOT1 (N5059, N5050);
not NOT1 (N5060, N5059);
nand NAND3 (N5061, N5055, N1254, N3912);
nand NAND4 (N5062, N5037, N4543, N1488, N3012);
nor NOR3 (N5063, N5051, N1926, N810);
xor XOR2 (N5064, N5060, N2347);
xor XOR2 (N5065, N5047, N2979);
nand NAND4 (N5066, N5062, N3888, N3574, N1210);
not NOT1 (N5067, N5066);
nand NAND4 (N5068, N5043, N4805, N1764, N1900);
nor NOR3 (N5069, N5049, N4901, N1030);
and AND3 (N5070, N5068, N4475, N4384);
xor XOR2 (N5071, N5058, N4205);
and AND2 (N5072, N5065, N960);
and AND4 (N5073, N5064, N3316, N3030, N1676);
not NOT1 (N5074, N5057);
or OR2 (N5075, N5061, N4807);
not NOT1 (N5076, N5069);
or OR2 (N5077, N5070, N1650);
and AND4 (N5078, N5054, N4171, N2299, N4741);
and AND2 (N5079, N5073, N237);
buf BUF1 (N5080, N5071);
nand NAND4 (N5081, N5063, N4440, N386, N93);
and AND3 (N5082, N5076, N3451, N1613);
nor NOR2 (N5083, N5079, N4084);
and AND3 (N5084, N5081, N1055, N3885);
buf BUF1 (N5085, N5067);
not NOT1 (N5086, N5072);
nor NOR3 (N5087, N5077, N1934, N2612);
xor XOR2 (N5088, N5075, N4752);
nand NAND3 (N5089, N5086, N3324, N1766);
nand NAND2 (N5090, N5085, N6);
xor XOR2 (N5091, N5089, N3525);
nor NOR2 (N5092, N5082, N4193);
xor XOR2 (N5093, N5092, N440);
nand NAND4 (N5094, N5087, N80, N669, N1211);
and AND3 (N5095, N5083, N2607, N3468);
xor XOR2 (N5096, N5078, N3995);
or OR2 (N5097, N5095, N1601);
buf BUF1 (N5098, N5080);
nor NOR3 (N5099, N5098, N3862, N4598);
and AND2 (N5100, N5074, N2599);
xor XOR2 (N5101, N5088, N2366);
not NOT1 (N5102, N5097);
not NOT1 (N5103, N5093);
xor XOR2 (N5104, N5094, N4638);
nor NOR4 (N5105, N5102, N2239, N2254, N3158);
or OR3 (N5106, N5103, N1574, N390);
buf BUF1 (N5107, N5084);
or OR4 (N5108, N5100, N3522, N2043, N4062);
not NOT1 (N5109, N5096);
nand NAND2 (N5110, N5107, N2182);
not NOT1 (N5111, N5110);
not NOT1 (N5112, N5109);
not NOT1 (N5113, N5090);
xor XOR2 (N5114, N5101, N327);
xor XOR2 (N5115, N5114, N2491);
xor XOR2 (N5116, N5115, N3467);
and AND2 (N5117, N5116, N3295);
buf BUF1 (N5118, N5108);
not NOT1 (N5119, N5105);
nand NAND3 (N5120, N5112, N3560, N4967);
and AND3 (N5121, N5113, N2937, N752);
xor XOR2 (N5122, N5120, N3384);
nor NOR2 (N5123, N5106, N1090);
not NOT1 (N5124, N5121);
and AND3 (N5125, N5122, N4662, N2401);
buf BUF1 (N5126, N5099);
nand NAND2 (N5127, N5124, N3043);
nor NOR2 (N5128, N5118, N1942);
xor XOR2 (N5129, N5119, N5008);
not NOT1 (N5130, N5126);
and AND2 (N5131, N5104, N922);
or OR4 (N5132, N5123, N314, N2356, N3252);
nor NOR3 (N5133, N5091, N3763, N2071);
and AND2 (N5134, N5125, N917);
xor XOR2 (N5135, N5131, N665);
or OR3 (N5136, N5128, N972, N3667);
nor NOR2 (N5137, N5134, N84);
xor XOR2 (N5138, N5137, N2715);
and AND4 (N5139, N5129, N4128, N2222, N3925);
or OR2 (N5140, N5135, N4524);
or OR2 (N5141, N5133, N5092);
and AND3 (N5142, N5130, N4725, N323);
and AND2 (N5143, N5138, N4603);
not NOT1 (N5144, N5136);
buf BUF1 (N5145, N5143);
nor NOR4 (N5146, N5144, N1818, N3359, N1036);
nand NAND3 (N5147, N5111, N901, N735);
and AND4 (N5148, N5142, N3523, N2815, N2760);
buf BUF1 (N5149, N5145);
or OR2 (N5150, N5139, N2615);
nand NAND3 (N5151, N5146, N2021, N3300);
or OR2 (N5152, N5151, N2939);
nor NOR2 (N5153, N5141, N1540);
not NOT1 (N5154, N5127);
buf BUF1 (N5155, N5147);
nand NAND4 (N5156, N5153, N3278, N2152, N2228);
xor XOR2 (N5157, N5117, N3292);
nand NAND2 (N5158, N5155, N4723);
buf BUF1 (N5159, N5149);
nand NAND4 (N5160, N5157, N4146, N5085, N1656);
nand NAND3 (N5161, N5158, N4049, N4837);
or OR3 (N5162, N5159, N2388, N751);
buf BUF1 (N5163, N5156);
not NOT1 (N5164, N5152);
xor XOR2 (N5165, N5163, N3429);
and AND4 (N5166, N5132, N2129, N5102, N1541);
nor NOR3 (N5167, N5154, N5151, N3153);
xor XOR2 (N5168, N5162, N4266);
nor NOR2 (N5169, N5140, N494);
nor NOR2 (N5170, N5161, N3952);
xor XOR2 (N5171, N5160, N891);
buf BUF1 (N5172, N5166);
nand NAND2 (N5173, N5170, N1440);
nand NAND4 (N5174, N5169, N3235, N1915, N4733);
xor XOR2 (N5175, N5171, N252);
and AND4 (N5176, N5148, N4500, N2781, N2410);
nand NAND4 (N5177, N5164, N1887, N3232, N3132);
nand NAND3 (N5178, N5150, N437, N3043);
nor NOR2 (N5179, N5176, N5127);
or OR4 (N5180, N5165, N2116, N1288, N3469);
nand NAND4 (N5181, N5175, N4389, N3354, N2115);
not NOT1 (N5182, N5180);
buf BUF1 (N5183, N5179);
or OR2 (N5184, N5174, N4991);
xor XOR2 (N5185, N5181, N2883);
xor XOR2 (N5186, N5172, N1478);
nand NAND3 (N5187, N5177, N1741, N2129);
nor NOR2 (N5188, N5183, N1508);
not NOT1 (N5189, N5188);
xor XOR2 (N5190, N5187, N2604);
and AND3 (N5191, N5182, N246, N890);
xor XOR2 (N5192, N5184, N1736);
and AND2 (N5193, N5189, N3789);
xor XOR2 (N5194, N5167, N634);
nand NAND4 (N5195, N5193, N3087, N307, N2042);
nor NOR2 (N5196, N5192, N4653);
nand NAND4 (N5197, N5194, N1456, N5082, N3444);
or OR2 (N5198, N5168, N2702);
nand NAND3 (N5199, N5178, N555, N649);
and AND2 (N5200, N5197, N1488);
nand NAND2 (N5201, N5200, N3228);
and AND4 (N5202, N5196, N2716, N1438, N4143);
and AND3 (N5203, N5195, N1180, N2765);
buf BUF1 (N5204, N5202);
nor NOR3 (N5205, N5190, N4107, N874);
xor XOR2 (N5206, N5191, N1051);
or OR3 (N5207, N5201, N475, N1815);
nor NOR2 (N5208, N5173, N2667);
buf BUF1 (N5209, N5204);
not NOT1 (N5210, N5199);
buf BUF1 (N5211, N5186);
xor XOR2 (N5212, N5208, N1604);
xor XOR2 (N5213, N5207, N3935);
or OR3 (N5214, N5211, N2449, N3895);
buf BUF1 (N5215, N5198);
not NOT1 (N5216, N5213);
nor NOR3 (N5217, N5185, N3715, N5039);
or OR3 (N5218, N5203, N4152, N3764);
xor XOR2 (N5219, N5218, N458);
and AND2 (N5220, N5215, N4432);
or OR3 (N5221, N5219, N3531, N1765);
xor XOR2 (N5222, N5210, N2572);
buf BUF1 (N5223, N5217);
buf BUF1 (N5224, N5205);
or OR2 (N5225, N5223, N2653);
xor XOR2 (N5226, N5225, N5216);
nand NAND4 (N5227, N731, N2434, N257, N1254);
nor NOR2 (N5228, N5221, N4516);
buf BUF1 (N5229, N5224);
not NOT1 (N5230, N5227);
nand NAND3 (N5231, N5222, N4502, N2772);
nand NAND2 (N5232, N5226, N2691);
nor NOR2 (N5233, N5212, N1164);
nor NOR3 (N5234, N5233, N120, N749);
or OR3 (N5235, N5232, N3071, N4707);
nand NAND2 (N5236, N5234, N2514);
not NOT1 (N5237, N5206);
nor NOR4 (N5238, N5229, N2454, N2785, N4887);
nor NOR4 (N5239, N5220, N1237, N1073, N991);
xor XOR2 (N5240, N5236, N468);
and AND4 (N5241, N5237, N1500, N216, N4371);
or OR4 (N5242, N5230, N990, N2991, N1128);
nor NOR3 (N5243, N5241, N815, N1162);
or OR2 (N5244, N5214, N1905);
not NOT1 (N5245, N5243);
nand NAND4 (N5246, N5244, N86, N526, N1899);
nor NOR4 (N5247, N5246, N1617, N3309, N4501);
or OR3 (N5248, N5238, N1442, N903);
or OR3 (N5249, N5245, N2078, N5084);
xor XOR2 (N5250, N5239, N4221);
nor NOR4 (N5251, N5248, N298, N1493, N2562);
buf BUF1 (N5252, N5242);
and AND2 (N5253, N5228, N3780);
and AND2 (N5254, N5240, N2077);
not NOT1 (N5255, N5209);
or OR2 (N5256, N5235, N61);
not NOT1 (N5257, N5247);
not NOT1 (N5258, N5256);
and AND3 (N5259, N5255, N4259, N317);
or OR3 (N5260, N5258, N5056, N4160);
not NOT1 (N5261, N5249);
not NOT1 (N5262, N5252);
buf BUF1 (N5263, N5250);
not NOT1 (N5264, N5231);
nor NOR3 (N5265, N5259, N182, N4055);
xor XOR2 (N5266, N5253, N3738);
nand NAND2 (N5267, N5261, N3905);
and AND2 (N5268, N5251, N3938);
buf BUF1 (N5269, N5257);
nand NAND2 (N5270, N5265, N4270);
not NOT1 (N5271, N5270);
nand NAND4 (N5272, N5263, N299, N1183, N3030);
buf BUF1 (N5273, N5254);
or OR3 (N5274, N5266, N3322, N4345);
not NOT1 (N5275, N5262);
not NOT1 (N5276, N5268);
buf BUF1 (N5277, N5274);
and AND3 (N5278, N5260, N4760, N279);
nor NOR4 (N5279, N5269, N3047, N4121, N3565);
nand NAND2 (N5280, N5275, N4620);
not NOT1 (N5281, N5280);
or OR4 (N5282, N5273, N3768, N3881, N1174);
nand NAND3 (N5283, N5276, N801, N4655);
and AND2 (N5284, N5281, N3935);
xor XOR2 (N5285, N5282, N198);
and AND3 (N5286, N5279, N929, N356);
buf BUF1 (N5287, N5283);
not NOT1 (N5288, N5267);
and AND3 (N5289, N5286, N1810, N3486);
not NOT1 (N5290, N5272);
not NOT1 (N5291, N5271);
nor NOR4 (N5292, N5264, N2631, N3729, N4260);
xor XOR2 (N5293, N5285, N651);
or OR4 (N5294, N5289, N4777, N3937, N586);
xor XOR2 (N5295, N5284, N3936);
xor XOR2 (N5296, N5295, N4107);
nand NAND4 (N5297, N5292, N2956, N3143, N746);
nand NAND4 (N5298, N5294, N1372, N4824, N3213);
nand NAND2 (N5299, N5297, N4845);
not NOT1 (N5300, N5293);
or OR3 (N5301, N5278, N649, N1835);
nand NAND2 (N5302, N5300, N1160);
buf BUF1 (N5303, N5302);
xor XOR2 (N5304, N5299, N146);
not NOT1 (N5305, N5287);
xor XOR2 (N5306, N5298, N827);
buf BUF1 (N5307, N5291);
nor NOR2 (N5308, N5301, N2901);
not NOT1 (N5309, N5296);
not NOT1 (N5310, N5305);
nand NAND3 (N5311, N5288, N1029, N1645);
buf BUF1 (N5312, N5308);
buf BUF1 (N5313, N5306);
buf BUF1 (N5314, N5309);
buf BUF1 (N5315, N5303);
xor XOR2 (N5316, N5290, N68);
buf BUF1 (N5317, N5315);
or OR2 (N5318, N5316, N3573);
nand NAND3 (N5319, N5312, N3179, N3595);
buf BUF1 (N5320, N5319);
or OR2 (N5321, N5320, N3250);
xor XOR2 (N5322, N5310, N1239);
not NOT1 (N5323, N5311);
not NOT1 (N5324, N5317);
nor NOR2 (N5325, N5314, N470);
not NOT1 (N5326, N5277);
not NOT1 (N5327, N5325);
and AND4 (N5328, N5321, N3515, N2809, N3687);
xor XOR2 (N5329, N5326, N1309);
buf BUF1 (N5330, N5322);
buf BUF1 (N5331, N5327);
nand NAND2 (N5332, N5331, N5006);
nor NOR3 (N5333, N5318, N3554, N4920);
buf BUF1 (N5334, N5323);
buf BUF1 (N5335, N5334);
nand NAND4 (N5336, N5307, N3466, N2307, N4859);
or OR4 (N5337, N5329, N2989, N3258, N5021);
not NOT1 (N5338, N5324);
or OR2 (N5339, N5333, N1114);
or OR2 (N5340, N5339, N2858);
or OR3 (N5341, N5330, N770, N3242);
xor XOR2 (N5342, N5336, N2311);
xor XOR2 (N5343, N5341, N2279);
buf BUF1 (N5344, N5340);
xor XOR2 (N5345, N5304, N3164);
nor NOR3 (N5346, N5338, N3419, N3065);
and AND2 (N5347, N5344, N4157);
nand NAND3 (N5348, N5345, N826, N3782);
and AND4 (N5349, N5313, N1296, N3245, N2680);
nor NOR2 (N5350, N5346, N4832);
nand NAND2 (N5351, N5347, N295);
and AND2 (N5352, N5343, N1078);
and AND4 (N5353, N5328, N5190, N1592, N1169);
nor NOR4 (N5354, N5352, N3937, N2764, N379);
not NOT1 (N5355, N5351);
nand NAND3 (N5356, N5349, N739, N301);
xor XOR2 (N5357, N5335, N3943);
or OR4 (N5358, N5353, N3065, N2467, N3302);
or OR2 (N5359, N5354, N3902);
and AND2 (N5360, N5348, N3855);
buf BUF1 (N5361, N5359);
not NOT1 (N5362, N5360);
nand NAND3 (N5363, N5357, N362, N864);
nand NAND4 (N5364, N5332, N3359, N1369, N1459);
or OR4 (N5365, N5356, N1758, N2291, N355);
and AND2 (N5366, N5355, N4043);
nor NOR4 (N5367, N5366, N2730, N19, N1032);
not NOT1 (N5368, N5362);
nor NOR3 (N5369, N5361, N2464, N3949);
or OR3 (N5370, N5350, N2913, N1409);
xor XOR2 (N5371, N5342, N1882);
not NOT1 (N5372, N5370);
and AND2 (N5373, N5367, N412);
or OR2 (N5374, N5363, N4076);
not NOT1 (N5375, N5371);
nor NOR3 (N5376, N5337, N867, N679);
and AND2 (N5377, N5364, N280);
buf BUF1 (N5378, N5375);
xor XOR2 (N5379, N5374, N219);
xor XOR2 (N5380, N5378, N1257);
and AND4 (N5381, N5365, N2001, N3556, N4708);
nor NOR2 (N5382, N5377, N2558);
xor XOR2 (N5383, N5381, N674);
nor NOR4 (N5384, N5372, N2718, N2264, N4386);
or OR4 (N5385, N5384, N699, N2775, N4082);
nand NAND2 (N5386, N5373, N4030);
buf BUF1 (N5387, N5386);
xor XOR2 (N5388, N5385, N2261);
buf BUF1 (N5389, N5388);
nand NAND3 (N5390, N5379, N2584, N1696);
buf BUF1 (N5391, N5390);
nand NAND2 (N5392, N5382, N3482);
not NOT1 (N5393, N5369);
not NOT1 (N5394, N5380);
xor XOR2 (N5395, N5393, N5134);
and AND4 (N5396, N5383, N1471, N4420, N2055);
xor XOR2 (N5397, N5368, N1346);
not NOT1 (N5398, N5394);
xor XOR2 (N5399, N5376, N1656);
not NOT1 (N5400, N5389);
not NOT1 (N5401, N5395);
xor XOR2 (N5402, N5387, N2407);
xor XOR2 (N5403, N5402, N2469);
nand NAND3 (N5404, N5399, N2270, N3321);
or OR4 (N5405, N5397, N1320, N3432, N1821);
xor XOR2 (N5406, N5391, N4607);
xor XOR2 (N5407, N5398, N5044);
nand NAND4 (N5408, N5405, N2680, N3768, N5186);
xor XOR2 (N5409, N5407, N1453);
and AND2 (N5410, N5358, N5398);
xor XOR2 (N5411, N5409, N527);
nor NOR2 (N5412, N5400, N3801);
buf BUF1 (N5413, N5392);
or OR4 (N5414, N5410, N704, N1065, N3499);
or OR3 (N5415, N5401, N4843, N2553);
nor NOR4 (N5416, N5415, N1100, N58, N1632);
not NOT1 (N5417, N5414);
xor XOR2 (N5418, N5416, N2166);
and AND3 (N5419, N5413, N1220, N2262);
and AND3 (N5420, N5404, N3847, N3794);
and AND2 (N5421, N5408, N4045);
or OR4 (N5422, N5411, N1601, N2582, N4076);
not NOT1 (N5423, N5412);
nand NAND4 (N5424, N5420, N4206, N1276, N3957);
nand NAND4 (N5425, N5406, N1386, N2345, N3285);
not NOT1 (N5426, N5419);
not NOT1 (N5427, N5396);
xor XOR2 (N5428, N5421, N3387);
or OR4 (N5429, N5424, N3116, N797, N1087);
xor XOR2 (N5430, N5426, N3511);
nor NOR3 (N5431, N5417, N4745, N2079);
buf BUF1 (N5432, N5428);
nor NOR2 (N5433, N5430, N4972);
or OR4 (N5434, N5427, N4247, N3180, N5284);
xor XOR2 (N5435, N5418, N4152);
buf BUF1 (N5436, N5431);
xor XOR2 (N5437, N5423, N1448);
or OR3 (N5438, N5429, N381, N4701);
xor XOR2 (N5439, N5432, N441);
buf BUF1 (N5440, N5433);
nor NOR4 (N5441, N5437, N1248, N4616, N4644);
nand NAND3 (N5442, N5435, N2773, N2009);
nand NAND2 (N5443, N5441, N931);
buf BUF1 (N5444, N5438);
nand NAND4 (N5445, N5439, N1438, N143, N4238);
nand NAND2 (N5446, N5434, N1716);
or OR2 (N5447, N5445, N1681);
or OR4 (N5448, N5443, N1587, N1845, N3048);
not NOT1 (N5449, N5444);
nor NOR2 (N5450, N5446, N358);
buf BUF1 (N5451, N5449);
nor NOR4 (N5452, N5425, N3495, N517, N5203);
not NOT1 (N5453, N5451);
xor XOR2 (N5454, N5422, N5171);
or OR4 (N5455, N5447, N685, N2171, N2309);
not NOT1 (N5456, N5442);
buf BUF1 (N5457, N5456);
nor NOR2 (N5458, N5450, N5318);
xor XOR2 (N5459, N5403, N2960);
nor NOR4 (N5460, N5436, N4451, N2035, N60);
not NOT1 (N5461, N5460);
xor XOR2 (N5462, N5452, N5370);
xor XOR2 (N5463, N5459, N190);
and AND2 (N5464, N5453, N3171);
not NOT1 (N5465, N5464);
nand NAND2 (N5466, N5440, N1829);
xor XOR2 (N5467, N5463, N1758);
xor XOR2 (N5468, N5467, N1350);
nand NAND2 (N5469, N5458, N3557);
not NOT1 (N5470, N5462);
buf BUF1 (N5471, N5448);
nor NOR3 (N5472, N5471, N1970, N2872);
not NOT1 (N5473, N5455);
not NOT1 (N5474, N5457);
and AND2 (N5475, N5472, N1636);
buf BUF1 (N5476, N5465);
and AND2 (N5477, N5476, N1440);
buf BUF1 (N5478, N5470);
or OR2 (N5479, N5468, N1581);
nor NOR3 (N5480, N5469, N3818, N2073);
not NOT1 (N5481, N5475);
buf BUF1 (N5482, N5481);
not NOT1 (N5483, N5479);
and AND2 (N5484, N5473, N3676);
xor XOR2 (N5485, N5461, N2272);
not NOT1 (N5486, N5484);
buf BUF1 (N5487, N5482);
not NOT1 (N5488, N5454);
xor XOR2 (N5489, N5466, N5406);
xor XOR2 (N5490, N5488, N1613);
buf BUF1 (N5491, N5477);
nand NAND4 (N5492, N5474, N2214, N266, N4857);
not NOT1 (N5493, N5480);
not NOT1 (N5494, N5489);
buf BUF1 (N5495, N5490);
and AND4 (N5496, N5493, N4028, N4894, N2679);
and AND2 (N5497, N5485, N341);
buf BUF1 (N5498, N5492);
not NOT1 (N5499, N5486);
not NOT1 (N5500, N5491);
buf BUF1 (N5501, N5496);
nor NOR4 (N5502, N5487, N4326, N4548, N3436);
xor XOR2 (N5503, N5497, N451);
nand NAND4 (N5504, N5495, N4759, N2794, N1145);
buf BUF1 (N5505, N5501);
nand NAND3 (N5506, N5503, N2541, N731);
xor XOR2 (N5507, N5502, N4264);
not NOT1 (N5508, N5504);
nor NOR4 (N5509, N5478, N543, N1007, N635);
buf BUF1 (N5510, N5498);
nor NOR2 (N5511, N5508, N851);
buf BUF1 (N5512, N5507);
not NOT1 (N5513, N5483);
nand NAND2 (N5514, N5505, N4603);
or OR3 (N5515, N5510, N2530, N2648);
or OR4 (N5516, N5506, N2099, N688, N595);
xor XOR2 (N5517, N5509, N4578);
buf BUF1 (N5518, N5516);
or OR2 (N5519, N5494, N2666);
nand NAND2 (N5520, N5511, N5152);
nor NOR3 (N5521, N5512, N3641, N5254);
not NOT1 (N5522, N5515);
nor NOR4 (N5523, N5518, N4559, N2235, N3609);
nand NAND2 (N5524, N5522, N1537);
buf BUF1 (N5525, N5513);
xor XOR2 (N5526, N5521, N3234);
xor XOR2 (N5527, N5525, N1309);
nor NOR4 (N5528, N5499, N2493, N133, N113);
nand NAND2 (N5529, N5528, N3089);
buf BUF1 (N5530, N5526);
or OR2 (N5531, N5520, N2038);
xor XOR2 (N5532, N5527, N4554);
nor NOR3 (N5533, N5514, N2519, N3899);
or OR4 (N5534, N5532, N2200, N5155, N35);
buf BUF1 (N5535, N5519);
nor NOR4 (N5536, N5500, N2115, N5125, N4533);
nor NOR2 (N5537, N5531, N1874);
or OR3 (N5538, N5534, N1365, N1106);
or OR3 (N5539, N5538, N879, N4543);
or OR4 (N5540, N5523, N3681, N1536, N3684);
nor NOR4 (N5541, N5530, N3682, N3905, N4805);
or OR2 (N5542, N5540, N4507);
nor NOR3 (N5543, N5535, N4307, N1967);
nor NOR3 (N5544, N5542, N1376, N5384);
or OR3 (N5545, N5517, N2803, N2449);
not NOT1 (N5546, N5533);
not NOT1 (N5547, N5524);
nor NOR4 (N5548, N5537, N1200, N2442, N5367);
xor XOR2 (N5549, N5536, N4853);
nand NAND4 (N5550, N5545, N1598, N2997, N4675);
xor XOR2 (N5551, N5529, N2944);
nor NOR3 (N5552, N5550, N824, N4735);
buf BUF1 (N5553, N5539);
not NOT1 (N5554, N5547);
or OR4 (N5555, N5546, N963, N1392, N4150);
xor XOR2 (N5556, N5554, N1630);
and AND3 (N5557, N5541, N4698, N498);
not NOT1 (N5558, N5543);
or OR2 (N5559, N5553, N3734);
not NOT1 (N5560, N5552);
nand NAND2 (N5561, N5556, N422);
xor XOR2 (N5562, N5555, N1658);
nand NAND2 (N5563, N5562, N3924);
nor NOR4 (N5564, N5544, N3491, N1271, N5319);
xor XOR2 (N5565, N5549, N2510);
not NOT1 (N5566, N5564);
buf BUF1 (N5567, N5563);
xor XOR2 (N5568, N5551, N1331);
or OR2 (N5569, N5567, N1428);
buf BUF1 (N5570, N5559);
xor XOR2 (N5571, N5561, N2709);
or OR4 (N5572, N5558, N433, N3371, N1615);
xor XOR2 (N5573, N5565, N1634);
nor NOR2 (N5574, N5569, N4563);
or OR4 (N5575, N5560, N5426, N1403, N1127);
and AND3 (N5576, N5575, N4028, N2312);
and AND3 (N5577, N5574, N2246, N3164);
nand NAND3 (N5578, N5573, N2321, N1063);
nand NAND4 (N5579, N5576, N1837, N1017, N5157);
nand NAND3 (N5580, N5579, N4264, N4186);
nand NAND3 (N5581, N5572, N3004, N5299);
xor XOR2 (N5582, N5557, N753);
or OR4 (N5583, N5580, N3306, N1634, N3212);
nand NAND2 (N5584, N5571, N3190);
and AND2 (N5585, N5578, N5174);
nor NOR3 (N5586, N5577, N3376, N3756);
nand NAND2 (N5587, N5581, N4025);
and AND3 (N5588, N5585, N1119, N5300);
buf BUF1 (N5589, N5588);
or OR2 (N5590, N5583, N2338);
or OR2 (N5591, N5566, N4892);
xor XOR2 (N5592, N5587, N4378);
or OR2 (N5593, N5582, N1419);
nand NAND2 (N5594, N5548, N2253);
xor XOR2 (N5595, N5592, N2616);
xor XOR2 (N5596, N5584, N2021);
or OR4 (N5597, N5570, N1811, N3000, N4024);
buf BUF1 (N5598, N5597);
not NOT1 (N5599, N5590);
nand NAND3 (N5600, N5586, N2298, N5429);
nand NAND4 (N5601, N5599, N5011, N3346, N3972);
nand NAND2 (N5602, N5594, N4183);
or OR2 (N5603, N5595, N4305);
nand NAND4 (N5604, N5593, N862, N5122, N1553);
or OR2 (N5605, N5596, N2764);
and AND4 (N5606, N5604, N2781, N3689, N1370);
and AND3 (N5607, N5600, N1167, N5138);
or OR4 (N5608, N5601, N5297, N2061, N5583);
not NOT1 (N5609, N5602);
not NOT1 (N5610, N5568);
and AND3 (N5611, N5605, N3854, N2210);
and AND4 (N5612, N5608, N2366, N501, N836);
xor XOR2 (N5613, N5609, N697);
and AND3 (N5614, N5606, N2725, N2312);
and AND3 (N5615, N5611, N463, N1141);
not NOT1 (N5616, N5615);
not NOT1 (N5617, N5610);
nor NOR4 (N5618, N5617, N4194, N4246, N973);
nand NAND3 (N5619, N5614, N383, N3842);
not NOT1 (N5620, N5607);
not NOT1 (N5621, N5616);
not NOT1 (N5622, N5603);
or OR2 (N5623, N5598, N812);
buf BUF1 (N5624, N5589);
nand NAND4 (N5625, N5618, N5385, N3300, N3073);
buf BUF1 (N5626, N5613);
not NOT1 (N5627, N5622);
or OR2 (N5628, N5591, N4808);
and AND2 (N5629, N5619, N227);
and AND4 (N5630, N5626, N3840, N513, N1598);
buf BUF1 (N5631, N5628);
or OR2 (N5632, N5612, N1908);
not NOT1 (N5633, N5632);
or OR4 (N5634, N5623, N1896, N5462, N2995);
not NOT1 (N5635, N5629);
buf BUF1 (N5636, N5634);
buf BUF1 (N5637, N5635);
nand NAND4 (N5638, N5627, N2833, N3064, N1329);
xor XOR2 (N5639, N5625, N4300);
nand NAND3 (N5640, N5633, N379, N188);
nor NOR4 (N5641, N5636, N881, N500, N472);
or OR3 (N5642, N5621, N356, N5572);
not NOT1 (N5643, N5624);
nor NOR2 (N5644, N5630, N126);
not NOT1 (N5645, N5640);
or OR3 (N5646, N5643, N4938, N244);
and AND4 (N5647, N5637, N3168, N2950, N1860);
nand NAND3 (N5648, N5647, N166, N2967);
buf BUF1 (N5649, N5620);
nand NAND3 (N5650, N5639, N4529, N4910);
nand NAND2 (N5651, N5648, N3705);
not NOT1 (N5652, N5646);
or OR4 (N5653, N5644, N4412, N1593, N235);
or OR4 (N5654, N5653, N3757, N1407, N2159);
nor NOR4 (N5655, N5641, N2252, N940, N2379);
or OR3 (N5656, N5654, N2910, N2310);
nand NAND4 (N5657, N5656, N2646, N4373, N1526);
and AND3 (N5658, N5638, N4309, N1593);
not NOT1 (N5659, N5650);
nand NAND2 (N5660, N5658, N4469);
or OR2 (N5661, N5645, N2248);
nand NAND2 (N5662, N5642, N2520);
xor XOR2 (N5663, N5655, N4622);
buf BUF1 (N5664, N5657);
buf BUF1 (N5665, N5651);
nand NAND2 (N5666, N5661, N434);
buf BUF1 (N5667, N5652);
nor NOR2 (N5668, N5660, N429);
buf BUF1 (N5669, N5667);
buf BUF1 (N5670, N5649);
not NOT1 (N5671, N5666);
not NOT1 (N5672, N5671);
or OR2 (N5673, N5662, N1657);
xor XOR2 (N5674, N5665, N4960);
xor XOR2 (N5675, N5664, N2753);
or OR3 (N5676, N5659, N4528, N4675);
xor XOR2 (N5677, N5676, N2659);
nand NAND2 (N5678, N5669, N3756);
nand NAND3 (N5679, N5673, N1724, N1909);
xor XOR2 (N5680, N5675, N4254);
nand NAND2 (N5681, N5672, N5397);
and AND3 (N5682, N5670, N3190, N740);
nor NOR2 (N5683, N5631, N4968);
xor XOR2 (N5684, N5680, N540);
xor XOR2 (N5685, N5683, N1616);
not NOT1 (N5686, N5681);
nand NAND2 (N5687, N5677, N1628);
buf BUF1 (N5688, N5674);
not NOT1 (N5689, N5686);
buf BUF1 (N5690, N5685);
nand NAND2 (N5691, N5682, N3532);
buf BUF1 (N5692, N5690);
buf BUF1 (N5693, N5687);
buf BUF1 (N5694, N5679);
buf BUF1 (N5695, N5668);
nor NOR4 (N5696, N5692, N603, N5128, N3637);
xor XOR2 (N5697, N5684, N714);
not NOT1 (N5698, N5678);
and AND3 (N5699, N5693, N3054, N4733);
nand NAND4 (N5700, N5691, N5555, N4419, N4822);
and AND3 (N5701, N5697, N5401, N2320);
buf BUF1 (N5702, N5688);
nor NOR4 (N5703, N5698, N1530, N1513, N887);
nand NAND2 (N5704, N5696, N1585);
not NOT1 (N5705, N5663);
or OR4 (N5706, N5701, N2087, N3982, N2231);
nor NOR4 (N5707, N5705, N3260, N4294, N2595);
or OR2 (N5708, N5695, N108);
and AND4 (N5709, N5706, N2170, N3342, N299);
or OR4 (N5710, N5707, N1214, N3268, N4269);
xor XOR2 (N5711, N5708, N682);
buf BUF1 (N5712, N5699);
not NOT1 (N5713, N5700);
or OR2 (N5714, N5712, N2607);
buf BUF1 (N5715, N5710);
buf BUF1 (N5716, N5714);
and AND3 (N5717, N5689, N256, N4938);
not NOT1 (N5718, N5713);
and AND4 (N5719, N5704, N4067, N1632, N2782);
and AND3 (N5720, N5719, N1622, N3212);
nand NAND3 (N5721, N5716, N4778, N3676);
nand NAND4 (N5722, N5715, N1770, N4024, N146);
not NOT1 (N5723, N5709);
buf BUF1 (N5724, N5717);
xor XOR2 (N5725, N5694, N2524);
or OR2 (N5726, N5723, N3860);
nor NOR2 (N5727, N5711, N4359);
not NOT1 (N5728, N5702);
not NOT1 (N5729, N5725);
buf BUF1 (N5730, N5728);
not NOT1 (N5731, N5726);
and AND2 (N5732, N5720, N1505);
nor NOR2 (N5733, N5729, N1809);
xor XOR2 (N5734, N5727, N4285);
xor XOR2 (N5735, N5733, N1322);
nand NAND4 (N5736, N5721, N4094, N5542, N799);
nor NOR2 (N5737, N5730, N4689);
xor XOR2 (N5738, N5724, N2896);
nor NOR4 (N5739, N5737, N137, N655, N216);
and AND4 (N5740, N5722, N3885, N3217, N4338);
xor XOR2 (N5741, N5734, N5186);
or OR4 (N5742, N5718, N1145, N2214, N3979);
nand NAND3 (N5743, N5732, N780, N1411);
and AND2 (N5744, N5738, N1631);
nand NAND3 (N5745, N5731, N1045, N494);
buf BUF1 (N5746, N5739);
and AND3 (N5747, N5742, N1547, N5249);
xor XOR2 (N5748, N5746, N3740);
and AND3 (N5749, N5748, N4466, N494);
or OR3 (N5750, N5743, N4623, N2441);
not NOT1 (N5751, N5750);
or OR3 (N5752, N5703, N3474, N5697);
xor XOR2 (N5753, N5751, N5184);
nor NOR3 (N5754, N5747, N1429, N924);
xor XOR2 (N5755, N5741, N1022);
nor NOR4 (N5756, N5753, N320, N1227, N5190);
buf BUF1 (N5757, N5752);
nor NOR2 (N5758, N5735, N3042);
xor XOR2 (N5759, N5744, N2127);
or OR4 (N5760, N5756, N4495, N4366, N3231);
not NOT1 (N5761, N5757);
nand NAND2 (N5762, N5758, N1024);
buf BUF1 (N5763, N5759);
and AND3 (N5764, N5754, N839, N3931);
nor NOR2 (N5765, N5749, N3603);
and AND4 (N5766, N5763, N1488, N5228, N3908);
or OR3 (N5767, N5764, N4683, N3926);
not NOT1 (N5768, N5765);
xor XOR2 (N5769, N5736, N4374);
nor NOR4 (N5770, N5769, N4617, N1125, N2826);
not NOT1 (N5771, N5760);
not NOT1 (N5772, N5761);
buf BUF1 (N5773, N5762);
xor XOR2 (N5774, N5770, N3883);
nor NOR2 (N5775, N5773, N4282);
not NOT1 (N5776, N5772);
xor XOR2 (N5777, N5740, N4199);
nor NOR4 (N5778, N5767, N5138, N4671, N2369);
buf BUF1 (N5779, N5776);
buf BUF1 (N5780, N5777);
nand NAND2 (N5781, N5778, N2823);
buf BUF1 (N5782, N5768);
and AND4 (N5783, N5771, N4488, N3524, N3692);
nand NAND2 (N5784, N5781, N358);
or OR3 (N5785, N5766, N1264, N2239);
and AND2 (N5786, N5775, N1329);
buf BUF1 (N5787, N5745);
nor NOR3 (N5788, N5784, N2191, N2007);
nand NAND4 (N5789, N5785, N3350, N5548, N1668);
or OR3 (N5790, N5755, N2547, N5445);
not NOT1 (N5791, N5783);
xor XOR2 (N5792, N5789, N1173);
nand NAND4 (N5793, N5786, N1536, N1915, N3719);
nor NOR3 (N5794, N5780, N5119, N5240);
not NOT1 (N5795, N5788);
xor XOR2 (N5796, N5793, N565);
nand NAND3 (N5797, N5779, N5120, N2797);
buf BUF1 (N5798, N5790);
xor XOR2 (N5799, N5797, N4137);
nand NAND2 (N5800, N5798, N1577);
and AND2 (N5801, N5787, N3065);
nor NOR2 (N5802, N5791, N3734);
nor NOR4 (N5803, N5774, N4520, N227, N1600);
and AND4 (N5804, N5795, N4528, N1942, N757);
nor NOR2 (N5805, N5792, N3641);
and AND2 (N5806, N5801, N1650);
buf BUF1 (N5807, N5794);
buf BUF1 (N5808, N5807);
not NOT1 (N5809, N5802);
or OR3 (N5810, N5796, N1831, N3504);
not NOT1 (N5811, N5782);
and AND3 (N5812, N5800, N4288, N698);
and AND3 (N5813, N5803, N3476, N4224);
buf BUF1 (N5814, N5805);
nand NAND3 (N5815, N5811, N2086, N233);
xor XOR2 (N5816, N5815, N562);
nor NOR3 (N5817, N5816, N4625, N1219);
not NOT1 (N5818, N5812);
nand NAND3 (N5819, N5806, N4856, N964);
not NOT1 (N5820, N5808);
nand NAND3 (N5821, N5818, N2901, N1376);
and AND2 (N5822, N5819, N5350);
xor XOR2 (N5823, N5822, N1602);
xor XOR2 (N5824, N5810, N80);
nand NAND3 (N5825, N5821, N4757, N4352);
nor NOR3 (N5826, N5809, N4875, N87);
buf BUF1 (N5827, N5814);
buf BUF1 (N5828, N5827);
buf BUF1 (N5829, N5825);
and AND4 (N5830, N5823, N3021, N3604, N5123);
and AND3 (N5831, N5830, N555, N5006);
buf BUF1 (N5832, N5826);
not NOT1 (N5833, N5813);
not NOT1 (N5834, N5833);
and AND2 (N5835, N5824, N4281);
xor XOR2 (N5836, N5828, N4517);
and AND4 (N5837, N5804, N3230, N3341, N3408);
or OR4 (N5838, N5837, N990, N1726, N1191);
nand NAND2 (N5839, N5835, N5120);
nand NAND4 (N5840, N5839, N828, N4797, N2950);
nor NOR2 (N5841, N5817, N2048);
nand NAND2 (N5842, N5829, N1154);
nor NOR4 (N5843, N5842, N5758, N3921, N5750);
or OR3 (N5844, N5831, N382, N5714);
xor XOR2 (N5845, N5838, N48);
or OR3 (N5846, N5840, N3016, N5153);
nand NAND3 (N5847, N5841, N1295, N866);
xor XOR2 (N5848, N5834, N978);
or OR3 (N5849, N5848, N5176, N5077);
or OR3 (N5850, N5847, N4662, N5321);
nor NOR4 (N5851, N5844, N3989, N1560, N5331);
buf BUF1 (N5852, N5845);
nor NOR2 (N5853, N5846, N1140);
nor NOR3 (N5854, N5852, N534, N701);
not NOT1 (N5855, N5854);
nor NOR4 (N5856, N5855, N1729, N2842, N1701);
nand NAND2 (N5857, N5851, N5362);
xor XOR2 (N5858, N5853, N5745);
xor XOR2 (N5859, N5836, N4470);
and AND3 (N5860, N5849, N4457, N514);
nor NOR2 (N5861, N5843, N3491);
nand NAND4 (N5862, N5799, N1981, N1040, N77);
nor NOR4 (N5863, N5857, N5262, N3550, N5032);
and AND3 (N5864, N5850, N301, N1133);
nand NAND3 (N5865, N5864, N4798, N4822);
nor NOR3 (N5866, N5863, N3223, N4975);
nand NAND2 (N5867, N5820, N3362);
nor NOR3 (N5868, N5865, N1678, N2377);
or OR3 (N5869, N5862, N425, N102);
xor XOR2 (N5870, N5869, N4901);
nor NOR2 (N5871, N5866, N986);
not NOT1 (N5872, N5868);
and AND3 (N5873, N5871, N908, N5776);
nor NOR4 (N5874, N5861, N1558, N1845, N4244);
and AND4 (N5875, N5870, N920, N5509, N5300);
nor NOR3 (N5876, N5874, N4748, N5869);
buf BUF1 (N5877, N5876);
nor NOR4 (N5878, N5875, N2852, N3796, N1927);
not NOT1 (N5879, N5872);
or OR3 (N5880, N5873, N1159, N242);
nand NAND4 (N5881, N5867, N2736, N1450, N2412);
or OR2 (N5882, N5880, N708);
or OR2 (N5883, N5879, N4381);
buf BUF1 (N5884, N5883);
buf BUF1 (N5885, N5858);
or OR2 (N5886, N5881, N4318);
and AND3 (N5887, N5832, N5289, N5477);
buf BUF1 (N5888, N5877);
not NOT1 (N5889, N5856);
not NOT1 (N5890, N5884);
not NOT1 (N5891, N5889);
xor XOR2 (N5892, N5860, N1804);
nor NOR4 (N5893, N5888, N4305, N2073, N2169);
nor NOR2 (N5894, N5878, N2897);
nor NOR2 (N5895, N5859, N2988);
buf BUF1 (N5896, N5891);
not NOT1 (N5897, N5890);
nand NAND4 (N5898, N5882, N3586, N2385, N2286);
not NOT1 (N5899, N5897);
not NOT1 (N5900, N5899);
not NOT1 (N5901, N5893);
xor XOR2 (N5902, N5896, N643);
nand NAND3 (N5903, N5885, N5353, N4804);
and AND3 (N5904, N5903, N2294, N300);
not NOT1 (N5905, N5886);
xor XOR2 (N5906, N5892, N3);
or OR2 (N5907, N5898, N3097);
or OR2 (N5908, N5894, N1306);
nand NAND3 (N5909, N5901, N1716, N2209);
buf BUF1 (N5910, N5887);
and AND3 (N5911, N5905, N4358, N1404);
or OR2 (N5912, N5907, N4184);
and AND3 (N5913, N5911, N4064, N3539);
and AND2 (N5914, N5900, N1504);
or OR3 (N5915, N5895, N534, N5592);
or OR3 (N5916, N5915, N4799, N3968);
buf BUF1 (N5917, N5913);
nor NOR2 (N5918, N5914, N2855);
nor NOR3 (N5919, N5910, N3976, N626);
or OR3 (N5920, N5904, N5464, N5536);
xor XOR2 (N5921, N5902, N2136);
nand NAND2 (N5922, N5921, N5242);
and AND4 (N5923, N5908, N1767, N496, N4906);
and AND2 (N5924, N5920, N254);
buf BUF1 (N5925, N5919);
nand NAND3 (N5926, N5909, N2322, N559);
nand NAND4 (N5927, N5918, N811, N3900, N102);
xor XOR2 (N5928, N5925, N4998);
nand NAND4 (N5929, N5916, N5271, N4971, N432);
nor NOR3 (N5930, N5926, N4721, N4088);
or OR4 (N5931, N5928, N1891, N3820, N2203);
not NOT1 (N5932, N5929);
nand NAND3 (N5933, N5930, N831, N5565);
nor NOR4 (N5934, N5923, N5798, N4668, N1362);
not NOT1 (N5935, N5931);
and AND3 (N5936, N5935, N895, N5117);
or OR3 (N5937, N5922, N1127, N4529);
or OR4 (N5938, N5906, N2045, N4842, N2);
nor NOR4 (N5939, N5936, N2906, N1706, N4920);
not NOT1 (N5940, N5934);
nor NOR3 (N5941, N5933, N1630, N5250);
nor NOR2 (N5942, N5940, N668);
and AND2 (N5943, N5924, N5357);
xor XOR2 (N5944, N5937, N828);
or OR4 (N5945, N5942, N3806, N1097, N916);
and AND2 (N5946, N5943, N4326);
or OR4 (N5947, N5938, N335, N1086, N5577);
buf BUF1 (N5948, N5947);
nor NOR4 (N5949, N5939, N2372, N678, N5132);
xor XOR2 (N5950, N5912, N3456);
xor XOR2 (N5951, N5946, N4228);
and AND4 (N5952, N5941, N5758, N1343, N5670);
and AND3 (N5953, N5949, N4410, N2602);
or OR2 (N5954, N5917, N5825);
nand NAND4 (N5955, N5954, N5594, N3367, N5109);
nand NAND2 (N5956, N5945, N3430);
xor XOR2 (N5957, N5927, N3031);
xor XOR2 (N5958, N5955, N4656);
xor XOR2 (N5959, N5956, N4633);
nand NAND3 (N5960, N5948, N2810, N2365);
buf BUF1 (N5961, N5932);
or OR4 (N5962, N5960, N2718, N2960, N2052);
and AND2 (N5963, N5952, N674);
and AND3 (N5964, N5951, N1933, N224);
xor XOR2 (N5965, N5961, N604);
or OR4 (N5966, N5959, N1012, N4740, N2068);
buf BUF1 (N5967, N5950);
nor NOR2 (N5968, N5944, N3418);
not NOT1 (N5969, N5957);
and AND3 (N5970, N5965, N1288, N484);
not NOT1 (N5971, N5964);
buf BUF1 (N5972, N5953);
and AND4 (N5973, N5969, N1995, N5553, N1507);
nand NAND2 (N5974, N5967, N5408);
xor XOR2 (N5975, N5970, N4438);
buf BUF1 (N5976, N5966);
buf BUF1 (N5977, N5962);
not NOT1 (N5978, N5958);
nor NOR3 (N5979, N5963, N3506, N2230);
and AND4 (N5980, N5974, N3968, N1446, N3186);
or OR3 (N5981, N5979, N412, N988);
and AND3 (N5982, N5971, N4335, N769);
xor XOR2 (N5983, N5976, N2864);
nand NAND3 (N5984, N5977, N2913, N3054);
not NOT1 (N5985, N5978);
or OR3 (N5986, N5985, N5464, N29);
or OR2 (N5987, N5981, N1938);
and AND2 (N5988, N5973, N2284);
xor XOR2 (N5989, N5968, N515);
or OR2 (N5990, N5982, N4026);
nor NOR3 (N5991, N5990, N2824, N3014);
or OR3 (N5992, N5983, N1713, N5507);
or OR3 (N5993, N5987, N4501, N4571);
nand NAND2 (N5994, N5988, N4225);
or OR3 (N5995, N5993, N1205, N221);
nand NAND4 (N5996, N5980, N651, N5006, N4005);
and AND4 (N5997, N5986, N3485, N718, N1908);
or OR2 (N5998, N5984, N51);
or OR3 (N5999, N5996, N4264, N4585);
nor NOR4 (N6000, N5989, N2026, N5570, N1007);
nand NAND3 (N6001, N5992, N5896, N1303);
nand NAND3 (N6002, N6001, N4154, N5809);
xor XOR2 (N6003, N5997, N5341);
nor NOR4 (N6004, N5999, N2912, N3757, N4975);
or OR3 (N6005, N5991, N1185, N4985);
xor XOR2 (N6006, N5995, N2694);
nor NOR2 (N6007, N6004, N2533);
xor XOR2 (N6008, N6000, N5207);
not NOT1 (N6009, N6006);
xor XOR2 (N6010, N5975, N4122);
xor XOR2 (N6011, N6007, N2001);
xor XOR2 (N6012, N6005, N2514);
or OR4 (N6013, N6002, N2856, N702, N5758);
nand NAND3 (N6014, N6009, N1303, N2522);
and AND3 (N6015, N6010, N2180, N4589);
not NOT1 (N6016, N6014);
not NOT1 (N6017, N6016);
nor NOR4 (N6018, N6017, N60, N60, N29);
nand NAND3 (N6019, N5998, N1121, N3763);
and AND3 (N6020, N6012, N955, N3217);
buf BUF1 (N6021, N6008);
xor XOR2 (N6022, N6020, N3123);
and AND4 (N6023, N6021, N4366, N319, N5293);
and AND4 (N6024, N5972, N2834, N3321, N1372);
or OR2 (N6025, N6024, N374);
and AND4 (N6026, N6023, N5347, N2183, N3673);
buf BUF1 (N6027, N6025);
xor XOR2 (N6028, N6015, N1504);
nor NOR3 (N6029, N6022, N685, N2122);
and AND2 (N6030, N6026, N911);
nor NOR3 (N6031, N6028, N1747, N239);
nand NAND4 (N6032, N6003, N4395, N900, N1614);
nand NAND2 (N6033, N6030, N5168);
not NOT1 (N6034, N6032);
nor NOR3 (N6035, N6018, N458, N4252);
nand NAND2 (N6036, N6033, N4080);
or OR4 (N6037, N6035, N1560, N4208, N4962);
nor NOR4 (N6038, N6037, N1731, N969, N1228);
nor NOR4 (N6039, N6029, N5221, N3921, N3334);
nor NOR2 (N6040, N6027, N735);
nor NOR3 (N6041, N6040, N1507, N972);
nand NAND3 (N6042, N6013, N5071, N5658);
xor XOR2 (N6043, N6038, N3064);
nand NAND3 (N6044, N6043, N2841, N1278);
xor XOR2 (N6045, N6019, N5068);
nor NOR3 (N6046, N6045, N2923, N959);
not NOT1 (N6047, N6044);
and AND4 (N6048, N6041, N2271, N4903, N1608);
buf BUF1 (N6049, N6046);
not NOT1 (N6050, N6047);
not NOT1 (N6051, N6048);
and AND3 (N6052, N6031, N5660, N2764);
not NOT1 (N6053, N6050);
or OR3 (N6054, N6053, N4805, N4168);
nor NOR4 (N6055, N6051, N606, N814, N2106);
buf BUF1 (N6056, N6039);
not NOT1 (N6057, N6011);
and AND4 (N6058, N6042, N2215, N5842, N4921);
and AND2 (N6059, N6034, N120);
buf BUF1 (N6060, N6036);
xor XOR2 (N6061, N6060, N4365);
or OR2 (N6062, N5994, N332);
nand NAND3 (N6063, N6058, N3564, N4215);
not NOT1 (N6064, N6057);
and AND3 (N6065, N6049, N4789, N4792);
nor NOR3 (N6066, N6052, N5758, N2406);
nor NOR3 (N6067, N6059, N2244, N5063);
or OR4 (N6068, N6061, N2977, N2991, N121);
xor XOR2 (N6069, N6062, N85);
and AND3 (N6070, N6055, N3100, N3463);
nor NOR3 (N6071, N6063, N2453, N5940);
nor NOR2 (N6072, N6070, N3212);
and AND3 (N6073, N6065, N5215, N3536);
nand NAND3 (N6074, N6069, N4500, N1466);
buf BUF1 (N6075, N6066);
nor NOR4 (N6076, N6071, N5508, N3927, N1742);
buf BUF1 (N6077, N6064);
nand NAND2 (N6078, N6074, N1689);
nand NAND3 (N6079, N6072, N2812, N1177);
buf BUF1 (N6080, N6077);
or OR3 (N6081, N6080, N1219, N3931);
nor NOR3 (N6082, N6067, N2128, N5647);
and AND3 (N6083, N6073, N3434, N1636);
buf BUF1 (N6084, N6068);
nor NOR3 (N6085, N6056, N2084, N10);
xor XOR2 (N6086, N6083, N720);
nand NAND2 (N6087, N6078, N5473);
and AND3 (N6088, N6054, N512, N2929);
or OR3 (N6089, N6088, N1397, N2467);
and AND4 (N6090, N6079, N4173, N4588, N4634);
xor XOR2 (N6091, N6084, N571);
xor XOR2 (N6092, N6085, N3277);
buf BUF1 (N6093, N6082);
or OR2 (N6094, N6076, N885);
or OR2 (N6095, N6093, N100);
nand NAND2 (N6096, N6094, N5786);
or OR3 (N6097, N6095, N3857, N462);
not NOT1 (N6098, N6089);
nor NOR3 (N6099, N6090, N4853, N5575);
or OR4 (N6100, N6096, N4220, N4305, N4873);
and AND2 (N6101, N6099, N4640);
not NOT1 (N6102, N6087);
or OR3 (N6103, N6091, N2541, N1209);
nand NAND4 (N6104, N6101, N923, N2025, N1299);
nand NAND4 (N6105, N6103, N4594, N525, N5767);
xor XOR2 (N6106, N6097, N2588);
or OR4 (N6107, N6086, N5365, N5460, N2733);
and AND2 (N6108, N6100, N5997);
not NOT1 (N6109, N6102);
or OR3 (N6110, N6109, N4548, N1212);
not NOT1 (N6111, N6104);
not NOT1 (N6112, N6106);
buf BUF1 (N6113, N6112);
nand NAND3 (N6114, N6107, N396, N3499);
and AND4 (N6115, N6114, N3723, N1528, N5548);
and AND4 (N6116, N6111, N5242, N601, N5439);
or OR3 (N6117, N6116, N66, N629);
not NOT1 (N6118, N6115);
and AND2 (N6119, N6108, N2630);
nand NAND2 (N6120, N6119, N299);
nand NAND4 (N6121, N6118, N6051, N1297, N4437);
xor XOR2 (N6122, N6075, N4089);
and AND2 (N6123, N6122, N2312);
buf BUF1 (N6124, N6092);
not NOT1 (N6125, N6124);
and AND4 (N6126, N6117, N4808, N686, N872);
nand NAND4 (N6127, N6098, N5323, N534, N1586);
buf BUF1 (N6128, N6123);
nand NAND3 (N6129, N6113, N4363, N1427);
not NOT1 (N6130, N6129);
xor XOR2 (N6131, N6130, N1866);
or OR2 (N6132, N6131, N6010);
not NOT1 (N6133, N6125);
and AND2 (N6134, N6105, N1966);
xor XOR2 (N6135, N6110, N2642);
or OR2 (N6136, N6128, N2592);
buf BUF1 (N6137, N6121);
nand NAND4 (N6138, N6126, N4881, N4888, N2456);
buf BUF1 (N6139, N6127);
or OR3 (N6140, N6133, N3458, N2414);
nor NOR2 (N6141, N6120, N2482);
nand NAND3 (N6142, N6141, N2836, N1449);
xor XOR2 (N6143, N6140, N2915);
nor NOR2 (N6144, N6081, N3453);
and AND3 (N6145, N6135, N2274, N4840);
nand NAND3 (N6146, N6137, N723, N2882);
nand NAND3 (N6147, N6145, N3402, N3609);
buf BUF1 (N6148, N6136);
not NOT1 (N6149, N6132);
or OR3 (N6150, N6142, N677, N5114);
nor NOR4 (N6151, N6147, N4849, N3274, N4106);
not NOT1 (N6152, N6139);
nand NAND2 (N6153, N6138, N5997);
or OR4 (N6154, N6153, N1187, N1021, N2707);
xor XOR2 (N6155, N6146, N4698);
or OR2 (N6156, N6149, N4842);
or OR2 (N6157, N6152, N3706);
and AND4 (N6158, N6143, N2942, N4296, N1234);
not NOT1 (N6159, N6144);
or OR4 (N6160, N6155, N6065, N203, N4494);
and AND2 (N6161, N6159, N673);
nor NOR3 (N6162, N6148, N4463, N5031);
and AND4 (N6163, N6160, N3155, N4770, N815);
or OR4 (N6164, N6157, N1193, N1101, N5532);
xor XOR2 (N6165, N6151, N3116);
and AND4 (N6166, N6162, N3427, N4819, N2077);
nor NOR2 (N6167, N6150, N1105);
not NOT1 (N6168, N6164);
not NOT1 (N6169, N6158);
nand NAND4 (N6170, N6166, N1522, N4451, N2885);
nor NOR4 (N6171, N6170, N5773, N5201, N3095);
buf BUF1 (N6172, N6161);
or OR3 (N6173, N6167, N2754, N5747);
and AND2 (N6174, N6165, N754);
not NOT1 (N6175, N6134);
not NOT1 (N6176, N6171);
buf BUF1 (N6177, N6174);
and AND2 (N6178, N6163, N1413);
not NOT1 (N6179, N6168);
and AND4 (N6180, N6176, N1619, N1374, N5377);
and AND3 (N6181, N6177, N2943, N2581);
nor NOR3 (N6182, N6175, N2502, N737);
or OR2 (N6183, N6172, N817);
xor XOR2 (N6184, N6154, N1851);
nand NAND2 (N6185, N6180, N398);
not NOT1 (N6186, N6181);
not NOT1 (N6187, N6179);
xor XOR2 (N6188, N6186, N2395);
buf BUF1 (N6189, N6185);
xor XOR2 (N6190, N6189, N1933);
nand NAND2 (N6191, N6173, N5857);
and AND2 (N6192, N6169, N1028);
not NOT1 (N6193, N6188);
nand NAND3 (N6194, N6190, N5196, N2354);
xor XOR2 (N6195, N6187, N2739);
and AND4 (N6196, N6194, N4970, N3451, N5203);
nand NAND4 (N6197, N6193, N5116, N2075, N2571);
buf BUF1 (N6198, N6183);
buf BUF1 (N6199, N6198);
or OR4 (N6200, N6156, N5023, N4565, N5808);
not NOT1 (N6201, N6192);
xor XOR2 (N6202, N6196, N5049);
or OR2 (N6203, N6182, N2502);
or OR3 (N6204, N6191, N5207, N1878);
or OR3 (N6205, N6178, N5550, N2000);
not NOT1 (N6206, N6205);
xor XOR2 (N6207, N6197, N1478);
not NOT1 (N6208, N6202);
or OR3 (N6209, N6207, N3148, N6126);
not NOT1 (N6210, N6208);
and AND4 (N6211, N6184, N72, N5020, N4845);
xor XOR2 (N6212, N6199, N1074);
not NOT1 (N6213, N6212);
nor NOR4 (N6214, N6211, N1566, N4019, N5276);
buf BUF1 (N6215, N6214);
nor NOR4 (N6216, N6210, N4487, N1480, N2191);
buf BUF1 (N6217, N6195);
buf BUF1 (N6218, N6204);
nor NOR2 (N6219, N6200, N723);
xor XOR2 (N6220, N6219, N4630);
not NOT1 (N6221, N6216);
nor NOR2 (N6222, N6206, N807);
nand NAND3 (N6223, N6217, N1634, N1355);
or OR2 (N6224, N6213, N3512);
xor XOR2 (N6225, N6223, N3862);
nand NAND4 (N6226, N6224, N5031, N5602, N1235);
buf BUF1 (N6227, N6226);
buf BUF1 (N6228, N6215);
nand NAND3 (N6229, N6203, N2867, N4663);
xor XOR2 (N6230, N6227, N4715);
or OR3 (N6231, N6229, N5091, N1115);
buf BUF1 (N6232, N6222);
and AND2 (N6233, N6201, N4520);
xor XOR2 (N6234, N6228, N63);
nor NOR4 (N6235, N6232, N821, N4874, N2367);
nand NAND2 (N6236, N6233, N2238);
and AND4 (N6237, N6218, N4562, N1816, N5434);
xor XOR2 (N6238, N6221, N5224);
nor NOR2 (N6239, N6234, N3836);
nor NOR2 (N6240, N6225, N2289);
nor NOR2 (N6241, N6230, N2178);
buf BUF1 (N6242, N6239);
or OR4 (N6243, N6242, N1593, N3305, N5131);
buf BUF1 (N6244, N6220);
buf BUF1 (N6245, N6238);
xor XOR2 (N6246, N6237, N4932);
nand NAND3 (N6247, N6231, N2190, N4676);
nor NOR3 (N6248, N6235, N3651, N5085);
not NOT1 (N6249, N6240);
nand NAND2 (N6250, N6243, N2324);
nand NAND4 (N6251, N6249, N4381, N5606, N1670);
buf BUF1 (N6252, N6250);
and AND2 (N6253, N6252, N4556);
not NOT1 (N6254, N6251);
or OR3 (N6255, N6248, N466, N5958);
xor XOR2 (N6256, N6247, N1766);
xor XOR2 (N6257, N6209, N1125);
and AND3 (N6258, N6257, N3873, N4119);
and AND4 (N6259, N6258, N3241, N2073, N5691);
buf BUF1 (N6260, N6256);
buf BUF1 (N6261, N6255);
and AND3 (N6262, N6236, N2891, N4289);
xor XOR2 (N6263, N6241, N507);
xor XOR2 (N6264, N6261, N5693);
not NOT1 (N6265, N6260);
nor NOR4 (N6266, N6254, N4639, N668, N3908);
buf BUF1 (N6267, N6253);
nor NOR4 (N6268, N6244, N2629, N4992, N5442);
nor NOR4 (N6269, N6259, N4540, N3313, N3486);
and AND2 (N6270, N6263, N1746);
nand NAND3 (N6271, N6266, N6025, N125);
or OR2 (N6272, N6268, N2270);
and AND3 (N6273, N6245, N5255, N1552);
nor NOR3 (N6274, N6271, N1703, N3135);
buf BUF1 (N6275, N6269);
xor XOR2 (N6276, N6274, N2639);
buf BUF1 (N6277, N6265);
nand NAND3 (N6278, N6264, N2125, N5169);
nor NOR4 (N6279, N6272, N1987, N385, N4494);
nor NOR2 (N6280, N6273, N2810);
or OR4 (N6281, N6275, N1703, N6020, N5293);
xor XOR2 (N6282, N6279, N1683);
buf BUF1 (N6283, N6262);
not NOT1 (N6284, N6277);
xor XOR2 (N6285, N6278, N1214);
buf BUF1 (N6286, N6285);
nor NOR3 (N6287, N6280, N3813, N1468);
nor NOR4 (N6288, N6246, N2117, N1485, N906);
nor NOR2 (N6289, N6267, N3606);
or OR3 (N6290, N6281, N3369, N5578);
buf BUF1 (N6291, N6286);
nor NOR2 (N6292, N6287, N5673);
xor XOR2 (N6293, N6276, N4090);
not NOT1 (N6294, N6289);
or OR3 (N6295, N6282, N5933, N1589);
xor XOR2 (N6296, N6288, N4308);
and AND3 (N6297, N6295, N2539, N1796);
and AND3 (N6298, N6292, N84, N2431);
nor NOR2 (N6299, N6290, N4284);
xor XOR2 (N6300, N6284, N2500);
or OR4 (N6301, N6297, N3400, N1946, N4888);
nand NAND4 (N6302, N6283, N1173, N2710, N2136);
nor NOR2 (N6303, N6293, N554);
not NOT1 (N6304, N6294);
buf BUF1 (N6305, N6298);
nand NAND4 (N6306, N6305, N5587, N2888, N6105);
buf BUF1 (N6307, N6304);
or OR3 (N6308, N6291, N6034, N438);
not NOT1 (N6309, N6306);
xor XOR2 (N6310, N6302, N1824);
xor XOR2 (N6311, N6299, N5531);
buf BUF1 (N6312, N6310);
nor NOR2 (N6313, N6296, N3202);
and AND2 (N6314, N6313, N2853);
xor XOR2 (N6315, N6301, N2970);
and AND2 (N6316, N6300, N6125);
nand NAND4 (N6317, N6307, N170, N5537, N1178);
xor XOR2 (N6318, N6314, N4384);
xor XOR2 (N6319, N6309, N3862);
not NOT1 (N6320, N6311);
xor XOR2 (N6321, N6315, N2353);
and AND2 (N6322, N6316, N3764);
or OR4 (N6323, N6321, N2799, N3900, N2448);
or OR2 (N6324, N6319, N6142);
nand NAND2 (N6325, N6308, N3618);
buf BUF1 (N6326, N6318);
and AND3 (N6327, N6325, N5910, N3597);
nand NAND3 (N6328, N6317, N4640, N4370);
xor XOR2 (N6329, N6303, N3499);
nor NOR4 (N6330, N6270, N5231, N994, N3188);
and AND2 (N6331, N6323, N1733);
xor XOR2 (N6332, N6328, N4048);
and AND4 (N6333, N6320, N5405, N5856, N3620);
nor NOR3 (N6334, N6329, N4474, N314);
not NOT1 (N6335, N6334);
and AND2 (N6336, N6324, N6187);
not NOT1 (N6337, N6336);
buf BUF1 (N6338, N6312);
nand NAND3 (N6339, N6337, N4912, N2376);
nor NOR3 (N6340, N6330, N1454, N3672);
nand NAND4 (N6341, N6327, N4313, N4902, N3650);
nor NOR3 (N6342, N6338, N1033, N4942);
and AND3 (N6343, N6342, N4513, N3425);
nand NAND3 (N6344, N6339, N5629, N699);
buf BUF1 (N6345, N6343);
buf BUF1 (N6346, N6335);
nor NOR4 (N6347, N6322, N6064, N2799, N4718);
nand NAND2 (N6348, N6332, N3087);
nand NAND3 (N6349, N6345, N365, N3655);
nor NOR3 (N6350, N6326, N2342, N2366);
buf BUF1 (N6351, N6348);
nor NOR3 (N6352, N6351, N213, N456);
and AND4 (N6353, N6341, N2461, N4494, N1832);
buf BUF1 (N6354, N6340);
and AND3 (N6355, N6353, N5769, N5858);
xor XOR2 (N6356, N6333, N4314);
buf BUF1 (N6357, N6355);
and AND3 (N6358, N6354, N466, N678);
nor NOR3 (N6359, N6347, N2065, N2357);
and AND4 (N6360, N6350, N4772, N3004, N1269);
nor NOR3 (N6361, N6359, N3650, N2951);
nand NAND3 (N6362, N6361, N4405, N5859);
or OR3 (N6363, N6357, N5269, N5225);
xor XOR2 (N6364, N6331, N2426);
buf BUF1 (N6365, N6362);
not NOT1 (N6366, N6349);
or OR4 (N6367, N6346, N3533, N2683, N4243);
not NOT1 (N6368, N6344);
xor XOR2 (N6369, N6368, N3374);
nand NAND4 (N6370, N6360, N4577, N2850, N4763);
nand NAND4 (N6371, N6356, N8, N3962, N2955);
not NOT1 (N6372, N6369);
xor XOR2 (N6373, N6363, N5873);
not NOT1 (N6374, N6358);
not NOT1 (N6375, N6352);
not NOT1 (N6376, N6374);
nor NOR3 (N6377, N6365, N5382, N4800);
nor NOR3 (N6378, N6366, N4473, N679);
not NOT1 (N6379, N6364);
or OR2 (N6380, N6377, N3367);
not NOT1 (N6381, N6380);
or OR3 (N6382, N6372, N1945, N1120);
xor XOR2 (N6383, N6371, N1222);
not NOT1 (N6384, N6382);
nor NOR3 (N6385, N6370, N6020, N1698);
nand NAND3 (N6386, N6383, N827, N2821);
and AND2 (N6387, N6384, N3416);
not NOT1 (N6388, N6375);
nor NOR3 (N6389, N6373, N2282, N1399);
nor NOR4 (N6390, N6387, N1377, N2288, N5995);
buf BUF1 (N6391, N6381);
or OR3 (N6392, N6379, N5396, N1551);
buf BUF1 (N6393, N6388);
nor NOR3 (N6394, N6378, N4631, N2784);
not NOT1 (N6395, N6376);
nand NAND2 (N6396, N6393, N3208);
and AND3 (N6397, N6391, N21, N666);
not NOT1 (N6398, N6392);
nor NOR2 (N6399, N6385, N5677);
xor XOR2 (N6400, N6367, N3124);
nor NOR3 (N6401, N6400, N451, N6335);
and AND4 (N6402, N6386, N2491, N2796, N3960);
buf BUF1 (N6403, N6394);
buf BUF1 (N6404, N6395);
and AND2 (N6405, N6404, N118);
and AND3 (N6406, N6402, N4631, N5017);
buf BUF1 (N6407, N6405);
buf BUF1 (N6408, N6399);
or OR4 (N6409, N6396, N2788, N1856, N2278);
not NOT1 (N6410, N6407);
buf BUF1 (N6411, N6403);
or OR2 (N6412, N6401, N4348);
buf BUF1 (N6413, N6397);
not NOT1 (N6414, N6390);
and AND4 (N6415, N6398, N4961, N4305, N4974);
nand NAND3 (N6416, N6389, N5425, N911);
not NOT1 (N6417, N6410);
not NOT1 (N6418, N6409);
or OR2 (N6419, N6406, N5794);
not NOT1 (N6420, N6417);
nor NOR2 (N6421, N6412, N2445);
not NOT1 (N6422, N6408);
xor XOR2 (N6423, N6420, N4075);
xor XOR2 (N6424, N6413, N5498);
not NOT1 (N6425, N6423);
nor NOR3 (N6426, N6418, N2454, N21);
xor XOR2 (N6427, N6416, N331);
and AND3 (N6428, N6419, N5987, N649);
xor XOR2 (N6429, N6411, N3253);
buf BUF1 (N6430, N6414);
or OR4 (N6431, N6415, N2516, N768, N4860);
not NOT1 (N6432, N6426);
nor NOR2 (N6433, N6432, N824);
buf BUF1 (N6434, N6421);
not NOT1 (N6435, N6422);
nand NAND4 (N6436, N6433, N3317, N249, N1381);
or OR4 (N6437, N6427, N2823, N6115, N3685);
nor NOR4 (N6438, N6424, N2902, N629, N5817);
not NOT1 (N6439, N6437);
nor NOR3 (N6440, N6434, N4286, N5162);
xor XOR2 (N6441, N6429, N5416);
buf BUF1 (N6442, N6425);
nand NAND4 (N6443, N6430, N4443, N1744, N4133);
xor XOR2 (N6444, N6440, N1678);
not NOT1 (N6445, N6438);
buf BUF1 (N6446, N6428);
and AND2 (N6447, N6431, N478);
buf BUF1 (N6448, N6441);
xor XOR2 (N6449, N6446, N5440);
xor XOR2 (N6450, N6443, N2811);
nand NAND2 (N6451, N6442, N2852);
nand NAND4 (N6452, N6451, N4079, N3839, N200);
buf BUF1 (N6453, N6445);
and AND4 (N6454, N6447, N2271, N2090, N2849);
buf BUF1 (N6455, N6444);
buf BUF1 (N6456, N6454);
or OR4 (N6457, N6453, N3247, N1512, N2461);
not NOT1 (N6458, N6457);
xor XOR2 (N6459, N6449, N2367);
or OR4 (N6460, N6448, N679, N4919, N3957);
nor NOR2 (N6461, N6456, N4373);
not NOT1 (N6462, N6452);
nor NOR4 (N6463, N6450, N4255, N4215, N3767);
or OR2 (N6464, N6435, N5845);
xor XOR2 (N6465, N6462, N3786);
nor NOR2 (N6466, N6436, N2294);
or OR4 (N6467, N6458, N5210, N4266, N1173);
nor NOR2 (N6468, N6467, N6431);
buf BUF1 (N6469, N6461);
and AND3 (N6470, N6468, N116, N6277);
xor XOR2 (N6471, N6464, N629);
xor XOR2 (N6472, N6471, N2559);
buf BUF1 (N6473, N6463);
not NOT1 (N6474, N6469);
or OR3 (N6475, N6473, N4274, N1829);
buf BUF1 (N6476, N6470);
not NOT1 (N6477, N6455);
nand NAND2 (N6478, N6460, N2012);
and AND2 (N6479, N6474, N5337);
or OR3 (N6480, N6477, N1159, N6119);
buf BUF1 (N6481, N6476);
or OR2 (N6482, N6479, N909);
xor XOR2 (N6483, N6482, N3761);
nand NAND4 (N6484, N6472, N4056, N5482, N718);
or OR4 (N6485, N6481, N4238, N4501, N6005);
nand NAND4 (N6486, N6459, N2388, N1289, N930);
and AND4 (N6487, N6483, N2799, N1136, N6085);
and AND4 (N6488, N6484, N5192, N5984, N2815);
nand NAND2 (N6489, N6488, N3751);
nor NOR3 (N6490, N6480, N230, N2255);
and AND4 (N6491, N6489, N2265, N3976, N762);
nand NAND2 (N6492, N6486, N5984);
nand NAND4 (N6493, N6487, N4790, N1172, N4792);
nor NOR3 (N6494, N6485, N419, N3563);
nor NOR4 (N6495, N6466, N6047, N2776, N878);
or OR4 (N6496, N6439, N3707, N701, N3875);
and AND4 (N6497, N6490, N2861, N1650, N4161);
buf BUF1 (N6498, N6492);
and AND3 (N6499, N6465, N672, N660);
buf BUF1 (N6500, N6496);
not NOT1 (N6501, N6475);
xor XOR2 (N6502, N6494, N174);
and AND4 (N6503, N6502, N603, N2052, N1538);
nor NOR4 (N6504, N6493, N4084, N2767, N2469);
not NOT1 (N6505, N6503);
xor XOR2 (N6506, N6500, N2008);
not NOT1 (N6507, N6495);
buf BUF1 (N6508, N6507);
nor NOR4 (N6509, N6491, N6106, N5062, N6282);
or OR2 (N6510, N6497, N4712);
xor XOR2 (N6511, N6505, N5015);
xor XOR2 (N6512, N6506, N598);
buf BUF1 (N6513, N6511);
nor NOR2 (N6514, N6513, N3904);
and AND3 (N6515, N6478, N1088, N619);
nand NAND3 (N6516, N6509, N3214, N3406);
xor XOR2 (N6517, N6515, N3127);
not NOT1 (N6518, N6510);
xor XOR2 (N6519, N6518, N5619);
and AND4 (N6520, N6519, N3471, N3072, N1948);
buf BUF1 (N6521, N6520);
nand NAND2 (N6522, N6501, N4545);
not NOT1 (N6523, N6521);
or OR2 (N6524, N6516, N4062);
nor NOR2 (N6525, N6498, N4072);
not NOT1 (N6526, N6523);
nor NOR2 (N6527, N6526, N916);
or OR3 (N6528, N6512, N413, N5258);
and AND3 (N6529, N6528, N1596, N4568);
and AND3 (N6530, N6508, N5708, N4063);
and AND4 (N6531, N6517, N3290, N2780, N4419);
not NOT1 (N6532, N6525);
xor XOR2 (N6533, N6532, N251);
nor NOR4 (N6534, N6533, N3993, N5645, N1355);
buf BUF1 (N6535, N6524);
or OR3 (N6536, N6535, N3280, N1178);
buf BUF1 (N6537, N6534);
nor NOR4 (N6538, N6527, N4110, N6, N929);
buf BUF1 (N6539, N6522);
xor XOR2 (N6540, N6539, N3750);
nor NOR4 (N6541, N6531, N1646, N2202, N986);
buf BUF1 (N6542, N6537);
not NOT1 (N6543, N6536);
or OR2 (N6544, N6499, N5125);
and AND2 (N6545, N6504, N1164);
or OR4 (N6546, N6530, N4316, N291, N558);
xor XOR2 (N6547, N6544, N1335);
nor NOR3 (N6548, N6543, N904, N164);
buf BUF1 (N6549, N6548);
xor XOR2 (N6550, N6529, N530);
xor XOR2 (N6551, N6549, N3020);
buf BUF1 (N6552, N6540);
nand NAND4 (N6553, N6551, N4667, N3317, N2016);
buf BUF1 (N6554, N6550);
buf BUF1 (N6555, N6541);
nand NAND4 (N6556, N6546, N1916, N5151, N1349);
or OR4 (N6557, N6538, N3527, N6522, N3581);
nor NOR2 (N6558, N6545, N2398);
buf BUF1 (N6559, N6547);
or OR2 (N6560, N6559, N5543);
nand NAND3 (N6561, N6555, N5379, N3175);
xor XOR2 (N6562, N6560, N267);
nor NOR4 (N6563, N6514, N1650, N1520, N2280);
xor XOR2 (N6564, N6552, N829);
and AND2 (N6565, N6553, N3253);
or OR4 (N6566, N6558, N4157, N1568, N6152);
buf BUF1 (N6567, N6554);
or OR2 (N6568, N6556, N1900);
buf BUF1 (N6569, N6564);
not NOT1 (N6570, N6565);
xor XOR2 (N6571, N6568, N916);
and AND4 (N6572, N6542, N113, N4916, N554);
nand NAND3 (N6573, N6561, N4119, N3480);
or OR2 (N6574, N6557, N2906);
not NOT1 (N6575, N6574);
and AND2 (N6576, N6566, N6417);
xor XOR2 (N6577, N6576, N4948);
nor NOR4 (N6578, N6572, N5552, N214, N6476);
nor NOR3 (N6579, N6563, N3398, N4031);
buf BUF1 (N6580, N6570);
and AND2 (N6581, N6579, N3782);
xor XOR2 (N6582, N6567, N6309);
nand NAND2 (N6583, N6571, N6450);
buf BUF1 (N6584, N6577);
buf BUF1 (N6585, N6575);
xor XOR2 (N6586, N6573, N3240);
and AND3 (N6587, N6583, N4776, N4938);
and AND2 (N6588, N6562, N3377);
nor NOR3 (N6589, N6581, N4473, N3627);
buf BUF1 (N6590, N6578);
or OR2 (N6591, N6589, N4185);
buf BUF1 (N6592, N6580);
buf BUF1 (N6593, N6584);
nor NOR2 (N6594, N6587, N5738);
nand NAND2 (N6595, N6585, N4566);
and AND3 (N6596, N6595, N3722, N6049);
or OR2 (N6597, N6593, N471);
xor XOR2 (N6598, N6597, N6590);
nor NOR2 (N6599, N768, N1176);
nand NAND4 (N6600, N6569, N4351, N1554, N1013);
or OR3 (N6601, N6598, N210, N598);
and AND4 (N6602, N6601, N2466, N6479, N4243);
nand NAND3 (N6603, N6591, N1478, N3407);
not NOT1 (N6604, N6596);
and AND2 (N6605, N6594, N5937);
nand NAND3 (N6606, N6605, N5945, N5699);
buf BUF1 (N6607, N6592);
and AND3 (N6608, N6599, N263, N5015);
not NOT1 (N6609, N6586);
nor NOR2 (N6610, N6607, N6059);
nor NOR4 (N6611, N6604, N3429, N5547, N78);
and AND2 (N6612, N6611, N4116);
buf BUF1 (N6613, N6603);
and AND3 (N6614, N6606, N2708, N3080);
buf BUF1 (N6615, N6610);
and AND2 (N6616, N6600, N4492);
xor XOR2 (N6617, N6588, N4942);
xor XOR2 (N6618, N6617, N2073);
buf BUF1 (N6619, N6616);
nand NAND4 (N6620, N6582, N4763, N2507, N5092);
nand NAND4 (N6621, N6602, N1676, N423, N6169);
nor NOR4 (N6622, N6609, N710, N3891, N665);
nand NAND4 (N6623, N6613, N6407, N4673, N5111);
nand NAND2 (N6624, N6622, N2335);
nand NAND4 (N6625, N6620, N2666, N2624, N4308);
buf BUF1 (N6626, N6619);
xor XOR2 (N6627, N6615, N5338);
or OR2 (N6628, N6621, N4492);
nor NOR4 (N6629, N6628, N1839, N2336, N4403);
not NOT1 (N6630, N6618);
nand NAND3 (N6631, N6608, N5795, N3628);
nand NAND2 (N6632, N6629, N6361);
nand NAND4 (N6633, N6614, N5779, N334, N3254);
not NOT1 (N6634, N6633);
buf BUF1 (N6635, N6612);
or OR2 (N6636, N6631, N3999);
not NOT1 (N6637, N6635);
nand NAND4 (N6638, N6630, N6168, N3407, N454);
xor XOR2 (N6639, N6624, N514);
xor XOR2 (N6640, N6637, N2414);
buf BUF1 (N6641, N6638);
or OR3 (N6642, N6640, N1763, N3041);
not NOT1 (N6643, N6634);
xor XOR2 (N6644, N6642, N159);
xor XOR2 (N6645, N6625, N5185);
buf BUF1 (N6646, N6627);
xor XOR2 (N6647, N6632, N5826);
buf BUF1 (N6648, N6623);
xor XOR2 (N6649, N6648, N1519);
not NOT1 (N6650, N6645);
not NOT1 (N6651, N6644);
nand NAND2 (N6652, N6636, N1135);
buf BUF1 (N6653, N6643);
or OR2 (N6654, N6646, N4807);
or OR2 (N6655, N6653, N1538);
xor XOR2 (N6656, N6641, N5975);
xor XOR2 (N6657, N6656, N4586);
not NOT1 (N6658, N6647);
nor NOR3 (N6659, N6658, N5948, N6468);
xor XOR2 (N6660, N6655, N3183);
or OR3 (N6661, N6649, N825, N1412);
nor NOR4 (N6662, N6661, N5747, N163, N2477);
and AND2 (N6663, N6626, N895);
nor NOR3 (N6664, N6650, N748, N3792);
xor XOR2 (N6665, N6654, N4967);
not NOT1 (N6666, N6664);
not NOT1 (N6667, N6662);
or OR3 (N6668, N6660, N3205, N4860);
buf BUF1 (N6669, N6666);
and AND3 (N6670, N6657, N1600, N3085);
not NOT1 (N6671, N6659);
or OR2 (N6672, N6668, N1138);
xor XOR2 (N6673, N6652, N3456);
buf BUF1 (N6674, N6651);
buf BUF1 (N6675, N6672);
nand NAND3 (N6676, N6671, N3177, N1038);
not NOT1 (N6677, N6669);
nand NAND4 (N6678, N6670, N3331, N5997, N1108);
not NOT1 (N6679, N6673);
not NOT1 (N6680, N6639);
buf BUF1 (N6681, N6680);
buf BUF1 (N6682, N6679);
xor XOR2 (N6683, N6677, N1369);
xor XOR2 (N6684, N6663, N1482);
nand NAND2 (N6685, N6667, N5678);
nor NOR2 (N6686, N6682, N4329);
buf BUF1 (N6687, N6675);
nand NAND2 (N6688, N6687, N1512);
xor XOR2 (N6689, N6686, N1285);
buf BUF1 (N6690, N6689);
and AND3 (N6691, N6681, N856, N4329);
nand NAND3 (N6692, N6678, N4696, N5876);
nor NOR2 (N6693, N6685, N5707);
xor XOR2 (N6694, N6665, N2088);
and AND4 (N6695, N6693, N4512, N666, N488);
and AND4 (N6696, N6691, N1596, N3315, N3107);
not NOT1 (N6697, N6692);
or OR3 (N6698, N6676, N633, N914);
or OR2 (N6699, N6674, N2687);
not NOT1 (N6700, N6695);
nor NOR2 (N6701, N6700, N2395);
buf BUF1 (N6702, N6694);
or OR3 (N6703, N6683, N6578, N1727);
nor NOR3 (N6704, N6697, N1982, N3968);
nor NOR4 (N6705, N6704, N4036, N4841, N2923);
not NOT1 (N6706, N6699);
and AND2 (N6707, N6705, N55);
and AND3 (N6708, N6688, N1039, N1417);
not NOT1 (N6709, N6702);
nand NAND3 (N6710, N6684, N2496, N5916);
xor XOR2 (N6711, N6706, N6250);
xor XOR2 (N6712, N6698, N4878);
not NOT1 (N6713, N6711);
buf BUF1 (N6714, N6701);
and AND2 (N6715, N6690, N216);
xor XOR2 (N6716, N6712, N5560);
not NOT1 (N6717, N6713);
buf BUF1 (N6718, N6715);
nor NOR3 (N6719, N6696, N2344, N6426);
and AND4 (N6720, N6707, N2840, N2027, N5433);
nand NAND2 (N6721, N6716, N1182);
nand NAND4 (N6722, N6708, N4523, N1822, N2127);
and AND3 (N6723, N6709, N2285, N6425);
buf BUF1 (N6724, N6718);
nand NAND4 (N6725, N6722, N3810, N14, N1972);
and AND4 (N6726, N6714, N6272, N484, N2255);
nand NAND4 (N6727, N6720, N2697, N234, N5237);
or OR2 (N6728, N6724, N77);
nand NAND3 (N6729, N6721, N4495, N4893);
nor NOR4 (N6730, N6717, N167, N1652, N2407);
xor XOR2 (N6731, N6723, N4313);
and AND3 (N6732, N6725, N2083, N593);
or OR2 (N6733, N6731, N3991);
nor NOR2 (N6734, N6730, N1352);
not NOT1 (N6735, N6734);
xor XOR2 (N6736, N6733, N771);
xor XOR2 (N6737, N6719, N6498);
nor NOR2 (N6738, N6736, N5579);
not NOT1 (N6739, N6710);
nor NOR2 (N6740, N6737, N3479);
and AND2 (N6741, N6740, N2);
buf BUF1 (N6742, N6703);
buf BUF1 (N6743, N6742);
or OR2 (N6744, N6743, N3855);
nand NAND3 (N6745, N6727, N3115, N4885);
nand NAND4 (N6746, N6728, N3038, N2574, N777);
buf BUF1 (N6747, N6746);
not NOT1 (N6748, N6745);
and AND2 (N6749, N6741, N5802);
buf BUF1 (N6750, N6749);
and AND3 (N6751, N6747, N2661, N2823);
nand NAND3 (N6752, N6739, N5742, N280);
nand NAND3 (N6753, N6735, N2910, N3385);
nand NAND4 (N6754, N6748, N1788, N1385, N2148);
not NOT1 (N6755, N6738);
nand NAND2 (N6756, N6754, N5625);
buf BUF1 (N6757, N6751);
nor NOR4 (N6758, N6752, N6511, N1410, N2451);
nor NOR4 (N6759, N6753, N1186, N6213, N277);
and AND4 (N6760, N6756, N3535, N408, N3416);
nand NAND2 (N6761, N6744, N3888);
or OR3 (N6762, N6729, N3750, N3425);
buf BUF1 (N6763, N6726);
not NOT1 (N6764, N6732);
or OR3 (N6765, N6759, N2753, N5622);
xor XOR2 (N6766, N6763, N3213);
and AND4 (N6767, N6757, N3213, N1661, N6432);
not NOT1 (N6768, N6758);
and AND2 (N6769, N6767, N4567);
xor XOR2 (N6770, N6766, N1391);
nor NOR3 (N6771, N6755, N4898, N2349);
not NOT1 (N6772, N6769);
or OR3 (N6773, N6760, N2653, N4575);
xor XOR2 (N6774, N6765, N4631);
or OR4 (N6775, N6761, N5639, N4857, N1438);
buf BUF1 (N6776, N6762);
nand NAND4 (N6777, N6750, N6179, N1233, N1409);
nand NAND3 (N6778, N6776, N1930, N1287);
or OR3 (N6779, N6775, N4390, N6467);
not NOT1 (N6780, N6773);
buf BUF1 (N6781, N6764);
nor NOR4 (N6782, N6771, N6000, N4109, N2275);
xor XOR2 (N6783, N6780, N4930);
nor NOR4 (N6784, N6779, N2475, N409, N4080);
not NOT1 (N6785, N6781);
and AND2 (N6786, N6770, N2433);
buf BUF1 (N6787, N6768);
nor NOR3 (N6788, N6774, N5690, N6781);
and AND3 (N6789, N6788, N4386, N361);
not NOT1 (N6790, N6784);
nor NOR4 (N6791, N6782, N3494, N125, N1111);
not NOT1 (N6792, N6791);
not NOT1 (N6793, N6772);
not NOT1 (N6794, N6778);
or OR4 (N6795, N6785, N4384, N4437, N1566);
nand NAND4 (N6796, N6793, N1400, N5471, N1989);
nor NOR2 (N6797, N6787, N4655);
xor XOR2 (N6798, N6797, N1993);
nor NOR2 (N6799, N6777, N4941);
xor XOR2 (N6800, N6799, N3311);
not NOT1 (N6801, N6800);
buf BUF1 (N6802, N6794);
nand NAND3 (N6803, N6792, N4470, N51);
xor XOR2 (N6804, N6803, N3579);
buf BUF1 (N6805, N6798);
nand NAND2 (N6806, N6783, N5059);
and AND3 (N6807, N6795, N2201, N4576);
not NOT1 (N6808, N6807);
nand NAND4 (N6809, N6804, N3308, N457, N2764);
and AND2 (N6810, N6802, N6705);
buf BUF1 (N6811, N6790);
nor NOR2 (N6812, N6806, N5720);
nand NAND2 (N6813, N6786, N6004);
nand NAND4 (N6814, N6805, N3238, N306, N707);
or OR3 (N6815, N6812, N5541, N822);
and AND2 (N6816, N6814, N5606);
nand NAND4 (N6817, N6811, N6611, N638, N388);
or OR3 (N6818, N6809, N38, N1925);
or OR4 (N6819, N6816, N3094, N192, N3791);
xor XOR2 (N6820, N6818, N2663);
nand NAND3 (N6821, N6813, N6104, N862);
xor XOR2 (N6822, N6808, N5349);
xor XOR2 (N6823, N6821, N1359);
nand NAND4 (N6824, N6796, N1411, N1707, N2100);
not NOT1 (N6825, N6801);
buf BUF1 (N6826, N6789);
buf BUF1 (N6827, N6820);
xor XOR2 (N6828, N6825, N5267);
xor XOR2 (N6829, N6819, N3241);
xor XOR2 (N6830, N6827, N3236);
xor XOR2 (N6831, N6830, N305);
not NOT1 (N6832, N6815);
nand NAND2 (N6833, N6817, N5955);
and AND2 (N6834, N6823, N5631);
and AND4 (N6835, N6831, N4852, N3352, N4312);
buf BUF1 (N6836, N6832);
not NOT1 (N6837, N6826);
nand NAND3 (N6838, N6837, N3457, N3420);
and AND2 (N6839, N6835, N951);
nand NAND3 (N6840, N6834, N4549, N5790);
not NOT1 (N6841, N6838);
buf BUF1 (N6842, N6829);
xor XOR2 (N6843, N6828, N6448);
not NOT1 (N6844, N6841);
not NOT1 (N6845, N6836);
xor XOR2 (N6846, N6824, N2102);
buf BUF1 (N6847, N6846);
xor XOR2 (N6848, N6843, N4754);
nor NOR3 (N6849, N6839, N4793, N1887);
xor XOR2 (N6850, N6810, N4961);
not NOT1 (N6851, N6840);
not NOT1 (N6852, N6845);
or OR2 (N6853, N6844, N3766);
and AND3 (N6854, N6851, N3753, N6468);
not NOT1 (N6855, N6850);
buf BUF1 (N6856, N6848);
not NOT1 (N6857, N6842);
xor XOR2 (N6858, N6822, N6246);
buf BUF1 (N6859, N6849);
xor XOR2 (N6860, N6833, N3377);
and AND2 (N6861, N6852, N288);
or OR3 (N6862, N6854, N6187, N5552);
xor XOR2 (N6863, N6862, N2565);
nand NAND2 (N6864, N6860, N2826);
nor NOR4 (N6865, N6857, N1353, N4088, N370);
buf BUF1 (N6866, N6858);
xor XOR2 (N6867, N6866, N2461);
xor XOR2 (N6868, N6847, N3167);
not NOT1 (N6869, N6859);
buf BUF1 (N6870, N6853);
buf BUF1 (N6871, N6867);
nor NOR3 (N6872, N6855, N3189, N354);
buf BUF1 (N6873, N6868);
and AND4 (N6874, N6870, N3692, N2137, N5902);
buf BUF1 (N6875, N6874);
and AND3 (N6876, N6863, N989, N1473);
and AND3 (N6877, N6856, N5029, N5877);
and AND4 (N6878, N6869, N3856, N6684, N6779);
buf BUF1 (N6879, N6877);
and AND3 (N6880, N6875, N4941, N518);
nand NAND4 (N6881, N6871, N5086, N1517, N2297);
nor NOR4 (N6882, N6864, N441, N3021, N3928);
nor NOR3 (N6883, N6872, N2206, N5517);
or OR2 (N6884, N6878, N1447);
or OR2 (N6885, N6879, N4401);
buf BUF1 (N6886, N6876);
and AND3 (N6887, N6883, N1843, N302);
buf BUF1 (N6888, N6873);
nor NOR3 (N6889, N6880, N4126, N554);
nand NAND2 (N6890, N6886, N6017);
not NOT1 (N6891, N6881);
buf BUF1 (N6892, N6889);
or OR2 (N6893, N6885, N3186);
nand NAND2 (N6894, N6861, N414);
and AND4 (N6895, N6884, N4424, N1889, N984);
not NOT1 (N6896, N6894);
or OR2 (N6897, N6888, N6153);
not NOT1 (N6898, N6895);
or OR4 (N6899, N6891, N4146, N3356, N4038);
nor NOR4 (N6900, N6890, N437, N1266, N1768);
and AND2 (N6901, N6898, N4629);
not NOT1 (N6902, N6882);
not NOT1 (N6903, N6865);
or OR3 (N6904, N6903, N2842, N4283);
xor XOR2 (N6905, N6892, N4615);
nand NAND3 (N6906, N6887, N863, N4660);
and AND3 (N6907, N6893, N1711, N1434);
buf BUF1 (N6908, N6896);
nand NAND3 (N6909, N6902, N2758, N6079);
nor NOR2 (N6910, N6899, N3043);
not NOT1 (N6911, N6906);
nand NAND4 (N6912, N6901, N325, N6452, N4285);
nand NAND3 (N6913, N6908, N1162, N2299);
not NOT1 (N6914, N6911);
and AND4 (N6915, N6904, N6458, N5518, N2517);
or OR3 (N6916, N6915, N6701, N1807);
or OR2 (N6917, N6914, N572);
buf BUF1 (N6918, N6907);
nor NOR4 (N6919, N6900, N1503, N3920, N6791);
xor XOR2 (N6920, N6909, N114);
nor NOR2 (N6921, N6913, N4483);
or OR3 (N6922, N6897, N880, N1608);
xor XOR2 (N6923, N6922, N6833);
nor NOR4 (N6924, N6918, N245, N4271, N6412);
xor XOR2 (N6925, N6924, N561);
xor XOR2 (N6926, N6912, N3292);
buf BUF1 (N6927, N6916);
nand NAND3 (N6928, N6917, N2380, N4881);
nor NOR3 (N6929, N6905, N5827, N6292);
xor XOR2 (N6930, N6929, N6896);
or OR4 (N6931, N6910, N6146, N2320, N3353);
not NOT1 (N6932, N6931);
xor XOR2 (N6933, N6927, N769);
buf BUF1 (N6934, N6930);
nor NOR4 (N6935, N6919, N2440, N4788, N2566);
xor XOR2 (N6936, N6935, N249);
nor NOR3 (N6937, N6928, N4923, N6814);
and AND4 (N6938, N6925, N768, N3245, N4739);
buf BUF1 (N6939, N6936);
nor NOR2 (N6940, N6932, N5155);
nand NAND4 (N6941, N6921, N3655, N6747, N6879);
xor XOR2 (N6942, N6941, N4186);
nor NOR3 (N6943, N6934, N5905, N74);
or OR3 (N6944, N6940, N936, N6499);
nor NOR2 (N6945, N6939, N3276);
nand NAND3 (N6946, N6942, N6380, N5444);
nand NAND4 (N6947, N6943, N5967, N1576, N3580);
nor NOR3 (N6948, N6938, N5440, N4814);
xor XOR2 (N6949, N6933, N2876);
buf BUF1 (N6950, N6948);
nand NAND2 (N6951, N6945, N5885);
xor XOR2 (N6952, N6926, N2075);
nand NAND3 (N6953, N6937, N152, N4022);
buf BUF1 (N6954, N6949);
nand NAND2 (N6955, N6947, N2883);
nand NAND3 (N6956, N6946, N1382, N5246);
not NOT1 (N6957, N6944);
or OR2 (N6958, N6954, N3921);
not NOT1 (N6959, N6958);
or OR2 (N6960, N6923, N1005);
nand NAND4 (N6961, N6959, N4168, N5871, N3959);
or OR4 (N6962, N6953, N3545, N6625, N4148);
nand NAND2 (N6963, N6955, N5097);
not NOT1 (N6964, N6963);
nor NOR3 (N6965, N6952, N1285, N4071);
nor NOR2 (N6966, N6960, N5505);
buf BUF1 (N6967, N6950);
nor NOR4 (N6968, N6956, N3715, N3478, N3544);
nor NOR2 (N6969, N6957, N5611);
and AND4 (N6970, N6951, N6120, N4565, N199);
and AND2 (N6971, N6920, N1747);
and AND4 (N6972, N6966, N6297, N390, N4379);
or OR2 (N6973, N6971, N5915);
nor NOR2 (N6974, N6967, N1699);
and AND4 (N6975, N6972, N6151, N858, N4274);
xor XOR2 (N6976, N6965, N4839);
nand NAND3 (N6977, N6969, N720, N4169);
not NOT1 (N6978, N6964);
or OR3 (N6979, N6961, N3607, N1547);
or OR4 (N6980, N6978, N3531, N3152, N2520);
buf BUF1 (N6981, N6968);
xor XOR2 (N6982, N6962, N2467);
buf BUF1 (N6983, N6982);
buf BUF1 (N6984, N6979);
not NOT1 (N6985, N6984);
nor NOR4 (N6986, N6974, N5541, N6130, N5542);
or OR3 (N6987, N6976, N2614, N4366);
nor NOR2 (N6988, N6985, N3515);
buf BUF1 (N6989, N6988);
buf BUF1 (N6990, N6987);
xor XOR2 (N6991, N6975, N5248);
buf BUF1 (N6992, N6980);
or OR2 (N6993, N6981, N3876);
or OR2 (N6994, N6973, N2070);
or OR4 (N6995, N6989, N6713, N3074, N3504);
or OR4 (N6996, N6977, N6318, N6903, N5970);
not NOT1 (N6997, N6996);
not NOT1 (N6998, N6983);
not NOT1 (N6999, N6986);
not NOT1 (N7000, N6999);
xor XOR2 (N7001, N6997, N4100);
or OR2 (N7002, N6992, N4674);
xor XOR2 (N7003, N6994, N3850);
or OR2 (N7004, N7000, N2323);
nor NOR3 (N7005, N7002, N4049, N5381);
nand NAND2 (N7006, N7003, N265);
nor NOR4 (N7007, N6998, N544, N5494, N682);
or OR2 (N7008, N7006, N4333);
nand NAND4 (N7009, N7004, N6999, N4491, N4963);
and AND2 (N7010, N7009, N5476);
nand NAND3 (N7011, N6991, N2697, N632);
and AND2 (N7012, N7008, N1247);
buf BUF1 (N7013, N7007);
xor XOR2 (N7014, N6970, N6303);
buf BUF1 (N7015, N7011);
xor XOR2 (N7016, N6993, N3838);
or OR2 (N7017, N7014, N1404);
nor NOR3 (N7018, N6995, N3052, N4693);
or OR3 (N7019, N7010, N1685, N2767);
nor NOR3 (N7020, N7012, N3029, N4907);
nor NOR4 (N7021, N7018, N1711, N4576, N3742);
not NOT1 (N7022, N7015);
xor XOR2 (N7023, N7005, N5960);
and AND2 (N7024, N7017, N2789);
not NOT1 (N7025, N7013);
not NOT1 (N7026, N7001);
xor XOR2 (N7027, N7022, N457);
buf BUF1 (N7028, N7025);
nor NOR2 (N7029, N7021, N1825);
or OR3 (N7030, N7016, N4866, N1105);
not NOT1 (N7031, N7023);
buf BUF1 (N7032, N7026);
and AND4 (N7033, N7024, N3311, N5739, N185);
xor XOR2 (N7034, N7029, N3660);
or OR2 (N7035, N7027, N4723);
or OR4 (N7036, N7019, N1887, N6960, N1997);
or OR3 (N7037, N6990, N1166, N2394);
nor NOR4 (N7038, N7031, N6042, N6925, N1831);
or OR3 (N7039, N7035, N6273, N6322);
nand NAND3 (N7040, N7033, N5805, N760);
or OR2 (N7041, N7028, N5938);
buf BUF1 (N7042, N7034);
nor NOR4 (N7043, N7041, N6416, N1649, N799);
nor NOR2 (N7044, N7032, N4276);
or OR3 (N7045, N7038, N2667, N1459);
xor XOR2 (N7046, N7036, N5140);
and AND3 (N7047, N7020, N4312, N3651);
buf BUF1 (N7048, N7043);
xor XOR2 (N7049, N7042, N3409);
xor XOR2 (N7050, N7044, N4125);
buf BUF1 (N7051, N7047);
nand NAND3 (N7052, N7045, N40, N1000);
or OR4 (N7053, N7040, N6817, N6681, N5069);
nor NOR4 (N7054, N7049, N1980, N2499, N5039);
nor NOR3 (N7055, N7052, N210, N2254);
and AND2 (N7056, N7055, N6274);
and AND3 (N7057, N7056, N4309, N4196);
and AND3 (N7058, N7053, N5623, N6823);
or OR4 (N7059, N7054, N325, N4488, N1898);
xor XOR2 (N7060, N7059, N4388);
nand NAND3 (N7061, N7057, N4597, N5910);
and AND4 (N7062, N7048, N6774, N2101, N4818);
not NOT1 (N7063, N7050);
nand NAND4 (N7064, N7060, N4421, N6314, N5433);
or OR3 (N7065, N7051, N1852, N2892);
nand NAND2 (N7066, N7046, N4065);
and AND3 (N7067, N7058, N963, N6002);
nand NAND2 (N7068, N7062, N6363);
xor XOR2 (N7069, N7039, N2728);
nand NAND2 (N7070, N7061, N160);
buf BUF1 (N7071, N7065);
xor XOR2 (N7072, N7030, N3715);
not NOT1 (N7073, N7071);
and AND4 (N7074, N7068, N841, N2952, N6327);
xor XOR2 (N7075, N7066, N1733);
nor NOR3 (N7076, N7072, N3568, N215);
buf BUF1 (N7077, N7074);
nor NOR4 (N7078, N7064, N2320, N2719, N6404);
or OR2 (N7079, N7037, N2121);
nor NOR2 (N7080, N7063, N6381);
nand NAND4 (N7081, N7080, N4200, N6316, N3430);
and AND2 (N7082, N7078, N4938);
xor XOR2 (N7083, N7073, N5753);
xor XOR2 (N7084, N7076, N4529);
buf BUF1 (N7085, N7070);
nand NAND2 (N7086, N7077, N556);
xor XOR2 (N7087, N7067, N1922);
xor XOR2 (N7088, N7083, N5568);
nand NAND2 (N7089, N7081, N3105);
buf BUF1 (N7090, N7086);
and AND2 (N7091, N7088, N7041);
not NOT1 (N7092, N7084);
xor XOR2 (N7093, N7085, N3113);
or OR4 (N7094, N7082, N4301, N5053, N6387);
or OR3 (N7095, N7069, N746, N2439);
nor NOR4 (N7096, N7095, N2748, N2145, N3974);
and AND2 (N7097, N7094, N4952);
buf BUF1 (N7098, N7092);
buf BUF1 (N7099, N7089);
nand NAND3 (N7100, N7079, N1797, N1593);
not NOT1 (N7101, N7096);
nand NAND3 (N7102, N7098, N1309, N701);
or OR3 (N7103, N7099, N2098, N5330);
nor NOR4 (N7104, N7093, N555, N3650, N2915);
not NOT1 (N7105, N7102);
not NOT1 (N7106, N7091);
buf BUF1 (N7107, N7105);
not NOT1 (N7108, N7075);
nor NOR2 (N7109, N7108, N2378);
and AND4 (N7110, N7107, N3425, N4981, N3969);
xor XOR2 (N7111, N7100, N6706);
and AND3 (N7112, N7103, N1144, N1591);
not NOT1 (N7113, N7110);
buf BUF1 (N7114, N7087);
nand NAND3 (N7115, N7111, N830, N64);
or OR2 (N7116, N7109, N519);
not NOT1 (N7117, N7106);
nor NOR2 (N7118, N7115, N5322);
nand NAND3 (N7119, N7104, N3956, N495);
and AND4 (N7120, N7112, N1111, N1815, N3117);
buf BUF1 (N7121, N7113);
xor XOR2 (N7122, N7097, N923);
or OR4 (N7123, N7118, N3857, N521, N1244);
or OR4 (N7124, N7116, N491, N3216, N5780);
xor XOR2 (N7125, N7121, N4311);
nand NAND4 (N7126, N7101, N1437, N2371, N1162);
buf BUF1 (N7127, N7122);
or OR4 (N7128, N7117, N7119, N3156, N1301);
nand NAND3 (N7129, N804, N2856, N4584);
or OR2 (N7130, N7090, N4499);
nand NAND2 (N7131, N7129, N4844);
not NOT1 (N7132, N7125);
nand NAND3 (N7133, N7120, N976, N578);
and AND3 (N7134, N7131, N1670, N3942);
xor XOR2 (N7135, N7123, N5104);
nor NOR2 (N7136, N7134, N889);
nor NOR4 (N7137, N7128, N4044, N4356, N1811);
and AND2 (N7138, N7124, N50);
and AND4 (N7139, N7135, N3628, N2531, N5973);
nor NOR3 (N7140, N7130, N2401, N1052);
buf BUF1 (N7141, N7132);
buf BUF1 (N7142, N7126);
buf BUF1 (N7143, N7133);
buf BUF1 (N7144, N7141);
buf BUF1 (N7145, N7143);
buf BUF1 (N7146, N7145);
not NOT1 (N7147, N7138);
and AND3 (N7148, N7137, N5129, N2163);
not NOT1 (N7149, N7148);
and AND2 (N7150, N7127, N2602);
and AND2 (N7151, N7142, N4382);
not NOT1 (N7152, N7147);
nand NAND4 (N7153, N7150, N6749, N6905, N4962);
xor XOR2 (N7154, N7139, N2747);
nor NOR4 (N7155, N7136, N3867, N4152, N2383);
or OR4 (N7156, N7153, N266, N5291, N376);
or OR2 (N7157, N7140, N3320);
xor XOR2 (N7158, N7151, N4700);
nand NAND4 (N7159, N7144, N2649, N2092, N5296);
nor NOR4 (N7160, N7152, N3400, N6194, N6307);
not NOT1 (N7161, N7154);
or OR2 (N7162, N7156, N3437);
or OR4 (N7163, N7149, N5092, N3278, N3743);
buf BUF1 (N7164, N7158);
not NOT1 (N7165, N7162);
buf BUF1 (N7166, N7160);
xor XOR2 (N7167, N7161, N4788);
nand NAND2 (N7168, N7159, N4343);
and AND3 (N7169, N7165, N2285, N6479);
buf BUF1 (N7170, N7168);
not NOT1 (N7171, N7155);
nand NAND3 (N7172, N7164, N6978, N1300);
nor NOR2 (N7173, N7167, N3677);
not NOT1 (N7174, N7169);
buf BUF1 (N7175, N7163);
or OR2 (N7176, N7171, N5285);
and AND3 (N7177, N7146, N2790, N6416);
xor XOR2 (N7178, N7172, N5252);
or OR3 (N7179, N7173, N1082, N2940);
nand NAND2 (N7180, N7174, N3324);
buf BUF1 (N7181, N7114);
or OR3 (N7182, N7166, N5370, N5538);
and AND4 (N7183, N7176, N4262, N625, N4413);
not NOT1 (N7184, N7179);
or OR4 (N7185, N7178, N375, N4524, N4684);
or OR4 (N7186, N7182, N5605, N3085, N1292);
nor NOR3 (N7187, N7157, N1179, N2079);
xor XOR2 (N7188, N7185, N6598);
xor XOR2 (N7189, N7184, N4348);
xor XOR2 (N7190, N7186, N3652);
nor NOR4 (N7191, N7181, N3325, N4868, N4513);
buf BUF1 (N7192, N7191);
nor NOR2 (N7193, N7175, N229);
and AND4 (N7194, N7192, N3956, N7064, N1575);
buf BUF1 (N7195, N7183);
and AND3 (N7196, N7190, N3308, N2146);
not NOT1 (N7197, N7189);
buf BUF1 (N7198, N7180);
or OR2 (N7199, N7198, N1592);
xor XOR2 (N7200, N7193, N807);
nor NOR2 (N7201, N7197, N4323);
nand NAND2 (N7202, N7194, N6647);
buf BUF1 (N7203, N7188);
buf BUF1 (N7204, N7203);
nand NAND4 (N7205, N7170, N116, N5059, N1569);
and AND3 (N7206, N7195, N6274, N6515);
or OR3 (N7207, N7205, N4242, N62);
not NOT1 (N7208, N7196);
nor NOR2 (N7209, N7177, N3898);
not NOT1 (N7210, N7202);
or OR3 (N7211, N7200, N915, N1201);
nor NOR3 (N7212, N7211, N3303, N5750);
nand NAND2 (N7213, N7212, N606);
buf BUF1 (N7214, N7204);
not NOT1 (N7215, N7213);
nand NAND2 (N7216, N7201, N4812);
and AND4 (N7217, N7187, N3765, N6366, N1739);
buf BUF1 (N7218, N7215);
and AND2 (N7219, N7214, N1880);
nand NAND3 (N7220, N7199, N2892, N6595);
and AND4 (N7221, N7217, N4607, N4898, N962);
buf BUF1 (N7222, N7210);
buf BUF1 (N7223, N7209);
nand NAND4 (N7224, N7222, N6983, N3983, N3554);
and AND2 (N7225, N7216, N888);
nor NOR2 (N7226, N7218, N5292);
not NOT1 (N7227, N7223);
not NOT1 (N7228, N7225);
buf BUF1 (N7229, N7227);
buf BUF1 (N7230, N7208);
or OR2 (N7231, N7229, N6115);
not NOT1 (N7232, N7231);
not NOT1 (N7233, N7207);
or OR3 (N7234, N7219, N1684, N6687);
nor NOR2 (N7235, N7232, N374);
nor NOR2 (N7236, N7224, N5628);
or OR4 (N7237, N7230, N5489, N5487, N71);
or OR2 (N7238, N7235, N4015);
nand NAND3 (N7239, N7238, N1336, N2231);
nand NAND4 (N7240, N7221, N255, N420, N5445);
buf BUF1 (N7241, N7228);
or OR3 (N7242, N7239, N1667, N2453);
not NOT1 (N7243, N7237);
xor XOR2 (N7244, N7241, N725);
or OR2 (N7245, N7226, N3711);
nand NAND3 (N7246, N7220, N6765, N3120);
nor NOR4 (N7247, N7240, N3102, N1210, N5731);
nor NOR3 (N7248, N7247, N1117, N6473);
and AND3 (N7249, N7206, N5421, N6216);
nand NAND3 (N7250, N7242, N6863, N2942);
xor XOR2 (N7251, N7246, N4605);
or OR4 (N7252, N7236, N1827, N1489, N6963);
buf BUF1 (N7253, N7250);
nand NAND2 (N7254, N7233, N3966);
not NOT1 (N7255, N7243);
and AND3 (N7256, N7254, N1747, N5843);
nor NOR3 (N7257, N7256, N3028, N258);
buf BUF1 (N7258, N7257);
or OR3 (N7259, N7245, N2617, N705);
not NOT1 (N7260, N7255);
nor NOR4 (N7261, N7248, N2758, N5157, N1087);
nor NOR3 (N7262, N7234, N1404, N3285);
or OR4 (N7263, N7261, N1326, N2271, N7082);
nor NOR3 (N7264, N7263, N4356, N3245);
nor NOR3 (N7265, N7252, N5231, N6429);
xor XOR2 (N7266, N7253, N5389);
or OR2 (N7267, N7249, N3200);
nand NAND4 (N7268, N7260, N457, N5685, N4990);
not NOT1 (N7269, N7264);
nor NOR2 (N7270, N7244, N6559);
xor XOR2 (N7271, N7266, N7146);
or OR2 (N7272, N7251, N1855);
buf BUF1 (N7273, N7271);
buf BUF1 (N7274, N7268);
not NOT1 (N7275, N7265);
xor XOR2 (N7276, N7269, N4893);
nand NAND2 (N7277, N7275, N3191);
buf BUF1 (N7278, N7277);
nor NOR2 (N7279, N7276, N5546);
nand NAND3 (N7280, N7267, N4744, N1475);
buf BUF1 (N7281, N7270);
and AND4 (N7282, N7274, N4444, N2345, N777);
nor NOR2 (N7283, N7262, N1379);
nor NOR3 (N7284, N7273, N3472, N3765);
or OR4 (N7285, N7272, N3524, N2948, N96);
buf BUF1 (N7286, N7283);
or OR4 (N7287, N7286, N1398, N1616, N969);
not NOT1 (N7288, N7284);
xor XOR2 (N7289, N7281, N5419);
nand NAND3 (N7290, N7279, N1017, N500);
buf BUF1 (N7291, N7285);
nand NAND4 (N7292, N7289, N6961, N2927, N3991);
not NOT1 (N7293, N7258);
buf BUF1 (N7294, N7292);
nor NOR2 (N7295, N7280, N4979);
buf BUF1 (N7296, N7259);
nand NAND2 (N7297, N7295, N3292);
not NOT1 (N7298, N7293);
buf BUF1 (N7299, N7296);
and AND2 (N7300, N7297, N5528);
nand NAND4 (N7301, N7298, N650, N1118, N5560);
buf BUF1 (N7302, N7290);
buf BUF1 (N7303, N7294);
and AND2 (N7304, N7300, N6529);
buf BUF1 (N7305, N7303);
nand NAND3 (N7306, N7305, N2939, N3306);
nand NAND3 (N7307, N7291, N177, N3906);
not NOT1 (N7308, N7306);
and AND4 (N7309, N7308, N1919, N289, N5028);
or OR3 (N7310, N7309, N1915, N7302);
nand NAND2 (N7311, N7082, N6802);
nand NAND4 (N7312, N7310, N6790, N3110, N5591);
buf BUF1 (N7313, N7304);
or OR3 (N7314, N7288, N3460, N5602);
or OR3 (N7315, N7287, N5746, N3518);
and AND3 (N7316, N7313, N3860, N4340);
xor XOR2 (N7317, N7312, N1647);
and AND2 (N7318, N7278, N1108);
nand NAND4 (N7319, N7317, N3802, N448, N4328);
nor NOR2 (N7320, N7307, N3896);
or OR2 (N7321, N7299, N6006);
not NOT1 (N7322, N7282);
nand NAND2 (N7323, N7322, N3666);
and AND2 (N7324, N7311, N3970);
and AND3 (N7325, N7316, N2918, N4437);
or OR4 (N7326, N7325, N2366, N4264, N4480);
and AND4 (N7327, N7315, N2494, N5368, N1519);
nor NOR4 (N7328, N7324, N2886, N7202, N4611);
or OR2 (N7329, N7301, N6154);
not NOT1 (N7330, N7319);
xor XOR2 (N7331, N7329, N2430);
not NOT1 (N7332, N7318);
xor XOR2 (N7333, N7320, N6001);
nor NOR2 (N7334, N7323, N2139);
not NOT1 (N7335, N7326);
not NOT1 (N7336, N7321);
not NOT1 (N7337, N7336);
or OR3 (N7338, N7330, N2521, N3353);
and AND4 (N7339, N7333, N1154, N1382, N2419);
nand NAND4 (N7340, N7338, N5121, N1774, N6120);
or OR3 (N7341, N7340, N7289, N7075);
nand NAND4 (N7342, N7328, N720, N2534, N2292);
or OR4 (N7343, N7327, N4622, N1655, N4381);
not NOT1 (N7344, N7335);
not NOT1 (N7345, N7314);
nand NAND2 (N7346, N7345, N3745);
nand NAND4 (N7347, N7343, N443, N4103, N6616);
or OR4 (N7348, N7332, N5495, N4349, N2612);
or OR3 (N7349, N7341, N4041, N2669);
xor XOR2 (N7350, N7337, N4415);
or OR4 (N7351, N7350, N4779, N4602, N2765);
xor XOR2 (N7352, N7342, N6883);
and AND4 (N7353, N7349, N778, N6289, N5165);
nor NOR2 (N7354, N7334, N5683);
and AND3 (N7355, N7352, N5343, N3754);
or OR3 (N7356, N7348, N3882, N3503);
buf BUF1 (N7357, N7354);
and AND2 (N7358, N7357, N5259);
buf BUF1 (N7359, N7344);
buf BUF1 (N7360, N7355);
nand NAND3 (N7361, N7353, N824, N1084);
or OR3 (N7362, N7347, N4868, N2837);
not NOT1 (N7363, N7361);
or OR2 (N7364, N7358, N6847);
xor XOR2 (N7365, N7364, N4267);
not NOT1 (N7366, N7351);
nand NAND3 (N7367, N7365, N5896, N3005);
nor NOR2 (N7368, N7360, N5472);
nand NAND4 (N7369, N7362, N1726, N285, N538);
nand NAND2 (N7370, N7331, N6444);
or OR3 (N7371, N7369, N4427, N3103);
buf BUF1 (N7372, N7368);
xor XOR2 (N7373, N7371, N7170);
not NOT1 (N7374, N7367);
buf BUF1 (N7375, N7370);
and AND3 (N7376, N7359, N5892, N2043);
and AND4 (N7377, N7346, N3923, N2631, N4653);
buf BUF1 (N7378, N7375);
nor NOR3 (N7379, N7378, N5647, N4029);
not NOT1 (N7380, N7363);
not NOT1 (N7381, N7374);
nor NOR3 (N7382, N7380, N3987, N1505);
or OR3 (N7383, N7356, N1213, N2948);
xor XOR2 (N7384, N7372, N214);
nor NOR4 (N7385, N7377, N1220, N4883, N4719);
not NOT1 (N7386, N7376);
or OR4 (N7387, N7384, N6621, N233, N3243);
nand NAND3 (N7388, N7383, N2197, N168);
and AND2 (N7389, N7385, N5162);
or OR4 (N7390, N7373, N3566, N5064, N5415);
nor NOR3 (N7391, N7386, N6884, N2272);
not NOT1 (N7392, N7391);
or OR3 (N7393, N7381, N4325, N6851);
xor XOR2 (N7394, N7390, N6874);
buf BUF1 (N7395, N7392);
not NOT1 (N7396, N7339);
or OR3 (N7397, N7366, N6029, N4712);
not NOT1 (N7398, N7394);
xor XOR2 (N7399, N7387, N1424);
xor XOR2 (N7400, N7379, N3222);
nor NOR4 (N7401, N7395, N6131, N3144, N5968);
nand NAND2 (N7402, N7401, N3677);
buf BUF1 (N7403, N7396);
not NOT1 (N7404, N7398);
not NOT1 (N7405, N7402);
xor XOR2 (N7406, N7397, N3108);
xor XOR2 (N7407, N7393, N1606);
nand NAND3 (N7408, N7388, N1932, N7375);
or OR2 (N7409, N7407, N7034);
nand NAND3 (N7410, N7400, N5521, N5950);
xor XOR2 (N7411, N7389, N6321);
buf BUF1 (N7412, N7406);
not NOT1 (N7413, N7408);
xor XOR2 (N7414, N7399, N6793);
xor XOR2 (N7415, N7403, N3666);
buf BUF1 (N7416, N7382);
or OR2 (N7417, N7410, N5415);
buf BUF1 (N7418, N7412);
nand NAND2 (N7419, N7414, N4075);
not NOT1 (N7420, N7418);
nand NAND3 (N7421, N7405, N7232, N3820);
or OR4 (N7422, N7409, N3330, N7240, N1351);
nor NOR4 (N7423, N7411, N4244, N5455, N5784);
buf BUF1 (N7424, N7417);
and AND2 (N7425, N7413, N1276);
or OR3 (N7426, N7421, N4790, N5095);
buf BUF1 (N7427, N7426);
not NOT1 (N7428, N7423);
not NOT1 (N7429, N7422);
nor NOR2 (N7430, N7416, N3541);
buf BUF1 (N7431, N7424);
nor NOR2 (N7432, N7404, N2123);
xor XOR2 (N7433, N7427, N3403);
or OR2 (N7434, N7433, N2295);
nor NOR2 (N7435, N7428, N5187);
or OR3 (N7436, N7430, N376, N3435);
buf BUF1 (N7437, N7415);
and AND2 (N7438, N7425, N5004);
nand NAND3 (N7439, N7432, N4844, N4736);
nor NOR3 (N7440, N7434, N6836, N278);
and AND4 (N7441, N7429, N4651, N5733, N4789);
nand NAND4 (N7442, N7431, N2287, N1925, N5899);
xor XOR2 (N7443, N7437, N1696);
xor XOR2 (N7444, N7443, N4943);
nor NOR3 (N7445, N7435, N1795, N4365);
and AND3 (N7446, N7442, N1117, N3733);
not NOT1 (N7447, N7446);
nand NAND2 (N7448, N7441, N3764);
xor XOR2 (N7449, N7436, N6211);
nor NOR2 (N7450, N7440, N3525);
or OR3 (N7451, N7447, N3604, N4549);
xor XOR2 (N7452, N7420, N4709);
xor XOR2 (N7453, N7452, N3638);
buf BUF1 (N7454, N7439);
and AND3 (N7455, N7451, N3427, N5663);
not NOT1 (N7456, N7438);
or OR3 (N7457, N7444, N6295, N7416);
nor NOR2 (N7458, N7450, N6308);
not NOT1 (N7459, N7454);
buf BUF1 (N7460, N7457);
or OR3 (N7461, N7445, N4864, N1646);
and AND4 (N7462, N7456, N5520, N982, N3079);
nor NOR4 (N7463, N7453, N2354, N2146, N5311);
buf BUF1 (N7464, N7461);
not NOT1 (N7465, N7460);
buf BUF1 (N7466, N7463);
or OR2 (N7467, N7462, N1512);
buf BUF1 (N7468, N7449);
or OR4 (N7469, N7419, N3718, N3722, N1202);
nor NOR2 (N7470, N7465, N2614);
nand NAND3 (N7471, N7459, N3893, N2587);
or OR2 (N7472, N7466, N6549);
buf BUF1 (N7473, N7455);
buf BUF1 (N7474, N7464);
nor NOR4 (N7475, N7469, N1287, N1438, N3804);
nor NOR2 (N7476, N7472, N6142);
buf BUF1 (N7477, N7476);
nor NOR2 (N7478, N7475, N7425);
xor XOR2 (N7479, N7448, N3808);
or OR3 (N7480, N7467, N1049, N3610);
or OR3 (N7481, N7479, N4875, N3537);
nor NOR2 (N7482, N7473, N6948);
nand NAND4 (N7483, N7471, N986, N1606, N1903);
or OR4 (N7484, N7470, N445, N2976, N4053);
not NOT1 (N7485, N7481);
xor XOR2 (N7486, N7458, N6746);
nand NAND3 (N7487, N7474, N2805, N4745);
nand NAND4 (N7488, N7477, N6462, N1715, N6965);
xor XOR2 (N7489, N7484, N6834);
and AND3 (N7490, N7482, N6854, N1087);
and AND2 (N7491, N7486, N3708);
nor NOR4 (N7492, N7483, N348, N386, N7261);
and AND4 (N7493, N7489, N6102, N4780, N3406);
nand NAND2 (N7494, N7493, N357);
not NOT1 (N7495, N7468);
nor NOR2 (N7496, N7490, N4651);
not NOT1 (N7497, N7480);
and AND3 (N7498, N7487, N6247, N1987);
not NOT1 (N7499, N7494);
or OR3 (N7500, N7499, N275, N562);
or OR2 (N7501, N7500, N6182);
and AND2 (N7502, N7495, N4290);
buf BUF1 (N7503, N7492);
or OR3 (N7504, N7478, N2123, N117);
xor XOR2 (N7505, N7497, N4877);
nor NOR3 (N7506, N7498, N5667, N3197);
nand NAND4 (N7507, N7506, N4409, N4052, N4927);
and AND2 (N7508, N7505, N2948);
and AND2 (N7509, N7488, N710);
xor XOR2 (N7510, N7509, N4689);
nand NAND4 (N7511, N7501, N6231, N2363, N3230);
and AND4 (N7512, N7507, N5691, N2766, N2867);
nor NOR4 (N7513, N7491, N7441, N1675, N4741);
buf BUF1 (N7514, N7513);
nor NOR3 (N7515, N7510, N6060, N553);
nand NAND3 (N7516, N7514, N3700, N1493);
and AND2 (N7517, N7503, N2162);
nor NOR3 (N7518, N7511, N7281, N5627);
nand NAND4 (N7519, N7516, N7360, N6224, N3699);
buf BUF1 (N7520, N7517);
xor XOR2 (N7521, N7485, N5639);
and AND2 (N7522, N7521, N6661);
not NOT1 (N7523, N7512);
not NOT1 (N7524, N7502);
buf BUF1 (N7525, N7508);
nor NOR2 (N7526, N7504, N2923);
and AND4 (N7527, N7526, N419, N4429, N4806);
not NOT1 (N7528, N7518);
and AND4 (N7529, N7525, N6526, N7373, N1826);
xor XOR2 (N7530, N7529, N484);
and AND2 (N7531, N7530, N4304);
buf BUF1 (N7532, N7524);
buf BUF1 (N7533, N7527);
nand NAND4 (N7534, N7531, N1111, N4124, N4594);
buf BUF1 (N7535, N7528);
nand NAND2 (N7536, N7535, N2398);
and AND2 (N7537, N7523, N205);
not NOT1 (N7538, N7496);
not NOT1 (N7539, N7534);
nand NAND2 (N7540, N7522, N6175);
not NOT1 (N7541, N7537);
xor XOR2 (N7542, N7533, N6566);
and AND2 (N7543, N7515, N5807);
nor NOR4 (N7544, N7536, N5048, N3277, N3644);
nor NOR2 (N7545, N7543, N1116);
nand NAND2 (N7546, N7545, N5437);
nor NOR3 (N7547, N7539, N1523, N2987);
or OR4 (N7548, N7520, N1765, N3104, N4714);
nor NOR3 (N7549, N7532, N852, N7469);
xor XOR2 (N7550, N7548, N6121);
nand NAND3 (N7551, N7519, N1441, N2906);
nor NOR3 (N7552, N7549, N2509, N7501);
not NOT1 (N7553, N7547);
and AND3 (N7554, N7553, N1502, N6849);
and AND4 (N7555, N7551, N4501, N2252, N4754);
and AND2 (N7556, N7552, N4029);
not NOT1 (N7557, N7540);
and AND3 (N7558, N7554, N1712, N2409);
nand NAND2 (N7559, N7555, N7005);
or OR4 (N7560, N7542, N3332, N1266, N1468);
xor XOR2 (N7561, N7550, N4609);
nor NOR2 (N7562, N7544, N4371);
or OR2 (N7563, N7538, N4593);
buf BUF1 (N7564, N7557);
nor NOR4 (N7565, N7559, N103, N2189, N4619);
and AND2 (N7566, N7541, N916);
and AND4 (N7567, N7562, N1731, N1618, N1117);
and AND2 (N7568, N7560, N4413);
xor XOR2 (N7569, N7568, N5148);
nor NOR2 (N7570, N7565, N4663);
not NOT1 (N7571, N7563);
and AND4 (N7572, N7564, N6282, N4504, N7241);
nand NAND4 (N7573, N7556, N7239, N2412, N309);
buf BUF1 (N7574, N7558);
and AND3 (N7575, N7566, N3414, N6420);
buf BUF1 (N7576, N7574);
and AND2 (N7577, N7576, N4049);
buf BUF1 (N7578, N7569);
buf BUF1 (N7579, N7570);
nand NAND4 (N7580, N7579, N3680, N7215, N5225);
nand NAND4 (N7581, N7567, N4602, N6540, N6838);
nand NAND2 (N7582, N7573, N1101);
nor NOR4 (N7583, N7581, N774, N2308, N4295);
xor XOR2 (N7584, N7571, N458);
not NOT1 (N7585, N7578);
buf BUF1 (N7586, N7580);
and AND4 (N7587, N7582, N1022, N5212, N642);
nand NAND2 (N7588, N7575, N4692);
not NOT1 (N7589, N7584);
nand NAND4 (N7590, N7589, N514, N861, N565);
xor XOR2 (N7591, N7572, N1625);
and AND2 (N7592, N7587, N3028);
not NOT1 (N7593, N7561);
nor NOR4 (N7594, N7590, N2251, N4918, N4745);
not NOT1 (N7595, N7583);
xor XOR2 (N7596, N7588, N1305);
nor NOR4 (N7597, N7596, N6732, N4409, N7565);
nand NAND3 (N7598, N7585, N3714, N4498);
xor XOR2 (N7599, N7591, N1803);
nor NOR4 (N7600, N7595, N932, N3950, N2973);
buf BUF1 (N7601, N7577);
xor XOR2 (N7602, N7593, N1592);
not NOT1 (N7603, N7600);
nor NOR2 (N7604, N7546, N5771);
and AND3 (N7605, N7597, N5360, N5507);
buf BUF1 (N7606, N7602);
nand NAND4 (N7607, N7603, N5491, N7162, N4278);
nor NOR2 (N7608, N7598, N816);
or OR2 (N7609, N7594, N294);
or OR2 (N7610, N7604, N3609);
and AND4 (N7611, N7601, N5277, N6150, N6222);
nor NOR2 (N7612, N7607, N817);
nor NOR2 (N7613, N7611, N6049);
not NOT1 (N7614, N7609);
buf BUF1 (N7615, N7612);
nand NAND3 (N7616, N7613, N7436, N3774);
xor XOR2 (N7617, N7605, N3948);
or OR2 (N7618, N7599, N1461);
buf BUF1 (N7619, N7617);
or OR3 (N7620, N7618, N2905, N6377);
not NOT1 (N7621, N7615);
or OR3 (N7622, N7621, N1412, N7033);
and AND2 (N7623, N7610, N2940);
nor NOR4 (N7624, N7616, N304, N836, N4373);
or OR4 (N7625, N7592, N324, N5381, N3401);
not NOT1 (N7626, N7608);
nor NOR2 (N7627, N7614, N4244);
nor NOR4 (N7628, N7619, N5504, N5688, N1651);
nand NAND4 (N7629, N7625, N509, N993, N7393);
nor NOR3 (N7630, N7622, N6877, N6033);
not NOT1 (N7631, N7627);
nor NOR2 (N7632, N7586, N5864);
not NOT1 (N7633, N7620);
xor XOR2 (N7634, N7631, N6754);
or OR4 (N7635, N7606, N5190, N7390, N8);
or OR4 (N7636, N7635, N4908, N7374, N6769);
not NOT1 (N7637, N7633);
nand NAND2 (N7638, N7630, N872);
or OR3 (N7639, N7624, N7609, N5965);
nor NOR3 (N7640, N7637, N6887, N851);
nand NAND2 (N7641, N7632, N1783);
xor XOR2 (N7642, N7623, N255);
and AND4 (N7643, N7628, N3882, N5453, N6586);
xor XOR2 (N7644, N7640, N3964);
nor NOR3 (N7645, N7641, N7234, N7347);
nand NAND3 (N7646, N7629, N7639, N7446);
or OR3 (N7647, N4655, N1584, N3690);
nor NOR4 (N7648, N7647, N4774, N3717, N1653);
and AND3 (N7649, N7648, N563, N4172);
not NOT1 (N7650, N7649);
xor XOR2 (N7651, N7645, N4007);
nor NOR4 (N7652, N7634, N966, N1463, N6818);
nand NAND2 (N7653, N7646, N6501);
and AND4 (N7654, N7651, N3386, N4676, N4384);
buf BUF1 (N7655, N7652);
and AND2 (N7656, N7638, N1596);
and AND2 (N7657, N7656, N1702);
xor XOR2 (N7658, N7642, N1475);
and AND3 (N7659, N7658, N544, N5445);
not NOT1 (N7660, N7650);
and AND2 (N7661, N7657, N818);
xor XOR2 (N7662, N7660, N951);
buf BUF1 (N7663, N7636);
nand NAND3 (N7664, N7659, N1648, N6815);
or OR2 (N7665, N7662, N7311);
buf BUF1 (N7666, N7664);
nor NOR3 (N7667, N7654, N5937, N5549);
xor XOR2 (N7668, N7653, N5666);
and AND4 (N7669, N7644, N3849, N5641, N3709);
or OR4 (N7670, N7668, N6660, N4595, N4243);
buf BUF1 (N7671, N7655);
and AND4 (N7672, N7665, N6790, N6512, N7023);
buf BUF1 (N7673, N7643);
buf BUF1 (N7674, N7670);
and AND2 (N7675, N7673, N1092);
xor XOR2 (N7676, N7666, N2905);
buf BUF1 (N7677, N7676);
and AND3 (N7678, N7675, N6811, N6854);
not NOT1 (N7679, N7672);
xor XOR2 (N7680, N7677, N2186);
or OR4 (N7681, N7674, N4038, N5169, N6800);
xor XOR2 (N7682, N7681, N831);
xor XOR2 (N7683, N7663, N4543);
nor NOR2 (N7684, N7626, N5423);
not NOT1 (N7685, N7661);
and AND2 (N7686, N7679, N2185);
nand NAND4 (N7687, N7680, N6129, N7296, N2024);
not NOT1 (N7688, N7669);
and AND3 (N7689, N7684, N2865, N7302);
and AND4 (N7690, N7667, N787, N7530, N5419);
nor NOR2 (N7691, N7688, N701);
not NOT1 (N7692, N7687);
buf BUF1 (N7693, N7690);
nand NAND4 (N7694, N7686, N6053, N1393, N6390);
not NOT1 (N7695, N7682);
or OR4 (N7696, N7691, N631, N2865, N6106);
not NOT1 (N7697, N7685);
and AND4 (N7698, N7678, N4393, N3206, N5770);
xor XOR2 (N7699, N7683, N5555);
xor XOR2 (N7700, N7697, N6670);
or OR3 (N7701, N7695, N5831, N2891);
or OR2 (N7702, N7700, N420);
nand NAND4 (N7703, N7701, N5552, N4740, N5292);
and AND4 (N7704, N7671, N3209, N4929, N3427);
not NOT1 (N7705, N7703);
buf BUF1 (N7706, N7699);
buf BUF1 (N7707, N7692);
and AND4 (N7708, N7706, N1006, N3146, N2984);
or OR2 (N7709, N7698, N6440);
nor NOR4 (N7710, N7696, N4702, N2302, N7415);
buf BUF1 (N7711, N7704);
nand NAND4 (N7712, N7689, N7351, N6788, N65);
nor NOR4 (N7713, N7710, N6411, N6887, N5697);
and AND4 (N7714, N7709, N6070, N6305, N2185);
nand NAND4 (N7715, N7714, N2154, N2469, N2636);
nand NAND2 (N7716, N7694, N3512);
buf BUF1 (N7717, N7705);
or OR3 (N7718, N7717, N2144, N6072);
buf BUF1 (N7719, N7702);
and AND2 (N7720, N7712, N6166);
nor NOR3 (N7721, N7711, N6268, N6592);
and AND4 (N7722, N7715, N7366, N5633, N6683);
not NOT1 (N7723, N7721);
xor XOR2 (N7724, N7716, N369);
nand NAND3 (N7725, N7720, N6768, N1278);
nand NAND4 (N7726, N7724, N2094, N5647, N1110);
or OR3 (N7727, N7719, N60, N6178);
not NOT1 (N7728, N7718);
not NOT1 (N7729, N7727);
not NOT1 (N7730, N7722);
or OR2 (N7731, N7723, N6082);
xor XOR2 (N7732, N7728, N4825);
nand NAND3 (N7733, N7708, N5577, N38);
and AND2 (N7734, N7726, N393);
xor XOR2 (N7735, N7713, N2042);
not NOT1 (N7736, N7732);
buf BUF1 (N7737, N7734);
and AND3 (N7738, N7733, N3408, N5881);
xor XOR2 (N7739, N7730, N4531);
buf BUF1 (N7740, N7739);
buf BUF1 (N7741, N7725);
not NOT1 (N7742, N7741);
nand NAND4 (N7743, N7707, N5569, N5423, N3630);
buf BUF1 (N7744, N7693);
buf BUF1 (N7745, N7735);
or OR3 (N7746, N7731, N7617, N6849);
buf BUF1 (N7747, N7743);
nand NAND3 (N7748, N7747, N3352, N3278);
nor NOR3 (N7749, N7746, N2168, N4729);
and AND3 (N7750, N7738, N6862, N7649);
and AND2 (N7751, N7737, N2103);
or OR4 (N7752, N7744, N4662, N6884, N5859);
nor NOR3 (N7753, N7740, N4110, N6974);
buf BUF1 (N7754, N7749);
xor XOR2 (N7755, N7752, N7456);
and AND2 (N7756, N7754, N4962);
nor NOR3 (N7757, N7756, N5574, N5375);
not NOT1 (N7758, N7753);
xor XOR2 (N7759, N7757, N1323);
nand NAND3 (N7760, N7745, N775, N744);
nor NOR4 (N7761, N7751, N4967, N870, N879);
or OR4 (N7762, N7729, N1737, N2443, N6627);
or OR4 (N7763, N7755, N6244, N3409, N64);
not NOT1 (N7764, N7759);
nor NOR4 (N7765, N7760, N6851, N3674, N558);
not NOT1 (N7766, N7762);
xor XOR2 (N7767, N7736, N200);
and AND2 (N7768, N7761, N4148);
buf BUF1 (N7769, N7758);
xor XOR2 (N7770, N7765, N3880);
nor NOR2 (N7771, N7764, N3252);
or OR2 (N7772, N7767, N4348);
or OR3 (N7773, N7770, N6570, N6703);
and AND3 (N7774, N7773, N3287, N5457);
buf BUF1 (N7775, N7766);
and AND4 (N7776, N7768, N2877, N4754, N7116);
not NOT1 (N7777, N7750);
nor NOR2 (N7778, N7772, N3353);
nand NAND3 (N7779, N7775, N1043, N591);
nor NOR2 (N7780, N7748, N1130);
not NOT1 (N7781, N7780);
and AND4 (N7782, N7769, N1282, N1243, N1848);
or OR3 (N7783, N7777, N4988, N872);
not NOT1 (N7784, N7771);
nor NOR4 (N7785, N7779, N4657, N4458, N6778);
or OR4 (N7786, N7742, N2376, N4713, N1516);
not NOT1 (N7787, N7763);
and AND4 (N7788, N7784, N7324, N932, N1589);
not NOT1 (N7789, N7786);
xor XOR2 (N7790, N7788, N1259);
nand NAND3 (N7791, N7776, N6399, N5280);
not NOT1 (N7792, N7781);
or OR3 (N7793, N7774, N5789, N664);
or OR3 (N7794, N7792, N3448, N7261);
xor XOR2 (N7795, N7783, N351);
nand NAND3 (N7796, N7791, N1535, N2505);
buf BUF1 (N7797, N7787);
nand NAND4 (N7798, N7794, N275, N6742, N6420);
or OR2 (N7799, N7797, N6140);
and AND4 (N7800, N7799, N2754, N179, N6879);
nor NOR2 (N7801, N7796, N7256);
nand NAND2 (N7802, N7793, N4439);
buf BUF1 (N7803, N7798);
buf BUF1 (N7804, N7802);
nor NOR3 (N7805, N7795, N1961, N3066);
nand NAND2 (N7806, N7789, N4704);
nand NAND2 (N7807, N7806, N6274);
nand NAND3 (N7808, N7807, N2568, N5909);
nor NOR4 (N7809, N7801, N2959, N5611, N1189);
not NOT1 (N7810, N7805);
xor XOR2 (N7811, N7785, N556);
not NOT1 (N7812, N7803);
nand NAND4 (N7813, N7809, N6941, N4379, N455);
not NOT1 (N7814, N7800);
buf BUF1 (N7815, N7810);
nor NOR4 (N7816, N7815, N2833, N7103, N4053);
not NOT1 (N7817, N7813);
or OR4 (N7818, N7814, N3855, N5707, N1476);
nand NAND4 (N7819, N7811, N4865, N241, N1670);
or OR2 (N7820, N7812, N3860);
or OR4 (N7821, N7820, N2108, N1486, N7420);
xor XOR2 (N7822, N7818, N3042);
nand NAND4 (N7823, N7819, N7704, N2898, N1527);
or OR4 (N7824, N7816, N6736, N6060, N902);
and AND2 (N7825, N7778, N214);
not NOT1 (N7826, N7790);
and AND3 (N7827, N7825, N4172, N836);
nor NOR4 (N7828, N7822, N1855, N4618, N5430);
nand NAND3 (N7829, N7821, N5158, N2625);
and AND3 (N7830, N7824, N7540, N1350);
not NOT1 (N7831, N7827);
not NOT1 (N7832, N7830);
or OR4 (N7833, N7808, N7814, N503, N5335);
not NOT1 (N7834, N7833);
or OR3 (N7835, N7826, N2058, N5427);
and AND4 (N7836, N7835, N4313, N5693, N5531);
nor NOR3 (N7837, N7836, N506, N3117);
or OR2 (N7838, N7829, N5439);
or OR3 (N7839, N7828, N6397, N7818);
not NOT1 (N7840, N7823);
nor NOR4 (N7841, N7782, N19, N6890, N7568);
nor NOR2 (N7842, N7831, N7657);
not NOT1 (N7843, N7804);
and AND3 (N7844, N7839, N5458, N6741);
nand NAND3 (N7845, N7840, N3207, N181);
nand NAND2 (N7846, N7832, N7160);
xor XOR2 (N7847, N7838, N2306);
not NOT1 (N7848, N7847);
and AND4 (N7849, N7834, N1399, N650, N3052);
not NOT1 (N7850, N7841);
nand NAND3 (N7851, N7850, N2178, N1610);
nand NAND4 (N7852, N7843, N4400, N1495, N3504);
nor NOR3 (N7853, N7848, N6471, N4325);
not NOT1 (N7854, N7842);
nand NAND3 (N7855, N7837, N3552, N1481);
buf BUF1 (N7856, N7855);
nand NAND4 (N7857, N7844, N5143, N3968, N4872);
nor NOR4 (N7858, N7852, N735, N7600, N778);
not NOT1 (N7859, N7845);
or OR4 (N7860, N7857, N2404, N3668, N529);
not NOT1 (N7861, N7856);
not NOT1 (N7862, N7849);
or OR4 (N7863, N7862, N805, N5180, N1057);
xor XOR2 (N7864, N7859, N6357);
and AND2 (N7865, N7858, N925);
or OR4 (N7866, N7860, N2782, N3916, N6656);
nand NAND2 (N7867, N7817, N7723);
nor NOR2 (N7868, N7863, N4653);
or OR3 (N7869, N7854, N2583, N6051);
and AND3 (N7870, N7853, N49, N589);
not NOT1 (N7871, N7864);
xor XOR2 (N7872, N7870, N5155);
nand NAND2 (N7873, N7865, N7196);
buf BUF1 (N7874, N7861);
nor NOR3 (N7875, N7866, N7767, N2424);
and AND3 (N7876, N7873, N681, N2454);
or OR2 (N7877, N7851, N7215);
nand NAND4 (N7878, N7846, N5410, N2910, N2222);
xor XOR2 (N7879, N7867, N1114);
xor XOR2 (N7880, N7879, N3089);
and AND2 (N7881, N7869, N845);
xor XOR2 (N7882, N7880, N684);
not NOT1 (N7883, N7877);
nor NOR3 (N7884, N7883, N3154, N1393);
buf BUF1 (N7885, N7884);
and AND4 (N7886, N7881, N7771, N148, N3305);
and AND2 (N7887, N7878, N4919);
nor NOR3 (N7888, N7875, N188, N5167);
buf BUF1 (N7889, N7885);
xor XOR2 (N7890, N7887, N3396);
nand NAND4 (N7891, N7876, N5134, N4494, N3438);
nor NOR4 (N7892, N7871, N2813, N3198, N4511);
not NOT1 (N7893, N7889);
buf BUF1 (N7894, N7891);
nor NOR3 (N7895, N7874, N5777, N942);
xor XOR2 (N7896, N7872, N4193);
nand NAND3 (N7897, N7886, N5052, N2079);
and AND3 (N7898, N7897, N6077, N14);
nand NAND3 (N7899, N7893, N1471, N1613);
not NOT1 (N7900, N7892);
or OR2 (N7901, N7898, N3564);
buf BUF1 (N7902, N7895);
or OR2 (N7903, N7902, N4141);
buf BUF1 (N7904, N7888);
buf BUF1 (N7905, N7899);
and AND3 (N7906, N7901, N7738, N4143);
nand NAND3 (N7907, N7894, N172, N6020);
nand NAND4 (N7908, N7900, N3886, N3703, N6094);
buf BUF1 (N7909, N7906);
nor NOR3 (N7910, N7908, N7168, N2238);
or OR3 (N7911, N7909, N7110, N6670);
and AND2 (N7912, N7868, N3796);
not NOT1 (N7913, N7911);
buf BUF1 (N7914, N7904);
not NOT1 (N7915, N7910);
not NOT1 (N7916, N7907);
and AND4 (N7917, N7916, N1463, N2960, N1508);
xor XOR2 (N7918, N7915, N6396);
and AND3 (N7919, N7890, N1771, N4150);
nor NOR4 (N7920, N7912, N5341, N1334, N7207);
or OR3 (N7921, N7919, N6500, N3622);
xor XOR2 (N7922, N7921, N4474);
buf BUF1 (N7923, N7922);
nand NAND4 (N7924, N7918, N3094, N7017, N4827);
or OR4 (N7925, N7905, N7459, N1354, N7674);
nand NAND3 (N7926, N7924, N3011, N5);
nand NAND3 (N7927, N7913, N5402, N4107);
nor NOR3 (N7928, N7925, N7663, N1645);
buf BUF1 (N7929, N7926);
xor XOR2 (N7930, N7923, N5744);
nand NAND2 (N7931, N7896, N5021);
nor NOR4 (N7932, N7929, N1329, N6047, N1220);
and AND4 (N7933, N7882, N1577, N5014, N6283);
and AND2 (N7934, N7903, N3923);
nand NAND4 (N7935, N7920, N3587, N3903, N4612);
not NOT1 (N7936, N7931);
nor NOR2 (N7937, N7934, N623);
buf BUF1 (N7938, N7935);
or OR4 (N7939, N7933, N7882, N3436, N791);
not NOT1 (N7940, N7930);
nand NAND4 (N7941, N7936, N7434, N1295, N4877);
and AND4 (N7942, N7927, N6338, N7941, N7167);
and AND2 (N7943, N3698, N591);
xor XOR2 (N7944, N7917, N7844);
not NOT1 (N7945, N7928);
xor XOR2 (N7946, N7940, N2317);
buf BUF1 (N7947, N7942);
xor XOR2 (N7948, N7946, N1506);
or OR4 (N7949, N7943, N3473, N4735, N7686);
or OR4 (N7950, N7947, N7809, N6830, N4438);
or OR4 (N7951, N7949, N5492, N524, N4929);
xor XOR2 (N7952, N7937, N1192);
nand NAND4 (N7953, N7939, N3562, N347, N3402);
nor NOR2 (N7954, N7945, N3886);
xor XOR2 (N7955, N7951, N2552);
and AND4 (N7956, N7948, N2075, N1117, N6460);
and AND3 (N7957, N7914, N2690, N7334);
and AND2 (N7958, N7954, N4962);
xor XOR2 (N7959, N7932, N5119);
buf BUF1 (N7960, N7958);
xor XOR2 (N7961, N7950, N5075);
xor XOR2 (N7962, N7959, N4410);
buf BUF1 (N7963, N7952);
nor NOR4 (N7964, N7953, N3136, N4190, N1715);
or OR3 (N7965, N7964, N4226, N3643);
not NOT1 (N7966, N7960);
xor XOR2 (N7967, N7963, N5750);
or OR3 (N7968, N7961, N6577, N2120);
buf BUF1 (N7969, N7956);
and AND4 (N7970, N7938, N1585, N706, N617);
not NOT1 (N7971, N7966);
nand NAND2 (N7972, N7969, N7836);
nand NAND4 (N7973, N7972, N1293, N3249, N4975);
nor NOR3 (N7974, N7955, N1361, N5393);
xor XOR2 (N7975, N7962, N3465);
buf BUF1 (N7976, N7944);
not NOT1 (N7977, N7971);
nor NOR4 (N7978, N7977, N6247, N4118, N3268);
xor XOR2 (N7979, N7978, N4458);
nor NOR2 (N7980, N7957, N1004);
nand NAND2 (N7981, N7965, N4061);
xor XOR2 (N7982, N7980, N6775);
nand NAND2 (N7983, N7976, N1183);
xor XOR2 (N7984, N7973, N6689);
not NOT1 (N7985, N7983);
buf BUF1 (N7986, N7985);
not NOT1 (N7987, N7968);
or OR2 (N7988, N7979, N5040);
buf BUF1 (N7989, N7967);
nand NAND2 (N7990, N7975, N937);
not NOT1 (N7991, N7989);
nand NAND3 (N7992, N7991, N6965, N5328);
nor NOR4 (N7993, N7987, N6435, N2161, N3993);
buf BUF1 (N7994, N7993);
nor NOR3 (N7995, N7986, N2816, N6055);
nor NOR2 (N7996, N7988, N7742);
or OR4 (N7997, N7990, N943, N3601, N5650);
or OR4 (N7998, N7994, N4989, N1979, N6984);
not NOT1 (N7999, N7996);
buf BUF1 (N8000, N7999);
nor NOR4 (N8001, N7982, N1711, N5051, N6638);
xor XOR2 (N8002, N8001, N2053);
and AND3 (N8003, N8002, N527, N1048);
buf BUF1 (N8004, N7992);
nor NOR4 (N8005, N7998, N3863, N7718, N3225);
nor NOR3 (N8006, N7997, N1892, N2414);
nor NOR4 (N8007, N8003, N4265, N1382, N6221);
not NOT1 (N8008, N7974);
nor NOR3 (N8009, N8007, N4932, N4747);
not NOT1 (N8010, N8000);
nor NOR2 (N8011, N8008, N632);
and AND2 (N8012, N8009, N1418);
nor NOR4 (N8013, N7995, N7297, N6204, N1920);
nand NAND4 (N8014, N8004, N1819, N7961, N6074);
or OR2 (N8015, N7970, N4464);
buf BUF1 (N8016, N8014);
nand NAND3 (N8017, N8006, N426, N4089);
nand NAND4 (N8018, N8013, N2752, N5503, N2628);
nor NOR2 (N8019, N8015, N4521);
and AND3 (N8020, N8016, N6036, N5893);
endmodule