// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18;

output N1003,N1014,N991,N1011,N1009,N1015,N1016,N1013,N986,N1018;

and AND3 (N19, N17, N17, N4);
not NOT1 (N20, N2);
not NOT1 (N21, N16);
or OR3 (N22, N4, N12, N13);
and AND3 (N23, N20, N3, N20);
and AND2 (N24, N19, N1);
or OR3 (N25, N14, N10, N13);
xor XOR2 (N26, N15, N9);
and AND4 (N27, N16, N5, N18, N8);
xor XOR2 (N28, N8, N18);
and AND3 (N29, N10, N28, N26);
not NOT1 (N30, N9);
not NOT1 (N31, N27);
buf BUF1 (N32, N26);
and AND2 (N33, N26, N13);
nor NOR4 (N34, N32, N2, N15, N21);
buf BUF1 (N35, N18);
or OR4 (N36, N25, N4, N11, N28);
nand NAND4 (N37, N29, N24, N12, N11);
nand NAND3 (N38, N10, N10, N32);
not NOT1 (N39, N38);
and AND3 (N40, N39, N29, N2);
nor NOR3 (N41, N31, N10, N15);
nor NOR2 (N42, N40, N8);
not NOT1 (N43, N34);
or OR3 (N44, N41, N19, N22);
nand NAND3 (N45, N8, N20, N5);
not NOT1 (N46, N33);
and AND2 (N47, N30, N23);
nand NAND4 (N48, N14, N46, N1, N8);
buf BUF1 (N49, N46);
and AND2 (N50, N36, N10);
buf BUF1 (N51, N43);
or OR2 (N52, N37, N11);
nand NAND3 (N53, N35, N45, N9);
nand NAND2 (N54, N25, N12);
or OR2 (N55, N51, N33);
nand NAND2 (N56, N50, N25);
nor NOR4 (N57, N44, N33, N17, N35);
nor NOR2 (N58, N47, N5);
nand NAND4 (N59, N54, N34, N45, N25);
nor NOR2 (N60, N49, N37);
and AND3 (N61, N59, N37, N51);
and AND2 (N62, N60, N43);
and AND3 (N63, N61, N44, N47);
nor NOR2 (N64, N42, N47);
and AND4 (N65, N64, N20, N30, N44);
not NOT1 (N66, N65);
not NOT1 (N67, N66);
and AND4 (N68, N67, N44, N39, N16);
or OR4 (N69, N55, N20, N27, N3);
not NOT1 (N70, N63);
buf BUF1 (N71, N53);
xor XOR2 (N72, N71, N25);
nand NAND4 (N73, N57, N36, N27, N46);
buf BUF1 (N74, N48);
xor XOR2 (N75, N70, N55);
not NOT1 (N76, N72);
or OR2 (N77, N76, N74);
and AND3 (N78, N29, N27, N12);
nand NAND4 (N79, N56, N45, N29, N15);
buf BUF1 (N80, N62);
or OR3 (N81, N78, N47, N31);
buf BUF1 (N82, N58);
nor NOR2 (N83, N52, N81);
or OR3 (N84, N70, N79, N56);
or OR2 (N85, N3, N42);
or OR4 (N86, N82, N1, N74, N31);
and AND2 (N87, N80, N85);
nor NOR4 (N88, N25, N71, N56, N5);
nand NAND2 (N89, N68, N66);
nand NAND3 (N90, N83, N35, N15);
nand NAND2 (N91, N88, N83);
buf BUF1 (N92, N73);
nand NAND4 (N93, N90, N36, N50, N64);
or OR4 (N94, N77, N75, N72, N67);
nand NAND4 (N95, N84, N21, N58, N10);
or OR4 (N96, N66, N61, N7, N72);
not NOT1 (N97, N96);
xor XOR2 (N98, N91, N13);
not NOT1 (N99, N93);
not NOT1 (N100, N69);
or OR2 (N101, N98, N10);
not NOT1 (N102, N89);
not NOT1 (N103, N94);
and AND3 (N104, N103, N20, N36);
not NOT1 (N105, N104);
and AND4 (N106, N95, N5, N97, N42);
nand NAND3 (N107, N61, N103, N28);
and AND3 (N108, N101, N100, N52);
and AND4 (N109, N37, N107, N34, N1);
or OR2 (N110, N32, N87);
or OR4 (N111, N95, N2, N3, N98);
not NOT1 (N112, N92);
or OR3 (N113, N102, N108, N50);
not NOT1 (N114, N19);
or OR2 (N115, N112, N107);
xor XOR2 (N116, N99, N43);
nand NAND3 (N117, N105, N10, N15);
or OR4 (N118, N117, N16, N70, N51);
and AND3 (N119, N109, N33, N51);
or OR3 (N120, N111, N46, N42);
or OR3 (N121, N120, N42, N1);
nor NOR2 (N122, N116, N119);
and AND4 (N123, N113, N14, N114, N109);
nor NOR2 (N124, N15, N36);
buf BUF1 (N125, N29);
xor XOR2 (N126, N125, N21);
xor XOR2 (N127, N123, N3);
not NOT1 (N128, N115);
not NOT1 (N129, N118);
and AND2 (N130, N128, N24);
xor XOR2 (N131, N130, N4);
buf BUF1 (N132, N106);
and AND4 (N133, N129, N3, N123, N24);
nor NOR2 (N134, N110, N23);
and AND2 (N135, N122, N105);
and AND4 (N136, N133, N49, N109, N35);
nor NOR3 (N137, N126, N74, N126);
nand NAND3 (N138, N132, N55, N74);
not NOT1 (N139, N121);
and AND4 (N140, N124, N81, N64, N61);
and AND2 (N141, N136, N103);
nor NOR3 (N142, N86, N57, N47);
buf BUF1 (N143, N139);
or OR3 (N144, N135, N126, N37);
not NOT1 (N145, N140);
and AND4 (N146, N143, N116, N45, N46);
nor NOR3 (N147, N131, N127, N128);
and AND3 (N148, N63, N140, N19);
or OR2 (N149, N146, N83);
buf BUF1 (N150, N141);
xor XOR2 (N151, N148, N42);
nand NAND4 (N152, N151, N136, N49, N143);
and AND4 (N153, N137, N64, N55, N138);
nand NAND2 (N154, N111, N47);
nand NAND4 (N155, N145, N105, N51, N83);
nor NOR3 (N156, N154, N42, N98);
and AND4 (N157, N153, N88, N128, N118);
buf BUF1 (N158, N149);
nand NAND4 (N159, N150, N61, N116, N151);
buf BUF1 (N160, N142);
buf BUF1 (N161, N158);
and AND3 (N162, N157, N157, N107);
nand NAND4 (N163, N162, N56, N158, N63);
xor XOR2 (N164, N160, N37);
buf BUF1 (N165, N164);
or OR3 (N166, N147, N27, N153);
not NOT1 (N167, N163);
or OR3 (N168, N134, N8, N41);
not NOT1 (N169, N155);
or OR2 (N170, N167, N159);
or OR2 (N171, N24, N168);
nand NAND3 (N172, N116, N34, N85);
or OR2 (N173, N161, N47);
not NOT1 (N174, N169);
and AND4 (N175, N152, N150, N30, N125);
buf BUF1 (N176, N170);
nand NAND4 (N177, N171, N156, N82, N109);
nor NOR4 (N178, N48, N132, N11, N42);
and AND3 (N179, N172, N124, N139);
not NOT1 (N180, N175);
nand NAND2 (N181, N166, N173);
xor XOR2 (N182, N143, N127);
not NOT1 (N183, N180);
nor NOR4 (N184, N165, N113, N24, N37);
or OR2 (N185, N177, N110);
nor NOR4 (N186, N176, N88, N180, N84);
xor XOR2 (N187, N183, N73);
and AND3 (N188, N186, N65, N40);
nand NAND2 (N189, N174, N156);
xor XOR2 (N190, N181, N180);
xor XOR2 (N191, N182, N186);
nand NAND2 (N192, N185, N111);
or OR4 (N193, N184, N181, N76, N71);
and AND3 (N194, N179, N143, N47);
not NOT1 (N195, N188);
nand NAND4 (N196, N178, N123, N78, N128);
xor XOR2 (N197, N194, N184);
or OR4 (N198, N189, N165, N1, N5);
not NOT1 (N199, N191);
xor XOR2 (N200, N197, N4);
not NOT1 (N201, N196);
nand NAND2 (N202, N198, N80);
or OR3 (N203, N200, N92, N99);
buf BUF1 (N204, N193);
and AND2 (N205, N201, N140);
or OR2 (N206, N187, N193);
buf BUF1 (N207, N202);
and AND4 (N208, N206, N184, N85, N22);
xor XOR2 (N209, N144, N10);
and AND3 (N210, N199, N27, N74);
not NOT1 (N211, N190);
not NOT1 (N212, N207);
not NOT1 (N213, N204);
nand NAND4 (N214, N211, N67, N56, N36);
nor NOR3 (N215, N212, N63, N139);
buf BUF1 (N216, N192);
not NOT1 (N217, N215);
not NOT1 (N218, N214);
xor XOR2 (N219, N205, N30);
and AND3 (N220, N219, N180, N189);
nor NOR2 (N221, N203, N33);
buf BUF1 (N222, N216);
or OR4 (N223, N213, N97, N83, N206);
xor XOR2 (N224, N217, N77);
buf BUF1 (N225, N210);
nor NOR4 (N226, N224, N27, N131, N69);
and AND4 (N227, N221, N8, N52, N68);
or OR3 (N228, N226, N29, N150);
or OR3 (N229, N220, N131, N8);
or OR2 (N230, N227, N220);
not NOT1 (N231, N209);
not NOT1 (N232, N225);
nand NAND4 (N233, N230, N117, N171, N184);
nor NOR2 (N234, N223, N2);
nand NAND2 (N235, N232, N53);
or OR3 (N236, N228, N187, N73);
or OR4 (N237, N234, N66, N194, N201);
and AND4 (N238, N208, N27, N137, N217);
not NOT1 (N239, N235);
buf BUF1 (N240, N195);
not NOT1 (N241, N240);
xor XOR2 (N242, N231, N87);
buf BUF1 (N243, N237);
and AND4 (N244, N242, N107, N150, N28);
not NOT1 (N245, N222);
or OR4 (N246, N244, N28, N60, N102);
not NOT1 (N247, N229);
xor XOR2 (N248, N233, N63);
buf BUF1 (N249, N239);
buf BUF1 (N250, N236);
nor NOR4 (N251, N241, N133, N25, N183);
nand NAND3 (N252, N243, N111, N134);
or OR4 (N253, N245, N208, N215, N72);
nor NOR3 (N254, N246, N167, N113);
xor XOR2 (N255, N252, N245);
xor XOR2 (N256, N254, N185);
xor XOR2 (N257, N218, N78);
nand NAND2 (N258, N249, N202);
buf BUF1 (N259, N251);
xor XOR2 (N260, N258, N247);
nand NAND3 (N261, N124, N3, N62);
or OR2 (N262, N259, N177);
nand NAND3 (N263, N248, N224, N68);
nand NAND2 (N264, N261, N39);
and AND2 (N265, N264, N106);
or OR2 (N266, N265, N150);
xor XOR2 (N267, N255, N107);
nor NOR3 (N268, N238, N98, N60);
or OR4 (N269, N263, N26, N59, N259);
buf BUF1 (N270, N269);
nor NOR3 (N271, N268, N220, N216);
buf BUF1 (N272, N266);
nand NAND4 (N273, N271, N27, N43, N152);
or OR2 (N274, N267, N195);
nor NOR2 (N275, N273, N227);
or OR4 (N276, N253, N251, N62, N110);
or OR2 (N277, N270, N119);
and AND3 (N278, N260, N169, N245);
nor NOR3 (N279, N274, N58, N51);
nor NOR3 (N280, N272, N49, N200);
nand NAND2 (N281, N262, N236);
and AND2 (N282, N250, N8);
and AND4 (N283, N279, N143, N212, N234);
or OR2 (N284, N275, N81);
xor XOR2 (N285, N278, N280);
and AND2 (N286, N95, N134);
nand NAND4 (N287, N285, N100, N210, N18);
buf BUF1 (N288, N283);
not NOT1 (N289, N281);
and AND3 (N290, N289, N278, N275);
or OR4 (N291, N287, N248, N156, N264);
not NOT1 (N292, N282);
buf BUF1 (N293, N256);
nand NAND3 (N294, N288, N290, N55);
nand NAND3 (N295, N110, N212, N131);
and AND3 (N296, N284, N50, N276);
nor NOR4 (N297, N296, N141, N80, N50);
xor XOR2 (N298, N154, N108);
nand NAND2 (N299, N257, N59);
buf BUF1 (N300, N286);
or OR3 (N301, N291, N11, N131);
or OR2 (N302, N293, N166);
not NOT1 (N303, N301);
nand NAND3 (N304, N277, N280, N182);
xor XOR2 (N305, N304, N113);
or OR2 (N306, N299, N165);
buf BUF1 (N307, N294);
nor NOR4 (N308, N302, N172, N105, N177);
xor XOR2 (N309, N307, N96);
xor XOR2 (N310, N300, N136);
or OR2 (N311, N292, N52);
xor XOR2 (N312, N306, N119);
nand NAND4 (N313, N308, N100, N79, N286);
not NOT1 (N314, N312);
buf BUF1 (N315, N298);
not NOT1 (N316, N310);
nor NOR4 (N317, N303, N265, N243, N274);
buf BUF1 (N318, N311);
nor NOR4 (N319, N309, N291, N121, N124);
nor NOR4 (N320, N314, N79, N35, N86);
and AND4 (N321, N320, N305, N150, N286);
or OR4 (N322, N139, N83, N316, N247);
xor XOR2 (N323, N161, N158);
not NOT1 (N324, N321);
and AND3 (N325, N323, N176, N305);
nand NAND4 (N326, N325, N204, N305, N248);
and AND2 (N327, N315, N270);
not NOT1 (N328, N327);
not NOT1 (N329, N328);
xor XOR2 (N330, N295, N96);
xor XOR2 (N331, N313, N34);
buf BUF1 (N332, N297);
not NOT1 (N333, N318);
xor XOR2 (N334, N319, N261);
buf BUF1 (N335, N331);
buf BUF1 (N336, N317);
nand NAND2 (N337, N330, N116);
not NOT1 (N338, N336);
buf BUF1 (N339, N324);
nor NOR3 (N340, N329, N196, N337);
buf BUF1 (N341, N202);
not NOT1 (N342, N332);
and AND3 (N343, N339, N256, N39);
xor XOR2 (N344, N334, N70);
not NOT1 (N345, N333);
and AND4 (N346, N326, N271, N286, N201);
or OR4 (N347, N346, N276, N227, N38);
or OR4 (N348, N322, N297, N14, N303);
nor NOR2 (N349, N342, N191);
xor XOR2 (N350, N341, N44);
nor NOR2 (N351, N345, N109);
not NOT1 (N352, N351);
not NOT1 (N353, N352);
xor XOR2 (N354, N349, N313);
nand NAND4 (N355, N348, N236, N20, N43);
and AND4 (N356, N353, N158, N169, N246);
nand NAND4 (N357, N356, N127, N73, N19);
not NOT1 (N358, N344);
not NOT1 (N359, N340);
xor XOR2 (N360, N338, N207);
nand NAND2 (N361, N359, N17);
nor NOR4 (N362, N335, N93, N318, N234);
buf BUF1 (N363, N361);
buf BUF1 (N364, N343);
or OR4 (N365, N357, N148, N19, N111);
or OR3 (N366, N354, N363, N119);
or OR4 (N367, N18, N93, N22, N38);
xor XOR2 (N368, N367, N303);
nor NOR2 (N369, N355, N271);
nand NAND2 (N370, N360, N220);
xor XOR2 (N371, N368, N227);
and AND3 (N372, N358, N64, N187);
and AND3 (N373, N364, N11, N321);
nand NAND2 (N374, N366, N248);
nor NOR4 (N375, N370, N202, N16, N300);
nand NAND2 (N376, N362, N365);
buf BUF1 (N377, N287);
nor NOR4 (N378, N369, N73, N360, N173);
or OR2 (N379, N376, N361);
buf BUF1 (N380, N372);
or OR4 (N381, N350, N171, N324, N2);
nor NOR4 (N382, N373, N364, N46, N111);
and AND3 (N383, N374, N105, N331);
xor XOR2 (N384, N371, N286);
nor NOR3 (N385, N380, N302, N250);
xor XOR2 (N386, N385, N381);
nand NAND3 (N387, N46, N149, N356);
or OR2 (N388, N379, N23);
nor NOR3 (N389, N375, N38, N203);
and AND2 (N390, N383, N228);
buf BUF1 (N391, N384);
or OR3 (N392, N391, N200, N300);
buf BUF1 (N393, N378);
or OR2 (N394, N382, N227);
buf BUF1 (N395, N389);
buf BUF1 (N396, N390);
and AND4 (N397, N347, N71, N335, N262);
nor NOR3 (N398, N396, N375, N298);
not NOT1 (N399, N395);
or OR3 (N400, N377, N146, N320);
xor XOR2 (N401, N393, N229);
not NOT1 (N402, N401);
and AND3 (N403, N400, N16, N151);
nor NOR2 (N404, N388, N61);
or OR2 (N405, N394, N271);
and AND2 (N406, N404, N369);
or OR2 (N407, N398, N235);
and AND3 (N408, N405, N262, N117);
and AND4 (N409, N403, N189, N39, N50);
not NOT1 (N410, N406);
or OR4 (N411, N397, N107, N332, N375);
buf BUF1 (N412, N408);
or OR4 (N413, N409, N66, N38, N254);
or OR3 (N414, N387, N322, N395);
xor XOR2 (N415, N412, N382);
and AND3 (N416, N410, N223, N84);
nand NAND2 (N417, N407, N275);
or OR2 (N418, N386, N264);
and AND4 (N419, N418, N417, N352, N418);
nand NAND3 (N420, N375, N285, N80);
xor XOR2 (N421, N402, N230);
buf BUF1 (N422, N415);
not NOT1 (N423, N420);
buf BUF1 (N424, N413);
not NOT1 (N425, N422);
buf BUF1 (N426, N419);
xor XOR2 (N427, N392, N198);
nor NOR2 (N428, N399, N262);
not NOT1 (N429, N427);
and AND3 (N430, N429, N37, N357);
buf BUF1 (N431, N411);
nand NAND2 (N432, N430, N22);
not NOT1 (N433, N426);
xor XOR2 (N434, N431, N209);
nand NAND2 (N435, N434, N153);
and AND3 (N436, N421, N199, N238);
and AND4 (N437, N428, N374, N275, N187);
xor XOR2 (N438, N416, N300);
and AND4 (N439, N438, N237, N24, N159);
nand NAND4 (N440, N435, N249, N272, N18);
nand NAND2 (N441, N436, N249);
or OR2 (N442, N423, N202);
or OR3 (N443, N442, N409, N199);
buf BUF1 (N444, N424);
and AND4 (N445, N432, N412, N294, N132);
buf BUF1 (N446, N440);
or OR3 (N447, N446, N164, N441);
buf BUF1 (N448, N123);
nor NOR3 (N449, N414, N48, N17);
nand NAND4 (N450, N425, N48, N162, N356);
or OR2 (N451, N450, N122);
nand NAND2 (N452, N448, N342);
nor NOR2 (N453, N445, N241);
nor NOR2 (N454, N447, N339);
and AND3 (N455, N451, N389, N405);
not NOT1 (N456, N452);
nand NAND2 (N457, N444, N190);
buf BUF1 (N458, N433);
not NOT1 (N459, N437);
or OR4 (N460, N457, N181, N443, N165);
xor XOR2 (N461, N335, N387);
or OR2 (N462, N458, N306);
not NOT1 (N463, N462);
xor XOR2 (N464, N461, N314);
nor NOR3 (N465, N449, N402, N384);
not NOT1 (N466, N456);
or OR3 (N467, N466, N149, N33);
nand NAND4 (N468, N454, N349, N245, N272);
not NOT1 (N469, N460);
and AND3 (N470, N459, N172, N240);
xor XOR2 (N471, N453, N34);
nand NAND3 (N472, N465, N345, N26);
nor NOR4 (N473, N455, N384, N441, N289);
nand NAND3 (N474, N467, N295, N90);
and AND3 (N475, N474, N402, N351);
nand NAND4 (N476, N439, N180, N409, N93);
not NOT1 (N477, N468);
and AND4 (N478, N469, N334, N324, N275);
nand NAND4 (N479, N477, N21, N101, N274);
and AND3 (N480, N476, N150, N169);
and AND3 (N481, N470, N421, N320);
nor NOR2 (N482, N472, N4);
nor NOR4 (N483, N463, N408, N375, N333);
buf BUF1 (N484, N471);
buf BUF1 (N485, N473);
buf BUF1 (N486, N483);
not NOT1 (N487, N481);
buf BUF1 (N488, N478);
and AND4 (N489, N479, N58, N279, N302);
nor NOR4 (N490, N485, N76, N448, N283);
buf BUF1 (N491, N475);
not NOT1 (N492, N482);
buf BUF1 (N493, N487);
and AND2 (N494, N480, N226);
not NOT1 (N495, N491);
and AND3 (N496, N484, N387, N215);
or OR4 (N497, N490, N190, N27, N492);
nor NOR4 (N498, N394, N341, N223, N57);
nand NAND2 (N499, N498, N362);
and AND2 (N500, N464, N308);
nand NAND3 (N501, N500, N160, N347);
not NOT1 (N502, N493);
buf BUF1 (N503, N501);
nand NAND3 (N504, N503, N389, N9);
xor XOR2 (N505, N504, N10);
not NOT1 (N506, N488);
or OR2 (N507, N499, N492);
buf BUF1 (N508, N507);
and AND4 (N509, N495, N150, N468, N197);
xor XOR2 (N510, N505, N318);
buf BUF1 (N511, N497);
not NOT1 (N512, N494);
and AND3 (N513, N511, N138, N441);
and AND2 (N514, N513, N98);
xor XOR2 (N515, N506, N255);
and AND3 (N516, N515, N213, N233);
or OR4 (N517, N489, N390, N229, N398);
not NOT1 (N518, N512);
and AND3 (N519, N516, N216, N354);
buf BUF1 (N520, N518);
buf BUF1 (N521, N509);
nand NAND4 (N522, N486, N213, N306, N296);
buf BUF1 (N523, N520);
and AND3 (N524, N502, N206, N437);
not NOT1 (N525, N519);
or OR4 (N526, N522, N233, N76, N86);
buf BUF1 (N527, N523);
xor XOR2 (N528, N521, N400);
not NOT1 (N529, N508);
buf BUF1 (N530, N514);
not NOT1 (N531, N528);
nor NOR4 (N532, N524, N366, N501, N490);
nand NAND3 (N533, N529, N24, N384);
or OR2 (N534, N532, N162);
not NOT1 (N535, N531);
nand NAND3 (N536, N517, N155, N246);
not NOT1 (N537, N526);
nor NOR2 (N538, N535, N173);
nand NAND3 (N539, N510, N328, N417);
or OR2 (N540, N534, N501);
and AND2 (N541, N536, N274);
or OR2 (N542, N533, N128);
xor XOR2 (N543, N496, N540);
buf BUF1 (N544, N279);
and AND4 (N545, N542, N180, N247, N179);
and AND4 (N546, N543, N31, N99, N153);
not NOT1 (N547, N539);
buf BUF1 (N548, N547);
nor NOR4 (N549, N544, N367, N259, N162);
not NOT1 (N550, N549);
nor NOR2 (N551, N546, N60);
and AND3 (N552, N525, N172, N208);
and AND4 (N553, N538, N474, N180, N258);
nor NOR3 (N554, N545, N294, N319);
or OR4 (N555, N553, N139, N381, N156);
and AND2 (N556, N541, N167);
nor NOR3 (N557, N551, N277, N4);
buf BUF1 (N558, N555);
not NOT1 (N559, N550);
or OR2 (N560, N554, N309);
xor XOR2 (N561, N560, N82);
xor XOR2 (N562, N561, N131);
nand NAND2 (N563, N556, N408);
xor XOR2 (N564, N530, N182);
nor NOR4 (N565, N552, N445, N91, N542);
buf BUF1 (N566, N558);
nand NAND2 (N567, N563, N561);
and AND4 (N568, N557, N560, N174, N259);
xor XOR2 (N569, N559, N286);
nand NAND2 (N570, N565, N490);
not NOT1 (N571, N562);
buf BUF1 (N572, N564);
xor XOR2 (N573, N537, N130);
or OR3 (N574, N572, N529, N495);
not NOT1 (N575, N568);
or OR3 (N576, N570, N575, N211);
xor XOR2 (N577, N405, N58);
nor NOR3 (N578, N571, N576, N152);
nor NOR4 (N579, N290, N203, N125, N104);
nand NAND4 (N580, N579, N570, N50, N242);
and AND4 (N581, N567, N60, N515, N539);
and AND3 (N582, N566, N73, N107);
nand NAND2 (N583, N573, N327);
or OR3 (N584, N574, N232, N407);
buf BUF1 (N585, N580);
buf BUF1 (N586, N584);
not NOT1 (N587, N577);
nor NOR4 (N588, N585, N433, N180, N544);
nand NAND3 (N589, N588, N417, N220);
nor NOR4 (N590, N548, N358, N178, N563);
and AND3 (N591, N589, N549, N408);
nand NAND4 (N592, N581, N406, N306, N354);
or OR4 (N593, N582, N48, N302, N103);
nor NOR3 (N594, N587, N556, N429);
or OR4 (N595, N527, N318, N292, N363);
and AND2 (N596, N583, N237);
xor XOR2 (N597, N586, N168);
and AND2 (N598, N592, N289);
or OR3 (N599, N595, N291, N340);
nand NAND2 (N600, N598, N348);
or OR4 (N601, N590, N282, N484, N392);
or OR3 (N602, N599, N123, N277);
not NOT1 (N603, N594);
xor XOR2 (N604, N597, N505);
not NOT1 (N605, N601);
and AND2 (N606, N569, N565);
xor XOR2 (N607, N604, N521);
xor XOR2 (N608, N591, N412);
buf BUF1 (N609, N596);
nor NOR4 (N610, N603, N262, N345, N139);
not NOT1 (N611, N605);
and AND2 (N612, N606, N220);
and AND4 (N613, N610, N508, N97, N212);
and AND3 (N614, N609, N88, N481);
nand NAND2 (N615, N593, N357);
nor NOR2 (N616, N600, N230);
nor NOR3 (N617, N578, N5, N313);
nor NOR4 (N618, N607, N448, N377, N305);
xor XOR2 (N619, N613, N28);
nand NAND4 (N620, N616, N254, N263, N512);
nand NAND2 (N621, N608, N156);
nor NOR2 (N622, N618, N301);
nand NAND3 (N623, N611, N264, N127);
not NOT1 (N624, N619);
not NOT1 (N625, N614);
not NOT1 (N626, N625);
and AND4 (N627, N623, N61, N183, N175);
not NOT1 (N628, N612);
nor NOR4 (N629, N621, N468, N234, N132);
nor NOR4 (N630, N628, N249, N66, N360);
xor XOR2 (N631, N626, N13);
nor NOR3 (N632, N620, N159, N63);
and AND3 (N633, N630, N534, N605);
nand NAND3 (N634, N602, N80, N143);
buf BUF1 (N635, N622);
and AND2 (N636, N615, N470);
buf BUF1 (N637, N627);
nand NAND4 (N638, N624, N585, N464, N261);
xor XOR2 (N639, N633, N463);
xor XOR2 (N640, N617, N81);
xor XOR2 (N641, N632, N566);
and AND4 (N642, N629, N636, N11, N390);
xor XOR2 (N643, N7, N469);
not NOT1 (N644, N641);
xor XOR2 (N645, N638, N352);
and AND4 (N646, N645, N188, N452, N76);
and AND2 (N647, N642, N490);
buf BUF1 (N648, N644);
nand NAND2 (N649, N646, N536);
not NOT1 (N650, N631);
and AND4 (N651, N649, N119, N298, N432);
not NOT1 (N652, N634);
not NOT1 (N653, N640);
nor NOR4 (N654, N647, N386, N391, N614);
or OR3 (N655, N637, N252, N259);
nand NAND2 (N656, N652, N51);
or OR2 (N657, N654, N328);
nor NOR3 (N658, N639, N335, N615);
xor XOR2 (N659, N635, N539);
nand NAND3 (N660, N659, N88, N196);
buf BUF1 (N661, N651);
buf BUF1 (N662, N656);
nor NOR3 (N663, N658, N431, N81);
not NOT1 (N664, N662);
not NOT1 (N665, N648);
not NOT1 (N666, N660);
or OR2 (N667, N657, N2);
nor NOR4 (N668, N655, N289, N610, N316);
not NOT1 (N669, N664);
nand NAND4 (N670, N667, N69, N154, N261);
nand NAND2 (N671, N668, N1);
not NOT1 (N672, N650);
nor NOR2 (N673, N663, N4);
nand NAND3 (N674, N666, N77, N415);
xor XOR2 (N675, N670, N648);
buf BUF1 (N676, N675);
buf BUF1 (N677, N672);
xor XOR2 (N678, N653, N538);
nand NAND3 (N679, N673, N102, N102);
nor NOR2 (N680, N669, N223);
not NOT1 (N681, N680);
xor XOR2 (N682, N677, N74);
and AND3 (N683, N681, N518, N616);
nand NAND2 (N684, N676, N491);
xor XOR2 (N685, N678, N192);
nor NOR3 (N686, N685, N386, N35);
nor NOR2 (N687, N671, N67);
not NOT1 (N688, N679);
not NOT1 (N689, N684);
nor NOR2 (N690, N689, N286);
xor XOR2 (N691, N661, N403);
nand NAND4 (N692, N688, N328, N688, N318);
not NOT1 (N693, N690);
nand NAND2 (N694, N691, N680);
and AND4 (N695, N674, N432, N107, N690);
or OR4 (N696, N693, N46, N540, N526);
buf BUF1 (N697, N683);
nor NOR4 (N698, N665, N200, N127, N577);
buf BUF1 (N699, N697);
xor XOR2 (N700, N686, N110);
nor NOR4 (N701, N700, N592, N631, N271);
nand NAND3 (N702, N696, N520, N552);
nor NOR2 (N703, N687, N418);
buf BUF1 (N704, N682);
or OR3 (N705, N701, N7, N56);
buf BUF1 (N706, N695);
nor NOR2 (N707, N702, N701);
nor NOR2 (N708, N705, N546);
buf BUF1 (N709, N704);
not NOT1 (N710, N706);
nand NAND3 (N711, N699, N353, N656);
not NOT1 (N712, N703);
not NOT1 (N713, N643);
or OR2 (N714, N692, N36);
not NOT1 (N715, N714);
and AND3 (N716, N711, N308, N332);
and AND2 (N717, N713, N104);
buf BUF1 (N718, N708);
and AND4 (N719, N710, N512, N294, N429);
xor XOR2 (N720, N719, N29);
not NOT1 (N721, N698);
xor XOR2 (N722, N715, N230);
or OR4 (N723, N716, N524, N609, N306);
not NOT1 (N724, N694);
or OR2 (N725, N718, N339);
nor NOR2 (N726, N722, N511);
or OR2 (N727, N707, N503);
not NOT1 (N728, N720);
or OR2 (N729, N724, N293);
and AND2 (N730, N729, N305);
and AND4 (N731, N723, N128, N728, N713);
buf BUF1 (N732, N289);
not NOT1 (N733, N712);
buf BUF1 (N734, N725);
buf BUF1 (N735, N726);
buf BUF1 (N736, N732);
nand NAND3 (N737, N709, N538, N636);
xor XOR2 (N738, N721, N577);
nand NAND2 (N739, N717, N469);
buf BUF1 (N740, N731);
nand NAND4 (N741, N736, N550, N520, N708);
xor XOR2 (N742, N737, N70);
xor XOR2 (N743, N727, N626);
or OR4 (N744, N740, N359, N18, N459);
or OR4 (N745, N739, N468, N62, N329);
nor NOR4 (N746, N738, N198, N546, N510);
not NOT1 (N747, N745);
and AND4 (N748, N735, N143, N584, N317);
xor XOR2 (N749, N734, N95);
xor XOR2 (N750, N747, N461);
buf BUF1 (N751, N733);
and AND2 (N752, N742, N552);
nor NOR3 (N753, N746, N71, N146);
not NOT1 (N754, N730);
and AND3 (N755, N743, N271, N660);
nand NAND3 (N756, N748, N731, N437);
not NOT1 (N757, N756);
nand NAND3 (N758, N750, N377, N509);
xor XOR2 (N759, N753, N259);
nand NAND3 (N760, N752, N49, N473);
xor XOR2 (N761, N759, N178);
buf BUF1 (N762, N760);
xor XOR2 (N763, N761, N425);
and AND4 (N764, N757, N324, N41, N562);
and AND3 (N765, N755, N176, N277);
and AND3 (N766, N758, N167, N177);
and AND3 (N767, N762, N241, N221);
nor NOR4 (N768, N765, N67, N184, N558);
not NOT1 (N769, N763);
nand NAND4 (N770, N766, N189, N668, N380);
xor XOR2 (N771, N769, N247);
nand NAND2 (N772, N749, N414);
not NOT1 (N773, N744);
nor NOR2 (N774, N772, N109);
xor XOR2 (N775, N768, N108);
xor XOR2 (N776, N771, N539);
nand NAND4 (N777, N754, N638, N443, N557);
not NOT1 (N778, N764);
xor XOR2 (N779, N778, N640);
or OR2 (N780, N777, N282);
not NOT1 (N781, N773);
xor XOR2 (N782, N779, N609);
or OR3 (N783, N770, N460, N515);
nor NOR4 (N784, N741, N212, N25, N534);
xor XOR2 (N785, N783, N558);
xor XOR2 (N786, N785, N434);
or OR3 (N787, N784, N280, N773);
buf BUF1 (N788, N767);
not NOT1 (N789, N776);
or OR4 (N790, N786, N25, N779, N553);
not NOT1 (N791, N774);
nor NOR2 (N792, N775, N744);
buf BUF1 (N793, N787);
nand NAND4 (N794, N791, N471, N462, N374);
not NOT1 (N795, N792);
buf BUF1 (N796, N751);
xor XOR2 (N797, N794, N662);
nand NAND4 (N798, N795, N4, N248, N12);
nand NAND4 (N799, N780, N399, N398, N28);
or OR2 (N800, N788, N358);
and AND2 (N801, N793, N117);
xor XOR2 (N802, N782, N2);
xor XOR2 (N803, N798, N499);
not NOT1 (N804, N803);
or OR2 (N805, N802, N708);
or OR4 (N806, N805, N402, N46, N193);
buf BUF1 (N807, N796);
buf BUF1 (N808, N781);
nor NOR2 (N809, N801, N206);
xor XOR2 (N810, N789, N382);
and AND4 (N811, N799, N262, N135, N577);
or OR4 (N812, N809, N40, N458, N154);
buf BUF1 (N813, N797);
xor XOR2 (N814, N812, N156);
nor NOR4 (N815, N813, N77, N769, N601);
nor NOR4 (N816, N790, N36, N171, N282);
xor XOR2 (N817, N810, N429);
and AND3 (N818, N811, N453, N254);
not NOT1 (N819, N814);
nor NOR4 (N820, N816, N215, N573, N687);
not NOT1 (N821, N820);
buf BUF1 (N822, N804);
buf BUF1 (N823, N817);
or OR2 (N824, N823, N453);
nor NOR2 (N825, N824, N444);
not NOT1 (N826, N807);
xor XOR2 (N827, N806, N274);
not NOT1 (N828, N827);
buf BUF1 (N829, N808);
not NOT1 (N830, N815);
or OR3 (N831, N818, N212, N722);
buf BUF1 (N832, N825);
or OR2 (N833, N829, N301);
or OR2 (N834, N828, N765);
or OR3 (N835, N819, N583, N34);
nor NOR2 (N836, N822, N407);
or OR3 (N837, N832, N612, N37);
xor XOR2 (N838, N831, N313);
or OR4 (N839, N800, N826, N800, N798);
not NOT1 (N840, N564);
not NOT1 (N841, N840);
nor NOR4 (N842, N835, N367, N774, N97);
and AND3 (N843, N838, N360, N325);
nor NOR3 (N844, N836, N46, N206);
xor XOR2 (N845, N830, N497);
xor XOR2 (N846, N821, N145);
and AND2 (N847, N833, N527);
nand NAND2 (N848, N846, N174);
nor NOR3 (N849, N844, N844, N119);
or OR2 (N850, N834, N831);
xor XOR2 (N851, N839, N505);
and AND3 (N852, N845, N545, N255);
buf BUF1 (N853, N848);
not NOT1 (N854, N853);
xor XOR2 (N855, N850, N10);
not NOT1 (N856, N837);
xor XOR2 (N857, N849, N558);
nor NOR3 (N858, N856, N709, N274);
or OR4 (N859, N858, N294, N792, N423);
not NOT1 (N860, N857);
and AND3 (N861, N847, N728, N285);
nand NAND3 (N862, N855, N182, N287);
not NOT1 (N863, N852);
and AND2 (N864, N862, N380);
or OR2 (N865, N842, N41);
or OR3 (N866, N854, N764, N463);
nand NAND3 (N867, N843, N725, N141);
buf BUF1 (N868, N859);
and AND2 (N869, N851, N56);
nor NOR2 (N870, N869, N287);
and AND3 (N871, N870, N669, N620);
or OR2 (N872, N863, N78);
xor XOR2 (N873, N861, N479);
not NOT1 (N874, N865);
not NOT1 (N875, N874);
nand NAND4 (N876, N875, N646, N590, N400);
xor XOR2 (N877, N872, N385);
or OR3 (N878, N841, N793, N783);
or OR3 (N879, N868, N120, N26);
buf BUF1 (N880, N877);
nand NAND4 (N881, N866, N724, N77, N441);
nand NAND4 (N882, N876, N835, N486, N607);
and AND4 (N883, N882, N546, N116, N310);
nand NAND3 (N884, N867, N604, N749);
not NOT1 (N885, N880);
not NOT1 (N886, N884);
or OR3 (N887, N883, N546, N288);
and AND2 (N888, N879, N256);
nand NAND3 (N889, N886, N670, N84);
and AND3 (N890, N871, N510, N472);
not NOT1 (N891, N864);
nand NAND3 (N892, N885, N94, N838);
buf BUF1 (N893, N888);
or OR3 (N894, N873, N856, N716);
or OR2 (N895, N889, N413);
not NOT1 (N896, N890);
nor NOR4 (N897, N881, N762, N609, N251);
not NOT1 (N898, N895);
and AND4 (N899, N860, N41, N301, N724);
or OR2 (N900, N893, N514);
nor NOR3 (N901, N897, N160, N425);
buf BUF1 (N902, N892);
nand NAND2 (N903, N887, N86);
nand NAND4 (N904, N903, N185, N682, N805);
nand NAND2 (N905, N904, N474);
and AND3 (N906, N901, N904, N300);
nand NAND2 (N907, N905, N572);
and AND3 (N908, N907, N76, N708);
not NOT1 (N909, N906);
not NOT1 (N910, N898);
or OR2 (N911, N899, N901);
and AND4 (N912, N894, N582, N7, N773);
nor NOR2 (N913, N908, N515);
or OR4 (N914, N913, N552, N57, N92);
and AND3 (N915, N896, N242, N304);
buf BUF1 (N916, N878);
nand NAND2 (N917, N912, N559);
nand NAND4 (N918, N910, N730, N643, N703);
and AND4 (N919, N909, N606, N103, N176);
not NOT1 (N920, N916);
or OR2 (N921, N911, N459);
nand NAND2 (N922, N915, N547);
and AND3 (N923, N914, N3, N114);
xor XOR2 (N924, N891, N510);
buf BUF1 (N925, N922);
not NOT1 (N926, N919);
and AND2 (N927, N926, N612);
nand NAND4 (N928, N918, N397, N208, N351);
nor NOR2 (N929, N925, N612);
and AND4 (N930, N924, N386, N607, N138);
xor XOR2 (N931, N902, N844);
and AND4 (N932, N928, N423, N161, N455);
buf BUF1 (N933, N930);
buf BUF1 (N934, N932);
nor NOR2 (N935, N931, N31);
and AND3 (N936, N917, N615, N158);
not NOT1 (N937, N921);
nand NAND4 (N938, N923, N180, N927, N378);
buf BUF1 (N939, N564);
and AND4 (N940, N939, N444, N912, N73);
nor NOR2 (N941, N935, N80);
not NOT1 (N942, N936);
and AND4 (N943, N929, N405, N709, N183);
buf BUF1 (N944, N937);
not NOT1 (N945, N933);
xor XOR2 (N946, N900, N759);
or OR2 (N947, N940, N732);
or OR4 (N948, N938, N257, N362, N60);
not NOT1 (N949, N942);
and AND2 (N950, N945, N408);
and AND2 (N951, N941, N210);
and AND4 (N952, N943, N147, N217, N104);
nand NAND3 (N953, N947, N856, N172);
not NOT1 (N954, N949);
not NOT1 (N955, N953);
or OR2 (N956, N946, N375);
nand NAND4 (N957, N956, N253, N469, N445);
or OR3 (N958, N957, N249, N781);
nand NAND2 (N959, N948, N750);
nor NOR2 (N960, N920, N34);
not NOT1 (N961, N954);
not NOT1 (N962, N934);
nor NOR2 (N963, N962, N377);
buf BUF1 (N964, N950);
or OR3 (N965, N955, N642, N527);
nand NAND3 (N966, N964, N308, N201);
or OR3 (N967, N958, N554, N248);
or OR2 (N968, N944, N863);
nor NOR2 (N969, N951, N16);
nand NAND4 (N970, N963, N198, N657, N654);
nor NOR4 (N971, N966, N438, N199, N232);
nand NAND4 (N972, N952, N213, N514, N539);
nand NAND2 (N973, N960, N612);
xor XOR2 (N974, N972, N13);
not NOT1 (N975, N971);
buf BUF1 (N976, N959);
and AND2 (N977, N967, N27);
and AND3 (N978, N974, N471, N312);
buf BUF1 (N979, N977);
buf BUF1 (N980, N961);
xor XOR2 (N981, N979, N535);
not NOT1 (N982, N973);
and AND3 (N983, N968, N861, N133);
nand NAND3 (N984, N970, N886, N837);
buf BUF1 (N985, N976);
and AND4 (N986, N982, N303, N733, N194);
xor XOR2 (N987, N981, N468);
or OR3 (N988, N983, N904, N705);
and AND3 (N989, N988, N133, N18);
or OR4 (N990, N975, N21, N837, N81);
buf BUF1 (N991, N987);
nor NOR3 (N992, N980, N136, N86);
or OR2 (N993, N984, N542);
nand NAND2 (N994, N969, N42);
xor XOR2 (N995, N990, N416);
nand NAND3 (N996, N989, N701, N478);
xor XOR2 (N997, N965, N769);
nor NOR3 (N998, N978, N801, N439);
not NOT1 (N999, N994);
buf BUF1 (N1000, N992);
buf BUF1 (N1001, N1000);
or OR4 (N1002, N997, N205, N988, N699);
not NOT1 (N1003, N985);
buf BUF1 (N1004, N1002);
not NOT1 (N1005, N995);
buf BUF1 (N1006, N999);
buf BUF1 (N1007, N1001);
nand NAND2 (N1008, N1005, N59);
nand NAND4 (N1009, N1008, N227, N106, N603);
nor NOR4 (N1010, N1004, N615, N906, N166);
xor XOR2 (N1011, N1007, N474);
not NOT1 (N1012, N1010);
nand NAND3 (N1013, N1006, N778, N80);
and AND3 (N1014, N996, N401, N532);
nand NAND3 (N1015, N1012, N155, N268);
and AND4 (N1016, N993, N138, N117, N179);
or OR4 (N1017, N998, N576, N324, N940);
not NOT1 (N1018, N1017);
endmodule