// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20;

output N3517,N3491,N3512,N3515,N3513,N3516,N3519,N3494,N3514,N3520;

or OR2 (N21, N11, N13);
nor NOR2 (N22, N5, N17);
nand NAND3 (N23, N9, N3, N19);
xor XOR2 (N24, N6, N14);
not NOT1 (N25, N23);
not NOT1 (N26, N5);
nor NOR3 (N27, N15, N21, N13);
and AND2 (N28, N26, N2);
xor XOR2 (N29, N4, N14);
xor XOR2 (N30, N7, N29);
nor NOR3 (N31, N16, N18, N26);
nand NAND3 (N32, N22, N22, N11);
nand NAND3 (N33, N9, N18, N9);
buf BUF1 (N34, N13);
nand NAND3 (N35, N23, N2, N10);
and AND2 (N36, N34, N17);
or OR3 (N37, N35, N17, N9);
xor XOR2 (N38, N32, N10);
xor XOR2 (N39, N31, N15);
nand NAND4 (N40, N33, N22, N36, N17);
or OR2 (N41, N39, N40);
nor NOR3 (N42, N20, N34, N33);
and AND4 (N43, N18, N35, N31, N28);
buf BUF1 (N44, N34);
nor NOR3 (N45, N38, N22, N22);
nor NOR3 (N46, N24, N40, N45);
buf BUF1 (N47, N39);
nor NOR4 (N48, N41, N37, N23, N37);
and AND4 (N49, N1, N5, N15, N27);
nor NOR3 (N50, N49, N25, N28);
xor XOR2 (N51, N13, N44);
xor XOR2 (N52, N15, N19);
buf BUF1 (N53, N11);
nand NAND3 (N54, N43, N14, N35);
nand NAND2 (N55, N42, N46);
or OR4 (N56, N48, N39, N53, N30);
buf BUF1 (N57, N5);
and AND4 (N58, N33, N33, N3, N13);
buf BUF1 (N59, N53);
xor XOR2 (N60, N51, N12);
nand NAND3 (N61, N58, N57, N26);
or OR2 (N62, N54, N57);
or OR3 (N63, N56, N13, N50);
xor XOR2 (N64, N24, N31);
nand NAND4 (N65, N10, N53, N50, N58);
nor NOR2 (N66, N47, N30);
nand NAND3 (N67, N65, N48, N1);
nand NAND3 (N68, N67, N49, N38);
xor XOR2 (N69, N60, N51);
not NOT1 (N70, N62);
not NOT1 (N71, N63);
nand NAND4 (N72, N71, N31, N40, N13);
buf BUF1 (N73, N55);
not NOT1 (N74, N73);
xor XOR2 (N75, N52, N53);
xor XOR2 (N76, N69, N27);
or OR3 (N77, N72, N74, N45);
not NOT1 (N78, N75);
xor XOR2 (N79, N42, N3);
nor NOR4 (N80, N76, N35, N10, N73);
not NOT1 (N81, N61);
nand NAND2 (N82, N64, N49);
nand NAND4 (N83, N82, N50, N32, N6);
buf BUF1 (N84, N78);
buf BUF1 (N85, N77);
not NOT1 (N86, N81);
nand NAND2 (N87, N79, N61);
or OR3 (N88, N59, N37, N68);
or OR2 (N89, N15, N44);
nor NOR3 (N90, N70, N13, N46);
nor NOR3 (N91, N87, N18, N11);
and AND2 (N92, N91, N13);
or OR3 (N93, N84, N74, N40);
not NOT1 (N94, N90);
not NOT1 (N95, N86);
nand NAND3 (N96, N93, N84, N87);
not NOT1 (N97, N85);
not NOT1 (N98, N97);
or OR2 (N99, N94, N84);
buf BUF1 (N100, N98);
nand NAND4 (N101, N66, N21, N25, N37);
not NOT1 (N102, N99);
or OR3 (N103, N100, N54, N80);
nand NAND4 (N104, N67, N97, N15, N6);
not NOT1 (N105, N103);
buf BUF1 (N106, N102);
nor NOR2 (N107, N106, N40);
nand NAND4 (N108, N101, N12, N30, N99);
xor XOR2 (N109, N104, N106);
xor XOR2 (N110, N83, N38);
nand NAND2 (N111, N95, N23);
nand NAND4 (N112, N108, N23, N65, N74);
buf BUF1 (N113, N89);
nand NAND4 (N114, N92, N58, N83, N14);
nand NAND3 (N115, N105, N31, N44);
and AND2 (N116, N88, N68);
xor XOR2 (N117, N109, N20);
and AND3 (N118, N115, N82, N28);
or OR2 (N119, N114, N32);
not NOT1 (N120, N107);
buf BUF1 (N121, N110);
xor XOR2 (N122, N121, N72);
buf BUF1 (N123, N120);
nand NAND4 (N124, N113, N84, N96, N48);
buf BUF1 (N125, N18);
or OR3 (N126, N119, N66, N18);
nor NOR2 (N127, N122, N93);
xor XOR2 (N128, N124, N36);
or OR3 (N129, N127, N109, N100);
nand NAND2 (N130, N116, N104);
not NOT1 (N131, N111);
nand NAND4 (N132, N112, N114, N32, N23);
buf BUF1 (N133, N128);
or OR4 (N134, N131, N112, N125, N124);
xor XOR2 (N135, N45, N64);
nor NOR3 (N136, N130, N125, N32);
and AND4 (N137, N133, N97, N67, N122);
nor NOR3 (N138, N129, N15, N52);
and AND2 (N139, N126, N50);
nand NAND2 (N140, N117, N109);
not NOT1 (N141, N136);
and AND4 (N142, N139, N22, N135, N78);
nand NAND3 (N143, N81, N72, N126);
and AND3 (N144, N134, N115, N105);
xor XOR2 (N145, N140, N93);
nand NAND2 (N146, N118, N51);
not NOT1 (N147, N144);
or OR2 (N148, N146, N23);
xor XOR2 (N149, N123, N144);
xor XOR2 (N150, N137, N117);
not NOT1 (N151, N147);
nor NOR2 (N152, N150, N39);
buf BUF1 (N153, N143);
buf BUF1 (N154, N141);
xor XOR2 (N155, N154, N33);
nor NOR4 (N156, N152, N37, N85, N7);
or OR4 (N157, N138, N33, N116, N132);
buf BUF1 (N158, N127);
buf BUF1 (N159, N145);
nor NOR3 (N160, N142, N147, N108);
buf BUF1 (N161, N155);
or OR2 (N162, N148, N50);
or OR3 (N163, N160, N72, N97);
nand NAND3 (N164, N149, N6, N154);
xor XOR2 (N165, N163, N12);
buf BUF1 (N166, N161);
and AND4 (N167, N162, N144, N116, N133);
and AND3 (N168, N158, N3, N32);
and AND2 (N169, N151, N11);
buf BUF1 (N170, N167);
nand NAND4 (N171, N170, N4, N6, N51);
xor XOR2 (N172, N171, N132);
nor NOR2 (N173, N168, N48);
buf BUF1 (N174, N164);
not NOT1 (N175, N159);
xor XOR2 (N176, N174, N137);
or OR2 (N177, N175, N82);
or OR4 (N178, N172, N48, N88, N7);
xor XOR2 (N179, N165, N7);
nor NOR2 (N180, N176, N177);
xor XOR2 (N181, N115, N87);
nor NOR2 (N182, N178, N21);
and AND3 (N183, N180, N19, N104);
not NOT1 (N184, N181);
and AND2 (N185, N183, N173);
buf BUF1 (N186, N176);
buf BUF1 (N187, N186);
and AND2 (N188, N184, N14);
nor NOR3 (N189, N166, N19, N188);
nand NAND4 (N190, N57, N135, N85, N108);
nand NAND2 (N191, N185, N187);
nor NOR2 (N192, N20, N164);
and AND3 (N193, N169, N131, N51);
or OR4 (N194, N192, N24, N3, N3);
and AND3 (N195, N156, N191, N52);
xor XOR2 (N196, N74, N111);
or OR2 (N197, N190, N191);
not NOT1 (N198, N157);
or OR4 (N199, N197, N60, N189, N171);
nand NAND2 (N200, N182, N144);
and AND3 (N201, N38, N112, N157);
not NOT1 (N202, N193);
nand NAND2 (N203, N153, N113);
and AND4 (N204, N200, N120, N65, N83);
nand NAND3 (N205, N199, N51, N122);
or OR3 (N206, N201, N64, N16);
or OR4 (N207, N205, N197, N124, N134);
or OR3 (N208, N179, N90, N77);
or OR4 (N209, N208, N128, N182, N146);
and AND4 (N210, N203, N8, N47, N172);
xor XOR2 (N211, N196, N115);
and AND4 (N212, N206, N192, N144, N97);
nor NOR4 (N213, N211, N110, N26, N70);
not NOT1 (N214, N204);
buf BUF1 (N215, N209);
buf BUF1 (N216, N214);
or OR2 (N217, N212, N59);
nor NOR4 (N218, N198, N33, N124, N87);
xor XOR2 (N219, N210, N39);
and AND2 (N220, N219, N63);
buf BUF1 (N221, N215);
and AND4 (N222, N202, N23, N196, N136);
nand NAND2 (N223, N218, N179);
nor NOR2 (N224, N217, N203);
nand NAND2 (N225, N195, N34);
nor NOR4 (N226, N224, N69, N6, N39);
xor XOR2 (N227, N225, N65);
not NOT1 (N228, N221);
xor XOR2 (N229, N223, N124);
and AND3 (N230, N213, N189, N190);
buf BUF1 (N231, N230);
nor NOR2 (N232, N228, N218);
xor XOR2 (N233, N226, N85);
nand NAND3 (N234, N233, N77, N36);
not NOT1 (N235, N234);
xor XOR2 (N236, N229, N97);
and AND3 (N237, N216, N88, N228);
or OR2 (N238, N237, N126);
nor NOR3 (N239, N238, N224, N181);
or OR3 (N240, N227, N219, N139);
xor XOR2 (N241, N220, N144);
and AND2 (N242, N222, N97);
buf BUF1 (N243, N194);
xor XOR2 (N244, N243, N105);
or OR4 (N245, N232, N80, N85, N233);
not NOT1 (N246, N241);
buf BUF1 (N247, N245);
nor NOR3 (N248, N242, N51, N244);
and AND2 (N249, N146, N246);
nor NOR3 (N250, N75, N89, N247);
buf BUF1 (N251, N100);
nand NAND2 (N252, N251, N112);
buf BUF1 (N253, N240);
xor XOR2 (N254, N239, N186);
buf BUF1 (N255, N248);
or OR2 (N256, N250, N197);
not NOT1 (N257, N236);
not NOT1 (N258, N207);
not NOT1 (N259, N258);
nor NOR2 (N260, N249, N238);
buf BUF1 (N261, N259);
xor XOR2 (N262, N235, N147);
or OR4 (N263, N253, N245, N245, N54);
nand NAND4 (N264, N257, N176, N75, N248);
xor XOR2 (N265, N252, N247);
buf BUF1 (N266, N265);
buf BUF1 (N267, N260);
and AND2 (N268, N266, N230);
or OR2 (N269, N263, N126);
and AND2 (N270, N268, N241);
and AND3 (N271, N256, N46, N60);
and AND2 (N272, N269, N188);
nand NAND3 (N273, N272, N67, N88);
nor NOR2 (N274, N273, N116);
xor XOR2 (N275, N254, N144);
buf BUF1 (N276, N262);
buf BUF1 (N277, N275);
not NOT1 (N278, N276);
not NOT1 (N279, N267);
not NOT1 (N280, N261);
or OR3 (N281, N279, N251, N208);
and AND2 (N282, N255, N67);
or OR4 (N283, N277, N62, N12, N193);
not NOT1 (N284, N274);
nand NAND3 (N285, N280, N194, N7);
and AND3 (N286, N231, N132, N133);
and AND3 (N287, N281, N142, N124);
nand NAND2 (N288, N271, N251);
buf BUF1 (N289, N286);
nor NOR4 (N290, N278, N268, N216, N37);
xor XOR2 (N291, N290, N19);
xor XOR2 (N292, N283, N261);
not NOT1 (N293, N284);
buf BUF1 (N294, N292);
buf BUF1 (N295, N282);
nor NOR2 (N296, N288, N66);
nor NOR3 (N297, N285, N102, N57);
or OR3 (N298, N270, N132, N247);
nor NOR4 (N299, N296, N230, N277, N81);
buf BUF1 (N300, N293);
buf BUF1 (N301, N287);
buf BUF1 (N302, N295);
and AND2 (N303, N302, N7);
or OR3 (N304, N300, N179, N101);
buf BUF1 (N305, N294);
not NOT1 (N306, N291);
buf BUF1 (N307, N303);
or OR2 (N308, N306, N245);
nand NAND4 (N309, N289, N137, N180, N160);
and AND3 (N310, N297, N112, N60);
nor NOR3 (N311, N305, N111, N204);
buf BUF1 (N312, N298);
buf BUF1 (N313, N301);
or OR4 (N314, N309, N101, N59, N139);
and AND4 (N315, N310, N195, N305, N220);
nor NOR3 (N316, N314, N161, N67);
or OR2 (N317, N299, N225);
nand NAND4 (N318, N317, N256, N150, N104);
not NOT1 (N319, N312);
xor XOR2 (N320, N316, N47);
nand NAND3 (N321, N318, N50, N37);
nand NAND3 (N322, N320, N123, N283);
buf BUF1 (N323, N307);
nand NAND4 (N324, N321, N279, N135, N132);
xor XOR2 (N325, N319, N316);
or OR3 (N326, N311, N96, N96);
and AND4 (N327, N322, N164, N223, N65);
nor NOR2 (N328, N327, N108);
or OR2 (N329, N326, N28);
xor XOR2 (N330, N264, N119);
nor NOR2 (N331, N324, N40);
nand NAND2 (N332, N328, N13);
nor NOR4 (N333, N323, N167, N252, N268);
or OR2 (N334, N313, N271);
and AND3 (N335, N315, N120, N14);
buf BUF1 (N336, N304);
nand NAND2 (N337, N332, N70);
or OR2 (N338, N308, N135);
xor XOR2 (N339, N325, N203);
not NOT1 (N340, N331);
xor XOR2 (N341, N338, N140);
buf BUF1 (N342, N330);
not NOT1 (N343, N329);
and AND3 (N344, N337, N102, N57);
buf BUF1 (N345, N344);
nand NAND3 (N346, N340, N171, N51);
xor XOR2 (N347, N343, N287);
xor XOR2 (N348, N347, N74);
nand NAND3 (N349, N341, N270, N247);
buf BUF1 (N350, N334);
not NOT1 (N351, N349);
xor XOR2 (N352, N345, N43);
or OR3 (N353, N333, N201, N125);
nor NOR4 (N354, N350, N289, N4, N65);
or OR4 (N355, N342, N3, N340, N305);
not NOT1 (N356, N354);
buf BUF1 (N357, N346);
not NOT1 (N358, N357);
xor XOR2 (N359, N339, N71);
buf BUF1 (N360, N353);
or OR4 (N361, N335, N269, N337, N308);
buf BUF1 (N362, N348);
nand NAND2 (N363, N336, N260);
xor XOR2 (N364, N363, N67);
or OR4 (N365, N352, N125, N300, N144);
not NOT1 (N366, N360);
xor XOR2 (N367, N351, N80);
nor NOR4 (N368, N359, N56, N263, N80);
or OR3 (N369, N361, N234, N180);
xor XOR2 (N370, N362, N322);
and AND3 (N371, N370, N256, N342);
or OR3 (N372, N371, N41, N295);
nor NOR4 (N373, N358, N218, N38, N149);
buf BUF1 (N374, N356);
xor XOR2 (N375, N364, N305);
nand NAND2 (N376, N372, N317);
buf BUF1 (N377, N376);
buf BUF1 (N378, N375);
not NOT1 (N379, N355);
and AND4 (N380, N365, N286, N207, N335);
nor NOR3 (N381, N368, N379, N197);
nand NAND4 (N382, N266, N138, N310, N287);
nand NAND2 (N383, N381, N213);
nor NOR2 (N384, N382, N284);
nand NAND2 (N385, N383, N309);
not NOT1 (N386, N378);
or OR2 (N387, N367, N174);
buf BUF1 (N388, N377);
and AND2 (N389, N388, N322);
nand NAND2 (N390, N389, N103);
xor XOR2 (N391, N380, N50);
or OR4 (N392, N390, N243, N83, N142);
nand NAND4 (N393, N385, N252, N92, N42);
not NOT1 (N394, N392);
not NOT1 (N395, N394);
and AND4 (N396, N369, N323, N275, N293);
nor NOR4 (N397, N395, N149, N379, N174);
xor XOR2 (N398, N374, N166);
not NOT1 (N399, N396);
xor XOR2 (N400, N397, N274);
or OR2 (N401, N400, N18);
or OR4 (N402, N393, N286, N18, N344);
or OR2 (N403, N391, N190);
or OR2 (N404, N403, N229);
xor XOR2 (N405, N399, N65);
buf BUF1 (N406, N386);
buf BUF1 (N407, N405);
not NOT1 (N408, N384);
not NOT1 (N409, N401);
buf BUF1 (N410, N366);
xor XOR2 (N411, N408, N382);
and AND3 (N412, N406, N166, N313);
or OR4 (N413, N398, N134, N335, N26);
nand NAND2 (N414, N407, N358);
and AND3 (N415, N412, N148, N214);
and AND2 (N416, N415, N227);
and AND4 (N417, N373, N96, N404, N323);
or OR3 (N418, N341, N385, N302);
or OR4 (N419, N416, N69, N168, N340);
xor XOR2 (N420, N413, N133);
nor NOR3 (N421, N411, N230, N51);
and AND3 (N422, N409, N8, N127);
nand NAND3 (N423, N422, N84, N99);
and AND4 (N424, N417, N279, N4, N295);
or OR2 (N425, N387, N190);
not NOT1 (N426, N423);
xor XOR2 (N427, N426, N82);
not NOT1 (N428, N421);
buf BUF1 (N429, N428);
nand NAND2 (N430, N429, N50);
or OR2 (N431, N424, N396);
not NOT1 (N432, N427);
nor NOR4 (N433, N410, N20, N175, N344);
nand NAND2 (N434, N402, N364);
nand NAND2 (N435, N433, N14);
nor NOR3 (N436, N419, N412, N15);
nor NOR4 (N437, N435, N196, N306, N342);
nor NOR2 (N438, N414, N193);
or OR3 (N439, N431, N421, N74);
or OR3 (N440, N432, N46, N304);
xor XOR2 (N441, N420, N11);
nand NAND3 (N442, N430, N148, N195);
nand NAND2 (N443, N437, N231);
nor NOR3 (N444, N425, N329, N223);
nand NAND3 (N445, N436, N344, N272);
xor XOR2 (N446, N434, N37);
buf BUF1 (N447, N445);
buf BUF1 (N448, N447);
nand NAND4 (N449, N440, N102, N347, N261);
not NOT1 (N450, N446);
or OR3 (N451, N450, N434, N295);
nor NOR4 (N452, N438, N367, N370, N273);
and AND2 (N453, N444, N233);
buf BUF1 (N454, N439);
xor XOR2 (N455, N449, N338);
or OR2 (N456, N452, N291);
buf BUF1 (N457, N454);
buf BUF1 (N458, N455);
or OR3 (N459, N456, N304, N412);
buf BUF1 (N460, N453);
buf BUF1 (N461, N457);
and AND4 (N462, N451, N32, N409, N77);
xor XOR2 (N463, N442, N456);
not NOT1 (N464, N460);
buf BUF1 (N465, N464);
buf BUF1 (N466, N461);
or OR3 (N467, N459, N288, N423);
xor XOR2 (N468, N467, N92);
nor NOR4 (N469, N463, N383, N363, N365);
xor XOR2 (N470, N468, N147);
not NOT1 (N471, N441);
and AND2 (N472, N443, N220);
nor NOR4 (N473, N462, N90, N304, N442);
xor XOR2 (N474, N458, N44);
nor NOR4 (N475, N470, N129, N183, N33);
nand NAND4 (N476, N418, N288, N300, N118);
nand NAND4 (N477, N469, N241, N124, N328);
not NOT1 (N478, N474);
or OR2 (N479, N465, N308);
nand NAND4 (N480, N473, N270, N138, N186);
xor XOR2 (N481, N475, N160);
not NOT1 (N482, N466);
nor NOR3 (N483, N481, N374, N278);
nor NOR3 (N484, N476, N263, N477);
nand NAND4 (N485, N5, N221, N474, N324);
and AND3 (N486, N485, N181, N141);
not NOT1 (N487, N478);
xor XOR2 (N488, N482, N353);
or OR4 (N489, N472, N422, N409, N405);
nor NOR2 (N490, N479, N357);
and AND3 (N491, N488, N69, N357);
buf BUF1 (N492, N484);
not NOT1 (N493, N489);
not NOT1 (N494, N493);
not NOT1 (N495, N487);
xor XOR2 (N496, N492, N79);
nor NOR3 (N497, N448, N49, N76);
or OR3 (N498, N480, N403, N234);
nor NOR3 (N499, N498, N285, N362);
or OR3 (N500, N471, N247, N442);
xor XOR2 (N501, N491, N257);
or OR2 (N502, N494, N500);
xor XOR2 (N503, N62, N98);
xor XOR2 (N504, N496, N87);
nor NOR3 (N505, N495, N203, N333);
and AND2 (N506, N486, N76);
not NOT1 (N507, N506);
buf BUF1 (N508, N504);
xor XOR2 (N509, N502, N53);
nor NOR2 (N510, N507, N82);
xor XOR2 (N511, N508, N218);
buf BUF1 (N512, N501);
nand NAND2 (N513, N497, N146);
and AND2 (N514, N490, N484);
xor XOR2 (N515, N510, N418);
xor XOR2 (N516, N515, N34);
buf BUF1 (N517, N512);
nor NOR2 (N518, N505, N361);
buf BUF1 (N519, N511);
not NOT1 (N520, N499);
nand NAND2 (N521, N520, N39);
nor NOR4 (N522, N517, N104, N509, N32);
nand NAND4 (N523, N6, N159, N100, N34);
not NOT1 (N524, N519);
nand NAND3 (N525, N483, N107, N342);
or OR3 (N526, N514, N158, N310);
or OR4 (N527, N526, N427, N442, N105);
not NOT1 (N528, N522);
or OR4 (N529, N516, N77, N100, N329);
nand NAND4 (N530, N525, N112, N459, N369);
nand NAND4 (N531, N528, N31, N235, N102);
and AND4 (N532, N527, N144, N150, N408);
and AND2 (N533, N530, N63);
buf BUF1 (N534, N529);
xor XOR2 (N535, N521, N14);
not NOT1 (N536, N534);
and AND4 (N537, N531, N492, N193, N372);
and AND3 (N538, N523, N187, N61);
nor NOR2 (N539, N538, N295);
buf BUF1 (N540, N537);
buf BUF1 (N541, N536);
or OR2 (N542, N540, N256);
not NOT1 (N543, N541);
and AND2 (N544, N539, N176);
nand NAND2 (N545, N513, N5);
or OR4 (N546, N543, N273, N36, N160);
nor NOR3 (N547, N545, N520, N1);
nor NOR4 (N548, N535, N191, N182, N77);
or OR2 (N549, N503, N31);
and AND4 (N550, N548, N248, N89, N442);
not NOT1 (N551, N547);
xor XOR2 (N552, N546, N151);
buf BUF1 (N553, N549);
not NOT1 (N554, N553);
and AND4 (N555, N542, N12, N374, N458);
and AND3 (N556, N555, N539, N370);
buf BUF1 (N557, N544);
and AND2 (N558, N532, N273);
and AND3 (N559, N554, N413, N333);
not NOT1 (N560, N556);
nor NOR3 (N561, N560, N474, N81);
and AND2 (N562, N559, N296);
nand NAND2 (N563, N550, N280);
and AND2 (N564, N518, N409);
or OR3 (N565, N558, N538, N338);
buf BUF1 (N566, N552);
and AND2 (N567, N551, N97);
xor XOR2 (N568, N524, N134);
nand NAND2 (N569, N563, N290);
nor NOR2 (N570, N568, N531);
nor NOR2 (N571, N533, N408);
xor XOR2 (N572, N569, N487);
not NOT1 (N573, N572);
and AND2 (N574, N562, N478);
buf BUF1 (N575, N574);
nor NOR4 (N576, N567, N387, N271, N546);
xor XOR2 (N577, N575, N239);
nor NOR2 (N578, N577, N453);
nor NOR2 (N579, N565, N501);
buf BUF1 (N580, N573);
nand NAND2 (N581, N578, N98);
or OR4 (N582, N561, N466, N367, N73);
nand NAND2 (N583, N566, N244);
nor NOR4 (N584, N570, N110, N198, N515);
or OR4 (N585, N580, N405, N429, N128);
or OR2 (N586, N564, N82);
nand NAND3 (N587, N576, N105, N18);
xor XOR2 (N588, N581, N300);
xor XOR2 (N589, N583, N555);
nand NAND3 (N590, N585, N310, N79);
xor XOR2 (N591, N557, N194);
xor XOR2 (N592, N584, N530);
xor XOR2 (N593, N590, N561);
nand NAND3 (N594, N571, N572, N68);
not NOT1 (N595, N586);
buf BUF1 (N596, N593);
buf BUF1 (N597, N587);
and AND3 (N598, N579, N349, N558);
nand NAND4 (N599, N594, N241, N541, N319);
nor NOR4 (N600, N599, N347, N197, N519);
or OR4 (N601, N596, N3, N20, N577);
xor XOR2 (N602, N598, N411);
buf BUF1 (N603, N592);
nor NOR3 (N604, N597, N560, N17);
xor XOR2 (N605, N603, N32);
nor NOR3 (N606, N591, N350, N89);
or OR4 (N607, N604, N579, N421, N408);
or OR3 (N608, N607, N337, N521);
nand NAND4 (N609, N608, N379, N128, N172);
buf BUF1 (N610, N606);
and AND3 (N611, N610, N440, N484);
buf BUF1 (N612, N602);
and AND2 (N613, N601, N403);
or OR2 (N614, N605, N555);
buf BUF1 (N615, N611);
or OR4 (N616, N582, N576, N408, N335);
and AND3 (N617, N600, N26, N42);
or OR2 (N618, N617, N550);
nor NOR3 (N619, N614, N276, N310);
nor NOR4 (N620, N613, N144, N86, N259);
xor XOR2 (N621, N589, N122);
or OR3 (N622, N609, N575, N614);
not NOT1 (N623, N595);
xor XOR2 (N624, N588, N447);
xor XOR2 (N625, N623, N275);
nor NOR3 (N626, N622, N101, N204);
not NOT1 (N627, N618);
buf BUF1 (N628, N626);
buf BUF1 (N629, N620);
and AND3 (N630, N627, N487, N166);
nor NOR2 (N631, N612, N160);
nand NAND4 (N632, N619, N221, N440, N83);
nor NOR4 (N633, N632, N184, N629, N273);
and AND3 (N634, N118, N112, N622);
and AND3 (N635, N625, N1, N515);
buf BUF1 (N636, N615);
or OR3 (N637, N635, N28, N441);
not NOT1 (N638, N633);
buf BUF1 (N639, N624);
xor XOR2 (N640, N639, N567);
xor XOR2 (N641, N631, N361);
nand NAND4 (N642, N628, N511, N11, N511);
not NOT1 (N643, N616);
or OR4 (N644, N621, N195, N281, N531);
not NOT1 (N645, N636);
nor NOR3 (N646, N640, N160, N246);
xor XOR2 (N647, N637, N30);
and AND4 (N648, N646, N455, N641, N479);
nor NOR3 (N649, N386, N423, N534);
or OR4 (N650, N647, N57, N449, N82);
buf BUF1 (N651, N630);
xor XOR2 (N652, N644, N521);
buf BUF1 (N653, N652);
or OR2 (N654, N643, N627);
xor XOR2 (N655, N634, N69);
buf BUF1 (N656, N642);
and AND4 (N657, N655, N602, N409, N615);
xor XOR2 (N658, N645, N604);
and AND3 (N659, N657, N84, N605);
not NOT1 (N660, N656);
and AND4 (N661, N651, N146, N311, N533);
nor NOR3 (N662, N654, N356, N165);
or OR3 (N663, N649, N57, N170);
or OR3 (N664, N658, N638, N119);
and AND3 (N665, N508, N249, N424);
or OR4 (N666, N663, N459, N167, N204);
or OR2 (N667, N659, N555);
and AND3 (N668, N665, N642, N121);
and AND3 (N669, N653, N510, N61);
nor NOR2 (N670, N660, N355);
not NOT1 (N671, N667);
nand NAND2 (N672, N666, N372);
not NOT1 (N673, N664);
xor XOR2 (N674, N648, N509);
nor NOR2 (N675, N661, N200);
nand NAND4 (N676, N669, N502, N245, N120);
buf BUF1 (N677, N674);
nand NAND4 (N678, N673, N273, N412, N238);
or OR2 (N679, N670, N545);
and AND3 (N680, N671, N553, N172);
or OR4 (N681, N676, N384, N172, N653);
nor NOR3 (N682, N677, N74, N295);
xor XOR2 (N683, N679, N655);
xor XOR2 (N684, N678, N643);
or OR4 (N685, N662, N385, N603, N25);
or OR4 (N686, N684, N134, N599, N446);
nor NOR4 (N687, N675, N335, N40, N7);
and AND2 (N688, N681, N279);
or OR2 (N689, N687, N568);
nand NAND2 (N690, N688, N228);
not NOT1 (N691, N680);
xor XOR2 (N692, N689, N255);
not NOT1 (N693, N686);
nor NOR2 (N694, N691, N119);
nand NAND2 (N695, N693, N62);
nor NOR3 (N696, N668, N462, N71);
buf BUF1 (N697, N690);
not NOT1 (N698, N697);
xor XOR2 (N699, N698, N149);
nand NAND2 (N700, N650, N68);
or OR2 (N701, N699, N102);
xor XOR2 (N702, N700, N52);
nand NAND2 (N703, N682, N477);
and AND3 (N704, N672, N499, N657);
and AND3 (N705, N696, N352, N197);
and AND2 (N706, N695, N11);
not NOT1 (N707, N702);
buf BUF1 (N708, N694);
not NOT1 (N709, N705);
nand NAND4 (N710, N709, N405, N81, N651);
or OR4 (N711, N692, N656, N209, N662);
buf BUF1 (N712, N707);
and AND3 (N713, N701, N174, N190);
or OR3 (N714, N703, N298, N365);
or OR3 (N715, N685, N694, N187);
xor XOR2 (N716, N712, N218);
not NOT1 (N717, N714);
nand NAND3 (N718, N706, N373, N145);
xor XOR2 (N719, N710, N193);
nand NAND4 (N720, N683, N319, N236, N67);
xor XOR2 (N721, N717, N168);
xor XOR2 (N722, N715, N586);
or OR3 (N723, N711, N280, N277);
or OR3 (N724, N716, N86, N395);
or OR3 (N725, N718, N400, N281);
nor NOR2 (N726, N719, N289);
or OR4 (N727, N704, N393, N15, N270);
xor XOR2 (N728, N726, N497);
nand NAND3 (N729, N728, N489, N516);
and AND2 (N730, N708, N267);
buf BUF1 (N731, N724);
buf BUF1 (N732, N731);
not NOT1 (N733, N727);
nor NOR4 (N734, N723, N276, N332, N319);
not NOT1 (N735, N730);
xor XOR2 (N736, N722, N612);
xor XOR2 (N737, N720, N551);
xor XOR2 (N738, N713, N522);
not NOT1 (N739, N737);
nand NAND2 (N740, N739, N363);
xor XOR2 (N741, N738, N697);
not NOT1 (N742, N733);
nor NOR4 (N743, N742, N366, N222, N533);
nor NOR2 (N744, N741, N73);
not NOT1 (N745, N732);
buf BUF1 (N746, N736);
buf BUF1 (N747, N734);
nand NAND2 (N748, N735, N256);
xor XOR2 (N749, N748, N722);
nor NOR3 (N750, N746, N380, N338);
xor XOR2 (N751, N721, N585);
nand NAND4 (N752, N745, N64, N601, N736);
xor XOR2 (N753, N750, N675);
and AND3 (N754, N753, N193, N700);
not NOT1 (N755, N754);
and AND3 (N756, N744, N553, N213);
buf BUF1 (N757, N729);
and AND2 (N758, N757, N224);
xor XOR2 (N759, N755, N639);
nand NAND2 (N760, N743, N258);
nand NAND4 (N761, N751, N281, N497, N350);
or OR4 (N762, N725, N463, N199, N511);
xor XOR2 (N763, N749, N523);
nor NOR3 (N764, N761, N6, N587);
not NOT1 (N765, N752);
or OR3 (N766, N747, N751, N718);
nor NOR2 (N767, N760, N53);
buf BUF1 (N768, N763);
nor NOR2 (N769, N758, N206);
not NOT1 (N770, N764);
not NOT1 (N771, N762);
and AND2 (N772, N766, N727);
nor NOR4 (N773, N767, N193, N407, N515);
xor XOR2 (N774, N740, N476);
nand NAND3 (N775, N773, N662, N66);
xor XOR2 (N776, N768, N360);
or OR4 (N777, N771, N603, N289, N414);
nand NAND2 (N778, N777, N362);
and AND2 (N779, N778, N471);
nand NAND3 (N780, N779, N76, N482);
and AND3 (N781, N780, N507, N334);
buf BUF1 (N782, N775);
not NOT1 (N783, N782);
nor NOR3 (N784, N756, N482, N720);
not NOT1 (N785, N781);
nor NOR3 (N786, N770, N34, N303);
nand NAND3 (N787, N772, N598, N185);
buf BUF1 (N788, N765);
xor XOR2 (N789, N776, N1);
xor XOR2 (N790, N769, N175);
and AND2 (N791, N789, N500);
and AND2 (N792, N790, N110);
xor XOR2 (N793, N759, N579);
and AND4 (N794, N784, N495, N438, N23);
nor NOR4 (N795, N788, N76, N592, N114);
not NOT1 (N796, N792);
nand NAND4 (N797, N783, N70, N310, N518);
nand NAND3 (N798, N794, N607, N667);
buf BUF1 (N799, N786);
buf BUF1 (N800, N791);
and AND3 (N801, N799, N312, N363);
nor NOR2 (N802, N785, N751);
and AND2 (N803, N796, N578);
and AND3 (N804, N798, N386, N171);
nor NOR4 (N805, N787, N67, N567, N381);
or OR4 (N806, N802, N136, N119, N362);
and AND3 (N807, N805, N753, N355);
not NOT1 (N808, N793);
or OR3 (N809, N797, N168, N411);
nand NAND3 (N810, N809, N789, N52);
or OR4 (N811, N774, N780, N285, N550);
or OR3 (N812, N811, N670, N260);
nor NOR4 (N813, N807, N95, N425, N165);
or OR3 (N814, N813, N143, N393);
and AND4 (N815, N803, N811, N505, N156);
nor NOR3 (N816, N801, N449, N781);
nor NOR3 (N817, N800, N695, N815);
nor NOR3 (N818, N243, N786, N614);
nand NAND3 (N819, N804, N12, N25);
nor NOR4 (N820, N816, N225, N536, N78);
xor XOR2 (N821, N812, N675);
xor XOR2 (N822, N819, N219);
nand NAND3 (N823, N810, N632, N268);
and AND4 (N824, N821, N575, N563, N298);
nand NAND2 (N825, N795, N55);
xor XOR2 (N826, N806, N173);
and AND4 (N827, N814, N750, N766, N674);
and AND3 (N828, N824, N313, N72);
buf BUF1 (N829, N808);
buf BUF1 (N830, N818);
nand NAND3 (N831, N830, N31, N392);
and AND2 (N832, N828, N771);
xor XOR2 (N833, N823, N670);
buf BUF1 (N834, N833);
buf BUF1 (N835, N817);
buf BUF1 (N836, N831);
xor XOR2 (N837, N836, N753);
nor NOR4 (N838, N820, N146, N314, N225);
xor XOR2 (N839, N826, N689);
buf BUF1 (N840, N822);
buf BUF1 (N841, N837);
or OR3 (N842, N825, N729, N781);
and AND4 (N843, N835, N403, N161, N776);
nor NOR4 (N844, N842, N400, N79, N559);
xor XOR2 (N845, N841, N224);
nand NAND2 (N846, N839, N332);
nor NOR4 (N847, N846, N248, N7, N830);
nand NAND2 (N848, N832, N273);
nor NOR4 (N849, N845, N154, N503, N687);
xor XOR2 (N850, N840, N491);
xor XOR2 (N851, N838, N799);
and AND4 (N852, N848, N155, N383, N591);
nor NOR2 (N853, N851, N721);
and AND3 (N854, N844, N68, N758);
or OR2 (N855, N829, N715);
buf BUF1 (N856, N850);
not NOT1 (N857, N834);
or OR4 (N858, N854, N803, N122, N265);
and AND2 (N859, N847, N264);
xor XOR2 (N860, N857, N620);
nand NAND4 (N861, N852, N113, N766, N13);
and AND4 (N862, N849, N634, N64, N810);
nand NAND2 (N863, N856, N648);
not NOT1 (N864, N860);
nand NAND4 (N865, N862, N335, N440, N524);
or OR3 (N866, N858, N712, N422);
buf BUF1 (N867, N863);
and AND4 (N868, N859, N865, N634, N311);
nand NAND3 (N869, N560, N563, N420);
buf BUF1 (N870, N866);
buf BUF1 (N871, N869);
nand NAND2 (N872, N868, N767);
not NOT1 (N873, N872);
not NOT1 (N874, N871);
buf BUF1 (N875, N867);
nand NAND2 (N876, N861, N404);
not NOT1 (N877, N874);
nor NOR3 (N878, N875, N122, N284);
not NOT1 (N879, N864);
nand NAND4 (N880, N827, N801, N552, N124);
xor XOR2 (N881, N880, N846);
xor XOR2 (N882, N870, N310);
xor XOR2 (N883, N878, N357);
and AND3 (N884, N882, N710, N38);
and AND4 (N885, N884, N802, N208, N22);
buf BUF1 (N886, N843);
and AND4 (N887, N873, N453, N520, N156);
not NOT1 (N888, N877);
xor XOR2 (N889, N879, N614);
xor XOR2 (N890, N889, N263);
not NOT1 (N891, N883);
nand NAND4 (N892, N853, N697, N398, N693);
or OR4 (N893, N886, N5, N643, N311);
xor XOR2 (N894, N876, N85);
buf BUF1 (N895, N887);
not NOT1 (N896, N893);
buf BUF1 (N897, N855);
xor XOR2 (N898, N897, N22);
buf BUF1 (N899, N894);
xor XOR2 (N900, N895, N781);
or OR3 (N901, N891, N193, N171);
and AND2 (N902, N898, N608);
nand NAND4 (N903, N900, N404, N286, N416);
or OR3 (N904, N892, N702, N770);
nand NAND3 (N905, N890, N41, N585);
or OR4 (N906, N902, N772, N577, N167);
buf BUF1 (N907, N903);
nor NOR3 (N908, N888, N136, N167);
nor NOR2 (N909, N905, N189);
xor XOR2 (N910, N896, N435);
nor NOR4 (N911, N908, N46, N201, N299);
not NOT1 (N912, N910);
nand NAND4 (N913, N912, N834, N769, N227);
or OR4 (N914, N906, N223, N436, N130);
xor XOR2 (N915, N901, N583);
nor NOR4 (N916, N915, N529, N905, N795);
nand NAND4 (N917, N911, N902, N228, N651);
buf BUF1 (N918, N899);
or OR4 (N919, N914, N821, N566, N547);
xor XOR2 (N920, N919, N397);
xor XOR2 (N921, N918, N216);
nor NOR2 (N922, N909, N409);
xor XOR2 (N923, N920, N783);
and AND3 (N924, N923, N705, N721);
or OR3 (N925, N881, N797, N463);
nor NOR4 (N926, N904, N303, N151, N344);
and AND4 (N927, N907, N311, N467, N711);
nand NAND3 (N928, N913, N410, N559);
buf BUF1 (N929, N926);
and AND3 (N930, N928, N625, N772);
buf BUF1 (N931, N924);
and AND2 (N932, N925, N661);
not NOT1 (N933, N921);
and AND3 (N934, N922, N360, N137);
not NOT1 (N935, N934);
buf BUF1 (N936, N929);
and AND4 (N937, N917, N5, N341, N777);
xor XOR2 (N938, N932, N852);
nand NAND4 (N939, N931, N173, N230, N13);
nand NAND2 (N940, N938, N797);
nand NAND2 (N941, N935, N857);
or OR3 (N942, N927, N42, N680);
and AND4 (N943, N916, N57, N235, N336);
not NOT1 (N944, N940);
xor XOR2 (N945, N943, N940);
buf BUF1 (N946, N942);
nor NOR2 (N947, N946, N773);
and AND4 (N948, N930, N286, N597, N940);
or OR4 (N949, N945, N162, N332, N6);
and AND4 (N950, N941, N530, N372, N852);
buf BUF1 (N951, N939);
buf BUF1 (N952, N944);
not NOT1 (N953, N936);
xor XOR2 (N954, N950, N765);
buf BUF1 (N955, N948);
and AND4 (N956, N949, N856, N143, N386);
and AND3 (N957, N937, N689, N560);
and AND3 (N958, N885, N714, N631);
nor NOR2 (N959, N954, N393);
or OR2 (N960, N951, N807);
buf BUF1 (N961, N947);
nand NAND4 (N962, N961, N613, N421, N52);
xor XOR2 (N963, N955, N773);
buf BUF1 (N964, N957);
buf BUF1 (N965, N964);
nor NOR2 (N966, N953, N908);
and AND2 (N967, N962, N303);
buf BUF1 (N968, N959);
nand NAND4 (N969, N956, N169, N29, N581);
not NOT1 (N970, N963);
not NOT1 (N971, N966);
nand NAND3 (N972, N933, N418, N6);
and AND2 (N973, N971, N761);
nor NOR2 (N974, N968, N370);
buf BUF1 (N975, N970);
nor NOR3 (N976, N973, N792, N386);
or OR2 (N977, N958, N862);
nand NAND2 (N978, N974, N61);
nor NOR3 (N979, N965, N395, N795);
or OR4 (N980, N960, N553, N119, N906);
nor NOR4 (N981, N978, N287, N524, N92);
nand NAND4 (N982, N952, N814, N835, N419);
not NOT1 (N983, N975);
and AND4 (N984, N983, N887, N446, N787);
nor NOR2 (N985, N984, N131);
nand NAND3 (N986, N972, N270, N792);
or OR2 (N987, N986, N697);
xor XOR2 (N988, N980, N14);
not NOT1 (N989, N982);
nor NOR3 (N990, N981, N830, N230);
buf BUF1 (N991, N988);
not NOT1 (N992, N985);
xor XOR2 (N993, N969, N820);
xor XOR2 (N994, N967, N737);
or OR4 (N995, N987, N134, N844, N526);
xor XOR2 (N996, N989, N477);
not NOT1 (N997, N977);
nand NAND2 (N998, N994, N804);
nand NAND2 (N999, N993, N897);
nand NAND2 (N1000, N991, N650);
xor XOR2 (N1001, N995, N998);
buf BUF1 (N1002, N794);
buf BUF1 (N1003, N999);
and AND4 (N1004, N1003, N163, N35, N35);
nand NAND3 (N1005, N979, N707, N512);
buf BUF1 (N1006, N996);
not NOT1 (N1007, N1000);
buf BUF1 (N1008, N990);
and AND3 (N1009, N1007, N816, N342);
or OR2 (N1010, N1005, N370);
or OR4 (N1011, N992, N890, N217, N479);
nor NOR2 (N1012, N1011, N505);
or OR3 (N1013, N1001, N427, N398);
not NOT1 (N1014, N997);
xor XOR2 (N1015, N1004, N567);
and AND2 (N1016, N1006, N207);
nand NAND2 (N1017, N1002, N796);
nor NOR2 (N1018, N1017, N855);
nor NOR2 (N1019, N1015, N41);
xor XOR2 (N1020, N976, N70);
xor XOR2 (N1021, N1020, N557);
or OR4 (N1022, N1016, N427, N687, N629);
and AND4 (N1023, N1019, N271, N153, N876);
and AND4 (N1024, N1023, N189, N1013, N678);
nand NAND3 (N1025, N834, N696, N422);
nand NAND2 (N1026, N1018, N763);
nor NOR4 (N1027, N1014, N134, N957, N687);
not NOT1 (N1028, N1024);
not NOT1 (N1029, N1028);
nand NAND3 (N1030, N1025, N886, N442);
nor NOR4 (N1031, N1012, N779, N108, N821);
nor NOR3 (N1032, N1031, N84, N243);
nor NOR3 (N1033, N1008, N501, N753);
xor XOR2 (N1034, N1032, N276);
nand NAND2 (N1035, N1030, N369);
and AND2 (N1036, N1026, N666);
nor NOR2 (N1037, N1033, N316);
not NOT1 (N1038, N1036);
buf BUF1 (N1039, N1037);
not NOT1 (N1040, N1022);
buf BUF1 (N1041, N1038);
or OR2 (N1042, N1035, N575);
nor NOR2 (N1043, N1039, N440);
or OR2 (N1044, N1042, N823);
or OR4 (N1045, N1040, N148, N300, N766);
not NOT1 (N1046, N1021);
not NOT1 (N1047, N1046);
xor XOR2 (N1048, N1010, N709);
or OR4 (N1049, N1034, N551, N437, N202);
buf BUF1 (N1050, N1041);
not NOT1 (N1051, N1043);
xor XOR2 (N1052, N1044, N259);
buf BUF1 (N1053, N1029);
xor XOR2 (N1054, N1051, N548);
buf BUF1 (N1055, N1009);
and AND4 (N1056, N1049, N150, N51, N35);
or OR3 (N1057, N1054, N1014, N420);
nor NOR4 (N1058, N1053, N402, N405, N157);
and AND3 (N1059, N1050, N481, N637);
nor NOR4 (N1060, N1059, N75, N982, N998);
and AND3 (N1061, N1027, N13, N617);
nand NAND3 (N1062, N1060, N775, N877);
nor NOR4 (N1063, N1048, N692, N660, N1056);
buf BUF1 (N1064, N625);
not NOT1 (N1065, N1052);
xor XOR2 (N1066, N1047, N281);
or OR4 (N1067, N1064, N273, N432, N80);
nor NOR3 (N1068, N1063, N711, N399);
or OR2 (N1069, N1065, N228);
nand NAND4 (N1070, N1067, N537, N339, N703);
buf BUF1 (N1071, N1058);
nor NOR3 (N1072, N1071, N747, N529);
and AND2 (N1073, N1069, N57);
nor NOR4 (N1074, N1066, N108, N760, N233);
and AND4 (N1075, N1073, N501, N118, N963);
and AND2 (N1076, N1074, N823);
nor NOR4 (N1077, N1070, N310, N227, N600);
and AND3 (N1078, N1062, N489, N859);
or OR4 (N1079, N1068, N1044, N596, N403);
or OR4 (N1080, N1061, N150, N1007, N332);
not NOT1 (N1081, N1080);
or OR2 (N1082, N1057, N766);
xor XOR2 (N1083, N1077, N249);
or OR4 (N1084, N1079, N472, N398, N295);
or OR3 (N1085, N1072, N326, N632);
nand NAND2 (N1086, N1078, N247);
nor NOR3 (N1087, N1084, N473, N255);
nor NOR3 (N1088, N1087, N603, N508);
or OR4 (N1089, N1075, N422, N555, N709);
buf BUF1 (N1090, N1083);
or OR3 (N1091, N1081, N892, N568);
or OR4 (N1092, N1045, N96, N930, N381);
xor XOR2 (N1093, N1088, N457);
nand NAND2 (N1094, N1092, N716);
and AND3 (N1095, N1085, N270, N763);
and AND3 (N1096, N1090, N203, N1054);
buf BUF1 (N1097, N1055);
nor NOR4 (N1098, N1097, N500, N1089, N388);
and AND2 (N1099, N648, N1019);
nand NAND4 (N1100, N1095, N1063, N1021, N315);
not NOT1 (N1101, N1086);
nor NOR3 (N1102, N1101, N697, N71);
and AND3 (N1103, N1102, N1052, N522);
xor XOR2 (N1104, N1096, N572);
nor NOR3 (N1105, N1091, N1067, N292);
not NOT1 (N1106, N1098);
xor XOR2 (N1107, N1099, N504);
nor NOR4 (N1108, N1106, N485, N21, N47);
buf BUF1 (N1109, N1108);
nand NAND4 (N1110, N1076, N17, N704, N13);
nand NAND3 (N1111, N1107, N133, N730);
buf BUF1 (N1112, N1103);
and AND2 (N1113, N1110, N295);
not NOT1 (N1114, N1112);
and AND2 (N1115, N1114, N577);
xor XOR2 (N1116, N1113, N392);
buf BUF1 (N1117, N1094);
and AND4 (N1118, N1104, N429, N985, N989);
not NOT1 (N1119, N1117);
or OR2 (N1120, N1111, N687);
or OR4 (N1121, N1118, N742, N101, N1113);
nand NAND3 (N1122, N1109, N70, N567);
nand NAND2 (N1123, N1119, N854);
xor XOR2 (N1124, N1100, N799);
or OR3 (N1125, N1105, N270, N405);
and AND3 (N1126, N1124, N1001, N941);
buf BUF1 (N1127, N1126);
and AND3 (N1128, N1115, N774, N682);
and AND3 (N1129, N1082, N1011, N422);
xor XOR2 (N1130, N1129, N349);
nor NOR2 (N1131, N1130, N270);
or OR4 (N1132, N1122, N1078, N1038, N932);
or OR4 (N1133, N1127, N365, N958, N492);
not NOT1 (N1134, N1123);
xor XOR2 (N1135, N1121, N691);
not NOT1 (N1136, N1133);
nand NAND4 (N1137, N1132, N551, N185, N888);
nor NOR2 (N1138, N1116, N1076);
xor XOR2 (N1139, N1135, N246);
or OR3 (N1140, N1137, N989, N1107);
or OR4 (N1141, N1125, N767, N967, N513);
and AND2 (N1142, N1141, N78);
nand NAND2 (N1143, N1134, N726);
buf BUF1 (N1144, N1136);
buf BUF1 (N1145, N1093);
xor XOR2 (N1146, N1144, N1066);
or OR2 (N1147, N1138, N64);
not NOT1 (N1148, N1131);
nand NAND4 (N1149, N1142, N113, N550, N547);
buf BUF1 (N1150, N1147);
nor NOR2 (N1151, N1145, N199);
not NOT1 (N1152, N1120);
or OR2 (N1153, N1148, N354);
nor NOR3 (N1154, N1139, N799, N329);
and AND2 (N1155, N1154, N648);
nand NAND2 (N1156, N1143, N749);
nand NAND4 (N1157, N1156, N903, N1100, N723);
or OR2 (N1158, N1128, N79);
not NOT1 (N1159, N1155);
and AND4 (N1160, N1140, N35, N180, N875);
nand NAND4 (N1161, N1153, N802, N1012, N558);
or OR4 (N1162, N1149, N819, N347, N485);
xor XOR2 (N1163, N1160, N691);
buf BUF1 (N1164, N1150);
nor NOR3 (N1165, N1164, N685, N189);
not NOT1 (N1166, N1162);
not NOT1 (N1167, N1161);
buf BUF1 (N1168, N1165);
nand NAND4 (N1169, N1168, N185, N495, N987);
or OR4 (N1170, N1157, N132, N18, N349);
not NOT1 (N1171, N1166);
not NOT1 (N1172, N1152);
nor NOR3 (N1173, N1172, N701, N309);
buf BUF1 (N1174, N1173);
buf BUF1 (N1175, N1159);
not NOT1 (N1176, N1169);
nor NOR3 (N1177, N1171, N629, N762);
nor NOR3 (N1178, N1146, N732, N906);
nand NAND2 (N1179, N1167, N875);
nand NAND4 (N1180, N1158, N462, N248, N660);
nor NOR2 (N1181, N1178, N1133);
nor NOR2 (N1182, N1174, N794);
nor NOR4 (N1183, N1177, N1065, N266, N1074);
xor XOR2 (N1184, N1176, N478);
nand NAND3 (N1185, N1182, N683, N1170);
or OR2 (N1186, N275, N811);
not NOT1 (N1187, N1179);
xor XOR2 (N1188, N1181, N768);
buf BUF1 (N1189, N1186);
not NOT1 (N1190, N1163);
buf BUF1 (N1191, N1185);
not NOT1 (N1192, N1184);
buf BUF1 (N1193, N1190);
and AND4 (N1194, N1180, N421, N619, N690);
xor XOR2 (N1195, N1191, N1083);
nor NOR3 (N1196, N1175, N892, N587);
not NOT1 (N1197, N1183);
nor NOR2 (N1198, N1195, N988);
not NOT1 (N1199, N1151);
nand NAND2 (N1200, N1198, N156);
nand NAND4 (N1201, N1200, N828, N324, N504);
and AND2 (N1202, N1188, N529);
or OR3 (N1203, N1193, N912, N515);
xor XOR2 (N1204, N1192, N515);
buf BUF1 (N1205, N1189);
and AND2 (N1206, N1187, N645);
xor XOR2 (N1207, N1199, N386);
and AND3 (N1208, N1194, N393, N601);
nand NAND2 (N1209, N1203, N923);
and AND4 (N1210, N1201, N495, N715, N646);
nor NOR4 (N1211, N1202, N388, N68, N869);
buf BUF1 (N1212, N1211);
not NOT1 (N1213, N1207);
or OR4 (N1214, N1197, N375, N1154, N170);
xor XOR2 (N1215, N1214, N115);
xor XOR2 (N1216, N1206, N334);
nand NAND2 (N1217, N1216, N1088);
buf BUF1 (N1218, N1217);
buf BUF1 (N1219, N1208);
buf BUF1 (N1220, N1196);
or OR4 (N1221, N1215, N1213, N317, N495);
xor XOR2 (N1222, N606, N1183);
xor XOR2 (N1223, N1220, N1101);
not NOT1 (N1224, N1205);
not NOT1 (N1225, N1222);
or OR4 (N1226, N1223, N1015, N417, N1198);
or OR2 (N1227, N1209, N701);
nand NAND2 (N1228, N1210, N623);
not NOT1 (N1229, N1218);
nor NOR2 (N1230, N1229, N926);
buf BUF1 (N1231, N1219);
buf BUF1 (N1232, N1212);
nor NOR2 (N1233, N1225, N832);
and AND3 (N1234, N1226, N1135, N929);
nor NOR4 (N1235, N1230, N139, N903, N816);
not NOT1 (N1236, N1228);
and AND3 (N1237, N1236, N244, N880);
buf BUF1 (N1238, N1233);
or OR2 (N1239, N1231, N564);
nand NAND4 (N1240, N1221, N774, N142, N1015);
nand NAND2 (N1241, N1240, N451);
nor NOR3 (N1242, N1238, N830, N1068);
nor NOR3 (N1243, N1234, N424, N222);
not NOT1 (N1244, N1235);
nor NOR2 (N1245, N1204, N1025);
or OR3 (N1246, N1242, N645, N103);
xor XOR2 (N1247, N1246, N162);
not NOT1 (N1248, N1239);
buf BUF1 (N1249, N1232);
nand NAND4 (N1250, N1249, N123, N709, N43);
buf BUF1 (N1251, N1224);
or OR3 (N1252, N1248, N412, N925);
nor NOR4 (N1253, N1237, N268, N313, N773);
xor XOR2 (N1254, N1245, N116);
and AND3 (N1255, N1254, N466, N627);
nand NAND3 (N1256, N1251, N799, N1075);
nand NAND3 (N1257, N1247, N1230, N810);
not NOT1 (N1258, N1227);
nor NOR2 (N1259, N1243, N1179);
nor NOR3 (N1260, N1259, N1237, N281);
nand NAND3 (N1261, N1255, N646, N143);
and AND3 (N1262, N1256, N865, N987);
nor NOR4 (N1263, N1241, N210, N707, N535);
nor NOR2 (N1264, N1253, N947);
nor NOR4 (N1265, N1260, N31, N473, N684);
nand NAND3 (N1266, N1264, N1244, N126);
xor XOR2 (N1267, N349, N1080);
not NOT1 (N1268, N1250);
buf BUF1 (N1269, N1266);
and AND2 (N1270, N1265, N1266);
nand NAND3 (N1271, N1262, N398, N465);
xor XOR2 (N1272, N1263, N227);
not NOT1 (N1273, N1261);
buf BUF1 (N1274, N1270);
xor XOR2 (N1275, N1267, N1265);
xor XOR2 (N1276, N1269, N389);
not NOT1 (N1277, N1272);
and AND4 (N1278, N1274, N566, N14, N1240);
nor NOR2 (N1279, N1271, N825);
and AND3 (N1280, N1257, N1253, N1083);
not NOT1 (N1281, N1276);
nor NOR3 (N1282, N1275, N955, N210);
or OR2 (N1283, N1273, N411);
or OR3 (N1284, N1281, N846, N709);
and AND3 (N1285, N1252, N297, N623);
xor XOR2 (N1286, N1280, N33);
or OR2 (N1287, N1279, N296);
not NOT1 (N1288, N1284);
xor XOR2 (N1289, N1286, N968);
nor NOR3 (N1290, N1289, N907, N456);
not NOT1 (N1291, N1277);
nor NOR4 (N1292, N1287, N668, N421, N4);
nor NOR2 (N1293, N1288, N899);
or OR2 (N1294, N1292, N1027);
or OR4 (N1295, N1291, N146, N345, N510);
and AND4 (N1296, N1293, N1023, N127, N564);
xor XOR2 (N1297, N1258, N446);
nor NOR2 (N1298, N1295, N961);
xor XOR2 (N1299, N1298, N108);
nand NAND2 (N1300, N1299, N267);
and AND4 (N1301, N1300, N108, N346, N275);
and AND3 (N1302, N1278, N1052, N804);
and AND3 (N1303, N1282, N97, N1236);
xor XOR2 (N1304, N1296, N613);
buf BUF1 (N1305, N1290);
buf BUF1 (N1306, N1285);
nor NOR2 (N1307, N1306, N993);
or OR2 (N1308, N1304, N2);
nand NAND2 (N1309, N1308, N656);
buf BUF1 (N1310, N1294);
buf BUF1 (N1311, N1268);
and AND3 (N1312, N1310, N1234, N82);
and AND4 (N1313, N1297, N794, N573, N704);
nand NAND3 (N1314, N1307, N920, N234);
nor NOR4 (N1315, N1303, N534, N721, N1091);
buf BUF1 (N1316, N1313);
buf BUF1 (N1317, N1315);
not NOT1 (N1318, N1317);
nor NOR4 (N1319, N1318, N730, N1179, N409);
buf BUF1 (N1320, N1309);
or OR3 (N1321, N1320, N640, N130);
nand NAND4 (N1322, N1283, N686, N483, N682);
and AND3 (N1323, N1319, N937, N725);
not NOT1 (N1324, N1311);
or OR2 (N1325, N1322, N483);
not NOT1 (N1326, N1314);
nor NOR3 (N1327, N1326, N167, N1050);
and AND2 (N1328, N1305, N982);
not NOT1 (N1329, N1328);
nor NOR3 (N1330, N1325, N1068, N38);
nand NAND3 (N1331, N1302, N1197, N950);
and AND3 (N1332, N1331, N310, N103);
xor XOR2 (N1333, N1327, N101);
nand NAND4 (N1334, N1321, N714, N1094, N700);
or OR4 (N1335, N1301, N568, N486, N398);
not NOT1 (N1336, N1330);
buf BUF1 (N1337, N1329);
nand NAND2 (N1338, N1336, N566);
xor XOR2 (N1339, N1337, N1114);
xor XOR2 (N1340, N1323, N624);
nor NOR3 (N1341, N1340, N878, N972);
or OR3 (N1342, N1334, N410, N152);
and AND3 (N1343, N1341, N725, N494);
nor NOR4 (N1344, N1312, N1145, N937, N624);
xor XOR2 (N1345, N1333, N478);
buf BUF1 (N1346, N1343);
and AND4 (N1347, N1345, N1187, N17, N742);
nand NAND3 (N1348, N1316, N348, N156);
nand NAND3 (N1349, N1338, N485, N987);
buf BUF1 (N1350, N1344);
nor NOR2 (N1351, N1332, N585);
and AND3 (N1352, N1339, N327, N672);
nand NAND3 (N1353, N1351, N690, N957);
buf BUF1 (N1354, N1324);
or OR3 (N1355, N1335, N605, N558);
or OR2 (N1356, N1350, N856);
buf BUF1 (N1357, N1346);
buf BUF1 (N1358, N1348);
nor NOR4 (N1359, N1353, N94, N975, N658);
xor XOR2 (N1360, N1342, N548);
nand NAND2 (N1361, N1358, N470);
or OR3 (N1362, N1359, N54, N424);
xor XOR2 (N1363, N1357, N911);
and AND3 (N1364, N1349, N657, N1213);
xor XOR2 (N1365, N1362, N953);
and AND3 (N1366, N1347, N41, N1202);
nor NOR3 (N1367, N1352, N513, N357);
nand NAND2 (N1368, N1365, N1359);
xor XOR2 (N1369, N1354, N1301);
nor NOR3 (N1370, N1356, N573, N597);
or OR2 (N1371, N1369, N336);
nand NAND2 (N1372, N1364, N882);
xor XOR2 (N1373, N1368, N1192);
nor NOR3 (N1374, N1371, N461, N1204);
and AND3 (N1375, N1360, N552, N472);
buf BUF1 (N1376, N1361);
not NOT1 (N1377, N1373);
buf BUF1 (N1378, N1376);
or OR2 (N1379, N1378, N1140);
nand NAND2 (N1380, N1372, N115);
not NOT1 (N1381, N1355);
nor NOR3 (N1382, N1370, N164, N682);
buf BUF1 (N1383, N1367);
buf BUF1 (N1384, N1374);
and AND3 (N1385, N1377, N1129, N725);
nor NOR3 (N1386, N1375, N190, N1011);
or OR3 (N1387, N1366, N1208, N807);
not NOT1 (N1388, N1384);
or OR3 (N1389, N1386, N1165, N109);
or OR3 (N1390, N1380, N639, N75);
nor NOR3 (N1391, N1387, N349, N891);
nor NOR3 (N1392, N1363, N578, N985);
or OR4 (N1393, N1382, N470, N424, N307);
not NOT1 (N1394, N1379);
and AND4 (N1395, N1391, N37, N337, N920);
nor NOR2 (N1396, N1381, N109);
xor XOR2 (N1397, N1388, N151);
xor XOR2 (N1398, N1396, N325);
and AND4 (N1399, N1390, N525, N1290, N34);
xor XOR2 (N1400, N1389, N33);
nor NOR4 (N1401, N1393, N631, N361, N310);
or OR2 (N1402, N1400, N1053);
nor NOR4 (N1403, N1394, N1139, N233, N813);
buf BUF1 (N1404, N1398);
and AND3 (N1405, N1383, N63, N1203);
not NOT1 (N1406, N1385);
not NOT1 (N1407, N1401);
buf BUF1 (N1408, N1406);
nor NOR2 (N1409, N1397, N1345);
or OR3 (N1410, N1407, N1099, N1275);
xor XOR2 (N1411, N1392, N758);
not NOT1 (N1412, N1403);
nand NAND2 (N1413, N1405, N1008);
buf BUF1 (N1414, N1412);
not NOT1 (N1415, N1410);
buf BUF1 (N1416, N1399);
not NOT1 (N1417, N1415);
buf BUF1 (N1418, N1411);
or OR2 (N1419, N1417, N769);
or OR2 (N1420, N1402, N1352);
and AND3 (N1421, N1408, N1351, N1213);
not NOT1 (N1422, N1418);
nor NOR4 (N1423, N1419, N252, N345, N614);
nand NAND2 (N1424, N1420, N974);
xor XOR2 (N1425, N1395, N695);
and AND4 (N1426, N1414, N860, N876, N1202);
or OR4 (N1427, N1423, N1169, N410, N686);
not NOT1 (N1428, N1426);
xor XOR2 (N1429, N1409, N1123);
buf BUF1 (N1430, N1427);
xor XOR2 (N1431, N1430, N424);
and AND3 (N1432, N1429, N358, N116);
and AND3 (N1433, N1413, N174, N760);
nor NOR4 (N1434, N1416, N1146, N1018, N76);
nor NOR4 (N1435, N1431, N200, N673, N287);
buf BUF1 (N1436, N1434);
xor XOR2 (N1437, N1421, N678);
nand NAND3 (N1438, N1428, N1170, N312);
xor XOR2 (N1439, N1425, N1047);
not NOT1 (N1440, N1438);
not NOT1 (N1441, N1422);
nand NAND4 (N1442, N1439, N1055, N294, N172);
xor XOR2 (N1443, N1432, N655);
and AND3 (N1444, N1443, N664, N1177);
or OR3 (N1445, N1424, N373, N1287);
not NOT1 (N1446, N1442);
xor XOR2 (N1447, N1404, N487);
xor XOR2 (N1448, N1436, N1292);
or OR3 (N1449, N1435, N1295, N183);
or OR4 (N1450, N1440, N1023, N856, N23);
buf BUF1 (N1451, N1447);
and AND3 (N1452, N1444, N1050, N30);
or OR3 (N1453, N1448, N1092, N341);
nand NAND4 (N1454, N1451, N839, N868, N510);
buf BUF1 (N1455, N1445);
nand NAND2 (N1456, N1437, N624);
nor NOR3 (N1457, N1452, N543, N9);
not NOT1 (N1458, N1449);
xor XOR2 (N1459, N1457, N44);
not NOT1 (N1460, N1446);
and AND2 (N1461, N1433, N1378);
nand NAND2 (N1462, N1461, N745);
buf BUF1 (N1463, N1450);
and AND3 (N1464, N1454, N166, N1337);
nor NOR2 (N1465, N1441, N1460);
not NOT1 (N1466, N962);
or OR4 (N1467, N1465, N128, N1408, N251);
buf BUF1 (N1468, N1463);
nand NAND3 (N1469, N1466, N995, N767);
and AND3 (N1470, N1468, N1142, N1400);
and AND3 (N1471, N1470, N471, N1099);
and AND4 (N1472, N1456, N1175, N1162, N1145);
xor XOR2 (N1473, N1458, N1057);
and AND3 (N1474, N1467, N276, N307);
not NOT1 (N1475, N1473);
not NOT1 (N1476, N1464);
buf BUF1 (N1477, N1474);
not NOT1 (N1478, N1453);
xor XOR2 (N1479, N1478, N301);
xor XOR2 (N1480, N1477, N224);
xor XOR2 (N1481, N1475, N479);
nand NAND3 (N1482, N1471, N800, N1053);
nor NOR3 (N1483, N1462, N560, N341);
and AND4 (N1484, N1480, N573, N472, N218);
not NOT1 (N1485, N1455);
nor NOR4 (N1486, N1476, N1005, N927, N889);
buf BUF1 (N1487, N1482);
nand NAND4 (N1488, N1459, N915, N967, N1361);
xor XOR2 (N1489, N1486, N1467);
xor XOR2 (N1490, N1484, N1077);
and AND4 (N1491, N1479, N89, N1291, N240);
not NOT1 (N1492, N1483);
and AND3 (N1493, N1488, N1403, N648);
buf BUF1 (N1494, N1472);
nor NOR4 (N1495, N1494, N728, N607, N1289);
or OR2 (N1496, N1495, N25);
and AND4 (N1497, N1490, N1387, N71, N241);
nand NAND4 (N1498, N1485, N1024, N886, N489);
or OR2 (N1499, N1497, N825);
and AND2 (N1500, N1493, N68);
nor NOR2 (N1501, N1496, N529);
nor NOR4 (N1502, N1492, N628, N262, N1081);
buf BUF1 (N1503, N1501);
nor NOR2 (N1504, N1498, N1466);
nor NOR4 (N1505, N1489, N1202, N1021, N1294);
and AND4 (N1506, N1491, N550, N219, N212);
and AND4 (N1507, N1504, N174, N208, N899);
nand NAND4 (N1508, N1499, N641, N887, N164);
xor XOR2 (N1509, N1505, N108);
and AND3 (N1510, N1503, N1232, N708);
and AND4 (N1511, N1509, N646, N1140, N356);
not NOT1 (N1512, N1500);
nand NAND3 (N1513, N1481, N1188, N1305);
nand NAND2 (N1514, N1508, N978);
xor XOR2 (N1515, N1510, N275);
buf BUF1 (N1516, N1514);
buf BUF1 (N1517, N1516);
xor XOR2 (N1518, N1512, N661);
buf BUF1 (N1519, N1487);
xor XOR2 (N1520, N1507, N974);
xor XOR2 (N1521, N1506, N298);
not NOT1 (N1522, N1520);
not NOT1 (N1523, N1502);
not NOT1 (N1524, N1513);
nor NOR3 (N1525, N1521, N1217, N1202);
or OR4 (N1526, N1517, N550, N214, N1394);
or OR4 (N1527, N1511, N421, N1045, N1327);
nor NOR4 (N1528, N1469, N697, N356, N1393);
and AND2 (N1529, N1528, N143);
or OR3 (N1530, N1524, N795, N592);
buf BUF1 (N1531, N1519);
xor XOR2 (N1532, N1526, N815);
and AND2 (N1533, N1522, N1346);
nor NOR4 (N1534, N1523, N919, N1477, N621);
xor XOR2 (N1535, N1525, N1259);
nand NAND2 (N1536, N1515, N181);
not NOT1 (N1537, N1529);
or OR3 (N1538, N1536, N855, N40);
nand NAND2 (N1539, N1530, N837);
buf BUF1 (N1540, N1537);
xor XOR2 (N1541, N1535, N398);
buf BUF1 (N1542, N1518);
buf BUF1 (N1543, N1533);
not NOT1 (N1544, N1531);
nor NOR3 (N1545, N1542, N1344, N592);
not NOT1 (N1546, N1544);
nand NAND3 (N1547, N1543, N1408, N757);
not NOT1 (N1548, N1540);
nand NAND3 (N1549, N1538, N539, N193);
nor NOR3 (N1550, N1549, N1198, N1303);
not NOT1 (N1551, N1547);
or OR3 (N1552, N1548, N824, N298);
buf BUF1 (N1553, N1552);
nor NOR3 (N1554, N1553, N177, N877);
nor NOR3 (N1555, N1539, N457, N1436);
buf BUF1 (N1556, N1545);
or OR3 (N1557, N1551, N541, N1008);
not NOT1 (N1558, N1534);
buf BUF1 (N1559, N1557);
xor XOR2 (N1560, N1550, N457);
nor NOR4 (N1561, N1560, N1423, N1341, N863);
nor NOR4 (N1562, N1532, N1482, N1385, N416);
and AND2 (N1563, N1559, N1016);
and AND4 (N1564, N1554, N102, N9, N374);
nand NAND2 (N1565, N1561, N912);
xor XOR2 (N1566, N1565, N233);
not NOT1 (N1567, N1564);
xor XOR2 (N1568, N1567, N405);
nand NAND4 (N1569, N1563, N273, N433, N470);
or OR3 (N1570, N1566, N323, N416);
not NOT1 (N1571, N1558);
xor XOR2 (N1572, N1546, N82);
and AND2 (N1573, N1541, N954);
xor XOR2 (N1574, N1572, N205);
xor XOR2 (N1575, N1569, N612);
nor NOR2 (N1576, N1527, N351);
or OR2 (N1577, N1556, N1465);
or OR4 (N1578, N1562, N219, N447, N783);
nor NOR4 (N1579, N1555, N506, N703, N1495);
and AND4 (N1580, N1573, N1145, N618, N250);
nand NAND4 (N1581, N1578, N904, N1184, N1483);
not NOT1 (N1582, N1570);
nand NAND3 (N1583, N1581, N437, N1089);
or OR3 (N1584, N1574, N812, N1054);
buf BUF1 (N1585, N1580);
and AND2 (N1586, N1575, N779);
and AND4 (N1587, N1583, N522, N1495, N1039);
or OR3 (N1588, N1571, N590, N1038);
and AND2 (N1589, N1588, N324);
nand NAND3 (N1590, N1584, N318, N337);
and AND2 (N1591, N1587, N1036);
not NOT1 (N1592, N1585);
xor XOR2 (N1593, N1568, N74);
not NOT1 (N1594, N1589);
and AND4 (N1595, N1577, N413, N313, N173);
nor NOR3 (N1596, N1590, N41, N82);
xor XOR2 (N1597, N1586, N1280);
nand NAND4 (N1598, N1595, N871, N1150, N644);
nor NOR4 (N1599, N1582, N1534, N152, N1023);
xor XOR2 (N1600, N1576, N1160);
buf BUF1 (N1601, N1594);
nor NOR4 (N1602, N1600, N1104, N1234, N28);
not NOT1 (N1603, N1597);
nor NOR3 (N1604, N1579, N983, N574);
buf BUF1 (N1605, N1598);
nand NAND2 (N1606, N1593, N223);
not NOT1 (N1607, N1602);
and AND4 (N1608, N1605, N1044, N199, N1183);
nor NOR4 (N1609, N1604, N504, N1462, N941);
buf BUF1 (N1610, N1607);
xor XOR2 (N1611, N1606, N1199);
not NOT1 (N1612, N1591);
and AND2 (N1613, N1612, N1529);
nand NAND4 (N1614, N1601, N940, N15, N619);
and AND3 (N1615, N1609, N425, N83);
not NOT1 (N1616, N1613);
nand NAND2 (N1617, N1592, N89);
or OR3 (N1618, N1611, N292, N856);
nor NOR2 (N1619, N1608, N611);
nand NAND2 (N1620, N1610, N1147);
nor NOR2 (N1621, N1615, N394);
or OR2 (N1622, N1619, N937);
nor NOR4 (N1623, N1616, N1089, N1080, N107);
or OR2 (N1624, N1620, N1145);
xor XOR2 (N1625, N1623, N1116);
xor XOR2 (N1626, N1618, N1293);
and AND4 (N1627, N1622, N1039, N1497, N20);
xor XOR2 (N1628, N1596, N758);
not NOT1 (N1629, N1626);
buf BUF1 (N1630, N1603);
and AND4 (N1631, N1624, N326, N501, N774);
or OR3 (N1632, N1625, N987, N1568);
nor NOR3 (N1633, N1614, N479, N1549);
nor NOR3 (N1634, N1621, N144, N282);
or OR4 (N1635, N1628, N482, N1588, N234);
and AND4 (N1636, N1634, N1138, N458, N414);
not NOT1 (N1637, N1617);
xor XOR2 (N1638, N1636, N1217);
or OR4 (N1639, N1599, N1380, N735, N93);
xor XOR2 (N1640, N1630, N921);
buf BUF1 (N1641, N1632);
not NOT1 (N1642, N1641);
nand NAND3 (N1643, N1642, N695, N476);
nor NOR3 (N1644, N1640, N1619, N1109);
xor XOR2 (N1645, N1639, N1231);
or OR2 (N1646, N1643, N169);
buf BUF1 (N1647, N1633);
or OR3 (N1648, N1647, N1428, N1226);
not NOT1 (N1649, N1629);
buf BUF1 (N1650, N1648);
nor NOR3 (N1651, N1650, N1023, N43);
xor XOR2 (N1652, N1627, N965);
nor NOR3 (N1653, N1638, N721, N875);
nor NOR2 (N1654, N1637, N1546);
and AND2 (N1655, N1644, N1543);
nand NAND4 (N1656, N1646, N348, N1488, N1405);
xor XOR2 (N1657, N1635, N223);
and AND2 (N1658, N1649, N1412);
xor XOR2 (N1659, N1631, N896);
buf BUF1 (N1660, N1658);
xor XOR2 (N1661, N1655, N794);
and AND3 (N1662, N1661, N107, N912);
and AND2 (N1663, N1659, N1497);
nand NAND4 (N1664, N1662, N405, N508, N1337);
nor NOR4 (N1665, N1656, N472, N1282, N1139);
xor XOR2 (N1666, N1657, N288);
and AND3 (N1667, N1665, N1379, N809);
xor XOR2 (N1668, N1660, N1376);
not NOT1 (N1669, N1668);
not NOT1 (N1670, N1664);
nor NOR3 (N1671, N1645, N143, N1551);
xor XOR2 (N1672, N1651, N175);
nor NOR4 (N1673, N1653, N358, N1412, N1138);
not NOT1 (N1674, N1652);
nand NAND3 (N1675, N1666, N1215, N1314);
not NOT1 (N1676, N1673);
buf BUF1 (N1677, N1672);
buf BUF1 (N1678, N1669);
buf BUF1 (N1679, N1654);
xor XOR2 (N1680, N1674, N1416);
not NOT1 (N1681, N1670);
xor XOR2 (N1682, N1675, N1099);
nand NAND4 (N1683, N1680, N871, N27, N189);
xor XOR2 (N1684, N1676, N220);
nor NOR2 (N1685, N1663, N337);
nand NAND2 (N1686, N1677, N1272);
buf BUF1 (N1687, N1679);
not NOT1 (N1688, N1683);
not NOT1 (N1689, N1686);
nand NAND2 (N1690, N1684, N1397);
and AND2 (N1691, N1667, N251);
and AND3 (N1692, N1678, N1640, N329);
nand NAND3 (N1693, N1685, N1330, N1040);
or OR3 (N1694, N1693, N1564, N1145);
or OR3 (N1695, N1682, N987, N221);
not NOT1 (N1696, N1690);
and AND4 (N1697, N1692, N1235, N760, N1573);
and AND2 (N1698, N1688, N305);
or OR2 (N1699, N1696, N1325);
or OR4 (N1700, N1694, N222, N890, N1039);
nor NOR3 (N1701, N1695, N908, N611);
nand NAND4 (N1702, N1687, N804, N408, N97);
and AND2 (N1703, N1702, N176);
not NOT1 (N1704, N1703);
nand NAND3 (N1705, N1701, N461, N1294);
not NOT1 (N1706, N1697);
xor XOR2 (N1707, N1689, N1251);
nor NOR2 (N1708, N1691, N1492);
and AND3 (N1709, N1700, N815, N1316);
or OR4 (N1710, N1707, N84, N560, N443);
or OR4 (N1711, N1708, N280, N1142, N1607);
xor XOR2 (N1712, N1705, N861);
not NOT1 (N1713, N1712);
not NOT1 (N1714, N1698);
nor NOR4 (N1715, N1713, N175, N841, N1040);
nand NAND3 (N1716, N1714, N537, N301);
or OR3 (N1717, N1711, N769, N688);
nor NOR3 (N1718, N1710, N1284, N914);
nor NOR3 (N1719, N1715, N41, N679);
nor NOR2 (N1720, N1706, N832);
and AND2 (N1721, N1717, N1050);
or OR4 (N1722, N1699, N1304, N751, N1425);
xor XOR2 (N1723, N1671, N1060);
nor NOR2 (N1724, N1721, N228);
nor NOR4 (N1725, N1704, N1039, N567, N1173);
and AND3 (N1726, N1722, N1260, N1405);
or OR4 (N1727, N1726, N727, N1396, N1430);
nor NOR3 (N1728, N1723, N1085, N1691);
buf BUF1 (N1729, N1716);
buf BUF1 (N1730, N1719);
or OR2 (N1731, N1727, N548);
nand NAND2 (N1732, N1718, N544);
nand NAND3 (N1733, N1725, N427, N453);
nor NOR4 (N1734, N1728, N1032, N711, N644);
or OR2 (N1735, N1729, N186);
nand NAND3 (N1736, N1732, N838, N1023);
and AND2 (N1737, N1681, N550);
not NOT1 (N1738, N1731);
xor XOR2 (N1739, N1733, N1022);
buf BUF1 (N1740, N1736);
or OR4 (N1741, N1737, N556, N1242, N1047);
nor NOR3 (N1742, N1724, N252, N1417);
not NOT1 (N1743, N1709);
buf BUF1 (N1744, N1740);
or OR4 (N1745, N1744, N1284, N60, N192);
nor NOR3 (N1746, N1734, N39, N846);
and AND4 (N1747, N1742, N1021, N1514, N303);
nor NOR3 (N1748, N1746, N1175, N1019);
and AND4 (N1749, N1720, N1563, N78, N106);
not NOT1 (N1750, N1741);
xor XOR2 (N1751, N1730, N314);
xor XOR2 (N1752, N1748, N1572);
xor XOR2 (N1753, N1735, N131);
and AND3 (N1754, N1747, N482, N610);
not NOT1 (N1755, N1753);
or OR3 (N1756, N1750, N1112, N912);
and AND2 (N1757, N1738, N1544);
nand NAND3 (N1758, N1743, N980, N217);
nand NAND2 (N1759, N1754, N574);
and AND3 (N1760, N1749, N596, N487);
and AND2 (N1761, N1757, N1057);
or OR4 (N1762, N1761, N1434, N479, N1495);
or OR2 (N1763, N1751, N376);
nor NOR4 (N1764, N1763, N1403, N462, N1547);
buf BUF1 (N1765, N1752);
or OR2 (N1766, N1764, N506);
nor NOR4 (N1767, N1765, N474, N1046, N1694);
not NOT1 (N1768, N1758);
buf BUF1 (N1769, N1755);
nand NAND3 (N1770, N1756, N367, N79);
xor XOR2 (N1771, N1768, N760);
nand NAND3 (N1772, N1767, N754, N1711);
and AND2 (N1773, N1759, N1360);
nand NAND3 (N1774, N1772, N198, N375);
buf BUF1 (N1775, N1762);
or OR3 (N1776, N1739, N610, N1167);
buf BUF1 (N1777, N1774);
or OR4 (N1778, N1775, N1032, N1759, N860);
or OR2 (N1779, N1745, N1380);
and AND3 (N1780, N1771, N255, N484);
xor XOR2 (N1781, N1780, N1316);
nand NAND4 (N1782, N1778, N1141, N715, N1254);
not NOT1 (N1783, N1782);
buf BUF1 (N1784, N1769);
xor XOR2 (N1785, N1783, N67);
and AND2 (N1786, N1781, N741);
xor XOR2 (N1787, N1760, N841);
or OR2 (N1788, N1786, N546);
and AND4 (N1789, N1779, N347, N932, N114);
or OR4 (N1790, N1789, N382, N240, N1234);
nor NOR2 (N1791, N1773, N1744);
and AND2 (N1792, N1791, N1750);
and AND3 (N1793, N1770, N1683, N574);
not NOT1 (N1794, N1793);
not NOT1 (N1795, N1790);
nor NOR4 (N1796, N1784, N1747, N731, N734);
nand NAND4 (N1797, N1796, N501, N352, N794);
or OR4 (N1798, N1795, N678, N1600, N844);
not NOT1 (N1799, N1785);
xor XOR2 (N1800, N1797, N55);
nand NAND2 (N1801, N1777, N1722);
nand NAND2 (N1802, N1801, N285);
nand NAND2 (N1803, N1794, N1061);
or OR3 (N1804, N1800, N291, N1780);
and AND4 (N1805, N1788, N662, N1142, N913);
and AND2 (N1806, N1787, N1553);
and AND4 (N1807, N1802, N699, N616, N1511);
xor XOR2 (N1808, N1792, N103);
or OR4 (N1809, N1766, N415, N1209, N1372);
and AND2 (N1810, N1806, N260);
and AND2 (N1811, N1809, N1461);
or OR3 (N1812, N1808, N1075, N265);
buf BUF1 (N1813, N1811);
and AND2 (N1814, N1812, N44);
or OR3 (N1815, N1810, N721, N1149);
nand NAND4 (N1816, N1814, N103, N851, N951);
xor XOR2 (N1817, N1776, N653);
buf BUF1 (N1818, N1799);
xor XOR2 (N1819, N1817, N476);
xor XOR2 (N1820, N1813, N349);
or OR4 (N1821, N1819, N672, N37, N1454);
nand NAND3 (N1822, N1816, N1297, N1291);
nor NOR3 (N1823, N1807, N143, N642);
or OR3 (N1824, N1805, N1800, N484);
not NOT1 (N1825, N1815);
nand NAND4 (N1826, N1821, N1461, N1181, N967);
not NOT1 (N1827, N1824);
or OR4 (N1828, N1826, N518, N1336, N195);
nor NOR4 (N1829, N1825, N110, N1434, N314);
xor XOR2 (N1830, N1820, N547);
buf BUF1 (N1831, N1822);
and AND3 (N1832, N1831, N259, N1726);
nand NAND3 (N1833, N1823, N1107, N901);
not NOT1 (N1834, N1829);
not NOT1 (N1835, N1803);
and AND3 (N1836, N1833, N1485, N546);
and AND4 (N1837, N1835, N263, N1198, N470);
xor XOR2 (N1838, N1834, N491);
and AND2 (N1839, N1837, N110);
not NOT1 (N1840, N1827);
or OR2 (N1841, N1804, N1367);
nor NOR2 (N1842, N1839, N1323);
or OR3 (N1843, N1830, N1698, N393);
nor NOR4 (N1844, N1841, N63, N157, N1516);
not NOT1 (N1845, N1842);
or OR2 (N1846, N1845, N1364);
not NOT1 (N1847, N1843);
and AND3 (N1848, N1840, N1553, N602);
not NOT1 (N1849, N1836);
buf BUF1 (N1850, N1848);
nand NAND4 (N1851, N1828, N1069, N814, N1650);
nor NOR3 (N1852, N1850, N702, N1045);
nor NOR3 (N1853, N1849, N19, N1767);
not NOT1 (N1854, N1853);
and AND2 (N1855, N1846, N104);
or OR2 (N1856, N1798, N1594);
buf BUF1 (N1857, N1832);
and AND4 (N1858, N1844, N1185, N1049, N1199);
and AND4 (N1859, N1855, N1044, N1402, N1615);
nand NAND2 (N1860, N1851, N1628);
buf BUF1 (N1861, N1857);
buf BUF1 (N1862, N1861);
and AND3 (N1863, N1854, N191, N900);
and AND2 (N1864, N1862, N508);
buf BUF1 (N1865, N1864);
not NOT1 (N1866, N1856);
not NOT1 (N1867, N1847);
nor NOR4 (N1868, N1866, N843, N723, N496);
not NOT1 (N1869, N1858);
or OR4 (N1870, N1859, N682, N1308, N1582);
not NOT1 (N1871, N1838);
and AND3 (N1872, N1870, N1348, N1560);
or OR2 (N1873, N1869, N151);
or OR4 (N1874, N1865, N1198, N1712, N819);
or OR2 (N1875, N1818, N327);
xor XOR2 (N1876, N1873, N1055);
xor XOR2 (N1877, N1852, N1870);
buf BUF1 (N1878, N1877);
and AND3 (N1879, N1875, N566, N1400);
xor XOR2 (N1880, N1878, N1837);
not NOT1 (N1881, N1860);
nand NAND3 (N1882, N1868, N888, N537);
not NOT1 (N1883, N1867);
buf BUF1 (N1884, N1881);
or OR2 (N1885, N1871, N1705);
buf BUF1 (N1886, N1880);
buf BUF1 (N1887, N1885);
xor XOR2 (N1888, N1887, N1840);
not NOT1 (N1889, N1876);
and AND3 (N1890, N1886, N1470, N1438);
buf BUF1 (N1891, N1872);
not NOT1 (N1892, N1884);
and AND2 (N1893, N1883, N1606);
or OR4 (N1894, N1889, N1598, N2, N137);
nor NOR4 (N1895, N1892, N1586, N857, N1592);
xor XOR2 (N1896, N1879, N212);
nor NOR2 (N1897, N1888, N530);
buf BUF1 (N1898, N1891);
and AND3 (N1899, N1863, N1534, N1691);
xor XOR2 (N1900, N1899, N1281);
buf BUF1 (N1901, N1900);
or OR2 (N1902, N1895, N1672);
and AND4 (N1903, N1890, N1738, N1231, N851);
or OR4 (N1904, N1902, N1586, N1768, N1853);
and AND2 (N1905, N1882, N1731);
or OR3 (N1906, N1904, N1769, N878);
nor NOR4 (N1907, N1874, N212, N1246, N41);
buf BUF1 (N1908, N1901);
xor XOR2 (N1909, N1898, N1592);
nor NOR4 (N1910, N1909, N1195, N1222, N1273);
not NOT1 (N1911, N1905);
nand NAND4 (N1912, N1911, N70, N257, N1769);
and AND3 (N1913, N1908, N1406, N1227);
or OR2 (N1914, N1907, N986);
nor NOR2 (N1915, N1894, N1111);
or OR4 (N1916, N1910, N1152, N282, N1788);
and AND3 (N1917, N1893, N970, N1892);
nor NOR2 (N1918, N1903, N772);
and AND4 (N1919, N1913, N954, N310, N941);
nor NOR3 (N1920, N1918, N1904, N1069);
nand NAND3 (N1921, N1897, N978, N739);
xor XOR2 (N1922, N1914, N1736);
buf BUF1 (N1923, N1917);
buf BUF1 (N1924, N1923);
nor NOR3 (N1925, N1915, N568, N1183);
and AND3 (N1926, N1921, N455, N1074);
xor XOR2 (N1927, N1912, N1918);
nand NAND4 (N1928, N1920, N1320, N1396, N1637);
nor NOR2 (N1929, N1919, N1395);
or OR2 (N1930, N1922, N1174);
not NOT1 (N1931, N1925);
buf BUF1 (N1932, N1924);
not NOT1 (N1933, N1932);
buf BUF1 (N1934, N1926);
xor XOR2 (N1935, N1930, N514);
and AND3 (N1936, N1935, N804, N905);
nor NOR3 (N1937, N1916, N1913, N38);
or OR4 (N1938, N1937, N1594, N158, N677);
not NOT1 (N1939, N1936);
nor NOR3 (N1940, N1906, N1661, N322);
nor NOR3 (N1941, N1938, N663, N1359);
or OR2 (N1942, N1939, N934);
xor XOR2 (N1943, N1942, N1330);
or OR2 (N1944, N1927, N711);
nor NOR4 (N1945, N1933, N263, N1821, N1197);
buf BUF1 (N1946, N1943);
or OR4 (N1947, N1944, N1775, N634, N1628);
not NOT1 (N1948, N1931);
not NOT1 (N1949, N1928);
xor XOR2 (N1950, N1929, N236);
nor NOR3 (N1951, N1945, N1142, N1222);
nor NOR2 (N1952, N1949, N157);
xor XOR2 (N1953, N1948, N1916);
or OR2 (N1954, N1951, N1859);
not NOT1 (N1955, N1954);
nand NAND2 (N1956, N1947, N538);
buf BUF1 (N1957, N1950);
buf BUF1 (N1958, N1952);
nor NOR2 (N1959, N1941, N409);
nor NOR2 (N1960, N1896, N92);
and AND4 (N1961, N1957, N356, N956, N1616);
or OR2 (N1962, N1960, N683);
nor NOR2 (N1963, N1959, N173);
nor NOR2 (N1964, N1934, N348);
not NOT1 (N1965, N1964);
not NOT1 (N1966, N1963);
and AND2 (N1967, N1965, N273);
buf BUF1 (N1968, N1967);
and AND3 (N1969, N1962, N1226, N918);
buf BUF1 (N1970, N1958);
not NOT1 (N1971, N1970);
not NOT1 (N1972, N1940);
not NOT1 (N1973, N1969);
xor XOR2 (N1974, N1956, N841);
and AND3 (N1975, N1968, N708, N1278);
and AND2 (N1976, N1961, N345);
xor XOR2 (N1977, N1966, N585);
or OR4 (N1978, N1971, N1119, N1268, N1937);
and AND2 (N1979, N1976, N1634);
and AND2 (N1980, N1973, N673);
not NOT1 (N1981, N1946);
buf BUF1 (N1982, N1981);
not NOT1 (N1983, N1978);
not NOT1 (N1984, N1974);
buf BUF1 (N1985, N1983);
or OR2 (N1986, N1972, N1658);
or OR3 (N1987, N1984, N1561, N1580);
not NOT1 (N1988, N1987);
not NOT1 (N1989, N1985);
and AND3 (N1990, N1982, N743, N194);
nor NOR4 (N1991, N1975, N244, N338, N96);
xor XOR2 (N1992, N1979, N427);
or OR2 (N1993, N1989, N1540);
nor NOR3 (N1994, N1977, N27, N745);
nand NAND4 (N1995, N1953, N369, N1646, N984);
or OR3 (N1996, N1986, N1848, N1922);
buf BUF1 (N1997, N1990);
or OR2 (N1998, N1993, N1092);
or OR2 (N1999, N1994, N1523);
not NOT1 (N2000, N1996);
nand NAND4 (N2001, N1991, N884, N1754, N1567);
nand NAND3 (N2002, N1955, N210, N572);
or OR4 (N2003, N1997, N1706, N1976, N1743);
buf BUF1 (N2004, N2002);
nand NAND4 (N2005, N2000, N1172, N1889, N1244);
or OR2 (N2006, N1998, N969);
and AND3 (N2007, N2005, N800, N1511);
nand NAND3 (N2008, N2004, N591, N664);
nor NOR3 (N2009, N1995, N756, N875);
nand NAND4 (N2010, N1992, N1824, N1023, N1029);
nand NAND3 (N2011, N2003, N1335, N1888);
xor XOR2 (N2012, N2011, N386);
xor XOR2 (N2013, N1999, N367);
buf BUF1 (N2014, N2001);
buf BUF1 (N2015, N2013);
xor XOR2 (N2016, N2007, N870);
xor XOR2 (N2017, N2006, N128);
nand NAND3 (N2018, N1980, N1988, N1891);
nand NAND3 (N2019, N1199, N1747, N1712);
nor NOR4 (N2020, N2018, N1856, N1258, N1019);
or OR4 (N2021, N2019, N1865, N660, N265);
not NOT1 (N2022, N2021);
xor XOR2 (N2023, N2017, N1522);
or OR4 (N2024, N2020, N246, N140, N1431);
nor NOR2 (N2025, N2023, N99);
nand NAND3 (N2026, N2022, N1859, N1838);
and AND4 (N2027, N2014, N1781, N818, N1012);
nor NOR4 (N2028, N2024, N880, N1402, N1767);
and AND4 (N2029, N2008, N1915, N1840, N205);
and AND3 (N2030, N2009, N139, N533);
or OR3 (N2031, N2029, N1156, N877);
nor NOR2 (N2032, N2010, N205);
xor XOR2 (N2033, N2031, N1532);
not NOT1 (N2034, N2012);
xor XOR2 (N2035, N2026, N280);
xor XOR2 (N2036, N2032, N547);
buf BUF1 (N2037, N2027);
buf BUF1 (N2038, N2035);
and AND2 (N2039, N2037, N164);
and AND4 (N2040, N2015, N143, N482, N601);
buf BUF1 (N2041, N2038);
or OR2 (N2042, N2028, N553);
or OR2 (N2043, N2040, N404);
and AND4 (N2044, N2042, N302, N146, N1117);
not NOT1 (N2045, N2025);
and AND4 (N2046, N2045, N875, N479, N1229);
buf BUF1 (N2047, N2043);
xor XOR2 (N2048, N2044, N646);
buf BUF1 (N2049, N2041);
xor XOR2 (N2050, N2034, N263);
xor XOR2 (N2051, N2016, N1930);
buf BUF1 (N2052, N2051);
buf BUF1 (N2053, N2047);
buf BUF1 (N2054, N2036);
not NOT1 (N2055, N2033);
xor XOR2 (N2056, N2046, N1630);
or OR3 (N2057, N2030, N1054, N458);
nand NAND2 (N2058, N2039, N426);
and AND3 (N2059, N2056, N1574, N1554);
buf BUF1 (N2060, N2052);
not NOT1 (N2061, N2060);
xor XOR2 (N2062, N2061, N836);
buf BUF1 (N2063, N2053);
xor XOR2 (N2064, N2058, N1573);
nand NAND3 (N2065, N2055, N712, N1505);
nand NAND4 (N2066, N2054, N469, N1655, N764);
xor XOR2 (N2067, N2059, N1206);
buf BUF1 (N2068, N2062);
nor NOR2 (N2069, N2066, N796);
xor XOR2 (N2070, N2049, N1218);
not NOT1 (N2071, N2067);
not NOT1 (N2072, N2069);
not NOT1 (N2073, N2071);
or OR4 (N2074, N2070, N1785, N1683, N1999);
nor NOR4 (N2075, N2068, N1437, N571, N903);
and AND4 (N2076, N2075, N1839, N1008, N1874);
nand NAND4 (N2077, N2048, N1668, N1952, N869);
xor XOR2 (N2078, N2057, N1931);
nand NAND3 (N2079, N2077, N817, N296);
or OR3 (N2080, N2064, N1668, N826);
and AND3 (N2081, N2076, N957, N1478);
or OR3 (N2082, N2081, N1924, N516);
nor NOR2 (N2083, N2073, N657);
buf BUF1 (N2084, N2050);
not NOT1 (N2085, N2072);
or OR4 (N2086, N2080, N1549, N119, N1034);
nand NAND3 (N2087, N2084, N177, N1321);
buf BUF1 (N2088, N2078);
xor XOR2 (N2089, N2063, N1743);
or OR3 (N2090, N2083, N493, N260);
nand NAND3 (N2091, N2089, N120, N301);
nor NOR2 (N2092, N2088, N1609);
nand NAND3 (N2093, N2090, N1690, N1559);
not NOT1 (N2094, N2092);
xor XOR2 (N2095, N2065, N117);
nor NOR3 (N2096, N2095, N146, N1750);
not NOT1 (N2097, N2079);
and AND4 (N2098, N2096, N1065, N50, N1497);
xor XOR2 (N2099, N2093, N1483);
and AND3 (N2100, N2098, N1743, N900);
or OR2 (N2101, N2074, N1);
nor NOR4 (N2102, N2086, N1764, N401, N1716);
or OR4 (N2103, N2099, N1409, N514, N869);
buf BUF1 (N2104, N2100);
and AND3 (N2105, N2082, N989, N279);
not NOT1 (N2106, N2094);
nor NOR4 (N2107, N2101, N1956, N634, N1121);
not NOT1 (N2108, N2106);
buf BUF1 (N2109, N2087);
buf BUF1 (N2110, N2097);
nor NOR4 (N2111, N2103, N1497, N858, N726);
xor XOR2 (N2112, N2102, N263);
buf BUF1 (N2113, N2110);
xor XOR2 (N2114, N2107, N2071);
not NOT1 (N2115, N2109);
xor XOR2 (N2116, N2091, N484);
buf BUF1 (N2117, N2115);
and AND2 (N2118, N2111, N854);
and AND2 (N2119, N2114, N435);
nand NAND2 (N2120, N2112, N1365);
and AND2 (N2121, N2116, N177);
or OR2 (N2122, N2105, N992);
or OR3 (N2123, N2121, N947, N1618);
nor NOR4 (N2124, N2120, N2025, N1841, N992);
and AND2 (N2125, N2113, N1082);
nand NAND4 (N2126, N2122, N124, N301, N139);
xor XOR2 (N2127, N2119, N261);
or OR3 (N2128, N2085, N1204, N573);
buf BUF1 (N2129, N2117);
nand NAND4 (N2130, N2125, N1279, N1474, N1909);
xor XOR2 (N2131, N2124, N1989);
nand NAND3 (N2132, N2130, N1872, N1794);
nor NOR2 (N2133, N2118, N1776);
buf BUF1 (N2134, N2126);
or OR4 (N2135, N2134, N544, N1598, N1371);
buf BUF1 (N2136, N2131);
and AND3 (N2137, N2127, N932, N394);
or OR4 (N2138, N2133, N546, N1634, N2029);
nand NAND3 (N2139, N2123, N213, N1367);
not NOT1 (N2140, N2138);
not NOT1 (N2141, N2135);
not NOT1 (N2142, N2136);
not NOT1 (N2143, N2132);
not NOT1 (N2144, N2140);
buf BUF1 (N2145, N2142);
or OR2 (N2146, N2128, N1633);
nand NAND2 (N2147, N2104, N1865);
not NOT1 (N2148, N2108);
buf BUF1 (N2149, N2147);
buf BUF1 (N2150, N2137);
not NOT1 (N2151, N2148);
or OR3 (N2152, N2139, N269, N1349);
not NOT1 (N2153, N2150);
nor NOR4 (N2154, N2129, N401, N1089, N956);
and AND3 (N2155, N2144, N124, N232);
nand NAND2 (N2156, N2141, N363);
nor NOR2 (N2157, N2143, N1958);
nand NAND2 (N2158, N2153, N800);
and AND3 (N2159, N2155, N2104, N1804);
and AND2 (N2160, N2145, N1320);
not NOT1 (N2161, N2149);
buf BUF1 (N2162, N2151);
buf BUF1 (N2163, N2159);
or OR2 (N2164, N2154, N540);
xor XOR2 (N2165, N2161, N511);
xor XOR2 (N2166, N2146, N724);
not NOT1 (N2167, N2165);
not NOT1 (N2168, N2158);
not NOT1 (N2169, N2164);
not NOT1 (N2170, N2169);
xor XOR2 (N2171, N2168, N1925);
xor XOR2 (N2172, N2152, N600);
not NOT1 (N2173, N2166);
not NOT1 (N2174, N2157);
nand NAND3 (N2175, N2167, N21, N2016);
buf BUF1 (N2176, N2173);
not NOT1 (N2177, N2160);
or OR4 (N2178, N2170, N2046, N1793, N1635);
nand NAND2 (N2179, N2163, N528);
nand NAND3 (N2180, N2179, N779, N1053);
nand NAND4 (N2181, N2176, N1262, N169, N247);
nand NAND3 (N2182, N2181, N1871, N1501);
or OR2 (N2183, N2172, N619);
or OR2 (N2184, N2156, N1398);
nand NAND2 (N2185, N2175, N2035);
xor XOR2 (N2186, N2180, N396);
xor XOR2 (N2187, N2184, N545);
buf BUF1 (N2188, N2186);
nor NOR3 (N2189, N2187, N810, N1528);
not NOT1 (N2190, N2183);
xor XOR2 (N2191, N2182, N1274);
and AND4 (N2192, N2177, N1373, N692, N1536);
nor NOR2 (N2193, N2178, N1932);
and AND2 (N2194, N2193, N1419);
not NOT1 (N2195, N2192);
buf BUF1 (N2196, N2191);
not NOT1 (N2197, N2188);
nor NOR4 (N2198, N2196, N1728, N1271, N1759);
nor NOR2 (N2199, N2194, N927);
buf BUF1 (N2200, N2197);
and AND4 (N2201, N2162, N996, N190, N663);
not NOT1 (N2202, N2190);
or OR2 (N2203, N2185, N404);
nand NAND3 (N2204, N2200, N1284, N524);
not NOT1 (N2205, N2199);
xor XOR2 (N2206, N2202, N130);
buf BUF1 (N2207, N2205);
nor NOR4 (N2208, N2174, N727, N502, N1705);
not NOT1 (N2209, N2203);
not NOT1 (N2210, N2207);
nand NAND4 (N2211, N2206, N1023, N697, N1594);
nor NOR4 (N2212, N2209, N1753, N1082, N426);
nor NOR2 (N2213, N2189, N653);
and AND2 (N2214, N2204, N1150);
not NOT1 (N2215, N2195);
or OR3 (N2216, N2201, N649, N253);
or OR3 (N2217, N2213, N1308, N1353);
not NOT1 (N2218, N2215);
xor XOR2 (N2219, N2217, N1919);
xor XOR2 (N2220, N2216, N1904);
xor XOR2 (N2221, N2220, N886);
buf BUF1 (N2222, N2221);
not NOT1 (N2223, N2214);
and AND3 (N2224, N2212, N1062, N2205);
xor XOR2 (N2225, N2198, N75);
nand NAND2 (N2226, N2210, N657);
nand NAND3 (N2227, N2208, N1846, N705);
xor XOR2 (N2228, N2224, N1679);
nand NAND3 (N2229, N2225, N1053, N2034);
xor XOR2 (N2230, N2229, N1521);
nand NAND4 (N2231, N2219, N1023, N532, N550);
not NOT1 (N2232, N2211);
nand NAND3 (N2233, N2230, N2021, N477);
not NOT1 (N2234, N2227);
buf BUF1 (N2235, N2171);
not NOT1 (N2236, N2222);
buf BUF1 (N2237, N2233);
buf BUF1 (N2238, N2236);
xor XOR2 (N2239, N2218, N416);
not NOT1 (N2240, N2235);
buf BUF1 (N2241, N2228);
nor NOR3 (N2242, N2240, N1353, N2015);
and AND3 (N2243, N2231, N2157, N648);
and AND3 (N2244, N2223, N1728, N2194);
not NOT1 (N2245, N2234);
or OR4 (N2246, N2232, N84, N1299, N2023);
and AND4 (N2247, N2237, N523, N1200, N1801);
or OR3 (N2248, N2238, N654, N2141);
nand NAND4 (N2249, N2239, N691, N1751, N790);
or OR4 (N2250, N2244, N1649, N1185, N1546);
not NOT1 (N2251, N2246);
nor NOR3 (N2252, N2249, N1922, N1853);
or OR4 (N2253, N2242, N1965, N1722, N456);
nor NOR3 (N2254, N2241, N1259, N1857);
not NOT1 (N2255, N2253);
nand NAND2 (N2256, N2252, N1891);
not NOT1 (N2257, N2247);
nor NOR4 (N2258, N2245, N606, N443, N1);
and AND2 (N2259, N2257, N103);
nor NOR3 (N2260, N2243, N686, N20);
nor NOR2 (N2261, N2258, N748);
nor NOR2 (N2262, N2254, N638);
and AND3 (N2263, N2262, N1575, N774);
nand NAND4 (N2264, N2248, N538, N1270, N70);
xor XOR2 (N2265, N2260, N2067);
nor NOR2 (N2266, N2264, N228);
nand NAND4 (N2267, N2255, N1771, N1728, N1193);
not NOT1 (N2268, N2263);
xor XOR2 (N2269, N2259, N746);
or OR3 (N2270, N2256, N646, N782);
not NOT1 (N2271, N2265);
nor NOR3 (N2272, N2268, N1991, N364);
or OR3 (N2273, N2270, N518, N1881);
xor XOR2 (N2274, N2266, N825);
nor NOR2 (N2275, N2272, N508);
buf BUF1 (N2276, N2269);
xor XOR2 (N2277, N2271, N1082);
nor NOR2 (N2278, N2261, N413);
not NOT1 (N2279, N2273);
nor NOR3 (N2280, N2275, N975, N2157);
not NOT1 (N2281, N2251);
nor NOR4 (N2282, N2250, N1244, N121, N27);
nand NAND2 (N2283, N2282, N2017);
or OR3 (N2284, N2278, N1135, N568);
nand NAND3 (N2285, N2284, N26, N1972);
not NOT1 (N2286, N2226);
not NOT1 (N2287, N2286);
and AND2 (N2288, N2276, N943);
buf BUF1 (N2289, N2281);
nor NOR4 (N2290, N2283, N908, N1380, N157);
not NOT1 (N2291, N2290);
xor XOR2 (N2292, N2289, N326);
and AND4 (N2293, N2274, N1617, N1566, N1360);
not NOT1 (N2294, N2267);
not NOT1 (N2295, N2287);
buf BUF1 (N2296, N2294);
and AND4 (N2297, N2279, N761, N1176, N23);
nand NAND4 (N2298, N2291, N1749, N1745, N1095);
nand NAND2 (N2299, N2296, N524);
nor NOR3 (N2300, N2288, N1408, N265);
nor NOR4 (N2301, N2299, N1731, N2150, N1343);
nand NAND2 (N2302, N2300, N1696);
xor XOR2 (N2303, N2277, N1825);
not NOT1 (N2304, N2297);
and AND4 (N2305, N2293, N822, N231, N2295);
buf BUF1 (N2306, N1426);
or OR4 (N2307, N2292, N24, N2210, N1896);
nor NOR2 (N2308, N2306, N1177);
or OR3 (N2309, N2301, N854, N1181);
nand NAND2 (N2310, N2303, N1867);
nand NAND2 (N2311, N2308, N2283);
nor NOR3 (N2312, N2280, N912, N2166);
xor XOR2 (N2313, N2310, N265);
xor XOR2 (N2314, N2312, N1712);
not NOT1 (N2315, N2314);
and AND2 (N2316, N2315, N928);
not NOT1 (N2317, N2304);
nor NOR3 (N2318, N2305, N836, N256);
nor NOR4 (N2319, N2307, N1664, N2205, N182);
or OR3 (N2320, N2311, N1794, N159);
xor XOR2 (N2321, N2320, N657);
and AND4 (N2322, N2316, N1186, N1220, N1958);
xor XOR2 (N2323, N2318, N954);
and AND2 (N2324, N2309, N1703);
or OR3 (N2325, N2321, N595, N159);
not NOT1 (N2326, N2323);
or OR2 (N2327, N2325, N239);
buf BUF1 (N2328, N2302);
and AND4 (N2329, N2319, N18, N492, N2266);
or OR3 (N2330, N2317, N199, N486);
and AND4 (N2331, N2329, N1144, N1828, N1517);
buf BUF1 (N2332, N2326);
and AND3 (N2333, N2332, N1275, N627);
and AND3 (N2334, N2328, N837, N1223);
xor XOR2 (N2335, N2327, N375);
and AND4 (N2336, N2324, N2187, N1665, N1635);
xor XOR2 (N2337, N2333, N1287);
xor XOR2 (N2338, N2334, N1612);
and AND4 (N2339, N2336, N301, N604, N382);
not NOT1 (N2340, N2322);
nor NOR2 (N2341, N2337, N1559);
or OR2 (N2342, N2338, N98);
not NOT1 (N2343, N2330);
and AND3 (N2344, N2331, N848, N1953);
xor XOR2 (N2345, N2335, N1269);
nand NAND3 (N2346, N2341, N1546, N598);
not NOT1 (N2347, N2345);
or OR3 (N2348, N2347, N2247, N413);
and AND4 (N2349, N2285, N1922, N931, N457);
buf BUF1 (N2350, N2346);
or OR3 (N2351, N2349, N1761, N833);
or OR4 (N2352, N2351, N1817, N19, N2037);
xor XOR2 (N2353, N2344, N1894);
or OR2 (N2354, N2350, N996);
or OR4 (N2355, N2353, N409, N443, N689);
or OR3 (N2356, N2354, N1225, N281);
and AND2 (N2357, N2313, N1614);
xor XOR2 (N2358, N2348, N428);
and AND4 (N2359, N2352, N1861, N422, N1835);
buf BUF1 (N2360, N2340);
and AND4 (N2361, N2357, N465, N482, N988);
or OR3 (N2362, N2359, N933, N217);
not NOT1 (N2363, N2361);
and AND2 (N2364, N2363, N1627);
nand NAND3 (N2365, N2342, N1433, N1262);
not NOT1 (N2366, N2343);
and AND3 (N2367, N2366, N1216, N114);
xor XOR2 (N2368, N2360, N1253);
or OR2 (N2369, N2367, N891);
xor XOR2 (N2370, N2355, N482);
and AND3 (N2371, N2369, N763, N637);
xor XOR2 (N2372, N2339, N1061);
or OR2 (N2373, N2298, N2213);
nor NOR4 (N2374, N2372, N1894, N1170, N1012);
nor NOR3 (N2375, N2374, N1049, N2094);
nand NAND2 (N2376, N2375, N1556);
buf BUF1 (N2377, N2373);
nand NAND3 (N2378, N2358, N48, N441);
or OR4 (N2379, N2364, N927, N1487, N1041);
and AND2 (N2380, N2377, N1682);
nand NAND4 (N2381, N2365, N1848, N332, N1107);
not NOT1 (N2382, N2381);
buf BUF1 (N2383, N2368);
xor XOR2 (N2384, N2356, N1140);
xor XOR2 (N2385, N2376, N2198);
nand NAND2 (N2386, N2378, N602);
not NOT1 (N2387, N2380);
nor NOR4 (N2388, N2385, N1272, N2057, N2382);
not NOT1 (N2389, N1508);
nand NAND3 (N2390, N2386, N557, N429);
nand NAND4 (N2391, N2362, N2325, N113, N1946);
and AND2 (N2392, N2370, N1794);
xor XOR2 (N2393, N2388, N131);
xor XOR2 (N2394, N2393, N367);
and AND2 (N2395, N2384, N722);
buf BUF1 (N2396, N2379);
and AND3 (N2397, N2371, N763, N530);
or OR2 (N2398, N2397, N1042);
xor XOR2 (N2399, N2392, N1285);
buf BUF1 (N2400, N2390);
nor NOR3 (N2401, N2391, N724, N2136);
and AND3 (N2402, N2387, N2122, N1776);
xor XOR2 (N2403, N2398, N1524);
nor NOR2 (N2404, N2394, N1374);
not NOT1 (N2405, N2396);
not NOT1 (N2406, N2389);
or OR2 (N2407, N2403, N1190);
xor XOR2 (N2408, N2404, N1032);
buf BUF1 (N2409, N2402);
and AND3 (N2410, N2408, N205, N1232);
xor XOR2 (N2411, N2383, N484);
and AND3 (N2412, N2405, N1166, N1274);
xor XOR2 (N2413, N2411, N752);
nor NOR2 (N2414, N2400, N1176);
xor XOR2 (N2415, N2407, N93);
and AND3 (N2416, N2413, N2320, N168);
not NOT1 (N2417, N2406);
and AND2 (N2418, N2415, N2088);
and AND4 (N2419, N2418, N2403, N303, N1076);
and AND2 (N2420, N2417, N1135);
nor NOR2 (N2421, N2399, N2318);
and AND2 (N2422, N2410, N948);
nand NAND2 (N2423, N2421, N464);
or OR4 (N2424, N2412, N1772, N665, N1580);
nor NOR2 (N2425, N2420, N1388);
and AND4 (N2426, N2419, N1742, N1165, N1843);
and AND4 (N2427, N2409, N876, N449, N580);
nand NAND4 (N2428, N2426, N2265, N2119, N421);
buf BUF1 (N2429, N2401);
nor NOR2 (N2430, N2416, N378);
or OR2 (N2431, N2424, N2128);
nand NAND2 (N2432, N2428, N115);
or OR2 (N2433, N2427, N182);
nor NOR3 (N2434, N2431, N911, N581);
and AND4 (N2435, N2429, N372, N1575, N1307);
or OR2 (N2436, N2434, N1163);
and AND3 (N2437, N2395, N2204, N32);
nand NAND3 (N2438, N2430, N691, N1591);
nand NAND3 (N2439, N2438, N1027, N2148);
and AND3 (N2440, N2423, N786, N328);
and AND3 (N2441, N2436, N1269, N1448);
not NOT1 (N2442, N2439);
and AND4 (N2443, N2435, N283, N2065, N1804);
nand NAND2 (N2444, N2442, N1496);
and AND2 (N2445, N2441, N1461);
xor XOR2 (N2446, N2437, N1635);
or OR3 (N2447, N2446, N968, N1882);
not NOT1 (N2448, N2433);
and AND3 (N2449, N2445, N2027, N1683);
nand NAND3 (N2450, N2422, N1166, N70);
or OR4 (N2451, N2432, N223, N93, N1086);
xor XOR2 (N2452, N2443, N153);
buf BUF1 (N2453, N2444);
nor NOR4 (N2454, N2450, N2265, N1385, N791);
and AND2 (N2455, N2448, N2120);
or OR3 (N2456, N2454, N736, N1085);
xor XOR2 (N2457, N2455, N1704);
buf BUF1 (N2458, N2440);
nand NAND3 (N2459, N2451, N2007, N1895);
buf BUF1 (N2460, N2447);
or OR2 (N2461, N2456, N1020);
nor NOR4 (N2462, N2457, N1442, N113, N2387);
buf BUF1 (N2463, N2425);
nor NOR3 (N2464, N2449, N540, N566);
nor NOR4 (N2465, N2463, N1787, N1211, N1229);
buf BUF1 (N2466, N2414);
or OR4 (N2467, N2453, N1257, N1611, N813);
nor NOR2 (N2468, N2460, N1549);
buf BUF1 (N2469, N2467);
not NOT1 (N2470, N2461);
nand NAND4 (N2471, N2465, N398, N1083, N1441);
not NOT1 (N2472, N2469);
nor NOR3 (N2473, N2464, N780, N2364);
xor XOR2 (N2474, N2470, N339);
nand NAND2 (N2475, N2472, N2154);
buf BUF1 (N2476, N2471);
and AND2 (N2477, N2466, N778);
nor NOR4 (N2478, N2473, N1605, N1810, N2352);
nor NOR2 (N2479, N2458, N212);
not NOT1 (N2480, N2474);
xor XOR2 (N2481, N2476, N160);
nor NOR4 (N2482, N2459, N2003, N2114, N1115);
and AND2 (N2483, N2452, N794);
buf BUF1 (N2484, N2483);
or OR2 (N2485, N2481, N781);
nor NOR2 (N2486, N2478, N1665);
xor XOR2 (N2487, N2484, N33);
nand NAND3 (N2488, N2487, N1256, N1284);
xor XOR2 (N2489, N2475, N1222);
not NOT1 (N2490, N2482);
nor NOR2 (N2491, N2486, N1896);
not NOT1 (N2492, N2490);
nor NOR4 (N2493, N2480, N168, N771, N720);
nand NAND4 (N2494, N2493, N233, N1972, N1691);
or OR2 (N2495, N2479, N1739);
buf BUF1 (N2496, N2491);
or OR2 (N2497, N2489, N2023);
or OR4 (N2498, N2494, N1808, N1359, N1210);
xor XOR2 (N2499, N2498, N2094);
buf BUF1 (N2500, N2499);
xor XOR2 (N2501, N2488, N2074);
nand NAND3 (N2502, N2497, N1541, N2396);
nand NAND3 (N2503, N2501, N2289, N1672);
nor NOR2 (N2504, N2495, N933);
buf BUF1 (N2505, N2492);
buf BUF1 (N2506, N2505);
buf BUF1 (N2507, N2504);
not NOT1 (N2508, N2503);
buf BUF1 (N2509, N2496);
or OR4 (N2510, N2506, N1820, N152, N1192);
buf BUF1 (N2511, N2510);
nand NAND4 (N2512, N2508, N177, N1078, N644);
buf BUF1 (N2513, N2477);
not NOT1 (N2514, N2468);
buf BUF1 (N2515, N2507);
and AND3 (N2516, N2512, N2363, N231);
nand NAND4 (N2517, N2515, N1302, N1188, N2352);
nor NOR4 (N2518, N2513, N244, N2343, N2404);
or OR3 (N2519, N2514, N1940, N652);
nor NOR3 (N2520, N2462, N646, N930);
and AND4 (N2521, N2485, N231, N1199, N2046);
nand NAND4 (N2522, N2521, N1046, N2186, N400);
and AND4 (N2523, N2502, N1261, N1270, N1142);
buf BUF1 (N2524, N2522);
and AND2 (N2525, N2509, N1971);
nor NOR4 (N2526, N2518, N291, N686, N1768);
nor NOR2 (N2527, N2511, N726);
nor NOR3 (N2528, N2519, N501, N250);
or OR2 (N2529, N2500, N2099);
not NOT1 (N2530, N2529);
xor XOR2 (N2531, N2517, N1675);
nor NOR2 (N2532, N2526, N988);
buf BUF1 (N2533, N2530);
or OR3 (N2534, N2524, N222, N1904);
or OR2 (N2535, N2523, N1329);
buf BUF1 (N2536, N2532);
nor NOR2 (N2537, N2520, N1317);
xor XOR2 (N2538, N2534, N65);
not NOT1 (N2539, N2536);
nand NAND2 (N2540, N2527, N760);
nand NAND3 (N2541, N2533, N1693, N349);
or OR2 (N2542, N2525, N345);
or OR4 (N2543, N2541, N1120, N1392, N1551);
not NOT1 (N2544, N2531);
xor XOR2 (N2545, N2537, N1463);
and AND2 (N2546, N2538, N1183);
nor NOR2 (N2547, N2544, N2463);
or OR3 (N2548, N2547, N1749, N1542);
and AND3 (N2549, N2528, N1639, N1393);
not NOT1 (N2550, N2545);
buf BUF1 (N2551, N2549);
nor NOR3 (N2552, N2551, N620, N271);
or OR2 (N2553, N2535, N1528);
not NOT1 (N2554, N2548);
not NOT1 (N2555, N2546);
not NOT1 (N2556, N2516);
xor XOR2 (N2557, N2555, N1511);
nand NAND4 (N2558, N2553, N562, N2278, N1757);
or OR4 (N2559, N2557, N430, N1663, N670);
nor NOR3 (N2560, N2540, N2525, N367);
nor NOR4 (N2561, N2554, N1312, N1295, N458);
xor XOR2 (N2562, N2556, N1824);
buf BUF1 (N2563, N2559);
buf BUF1 (N2564, N2561);
or OR3 (N2565, N2542, N1133, N766);
and AND3 (N2566, N2562, N1386, N2132);
and AND2 (N2567, N2563, N59);
or OR3 (N2568, N2564, N2431, N668);
or OR4 (N2569, N2566, N1312, N32, N832);
nor NOR2 (N2570, N2568, N1055);
not NOT1 (N2571, N2543);
buf BUF1 (N2572, N2569);
and AND3 (N2573, N2565, N69, N1090);
not NOT1 (N2574, N2550);
not NOT1 (N2575, N2573);
and AND3 (N2576, N2539, N2093, N1302);
nor NOR2 (N2577, N2567, N2001);
nor NOR2 (N2578, N2552, N1387);
buf BUF1 (N2579, N2574);
nand NAND3 (N2580, N2579, N249, N1308);
buf BUF1 (N2581, N2580);
nor NOR4 (N2582, N2558, N2475, N2409, N1478);
nand NAND3 (N2583, N2578, N1974, N738);
xor XOR2 (N2584, N2583, N849);
buf BUF1 (N2585, N2572);
not NOT1 (N2586, N2577);
not NOT1 (N2587, N2560);
not NOT1 (N2588, N2584);
buf BUF1 (N2589, N2571);
nand NAND2 (N2590, N2589, N1978);
buf BUF1 (N2591, N2588);
buf BUF1 (N2592, N2576);
not NOT1 (N2593, N2586);
nand NAND4 (N2594, N2587, N126, N94, N946);
nor NOR3 (N2595, N2581, N795, N754);
xor XOR2 (N2596, N2595, N2161);
nand NAND4 (N2597, N2575, N1498, N2083, N2562);
or OR4 (N2598, N2594, N1593, N416, N382);
not NOT1 (N2599, N2590);
nor NOR3 (N2600, N2570, N2003, N1090);
buf BUF1 (N2601, N2596);
not NOT1 (N2602, N2600);
and AND2 (N2603, N2585, N1358);
not NOT1 (N2604, N2603);
or OR4 (N2605, N2602, N643, N717, N61);
buf BUF1 (N2606, N2601);
nand NAND4 (N2607, N2598, N2196, N1374, N770);
nor NOR2 (N2608, N2597, N258);
and AND2 (N2609, N2608, N536);
buf BUF1 (N2610, N2582);
nand NAND2 (N2611, N2599, N1829);
buf BUF1 (N2612, N2611);
and AND3 (N2613, N2607, N1509, N1152);
not NOT1 (N2614, N2593);
nor NOR4 (N2615, N2614, N752, N981, N2450);
buf BUF1 (N2616, N2592);
nor NOR2 (N2617, N2610, N1704);
and AND3 (N2618, N2615, N2019, N128);
not NOT1 (N2619, N2604);
and AND2 (N2620, N2618, N2545);
or OR2 (N2621, N2612, N199);
not NOT1 (N2622, N2609);
xor XOR2 (N2623, N2619, N533);
not NOT1 (N2624, N2617);
or OR4 (N2625, N2605, N220, N2594, N2226);
not NOT1 (N2626, N2613);
or OR3 (N2627, N2626, N46, N2104);
buf BUF1 (N2628, N2627);
buf BUF1 (N2629, N2621);
nor NOR2 (N2630, N2591, N2259);
not NOT1 (N2631, N2606);
xor XOR2 (N2632, N2623, N485);
xor XOR2 (N2633, N2631, N2462);
and AND2 (N2634, N2632, N31);
buf BUF1 (N2635, N2629);
nand NAND3 (N2636, N2628, N1614, N508);
nand NAND2 (N2637, N2630, N2586);
or OR3 (N2638, N2636, N1499, N871);
xor XOR2 (N2639, N2635, N1403);
nand NAND4 (N2640, N2624, N2274, N2328, N1052);
xor XOR2 (N2641, N2616, N1867);
not NOT1 (N2642, N2622);
or OR2 (N2643, N2634, N172);
and AND2 (N2644, N2637, N2584);
buf BUF1 (N2645, N2633);
not NOT1 (N2646, N2640);
or OR3 (N2647, N2643, N158, N2507);
or OR3 (N2648, N2625, N763, N1809);
or OR2 (N2649, N2647, N1979);
and AND2 (N2650, N2644, N634);
buf BUF1 (N2651, N2648);
buf BUF1 (N2652, N2641);
nor NOR3 (N2653, N2620, N777, N1238);
nand NAND2 (N2654, N2651, N1117);
nand NAND3 (N2655, N2653, N1166, N1498);
nand NAND4 (N2656, N2639, N1963, N671, N2065);
nor NOR2 (N2657, N2649, N914);
buf BUF1 (N2658, N2650);
xor XOR2 (N2659, N2655, N1620);
and AND3 (N2660, N2638, N1458, N1300);
buf BUF1 (N2661, N2654);
and AND4 (N2662, N2652, N536, N1245, N1455);
or OR4 (N2663, N2645, N196, N694, N43);
xor XOR2 (N2664, N2656, N693);
or OR4 (N2665, N2659, N1113, N2160, N1641);
nor NOR3 (N2666, N2661, N293, N1539);
not NOT1 (N2667, N2664);
or OR2 (N2668, N2663, N2628);
buf BUF1 (N2669, N2657);
not NOT1 (N2670, N2660);
and AND3 (N2671, N2658, N685, N389);
buf BUF1 (N2672, N2671);
not NOT1 (N2673, N2646);
buf BUF1 (N2674, N2670);
and AND4 (N2675, N2672, N68, N624, N1654);
xor XOR2 (N2676, N2673, N70);
or OR2 (N2677, N2676, N589);
nor NOR2 (N2678, N2668, N1046);
nand NAND2 (N2679, N2675, N1939);
and AND4 (N2680, N2677, N500, N139, N2253);
nor NOR4 (N2681, N2679, N1933, N476, N1315);
buf BUF1 (N2682, N2662);
nor NOR3 (N2683, N2682, N948, N2407);
nor NOR3 (N2684, N2667, N900, N1248);
buf BUF1 (N2685, N2678);
buf BUF1 (N2686, N2674);
and AND3 (N2687, N2666, N1829, N722);
xor XOR2 (N2688, N2687, N919);
buf BUF1 (N2689, N2642);
nand NAND4 (N2690, N2681, N628, N37, N1767);
xor XOR2 (N2691, N2688, N1268);
or OR3 (N2692, N2690, N2235, N1748);
or OR4 (N2693, N2686, N767, N1174, N2277);
or OR4 (N2694, N2669, N2676, N1371, N909);
nor NOR2 (N2695, N2684, N2175);
nor NOR3 (N2696, N2695, N2324, N166);
and AND3 (N2697, N2665, N985, N768);
buf BUF1 (N2698, N2689);
xor XOR2 (N2699, N2692, N486);
or OR4 (N2700, N2696, N1379, N2288, N734);
not NOT1 (N2701, N2698);
buf BUF1 (N2702, N2685);
nand NAND3 (N2703, N2694, N949, N2375);
xor XOR2 (N2704, N2691, N2563);
buf BUF1 (N2705, N2680);
nor NOR4 (N2706, N2700, N1503, N1329, N2023);
or OR2 (N2707, N2701, N1618);
or OR3 (N2708, N2693, N1202, N2570);
and AND4 (N2709, N2705, N1136, N200, N2641);
xor XOR2 (N2710, N2697, N2347);
or OR4 (N2711, N2699, N666, N2340, N42);
buf BUF1 (N2712, N2683);
buf BUF1 (N2713, N2708);
and AND2 (N2714, N2704, N372);
and AND2 (N2715, N2707, N279);
buf BUF1 (N2716, N2713);
nor NOR4 (N2717, N2714, N2609, N2200, N2151);
and AND2 (N2718, N2710, N924);
or OR4 (N2719, N2716, N768, N647, N175);
not NOT1 (N2720, N2719);
xor XOR2 (N2721, N2718, N2395);
buf BUF1 (N2722, N2715);
nor NOR2 (N2723, N2709, N1547);
and AND4 (N2724, N2717, N2389, N2593, N2228);
and AND4 (N2725, N2724, N277, N688, N2111);
or OR2 (N2726, N2721, N435);
and AND3 (N2727, N2703, N1974, N1480);
buf BUF1 (N2728, N2723);
buf BUF1 (N2729, N2726);
nor NOR4 (N2730, N2712, N2065, N1772, N1254);
buf BUF1 (N2731, N2706);
nor NOR4 (N2732, N2730, N1978, N1053, N2731);
not NOT1 (N2733, N1770);
and AND3 (N2734, N2720, N201, N267);
or OR3 (N2735, N2702, N1405, N2494);
not NOT1 (N2736, N2734);
xor XOR2 (N2737, N2722, N1076);
and AND3 (N2738, N2737, N2041, N1993);
and AND4 (N2739, N2738, N1932, N1347, N2460);
xor XOR2 (N2740, N2739, N1083);
not NOT1 (N2741, N2727);
buf BUF1 (N2742, N2711);
or OR2 (N2743, N2725, N1786);
and AND2 (N2744, N2735, N2483);
not NOT1 (N2745, N2740);
buf BUF1 (N2746, N2743);
not NOT1 (N2747, N2746);
or OR4 (N2748, N2747, N1583, N988, N2177);
and AND2 (N2749, N2744, N2684);
and AND3 (N2750, N2748, N1243, N1609);
and AND4 (N2751, N2728, N1894, N1738, N250);
nand NAND4 (N2752, N2745, N2008, N923, N34);
xor XOR2 (N2753, N2733, N297);
nor NOR4 (N2754, N2732, N2500, N2490, N335);
buf BUF1 (N2755, N2729);
nor NOR3 (N2756, N2752, N216, N1378);
xor XOR2 (N2757, N2742, N691);
xor XOR2 (N2758, N2754, N147);
nand NAND3 (N2759, N2741, N657, N2176);
nor NOR2 (N2760, N2753, N2687);
and AND4 (N2761, N2751, N754, N1225, N2332);
nor NOR3 (N2762, N2759, N1374, N2085);
buf BUF1 (N2763, N2756);
nand NAND3 (N2764, N2760, N505, N3);
or OR3 (N2765, N2750, N174, N1598);
or OR2 (N2766, N2758, N2321);
nand NAND4 (N2767, N2736, N619, N616, N2208);
or OR2 (N2768, N2766, N2373);
nand NAND3 (N2769, N2763, N2113, N1194);
xor XOR2 (N2770, N2769, N1894);
nor NOR3 (N2771, N2757, N1088, N1935);
and AND3 (N2772, N2764, N1600, N318);
xor XOR2 (N2773, N2749, N1953);
and AND3 (N2774, N2771, N1631, N1260);
and AND4 (N2775, N2772, N1978, N2205, N2610);
or OR4 (N2776, N2775, N2312, N2741, N1983);
not NOT1 (N2777, N2773);
and AND4 (N2778, N2755, N2631, N900, N2078);
xor XOR2 (N2779, N2770, N2066);
buf BUF1 (N2780, N2767);
buf BUF1 (N2781, N2779);
nand NAND2 (N2782, N2774, N2102);
xor XOR2 (N2783, N2762, N1718);
or OR4 (N2784, N2783, N2680, N1571, N2156);
nand NAND4 (N2785, N2780, N140, N2526, N1411);
xor XOR2 (N2786, N2785, N2246);
nor NOR2 (N2787, N2768, N196);
buf BUF1 (N2788, N2781);
not NOT1 (N2789, N2761);
nand NAND3 (N2790, N2776, N1092, N2115);
buf BUF1 (N2791, N2777);
or OR2 (N2792, N2788, N376);
nor NOR2 (N2793, N2791, N1404);
not NOT1 (N2794, N2782);
and AND3 (N2795, N2786, N2151, N2627);
nor NOR3 (N2796, N2790, N1414, N1499);
nand NAND3 (N2797, N2784, N750, N1274);
xor XOR2 (N2798, N2797, N2675);
buf BUF1 (N2799, N2787);
xor XOR2 (N2800, N2765, N2068);
and AND3 (N2801, N2778, N1280, N288);
xor XOR2 (N2802, N2798, N456);
nand NAND2 (N2803, N2799, N1414);
or OR3 (N2804, N2800, N2413, N2430);
or OR2 (N2805, N2803, N2170);
buf BUF1 (N2806, N2794);
not NOT1 (N2807, N2804);
xor XOR2 (N2808, N2806, N178);
buf BUF1 (N2809, N2796);
and AND2 (N2810, N2792, N1898);
and AND2 (N2811, N2793, N850);
buf BUF1 (N2812, N2808);
nor NOR3 (N2813, N2810, N251, N1288);
and AND3 (N2814, N2802, N284, N1732);
or OR2 (N2815, N2807, N2127);
nand NAND3 (N2816, N2789, N2344, N749);
and AND4 (N2817, N2815, N2797, N2681, N98);
not NOT1 (N2818, N2813);
and AND2 (N2819, N2805, N2180);
and AND2 (N2820, N2818, N1973);
and AND3 (N2821, N2817, N1313, N268);
buf BUF1 (N2822, N2816);
not NOT1 (N2823, N2822);
or OR4 (N2824, N2809, N1760, N211, N380);
buf BUF1 (N2825, N2821);
buf BUF1 (N2826, N2812);
buf BUF1 (N2827, N2825);
xor XOR2 (N2828, N2819, N280);
and AND3 (N2829, N2814, N338, N440);
xor XOR2 (N2830, N2811, N2160);
nor NOR3 (N2831, N2801, N1257, N93);
and AND2 (N2832, N2828, N1560);
not NOT1 (N2833, N2827);
buf BUF1 (N2834, N2824);
not NOT1 (N2835, N2833);
nand NAND2 (N2836, N2831, N1897);
nand NAND4 (N2837, N2823, N1580, N1244, N1915);
xor XOR2 (N2838, N2834, N2606);
xor XOR2 (N2839, N2795, N75);
buf BUF1 (N2840, N2838);
not NOT1 (N2841, N2829);
or OR3 (N2842, N2837, N1200, N619);
or OR2 (N2843, N2841, N7);
not NOT1 (N2844, N2842);
nor NOR4 (N2845, N2836, N1362, N797, N1089);
nor NOR4 (N2846, N2830, N2188, N2661, N1855);
nand NAND2 (N2847, N2844, N27);
not NOT1 (N2848, N2820);
nor NOR4 (N2849, N2848, N1985, N2588, N114);
xor XOR2 (N2850, N2840, N2457);
and AND3 (N2851, N2835, N896, N2079);
nand NAND2 (N2852, N2826, N2716);
and AND4 (N2853, N2843, N2700, N1096, N222);
buf BUF1 (N2854, N2839);
or OR4 (N2855, N2852, N1630, N653, N2258);
or OR2 (N2856, N2855, N2159);
or OR4 (N2857, N2854, N2292, N168, N961);
nor NOR3 (N2858, N2856, N1877, N163);
nand NAND3 (N2859, N2846, N1929, N643);
buf BUF1 (N2860, N2849);
nand NAND4 (N2861, N2853, N546, N2608, N406);
nor NOR4 (N2862, N2847, N687, N672, N1699);
nor NOR2 (N2863, N2832, N1855);
or OR2 (N2864, N2861, N1184);
nor NOR4 (N2865, N2850, N279, N812, N1549);
nor NOR3 (N2866, N2860, N2445, N2310);
xor XOR2 (N2867, N2857, N131);
xor XOR2 (N2868, N2866, N2397);
nor NOR4 (N2869, N2845, N161, N231, N2212);
xor XOR2 (N2870, N2864, N392);
and AND4 (N2871, N2858, N1259, N2793, N587);
not NOT1 (N2872, N2871);
not NOT1 (N2873, N2851);
or OR4 (N2874, N2873, N2296, N715, N726);
or OR4 (N2875, N2863, N1321, N1832, N2028);
nand NAND3 (N2876, N2870, N2707, N257);
not NOT1 (N2877, N2867);
xor XOR2 (N2878, N2875, N392);
buf BUF1 (N2879, N2874);
not NOT1 (N2880, N2869);
nand NAND4 (N2881, N2862, N610, N2708, N951);
and AND4 (N2882, N2877, N2395, N873, N1980);
buf BUF1 (N2883, N2876);
buf BUF1 (N2884, N2865);
or OR3 (N2885, N2859, N216, N2181);
nor NOR2 (N2886, N2879, N2579);
or OR2 (N2887, N2882, N102);
not NOT1 (N2888, N2881);
nand NAND3 (N2889, N2883, N1681, N2454);
not NOT1 (N2890, N2888);
not NOT1 (N2891, N2878);
nor NOR2 (N2892, N2886, N1155);
nor NOR3 (N2893, N2889, N2229, N1073);
nand NAND3 (N2894, N2880, N1165, N2251);
and AND4 (N2895, N2893, N73, N1476, N377);
xor XOR2 (N2896, N2891, N2837);
nand NAND2 (N2897, N2885, N198);
buf BUF1 (N2898, N2872);
xor XOR2 (N2899, N2898, N2165);
xor XOR2 (N2900, N2884, N606);
buf BUF1 (N2901, N2887);
nand NAND3 (N2902, N2899, N52, N644);
not NOT1 (N2903, N2896);
not NOT1 (N2904, N2902);
xor XOR2 (N2905, N2900, N1822);
nor NOR2 (N2906, N2892, N1042);
not NOT1 (N2907, N2868);
nor NOR4 (N2908, N2894, N494, N2164, N2890);
buf BUF1 (N2909, N2204);
or OR3 (N2910, N2895, N1283, N878);
nand NAND4 (N2911, N2897, N1150, N1619, N1142);
xor XOR2 (N2912, N2905, N1006);
xor XOR2 (N2913, N2901, N543);
buf BUF1 (N2914, N2913);
nand NAND2 (N2915, N2914, N1459);
not NOT1 (N2916, N2911);
and AND2 (N2917, N2910, N2646);
or OR2 (N2918, N2909, N1813);
xor XOR2 (N2919, N2912, N1603);
or OR3 (N2920, N2918, N1235, N1188);
nor NOR2 (N2921, N2907, N2315);
and AND2 (N2922, N2903, N225);
or OR4 (N2923, N2920, N1549, N1314, N2602);
and AND3 (N2924, N2923, N191, N922);
buf BUF1 (N2925, N2908);
or OR4 (N2926, N2915, N1909, N932, N2053);
nor NOR3 (N2927, N2926, N771, N585);
not NOT1 (N2928, N2919);
nor NOR3 (N2929, N2925, N634, N2399);
xor XOR2 (N2930, N2927, N1774);
buf BUF1 (N2931, N2904);
xor XOR2 (N2932, N2906, N840);
or OR3 (N2933, N2922, N2272, N1424);
not NOT1 (N2934, N2916);
or OR3 (N2935, N2928, N1914, N1897);
and AND3 (N2936, N2935, N1112, N2556);
and AND2 (N2937, N2930, N330);
and AND4 (N2938, N2931, N299, N2650, N1504);
buf BUF1 (N2939, N2933);
nor NOR2 (N2940, N2929, N1315);
not NOT1 (N2941, N2917);
buf BUF1 (N2942, N2937);
xor XOR2 (N2943, N2940, N508);
and AND3 (N2944, N2943, N2005, N2735);
and AND2 (N2945, N2941, N784);
and AND4 (N2946, N2934, N2052, N1768, N846);
nor NOR4 (N2947, N2946, N399, N2345, N230);
buf BUF1 (N2948, N2921);
or OR4 (N2949, N2944, N1802, N2307, N2001);
nor NOR3 (N2950, N2949, N2058, N2839);
or OR3 (N2951, N2938, N1038, N289);
buf BUF1 (N2952, N2947);
nand NAND4 (N2953, N2932, N680, N92, N625);
not NOT1 (N2954, N2948);
buf BUF1 (N2955, N2950);
xor XOR2 (N2956, N2924, N2905);
nand NAND4 (N2957, N2954, N2500, N2924, N1084);
xor XOR2 (N2958, N2936, N449);
buf BUF1 (N2959, N2957);
or OR2 (N2960, N2945, N1015);
xor XOR2 (N2961, N2959, N2891);
xor XOR2 (N2962, N2952, N1020);
nand NAND4 (N2963, N2961, N1881, N978, N68);
and AND4 (N2964, N2955, N1031, N2818, N2261);
or OR3 (N2965, N2942, N900, N2000);
xor XOR2 (N2966, N2964, N2720);
nor NOR2 (N2967, N2960, N402);
nand NAND4 (N2968, N2956, N1659, N1547, N1911);
nor NOR4 (N2969, N2962, N465, N2011, N1808);
and AND2 (N2970, N2967, N1762);
and AND2 (N2971, N2968, N363);
and AND3 (N2972, N2970, N2897, N2113);
not NOT1 (N2973, N2971);
or OR3 (N2974, N2973, N713, N527);
not NOT1 (N2975, N2953);
nand NAND2 (N2976, N2939, N2725);
nand NAND2 (N2977, N2965, N797);
buf BUF1 (N2978, N2966);
xor XOR2 (N2979, N2972, N1953);
and AND2 (N2980, N2963, N2039);
nor NOR2 (N2981, N2958, N1700);
nor NOR4 (N2982, N2951, N395, N1077, N2363);
not NOT1 (N2983, N2981);
buf BUF1 (N2984, N2979);
or OR2 (N2985, N2976, N1508);
xor XOR2 (N2986, N2978, N1960);
and AND2 (N2987, N2975, N2811);
and AND4 (N2988, N2984, N1778, N2595, N1852);
not NOT1 (N2989, N2982);
nor NOR4 (N2990, N2985, N781, N147, N87);
and AND2 (N2991, N2987, N1738);
buf BUF1 (N2992, N2977);
and AND3 (N2993, N2974, N2391, N427);
and AND3 (N2994, N2989, N2012, N2459);
or OR4 (N2995, N2983, N2413, N1611, N2293);
nor NOR4 (N2996, N2986, N1285, N2497, N548);
xor XOR2 (N2997, N2980, N2950);
nand NAND4 (N2998, N2992, N2686, N1242, N1851);
buf BUF1 (N2999, N2997);
and AND3 (N3000, N2995, N1810, N2648);
and AND4 (N3001, N2994, N77, N2403, N412);
buf BUF1 (N3002, N2991);
and AND4 (N3003, N2998, N265, N2491, N2497);
buf BUF1 (N3004, N2969);
not NOT1 (N3005, N3001);
and AND2 (N3006, N3005, N252);
or OR2 (N3007, N2996, N143);
xor XOR2 (N3008, N3003, N1062);
xor XOR2 (N3009, N3000, N942);
nand NAND4 (N3010, N3007, N1269, N254, N1947);
and AND2 (N3011, N2999, N594);
or OR3 (N3012, N3009, N2592, N334);
and AND3 (N3013, N3002, N2120, N581);
xor XOR2 (N3014, N3013, N2641);
and AND3 (N3015, N3006, N385, N2043);
nor NOR2 (N3016, N2988, N2347);
or OR2 (N3017, N3014, N2950);
xor XOR2 (N3018, N3016, N1988);
nor NOR4 (N3019, N3017, N1941, N27, N165);
nand NAND3 (N3020, N3004, N1170, N240);
and AND2 (N3021, N3018, N1610);
nand NAND3 (N3022, N3020, N1756, N1734);
not NOT1 (N3023, N3010);
or OR2 (N3024, N3022, N1661);
buf BUF1 (N3025, N3012);
xor XOR2 (N3026, N2993, N771);
and AND2 (N3027, N3024, N448);
xor XOR2 (N3028, N2990, N2214);
buf BUF1 (N3029, N3008);
buf BUF1 (N3030, N3015);
or OR2 (N3031, N3019, N1888);
xor XOR2 (N3032, N3023, N1848);
xor XOR2 (N3033, N3021, N71);
nand NAND4 (N3034, N3011, N731, N2419, N1948);
nor NOR3 (N3035, N3029, N870, N2);
buf BUF1 (N3036, N3033);
nand NAND3 (N3037, N3032, N1482, N2941);
not NOT1 (N3038, N3036);
nor NOR2 (N3039, N3031, N158);
nand NAND2 (N3040, N3035, N480);
nand NAND4 (N3041, N3030, N3023, N596, N2167);
nor NOR3 (N3042, N3026, N1560, N781);
buf BUF1 (N3043, N3037);
and AND3 (N3044, N3039, N2014, N2164);
nor NOR2 (N3045, N3043, N471);
not NOT1 (N3046, N3044);
nor NOR3 (N3047, N3038, N1549, N2118);
not NOT1 (N3048, N3025);
buf BUF1 (N3049, N3046);
or OR3 (N3050, N3045, N1857, N2879);
nand NAND3 (N3051, N3047, N129, N2895);
or OR3 (N3052, N3048, N823, N1792);
not NOT1 (N3053, N3051);
nand NAND2 (N3054, N3050, N346);
or OR2 (N3055, N3040, N2349);
nand NAND4 (N3056, N3027, N2717, N1563, N2551);
nand NAND3 (N3057, N3056, N1164, N796);
not NOT1 (N3058, N3057);
nand NAND4 (N3059, N3052, N1982, N525, N901);
xor XOR2 (N3060, N3034, N2104);
or OR2 (N3061, N3042, N1827);
nor NOR4 (N3062, N3053, N541, N1496, N1271);
nor NOR4 (N3063, N3059, N2572, N291, N228);
or OR3 (N3064, N3055, N1454, N2930);
or OR4 (N3065, N3054, N2310, N1534, N116);
xor XOR2 (N3066, N3063, N2167);
not NOT1 (N3067, N3066);
or OR3 (N3068, N3049, N772, N1733);
not NOT1 (N3069, N3041);
nand NAND3 (N3070, N3065, N2615, N28);
or OR3 (N3071, N3068, N1959, N2247);
nor NOR3 (N3072, N3071, N1713, N2224);
buf BUF1 (N3073, N3061);
xor XOR2 (N3074, N3072, N2179);
not NOT1 (N3075, N3074);
nand NAND4 (N3076, N3028, N2809, N72, N1088);
not NOT1 (N3077, N3069);
xor XOR2 (N3078, N3062, N564);
not NOT1 (N3079, N3058);
xor XOR2 (N3080, N3067, N2108);
nand NAND2 (N3081, N3060, N348);
and AND2 (N3082, N3075, N818);
or OR3 (N3083, N3078, N2198, N2822);
xor XOR2 (N3084, N3083, N1982);
and AND2 (N3085, N3064, N504);
nor NOR3 (N3086, N3070, N102, N1996);
not NOT1 (N3087, N3073);
or OR4 (N3088, N3082, N2273, N2976, N901);
and AND2 (N3089, N3088, N493);
buf BUF1 (N3090, N3089);
nor NOR3 (N3091, N3079, N1987, N1504);
nor NOR4 (N3092, N3087, N2379, N272, N1382);
and AND4 (N3093, N3085, N49, N535, N355);
xor XOR2 (N3094, N3076, N412);
not NOT1 (N3095, N3092);
xor XOR2 (N3096, N3095, N3045);
and AND3 (N3097, N3090, N592, N3034);
and AND3 (N3098, N3081, N371, N1497);
not NOT1 (N3099, N3077);
nand NAND4 (N3100, N3084, N1587, N2236, N2824);
nor NOR4 (N3101, N3091, N736, N360, N1922);
nand NAND4 (N3102, N3096, N2302, N2375, N94);
not NOT1 (N3103, N3086);
nor NOR2 (N3104, N3094, N1997);
nor NOR3 (N3105, N3102, N1719, N3100);
not NOT1 (N3106, N2989);
buf BUF1 (N3107, N3097);
buf BUF1 (N3108, N3099);
and AND4 (N3109, N3108, N2032, N2316, N2955);
xor XOR2 (N3110, N3080, N983);
not NOT1 (N3111, N3107);
or OR4 (N3112, N3111, N914, N367, N2212);
buf BUF1 (N3113, N3110);
nand NAND4 (N3114, N3109, N2903, N3019, N1367);
not NOT1 (N3115, N3112);
nor NOR3 (N3116, N3098, N885, N2416);
not NOT1 (N3117, N3105);
and AND2 (N3118, N3093, N2339);
buf BUF1 (N3119, N3114);
not NOT1 (N3120, N3115);
buf BUF1 (N3121, N3113);
nand NAND2 (N3122, N3116, N954);
xor XOR2 (N3123, N3120, N551);
not NOT1 (N3124, N3123);
nor NOR2 (N3125, N3121, N2972);
not NOT1 (N3126, N3106);
or OR2 (N3127, N3124, N266);
not NOT1 (N3128, N3104);
not NOT1 (N3129, N3117);
nor NOR2 (N3130, N3118, N2284);
nor NOR4 (N3131, N3103, N226, N1397, N2819);
nand NAND2 (N3132, N3127, N1046);
xor XOR2 (N3133, N3119, N311);
nor NOR4 (N3134, N3101, N2555, N769, N803);
and AND3 (N3135, N3133, N2315, N1588);
not NOT1 (N3136, N3129);
nor NOR4 (N3137, N3132, N1358, N3011, N1395);
xor XOR2 (N3138, N3136, N2057);
nand NAND3 (N3139, N3131, N2455, N147);
nand NAND3 (N3140, N3130, N851, N2815);
not NOT1 (N3141, N3140);
and AND2 (N3142, N3134, N1277);
nand NAND2 (N3143, N3128, N1486);
xor XOR2 (N3144, N3141, N2700);
not NOT1 (N3145, N3126);
buf BUF1 (N3146, N3137);
nor NOR2 (N3147, N3139, N3113);
nor NOR4 (N3148, N3144, N2254, N241, N793);
nand NAND3 (N3149, N3145, N1117, N1097);
or OR4 (N3150, N3135, N2386, N1863, N2737);
or OR2 (N3151, N3147, N261);
xor XOR2 (N3152, N3138, N2569);
nand NAND2 (N3153, N3143, N192);
xor XOR2 (N3154, N3146, N996);
buf BUF1 (N3155, N3148);
xor XOR2 (N3156, N3125, N104);
nor NOR3 (N3157, N3155, N618, N2448);
xor XOR2 (N3158, N3157, N802);
nand NAND2 (N3159, N3150, N1911);
nand NAND4 (N3160, N3152, N706, N1105, N1343);
not NOT1 (N3161, N3160);
buf BUF1 (N3162, N3142);
and AND3 (N3163, N3158, N18, N2130);
buf BUF1 (N3164, N3163);
nor NOR4 (N3165, N3162, N3045, N905, N2182);
and AND4 (N3166, N3165, N208, N477, N357);
and AND4 (N3167, N3156, N322, N1139, N984);
nor NOR2 (N3168, N3149, N923);
and AND3 (N3169, N3153, N2312, N45);
nor NOR3 (N3170, N3122, N2107, N1074);
xor XOR2 (N3171, N3167, N2827);
buf BUF1 (N3172, N3151);
buf BUF1 (N3173, N3169);
buf BUF1 (N3174, N3168);
and AND2 (N3175, N3154, N988);
buf BUF1 (N3176, N3164);
nor NOR3 (N3177, N3170, N556, N2142);
nand NAND2 (N3178, N3159, N843);
or OR4 (N3179, N3175, N2185, N2336, N1520);
nor NOR4 (N3180, N3172, N2744, N718, N575);
buf BUF1 (N3181, N3180);
and AND4 (N3182, N3166, N39, N850, N2385);
nand NAND2 (N3183, N3171, N1460);
not NOT1 (N3184, N3183);
and AND3 (N3185, N3177, N68, N2111);
or OR2 (N3186, N3179, N2349);
and AND2 (N3187, N3185, N1141);
nor NOR4 (N3188, N3173, N2289, N2208, N387);
not NOT1 (N3189, N3186);
or OR2 (N3190, N3182, N1698);
buf BUF1 (N3191, N3189);
or OR2 (N3192, N3184, N2048);
and AND2 (N3193, N3192, N2635);
nand NAND2 (N3194, N3187, N726);
and AND2 (N3195, N3181, N1490);
buf BUF1 (N3196, N3174);
or OR3 (N3197, N3188, N771, N2412);
not NOT1 (N3198, N3197);
or OR2 (N3199, N3161, N940);
nand NAND2 (N3200, N3176, N1897);
and AND4 (N3201, N3195, N324, N208, N812);
or OR2 (N3202, N3193, N473);
and AND3 (N3203, N3191, N1189, N2137);
or OR4 (N3204, N3202, N2231, N2450, N1049);
not NOT1 (N3205, N3198);
or OR3 (N3206, N3201, N1947, N679);
and AND3 (N3207, N3206, N1866, N1765);
xor XOR2 (N3208, N3200, N2062);
nor NOR3 (N3209, N3204, N1452, N989);
not NOT1 (N3210, N3203);
and AND4 (N3211, N3208, N1590, N782, N38);
not NOT1 (N3212, N3209);
nor NOR4 (N3213, N3178, N1941, N19, N811);
xor XOR2 (N3214, N3213, N1809);
or OR2 (N3215, N3214, N1013);
xor XOR2 (N3216, N3212, N2525);
not NOT1 (N3217, N3215);
nand NAND4 (N3218, N3205, N2984, N1015, N657);
nor NOR4 (N3219, N3207, N1150, N2253, N999);
or OR2 (N3220, N3216, N2216);
and AND4 (N3221, N3190, N1007, N1420, N1948);
nand NAND3 (N3222, N3210, N1815, N466);
or OR3 (N3223, N3219, N2893, N2472);
nor NOR3 (N3224, N3211, N430, N2708);
buf BUF1 (N3225, N3217);
nand NAND4 (N3226, N3218, N9, N216, N1582);
nand NAND3 (N3227, N3225, N1793, N59);
buf BUF1 (N3228, N3221);
buf BUF1 (N3229, N3196);
nand NAND2 (N3230, N3194, N1723);
nor NOR3 (N3231, N3220, N2870, N1884);
or OR3 (N3232, N3222, N851, N2295);
nand NAND4 (N3233, N3224, N215, N595, N353);
and AND3 (N3234, N3230, N1820, N792);
nor NOR4 (N3235, N3231, N1624, N1067, N259);
not NOT1 (N3236, N3199);
or OR3 (N3237, N3229, N3162, N885);
buf BUF1 (N3238, N3236);
or OR3 (N3239, N3237, N1504, N705);
buf BUF1 (N3240, N3226);
buf BUF1 (N3241, N3234);
not NOT1 (N3242, N3241);
not NOT1 (N3243, N3235);
buf BUF1 (N3244, N3227);
or OR2 (N3245, N3239, N1355);
not NOT1 (N3246, N3223);
or OR4 (N3247, N3240, N2529, N1170, N219);
xor XOR2 (N3248, N3238, N671);
nor NOR4 (N3249, N3232, N1120, N14, N2812);
not NOT1 (N3250, N3242);
buf BUF1 (N3251, N3233);
xor XOR2 (N3252, N3244, N251);
nor NOR4 (N3253, N3228, N2157, N2395, N2570);
and AND2 (N3254, N3250, N1829);
not NOT1 (N3255, N3254);
nor NOR3 (N3256, N3246, N544, N81);
and AND3 (N3257, N3252, N2038, N59);
or OR4 (N3258, N3256, N2657, N2364, N306);
xor XOR2 (N3259, N3243, N833);
and AND4 (N3260, N3245, N2012, N2045, N157);
nand NAND4 (N3261, N3248, N1481, N752, N1090);
nand NAND2 (N3262, N3253, N3188);
not NOT1 (N3263, N3249);
or OR2 (N3264, N3263, N342);
nand NAND2 (N3265, N3247, N652);
xor XOR2 (N3266, N3262, N1915);
or OR2 (N3267, N3265, N1040);
nand NAND3 (N3268, N3261, N3045, N1606);
buf BUF1 (N3269, N3260);
not NOT1 (N3270, N3267);
xor XOR2 (N3271, N3255, N1121);
xor XOR2 (N3272, N3266, N2908);
nor NOR4 (N3273, N3259, N1714, N1, N1771);
not NOT1 (N3274, N3270);
not NOT1 (N3275, N3271);
buf BUF1 (N3276, N3251);
xor XOR2 (N3277, N3276, N1791);
xor XOR2 (N3278, N3269, N3037);
not NOT1 (N3279, N3268);
buf BUF1 (N3280, N3273);
not NOT1 (N3281, N3272);
nor NOR3 (N3282, N3280, N1208, N1668);
nand NAND2 (N3283, N3279, N2567);
or OR4 (N3284, N3264, N1416, N741, N1869);
and AND4 (N3285, N3257, N2956, N214, N2088);
xor XOR2 (N3286, N3278, N2812);
or OR3 (N3287, N3275, N210, N1797);
or OR3 (N3288, N3285, N1081, N265);
nor NOR2 (N3289, N3282, N795);
nand NAND3 (N3290, N3286, N1176, N1210);
buf BUF1 (N3291, N3287);
xor XOR2 (N3292, N3288, N3061);
not NOT1 (N3293, N3292);
not NOT1 (N3294, N3277);
or OR3 (N3295, N3291, N2239, N2174);
buf BUF1 (N3296, N3289);
or OR4 (N3297, N3284, N1739, N3198, N2327);
nand NAND4 (N3298, N3295, N974, N906, N1843);
nor NOR4 (N3299, N3298, N2141, N3285, N1999);
or OR3 (N3300, N3258, N2329, N2488);
not NOT1 (N3301, N3299);
not NOT1 (N3302, N3301);
buf BUF1 (N3303, N3296);
or OR4 (N3304, N3283, N1003, N2179, N1140);
buf BUF1 (N3305, N3304);
nand NAND3 (N3306, N3303, N3301, N1827);
xor XOR2 (N3307, N3305, N3123);
xor XOR2 (N3308, N3307, N885);
xor XOR2 (N3309, N3293, N2785);
buf BUF1 (N3310, N3274);
or OR4 (N3311, N3294, N2374, N2930, N40);
and AND2 (N3312, N3290, N179);
and AND2 (N3313, N3312, N2900);
nand NAND4 (N3314, N3302, N1629, N1098, N1785);
xor XOR2 (N3315, N3281, N233);
not NOT1 (N3316, N3315);
nand NAND2 (N3317, N3311, N1463);
and AND4 (N3318, N3310, N580, N107, N1907);
not NOT1 (N3319, N3316);
xor XOR2 (N3320, N3306, N505);
buf BUF1 (N3321, N3317);
not NOT1 (N3322, N3313);
nand NAND4 (N3323, N3322, N436, N1191, N2726);
or OR3 (N3324, N3314, N944, N2259);
and AND3 (N3325, N3320, N2011, N2080);
xor XOR2 (N3326, N3300, N2593);
nand NAND3 (N3327, N3318, N1964, N1697);
not NOT1 (N3328, N3308);
nor NOR3 (N3329, N3309, N840, N1564);
and AND3 (N3330, N3297, N1351, N1227);
buf BUF1 (N3331, N3319);
nand NAND3 (N3332, N3328, N1710, N172);
xor XOR2 (N3333, N3321, N770);
xor XOR2 (N3334, N3332, N2684);
not NOT1 (N3335, N3331);
nor NOR4 (N3336, N3333, N1253, N1291, N1028);
nor NOR4 (N3337, N3334, N2750, N1665, N3031);
and AND4 (N3338, N3323, N2337, N1098, N1700);
buf BUF1 (N3339, N3338);
xor XOR2 (N3340, N3339, N890);
xor XOR2 (N3341, N3336, N256);
not NOT1 (N3342, N3341);
not NOT1 (N3343, N3324);
nand NAND4 (N3344, N3343, N167, N772, N830);
nor NOR4 (N3345, N3337, N463, N2328, N3275);
buf BUF1 (N3346, N3325);
nand NAND3 (N3347, N3327, N2904, N1970);
not NOT1 (N3348, N3329);
not NOT1 (N3349, N3335);
nor NOR2 (N3350, N3342, N24);
and AND4 (N3351, N3330, N233, N1137, N2384);
or OR3 (N3352, N3351, N828, N1914);
xor XOR2 (N3353, N3347, N2911);
not NOT1 (N3354, N3349);
not NOT1 (N3355, N3344);
xor XOR2 (N3356, N3352, N1080);
and AND2 (N3357, N3348, N353);
not NOT1 (N3358, N3346);
or OR3 (N3359, N3356, N1789, N3155);
xor XOR2 (N3360, N3357, N1763);
nor NOR2 (N3361, N3350, N3050);
or OR2 (N3362, N3355, N491);
nand NAND4 (N3363, N3345, N1336, N2185, N2108);
xor XOR2 (N3364, N3326, N720);
or OR2 (N3365, N3354, N1677);
nand NAND4 (N3366, N3358, N722, N29, N898);
nand NAND2 (N3367, N3363, N168);
not NOT1 (N3368, N3340);
xor XOR2 (N3369, N3359, N1357);
xor XOR2 (N3370, N3360, N784);
nand NAND2 (N3371, N3366, N2609);
nand NAND4 (N3372, N3365, N2572, N2823, N1768);
buf BUF1 (N3373, N3368);
xor XOR2 (N3374, N3371, N315);
buf BUF1 (N3375, N3373);
nand NAND4 (N3376, N3370, N2694, N3164, N2890);
nand NAND4 (N3377, N3364, N1632, N2003, N31);
xor XOR2 (N3378, N3376, N1326);
nand NAND2 (N3379, N3377, N2332);
nor NOR2 (N3380, N3367, N3043);
nor NOR4 (N3381, N3379, N761, N3332, N2952);
nor NOR2 (N3382, N3369, N66);
not NOT1 (N3383, N3382);
xor XOR2 (N3384, N3380, N2072);
xor XOR2 (N3385, N3374, N1701);
nand NAND2 (N3386, N3362, N1849);
not NOT1 (N3387, N3375);
and AND4 (N3388, N3384, N971, N2051, N3046);
not NOT1 (N3389, N3381);
nor NOR2 (N3390, N3389, N1181);
nor NOR4 (N3391, N3361, N2390, N1045, N376);
and AND4 (N3392, N3391, N2919, N3064, N448);
xor XOR2 (N3393, N3385, N2403);
or OR3 (N3394, N3388, N1688, N3284);
nand NAND4 (N3395, N3383, N2392, N1816, N1099);
not NOT1 (N3396, N3392);
or OR4 (N3397, N3353, N430, N2828, N590);
nor NOR2 (N3398, N3378, N3245);
nand NAND4 (N3399, N3393, N2680, N1651, N3185);
nor NOR4 (N3400, N3386, N2057, N230, N2183);
and AND3 (N3401, N3398, N1076, N3100);
buf BUF1 (N3402, N3390);
or OR4 (N3403, N3395, N342, N2421, N1483);
xor XOR2 (N3404, N3400, N2058);
and AND3 (N3405, N3402, N2488, N1582);
and AND4 (N3406, N3397, N2940, N693, N1937);
nor NOR2 (N3407, N3394, N2333);
not NOT1 (N3408, N3407);
not NOT1 (N3409, N3405);
or OR4 (N3410, N3399, N1166, N1103, N1842);
xor XOR2 (N3411, N3410, N722);
not NOT1 (N3412, N3401);
nor NOR4 (N3413, N3406, N482, N469, N53);
or OR3 (N3414, N3412, N713, N3227);
and AND2 (N3415, N3408, N1038);
nand NAND4 (N3416, N3403, N802, N1408, N3334);
not NOT1 (N3417, N3415);
nand NAND2 (N3418, N3409, N1572);
buf BUF1 (N3419, N3404);
buf BUF1 (N3420, N3416);
buf BUF1 (N3421, N3420);
or OR3 (N3422, N3418, N3137, N94);
and AND2 (N3423, N3417, N1969);
buf BUF1 (N3424, N3411);
and AND3 (N3425, N3413, N806, N2024);
xor XOR2 (N3426, N3387, N2787);
or OR2 (N3427, N3425, N341);
or OR4 (N3428, N3396, N183, N208, N1144);
xor XOR2 (N3429, N3428, N1861);
nand NAND2 (N3430, N3424, N2568);
not NOT1 (N3431, N3430);
and AND3 (N3432, N3414, N1386, N681);
buf BUF1 (N3433, N3427);
nand NAND4 (N3434, N3422, N1042, N1666, N2920);
buf BUF1 (N3435, N3434);
buf BUF1 (N3436, N3432);
or OR3 (N3437, N3436, N2089, N2137);
nor NOR2 (N3438, N3437, N3272);
and AND4 (N3439, N3431, N2370, N541, N2226);
not NOT1 (N3440, N3419);
and AND3 (N3441, N3439, N3277, N2774);
not NOT1 (N3442, N3433);
nand NAND4 (N3443, N3438, N1217, N617, N3);
xor XOR2 (N3444, N3372, N1943);
and AND3 (N3445, N3429, N2025, N1960);
and AND4 (N3446, N3426, N3391, N1892, N2175);
nor NOR3 (N3447, N3443, N209, N1369);
or OR2 (N3448, N3440, N863);
xor XOR2 (N3449, N3421, N2745);
buf BUF1 (N3450, N3449);
and AND4 (N3451, N3423, N692, N3245, N413);
buf BUF1 (N3452, N3445);
or OR2 (N3453, N3446, N1145);
not NOT1 (N3454, N3453);
buf BUF1 (N3455, N3444);
nor NOR3 (N3456, N3442, N2052, N374);
not NOT1 (N3457, N3451);
not NOT1 (N3458, N3450);
nand NAND2 (N3459, N3454, N1312);
and AND4 (N3460, N3458, N1401, N341, N1697);
and AND4 (N3461, N3447, N373, N666, N2618);
nand NAND3 (N3462, N3452, N2696, N1627);
nor NOR3 (N3463, N3459, N709, N2320);
xor XOR2 (N3464, N3457, N236);
xor XOR2 (N3465, N3460, N3201);
or OR2 (N3466, N3463, N2088);
buf BUF1 (N3467, N3464);
xor XOR2 (N3468, N3455, N1072);
buf BUF1 (N3469, N3461);
nand NAND3 (N3470, N3448, N1215, N2392);
not NOT1 (N3471, N3468);
or OR2 (N3472, N3465, N2365);
nand NAND3 (N3473, N3467, N326, N2097);
or OR2 (N3474, N3441, N3150);
xor XOR2 (N3475, N3473, N3311);
buf BUF1 (N3476, N3462);
buf BUF1 (N3477, N3475);
nor NOR3 (N3478, N3469, N101, N3237);
xor XOR2 (N3479, N3477, N1480);
xor XOR2 (N3480, N3474, N3343);
or OR3 (N3481, N3466, N2956, N927);
or OR2 (N3482, N3456, N730);
xor XOR2 (N3483, N3470, N1080);
or OR3 (N3484, N3472, N638, N1324);
not NOT1 (N3485, N3482);
xor XOR2 (N3486, N3435, N1209);
and AND2 (N3487, N3485, N1299);
or OR2 (N3488, N3479, N1369);
xor XOR2 (N3489, N3486, N496);
or OR2 (N3490, N3487, N666);
not NOT1 (N3491, N3478);
or OR4 (N3492, N3488, N3012, N553, N2517);
nor NOR3 (N3493, N3480, N2979, N3323);
nand NAND4 (N3494, N3471, N2080, N399, N2505);
nand NAND3 (N3495, N3484, N2560, N311);
nand NAND2 (N3496, N3481, N1246);
not NOT1 (N3497, N3476);
nor NOR3 (N3498, N3497, N2778, N1548);
or OR4 (N3499, N3495, N534, N88, N712);
or OR3 (N3500, N3499, N791, N2457);
not NOT1 (N3501, N3490);
not NOT1 (N3502, N3489);
nor NOR3 (N3503, N3483, N2935, N1152);
xor XOR2 (N3504, N3498, N1894);
nor NOR4 (N3505, N3501, N775, N2584, N738);
nor NOR3 (N3506, N3505, N1191, N2527);
buf BUF1 (N3507, N3502);
xor XOR2 (N3508, N3492, N2796);
and AND2 (N3509, N3504, N3442);
buf BUF1 (N3510, N3496);
not NOT1 (N3511, N3509);
xor XOR2 (N3512, N3500, N3409);
nand NAND2 (N3513, N3503, N2899);
or OR4 (N3514, N3493, N2717, N3006, N1441);
or OR4 (N3515, N3511, N1437, N1359, N116);
and AND3 (N3516, N3506, N601, N1957);
and AND2 (N3517, N3508, N449);
nand NAND4 (N3518, N3507, N1571, N3031, N2955);
or OR4 (N3519, N3510, N518, N77, N3044);
not NOT1 (N3520, N3518);
endmodule