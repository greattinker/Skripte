// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15;

output N810,N796,N812,N808,N807,N811,N814,N805,N806,N815;

not NOT1 (N16, N13);
not NOT1 (N17, N8);
xor XOR2 (N18, N1, N9);
nor NOR4 (N19, N15, N5, N10, N4);
nand NAND3 (N20, N4, N1, N7);
not NOT1 (N21, N11);
nand NAND3 (N22, N11, N1, N18);
or OR2 (N23, N2, N5);
nor NOR2 (N24, N13, N10);
nor NOR2 (N25, N8, N17);
not NOT1 (N26, N6);
and AND3 (N27, N11, N11, N18);
not NOT1 (N28, N25);
buf BUF1 (N29, N28);
xor XOR2 (N30, N16, N10);
nor NOR2 (N31, N20, N13);
and AND2 (N32, N27, N8);
nor NOR2 (N33, N29, N32);
not NOT1 (N34, N32);
nor NOR4 (N35, N23, N8, N17, N4);
or OR3 (N36, N19, N10, N25);
or OR3 (N37, N31, N28, N13);
buf BUF1 (N38, N24);
nor NOR2 (N39, N30, N8);
nor NOR2 (N40, N22, N2);
xor XOR2 (N41, N37, N37);
or OR4 (N42, N21, N6, N40, N11);
nand NAND2 (N43, N7, N10);
xor XOR2 (N44, N43, N12);
not NOT1 (N45, N26);
xor XOR2 (N46, N44, N12);
not NOT1 (N47, N38);
buf BUF1 (N48, N33);
and AND2 (N49, N46, N4);
not NOT1 (N50, N42);
buf BUF1 (N51, N50);
xor XOR2 (N52, N35, N17);
nand NAND3 (N53, N48, N27, N17);
and AND3 (N54, N49, N18, N43);
or OR4 (N55, N53, N27, N41, N45);
nor NOR2 (N56, N13, N21);
not NOT1 (N57, N30);
and AND2 (N58, N57, N4);
or OR3 (N59, N54, N26, N2);
xor XOR2 (N60, N51, N38);
nor NOR2 (N61, N58, N15);
or OR3 (N62, N56, N13, N9);
buf BUF1 (N63, N61);
or OR3 (N64, N60, N14, N23);
not NOT1 (N65, N59);
or OR3 (N66, N52, N41, N49);
not NOT1 (N67, N62);
or OR3 (N68, N64, N1, N40);
buf BUF1 (N69, N66);
not NOT1 (N70, N65);
and AND4 (N71, N39, N13, N29, N61);
nand NAND3 (N72, N69, N39, N55);
nor NOR4 (N73, N72, N1, N58, N34);
nor NOR3 (N74, N29, N46, N57);
and AND4 (N75, N36, N30, N68, N49);
and AND3 (N76, N26, N47, N40);
xor XOR2 (N77, N33, N44);
or OR4 (N78, N42, N48, N8, N39);
nor NOR2 (N79, N74, N61);
buf BUF1 (N80, N71);
nand NAND4 (N81, N79, N41, N25, N52);
or OR4 (N82, N76, N44, N54, N33);
buf BUF1 (N83, N77);
nor NOR4 (N84, N63, N42, N60, N38);
nor NOR2 (N85, N81, N35);
xor XOR2 (N86, N70, N85);
not NOT1 (N87, N9);
xor XOR2 (N88, N86, N7);
nor NOR4 (N89, N78, N28, N85, N75);
nand NAND3 (N90, N45, N71, N59);
and AND2 (N91, N88, N18);
or OR4 (N92, N83, N55, N10, N8);
buf BUF1 (N93, N90);
not NOT1 (N94, N84);
or OR4 (N95, N93, N1, N35, N34);
or OR3 (N96, N82, N57, N6);
xor XOR2 (N97, N96, N90);
nor NOR4 (N98, N67, N31, N96, N28);
and AND4 (N99, N73, N28, N73, N78);
nand NAND4 (N100, N87, N65, N21, N86);
buf BUF1 (N101, N98);
or OR3 (N102, N99, N3, N18);
and AND2 (N103, N89, N40);
and AND3 (N104, N102, N96, N89);
nor NOR2 (N105, N94, N34);
xor XOR2 (N106, N91, N1);
buf BUF1 (N107, N95);
not NOT1 (N108, N107);
nor NOR2 (N109, N97, N18);
nor NOR2 (N110, N106, N97);
buf BUF1 (N111, N104);
and AND4 (N112, N108, N35, N95, N85);
not NOT1 (N113, N112);
nor NOR4 (N114, N100, N85, N8, N58);
buf BUF1 (N115, N103);
buf BUF1 (N116, N111);
nand NAND4 (N117, N114, N45, N109, N9);
xor XOR2 (N118, N28, N84);
or OR3 (N119, N117, N69, N25);
nand NAND4 (N120, N119, N16, N94, N80);
xor XOR2 (N121, N55, N21);
nor NOR3 (N122, N92, N108, N63);
and AND3 (N123, N110, N117, N73);
nor NOR2 (N124, N101, N19);
not NOT1 (N125, N105);
nand NAND3 (N126, N124, N66, N62);
not NOT1 (N127, N121);
xor XOR2 (N128, N115, N27);
nand NAND4 (N129, N118, N102, N54, N79);
not NOT1 (N130, N122);
not NOT1 (N131, N120);
or OR4 (N132, N131, N14, N128, N18);
xor XOR2 (N133, N100, N95);
not NOT1 (N134, N125);
nand NAND2 (N135, N127, N125);
xor XOR2 (N136, N129, N117);
not NOT1 (N137, N116);
xor XOR2 (N138, N126, N35);
nand NAND2 (N139, N132, N98);
nand NAND2 (N140, N139, N94);
not NOT1 (N141, N134);
nand NAND2 (N142, N136, N16);
and AND4 (N143, N133, N107, N92, N61);
and AND4 (N144, N123, N132, N134, N77);
or OR4 (N145, N143, N138, N22, N38);
xor XOR2 (N146, N92, N21);
buf BUF1 (N147, N113);
and AND4 (N148, N140, N53, N46, N128);
or OR3 (N149, N142, N24, N123);
nand NAND4 (N150, N141, N21, N75, N110);
xor XOR2 (N151, N149, N95);
buf BUF1 (N152, N145);
buf BUF1 (N153, N144);
buf BUF1 (N154, N146);
buf BUF1 (N155, N150);
xor XOR2 (N156, N137, N100);
and AND4 (N157, N130, N120, N99, N50);
buf BUF1 (N158, N135);
or OR2 (N159, N153, N138);
xor XOR2 (N160, N157, N58);
and AND2 (N161, N160, N13);
buf BUF1 (N162, N152);
xor XOR2 (N163, N158, N72);
not NOT1 (N164, N161);
xor XOR2 (N165, N159, N81);
nor NOR4 (N166, N164, N103, N138, N73);
not NOT1 (N167, N156);
nand NAND2 (N168, N148, N161);
nand NAND2 (N169, N154, N156);
xor XOR2 (N170, N163, N6);
xor XOR2 (N171, N147, N28);
nand NAND3 (N172, N168, N31, N24);
not NOT1 (N173, N165);
or OR4 (N174, N151, N117, N161, N31);
and AND4 (N175, N162, N108, N19, N7);
xor XOR2 (N176, N155, N130);
not NOT1 (N177, N175);
and AND2 (N178, N171, N15);
nor NOR2 (N179, N177, N48);
not NOT1 (N180, N170);
not NOT1 (N181, N172);
xor XOR2 (N182, N180, N4);
xor XOR2 (N183, N174, N69);
nand NAND3 (N184, N181, N85, N79);
or OR4 (N185, N166, N167, N142, N47);
not NOT1 (N186, N18);
nor NOR2 (N187, N178, N58);
nor NOR2 (N188, N169, N62);
or OR2 (N189, N188, N99);
not NOT1 (N190, N189);
nand NAND2 (N191, N187, N124);
xor XOR2 (N192, N176, N129);
or OR2 (N193, N191, N4);
not NOT1 (N194, N193);
nand NAND3 (N195, N173, N81, N123);
nor NOR4 (N196, N185, N192, N97, N25);
nand NAND3 (N197, N50, N22, N56);
buf BUF1 (N198, N184);
xor XOR2 (N199, N183, N7);
nor NOR3 (N200, N197, N171, N25);
not NOT1 (N201, N179);
not NOT1 (N202, N196);
and AND4 (N203, N190, N134, N79, N140);
xor XOR2 (N204, N200, N136);
not NOT1 (N205, N203);
xor XOR2 (N206, N204, N26);
buf BUF1 (N207, N199);
and AND3 (N208, N202, N121, N107);
or OR3 (N209, N198, N176, N30);
not NOT1 (N210, N207);
not NOT1 (N211, N182);
buf BUF1 (N212, N210);
xor XOR2 (N213, N206, N55);
nand NAND2 (N214, N209, N18);
and AND2 (N215, N208, N185);
nand NAND3 (N216, N213, N102, N28);
xor XOR2 (N217, N215, N179);
buf BUF1 (N218, N201);
nor NOR2 (N219, N214, N16);
and AND3 (N220, N194, N219, N27);
not NOT1 (N221, N116);
nand NAND4 (N222, N218, N71, N139, N73);
nor NOR2 (N223, N205, N90);
or OR2 (N224, N222, N53);
and AND2 (N225, N223, N67);
xor XOR2 (N226, N221, N115);
buf BUF1 (N227, N217);
xor XOR2 (N228, N211, N17);
not NOT1 (N229, N225);
and AND4 (N230, N220, N85, N162, N175);
xor XOR2 (N231, N227, N223);
not NOT1 (N232, N224);
nand NAND4 (N233, N230, N139, N118, N102);
and AND3 (N234, N232, N30, N91);
nor NOR3 (N235, N228, N44, N94);
or OR4 (N236, N231, N222, N65, N171);
buf BUF1 (N237, N235);
nand NAND4 (N238, N229, N129, N141, N148);
nand NAND3 (N239, N212, N86, N2);
not NOT1 (N240, N186);
not NOT1 (N241, N234);
nor NOR4 (N242, N240, N164, N110, N229);
buf BUF1 (N243, N236);
xor XOR2 (N244, N216, N229);
nor NOR4 (N245, N238, N148, N165, N120);
and AND4 (N246, N239, N155, N35, N215);
nand NAND4 (N247, N237, N135, N68, N109);
buf BUF1 (N248, N243);
and AND3 (N249, N244, N17, N109);
and AND2 (N250, N247, N93);
or OR4 (N251, N241, N186, N223, N169);
nand NAND3 (N252, N226, N5, N222);
xor XOR2 (N253, N251, N98);
and AND2 (N254, N249, N230);
or OR2 (N255, N242, N6);
nor NOR3 (N256, N254, N160, N172);
not NOT1 (N257, N233);
buf BUF1 (N258, N195);
xor XOR2 (N259, N255, N150);
not NOT1 (N260, N250);
not NOT1 (N261, N258);
not NOT1 (N262, N252);
xor XOR2 (N263, N248, N43);
not NOT1 (N264, N245);
buf BUF1 (N265, N259);
or OR4 (N266, N262, N45, N195, N177);
nand NAND2 (N267, N260, N155);
nand NAND2 (N268, N256, N207);
nor NOR2 (N269, N265, N70);
or OR2 (N270, N261, N225);
and AND4 (N271, N266, N8, N198, N123);
or OR3 (N272, N253, N32, N139);
xor XOR2 (N273, N263, N185);
and AND3 (N274, N268, N269, N132);
nand NAND2 (N275, N103, N136);
buf BUF1 (N276, N267);
or OR4 (N277, N271, N216, N20, N167);
nor NOR3 (N278, N277, N169, N258);
and AND4 (N279, N264, N265, N55, N92);
nor NOR4 (N280, N276, N63, N234, N237);
or OR3 (N281, N280, N128, N26);
nand NAND3 (N282, N278, N221, N243);
not NOT1 (N283, N270);
or OR4 (N284, N282, N25, N163, N134);
nor NOR4 (N285, N284, N2, N274, N123);
xor XOR2 (N286, N229, N13);
not NOT1 (N287, N275);
nor NOR3 (N288, N285, N232, N205);
and AND4 (N289, N273, N155, N189, N59);
not NOT1 (N290, N289);
nor NOR2 (N291, N290, N149);
buf BUF1 (N292, N288);
buf BUF1 (N293, N246);
nand NAND4 (N294, N292, N47, N172, N225);
nand NAND2 (N295, N291, N78);
buf BUF1 (N296, N281);
buf BUF1 (N297, N293);
not NOT1 (N298, N297);
or OR4 (N299, N287, N226, N110, N111);
nand NAND2 (N300, N257, N270);
or OR3 (N301, N298, N83, N273);
buf BUF1 (N302, N279);
or OR2 (N303, N283, N286);
xor XOR2 (N304, N68, N234);
nor NOR2 (N305, N295, N79);
and AND4 (N306, N272, N144, N7, N160);
or OR4 (N307, N302, N172, N151, N142);
not NOT1 (N308, N299);
and AND3 (N309, N308, N161, N41);
xor XOR2 (N310, N307, N155);
not NOT1 (N311, N296);
nor NOR4 (N312, N300, N69, N270, N28);
buf BUF1 (N313, N305);
buf BUF1 (N314, N301);
xor XOR2 (N315, N306, N84);
and AND2 (N316, N294, N183);
nand NAND2 (N317, N316, N20);
nor NOR4 (N318, N314, N133, N234, N297);
nand NAND3 (N319, N318, N77, N162);
nand NAND3 (N320, N309, N259, N191);
buf BUF1 (N321, N319);
not NOT1 (N322, N320);
xor XOR2 (N323, N312, N266);
nand NAND3 (N324, N304, N251, N16);
xor XOR2 (N325, N324, N271);
and AND3 (N326, N323, N203, N56);
and AND3 (N327, N321, N181, N127);
nor NOR3 (N328, N303, N252, N150);
and AND3 (N329, N315, N137, N280);
nand NAND2 (N330, N329, N217);
or OR3 (N331, N325, N297, N131);
nor NOR4 (N332, N311, N251, N124, N131);
buf BUF1 (N333, N331);
not NOT1 (N334, N333);
buf BUF1 (N335, N332);
buf BUF1 (N336, N326);
nor NOR2 (N337, N336, N234);
nand NAND2 (N338, N317, N252);
xor XOR2 (N339, N322, N48);
buf BUF1 (N340, N334);
and AND4 (N341, N328, N200, N80, N124);
nand NAND2 (N342, N310, N193);
nor NOR3 (N343, N335, N228, N35);
buf BUF1 (N344, N313);
nand NAND4 (N345, N339, N210, N68, N122);
nor NOR2 (N346, N341, N65);
or OR4 (N347, N345, N271, N212, N277);
xor XOR2 (N348, N338, N249);
not NOT1 (N349, N347);
nor NOR3 (N350, N337, N77, N226);
nor NOR2 (N351, N344, N86);
nand NAND3 (N352, N348, N209, N93);
or OR2 (N353, N352, N298);
xor XOR2 (N354, N342, N201);
xor XOR2 (N355, N330, N113);
buf BUF1 (N356, N327);
buf BUF1 (N357, N340);
nor NOR3 (N358, N346, N242, N272);
and AND2 (N359, N358, N266);
nor NOR3 (N360, N349, N137, N296);
and AND3 (N361, N360, N134, N106);
xor XOR2 (N362, N343, N306);
or OR2 (N363, N357, N292);
xor XOR2 (N364, N362, N124);
not NOT1 (N365, N353);
nand NAND2 (N366, N350, N97);
xor XOR2 (N367, N364, N100);
nor NOR4 (N368, N366, N240, N268, N156);
buf BUF1 (N369, N365);
buf BUF1 (N370, N351);
or OR3 (N371, N368, N305, N189);
and AND4 (N372, N370, N14, N87, N87);
and AND2 (N373, N354, N127);
buf BUF1 (N374, N359);
nor NOR2 (N375, N369, N283);
not NOT1 (N376, N371);
and AND3 (N377, N373, N232, N119);
nand NAND3 (N378, N356, N65, N23);
or OR2 (N379, N367, N143);
and AND4 (N380, N363, N132, N225, N97);
and AND4 (N381, N355, N139, N286, N115);
xor XOR2 (N382, N372, N323);
nand NAND4 (N383, N380, N76, N10, N360);
and AND4 (N384, N383, N57, N202, N112);
not NOT1 (N385, N361);
xor XOR2 (N386, N375, N65);
or OR2 (N387, N378, N77);
nand NAND2 (N388, N374, N211);
or OR3 (N389, N377, N249, N74);
nand NAND4 (N390, N376, N131, N120, N164);
nor NOR4 (N391, N381, N348, N237, N164);
and AND4 (N392, N379, N16, N259, N285);
not NOT1 (N393, N390);
nand NAND4 (N394, N391, N274, N222, N268);
or OR4 (N395, N382, N180, N161, N165);
buf BUF1 (N396, N384);
nor NOR3 (N397, N385, N360, N15);
nand NAND3 (N398, N392, N115, N266);
nand NAND2 (N399, N393, N77);
not NOT1 (N400, N394);
xor XOR2 (N401, N399, N190);
nor NOR3 (N402, N400, N207, N241);
nor NOR4 (N403, N398, N207, N381, N85);
nor NOR3 (N404, N387, N100, N62);
buf BUF1 (N405, N403);
nor NOR3 (N406, N388, N337, N178);
buf BUF1 (N407, N402);
or OR2 (N408, N406, N91);
or OR3 (N409, N401, N155, N324);
nor NOR3 (N410, N396, N178, N130);
or OR3 (N411, N404, N63, N40);
nor NOR3 (N412, N410, N68, N297);
and AND4 (N413, N411, N236, N88, N38);
xor XOR2 (N414, N408, N257);
or OR3 (N415, N386, N400, N186);
xor XOR2 (N416, N415, N11);
and AND4 (N417, N416, N414, N101, N107);
not NOT1 (N418, N1);
nor NOR4 (N419, N389, N61, N384, N374);
or OR2 (N420, N418, N173);
nor NOR2 (N421, N409, N42);
xor XOR2 (N422, N412, N203);
nand NAND3 (N423, N422, N324, N238);
or OR3 (N424, N407, N210, N368);
not NOT1 (N425, N421);
and AND2 (N426, N405, N329);
nand NAND2 (N427, N417, N164);
and AND2 (N428, N424, N237);
buf BUF1 (N429, N419);
buf BUF1 (N430, N429);
xor XOR2 (N431, N430, N270);
buf BUF1 (N432, N420);
nand NAND2 (N433, N423, N369);
or OR4 (N434, N427, N45, N433, N100);
buf BUF1 (N435, N231);
xor XOR2 (N436, N432, N329);
and AND4 (N437, N425, N89, N140, N193);
nand NAND2 (N438, N437, N111);
and AND4 (N439, N397, N212, N432, N433);
or OR2 (N440, N438, N196);
and AND3 (N441, N395, N108, N45);
not NOT1 (N442, N426);
or OR4 (N443, N434, N5, N202, N150);
not NOT1 (N444, N435);
nor NOR4 (N445, N428, N433, N78, N339);
or OR3 (N446, N431, N379, N77);
or OR2 (N447, N442, N228);
not NOT1 (N448, N445);
not NOT1 (N449, N436);
nor NOR4 (N450, N439, N76, N382, N155);
nand NAND4 (N451, N450, N56, N441, N433);
or OR2 (N452, N430, N157);
not NOT1 (N453, N443);
buf BUF1 (N454, N444);
or OR4 (N455, N448, N145, N99, N129);
and AND2 (N456, N440, N169);
buf BUF1 (N457, N454);
nor NOR2 (N458, N447, N37);
or OR2 (N459, N451, N61);
xor XOR2 (N460, N452, N370);
buf BUF1 (N461, N455);
nand NAND3 (N462, N446, N73, N191);
buf BUF1 (N463, N453);
xor XOR2 (N464, N459, N319);
nand NAND2 (N465, N462, N87);
not NOT1 (N466, N464);
and AND3 (N467, N460, N275, N204);
xor XOR2 (N468, N413, N281);
and AND3 (N469, N461, N329, N109);
or OR4 (N470, N467, N4, N102, N296);
xor XOR2 (N471, N469, N24);
not NOT1 (N472, N465);
buf BUF1 (N473, N449);
xor XOR2 (N474, N466, N206);
nor NOR3 (N475, N473, N407, N257);
and AND3 (N476, N471, N236, N269);
nor NOR2 (N477, N468, N395);
xor XOR2 (N478, N463, N103);
buf BUF1 (N479, N476);
nand NAND4 (N480, N456, N67, N348, N375);
or OR2 (N481, N480, N219);
and AND4 (N482, N470, N191, N459, N407);
buf BUF1 (N483, N481);
xor XOR2 (N484, N475, N54);
buf BUF1 (N485, N479);
not NOT1 (N486, N484);
buf BUF1 (N487, N474);
or OR3 (N488, N483, N181, N434);
nor NOR3 (N489, N488, N385, N258);
or OR3 (N490, N482, N303, N401);
not NOT1 (N491, N487);
nor NOR3 (N492, N472, N392, N209);
xor XOR2 (N493, N489, N380);
nand NAND2 (N494, N490, N86);
xor XOR2 (N495, N478, N493);
nand NAND2 (N496, N180, N423);
not NOT1 (N497, N458);
and AND2 (N498, N477, N114);
not NOT1 (N499, N495);
nor NOR2 (N500, N491, N492);
and AND4 (N501, N438, N434, N110, N162);
xor XOR2 (N502, N500, N52);
or OR2 (N503, N494, N393);
xor XOR2 (N504, N485, N421);
xor XOR2 (N505, N486, N266);
nand NAND3 (N506, N504, N499, N111);
or OR4 (N507, N484, N291, N457, N504);
or OR2 (N508, N110, N51);
and AND3 (N509, N503, N185, N138);
nand NAND2 (N510, N509, N372);
nand NAND2 (N511, N505, N450);
nand NAND2 (N512, N498, N484);
nand NAND4 (N513, N512, N394, N129, N303);
and AND2 (N514, N501, N365);
xor XOR2 (N515, N496, N52);
and AND2 (N516, N511, N72);
xor XOR2 (N517, N516, N508);
buf BUF1 (N518, N103);
nor NOR4 (N519, N506, N56, N382, N458);
and AND4 (N520, N502, N236, N288, N402);
nor NOR2 (N521, N519, N97);
not NOT1 (N522, N518);
nor NOR3 (N523, N517, N338, N188);
or OR3 (N524, N523, N202, N124);
buf BUF1 (N525, N507);
buf BUF1 (N526, N522);
buf BUF1 (N527, N526);
xor XOR2 (N528, N513, N522);
and AND3 (N529, N514, N277, N453);
and AND4 (N530, N527, N200, N153, N206);
not NOT1 (N531, N530);
or OR4 (N532, N529, N285, N382, N365);
and AND2 (N533, N524, N355);
nand NAND3 (N534, N531, N255, N394);
xor XOR2 (N535, N515, N417);
not NOT1 (N536, N525);
buf BUF1 (N537, N534);
xor XOR2 (N538, N497, N217);
xor XOR2 (N539, N536, N301);
or OR4 (N540, N521, N471, N382, N447);
not NOT1 (N541, N539);
xor XOR2 (N542, N533, N333);
and AND3 (N543, N510, N2, N280);
nand NAND3 (N544, N542, N427, N126);
nand NAND4 (N545, N544, N268, N306, N63);
buf BUF1 (N546, N528);
and AND2 (N547, N546, N376);
buf BUF1 (N548, N543);
buf BUF1 (N549, N520);
nor NOR4 (N550, N537, N257, N328, N295);
and AND3 (N551, N541, N489, N130);
not NOT1 (N552, N551);
not NOT1 (N553, N535);
xor XOR2 (N554, N553, N539);
nand NAND4 (N555, N547, N369, N435, N93);
or OR2 (N556, N548, N207);
xor XOR2 (N557, N556, N101);
or OR2 (N558, N549, N223);
and AND2 (N559, N555, N358);
xor XOR2 (N560, N538, N458);
nor NOR4 (N561, N545, N171, N326, N514);
xor XOR2 (N562, N550, N147);
nand NAND2 (N563, N562, N493);
xor XOR2 (N564, N559, N165);
not NOT1 (N565, N564);
not NOT1 (N566, N563);
nor NOR4 (N567, N540, N415, N348, N222);
nor NOR4 (N568, N558, N262, N15, N131);
nand NAND4 (N569, N566, N26, N447, N272);
nand NAND4 (N570, N557, N505, N142, N221);
or OR4 (N571, N569, N44, N288, N229);
nand NAND3 (N572, N554, N399, N278);
or OR3 (N573, N568, N358, N193);
and AND2 (N574, N567, N127);
nor NOR4 (N575, N552, N167, N500, N503);
nand NAND4 (N576, N561, N19, N362, N271);
xor XOR2 (N577, N565, N228);
buf BUF1 (N578, N570);
not NOT1 (N579, N560);
nor NOR2 (N580, N577, N372);
buf BUF1 (N581, N573);
not NOT1 (N582, N581);
not NOT1 (N583, N532);
buf BUF1 (N584, N578);
xor XOR2 (N585, N575, N263);
nand NAND4 (N586, N582, N351, N119, N547);
not NOT1 (N587, N584);
nor NOR3 (N588, N571, N222, N498);
nand NAND2 (N589, N572, N496);
not NOT1 (N590, N586);
nor NOR2 (N591, N590, N581);
nor NOR3 (N592, N591, N108, N480);
or OR3 (N593, N589, N32, N229);
or OR3 (N594, N580, N261, N488);
nand NAND2 (N595, N592, N18);
and AND4 (N596, N579, N358, N570, N209);
or OR2 (N597, N583, N12);
xor XOR2 (N598, N597, N238);
nand NAND4 (N599, N594, N534, N89, N398);
buf BUF1 (N600, N598);
xor XOR2 (N601, N593, N341);
and AND2 (N602, N576, N78);
nor NOR4 (N603, N585, N7, N19, N469);
nor NOR3 (N604, N599, N132, N21);
not NOT1 (N605, N574);
xor XOR2 (N606, N602, N460);
or OR2 (N607, N596, N38);
buf BUF1 (N608, N595);
and AND2 (N609, N588, N38);
nor NOR3 (N610, N606, N171, N453);
xor XOR2 (N611, N601, N86);
xor XOR2 (N612, N611, N20);
or OR4 (N613, N587, N276, N586, N22);
and AND3 (N614, N609, N606, N269);
and AND4 (N615, N604, N30, N603, N117);
nor NOR2 (N616, N356, N115);
and AND3 (N617, N607, N95, N54);
xor XOR2 (N618, N615, N417);
buf BUF1 (N619, N617);
and AND2 (N620, N619, N587);
or OR3 (N621, N613, N545, N393);
xor XOR2 (N622, N612, N236);
buf BUF1 (N623, N618);
and AND3 (N624, N614, N32, N153);
not NOT1 (N625, N620);
nor NOR4 (N626, N624, N471, N356, N130);
not NOT1 (N627, N621);
nand NAND2 (N628, N616, N609);
and AND3 (N629, N623, N171, N32);
nand NAND2 (N630, N628, N117);
not NOT1 (N631, N630);
not NOT1 (N632, N625);
xor XOR2 (N633, N632, N323);
and AND3 (N634, N626, N513, N442);
and AND2 (N635, N608, N224);
and AND2 (N636, N605, N366);
xor XOR2 (N637, N635, N540);
or OR2 (N638, N627, N145);
nand NAND2 (N639, N637, N217);
and AND4 (N640, N639, N435, N510, N375);
xor XOR2 (N641, N638, N76);
not NOT1 (N642, N622);
or OR2 (N643, N631, N197);
xor XOR2 (N644, N640, N57);
buf BUF1 (N645, N634);
xor XOR2 (N646, N644, N233);
or OR3 (N647, N600, N209, N432);
xor XOR2 (N648, N642, N91);
nand NAND3 (N649, N641, N493, N161);
or OR4 (N650, N649, N488, N646, N420);
and AND2 (N651, N287, N619);
xor XOR2 (N652, N643, N548);
xor XOR2 (N653, N636, N609);
buf BUF1 (N654, N633);
nand NAND2 (N655, N650, N447);
nand NAND2 (N656, N629, N145);
and AND2 (N657, N655, N278);
or OR2 (N658, N651, N620);
and AND3 (N659, N653, N380, N434);
xor XOR2 (N660, N659, N427);
nor NOR3 (N661, N656, N180, N201);
nor NOR4 (N662, N647, N409, N440, N10);
nor NOR3 (N663, N661, N44, N602);
and AND4 (N664, N648, N539, N388, N517);
not NOT1 (N665, N645);
and AND3 (N666, N657, N144, N340);
and AND3 (N667, N666, N654, N581);
and AND3 (N668, N127, N241, N540);
and AND4 (N669, N662, N555, N630, N388);
and AND4 (N670, N669, N568, N403, N368);
not NOT1 (N671, N664);
nand NAND2 (N672, N658, N570);
xor XOR2 (N673, N668, N356);
xor XOR2 (N674, N665, N669);
or OR2 (N675, N663, N657);
nand NAND4 (N676, N610, N166, N276, N185);
nand NAND4 (N677, N674, N379, N91, N345);
and AND2 (N678, N677, N347);
not NOT1 (N679, N671);
nand NAND4 (N680, N679, N8, N514, N81);
not NOT1 (N681, N672);
xor XOR2 (N682, N676, N49);
nand NAND3 (N683, N678, N287, N31);
not NOT1 (N684, N682);
xor XOR2 (N685, N681, N116);
buf BUF1 (N686, N652);
buf BUF1 (N687, N667);
buf BUF1 (N688, N683);
nand NAND4 (N689, N660, N304, N402, N253);
buf BUF1 (N690, N688);
nor NOR3 (N691, N673, N47, N132);
and AND4 (N692, N686, N614, N555, N496);
buf BUF1 (N693, N684);
nor NOR2 (N694, N670, N158);
nor NOR2 (N695, N689, N315);
buf BUF1 (N696, N694);
and AND3 (N697, N680, N356, N646);
buf BUF1 (N698, N695);
nand NAND3 (N699, N685, N642, N692);
or OR2 (N700, N609, N124);
or OR3 (N701, N687, N184, N192);
xor XOR2 (N702, N697, N645);
nand NAND4 (N703, N701, N162, N512, N147);
not NOT1 (N704, N700);
nor NOR3 (N705, N698, N355, N12);
not NOT1 (N706, N675);
buf BUF1 (N707, N693);
not NOT1 (N708, N706);
not NOT1 (N709, N702);
nor NOR4 (N710, N703, N420, N664, N424);
not NOT1 (N711, N699);
and AND2 (N712, N691, N619);
and AND3 (N713, N705, N119, N256);
or OR2 (N714, N712, N303);
nand NAND4 (N715, N709, N293, N95, N290);
buf BUF1 (N716, N707);
not NOT1 (N717, N704);
or OR3 (N718, N716, N682, N566);
and AND2 (N719, N718, N13);
and AND2 (N720, N715, N452);
buf BUF1 (N721, N713);
nor NOR4 (N722, N711, N221, N134, N315);
buf BUF1 (N723, N721);
xor XOR2 (N724, N719, N419);
buf BUF1 (N725, N723);
buf BUF1 (N726, N717);
not NOT1 (N727, N696);
and AND4 (N728, N725, N298, N592, N476);
xor XOR2 (N729, N722, N295);
and AND4 (N730, N728, N590, N406, N439);
xor XOR2 (N731, N727, N19);
buf BUF1 (N732, N720);
nand NAND2 (N733, N730, N370);
not NOT1 (N734, N732);
not NOT1 (N735, N731);
buf BUF1 (N736, N726);
nor NOR4 (N737, N690, N377, N560, N99);
nand NAND3 (N738, N737, N670, N491);
nor NOR2 (N739, N710, N214);
nor NOR4 (N740, N739, N316, N588, N283);
or OR2 (N741, N735, N240);
nor NOR2 (N742, N729, N134);
buf BUF1 (N743, N742);
nor NOR3 (N744, N714, N427, N85);
nor NOR2 (N745, N733, N194);
or OR3 (N746, N741, N557, N471);
buf BUF1 (N747, N734);
and AND4 (N748, N724, N134, N63, N668);
xor XOR2 (N749, N744, N3);
xor XOR2 (N750, N748, N111);
or OR4 (N751, N746, N660, N428, N715);
not NOT1 (N752, N749);
xor XOR2 (N753, N740, N312);
or OR3 (N754, N750, N363, N427);
not NOT1 (N755, N753);
xor XOR2 (N756, N708, N389);
and AND4 (N757, N743, N571, N447, N280);
and AND2 (N758, N736, N710);
buf BUF1 (N759, N755);
nand NAND3 (N760, N759, N474, N142);
nor NOR3 (N761, N756, N256, N355);
buf BUF1 (N762, N745);
nor NOR4 (N763, N761, N493, N753, N59);
xor XOR2 (N764, N752, N544);
not NOT1 (N765, N757);
xor XOR2 (N766, N758, N465);
xor XOR2 (N767, N754, N117);
and AND4 (N768, N738, N419, N644, N95);
buf BUF1 (N769, N763);
not NOT1 (N770, N760);
not NOT1 (N771, N770);
or OR3 (N772, N766, N171, N493);
and AND2 (N773, N768, N72);
nor NOR4 (N774, N772, N725, N191, N98);
or OR3 (N775, N751, N585, N552);
nor NOR4 (N776, N764, N729, N590, N421);
and AND3 (N777, N747, N304, N684);
nand NAND2 (N778, N769, N232);
not NOT1 (N779, N778);
and AND4 (N780, N771, N134, N45, N20);
xor XOR2 (N781, N780, N302);
nor NOR2 (N782, N779, N761);
and AND2 (N783, N781, N255);
xor XOR2 (N784, N773, N311);
xor XOR2 (N785, N776, N343);
not NOT1 (N786, N783);
and AND4 (N787, N765, N56, N195, N619);
xor XOR2 (N788, N767, N321);
buf BUF1 (N789, N762);
nor NOR3 (N790, N782, N261, N570);
not NOT1 (N791, N788);
nor NOR3 (N792, N791, N56, N34);
nand NAND4 (N793, N784, N425, N76, N146);
or OR4 (N794, N775, N58, N501, N125);
xor XOR2 (N795, N793, N487);
or OR2 (N796, N789, N184);
and AND3 (N797, N786, N757, N328);
buf BUF1 (N798, N792);
nor NOR2 (N799, N795, N147);
buf BUF1 (N800, N785);
not NOT1 (N801, N787);
nor NOR2 (N802, N798, N477);
not NOT1 (N803, N802);
not NOT1 (N804, N777);
and AND3 (N805, N801, N73, N527);
nand NAND2 (N806, N790, N657);
and AND2 (N807, N794, N539);
or OR2 (N808, N797, N261);
nand NAND4 (N809, N799, N50, N20, N184);
not NOT1 (N810, N800);
buf BUF1 (N811, N804);
or OR4 (N812, N809, N719, N104, N302);
nor NOR4 (N813, N803, N193, N662, N614);
nand NAND2 (N814, N813, N642);
or OR4 (N815, N774, N444, N26, N387);
endmodule