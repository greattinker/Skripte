// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11;

output N1510,N1470,N1503,N1506,N1502,N1508,N1509,N1497,N1504,N1511;

not NOT1 (N12, N3);
xor XOR2 (N13, N8, N11);
buf BUF1 (N14, N7);
not NOT1 (N15, N1);
nor NOR3 (N16, N14, N2, N3);
or OR3 (N17, N2, N9, N13);
not NOT1 (N18, N14);
and AND4 (N19, N13, N9, N5, N11);
xor XOR2 (N20, N6, N5);
and AND3 (N21, N13, N16, N17);
nor NOR3 (N22, N4, N3, N15);
buf BUF1 (N23, N21);
or OR3 (N24, N21, N16, N23);
or OR3 (N25, N12, N14, N24);
or OR2 (N26, N18, N9);
and AND2 (N27, N6, N10);
not NOT1 (N28, N13);
and AND2 (N29, N5, N16);
buf BUF1 (N30, N22);
xor XOR2 (N31, N3, N7);
not NOT1 (N32, N12);
buf BUF1 (N33, N31);
and AND4 (N34, N29, N18, N30, N1);
nor NOR4 (N35, N22, N32, N1, N20);
xor XOR2 (N36, N20, N31);
nor NOR4 (N37, N21, N34, N21, N15);
or OR2 (N38, N21, N23);
xor XOR2 (N39, N27, N28);
buf BUF1 (N40, N33);
nor NOR2 (N41, N32, N1);
and AND3 (N42, N19, N27, N18);
nand NAND2 (N43, N41, N39);
buf BUF1 (N44, N5);
nor NOR4 (N45, N36, N35, N39, N25);
nand NAND2 (N46, N7, N27);
or OR2 (N47, N32, N8);
not NOT1 (N48, N38);
xor XOR2 (N49, N48, N30);
nor NOR3 (N50, N42, N46, N5);
xor XOR2 (N51, N18, N31);
nor NOR2 (N52, N49, N38);
not NOT1 (N53, N26);
xor XOR2 (N54, N43, N40);
not NOT1 (N55, N49);
xor XOR2 (N56, N54, N53);
nand NAND2 (N57, N48, N2);
not NOT1 (N58, N44);
nand NAND2 (N59, N37, N1);
nand NAND2 (N60, N51, N53);
nor NOR2 (N61, N45, N54);
nor NOR3 (N62, N50, N11, N6);
not NOT1 (N63, N61);
xor XOR2 (N64, N47, N41);
nor NOR2 (N65, N64, N61);
or OR3 (N66, N57, N35, N50);
and AND4 (N67, N62, N64, N57, N4);
xor XOR2 (N68, N55, N37);
nor NOR2 (N69, N58, N58);
nor NOR4 (N70, N59, N50, N55, N62);
buf BUF1 (N71, N56);
or OR3 (N72, N69, N10, N20);
and AND3 (N73, N71, N16, N17);
and AND3 (N74, N73, N38, N1);
xor XOR2 (N75, N66, N34);
nor NOR4 (N76, N60, N21, N43, N58);
not NOT1 (N77, N52);
and AND4 (N78, N76, N7, N73, N60);
and AND4 (N79, N74, N64, N68, N68);
nand NAND2 (N80, N74, N61);
nand NAND2 (N81, N72, N43);
not NOT1 (N82, N67);
and AND3 (N83, N78, N52, N79);
and AND4 (N84, N78, N37, N19, N32);
and AND3 (N85, N77, N73, N37);
nand NAND3 (N86, N83, N6, N44);
not NOT1 (N87, N63);
or OR2 (N88, N81, N2);
and AND2 (N89, N88, N7);
not NOT1 (N90, N85);
and AND2 (N91, N75, N63);
not NOT1 (N92, N82);
nor NOR3 (N93, N87, N53, N72);
or OR4 (N94, N80, N29, N22, N22);
nand NAND3 (N95, N70, N20, N91);
buf BUF1 (N96, N41);
or OR3 (N97, N93, N82, N58);
or OR4 (N98, N97, N9, N3, N91);
nand NAND2 (N99, N86, N75);
not NOT1 (N100, N92);
nand NAND2 (N101, N95, N3);
nor NOR3 (N102, N84, N45, N100);
or OR4 (N103, N75, N21, N71, N57);
not NOT1 (N104, N96);
and AND2 (N105, N103, N99);
buf BUF1 (N106, N72);
nand NAND3 (N107, N94, N73, N84);
nand NAND3 (N108, N107, N40, N100);
or OR4 (N109, N104, N49, N25, N103);
nor NOR4 (N110, N90, N52, N54, N92);
nand NAND3 (N111, N106, N82, N36);
nand NAND4 (N112, N98, N87, N6, N2);
or OR3 (N113, N102, N79, N86);
nor NOR2 (N114, N109, N88);
xor XOR2 (N115, N111, N96);
nor NOR3 (N116, N108, N27, N52);
nor NOR3 (N117, N116, N23, N71);
not NOT1 (N118, N65);
nor NOR4 (N119, N112, N14, N24, N92);
or OR3 (N120, N119, N75, N76);
or OR4 (N121, N110, N96, N37, N117);
or OR4 (N122, N68, N95, N106, N80);
and AND2 (N123, N113, N92);
nand NAND3 (N124, N120, N81, N39);
buf BUF1 (N125, N101);
or OR4 (N126, N89, N97, N51, N42);
or OR3 (N127, N105, N76, N18);
and AND3 (N128, N114, N119, N23);
nor NOR3 (N129, N128, N128, N122);
and AND4 (N130, N101, N106, N29, N36);
nor NOR3 (N131, N121, N41, N18);
xor XOR2 (N132, N123, N107);
and AND3 (N133, N125, N25, N56);
xor XOR2 (N134, N131, N66);
xor XOR2 (N135, N134, N78);
buf BUF1 (N136, N115);
or OR4 (N137, N124, N133, N111, N57);
xor XOR2 (N138, N117, N32);
xor XOR2 (N139, N138, N123);
nand NAND4 (N140, N130, N43, N75, N76);
and AND4 (N141, N136, N46, N61, N21);
or OR4 (N142, N129, N87, N60, N118);
nor NOR3 (N143, N61, N80, N57);
xor XOR2 (N144, N137, N117);
nor NOR2 (N145, N139, N57);
or OR3 (N146, N140, N137, N139);
xor XOR2 (N147, N143, N118);
xor XOR2 (N148, N127, N27);
or OR3 (N149, N142, N145, N47);
not NOT1 (N150, N54);
nand NAND4 (N151, N132, N107, N23, N110);
not NOT1 (N152, N126);
nor NOR3 (N153, N141, N6, N148);
nand NAND4 (N154, N33, N43, N81, N24);
nand NAND4 (N155, N149, N132, N9, N29);
buf BUF1 (N156, N147);
or OR2 (N157, N153, N78);
xor XOR2 (N158, N155, N40);
not NOT1 (N159, N144);
nor NOR3 (N160, N146, N145, N123);
nand NAND4 (N161, N157, N41, N66, N159);
nand NAND3 (N162, N94, N53, N155);
nor NOR2 (N163, N161, N141);
buf BUF1 (N164, N154);
nand NAND4 (N165, N156, N82, N46, N64);
nand NAND3 (N166, N165, N18, N77);
not NOT1 (N167, N152);
xor XOR2 (N168, N160, N147);
buf BUF1 (N169, N151);
nand NAND4 (N170, N166, N137, N143, N7);
xor XOR2 (N171, N169, N65);
nand NAND3 (N172, N164, N62, N12);
or OR3 (N173, N163, N66, N161);
not NOT1 (N174, N170);
not NOT1 (N175, N135);
or OR4 (N176, N167, N171, N96, N132);
or OR2 (N177, N89, N119);
not NOT1 (N178, N162);
or OR4 (N179, N150, N149, N4, N110);
nor NOR3 (N180, N158, N144, N62);
nand NAND2 (N181, N177, N22);
buf BUF1 (N182, N175);
and AND4 (N183, N168, N126, N23, N64);
buf BUF1 (N184, N172);
nor NOR2 (N185, N181, N111);
nand NAND4 (N186, N176, N107, N169, N13);
xor XOR2 (N187, N183, N71);
and AND2 (N188, N185, N149);
buf BUF1 (N189, N178);
not NOT1 (N190, N173);
buf BUF1 (N191, N180);
nand NAND4 (N192, N186, N107, N55, N118);
or OR4 (N193, N191, N168, N116, N112);
nand NAND2 (N194, N188, N103);
nor NOR3 (N195, N184, N121, N72);
buf BUF1 (N196, N182);
nand NAND2 (N197, N194, N111);
not NOT1 (N198, N174);
nor NOR2 (N199, N189, N176);
buf BUF1 (N200, N190);
or OR2 (N201, N200, N18);
xor XOR2 (N202, N179, N70);
and AND2 (N203, N196, N164);
or OR2 (N204, N187, N137);
xor XOR2 (N205, N195, N79);
nand NAND3 (N206, N203, N44, N126);
and AND2 (N207, N204, N129);
nand NAND2 (N208, N192, N110);
nand NAND2 (N209, N207, N144);
xor XOR2 (N210, N201, N125);
buf BUF1 (N211, N202);
buf BUF1 (N212, N211);
not NOT1 (N213, N209);
xor XOR2 (N214, N212, N33);
nand NAND4 (N215, N213, N46, N34, N102);
or OR2 (N216, N193, N64);
and AND3 (N217, N208, N12, N63);
buf BUF1 (N218, N197);
nand NAND4 (N219, N218, N68, N120, N72);
not NOT1 (N220, N198);
and AND2 (N221, N217, N170);
xor XOR2 (N222, N199, N191);
not NOT1 (N223, N220);
buf BUF1 (N224, N215);
nor NOR4 (N225, N214, N177, N182, N22);
xor XOR2 (N226, N225, N198);
and AND3 (N227, N224, N81, N58);
or OR2 (N228, N223, N19);
nor NOR4 (N229, N222, N169, N104, N37);
xor XOR2 (N230, N210, N73);
nor NOR2 (N231, N226, N132);
xor XOR2 (N232, N230, N210);
xor XOR2 (N233, N219, N113);
and AND4 (N234, N229, N189, N174, N76);
or OR3 (N235, N227, N140, N98);
xor XOR2 (N236, N206, N118);
and AND4 (N237, N233, N22, N112, N103);
not NOT1 (N238, N216);
nor NOR4 (N239, N221, N97, N41, N191);
xor XOR2 (N240, N234, N53);
xor XOR2 (N241, N236, N137);
not NOT1 (N242, N235);
not NOT1 (N243, N205);
nor NOR2 (N244, N232, N71);
buf BUF1 (N245, N244);
and AND3 (N246, N242, N158, N138);
nand NAND3 (N247, N241, N245, N66);
not NOT1 (N248, N104);
buf BUF1 (N249, N248);
or OR3 (N250, N231, N185, N67);
buf BUF1 (N251, N243);
or OR2 (N252, N239, N242);
nor NOR2 (N253, N240, N3);
and AND4 (N254, N250, N137, N68, N48);
buf BUF1 (N255, N237);
buf BUF1 (N256, N255);
xor XOR2 (N257, N256, N179);
buf BUF1 (N258, N228);
or OR2 (N259, N247, N63);
xor XOR2 (N260, N252, N105);
and AND3 (N261, N257, N31, N113);
and AND4 (N262, N258, N148, N174, N121);
nor NOR3 (N263, N238, N127, N169);
nor NOR4 (N264, N260, N139, N166, N77);
xor XOR2 (N265, N249, N71);
and AND2 (N266, N253, N229);
and AND2 (N267, N264, N10);
nand NAND2 (N268, N254, N47);
not NOT1 (N269, N268);
nand NAND4 (N270, N246, N212, N269, N42);
nor NOR4 (N271, N186, N146, N266, N9);
xor XOR2 (N272, N8, N56);
nor NOR4 (N273, N271, N183, N53, N178);
not NOT1 (N274, N262);
buf BUF1 (N275, N265);
not NOT1 (N276, N259);
nand NAND4 (N277, N272, N161, N253, N135);
and AND4 (N278, N261, N34, N160, N107);
xor XOR2 (N279, N267, N170);
nor NOR4 (N280, N270, N94, N78, N146);
buf BUF1 (N281, N279);
nand NAND2 (N282, N274, N88);
not NOT1 (N283, N281);
and AND3 (N284, N277, N66, N38);
nor NOR2 (N285, N263, N259);
nand NAND4 (N286, N273, N87, N222, N89);
xor XOR2 (N287, N280, N257);
xor XOR2 (N288, N284, N249);
buf BUF1 (N289, N283);
nor NOR2 (N290, N285, N65);
nand NAND2 (N291, N290, N82);
buf BUF1 (N292, N291);
nor NOR4 (N293, N282, N96, N287, N76);
xor XOR2 (N294, N64, N245);
nand NAND3 (N295, N286, N165, N27);
nor NOR3 (N296, N293, N67, N98);
and AND3 (N297, N296, N142, N36);
buf BUF1 (N298, N278);
or OR3 (N299, N275, N150, N219);
and AND2 (N300, N299, N209);
nand NAND4 (N301, N251, N209, N294, N36);
buf BUF1 (N302, N271);
and AND3 (N303, N295, N228, N179);
not NOT1 (N304, N301);
and AND3 (N305, N289, N221, N154);
nor NOR4 (N306, N302, N48, N87, N118);
buf BUF1 (N307, N306);
or OR3 (N308, N303, N147, N139);
or OR3 (N309, N308, N220, N44);
buf BUF1 (N310, N297);
xor XOR2 (N311, N310, N95);
nand NAND2 (N312, N298, N78);
or OR3 (N313, N276, N242, N63);
nand NAND4 (N314, N307, N227, N49, N124);
and AND4 (N315, N300, N43, N57, N123);
nand NAND3 (N316, N312, N127, N166);
and AND3 (N317, N305, N1, N80);
not NOT1 (N318, N317);
xor XOR2 (N319, N288, N161);
not NOT1 (N320, N292);
nor NOR4 (N321, N319, N43, N115, N294);
not NOT1 (N322, N304);
or OR3 (N323, N314, N91, N259);
nor NOR4 (N324, N318, N162, N173, N216);
xor XOR2 (N325, N324, N206);
buf BUF1 (N326, N311);
or OR3 (N327, N321, N298, N297);
nor NOR2 (N328, N327, N113);
not NOT1 (N329, N315);
nor NOR2 (N330, N322, N6);
and AND2 (N331, N329, N20);
buf BUF1 (N332, N331);
buf BUF1 (N333, N323);
nor NOR3 (N334, N313, N320, N282);
nor NOR2 (N335, N241, N108);
not NOT1 (N336, N330);
nor NOR2 (N337, N309, N69);
and AND4 (N338, N326, N334, N111, N15);
or OR4 (N339, N75, N242, N7, N110);
nand NAND2 (N340, N338, N79);
xor XOR2 (N341, N332, N5);
xor XOR2 (N342, N340, N149);
buf BUF1 (N343, N342);
xor XOR2 (N344, N343, N81);
nor NOR4 (N345, N328, N221, N313, N293);
not NOT1 (N346, N341);
or OR2 (N347, N344, N115);
not NOT1 (N348, N333);
buf BUF1 (N349, N336);
nor NOR3 (N350, N347, N285, N281);
buf BUF1 (N351, N316);
or OR4 (N352, N350, N178, N157, N315);
buf BUF1 (N353, N345);
xor XOR2 (N354, N346, N18);
not NOT1 (N355, N352);
nand NAND4 (N356, N351, N321, N260, N54);
and AND2 (N357, N348, N307);
xor XOR2 (N358, N356, N277);
nand NAND4 (N359, N353, N79, N171, N318);
nor NOR2 (N360, N337, N184);
or OR3 (N361, N339, N208, N156);
nor NOR3 (N362, N355, N192, N146);
xor XOR2 (N363, N349, N180);
nor NOR2 (N364, N359, N46);
xor XOR2 (N365, N358, N217);
and AND2 (N366, N335, N325);
not NOT1 (N367, N152);
nor NOR2 (N368, N363, N41);
not NOT1 (N369, N354);
and AND3 (N370, N365, N154, N340);
nor NOR4 (N371, N370, N106, N60, N321);
xor XOR2 (N372, N368, N11);
not NOT1 (N373, N366);
not NOT1 (N374, N362);
nor NOR4 (N375, N364, N32, N64, N69);
buf BUF1 (N376, N372);
xor XOR2 (N377, N375, N92);
and AND3 (N378, N369, N146, N104);
nor NOR3 (N379, N371, N336, N236);
buf BUF1 (N380, N379);
nand NAND4 (N381, N357, N226, N100, N126);
and AND4 (N382, N380, N100, N171, N199);
or OR4 (N383, N367, N175, N167, N373);
and AND2 (N384, N142, N180);
or OR2 (N385, N377, N15);
and AND3 (N386, N378, N50, N130);
or OR4 (N387, N381, N80, N79, N261);
and AND4 (N388, N361, N360, N229, N238);
and AND2 (N389, N241, N65);
nor NOR4 (N390, N376, N127, N299, N129);
not NOT1 (N391, N388);
nor NOR4 (N392, N391, N46, N382, N375);
xor XOR2 (N393, N135, N322);
or OR4 (N394, N385, N382, N42, N89);
or OR2 (N395, N384, N163);
and AND3 (N396, N393, N337, N116);
not NOT1 (N397, N392);
not NOT1 (N398, N394);
not NOT1 (N399, N374);
xor XOR2 (N400, N395, N230);
nand NAND2 (N401, N399, N208);
not NOT1 (N402, N398);
buf BUF1 (N403, N401);
xor XOR2 (N404, N400, N170);
or OR2 (N405, N397, N129);
or OR4 (N406, N405, N230, N325, N395);
or OR2 (N407, N404, N60);
buf BUF1 (N408, N407);
xor XOR2 (N409, N390, N344);
buf BUF1 (N410, N389);
not NOT1 (N411, N396);
nor NOR3 (N412, N408, N409, N330);
not NOT1 (N413, N144);
buf BUF1 (N414, N411);
and AND4 (N415, N403, N48, N327, N150);
not NOT1 (N416, N410);
or OR4 (N417, N386, N49, N181, N314);
not NOT1 (N418, N417);
buf BUF1 (N419, N415);
and AND2 (N420, N406, N211);
and AND3 (N421, N414, N57, N267);
xor XOR2 (N422, N420, N340);
not NOT1 (N423, N402);
nand NAND4 (N424, N413, N59, N327, N126);
buf BUF1 (N425, N423);
buf BUF1 (N426, N412);
xor XOR2 (N427, N419, N345);
or OR3 (N428, N421, N123, N410);
or OR4 (N429, N428, N232, N81, N61);
or OR3 (N430, N429, N280, N339);
nor NOR2 (N431, N430, N358);
nor NOR3 (N432, N426, N54, N355);
xor XOR2 (N433, N387, N295);
buf BUF1 (N434, N424);
nand NAND4 (N435, N383, N276, N337, N47);
xor XOR2 (N436, N425, N207);
nand NAND4 (N437, N418, N257, N348, N174);
or OR4 (N438, N432, N383, N298, N142);
nand NAND2 (N439, N435, N92);
buf BUF1 (N440, N436);
nand NAND3 (N441, N440, N141, N316);
xor XOR2 (N442, N437, N371);
not NOT1 (N443, N422);
buf BUF1 (N444, N427);
nand NAND2 (N445, N443, N290);
nand NAND2 (N446, N431, N233);
nor NOR3 (N447, N416, N221, N154);
nand NAND2 (N448, N439, N138);
and AND3 (N449, N448, N364, N302);
buf BUF1 (N450, N449);
or OR3 (N451, N434, N223, N163);
nand NAND3 (N452, N442, N279, N105);
and AND4 (N453, N444, N402, N380, N170);
nor NOR3 (N454, N433, N436, N254);
xor XOR2 (N455, N441, N209);
xor XOR2 (N456, N447, N268);
or OR3 (N457, N445, N344, N62);
or OR3 (N458, N451, N211, N426);
xor XOR2 (N459, N452, N378);
nor NOR4 (N460, N458, N186, N215, N367);
buf BUF1 (N461, N453);
or OR2 (N462, N450, N426);
xor XOR2 (N463, N461, N66);
and AND3 (N464, N454, N243, N372);
or OR2 (N465, N446, N414);
buf BUF1 (N466, N459);
not NOT1 (N467, N455);
xor XOR2 (N468, N457, N193);
or OR2 (N469, N466, N155);
xor XOR2 (N470, N465, N408);
nor NOR3 (N471, N462, N37, N191);
nand NAND4 (N472, N471, N145, N382, N396);
and AND2 (N473, N472, N131);
xor XOR2 (N474, N467, N271);
not NOT1 (N475, N469);
nor NOR2 (N476, N456, N433);
or OR3 (N477, N470, N84, N276);
and AND4 (N478, N477, N88, N26, N111);
nand NAND4 (N479, N476, N153, N232, N117);
xor XOR2 (N480, N474, N122);
and AND3 (N481, N475, N382, N438);
not NOT1 (N482, N202);
not NOT1 (N483, N482);
not NOT1 (N484, N479);
not NOT1 (N485, N460);
and AND3 (N486, N473, N282, N37);
xor XOR2 (N487, N478, N158);
not NOT1 (N488, N487);
buf BUF1 (N489, N488);
not NOT1 (N490, N481);
not NOT1 (N491, N486);
not NOT1 (N492, N464);
and AND3 (N493, N484, N292, N275);
and AND3 (N494, N491, N430, N205);
buf BUF1 (N495, N468);
not NOT1 (N496, N490);
xor XOR2 (N497, N495, N464);
and AND3 (N498, N480, N322, N444);
nor NOR2 (N499, N494, N280);
and AND2 (N500, N492, N379);
nor NOR4 (N501, N496, N386, N498, N420);
nand NAND3 (N502, N239, N175, N363);
nor NOR2 (N503, N463, N124);
or OR4 (N504, N483, N368, N103, N275);
buf BUF1 (N505, N485);
or OR3 (N506, N493, N293, N1);
buf BUF1 (N507, N506);
buf BUF1 (N508, N499);
xor XOR2 (N509, N504, N247);
and AND2 (N510, N497, N145);
and AND4 (N511, N500, N249, N95, N113);
buf BUF1 (N512, N503);
not NOT1 (N513, N507);
buf BUF1 (N514, N505);
nand NAND4 (N515, N508, N250, N457, N513);
buf BUF1 (N516, N157);
nand NAND2 (N517, N501, N11);
buf BUF1 (N518, N510);
buf BUF1 (N519, N489);
nor NOR3 (N520, N518, N389, N359);
xor XOR2 (N521, N519, N62);
xor XOR2 (N522, N515, N344);
xor XOR2 (N523, N517, N166);
or OR2 (N524, N523, N193);
or OR4 (N525, N522, N385, N428, N178);
nor NOR4 (N526, N514, N395, N65, N288);
nand NAND3 (N527, N526, N297, N138);
not NOT1 (N528, N502);
nor NOR2 (N529, N525, N261);
nand NAND4 (N530, N521, N52, N419, N41);
nor NOR4 (N531, N516, N349, N251, N60);
xor XOR2 (N532, N528, N367);
or OR3 (N533, N512, N429, N210);
or OR4 (N534, N529, N68, N162, N516);
buf BUF1 (N535, N530);
nor NOR4 (N536, N509, N320, N522, N421);
not NOT1 (N537, N533);
nor NOR3 (N538, N534, N95, N130);
xor XOR2 (N539, N535, N16);
or OR4 (N540, N539, N130, N52, N399);
and AND2 (N541, N531, N158);
xor XOR2 (N542, N540, N527);
or OR3 (N543, N410, N226, N445);
nor NOR3 (N544, N538, N69, N51);
or OR2 (N545, N511, N229);
or OR3 (N546, N537, N173, N168);
buf BUF1 (N547, N543);
and AND2 (N548, N541, N405);
nand NAND4 (N549, N520, N101, N100, N69);
not NOT1 (N550, N536);
and AND4 (N551, N542, N533, N81, N365);
or OR3 (N552, N551, N132, N492);
and AND3 (N553, N547, N20, N21);
buf BUF1 (N554, N524);
xor XOR2 (N555, N546, N81);
buf BUF1 (N556, N554);
and AND2 (N557, N548, N407);
nor NOR3 (N558, N553, N29, N254);
nand NAND3 (N559, N544, N429, N340);
xor XOR2 (N560, N558, N179);
or OR4 (N561, N555, N345, N512, N556);
and AND3 (N562, N382, N368, N424);
nor NOR2 (N563, N549, N509);
xor XOR2 (N564, N563, N560);
xor XOR2 (N565, N405, N241);
xor XOR2 (N566, N557, N539);
nand NAND4 (N567, N562, N346, N229, N276);
nand NAND2 (N568, N564, N289);
nand NAND3 (N569, N545, N355, N64);
not NOT1 (N570, N565);
nand NAND2 (N571, N561, N512);
not NOT1 (N572, N532);
or OR3 (N573, N566, N416, N444);
nand NAND3 (N574, N571, N280, N417);
xor XOR2 (N575, N552, N419);
not NOT1 (N576, N559);
or OR2 (N577, N574, N425);
not NOT1 (N578, N567);
buf BUF1 (N579, N573);
not NOT1 (N580, N577);
and AND2 (N581, N550, N249);
or OR4 (N582, N570, N412, N223, N225);
and AND4 (N583, N568, N43, N96, N342);
nor NOR2 (N584, N575, N485);
nand NAND3 (N585, N569, N248, N399);
nor NOR2 (N586, N580, N266);
buf BUF1 (N587, N586);
nor NOR3 (N588, N578, N299, N203);
xor XOR2 (N589, N588, N256);
buf BUF1 (N590, N589);
nor NOR3 (N591, N581, N1, N34);
nand NAND2 (N592, N576, N295);
or OR4 (N593, N582, N119, N340, N142);
buf BUF1 (N594, N592);
nand NAND3 (N595, N584, N486, N80);
xor XOR2 (N596, N585, N214);
or OR3 (N597, N591, N321, N334);
nand NAND3 (N598, N597, N212, N141);
not NOT1 (N599, N598);
and AND4 (N600, N593, N491, N340, N595);
and AND3 (N601, N461, N498, N102);
buf BUF1 (N602, N601);
or OR3 (N603, N587, N217, N249);
nand NAND3 (N604, N600, N539, N54);
nor NOR4 (N605, N594, N362, N62, N581);
not NOT1 (N606, N602);
nor NOR4 (N607, N605, N225, N202, N468);
and AND3 (N608, N572, N453, N224);
not NOT1 (N609, N604);
or OR2 (N610, N607, N30);
or OR3 (N611, N603, N242, N362);
and AND4 (N612, N599, N324, N169, N591);
nand NAND3 (N613, N590, N131, N282);
buf BUF1 (N614, N610);
nand NAND2 (N615, N596, N175);
buf BUF1 (N616, N611);
xor XOR2 (N617, N615, N603);
xor XOR2 (N618, N617, N78);
xor XOR2 (N619, N616, N39);
or OR3 (N620, N606, N208, N577);
not NOT1 (N621, N612);
buf BUF1 (N622, N620);
nand NAND2 (N623, N583, N193);
not NOT1 (N624, N579);
or OR2 (N625, N619, N149);
buf BUF1 (N626, N623);
or OR4 (N627, N624, N6, N533, N308);
not NOT1 (N628, N618);
xor XOR2 (N629, N613, N465);
nand NAND3 (N630, N627, N205, N115);
not NOT1 (N631, N625);
xor XOR2 (N632, N621, N391);
or OR4 (N633, N608, N256, N376, N446);
xor XOR2 (N634, N629, N599);
nand NAND3 (N635, N634, N495, N517);
nor NOR2 (N636, N635, N590);
not NOT1 (N637, N626);
nor NOR3 (N638, N609, N129, N40);
nand NAND4 (N639, N638, N29, N36, N185);
not NOT1 (N640, N632);
and AND4 (N641, N622, N589, N246, N507);
xor XOR2 (N642, N614, N325);
buf BUF1 (N643, N639);
not NOT1 (N644, N636);
nand NAND2 (N645, N631, N441);
or OR4 (N646, N630, N396, N534, N638);
nor NOR3 (N647, N645, N489, N134);
and AND2 (N648, N647, N106);
and AND3 (N649, N641, N250, N63);
and AND2 (N650, N646, N266);
xor XOR2 (N651, N642, N270);
nand NAND3 (N652, N650, N383, N98);
and AND4 (N653, N651, N525, N147, N134);
nand NAND4 (N654, N648, N554, N496, N457);
nor NOR3 (N655, N644, N527, N349);
nor NOR2 (N656, N653, N128);
not NOT1 (N657, N654);
xor XOR2 (N658, N649, N501);
or OR4 (N659, N628, N485, N583, N623);
and AND2 (N660, N643, N358);
not NOT1 (N661, N655);
not NOT1 (N662, N660);
or OR2 (N663, N656, N307);
nor NOR3 (N664, N659, N403, N276);
buf BUF1 (N665, N663);
xor XOR2 (N666, N658, N661);
not NOT1 (N667, N250);
nand NAND4 (N668, N633, N477, N113, N494);
nor NOR3 (N669, N657, N560, N197);
xor XOR2 (N670, N640, N373);
not NOT1 (N671, N667);
not NOT1 (N672, N662);
or OR4 (N673, N665, N360, N429, N169);
buf BUF1 (N674, N666);
or OR3 (N675, N668, N455, N134);
nor NOR3 (N676, N637, N105, N32);
nand NAND3 (N677, N672, N103, N258);
buf BUF1 (N678, N677);
nor NOR3 (N679, N675, N76, N268);
nor NOR4 (N680, N673, N357, N269, N43);
xor XOR2 (N681, N670, N111);
and AND4 (N682, N680, N456, N50, N623);
xor XOR2 (N683, N682, N546);
xor XOR2 (N684, N683, N227);
not NOT1 (N685, N676);
not NOT1 (N686, N669);
and AND4 (N687, N684, N165, N343, N375);
nor NOR2 (N688, N652, N632);
nor NOR2 (N689, N688, N106);
and AND2 (N690, N689, N287);
nand NAND3 (N691, N671, N582, N20);
buf BUF1 (N692, N679);
or OR2 (N693, N674, N412);
buf BUF1 (N694, N686);
or OR3 (N695, N693, N617, N341);
nand NAND2 (N696, N692, N19);
buf BUF1 (N697, N685);
xor XOR2 (N698, N681, N695);
xor XOR2 (N699, N394, N661);
nand NAND3 (N700, N699, N194, N688);
xor XOR2 (N701, N698, N463);
buf BUF1 (N702, N696);
and AND3 (N703, N701, N202, N211);
nor NOR2 (N704, N694, N677);
or OR2 (N705, N678, N371);
xor XOR2 (N706, N687, N620);
not NOT1 (N707, N664);
buf BUF1 (N708, N707);
not NOT1 (N709, N700);
buf BUF1 (N710, N690);
xor XOR2 (N711, N705, N196);
not NOT1 (N712, N709);
nor NOR3 (N713, N691, N686, N658);
or OR2 (N714, N697, N441);
buf BUF1 (N715, N708);
xor XOR2 (N716, N710, N212);
xor XOR2 (N717, N702, N86);
nor NOR3 (N718, N715, N374, N361);
buf BUF1 (N719, N713);
nand NAND4 (N720, N711, N389, N280, N508);
xor XOR2 (N721, N703, N197);
nand NAND2 (N722, N720, N629);
xor XOR2 (N723, N721, N70);
or OR4 (N724, N716, N176, N362, N343);
xor XOR2 (N725, N719, N188);
and AND2 (N726, N722, N350);
xor XOR2 (N727, N725, N654);
nand NAND2 (N728, N718, N273);
buf BUF1 (N729, N727);
buf BUF1 (N730, N729);
and AND4 (N731, N726, N685, N554, N332);
not NOT1 (N732, N730);
and AND3 (N733, N732, N263, N575);
or OR3 (N734, N704, N541, N47);
buf BUF1 (N735, N712);
not NOT1 (N736, N731);
buf BUF1 (N737, N734);
and AND3 (N738, N728, N640, N51);
not NOT1 (N739, N706);
not NOT1 (N740, N724);
or OR3 (N741, N738, N459, N267);
not NOT1 (N742, N737);
nor NOR3 (N743, N714, N538, N169);
buf BUF1 (N744, N743);
or OR2 (N745, N735, N85);
and AND3 (N746, N740, N406, N438);
nor NOR2 (N747, N741, N242);
xor XOR2 (N748, N745, N128);
nand NAND4 (N749, N717, N620, N640, N717);
nand NAND3 (N750, N742, N706, N440);
and AND3 (N751, N748, N461, N99);
and AND3 (N752, N749, N281, N739);
and AND2 (N753, N331, N352);
not NOT1 (N754, N733);
nand NAND2 (N755, N744, N232);
nor NOR4 (N756, N751, N56, N745, N517);
not NOT1 (N757, N753);
nand NAND4 (N758, N723, N307, N711, N657);
buf BUF1 (N759, N757);
and AND3 (N760, N756, N474, N136);
and AND4 (N761, N736, N401, N755, N207);
and AND3 (N762, N605, N343, N74);
buf BUF1 (N763, N758);
nand NAND2 (N764, N750, N52);
nor NOR3 (N765, N759, N368, N678);
buf BUF1 (N766, N765);
xor XOR2 (N767, N752, N117);
nor NOR2 (N768, N767, N282);
nor NOR2 (N769, N768, N581);
xor XOR2 (N770, N760, N640);
nor NOR3 (N771, N766, N727, N565);
and AND2 (N772, N764, N584);
nand NAND2 (N773, N754, N367);
not NOT1 (N774, N762);
nand NAND2 (N775, N774, N602);
or OR4 (N776, N770, N234, N709, N555);
not NOT1 (N777, N773);
buf BUF1 (N778, N772);
nor NOR3 (N779, N746, N734, N381);
not NOT1 (N780, N777);
not NOT1 (N781, N761);
and AND4 (N782, N781, N339, N672, N708);
and AND4 (N783, N747, N200, N211, N689);
nor NOR2 (N784, N782, N543);
buf BUF1 (N785, N780);
or OR3 (N786, N779, N419, N662);
xor XOR2 (N787, N778, N111);
nand NAND2 (N788, N771, N561);
buf BUF1 (N789, N763);
nor NOR3 (N790, N783, N729, N17);
or OR2 (N791, N786, N250);
or OR4 (N792, N785, N562, N144, N233);
not NOT1 (N793, N784);
buf BUF1 (N794, N793);
nor NOR2 (N795, N790, N747);
and AND4 (N796, N776, N146, N545, N697);
xor XOR2 (N797, N795, N110);
or OR3 (N798, N791, N155, N279);
nor NOR4 (N799, N775, N34, N161, N463);
nor NOR2 (N800, N787, N797);
and AND3 (N801, N653, N578, N773);
nor NOR4 (N802, N792, N334, N372, N331);
nor NOR4 (N803, N802, N747, N506, N635);
or OR3 (N804, N801, N218, N119);
nand NAND3 (N805, N788, N656, N132);
nor NOR3 (N806, N796, N24, N259);
nand NAND2 (N807, N805, N806);
xor XOR2 (N808, N315, N266);
or OR2 (N809, N800, N480);
nand NAND2 (N810, N769, N48);
or OR3 (N811, N809, N332, N348);
xor XOR2 (N812, N794, N749);
xor XOR2 (N813, N803, N437);
or OR3 (N814, N798, N507, N19);
xor XOR2 (N815, N804, N635);
xor XOR2 (N816, N815, N476);
nor NOR3 (N817, N814, N301, N709);
buf BUF1 (N818, N807);
nor NOR3 (N819, N789, N639, N195);
and AND4 (N820, N817, N768, N359, N106);
nand NAND2 (N821, N810, N370);
buf BUF1 (N822, N813);
buf BUF1 (N823, N820);
xor XOR2 (N824, N812, N259);
nand NAND2 (N825, N818, N753);
buf BUF1 (N826, N816);
and AND2 (N827, N824, N138);
or OR3 (N828, N821, N730, N291);
xor XOR2 (N829, N823, N285);
nand NAND2 (N830, N828, N408);
buf BUF1 (N831, N827);
nor NOR2 (N832, N825, N253);
buf BUF1 (N833, N819);
nand NAND2 (N834, N829, N226);
or OR3 (N835, N811, N359, N780);
buf BUF1 (N836, N830);
and AND4 (N837, N808, N111, N350, N9);
nor NOR3 (N838, N833, N207, N308);
or OR2 (N839, N831, N620);
buf BUF1 (N840, N832);
buf BUF1 (N841, N835);
not NOT1 (N842, N822);
not NOT1 (N843, N799);
xor XOR2 (N844, N843, N41);
xor XOR2 (N845, N844, N700);
nor NOR3 (N846, N838, N51, N246);
buf BUF1 (N847, N826);
nor NOR3 (N848, N847, N581, N406);
or OR3 (N849, N845, N14, N562);
not NOT1 (N850, N837);
nand NAND2 (N851, N850, N628);
and AND2 (N852, N851, N150);
buf BUF1 (N853, N848);
buf BUF1 (N854, N836);
or OR4 (N855, N849, N440, N801, N734);
buf BUF1 (N856, N852);
and AND4 (N857, N855, N664, N846, N826);
nand NAND4 (N858, N634, N376, N491, N13);
nand NAND2 (N859, N853, N560);
nand NAND3 (N860, N834, N558, N256);
and AND2 (N861, N854, N455);
not NOT1 (N862, N840);
nor NOR4 (N863, N856, N512, N531, N54);
nand NAND3 (N864, N842, N860, N240);
nand NAND2 (N865, N700, N65);
and AND4 (N866, N839, N355, N134, N664);
nand NAND3 (N867, N866, N830, N44);
buf BUF1 (N868, N863);
not NOT1 (N869, N868);
buf BUF1 (N870, N862);
xor XOR2 (N871, N865, N38);
or OR2 (N872, N859, N314);
xor XOR2 (N873, N841, N22);
not NOT1 (N874, N864);
buf BUF1 (N875, N872);
nor NOR2 (N876, N858, N114);
or OR4 (N877, N870, N122, N546, N667);
nand NAND3 (N878, N877, N624, N685);
not NOT1 (N879, N857);
xor XOR2 (N880, N861, N146);
not NOT1 (N881, N875);
xor XOR2 (N882, N878, N861);
nand NAND2 (N883, N881, N736);
or OR2 (N884, N867, N851);
and AND4 (N885, N871, N853, N496, N481);
not NOT1 (N886, N883);
and AND2 (N887, N873, N473);
xor XOR2 (N888, N879, N81);
nand NAND2 (N889, N876, N547);
nand NAND3 (N890, N882, N490, N502);
buf BUF1 (N891, N874);
and AND3 (N892, N869, N563, N4);
nand NAND3 (N893, N884, N356, N138);
nor NOR3 (N894, N891, N123, N342);
buf BUF1 (N895, N889);
and AND2 (N896, N888, N457);
buf BUF1 (N897, N892);
and AND2 (N898, N897, N746);
nor NOR2 (N899, N880, N500);
and AND3 (N900, N893, N116, N533);
and AND4 (N901, N900, N4, N83, N533);
or OR2 (N902, N885, N612);
and AND4 (N903, N901, N499, N371, N429);
or OR4 (N904, N886, N284, N274, N726);
not NOT1 (N905, N887);
nand NAND3 (N906, N905, N205, N622);
buf BUF1 (N907, N898);
xor XOR2 (N908, N904, N686);
or OR3 (N909, N894, N356, N62);
nor NOR4 (N910, N890, N17, N355, N200);
buf BUF1 (N911, N903);
not NOT1 (N912, N895);
or OR2 (N913, N906, N205);
not NOT1 (N914, N912);
xor XOR2 (N915, N909, N107);
and AND2 (N916, N914, N632);
buf BUF1 (N917, N907);
nand NAND3 (N918, N916, N157, N823);
not NOT1 (N919, N911);
buf BUF1 (N920, N910);
buf BUF1 (N921, N896);
xor XOR2 (N922, N902, N852);
not NOT1 (N923, N908);
not NOT1 (N924, N922);
or OR3 (N925, N923, N79, N422);
buf BUF1 (N926, N919);
not NOT1 (N927, N917);
buf BUF1 (N928, N924);
and AND2 (N929, N918, N424);
or OR3 (N930, N913, N715, N774);
or OR3 (N931, N929, N713, N286);
buf BUF1 (N932, N899);
nor NOR2 (N933, N930, N640);
nand NAND3 (N934, N915, N738, N35);
nor NOR4 (N935, N934, N707, N225, N831);
or OR3 (N936, N928, N45, N32);
nor NOR3 (N937, N936, N80, N482);
nor NOR2 (N938, N935, N874);
and AND3 (N939, N931, N352, N594);
nand NAND3 (N940, N921, N876, N471);
not NOT1 (N941, N932);
xor XOR2 (N942, N925, N741);
or OR2 (N943, N940, N382);
xor XOR2 (N944, N939, N704);
nor NOR4 (N945, N933, N670, N2, N724);
buf BUF1 (N946, N937);
nand NAND2 (N947, N938, N779);
nand NAND4 (N948, N942, N907, N437, N133);
nor NOR4 (N949, N941, N487, N71, N695);
nand NAND4 (N950, N927, N684, N842, N637);
not NOT1 (N951, N949);
nor NOR2 (N952, N948, N370);
nand NAND4 (N953, N947, N285, N768, N205);
buf BUF1 (N954, N926);
or OR4 (N955, N945, N263, N381, N150);
and AND3 (N956, N954, N281, N825);
nor NOR4 (N957, N950, N693, N951, N655);
and AND4 (N958, N388, N902, N660, N875);
or OR3 (N959, N957, N405, N879);
not NOT1 (N960, N920);
and AND3 (N961, N952, N816, N671);
buf BUF1 (N962, N944);
nor NOR3 (N963, N958, N69, N538);
or OR3 (N964, N946, N949, N551);
nor NOR3 (N965, N959, N473, N80);
nor NOR2 (N966, N953, N35);
or OR2 (N967, N955, N742);
xor XOR2 (N968, N962, N9);
nand NAND2 (N969, N964, N123);
or OR4 (N970, N943, N509, N486, N652);
buf BUF1 (N971, N970);
or OR2 (N972, N967, N175);
buf BUF1 (N973, N961);
or OR4 (N974, N972, N735, N957, N322);
or OR2 (N975, N973, N84);
not NOT1 (N976, N960);
and AND3 (N977, N975, N820, N647);
buf BUF1 (N978, N969);
and AND2 (N979, N965, N629);
nor NOR2 (N980, N977, N585);
or OR4 (N981, N974, N541, N738, N770);
and AND3 (N982, N978, N111, N373);
not NOT1 (N983, N963);
nand NAND2 (N984, N982, N305);
or OR2 (N985, N979, N893);
not NOT1 (N986, N981);
nand NAND2 (N987, N966, N707);
or OR4 (N988, N956, N877, N629, N6);
or OR2 (N989, N971, N659);
or OR3 (N990, N989, N940, N125);
nand NAND4 (N991, N980, N361, N836, N834);
or OR3 (N992, N990, N714, N506);
xor XOR2 (N993, N968, N961);
xor XOR2 (N994, N993, N122);
nand NAND3 (N995, N986, N514, N534);
nand NAND2 (N996, N994, N619);
xor XOR2 (N997, N988, N36);
xor XOR2 (N998, N997, N703);
buf BUF1 (N999, N998);
buf BUF1 (N1000, N992);
and AND4 (N1001, N987, N411, N424, N540);
nand NAND2 (N1002, N991, N922);
or OR4 (N1003, N1001, N383, N804, N229);
not NOT1 (N1004, N996);
nor NOR2 (N1005, N1003, N573);
and AND4 (N1006, N1002, N819, N93, N649);
nand NAND3 (N1007, N1000, N587, N505);
xor XOR2 (N1008, N985, N840);
buf BUF1 (N1009, N1005);
or OR3 (N1010, N976, N263, N309);
buf BUF1 (N1011, N1007);
not NOT1 (N1012, N1011);
buf BUF1 (N1013, N1008);
or OR2 (N1014, N983, N314);
not NOT1 (N1015, N999);
nor NOR2 (N1016, N1004, N854);
not NOT1 (N1017, N1009);
and AND2 (N1018, N1015, N113);
buf BUF1 (N1019, N1018);
and AND4 (N1020, N1010, N677, N254, N192);
not NOT1 (N1021, N1017);
or OR3 (N1022, N1016, N204, N478);
buf BUF1 (N1023, N1022);
nand NAND4 (N1024, N1013, N109, N359, N432);
nor NOR4 (N1025, N1020, N216, N1014, N38);
or OR3 (N1026, N238, N352, N694);
and AND3 (N1027, N1026, N204, N364);
nor NOR2 (N1028, N1025, N890);
xor XOR2 (N1029, N1012, N106);
not NOT1 (N1030, N1006);
nor NOR4 (N1031, N1023, N245, N674, N582);
buf BUF1 (N1032, N1024);
or OR4 (N1033, N1030, N382, N334, N435);
nand NAND2 (N1034, N1029, N348);
or OR2 (N1035, N1021, N942);
or OR3 (N1036, N1027, N299, N477);
xor XOR2 (N1037, N1028, N608);
nand NAND4 (N1038, N1034, N374, N995, N189);
xor XOR2 (N1039, N850, N69);
nand NAND4 (N1040, N1031, N844, N266, N439);
not NOT1 (N1041, N1035);
or OR2 (N1042, N1019, N768);
nand NAND4 (N1043, N1039, N221, N1009, N376);
not NOT1 (N1044, N1036);
or OR4 (N1045, N1038, N22, N354, N902);
xor XOR2 (N1046, N1042, N661);
buf BUF1 (N1047, N1033);
buf BUF1 (N1048, N1045);
nor NOR3 (N1049, N1044, N522, N1007);
nor NOR4 (N1050, N984, N315, N994, N375);
nand NAND4 (N1051, N1050, N714, N414, N958);
and AND3 (N1052, N1048, N217, N673);
xor XOR2 (N1053, N1049, N192);
and AND4 (N1054, N1052, N607, N389, N180);
xor XOR2 (N1055, N1047, N744);
nand NAND2 (N1056, N1043, N941);
and AND2 (N1057, N1037, N967);
not NOT1 (N1058, N1053);
not NOT1 (N1059, N1058);
or OR3 (N1060, N1051, N821, N403);
and AND4 (N1061, N1046, N503, N798, N422);
nor NOR2 (N1062, N1061, N406);
xor XOR2 (N1063, N1056, N397);
not NOT1 (N1064, N1041);
xor XOR2 (N1065, N1060, N508);
or OR3 (N1066, N1065, N115, N226);
or OR4 (N1067, N1066, N840, N76, N765);
or OR3 (N1068, N1032, N106, N931);
xor XOR2 (N1069, N1068, N1002);
nand NAND4 (N1070, N1064, N232, N276, N326);
or OR3 (N1071, N1067, N627, N172);
nand NAND3 (N1072, N1062, N373, N29);
not NOT1 (N1073, N1055);
xor XOR2 (N1074, N1070, N838);
or OR2 (N1075, N1059, N814);
nand NAND2 (N1076, N1057, N820);
nand NAND4 (N1077, N1074, N1037, N459, N327);
and AND3 (N1078, N1075, N968, N251);
or OR3 (N1079, N1063, N228, N107);
nand NAND3 (N1080, N1077, N139, N413);
xor XOR2 (N1081, N1072, N119);
nand NAND4 (N1082, N1040, N775, N852, N904);
buf BUF1 (N1083, N1073);
nand NAND4 (N1084, N1071, N637, N646, N550);
buf BUF1 (N1085, N1080);
and AND3 (N1086, N1069, N994, N131);
not NOT1 (N1087, N1076);
nor NOR2 (N1088, N1084, N325);
not NOT1 (N1089, N1088);
and AND3 (N1090, N1079, N794, N484);
or OR4 (N1091, N1085, N695, N674, N1026);
nor NOR4 (N1092, N1091, N778, N983, N622);
nand NAND2 (N1093, N1081, N900);
xor XOR2 (N1094, N1092, N1085);
nand NAND2 (N1095, N1093, N852);
not NOT1 (N1096, N1054);
and AND3 (N1097, N1087, N905, N1025);
xor XOR2 (N1098, N1095, N416);
not NOT1 (N1099, N1078);
nor NOR4 (N1100, N1089, N732, N1087, N729);
nor NOR3 (N1101, N1100, N89, N926);
buf BUF1 (N1102, N1097);
and AND2 (N1103, N1099, N149);
nand NAND3 (N1104, N1101, N1027, N687);
nor NOR2 (N1105, N1102, N508);
xor XOR2 (N1106, N1096, N780);
xor XOR2 (N1107, N1094, N900);
not NOT1 (N1108, N1083);
and AND2 (N1109, N1103, N140);
not NOT1 (N1110, N1104);
or OR3 (N1111, N1110, N245, N49);
or OR3 (N1112, N1090, N541, N988);
nand NAND3 (N1113, N1111, N473, N1111);
nand NAND4 (N1114, N1112, N37, N954, N459);
xor XOR2 (N1115, N1114, N928);
nand NAND4 (N1116, N1106, N805, N255, N300);
buf BUF1 (N1117, N1108);
buf BUF1 (N1118, N1109);
xor XOR2 (N1119, N1118, N1018);
not NOT1 (N1120, N1105);
xor XOR2 (N1121, N1107, N990);
not NOT1 (N1122, N1098);
or OR4 (N1123, N1119, N851, N135, N997);
not NOT1 (N1124, N1082);
buf BUF1 (N1125, N1121);
not NOT1 (N1126, N1113);
nor NOR4 (N1127, N1123, N823, N447, N804);
not NOT1 (N1128, N1127);
not NOT1 (N1129, N1125);
xor XOR2 (N1130, N1128, N581);
or OR4 (N1131, N1129, N450, N972, N594);
xor XOR2 (N1132, N1120, N369);
xor XOR2 (N1133, N1126, N940);
xor XOR2 (N1134, N1116, N1006);
and AND2 (N1135, N1086, N805);
xor XOR2 (N1136, N1133, N473);
nor NOR4 (N1137, N1134, N895, N986, N928);
or OR3 (N1138, N1115, N602, N148);
or OR2 (N1139, N1136, N318);
xor XOR2 (N1140, N1117, N311);
xor XOR2 (N1141, N1139, N263);
not NOT1 (N1142, N1137);
nor NOR4 (N1143, N1142, N495, N1032, N258);
or OR2 (N1144, N1140, N39);
nor NOR3 (N1145, N1122, N84, N1129);
and AND2 (N1146, N1130, N907);
buf BUF1 (N1147, N1138);
and AND4 (N1148, N1146, N1080, N911, N1056);
and AND3 (N1149, N1144, N1037, N383);
not NOT1 (N1150, N1147);
xor XOR2 (N1151, N1124, N249);
xor XOR2 (N1152, N1150, N972);
and AND3 (N1153, N1145, N866, N1070);
not NOT1 (N1154, N1151);
nand NAND4 (N1155, N1148, N376, N347, N739);
buf BUF1 (N1156, N1135);
nand NAND2 (N1157, N1152, N382);
or OR2 (N1158, N1155, N642);
xor XOR2 (N1159, N1141, N468);
xor XOR2 (N1160, N1131, N990);
nand NAND4 (N1161, N1153, N390, N731, N38);
and AND4 (N1162, N1159, N502, N627, N637);
and AND4 (N1163, N1157, N990, N557, N371);
buf BUF1 (N1164, N1162);
xor XOR2 (N1165, N1156, N57);
and AND2 (N1166, N1149, N494);
and AND3 (N1167, N1163, N835, N921);
and AND2 (N1168, N1154, N18);
and AND4 (N1169, N1160, N474, N491, N735);
and AND4 (N1170, N1168, N1015, N559, N96);
and AND3 (N1171, N1132, N71, N951);
not NOT1 (N1172, N1166);
and AND3 (N1173, N1169, N100, N907);
nand NAND3 (N1174, N1171, N169, N1103);
not NOT1 (N1175, N1174);
xor XOR2 (N1176, N1164, N954);
not NOT1 (N1177, N1175);
and AND4 (N1178, N1172, N871, N337, N101);
nor NOR3 (N1179, N1161, N1061, N354);
nand NAND4 (N1180, N1176, N663, N747, N345);
buf BUF1 (N1181, N1173);
nand NAND2 (N1182, N1178, N130);
nand NAND2 (N1183, N1165, N420);
nor NOR3 (N1184, N1158, N779, N939);
and AND4 (N1185, N1181, N864, N786, N917);
and AND4 (N1186, N1184, N1101, N1025, N295);
xor XOR2 (N1187, N1167, N839);
not NOT1 (N1188, N1177);
and AND4 (N1189, N1188, N758, N546, N910);
and AND3 (N1190, N1170, N804, N971);
nand NAND2 (N1191, N1180, N570);
or OR4 (N1192, N1179, N948, N1161, N1155);
xor XOR2 (N1193, N1191, N569);
nor NOR4 (N1194, N1185, N497, N969, N977);
nand NAND4 (N1195, N1186, N300, N964, N872);
and AND3 (N1196, N1189, N275, N623);
or OR2 (N1197, N1192, N570);
and AND3 (N1198, N1182, N137, N906);
buf BUF1 (N1199, N1194);
buf BUF1 (N1200, N1197);
nand NAND4 (N1201, N1199, N497, N305, N168);
or OR3 (N1202, N1190, N986, N103);
xor XOR2 (N1203, N1143, N939);
not NOT1 (N1204, N1193);
nor NOR3 (N1205, N1201, N101, N249);
nor NOR4 (N1206, N1198, N269, N913, N438);
and AND4 (N1207, N1205, N518, N1000, N144);
xor XOR2 (N1208, N1203, N921);
and AND3 (N1209, N1208, N743, N1193);
nor NOR3 (N1210, N1209, N345, N790);
and AND4 (N1211, N1206, N1130, N918, N728);
not NOT1 (N1212, N1200);
nand NAND2 (N1213, N1212, N456);
nand NAND2 (N1214, N1187, N965);
xor XOR2 (N1215, N1207, N195);
nand NAND4 (N1216, N1215, N574, N824, N150);
nor NOR2 (N1217, N1216, N539);
buf BUF1 (N1218, N1202);
nand NAND3 (N1219, N1213, N115, N844);
and AND3 (N1220, N1219, N77, N638);
nor NOR4 (N1221, N1204, N519, N560, N1112);
not NOT1 (N1222, N1195);
and AND4 (N1223, N1221, N553, N670, N968);
nor NOR4 (N1224, N1222, N443, N1176, N294);
or OR4 (N1225, N1196, N66, N407, N506);
nor NOR2 (N1226, N1218, N661);
nor NOR2 (N1227, N1217, N351);
and AND4 (N1228, N1226, N637, N184, N83);
and AND4 (N1229, N1223, N1118, N979, N726);
or OR3 (N1230, N1210, N496, N1126);
or OR2 (N1231, N1227, N564);
nor NOR3 (N1232, N1228, N75, N1015);
nand NAND3 (N1233, N1232, N649, N90);
or OR4 (N1234, N1233, N1178, N853, N536);
not NOT1 (N1235, N1231);
xor XOR2 (N1236, N1183, N742);
buf BUF1 (N1237, N1220);
not NOT1 (N1238, N1214);
and AND3 (N1239, N1211, N457, N612);
nand NAND4 (N1240, N1236, N465, N27, N818);
nand NAND4 (N1241, N1234, N1212, N540, N507);
not NOT1 (N1242, N1224);
nor NOR3 (N1243, N1237, N888, N282);
not NOT1 (N1244, N1239);
nand NAND3 (N1245, N1240, N975, N1201);
or OR3 (N1246, N1229, N1028, N1053);
not NOT1 (N1247, N1230);
nor NOR3 (N1248, N1244, N216, N1172);
buf BUF1 (N1249, N1238);
nor NOR3 (N1250, N1243, N1087, N639);
nand NAND3 (N1251, N1245, N805, N371);
not NOT1 (N1252, N1235);
and AND2 (N1253, N1250, N242);
or OR4 (N1254, N1249, N403, N25, N817);
not NOT1 (N1255, N1253);
and AND3 (N1256, N1247, N856, N1135);
xor XOR2 (N1257, N1252, N181);
and AND4 (N1258, N1251, N572, N1090, N79);
or OR3 (N1259, N1258, N1155, N1153);
and AND4 (N1260, N1257, N221, N709, N841);
xor XOR2 (N1261, N1246, N107);
buf BUF1 (N1262, N1248);
and AND2 (N1263, N1241, N953);
buf BUF1 (N1264, N1255);
nor NOR3 (N1265, N1263, N1220, N47);
buf BUF1 (N1266, N1265);
nor NOR2 (N1267, N1266, N1203);
and AND4 (N1268, N1262, N891, N757, N550);
buf BUF1 (N1269, N1225);
and AND4 (N1270, N1268, N747, N1176, N802);
or OR3 (N1271, N1254, N329, N71);
xor XOR2 (N1272, N1267, N888);
and AND4 (N1273, N1260, N590, N508, N1172);
not NOT1 (N1274, N1270);
xor XOR2 (N1275, N1256, N896);
buf BUF1 (N1276, N1271);
nand NAND3 (N1277, N1242, N644, N771);
or OR3 (N1278, N1274, N179, N141);
and AND2 (N1279, N1261, N401);
or OR3 (N1280, N1264, N796, N373);
xor XOR2 (N1281, N1269, N1159);
not NOT1 (N1282, N1259);
nor NOR2 (N1283, N1278, N428);
nand NAND4 (N1284, N1283, N1209, N602, N463);
nor NOR4 (N1285, N1280, N852, N631, N961);
not NOT1 (N1286, N1272);
not NOT1 (N1287, N1282);
buf BUF1 (N1288, N1285);
and AND2 (N1289, N1281, N168);
and AND2 (N1290, N1289, N1168);
or OR3 (N1291, N1279, N750, N30);
or OR3 (N1292, N1291, N1164, N166);
or OR3 (N1293, N1275, N693, N1289);
nor NOR4 (N1294, N1284, N1115, N3, N214);
and AND4 (N1295, N1286, N995, N1260, N1216);
buf BUF1 (N1296, N1287);
nand NAND3 (N1297, N1288, N211, N506);
xor XOR2 (N1298, N1277, N1098);
not NOT1 (N1299, N1295);
and AND4 (N1300, N1273, N688, N177, N601);
buf BUF1 (N1301, N1290);
nor NOR2 (N1302, N1297, N225);
nor NOR4 (N1303, N1296, N609, N1219, N126);
buf BUF1 (N1304, N1298);
and AND2 (N1305, N1294, N55);
not NOT1 (N1306, N1304);
not NOT1 (N1307, N1293);
nand NAND4 (N1308, N1292, N1223, N1295, N1229);
xor XOR2 (N1309, N1301, N1251);
nor NOR2 (N1310, N1300, N1153);
or OR3 (N1311, N1299, N1011, N904);
and AND4 (N1312, N1306, N717, N473, N1306);
not NOT1 (N1313, N1312);
nor NOR3 (N1314, N1313, N831, N268);
buf BUF1 (N1315, N1302);
nand NAND2 (N1316, N1307, N148);
nand NAND4 (N1317, N1315, N947, N988, N1248);
buf BUF1 (N1318, N1308);
xor XOR2 (N1319, N1276, N266);
xor XOR2 (N1320, N1311, N506);
nor NOR4 (N1321, N1317, N770, N893, N681);
xor XOR2 (N1322, N1314, N1209);
not NOT1 (N1323, N1310);
xor XOR2 (N1324, N1321, N1212);
not NOT1 (N1325, N1316);
nor NOR3 (N1326, N1309, N433, N406);
nand NAND2 (N1327, N1318, N210);
xor XOR2 (N1328, N1303, N628);
buf BUF1 (N1329, N1327);
not NOT1 (N1330, N1320);
xor XOR2 (N1331, N1322, N551);
nand NAND3 (N1332, N1323, N24, N701);
buf BUF1 (N1333, N1324);
not NOT1 (N1334, N1329);
xor XOR2 (N1335, N1330, N442);
buf BUF1 (N1336, N1334);
nand NAND2 (N1337, N1305, N1335);
or OR3 (N1338, N1015, N488, N383);
nor NOR2 (N1339, N1319, N766);
buf BUF1 (N1340, N1331);
nand NAND2 (N1341, N1337, N410);
xor XOR2 (N1342, N1325, N439);
xor XOR2 (N1343, N1338, N796);
or OR3 (N1344, N1339, N806, N514);
and AND4 (N1345, N1336, N288, N597, N824);
or OR2 (N1346, N1332, N1193);
not NOT1 (N1347, N1343);
or OR2 (N1348, N1326, N639);
xor XOR2 (N1349, N1333, N197);
xor XOR2 (N1350, N1342, N1082);
or OR4 (N1351, N1347, N300, N900, N1147);
xor XOR2 (N1352, N1344, N361);
not NOT1 (N1353, N1350);
and AND3 (N1354, N1353, N1276, N1221);
and AND3 (N1355, N1354, N1292, N1255);
nor NOR3 (N1356, N1340, N899, N1223);
or OR4 (N1357, N1351, N623, N475, N179);
nor NOR2 (N1358, N1357, N1309);
and AND4 (N1359, N1349, N73, N1337, N672);
nand NAND4 (N1360, N1359, N914, N802, N215);
and AND4 (N1361, N1346, N317, N651, N375);
buf BUF1 (N1362, N1355);
and AND2 (N1363, N1356, N1053);
or OR2 (N1364, N1361, N1344);
or OR3 (N1365, N1341, N168, N71);
or OR3 (N1366, N1352, N646, N269);
buf BUF1 (N1367, N1358);
buf BUF1 (N1368, N1366);
nor NOR3 (N1369, N1363, N627, N347);
nand NAND4 (N1370, N1367, N51, N965, N132);
xor XOR2 (N1371, N1365, N443);
nor NOR4 (N1372, N1370, N880, N597, N505);
not NOT1 (N1373, N1369);
or OR3 (N1374, N1364, N1017, N974);
buf BUF1 (N1375, N1371);
not NOT1 (N1376, N1372);
and AND2 (N1377, N1368, N772);
nor NOR2 (N1378, N1362, N514);
nor NOR2 (N1379, N1375, N476);
nor NOR2 (N1380, N1378, N690);
or OR4 (N1381, N1348, N431, N499, N629);
not NOT1 (N1382, N1380);
or OR3 (N1383, N1376, N669, N650);
and AND3 (N1384, N1360, N136, N769);
or OR4 (N1385, N1374, N551, N97, N826);
buf BUF1 (N1386, N1381);
nand NAND2 (N1387, N1345, N1376);
and AND2 (N1388, N1377, N676);
not NOT1 (N1389, N1328);
not NOT1 (N1390, N1387);
nor NOR2 (N1391, N1386, N1129);
or OR4 (N1392, N1382, N23, N609, N413);
nor NOR2 (N1393, N1379, N807);
or OR2 (N1394, N1384, N599);
nor NOR2 (N1395, N1383, N1027);
not NOT1 (N1396, N1385);
and AND2 (N1397, N1388, N1245);
nor NOR3 (N1398, N1394, N871, N8);
or OR3 (N1399, N1392, N578, N1119);
and AND2 (N1400, N1395, N876);
nor NOR3 (N1401, N1393, N528, N1095);
nor NOR2 (N1402, N1373, N913);
and AND4 (N1403, N1397, N684, N16, N135);
nand NAND4 (N1404, N1389, N1050, N30, N1177);
nor NOR3 (N1405, N1404, N608, N621);
nor NOR2 (N1406, N1401, N828);
nor NOR4 (N1407, N1391, N153, N1284, N1351);
nand NAND2 (N1408, N1402, N1329);
or OR4 (N1409, N1396, N50, N1376, N1296);
nor NOR3 (N1410, N1399, N233, N38);
or OR2 (N1411, N1390, N1141);
nand NAND2 (N1412, N1410, N247);
and AND3 (N1413, N1407, N1347, N1137);
xor XOR2 (N1414, N1406, N747);
not NOT1 (N1415, N1405);
xor XOR2 (N1416, N1398, N1333);
buf BUF1 (N1417, N1409);
xor XOR2 (N1418, N1403, N10);
buf BUF1 (N1419, N1413);
xor XOR2 (N1420, N1416, N412);
nand NAND3 (N1421, N1414, N1398, N792);
nand NAND4 (N1422, N1421, N1140, N254, N1201);
buf BUF1 (N1423, N1422);
nor NOR4 (N1424, N1423, N1337, N23, N717);
not NOT1 (N1425, N1419);
or OR4 (N1426, N1420, N114, N1423, N486);
and AND2 (N1427, N1408, N1258);
and AND4 (N1428, N1415, N1424, N41, N1188);
buf BUF1 (N1429, N12);
or OR3 (N1430, N1429, N636, N249);
nor NOR3 (N1431, N1411, N401, N963);
and AND2 (N1432, N1425, N507);
xor XOR2 (N1433, N1417, N690);
or OR2 (N1434, N1418, N202);
nor NOR2 (N1435, N1433, N929);
nor NOR4 (N1436, N1430, N668, N1006, N482);
or OR2 (N1437, N1412, N1315);
nand NAND2 (N1438, N1435, N6);
nor NOR3 (N1439, N1428, N153, N737);
nor NOR2 (N1440, N1400, N1242);
not NOT1 (N1441, N1439);
and AND2 (N1442, N1440, N802);
buf BUF1 (N1443, N1431);
nand NAND3 (N1444, N1427, N1077, N897);
or OR3 (N1445, N1437, N1086, N231);
xor XOR2 (N1446, N1445, N762);
not NOT1 (N1447, N1438);
not NOT1 (N1448, N1443);
not NOT1 (N1449, N1447);
or OR3 (N1450, N1432, N303, N1360);
xor XOR2 (N1451, N1426, N889);
nand NAND4 (N1452, N1444, N724, N234, N1105);
xor XOR2 (N1453, N1442, N87);
not NOT1 (N1454, N1446);
buf BUF1 (N1455, N1451);
nor NOR4 (N1456, N1453, N1445, N614, N978);
not NOT1 (N1457, N1436);
not NOT1 (N1458, N1455);
and AND2 (N1459, N1450, N1086);
and AND2 (N1460, N1434, N1334);
nand NAND4 (N1461, N1454, N1035, N1261, N296);
xor XOR2 (N1462, N1448, N146);
or OR2 (N1463, N1458, N207);
buf BUF1 (N1464, N1449);
buf BUF1 (N1465, N1441);
nor NOR4 (N1466, N1461, N966, N379, N876);
buf BUF1 (N1467, N1462);
nor NOR4 (N1468, N1457, N611, N770, N1014);
nor NOR2 (N1469, N1466, N136);
buf BUF1 (N1470, N1465);
nor NOR3 (N1471, N1464, N529, N958);
xor XOR2 (N1472, N1469, N795);
nand NAND2 (N1473, N1452, N967);
nand NAND3 (N1474, N1472, N877, N547);
and AND3 (N1475, N1460, N1004, N485);
buf BUF1 (N1476, N1459);
not NOT1 (N1477, N1475);
or OR2 (N1478, N1473, N380);
and AND4 (N1479, N1476, N1241, N939, N307);
xor XOR2 (N1480, N1477, N1311);
and AND3 (N1481, N1456, N1304, N706);
nand NAND3 (N1482, N1463, N21, N606);
nand NAND4 (N1483, N1474, N776, N1350, N1466);
or OR4 (N1484, N1471, N894, N518, N1232);
nor NOR4 (N1485, N1467, N554, N198, N570);
not NOT1 (N1486, N1484);
not NOT1 (N1487, N1486);
or OR2 (N1488, N1483, N105);
or OR2 (N1489, N1480, N403);
not NOT1 (N1490, N1489);
nor NOR2 (N1491, N1482, N825);
not NOT1 (N1492, N1490);
not NOT1 (N1493, N1488);
buf BUF1 (N1494, N1487);
nand NAND2 (N1495, N1492, N449);
or OR4 (N1496, N1468, N1028, N860, N637);
and AND3 (N1497, N1485, N163, N515);
xor XOR2 (N1498, N1495, N456);
xor XOR2 (N1499, N1498, N244);
xor XOR2 (N1500, N1499, N826);
and AND2 (N1501, N1479, N635);
not NOT1 (N1502, N1496);
xor XOR2 (N1503, N1478, N1334);
xor XOR2 (N1504, N1493, N1255);
and AND2 (N1505, N1481, N1028);
xor XOR2 (N1506, N1500, N1273);
not NOT1 (N1507, N1494);
and AND4 (N1508, N1491, N373, N938, N793);
buf BUF1 (N1509, N1507);
and AND2 (N1510, N1505, N104);
buf BUF1 (N1511, N1501);
endmodule