// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20;

output N1515,N1509,N1500,N1517,N1516,N1519,N1510,N1508,N1490,N1520;

not NOT1 (N21, N3);
not NOT1 (N22, N13);
or OR3 (N23, N22, N6, N8);
buf BUF1 (N24, N11);
nor NOR2 (N25, N10, N5);
and AND2 (N26, N23, N25);
nand NAND2 (N27, N26, N20);
nor NOR2 (N28, N21, N11);
or OR3 (N29, N19, N13, N2);
not NOT1 (N30, N20);
nor NOR4 (N31, N30, N11, N4, N7);
xor XOR2 (N32, N19, N23);
xor XOR2 (N33, N1, N7);
xor XOR2 (N34, N15, N31);
nor NOR4 (N35, N27, N4, N6, N2);
not NOT1 (N36, N29);
and AND4 (N37, N24, N15, N25, N7);
and AND2 (N38, N11, N26);
not NOT1 (N39, N35);
nand NAND4 (N40, N38, N1, N8, N12);
or OR2 (N41, N8, N14);
nor NOR3 (N42, N30, N14, N4);
nor NOR3 (N43, N34, N20, N29);
or OR4 (N44, N43, N23, N28, N26);
buf BUF1 (N45, N40);
or OR3 (N46, N42, N39, N1);
and AND2 (N47, N26, N23);
xor XOR2 (N48, N39, N46);
and AND2 (N49, N18, N22);
nand NAND3 (N50, N32, N46, N48);
or OR4 (N51, N7, N36, N14, N29);
buf BUF1 (N52, N15);
nor NOR2 (N53, N33, N44);
buf BUF1 (N54, N36);
xor XOR2 (N55, N53, N33);
xor XOR2 (N56, N50, N14);
xor XOR2 (N57, N47, N32);
nor NOR3 (N58, N54, N51, N15);
or OR4 (N59, N47, N22, N29, N7);
nand NAND4 (N60, N52, N5, N55, N48);
not NOT1 (N61, N56);
nand NAND3 (N62, N30, N27, N50);
buf BUF1 (N63, N45);
nand NAND4 (N64, N59, N22, N27, N51);
xor XOR2 (N65, N41, N33);
or OR2 (N66, N63, N2);
xor XOR2 (N67, N60, N9);
nor NOR2 (N68, N67, N29);
not NOT1 (N69, N64);
buf BUF1 (N70, N58);
nor NOR4 (N71, N70, N10, N14, N12);
buf BUF1 (N72, N71);
and AND4 (N73, N37, N5, N67, N46);
or OR2 (N74, N66, N20);
not NOT1 (N75, N73);
buf BUF1 (N76, N49);
or OR4 (N77, N74, N62, N71, N68);
nand NAND3 (N78, N50, N21, N42);
or OR3 (N79, N28, N22, N11);
nand NAND2 (N80, N65, N47);
xor XOR2 (N81, N78, N66);
buf BUF1 (N82, N57);
xor XOR2 (N83, N72, N31);
nand NAND3 (N84, N82, N2, N75);
xor XOR2 (N85, N33, N15);
nand NAND4 (N86, N85, N74, N71, N43);
xor XOR2 (N87, N69, N20);
not NOT1 (N88, N61);
nor NOR3 (N89, N83, N56, N80);
nor NOR4 (N90, N12, N27, N45, N37);
nor NOR3 (N91, N76, N55, N74);
nor NOR3 (N92, N91, N75, N28);
not NOT1 (N93, N79);
xor XOR2 (N94, N84, N57);
not NOT1 (N95, N87);
and AND2 (N96, N88, N3);
buf BUF1 (N97, N95);
nor NOR2 (N98, N90, N8);
not NOT1 (N99, N81);
buf BUF1 (N100, N98);
not NOT1 (N101, N89);
xor XOR2 (N102, N99, N13);
buf BUF1 (N103, N101);
xor XOR2 (N104, N86, N29);
nand NAND3 (N105, N97, N86, N55);
and AND2 (N106, N100, N26);
nor NOR4 (N107, N106, N15, N72, N50);
not NOT1 (N108, N96);
nor NOR4 (N109, N105, N73, N96, N31);
or OR3 (N110, N77, N57, N94);
or OR2 (N111, N52, N90);
nand NAND3 (N112, N111, N29, N70);
nand NAND3 (N113, N107, N30, N101);
or OR4 (N114, N108, N46, N66, N59);
and AND2 (N115, N112, N16);
xor XOR2 (N116, N92, N68);
not NOT1 (N117, N102);
nand NAND4 (N118, N115, N6, N105, N107);
nand NAND2 (N119, N109, N20);
nand NAND2 (N120, N113, N84);
nand NAND3 (N121, N119, N49, N58);
or OR2 (N122, N118, N77);
buf BUF1 (N123, N120);
or OR4 (N124, N110, N21, N16, N104);
buf BUF1 (N125, N12);
or OR3 (N126, N103, N29, N118);
or OR4 (N127, N125, N31, N29, N103);
and AND3 (N128, N116, N46, N20);
nand NAND2 (N129, N123, N32);
not NOT1 (N130, N129);
not NOT1 (N131, N128);
nand NAND3 (N132, N131, N11, N43);
and AND2 (N133, N124, N125);
xor XOR2 (N134, N122, N130);
not NOT1 (N135, N68);
not NOT1 (N136, N93);
and AND3 (N137, N126, N68, N50);
xor XOR2 (N138, N135, N128);
and AND3 (N139, N134, N56, N83);
nand NAND2 (N140, N114, N19);
or OR4 (N141, N140, N124, N52, N45);
not NOT1 (N142, N127);
or OR4 (N143, N121, N56, N45, N38);
not NOT1 (N144, N137);
and AND3 (N145, N139, N64, N5);
xor XOR2 (N146, N144, N23);
buf BUF1 (N147, N142);
xor XOR2 (N148, N136, N143);
nand NAND4 (N149, N60, N20, N122, N89);
or OR4 (N150, N147, N39, N74, N44);
and AND3 (N151, N138, N130, N135);
xor XOR2 (N152, N146, N111);
and AND2 (N153, N151, N108);
or OR4 (N154, N117, N102, N111, N106);
nand NAND3 (N155, N150, N149, N123);
or OR4 (N156, N16, N19, N10, N10);
buf BUF1 (N157, N155);
nor NOR4 (N158, N156, N141, N5, N148);
buf BUF1 (N159, N132);
buf BUF1 (N160, N58);
or OR3 (N161, N8, N76, N148);
and AND4 (N162, N145, N5, N45, N138);
not NOT1 (N163, N152);
not NOT1 (N164, N163);
xor XOR2 (N165, N161, N57);
nand NAND2 (N166, N157, N38);
nor NOR4 (N167, N162, N110, N164, N103);
or OR2 (N168, N97, N61);
or OR4 (N169, N167, N89, N67, N65);
or OR4 (N170, N168, N95, N71, N159);
and AND2 (N171, N50, N48);
nand NAND4 (N172, N158, N27, N98, N121);
not NOT1 (N173, N160);
nor NOR4 (N174, N154, N119, N9, N70);
xor XOR2 (N175, N153, N111);
not NOT1 (N176, N169);
not NOT1 (N177, N176);
not NOT1 (N178, N171);
or OR3 (N179, N165, N82, N16);
buf BUF1 (N180, N173);
xor XOR2 (N181, N180, N137);
buf BUF1 (N182, N177);
and AND3 (N183, N170, N13, N36);
and AND3 (N184, N172, N77, N74);
xor XOR2 (N185, N182, N55);
not NOT1 (N186, N178);
xor XOR2 (N187, N184, N7);
or OR2 (N188, N183, N63);
nand NAND3 (N189, N187, N176, N51);
buf BUF1 (N190, N133);
not NOT1 (N191, N190);
or OR4 (N192, N186, N95, N123, N184);
and AND2 (N193, N175, N10);
buf BUF1 (N194, N193);
xor XOR2 (N195, N174, N22);
nor NOR2 (N196, N189, N141);
xor XOR2 (N197, N179, N107);
xor XOR2 (N198, N185, N4);
nor NOR3 (N199, N195, N174, N186);
buf BUF1 (N200, N192);
not NOT1 (N201, N194);
nor NOR2 (N202, N188, N4);
or OR2 (N203, N199, N86);
nand NAND2 (N204, N166, N44);
not NOT1 (N205, N203);
or OR3 (N206, N191, N92, N97);
and AND2 (N207, N204, N23);
xor XOR2 (N208, N181, N169);
xor XOR2 (N209, N201, N195);
or OR4 (N210, N196, N73, N112, N130);
nand NAND2 (N211, N202, N100);
and AND3 (N212, N200, N43, N174);
and AND2 (N213, N212, N159);
not NOT1 (N214, N209);
xor XOR2 (N215, N211, N59);
xor XOR2 (N216, N206, N194);
xor XOR2 (N217, N214, N140);
or OR2 (N218, N207, N7);
buf BUF1 (N219, N210);
or OR2 (N220, N205, N94);
not NOT1 (N221, N197);
xor XOR2 (N222, N216, N70);
nand NAND4 (N223, N208, N35, N14, N162);
xor XOR2 (N224, N219, N7);
nand NAND3 (N225, N218, N186, N127);
nand NAND3 (N226, N224, N15, N57);
or OR2 (N227, N222, N17);
buf BUF1 (N228, N225);
nor NOR2 (N229, N226, N188);
not NOT1 (N230, N215);
or OR4 (N231, N213, N173, N101, N201);
buf BUF1 (N232, N223);
nor NOR3 (N233, N220, N33, N168);
nand NAND2 (N234, N227, N16);
nor NOR4 (N235, N234, N194, N31, N21);
or OR3 (N236, N230, N225, N213);
not NOT1 (N237, N229);
not NOT1 (N238, N233);
and AND4 (N239, N231, N46, N75, N188);
buf BUF1 (N240, N228);
nor NOR3 (N241, N217, N84, N68);
nor NOR3 (N242, N237, N165, N162);
or OR4 (N243, N238, N102, N185, N25);
nor NOR2 (N244, N243, N50);
and AND2 (N245, N239, N40);
nor NOR4 (N246, N236, N13, N187, N89);
buf BUF1 (N247, N241);
xor XOR2 (N248, N245, N84);
nor NOR2 (N249, N221, N171);
xor XOR2 (N250, N232, N33);
not NOT1 (N251, N250);
xor XOR2 (N252, N248, N204);
nor NOR4 (N253, N251, N252, N13, N176);
nor NOR2 (N254, N27, N78);
xor XOR2 (N255, N249, N44);
buf BUF1 (N256, N235);
nand NAND4 (N257, N240, N57, N43, N244);
nand NAND4 (N258, N93, N192, N99, N223);
buf BUF1 (N259, N257);
not NOT1 (N260, N256);
xor XOR2 (N261, N247, N87);
xor XOR2 (N262, N255, N165);
nand NAND4 (N263, N198, N92, N152, N17);
nor NOR4 (N264, N246, N91, N254, N29);
nor NOR4 (N265, N138, N191, N215, N125);
or OR2 (N266, N242, N74);
buf BUF1 (N267, N259);
xor XOR2 (N268, N258, N168);
or OR2 (N269, N253, N165);
and AND4 (N270, N261, N4, N13, N76);
xor XOR2 (N271, N263, N223);
buf BUF1 (N272, N265);
and AND4 (N273, N267, N65, N36, N70);
buf BUF1 (N274, N264);
xor XOR2 (N275, N266, N111);
nand NAND4 (N276, N271, N158, N49, N7);
or OR2 (N277, N273, N163);
xor XOR2 (N278, N274, N139);
nor NOR3 (N279, N268, N33, N85);
not NOT1 (N280, N260);
nor NOR3 (N281, N277, N239, N166);
xor XOR2 (N282, N272, N156);
not NOT1 (N283, N278);
nand NAND4 (N284, N269, N49, N123, N267);
and AND4 (N285, N281, N72, N80, N197);
nand NAND3 (N286, N283, N264, N36);
and AND4 (N287, N275, N63, N281, N157);
nor NOR4 (N288, N276, N90, N107, N214);
nor NOR4 (N289, N279, N220, N183, N275);
or OR3 (N290, N262, N286, N201);
not NOT1 (N291, N91);
nand NAND2 (N292, N288, N162);
buf BUF1 (N293, N292);
nand NAND2 (N294, N293, N48);
not NOT1 (N295, N282);
not NOT1 (N296, N287);
or OR2 (N297, N284, N255);
or OR4 (N298, N296, N85, N8, N80);
nand NAND4 (N299, N280, N267, N125, N123);
or OR4 (N300, N299, N42, N241, N166);
buf BUF1 (N301, N297);
xor XOR2 (N302, N295, N6);
or OR4 (N303, N301, N291, N178, N148);
xor XOR2 (N304, N151, N266);
or OR2 (N305, N298, N11);
nand NAND2 (N306, N294, N44);
nor NOR2 (N307, N306, N129);
nand NAND2 (N308, N304, N120);
buf BUF1 (N309, N285);
and AND4 (N310, N303, N147, N228, N154);
and AND4 (N311, N305, N167, N283, N184);
buf BUF1 (N312, N270);
nand NAND4 (N313, N307, N22, N245, N162);
buf BUF1 (N314, N311);
xor XOR2 (N315, N308, N122);
and AND2 (N316, N290, N221);
buf BUF1 (N317, N315);
not NOT1 (N318, N316);
xor XOR2 (N319, N302, N225);
nand NAND2 (N320, N319, N200);
not NOT1 (N321, N310);
or OR3 (N322, N312, N119, N46);
buf BUF1 (N323, N318);
not NOT1 (N324, N314);
buf BUF1 (N325, N320);
xor XOR2 (N326, N289, N55);
and AND4 (N327, N325, N28, N124, N308);
and AND3 (N328, N323, N85, N155);
nand NAND2 (N329, N326, N164);
nor NOR4 (N330, N313, N277, N37, N48);
nor NOR2 (N331, N309, N105);
or OR2 (N332, N330, N286);
nor NOR4 (N333, N327, N282, N194, N58);
or OR4 (N334, N324, N318, N45, N25);
nand NAND4 (N335, N329, N174, N165, N26);
and AND2 (N336, N335, N178);
nand NAND2 (N337, N336, N45);
nor NOR3 (N338, N321, N202, N172);
and AND3 (N339, N328, N316, N1);
buf BUF1 (N340, N317);
and AND3 (N341, N338, N223, N204);
and AND3 (N342, N334, N16, N42);
nand NAND4 (N343, N333, N341, N109, N100);
nor NOR3 (N344, N301, N6, N53);
or OR2 (N345, N300, N160);
nor NOR4 (N346, N331, N167, N179, N342);
xor XOR2 (N347, N82, N103);
nand NAND4 (N348, N346, N3, N207, N209);
buf BUF1 (N349, N332);
nand NAND4 (N350, N322, N244, N51, N117);
nor NOR4 (N351, N343, N72, N136, N306);
xor XOR2 (N352, N348, N326);
xor XOR2 (N353, N340, N113);
and AND3 (N354, N339, N285, N193);
not NOT1 (N355, N344);
buf BUF1 (N356, N350);
xor XOR2 (N357, N354, N95);
and AND3 (N358, N355, N324, N67);
not NOT1 (N359, N347);
xor XOR2 (N360, N352, N78);
nor NOR4 (N361, N357, N334, N161, N286);
nor NOR2 (N362, N353, N164);
nor NOR4 (N363, N356, N25, N15, N266);
and AND4 (N364, N349, N160, N242, N269);
or OR4 (N365, N345, N249, N163, N220);
not NOT1 (N366, N359);
not NOT1 (N367, N366);
xor XOR2 (N368, N364, N54);
buf BUF1 (N369, N358);
nand NAND4 (N370, N368, N95, N126, N295);
or OR4 (N371, N363, N185, N82, N60);
nor NOR2 (N372, N337, N122);
nand NAND4 (N373, N367, N354, N366, N308);
xor XOR2 (N374, N370, N185);
buf BUF1 (N375, N373);
nand NAND2 (N376, N365, N74);
nor NOR3 (N377, N351, N24, N272);
and AND2 (N378, N369, N127);
nand NAND2 (N379, N362, N207);
not NOT1 (N380, N378);
nand NAND4 (N381, N375, N98, N118, N72);
not NOT1 (N382, N380);
nor NOR3 (N383, N361, N168, N375);
not NOT1 (N384, N381);
nand NAND3 (N385, N383, N88, N43);
xor XOR2 (N386, N360, N203);
not NOT1 (N387, N371);
xor XOR2 (N388, N372, N352);
or OR3 (N389, N388, N104, N159);
nand NAND3 (N390, N379, N201, N172);
nand NAND2 (N391, N386, N245);
or OR4 (N392, N389, N180, N194, N113);
and AND3 (N393, N377, N352, N334);
nand NAND3 (N394, N384, N294, N198);
buf BUF1 (N395, N374);
buf BUF1 (N396, N392);
xor XOR2 (N397, N385, N344);
and AND4 (N398, N393, N317, N202, N209);
not NOT1 (N399, N397);
nor NOR2 (N400, N387, N131);
buf BUF1 (N401, N400);
or OR3 (N402, N398, N180, N8);
xor XOR2 (N403, N402, N308);
buf BUF1 (N404, N390);
or OR4 (N405, N404, N260, N60, N124);
or OR2 (N406, N394, N256);
nand NAND2 (N407, N395, N170);
nand NAND4 (N408, N396, N215, N312, N306);
and AND4 (N409, N391, N102, N95, N333);
buf BUF1 (N410, N407);
and AND4 (N411, N376, N296, N70, N118);
xor XOR2 (N412, N405, N259);
nor NOR2 (N413, N412, N241);
or OR2 (N414, N399, N122);
nand NAND4 (N415, N406, N14, N171, N271);
buf BUF1 (N416, N409);
not NOT1 (N417, N413);
nor NOR4 (N418, N401, N377, N411, N303);
and AND4 (N419, N146, N387, N328, N74);
and AND3 (N420, N419, N365, N109);
or OR4 (N421, N382, N19, N352, N270);
buf BUF1 (N422, N420);
xor XOR2 (N423, N414, N281);
and AND4 (N424, N415, N416, N392, N203);
not NOT1 (N425, N363);
nor NOR2 (N426, N425, N293);
and AND4 (N427, N426, N276, N48, N329);
and AND4 (N428, N403, N24, N171, N264);
or OR2 (N429, N422, N72);
buf BUF1 (N430, N423);
not NOT1 (N431, N430);
and AND4 (N432, N417, N350, N17, N396);
and AND2 (N433, N424, N143);
nand NAND3 (N434, N428, N122, N389);
nor NOR2 (N435, N427, N299);
not NOT1 (N436, N432);
nand NAND2 (N437, N434, N89);
buf BUF1 (N438, N429);
buf BUF1 (N439, N435);
or OR2 (N440, N421, N227);
buf BUF1 (N441, N439);
or OR4 (N442, N418, N156, N265, N356);
xor XOR2 (N443, N433, N190);
nand NAND4 (N444, N443, N402, N14, N295);
or OR2 (N445, N410, N292);
and AND2 (N446, N444, N426);
nor NOR3 (N447, N408, N375, N107);
xor XOR2 (N448, N437, N230);
and AND4 (N449, N441, N442, N16, N326);
or OR2 (N450, N419, N243);
or OR4 (N451, N446, N249, N387, N419);
and AND2 (N452, N449, N190);
or OR4 (N453, N436, N95, N108, N177);
xor XOR2 (N454, N431, N419);
and AND2 (N455, N450, N305);
nand NAND4 (N456, N455, N40, N37, N160);
and AND2 (N457, N440, N243);
xor XOR2 (N458, N452, N240);
nand NAND2 (N459, N453, N227);
buf BUF1 (N460, N459);
not NOT1 (N461, N451);
nand NAND3 (N462, N438, N185, N390);
or OR2 (N463, N448, N307);
buf BUF1 (N464, N456);
nor NOR2 (N465, N460, N14);
nor NOR2 (N466, N461, N435);
xor XOR2 (N467, N447, N216);
and AND2 (N468, N464, N360);
or OR4 (N469, N458, N438, N185, N33);
nor NOR2 (N470, N466, N9);
and AND2 (N471, N467, N283);
or OR4 (N472, N470, N435, N124, N82);
and AND4 (N473, N465, N36, N248, N232);
not NOT1 (N474, N445);
buf BUF1 (N475, N463);
xor XOR2 (N476, N468, N291);
nand NAND3 (N477, N469, N459, N360);
or OR4 (N478, N473, N384, N161, N208);
nand NAND4 (N479, N454, N446, N253, N125);
nor NOR3 (N480, N471, N447, N173);
and AND3 (N481, N477, N468, N248);
buf BUF1 (N482, N474);
nor NOR4 (N483, N481, N154, N424, N50);
nand NAND2 (N484, N457, N144);
or OR4 (N485, N484, N37, N468, N61);
xor XOR2 (N486, N478, N231);
and AND4 (N487, N479, N214, N348, N376);
xor XOR2 (N488, N480, N27);
nor NOR4 (N489, N462, N444, N185, N152);
and AND3 (N490, N486, N14, N196);
nand NAND2 (N491, N485, N465);
or OR4 (N492, N488, N308, N131, N89);
nor NOR2 (N493, N492, N351);
not NOT1 (N494, N489);
not NOT1 (N495, N483);
nor NOR3 (N496, N476, N76, N314);
or OR3 (N497, N493, N44, N138);
nand NAND4 (N498, N472, N145, N231, N211);
nand NAND2 (N499, N495, N204);
nand NAND4 (N500, N491, N100, N235, N406);
and AND4 (N501, N500, N248, N238, N66);
or OR2 (N502, N490, N38);
and AND3 (N503, N501, N393, N248);
nor NOR3 (N504, N482, N423, N478);
or OR4 (N505, N504, N483, N254, N156);
nor NOR2 (N506, N498, N161);
and AND2 (N507, N506, N270);
nand NAND4 (N508, N503, N188, N93, N103);
or OR3 (N509, N487, N347, N478);
or OR4 (N510, N505, N152, N277, N505);
or OR4 (N511, N508, N188, N385, N485);
and AND3 (N512, N507, N60, N460);
nand NAND4 (N513, N511, N427, N157, N356);
and AND2 (N514, N509, N61);
nor NOR3 (N515, N513, N41, N263);
xor XOR2 (N516, N496, N343);
buf BUF1 (N517, N514);
xor XOR2 (N518, N517, N486);
nor NOR4 (N519, N494, N258, N511, N175);
not NOT1 (N520, N512);
nor NOR4 (N521, N519, N132, N158, N347);
not NOT1 (N522, N515);
and AND3 (N523, N502, N402, N512);
or OR2 (N524, N499, N102);
buf BUF1 (N525, N520);
nor NOR4 (N526, N523, N2, N406, N521);
and AND2 (N527, N214, N414);
not NOT1 (N528, N516);
and AND3 (N529, N528, N268, N514);
or OR2 (N530, N526, N446);
xor XOR2 (N531, N530, N140);
buf BUF1 (N532, N522);
not NOT1 (N533, N510);
nor NOR4 (N534, N525, N63, N110, N299);
nor NOR2 (N535, N533, N34);
and AND3 (N536, N531, N82, N406);
buf BUF1 (N537, N518);
not NOT1 (N538, N536);
or OR3 (N539, N535, N449, N55);
buf BUF1 (N540, N524);
nor NOR2 (N541, N497, N40);
xor XOR2 (N542, N538, N86);
xor XOR2 (N543, N540, N270);
not NOT1 (N544, N527);
nor NOR4 (N545, N539, N116, N420, N183);
not NOT1 (N546, N541);
buf BUF1 (N547, N537);
nand NAND2 (N548, N542, N130);
buf BUF1 (N549, N534);
or OR3 (N550, N529, N50, N42);
nor NOR2 (N551, N548, N407);
nor NOR2 (N552, N544, N211);
nand NAND2 (N553, N543, N124);
nor NOR4 (N554, N532, N301, N93, N524);
not NOT1 (N555, N553);
and AND2 (N556, N545, N448);
xor XOR2 (N557, N475, N457);
nor NOR3 (N558, N552, N11, N423);
nand NAND4 (N559, N551, N215, N230, N305);
buf BUF1 (N560, N558);
or OR4 (N561, N555, N180, N182, N212);
not NOT1 (N562, N554);
xor XOR2 (N563, N561, N434);
nand NAND4 (N564, N559, N265, N124, N323);
or OR2 (N565, N547, N223);
nand NAND4 (N566, N563, N145, N521, N181);
or OR4 (N567, N564, N245, N100, N27);
nand NAND4 (N568, N546, N393, N476, N251);
nand NAND3 (N569, N567, N509, N272);
xor XOR2 (N570, N569, N398);
nand NAND2 (N571, N556, N263);
buf BUF1 (N572, N562);
not NOT1 (N573, N549);
buf BUF1 (N574, N568);
or OR2 (N575, N550, N6);
nor NOR2 (N576, N572, N42);
xor XOR2 (N577, N557, N287);
not NOT1 (N578, N574);
and AND2 (N579, N573, N517);
not NOT1 (N580, N579);
xor XOR2 (N581, N575, N334);
buf BUF1 (N582, N571);
not NOT1 (N583, N576);
and AND2 (N584, N566, N25);
or OR4 (N585, N577, N61, N401, N229);
buf BUF1 (N586, N570);
or OR3 (N587, N581, N412, N515);
or OR2 (N588, N586, N269);
not NOT1 (N589, N582);
nand NAND4 (N590, N560, N439, N179, N414);
not NOT1 (N591, N580);
xor XOR2 (N592, N584, N170);
nor NOR3 (N593, N588, N99, N258);
and AND3 (N594, N585, N298, N27);
nand NAND2 (N595, N589, N234);
xor XOR2 (N596, N590, N498);
nor NOR4 (N597, N587, N494, N422, N231);
buf BUF1 (N598, N594);
xor XOR2 (N599, N565, N187);
xor XOR2 (N600, N592, N303);
and AND2 (N601, N591, N520);
or OR3 (N602, N578, N465, N524);
nand NAND2 (N603, N593, N273);
xor XOR2 (N604, N601, N425);
not NOT1 (N605, N598);
or OR4 (N606, N600, N145, N182, N283);
nand NAND4 (N607, N595, N276, N198, N109);
not NOT1 (N608, N597);
xor XOR2 (N609, N583, N581);
nand NAND3 (N610, N606, N71, N596);
buf BUF1 (N611, N6);
xor XOR2 (N612, N607, N124);
nor NOR4 (N613, N612, N605, N51, N14);
or OR4 (N614, N53, N121, N537, N177);
nand NAND2 (N615, N602, N532);
buf BUF1 (N616, N604);
buf BUF1 (N617, N609);
and AND4 (N618, N608, N25, N158, N134);
xor XOR2 (N619, N616, N172);
not NOT1 (N620, N611);
nor NOR2 (N621, N620, N339);
xor XOR2 (N622, N618, N400);
nand NAND2 (N623, N613, N568);
and AND4 (N624, N619, N349, N521, N103);
xor XOR2 (N625, N615, N400);
buf BUF1 (N626, N617);
and AND3 (N627, N626, N474, N107);
buf BUF1 (N628, N599);
and AND4 (N629, N624, N126, N531, N82);
and AND3 (N630, N603, N589, N309);
xor XOR2 (N631, N628, N412);
buf BUF1 (N632, N630);
or OR4 (N633, N625, N234, N281, N379);
buf BUF1 (N634, N627);
buf BUF1 (N635, N610);
and AND2 (N636, N614, N227);
and AND4 (N637, N621, N362, N187, N385);
nand NAND3 (N638, N629, N145, N522);
and AND4 (N639, N638, N302, N81, N472);
or OR2 (N640, N632, N561);
buf BUF1 (N641, N631);
or OR2 (N642, N634, N298);
nand NAND2 (N643, N633, N187);
not NOT1 (N644, N642);
nor NOR3 (N645, N636, N288, N297);
or OR3 (N646, N623, N630, N128);
and AND2 (N647, N622, N586);
nor NOR4 (N648, N646, N384, N596, N618);
xor XOR2 (N649, N637, N190);
xor XOR2 (N650, N645, N386);
buf BUF1 (N651, N643);
and AND3 (N652, N651, N160, N627);
nand NAND3 (N653, N639, N14, N450);
nand NAND3 (N654, N640, N32, N444);
not NOT1 (N655, N649);
or OR2 (N656, N650, N302);
nand NAND2 (N657, N648, N381);
buf BUF1 (N658, N655);
not NOT1 (N659, N635);
nand NAND2 (N660, N647, N492);
nand NAND2 (N661, N653, N473);
not NOT1 (N662, N657);
or OR4 (N663, N654, N466, N163, N241);
buf BUF1 (N664, N662);
not NOT1 (N665, N664);
buf BUF1 (N666, N665);
buf BUF1 (N667, N660);
and AND3 (N668, N656, N369, N443);
nor NOR4 (N669, N644, N152, N231, N252);
xor XOR2 (N670, N663, N445);
nor NOR3 (N671, N669, N546, N22);
and AND2 (N672, N658, N240);
or OR2 (N673, N670, N52);
xor XOR2 (N674, N673, N382);
and AND4 (N675, N667, N297, N358, N650);
xor XOR2 (N676, N668, N378);
not NOT1 (N677, N672);
and AND2 (N678, N671, N347);
xor XOR2 (N679, N676, N179);
not NOT1 (N680, N679);
not NOT1 (N681, N659);
not NOT1 (N682, N666);
nor NOR4 (N683, N674, N372, N465, N594);
or OR2 (N684, N681, N535);
not NOT1 (N685, N680);
nor NOR2 (N686, N675, N249);
xor XOR2 (N687, N682, N64);
and AND4 (N688, N684, N659, N387, N260);
or OR4 (N689, N685, N271, N596, N82);
nor NOR3 (N690, N677, N177, N2);
xor XOR2 (N691, N689, N431);
or OR3 (N692, N661, N516, N196);
nor NOR3 (N693, N692, N409, N75);
not NOT1 (N694, N690);
and AND2 (N695, N694, N94);
nand NAND4 (N696, N686, N172, N481, N485);
not NOT1 (N697, N688);
nor NOR4 (N698, N691, N177, N652, N65);
buf BUF1 (N699, N98);
nor NOR4 (N700, N678, N288, N481, N337);
nor NOR3 (N701, N697, N389, N266);
buf BUF1 (N702, N699);
and AND4 (N703, N702, N76, N483, N373);
not NOT1 (N704, N696);
nor NOR4 (N705, N703, N627, N235, N652);
nor NOR4 (N706, N704, N665, N476, N58);
and AND4 (N707, N698, N200, N305, N202);
and AND2 (N708, N706, N536);
nor NOR4 (N709, N708, N163, N354, N98);
nor NOR4 (N710, N687, N32, N140, N575);
and AND4 (N711, N695, N355, N359, N690);
and AND3 (N712, N711, N589, N599);
buf BUF1 (N713, N700);
or OR2 (N714, N713, N209);
nor NOR2 (N715, N712, N683);
not NOT1 (N716, N297);
not NOT1 (N717, N705);
buf BUF1 (N718, N641);
nor NOR4 (N719, N710, N113, N336, N561);
not NOT1 (N720, N709);
nor NOR4 (N721, N701, N499, N393, N45);
buf BUF1 (N722, N717);
or OR2 (N723, N719, N705);
not NOT1 (N724, N718);
nand NAND2 (N725, N724, N470);
xor XOR2 (N726, N720, N373);
or OR3 (N727, N714, N188, N450);
not NOT1 (N728, N693);
or OR2 (N729, N727, N13);
nand NAND4 (N730, N722, N680, N169, N228);
xor XOR2 (N731, N715, N423);
xor XOR2 (N732, N707, N434);
nor NOR3 (N733, N728, N123, N620);
or OR2 (N734, N726, N642);
xor XOR2 (N735, N733, N688);
not NOT1 (N736, N734);
buf BUF1 (N737, N725);
and AND2 (N738, N731, N615);
not NOT1 (N739, N721);
buf BUF1 (N740, N729);
not NOT1 (N741, N737);
nor NOR2 (N742, N723, N310);
nand NAND2 (N743, N730, N608);
nor NOR4 (N744, N742, N715, N174, N499);
not NOT1 (N745, N732);
xor XOR2 (N746, N740, N536);
xor XOR2 (N747, N745, N15);
xor XOR2 (N748, N739, N23);
buf BUF1 (N749, N743);
xor XOR2 (N750, N716, N19);
buf BUF1 (N751, N746);
xor XOR2 (N752, N750, N425);
and AND4 (N753, N752, N255, N479, N739);
xor XOR2 (N754, N736, N617);
and AND2 (N755, N754, N519);
xor XOR2 (N756, N744, N139);
nand NAND2 (N757, N747, N233);
or OR2 (N758, N738, N383);
nor NOR3 (N759, N735, N696, N52);
not NOT1 (N760, N748);
xor XOR2 (N761, N758, N286);
nand NAND4 (N762, N761, N646, N666, N452);
not NOT1 (N763, N753);
nand NAND3 (N764, N759, N168, N62);
xor XOR2 (N765, N756, N71);
xor XOR2 (N766, N765, N539);
buf BUF1 (N767, N755);
nand NAND4 (N768, N766, N16, N516, N23);
or OR3 (N769, N764, N612, N204);
or OR3 (N770, N763, N644, N229);
xor XOR2 (N771, N751, N743);
xor XOR2 (N772, N760, N466);
and AND2 (N773, N772, N79);
or OR3 (N774, N762, N533, N459);
xor XOR2 (N775, N749, N377);
and AND3 (N776, N773, N443, N30);
nor NOR2 (N777, N771, N699);
nand NAND3 (N778, N741, N661, N577);
nor NOR4 (N779, N757, N600, N763, N671);
nand NAND4 (N780, N768, N366, N260, N621);
not NOT1 (N781, N769);
xor XOR2 (N782, N776, N594);
or OR4 (N783, N779, N158, N619, N638);
buf BUF1 (N784, N781);
xor XOR2 (N785, N777, N295);
xor XOR2 (N786, N785, N418);
nand NAND3 (N787, N783, N623, N579);
or OR2 (N788, N782, N351);
not NOT1 (N789, N767);
nand NAND4 (N790, N770, N780, N32, N347);
xor XOR2 (N791, N268, N348);
or OR2 (N792, N786, N364);
buf BUF1 (N793, N792);
not NOT1 (N794, N789);
buf BUF1 (N795, N788);
xor XOR2 (N796, N793, N173);
or OR3 (N797, N775, N126, N235);
and AND4 (N798, N797, N217, N78, N16);
nand NAND2 (N799, N790, N9);
and AND3 (N800, N778, N615, N537);
nor NOR3 (N801, N791, N558, N763);
not NOT1 (N802, N798);
nor NOR2 (N803, N799, N131);
or OR3 (N804, N803, N562, N632);
and AND3 (N805, N801, N588, N207);
or OR2 (N806, N774, N687);
nand NAND2 (N807, N804, N177);
buf BUF1 (N808, N805);
and AND3 (N809, N796, N461, N177);
not NOT1 (N810, N806);
xor XOR2 (N811, N784, N566);
or OR2 (N812, N794, N768);
not NOT1 (N813, N807);
nor NOR4 (N814, N795, N299, N121, N573);
xor XOR2 (N815, N802, N455);
buf BUF1 (N816, N800);
xor XOR2 (N817, N814, N593);
and AND2 (N818, N811, N314);
or OR2 (N819, N787, N386);
or OR4 (N820, N817, N497, N391, N683);
not NOT1 (N821, N813);
not NOT1 (N822, N818);
buf BUF1 (N823, N822);
nor NOR2 (N824, N816, N408);
xor XOR2 (N825, N812, N702);
not NOT1 (N826, N821);
or OR3 (N827, N810, N576, N281);
not NOT1 (N828, N825);
not NOT1 (N829, N824);
xor XOR2 (N830, N819, N789);
buf BUF1 (N831, N823);
buf BUF1 (N832, N829);
nand NAND2 (N833, N826, N728);
nand NAND2 (N834, N808, N541);
and AND3 (N835, N809, N348, N4);
nor NOR4 (N836, N827, N337, N242, N293);
not NOT1 (N837, N833);
and AND3 (N838, N830, N655, N697);
not NOT1 (N839, N831);
xor XOR2 (N840, N837, N627);
xor XOR2 (N841, N836, N81);
nand NAND3 (N842, N828, N680, N125);
xor XOR2 (N843, N834, N825);
nor NOR3 (N844, N820, N144, N701);
and AND4 (N845, N842, N87, N509, N579);
xor XOR2 (N846, N840, N306);
xor XOR2 (N847, N846, N358);
nor NOR2 (N848, N815, N395);
xor XOR2 (N849, N832, N294);
nand NAND2 (N850, N849, N60);
buf BUF1 (N851, N847);
buf BUF1 (N852, N851);
nand NAND3 (N853, N845, N351, N573);
not NOT1 (N854, N839);
nor NOR2 (N855, N853, N196);
and AND4 (N856, N843, N98, N94, N737);
and AND4 (N857, N835, N520, N711, N17);
nor NOR4 (N858, N856, N355, N502, N176);
or OR3 (N859, N857, N749, N237);
or OR2 (N860, N852, N68);
buf BUF1 (N861, N844);
not NOT1 (N862, N850);
not NOT1 (N863, N860);
xor XOR2 (N864, N861, N386);
xor XOR2 (N865, N859, N796);
not NOT1 (N866, N854);
not NOT1 (N867, N858);
xor XOR2 (N868, N838, N160);
xor XOR2 (N869, N855, N87);
and AND2 (N870, N863, N824);
buf BUF1 (N871, N862);
or OR3 (N872, N867, N144, N461);
buf BUF1 (N873, N868);
or OR4 (N874, N871, N633, N225, N586);
xor XOR2 (N875, N864, N90);
nand NAND4 (N876, N841, N234, N102, N710);
nor NOR4 (N877, N848, N2, N734, N124);
nor NOR3 (N878, N865, N634, N88);
not NOT1 (N879, N876);
xor XOR2 (N880, N873, N875);
nor NOR3 (N881, N166, N820, N196);
and AND2 (N882, N879, N224);
nor NOR2 (N883, N880, N624);
nand NAND2 (N884, N881, N871);
or OR2 (N885, N874, N817);
and AND4 (N886, N883, N605, N736, N879);
xor XOR2 (N887, N878, N670);
nand NAND4 (N888, N885, N45, N310, N169);
buf BUF1 (N889, N887);
nor NOR4 (N890, N872, N882, N204, N670);
or OR4 (N891, N87, N855, N349, N669);
nand NAND2 (N892, N889, N273);
and AND4 (N893, N890, N338, N341, N594);
xor XOR2 (N894, N866, N199);
or OR3 (N895, N891, N20, N112);
or OR4 (N896, N884, N444, N661, N835);
or OR4 (N897, N892, N296, N661, N303);
xor XOR2 (N898, N869, N619);
or OR4 (N899, N886, N59, N762, N339);
nor NOR2 (N900, N894, N114);
nand NAND3 (N901, N897, N465, N691);
not NOT1 (N902, N893);
or OR2 (N903, N898, N29);
xor XOR2 (N904, N901, N483);
nand NAND4 (N905, N899, N890, N722, N354);
nand NAND3 (N906, N870, N746, N456);
buf BUF1 (N907, N905);
or OR2 (N908, N888, N852);
xor XOR2 (N909, N907, N549);
nand NAND4 (N910, N906, N224, N551, N481);
and AND4 (N911, N910, N829, N877, N77);
or OR3 (N912, N418, N387, N226);
and AND4 (N913, N902, N241, N98, N678);
xor XOR2 (N914, N909, N211);
buf BUF1 (N915, N911);
nand NAND3 (N916, N913, N83, N588);
or OR3 (N917, N900, N613, N112);
or OR2 (N918, N912, N789);
xor XOR2 (N919, N917, N68);
buf BUF1 (N920, N903);
nand NAND2 (N921, N896, N245);
or OR3 (N922, N914, N76, N873);
and AND3 (N923, N920, N428, N533);
buf BUF1 (N924, N908);
nor NOR3 (N925, N915, N315, N123);
not NOT1 (N926, N918);
or OR2 (N927, N925, N195);
xor XOR2 (N928, N895, N730);
or OR3 (N929, N927, N840, N763);
and AND3 (N930, N904, N694, N283);
buf BUF1 (N931, N930);
nand NAND4 (N932, N916, N540, N446, N889);
nand NAND3 (N933, N921, N777, N596);
xor XOR2 (N934, N928, N226);
and AND2 (N935, N932, N399);
or OR4 (N936, N924, N845, N615, N921);
xor XOR2 (N937, N935, N732);
nor NOR3 (N938, N936, N547, N227);
and AND2 (N939, N934, N655);
or OR3 (N940, N933, N182, N595);
or OR2 (N941, N937, N568);
buf BUF1 (N942, N926);
nand NAND3 (N943, N940, N248, N315);
buf BUF1 (N944, N943);
xor XOR2 (N945, N938, N579);
xor XOR2 (N946, N942, N551);
not NOT1 (N947, N931);
xor XOR2 (N948, N947, N319);
buf BUF1 (N949, N948);
buf BUF1 (N950, N945);
buf BUF1 (N951, N929);
xor XOR2 (N952, N951, N325);
nand NAND3 (N953, N923, N182, N692);
xor XOR2 (N954, N939, N937);
not NOT1 (N955, N950);
not NOT1 (N956, N946);
xor XOR2 (N957, N955, N244);
or OR2 (N958, N944, N908);
or OR3 (N959, N952, N415, N247);
or OR3 (N960, N949, N83, N113);
and AND3 (N961, N922, N99, N842);
xor XOR2 (N962, N957, N373);
nor NOR2 (N963, N962, N936);
or OR4 (N964, N959, N809, N360, N215);
nor NOR2 (N965, N964, N579);
or OR4 (N966, N963, N588, N226, N676);
or OR2 (N967, N941, N107);
buf BUF1 (N968, N956);
buf BUF1 (N969, N954);
not NOT1 (N970, N967);
or OR3 (N971, N953, N238, N138);
or OR2 (N972, N958, N612);
xor XOR2 (N973, N969, N284);
and AND4 (N974, N971, N267, N959, N763);
and AND2 (N975, N968, N594);
not NOT1 (N976, N965);
and AND4 (N977, N973, N436, N569, N130);
nand NAND3 (N978, N972, N478, N173);
xor XOR2 (N979, N977, N375);
not NOT1 (N980, N970);
xor XOR2 (N981, N980, N457);
nor NOR2 (N982, N966, N333);
or OR3 (N983, N976, N322, N23);
buf BUF1 (N984, N961);
or OR4 (N985, N979, N840, N10, N55);
nand NAND2 (N986, N960, N482);
xor XOR2 (N987, N985, N606);
or OR4 (N988, N984, N248, N951, N12);
and AND4 (N989, N919, N152, N227, N689);
buf BUF1 (N990, N987);
or OR2 (N991, N989, N804);
or OR2 (N992, N975, N256);
not NOT1 (N993, N988);
or OR2 (N994, N991, N651);
or OR4 (N995, N992, N344, N220, N742);
nor NOR4 (N996, N982, N804, N519, N729);
nand NAND3 (N997, N996, N157, N935);
buf BUF1 (N998, N990);
not NOT1 (N999, N995);
not NOT1 (N1000, N999);
buf BUF1 (N1001, N997);
nor NOR2 (N1002, N993, N269);
nor NOR2 (N1003, N1000, N694);
xor XOR2 (N1004, N998, N72);
not NOT1 (N1005, N978);
and AND3 (N1006, N994, N369, N984);
not NOT1 (N1007, N986);
xor XOR2 (N1008, N1007, N574);
buf BUF1 (N1009, N974);
nor NOR2 (N1010, N1005, N766);
nand NAND3 (N1011, N983, N666, N18);
xor XOR2 (N1012, N1004, N354);
buf BUF1 (N1013, N1010);
nand NAND3 (N1014, N1013, N273, N214);
or OR4 (N1015, N1011, N116, N220, N121);
buf BUF1 (N1016, N1006);
and AND2 (N1017, N1012, N109);
buf BUF1 (N1018, N1001);
nor NOR4 (N1019, N1017, N328, N933, N764);
buf BUF1 (N1020, N1015);
nor NOR4 (N1021, N1002, N246, N550, N1008);
and AND2 (N1022, N639, N834);
buf BUF1 (N1023, N981);
nand NAND2 (N1024, N1018, N137);
buf BUF1 (N1025, N1019);
or OR2 (N1026, N1024, N785);
not NOT1 (N1027, N1003);
and AND2 (N1028, N1014, N189);
not NOT1 (N1029, N1026);
xor XOR2 (N1030, N1028, N719);
or OR2 (N1031, N1020, N37);
buf BUF1 (N1032, N1021);
nor NOR2 (N1033, N1030, N615);
not NOT1 (N1034, N1023);
buf BUF1 (N1035, N1032);
nor NOR2 (N1036, N1009, N189);
not NOT1 (N1037, N1034);
nor NOR4 (N1038, N1035, N200, N610, N747);
nor NOR3 (N1039, N1025, N662, N796);
not NOT1 (N1040, N1029);
not NOT1 (N1041, N1039);
buf BUF1 (N1042, N1041);
buf BUF1 (N1043, N1042);
xor XOR2 (N1044, N1040, N206);
not NOT1 (N1045, N1022);
xor XOR2 (N1046, N1036, N903);
xor XOR2 (N1047, N1043, N288);
xor XOR2 (N1048, N1016, N305);
nor NOR4 (N1049, N1031, N554, N102, N120);
and AND3 (N1050, N1033, N21, N833);
buf BUF1 (N1051, N1050);
buf BUF1 (N1052, N1046);
nor NOR2 (N1053, N1049, N282);
and AND3 (N1054, N1044, N174, N1022);
not NOT1 (N1055, N1037);
not NOT1 (N1056, N1027);
and AND2 (N1057, N1048, N403);
and AND2 (N1058, N1038, N249);
not NOT1 (N1059, N1058);
nor NOR3 (N1060, N1052, N1018, N399);
nor NOR3 (N1061, N1053, N352, N517);
not NOT1 (N1062, N1061);
buf BUF1 (N1063, N1055);
nand NAND3 (N1064, N1051, N746, N256);
buf BUF1 (N1065, N1054);
nor NOR3 (N1066, N1045, N402, N224);
buf BUF1 (N1067, N1047);
and AND3 (N1068, N1060, N768, N984);
xor XOR2 (N1069, N1063, N911);
nand NAND3 (N1070, N1065, N1027, N447);
and AND2 (N1071, N1057, N748);
xor XOR2 (N1072, N1069, N634);
xor XOR2 (N1073, N1066, N352);
or OR3 (N1074, N1064, N440, N770);
nand NAND3 (N1075, N1056, N985, N277);
and AND3 (N1076, N1067, N159, N744);
xor XOR2 (N1077, N1073, N270);
nor NOR3 (N1078, N1070, N381, N576);
not NOT1 (N1079, N1068);
nand NAND4 (N1080, N1072, N873, N294, N444);
nand NAND4 (N1081, N1076, N82, N1064, N862);
not NOT1 (N1082, N1059);
xor XOR2 (N1083, N1080, N626);
and AND3 (N1084, N1078, N778, N385);
xor XOR2 (N1085, N1077, N967);
nor NOR3 (N1086, N1082, N195, N515);
nor NOR3 (N1087, N1062, N496, N677);
buf BUF1 (N1088, N1083);
nor NOR4 (N1089, N1079, N1069, N422, N964);
buf BUF1 (N1090, N1081);
and AND2 (N1091, N1085, N118);
buf BUF1 (N1092, N1088);
and AND3 (N1093, N1071, N622, N246);
xor XOR2 (N1094, N1092, N655);
nand NAND3 (N1095, N1086, N538, N70);
and AND2 (N1096, N1089, N792);
nor NOR4 (N1097, N1095, N211, N308, N948);
xor XOR2 (N1098, N1093, N577);
or OR4 (N1099, N1074, N952, N718, N316);
nand NAND2 (N1100, N1099, N876);
nor NOR3 (N1101, N1075, N657, N16);
buf BUF1 (N1102, N1096);
not NOT1 (N1103, N1087);
not NOT1 (N1104, N1084);
not NOT1 (N1105, N1097);
buf BUF1 (N1106, N1091);
buf BUF1 (N1107, N1106);
buf BUF1 (N1108, N1107);
and AND3 (N1109, N1103, N46, N1072);
and AND4 (N1110, N1100, N642, N765, N192);
and AND2 (N1111, N1098, N1023);
xor XOR2 (N1112, N1110, N1067);
nor NOR4 (N1113, N1102, N206, N321, N864);
not NOT1 (N1114, N1109);
xor XOR2 (N1115, N1090, N874);
xor XOR2 (N1116, N1115, N1029);
nor NOR3 (N1117, N1114, N96, N242);
not NOT1 (N1118, N1111);
xor XOR2 (N1119, N1101, N918);
buf BUF1 (N1120, N1108);
nor NOR2 (N1121, N1113, N322);
xor XOR2 (N1122, N1104, N314);
nand NAND2 (N1123, N1119, N959);
not NOT1 (N1124, N1123);
and AND4 (N1125, N1120, N97, N923, N575);
xor XOR2 (N1126, N1117, N130);
or OR2 (N1127, N1125, N102);
xor XOR2 (N1128, N1105, N18);
xor XOR2 (N1129, N1116, N460);
nand NAND2 (N1130, N1094, N881);
xor XOR2 (N1131, N1122, N347);
and AND3 (N1132, N1129, N791, N692);
and AND2 (N1133, N1128, N1044);
and AND2 (N1134, N1130, N548);
nand NAND2 (N1135, N1124, N984);
not NOT1 (N1136, N1112);
or OR4 (N1137, N1136, N50, N969, N545);
not NOT1 (N1138, N1131);
not NOT1 (N1139, N1135);
xor XOR2 (N1140, N1138, N47);
not NOT1 (N1141, N1126);
and AND2 (N1142, N1133, N339);
not NOT1 (N1143, N1139);
nor NOR2 (N1144, N1132, N463);
xor XOR2 (N1145, N1144, N649);
and AND3 (N1146, N1141, N862, N990);
buf BUF1 (N1147, N1142);
or OR3 (N1148, N1140, N1064, N228);
nand NAND2 (N1149, N1118, N97);
and AND4 (N1150, N1149, N395, N688, N135);
nand NAND2 (N1151, N1143, N985);
nand NAND4 (N1152, N1121, N749, N31, N943);
not NOT1 (N1153, N1134);
nor NOR4 (N1154, N1150, N15, N323, N7);
nand NAND3 (N1155, N1146, N250, N483);
nor NOR4 (N1156, N1154, N1031, N1058, N561);
and AND4 (N1157, N1152, N1086, N1046, N1144);
not NOT1 (N1158, N1155);
buf BUF1 (N1159, N1158);
nor NOR2 (N1160, N1156, N143);
buf BUF1 (N1161, N1145);
buf BUF1 (N1162, N1160);
buf BUF1 (N1163, N1148);
not NOT1 (N1164, N1157);
or OR3 (N1165, N1137, N249, N159);
nand NAND2 (N1166, N1159, N1134);
nor NOR2 (N1167, N1162, N1116);
or OR4 (N1168, N1163, N28, N215, N16);
buf BUF1 (N1169, N1168);
nand NAND2 (N1170, N1147, N576);
xor XOR2 (N1171, N1169, N1014);
or OR3 (N1172, N1170, N1109, N538);
nor NOR2 (N1173, N1167, N569);
nor NOR3 (N1174, N1164, N538, N11);
nor NOR2 (N1175, N1165, N1119);
and AND2 (N1176, N1173, N889);
not NOT1 (N1177, N1151);
and AND3 (N1178, N1177, N345, N1018);
xor XOR2 (N1179, N1176, N206);
and AND2 (N1180, N1161, N1168);
xor XOR2 (N1181, N1172, N191);
nor NOR3 (N1182, N1153, N924, N785);
and AND3 (N1183, N1166, N1174, N195);
xor XOR2 (N1184, N806, N853);
not NOT1 (N1185, N1127);
not NOT1 (N1186, N1175);
or OR4 (N1187, N1183, N912, N634, N627);
nand NAND3 (N1188, N1187, N753, N1144);
or OR4 (N1189, N1180, N505, N139, N770);
not NOT1 (N1190, N1184);
buf BUF1 (N1191, N1185);
nor NOR4 (N1192, N1179, N205, N471, N534);
or OR3 (N1193, N1178, N1155, N1122);
not NOT1 (N1194, N1182);
or OR4 (N1195, N1191, N72, N438, N545);
and AND3 (N1196, N1181, N56, N676);
nor NOR4 (N1197, N1194, N213, N969, N831);
and AND3 (N1198, N1188, N44, N54);
nand NAND4 (N1199, N1195, N311, N166, N1056);
xor XOR2 (N1200, N1189, N1012);
nand NAND4 (N1201, N1192, N18, N420, N448);
nand NAND2 (N1202, N1196, N735);
or OR2 (N1203, N1171, N570);
buf BUF1 (N1204, N1202);
xor XOR2 (N1205, N1197, N1059);
and AND4 (N1206, N1205, N226, N812, N623);
or OR4 (N1207, N1204, N1167, N498, N873);
buf BUF1 (N1208, N1206);
buf BUF1 (N1209, N1200);
or OR2 (N1210, N1193, N873);
nand NAND2 (N1211, N1208, N826);
or OR4 (N1212, N1211, N136, N380, N782);
nor NOR3 (N1213, N1212, N461, N962);
not NOT1 (N1214, N1201);
nor NOR4 (N1215, N1199, N98, N1040, N364);
and AND4 (N1216, N1214, N159, N782, N174);
nand NAND2 (N1217, N1210, N888);
not NOT1 (N1218, N1217);
buf BUF1 (N1219, N1213);
nor NOR2 (N1220, N1215, N1204);
and AND2 (N1221, N1190, N1075);
and AND2 (N1222, N1219, N491);
not NOT1 (N1223, N1220);
not NOT1 (N1224, N1203);
xor XOR2 (N1225, N1218, N151);
or OR4 (N1226, N1186, N1128, N536, N951);
nor NOR2 (N1227, N1226, N1107);
and AND2 (N1228, N1221, N560);
xor XOR2 (N1229, N1223, N1110);
nand NAND4 (N1230, N1216, N1157, N925, N803);
nand NAND3 (N1231, N1222, N254, N1101);
nand NAND3 (N1232, N1198, N820, N417);
and AND2 (N1233, N1229, N343);
not NOT1 (N1234, N1230);
buf BUF1 (N1235, N1209);
not NOT1 (N1236, N1232);
or OR2 (N1237, N1233, N290);
or OR4 (N1238, N1235, N170, N626, N956);
xor XOR2 (N1239, N1237, N461);
and AND4 (N1240, N1239, N54, N842, N1071);
buf BUF1 (N1241, N1240);
not NOT1 (N1242, N1236);
xor XOR2 (N1243, N1234, N660);
nor NOR2 (N1244, N1228, N711);
and AND4 (N1245, N1244, N465, N755, N3);
buf BUF1 (N1246, N1245);
buf BUF1 (N1247, N1224);
nor NOR2 (N1248, N1243, N1243);
or OR4 (N1249, N1238, N1110, N960, N533);
xor XOR2 (N1250, N1227, N903);
xor XOR2 (N1251, N1207, N196);
and AND2 (N1252, N1247, N722);
or OR4 (N1253, N1251, N386, N72, N191);
or OR2 (N1254, N1253, N1225);
and AND4 (N1255, N1177, N1089, N1189, N925);
and AND3 (N1256, N1248, N349, N1251);
xor XOR2 (N1257, N1242, N878);
or OR4 (N1258, N1250, N928, N1196, N837);
buf BUF1 (N1259, N1258);
nand NAND3 (N1260, N1241, N1164, N742);
buf BUF1 (N1261, N1246);
nor NOR2 (N1262, N1256, N1101);
buf BUF1 (N1263, N1261);
and AND3 (N1264, N1257, N316, N1230);
nor NOR4 (N1265, N1260, N723, N549, N683);
buf BUF1 (N1266, N1255);
and AND2 (N1267, N1264, N516);
and AND3 (N1268, N1252, N1116, N1075);
nand NAND2 (N1269, N1231, N448);
nand NAND4 (N1270, N1268, N808, N1001, N362);
xor XOR2 (N1271, N1267, N826);
nand NAND3 (N1272, N1259, N288, N201);
buf BUF1 (N1273, N1272);
not NOT1 (N1274, N1273);
and AND2 (N1275, N1271, N4);
nor NOR4 (N1276, N1263, N1001, N863, N460);
or OR2 (N1277, N1266, N895);
nor NOR4 (N1278, N1270, N115, N236, N603);
buf BUF1 (N1279, N1265);
and AND2 (N1280, N1274, N474);
buf BUF1 (N1281, N1269);
nand NAND4 (N1282, N1254, N945, N114, N1074);
not NOT1 (N1283, N1249);
and AND4 (N1284, N1278, N679, N216, N989);
xor XOR2 (N1285, N1281, N1060);
and AND3 (N1286, N1280, N129, N76);
or OR4 (N1287, N1284, N767, N560, N367);
and AND2 (N1288, N1285, N752);
and AND3 (N1289, N1287, N496, N622);
nand NAND2 (N1290, N1288, N123);
nor NOR4 (N1291, N1279, N1272, N124, N1287);
buf BUF1 (N1292, N1286);
nor NOR4 (N1293, N1291, N500, N248, N983);
nand NAND3 (N1294, N1277, N34, N404);
or OR2 (N1295, N1294, N910);
nor NOR2 (N1296, N1262, N1029);
nor NOR2 (N1297, N1293, N677);
nand NAND4 (N1298, N1295, N737, N1208, N684);
nand NAND3 (N1299, N1297, N1189, N1091);
xor XOR2 (N1300, N1282, N152);
nand NAND3 (N1301, N1300, N462, N1131);
not NOT1 (N1302, N1292);
and AND4 (N1303, N1299, N10, N132, N395);
and AND3 (N1304, N1298, N893, N1214);
xor XOR2 (N1305, N1275, N864);
nor NOR3 (N1306, N1303, N457, N214);
buf BUF1 (N1307, N1305);
xor XOR2 (N1308, N1289, N65);
or OR2 (N1309, N1283, N1255);
buf BUF1 (N1310, N1302);
xor XOR2 (N1311, N1301, N274);
buf BUF1 (N1312, N1296);
or OR4 (N1313, N1276, N131, N683, N545);
or OR2 (N1314, N1306, N917);
nor NOR2 (N1315, N1313, N916);
not NOT1 (N1316, N1307);
nor NOR2 (N1317, N1316, N866);
or OR4 (N1318, N1315, N652, N753, N1256);
or OR2 (N1319, N1312, N1098);
nor NOR4 (N1320, N1318, N370, N1269, N157);
and AND4 (N1321, N1308, N542, N1128, N522);
xor XOR2 (N1322, N1319, N408);
or OR4 (N1323, N1290, N433, N148, N24);
nand NAND3 (N1324, N1317, N35, N1161);
or OR2 (N1325, N1324, N541);
buf BUF1 (N1326, N1311);
nand NAND3 (N1327, N1321, N799, N292);
nor NOR3 (N1328, N1327, N1024, N1140);
xor XOR2 (N1329, N1320, N854);
not NOT1 (N1330, N1328);
buf BUF1 (N1331, N1325);
buf BUF1 (N1332, N1314);
buf BUF1 (N1333, N1304);
not NOT1 (N1334, N1310);
nor NOR4 (N1335, N1332, N319, N684, N467);
and AND4 (N1336, N1331, N314, N1097, N878);
nor NOR4 (N1337, N1322, N317, N738, N332);
and AND3 (N1338, N1329, N1069, N1336);
not NOT1 (N1339, N1074);
buf BUF1 (N1340, N1309);
and AND4 (N1341, N1323, N299, N459, N1142);
xor XOR2 (N1342, N1335, N357);
buf BUF1 (N1343, N1341);
nor NOR4 (N1344, N1340, N1224, N321, N856);
not NOT1 (N1345, N1333);
not NOT1 (N1346, N1334);
or OR4 (N1347, N1330, N612, N948, N520);
not NOT1 (N1348, N1342);
or OR4 (N1349, N1348, N189, N63, N496);
buf BUF1 (N1350, N1338);
not NOT1 (N1351, N1346);
not NOT1 (N1352, N1349);
not NOT1 (N1353, N1350);
nand NAND2 (N1354, N1344, N818);
not NOT1 (N1355, N1337);
nor NOR4 (N1356, N1347, N1310, N621, N173);
and AND2 (N1357, N1352, N744);
nand NAND3 (N1358, N1356, N388, N600);
not NOT1 (N1359, N1353);
and AND3 (N1360, N1357, N1359, N1325);
nor NOR3 (N1361, N865, N671, N475);
or OR2 (N1362, N1345, N1024);
buf BUF1 (N1363, N1362);
not NOT1 (N1364, N1351);
not NOT1 (N1365, N1326);
and AND3 (N1366, N1363, N1085, N158);
nor NOR2 (N1367, N1366, N487);
xor XOR2 (N1368, N1343, N114);
xor XOR2 (N1369, N1367, N973);
buf BUF1 (N1370, N1339);
or OR4 (N1371, N1364, N760, N663, N593);
not NOT1 (N1372, N1371);
and AND4 (N1373, N1368, N505, N760, N531);
buf BUF1 (N1374, N1358);
and AND3 (N1375, N1370, N500, N1280);
xor XOR2 (N1376, N1355, N1353);
nor NOR2 (N1377, N1372, N1341);
buf BUF1 (N1378, N1376);
buf BUF1 (N1379, N1354);
not NOT1 (N1380, N1375);
xor XOR2 (N1381, N1361, N870);
buf BUF1 (N1382, N1365);
nor NOR4 (N1383, N1380, N467, N667, N867);
not NOT1 (N1384, N1379);
nor NOR4 (N1385, N1382, N667, N671, N654);
not NOT1 (N1386, N1381);
nand NAND4 (N1387, N1369, N1181, N382, N1365);
nand NAND4 (N1388, N1386, N876, N11, N1062);
xor XOR2 (N1389, N1373, N1193);
buf BUF1 (N1390, N1377);
nor NOR2 (N1391, N1388, N870);
xor XOR2 (N1392, N1374, N315);
not NOT1 (N1393, N1391);
buf BUF1 (N1394, N1387);
buf BUF1 (N1395, N1390);
nor NOR3 (N1396, N1384, N523, N889);
nor NOR2 (N1397, N1389, N194);
and AND2 (N1398, N1394, N128);
or OR2 (N1399, N1383, N1086);
buf BUF1 (N1400, N1360);
nand NAND3 (N1401, N1392, N1124, N453);
nand NAND3 (N1402, N1378, N1243, N1365);
or OR4 (N1403, N1400, N994, N108, N588);
nand NAND4 (N1404, N1385, N1336, N733, N703);
or OR2 (N1405, N1399, N727);
nor NOR3 (N1406, N1396, N1278, N1117);
buf BUF1 (N1407, N1403);
xor XOR2 (N1408, N1398, N1243);
xor XOR2 (N1409, N1402, N1006);
nand NAND3 (N1410, N1393, N1102, N480);
buf BUF1 (N1411, N1401);
not NOT1 (N1412, N1411);
xor XOR2 (N1413, N1404, N35);
buf BUF1 (N1414, N1407);
or OR4 (N1415, N1410, N556, N1259, N896);
buf BUF1 (N1416, N1405);
nand NAND4 (N1417, N1413, N111, N666, N171);
and AND3 (N1418, N1415, N795, N267);
not NOT1 (N1419, N1397);
nand NAND4 (N1420, N1412, N84, N444, N906);
or OR4 (N1421, N1409, N920, N119, N266);
not NOT1 (N1422, N1418);
and AND4 (N1423, N1421, N300, N382, N77);
or OR3 (N1424, N1417, N57, N555);
and AND4 (N1425, N1420, N493, N302, N654);
nor NOR3 (N1426, N1425, N993, N522);
or OR4 (N1427, N1406, N821, N195, N1184);
and AND2 (N1428, N1408, N356);
nand NAND3 (N1429, N1424, N561, N368);
nor NOR2 (N1430, N1423, N757);
not NOT1 (N1431, N1419);
nor NOR4 (N1432, N1422, N538, N1151, N1296);
xor XOR2 (N1433, N1416, N1122);
nand NAND2 (N1434, N1395, N173);
and AND2 (N1435, N1433, N883);
and AND2 (N1436, N1432, N1040);
or OR3 (N1437, N1434, N1248, N457);
or OR3 (N1438, N1436, N782, N338);
buf BUF1 (N1439, N1414);
or OR4 (N1440, N1426, N771, N1031, N751);
buf BUF1 (N1441, N1435);
nor NOR4 (N1442, N1438, N1133, N1046, N1104);
xor XOR2 (N1443, N1428, N467);
nand NAND3 (N1444, N1427, N104, N867);
nor NOR3 (N1445, N1444, N242, N1184);
or OR4 (N1446, N1439, N737, N819, N1271);
nand NAND3 (N1447, N1445, N210, N1132);
not NOT1 (N1448, N1429);
buf BUF1 (N1449, N1442);
xor XOR2 (N1450, N1431, N261);
nor NOR4 (N1451, N1450, N649, N13, N254);
buf BUF1 (N1452, N1446);
nand NAND2 (N1453, N1440, N607);
buf BUF1 (N1454, N1448);
nor NOR4 (N1455, N1441, N979, N1066, N62);
nor NOR2 (N1456, N1453, N435);
and AND4 (N1457, N1447, N913, N1040, N655);
and AND3 (N1458, N1437, N740, N1121);
buf BUF1 (N1459, N1449);
buf BUF1 (N1460, N1457);
or OR2 (N1461, N1454, N1380);
and AND2 (N1462, N1460, N1350);
nand NAND3 (N1463, N1459, N427, N1175);
buf BUF1 (N1464, N1430);
and AND3 (N1465, N1456, N724, N306);
not NOT1 (N1466, N1464);
or OR4 (N1467, N1451, N220, N464, N1312);
nand NAND2 (N1468, N1452, N140);
nor NOR2 (N1469, N1458, N833);
not NOT1 (N1470, N1463);
not NOT1 (N1471, N1462);
buf BUF1 (N1472, N1470);
or OR4 (N1473, N1468, N805, N826, N1259);
not NOT1 (N1474, N1469);
nand NAND4 (N1475, N1443, N942, N297, N720);
and AND2 (N1476, N1474, N510);
buf BUF1 (N1477, N1455);
or OR2 (N1478, N1472, N1105);
buf BUF1 (N1479, N1466);
nor NOR3 (N1480, N1476, N1432, N1182);
and AND4 (N1481, N1465, N813, N1079, N505);
or OR2 (N1482, N1475, N535);
not NOT1 (N1483, N1482);
or OR2 (N1484, N1461, N4);
or OR3 (N1485, N1478, N1042, N495);
xor XOR2 (N1486, N1479, N1365);
xor XOR2 (N1487, N1467, N793);
nor NOR2 (N1488, N1481, N358);
buf BUF1 (N1489, N1471);
buf BUF1 (N1490, N1477);
xor XOR2 (N1491, N1473, N638);
nand NAND3 (N1492, N1485, N1239, N428);
xor XOR2 (N1493, N1486, N354);
and AND2 (N1494, N1492, N497);
or OR4 (N1495, N1483, N864, N1014, N678);
not NOT1 (N1496, N1487);
not NOT1 (N1497, N1491);
and AND2 (N1498, N1496, N1041);
buf BUF1 (N1499, N1494);
and AND4 (N1500, N1493, N1018, N1086, N730);
xor XOR2 (N1501, N1495, N31);
not NOT1 (N1502, N1480);
buf BUF1 (N1503, N1488);
not NOT1 (N1504, N1501);
nand NAND4 (N1505, N1497, N400, N1393, N569);
nand NAND3 (N1506, N1484, N671, N448);
not NOT1 (N1507, N1506);
or OR2 (N1508, N1502, N699);
and AND2 (N1509, N1499, N605);
xor XOR2 (N1510, N1498, N373);
nor NOR4 (N1511, N1507, N1344, N899, N1375);
and AND2 (N1512, N1511, N827);
or OR3 (N1513, N1489, N258, N943);
and AND3 (N1514, N1513, N1203, N1133);
xor XOR2 (N1515, N1505, N1297);
xor XOR2 (N1516, N1504, N1314);
not NOT1 (N1517, N1514);
and AND2 (N1518, N1503, N149);
nor NOR3 (N1519, N1512, N1301, N477);
or OR3 (N1520, N1518, N1225, N278);
endmodule