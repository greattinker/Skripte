// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21;

output N511,N515,N508,N518,N513,N506,N520,N493,N507,N521;

xor XOR2 (N22, N5, N18);
and AND3 (N23, N13, N4, N21);
buf BUF1 (N24, N11);
buf BUF1 (N25, N20);
xor XOR2 (N26, N4, N2);
not NOT1 (N27, N17);
nand NAND4 (N28, N21, N13, N22, N19);
nor NOR3 (N29, N25, N19, N19);
not NOT1 (N30, N24);
xor XOR2 (N31, N17, N29);
buf BUF1 (N32, N6);
or OR2 (N33, N21, N23);
xor XOR2 (N34, N16, N7);
nand NAND2 (N35, N1, N19);
not NOT1 (N36, N24);
not NOT1 (N37, N36);
or OR3 (N38, N34, N37, N19);
buf BUF1 (N39, N30);
or OR3 (N40, N25, N5, N26);
nand NAND3 (N41, N15, N30, N11);
and AND4 (N42, N39, N2, N36, N2);
not NOT1 (N43, N31);
xor XOR2 (N44, N28, N4);
not NOT1 (N45, N42);
nor NOR2 (N46, N41, N7);
buf BUF1 (N47, N33);
or OR3 (N48, N46, N26, N44);
or OR2 (N49, N36, N40);
not NOT1 (N50, N47);
buf BUF1 (N51, N37);
xor XOR2 (N52, N43, N37);
buf BUF1 (N53, N49);
buf BUF1 (N54, N50);
or OR4 (N55, N52, N47, N52, N33);
or OR3 (N56, N38, N45, N55);
xor XOR2 (N57, N16, N26);
and AND4 (N58, N9, N12, N40, N29);
xor XOR2 (N59, N51, N3);
not NOT1 (N60, N59);
not NOT1 (N61, N32);
xor XOR2 (N62, N54, N21);
not NOT1 (N63, N57);
nor NOR3 (N64, N53, N63, N28);
not NOT1 (N65, N59);
nand NAND4 (N66, N58, N41, N61, N47);
and AND3 (N67, N60, N26, N53);
nor NOR3 (N68, N21, N59, N57);
nand NAND3 (N69, N68, N32, N33);
nand NAND2 (N70, N35, N48);
and AND3 (N71, N3, N46, N70);
and AND3 (N72, N37, N45, N58);
nor NOR4 (N73, N65, N39, N41, N48);
nor NOR4 (N74, N73, N58, N38, N8);
buf BUF1 (N75, N71);
not NOT1 (N76, N67);
buf BUF1 (N77, N74);
nor NOR2 (N78, N64, N51);
nand NAND4 (N79, N27, N49, N72, N60);
buf BUF1 (N80, N30);
xor XOR2 (N81, N77, N9);
xor XOR2 (N82, N78, N22);
xor XOR2 (N83, N66, N20);
or OR4 (N84, N56, N55, N3, N61);
or OR4 (N85, N76, N6, N41, N47);
nand NAND4 (N86, N80, N46, N29, N64);
and AND4 (N87, N79, N46, N26, N44);
or OR3 (N88, N85, N49, N1);
nor NOR2 (N89, N75, N10);
nor NOR4 (N90, N87, N29, N38, N11);
nor NOR2 (N91, N84, N84);
buf BUF1 (N92, N69);
and AND3 (N93, N90, N13, N20);
buf BUF1 (N94, N88);
nand NAND4 (N95, N94, N92, N25, N64);
not NOT1 (N96, N60);
and AND3 (N97, N93, N40, N67);
or OR3 (N98, N62, N90, N60);
buf BUF1 (N99, N91);
or OR4 (N100, N82, N5, N60, N66);
not NOT1 (N101, N81);
xor XOR2 (N102, N101, N61);
xor XOR2 (N103, N97, N90);
nand NAND2 (N104, N100, N22);
not NOT1 (N105, N96);
and AND4 (N106, N105, N95, N79, N34);
buf BUF1 (N107, N46);
or OR4 (N108, N102, N75, N101, N72);
xor XOR2 (N109, N103, N50);
buf BUF1 (N110, N99);
nand NAND2 (N111, N86, N106);
or OR3 (N112, N46, N76, N95);
or OR4 (N113, N111, N108, N30, N64);
nor NOR4 (N114, N31, N77, N97, N67);
not NOT1 (N115, N114);
buf BUF1 (N116, N112);
not NOT1 (N117, N110);
or OR4 (N118, N107, N85, N115, N90);
not NOT1 (N119, N95);
nor NOR2 (N120, N113, N94);
xor XOR2 (N121, N109, N60);
not NOT1 (N122, N119);
xor XOR2 (N123, N104, N85);
and AND2 (N124, N123, N86);
or OR3 (N125, N98, N71, N19);
and AND3 (N126, N83, N125, N94);
nor NOR2 (N127, N116, N81);
not NOT1 (N128, N29);
xor XOR2 (N129, N89, N70);
nand NAND2 (N130, N117, N96);
not NOT1 (N131, N124);
nand NAND2 (N132, N126, N53);
xor XOR2 (N133, N122, N102);
buf BUF1 (N134, N132);
buf BUF1 (N135, N130);
not NOT1 (N136, N135);
or OR3 (N137, N120, N50, N114);
and AND2 (N138, N128, N68);
not NOT1 (N139, N137);
xor XOR2 (N140, N118, N23);
xor XOR2 (N141, N133, N70);
or OR2 (N142, N141, N141);
not NOT1 (N143, N129);
xor XOR2 (N144, N143, N125);
buf BUF1 (N145, N121);
or OR3 (N146, N134, N48, N119);
and AND3 (N147, N140, N73, N82);
or OR3 (N148, N127, N29, N147);
and AND2 (N149, N104, N62);
nor NOR4 (N150, N138, N71, N54, N64);
nand NAND4 (N151, N146, N106, N79, N143);
nand NAND2 (N152, N142, N119);
xor XOR2 (N153, N150, N33);
xor XOR2 (N154, N148, N143);
nand NAND2 (N155, N151, N31);
or OR2 (N156, N154, N84);
nor NOR4 (N157, N155, N81, N119, N98);
or OR4 (N158, N153, N35, N80, N85);
nor NOR2 (N159, N145, N30);
not NOT1 (N160, N152);
or OR2 (N161, N160, N28);
and AND2 (N162, N156, N25);
nor NOR2 (N163, N161, N130);
xor XOR2 (N164, N136, N17);
xor XOR2 (N165, N131, N137);
not NOT1 (N166, N163);
and AND2 (N167, N158, N151);
or OR4 (N168, N159, N2, N123, N120);
xor XOR2 (N169, N144, N62);
xor XOR2 (N170, N139, N128);
nand NAND3 (N171, N164, N43, N118);
buf BUF1 (N172, N171);
and AND3 (N173, N166, N81, N85);
xor XOR2 (N174, N157, N40);
not NOT1 (N175, N170);
or OR2 (N176, N173, N71);
buf BUF1 (N177, N176);
buf BUF1 (N178, N165);
or OR2 (N179, N167, N148);
nand NAND3 (N180, N175, N76, N162);
nand NAND3 (N181, N47, N129, N1);
not NOT1 (N182, N172);
not NOT1 (N183, N174);
nand NAND4 (N184, N183, N18, N81, N171);
xor XOR2 (N185, N181, N121);
and AND2 (N186, N182, N38);
nand NAND4 (N187, N180, N79, N4, N47);
or OR3 (N188, N149, N148, N106);
nor NOR4 (N189, N188, N37, N136, N33);
and AND4 (N190, N187, N83, N111, N187);
not NOT1 (N191, N178);
or OR3 (N192, N179, N143, N62);
nand NAND2 (N193, N190, N156);
xor XOR2 (N194, N177, N48);
xor XOR2 (N195, N192, N183);
nor NOR3 (N196, N186, N128, N128);
or OR2 (N197, N169, N66);
xor XOR2 (N198, N196, N148);
nand NAND3 (N199, N197, N102, N61);
or OR4 (N200, N191, N9, N160, N199);
and AND2 (N201, N26, N186);
and AND4 (N202, N185, N162, N152, N161);
buf BUF1 (N203, N168);
xor XOR2 (N204, N200, N149);
or OR4 (N205, N201, N156, N65, N146);
nand NAND2 (N206, N205, N2);
and AND3 (N207, N194, N144, N50);
nand NAND3 (N208, N193, N120, N157);
not NOT1 (N209, N202);
not NOT1 (N210, N203);
and AND4 (N211, N208, N140, N36, N208);
or OR4 (N212, N209, N77, N189, N65);
buf BUF1 (N213, N108);
nor NOR3 (N214, N206, N86, N163);
and AND2 (N215, N204, N173);
nor NOR2 (N216, N214, N111);
nand NAND4 (N217, N207, N48, N141, N2);
nand NAND4 (N218, N212, N165, N28, N126);
nor NOR2 (N219, N211, N218);
not NOT1 (N220, N67);
nor NOR4 (N221, N220, N195, N62, N111);
nand NAND3 (N222, N22, N75, N181);
and AND4 (N223, N216, N36, N57, N189);
not NOT1 (N224, N223);
not NOT1 (N225, N217);
nor NOR2 (N226, N213, N204);
or OR2 (N227, N198, N14);
buf BUF1 (N228, N184);
nor NOR3 (N229, N215, N218, N205);
nand NAND2 (N230, N221, N58);
buf BUF1 (N231, N219);
nor NOR4 (N232, N227, N224, N99, N98);
or OR3 (N233, N148, N95, N170);
nand NAND4 (N234, N226, N156, N90, N187);
not NOT1 (N235, N228);
or OR2 (N236, N231, N67);
and AND2 (N237, N230, N5);
or OR4 (N238, N236, N135, N24, N230);
buf BUF1 (N239, N237);
or OR2 (N240, N233, N226);
or OR4 (N241, N234, N21, N138, N101);
nor NOR4 (N242, N238, N176, N44, N149);
nor NOR3 (N243, N222, N220, N176);
xor XOR2 (N244, N243, N133);
nor NOR4 (N245, N232, N203, N162, N216);
buf BUF1 (N246, N235);
nor NOR3 (N247, N229, N224, N14);
or OR2 (N248, N225, N159);
nand NAND3 (N249, N245, N103, N205);
buf BUF1 (N250, N240);
xor XOR2 (N251, N248, N200);
buf BUF1 (N252, N246);
buf BUF1 (N253, N250);
not NOT1 (N254, N252);
or OR3 (N255, N244, N169, N114);
or OR3 (N256, N253, N49, N155);
and AND3 (N257, N242, N175, N211);
not NOT1 (N258, N254);
nand NAND3 (N259, N256, N45, N212);
buf BUF1 (N260, N258);
or OR2 (N261, N257, N121);
and AND3 (N262, N210, N103, N29);
and AND3 (N263, N261, N196, N27);
xor XOR2 (N264, N247, N165);
not NOT1 (N265, N241);
and AND2 (N266, N255, N211);
and AND3 (N267, N251, N44, N42);
not NOT1 (N268, N265);
or OR4 (N269, N266, N118, N6, N124);
and AND4 (N270, N239, N204, N216, N224);
buf BUF1 (N271, N260);
or OR3 (N272, N271, N85, N256);
nand NAND2 (N273, N262, N67);
or OR2 (N274, N270, N73);
nand NAND2 (N275, N259, N119);
buf BUF1 (N276, N263);
buf BUF1 (N277, N273);
not NOT1 (N278, N249);
nand NAND2 (N279, N278, N176);
nor NOR2 (N280, N277, N42);
xor XOR2 (N281, N280, N51);
nor NOR3 (N282, N276, N154, N91);
xor XOR2 (N283, N279, N267);
nor NOR2 (N284, N236, N150);
buf BUF1 (N285, N275);
and AND4 (N286, N269, N115, N200, N119);
and AND2 (N287, N268, N181);
not NOT1 (N288, N286);
not NOT1 (N289, N288);
buf BUF1 (N290, N289);
buf BUF1 (N291, N281);
or OR2 (N292, N283, N193);
or OR4 (N293, N290, N25, N251, N3);
and AND4 (N294, N285, N211, N104, N258);
or OR2 (N295, N293, N161);
not NOT1 (N296, N292);
buf BUF1 (N297, N291);
buf BUF1 (N298, N297);
nor NOR4 (N299, N294, N129, N216, N247);
or OR3 (N300, N282, N76, N286);
nor NOR4 (N301, N296, N37, N227, N71);
buf BUF1 (N302, N284);
nor NOR2 (N303, N300, N236);
or OR4 (N304, N274, N224, N242, N244);
not NOT1 (N305, N301);
xor XOR2 (N306, N299, N224);
buf BUF1 (N307, N304);
or OR2 (N308, N287, N219);
or OR4 (N309, N306, N129, N118, N283);
and AND4 (N310, N302, N269, N1, N250);
nor NOR4 (N311, N307, N143, N49, N87);
nand NAND2 (N312, N298, N111);
xor XOR2 (N313, N264, N81);
nor NOR2 (N314, N309, N233);
nor NOR3 (N315, N312, N81, N126);
or OR4 (N316, N272, N196, N122, N284);
nand NAND3 (N317, N311, N206, N239);
xor XOR2 (N318, N313, N238);
xor XOR2 (N319, N317, N82);
nor NOR3 (N320, N303, N250, N188);
and AND2 (N321, N318, N71);
nor NOR3 (N322, N305, N242, N237);
nand NAND3 (N323, N295, N152, N79);
buf BUF1 (N324, N308);
or OR3 (N325, N323, N222, N227);
or OR3 (N326, N322, N116, N307);
and AND4 (N327, N325, N129, N144, N119);
nor NOR3 (N328, N321, N193, N271);
not NOT1 (N329, N315);
not NOT1 (N330, N319);
or OR3 (N331, N310, N322, N258);
buf BUF1 (N332, N320);
buf BUF1 (N333, N326);
nor NOR3 (N334, N329, N210, N281);
nand NAND4 (N335, N331, N245, N100, N296);
xor XOR2 (N336, N332, N153);
nor NOR2 (N337, N316, N275);
nand NAND2 (N338, N324, N325);
nor NOR2 (N339, N337, N283);
nor NOR3 (N340, N334, N335, N123);
and AND4 (N341, N2, N263, N134, N337);
nor NOR3 (N342, N333, N311, N337);
xor XOR2 (N343, N341, N32);
nor NOR2 (N344, N339, N261);
or OR2 (N345, N340, N261);
and AND3 (N346, N338, N160, N208);
not NOT1 (N347, N343);
not NOT1 (N348, N345);
nor NOR4 (N349, N347, N123, N78, N112);
nand NAND2 (N350, N349, N312);
or OR2 (N351, N328, N304);
and AND4 (N352, N330, N133, N285, N265);
or OR4 (N353, N342, N52, N203, N207);
nand NAND4 (N354, N314, N118, N277, N88);
nand NAND2 (N355, N351, N105);
or OR4 (N356, N350, N28, N1, N214);
nor NOR3 (N357, N348, N95, N19);
and AND3 (N358, N354, N309, N175);
and AND4 (N359, N358, N197, N152, N179);
xor XOR2 (N360, N357, N148);
or OR4 (N361, N356, N190, N86, N8);
and AND2 (N362, N336, N242);
or OR3 (N363, N361, N199, N228);
nand NAND2 (N364, N353, N87);
xor XOR2 (N365, N327, N344);
nor NOR4 (N366, N215, N238, N307, N88);
and AND4 (N367, N364, N266, N348, N312);
xor XOR2 (N368, N366, N56);
not NOT1 (N369, N367);
xor XOR2 (N370, N363, N169);
or OR4 (N371, N362, N5, N255, N113);
nor NOR4 (N372, N352, N221, N107, N110);
nor NOR3 (N373, N372, N239, N177);
not NOT1 (N374, N346);
and AND2 (N375, N369, N118);
xor XOR2 (N376, N355, N170);
nand NAND4 (N377, N360, N358, N170, N1);
buf BUF1 (N378, N374);
and AND3 (N379, N368, N10, N316);
nand NAND3 (N380, N377, N235, N329);
not NOT1 (N381, N375);
xor XOR2 (N382, N378, N171);
or OR4 (N383, N370, N121, N344, N314);
nor NOR4 (N384, N383, N329, N44, N365);
not NOT1 (N385, N380);
and AND2 (N386, N179, N256);
or OR3 (N387, N386, N202, N286);
nor NOR4 (N388, N379, N39, N105, N257);
nand NAND4 (N389, N385, N8, N368, N89);
and AND4 (N390, N382, N242, N19, N67);
not NOT1 (N391, N373);
or OR3 (N392, N391, N76, N171);
xor XOR2 (N393, N387, N373);
and AND3 (N394, N393, N6, N164);
xor XOR2 (N395, N389, N324);
nand NAND3 (N396, N376, N288, N328);
nand NAND4 (N397, N381, N124, N52, N301);
buf BUF1 (N398, N384);
not NOT1 (N399, N395);
xor XOR2 (N400, N371, N101);
xor XOR2 (N401, N398, N28);
and AND2 (N402, N397, N7);
nand NAND2 (N403, N399, N8);
xor XOR2 (N404, N396, N144);
xor XOR2 (N405, N401, N242);
nor NOR2 (N406, N400, N161);
not NOT1 (N407, N402);
and AND3 (N408, N359, N44, N25);
not NOT1 (N409, N390);
not NOT1 (N410, N405);
or OR2 (N411, N406, N46);
not NOT1 (N412, N407);
and AND2 (N413, N409, N34);
not NOT1 (N414, N388);
not NOT1 (N415, N404);
and AND2 (N416, N413, N253);
xor XOR2 (N417, N408, N331);
xor XOR2 (N418, N411, N213);
nand NAND4 (N419, N403, N223, N220, N211);
not NOT1 (N420, N418);
nand NAND2 (N421, N420, N210);
xor XOR2 (N422, N412, N67);
nand NAND2 (N423, N414, N58);
buf BUF1 (N424, N416);
xor XOR2 (N425, N410, N250);
nand NAND2 (N426, N423, N239);
buf BUF1 (N427, N424);
xor XOR2 (N428, N419, N23);
nor NOR2 (N429, N421, N173);
and AND4 (N430, N415, N155, N315, N252);
xor XOR2 (N431, N392, N424);
or OR4 (N432, N430, N340, N48, N332);
and AND2 (N433, N394, N77);
and AND4 (N434, N431, N123, N46, N175);
nor NOR3 (N435, N425, N11, N66);
xor XOR2 (N436, N432, N194);
and AND3 (N437, N428, N114, N307);
nor NOR4 (N438, N429, N123, N263, N326);
not NOT1 (N439, N427);
xor XOR2 (N440, N433, N118);
xor XOR2 (N441, N436, N343);
or OR3 (N442, N437, N415, N265);
buf BUF1 (N443, N422);
nor NOR3 (N444, N434, N55, N293);
or OR4 (N445, N439, N44, N66, N290);
nor NOR2 (N446, N417, N336);
not NOT1 (N447, N441);
buf BUF1 (N448, N442);
xor XOR2 (N449, N448, N414);
buf BUF1 (N450, N444);
or OR4 (N451, N440, N296, N212, N211);
xor XOR2 (N452, N435, N28);
nand NAND2 (N453, N443, N215);
buf BUF1 (N454, N449);
xor XOR2 (N455, N453, N411);
nand NAND3 (N456, N451, N41, N65);
or OR2 (N457, N446, N247);
buf BUF1 (N458, N450);
not NOT1 (N459, N438);
xor XOR2 (N460, N454, N438);
xor XOR2 (N461, N458, N3);
not NOT1 (N462, N447);
xor XOR2 (N463, N461, N252);
and AND2 (N464, N463, N15);
nand NAND4 (N465, N456, N237, N281, N161);
or OR3 (N466, N459, N143, N75);
or OR4 (N467, N464, N110, N263, N261);
xor XOR2 (N468, N426, N18);
nand NAND2 (N469, N466, N47);
buf BUF1 (N470, N468);
or OR2 (N471, N470, N330);
nand NAND4 (N472, N465, N195, N185, N347);
or OR3 (N473, N445, N463, N186);
buf BUF1 (N474, N455);
or OR3 (N475, N474, N429, N392);
nand NAND2 (N476, N472, N277);
xor XOR2 (N477, N471, N306);
buf BUF1 (N478, N462);
buf BUF1 (N479, N467);
xor XOR2 (N480, N478, N21);
xor XOR2 (N481, N452, N477);
nor NOR2 (N482, N382, N217);
nand NAND3 (N483, N469, N165, N379);
nand NAND2 (N484, N479, N440);
buf BUF1 (N485, N457);
and AND4 (N486, N483, N206, N245, N414);
nand NAND3 (N487, N485, N132, N383);
and AND3 (N488, N475, N132, N456);
or OR2 (N489, N484, N457);
and AND4 (N490, N480, N289, N367, N86);
nand NAND2 (N491, N482, N220);
nand NAND4 (N492, N486, N67, N470, N188);
nand NAND3 (N493, N492, N396, N314);
buf BUF1 (N494, N460);
buf BUF1 (N495, N476);
nand NAND2 (N496, N488, N389);
and AND4 (N497, N491, N437, N382, N336);
nor NOR2 (N498, N495, N323);
nor NOR4 (N499, N473, N383, N196, N321);
xor XOR2 (N500, N481, N114);
nor NOR2 (N501, N494, N131);
xor XOR2 (N502, N489, N483);
nand NAND3 (N503, N498, N282, N346);
nor NOR3 (N504, N487, N91, N432);
xor XOR2 (N505, N499, N40);
and AND2 (N506, N504, N103);
not NOT1 (N507, N497);
nand NAND2 (N508, N503, N231);
and AND4 (N509, N490, N233, N197, N124);
not NOT1 (N510, N509);
and AND2 (N511, N500, N477);
nor NOR4 (N512, N510, N393, N304, N463);
buf BUF1 (N513, N501);
nor NOR2 (N514, N505, N97);
or OR2 (N515, N496, N60);
nor NOR3 (N516, N502, N462, N97);
nor NOR2 (N517, N512, N378);
xor XOR2 (N518, N516, N447);
not NOT1 (N519, N514);
buf BUF1 (N520, N517);
nand NAND2 (N521, N519, N276);
endmodule