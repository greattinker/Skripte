// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22;

output N3215,N3219,N3221,N3213,N3208,N3218,N3220,N3205,N3216,N3222;

buf BUF1 (N23, N3);
nand NAND2 (N24, N20, N7);
or OR4 (N25, N13, N1, N8, N16);
xor XOR2 (N26, N18, N13);
xor XOR2 (N27, N8, N21);
or OR2 (N28, N17, N19);
nand NAND2 (N29, N15, N22);
buf BUF1 (N30, N7);
nor NOR2 (N31, N2, N24);
xor XOR2 (N32, N12, N2);
or OR2 (N33, N10, N26);
and AND3 (N34, N24, N17, N4);
buf BUF1 (N35, N29);
xor XOR2 (N36, N35, N2);
and AND3 (N37, N33, N19, N7);
nand NAND2 (N38, N31, N14);
or OR2 (N39, N23, N38);
not NOT1 (N40, N35);
or OR4 (N41, N27, N33, N4, N19);
nor NOR4 (N42, N40, N36, N34, N19);
nor NOR3 (N43, N26, N10, N9);
or OR2 (N44, N11, N24);
xor XOR2 (N45, N43, N28);
nor NOR2 (N46, N3, N2);
nor NOR2 (N47, N39, N5);
not NOT1 (N48, N42);
buf BUF1 (N49, N48);
nand NAND3 (N50, N46, N40, N39);
and AND3 (N51, N30, N2, N1);
nand NAND3 (N52, N49, N7, N3);
not NOT1 (N53, N47);
not NOT1 (N54, N53);
buf BUF1 (N55, N44);
and AND2 (N56, N45, N40);
nor NOR4 (N57, N50, N18, N54, N26);
buf BUF1 (N58, N50);
and AND2 (N59, N56, N29);
or OR3 (N60, N55, N7, N26);
or OR3 (N61, N59, N32, N17);
buf BUF1 (N62, N24);
not NOT1 (N63, N57);
nor NOR2 (N64, N61, N36);
not NOT1 (N65, N51);
nand NAND4 (N66, N63, N13, N19, N12);
or OR3 (N67, N60, N59, N47);
nor NOR4 (N68, N64, N51, N55, N12);
nand NAND4 (N69, N58, N65, N31, N63);
xor XOR2 (N70, N53, N32);
not NOT1 (N71, N67);
nand NAND3 (N72, N69, N49, N53);
nand NAND4 (N73, N71, N42, N58, N65);
nor NOR2 (N74, N52, N41);
nand NAND4 (N75, N4, N34, N57, N42);
buf BUF1 (N76, N37);
nor NOR2 (N77, N73, N56);
or OR2 (N78, N76, N74);
buf BUF1 (N79, N14);
or OR4 (N80, N79, N34, N5, N14);
xor XOR2 (N81, N77, N50);
and AND2 (N82, N75, N6);
not NOT1 (N83, N81);
buf BUF1 (N84, N82);
xor XOR2 (N85, N68, N52);
nor NOR2 (N86, N83, N57);
nand NAND2 (N87, N84, N10);
xor XOR2 (N88, N85, N53);
buf BUF1 (N89, N25);
xor XOR2 (N90, N89, N60);
not NOT1 (N91, N87);
nor NOR3 (N92, N90, N79, N66);
nor NOR2 (N93, N12, N68);
nor NOR2 (N94, N86, N90);
xor XOR2 (N95, N72, N57);
not NOT1 (N96, N92);
buf BUF1 (N97, N80);
nand NAND3 (N98, N91, N29, N85);
and AND2 (N99, N70, N16);
or OR3 (N100, N95, N75, N4);
not NOT1 (N101, N99);
xor XOR2 (N102, N88, N3);
or OR4 (N103, N96, N44, N94, N93);
xor XOR2 (N104, N65, N41);
nor NOR3 (N105, N25, N89, N83);
nor NOR2 (N106, N102, N8);
or OR4 (N107, N101, N64, N74, N84);
nor NOR3 (N108, N107, N85, N94);
nand NAND3 (N109, N104, N95, N17);
and AND4 (N110, N78, N20, N84, N82);
not NOT1 (N111, N100);
and AND2 (N112, N97, N89);
or OR3 (N113, N111, N30, N83);
or OR4 (N114, N98, N37, N16, N43);
xor XOR2 (N115, N108, N88);
not NOT1 (N116, N105);
not NOT1 (N117, N62);
and AND4 (N118, N114, N74, N99, N1);
xor XOR2 (N119, N110, N8);
buf BUF1 (N120, N115);
or OR3 (N121, N109, N72, N48);
nand NAND3 (N122, N120, N28, N54);
buf BUF1 (N123, N116);
buf BUF1 (N124, N121);
xor XOR2 (N125, N106, N28);
not NOT1 (N126, N112);
not NOT1 (N127, N119);
xor XOR2 (N128, N126, N79);
and AND4 (N129, N127, N94, N84, N76);
nor NOR2 (N130, N128, N117);
or OR2 (N131, N127, N15);
nand NAND4 (N132, N125, N38, N71, N75);
or OR3 (N133, N132, N59, N78);
not NOT1 (N134, N123);
xor XOR2 (N135, N134, N97);
buf BUF1 (N136, N118);
nand NAND4 (N137, N136, N116, N103, N16);
and AND4 (N138, N102, N2, N55, N4);
buf BUF1 (N139, N113);
nor NOR2 (N140, N135, N57);
buf BUF1 (N141, N140);
and AND2 (N142, N122, N15);
not NOT1 (N143, N133);
nand NAND3 (N144, N141, N77, N12);
nor NOR2 (N145, N129, N23);
and AND4 (N146, N138, N138, N98, N72);
not NOT1 (N147, N124);
and AND3 (N148, N146, N24, N132);
nor NOR4 (N149, N148, N66, N95, N45);
xor XOR2 (N150, N137, N84);
nand NAND2 (N151, N139, N86);
xor XOR2 (N152, N130, N54);
and AND4 (N153, N152, N28, N147, N110);
xor XOR2 (N154, N40, N146);
xor XOR2 (N155, N143, N89);
or OR2 (N156, N155, N10);
or OR2 (N157, N145, N95);
xor XOR2 (N158, N157, N12);
not NOT1 (N159, N156);
xor XOR2 (N160, N144, N33);
buf BUF1 (N161, N158);
nand NAND2 (N162, N151, N158);
nand NAND4 (N163, N159, N124, N51, N143);
xor XOR2 (N164, N154, N129);
nand NAND2 (N165, N164, N55);
buf BUF1 (N166, N165);
and AND3 (N167, N131, N163, N119);
xor XOR2 (N168, N28, N101);
or OR4 (N169, N153, N84, N140, N154);
xor XOR2 (N170, N167, N94);
nor NOR4 (N171, N142, N103, N96, N71);
buf BUF1 (N172, N169);
buf BUF1 (N173, N170);
xor XOR2 (N174, N168, N161);
xor XOR2 (N175, N133, N96);
and AND3 (N176, N166, N71, N20);
not NOT1 (N177, N175);
or OR2 (N178, N162, N42);
xor XOR2 (N179, N176, N38);
xor XOR2 (N180, N171, N177);
xor XOR2 (N181, N139, N43);
xor XOR2 (N182, N179, N127);
or OR2 (N183, N174, N7);
and AND3 (N184, N178, N126, N110);
nor NOR2 (N185, N181, N48);
buf BUF1 (N186, N172);
and AND3 (N187, N182, N94, N124);
nor NOR4 (N188, N150, N177, N79, N87);
nand NAND4 (N189, N180, N124, N133, N26);
or OR2 (N190, N183, N87);
not NOT1 (N191, N184);
nand NAND4 (N192, N190, N182, N120, N76);
nand NAND2 (N193, N149, N144);
and AND4 (N194, N185, N152, N18, N163);
nor NOR4 (N195, N193, N134, N113, N129);
not NOT1 (N196, N173);
xor XOR2 (N197, N196, N89);
or OR3 (N198, N195, N20, N123);
nand NAND3 (N199, N191, N58, N180);
not NOT1 (N200, N188);
nor NOR4 (N201, N197, N176, N177, N103);
nand NAND4 (N202, N201, N79, N187, N62);
buf BUF1 (N203, N153);
nand NAND2 (N204, N194, N112);
xor XOR2 (N205, N189, N20);
and AND2 (N206, N202, N71);
nand NAND2 (N207, N198, N161);
xor XOR2 (N208, N160, N3);
not NOT1 (N209, N203);
buf BUF1 (N210, N206);
not NOT1 (N211, N186);
or OR2 (N212, N200, N61);
xor XOR2 (N213, N209, N119);
and AND4 (N214, N199, N29, N79, N17);
not NOT1 (N215, N210);
xor XOR2 (N216, N211, N188);
xor XOR2 (N217, N213, N90);
nand NAND3 (N218, N205, N22, N34);
nor NOR3 (N219, N204, N166, N183);
nor NOR3 (N220, N217, N12, N156);
nor NOR2 (N221, N219, N44);
not NOT1 (N222, N207);
nor NOR3 (N223, N220, N202, N114);
not NOT1 (N224, N212);
nand NAND2 (N225, N192, N67);
or OR2 (N226, N222, N28);
buf BUF1 (N227, N214);
and AND2 (N228, N226, N71);
and AND3 (N229, N215, N223, N30);
buf BUF1 (N230, N23);
buf BUF1 (N231, N224);
buf BUF1 (N232, N227);
or OR2 (N233, N208, N90);
xor XOR2 (N234, N228, N190);
and AND2 (N235, N229, N180);
not NOT1 (N236, N230);
nor NOR2 (N237, N234, N232);
nand NAND3 (N238, N209, N27, N34);
buf BUF1 (N239, N237);
and AND4 (N240, N236, N135, N192, N96);
and AND4 (N241, N231, N212, N217, N167);
and AND3 (N242, N225, N63, N113);
nand NAND4 (N243, N235, N97, N51, N46);
not NOT1 (N244, N242);
nor NOR4 (N245, N239, N158, N199, N132);
nand NAND3 (N246, N243, N153, N36);
and AND4 (N247, N221, N156, N136, N233);
or OR2 (N248, N237, N198);
buf BUF1 (N249, N246);
nand NAND4 (N250, N241, N42, N226, N176);
not NOT1 (N251, N245);
not NOT1 (N252, N244);
or OR3 (N253, N238, N176, N47);
nand NAND3 (N254, N251, N248, N110);
not NOT1 (N255, N82);
nand NAND2 (N256, N249, N80);
and AND3 (N257, N252, N147, N233);
or OR3 (N258, N255, N136, N48);
nor NOR2 (N259, N218, N37);
xor XOR2 (N260, N259, N245);
nand NAND3 (N261, N216, N63, N177);
nor NOR2 (N262, N247, N171);
and AND3 (N263, N261, N164, N56);
and AND4 (N264, N257, N17, N228, N35);
nor NOR2 (N265, N254, N139);
and AND2 (N266, N256, N201);
nor NOR2 (N267, N240, N22);
nor NOR4 (N268, N250, N128, N205, N260);
not NOT1 (N269, N152);
nor NOR3 (N270, N263, N91, N55);
buf BUF1 (N271, N269);
buf BUF1 (N272, N266);
xor XOR2 (N273, N265, N159);
nor NOR4 (N274, N253, N13, N88, N64);
buf BUF1 (N275, N267);
nor NOR4 (N276, N275, N121, N159, N231);
xor XOR2 (N277, N268, N107);
and AND2 (N278, N264, N265);
xor XOR2 (N279, N278, N198);
nand NAND2 (N280, N277, N123);
or OR2 (N281, N272, N272);
nor NOR2 (N282, N276, N26);
not NOT1 (N283, N271);
and AND2 (N284, N262, N189);
or OR4 (N285, N280, N51, N233, N8);
not NOT1 (N286, N285);
nor NOR3 (N287, N281, N53, N40);
not NOT1 (N288, N258);
nor NOR4 (N289, N288, N124, N233, N242);
not NOT1 (N290, N286);
buf BUF1 (N291, N274);
and AND4 (N292, N270, N281, N251, N241);
or OR3 (N293, N284, N281, N231);
and AND3 (N294, N287, N126, N255);
nor NOR3 (N295, N293, N266, N44);
or OR2 (N296, N279, N87);
xor XOR2 (N297, N294, N129);
not NOT1 (N298, N295);
nor NOR3 (N299, N291, N235, N167);
nor NOR4 (N300, N298, N215, N45, N60);
buf BUF1 (N301, N297);
nand NAND3 (N302, N301, N6, N269);
nand NAND4 (N303, N292, N246, N71, N17);
not NOT1 (N304, N282);
and AND4 (N305, N290, N236, N118, N70);
or OR4 (N306, N289, N261, N146, N262);
or OR4 (N307, N306, N199, N206, N288);
nand NAND4 (N308, N273, N295, N261, N94);
buf BUF1 (N309, N300);
nand NAND4 (N310, N307, N266, N297, N75);
or OR2 (N311, N305, N136);
buf BUF1 (N312, N299);
not NOT1 (N313, N310);
nand NAND3 (N314, N309, N19, N232);
buf BUF1 (N315, N314);
not NOT1 (N316, N312);
or OR4 (N317, N302, N155, N42, N210);
xor XOR2 (N318, N303, N297);
not NOT1 (N319, N311);
nand NAND3 (N320, N296, N140, N81);
or OR2 (N321, N317, N225);
buf BUF1 (N322, N308);
buf BUF1 (N323, N321);
nor NOR3 (N324, N322, N37, N125);
not NOT1 (N325, N323);
xor XOR2 (N326, N316, N201);
xor XOR2 (N327, N320, N2);
buf BUF1 (N328, N315);
nand NAND2 (N329, N324, N199);
and AND3 (N330, N318, N74, N290);
buf BUF1 (N331, N283);
not NOT1 (N332, N327);
xor XOR2 (N333, N319, N65);
buf BUF1 (N334, N332);
or OR4 (N335, N313, N23, N31, N37);
not NOT1 (N336, N326);
xor XOR2 (N337, N331, N71);
nor NOR2 (N338, N325, N228);
xor XOR2 (N339, N330, N267);
nand NAND2 (N340, N337, N293);
nand NAND2 (N341, N304, N180);
nor NOR2 (N342, N338, N259);
not NOT1 (N343, N328);
and AND4 (N344, N329, N193, N268, N15);
nor NOR4 (N345, N342, N253, N102, N186);
nand NAND4 (N346, N345, N336, N200, N221);
xor XOR2 (N347, N71, N36);
and AND2 (N348, N333, N201);
and AND2 (N349, N346, N80);
buf BUF1 (N350, N334);
or OR4 (N351, N349, N339, N170, N222);
not NOT1 (N352, N296);
and AND3 (N353, N343, N99, N347);
xor XOR2 (N354, N44, N234);
or OR4 (N355, N351, N343, N347, N111);
nor NOR4 (N356, N344, N75, N280, N314);
nand NAND4 (N357, N356, N118, N339, N40);
nor NOR4 (N358, N354, N183, N131, N280);
nor NOR2 (N359, N352, N330);
nand NAND4 (N360, N341, N201, N88, N64);
or OR4 (N361, N355, N303, N36, N184);
xor XOR2 (N362, N335, N275);
and AND2 (N363, N359, N230);
or OR4 (N364, N340, N110, N126, N42);
or OR2 (N365, N363, N331);
buf BUF1 (N366, N350);
nor NOR3 (N367, N366, N254, N254);
or OR2 (N368, N358, N310);
not NOT1 (N369, N360);
nand NAND3 (N370, N368, N24, N21);
and AND4 (N371, N367, N309, N138, N252);
not NOT1 (N372, N348);
and AND3 (N373, N357, N134, N231);
not NOT1 (N374, N373);
nor NOR4 (N375, N370, N2, N123, N29);
nand NAND4 (N376, N369, N192, N189, N353);
buf BUF1 (N377, N92);
not NOT1 (N378, N364);
not NOT1 (N379, N372);
or OR3 (N380, N376, N290, N315);
buf BUF1 (N381, N377);
or OR4 (N382, N374, N50, N110, N156);
and AND4 (N383, N379, N179, N48, N334);
nand NAND2 (N384, N383, N3);
xor XOR2 (N385, N375, N367);
or OR2 (N386, N380, N341);
not NOT1 (N387, N361);
nor NOR3 (N388, N362, N107, N124);
or OR2 (N389, N381, N365);
or OR4 (N390, N379, N216, N88, N243);
xor XOR2 (N391, N390, N228);
nor NOR2 (N392, N385, N374);
not NOT1 (N393, N392);
not NOT1 (N394, N382);
and AND4 (N395, N384, N154, N226, N296);
nand NAND4 (N396, N386, N116, N51, N242);
xor XOR2 (N397, N387, N48);
nor NOR3 (N398, N395, N152, N244);
nor NOR3 (N399, N378, N21, N236);
nand NAND2 (N400, N371, N240);
nor NOR2 (N401, N396, N275);
not NOT1 (N402, N393);
not NOT1 (N403, N391);
not NOT1 (N404, N389);
nor NOR4 (N405, N402, N99, N166, N356);
not NOT1 (N406, N405);
xor XOR2 (N407, N399, N240);
buf BUF1 (N408, N406);
or OR2 (N409, N407, N251);
or OR3 (N410, N403, N279, N19);
nand NAND3 (N411, N400, N334, N373);
buf BUF1 (N412, N410);
buf BUF1 (N413, N398);
or OR3 (N414, N397, N378, N21);
xor XOR2 (N415, N412, N70);
not NOT1 (N416, N404);
nand NAND3 (N417, N409, N404, N124);
nor NOR4 (N418, N415, N106, N350, N162);
nor NOR3 (N419, N408, N251, N178);
not NOT1 (N420, N418);
nand NAND3 (N421, N411, N218, N206);
buf BUF1 (N422, N413);
and AND3 (N423, N422, N363, N187);
or OR2 (N424, N416, N421);
not NOT1 (N425, N297);
xor XOR2 (N426, N388, N184);
nand NAND3 (N427, N394, N191, N387);
and AND2 (N428, N414, N394);
nand NAND4 (N429, N423, N212, N276, N278);
buf BUF1 (N430, N428);
or OR2 (N431, N429, N171);
nor NOR2 (N432, N420, N82);
nand NAND4 (N433, N431, N190, N20, N249);
nor NOR4 (N434, N426, N408, N151, N140);
nor NOR4 (N435, N419, N110, N180, N62);
or OR2 (N436, N427, N417);
or OR4 (N437, N155, N66, N213, N20);
nand NAND4 (N438, N425, N407, N124, N369);
nand NAND2 (N439, N432, N302);
nor NOR2 (N440, N439, N392);
buf BUF1 (N441, N436);
nand NAND2 (N442, N433, N135);
nand NAND4 (N443, N442, N305, N434, N51);
nor NOR3 (N444, N206, N262, N313);
xor XOR2 (N445, N443, N218);
or OR3 (N446, N401, N110, N150);
and AND3 (N447, N435, N152, N413);
nor NOR3 (N448, N440, N391, N239);
nor NOR2 (N449, N444, N11);
xor XOR2 (N450, N447, N327);
xor XOR2 (N451, N445, N394);
not NOT1 (N452, N437);
nor NOR3 (N453, N424, N216, N26);
not NOT1 (N454, N451);
not NOT1 (N455, N438);
nor NOR3 (N456, N441, N417, N418);
buf BUF1 (N457, N452);
not NOT1 (N458, N448);
buf BUF1 (N459, N454);
xor XOR2 (N460, N456, N192);
nor NOR4 (N461, N460, N430, N221, N178);
not NOT1 (N462, N107);
or OR3 (N463, N450, N299, N157);
nor NOR4 (N464, N446, N428, N184, N255);
xor XOR2 (N465, N457, N174);
nor NOR3 (N466, N453, N355, N1);
nand NAND4 (N467, N455, N131, N303, N215);
nand NAND3 (N468, N462, N250, N33);
not NOT1 (N469, N459);
nand NAND2 (N470, N449, N413);
and AND3 (N471, N461, N234, N18);
not NOT1 (N472, N465);
and AND4 (N473, N469, N469, N449, N242);
not NOT1 (N474, N458);
or OR3 (N475, N474, N270, N343);
buf BUF1 (N476, N472);
or OR2 (N477, N471, N436);
nor NOR3 (N478, N477, N238, N37);
xor XOR2 (N479, N468, N17);
and AND3 (N480, N466, N344, N389);
and AND4 (N481, N479, N142, N97, N9);
not NOT1 (N482, N463);
or OR3 (N483, N475, N333, N469);
and AND3 (N484, N480, N377, N419);
buf BUF1 (N485, N483);
or OR3 (N486, N476, N141, N434);
not NOT1 (N487, N478);
nor NOR4 (N488, N470, N450, N213, N169);
or OR3 (N489, N486, N408, N404);
xor XOR2 (N490, N485, N289);
buf BUF1 (N491, N490);
nand NAND2 (N492, N487, N146);
buf BUF1 (N493, N491);
buf BUF1 (N494, N492);
xor XOR2 (N495, N489, N396);
nand NAND2 (N496, N464, N261);
or OR2 (N497, N495, N430);
nor NOR2 (N498, N482, N466);
xor XOR2 (N499, N467, N427);
or OR2 (N500, N496, N284);
and AND4 (N501, N498, N442, N32, N474);
not NOT1 (N502, N493);
and AND2 (N503, N494, N392);
xor XOR2 (N504, N484, N3);
nor NOR4 (N505, N502, N138, N463, N128);
buf BUF1 (N506, N500);
or OR3 (N507, N481, N82, N275);
or OR3 (N508, N505, N353, N57);
nor NOR4 (N509, N504, N308, N361, N152);
not NOT1 (N510, N501);
nand NAND2 (N511, N506, N226);
and AND3 (N512, N499, N193, N298);
xor XOR2 (N513, N512, N450);
or OR3 (N514, N513, N259, N52);
not NOT1 (N515, N509);
not NOT1 (N516, N508);
or OR4 (N517, N497, N443, N270, N260);
nor NOR3 (N518, N516, N445, N152);
buf BUF1 (N519, N510);
and AND3 (N520, N519, N146, N21);
xor XOR2 (N521, N517, N303);
not NOT1 (N522, N521);
nor NOR2 (N523, N473, N265);
nand NAND2 (N524, N520, N278);
xor XOR2 (N525, N488, N505);
buf BUF1 (N526, N522);
nand NAND3 (N527, N525, N20, N411);
buf BUF1 (N528, N507);
not NOT1 (N529, N518);
xor XOR2 (N530, N526, N260);
nor NOR2 (N531, N515, N258);
xor XOR2 (N532, N503, N423);
buf BUF1 (N533, N532);
not NOT1 (N534, N528);
not NOT1 (N535, N514);
or OR4 (N536, N531, N376, N39, N437);
nor NOR4 (N537, N527, N341, N326, N327);
and AND2 (N538, N530, N227);
nor NOR2 (N539, N538, N493);
or OR2 (N540, N511, N17);
buf BUF1 (N541, N534);
xor XOR2 (N542, N524, N290);
buf BUF1 (N543, N529);
buf BUF1 (N544, N540);
buf BUF1 (N545, N523);
nand NAND2 (N546, N542, N87);
or OR2 (N547, N535, N172);
xor XOR2 (N548, N547, N497);
and AND3 (N549, N548, N547, N401);
xor XOR2 (N550, N543, N100);
nor NOR2 (N551, N533, N76);
or OR2 (N552, N549, N130);
or OR2 (N553, N537, N159);
or OR3 (N554, N539, N321, N392);
xor XOR2 (N555, N553, N170);
not NOT1 (N556, N554);
nand NAND2 (N557, N546, N329);
nand NAND2 (N558, N550, N207);
nand NAND2 (N559, N544, N16);
nor NOR3 (N560, N545, N3, N554);
not NOT1 (N561, N559);
nor NOR2 (N562, N557, N304);
nand NAND2 (N563, N560, N302);
nand NAND4 (N564, N536, N227, N355, N5);
nor NOR4 (N565, N558, N537, N58, N486);
or OR4 (N566, N551, N459, N329, N120);
not NOT1 (N567, N563);
nor NOR4 (N568, N561, N84, N6, N77);
and AND4 (N569, N552, N64, N200, N391);
nor NOR2 (N570, N556, N312);
nand NAND2 (N571, N541, N481);
xor XOR2 (N572, N566, N452);
nand NAND4 (N573, N570, N406, N211, N348);
and AND3 (N574, N573, N263, N397);
not NOT1 (N575, N565);
nor NOR3 (N576, N575, N14, N558);
xor XOR2 (N577, N562, N273);
nand NAND3 (N578, N572, N167, N35);
and AND4 (N579, N578, N172, N192, N385);
not NOT1 (N580, N564);
nor NOR4 (N581, N580, N195, N163, N404);
not NOT1 (N582, N567);
and AND2 (N583, N582, N581);
and AND4 (N584, N328, N163, N230, N46);
xor XOR2 (N585, N584, N564);
and AND2 (N586, N585, N377);
and AND2 (N587, N571, N21);
nor NOR4 (N588, N577, N187, N520, N257);
nand NAND2 (N589, N576, N107);
xor XOR2 (N590, N555, N557);
or OR2 (N591, N588, N521);
xor XOR2 (N592, N589, N36);
or OR2 (N593, N586, N298);
xor XOR2 (N594, N568, N224);
nand NAND3 (N595, N594, N219, N73);
nor NOR4 (N596, N579, N492, N80, N336);
buf BUF1 (N597, N591);
xor XOR2 (N598, N590, N154);
nor NOR2 (N599, N595, N370);
buf BUF1 (N600, N596);
not NOT1 (N601, N598);
and AND3 (N602, N574, N404, N327);
xor XOR2 (N603, N599, N90);
and AND4 (N604, N592, N586, N524, N356);
buf BUF1 (N605, N604);
nor NOR4 (N606, N593, N477, N159, N451);
or OR3 (N607, N597, N340, N245);
or OR2 (N608, N587, N489);
not NOT1 (N609, N601);
or OR4 (N610, N569, N147, N360, N282);
and AND3 (N611, N603, N494, N203);
and AND4 (N612, N610, N243, N124, N582);
or OR4 (N613, N605, N112, N19, N363);
or OR2 (N614, N583, N59);
nor NOR4 (N615, N600, N328, N69, N95);
buf BUF1 (N616, N614);
xor XOR2 (N617, N608, N484);
and AND4 (N618, N613, N36, N154, N159);
not NOT1 (N619, N611);
xor XOR2 (N620, N612, N114);
not NOT1 (N621, N617);
or OR4 (N622, N606, N579, N404, N284);
xor XOR2 (N623, N607, N380);
not NOT1 (N624, N616);
xor XOR2 (N625, N619, N173);
xor XOR2 (N626, N622, N538);
nor NOR2 (N627, N615, N576);
or OR3 (N628, N623, N603, N424);
or OR3 (N629, N620, N125, N21);
buf BUF1 (N630, N624);
xor XOR2 (N631, N627, N557);
or OR4 (N632, N630, N435, N460, N359);
and AND2 (N633, N602, N124);
or OR3 (N634, N631, N299, N413);
nand NAND2 (N635, N629, N328);
buf BUF1 (N636, N626);
xor XOR2 (N637, N636, N489);
nor NOR3 (N638, N625, N155, N154);
xor XOR2 (N639, N633, N172);
nor NOR4 (N640, N638, N135, N299, N546);
nand NAND2 (N641, N634, N457);
not NOT1 (N642, N632);
not NOT1 (N643, N642);
or OR3 (N644, N635, N448, N135);
xor XOR2 (N645, N621, N547);
nor NOR3 (N646, N628, N25, N125);
not NOT1 (N647, N639);
or OR4 (N648, N637, N289, N638, N76);
and AND3 (N649, N618, N74, N526);
or OR4 (N650, N645, N114, N227, N30);
and AND3 (N651, N609, N512, N403);
xor XOR2 (N652, N651, N83);
xor XOR2 (N653, N648, N439);
nand NAND2 (N654, N640, N551);
xor XOR2 (N655, N641, N67);
nand NAND3 (N656, N655, N549, N621);
buf BUF1 (N657, N649);
buf BUF1 (N658, N650);
xor XOR2 (N659, N658, N88);
or OR2 (N660, N646, N67);
or OR3 (N661, N660, N50, N215);
or OR3 (N662, N644, N537, N263);
not NOT1 (N663, N652);
nand NAND4 (N664, N659, N185, N470, N558);
xor XOR2 (N665, N656, N164);
buf BUF1 (N666, N661);
or OR3 (N667, N663, N80, N32);
or OR4 (N668, N666, N56, N62, N533);
and AND4 (N669, N664, N456, N243, N634);
buf BUF1 (N670, N668);
xor XOR2 (N671, N643, N455);
and AND3 (N672, N665, N411, N389);
or OR4 (N673, N670, N541, N586, N172);
not NOT1 (N674, N647);
nand NAND4 (N675, N657, N334, N528, N358);
buf BUF1 (N676, N674);
and AND2 (N677, N662, N570);
buf BUF1 (N678, N654);
xor XOR2 (N679, N653, N561);
xor XOR2 (N680, N677, N14);
or OR2 (N681, N667, N564);
buf BUF1 (N682, N680);
and AND4 (N683, N675, N597, N592, N414);
not NOT1 (N684, N682);
or OR4 (N685, N684, N260, N542, N412);
and AND2 (N686, N681, N137);
or OR3 (N687, N685, N312, N482);
or OR2 (N688, N669, N543);
xor XOR2 (N689, N673, N270);
xor XOR2 (N690, N686, N400);
buf BUF1 (N691, N690);
nand NAND4 (N692, N683, N102, N267, N358);
xor XOR2 (N693, N671, N189);
buf BUF1 (N694, N678);
xor XOR2 (N695, N692, N635);
buf BUF1 (N696, N691);
xor XOR2 (N697, N694, N571);
xor XOR2 (N698, N679, N481);
and AND2 (N699, N697, N470);
xor XOR2 (N700, N688, N499);
not NOT1 (N701, N687);
nand NAND2 (N702, N689, N454);
buf BUF1 (N703, N702);
xor XOR2 (N704, N695, N343);
xor XOR2 (N705, N676, N341);
or OR2 (N706, N672, N328);
xor XOR2 (N707, N699, N166);
xor XOR2 (N708, N700, N478);
and AND2 (N709, N693, N127);
and AND2 (N710, N705, N583);
xor XOR2 (N711, N706, N653);
buf BUF1 (N712, N707);
or OR2 (N713, N712, N360);
and AND3 (N714, N696, N610, N541);
nand NAND4 (N715, N714, N126, N648, N238);
buf BUF1 (N716, N704);
xor XOR2 (N717, N716, N174);
buf BUF1 (N718, N703);
and AND4 (N719, N711, N443, N425, N495);
or OR3 (N720, N717, N605, N577);
or OR3 (N721, N708, N571, N560);
and AND4 (N722, N710, N674, N446, N531);
and AND2 (N723, N722, N672);
not NOT1 (N724, N698);
nand NAND3 (N725, N720, N706, N181);
nor NOR3 (N726, N721, N122, N218);
nand NAND2 (N727, N715, N704);
nand NAND3 (N728, N701, N149, N518);
xor XOR2 (N729, N723, N402);
not NOT1 (N730, N726);
nor NOR3 (N731, N713, N176, N489);
nor NOR4 (N732, N718, N208, N490, N313);
or OR3 (N733, N729, N711, N546);
buf BUF1 (N734, N732);
nand NAND2 (N735, N733, N567);
or OR4 (N736, N719, N579, N313, N694);
or OR2 (N737, N731, N15);
xor XOR2 (N738, N727, N187);
nand NAND2 (N739, N709, N155);
xor XOR2 (N740, N738, N20);
xor XOR2 (N741, N725, N13);
buf BUF1 (N742, N741);
buf BUF1 (N743, N742);
buf BUF1 (N744, N740);
or OR4 (N745, N724, N172, N375, N405);
not NOT1 (N746, N736);
nor NOR2 (N747, N744, N185);
xor XOR2 (N748, N737, N289);
xor XOR2 (N749, N747, N579);
nor NOR4 (N750, N749, N384, N466, N205);
xor XOR2 (N751, N748, N47);
nor NOR3 (N752, N746, N94, N48);
nor NOR4 (N753, N730, N481, N105, N133);
xor XOR2 (N754, N752, N588);
nand NAND4 (N755, N728, N15, N530, N717);
nand NAND2 (N756, N734, N726);
not NOT1 (N757, N743);
or OR3 (N758, N754, N754, N680);
and AND4 (N759, N739, N96, N130, N576);
xor XOR2 (N760, N751, N509);
and AND3 (N761, N753, N186, N713);
xor XOR2 (N762, N758, N256);
xor XOR2 (N763, N755, N246);
and AND2 (N764, N750, N639);
nor NOR3 (N765, N756, N188, N686);
nand NAND4 (N766, N757, N379, N40, N579);
nor NOR4 (N767, N765, N42, N292, N763);
and AND3 (N768, N668, N379, N223);
xor XOR2 (N769, N760, N108);
buf BUF1 (N770, N745);
not NOT1 (N771, N769);
nor NOR2 (N772, N735, N619);
buf BUF1 (N773, N768);
nand NAND4 (N774, N764, N216, N755, N347);
not NOT1 (N775, N770);
buf BUF1 (N776, N773);
buf BUF1 (N777, N759);
and AND3 (N778, N766, N353, N365);
and AND4 (N779, N775, N17, N344, N158);
and AND4 (N780, N778, N83, N256, N373);
nor NOR3 (N781, N780, N236, N381);
nor NOR3 (N782, N774, N293, N129);
or OR4 (N783, N782, N673, N769, N199);
not NOT1 (N784, N776);
not NOT1 (N785, N761);
nor NOR2 (N786, N767, N268);
nor NOR4 (N787, N779, N263, N538, N279);
not NOT1 (N788, N762);
buf BUF1 (N789, N786);
and AND4 (N790, N789, N768, N673, N769);
nor NOR2 (N791, N790, N98);
nor NOR4 (N792, N785, N545, N258, N435);
nand NAND4 (N793, N783, N222, N204, N189);
nor NOR4 (N794, N788, N464, N128, N85);
not NOT1 (N795, N787);
or OR4 (N796, N793, N665, N25, N587);
buf BUF1 (N797, N792);
nor NOR3 (N798, N777, N223, N231);
nor NOR4 (N799, N794, N244, N474, N226);
or OR4 (N800, N797, N732, N437, N258);
buf BUF1 (N801, N791);
buf BUF1 (N802, N801);
or OR2 (N803, N798, N632);
xor XOR2 (N804, N795, N702);
and AND4 (N805, N784, N336, N472, N611);
or OR2 (N806, N771, N421);
xor XOR2 (N807, N803, N632);
nor NOR2 (N808, N772, N194);
buf BUF1 (N809, N802);
not NOT1 (N810, N799);
nor NOR4 (N811, N808, N502, N267, N634);
and AND4 (N812, N809, N199, N61, N565);
or OR2 (N813, N805, N334);
xor XOR2 (N814, N812, N35);
buf BUF1 (N815, N811);
not NOT1 (N816, N804);
xor XOR2 (N817, N814, N351);
xor XOR2 (N818, N781, N449);
not NOT1 (N819, N817);
nand NAND4 (N820, N813, N193, N35, N321);
nor NOR3 (N821, N816, N557, N266);
or OR2 (N822, N820, N670);
xor XOR2 (N823, N800, N631);
and AND3 (N824, N815, N583, N95);
not NOT1 (N825, N824);
and AND2 (N826, N819, N159);
not NOT1 (N827, N807);
not NOT1 (N828, N823);
or OR3 (N829, N822, N429, N246);
and AND2 (N830, N796, N215);
and AND2 (N831, N810, N294);
nand NAND4 (N832, N828, N269, N830, N331);
buf BUF1 (N833, N67);
buf BUF1 (N834, N833);
not NOT1 (N835, N821);
and AND4 (N836, N806, N716, N329, N669);
buf BUF1 (N837, N834);
buf BUF1 (N838, N836);
nand NAND3 (N839, N838, N535, N249);
or OR3 (N840, N825, N448, N443);
and AND2 (N841, N835, N523);
nor NOR3 (N842, N818, N584, N285);
buf BUF1 (N843, N827);
nor NOR2 (N844, N840, N488);
or OR3 (N845, N837, N756, N700);
xor XOR2 (N846, N832, N647);
and AND2 (N847, N839, N86);
not NOT1 (N848, N844);
or OR4 (N849, N826, N693, N142, N463);
or OR3 (N850, N848, N220, N479);
not NOT1 (N851, N831);
or OR4 (N852, N829, N835, N130, N212);
buf BUF1 (N853, N843);
and AND4 (N854, N851, N193, N610, N819);
or OR3 (N855, N845, N641, N498);
not NOT1 (N856, N847);
and AND3 (N857, N849, N71, N608);
and AND2 (N858, N852, N590);
not NOT1 (N859, N857);
or OR4 (N860, N858, N289, N547, N13);
or OR3 (N861, N855, N81, N517);
buf BUF1 (N862, N846);
or OR3 (N863, N856, N438, N833);
nor NOR4 (N864, N842, N200, N190, N760);
xor XOR2 (N865, N861, N186);
and AND4 (N866, N860, N555, N23, N241);
and AND4 (N867, N841, N822, N308, N576);
xor XOR2 (N868, N862, N306);
xor XOR2 (N869, N867, N403);
buf BUF1 (N870, N864);
xor XOR2 (N871, N863, N336);
xor XOR2 (N872, N869, N103);
nor NOR4 (N873, N854, N488, N220, N758);
nor NOR2 (N874, N870, N278);
nor NOR4 (N875, N850, N8, N335, N297);
buf BUF1 (N876, N874);
not NOT1 (N877, N866);
nand NAND4 (N878, N877, N193, N377, N876);
nor NOR4 (N879, N522, N511, N169, N503);
not NOT1 (N880, N871);
xor XOR2 (N881, N875, N241);
and AND2 (N882, N873, N442);
xor XOR2 (N883, N868, N313);
nor NOR2 (N884, N865, N110);
or OR2 (N885, N882, N204);
or OR4 (N886, N859, N503, N789, N87);
and AND3 (N887, N880, N161, N665);
nor NOR4 (N888, N879, N23, N482, N67);
and AND4 (N889, N883, N784, N446, N89);
nand NAND3 (N890, N887, N754, N478);
and AND3 (N891, N886, N518, N359);
xor XOR2 (N892, N891, N286);
xor XOR2 (N893, N884, N501);
xor XOR2 (N894, N892, N542);
and AND3 (N895, N878, N762, N288);
not NOT1 (N896, N853);
nand NAND4 (N897, N885, N134, N380, N7);
buf BUF1 (N898, N893);
nand NAND2 (N899, N872, N274);
and AND3 (N900, N898, N511, N757);
nor NOR4 (N901, N895, N563, N235, N593);
and AND3 (N902, N900, N621, N9);
nor NOR2 (N903, N902, N418);
and AND2 (N904, N888, N83);
xor XOR2 (N905, N894, N280);
not NOT1 (N906, N881);
nand NAND2 (N907, N903, N161);
nand NAND3 (N908, N897, N824, N83);
nand NAND2 (N909, N896, N856);
and AND3 (N910, N904, N383, N504);
buf BUF1 (N911, N899);
buf BUF1 (N912, N905);
nand NAND2 (N913, N890, N78);
buf BUF1 (N914, N906);
not NOT1 (N915, N910);
not NOT1 (N916, N901);
or OR2 (N917, N914, N569);
not NOT1 (N918, N889);
not NOT1 (N919, N916);
buf BUF1 (N920, N919);
xor XOR2 (N921, N917, N138);
nor NOR3 (N922, N913, N438, N99);
not NOT1 (N923, N915);
not NOT1 (N924, N911);
nor NOR3 (N925, N922, N154, N125);
not NOT1 (N926, N908);
not NOT1 (N927, N920);
nand NAND2 (N928, N918, N847);
and AND4 (N929, N926, N270, N753, N571);
or OR2 (N930, N923, N492);
not NOT1 (N931, N925);
nand NAND3 (N932, N931, N252, N142);
xor XOR2 (N933, N930, N591);
or OR4 (N934, N929, N927, N707, N624);
and AND3 (N935, N880, N639, N437);
or OR4 (N936, N928, N280, N364, N234);
nand NAND3 (N937, N934, N715, N923);
or OR3 (N938, N907, N288, N560);
nor NOR3 (N939, N938, N282, N772);
buf BUF1 (N940, N936);
not NOT1 (N941, N912);
buf BUF1 (N942, N924);
or OR2 (N943, N921, N772);
or OR2 (N944, N933, N104);
nand NAND4 (N945, N932, N188, N536, N934);
or OR4 (N946, N940, N324, N543, N714);
or OR2 (N947, N946, N866);
nand NAND2 (N948, N937, N293);
nand NAND3 (N949, N948, N867, N413);
or OR3 (N950, N945, N312, N413);
not NOT1 (N951, N942);
nand NAND2 (N952, N943, N104);
or OR3 (N953, N909, N654, N772);
and AND4 (N954, N952, N526, N295, N110);
nand NAND3 (N955, N949, N686, N598);
nand NAND3 (N956, N939, N434, N439);
buf BUF1 (N957, N951);
xor XOR2 (N958, N955, N490);
or OR4 (N959, N941, N684, N182, N649);
not NOT1 (N960, N957);
buf BUF1 (N961, N956);
or OR2 (N962, N958, N605);
nor NOR4 (N963, N959, N338, N397, N58);
and AND3 (N964, N947, N455, N298);
not NOT1 (N965, N954);
and AND3 (N966, N963, N270, N521);
nand NAND2 (N967, N950, N516);
and AND2 (N968, N965, N874);
and AND4 (N969, N967, N615, N840, N685);
not NOT1 (N970, N962);
nand NAND4 (N971, N966, N920, N711, N755);
not NOT1 (N972, N971);
nor NOR3 (N973, N935, N923, N551);
not NOT1 (N974, N964);
xor XOR2 (N975, N973, N692);
or OR4 (N976, N969, N566, N596, N309);
and AND4 (N977, N968, N587, N721, N442);
and AND4 (N978, N976, N52, N184, N846);
or OR4 (N979, N978, N968, N428, N305);
or OR2 (N980, N979, N824);
nor NOR2 (N981, N961, N495);
nor NOR2 (N982, N980, N517);
nor NOR3 (N983, N953, N255, N274);
nand NAND2 (N984, N977, N429);
and AND4 (N985, N944, N214, N707, N877);
not NOT1 (N986, N975);
nor NOR3 (N987, N972, N260, N105);
or OR4 (N988, N982, N700, N155, N947);
and AND4 (N989, N988, N977, N186, N419);
or OR4 (N990, N983, N373, N94, N570);
not NOT1 (N991, N970);
nor NOR4 (N992, N990, N775, N872, N306);
nand NAND2 (N993, N986, N973);
or OR4 (N994, N989, N868, N566, N477);
xor XOR2 (N995, N992, N18);
nand NAND4 (N996, N995, N950, N63, N692);
nand NAND3 (N997, N981, N554, N568);
or OR3 (N998, N993, N705, N644);
not NOT1 (N999, N987);
nor NOR4 (N1000, N994, N962, N221, N764);
buf BUF1 (N1001, N1000);
buf BUF1 (N1002, N974);
xor XOR2 (N1003, N985, N293);
nand NAND3 (N1004, N1001, N612, N254);
buf BUF1 (N1005, N1002);
nand NAND3 (N1006, N1003, N523, N276);
or OR2 (N1007, N1004, N378);
and AND3 (N1008, N1007, N568, N486);
not NOT1 (N1009, N999);
nor NOR4 (N1010, N984, N330, N600, N606);
nor NOR3 (N1011, N1006, N998, N100);
and AND4 (N1012, N864, N689, N791, N722);
buf BUF1 (N1013, N1008);
and AND4 (N1014, N997, N52, N478, N634);
nor NOR4 (N1015, N991, N278, N320, N637);
buf BUF1 (N1016, N1011);
xor XOR2 (N1017, N1010, N85);
and AND3 (N1018, N1012, N429, N54);
nor NOR4 (N1019, N960, N792, N804, N463);
not NOT1 (N1020, N1018);
or OR2 (N1021, N996, N803);
nor NOR4 (N1022, N1017, N805, N295, N275);
nor NOR4 (N1023, N1014, N805, N685, N802);
or OR3 (N1024, N1022, N523, N266);
not NOT1 (N1025, N1016);
and AND3 (N1026, N1019, N393, N611);
not NOT1 (N1027, N1024);
buf BUF1 (N1028, N1021);
buf BUF1 (N1029, N1020);
and AND3 (N1030, N1027, N778, N188);
buf BUF1 (N1031, N1023);
buf BUF1 (N1032, N1013);
and AND3 (N1033, N1030, N383, N670);
buf BUF1 (N1034, N1025);
nor NOR4 (N1035, N1028, N674, N209, N665);
and AND3 (N1036, N1033, N793, N258);
or OR2 (N1037, N1032, N328);
buf BUF1 (N1038, N1031);
buf BUF1 (N1039, N1036);
nor NOR2 (N1040, N1005, N16);
not NOT1 (N1041, N1035);
or OR2 (N1042, N1041, N466);
nand NAND4 (N1043, N1034, N920, N910, N704);
xor XOR2 (N1044, N1037, N479);
and AND4 (N1045, N1026, N980, N828, N53);
or OR3 (N1046, N1029, N878, N319);
not NOT1 (N1047, N1040);
nand NAND2 (N1048, N1042, N18);
or OR3 (N1049, N1039, N474, N462);
nor NOR2 (N1050, N1046, N828);
buf BUF1 (N1051, N1050);
or OR2 (N1052, N1047, N802);
buf BUF1 (N1053, N1048);
nor NOR3 (N1054, N1038, N758, N649);
nor NOR3 (N1055, N1053, N815, N593);
or OR3 (N1056, N1045, N781, N457);
or OR4 (N1057, N1009, N343, N610, N610);
not NOT1 (N1058, N1043);
buf BUF1 (N1059, N1015);
nor NOR3 (N1060, N1054, N537, N280);
buf BUF1 (N1061, N1056);
or OR3 (N1062, N1051, N796, N693);
nand NAND3 (N1063, N1058, N1019, N449);
or OR4 (N1064, N1063, N169, N478, N457);
or OR4 (N1065, N1044, N748, N445, N669);
nor NOR4 (N1066, N1062, N291, N54, N14);
buf BUF1 (N1067, N1060);
nand NAND2 (N1068, N1066, N599);
and AND4 (N1069, N1052, N288, N123, N972);
and AND4 (N1070, N1061, N13, N147, N594);
not NOT1 (N1071, N1065);
or OR4 (N1072, N1069, N882, N440, N648);
buf BUF1 (N1073, N1064);
not NOT1 (N1074, N1073);
nand NAND2 (N1075, N1049, N877);
xor XOR2 (N1076, N1071, N437);
nor NOR3 (N1077, N1059, N699, N922);
xor XOR2 (N1078, N1074, N834);
or OR3 (N1079, N1070, N783, N1029);
or OR3 (N1080, N1076, N449, N135);
xor XOR2 (N1081, N1055, N1042);
nand NAND3 (N1082, N1075, N81, N859);
and AND3 (N1083, N1068, N94, N975);
not NOT1 (N1084, N1067);
nor NOR4 (N1085, N1078, N595, N803, N317);
nor NOR2 (N1086, N1079, N186);
and AND3 (N1087, N1085, N901, N714);
and AND2 (N1088, N1084, N324);
not NOT1 (N1089, N1086);
nor NOR2 (N1090, N1088, N801);
not NOT1 (N1091, N1077);
nor NOR3 (N1092, N1080, N1041, N574);
not NOT1 (N1093, N1087);
nand NAND2 (N1094, N1082, N118);
and AND4 (N1095, N1092, N219, N19, N190);
and AND4 (N1096, N1083, N167, N330, N240);
and AND4 (N1097, N1095, N877, N966, N448);
buf BUF1 (N1098, N1090);
buf BUF1 (N1099, N1089);
and AND3 (N1100, N1094, N350, N989);
nor NOR3 (N1101, N1100, N849, N1012);
buf BUF1 (N1102, N1097);
or OR4 (N1103, N1081, N1087, N1041, N6);
not NOT1 (N1104, N1057);
buf BUF1 (N1105, N1102);
or OR4 (N1106, N1103, N207, N5, N1030);
nor NOR3 (N1107, N1091, N769, N555);
buf BUF1 (N1108, N1105);
xor XOR2 (N1109, N1107, N228);
buf BUF1 (N1110, N1101);
not NOT1 (N1111, N1072);
and AND4 (N1112, N1099, N945, N256, N1047);
or OR2 (N1113, N1106, N972);
nor NOR2 (N1114, N1108, N361);
nand NAND4 (N1115, N1096, N870, N251, N964);
nand NAND4 (N1116, N1104, N456, N858, N478);
or OR2 (N1117, N1110, N225);
nor NOR3 (N1118, N1117, N1080, N172);
or OR4 (N1119, N1114, N148, N178, N772);
not NOT1 (N1120, N1115);
nand NAND4 (N1121, N1112, N967, N704, N423);
not NOT1 (N1122, N1111);
and AND3 (N1123, N1120, N450, N201);
not NOT1 (N1124, N1119);
nand NAND3 (N1125, N1121, N889, N568);
nor NOR2 (N1126, N1118, N1067);
xor XOR2 (N1127, N1123, N532);
nor NOR3 (N1128, N1093, N505, N500);
buf BUF1 (N1129, N1109);
xor XOR2 (N1130, N1127, N154);
xor XOR2 (N1131, N1098, N993);
nor NOR2 (N1132, N1129, N587);
xor XOR2 (N1133, N1130, N217);
nor NOR4 (N1134, N1133, N772, N492, N31);
not NOT1 (N1135, N1124);
nand NAND2 (N1136, N1134, N717);
nor NOR3 (N1137, N1113, N698, N620);
buf BUF1 (N1138, N1132);
not NOT1 (N1139, N1131);
buf BUF1 (N1140, N1139);
nor NOR3 (N1141, N1137, N191, N599);
and AND3 (N1142, N1128, N283, N712);
not NOT1 (N1143, N1135);
buf BUF1 (N1144, N1138);
buf BUF1 (N1145, N1126);
buf BUF1 (N1146, N1141);
xor XOR2 (N1147, N1125, N460);
or OR3 (N1148, N1143, N720, N710);
or OR3 (N1149, N1136, N799, N219);
buf BUF1 (N1150, N1122);
not NOT1 (N1151, N1148);
buf BUF1 (N1152, N1150);
buf BUF1 (N1153, N1145);
and AND3 (N1154, N1152, N1017, N379);
and AND3 (N1155, N1146, N502, N666);
nand NAND3 (N1156, N1142, N118, N251);
or OR2 (N1157, N1140, N921);
not NOT1 (N1158, N1153);
and AND2 (N1159, N1149, N1146);
buf BUF1 (N1160, N1158);
nor NOR3 (N1161, N1147, N389, N1037);
not NOT1 (N1162, N1156);
nor NOR3 (N1163, N1161, N1059, N182);
not NOT1 (N1164, N1163);
nand NAND2 (N1165, N1164, N907);
and AND4 (N1166, N1144, N846, N1126, N415);
xor XOR2 (N1167, N1165, N232);
buf BUF1 (N1168, N1155);
not NOT1 (N1169, N1166);
and AND4 (N1170, N1162, N399, N460, N892);
nor NOR4 (N1171, N1160, N1141, N781, N350);
or OR3 (N1172, N1159, N1087, N1120);
nor NOR2 (N1173, N1171, N153);
nand NAND2 (N1174, N1172, N1108);
and AND3 (N1175, N1169, N1051, N88);
or OR4 (N1176, N1116, N728, N58, N506);
xor XOR2 (N1177, N1154, N748);
and AND3 (N1178, N1173, N253, N680);
xor XOR2 (N1179, N1175, N1141);
nor NOR2 (N1180, N1176, N657);
or OR4 (N1181, N1167, N525, N135, N923);
or OR3 (N1182, N1168, N261, N46);
or OR3 (N1183, N1177, N127, N602);
not NOT1 (N1184, N1181);
xor XOR2 (N1185, N1184, N366);
or OR3 (N1186, N1185, N582, N221);
and AND4 (N1187, N1183, N24, N77, N657);
and AND2 (N1188, N1174, N392);
nor NOR4 (N1189, N1188, N739, N517, N296);
not NOT1 (N1190, N1157);
or OR4 (N1191, N1179, N368, N288, N991);
and AND3 (N1192, N1180, N1058, N1191);
nand NAND3 (N1193, N839, N894, N186);
nor NOR3 (N1194, N1186, N734, N1002);
buf BUF1 (N1195, N1190);
xor XOR2 (N1196, N1182, N906);
not NOT1 (N1197, N1196);
and AND2 (N1198, N1178, N708);
buf BUF1 (N1199, N1187);
nor NOR4 (N1200, N1189, N770, N1165, N1165);
nand NAND3 (N1201, N1198, N867, N380);
nand NAND2 (N1202, N1170, N585);
buf BUF1 (N1203, N1194);
xor XOR2 (N1204, N1192, N815);
buf BUF1 (N1205, N1201);
xor XOR2 (N1206, N1193, N753);
nand NAND2 (N1207, N1202, N209);
buf BUF1 (N1208, N1151);
and AND2 (N1209, N1203, N158);
and AND3 (N1210, N1207, N879, N119);
and AND3 (N1211, N1208, N275, N906);
and AND4 (N1212, N1210, N868, N19, N71);
xor XOR2 (N1213, N1197, N1169);
nor NOR4 (N1214, N1200, N1171, N759, N810);
xor XOR2 (N1215, N1211, N158);
or OR2 (N1216, N1209, N157);
nor NOR2 (N1217, N1214, N1194);
or OR3 (N1218, N1205, N542, N1056);
or OR4 (N1219, N1195, N1101, N281, N831);
nand NAND2 (N1220, N1218, N829);
not NOT1 (N1221, N1216);
or OR2 (N1222, N1215, N1144);
or OR3 (N1223, N1221, N534, N571);
not NOT1 (N1224, N1223);
not NOT1 (N1225, N1204);
xor XOR2 (N1226, N1217, N859);
buf BUF1 (N1227, N1222);
or OR2 (N1228, N1199, N768);
xor XOR2 (N1229, N1227, N605);
or OR4 (N1230, N1226, N910, N780, N584);
buf BUF1 (N1231, N1224);
nand NAND4 (N1232, N1212, N593, N1035, N867);
xor XOR2 (N1233, N1229, N915);
not NOT1 (N1234, N1213);
not NOT1 (N1235, N1231);
buf BUF1 (N1236, N1219);
nor NOR2 (N1237, N1220, N256);
or OR3 (N1238, N1237, N882, N613);
nand NAND4 (N1239, N1233, N947, N358, N1230);
nand NAND4 (N1240, N684, N624, N622, N386);
xor XOR2 (N1241, N1228, N267);
nand NAND4 (N1242, N1206, N1166, N255, N425);
or OR4 (N1243, N1235, N217, N186, N723);
not NOT1 (N1244, N1236);
not NOT1 (N1245, N1238);
buf BUF1 (N1246, N1232);
not NOT1 (N1247, N1241);
buf BUF1 (N1248, N1240);
and AND2 (N1249, N1243, N1232);
nand NAND2 (N1250, N1248, N589);
nor NOR2 (N1251, N1246, N193);
nand NAND3 (N1252, N1242, N187, N937);
nor NOR4 (N1253, N1239, N739, N504, N1132);
and AND2 (N1254, N1251, N407);
xor XOR2 (N1255, N1250, N773);
and AND3 (N1256, N1234, N321, N426);
or OR2 (N1257, N1247, N1111);
not NOT1 (N1258, N1257);
nand NAND3 (N1259, N1258, N869, N822);
nor NOR3 (N1260, N1255, N726, N1109);
nor NOR2 (N1261, N1256, N623);
nand NAND4 (N1262, N1252, N1172, N970, N518);
nand NAND4 (N1263, N1259, N227, N878, N481);
not NOT1 (N1264, N1261);
buf BUF1 (N1265, N1264);
not NOT1 (N1266, N1225);
not NOT1 (N1267, N1244);
not NOT1 (N1268, N1245);
or OR2 (N1269, N1267, N1216);
or OR2 (N1270, N1266, N876);
or OR3 (N1271, N1269, N734, N747);
or OR4 (N1272, N1254, N372, N57, N764);
and AND3 (N1273, N1268, N243, N906);
buf BUF1 (N1274, N1253);
and AND2 (N1275, N1263, N356);
and AND2 (N1276, N1265, N504);
buf BUF1 (N1277, N1260);
nand NAND4 (N1278, N1271, N860, N358, N604);
buf BUF1 (N1279, N1277);
xor XOR2 (N1280, N1278, N1106);
or OR4 (N1281, N1274, N404, N340, N1112);
nand NAND2 (N1282, N1280, N1232);
nand NAND4 (N1283, N1281, N636, N1164, N536);
and AND2 (N1284, N1282, N250);
or OR3 (N1285, N1275, N1224, N565);
xor XOR2 (N1286, N1272, N111);
xor XOR2 (N1287, N1283, N756);
and AND2 (N1288, N1273, N1199);
not NOT1 (N1289, N1249);
or OR3 (N1290, N1262, N1232, N181);
or OR3 (N1291, N1285, N438, N631);
and AND2 (N1292, N1291, N870);
or OR3 (N1293, N1279, N499, N744);
and AND3 (N1294, N1276, N868, N353);
and AND3 (N1295, N1288, N571, N197);
nand NAND4 (N1296, N1293, N945, N107, N402);
and AND4 (N1297, N1286, N214, N908, N987);
buf BUF1 (N1298, N1290);
xor XOR2 (N1299, N1296, N1209);
nor NOR2 (N1300, N1287, N1194);
and AND3 (N1301, N1299, N481, N686);
or OR2 (N1302, N1284, N386);
xor XOR2 (N1303, N1300, N67);
and AND4 (N1304, N1303, N1205, N1113, N1050);
or OR3 (N1305, N1270, N995, N1150);
nand NAND4 (N1306, N1304, N1241, N572, N303);
nor NOR3 (N1307, N1301, N1129, N463);
and AND2 (N1308, N1295, N1157);
not NOT1 (N1309, N1297);
and AND3 (N1310, N1289, N1066, N1055);
buf BUF1 (N1311, N1309);
nor NOR2 (N1312, N1305, N601);
xor XOR2 (N1313, N1302, N1301);
nand NAND3 (N1314, N1307, N145, N117);
nor NOR2 (N1315, N1292, N486);
or OR4 (N1316, N1294, N672, N883, N935);
xor XOR2 (N1317, N1310, N652);
nand NAND3 (N1318, N1315, N485, N357);
nand NAND4 (N1319, N1298, N1140, N665, N30);
xor XOR2 (N1320, N1314, N1247);
or OR2 (N1321, N1318, N868);
or OR4 (N1322, N1311, N167, N661, N735);
and AND2 (N1323, N1321, N1219);
or OR4 (N1324, N1323, N482, N400, N1296);
or OR2 (N1325, N1319, N1277);
and AND2 (N1326, N1322, N1299);
and AND2 (N1327, N1326, N911);
nand NAND3 (N1328, N1313, N888, N846);
or OR4 (N1329, N1306, N664, N888, N1159);
nor NOR2 (N1330, N1324, N282);
and AND3 (N1331, N1308, N254, N177);
nor NOR3 (N1332, N1325, N580, N676);
nand NAND2 (N1333, N1330, N308);
and AND4 (N1334, N1328, N183, N396, N1072);
not NOT1 (N1335, N1316);
nand NAND3 (N1336, N1334, N994, N777);
or OR2 (N1337, N1327, N638);
and AND2 (N1338, N1337, N329);
nor NOR3 (N1339, N1332, N1269, N1114);
xor XOR2 (N1340, N1329, N727);
and AND2 (N1341, N1336, N264);
buf BUF1 (N1342, N1320);
and AND4 (N1343, N1341, N826, N935, N391);
buf BUF1 (N1344, N1317);
and AND3 (N1345, N1340, N1229, N802);
or OR4 (N1346, N1339, N13, N16, N1138);
buf BUF1 (N1347, N1345);
or OR2 (N1348, N1342, N1315);
and AND4 (N1349, N1312, N52, N899, N1164);
nand NAND3 (N1350, N1331, N535, N422);
and AND3 (N1351, N1344, N1270, N317);
or OR4 (N1352, N1346, N370, N1162, N1108);
xor XOR2 (N1353, N1348, N153);
nand NAND2 (N1354, N1333, N155);
not NOT1 (N1355, N1353);
nor NOR2 (N1356, N1351, N273);
or OR4 (N1357, N1347, N420, N670, N584);
not NOT1 (N1358, N1357);
nand NAND2 (N1359, N1349, N602);
and AND4 (N1360, N1343, N459, N303, N1111);
and AND4 (N1361, N1359, N5, N534, N614);
nor NOR2 (N1362, N1361, N583);
or OR2 (N1363, N1352, N729);
xor XOR2 (N1364, N1356, N738);
buf BUF1 (N1365, N1362);
nand NAND3 (N1366, N1358, N1291, N839);
and AND3 (N1367, N1354, N1243, N285);
and AND4 (N1368, N1367, N73, N1147, N856);
and AND4 (N1369, N1360, N361, N1340, N805);
not NOT1 (N1370, N1368);
or OR2 (N1371, N1365, N1352);
nand NAND4 (N1372, N1350, N208, N65, N790);
nand NAND2 (N1373, N1369, N458);
nor NOR2 (N1374, N1371, N1051);
or OR4 (N1375, N1363, N458, N588, N259);
xor XOR2 (N1376, N1374, N1260);
xor XOR2 (N1377, N1338, N35);
nor NOR2 (N1378, N1364, N1032);
xor XOR2 (N1379, N1335, N817);
or OR3 (N1380, N1375, N271, N65);
xor XOR2 (N1381, N1380, N753);
not NOT1 (N1382, N1370);
xor XOR2 (N1383, N1377, N108);
and AND4 (N1384, N1382, N1171, N989, N585);
nor NOR4 (N1385, N1366, N406, N893, N638);
nor NOR3 (N1386, N1384, N1057, N283);
nor NOR4 (N1387, N1383, N123, N141, N1065);
nor NOR4 (N1388, N1385, N1118, N637, N432);
or OR3 (N1389, N1373, N998, N556);
buf BUF1 (N1390, N1378);
xor XOR2 (N1391, N1388, N361);
and AND3 (N1392, N1387, N887, N897);
nand NAND4 (N1393, N1392, N652, N580, N209);
buf BUF1 (N1394, N1390);
not NOT1 (N1395, N1393);
nand NAND3 (N1396, N1394, N239, N1328);
xor XOR2 (N1397, N1389, N452);
nor NOR3 (N1398, N1355, N1226, N1366);
nand NAND3 (N1399, N1398, N1283, N1325);
xor XOR2 (N1400, N1372, N718);
buf BUF1 (N1401, N1400);
xor XOR2 (N1402, N1395, N1268);
nand NAND3 (N1403, N1396, N226, N1316);
xor XOR2 (N1404, N1403, N103);
buf BUF1 (N1405, N1401);
not NOT1 (N1406, N1397);
not NOT1 (N1407, N1376);
xor XOR2 (N1408, N1399, N1055);
nor NOR3 (N1409, N1404, N1023, N25);
not NOT1 (N1410, N1408);
buf BUF1 (N1411, N1406);
buf BUF1 (N1412, N1407);
nor NOR3 (N1413, N1405, N901, N1219);
nand NAND3 (N1414, N1411, N1389, N19);
or OR4 (N1415, N1413, N970, N206, N971);
nand NAND3 (N1416, N1381, N427, N29);
buf BUF1 (N1417, N1402);
nand NAND4 (N1418, N1410, N1020, N522, N146);
nand NAND4 (N1419, N1417, N697, N4, N255);
nor NOR4 (N1420, N1415, N1231, N532, N1402);
nor NOR4 (N1421, N1416, N1344, N1387, N545);
nand NAND2 (N1422, N1386, N960);
not NOT1 (N1423, N1412);
nor NOR3 (N1424, N1423, N1006, N705);
not NOT1 (N1425, N1391);
xor XOR2 (N1426, N1424, N1232);
or OR4 (N1427, N1414, N544, N1391, N652);
nor NOR2 (N1428, N1427, N342);
nor NOR4 (N1429, N1425, N1403, N754, N699);
buf BUF1 (N1430, N1426);
xor XOR2 (N1431, N1421, N747);
xor XOR2 (N1432, N1429, N742);
or OR3 (N1433, N1430, N626, N1327);
or OR3 (N1434, N1431, N970, N97);
and AND2 (N1435, N1409, N451);
or OR4 (N1436, N1433, N569, N203, N814);
or OR2 (N1437, N1419, N393);
and AND3 (N1438, N1422, N171, N572);
not NOT1 (N1439, N1420);
xor XOR2 (N1440, N1436, N622);
buf BUF1 (N1441, N1428);
not NOT1 (N1442, N1438);
not NOT1 (N1443, N1434);
not NOT1 (N1444, N1418);
and AND4 (N1445, N1432, N647, N1374, N132);
not NOT1 (N1446, N1440);
nand NAND4 (N1447, N1442, N570, N219, N638);
xor XOR2 (N1448, N1445, N955);
nand NAND2 (N1449, N1446, N540);
nand NAND2 (N1450, N1448, N325);
nand NAND3 (N1451, N1450, N686, N910);
not NOT1 (N1452, N1379);
and AND3 (N1453, N1447, N469, N991);
nor NOR4 (N1454, N1449, N191, N770, N799);
buf BUF1 (N1455, N1439);
not NOT1 (N1456, N1451);
xor XOR2 (N1457, N1443, N342);
nor NOR4 (N1458, N1453, N968, N828, N591);
nor NOR2 (N1459, N1454, N624);
not NOT1 (N1460, N1452);
nand NAND3 (N1461, N1444, N1311, N747);
nand NAND2 (N1462, N1460, N273);
nor NOR2 (N1463, N1462, N163);
not NOT1 (N1464, N1435);
or OR2 (N1465, N1455, N238);
and AND3 (N1466, N1456, N461, N931);
nand NAND3 (N1467, N1465, N951, N1123);
nor NOR2 (N1468, N1467, N287);
nor NOR4 (N1469, N1464, N601, N597, N560);
and AND2 (N1470, N1437, N1388);
and AND4 (N1471, N1469, N1420, N437, N1343);
not NOT1 (N1472, N1461);
or OR3 (N1473, N1471, N245, N944);
or OR4 (N1474, N1468, N495, N208, N1263);
and AND4 (N1475, N1459, N846, N952, N804);
buf BUF1 (N1476, N1458);
buf BUF1 (N1477, N1466);
not NOT1 (N1478, N1474);
and AND3 (N1479, N1475, N916, N479);
or OR3 (N1480, N1457, N753, N113);
buf BUF1 (N1481, N1463);
or OR4 (N1482, N1470, N1244, N353, N512);
nand NAND3 (N1483, N1473, N773, N1171);
not NOT1 (N1484, N1476);
and AND4 (N1485, N1479, N554, N220, N443);
nor NOR3 (N1486, N1483, N1436, N923);
not NOT1 (N1487, N1481);
or OR4 (N1488, N1472, N820, N751, N1033);
not NOT1 (N1489, N1484);
not NOT1 (N1490, N1487);
xor XOR2 (N1491, N1490, N465);
nand NAND3 (N1492, N1485, N1113, N1059);
and AND3 (N1493, N1488, N550, N793);
and AND3 (N1494, N1491, N1346, N996);
nor NOR2 (N1495, N1489, N134);
not NOT1 (N1496, N1480);
not NOT1 (N1497, N1478);
or OR3 (N1498, N1477, N106, N1269);
or OR4 (N1499, N1441, N1489, N384, N1286);
and AND4 (N1500, N1497, N137, N84, N1173);
not NOT1 (N1501, N1499);
or OR2 (N1502, N1486, N570);
nor NOR3 (N1503, N1498, N87, N558);
xor XOR2 (N1504, N1495, N1400);
nor NOR3 (N1505, N1504, N903, N635);
or OR4 (N1506, N1505, N7, N311, N415);
not NOT1 (N1507, N1493);
nor NOR4 (N1508, N1492, N1177, N881, N323);
nand NAND3 (N1509, N1507, N1469, N162);
buf BUF1 (N1510, N1501);
not NOT1 (N1511, N1496);
nor NOR2 (N1512, N1511, N815);
nor NOR4 (N1513, N1494, N922, N1489, N627);
buf BUF1 (N1514, N1513);
or OR3 (N1515, N1482, N1440, N279);
nor NOR4 (N1516, N1506, N267, N24, N255);
xor XOR2 (N1517, N1508, N1025);
not NOT1 (N1518, N1515);
or OR4 (N1519, N1512, N1370, N329, N935);
nor NOR2 (N1520, N1500, N610);
and AND3 (N1521, N1510, N379, N794);
nand NAND2 (N1522, N1520, N1238);
not NOT1 (N1523, N1518);
nor NOR2 (N1524, N1521, N202);
nor NOR3 (N1525, N1523, N816, N1157);
nand NAND4 (N1526, N1502, N531, N873, N584);
nor NOR3 (N1527, N1516, N254, N1190);
nand NAND2 (N1528, N1514, N134);
not NOT1 (N1529, N1517);
xor XOR2 (N1530, N1529, N39);
xor XOR2 (N1531, N1503, N1023);
xor XOR2 (N1532, N1509, N1489);
nand NAND2 (N1533, N1527, N353);
nand NAND3 (N1534, N1531, N1372, N839);
nor NOR2 (N1535, N1534, N578);
or OR2 (N1536, N1530, N22);
not NOT1 (N1537, N1532);
buf BUF1 (N1538, N1537);
nand NAND3 (N1539, N1524, N241, N970);
nand NAND3 (N1540, N1539, N1504, N13);
and AND3 (N1541, N1536, N1534, N553);
not NOT1 (N1542, N1525);
xor XOR2 (N1543, N1519, N886);
buf BUF1 (N1544, N1542);
buf BUF1 (N1545, N1522);
buf BUF1 (N1546, N1528);
not NOT1 (N1547, N1538);
not NOT1 (N1548, N1547);
buf BUF1 (N1549, N1526);
xor XOR2 (N1550, N1540, N418);
buf BUF1 (N1551, N1544);
buf BUF1 (N1552, N1541);
buf BUF1 (N1553, N1552);
buf BUF1 (N1554, N1546);
or OR3 (N1555, N1548, N320, N1513);
not NOT1 (N1556, N1555);
nand NAND4 (N1557, N1543, N1258, N1507, N147);
not NOT1 (N1558, N1556);
or OR4 (N1559, N1545, N632, N727, N329);
buf BUF1 (N1560, N1559);
nor NOR4 (N1561, N1533, N276, N918, N411);
buf BUF1 (N1562, N1561);
nand NAND2 (N1563, N1551, N1530);
nor NOR4 (N1564, N1562, N1415, N1149, N1255);
buf BUF1 (N1565, N1558);
xor XOR2 (N1566, N1565, N1499);
or OR4 (N1567, N1554, N439, N452, N582);
nor NOR2 (N1568, N1535, N1283);
buf BUF1 (N1569, N1549);
nor NOR4 (N1570, N1564, N1031, N183, N1120);
or OR3 (N1571, N1566, N1448, N655);
not NOT1 (N1572, N1560);
buf BUF1 (N1573, N1572);
nor NOR3 (N1574, N1570, N1094, N1422);
buf BUF1 (N1575, N1557);
buf BUF1 (N1576, N1553);
nor NOR2 (N1577, N1575, N30);
and AND3 (N1578, N1569, N744, N1305);
and AND3 (N1579, N1550, N215, N614);
xor XOR2 (N1580, N1571, N187);
nand NAND3 (N1581, N1576, N186, N1012);
or OR3 (N1582, N1578, N1551, N805);
or OR4 (N1583, N1580, N366, N183, N288);
xor XOR2 (N1584, N1574, N1453);
not NOT1 (N1585, N1583);
and AND2 (N1586, N1567, N1512);
buf BUF1 (N1587, N1573);
not NOT1 (N1588, N1587);
and AND3 (N1589, N1585, N1044, N624);
or OR4 (N1590, N1584, N51, N640, N1264);
nor NOR2 (N1591, N1590, N1379);
nand NAND2 (N1592, N1586, N993);
not NOT1 (N1593, N1579);
not NOT1 (N1594, N1563);
nor NOR4 (N1595, N1593, N804, N316, N773);
not NOT1 (N1596, N1581);
nand NAND4 (N1597, N1594, N1148, N119, N435);
xor XOR2 (N1598, N1588, N472);
and AND4 (N1599, N1596, N288, N624, N1032);
xor XOR2 (N1600, N1599, N1318);
not NOT1 (N1601, N1577);
and AND2 (N1602, N1592, N866);
or OR4 (N1603, N1602, N389, N167, N83);
xor XOR2 (N1604, N1568, N1516);
or OR2 (N1605, N1604, N127);
xor XOR2 (N1606, N1589, N1403);
and AND2 (N1607, N1595, N1404);
or OR4 (N1608, N1598, N650, N1128, N189);
buf BUF1 (N1609, N1606);
nor NOR3 (N1610, N1609, N941, N256);
buf BUF1 (N1611, N1582);
not NOT1 (N1612, N1608);
xor XOR2 (N1613, N1601, N21);
buf BUF1 (N1614, N1605);
buf BUF1 (N1615, N1610);
xor XOR2 (N1616, N1612, N1186);
not NOT1 (N1617, N1611);
or OR4 (N1618, N1597, N41, N235, N1023);
or OR2 (N1619, N1614, N1258);
nand NAND3 (N1620, N1615, N222, N1007);
buf BUF1 (N1621, N1613);
xor XOR2 (N1622, N1620, N1443);
nor NOR4 (N1623, N1603, N635, N1503, N90);
not NOT1 (N1624, N1617);
xor XOR2 (N1625, N1618, N630);
and AND2 (N1626, N1591, N226);
nand NAND4 (N1627, N1600, N147, N974, N255);
not NOT1 (N1628, N1619);
nand NAND4 (N1629, N1621, N1437, N852, N1233);
nand NAND3 (N1630, N1627, N1236, N1375);
and AND3 (N1631, N1624, N225, N1599);
and AND2 (N1632, N1616, N846);
nand NAND4 (N1633, N1623, N637, N640, N547);
buf BUF1 (N1634, N1625);
buf BUF1 (N1635, N1628);
xor XOR2 (N1636, N1631, N1354);
not NOT1 (N1637, N1633);
nand NAND4 (N1638, N1632, N680, N731, N1626);
nand NAND2 (N1639, N365, N1364);
xor XOR2 (N1640, N1629, N575);
buf BUF1 (N1641, N1636);
not NOT1 (N1642, N1638);
nor NOR3 (N1643, N1635, N711, N536);
nand NAND3 (N1644, N1630, N1089, N781);
or OR3 (N1645, N1642, N1429, N1239);
xor XOR2 (N1646, N1645, N1205);
nor NOR3 (N1647, N1643, N820, N792);
xor XOR2 (N1648, N1640, N1493);
not NOT1 (N1649, N1639);
and AND2 (N1650, N1646, N90);
xor XOR2 (N1651, N1648, N1176);
xor XOR2 (N1652, N1644, N708);
xor XOR2 (N1653, N1637, N816);
nand NAND2 (N1654, N1622, N873);
or OR2 (N1655, N1652, N1521);
not NOT1 (N1656, N1649);
and AND3 (N1657, N1654, N1192, N781);
and AND3 (N1658, N1607, N43, N415);
and AND3 (N1659, N1647, N179, N912);
and AND2 (N1660, N1656, N1429);
xor XOR2 (N1661, N1650, N1384);
nand NAND3 (N1662, N1657, N1499, N712);
or OR2 (N1663, N1660, N988);
xor XOR2 (N1664, N1659, N623);
buf BUF1 (N1665, N1662);
not NOT1 (N1666, N1665);
and AND4 (N1667, N1658, N1277, N401, N1654);
nand NAND2 (N1668, N1666, N663);
xor XOR2 (N1669, N1655, N80);
nor NOR2 (N1670, N1664, N415);
not NOT1 (N1671, N1634);
nor NOR2 (N1672, N1661, N583);
buf BUF1 (N1673, N1667);
nand NAND2 (N1674, N1673, N676);
nor NOR3 (N1675, N1663, N585, N781);
buf BUF1 (N1676, N1669);
nor NOR3 (N1677, N1670, N539, N1382);
not NOT1 (N1678, N1672);
and AND4 (N1679, N1677, N1150, N994, N1315);
buf BUF1 (N1680, N1668);
not NOT1 (N1681, N1678);
nor NOR3 (N1682, N1651, N1546, N1017);
xor XOR2 (N1683, N1679, N924);
nand NAND2 (N1684, N1676, N1078);
nor NOR4 (N1685, N1641, N31, N1525, N470);
and AND3 (N1686, N1683, N776, N874);
nand NAND4 (N1687, N1682, N1236, N1394, N1359);
or OR3 (N1688, N1684, N440, N280);
nand NAND2 (N1689, N1675, N627);
buf BUF1 (N1690, N1688);
not NOT1 (N1691, N1689);
nand NAND3 (N1692, N1687, N1638, N543);
not NOT1 (N1693, N1671);
and AND2 (N1694, N1690, N414);
not NOT1 (N1695, N1686);
buf BUF1 (N1696, N1680);
nor NOR2 (N1697, N1694, N426);
not NOT1 (N1698, N1697);
buf BUF1 (N1699, N1685);
nor NOR4 (N1700, N1699, N1195, N928, N876);
xor XOR2 (N1701, N1691, N813);
nor NOR4 (N1702, N1695, N1595, N499, N1098);
or OR2 (N1703, N1693, N692);
nor NOR4 (N1704, N1700, N1112, N1633, N507);
nand NAND3 (N1705, N1698, N1520, N626);
or OR3 (N1706, N1653, N790, N34);
and AND3 (N1707, N1705, N857, N499);
nor NOR4 (N1708, N1704, N447, N145, N48);
and AND4 (N1709, N1696, N1459, N848, N323);
buf BUF1 (N1710, N1701);
not NOT1 (N1711, N1703);
not NOT1 (N1712, N1692);
nor NOR4 (N1713, N1674, N1304, N1151, N1304);
xor XOR2 (N1714, N1713, N226);
xor XOR2 (N1715, N1710, N168);
not NOT1 (N1716, N1711);
xor XOR2 (N1717, N1681, N981);
nor NOR3 (N1718, N1707, N1353, N1211);
nor NOR2 (N1719, N1702, N598);
and AND4 (N1720, N1715, N1341, N191, N546);
nor NOR2 (N1721, N1714, N606);
nor NOR4 (N1722, N1716, N107, N802, N1512);
xor XOR2 (N1723, N1722, N777);
nor NOR3 (N1724, N1723, N1695, N995);
not NOT1 (N1725, N1709);
buf BUF1 (N1726, N1708);
nor NOR2 (N1727, N1721, N887);
xor XOR2 (N1728, N1727, N1421);
or OR4 (N1729, N1728, N1128, N1670, N293);
or OR2 (N1730, N1717, N1235);
buf BUF1 (N1731, N1729);
and AND2 (N1732, N1726, N1096);
buf BUF1 (N1733, N1720);
buf BUF1 (N1734, N1718);
and AND4 (N1735, N1725, N392, N537, N742);
nor NOR2 (N1736, N1734, N92);
not NOT1 (N1737, N1712);
or OR3 (N1738, N1736, N1100, N560);
xor XOR2 (N1739, N1724, N189);
or OR2 (N1740, N1735, N645);
and AND4 (N1741, N1719, N915, N803, N508);
nand NAND3 (N1742, N1733, N78, N1568);
buf BUF1 (N1743, N1738);
nand NAND4 (N1744, N1730, N1724, N328, N294);
nand NAND2 (N1745, N1732, N911);
or OR2 (N1746, N1740, N306);
nand NAND3 (N1747, N1737, N326, N136);
nor NOR4 (N1748, N1731, N1698, N1517, N1126);
xor XOR2 (N1749, N1739, N119);
xor XOR2 (N1750, N1741, N1661);
nand NAND4 (N1751, N1749, N1121, N1266, N1456);
xor XOR2 (N1752, N1750, N1658);
nand NAND3 (N1753, N1745, N1557, N950);
nor NOR2 (N1754, N1747, N1023);
nor NOR4 (N1755, N1751, N497, N706, N422);
nand NAND2 (N1756, N1755, N883);
xor XOR2 (N1757, N1744, N303);
or OR4 (N1758, N1746, N377, N740, N75);
xor XOR2 (N1759, N1756, N328);
buf BUF1 (N1760, N1706);
nand NAND3 (N1761, N1753, N814, N497);
not NOT1 (N1762, N1759);
nand NAND2 (N1763, N1754, N1498);
or OR3 (N1764, N1760, N904, N1670);
buf BUF1 (N1765, N1761);
not NOT1 (N1766, N1765);
buf BUF1 (N1767, N1748);
nand NAND3 (N1768, N1742, N1055, N1685);
or OR4 (N1769, N1768, N1145, N255, N703);
buf BUF1 (N1770, N1763);
nor NOR2 (N1771, N1752, N254);
nand NAND2 (N1772, N1758, N1137);
nor NOR2 (N1773, N1772, N1558);
buf BUF1 (N1774, N1770);
buf BUF1 (N1775, N1757);
xor XOR2 (N1776, N1774, N308);
not NOT1 (N1777, N1764);
xor XOR2 (N1778, N1776, N1279);
buf BUF1 (N1779, N1778);
xor XOR2 (N1780, N1775, N1273);
xor XOR2 (N1781, N1771, N262);
xor XOR2 (N1782, N1777, N720);
nand NAND2 (N1783, N1769, N1167);
and AND4 (N1784, N1781, N206, N578, N1405);
nor NOR4 (N1785, N1762, N1138, N922, N1213);
nand NAND2 (N1786, N1743, N977);
nand NAND2 (N1787, N1779, N455);
nor NOR2 (N1788, N1773, N681);
nor NOR3 (N1789, N1784, N22, N566);
and AND2 (N1790, N1783, N1760);
xor XOR2 (N1791, N1788, N1748);
and AND4 (N1792, N1780, N170, N715, N1246);
or OR2 (N1793, N1791, N1411);
buf BUF1 (N1794, N1790);
not NOT1 (N1795, N1787);
buf BUF1 (N1796, N1767);
nand NAND3 (N1797, N1786, N512, N1178);
nand NAND4 (N1798, N1793, N1331, N1525, N665);
or OR3 (N1799, N1798, N638, N353);
and AND2 (N1800, N1794, N88);
not NOT1 (N1801, N1800);
nand NAND2 (N1802, N1789, N11);
nor NOR2 (N1803, N1795, N1272);
not NOT1 (N1804, N1782);
and AND3 (N1805, N1803, N1300, N690);
or OR4 (N1806, N1804, N246, N666, N1745);
xor XOR2 (N1807, N1796, N1530);
nand NAND2 (N1808, N1802, N1568);
and AND2 (N1809, N1785, N113);
nor NOR4 (N1810, N1799, N976, N1205, N1685);
not NOT1 (N1811, N1810);
nor NOR4 (N1812, N1811, N51, N635, N1330);
or OR4 (N1813, N1807, N1556, N1338, N938);
or OR3 (N1814, N1806, N1529, N1291);
buf BUF1 (N1815, N1814);
nor NOR2 (N1816, N1797, N485);
xor XOR2 (N1817, N1801, N1727);
xor XOR2 (N1818, N1815, N1547);
and AND3 (N1819, N1792, N1391, N620);
and AND3 (N1820, N1812, N720, N526);
nor NOR2 (N1821, N1816, N140);
not NOT1 (N1822, N1817);
nor NOR2 (N1823, N1821, N1732);
nor NOR4 (N1824, N1818, N539, N275, N1785);
nor NOR3 (N1825, N1808, N1538, N943);
xor XOR2 (N1826, N1766, N500);
and AND2 (N1827, N1826, N1274);
nor NOR3 (N1828, N1822, N1822, N869);
not NOT1 (N1829, N1823);
or OR4 (N1830, N1824, N1034, N737, N444);
or OR2 (N1831, N1828, N1676);
nand NAND3 (N1832, N1805, N1671, N785);
nor NOR2 (N1833, N1831, N371);
nor NOR4 (N1834, N1832, N459, N369, N904);
buf BUF1 (N1835, N1829);
nand NAND4 (N1836, N1835, N616, N238, N1068);
nand NAND3 (N1837, N1825, N872, N285);
or OR4 (N1838, N1833, N1788, N249, N217);
and AND2 (N1839, N1827, N977);
xor XOR2 (N1840, N1839, N1166);
and AND4 (N1841, N1836, N1577, N1075, N1479);
buf BUF1 (N1842, N1834);
not NOT1 (N1843, N1840);
buf BUF1 (N1844, N1842);
and AND3 (N1845, N1837, N1777, N295);
nor NOR4 (N1846, N1819, N1552, N159, N1816);
nand NAND4 (N1847, N1844, N362, N1231, N1787);
xor XOR2 (N1848, N1845, N630);
buf BUF1 (N1849, N1830);
not NOT1 (N1850, N1848);
xor XOR2 (N1851, N1813, N1573);
or OR4 (N1852, N1820, N1090, N1308, N766);
buf BUF1 (N1853, N1838);
nand NAND2 (N1854, N1849, N521);
xor XOR2 (N1855, N1841, N1128);
buf BUF1 (N1856, N1855);
xor XOR2 (N1857, N1856, N903);
not NOT1 (N1858, N1851);
buf BUF1 (N1859, N1852);
xor XOR2 (N1860, N1809, N1597);
or OR2 (N1861, N1847, N746);
nand NAND2 (N1862, N1843, N279);
xor XOR2 (N1863, N1854, N1372);
nor NOR3 (N1864, N1859, N1782, N910);
buf BUF1 (N1865, N1864);
buf BUF1 (N1866, N1853);
nand NAND4 (N1867, N1866, N1794, N70, N253);
nor NOR3 (N1868, N1865, N730, N533);
or OR4 (N1869, N1863, N1480, N1407, N1580);
nor NOR3 (N1870, N1850, N1033, N531);
buf BUF1 (N1871, N1870);
nor NOR3 (N1872, N1867, N916, N1665);
not NOT1 (N1873, N1871);
xor XOR2 (N1874, N1873, N920);
nor NOR2 (N1875, N1857, N345);
not NOT1 (N1876, N1846);
and AND4 (N1877, N1872, N958, N506, N809);
xor XOR2 (N1878, N1860, N973);
xor XOR2 (N1879, N1876, N1383);
not NOT1 (N1880, N1858);
buf BUF1 (N1881, N1879);
and AND2 (N1882, N1877, N1323);
buf BUF1 (N1883, N1881);
nor NOR4 (N1884, N1862, N51, N735, N863);
xor XOR2 (N1885, N1880, N773);
or OR2 (N1886, N1861, N794);
nand NAND3 (N1887, N1878, N648, N1633);
or OR4 (N1888, N1875, N1827, N1204, N303);
xor XOR2 (N1889, N1887, N845);
xor XOR2 (N1890, N1889, N801);
nand NAND2 (N1891, N1886, N1763);
and AND4 (N1892, N1885, N402, N1427, N1584);
nor NOR4 (N1893, N1890, N107, N1319, N909);
nand NAND2 (N1894, N1884, N1809);
buf BUF1 (N1895, N1888);
not NOT1 (N1896, N1883);
nand NAND4 (N1897, N1891, N1468, N1722, N1394);
nor NOR3 (N1898, N1893, N774, N624);
and AND4 (N1899, N1869, N634, N1100, N221);
xor XOR2 (N1900, N1892, N852);
and AND4 (N1901, N1868, N835, N1832, N912);
or OR2 (N1902, N1882, N837);
not NOT1 (N1903, N1896);
not NOT1 (N1904, N1895);
nor NOR4 (N1905, N1897, N1807, N1682, N242);
not NOT1 (N1906, N1905);
xor XOR2 (N1907, N1898, N1068);
not NOT1 (N1908, N1894);
nor NOR3 (N1909, N1902, N547, N971);
and AND3 (N1910, N1907, N969, N753);
or OR4 (N1911, N1910, N520, N569, N1382);
not NOT1 (N1912, N1911);
and AND3 (N1913, N1912, N1367, N144);
not NOT1 (N1914, N1906);
nor NOR3 (N1915, N1908, N1673, N1245);
nand NAND4 (N1916, N1914, N984, N1845, N1015);
buf BUF1 (N1917, N1916);
not NOT1 (N1918, N1913);
and AND3 (N1919, N1917, N1603, N86);
and AND4 (N1920, N1904, N917, N1610, N1163);
nand NAND3 (N1921, N1903, N1154, N1514);
xor XOR2 (N1922, N1900, N219);
xor XOR2 (N1923, N1919, N883);
buf BUF1 (N1924, N1909);
nand NAND4 (N1925, N1899, N566, N619, N63);
nand NAND4 (N1926, N1901, N1367, N135, N72);
or OR4 (N1927, N1874, N891, N138, N364);
not NOT1 (N1928, N1923);
or OR4 (N1929, N1928, N727, N786, N1187);
or OR2 (N1930, N1924, N1196);
and AND3 (N1931, N1918, N557, N1408);
buf BUF1 (N1932, N1926);
nand NAND2 (N1933, N1927, N380);
nand NAND2 (N1934, N1930, N460);
and AND2 (N1935, N1925, N1884);
and AND2 (N1936, N1929, N155);
nor NOR3 (N1937, N1922, N1254, N562);
xor XOR2 (N1938, N1920, N555);
buf BUF1 (N1939, N1915);
nor NOR2 (N1940, N1934, N694);
not NOT1 (N1941, N1931);
or OR3 (N1942, N1937, N1417, N1923);
xor XOR2 (N1943, N1942, N1885);
or OR2 (N1944, N1933, N1172);
and AND3 (N1945, N1921, N361, N268);
or OR2 (N1946, N1940, N1449);
buf BUF1 (N1947, N1946);
nand NAND3 (N1948, N1936, N1263, N1780);
nand NAND3 (N1949, N1943, N693, N1242);
xor XOR2 (N1950, N1949, N254);
xor XOR2 (N1951, N1948, N1421);
or OR2 (N1952, N1935, N823);
not NOT1 (N1953, N1944);
not NOT1 (N1954, N1953);
or OR4 (N1955, N1939, N731, N488, N181);
not NOT1 (N1956, N1932);
nand NAND3 (N1957, N1951, N844, N490);
xor XOR2 (N1958, N1955, N1777);
xor XOR2 (N1959, N1954, N1557);
xor XOR2 (N1960, N1950, N240);
buf BUF1 (N1961, N1957);
xor XOR2 (N1962, N1961, N1584);
nor NOR3 (N1963, N1960, N412, N1008);
or OR2 (N1964, N1945, N1312);
nand NAND2 (N1965, N1956, N60);
nor NOR2 (N1966, N1965, N1184);
nor NOR4 (N1967, N1964, N242, N166, N236);
nand NAND3 (N1968, N1952, N1637, N1754);
buf BUF1 (N1969, N1941);
nand NAND2 (N1970, N1947, N622);
and AND2 (N1971, N1962, N1843);
buf BUF1 (N1972, N1969);
not NOT1 (N1973, N1968);
xor XOR2 (N1974, N1971, N1164);
nand NAND3 (N1975, N1974, N1100, N296);
nor NOR3 (N1976, N1973, N752, N1962);
xor XOR2 (N1977, N1958, N35);
or OR3 (N1978, N1976, N1787, N571);
nor NOR2 (N1979, N1970, N765);
nor NOR2 (N1980, N1972, N701);
xor XOR2 (N1981, N1975, N1451);
and AND2 (N1982, N1967, N737);
and AND2 (N1983, N1963, N486);
and AND2 (N1984, N1977, N1019);
or OR3 (N1985, N1983, N1574, N361);
nand NAND2 (N1986, N1985, N1644);
not NOT1 (N1987, N1938);
xor XOR2 (N1988, N1987, N1342);
or OR2 (N1989, N1984, N647);
or OR3 (N1990, N1980, N1127, N1896);
or OR3 (N1991, N1959, N445, N736);
and AND4 (N1992, N1986, N747, N737, N1650);
or OR3 (N1993, N1982, N275, N1909);
nand NAND3 (N1994, N1992, N935, N512);
or OR2 (N1995, N1966, N923);
nor NOR2 (N1996, N1991, N360);
or OR2 (N1997, N1989, N689);
nor NOR2 (N1998, N1988, N887);
nand NAND4 (N1999, N1995, N369, N1352, N658);
and AND4 (N2000, N1997, N962, N713, N1091);
and AND2 (N2001, N1993, N217);
nor NOR3 (N2002, N1998, N1948, N1156);
nand NAND3 (N2003, N2001, N1939, N346);
nand NAND2 (N2004, N1996, N718);
not NOT1 (N2005, N1979);
not NOT1 (N2006, N2000);
xor XOR2 (N2007, N2005, N118);
not NOT1 (N2008, N1994);
nor NOR3 (N2009, N1990, N1703, N635);
nand NAND4 (N2010, N1999, N1484, N918, N1929);
or OR2 (N2011, N2006, N1108);
nand NAND2 (N2012, N2011, N1034);
and AND4 (N2013, N1978, N75, N995, N200);
and AND4 (N2014, N1981, N440, N875, N217);
nor NOR2 (N2015, N2014, N1705);
nand NAND3 (N2016, N2008, N40, N1985);
or OR3 (N2017, N2004, N460, N1980);
xor XOR2 (N2018, N2015, N1234);
nor NOR3 (N2019, N2009, N571, N171);
nor NOR2 (N2020, N2010, N184);
nand NAND3 (N2021, N2002, N1422, N760);
buf BUF1 (N2022, N2003);
xor XOR2 (N2023, N2019, N1664);
buf BUF1 (N2024, N2018);
or OR4 (N2025, N2023, N1088, N354, N1295);
xor XOR2 (N2026, N2025, N694);
nor NOR3 (N2027, N2013, N9, N134);
not NOT1 (N2028, N2012);
and AND2 (N2029, N2026, N792);
nand NAND2 (N2030, N2021, N1486);
or OR2 (N2031, N2029, N1983);
or OR4 (N2032, N2028, N271, N958, N426);
and AND4 (N2033, N2031, N1315, N1487, N1348);
buf BUF1 (N2034, N2017);
and AND2 (N2035, N2032, N134);
or OR2 (N2036, N2022, N1565);
not NOT1 (N2037, N2030);
and AND3 (N2038, N2033, N1578, N1911);
buf BUF1 (N2039, N2034);
and AND3 (N2040, N2038, N1312, N1700);
nand NAND3 (N2041, N2040, N1185, N1718);
nand NAND4 (N2042, N2027, N1513, N685, N96);
or OR4 (N2043, N2024, N1905, N1290, N1773);
or OR2 (N2044, N2037, N923);
and AND4 (N2045, N2039, N836, N1056, N1046);
nor NOR4 (N2046, N2036, N524, N1039, N122);
nand NAND4 (N2047, N2035, N306, N369, N1745);
xor XOR2 (N2048, N2020, N1540);
nor NOR3 (N2049, N2041, N121, N1731);
not NOT1 (N2050, N2047);
nand NAND4 (N2051, N2050, N934, N1997, N1390);
xor XOR2 (N2052, N2044, N882);
not NOT1 (N2053, N2051);
not NOT1 (N2054, N2042);
not NOT1 (N2055, N2046);
not NOT1 (N2056, N2048);
buf BUF1 (N2057, N2056);
not NOT1 (N2058, N2054);
and AND3 (N2059, N2045, N633, N1100);
not NOT1 (N2060, N2043);
buf BUF1 (N2061, N2057);
and AND2 (N2062, N2053, N949);
not NOT1 (N2063, N2058);
nand NAND4 (N2064, N2060, N1996, N1170, N412);
or OR3 (N2065, N2016, N530, N461);
buf BUF1 (N2066, N2049);
not NOT1 (N2067, N2063);
buf BUF1 (N2068, N2062);
or OR2 (N2069, N2065, N1122);
nand NAND2 (N2070, N2052, N194);
and AND3 (N2071, N2070, N1711, N1287);
or OR2 (N2072, N2059, N647);
or OR4 (N2073, N2072, N1793, N1791, N1269);
or OR4 (N2074, N2067, N671, N1120, N360);
nand NAND2 (N2075, N2055, N1258);
xor XOR2 (N2076, N2069, N1092);
xor XOR2 (N2077, N2071, N379);
not NOT1 (N2078, N2064);
nand NAND2 (N2079, N2068, N1751);
buf BUF1 (N2080, N2066);
buf BUF1 (N2081, N2073);
and AND4 (N2082, N2081, N15, N172, N580);
and AND2 (N2083, N2061, N969);
nand NAND4 (N2084, N2077, N1575, N1543, N4);
buf BUF1 (N2085, N2076);
or OR3 (N2086, N2074, N1786, N1475);
nand NAND3 (N2087, N2086, N340, N1802);
or OR2 (N2088, N2080, N838);
buf BUF1 (N2089, N2088);
buf BUF1 (N2090, N2082);
not NOT1 (N2091, N2083);
xor XOR2 (N2092, N2084, N1264);
buf BUF1 (N2093, N2090);
not NOT1 (N2094, N2093);
not NOT1 (N2095, N2085);
nor NOR2 (N2096, N2007, N106);
xor XOR2 (N2097, N2092, N256);
or OR4 (N2098, N2075, N842, N1485, N15);
nor NOR2 (N2099, N2094, N1496);
or OR2 (N2100, N2097, N834);
buf BUF1 (N2101, N2087);
and AND4 (N2102, N2078, N2039, N774, N1879);
buf BUF1 (N2103, N2098);
nand NAND2 (N2104, N2089, N243);
xor XOR2 (N2105, N2079, N1813);
or OR4 (N2106, N2095, N1516, N689, N373);
nand NAND4 (N2107, N2105, N1660, N191, N318);
and AND4 (N2108, N2099, N240, N1628, N1491);
not NOT1 (N2109, N2107);
or OR3 (N2110, N2108, N1994, N1504);
xor XOR2 (N2111, N2110, N1921);
nor NOR2 (N2112, N2111, N1002);
and AND2 (N2113, N2091, N862);
nand NAND2 (N2114, N2103, N1854);
not NOT1 (N2115, N2113);
buf BUF1 (N2116, N2106);
nor NOR4 (N2117, N2109, N1178, N586, N1578);
buf BUF1 (N2118, N2104);
or OR4 (N2119, N2114, N994, N1204, N1598);
xor XOR2 (N2120, N2096, N879);
or OR4 (N2121, N2118, N1818, N1387, N656);
xor XOR2 (N2122, N2121, N1508);
buf BUF1 (N2123, N2102);
buf BUF1 (N2124, N2122);
nand NAND4 (N2125, N2124, N1508, N2083, N73);
nor NOR3 (N2126, N2112, N700, N1370);
xor XOR2 (N2127, N2100, N2096);
nor NOR4 (N2128, N2126, N2125, N2126, N1813);
nand NAND3 (N2129, N1402, N1580, N384);
buf BUF1 (N2130, N2117);
not NOT1 (N2131, N2128);
and AND4 (N2132, N2127, N133, N439, N1073);
buf BUF1 (N2133, N2132);
xor XOR2 (N2134, N2129, N1542);
nand NAND2 (N2135, N2131, N1487);
xor XOR2 (N2136, N2119, N1258);
and AND3 (N2137, N2133, N1494, N2112);
nand NAND2 (N2138, N2135, N1352);
xor XOR2 (N2139, N2115, N1466);
nand NAND3 (N2140, N2138, N1866, N1970);
nor NOR3 (N2141, N2123, N420, N421);
xor XOR2 (N2142, N2139, N870);
nor NOR2 (N2143, N2137, N557);
and AND4 (N2144, N2134, N201, N19, N321);
xor XOR2 (N2145, N2141, N2036);
xor XOR2 (N2146, N2101, N93);
nor NOR3 (N2147, N2130, N514, N550);
nand NAND4 (N2148, N2120, N937, N23, N2034);
nand NAND2 (N2149, N2144, N1653);
buf BUF1 (N2150, N2147);
xor XOR2 (N2151, N2143, N1301);
buf BUF1 (N2152, N2150);
buf BUF1 (N2153, N2146);
not NOT1 (N2154, N2148);
buf BUF1 (N2155, N2152);
buf BUF1 (N2156, N2142);
buf BUF1 (N2157, N2116);
buf BUF1 (N2158, N2157);
or OR3 (N2159, N2136, N561, N1528);
nor NOR2 (N2160, N2159, N159);
buf BUF1 (N2161, N2155);
nand NAND3 (N2162, N2161, N184, N1013);
xor XOR2 (N2163, N2140, N839);
nand NAND2 (N2164, N2153, N966);
nand NAND4 (N2165, N2164, N2042, N428, N359);
xor XOR2 (N2166, N2149, N1887);
buf BUF1 (N2167, N2156);
or OR2 (N2168, N2160, N1190);
not NOT1 (N2169, N2162);
or OR4 (N2170, N2163, N662, N932, N2094);
nand NAND3 (N2171, N2154, N36, N937);
xor XOR2 (N2172, N2166, N122);
nor NOR4 (N2173, N2167, N2104, N2097, N40);
xor XOR2 (N2174, N2172, N1980);
nand NAND4 (N2175, N2145, N1327, N2012, N2155);
nor NOR2 (N2176, N2168, N1742);
nor NOR4 (N2177, N2158, N1154, N1297, N875);
and AND4 (N2178, N2174, N580, N194, N481);
buf BUF1 (N2179, N2165);
not NOT1 (N2180, N2151);
buf BUF1 (N2181, N2171);
buf BUF1 (N2182, N2169);
nand NAND3 (N2183, N2177, N1904, N1927);
not NOT1 (N2184, N2183);
xor XOR2 (N2185, N2175, N1480);
xor XOR2 (N2186, N2185, N228);
nor NOR4 (N2187, N2176, N1590, N2004, N1652);
nor NOR3 (N2188, N2186, N512, N1263);
not NOT1 (N2189, N2187);
nand NAND4 (N2190, N2173, N1703, N2034, N1953);
nor NOR4 (N2191, N2184, N1256, N1935, N1851);
xor XOR2 (N2192, N2182, N32);
xor XOR2 (N2193, N2180, N988);
xor XOR2 (N2194, N2188, N1239);
nor NOR2 (N2195, N2178, N1530);
xor XOR2 (N2196, N2181, N1183);
nor NOR4 (N2197, N2195, N592, N1289, N973);
or OR4 (N2198, N2170, N1668, N901, N1219);
nor NOR2 (N2199, N2189, N851);
nand NAND4 (N2200, N2191, N1077, N1050, N20);
not NOT1 (N2201, N2194);
nor NOR4 (N2202, N2190, N1836, N1601, N716);
buf BUF1 (N2203, N2197);
not NOT1 (N2204, N2192);
nand NAND2 (N2205, N2203, N1418);
or OR4 (N2206, N2198, N395, N672, N1962);
buf BUF1 (N2207, N2205);
or OR4 (N2208, N2201, N1318, N440, N977);
buf BUF1 (N2209, N2179);
xor XOR2 (N2210, N2200, N1008);
buf BUF1 (N2211, N2202);
xor XOR2 (N2212, N2193, N972);
nor NOR3 (N2213, N2212, N1048, N1883);
buf BUF1 (N2214, N2211);
or OR3 (N2215, N2207, N1693, N492);
or OR3 (N2216, N2199, N302, N711);
buf BUF1 (N2217, N2210);
and AND2 (N2218, N2208, N221);
buf BUF1 (N2219, N2204);
and AND3 (N2220, N2218, N1549, N906);
and AND3 (N2221, N2219, N334, N1975);
nand NAND3 (N2222, N2213, N1316, N2111);
not NOT1 (N2223, N2220);
or OR4 (N2224, N2221, N87, N1274, N1921);
xor XOR2 (N2225, N2217, N646);
xor XOR2 (N2226, N2206, N820);
nor NOR4 (N2227, N2196, N1435, N2156, N1039);
not NOT1 (N2228, N2225);
and AND4 (N2229, N2209, N934, N1936, N831);
nor NOR3 (N2230, N2228, N1382, N1439);
and AND4 (N2231, N2222, N466, N890, N924);
or OR3 (N2232, N2229, N1097, N920);
and AND3 (N2233, N2224, N1827, N1521);
buf BUF1 (N2234, N2216);
and AND4 (N2235, N2231, N219, N2160, N1898);
nor NOR3 (N2236, N2233, N358, N1916);
and AND4 (N2237, N2236, N170, N36, N190);
buf BUF1 (N2238, N2215);
buf BUF1 (N2239, N2238);
or OR4 (N2240, N2230, N592, N788, N542);
xor XOR2 (N2241, N2232, N1221);
buf BUF1 (N2242, N2241);
xor XOR2 (N2243, N2227, N728);
nor NOR4 (N2244, N2226, N1847, N884, N387);
nor NOR4 (N2245, N2239, N65, N389, N111);
and AND4 (N2246, N2223, N139, N1691, N1380);
buf BUF1 (N2247, N2242);
or OR3 (N2248, N2244, N255, N894);
buf BUF1 (N2249, N2234);
and AND4 (N2250, N2246, N1965, N847, N850);
or OR4 (N2251, N2249, N1081, N888, N1377);
nor NOR2 (N2252, N2235, N2159);
nor NOR2 (N2253, N2237, N1153);
nor NOR2 (N2254, N2251, N160);
and AND3 (N2255, N2214, N1304, N458);
nand NAND4 (N2256, N2253, N1047, N615, N595);
xor XOR2 (N2257, N2255, N1568);
or OR4 (N2258, N2250, N1207, N488, N1898);
or OR3 (N2259, N2252, N1522, N448);
xor XOR2 (N2260, N2256, N1379);
nor NOR4 (N2261, N2240, N952, N867, N2127);
xor XOR2 (N2262, N2257, N1410);
buf BUF1 (N2263, N2259);
and AND3 (N2264, N2262, N2078, N237);
not NOT1 (N2265, N2248);
not NOT1 (N2266, N2260);
buf BUF1 (N2267, N2245);
xor XOR2 (N2268, N2254, N1631);
and AND2 (N2269, N2258, N1506);
nor NOR2 (N2270, N2268, N1082);
nand NAND2 (N2271, N2265, N1488);
or OR3 (N2272, N2264, N2226, N1707);
or OR3 (N2273, N2272, N1429, N23);
nor NOR3 (N2274, N2270, N1862, N664);
buf BUF1 (N2275, N2274);
or OR4 (N2276, N2247, N1158, N741, N2050);
nor NOR3 (N2277, N2243, N2069, N681);
not NOT1 (N2278, N2263);
not NOT1 (N2279, N2277);
xor XOR2 (N2280, N2278, N1910);
not NOT1 (N2281, N2267);
and AND3 (N2282, N2269, N1683, N327);
or OR2 (N2283, N2280, N858);
or OR4 (N2284, N2279, N1547, N1289, N585);
xor XOR2 (N2285, N2281, N2083);
not NOT1 (N2286, N2282);
xor XOR2 (N2287, N2285, N785);
not NOT1 (N2288, N2266);
nor NOR2 (N2289, N2261, N1193);
or OR3 (N2290, N2284, N1282, N59);
not NOT1 (N2291, N2287);
nor NOR3 (N2292, N2271, N288, N257);
not NOT1 (N2293, N2276);
and AND4 (N2294, N2275, N142, N141, N567);
not NOT1 (N2295, N2288);
nand NAND2 (N2296, N2289, N47);
not NOT1 (N2297, N2291);
nor NOR2 (N2298, N2296, N1272);
buf BUF1 (N2299, N2294);
or OR4 (N2300, N2290, N150, N2004, N2237);
nor NOR3 (N2301, N2292, N1749, N771);
buf BUF1 (N2302, N2301);
xor XOR2 (N2303, N2283, N1227);
and AND4 (N2304, N2300, N373, N1377, N1750);
xor XOR2 (N2305, N2302, N432);
nor NOR2 (N2306, N2295, N727);
nor NOR3 (N2307, N2293, N598, N2272);
nand NAND2 (N2308, N2305, N445);
or OR3 (N2309, N2303, N282, N1068);
xor XOR2 (N2310, N2309, N850);
and AND4 (N2311, N2298, N1913, N1091, N1555);
nand NAND3 (N2312, N2306, N2029, N61);
not NOT1 (N2313, N2312);
and AND4 (N2314, N2313, N882, N928, N692);
nand NAND2 (N2315, N2311, N1926);
nand NAND2 (N2316, N2315, N1105);
not NOT1 (N2317, N2316);
nand NAND2 (N2318, N2317, N1268);
xor XOR2 (N2319, N2297, N39);
xor XOR2 (N2320, N2314, N853);
nor NOR3 (N2321, N2286, N1566, N2092);
nor NOR2 (N2322, N2307, N1740);
nor NOR2 (N2323, N2319, N380);
not NOT1 (N2324, N2321);
xor XOR2 (N2325, N2304, N403);
or OR3 (N2326, N2323, N436, N2154);
buf BUF1 (N2327, N2320);
buf BUF1 (N2328, N2327);
or OR3 (N2329, N2326, N104, N1030);
buf BUF1 (N2330, N2310);
xor XOR2 (N2331, N2330, N2072);
not NOT1 (N2332, N2329);
and AND4 (N2333, N2324, N436, N13, N1750);
and AND4 (N2334, N2299, N2116, N400, N143);
not NOT1 (N2335, N2333);
xor XOR2 (N2336, N2334, N684);
buf BUF1 (N2337, N2322);
buf BUF1 (N2338, N2318);
nor NOR2 (N2339, N2273, N1413);
not NOT1 (N2340, N2335);
not NOT1 (N2341, N2336);
buf BUF1 (N2342, N2341);
and AND4 (N2343, N2331, N698, N1722, N476);
or OR2 (N2344, N2337, N1392);
and AND2 (N2345, N2332, N595);
or OR3 (N2346, N2325, N630, N106);
or OR3 (N2347, N2342, N1582, N384);
nand NAND4 (N2348, N2345, N1426, N519, N2151);
and AND4 (N2349, N2338, N2217, N1468, N1649);
and AND4 (N2350, N2343, N1629, N676, N2269);
buf BUF1 (N2351, N2347);
and AND2 (N2352, N2328, N1411);
nand NAND3 (N2353, N2351, N1979, N2030);
and AND3 (N2354, N2346, N1967, N621);
nor NOR4 (N2355, N2352, N439, N487, N354);
buf BUF1 (N2356, N2340);
or OR4 (N2357, N2349, N1786, N1107, N2190);
buf BUF1 (N2358, N2357);
xor XOR2 (N2359, N2356, N1652);
and AND4 (N2360, N2348, N1156, N477, N344);
or OR2 (N2361, N2350, N1504);
nand NAND2 (N2362, N2360, N810);
or OR3 (N2363, N2362, N2199, N1380);
xor XOR2 (N2364, N2355, N2082);
or OR2 (N2365, N2339, N620);
xor XOR2 (N2366, N2344, N2201);
nor NOR3 (N2367, N2354, N356, N1104);
or OR4 (N2368, N2364, N2044, N60, N2114);
xor XOR2 (N2369, N2363, N1752);
and AND3 (N2370, N2361, N862, N1994);
nand NAND4 (N2371, N2366, N33, N108, N852);
not NOT1 (N2372, N2359);
nand NAND4 (N2373, N2353, N800, N1495, N296);
or OR4 (N2374, N2367, N1641, N2025, N1417);
not NOT1 (N2375, N2374);
nand NAND3 (N2376, N2370, N468, N1736);
and AND3 (N2377, N2358, N1878, N184);
xor XOR2 (N2378, N2368, N870);
nand NAND4 (N2379, N2372, N1699, N471, N1654);
nor NOR3 (N2380, N2308, N1089, N2300);
not NOT1 (N2381, N2376);
nor NOR3 (N2382, N2373, N1608, N936);
or OR4 (N2383, N2369, N1445, N190, N1940);
nand NAND3 (N2384, N2380, N306, N1239);
and AND2 (N2385, N2375, N2051);
or OR2 (N2386, N2385, N701);
xor XOR2 (N2387, N2365, N855);
nor NOR3 (N2388, N2377, N2064, N44);
nand NAND3 (N2389, N2382, N307, N684);
not NOT1 (N2390, N2386);
nand NAND2 (N2391, N2383, N1705);
or OR3 (N2392, N2381, N846, N1293);
or OR3 (N2393, N2378, N2033, N1317);
buf BUF1 (N2394, N2371);
nor NOR3 (N2395, N2389, N280, N708);
buf BUF1 (N2396, N2392);
nor NOR2 (N2397, N2395, N469);
nand NAND2 (N2398, N2393, N2314);
nand NAND2 (N2399, N2397, N166);
nand NAND4 (N2400, N2388, N1288, N2309, N1376);
nand NAND3 (N2401, N2396, N854, N501);
buf BUF1 (N2402, N2401);
not NOT1 (N2403, N2379);
nor NOR2 (N2404, N2391, N821);
buf BUF1 (N2405, N2403);
nand NAND3 (N2406, N2404, N1481, N273);
nand NAND3 (N2407, N2390, N500, N1670);
not NOT1 (N2408, N2398);
nand NAND4 (N2409, N2405, N599, N912, N9);
nand NAND3 (N2410, N2399, N78, N1330);
nand NAND4 (N2411, N2408, N2053, N1095, N2050);
buf BUF1 (N2412, N2402);
xor XOR2 (N2413, N2407, N801);
or OR2 (N2414, N2400, N291);
or OR4 (N2415, N2384, N839, N1175, N1281);
xor XOR2 (N2416, N2412, N1594);
nor NOR2 (N2417, N2406, N1936);
not NOT1 (N2418, N2409);
nor NOR3 (N2419, N2415, N1877, N982);
buf BUF1 (N2420, N2410);
buf BUF1 (N2421, N2419);
nor NOR4 (N2422, N2417, N2272, N278, N84);
and AND2 (N2423, N2416, N1392);
nand NAND4 (N2424, N2414, N2419, N1796, N1224);
xor XOR2 (N2425, N2422, N477);
nand NAND4 (N2426, N2413, N2421, N1949, N976);
not NOT1 (N2427, N324);
nor NOR3 (N2428, N2427, N2254, N2342);
buf BUF1 (N2429, N2394);
nand NAND4 (N2430, N2425, N672, N834, N2016);
and AND4 (N2431, N2430, N1273, N868, N2188);
not NOT1 (N2432, N2431);
or OR2 (N2433, N2432, N1685);
and AND3 (N2434, N2418, N241, N699);
and AND2 (N2435, N2434, N288);
nor NOR4 (N2436, N2433, N2329, N2304, N2422);
buf BUF1 (N2437, N2436);
not NOT1 (N2438, N2426);
buf BUF1 (N2439, N2424);
not NOT1 (N2440, N2435);
not NOT1 (N2441, N2429);
xor XOR2 (N2442, N2423, N754);
not NOT1 (N2443, N2441);
nor NOR4 (N2444, N2437, N1807, N2440, N1496);
xor XOR2 (N2445, N2257, N2235);
and AND3 (N2446, N2445, N106, N753);
buf BUF1 (N2447, N2411);
nor NOR2 (N2448, N2443, N1051);
not NOT1 (N2449, N2428);
and AND3 (N2450, N2420, N355, N60);
not NOT1 (N2451, N2438);
not NOT1 (N2452, N2450);
nand NAND4 (N2453, N2439, N485, N1280, N474);
nand NAND2 (N2454, N2451, N110);
not NOT1 (N2455, N2444);
not NOT1 (N2456, N2447);
and AND4 (N2457, N2452, N1381, N2153, N1381);
xor XOR2 (N2458, N2453, N524);
and AND4 (N2459, N2457, N1283, N2307, N2094);
nand NAND4 (N2460, N2448, N977, N2167, N1840);
nand NAND2 (N2461, N2446, N2023);
xor XOR2 (N2462, N2456, N1393);
not NOT1 (N2463, N2461);
not NOT1 (N2464, N2460);
nor NOR4 (N2465, N2455, N602, N1453, N1957);
xor XOR2 (N2466, N2462, N1310);
nor NOR3 (N2467, N2387, N1425, N1440);
buf BUF1 (N2468, N2458);
nor NOR4 (N2469, N2459, N729, N2373, N1941);
or OR3 (N2470, N2469, N1265, N508);
xor XOR2 (N2471, N2466, N2277);
or OR2 (N2472, N2454, N2309);
nor NOR3 (N2473, N2464, N661, N1312);
not NOT1 (N2474, N2471);
or OR3 (N2475, N2474, N2187, N317);
not NOT1 (N2476, N2470);
xor XOR2 (N2477, N2449, N599);
and AND3 (N2478, N2475, N2198, N2415);
not NOT1 (N2479, N2468);
nand NAND2 (N2480, N2477, N305);
and AND4 (N2481, N2472, N221, N1764, N204);
and AND4 (N2482, N2479, N1995, N651, N2289);
buf BUF1 (N2483, N2478);
and AND4 (N2484, N2482, N502, N1650, N2369);
nand NAND2 (N2485, N2484, N1059);
not NOT1 (N2486, N2483);
xor XOR2 (N2487, N2486, N628);
not NOT1 (N2488, N2487);
xor XOR2 (N2489, N2481, N2396);
not NOT1 (N2490, N2488);
not NOT1 (N2491, N2473);
buf BUF1 (N2492, N2490);
nand NAND4 (N2493, N2492, N1899, N1254, N991);
not NOT1 (N2494, N2480);
nand NAND3 (N2495, N2442, N652, N952);
not NOT1 (N2496, N2476);
buf BUF1 (N2497, N2465);
or OR3 (N2498, N2493, N1237, N2444);
not NOT1 (N2499, N2494);
buf BUF1 (N2500, N2497);
xor XOR2 (N2501, N2498, N521);
not NOT1 (N2502, N2489);
nor NOR2 (N2503, N2495, N1084);
and AND3 (N2504, N2503, N1581, N180);
or OR2 (N2505, N2502, N1770);
not NOT1 (N2506, N2467);
or OR2 (N2507, N2504, N501);
and AND4 (N2508, N2500, N732, N672, N2320);
not NOT1 (N2509, N2506);
or OR4 (N2510, N2491, N1759, N57, N1980);
not NOT1 (N2511, N2505);
or OR3 (N2512, N2463, N303, N1315);
and AND2 (N2513, N2501, N2389);
not NOT1 (N2514, N2507);
not NOT1 (N2515, N2496);
buf BUF1 (N2516, N2512);
nand NAND4 (N2517, N2516, N614, N1334, N1671);
not NOT1 (N2518, N2509);
or OR4 (N2519, N2517, N363, N290, N1709);
buf BUF1 (N2520, N2515);
buf BUF1 (N2521, N2510);
or OR3 (N2522, N2485, N2068, N1110);
nand NAND3 (N2523, N2519, N165, N1893);
buf BUF1 (N2524, N2499);
nor NOR3 (N2525, N2508, N1578, N1002);
buf BUF1 (N2526, N2518);
buf BUF1 (N2527, N2526);
buf BUF1 (N2528, N2523);
or OR4 (N2529, N2520, N702, N345, N1767);
or OR4 (N2530, N2525, N1539, N906, N1799);
nor NOR3 (N2531, N2522, N508, N1816);
xor XOR2 (N2532, N2511, N1008);
nor NOR4 (N2533, N2531, N220, N962, N785);
and AND4 (N2534, N2530, N950, N578, N1760);
and AND3 (N2535, N2514, N1987, N2327);
buf BUF1 (N2536, N2524);
and AND2 (N2537, N2532, N1048);
nand NAND2 (N2538, N2535, N2392);
xor XOR2 (N2539, N2528, N483);
or OR4 (N2540, N2534, N1388, N610, N1790);
buf BUF1 (N2541, N2536);
and AND4 (N2542, N2533, N1542, N1906, N1087);
xor XOR2 (N2543, N2537, N1948);
and AND4 (N2544, N2539, N1649, N1318, N2366);
nor NOR4 (N2545, N2521, N1693, N1340, N1252);
nor NOR2 (N2546, N2543, N5);
or OR4 (N2547, N2538, N880, N1999, N1374);
not NOT1 (N2548, N2545);
not NOT1 (N2549, N2541);
nor NOR2 (N2550, N2544, N2402);
nand NAND3 (N2551, N2546, N1851, N925);
nand NAND2 (N2552, N2542, N2269);
xor XOR2 (N2553, N2548, N1932);
nor NOR2 (N2554, N2547, N655);
or OR4 (N2555, N2540, N1529, N1827, N1051);
nor NOR2 (N2556, N2553, N1906);
and AND4 (N2557, N2527, N1479, N982, N801);
nand NAND2 (N2558, N2554, N1191);
or OR4 (N2559, N2555, N2208, N700, N2453);
xor XOR2 (N2560, N2559, N96);
or OR4 (N2561, N2560, N1210, N1872, N1725);
buf BUF1 (N2562, N2513);
buf BUF1 (N2563, N2557);
nand NAND3 (N2564, N2549, N1400, N2355);
nor NOR3 (N2565, N2529, N1124, N607);
or OR3 (N2566, N2564, N2464, N689);
buf BUF1 (N2567, N2550);
not NOT1 (N2568, N2561);
and AND4 (N2569, N2552, N342, N98, N2175);
not NOT1 (N2570, N2567);
and AND4 (N2571, N2562, N956, N65, N1817);
nand NAND4 (N2572, N2571, N1392, N1110, N1462);
nand NAND2 (N2573, N2570, N937);
not NOT1 (N2574, N2566);
and AND3 (N2575, N2551, N2027, N1317);
xor XOR2 (N2576, N2575, N889);
nand NAND4 (N2577, N2568, N172, N298, N2164);
nor NOR2 (N2578, N2572, N2256);
xor XOR2 (N2579, N2558, N224);
and AND4 (N2580, N2578, N1857, N575, N802);
and AND3 (N2581, N2563, N135, N2070);
not NOT1 (N2582, N2573);
and AND3 (N2583, N2579, N1941, N1648);
not NOT1 (N2584, N2574);
and AND2 (N2585, N2565, N1161);
not NOT1 (N2586, N2582);
nand NAND2 (N2587, N2585, N389);
or OR3 (N2588, N2587, N1335, N1679);
nor NOR2 (N2589, N2581, N184);
nand NAND3 (N2590, N2588, N436, N1387);
not NOT1 (N2591, N2589);
and AND2 (N2592, N2586, N1561);
buf BUF1 (N2593, N2576);
nor NOR4 (N2594, N2577, N664, N2572, N2086);
not NOT1 (N2595, N2592);
buf BUF1 (N2596, N2580);
xor XOR2 (N2597, N2556, N550);
buf BUF1 (N2598, N2595);
buf BUF1 (N2599, N2583);
nand NAND4 (N2600, N2599, N1511, N1022, N1644);
or OR3 (N2601, N2593, N2028, N1384);
xor XOR2 (N2602, N2591, N1833);
and AND3 (N2603, N2598, N522, N962);
or OR2 (N2604, N2600, N1357);
nand NAND2 (N2605, N2603, N1855);
nor NOR4 (N2606, N2601, N2103, N2415, N1991);
xor XOR2 (N2607, N2597, N789);
xor XOR2 (N2608, N2569, N2010);
not NOT1 (N2609, N2590);
nor NOR3 (N2610, N2608, N325, N579);
buf BUF1 (N2611, N2584);
or OR2 (N2612, N2607, N1351);
not NOT1 (N2613, N2594);
or OR2 (N2614, N2611, N107);
not NOT1 (N2615, N2606);
nand NAND2 (N2616, N2605, N1792);
xor XOR2 (N2617, N2612, N1753);
nand NAND4 (N2618, N2609, N1988, N116, N2562);
buf BUF1 (N2619, N2610);
nand NAND3 (N2620, N2604, N2357, N230);
xor XOR2 (N2621, N2617, N2344);
xor XOR2 (N2622, N2620, N2492);
and AND2 (N2623, N2616, N2439);
xor XOR2 (N2624, N2623, N2503);
nand NAND4 (N2625, N2621, N571, N2533, N2511);
not NOT1 (N2626, N2618);
nor NOR4 (N2627, N2613, N1884, N1084, N1660);
nor NOR3 (N2628, N2596, N2080, N1917);
xor XOR2 (N2629, N2619, N218);
xor XOR2 (N2630, N2602, N1174);
nor NOR2 (N2631, N2628, N2076);
or OR4 (N2632, N2629, N285, N1646, N1387);
nand NAND4 (N2633, N2627, N1419, N2543, N545);
xor XOR2 (N2634, N2625, N1982);
nor NOR3 (N2635, N2626, N639, N2477);
or OR2 (N2636, N2624, N275);
buf BUF1 (N2637, N2615);
nand NAND3 (N2638, N2633, N1658, N1298);
or OR4 (N2639, N2614, N419, N974, N1343);
nor NOR2 (N2640, N2637, N961);
nand NAND3 (N2641, N2636, N545, N2224);
buf BUF1 (N2642, N2632);
nor NOR2 (N2643, N2622, N2569);
nor NOR3 (N2644, N2635, N362, N438);
xor XOR2 (N2645, N2643, N424);
buf BUF1 (N2646, N2639);
and AND4 (N2647, N2640, N1364, N1151, N1849);
buf BUF1 (N2648, N2642);
and AND4 (N2649, N2645, N1281, N1151, N447);
or OR4 (N2650, N2638, N2266, N1467, N1019);
nor NOR3 (N2651, N2647, N1464, N2048);
buf BUF1 (N2652, N2646);
not NOT1 (N2653, N2630);
buf BUF1 (N2654, N2648);
and AND4 (N2655, N2634, N1018, N1728, N377);
buf BUF1 (N2656, N2653);
or OR4 (N2657, N2644, N1573, N1996, N2523);
not NOT1 (N2658, N2655);
nor NOR2 (N2659, N2650, N1628);
not NOT1 (N2660, N2651);
nand NAND4 (N2661, N2659, N1902, N2269, N630);
xor XOR2 (N2662, N2661, N239);
nor NOR3 (N2663, N2656, N417, N241);
not NOT1 (N2664, N2657);
nor NOR4 (N2665, N2660, N404, N1990, N2039);
and AND3 (N2666, N2652, N2291, N595);
or OR3 (N2667, N2654, N1823, N2585);
or OR3 (N2668, N2664, N1580, N814);
xor XOR2 (N2669, N2663, N1703);
buf BUF1 (N2670, N2669);
nand NAND3 (N2671, N2668, N2030, N1232);
buf BUF1 (N2672, N2631);
and AND3 (N2673, N2662, N141, N1790);
nand NAND2 (N2674, N2666, N236);
nand NAND4 (N2675, N2641, N996, N199, N1102);
nand NAND2 (N2676, N2675, N482);
xor XOR2 (N2677, N2667, N2589);
not NOT1 (N2678, N2674);
buf BUF1 (N2679, N2658);
xor XOR2 (N2680, N2677, N1368);
or OR2 (N2681, N2673, N867);
buf BUF1 (N2682, N2670);
nor NOR2 (N2683, N2649, N1940);
not NOT1 (N2684, N2681);
nand NAND2 (N2685, N2684, N1548);
nand NAND2 (N2686, N2665, N1424);
nand NAND4 (N2687, N2685, N485, N279, N1420);
not NOT1 (N2688, N2671);
or OR3 (N2689, N2678, N1884, N2403);
xor XOR2 (N2690, N2682, N1725);
buf BUF1 (N2691, N2689);
and AND3 (N2692, N2683, N1139, N1102);
and AND3 (N2693, N2688, N1734, N304);
xor XOR2 (N2694, N2679, N1498);
and AND3 (N2695, N2676, N830, N1904);
xor XOR2 (N2696, N2693, N911);
nand NAND3 (N2697, N2696, N355, N282);
and AND4 (N2698, N2680, N888, N272, N2011);
and AND3 (N2699, N2687, N2246, N2532);
nand NAND4 (N2700, N2697, N2402, N1947, N1767);
nor NOR3 (N2701, N2672, N2183, N1193);
nand NAND2 (N2702, N2694, N673);
or OR4 (N2703, N2690, N1154, N1784, N2015);
nand NAND3 (N2704, N2700, N1683, N2633);
nand NAND3 (N2705, N2691, N18, N2130);
nand NAND3 (N2706, N2702, N627, N2615);
xor XOR2 (N2707, N2686, N2167);
and AND4 (N2708, N2695, N2519, N2065, N1432);
nand NAND4 (N2709, N2703, N169, N863, N827);
and AND4 (N2710, N2708, N1511, N727, N796);
nand NAND3 (N2711, N2709, N2049, N1330);
and AND3 (N2712, N2710, N1296, N1515);
or OR3 (N2713, N2706, N1123, N218);
and AND4 (N2714, N2713, N1690, N896, N2710);
buf BUF1 (N2715, N2692);
not NOT1 (N2716, N2707);
nor NOR3 (N2717, N2699, N487, N285);
or OR4 (N2718, N2698, N1577, N938, N1482);
not NOT1 (N2719, N2712);
not NOT1 (N2720, N2718);
not NOT1 (N2721, N2720);
and AND4 (N2722, N2701, N2435, N1343, N2386);
not NOT1 (N2723, N2719);
xor XOR2 (N2724, N2705, N836);
xor XOR2 (N2725, N2704, N2053);
buf BUF1 (N2726, N2715);
buf BUF1 (N2727, N2711);
nor NOR3 (N2728, N2724, N2139, N723);
not NOT1 (N2729, N2714);
buf BUF1 (N2730, N2725);
buf BUF1 (N2731, N2723);
not NOT1 (N2732, N2730);
nor NOR2 (N2733, N2732, N1367);
xor XOR2 (N2734, N2717, N164);
xor XOR2 (N2735, N2728, N1322);
xor XOR2 (N2736, N2729, N963);
nor NOR4 (N2737, N2716, N945, N1381, N1418);
and AND2 (N2738, N2737, N2034);
and AND2 (N2739, N2733, N308);
nand NAND3 (N2740, N2721, N616, N2623);
buf BUF1 (N2741, N2735);
or OR4 (N2742, N2738, N1042, N1141, N2215);
and AND4 (N2743, N2741, N1751, N1835, N1598);
nor NOR2 (N2744, N2734, N1463);
nor NOR2 (N2745, N2739, N1893);
nand NAND4 (N2746, N2743, N2633, N1214, N1422);
nand NAND4 (N2747, N2742, N1624, N1138, N1040);
and AND4 (N2748, N2731, N2348, N650, N2389);
nand NAND4 (N2749, N2727, N1930, N1009, N300);
not NOT1 (N2750, N2722);
xor XOR2 (N2751, N2744, N598);
or OR2 (N2752, N2726, N365);
buf BUF1 (N2753, N2751);
not NOT1 (N2754, N2746);
buf BUF1 (N2755, N2752);
and AND4 (N2756, N2736, N554, N1229, N2684);
and AND3 (N2757, N2740, N1089, N2480);
xor XOR2 (N2758, N2757, N1131);
nand NAND3 (N2759, N2755, N763, N1523);
and AND3 (N2760, N2748, N2165, N1924);
nor NOR2 (N2761, N2749, N2512);
xor XOR2 (N2762, N2760, N1771);
buf BUF1 (N2763, N2750);
xor XOR2 (N2764, N2762, N839);
not NOT1 (N2765, N2756);
or OR3 (N2766, N2763, N995, N1817);
or OR4 (N2767, N2747, N2597, N1876, N2064);
or OR2 (N2768, N2758, N1408);
buf BUF1 (N2769, N2745);
xor XOR2 (N2770, N2764, N493);
not NOT1 (N2771, N2770);
nand NAND2 (N2772, N2765, N2344);
or OR4 (N2773, N2768, N584, N1585, N132);
not NOT1 (N2774, N2753);
buf BUF1 (N2775, N2774);
nand NAND2 (N2776, N2773, N1059);
not NOT1 (N2777, N2771);
nand NAND2 (N2778, N2776, N2644);
not NOT1 (N2779, N2761);
or OR3 (N2780, N2775, N1561, N1243);
nand NAND4 (N2781, N2759, N1034, N2167, N382);
xor XOR2 (N2782, N2772, N2584);
nor NOR3 (N2783, N2767, N1570, N1813);
xor XOR2 (N2784, N2781, N1194);
or OR2 (N2785, N2784, N269);
nand NAND3 (N2786, N2766, N1485, N2460);
buf BUF1 (N2787, N2754);
not NOT1 (N2788, N2787);
nand NAND3 (N2789, N2778, N2099, N1225);
nor NOR2 (N2790, N2769, N402);
not NOT1 (N2791, N2789);
not NOT1 (N2792, N2790);
and AND2 (N2793, N2779, N1628);
nor NOR2 (N2794, N2783, N449);
not NOT1 (N2795, N2791);
and AND4 (N2796, N2795, N1717, N720, N1464);
xor XOR2 (N2797, N2780, N19);
nand NAND3 (N2798, N2782, N976, N795);
and AND4 (N2799, N2788, N1616, N578, N892);
buf BUF1 (N2800, N2777);
and AND2 (N2801, N2786, N2564);
nand NAND2 (N2802, N2797, N2556);
and AND3 (N2803, N2800, N2458, N628);
nor NOR3 (N2804, N2803, N494, N1909);
buf BUF1 (N2805, N2802);
not NOT1 (N2806, N2794);
nand NAND3 (N2807, N2793, N2666, N73);
not NOT1 (N2808, N2796);
buf BUF1 (N2809, N2805);
buf BUF1 (N2810, N2799);
buf BUF1 (N2811, N2792);
not NOT1 (N2812, N2804);
nand NAND4 (N2813, N2806, N1488, N2770, N2248);
buf BUF1 (N2814, N2811);
buf BUF1 (N2815, N2809);
xor XOR2 (N2816, N2785, N2042);
buf BUF1 (N2817, N2812);
or OR4 (N2818, N2810, N300, N375, N583);
buf BUF1 (N2819, N2818);
nand NAND4 (N2820, N2816, N1692, N269, N1423);
not NOT1 (N2821, N2807);
or OR2 (N2822, N2815, N952);
xor XOR2 (N2823, N2820, N2644);
xor XOR2 (N2824, N2822, N2600);
nor NOR3 (N2825, N2823, N2601, N2262);
xor XOR2 (N2826, N2801, N1926);
buf BUF1 (N2827, N2814);
not NOT1 (N2828, N2808);
buf BUF1 (N2829, N2824);
not NOT1 (N2830, N2819);
buf BUF1 (N2831, N2798);
not NOT1 (N2832, N2829);
or OR4 (N2833, N2813, N1060, N1830, N2144);
nand NAND2 (N2834, N2828, N197);
buf BUF1 (N2835, N2832);
nand NAND3 (N2836, N2821, N547, N1778);
buf BUF1 (N2837, N2826);
and AND3 (N2838, N2831, N165, N1326);
or OR4 (N2839, N2838, N1758, N2427, N2684);
nor NOR2 (N2840, N2833, N2786);
not NOT1 (N2841, N2825);
nor NOR4 (N2842, N2835, N1357, N1977, N416);
or OR3 (N2843, N2817, N223, N2809);
and AND2 (N2844, N2830, N1274);
buf BUF1 (N2845, N2827);
or OR4 (N2846, N2839, N2736, N2366, N1644);
buf BUF1 (N2847, N2846);
or OR2 (N2848, N2837, N71);
xor XOR2 (N2849, N2840, N2292);
and AND4 (N2850, N2843, N2563, N838, N869);
xor XOR2 (N2851, N2850, N1104);
buf BUF1 (N2852, N2851);
or OR3 (N2853, N2841, N2631, N2477);
xor XOR2 (N2854, N2848, N1279);
and AND2 (N2855, N2849, N1220);
nand NAND4 (N2856, N2836, N1722, N2082, N2732);
nor NOR2 (N2857, N2856, N1776);
or OR3 (N2858, N2847, N1850, N930);
buf BUF1 (N2859, N2854);
not NOT1 (N2860, N2853);
nor NOR2 (N2861, N2844, N1043);
xor XOR2 (N2862, N2859, N1049);
not NOT1 (N2863, N2862);
nand NAND2 (N2864, N2845, N1377);
nor NOR4 (N2865, N2852, N1494, N1368, N2104);
buf BUF1 (N2866, N2864);
nand NAND2 (N2867, N2858, N111);
or OR2 (N2868, N2834, N2485);
and AND2 (N2869, N2855, N801);
not NOT1 (N2870, N2869);
nand NAND4 (N2871, N2857, N1277, N1538, N963);
nand NAND3 (N2872, N2866, N1819, N1037);
not NOT1 (N2873, N2842);
nand NAND4 (N2874, N2871, N2567, N1153, N1462);
nand NAND2 (N2875, N2870, N2119);
not NOT1 (N2876, N2861);
and AND4 (N2877, N2872, N1396, N1300, N272);
not NOT1 (N2878, N2865);
and AND2 (N2879, N2876, N232);
nand NAND2 (N2880, N2868, N2617);
nand NAND2 (N2881, N2860, N159);
and AND4 (N2882, N2867, N683, N1897, N1328);
not NOT1 (N2883, N2863);
or OR2 (N2884, N2883, N2302);
and AND3 (N2885, N2884, N892, N910);
nand NAND3 (N2886, N2874, N1348, N1467);
xor XOR2 (N2887, N2885, N2837);
not NOT1 (N2888, N2879);
buf BUF1 (N2889, N2875);
and AND2 (N2890, N2877, N1006);
not NOT1 (N2891, N2888);
xor XOR2 (N2892, N2881, N1396);
xor XOR2 (N2893, N2880, N769);
nand NAND3 (N2894, N2891, N2657, N1577);
or OR3 (N2895, N2892, N1756, N62);
not NOT1 (N2896, N2887);
buf BUF1 (N2897, N2873);
and AND2 (N2898, N2894, N2237);
and AND3 (N2899, N2897, N226, N266);
and AND2 (N2900, N2882, N35);
and AND2 (N2901, N2886, N2090);
nand NAND3 (N2902, N2901, N654, N2446);
or OR4 (N2903, N2899, N26, N2488, N805);
nor NOR3 (N2904, N2893, N2129, N2358);
and AND2 (N2905, N2898, N1510);
buf BUF1 (N2906, N2905);
or OR4 (N2907, N2896, N957, N88, N1790);
buf BUF1 (N2908, N2900);
not NOT1 (N2909, N2906);
or OR4 (N2910, N2878, N1980, N2090, N1594);
nor NOR4 (N2911, N2907, N2835, N992, N1937);
buf BUF1 (N2912, N2903);
and AND4 (N2913, N2889, N2765, N1698, N1549);
buf BUF1 (N2914, N2912);
nor NOR2 (N2915, N2913, N2607);
not NOT1 (N2916, N2909);
nand NAND3 (N2917, N2910, N1112, N623);
xor XOR2 (N2918, N2915, N736);
or OR3 (N2919, N2916, N400, N1110);
nor NOR2 (N2920, N2919, N1932);
and AND4 (N2921, N2917, N2787, N11, N1165);
xor XOR2 (N2922, N2920, N1889);
buf BUF1 (N2923, N2918);
not NOT1 (N2924, N2908);
or OR4 (N2925, N2895, N2244, N2668, N1812);
buf BUF1 (N2926, N2923);
or OR4 (N2927, N2924, N35, N1510, N1530);
and AND3 (N2928, N2926, N2448, N1137);
not NOT1 (N2929, N2927);
nor NOR4 (N2930, N2922, N1282, N1189, N215);
or OR2 (N2931, N2890, N1868);
xor XOR2 (N2932, N2904, N2890);
buf BUF1 (N2933, N2925);
not NOT1 (N2934, N2930);
not NOT1 (N2935, N2902);
buf BUF1 (N2936, N2921);
and AND2 (N2937, N2911, N774);
and AND3 (N2938, N2933, N2884, N123);
buf BUF1 (N2939, N2936);
nor NOR4 (N2940, N2935, N1181, N1082, N205);
and AND3 (N2941, N2937, N1125, N111);
or OR4 (N2942, N2934, N1552, N2094, N719);
xor XOR2 (N2943, N2914, N2462);
not NOT1 (N2944, N2928);
not NOT1 (N2945, N2931);
and AND4 (N2946, N2941, N2755, N605, N1022);
not NOT1 (N2947, N2945);
nor NOR3 (N2948, N2939, N1008, N940);
buf BUF1 (N2949, N2944);
buf BUF1 (N2950, N2932);
or OR4 (N2951, N2943, N2879, N960, N1085);
xor XOR2 (N2952, N2950, N462);
xor XOR2 (N2953, N2951, N1209);
nor NOR2 (N2954, N2949, N1560);
nand NAND2 (N2955, N2952, N2910);
and AND2 (N2956, N2938, N1285);
buf BUF1 (N2957, N2953);
nor NOR2 (N2958, N2954, N532);
xor XOR2 (N2959, N2948, N2952);
xor XOR2 (N2960, N2940, N1578);
not NOT1 (N2961, N2958);
not NOT1 (N2962, N2957);
or OR4 (N2963, N2947, N1085, N1112, N1699);
nand NAND2 (N2964, N2955, N1124);
and AND2 (N2965, N2961, N2632);
not NOT1 (N2966, N2946);
nor NOR3 (N2967, N2942, N555, N2596);
not NOT1 (N2968, N2960);
nor NOR2 (N2969, N2956, N91);
xor XOR2 (N2970, N2962, N737);
not NOT1 (N2971, N2959);
or OR2 (N2972, N2969, N421);
buf BUF1 (N2973, N2968);
not NOT1 (N2974, N2967);
nor NOR3 (N2975, N2963, N2250, N1784);
not NOT1 (N2976, N2929);
nand NAND4 (N2977, N2964, N2441, N455, N2884);
buf BUF1 (N2978, N2971);
buf BUF1 (N2979, N2966);
buf BUF1 (N2980, N2973);
nand NAND3 (N2981, N2977, N1728, N2691);
xor XOR2 (N2982, N2978, N2470);
buf BUF1 (N2983, N2979);
or OR4 (N2984, N2965, N2971, N2651, N2869);
and AND2 (N2985, N2982, N527);
not NOT1 (N2986, N2981);
and AND4 (N2987, N2974, N1335, N1185, N8);
nand NAND3 (N2988, N2985, N1158, N2929);
nor NOR2 (N2989, N2975, N119);
and AND2 (N2990, N2989, N1899);
nand NAND4 (N2991, N2987, N1971, N2491, N668);
nand NAND4 (N2992, N2980, N975, N2271, N2783);
not NOT1 (N2993, N2970);
nand NAND3 (N2994, N2992, N679, N324);
xor XOR2 (N2995, N2986, N2954);
not NOT1 (N2996, N2990);
or OR2 (N2997, N2976, N1865);
or OR4 (N2998, N2972, N2160, N1155, N1849);
or OR3 (N2999, N2995, N2148, N1499);
buf BUF1 (N3000, N2991);
xor XOR2 (N3001, N2996, N1969);
nand NAND2 (N3002, N3000, N128);
xor XOR2 (N3003, N2988, N2083);
or OR2 (N3004, N2984, N740);
or OR3 (N3005, N3004, N1062, N1378);
or OR2 (N3006, N2994, N2248);
xor XOR2 (N3007, N3001, N1911);
xor XOR2 (N3008, N2993, N2590);
xor XOR2 (N3009, N3006, N16);
nor NOR3 (N3010, N3008, N845, N355);
not NOT1 (N3011, N3010);
nand NAND4 (N3012, N3007, N134, N2909, N1177);
nand NAND4 (N3013, N2999, N5, N310, N919);
not NOT1 (N3014, N3013);
and AND2 (N3015, N3012, N2143);
nand NAND2 (N3016, N3011, N1156);
nor NOR2 (N3017, N2983, N2096);
nand NAND3 (N3018, N2998, N2624, N802);
and AND2 (N3019, N3017, N1640);
buf BUF1 (N3020, N3016);
nand NAND4 (N3021, N3020, N2119, N522, N2381);
buf BUF1 (N3022, N3005);
nor NOR2 (N3023, N3022, N345);
or OR2 (N3024, N3014, N174);
nor NOR3 (N3025, N3002, N575, N512);
nand NAND4 (N3026, N3019, N1339, N1767, N1912);
nor NOR3 (N3027, N2997, N306, N2806);
not NOT1 (N3028, N3015);
nand NAND2 (N3029, N3028, N1712);
xor XOR2 (N3030, N3024, N1855);
or OR2 (N3031, N3009, N1148);
xor XOR2 (N3032, N3031, N996);
xor XOR2 (N3033, N3003, N1515);
xor XOR2 (N3034, N3032, N2387);
or OR2 (N3035, N3021, N367);
and AND4 (N3036, N3027, N1018, N651, N1581);
not NOT1 (N3037, N3023);
or OR3 (N3038, N3033, N3008, N2593);
nor NOR3 (N3039, N3036, N2484, N822);
or OR3 (N3040, N3030, N1646, N2226);
buf BUF1 (N3041, N3040);
nand NAND2 (N3042, N3029, N2080);
or OR3 (N3043, N3041, N251, N450);
buf BUF1 (N3044, N3038);
xor XOR2 (N3045, N3035, N2513);
or OR2 (N3046, N3043, N55);
and AND4 (N3047, N3034, N882, N2283, N1529);
buf BUF1 (N3048, N3039);
not NOT1 (N3049, N3026);
xor XOR2 (N3050, N3048, N359);
nor NOR2 (N3051, N3045, N1298);
and AND2 (N3052, N3046, N1669);
nand NAND3 (N3053, N3018, N2765, N482);
or OR2 (N3054, N3042, N2028);
or OR3 (N3055, N3044, N2778, N377);
nand NAND4 (N3056, N3051, N152, N2411, N696);
nor NOR2 (N3057, N3053, N2011);
and AND3 (N3058, N3052, N1188, N2004);
not NOT1 (N3059, N3054);
or OR3 (N3060, N3025, N2810, N2855);
and AND4 (N3061, N3059, N530, N1037, N2726);
xor XOR2 (N3062, N3049, N2006);
or OR4 (N3063, N3058, N3018, N859, N143);
nor NOR4 (N3064, N3062, N396, N122, N472);
nand NAND2 (N3065, N3061, N2900);
or OR4 (N3066, N3064, N3017, N2323, N1281);
buf BUF1 (N3067, N3065);
nor NOR4 (N3068, N3067, N1433, N1067, N737);
nand NAND2 (N3069, N3057, N194);
nand NAND3 (N3070, N3068, N2442, N904);
nand NAND4 (N3071, N3060, N3018, N2556, N1993);
not NOT1 (N3072, N3055);
nor NOR3 (N3073, N3066, N997, N476);
not NOT1 (N3074, N3063);
nor NOR2 (N3075, N3074, N2418);
nor NOR3 (N3076, N3050, N161, N1185);
xor XOR2 (N3077, N3037, N379);
or OR4 (N3078, N3070, N3069, N1962, N439);
nor NOR3 (N3079, N561, N831, N624);
nand NAND3 (N3080, N3047, N2637, N560);
and AND2 (N3081, N3056, N2929);
and AND4 (N3082, N3076, N2735, N1438, N1499);
or OR3 (N3083, N3073, N1425, N1549);
nand NAND3 (N3084, N3082, N1560, N1556);
not NOT1 (N3085, N3075);
not NOT1 (N3086, N3084);
buf BUF1 (N3087, N3085);
nor NOR4 (N3088, N3077, N2960, N1995, N646);
or OR4 (N3089, N3071, N1620, N1366, N729);
buf BUF1 (N3090, N3087);
nor NOR2 (N3091, N3080, N990);
and AND4 (N3092, N3081, N410, N908, N2313);
not NOT1 (N3093, N3088);
buf BUF1 (N3094, N3089);
buf BUF1 (N3095, N3079);
nor NOR4 (N3096, N3091, N1456, N1828, N2933);
xor XOR2 (N3097, N3092, N1361);
nand NAND3 (N3098, N3086, N2431, N70);
buf BUF1 (N3099, N3093);
or OR4 (N3100, N3096, N882, N273, N2755);
and AND4 (N3101, N3097, N1243, N1608, N1576);
xor XOR2 (N3102, N3090, N2325);
or OR4 (N3103, N3072, N2984, N2312, N1802);
buf BUF1 (N3104, N3103);
and AND3 (N3105, N3083, N1063, N2747);
or OR4 (N3106, N3094, N2424, N305, N614);
nor NOR4 (N3107, N3078, N2688, N2576, N538);
nor NOR3 (N3108, N3105, N198, N2799);
nand NAND4 (N3109, N3102, N1340, N1813, N66);
or OR3 (N3110, N3098, N1332, N1614);
xor XOR2 (N3111, N3106, N614);
nand NAND2 (N3112, N3110, N1211);
not NOT1 (N3113, N3104);
nand NAND4 (N3114, N3107, N598, N203, N1232);
nor NOR4 (N3115, N3095, N595, N2344, N2465);
and AND4 (N3116, N3100, N1040, N83, N1530);
buf BUF1 (N3117, N3111);
xor XOR2 (N3118, N3113, N542);
not NOT1 (N3119, N3112);
xor XOR2 (N3120, N3117, N613);
or OR2 (N3121, N3114, N1139);
xor XOR2 (N3122, N3120, N875);
nor NOR3 (N3123, N3108, N736, N1989);
nor NOR2 (N3124, N3123, N1407);
nand NAND3 (N3125, N3101, N2876, N539);
or OR4 (N3126, N3099, N2847, N536, N1086);
not NOT1 (N3127, N3121);
buf BUF1 (N3128, N3119);
not NOT1 (N3129, N3116);
or OR3 (N3130, N3125, N331, N1019);
not NOT1 (N3131, N3109);
buf BUF1 (N3132, N3128);
or OR4 (N3133, N3124, N2432, N2796, N2596);
nand NAND4 (N3134, N3122, N2747, N2201, N2858);
xor XOR2 (N3135, N3127, N1027);
and AND4 (N3136, N3129, N1409, N2476, N823);
nor NOR4 (N3137, N3118, N2846, N2789, N1977);
buf BUF1 (N3138, N3133);
xor XOR2 (N3139, N3134, N718);
not NOT1 (N3140, N3139);
buf BUF1 (N3141, N3132);
not NOT1 (N3142, N3126);
xor XOR2 (N3143, N3142, N1124);
nand NAND3 (N3144, N3137, N443, N273);
and AND2 (N3145, N3141, N743);
nand NAND3 (N3146, N3115, N2518, N1107);
or OR4 (N3147, N3138, N3075, N1531, N2046);
and AND2 (N3148, N3144, N1913);
nand NAND3 (N3149, N3135, N1772, N604);
or OR4 (N3150, N3130, N3021, N1958, N1938);
and AND3 (N3151, N3136, N574, N274);
buf BUF1 (N3152, N3148);
xor XOR2 (N3153, N3145, N970);
nand NAND2 (N3154, N3153, N2942);
nand NAND4 (N3155, N3152, N436, N510, N452);
xor XOR2 (N3156, N3154, N2347);
nor NOR3 (N3157, N3150, N2938, N2624);
xor XOR2 (N3158, N3140, N1807);
xor XOR2 (N3159, N3151, N1244);
nor NOR2 (N3160, N3159, N1461);
not NOT1 (N3161, N3149);
buf BUF1 (N3162, N3131);
xor XOR2 (N3163, N3160, N91);
or OR3 (N3164, N3161, N2821, N1126);
or OR4 (N3165, N3146, N2149, N1155, N1344);
or OR2 (N3166, N3147, N530);
xor XOR2 (N3167, N3143, N1240);
not NOT1 (N3168, N3156);
not NOT1 (N3169, N3162);
and AND3 (N3170, N3164, N3091, N122);
xor XOR2 (N3171, N3170, N1998);
nand NAND4 (N3172, N3163, N691, N1560, N745);
and AND2 (N3173, N3165, N1315);
and AND2 (N3174, N3167, N1373);
or OR2 (N3175, N3157, N2677);
xor XOR2 (N3176, N3158, N2058);
buf BUF1 (N3177, N3175);
nand NAND3 (N3178, N3168, N851, N559);
not NOT1 (N3179, N3173);
nor NOR2 (N3180, N3172, N2408);
xor XOR2 (N3181, N3177, N489);
nor NOR2 (N3182, N3176, N2063);
buf BUF1 (N3183, N3155);
buf BUF1 (N3184, N3169);
not NOT1 (N3185, N3166);
xor XOR2 (N3186, N3174, N2036);
buf BUF1 (N3187, N3185);
xor XOR2 (N3188, N3186, N2130);
xor XOR2 (N3189, N3187, N1730);
nor NOR3 (N3190, N3179, N1110, N2049);
nand NAND4 (N3191, N3181, N2928, N1571, N1211);
not NOT1 (N3192, N3184);
nor NOR4 (N3193, N3171, N1638, N1459, N1091);
and AND2 (N3194, N3188, N147);
xor XOR2 (N3195, N3182, N2052);
nor NOR3 (N3196, N3183, N1767, N480);
not NOT1 (N3197, N3180);
xor XOR2 (N3198, N3189, N2578);
and AND3 (N3199, N3196, N3015, N1581);
xor XOR2 (N3200, N3191, N2769);
nand NAND4 (N3201, N3198, N785, N2985, N2798);
and AND4 (N3202, N3192, N780, N1347, N2215);
nor NOR3 (N3203, N3201, N501, N1882);
xor XOR2 (N3204, N3199, N1414);
nor NOR3 (N3205, N3204, N2702, N2991);
or OR3 (N3206, N3195, N1096, N2440);
nand NAND3 (N3207, N3203, N1848, N2476);
not NOT1 (N3208, N3194);
or OR3 (N3209, N3190, N1466, N1336);
not NOT1 (N3210, N3209);
not NOT1 (N3211, N3202);
not NOT1 (N3212, N3197);
buf BUF1 (N3213, N3211);
xor XOR2 (N3214, N3193, N207);
nor NOR3 (N3215, N3210, N1687, N1041);
nor NOR4 (N3216, N3206, N1057, N662, N3036);
or OR3 (N3217, N3212, N1509, N512);
buf BUF1 (N3218, N3178);
buf BUF1 (N3219, N3200);
not NOT1 (N3220, N3217);
or OR4 (N3221, N3207, N93, N2308, N1360);
not NOT1 (N3222, N3214);
endmodule