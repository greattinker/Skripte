// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14;

output N3010,N3011,N3002,N2990,N3013,N2981,N2997,N2987,N3012,N3014;

not NOT1 (N15, N14);
or OR3 (N16, N4, N1, N5);
nor NOR4 (N17, N1, N12, N12, N8);
buf BUF1 (N18, N10);
not NOT1 (N19, N17);
nor NOR2 (N20, N7, N14);
not NOT1 (N21, N9);
buf BUF1 (N22, N14);
buf BUF1 (N23, N15);
not NOT1 (N24, N22);
and AND2 (N25, N10, N13);
nand NAND3 (N26, N8, N10, N1);
xor XOR2 (N27, N1, N9);
or OR4 (N28, N19, N22, N26, N18);
not NOT1 (N29, N15);
xor XOR2 (N30, N24, N26);
not NOT1 (N31, N7);
xor XOR2 (N32, N29, N28);
not NOT1 (N33, N11);
buf BUF1 (N34, N33);
nand NAND4 (N35, N31, N25, N24, N3);
xor XOR2 (N36, N25, N13);
and AND4 (N37, N20, N14, N12, N22);
not NOT1 (N38, N16);
xor XOR2 (N39, N27, N23);
or OR3 (N40, N31, N2, N7);
not NOT1 (N41, N21);
nand NAND2 (N42, N39, N39);
and AND4 (N43, N36, N11, N10, N19);
nor NOR3 (N44, N30, N41, N43);
or OR3 (N45, N8, N39, N18);
or OR4 (N46, N17, N6, N41, N31);
nand NAND4 (N47, N45, N1, N4, N30);
buf BUF1 (N48, N37);
or OR4 (N49, N40, N31, N6, N11);
nand NAND4 (N50, N46, N3, N44, N46);
nand NAND2 (N51, N16, N21);
or OR2 (N52, N51, N1);
buf BUF1 (N53, N52);
nor NOR2 (N54, N53, N15);
buf BUF1 (N55, N47);
xor XOR2 (N56, N48, N35);
nor NOR4 (N57, N29, N40, N44, N30);
buf BUF1 (N58, N55);
or OR3 (N59, N38, N52, N36);
and AND3 (N60, N57, N59, N14);
not NOT1 (N61, N42);
and AND3 (N62, N20, N53, N59);
and AND4 (N63, N58, N51, N24, N31);
and AND3 (N64, N49, N28, N1);
or OR3 (N65, N32, N55, N23);
buf BUF1 (N66, N60);
buf BUF1 (N67, N56);
and AND2 (N68, N65, N62);
not NOT1 (N69, N68);
buf BUF1 (N70, N48);
buf BUF1 (N71, N61);
nand NAND4 (N72, N71, N1, N38, N57);
nor NOR3 (N73, N69, N36, N31);
or OR3 (N74, N66, N58, N69);
nor NOR2 (N75, N34, N3);
or OR4 (N76, N54, N44, N71, N59);
not NOT1 (N77, N74);
nand NAND2 (N78, N64, N28);
or OR4 (N79, N63, N63, N58, N54);
nor NOR2 (N80, N73, N13);
nor NOR3 (N81, N76, N10, N74);
buf BUF1 (N82, N75);
not NOT1 (N83, N82);
and AND4 (N84, N79, N22, N63, N74);
not NOT1 (N85, N80);
nor NOR2 (N86, N72, N58);
or OR2 (N87, N83, N20);
not NOT1 (N88, N81);
nor NOR3 (N89, N86, N51, N14);
or OR2 (N90, N78, N65);
nor NOR3 (N91, N90, N89, N20);
or OR2 (N92, N90, N49);
and AND4 (N93, N85, N66, N51, N30);
or OR4 (N94, N88, N7, N55, N13);
nand NAND4 (N95, N77, N91, N7, N61);
and AND4 (N96, N8, N46, N51, N60);
xor XOR2 (N97, N96, N14);
not NOT1 (N98, N67);
or OR3 (N99, N94, N87, N18);
buf BUF1 (N100, N46);
nor NOR3 (N101, N50, N91, N44);
buf BUF1 (N102, N84);
buf BUF1 (N103, N100);
nand NAND2 (N104, N93, N76);
xor XOR2 (N105, N92, N51);
or OR2 (N106, N98, N51);
buf BUF1 (N107, N97);
xor XOR2 (N108, N106, N9);
and AND4 (N109, N99, N81, N27, N36);
buf BUF1 (N110, N104);
not NOT1 (N111, N101);
and AND2 (N112, N105, N76);
xor XOR2 (N113, N95, N3);
not NOT1 (N114, N111);
xor XOR2 (N115, N113, N93);
nand NAND4 (N116, N108, N41, N52, N69);
xor XOR2 (N117, N116, N45);
or OR3 (N118, N70, N116, N72);
not NOT1 (N119, N110);
and AND2 (N120, N117, N79);
and AND3 (N121, N120, N11, N39);
not NOT1 (N122, N114);
or OR3 (N123, N115, N87, N21);
xor XOR2 (N124, N122, N118);
nor NOR4 (N125, N32, N54, N52, N65);
nor NOR4 (N126, N112, N93, N83, N1);
or OR4 (N127, N123, N38, N71, N27);
xor XOR2 (N128, N102, N70);
not NOT1 (N129, N119);
not NOT1 (N130, N107);
buf BUF1 (N131, N124);
buf BUF1 (N132, N129);
or OR2 (N133, N132, N43);
or OR2 (N134, N121, N7);
and AND3 (N135, N109, N113, N79);
and AND3 (N136, N130, N84, N126);
buf BUF1 (N137, N99);
not NOT1 (N138, N103);
nor NOR4 (N139, N137, N28, N105, N14);
buf BUF1 (N140, N135);
nor NOR3 (N141, N134, N47, N64);
or OR2 (N142, N131, N50);
nand NAND4 (N143, N127, N65, N13, N96);
xor XOR2 (N144, N139, N9);
xor XOR2 (N145, N140, N104);
xor XOR2 (N146, N128, N88);
buf BUF1 (N147, N133);
nor NOR4 (N148, N141, N135, N104, N105);
or OR4 (N149, N148, N63, N58, N64);
or OR3 (N150, N125, N44, N70);
buf BUF1 (N151, N145);
nor NOR2 (N152, N150, N82);
xor XOR2 (N153, N152, N54);
xor XOR2 (N154, N146, N142);
xor XOR2 (N155, N39, N128);
buf BUF1 (N156, N153);
nand NAND3 (N157, N144, N150, N39);
not NOT1 (N158, N157);
nand NAND4 (N159, N151, N134, N83, N14);
or OR2 (N160, N156, N22);
xor XOR2 (N161, N149, N7);
not NOT1 (N162, N136);
xor XOR2 (N163, N162, N29);
nor NOR4 (N164, N161, N121, N106, N147);
not NOT1 (N165, N109);
or OR3 (N166, N160, N100, N108);
nand NAND3 (N167, N138, N148, N137);
or OR4 (N168, N167, N18, N124, N105);
or OR4 (N169, N163, N61, N155, N80);
xor XOR2 (N170, N136, N94);
or OR2 (N171, N158, N89);
not NOT1 (N172, N165);
or OR4 (N173, N143, N42, N78, N68);
not NOT1 (N174, N159);
not NOT1 (N175, N166);
and AND2 (N176, N168, N52);
buf BUF1 (N177, N175);
nor NOR3 (N178, N176, N41, N51);
buf BUF1 (N179, N164);
and AND2 (N180, N171, N16);
nand NAND3 (N181, N179, N45, N140);
not NOT1 (N182, N177);
nand NAND3 (N183, N180, N10, N54);
and AND2 (N184, N173, N16);
nor NOR4 (N185, N169, N99, N157, N106);
xor XOR2 (N186, N183, N26);
and AND3 (N187, N170, N131, N24);
and AND3 (N188, N181, N161, N111);
nor NOR4 (N189, N184, N51, N15, N120);
buf BUF1 (N190, N185);
not NOT1 (N191, N188);
or OR3 (N192, N189, N177, N130);
buf BUF1 (N193, N186);
nor NOR3 (N194, N172, N133, N41);
not NOT1 (N195, N190);
buf BUF1 (N196, N154);
nor NOR2 (N197, N196, N76);
nand NAND4 (N198, N182, N131, N33, N155);
xor XOR2 (N199, N198, N197);
not NOT1 (N200, N188);
nand NAND3 (N201, N199, N10, N60);
not NOT1 (N202, N191);
and AND4 (N203, N178, N37, N19, N192);
and AND2 (N204, N177, N162);
not NOT1 (N205, N203);
nand NAND2 (N206, N204, N30);
not NOT1 (N207, N206);
buf BUF1 (N208, N202);
or OR4 (N209, N208, N143, N8, N174);
and AND2 (N210, N169, N114);
xor XOR2 (N211, N210, N114);
and AND3 (N212, N200, N183, N23);
nor NOR4 (N213, N193, N196, N1, N14);
or OR4 (N214, N195, N13, N120, N148);
and AND2 (N215, N211, N89);
buf BUF1 (N216, N205);
nor NOR4 (N217, N207, N212, N68, N94);
nand NAND2 (N218, N202, N9);
nand NAND4 (N219, N194, N108, N79, N160);
or OR2 (N220, N218, N147);
xor XOR2 (N221, N215, N22);
nand NAND2 (N222, N216, N11);
and AND4 (N223, N220, N151, N49, N154);
xor XOR2 (N224, N221, N124);
nor NOR3 (N225, N201, N64, N192);
nand NAND3 (N226, N217, N81, N118);
or OR2 (N227, N222, N116);
buf BUF1 (N228, N187);
and AND2 (N229, N209, N106);
or OR2 (N230, N224, N35);
not NOT1 (N231, N228);
or OR4 (N232, N231, N196, N126, N106);
or OR3 (N233, N223, N154, N128);
xor XOR2 (N234, N230, N143);
or OR2 (N235, N229, N94);
buf BUF1 (N236, N232);
and AND2 (N237, N227, N171);
or OR4 (N238, N235, N227, N141, N77);
and AND4 (N239, N225, N39, N13, N222);
not NOT1 (N240, N237);
nand NAND3 (N241, N213, N70, N230);
or OR4 (N242, N219, N51, N151, N90);
xor XOR2 (N243, N241, N175);
not NOT1 (N244, N233);
xor XOR2 (N245, N236, N4);
xor XOR2 (N246, N214, N136);
xor XOR2 (N247, N234, N52);
xor XOR2 (N248, N244, N151);
buf BUF1 (N249, N243);
xor XOR2 (N250, N242, N209);
nand NAND3 (N251, N246, N187, N162);
and AND4 (N252, N248, N51, N167, N89);
nand NAND3 (N253, N245, N95, N244);
nand NAND2 (N254, N252, N134);
nor NOR4 (N255, N253, N66, N102, N88);
and AND4 (N256, N250, N61, N141, N138);
and AND3 (N257, N240, N28, N163);
and AND3 (N258, N257, N9, N2);
nand NAND2 (N259, N256, N45);
and AND2 (N260, N238, N253);
xor XOR2 (N261, N239, N17);
not NOT1 (N262, N261);
nand NAND3 (N263, N249, N237, N108);
not NOT1 (N264, N262);
and AND3 (N265, N263, N23, N157);
nand NAND4 (N266, N259, N117, N126, N186);
nand NAND2 (N267, N260, N134);
buf BUF1 (N268, N265);
nor NOR2 (N269, N267, N121);
or OR2 (N270, N264, N186);
not NOT1 (N271, N255);
nand NAND4 (N272, N269, N204, N1, N204);
nor NOR4 (N273, N268, N139, N12, N181);
buf BUF1 (N274, N251);
and AND2 (N275, N258, N123);
buf BUF1 (N276, N247);
xor XOR2 (N277, N276, N257);
buf BUF1 (N278, N275);
and AND3 (N279, N273, N68, N108);
nand NAND4 (N280, N278, N128, N163, N160);
or OR2 (N281, N277, N28);
or OR3 (N282, N281, N92, N186);
and AND2 (N283, N271, N231);
buf BUF1 (N284, N254);
or OR2 (N285, N270, N140);
buf BUF1 (N286, N226);
or OR2 (N287, N274, N159);
not NOT1 (N288, N279);
not NOT1 (N289, N283);
buf BUF1 (N290, N284);
nor NOR3 (N291, N289, N17, N159);
nand NAND4 (N292, N280, N143, N44, N160);
buf BUF1 (N293, N288);
xor XOR2 (N294, N286, N2);
and AND3 (N295, N292, N235, N222);
nand NAND2 (N296, N285, N51);
not NOT1 (N297, N287);
nor NOR3 (N298, N294, N271, N105);
not NOT1 (N299, N295);
buf BUF1 (N300, N266);
or OR2 (N301, N293, N252);
xor XOR2 (N302, N301, N258);
buf BUF1 (N303, N291);
buf BUF1 (N304, N272);
or OR3 (N305, N296, N228, N124);
xor XOR2 (N306, N302, N68);
and AND3 (N307, N290, N301, N148);
not NOT1 (N308, N297);
or OR2 (N309, N300, N25);
and AND3 (N310, N298, N210, N95);
and AND3 (N311, N282, N104, N219);
buf BUF1 (N312, N306);
buf BUF1 (N313, N299);
or OR2 (N314, N312, N121);
xor XOR2 (N315, N314, N184);
nor NOR3 (N316, N308, N302, N217);
xor XOR2 (N317, N309, N102);
or OR3 (N318, N317, N78, N67);
buf BUF1 (N319, N315);
nand NAND2 (N320, N313, N293);
not NOT1 (N321, N318);
xor XOR2 (N322, N316, N66);
nor NOR3 (N323, N305, N13, N311);
or OR3 (N324, N256, N102, N192);
or OR3 (N325, N322, N116, N199);
nand NAND4 (N326, N323, N203, N153, N115);
and AND3 (N327, N326, N234, N170);
and AND2 (N328, N327, N259);
and AND4 (N329, N320, N192, N192, N161);
buf BUF1 (N330, N307);
nor NOR2 (N331, N310, N132);
nor NOR4 (N332, N330, N86, N228, N299);
or OR3 (N333, N324, N58, N284);
buf BUF1 (N334, N331);
or OR4 (N335, N334, N80, N17, N148);
buf BUF1 (N336, N303);
and AND2 (N337, N335, N99);
nor NOR3 (N338, N329, N180, N74);
not NOT1 (N339, N325);
or OR4 (N340, N332, N263, N103, N300);
nor NOR3 (N341, N321, N268, N85);
buf BUF1 (N342, N339);
nand NAND4 (N343, N337, N152, N22, N232);
not NOT1 (N344, N336);
and AND4 (N345, N343, N177, N19, N215);
xor XOR2 (N346, N333, N3);
or OR3 (N347, N341, N56, N43);
xor XOR2 (N348, N346, N262);
buf BUF1 (N349, N319);
nor NOR3 (N350, N348, N63, N50);
and AND3 (N351, N344, N334, N134);
nand NAND2 (N352, N328, N212);
xor XOR2 (N353, N351, N75);
xor XOR2 (N354, N350, N127);
nand NAND4 (N355, N352, N106, N51, N210);
buf BUF1 (N356, N347);
nand NAND3 (N357, N356, N136, N116);
and AND2 (N358, N353, N45);
not NOT1 (N359, N345);
buf BUF1 (N360, N304);
and AND4 (N361, N354, N212, N7, N27);
and AND2 (N362, N340, N180);
buf BUF1 (N363, N342);
nand NAND2 (N364, N358, N361);
xor XOR2 (N365, N285, N104);
nand NAND3 (N366, N362, N238, N345);
xor XOR2 (N367, N363, N32);
nor NOR4 (N368, N365, N307, N181, N239);
nand NAND3 (N369, N360, N223, N131);
not NOT1 (N370, N366);
buf BUF1 (N371, N369);
xor XOR2 (N372, N368, N246);
and AND4 (N373, N364, N119, N27, N217);
or OR3 (N374, N371, N187, N236);
not NOT1 (N375, N355);
xor XOR2 (N376, N349, N131);
nor NOR2 (N377, N367, N223);
or OR4 (N378, N374, N209, N129, N260);
not NOT1 (N379, N377);
nand NAND4 (N380, N378, N109, N327, N232);
or OR3 (N381, N359, N197, N326);
xor XOR2 (N382, N379, N339);
xor XOR2 (N383, N375, N252);
not NOT1 (N384, N381);
buf BUF1 (N385, N384);
or OR4 (N386, N372, N127, N274, N271);
nor NOR3 (N387, N370, N280, N355);
nor NOR4 (N388, N383, N338, N353, N317);
nand NAND3 (N389, N12, N135, N183);
nor NOR3 (N390, N380, N233, N238);
nand NAND2 (N391, N385, N33);
not NOT1 (N392, N373);
nand NAND3 (N393, N382, N141, N103);
xor XOR2 (N394, N392, N255);
nor NOR4 (N395, N388, N26, N21, N225);
or OR4 (N396, N357, N222, N129, N45);
buf BUF1 (N397, N393);
buf BUF1 (N398, N386);
xor XOR2 (N399, N376, N136);
nor NOR3 (N400, N397, N390, N99);
buf BUF1 (N401, N383);
and AND2 (N402, N396, N187);
not NOT1 (N403, N389);
xor XOR2 (N404, N387, N72);
buf BUF1 (N405, N399);
nand NAND4 (N406, N400, N258, N242, N138);
nand NAND3 (N407, N401, N159, N309);
xor XOR2 (N408, N403, N395);
nand NAND3 (N409, N91, N257, N74);
nand NAND3 (N410, N405, N394, N406);
or OR2 (N411, N9, N324);
not NOT1 (N412, N162);
and AND4 (N413, N410, N189, N52, N251);
buf BUF1 (N414, N412);
buf BUF1 (N415, N398);
nor NOR4 (N416, N415, N312, N349, N1);
buf BUF1 (N417, N408);
nor NOR2 (N418, N402, N329);
nor NOR3 (N419, N391, N101, N358);
nand NAND4 (N420, N417, N312, N5, N307);
nand NAND3 (N421, N409, N290, N201);
or OR4 (N422, N414, N64, N37, N132);
nor NOR3 (N423, N419, N301, N326);
nor NOR2 (N424, N421, N157);
and AND3 (N425, N413, N421, N90);
buf BUF1 (N426, N404);
buf BUF1 (N427, N420);
nor NOR3 (N428, N422, N427, N353);
not NOT1 (N429, N86);
nand NAND3 (N430, N428, N79, N421);
and AND3 (N431, N423, N323, N115);
nand NAND4 (N432, N411, N100, N145, N14);
nor NOR2 (N433, N426, N385);
or OR2 (N434, N418, N386);
buf BUF1 (N435, N434);
not NOT1 (N436, N429);
buf BUF1 (N437, N416);
nand NAND4 (N438, N435, N18, N280, N358);
and AND4 (N439, N438, N7, N216, N136);
not NOT1 (N440, N430);
xor XOR2 (N441, N425, N357);
nor NOR3 (N442, N433, N161, N56);
xor XOR2 (N443, N432, N284);
not NOT1 (N444, N442);
and AND2 (N445, N441, N391);
not NOT1 (N446, N407);
not NOT1 (N447, N446);
and AND2 (N448, N436, N274);
not NOT1 (N449, N445);
and AND3 (N450, N443, N152, N245);
buf BUF1 (N451, N431);
buf BUF1 (N452, N449);
nor NOR4 (N453, N437, N21, N320, N211);
and AND3 (N454, N452, N135, N30);
not NOT1 (N455, N453);
nand NAND2 (N456, N454, N351);
xor XOR2 (N457, N444, N169);
not NOT1 (N458, N439);
buf BUF1 (N459, N456);
nand NAND2 (N460, N440, N234);
buf BUF1 (N461, N451);
nor NOR3 (N462, N461, N8, N399);
xor XOR2 (N463, N450, N31);
xor XOR2 (N464, N460, N210);
xor XOR2 (N465, N458, N446);
nand NAND3 (N466, N465, N207, N445);
and AND4 (N467, N455, N305, N451, N208);
not NOT1 (N468, N457);
and AND2 (N469, N463, N90);
not NOT1 (N470, N462);
or OR4 (N471, N467, N175, N41, N315);
nand NAND2 (N472, N469, N133);
not NOT1 (N473, N472);
buf BUF1 (N474, N466);
nand NAND4 (N475, N474, N471, N367, N59);
or OR2 (N476, N204, N364);
and AND4 (N477, N468, N411, N32, N350);
and AND4 (N478, N459, N8, N430, N362);
buf BUF1 (N479, N448);
buf BUF1 (N480, N479);
xor XOR2 (N481, N477, N107);
or OR3 (N482, N476, N50, N458);
buf BUF1 (N483, N464);
or OR3 (N484, N424, N218, N467);
not NOT1 (N485, N483);
xor XOR2 (N486, N473, N240);
not NOT1 (N487, N480);
not NOT1 (N488, N485);
and AND4 (N489, N470, N65, N376, N231);
or OR3 (N490, N489, N61, N88);
and AND4 (N491, N488, N129, N373, N382);
not NOT1 (N492, N487);
xor XOR2 (N493, N491, N230);
buf BUF1 (N494, N484);
xor XOR2 (N495, N490, N51);
buf BUF1 (N496, N475);
xor XOR2 (N497, N447, N486);
not NOT1 (N498, N496);
buf BUF1 (N499, N105);
buf BUF1 (N500, N492);
or OR2 (N501, N500, N286);
nor NOR3 (N502, N493, N195, N63);
nand NAND4 (N503, N495, N286, N481, N44);
buf BUF1 (N504, N400);
or OR2 (N505, N478, N330);
and AND3 (N506, N501, N221, N439);
or OR3 (N507, N506, N478, N33);
buf BUF1 (N508, N482);
xor XOR2 (N509, N504, N261);
or OR4 (N510, N503, N282, N392, N449);
xor XOR2 (N511, N508, N53);
buf BUF1 (N512, N507);
nor NOR2 (N513, N510, N31);
buf BUF1 (N514, N494);
and AND3 (N515, N509, N23, N127);
not NOT1 (N516, N499);
and AND3 (N517, N514, N147, N396);
buf BUF1 (N518, N505);
or OR4 (N519, N516, N354, N63, N499);
or OR2 (N520, N513, N497);
not NOT1 (N521, N367);
not NOT1 (N522, N521);
not NOT1 (N523, N519);
and AND4 (N524, N515, N274, N499, N158);
nor NOR2 (N525, N498, N366);
buf BUF1 (N526, N518);
not NOT1 (N527, N524);
xor XOR2 (N528, N520, N228);
nor NOR3 (N529, N525, N523, N303);
and AND4 (N530, N330, N63, N53, N504);
or OR3 (N531, N522, N295, N402);
and AND2 (N532, N517, N478);
or OR3 (N533, N512, N523, N179);
and AND3 (N534, N529, N206, N164);
or OR3 (N535, N532, N492, N326);
nor NOR3 (N536, N534, N362, N427);
buf BUF1 (N537, N531);
not NOT1 (N538, N537);
or OR2 (N539, N536, N83);
nor NOR2 (N540, N538, N249);
nor NOR4 (N541, N533, N91, N17, N5);
or OR4 (N542, N502, N113, N403, N4);
or OR2 (N543, N527, N422);
or OR2 (N544, N541, N494);
and AND4 (N545, N539, N9, N358, N398);
xor XOR2 (N546, N544, N235);
and AND3 (N547, N540, N442, N31);
xor XOR2 (N548, N511, N544);
xor XOR2 (N549, N546, N92);
nand NAND2 (N550, N530, N286);
not NOT1 (N551, N547);
or OR2 (N552, N528, N97);
nor NOR4 (N553, N551, N66, N333, N14);
xor XOR2 (N554, N543, N338);
nand NAND2 (N555, N549, N430);
buf BUF1 (N556, N552);
or OR4 (N557, N526, N459, N160, N404);
and AND3 (N558, N550, N167, N420);
buf BUF1 (N559, N553);
nand NAND3 (N560, N548, N143, N51);
and AND3 (N561, N555, N210, N324);
nand NAND4 (N562, N561, N496, N480, N170);
xor XOR2 (N563, N554, N290);
buf BUF1 (N564, N559);
or OR2 (N565, N557, N268);
and AND4 (N566, N535, N19, N470, N541);
buf BUF1 (N567, N564);
or OR2 (N568, N560, N68);
nor NOR3 (N569, N542, N128, N518);
not NOT1 (N570, N568);
buf BUF1 (N571, N565);
xor XOR2 (N572, N566, N239);
or OR3 (N573, N572, N477, N413);
and AND3 (N574, N569, N207, N139);
nand NAND2 (N575, N545, N145);
buf BUF1 (N576, N556);
buf BUF1 (N577, N576);
buf BUF1 (N578, N567);
nand NAND2 (N579, N578, N140);
not NOT1 (N580, N562);
or OR4 (N581, N577, N61, N258, N532);
and AND4 (N582, N573, N346, N99, N534);
and AND2 (N583, N571, N487);
nand NAND3 (N584, N583, N474, N126);
buf BUF1 (N585, N563);
buf BUF1 (N586, N582);
not NOT1 (N587, N581);
or OR4 (N588, N586, N400, N547, N109);
xor XOR2 (N589, N587, N377);
nand NAND2 (N590, N574, N261);
nor NOR4 (N591, N558, N208, N8, N502);
xor XOR2 (N592, N575, N112);
nor NOR4 (N593, N590, N21, N39, N525);
buf BUF1 (N594, N570);
xor XOR2 (N595, N579, N169);
xor XOR2 (N596, N588, N78);
nor NOR2 (N597, N595, N34);
nor NOR3 (N598, N597, N180, N208);
and AND3 (N599, N585, N290, N529);
nand NAND2 (N600, N598, N575);
and AND3 (N601, N580, N404, N242);
or OR2 (N602, N589, N538);
buf BUF1 (N603, N602);
nand NAND3 (N604, N596, N579, N52);
nor NOR4 (N605, N600, N516, N300, N210);
xor XOR2 (N606, N594, N381);
and AND3 (N607, N584, N341, N104);
xor XOR2 (N608, N606, N188);
nor NOR3 (N609, N605, N51, N118);
buf BUF1 (N610, N603);
nand NAND2 (N611, N607, N591);
and AND4 (N612, N65, N452, N14, N168);
buf BUF1 (N613, N592);
not NOT1 (N614, N609);
or OR2 (N615, N614, N227);
xor XOR2 (N616, N615, N162);
nand NAND3 (N617, N601, N461, N473);
or OR2 (N618, N599, N55);
nand NAND4 (N619, N611, N71, N87, N202);
nand NAND3 (N620, N612, N259, N340);
or OR2 (N621, N608, N335);
xor XOR2 (N622, N593, N608);
nand NAND3 (N623, N604, N457, N74);
buf BUF1 (N624, N621);
xor XOR2 (N625, N617, N61);
not NOT1 (N626, N610);
and AND2 (N627, N622, N518);
or OR2 (N628, N623, N468);
nor NOR2 (N629, N616, N512);
and AND4 (N630, N624, N357, N317, N32);
or OR3 (N631, N628, N270, N44);
and AND3 (N632, N626, N333, N484);
nand NAND2 (N633, N630, N108);
xor XOR2 (N634, N625, N417);
nand NAND3 (N635, N627, N402, N468);
or OR4 (N636, N618, N536, N26, N622);
nor NOR3 (N637, N629, N79, N305);
or OR2 (N638, N633, N547);
nor NOR2 (N639, N637, N91);
nor NOR2 (N640, N638, N363);
nor NOR2 (N641, N635, N550);
nor NOR2 (N642, N620, N276);
xor XOR2 (N643, N631, N59);
nor NOR2 (N644, N642, N303);
nand NAND3 (N645, N632, N23, N178);
nand NAND4 (N646, N639, N188, N136, N562);
xor XOR2 (N647, N640, N319);
xor XOR2 (N648, N645, N364);
nor NOR3 (N649, N647, N363, N178);
and AND4 (N650, N636, N293, N471, N274);
nor NOR4 (N651, N648, N633, N121, N581);
nand NAND2 (N652, N619, N641);
not NOT1 (N653, N556);
nor NOR2 (N654, N644, N222);
nor NOR2 (N655, N643, N632);
nand NAND2 (N656, N652, N470);
and AND2 (N657, N656, N598);
nor NOR4 (N658, N634, N109, N567, N432);
buf BUF1 (N659, N653);
not NOT1 (N660, N655);
nand NAND2 (N661, N649, N443);
nand NAND3 (N662, N651, N363, N86);
or OR2 (N663, N646, N6);
or OR2 (N664, N654, N599);
nand NAND3 (N665, N658, N638, N510);
nor NOR4 (N666, N662, N301, N357, N266);
not NOT1 (N667, N666);
nor NOR2 (N668, N660, N77);
and AND3 (N669, N667, N213, N572);
nor NOR4 (N670, N659, N261, N218, N4);
not NOT1 (N671, N670);
buf BUF1 (N672, N663);
or OR2 (N673, N661, N619);
nor NOR2 (N674, N671, N402);
and AND2 (N675, N613, N91);
and AND3 (N676, N657, N669, N433);
xor XOR2 (N677, N164, N520);
and AND4 (N678, N673, N309, N6, N381);
xor XOR2 (N679, N665, N437);
and AND4 (N680, N650, N590, N235, N245);
or OR2 (N681, N679, N405);
nor NOR3 (N682, N678, N26, N653);
buf BUF1 (N683, N680);
and AND3 (N684, N664, N119, N40);
nor NOR4 (N685, N672, N630, N122, N680);
and AND4 (N686, N674, N367, N258, N161);
nand NAND2 (N687, N668, N162);
and AND3 (N688, N682, N574, N115);
buf BUF1 (N689, N683);
nand NAND4 (N690, N689, N373, N410, N289);
not NOT1 (N691, N690);
not NOT1 (N692, N681);
nand NAND3 (N693, N675, N377, N420);
nor NOR3 (N694, N684, N456, N567);
nand NAND3 (N695, N691, N51, N279);
nor NOR4 (N696, N692, N516, N556, N672);
and AND4 (N697, N693, N519, N273, N24);
buf BUF1 (N698, N694);
nand NAND2 (N699, N695, N389);
nand NAND4 (N700, N698, N232, N491, N682);
not NOT1 (N701, N676);
or OR3 (N702, N688, N495, N398);
nor NOR3 (N703, N700, N457, N163);
and AND4 (N704, N677, N536, N241, N375);
xor XOR2 (N705, N697, N288);
and AND2 (N706, N703, N423);
nand NAND3 (N707, N699, N185, N260);
not NOT1 (N708, N686);
or OR4 (N709, N701, N266, N254, N183);
or OR2 (N710, N706, N58);
not NOT1 (N711, N705);
nand NAND3 (N712, N687, N108, N546);
xor XOR2 (N713, N712, N238);
and AND3 (N714, N702, N532, N576);
nand NAND2 (N715, N713, N229);
or OR2 (N716, N715, N351);
and AND4 (N717, N711, N224, N56, N606);
not NOT1 (N718, N716);
xor XOR2 (N719, N710, N544);
buf BUF1 (N720, N708);
or OR4 (N721, N704, N15, N330, N447);
or OR4 (N722, N721, N621, N184, N629);
nor NOR3 (N723, N696, N669, N402);
xor XOR2 (N724, N722, N370);
nand NAND4 (N725, N707, N681, N124, N83);
or OR2 (N726, N719, N509);
and AND4 (N727, N717, N717, N554, N31);
buf BUF1 (N728, N724);
xor XOR2 (N729, N720, N306);
buf BUF1 (N730, N723);
or OR2 (N731, N709, N379);
nor NOR2 (N732, N725, N643);
nand NAND2 (N733, N727, N731);
xor XOR2 (N734, N567, N677);
nand NAND3 (N735, N730, N212, N133);
or OR2 (N736, N718, N22);
and AND2 (N737, N726, N131);
or OR3 (N738, N728, N670, N356);
and AND3 (N739, N732, N631, N447);
buf BUF1 (N740, N736);
or OR4 (N741, N740, N40, N232, N471);
nor NOR2 (N742, N741, N554);
not NOT1 (N743, N737);
buf BUF1 (N744, N739);
nand NAND4 (N745, N743, N250, N470, N715);
and AND4 (N746, N733, N56, N496, N628);
or OR2 (N747, N738, N656);
buf BUF1 (N748, N734);
xor XOR2 (N749, N685, N440);
and AND3 (N750, N747, N118, N166);
nand NAND4 (N751, N750, N598, N186, N88);
buf BUF1 (N752, N729);
xor XOR2 (N753, N752, N208);
and AND4 (N754, N714, N730, N676, N405);
or OR3 (N755, N751, N475, N396);
nor NOR2 (N756, N753, N176);
not NOT1 (N757, N754);
not NOT1 (N758, N748);
and AND3 (N759, N755, N160, N295);
nor NOR2 (N760, N759, N586);
not NOT1 (N761, N758);
not NOT1 (N762, N749);
nor NOR3 (N763, N761, N62, N411);
nand NAND3 (N764, N756, N598, N362);
buf BUF1 (N765, N763);
or OR4 (N766, N765, N709, N352, N603);
nor NOR2 (N767, N744, N405);
not NOT1 (N768, N766);
nand NAND2 (N769, N762, N203);
and AND4 (N770, N742, N563, N385, N379);
buf BUF1 (N771, N767);
and AND3 (N772, N745, N360, N213);
buf BUF1 (N773, N735);
or OR2 (N774, N757, N639);
xor XOR2 (N775, N746, N689);
nor NOR4 (N776, N773, N701, N45, N497);
and AND4 (N777, N771, N590, N272, N281);
nor NOR4 (N778, N777, N206, N320, N770);
nor NOR2 (N779, N32, N364);
xor XOR2 (N780, N772, N37);
xor XOR2 (N781, N774, N424);
not NOT1 (N782, N768);
xor XOR2 (N783, N778, N442);
or OR3 (N784, N783, N667, N721);
xor XOR2 (N785, N776, N628);
or OR2 (N786, N764, N175);
not NOT1 (N787, N786);
buf BUF1 (N788, N782);
not NOT1 (N789, N780);
and AND2 (N790, N788, N562);
nand NAND4 (N791, N779, N192, N430, N449);
nand NAND4 (N792, N789, N495, N169, N612);
or OR3 (N793, N785, N459, N92);
and AND2 (N794, N760, N748);
and AND3 (N795, N769, N402, N157);
nand NAND2 (N796, N791, N477);
xor XOR2 (N797, N796, N324);
not NOT1 (N798, N781);
xor XOR2 (N799, N797, N485);
not NOT1 (N800, N787);
and AND3 (N801, N792, N285, N506);
xor XOR2 (N802, N775, N412);
xor XOR2 (N803, N800, N796);
buf BUF1 (N804, N798);
xor XOR2 (N805, N790, N353);
or OR4 (N806, N793, N130, N160, N521);
nand NAND3 (N807, N804, N652, N59);
buf BUF1 (N808, N801);
buf BUF1 (N809, N807);
and AND3 (N810, N806, N617, N330);
nand NAND3 (N811, N802, N776, N370);
nor NOR3 (N812, N799, N439, N750);
not NOT1 (N813, N805);
not NOT1 (N814, N811);
xor XOR2 (N815, N813, N559);
xor XOR2 (N816, N794, N76);
not NOT1 (N817, N809);
not NOT1 (N818, N808);
buf BUF1 (N819, N803);
not NOT1 (N820, N814);
buf BUF1 (N821, N810);
not NOT1 (N822, N817);
or OR4 (N823, N821, N735, N492, N815);
buf BUF1 (N824, N698);
nor NOR2 (N825, N820, N39);
xor XOR2 (N826, N816, N342);
nor NOR4 (N827, N823, N181, N603, N701);
not NOT1 (N828, N824);
nor NOR4 (N829, N795, N525, N427, N497);
not NOT1 (N830, N829);
xor XOR2 (N831, N826, N506);
or OR2 (N832, N825, N812);
buf BUF1 (N833, N281);
xor XOR2 (N834, N784, N17);
nor NOR2 (N835, N818, N283);
not NOT1 (N836, N827);
buf BUF1 (N837, N831);
nand NAND4 (N838, N835, N725, N832, N302);
xor XOR2 (N839, N757, N315);
nor NOR4 (N840, N839, N140, N774, N379);
nor NOR4 (N841, N828, N327, N34, N283);
and AND3 (N842, N822, N788, N512);
and AND3 (N843, N841, N126, N738);
or OR2 (N844, N843, N639);
xor XOR2 (N845, N833, N458);
xor XOR2 (N846, N837, N804);
nand NAND4 (N847, N819, N267, N616, N548);
and AND3 (N848, N844, N773, N728);
or OR4 (N849, N847, N316, N472, N497);
nor NOR2 (N850, N834, N579);
buf BUF1 (N851, N838);
nand NAND4 (N852, N836, N748, N254, N470);
nor NOR2 (N853, N848, N728);
and AND4 (N854, N853, N552, N821, N272);
xor XOR2 (N855, N854, N439);
nand NAND4 (N856, N840, N33, N51, N595);
not NOT1 (N857, N846);
not NOT1 (N858, N842);
not NOT1 (N859, N851);
xor XOR2 (N860, N852, N762);
buf BUF1 (N861, N845);
not NOT1 (N862, N830);
not NOT1 (N863, N859);
xor XOR2 (N864, N856, N206);
buf BUF1 (N865, N857);
or OR2 (N866, N849, N805);
not NOT1 (N867, N865);
xor XOR2 (N868, N862, N482);
or OR2 (N869, N860, N693);
and AND2 (N870, N861, N176);
xor XOR2 (N871, N870, N394);
and AND3 (N872, N866, N822, N762);
not NOT1 (N873, N868);
and AND3 (N874, N869, N171, N251);
not NOT1 (N875, N872);
not NOT1 (N876, N871);
buf BUF1 (N877, N875);
xor XOR2 (N878, N863, N343);
not NOT1 (N879, N858);
xor XOR2 (N880, N873, N620);
buf BUF1 (N881, N879);
nand NAND2 (N882, N877, N488);
and AND2 (N883, N882, N213);
buf BUF1 (N884, N855);
buf BUF1 (N885, N881);
not NOT1 (N886, N867);
xor XOR2 (N887, N876, N323);
not NOT1 (N888, N887);
not NOT1 (N889, N874);
not NOT1 (N890, N885);
xor XOR2 (N891, N888, N604);
or OR2 (N892, N889, N66);
nand NAND4 (N893, N891, N15, N578, N694);
or OR4 (N894, N850, N69, N731, N44);
buf BUF1 (N895, N892);
not NOT1 (N896, N864);
nand NAND3 (N897, N890, N269, N4);
nand NAND3 (N898, N883, N690, N74);
buf BUF1 (N899, N893);
not NOT1 (N900, N896);
nand NAND2 (N901, N894, N463);
xor XOR2 (N902, N901, N859);
xor XOR2 (N903, N880, N478);
nor NOR3 (N904, N902, N457, N560);
and AND2 (N905, N904, N136);
nor NOR3 (N906, N900, N598, N817);
and AND2 (N907, N905, N683);
nand NAND4 (N908, N897, N367, N678, N665);
nor NOR4 (N909, N906, N221, N875, N273);
nand NAND3 (N910, N895, N481, N644);
nand NAND2 (N911, N899, N202);
nand NAND4 (N912, N910, N603, N438, N215);
or OR4 (N913, N912, N731, N484, N432);
or OR4 (N914, N878, N199, N323, N392);
xor XOR2 (N915, N911, N508);
and AND4 (N916, N913, N177, N234, N647);
and AND3 (N917, N903, N750, N628);
xor XOR2 (N918, N884, N875);
and AND4 (N919, N908, N411, N846, N610);
nor NOR2 (N920, N914, N299);
xor XOR2 (N921, N916, N216);
or OR2 (N922, N915, N893);
or OR2 (N923, N909, N791);
nand NAND2 (N924, N921, N853);
nand NAND3 (N925, N924, N888, N316);
buf BUF1 (N926, N920);
and AND2 (N927, N886, N910);
xor XOR2 (N928, N922, N23);
and AND3 (N929, N917, N706, N553);
nand NAND4 (N930, N919, N769, N867, N831);
nor NOR2 (N931, N928, N767);
nor NOR3 (N932, N931, N332, N428);
nand NAND2 (N933, N932, N329);
or OR3 (N934, N926, N101, N355);
nand NAND4 (N935, N927, N845, N895, N598);
or OR2 (N936, N925, N305);
not NOT1 (N937, N934);
buf BUF1 (N938, N930);
nor NOR3 (N939, N898, N531, N668);
and AND4 (N940, N937, N619, N262, N175);
nor NOR3 (N941, N938, N519, N42);
nand NAND2 (N942, N939, N378);
not NOT1 (N943, N907);
buf BUF1 (N944, N942);
xor XOR2 (N945, N918, N342);
and AND4 (N946, N933, N1, N935, N265);
nand NAND4 (N947, N815, N213, N715, N803);
buf BUF1 (N948, N945);
or OR4 (N949, N946, N696, N521, N178);
and AND2 (N950, N943, N58);
xor XOR2 (N951, N949, N893);
xor XOR2 (N952, N944, N777);
and AND3 (N953, N947, N584, N878);
and AND3 (N954, N948, N431, N794);
or OR2 (N955, N936, N597);
nor NOR3 (N956, N955, N557, N196);
nor NOR2 (N957, N951, N664);
nor NOR2 (N958, N929, N404);
xor XOR2 (N959, N958, N891);
nor NOR4 (N960, N957, N355, N673, N655);
xor XOR2 (N961, N923, N129);
not NOT1 (N962, N940);
nand NAND3 (N963, N950, N938, N565);
nor NOR3 (N964, N956, N947, N709);
or OR3 (N965, N953, N564, N863);
buf BUF1 (N966, N941);
or OR2 (N967, N961, N157);
xor XOR2 (N968, N965, N394);
not NOT1 (N969, N959);
nand NAND3 (N970, N960, N672, N460);
buf BUF1 (N971, N966);
not NOT1 (N972, N967);
xor XOR2 (N973, N963, N218);
or OR3 (N974, N973, N621, N455);
nor NOR4 (N975, N964, N64, N800, N211);
and AND3 (N976, N970, N464, N431);
xor XOR2 (N977, N969, N652);
buf BUF1 (N978, N952);
nand NAND4 (N979, N976, N332, N56, N781);
nand NAND3 (N980, N972, N567, N183);
and AND4 (N981, N971, N414, N626, N589);
or OR3 (N982, N975, N756, N675);
nor NOR3 (N983, N954, N95, N156);
xor XOR2 (N984, N982, N629);
buf BUF1 (N985, N984);
or OR4 (N986, N981, N398, N124, N818);
nand NAND4 (N987, N978, N258, N458, N692);
or OR2 (N988, N985, N771);
xor XOR2 (N989, N980, N970);
xor XOR2 (N990, N962, N421);
nor NOR4 (N991, N979, N557, N922, N877);
not NOT1 (N992, N977);
nand NAND4 (N993, N991, N290, N303, N621);
buf BUF1 (N994, N988);
nor NOR2 (N995, N968, N576);
nand NAND4 (N996, N990, N411, N801, N3);
nand NAND3 (N997, N992, N658, N430);
xor XOR2 (N998, N995, N787);
or OR2 (N999, N998, N198);
buf BUF1 (N1000, N986);
or OR2 (N1001, N994, N54);
or OR3 (N1002, N999, N728, N290);
and AND4 (N1003, N1002, N490, N606, N407);
or OR3 (N1004, N1001, N112, N382);
xor XOR2 (N1005, N983, N716);
xor XOR2 (N1006, N1005, N528);
and AND3 (N1007, N1003, N932, N58);
nor NOR3 (N1008, N993, N137, N697);
or OR3 (N1009, N989, N184, N392);
xor XOR2 (N1010, N1006, N61);
buf BUF1 (N1011, N1004);
or OR3 (N1012, N987, N370, N707);
nor NOR3 (N1013, N1008, N594, N779);
xor XOR2 (N1014, N1013, N668);
or OR2 (N1015, N1000, N335);
not NOT1 (N1016, N1010);
buf BUF1 (N1017, N974);
not NOT1 (N1018, N1012);
nor NOR2 (N1019, N996, N832);
nand NAND4 (N1020, N1019, N889, N858, N635);
xor XOR2 (N1021, N1020, N2);
xor XOR2 (N1022, N1011, N376);
nor NOR2 (N1023, N1017, N401);
not NOT1 (N1024, N1021);
or OR3 (N1025, N1016, N596, N629);
nand NAND2 (N1026, N997, N704);
xor XOR2 (N1027, N1009, N931);
xor XOR2 (N1028, N1026, N866);
buf BUF1 (N1029, N1015);
nor NOR2 (N1030, N1024, N633);
buf BUF1 (N1031, N1023);
nor NOR3 (N1032, N1030, N886, N124);
buf BUF1 (N1033, N1031);
buf BUF1 (N1034, N1007);
and AND2 (N1035, N1018, N76);
not NOT1 (N1036, N1027);
and AND3 (N1037, N1014, N294, N735);
or OR3 (N1038, N1034, N604, N533);
or OR2 (N1039, N1029, N896);
nor NOR4 (N1040, N1033, N985, N688, N862);
nand NAND4 (N1041, N1037, N275, N270, N539);
nand NAND2 (N1042, N1022, N531);
or OR3 (N1043, N1038, N28, N751);
or OR3 (N1044, N1035, N170, N675);
nand NAND4 (N1045, N1025, N1002, N222, N471);
nand NAND4 (N1046, N1045, N493, N400, N760);
and AND3 (N1047, N1043, N400, N567);
and AND4 (N1048, N1036, N393, N152, N793);
not NOT1 (N1049, N1044);
or OR3 (N1050, N1040, N422, N587);
buf BUF1 (N1051, N1047);
xor XOR2 (N1052, N1039, N1004);
not NOT1 (N1053, N1049);
xor XOR2 (N1054, N1052, N1035);
nor NOR3 (N1055, N1050, N711, N594);
buf BUF1 (N1056, N1051);
and AND3 (N1057, N1048, N1028, N549);
nor NOR2 (N1058, N300, N131);
xor XOR2 (N1059, N1041, N950);
and AND3 (N1060, N1046, N536, N69);
buf BUF1 (N1061, N1056);
xor XOR2 (N1062, N1061, N866);
not NOT1 (N1063, N1055);
not NOT1 (N1064, N1062);
and AND2 (N1065, N1058, N234);
buf BUF1 (N1066, N1042);
xor XOR2 (N1067, N1065, N557);
nor NOR2 (N1068, N1063, N839);
nor NOR3 (N1069, N1054, N651, N866);
nor NOR2 (N1070, N1067, N652);
not NOT1 (N1071, N1066);
and AND2 (N1072, N1053, N228);
xor XOR2 (N1073, N1070, N8);
nor NOR3 (N1074, N1057, N834, N681);
buf BUF1 (N1075, N1069);
nor NOR3 (N1076, N1064, N615, N932);
nand NAND4 (N1077, N1071, N458, N1011, N200);
not NOT1 (N1078, N1068);
xor XOR2 (N1079, N1072, N137);
buf BUF1 (N1080, N1075);
and AND4 (N1081, N1073, N770, N489, N139);
buf BUF1 (N1082, N1077);
not NOT1 (N1083, N1080);
xor XOR2 (N1084, N1076, N486);
buf BUF1 (N1085, N1083);
xor XOR2 (N1086, N1079, N965);
nand NAND4 (N1087, N1085, N212, N644, N1037);
buf BUF1 (N1088, N1074);
or OR3 (N1089, N1081, N326, N1077);
or OR2 (N1090, N1084, N590);
and AND3 (N1091, N1032, N682, N730);
nor NOR4 (N1092, N1091, N292, N517, N446);
buf BUF1 (N1093, N1092);
nand NAND2 (N1094, N1059, N464);
nand NAND4 (N1095, N1086, N754, N850, N1000);
nor NOR3 (N1096, N1090, N12, N360);
not NOT1 (N1097, N1096);
nor NOR2 (N1098, N1093, N460);
nor NOR3 (N1099, N1098, N702, N1086);
or OR4 (N1100, N1078, N544, N594, N296);
not NOT1 (N1101, N1060);
and AND3 (N1102, N1100, N774, N183);
and AND2 (N1103, N1095, N354);
xor XOR2 (N1104, N1101, N616);
nor NOR4 (N1105, N1099, N429, N541, N11);
xor XOR2 (N1106, N1104, N395);
nand NAND2 (N1107, N1094, N348);
or OR2 (N1108, N1107, N1010);
or OR2 (N1109, N1088, N60);
and AND4 (N1110, N1106, N89, N425, N248);
nor NOR3 (N1111, N1089, N823, N1053);
nor NOR4 (N1112, N1111, N408, N664, N634);
xor XOR2 (N1113, N1082, N837);
nor NOR3 (N1114, N1097, N49, N1028);
nor NOR4 (N1115, N1102, N454, N294, N660);
nand NAND3 (N1116, N1113, N226, N930);
buf BUF1 (N1117, N1105);
nor NOR3 (N1118, N1114, N212, N602);
not NOT1 (N1119, N1109);
nand NAND2 (N1120, N1116, N926);
or OR4 (N1121, N1112, N877, N22, N792);
not NOT1 (N1122, N1121);
buf BUF1 (N1123, N1087);
nand NAND4 (N1124, N1115, N527, N553, N980);
buf BUF1 (N1125, N1122);
or OR3 (N1126, N1124, N179, N74);
nor NOR3 (N1127, N1126, N152, N479);
nand NAND3 (N1128, N1119, N31, N196);
nor NOR2 (N1129, N1128, N40);
nand NAND4 (N1130, N1108, N545, N728, N1010);
xor XOR2 (N1131, N1125, N914);
nor NOR2 (N1132, N1127, N117);
not NOT1 (N1133, N1129);
and AND3 (N1134, N1132, N407, N591);
not NOT1 (N1135, N1110);
nand NAND2 (N1136, N1135, N1078);
nor NOR3 (N1137, N1134, N650, N792);
nor NOR4 (N1138, N1118, N687, N365, N704);
or OR3 (N1139, N1131, N543, N31);
xor XOR2 (N1140, N1120, N1037);
nor NOR2 (N1141, N1103, N634);
nand NAND2 (N1142, N1117, N483);
xor XOR2 (N1143, N1130, N145);
buf BUF1 (N1144, N1123);
nand NAND4 (N1145, N1139, N913, N214, N103);
xor XOR2 (N1146, N1136, N326);
xor XOR2 (N1147, N1133, N740);
nor NOR3 (N1148, N1146, N63, N928);
not NOT1 (N1149, N1137);
not NOT1 (N1150, N1140);
not NOT1 (N1151, N1142);
xor XOR2 (N1152, N1144, N728);
nand NAND2 (N1153, N1138, N832);
buf BUF1 (N1154, N1153);
buf BUF1 (N1155, N1152);
xor XOR2 (N1156, N1148, N374);
nand NAND2 (N1157, N1145, N924);
not NOT1 (N1158, N1143);
buf BUF1 (N1159, N1156);
nor NOR4 (N1160, N1157, N760, N974, N88);
or OR3 (N1161, N1149, N218, N1097);
nor NOR3 (N1162, N1150, N540, N92);
xor XOR2 (N1163, N1160, N1104);
or OR2 (N1164, N1159, N854);
buf BUF1 (N1165, N1162);
or OR3 (N1166, N1161, N1024, N444);
or OR2 (N1167, N1158, N1093);
xor XOR2 (N1168, N1151, N864);
nor NOR4 (N1169, N1168, N563, N1044, N243);
or OR2 (N1170, N1164, N973);
xor XOR2 (N1171, N1165, N1092);
or OR2 (N1172, N1155, N762);
nor NOR2 (N1173, N1163, N628);
not NOT1 (N1174, N1170);
not NOT1 (N1175, N1174);
nand NAND2 (N1176, N1141, N615);
nor NOR3 (N1177, N1172, N1113, N34);
buf BUF1 (N1178, N1171);
or OR3 (N1179, N1169, N835, N44);
and AND2 (N1180, N1166, N909);
buf BUF1 (N1181, N1147);
nand NAND2 (N1182, N1179, N1062);
xor XOR2 (N1183, N1180, N173);
nand NAND3 (N1184, N1181, N1116, N62);
xor XOR2 (N1185, N1183, N181);
xor XOR2 (N1186, N1173, N259);
and AND3 (N1187, N1175, N138, N633);
nor NOR3 (N1188, N1182, N1109, N75);
nor NOR4 (N1189, N1187, N93, N854, N596);
buf BUF1 (N1190, N1178);
or OR2 (N1191, N1167, N583);
and AND3 (N1192, N1186, N731, N675);
buf BUF1 (N1193, N1176);
xor XOR2 (N1194, N1185, N913);
nor NOR2 (N1195, N1177, N65);
nor NOR3 (N1196, N1193, N899, N409);
xor XOR2 (N1197, N1195, N375);
or OR4 (N1198, N1192, N1059, N989, N1076);
not NOT1 (N1199, N1197);
nor NOR3 (N1200, N1199, N97, N1032);
and AND2 (N1201, N1198, N523);
nand NAND2 (N1202, N1184, N1103);
buf BUF1 (N1203, N1196);
nor NOR3 (N1204, N1190, N138, N437);
nor NOR4 (N1205, N1202, N203, N1192, N537);
and AND4 (N1206, N1203, N1009, N713, N1073);
or OR2 (N1207, N1194, N1057);
or OR3 (N1208, N1207, N1117, N1053);
buf BUF1 (N1209, N1188);
nand NAND4 (N1210, N1204, N797, N203, N690);
not NOT1 (N1211, N1189);
or OR3 (N1212, N1211, N85, N581);
buf BUF1 (N1213, N1209);
or OR4 (N1214, N1191, N513, N230, N618);
buf BUF1 (N1215, N1212);
nand NAND2 (N1216, N1215, N932);
and AND3 (N1217, N1214, N923, N856);
or OR2 (N1218, N1216, N1095);
xor XOR2 (N1219, N1213, N391);
buf BUF1 (N1220, N1218);
and AND3 (N1221, N1200, N1169, N363);
and AND3 (N1222, N1220, N584, N71);
buf BUF1 (N1223, N1154);
or OR4 (N1224, N1201, N1144, N639, N306);
buf BUF1 (N1225, N1224);
nand NAND4 (N1226, N1208, N47, N1155, N488);
xor XOR2 (N1227, N1206, N1132);
not NOT1 (N1228, N1223);
not NOT1 (N1229, N1227);
nand NAND4 (N1230, N1222, N892, N183, N764);
nor NOR3 (N1231, N1210, N3, N856);
xor XOR2 (N1232, N1221, N704);
and AND4 (N1233, N1217, N269, N295, N26);
and AND2 (N1234, N1228, N837);
or OR2 (N1235, N1230, N394);
xor XOR2 (N1236, N1235, N500);
nor NOR3 (N1237, N1225, N250, N588);
nand NAND2 (N1238, N1237, N604);
and AND2 (N1239, N1231, N1202);
xor XOR2 (N1240, N1205, N229);
xor XOR2 (N1241, N1229, N149);
nor NOR2 (N1242, N1236, N1045);
not NOT1 (N1243, N1240);
xor XOR2 (N1244, N1238, N412);
not NOT1 (N1245, N1234);
buf BUF1 (N1246, N1233);
nor NOR3 (N1247, N1245, N311, N974);
nand NAND2 (N1248, N1241, N499);
nand NAND2 (N1249, N1244, N896);
nand NAND4 (N1250, N1248, N914, N540, N865);
nand NAND4 (N1251, N1247, N1214, N69, N1096);
buf BUF1 (N1252, N1219);
not NOT1 (N1253, N1246);
or OR2 (N1254, N1251, N588);
nor NOR3 (N1255, N1243, N395, N203);
not NOT1 (N1256, N1253);
xor XOR2 (N1257, N1250, N879);
buf BUF1 (N1258, N1226);
not NOT1 (N1259, N1254);
not NOT1 (N1260, N1249);
or OR3 (N1261, N1239, N581, N134);
not NOT1 (N1262, N1260);
and AND4 (N1263, N1255, N185, N559, N4);
not NOT1 (N1264, N1232);
or OR4 (N1265, N1264, N1067, N1210, N628);
and AND4 (N1266, N1263, N522, N762, N1033);
or OR2 (N1267, N1262, N767);
nor NOR3 (N1268, N1265, N717, N1167);
xor XOR2 (N1269, N1267, N1147);
xor XOR2 (N1270, N1258, N771);
nand NAND2 (N1271, N1257, N1114);
and AND3 (N1272, N1261, N1199, N893);
buf BUF1 (N1273, N1269);
or OR2 (N1274, N1272, N514);
not NOT1 (N1275, N1271);
and AND3 (N1276, N1252, N409, N252);
or OR2 (N1277, N1276, N571);
or OR4 (N1278, N1275, N676, N1050, N794);
nand NAND2 (N1279, N1273, N1083);
nand NAND3 (N1280, N1274, N891, N324);
and AND2 (N1281, N1279, N471);
and AND3 (N1282, N1280, N807, N1150);
buf BUF1 (N1283, N1281);
or OR4 (N1284, N1268, N1167, N1079, N622);
and AND2 (N1285, N1256, N1173);
and AND4 (N1286, N1285, N557, N998, N1108);
buf BUF1 (N1287, N1277);
and AND4 (N1288, N1283, N45, N205, N493);
not NOT1 (N1289, N1282);
nand NAND3 (N1290, N1289, N984, N961);
or OR3 (N1291, N1242, N1278, N227);
nor NOR3 (N1292, N1125, N501, N316);
or OR2 (N1293, N1259, N647);
or OR3 (N1294, N1287, N1047, N374);
and AND2 (N1295, N1266, N658);
or OR3 (N1296, N1293, N376, N240);
or OR2 (N1297, N1288, N308);
nand NAND4 (N1298, N1295, N110, N81, N991);
xor XOR2 (N1299, N1291, N389);
not NOT1 (N1300, N1292);
nor NOR2 (N1301, N1297, N510);
and AND2 (N1302, N1296, N35);
or OR4 (N1303, N1290, N39, N517, N876);
and AND3 (N1304, N1301, N554, N650);
xor XOR2 (N1305, N1286, N498);
not NOT1 (N1306, N1284);
or OR2 (N1307, N1302, N485);
buf BUF1 (N1308, N1306);
buf BUF1 (N1309, N1308);
buf BUF1 (N1310, N1270);
or OR3 (N1311, N1305, N1153, N565);
not NOT1 (N1312, N1299);
nand NAND3 (N1313, N1294, N201, N1046);
nor NOR4 (N1314, N1300, N140, N1246, N1292);
or OR4 (N1315, N1314, N533, N205, N965);
buf BUF1 (N1316, N1315);
or OR2 (N1317, N1298, N122);
not NOT1 (N1318, N1307);
not NOT1 (N1319, N1318);
nand NAND2 (N1320, N1313, N661);
nor NOR3 (N1321, N1310, N138, N500);
nand NAND2 (N1322, N1303, N391);
and AND3 (N1323, N1317, N692, N192);
or OR3 (N1324, N1304, N1309, N113);
nand NAND3 (N1325, N551, N337, N1151);
or OR4 (N1326, N1321, N128, N228, N252);
and AND3 (N1327, N1324, N1008, N823);
not NOT1 (N1328, N1316);
xor XOR2 (N1329, N1327, N862);
not NOT1 (N1330, N1311);
nand NAND4 (N1331, N1320, N863, N1323, N144);
not NOT1 (N1332, N994);
nor NOR2 (N1333, N1319, N592);
or OR2 (N1334, N1329, N645);
xor XOR2 (N1335, N1326, N829);
buf BUF1 (N1336, N1331);
buf BUF1 (N1337, N1334);
xor XOR2 (N1338, N1332, N542);
xor XOR2 (N1339, N1337, N1152);
nor NOR3 (N1340, N1338, N327, N502);
or OR4 (N1341, N1333, N378, N977, N774);
nor NOR2 (N1342, N1339, N512);
xor XOR2 (N1343, N1336, N284);
not NOT1 (N1344, N1335);
nor NOR4 (N1345, N1340, N1302, N1227, N672);
nor NOR2 (N1346, N1344, N1162);
nor NOR3 (N1347, N1330, N22, N1046);
nand NAND2 (N1348, N1346, N552);
and AND2 (N1349, N1328, N165);
xor XOR2 (N1350, N1348, N34);
nand NAND2 (N1351, N1347, N118);
or OR4 (N1352, N1325, N1081, N1178, N1098);
nor NOR2 (N1353, N1343, N238);
or OR4 (N1354, N1312, N103, N992, N409);
and AND2 (N1355, N1341, N725);
and AND2 (N1356, N1352, N181);
nor NOR3 (N1357, N1354, N1281, N354);
nand NAND3 (N1358, N1351, N456, N12);
not NOT1 (N1359, N1353);
xor XOR2 (N1360, N1358, N323);
nand NAND4 (N1361, N1345, N882, N94, N981);
nor NOR2 (N1362, N1361, N359);
or OR4 (N1363, N1349, N592, N1188, N1213);
not NOT1 (N1364, N1357);
buf BUF1 (N1365, N1350);
nand NAND4 (N1366, N1359, N246, N351, N367);
xor XOR2 (N1367, N1355, N700);
nand NAND4 (N1368, N1342, N680, N1330, N309);
nand NAND2 (N1369, N1364, N926);
and AND3 (N1370, N1365, N384, N321);
not NOT1 (N1371, N1369);
buf BUF1 (N1372, N1322);
or OR4 (N1373, N1363, N899, N404, N12);
not NOT1 (N1374, N1366);
and AND2 (N1375, N1368, N81);
nor NOR3 (N1376, N1360, N634, N952);
xor XOR2 (N1377, N1362, N209);
or OR4 (N1378, N1370, N147, N969, N607);
nand NAND3 (N1379, N1378, N127, N820);
buf BUF1 (N1380, N1375);
or OR2 (N1381, N1372, N802);
or OR4 (N1382, N1377, N1380, N366, N826);
nand NAND2 (N1383, N89, N878);
or OR2 (N1384, N1367, N270);
buf BUF1 (N1385, N1356);
nand NAND4 (N1386, N1374, N818, N518, N934);
buf BUF1 (N1387, N1373);
xor XOR2 (N1388, N1385, N395);
not NOT1 (N1389, N1381);
or OR2 (N1390, N1383, N852);
not NOT1 (N1391, N1382);
nor NOR2 (N1392, N1384, N240);
nor NOR3 (N1393, N1388, N907, N204);
nand NAND2 (N1394, N1376, N122);
or OR3 (N1395, N1393, N793, N122);
nor NOR4 (N1396, N1389, N447, N261, N748);
nor NOR4 (N1397, N1379, N890, N915, N569);
xor XOR2 (N1398, N1397, N791);
xor XOR2 (N1399, N1387, N615);
nand NAND4 (N1400, N1386, N1142, N377, N588);
not NOT1 (N1401, N1394);
not NOT1 (N1402, N1390);
xor XOR2 (N1403, N1401, N490);
nor NOR2 (N1404, N1403, N1323);
or OR2 (N1405, N1399, N121);
nand NAND3 (N1406, N1371, N1317, N987);
buf BUF1 (N1407, N1392);
not NOT1 (N1408, N1398);
not NOT1 (N1409, N1396);
and AND2 (N1410, N1391, N1209);
or OR3 (N1411, N1408, N745, N904);
not NOT1 (N1412, N1410);
or OR2 (N1413, N1406, N1284);
nor NOR3 (N1414, N1407, N358, N425);
buf BUF1 (N1415, N1405);
and AND2 (N1416, N1402, N12);
nand NAND3 (N1417, N1409, N984, N194);
xor XOR2 (N1418, N1411, N803);
buf BUF1 (N1419, N1415);
xor XOR2 (N1420, N1400, N620);
buf BUF1 (N1421, N1420);
and AND2 (N1422, N1418, N1007);
xor XOR2 (N1423, N1414, N1319);
nor NOR2 (N1424, N1413, N1163);
xor XOR2 (N1425, N1421, N122);
buf BUF1 (N1426, N1412);
nor NOR4 (N1427, N1416, N844, N30, N152);
buf BUF1 (N1428, N1404);
not NOT1 (N1429, N1419);
not NOT1 (N1430, N1423);
or OR3 (N1431, N1395, N1092, N777);
not NOT1 (N1432, N1430);
xor XOR2 (N1433, N1426, N609);
buf BUF1 (N1434, N1417);
or OR4 (N1435, N1433, N837, N558, N920);
and AND2 (N1436, N1435, N330);
nand NAND2 (N1437, N1424, N438);
nand NAND2 (N1438, N1434, N391);
buf BUF1 (N1439, N1432);
nand NAND2 (N1440, N1437, N166);
or OR3 (N1441, N1431, N455, N839);
nor NOR3 (N1442, N1422, N868, N993);
and AND2 (N1443, N1438, N1370);
nand NAND3 (N1444, N1429, N325, N204);
nand NAND2 (N1445, N1439, N404);
and AND3 (N1446, N1440, N769, N414);
and AND2 (N1447, N1443, N963);
buf BUF1 (N1448, N1445);
xor XOR2 (N1449, N1448, N574);
nand NAND4 (N1450, N1444, N743, N1159, N1136);
xor XOR2 (N1451, N1441, N522);
nor NOR2 (N1452, N1425, N223);
xor XOR2 (N1453, N1446, N731);
not NOT1 (N1454, N1449);
and AND4 (N1455, N1436, N791, N171, N257);
xor XOR2 (N1456, N1427, N675);
not NOT1 (N1457, N1450);
and AND2 (N1458, N1452, N436);
and AND2 (N1459, N1451, N1339);
nand NAND2 (N1460, N1458, N822);
buf BUF1 (N1461, N1460);
or OR4 (N1462, N1461, N776, N589, N1150);
nor NOR4 (N1463, N1447, N581, N797, N1153);
nand NAND2 (N1464, N1428, N1329);
nor NOR2 (N1465, N1457, N780);
buf BUF1 (N1466, N1464);
and AND4 (N1467, N1459, N384, N137, N936);
or OR2 (N1468, N1454, N958);
xor XOR2 (N1469, N1468, N1277);
not NOT1 (N1470, N1467);
xor XOR2 (N1471, N1462, N657);
xor XOR2 (N1472, N1442, N1190);
buf BUF1 (N1473, N1463);
xor XOR2 (N1474, N1473, N1372);
xor XOR2 (N1475, N1470, N1350);
not NOT1 (N1476, N1475);
and AND3 (N1477, N1469, N1168, N728);
buf BUF1 (N1478, N1466);
and AND3 (N1479, N1474, N688, N1270);
xor XOR2 (N1480, N1478, N692);
not NOT1 (N1481, N1476);
or OR4 (N1482, N1456, N1457, N1422, N737);
nand NAND3 (N1483, N1471, N400, N1169);
or OR3 (N1484, N1472, N434, N703);
xor XOR2 (N1485, N1483, N81);
or OR4 (N1486, N1477, N990, N569, N1358);
buf BUF1 (N1487, N1485);
buf BUF1 (N1488, N1487);
nor NOR2 (N1489, N1480, N595);
xor XOR2 (N1490, N1488, N188);
nand NAND4 (N1491, N1486, N86, N1428, N393);
nand NAND3 (N1492, N1455, N810, N1140);
and AND2 (N1493, N1465, N1362);
buf BUF1 (N1494, N1481);
or OR3 (N1495, N1491, N547, N604);
xor XOR2 (N1496, N1453, N221);
xor XOR2 (N1497, N1484, N554);
or OR2 (N1498, N1496, N253);
or OR4 (N1499, N1494, N965, N1307, N1428);
nand NAND2 (N1500, N1482, N1415);
nand NAND4 (N1501, N1499, N1430, N695, N771);
or OR2 (N1502, N1501, N927);
nor NOR3 (N1503, N1479, N419, N1204);
not NOT1 (N1504, N1489);
not NOT1 (N1505, N1504);
not NOT1 (N1506, N1505);
and AND4 (N1507, N1490, N640, N1074, N626);
nand NAND3 (N1508, N1497, N50, N1102);
nand NAND4 (N1509, N1495, N199, N1338, N378);
or OR4 (N1510, N1498, N875, N999, N444);
nand NAND4 (N1511, N1506, N4, N1182, N316);
xor XOR2 (N1512, N1511, N647);
xor XOR2 (N1513, N1493, N1342);
and AND2 (N1514, N1507, N354);
nor NOR3 (N1515, N1508, N532, N1064);
xor XOR2 (N1516, N1512, N827);
xor XOR2 (N1517, N1510, N476);
xor XOR2 (N1518, N1502, N1049);
buf BUF1 (N1519, N1516);
nand NAND3 (N1520, N1509, N619, N1505);
not NOT1 (N1521, N1520);
not NOT1 (N1522, N1492);
nor NOR4 (N1523, N1500, N879, N40, N788);
and AND2 (N1524, N1523, N405);
not NOT1 (N1525, N1519);
nand NAND2 (N1526, N1522, N845);
not NOT1 (N1527, N1521);
or OR2 (N1528, N1527, N179);
not NOT1 (N1529, N1518);
buf BUF1 (N1530, N1503);
not NOT1 (N1531, N1515);
buf BUF1 (N1532, N1517);
nor NOR4 (N1533, N1525, N995, N1482, N930);
or OR4 (N1534, N1528, N74, N537, N673);
not NOT1 (N1535, N1529);
and AND2 (N1536, N1532, N1456);
nand NAND4 (N1537, N1534, N750, N1050, N1027);
not NOT1 (N1538, N1536);
nor NOR4 (N1539, N1514, N1472, N1215, N601);
or OR2 (N1540, N1535, N1118);
buf BUF1 (N1541, N1533);
not NOT1 (N1542, N1540);
and AND4 (N1543, N1541, N4, N545, N1239);
and AND4 (N1544, N1530, N1039, N756, N939);
nor NOR2 (N1545, N1537, N873);
and AND4 (N1546, N1524, N758, N1034, N893);
or OR2 (N1547, N1513, N632);
nor NOR2 (N1548, N1546, N928);
and AND3 (N1549, N1547, N99, N377);
xor XOR2 (N1550, N1538, N63);
and AND3 (N1551, N1548, N246, N14);
nand NAND2 (N1552, N1545, N764);
not NOT1 (N1553, N1531);
or OR3 (N1554, N1550, N404, N126);
nor NOR3 (N1555, N1542, N655, N1102);
xor XOR2 (N1556, N1553, N287);
and AND2 (N1557, N1543, N132);
buf BUF1 (N1558, N1539);
or OR2 (N1559, N1551, N291);
and AND2 (N1560, N1526, N230);
nand NAND3 (N1561, N1549, N253, N1);
not NOT1 (N1562, N1559);
not NOT1 (N1563, N1554);
and AND2 (N1564, N1562, N692);
buf BUF1 (N1565, N1561);
nor NOR3 (N1566, N1544, N519, N1098);
and AND3 (N1567, N1552, N319, N340);
or OR4 (N1568, N1556, N594, N24, N930);
buf BUF1 (N1569, N1564);
nand NAND2 (N1570, N1569, N282);
xor XOR2 (N1571, N1568, N615);
nor NOR4 (N1572, N1566, N696, N59, N1184);
and AND3 (N1573, N1560, N1155, N23);
or OR4 (N1574, N1558, N1366, N111, N815);
nor NOR3 (N1575, N1572, N865, N41);
not NOT1 (N1576, N1557);
not NOT1 (N1577, N1555);
and AND4 (N1578, N1571, N721, N222, N866);
buf BUF1 (N1579, N1574);
nand NAND2 (N1580, N1577, N812);
and AND3 (N1581, N1579, N762, N1557);
nand NAND4 (N1582, N1578, N23, N969, N500);
nand NAND3 (N1583, N1576, N671, N951);
nand NAND3 (N1584, N1567, N1378, N152);
buf BUF1 (N1585, N1565);
or OR2 (N1586, N1575, N168);
or OR3 (N1587, N1583, N1480, N1352);
not NOT1 (N1588, N1581);
not NOT1 (N1589, N1582);
or OR4 (N1590, N1580, N861, N1561, N384);
buf BUF1 (N1591, N1589);
buf BUF1 (N1592, N1590);
xor XOR2 (N1593, N1563, N824);
nand NAND4 (N1594, N1584, N1135, N1067, N582);
xor XOR2 (N1595, N1570, N975);
xor XOR2 (N1596, N1573, N1251);
xor XOR2 (N1597, N1594, N448);
not NOT1 (N1598, N1596);
buf BUF1 (N1599, N1593);
and AND3 (N1600, N1591, N379, N711);
and AND4 (N1601, N1597, N67, N250, N696);
not NOT1 (N1602, N1588);
buf BUF1 (N1603, N1599);
nand NAND3 (N1604, N1601, N377, N987);
xor XOR2 (N1605, N1600, N412);
or OR2 (N1606, N1602, N697);
not NOT1 (N1607, N1606);
buf BUF1 (N1608, N1587);
not NOT1 (N1609, N1598);
and AND3 (N1610, N1585, N565, N907);
or OR3 (N1611, N1610, N647, N1337);
nand NAND2 (N1612, N1607, N163);
or OR2 (N1613, N1586, N30);
not NOT1 (N1614, N1603);
nor NOR3 (N1615, N1611, N461, N235);
and AND4 (N1616, N1615, N331, N695, N546);
or OR4 (N1617, N1616, N209, N182, N630);
not NOT1 (N1618, N1605);
and AND2 (N1619, N1595, N34);
nor NOR3 (N1620, N1604, N843, N1220);
nor NOR4 (N1621, N1619, N737, N5, N856);
or OR3 (N1622, N1620, N492, N264);
nor NOR3 (N1623, N1618, N1563, N410);
nor NOR3 (N1624, N1612, N1557, N768);
xor XOR2 (N1625, N1613, N790);
not NOT1 (N1626, N1621);
nand NAND2 (N1627, N1626, N876);
or OR3 (N1628, N1625, N1464, N322);
buf BUF1 (N1629, N1622);
or OR3 (N1630, N1592, N1614, N746);
xor XOR2 (N1631, N103, N1118);
or OR3 (N1632, N1630, N195, N800);
nand NAND4 (N1633, N1608, N1180, N1384, N1059);
not NOT1 (N1634, N1624);
xor XOR2 (N1635, N1609, N452);
buf BUF1 (N1636, N1627);
buf BUF1 (N1637, N1633);
nand NAND4 (N1638, N1628, N1094, N480, N44);
xor XOR2 (N1639, N1634, N731);
nor NOR3 (N1640, N1631, N45, N433);
nor NOR3 (N1641, N1635, N455, N996);
or OR2 (N1642, N1632, N512);
xor XOR2 (N1643, N1638, N596);
xor XOR2 (N1644, N1617, N820);
buf BUF1 (N1645, N1640);
and AND4 (N1646, N1645, N507, N895, N1562);
nor NOR4 (N1647, N1637, N873, N1381, N745);
or OR2 (N1648, N1644, N92);
not NOT1 (N1649, N1641);
nor NOR3 (N1650, N1647, N271, N107);
or OR3 (N1651, N1648, N783, N1464);
and AND3 (N1652, N1646, N38, N591);
buf BUF1 (N1653, N1652);
nand NAND3 (N1654, N1629, N506, N247);
nand NAND4 (N1655, N1649, N1301, N9, N1359);
xor XOR2 (N1656, N1650, N607);
xor XOR2 (N1657, N1639, N836);
and AND4 (N1658, N1656, N798, N1167, N582);
xor XOR2 (N1659, N1657, N427);
xor XOR2 (N1660, N1643, N371);
buf BUF1 (N1661, N1636);
nand NAND4 (N1662, N1659, N1651, N1628, N62);
nand NAND2 (N1663, N1087, N207);
nand NAND2 (N1664, N1661, N234);
nand NAND3 (N1665, N1658, N1023, N123);
xor XOR2 (N1666, N1662, N1445);
and AND3 (N1667, N1654, N1051, N389);
buf BUF1 (N1668, N1664);
nor NOR3 (N1669, N1663, N956, N1057);
buf BUF1 (N1670, N1655);
nor NOR3 (N1671, N1669, N429, N1571);
nor NOR3 (N1672, N1667, N1292, N619);
nor NOR4 (N1673, N1665, N649, N1589, N553);
or OR3 (N1674, N1668, N671, N1141);
buf BUF1 (N1675, N1672);
and AND2 (N1676, N1670, N492);
nor NOR2 (N1677, N1653, N1237);
nand NAND4 (N1678, N1677, N532, N835, N917);
buf BUF1 (N1679, N1674);
xor XOR2 (N1680, N1666, N900);
nand NAND3 (N1681, N1671, N496, N1592);
buf BUF1 (N1682, N1642);
not NOT1 (N1683, N1678);
and AND2 (N1684, N1673, N1027);
nand NAND2 (N1685, N1682, N1597);
xor XOR2 (N1686, N1679, N1139);
buf BUF1 (N1687, N1623);
nor NOR3 (N1688, N1680, N368, N330);
and AND3 (N1689, N1687, N339, N213);
nor NOR2 (N1690, N1688, N754);
or OR3 (N1691, N1685, N1498, N1610);
nor NOR3 (N1692, N1686, N1549, N1172);
nand NAND4 (N1693, N1689, N402, N1408, N1035);
nor NOR4 (N1694, N1681, N888, N1646, N1206);
and AND4 (N1695, N1660, N1057, N315, N1205);
buf BUF1 (N1696, N1676);
nand NAND4 (N1697, N1684, N903, N1549, N276);
xor XOR2 (N1698, N1691, N1331);
nor NOR4 (N1699, N1698, N154, N1105, N1283);
buf BUF1 (N1700, N1675);
nand NAND2 (N1701, N1696, N100);
nor NOR3 (N1702, N1683, N789, N896);
xor XOR2 (N1703, N1690, N184);
nand NAND2 (N1704, N1693, N1390);
nor NOR2 (N1705, N1695, N1057);
or OR4 (N1706, N1705, N1167, N147, N1093);
and AND3 (N1707, N1699, N970, N1345);
and AND2 (N1708, N1704, N89);
nor NOR2 (N1709, N1706, N1163);
buf BUF1 (N1710, N1694);
or OR2 (N1711, N1710, N108);
or OR3 (N1712, N1707, N737, N652);
or OR3 (N1713, N1712, N252, N64);
nor NOR2 (N1714, N1700, N209);
not NOT1 (N1715, N1703);
nand NAND4 (N1716, N1702, N1302, N1424, N668);
or OR4 (N1717, N1692, N1167, N412, N1634);
nand NAND3 (N1718, N1716, N685, N1377);
xor XOR2 (N1719, N1717, N1556);
or OR2 (N1720, N1708, N626);
and AND2 (N1721, N1720, N1058);
buf BUF1 (N1722, N1711);
not NOT1 (N1723, N1714);
nand NAND3 (N1724, N1715, N1649, N105);
nor NOR2 (N1725, N1723, N1678);
and AND4 (N1726, N1713, N1259, N1123, N442);
xor XOR2 (N1727, N1701, N409);
nand NAND4 (N1728, N1721, N1589, N1078, N966);
not NOT1 (N1729, N1722);
xor XOR2 (N1730, N1719, N1311);
not NOT1 (N1731, N1724);
xor XOR2 (N1732, N1731, N1092);
not NOT1 (N1733, N1727);
or OR2 (N1734, N1730, N1277);
buf BUF1 (N1735, N1732);
and AND2 (N1736, N1697, N1490);
xor XOR2 (N1737, N1725, N995);
not NOT1 (N1738, N1729);
nand NAND2 (N1739, N1718, N451);
xor XOR2 (N1740, N1737, N1304);
nand NAND4 (N1741, N1740, N413, N1246, N136);
buf BUF1 (N1742, N1709);
buf BUF1 (N1743, N1735);
or OR2 (N1744, N1726, N794);
or OR2 (N1745, N1743, N907);
xor XOR2 (N1746, N1738, N1203);
and AND4 (N1747, N1733, N589, N456, N1582);
or OR4 (N1748, N1736, N1121, N504, N1180);
nor NOR4 (N1749, N1746, N1172, N554, N1527);
and AND2 (N1750, N1742, N580);
nand NAND4 (N1751, N1728, N200, N1218, N820);
nand NAND2 (N1752, N1739, N1216);
buf BUF1 (N1753, N1750);
and AND4 (N1754, N1741, N939, N943, N1753);
xor XOR2 (N1755, N544, N1535);
xor XOR2 (N1756, N1755, N596);
buf BUF1 (N1757, N1745);
buf BUF1 (N1758, N1747);
xor XOR2 (N1759, N1757, N1500);
xor XOR2 (N1760, N1734, N1371);
nor NOR4 (N1761, N1754, N598, N1253, N951);
or OR4 (N1762, N1744, N629, N1186, N782);
and AND3 (N1763, N1749, N1762, N857);
buf BUF1 (N1764, N1126);
nor NOR4 (N1765, N1760, N169, N673, N1541);
nand NAND3 (N1766, N1751, N806, N344);
xor XOR2 (N1767, N1765, N1079);
buf BUF1 (N1768, N1756);
and AND3 (N1769, N1766, N1744, N1417);
not NOT1 (N1770, N1768);
buf BUF1 (N1771, N1752);
not NOT1 (N1772, N1770);
and AND3 (N1773, N1758, N1276, N1028);
nand NAND4 (N1774, N1773, N1351, N500, N856);
and AND2 (N1775, N1761, N1726);
nand NAND4 (N1776, N1759, N72, N1182, N788);
and AND2 (N1777, N1774, N1559);
or OR2 (N1778, N1763, N310);
nor NOR3 (N1779, N1771, N1099, N806);
or OR4 (N1780, N1748, N459, N1100, N1535);
not NOT1 (N1781, N1777);
xor XOR2 (N1782, N1779, N1660);
nor NOR4 (N1783, N1767, N727, N1231, N28);
nor NOR2 (N1784, N1772, N540);
nand NAND2 (N1785, N1784, N343);
or OR4 (N1786, N1782, N1294, N477, N1621);
buf BUF1 (N1787, N1778);
buf BUF1 (N1788, N1786);
not NOT1 (N1789, N1787);
not NOT1 (N1790, N1769);
buf BUF1 (N1791, N1776);
buf BUF1 (N1792, N1775);
nand NAND4 (N1793, N1764, N106, N159, N642);
and AND4 (N1794, N1781, N179, N1597, N1653);
buf BUF1 (N1795, N1789);
not NOT1 (N1796, N1788);
nor NOR2 (N1797, N1795, N162);
nand NAND3 (N1798, N1793, N719, N243);
or OR4 (N1799, N1797, N32, N516, N1327);
buf BUF1 (N1800, N1799);
xor XOR2 (N1801, N1794, N1448);
and AND3 (N1802, N1790, N73, N656);
not NOT1 (N1803, N1792);
nand NAND3 (N1804, N1785, N1159, N31);
nor NOR3 (N1805, N1780, N1605, N1031);
not NOT1 (N1806, N1783);
nand NAND2 (N1807, N1805, N797);
xor XOR2 (N1808, N1807, N1334);
buf BUF1 (N1809, N1798);
xor XOR2 (N1810, N1809, N792);
nand NAND3 (N1811, N1796, N1472, N1467);
not NOT1 (N1812, N1804);
and AND4 (N1813, N1801, N251, N1472, N1707);
or OR4 (N1814, N1811, N429, N187, N787);
nor NOR4 (N1815, N1806, N1720, N1758, N1121);
and AND4 (N1816, N1800, N541, N814, N317);
and AND2 (N1817, N1791, N765);
buf BUF1 (N1818, N1812);
or OR2 (N1819, N1818, N1018);
xor XOR2 (N1820, N1810, N1640);
xor XOR2 (N1821, N1802, N752);
or OR4 (N1822, N1808, N856, N1771, N948);
nand NAND3 (N1823, N1817, N1008, N1005);
xor XOR2 (N1824, N1815, N332);
xor XOR2 (N1825, N1822, N428);
or OR4 (N1826, N1819, N1785, N1206, N1509);
xor XOR2 (N1827, N1816, N406);
or OR2 (N1828, N1823, N1);
buf BUF1 (N1829, N1813);
nand NAND2 (N1830, N1829, N451);
nor NOR3 (N1831, N1830, N1761, N1281);
or OR3 (N1832, N1824, N1185, N650);
buf BUF1 (N1833, N1803);
or OR3 (N1834, N1827, N954, N602);
not NOT1 (N1835, N1834);
xor XOR2 (N1836, N1828, N1662);
nor NOR3 (N1837, N1825, N1824, N689);
xor XOR2 (N1838, N1821, N1561);
or OR2 (N1839, N1826, N232);
or OR3 (N1840, N1838, N302, N1285);
nand NAND3 (N1841, N1836, N1666, N1147);
and AND4 (N1842, N1839, N1027, N458, N1651);
xor XOR2 (N1843, N1840, N363);
buf BUF1 (N1844, N1814);
not NOT1 (N1845, N1833);
nor NOR3 (N1846, N1835, N989, N529);
xor XOR2 (N1847, N1843, N54);
nand NAND4 (N1848, N1831, N1691, N581, N1118);
buf BUF1 (N1849, N1842);
or OR3 (N1850, N1849, N278, N788);
xor XOR2 (N1851, N1844, N1685);
or OR4 (N1852, N1848, N1337, N518, N717);
buf BUF1 (N1853, N1852);
not NOT1 (N1854, N1850);
buf BUF1 (N1855, N1846);
nand NAND4 (N1856, N1845, N438, N1054, N388);
xor XOR2 (N1857, N1820, N315);
or OR3 (N1858, N1857, N241, N448);
buf BUF1 (N1859, N1855);
buf BUF1 (N1860, N1851);
or OR3 (N1861, N1832, N17, N387);
buf BUF1 (N1862, N1860);
or OR3 (N1863, N1859, N425, N1027);
and AND4 (N1864, N1853, N730, N178, N1482);
xor XOR2 (N1865, N1854, N1469);
and AND3 (N1866, N1837, N1312, N1865);
buf BUF1 (N1867, N145);
nand NAND3 (N1868, N1847, N93, N1319);
nand NAND3 (N1869, N1841, N1840, N538);
not NOT1 (N1870, N1866);
nor NOR2 (N1871, N1870, N1240);
not NOT1 (N1872, N1864);
not NOT1 (N1873, N1861);
and AND4 (N1874, N1868, N53, N151, N389);
not NOT1 (N1875, N1863);
nor NOR3 (N1876, N1869, N176, N1636);
or OR3 (N1877, N1871, N172, N1635);
xor XOR2 (N1878, N1867, N729);
not NOT1 (N1879, N1862);
xor XOR2 (N1880, N1879, N800);
nor NOR3 (N1881, N1877, N766, N221);
nor NOR3 (N1882, N1873, N1553, N1131);
not NOT1 (N1883, N1878);
nand NAND2 (N1884, N1858, N182);
not NOT1 (N1885, N1875);
nand NAND3 (N1886, N1856, N519, N1351);
or OR2 (N1887, N1876, N662);
or OR2 (N1888, N1884, N1726);
or OR4 (N1889, N1885, N128, N26, N1312);
or OR3 (N1890, N1888, N1330, N291);
or OR3 (N1891, N1883, N351, N487);
not NOT1 (N1892, N1890);
xor XOR2 (N1893, N1881, N220);
and AND4 (N1894, N1893, N1217, N828, N1382);
nor NOR4 (N1895, N1894, N1350, N779, N1725);
nand NAND3 (N1896, N1886, N158, N594);
buf BUF1 (N1897, N1882);
nor NOR3 (N1898, N1874, N1670, N375);
and AND4 (N1899, N1887, N1017, N1240, N1380);
xor XOR2 (N1900, N1895, N894);
xor XOR2 (N1901, N1900, N1342);
and AND3 (N1902, N1880, N1191, N1800);
nand NAND3 (N1903, N1902, N178, N537);
or OR4 (N1904, N1898, N776, N418, N862);
xor XOR2 (N1905, N1901, N1148);
and AND2 (N1906, N1892, N204);
nor NOR4 (N1907, N1891, N1182, N1236, N877);
xor XOR2 (N1908, N1903, N1381);
xor XOR2 (N1909, N1907, N970);
nand NAND4 (N1910, N1904, N162, N1455, N893);
nand NAND2 (N1911, N1910, N1236);
nor NOR2 (N1912, N1909, N939);
nor NOR4 (N1913, N1872, N767, N404, N1634);
and AND2 (N1914, N1905, N1765);
not NOT1 (N1915, N1908);
not NOT1 (N1916, N1913);
or OR2 (N1917, N1915, N1868);
not NOT1 (N1918, N1906);
xor XOR2 (N1919, N1914, N1058);
nor NOR2 (N1920, N1889, N609);
nor NOR4 (N1921, N1896, N648, N687, N314);
nor NOR2 (N1922, N1918, N305);
nor NOR2 (N1923, N1921, N124);
or OR4 (N1924, N1917, N1098, N368, N1791);
or OR3 (N1925, N1922, N280, N1380);
nand NAND2 (N1926, N1897, N758);
or OR2 (N1927, N1919, N1585);
xor XOR2 (N1928, N1912, N1694);
not NOT1 (N1929, N1923);
xor XOR2 (N1930, N1899, N1171);
nor NOR3 (N1931, N1924, N1237, N283);
nor NOR3 (N1932, N1925, N862, N1180);
or OR3 (N1933, N1916, N249, N1821);
not NOT1 (N1934, N1911);
not NOT1 (N1935, N1933);
and AND4 (N1936, N1931, N581, N1931, N1672);
buf BUF1 (N1937, N1932);
xor XOR2 (N1938, N1936, N1841);
and AND2 (N1939, N1930, N205);
buf BUF1 (N1940, N1935);
nor NOR2 (N1941, N1937, N805);
and AND3 (N1942, N1927, N427, N633);
nor NOR4 (N1943, N1929, N326, N1850, N1589);
buf BUF1 (N1944, N1920);
not NOT1 (N1945, N1940);
nand NAND3 (N1946, N1939, N147, N608);
nor NOR4 (N1947, N1941, N847, N964, N1660);
nor NOR3 (N1948, N1938, N884, N247);
buf BUF1 (N1949, N1948);
not NOT1 (N1950, N1946);
xor XOR2 (N1951, N1945, N1184);
and AND4 (N1952, N1926, N1195, N442, N1200);
or OR3 (N1953, N1928, N181, N1296);
nand NAND2 (N1954, N1947, N896);
nand NAND4 (N1955, N1934, N339, N173, N1037);
or OR3 (N1956, N1942, N817, N301);
not NOT1 (N1957, N1956);
nand NAND4 (N1958, N1952, N1585, N941, N1055);
buf BUF1 (N1959, N1954);
nand NAND2 (N1960, N1959, N1906);
nor NOR4 (N1961, N1960, N1716, N537, N395);
nand NAND3 (N1962, N1953, N575, N1133);
nor NOR4 (N1963, N1943, N526, N1486, N1669);
nor NOR3 (N1964, N1955, N107, N918);
buf BUF1 (N1965, N1962);
xor XOR2 (N1966, N1963, N1555);
or OR2 (N1967, N1961, N875);
and AND4 (N1968, N1966, N930, N68, N1671);
and AND4 (N1969, N1958, N960, N774, N897);
nor NOR2 (N1970, N1950, N1912);
not NOT1 (N1971, N1944);
and AND4 (N1972, N1967, N714, N175, N1867);
buf BUF1 (N1973, N1965);
nor NOR2 (N1974, N1949, N1861);
buf BUF1 (N1975, N1969);
nor NOR4 (N1976, N1951, N1787, N365, N1712);
nand NAND3 (N1977, N1975, N1853, N868);
or OR3 (N1978, N1964, N916, N1547);
or OR4 (N1979, N1972, N835, N519, N1343);
xor XOR2 (N1980, N1978, N356);
nor NOR4 (N1981, N1979, N1910, N892, N1188);
or OR4 (N1982, N1968, N1925, N1764, N247);
nand NAND2 (N1983, N1976, N1020);
and AND2 (N1984, N1982, N1980);
not NOT1 (N1985, N1597);
and AND3 (N1986, N1957, N453, N1153);
xor XOR2 (N1987, N1985, N1276);
nand NAND3 (N1988, N1983, N71, N135);
not NOT1 (N1989, N1984);
not NOT1 (N1990, N1971);
nor NOR3 (N1991, N1986, N1025, N1844);
nor NOR3 (N1992, N1973, N331, N1061);
buf BUF1 (N1993, N1970);
and AND4 (N1994, N1990, N818, N1504, N499);
not NOT1 (N1995, N1987);
nor NOR2 (N1996, N1981, N854);
buf BUF1 (N1997, N1992);
buf BUF1 (N1998, N1991);
xor XOR2 (N1999, N1997, N1012);
xor XOR2 (N2000, N1993, N1019);
and AND3 (N2001, N1996, N1138, N1729);
nor NOR4 (N2002, N1977, N1521, N601, N1198);
and AND4 (N2003, N1989, N325, N1696, N1520);
and AND3 (N2004, N2000, N1554, N226);
not NOT1 (N2005, N1988);
not NOT1 (N2006, N1995);
or OR2 (N2007, N2001, N1580);
not NOT1 (N2008, N2005);
nor NOR3 (N2009, N2003, N454, N613);
xor XOR2 (N2010, N2008, N1619);
not NOT1 (N2011, N2007);
buf BUF1 (N2012, N2006);
nand NAND2 (N2013, N2002, N655);
not NOT1 (N2014, N1974);
buf BUF1 (N2015, N2011);
nor NOR2 (N2016, N2014, N86);
not NOT1 (N2017, N1999);
xor XOR2 (N2018, N2017, N1224);
nand NAND4 (N2019, N2015, N1590, N1025, N118);
nand NAND2 (N2020, N2016, N3);
and AND3 (N2021, N2019, N1640, N1659);
not NOT1 (N2022, N2018);
not NOT1 (N2023, N2010);
or OR3 (N2024, N2012, N1549, N28);
nand NAND3 (N2025, N1998, N685, N222);
xor XOR2 (N2026, N2013, N1307);
not NOT1 (N2027, N2020);
and AND4 (N2028, N2024, N1936, N9, N793);
xor XOR2 (N2029, N2025, N1675);
or OR3 (N2030, N2028, N1140, N818);
xor XOR2 (N2031, N2023, N315);
nand NAND4 (N2032, N2009, N856, N1633, N390);
xor XOR2 (N2033, N2027, N872);
xor XOR2 (N2034, N2022, N251);
nand NAND4 (N2035, N2004, N855, N186, N1154);
xor XOR2 (N2036, N2030, N1344);
and AND4 (N2037, N1994, N855, N560, N126);
and AND2 (N2038, N2033, N14);
or OR3 (N2039, N2035, N316, N391);
buf BUF1 (N2040, N2021);
or OR4 (N2041, N2031, N138, N440, N184);
not NOT1 (N2042, N2032);
buf BUF1 (N2043, N2029);
nand NAND4 (N2044, N2039, N1383, N1420, N1054);
nor NOR4 (N2045, N2036, N550, N1758, N1394);
buf BUF1 (N2046, N2042);
nor NOR4 (N2047, N2034, N142, N797, N206);
nand NAND4 (N2048, N2047, N983, N1010, N700);
or OR3 (N2049, N2026, N1250, N1895);
or OR4 (N2050, N2046, N1719, N1157, N1284);
buf BUF1 (N2051, N2040);
nor NOR2 (N2052, N2041, N1294);
not NOT1 (N2053, N2037);
and AND4 (N2054, N2044, N145, N444, N803);
not NOT1 (N2055, N2054);
or OR3 (N2056, N2049, N505, N67);
nor NOR2 (N2057, N2038, N1657);
nor NOR3 (N2058, N2055, N133, N1936);
nand NAND2 (N2059, N2045, N327);
xor XOR2 (N2060, N2048, N1080);
nor NOR3 (N2061, N2056, N622, N1530);
xor XOR2 (N2062, N2053, N1702);
or OR4 (N2063, N2043, N16, N201, N195);
xor XOR2 (N2064, N2063, N689);
or OR3 (N2065, N2057, N1451, N673);
xor XOR2 (N2066, N2052, N754);
buf BUF1 (N2067, N2061);
not NOT1 (N2068, N2050);
buf BUF1 (N2069, N2065);
not NOT1 (N2070, N2069);
and AND2 (N2071, N2068, N1873);
not NOT1 (N2072, N2070);
nand NAND3 (N2073, N2059, N811, N1479);
nand NAND4 (N2074, N2058, N1687, N1271, N1940);
nand NAND3 (N2075, N2067, N506, N811);
or OR3 (N2076, N2074, N309, N457);
buf BUF1 (N2077, N2071);
nand NAND3 (N2078, N2064, N950, N2071);
xor XOR2 (N2079, N2076, N1509);
xor XOR2 (N2080, N2066, N1156);
nand NAND2 (N2081, N2051, N833);
nand NAND3 (N2082, N2077, N2076, N1503);
and AND4 (N2083, N2079, N480, N2043, N1659);
not NOT1 (N2084, N2081);
nor NOR3 (N2085, N2075, N309, N1560);
nand NAND3 (N2086, N2080, N116, N1724);
nor NOR3 (N2087, N2083, N1737, N816);
or OR4 (N2088, N2073, N963, N55, N636);
and AND4 (N2089, N2087, N1016, N1550, N76);
or OR3 (N2090, N2072, N1310, N1514);
not NOT1 (N2091, N2088);
nand NAND2 (N2092, N2062, N1016);
nor NOR3 (N2093, N2085, N1550, N699);
or OR2 (N2094, N2092, N462);
nand NAND2 (N2095, N2089, N527);
and AND3 (N2096, N2082, N89, N754);
not NOT1 (N2097, N2078);
and AND2 (N2098, N2090, N679);
not NOT1 (N2099, N2097);
and AND4 (N2100, N2094, N1281, N740, N1766);
xor XOR2 (N2101, N2100, N1226);
or OR3 (N2102, N2095, N728, N435);
nor NOR2 (N2103, N2060, N1984);
not NOT1 (N2104, N2086);
nor NOR4 (N2105, N2096, N1172, N1721, N1221);
xor XOR2 (N2106, N2102, N804);
nor NOR4 (N2107, N2098, N56, N348, N1228);
nand NAND2 (N2108, N2105, N1107);
or OR2 (N2109, N2103, N1259);
not NOT1 (N2110, N2106);
xor XOR2 (N2111, N2110, N1742);
nor NOR3 (N2112, N2108, N1814, N913);
nor NOR2 (N2113, N2107, N1150);
nand NAND3 (N2114, N2109, N1902, N814);
nand NAND2 (N2115, N2099, N690);
nand NAND2 (N2116, N2113, N1693);
nor NOR3 (N2117, N2114, N1454, N414);
nor NOR3 (N2118, N2111, N918, N356);
buf BUF1 (N2119, N2091);
and AND3 (N2120, N2101, N1549, N343);
xor XOR2 (N2121, N2120, N1922);
nor NOR3 (N2122, N2121, N1876, N1730);
not NOT1 (N2123, N2118);
xor XOR2 (N2124, N2093, N766);
or OR3 (N2125, N2123, N2049, N923);
nor NOR2 (N2126, N2117, N176);
buf BUF1 (N2127, N2119);
xor XOR2 (N2128, N2115, N1150);
buf BUF1 (N2129, N2104);
not NOT1 (N2130, N2084);
nand NAND2 (N2131, N2129, N1002);
nand NAND2 (N2132, N2128, N1676);
and AND2 (N2133, N2130, N759);
and AND3 (N2134, N2122, N1026, N1388);
xor XOR2 (N2135, N2127, N1179);
xor XOR2 (N2136, N2112, N594);
xor XOR2 (N2137, N2126, N1848);
buf BUF1 (N2138, N2132);
nor NOR3 (N2139, N2124, N1352, N12);
not NOT1 (N2140, N2138);
not NOT1 (N2141, N2139);
nor NOR3 (N2142, N2141, N269, N1831);
and AND4 (N2143, N2136, N354, N231, N1563);
or OR2 (N2144, N2135, N362);
xor XOR2 (N2145, N2142, N588);
nor NOR2 (N2146, N2125, N1754);
and AND4 (N2147, N2145, N1602, N1860, N237);
and AND3 (N2148, N2146, N275, N776);
buf BUF1 (N2149, N2137);
not NOT1 (N2150, N2149);
or OR2 (N2151, N2116, N1191);
and AND2 (N2152, N2133, N667);
not NOT1 (N2153, N2140);
xor XOR2 (N2154, N2144, N823);
xor XOR2 (N2155, N2134, N103);
not NOT1 (N2156, N2147);
not NOT1 (N2157, N2155);
not NOT1 (N2158, N2153);
buf BUF1 (N2159, N2151);
xor XOR2 (N2160, N2157, N761);
not NOT1 (N2161, N2159);
and AND3 (N2162, N2154, N412, N560);
not NOT1 (N2163, N2160);
nor NOR3 (N2164, N2152, N1863, N1318);
nand NAND3 (N2165, N2163, N1105, N1103);
nand NAND4 (N2166, N2148, N1831, N1787, N1642);
and AND2 (N2167, N2131, N1079);
or OR3 (N2168, N2167, N718, N393);
and AND4 (N2169, N2165, N1298, N129, N2064);
nand NAND2 (N2170, N2158, N1087);
and AND3 (N2171, N2161, N46, N1483);
nor NOR3 (N2172, N2164, N1633, N1940);
not NOT1 (N2173, N2162);
buf BUF1 (N2174, N2150);
not NOT1 (N2175, N2156);
or OR2 (N2176, N2143, N1158);
buf BUF1 (N2177, N2172);
or OR4 (N2178, N2171, N496, N1986, N1437);
buf BUF1 (N2179, N2170);
nand NAND4 (N2180, N2169, N29, N1798, N423);
buf BUF1 (N2181, N2178);
xor XOR2 (N2182, N2179, N1742);
nor NOR3 (N2183, N2177, N623, N1660);
xor XOR2 (N2184, N2166, N1010);
and AND3 (N2185, N2168, N603, N229);
or OR4 (N2186, N2174, N560, N593, N2034);
buf BUF1 (N2187, N2185);
not NOT1 (N2188, N2176);
nor NOR4 (N2189, N2187, N1436, N78, N948);
nor NOR4 (N2190, N2175, N1132, N1582, N1031);
buf BUF1 (N2191, N2190);
nand NAND2 (N2192, N2191, N653);
and AND2 (N2193, N2173, N1326);
or OR3 (N2194, N2182, N2010, N504);
nand NAND4 (N2195, N2180, N1381, N120, N220);
and AND2 (N2196, N2184, N1908);
nor NOR3 (N2197, N2189, N2138, N2057);
or OR3 (N2198, N2183, N1276, N1851);
not NOT1 (N2199, N2194);
not NOT1 (N2200, N2195);
nor NOR4 (N2201, N2196, N388, N618, N591);
not NOT1 (N2202, N2201);
nand NAND2 (N2203, N2199, N484);
not NOT1 (N2204, N2202);
and AND2 (N2205, N2203, N2159);
not NOT1 (N2206, N2192);
nand NAND4 (N2207, N2193, N1333, N1063, N1392);
nor NOR3 (N2208, N2186, N631, N1946);
nor NOR4 (N2209, N2206, N1685, N1472, N2121);
xor XOR2 (N2210, N2205, N291);
nor NOR4 (N2211, N2207, N826, N586, N435);
nor NOR4 (N2212, N2208, N1401, N2190, N2061);
buf BUF1 (N2213, N2198);
xor XOR2 (N2214, N2211, N2180);
xor XOR2 (N2215, N2213, N701);
xor XOR2 (N2216, N2197, N1266);
or OR3 (N2217, N2181, N1282, N1078);
or OR2 (N2218, N2216, N2203);
nor NOR4 (N2219, N2212, N1879, N142, N718);
nand NAND3 (N2220, N2217, N1295, N544);
nor NOR3 (N2221, N2214, N559, N566);
nand NAND3 (N2222, N2219, N94, N1766);
buf BUF1 (N2223, N2188);
and AND4 (N2224, N2218, N1688, N2048, N1982);
or OR4 (N2225, N2209, N659, N1742, N1054);
nor NOR2 (N2226, N2224, N2194);
nand NAND4 (N2227, N2225, N989, N2158, N805);
nand NAND3 (N2228, N2210, N1701, N1347);
and AND2 (N2229, N2226, N1120);
or OR3 (N2230, N2220, N2032, N2084);
xor XOR2 (N2231, N2228, N1922);
or OR2 (N2232, N2231, N431);
xor XOR2 (N2233, N2221, N221);
buf BUF1 (N2234, N2215);
nor NOR4 (N2235, N2200, N547, N96, N1107);
nor NOR4 (N2236, N2227, N2093, N120, N1212);
nor NOR2 (N2237, N2235, N671);
nand NAND2 (N2238, N2229, N1127);
xor XOR2 (N2239, N2233, N1982);
or OR4 (N2240, N2238, N742, N1717, N1573);
not NOT1 (N2241, N2239);
buf BUF1 (N2242, N2222);
buf BUF1 (N2243, N2223);
and AND4 (N2244, N2236, N1229, N1554, N1889);
nor NOR2 (N2245, N2232, N1691);
and AND4 (N2246, N2241, N1718, N1717, N339);
xor XOR2 (N2247, N2242, N580);
buf BUF1 (N2248, N2245);
buf BUF1 (N2249, N2234);
or OR3 (N2250, N2204, N2185, N1347);
nor NOR3 (N2251, N2250, N883, N1114);
nor NOR2 (N2252, N2240, N1548);
not NOT1 (N2253, N2251);
buf BUF1 (N2254, N2248);
buf BUF1 (N2255, N2253);
and AND3 (N2256, N2252, N1476, N2035);
and AND3 (N2257, N2249, N735, N1693);
buf BUF1 (N2258, N2256);
buf BUF1 (N2259, N2244);
xor XOR2 (N2260, N2230, N1090);
not NOT1 (N2261, N2255);
buf BUF1 (N2262, N2258);
nor NOR4 (N2263, N2237, N1537, N1782, N157);
or OR3 (N2264, N2247, N2, N1757);
not NOT1 (N2265, N2262);
and AND4 (N2266, N2246, N2157, N2023, N758);
buf BUF1 (N2267, N2257);
or OR2 (N2268, N2254, N1585);
buf BUF1 (N2269, N2268);
not NOT1 (N2270, N2261);
buf BUF1 (N2271, N2259);
xor XOR2 (N2272, N2265, N1413);
or OR2 (N2273, N2243, N1951);
xor XOR2 (N2274, N2270, N1115);
xor XOR2 (N2275, N2267, N1667);
buf BUF1 (N2276, N2263);
xor XOR2 (N2277, N2271, N484);
not NOT1 (N2278, N2277);
xor XOR2 (N2279, N2276, N1718);
xor XOR2 (N2280, N2260, N1415);
xor XOR2 (N2281, N2264, N996);
nor NOR2 (N2282, N2275, N34);
and AND2 (N2283, N2274, N1946);
not NOT1 (N2284, N2266);
buf BUF1 (N2285, N2273);
and AND3 (N2286, N2281, N761, N1428);
buf BUF1 (N2287, N2286);
or OR4 (N2288, N2282, N909, N2186, N855);
buf BUF1 (N2289, N2288);
nor NOR3 (N2290, N2284, N1796, N132);
xor XOR2 (N2291, N2272, N659);
or OR2 (N2292, N2287, N169);
nand NAND4 (N2293, N2269, N1571, N2035, N1792);
or OR3 (N2294, N2283, N1431, N887);
nor NOR4 (N2295, N2279, N2097, N1524, N461);
buf BUF1 (N2296, N2280);
or OR4 (N2297, N2295, N1103, N379, N1546);
buf BUF1 (N2298, N2278);
buf BUF1 (N2299, N2297);
buf BUF1 (N2300, N2293);
buf BUF1 (N2301, N2290);
buf BUF1 (N2302, N2301);
and AND2 (N2303, N2292, N1133);
xor XOR2 (N2304, N2285, N273);
xor XOR2 (N2305, N2289, N1122);
and AND2 (N2306, N2294, N1845);
and AND2 (N2307, N2300, N1410);
buf BUF1 (N2308, N2291);
not NOT1 (N2309, N2299);
nor NOR2 (N2310, N2305, N1155);
or OR3 (N2311, N2298, N967, N2233);
and AND3 (N2312, N2310, N985, N1874);
and AND2 (N2313, N2302, N1778);
or OR4 (N2314, N2312, N1895, N1556, N927);
or OR2 (N2315, N2308, N2002);
and AND3 (N2316, N2306, N918, N179);
and AND2 (N2317, N2307, N343);
nor NOR4 (N2318, N2303, N635, N1964, N506);
xor XOR2 (N2319, N2313, N1675);
nor NOR3 (N2320, N2311, N2101, N1455);
nand NAND3 (N2321, N2314, N557, N1029);
nor NOR3 (N2322, N2315, N160, N926);
nand NAND4 (N2323, N2318, N1854, N335, N649);
and AND4 (N2324, N2296, N1247, N10, N2300);
not NOT1 (N2325, N2324);
or OR3 (N2326, N2317, N86, N2265);
or OR4 (N2327, N2325, N1459, N808, N480);
nor NOR3 (N2328, N2319, N1378, N1921);
not NOT1 (N2329, N2323);
xor XOR2 (N2330, N2316, N2109);
nand NAND3 (N2331, N2309, N547, N1344);
not NOT1 (N2332, N2329);
nand NAND4 (N2333, N2327, N1320, N2145, N963);
xor XOR2 (N2334, N2328, N931);
buf BUF1 (N2335, N2304);
nor NOR3 (N2336, N2321, N2180, N208);
xor XOR2 (N2337, N2320, N890);
and AND4 (N2338, N2334, N1754, N82, N400);
nor NOR3 (N2339, N2338, N1409, N1521);
buf BUF1 (N2340, N2332);
or OR2 (N2341, N2330, N2245);
not NOT1 (N2342, N2337);
not NOT1 (N2343, N2336);
nor NOR3 (N2344, N2326, N948, N1737);
xor XOR2 (N2345, N2341, N1333);
not NOT1 (N2346, N2335);
xor XOR2 (N2347, N2333, N285);
nor NOR2 (N2348, N2345, N2067);
xor XOR2 (N2349, N2331, N57);
and AND3 (N2350, N2346, N1954, N1206);
buf BUF1 (N2351, N2347);
buf BUF1 (N2352, N2339);
buf BUF1 (N2353, N2340);
nor NOR4 (N2354, N2353, N1882, N692, N1301);
nor NOR2 (N2355, N2322, N2121);
xor XOR2 (N2356, N2349, N774);
or OR2 (N2357, N2355, N1700);
or OR2 (N2358, N2343, N153);
xor XOR2 (N2359, N2350, N939);
or OR2 (N2360, N2359, N870);
nor NOR3 (N2361, N2354, N1702, N159);
nor NOR4 (N2362, N2356, N327, N374, N187);
buf BUF1 (N2363, N2357);
buf BUF1 (N2364, N2351);
and AND4 (N2365, N2362, N1799, N2127, N1997);
nor NOR2 (N2366, N2361, N343);
nand NAND4 (N2367, N2363, N1360, N46, N104);
buf BUF1 (N2368, N2348);
or OR4 (N2369, N2352, N1362, N1609, N691);
or OR3 (N2370, N2344, N720, N455);
not NOT1 (N2371, N2367);
not NOT1 (N2372, N2369);
buf BUF1 (N2373, N2366);
xor XOR2 (N2374, N2372, N902);
not NOT1 (N2375, N2360);
and AND3 (N2376, N2374, N393, N993);
nand NAND2 (N2377, N2358, N2279);
xor XOR2 (N2378, N2342, N1784);
or OR2 (N2379, N2376, N2076);
not NOT1 (N2380, N2365);
or OR4 (N2381, N2379, N944, N994, N1911);
nand NAND2 (N2382, N2380, N1679);
nor NOR4 (N2383, N2370, N725, N2353, N2355);
not NOT1 (N2384, N2383);
and AND2 (N2385, N2378, N2272);
not NOT1 (N2386, N2364);
not NOT1 (N2387, N2385);
xor XOR2 (N2388, N2387, N1333);
and AND4 (N2389, N2377, N2178, N378, N1139);
xor XOR2 (N2390, N2373, N183);
buf BUF1 (N2391, N2388);
and AND2 (N2392, N2371, N1707);
or OR4 (N2393, N2389, N2341, N767, N25);
not NOT1 (N2394, N2390);
or OR4 (N2395, N2391, N1042, N566, N476);
xor XOR2 (N2396, N2395, N2361);
xor XOR2 (N2397, N2381, N941);
and AND2 (N2398, N2396, N1843);
nor NOR2 (N2399, N2392, N1638);
or OR2 (N2400, N2393, N21);
and AND4 (N2401, N2368, N337, N2117, N1187);
nand NAND4 (N2402, N2384, N2327, N166, N1929);
and AND2 (N2403, N2375, N1159);
nand NAND4 (N2404, N2398, N179, N1342, N1528);
or OR4 (N2405, N2403, N2019, N780, N25);
nor NOR2 (N2406, N2382, N2303);
nor NOR4 (N2407, N2386, N879, N2191, N1013);
xor XOR2 (N2408, N2397, N82);
or OR3 (N2409, N2406, N1574, N432);
and AND2 (N2410, N2404, N174);
nor NOR4 (N2411, N2410, N2183, N384, N1538);
nor NOR2 (N2412, N2411, N2049);
and AND3 (N2413, N2400, N2087, N1712);
and AND4 (N2414, N2409, N764, N1061, N420);
buf BUF1 (N2415, N2394);
nor NOR2 (N2416, N2412, N380);
buf BUF1 (N2417, N2405);
and AND2 (N2418, N2413, N418);
nand NAND4 (N2419, N2416, N395, N1251, N1656);
xor XOR2 (N2420, N2401, N86);
xor XOR2 (N2421, N2399, N711);
and AND4 (N2422, N2414, N2389, N688, N1207);
or OR3 (N2423, N2415, N201, N1725);
buf BUF1 (N2424, N2402);
buf BUF1 (N2425, N2424);
or OR4 (N2426, N2420, N691, N235, N689);
nand NAND2 (N2427, N2417, N1907);
not NOT1 (N2428, N2419);
and AND4 (N2429, N2422, N1834, N2043, N1758);
or OR4 (N2430, N2428, N2143, N548, N750);
and AND4 (N2431, N2408, N1845, N1475, N1067);
buf BUF1 (N2432, N2418);
nand NAND3 (N2433, N2407, N1202, N214);
and AND2 (N2434, N2421, N1207);
and AND4 (N2435, N2425, N1922, N1747, N2278);
or OR4 (N2436, N2432, N1204, N178, N1055);
or OR4 (N2437, N2429, N1901, N1214, N169);
nor NOR3 (N2438, N2434, N1976, N35);
and AND4 (N2439, N2431, N2046, N804, N1649);
or OR3 (N2440, N2433, N711, N1792);
nand NAND4 (N2441, N2426, N534, N855, N252);
nand NAND2 (N2442, N2441, N1811);
or OR3 (N2443, N2430, N1493, N1648);
nand NAND3 (N2444, N2427, N73, N389);
or OR3 (N2445, N2444, N2122, N423);
buf BUF1 (N2446, N2445);
nand NAND3 (N2447, N2439, N178, N1006);
xor XOR2 (N2448, N2442, N435);
not NOT1 (N2449, N2440);
and AND3 (N2450, N2449, N1881, N2413);
not NOT1 (N2451, N2443);
nand NAND2 (N2452, N2436, N1713);
nor NOR3 (N2453, N2451, N1417, N1235);
not NOT1 (N2454, N2446);
nand NAND3 (N2455, N2437, N1869, N1522);
or OR2 (N2456, N2455, N615);
nor NOR3 (N2457, N2435, N2417, N597);
or OR4 (N2458, N2423, N342, N891, N1684);
not NOT1 (N2459, N2453);
not NOT1 (N2460, N2452);
and AND2 (N2461, N2447, N307);
buf BUF1 (N2462, N2460);
nor NOR2 (N2463, N2461, N21);
nand NAND2 (N2464, N2438, N27);
nor NOR4 (N2465, N2456, N1457, N1245, N497);
not NOT1 (N2466, N2465);
buf BUF1 (N2467, N2448);
nand NAND4 (N2468, N2459, N1408, N1594, N2236);
not NOT1 (N2469, N2463);
xor XOR2 (N2470, N2466, N2459);
or OR3 (N2471, N2470, N1631, N863);
buf BUF1 (N2472, N2458);
xor XOR2 (N2473, N2471, N2173);
xor XOR2 (N2474, N2464, N273);
xor XOR2 (N2475, N2457, N472);
nor NOR3 (N2476, N2450, N1934, N208);
not NOT1 (N2477, N2454);
and AND3 (N2478, N2473, N2066, N437);
nand NAND4 (N2479, N2467, N261, N348, N1826);
and AND4 (N2480, N2475, N1286, N1964, N2424);
and AND2 (N2481, N2472, N1841);
xor XOR2 (N2482, N2478, N37);
and AND3 (N2483, N2480, N799, N1985);
and AND3 (N2484, N2477, N1579, N2416);
not NOT1 (N2485, N2469);
and AND2 (N2486, N2484, N945);
buf BUF1 (N2487, N2479);
xor XOR2 (N2488, N2468, N1722);
xor XOR2 (N2489, N2476, N252);
or OR3 (N2490, N2486, N1806, N2214);
buf BUF1 (N2491, N2474);
not NOT1 (N2492, N2489);
nand NAND2 (N2493, N2491, N1382);
nand NAND3 (N2494, N2481, N2312, N21);
not NOT1 (N2495, N2462);
not NOT1 (N2496, N2483);
nand NAND4 (N2497, N2490, N701, N2114, N1895);
not NOT1 (N2498, N2482);
not NOT1 (N2499, N2497);
nand NAND2 (N2500, N2492, N610);
and AND3 (N2501, N2500, N1033, N1396);
nand NAND4 (N2502, N2499, N1321, N1278, N882);
and AND2 (N2503, N2493, N972);
or OR3 (N2504, N2502, N414, N2230);
nor NOR4 (N2505, N2495, N2205, N545, N577);
nor NOR3 (N2506, N2494, N1974, N2431);
nand NAND4 (N2507, N2498, N1392, N2112, N620);
nand NAND3 (N2508, N2507, N1529, N1206);
xor XOR2 (N2509, N2506, N1021);
nor NOR2 (N2510, N2509, N1262);
buf BUF1 (N2511, N2503);
nand NAND2 (N2512, N2511, N604);
and AND3 (N2513, N2512, N1024, N886);
xor XOR2 (N2514, N2504, N1239);
xor XOR2 (N2515, N2508, N1760);
xor XOR2 (N2516, N2501, N1947);
nor NOR3 (N2517, N2488, N2115, N21);
xor XOR2 (N2518, N2514, N1224);
or OR4 (N2519, N2510, N1488, N1589, N654);
or OR4 (N2520, N2485, N1264, N328, N319);
and AND4 (N2521, N2518, N385, N1518, N1323);
xor XOR2 (N2522, N2521, N724);
nand NAND4 (N2523, N2496, N884, N66, N2106);
not NOT1 (N2524, N2519);
or OR2 (N2525, N2517, N1715);
nor NOR3 (N2526, N2513, N1515, N1029);
not NOT1 (N2527, N2522);
nor NOR2 (N2528, N2520, N210);
xor XOR2 (N2529, N2523, N1062);
xor XOR2 (N2530, N2515, N1200);
and AND4 (N2531, N2528, N1077, N1958, N558);
xor XOR2 (N2532, N2487, N565);
xor XOR2 (N2533, N2516, N1408);
not NOT1 (N2534, N2531);
not NOT1 (N2535, N2530);
buf BUF1 (N2536, N2532);
nand NAND4 (N2537, N2534, N491, N1411, N661);
nand NAND4 (N2538, N2535, N249, N2011, N798);
and AND4 (N2539, N2533, N635, N2244, N947);
buf BUF1 (N2540, N2525);
xor XOR2 (N2541, N2527, N857);
or OR4 (N2542, N2538, N2319, N2307, N1559);
and AND3 (N2543, N2526, N1315, N652);
not NOT1 (N2544, N2529);
xor XOR2 (N2545, N2544, N2382);
buf BUF1 (N2546, N2505);
and AND2 (N2547, N2540, N27);
nor NOR4 (N2548, N2543, N2075, N2479, N1311);
xor XOR2 (N2549, N2537, N2398);
or OR2 (N2550, N2542, N679);
nor NOR3 (N2551, N2536, N1233, N985);
buf BUF1 (N2552, N2551);
or OR2 (N2553, N2524, N2295);
buf BUF1 (N2554, N2549);
not NOT1 (N2555, N2541);
buf BUF1 (N2556, N2550);
or OR3 (N2557, N2545, N1146, N2373);
not NOT1 (N2558, N2556);
and AND2 (N2559, N2539, N1843);
xor XOR2 (N2560, N2558, N202);
or OR3 (N2561, N2548, N2435, N679);
not NOT1 (N2562, N2560);
xor XOR2 (N2563, N2557, N756);
buf BUF1 (N2564, N2563);
nand NAND2 (N2565, N2553, N492);
xor XOR2 (N2566, N2554, N491);
xor XOR2 (N2567, N2562, N1541);
and AND2 (N2568, N2546, N640);
or OR4 (N2569, N2559, N1305, N1253, N1403);
nand NAND4 (N2570, N2566, N487, N1749, N619);
xor XOR2 (N2571, N2564, N2328);
buf BUF1 (N2572, N2555);
not NOT1 (N2573, N2561);
not NOT1 (N2574, N2567);
or OR2 (N2575, N2574, N1369);
and AND4 (N2576, N2575, N230, N329, N1198);
and AND4 (N2577, N2547, N2512, N204, N171);
or OR4 (N2578, N2568, N950, N166, N1389);
and AND4 (N2579, N2571, N1285, N2007, N1503);
and AND4 (N2580, N2565, N839, N992, N2088);
xor XOR2 (N2581, N2569, N1018);
xor XOR2 (N2582, N2572, N1962);
buf BUF1 (N2583, N2581);
nand NAND4 (N2584, N2578, N2125, N2556, N763);
nor NOR3 (N2585, N2580, N499, N1915);
xor XOR2 (N2586, N2584, N1944);
nor NOR2 (N2587, N2585, N280);
nor NOR3 (N2588, N2552, N755, N458);
not NOT1 (N2589, N2588);
nor NOR3 (N2590, N2576, N2260, N33);
not NOT1 (N2591, N2579);
buf BUF1 (N2592, N2577);
not NOT1 (N2593, N2587);
xor XOR2 (N2594, N2586, N523);
xor XOR2 (N2595, N2594, N550);
not NOT1 (N2596, N2589);
nand NAND2 (N2597, N2592, N464);
not NOT1 (N2598, N2591);
xor XOR2 (N2599, N2597, N1848);
buf BUF1 (N2600, N2582);
not NOT1 (N2601, N2599);
not NOT1 (N2602, N2573);
nand NAND2 (N2603, N2593, N740);
nand NAND4 (N2604, N2570, N1180, N2404, N1540);
or OR2 (N2605, N2603, N1182);
and AND2 (N2606, N2605, N215);
nor NOR3 (N2607, N2601, N1185, N2101);
nand NAND3 (N2608, N2604, N791, N126);
and AND4 (N2609, N2608, N1504, N600, N2033);
not NOT1 (N2610, N2602);
not NOT1 (N2611, N2590);
not NOT1 (N2612, N2610);
not NOT1 (N2613, N2598);
and AND2 (N2614, N2607, N601);
nand NAND4 (N2615, N2609, N564, N1033, N1539);
or OR3 (N2616, N2596, N849, N254);
nand NAND2 (N2617, N2616, N2220);
nand NAND3 (N2618, N2583, N2545, N1258);
or OR3 (N2619, N2617, N399, N1668);
not NOT1 (N2620, N2615);
not NOT1 (N2621, N2612);
not NOT1 (N2622, N2613);
or OR4 (N2623, N2618, N843, N2254, N1447);
nor NOR2 (N2624, N2622, N2081);
or OR2 (N2625, N2611, N2404);
buf BUF1 (N2626, N2623);
nand NAND3 (N2627, N2606, N1882, N937);
or OR2 (N2628, N2620, N2294);
not NOT1 (N2629, N2595);
xor XOR2 (N2630, N2619, N1935);
nor NOR2 (N2631, N2614, N598);
or OR2 (N2632, N2627, N2041);
and AND4 (N2633, N2629, N117, N29, N140);
and AND4 (N2634, N2625, N549, N774, N2454);
or OR2 (N2635, N2626, N1142);
buf BUF1 (N2636, N2621);
and AND2 (N2637, N2630, N1273);
buf BUF1 (N2638, N2634);
not NOT1 (N2639, N2632);
nor NOR3 (N2640, N2638, N32, N993);
nand NAND3 (N2641, N2628, N541, N1748);
and AND3 (N2642, N2637, N1087, N142);
not NOT1 (N2643, N2636);
nand NAND3 (N2644, N2642, N283, N521);
nor NOR2 (N2645, N2635, N211);
or OR2 (N2646, N2631, N1373);
nor NOR4 (N2647, N2645, N2102, N1335, N2070);
buf BUF1 (N2648, N2646);
nor NOR4 (N2649, N2624, N1336, N1327, N243);
buf BUF1 (N2650, N2600);
and AND2 (N2651, N2649, N2156);
nor NOR3 (N2652, N2647, N1553, N1486);
nand NAND4 (N2653, N2643, N1569, N433, N936);
not NOT1 (N2654, N2644);
not NOT1 (N2655, N2653);
nor NOR4 (N2656, N2639, N55, N1372, N958);
and AND4 (N2657, N2652, N411, N353, N1214);
or OR4 (N2658, N2654, N79, N1187, N1973);
nand NAND3 (N2659, N2641, N874, N1);
xor XOR2 (N2660, N2648, N105);
nor NOR4 (N2661, N2657, N340, N408, N1148);
nand NAND3 (N2662, N2659, N2416, N2177);
not NOT1 (N2663, N2656);
or OR2 (N2664, N2650, N870);
xor XOR2 (N2665, N2663, N1774);
or OR4 (N2666, N2651, N2327, N384, N1694);
nand NAND3 (N2667, N2662, N1747, N1742);
buf BUF1 (N2668, N2665);
buf BUF1 (N2669, N2666);
xor XOR2 (N2670, N2667, N2252);
or OR2 (N2671, N2670, N577);
nor NOR2 (N2672, N2671, N1903);
xor XOR2 (N2673, N2655, N745);
not NOT1 (N2674, N2669);
buf BUF1 (N2675, N2640);
xor XOR2 (N2676, N2658, N2157);
nor NOR4 (N2677, N2660, N794, N1538, N2294);
not NOT1 (N2678, N2661);
and AND2 (N2679, N2675, N1314);
xor XOR2 (N2680, N2633, N202);
and AND4 (N2681, N2673, N1186, N741, N1249);
buf BUF1 (N2682, N2672);
not NOT1 (N2683, N2664);
and AND3 (N2684, N2682, N2362, N1354);
buf BUF1 (N2685, N2680);
or OR3 (N2686, N2676, N2551, N1319);
nor NOR2 (N2687, N2681, N1306);
or OR4 (N2688, N2683, N2559, N2188, N2203);
not NOT1 (N2689, N2678);
nor NOR2 (N2690, N2687, N1841);
buf BUF1 (N2691, N2690);
nor NOR2 (N2692, N2686, N1587);
not NOT1 (N2693, N2668);
nand NAND3 (N2694, N2692, N1323, N2024);
not NOT1 (N2695, N2694);
or OR2 (N2696, N2688, N1411);
nand NAND4 (N2697, N2691, N1991, N1273, N2692);
xor XOR2 (N2698, N2689, N316);
and AND4 (N2699, N2685, N2644, N1300, N2194);
buf BUF1 (N2700, N2697);
nor NOR2 (N2701, N2696, N2520);
not NOT1 (N2702, N2679);
nor NOR2 (N2703, N2677, N1544);
nor NOR2 (N2704, N2684, N1673);
nand NAND3 (N2705, N2699, N2206, N2596);
not NOT1 (N2706, N2693);
buf BUF1 (N2707, N2703);
nand NAND3 (N2708, N2705, N1904, N1264);
nand NAND2 (N2709, N2674, N738);
not NOT1 (N2710, N2706);
and AND3 (N2711, N2708, N1917, N2160);
or OR2 (N2712, N2707, N1134);
not NOT1 (N2713, N2695);
nor NOR3 (N2714, N2698, N2698, N814);
nor NOR3 (N2715, N2704, N1786, N1687);
buf BUF1 (N2716, N2710);
nand NAND3 (N2717, N2709, N2555, N164);
nand NAND3 (N2718, N2716, N862, N1411);
nand NAND3 (N2719, N2711, N2199, N895);
nor NOR3 (N2720, N2714, N383, N2232);
or OR3 (N2721, N2715, N271, N1340);
buf BUF1 (N2722, N2717);
not NOT1 (N2723, N2701);
or OR4 (N2724, N2719, N932, N2279, N1159);
or OR3 (N2725, N2723, N273, N1740);
or OR4 (N2726, N2712, N329, N1507, N505);
or OR2 (N2727, N2722, N1256);
not NOT1 (N2728, N2725);
and AND4 (N2729, N2724, N1807, N714, N2364);
nor NOR2 (N2730, N2713, N2562);
nor NOR4 (N2731, N2700, N1534, N2636, N28);
or OR4 (N2732, N2729, N350, N1576, N2423);
or OR3 (N2733, N2731, N50, N1842);
xor XOR2 (N2734, N2702, N1232);
xor XOR2 (N2735, N2732, N461);
xor XOR2 (N2736, N2718, N2709);
or OR3 (N2737, N2728, N1842, N2016);
and AND2 (N2738, N2726, N1808);
nor NOR2 (N2739, N2733, N2519);
xor XOR2 (N2740, N2736, N695);
xor XOR2 (N2741, N2735, N1082);
not NOT1 (N2742, N2734);
buf BUF1 (N2743, N2741);
nand NAND3 (N2744, N2730, N1406, N419);
nand NAND4 (N2745, N2738, N559, N555, N739);
nand NAND4 (N2746, N2721, N984, N2271, N2123);
xor XOR2 (N2747, N2744, N1438);
nor NOR4 (N2748, N2727, N2206, N794, N1557);
nor NOR2 (N2749, N2747, N1957);
or OR3 (N2750, N2748, N161, N972);
nor NOR4 (N2751, N2743, N1070, N1858, N1921);
nor NOR2 (N2752, N2751, N1320);
nand NAND2 (N2753, N2752, N905);
buf BUF1 (N2754, N2739);
and AND3 (N2755, N2746, N2638, N344);
or OR3 (N2756, N2755, N1344, N1826);
nand NAND3 (N2757, N2754, N570, N1439);
or OR3 (N2758, N2740, N2275, N2677);
and AND3 (N2759, N2750, N137, N10);
and AND4 (N2760, N2756, N1439, N2483, N1253);
nor NOR4 (N2761, N2760, N2040, N1539, N1529);
and AND2 (N2762, N2745, N2101);
nor NOR3 (N2763, N2720, N1457, N1384);
buf BUF1 (N2764, N2757);
and AND4 (N2765, N2758, N42, N873, N521);
xor XOR2 (N2766, N2753, N1665);
or OR4 (N2767, N2761, N2164, N2750, N1407);
xor XOR2 (N2768, N2737, N2652);
and AND2 (N2769, N2768, N1830);
xor XOR2 (N2770, N2742, N2);
nor NOR2 (N2771, N2770, N1381);
buf BUF1 (N2772, N2765);
or OR4 (N2773, N2764, N727, N673, N368);
xor XOR2 (N2774, N2769, N2756);
and AND3 (N2775, N2763, N480, N439);
nand NAND4 (N2776, N2775, N67, N2687, N2069);
buf BUF1 (N2777, N2762);
or OR4 (N2778, N2749, N2542, N2618, N2228);
nor NOR2 (N2779, N2778, N358);
nor NOR3 (N2780, N2759, N910, N35);
buf BUF1 (N2781, N2777);
or OR2 (N2782, N2776, N2047);
nor NOR2 (N2783, N2781, N949);
and AND4 (N2784, N2783, N428, N706, N1480);
or OR2 (N2785, N2773, N752);
nor NOR2 (N2786, N2785, N2524);
buf BUF1 (N2787, N2780);
xor XOR2 (N2788, N2782, N126);
xor XOR2 (N2789, N2774, N1744);
buf BUF1 (N2790, N2787);
buf BUF1 (N2791, N2766);
and AND2 (N2792, N2791, N2373);
nand NAND4 (N2793, N2790, N870, N629, N2117);
buf BUF1 (N2794, N2784);
and AND3 (N2795, N2794, N835, N2278);
nand NAND3 (N2796, N2772, N798, N916);
and AND3 (N2797, N2792, N1197, N1222);
nand NAND4 (N2798, N2793, N2150, N1108, N808);
nand NAND3 (N2799, N2779, N847, N1706);
xor XOR2 (N2800, N2786, N1373);
not NOT1 (N2801, N2788);
buf BUF1 (N2802, N2795);
or OR2 (N2803, N2798, N2621);
nand NAND2 (N2804, N2800, N656);
buf BUF1 (N2805, N2771);
xor XOR2 (N2806, N2805, N683);
or OR4 (N2807, N2802, N1663, N1476, N2105);
or OR2 (N2808, N2797, N2508);
not NOT1 (N2809, N2808);
not NOT1 (N2810, N2801);
and AND3 (N2811, N2804, N1713, N1760);
nand NAND2 (N2812, N2789, N1648);
xor XOR2 (N2813, N2807, N963);
xor XOR2 (N2814, N2813, N704);
or OR2 (N2815, N2803, N490);
nand NAND4 (N2816, N2812, N1532, N1246, N484);
xor XOR2 (N2817, N2814, N2395);
xor XOR2 (N2818, N2817, N794);
not NOT1 (N2819, N2767);
and AND4 (N2820, N2811, N1485, N47, N1124);
nand NAND2 (N2821, N2809, N903);
buf BUF1 (N2822, N2816);
not NOT1 (N2823, N2796);
nor NOR3 (N2824, N2799, N1821, N1183);
xor XOR2 (N2825, N2822, N2044);
not NOT1 (N2826, N2818);
and AND4 (N2827, N2819, N1671, N751, N2319);
xor XOR2 (N2828, N2806, N2643);
not NOT1 (N2829, N2824);
xor XOR2 (N2830, N2828, N1713);
and AND4 (N2831, N2821, N2012, N1536, N1702);
not NOT1 (N2832, N2810);
buf BUF1 (N2833, N2831);
not NOT1 (N2834, N2823);
or OR3 (N2835, N2825, N1240, N909);
not NOT1 (N2836, N2827);
or OR3 (N2837, N2815, N1282, N733);
not NOT1 (N2838, N2837);
nor NOR2 (N2839, N2826, N2639);
nor NOR2 (N2840, N2833, N1953);
buf BUF1 (N2841, N2820);
nand NAND2 (N2842, N2841, N1906);
buf BUF1 (N2843, N2834);
or OR4 (N2844, N2843, N2426, N777, N302);
nor NOR3 (N2845, N2835, N229, N2077);
buf BUF1 (N2846, N2840);
nor NOR2 (N2847, N2838, N1177);
and AND4 (N2848, N2846, N1571, N1429, N1676);
nand NAND4 (N2849, N2845, N448, N1314, N66);
and AND4 (N2850, N2830, N1911, N409, N2516);
and AND2 (N2851, N2832, N1945);
nand NAND2 (N2852, N2829, N2261);
xor XOR2 (N2853, N2839, N1732);
not NOT1 (N2854, N2836);
not NOT1 (N2855, N2854);
nand NAND2 (N2856, N2842, N1310);
buf BUF1 (N2857, N2844);
buf BUF1 (N2858, N2848);
or OR3 (N2859, N2857, N1779, N1672);
not NOT1 (N2860, N2858);
xor XOR2 (N2861, N2847, N752);
and AND3 (N2862, N2856, N521, N2189);
and AND3 (N2863, N2850, N2664, N2282);
nand NAND4 (N2864, N2849, N886, N905, N574);
buf BUF1 (N2865, N2860);
buf BUF1 (N2866, N2853);
nand NAND2 (N2867, N2865, N1497);
not NOT1 (N2868, N2863);
not NOT1 (N2869, N2864);
buf BUF1 (N2870, N2868);
nand NAND4 (N2871, N2862, N115, N1327, N468);
buf BUF1 (N2872, N2861);
xor XOR2 (N2873, N2851, N692);
or OR3 (N2874, N2866, N764, N422);
buf BUF1 (N2875, N2859);
nor NOR4 (N2876, N2867, N1687, N1180, N1681);
buf BUF1 (N2877, N2855);
and AND3 (N2878, N2852, N1170, N9);
buf BUF1 (N2879, N2874);
not NOT1 (N2880, N2872);
not NOT1 (N2881, N2879);
xor XOR2 (N2882, N2877, N980);
nor NOR2 (N2883, N2880, N2262);
nand NAND4 (N2884, N2883, N629, N2138, N925);
not NOT1 (N2885, N2881);
and AND2 (N2886, N2871, N348);
not NOT1 (N2887, N2870);
nor NOR3 (N2888, N2884, N1878, N647);
xor XOR2 (N2889, N2882, N2498);
nor NOR2 (N2890, N2887, N702);
nor NOR3 (N2891, N2869, N2628, N2724);
xor XOR2 (N2892, N2873, N1040);
nand NAND2 (N2893, N2886, N2475);
buf BUF1 (N2894, N2893);
or OR3 (N2895, N2875, N1988, N1106);
buf BUF1 (N2896, N2891);
nor NOR4 (N2897, N2885, N1383, N1377, N632);
buf BUF1 (N2898, N2890);
nor NOR2 (N2899, N2889, N1101);
nand NAND4 (N2900, N2878, N1497, N376, N2517);
and AND4 (N2901, N2892, N1099, N583, N2844);
not NOT1 (N2902, N2876);
or OR3 (N2903, N2902, N1449, N2529);
xor XOR2 (N2904, N2894, N307);
xor XOR2 (N2905, N2899, N2209);
nand NAND2 (N2906, N2888, N280);
or OR4 (N2907, N2901, N301, N2393, N505);
not NOT1 (N2908, N2907);
buf BUF1 (N2909, N2898);
nor NOR3 (N2910, N2906, N857, N1868);
nand NAND4 (N2911, N2896, N2160, N2889, N2046);
buf BUF1 (N2912, N2904);
and AND3 (N2913, N2908, N2667, N2040);
and AND3 (N2914, N2903, N2831, N1391);
buf BUF1 (N2915, N2911);
and AND4 (N2916, N2909, N2398, N855, N679);
nand NAND4 (N2917, N2914, N31, N663, N2780);
buf BUF1 (N2918, N2905);
nor NOR4 (N2919, N2897, N2885, N469, N1179);
not NOT1 (N2920, N2900);
not NOT1 (N2921, N2918);
and AND4 (N2922, N2919, N2511, N2324, N355);
nand NAND2 (N2923, N2922, N2377);
and AND4 (N2924, N2921, N2614, N1296, N1696);
xor XOR2 (N2925, N2917, N1974);
nand NAND2 (N2926, N2910, N1917);
buf BUF1 (N2927, N2925);
and AND4 (N2928, N2916, N2163, N934, N2403);
or OR4 (N2929, N2913, N2342, N1634, N1557);
or OR4 (N2930, N2927, N2388, N574, N1904);
buf BUF1 (N2931, N2924);
not NOT1 (N2932, N2928);
nand NAND2 (N2933, N2915, N395);
nand NAND4 (N2934, N2931, N832, N977, N184);
and AND3 (N2935, N2934, N2910, N573);
xor XOR2 (N2936, N2929, N2371);
not NOT1 (N2937, N2895);
and AND2 (N2938, N2912, N1963);
nand NAND2 (N2939, N2920, N308);
or OR3 (N2940, N2926, N2819, N2186);
and AND3 (N2941, N2940, N769, N1004);
not NOT1 (N2942, N2933);
nor NOR2 (N2943, N2937, N2014);
nand NAND4 (N2944, N2939, N1371, N401, N2313);
nor NOR3 (N2945, N2942, N2589, N2609);
nor NOR3 (N2946, N2943, N2741, N1363);
xor XOR2 (N2947, N2944, N142);
and AND3 (N2948, N2941, N241, N1235);
nand NAND4 (N2949, N2938, N1776, N492, N77);
buf BUF1 (N2950, N2947);
xor XOR2 (N2951, N2935, N2124);
nor NOR2 (N2952, N2936, N1253);
xor XOR2 (N2953, N2923, N2575);
or OR4 (N2954, N2946, N1527, N1907, N1181);
not NOT1 (N2955, N2949);
nand NAND3 (N2956, N2952, N603, N2921);
nor NOR4 (N2957, N2951, N2844, N46, N1135);
nand NAND3 (N2958, N2948, N2088, N128);
xor XOR2 (N2959, N2930, N2937);
xor XOR2 (N2960, N2956, N1284);
not NOT1 (N2961, N2954);
buf BUF1 (N2962, N2950);
nor NOR2 (N2963, N2961, N154);
or OR2 (N2964, N2932, N818);
buf BUF1 (N2965, N2960);
xor XOR2 (N2966, N2959, N1112);
xor XOR2 (N2967, N2945, N2177);
not NOT1 (N2968, N2955);
not NOT1 (N2969, N2958);
xor XOR2 (N2970, N2963, N1442);
nor NOR2 (N2971, N2962, N2794);
nor NOR3 (N2972, N2957, N314, N930);
not NOT1 (N2973, N2965);
and AND2 (N2974, N2968, N1488);
xor XOR2 (N2975, N2967, N475);
not NOT1 (N2976, N2972);
nand NAND2 (N2977, N2973, N1340);
and AND3 (N2978, N2975, N615, N1906);
buf BUF1 (N2979, N2953);
and AND4 (N2980, N2964, N1779, N2658, N1881);
and AND3 (N2981, N2977, N694, N1779);
nor NOR4 (N2982, N2976, N2857, N1928, N1815);
not NOT1 (N2983, N2978);
nor NOR4 (N2984, N2982, N661, N1302, N1865);
xor XOR2 (N2985, N2984, N392);
or OR4 (N2986, N2980, N2681, N1344, N2265);
nand NAND3 (N2987, N2969, N2229, N1145);
not NOT1 (N2988, N2971);
buf BUF1 (N2989, N2979);
not NOT1 (N2990, N2988);
nor NOR3 (N2991, N2985, N896, N602);
buf BUF1 (N2992, N2974);
nor NOR4 (N2993, N2986, N2021, N1873, N781);
not NOT1 (N2994, N2989);
xor XOR2 (N2995, N2983, N2948);
buf BUF1 (N2996, N2966);
nor NOR3 (N2997, N2994, N2008, N559);
nand NAND3 (N2998, N2970, N598, N2736);
nor NOR4 (N2999, N2998, N1363, N1677, N939);
and AND4 (N3000, N2995, N1637, N2372, N138);
and AND3 (N3001, N2991, N2784, N1979);
and AND3 (N3002, N2993, N49, N948);
buf BUF1 (N3003, N2996);
nor NOR2 (N3004, N3003, N306);
xor XOR2 (N3005, N3000, N1691);
xor XOR2 (N3006, N3005, N1311);
nor NOR3 (N3007, N2999, N1404, N2768);
not NOT1 (N3008, N3006);
xor XOR2 (N3009, N3004, N989);
xor XOR2 (N3010, N3007, N2130);
or OR3 (N3011, N3008, N2218, N54);
xor XOR2 (N3012, N2992, N2166);
xor XOR2 (N3013, N3001, N1858);
nor NOR3 (N3014, N3009, N2827, N2633);
endmodule