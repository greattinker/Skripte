// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19;

output N2510,N2516,N2511,N2518,N2513,N2508,N2506,N2514,N2505,N2519;

buf BUF1 (N20, N13);
or OR3 (N21, N11, N13, N7);
nor NOR3 (N22, N1, N7, N4);
buf BUF1 (N23, N14);
nand NAND2 (N24, N16, N15);
nand NAND3 (N25, N1, N6, N4);
nand NAND4 (N26, N24, N7, N5, N3);
nor NOR4 (N27, N25, N3, N4, N4);
or OR2 (N28, N18, N11);
nor NOR4 (N29, N18, N9, N11, N11);
buf BUF1 (N30, N11);
buf BUF1 (N31, N27);
nand NAND3 (N32, N12, N8, N14);
or OR3 (N33, N30, N13, N21);
nor NOR2 (N34, N8, N5);
buf BUF1 (N35, N22);
buf BUF1 (N36, N26);
not NOT1 (N37, N28);
or OR3 (N38, N37, N35, N14);
xor XOR2 (N39, N23, N22);
nor NOR2 (N40, N9, N8);
xor XOR2 (N41, N29, N13);
and AND3 (N42, N39, N11, N1);
or OR3 (N43, N32, N17, N21);
not NOT1 (N44, N43);
and AND4 (N45, N41, N39, N20, N17);
not NOT1 (N46, N19);
nor NOR2 (N47, N46, N19);
nand NAND4 (N48, N42, N5, N40, N16);
nand NAND2 (N49, N44, N41);
nor NOR2 (N50, N18, N17);
not NOT1 (N51, N34);
nand NAND3 (N52, N38, N28, N3);
and AND2 (N53, N33, N44);
buf BUF1 (N54, N31);
nand NAND4 (N55, N45, N29, N44, N53);
and AND4 (N56, N44, N49, N27, N3);
not NOT1 (N57, N47);
or OR2 (N58, N5, N10);
nor NOR3 (N59, N48, N30, N51);
nand NAND3 (N60, N5, N2, N51);
and AND2 (N61, N55, N19);
xor XOR2 (N62, N54, N6);
or OR3 (N63, N36, N8, N21);
not NOT1 (N64, N50);
buf BUF1 (N65, N52);
nand NAND3 (N66, N62, N13, N24);
nor NOR4 (N67, N66, N3, N36, N32);
xor XOR2 (N68, N60, N20);
nor NOR4 (N69, N56, N42, N68, N57);
or OR3 (N70, N18, N48, N57);
and AND4 (N71, N53, N64, N9, N63);
nand NAND2 (N72, N10, N11);
xor XOR2 (N73, N13, N27);
xor XOR2 (N74, N69, N26);
nand NAND4 (N75, N67, N44, N68, N10);
not NOT1 (N76, N59);
nor NOR3 (N77, N71, N74, N66);
xor XOR2 (N78, N7, N27);
not NOT1 (N79, N61);
nand NAND4 (N80, N73, N38, N24, N36);
buf BUF1 (N81, N70);
buf BUF1 (N82, N81);
and AND3 (N83, N79, N14, N13);
nand NAND2 (N84, N80, N59);
not NOT1 (N85, N72);
xor XOR2 (N86, N65, N33);
xor XOR2 (N87, N78, N85);
nor NOR4 (N88, N37, N52, N76, N71);
or OR3 (N89, N23, N51, N64);
and AND4 (N90, N82, N88, N7, N49);
buf BUF1 (N91, N33);
xor XOR2 (N92, N75, N2);
not NOT1 (N93, N92);
buf BUF1 (N94, N90);
buf BUF1 (N95, N83);
not NOT1 (N96, N95);
xor XOR2 (N97, N84, N81);
and AND4 (N98, N94, N94, N55, N74);
buf BUF1 (N99, N89);
nand NAND4 (N100, N77, N43, N6, N18);
xor XOR2 (N101, N58, N68);
nand NAND2 (N102, N98, N61);
or OR3 (N103, N99, N54, N44);
or OR3 (N104, N101, N77, N87);
and AND4 (N105, N72, N87, N101, N51);
nor NOR3 (N106, N102, N100, N88);
or OR2 (N107, N80, N17);
and AND3 (N108, N104, N69, N8);
and AND3 (N109, N105, N46, N55);
nor NOR4 (N110, N91, N72, N10, N20);
not NOT1 (N111, N93);
nand NAND2 (N112, N111, N70);
not NOT1 (N113, N106);
nand NAND2 (N114, N113, N60);
xor XOR2 (N115, N114, N28);
xor XOR2 (N116, N108, N107);
not NOT1 (N117, N19);
nor NOR3 (N118, N110, N6, N65);
nand NAND3 (N119, N109, N92, N37);
buf BUF1 (N120, N115);
not NOT1 (N121, N117);
buf BUF1 (N122, N97);
buf BUF1 (N123, N86);
xor XOR2 (N124, N120, N115);
nand NAND2 (N125, N116, N82);
nand NAND2 (N126, N96, N54);
nand NAND2 (N127, N124, N19);
nand NAND2 (N128, N118, N116);
and AND2 (N129, N122, N97);
or OR4 (N130, N127, N49, N93, N129);
or OR2 (N131, N121, N118);
buf BUF1 (N132, N70);
nand NAND2 (N133, N123, N88);
nand NAND2 (N134, N103, N26);
not NOT1 (N135, N119);
and AND3 (N136, N126, N6, N120);
xor XOR2 (N137, N133, N39);
nand NAND3 (N138, N137, N120, N9);
nor NOR4 (N139, N136, N30, N42, N45);
and AND4 (N140, N135, N117, N40, N94);
xor XOR2 (N141, N131, N80);
nand NAND4 (N142, N125, N123, N11, N130);
or OR4 (N143, N74, N3, N93, N21);
xor XOR2 (N144, N143, N60);
or OR3 (N145, N144, N64, N9);
not NOT1 (N146, N132);
buf BUF1 (N147, N128);
nand NAND3 (N148, N141, N112, N43);
nand NAND3 (N149, N25, N79, N71);
nor NOR2 (N150, N138, N32);
nand NAND4 (N151, N139, N76, N148, N136);
nor NOR2 (N152, N35, N4);
or OR4 (N153, N152, N114, N136, N150);
nand NAND3 (N154, N61, N73, N52);
not NOT1 (N155, N154);
nor NOR2 (N156, N146, N137);
not NOT1 (N157, N134);
nand NAND2 (N158, N153, N23);
xor XOR2 (N159, N158, N79);
nand NAND2 (N160, N149, N79);
buf BUF1 (N161, N156);
not NOT1 (N162, N161);
not NOT1 (N163, N157);
buf BUF1 (N164, N162);
not NOT1 (N165, N164);
xor XOR2 (N166, N155, N70);
not NOT1 (N167, N159);
not NOT1 (N168, N145);
nor NOR2 (N169, N165, N14);
and AND3 (N170, N142, N64, N147);
buf BUF1 (N171, N31);
xor XOR2 (N172, N140, N30);
not NOT1 (N173, N172);
xor XOR2 (N174, N163, N62);
xor XOR2 (N175, N151, N129);
and AND4 (N176, N160, N34, N23, N7);
or OR4 (N177, N170, N45, N69, N12);
nor NOR2 (N178, N177, N136);
not NOT1 (N179, N167);
not NOT1 (N180, N176);
buf BUF1 (N181, N180);
and AND2 (N182, N181, N7);
xor XOR2 (N183, N171, N139);
and AND3 (N184, N169, N181, N136);
not NOT1 (N185, N184);
not NOT1 (N186, N182);
xor XOR2 (N187, N185, N60);
nand NAND4 (N188, N166, N175, N121, N43);
nand NAND4 (N189, N86, N127, N83, N153);
and AND4 (N190, N183, N63, N155, N56);
xor XOR2 (N191, N168, N190);
buf BUF1 (N192, N10);
xor XOR2 (N193, N179, N140);
nand NAND2 (N194, N187, N136);
buf BUF1 (N195, N191);
and AND3 (N196, N178, N124, N140);
nand NAND4 (N197, N188, N27, N28, N52);
or OR4 (N198, N186, N148, N68, N108);
nor NOR2 (N199, N195, N62);
not NOT1 (N200, N173);
or OR3 (N201, N193, N25, N109);
nor NOR2 (N202, N197, N54);
and AND2 (N203, N194, N3);
xor XOR2 (N204, N200, N148);
buf BUF1 (N205, N196);
not NOT1 (N206, N192);
or OR4 (N207, N201, N204, N116, N109);
nand NAND4 (N208, N178, N15, N18, N144);
xor XOR2 (N209, N202, N38);
nor NOR4 (N210, N199, N34, N73, N65);
nand NAND4 (N211, N189, N123, N82, N168);
and AND2 (N212, N174, N68);
xor XOR2 (N213, N210, N83);
or OR4 (N214, N207, N121, N15, N99);
nand NAND3 (N215, N203, N174, N176);
or OR4 (N216, N212, N121, N38, N138);
nor NOR3 (N217, N215, N156, N19);
xor XOR2 (N218, N198, N153);
or OR2 (N219, N211, N55);
nand NAND4 (N220, N217, N6, N218, N7);
or OR2 (N221, N212, N203);
xor XOR2 (N222, N208, N14);
buf BUF1 (N223, N222);
buf BUF1 (N224, N223);
nand NAND3 (N225, N216, N196, N61);
nor NOR2 (N226, N214, N31);
not NOT1 (N227, N209);
or OR4 (N228, N221, N211, N59, N140);
nand NAND3 (N229, N226, N82, N161);
nor NOR3 (N230, N227, N188, N88);
nor NOR4 (N231, N230, N98, N13, N204);
and AND3 (N232, N219, N135, N107);
or OR4 (N233, N205, N209, N217, N88);
and AND3 (N234, N224, N166, N68);
nor NOR2 (N235, N213, N89);
not NOT1 (N236, N231);
and AND2 (N237, N225, N184);
nand NAND2 (N238, N220, N113);
not NOT1 (N239, N206);
nand NAND2 (N240, N238, N194);
buf BUF1 (N241, N234);
nor NOR4 (N242, N237, N24, N10, N68);
nor NOR2 (N243, N239, N173);
or OR2 (N244, N228, N90);
nand NAND4 (N245, N241, N73, N23, N201);
buf BUF1 (N246, N242);
nor NOR4 (N247, N233, N132, N180, N121);
nand NAND3 (N248, N243, N16, N121);
not NOT1 (N249, N246);
not NOT1 (N250, N244);
buf BUF1 (N251, N250);
nand NAND3 (N252, N240, N105, N10);
not NOT1 (N253, N245);
buf BUF1 (N254, N247);
nor NOR3 (N255, N236, N5, N177);
xor XOR2 (N256, N235, N249);
or OR4 (N257, N27, N163, N29, N23);
nor NOR2 (N258, N254, N34);
nand NAND4 (N259, N257, N33, N23, N79);
not NOT1 (N260, N229);
not NOT1 (N261, N255);
xor XOR2 (N262, N248, N80);
nor NOR2 (N263, N251, N91);
xor XOR2 (N264, N259, N101);
nand NAND4 (N265, N262, N212, N258, N141);
xor XOR2 (N266, N164, N33);
and AND3 (N267, N260, N199, N16);
and AND3 (N268, N253, N5, N51);
xor XOR2 (N269, N264, N154);
nand NAND2 (N270, N266, N173);
buf BUF1 (N271, N268);
or OR3 (N272, N256, N60, N155);
nor NOR3 (N273, N265, N188, N265);
nor NOR2 (N274, N270, N166);
nor NOR4 (N275, N252, N157, N233, N245);
nand NAND3 (N276, N274, N85, N22);
buf BUF1 (N277, N273);
not NOT1 (N278, N272);
buf BUF1 (N279, N261);
or OR3 (N280, N267, N33, N154);
buf BUF1 (N281, N278);
nor NOR2 (N282, N277, N165);
xor XOR2 (N283, N281, N198);
xor XOR2 (N284, N282, N135);
not NOT1 (N285, N275);
or OR3 (N286, N279, N271, N154);
and AND4 (N287, N167, N29, N198, N68);
and AND3 (N288, N283, N244, N250);
nor NOR2 (N289, N287, N140);
or OR3 (N290, N232, N6, N60);
or OR3 (N291, N263, N257, N111);
nor NOR2 (N292, N288, N71);
not NOT1 (N293, N276);
or OR2 (N294, N292, N18);
xor XOR2 (N295, N291, N29);
and AND3 (N296, N285, N130, N43);
and AND2 (N297, N269, N105);
or OR3 (N298, N290, N84, N273);
xor XOR2 (N299, N284, N187);
nand NAND3 (N300, N298, N140, N144);
nor NOR2 (N301, N293, N266);
buf BUF1 (N302, N297);
nand NAND2 (N303, N301, N216);
xor XOR2 (N304, N303, N146);
not NOT1 (N305, N289);
xor XOR2 (N306, N305, N208);
or OR4 (N307, N294, N44, N18, N293);
or OR4 (N308, N304, N10, N269, N127);
xor XOR2 (N309, N296, N304);
xor XOR2 (N310, N300, N51);
buf BUF1 (N311, N308);
or OR4 (N312, N307, N302, N176, N240);
buf BUF1 (N313, N216);
and AND4 (N314, N310, N51, N25, N147);
xor XOR2 (N315, N309, N155);
and AND4 (N316, N314, N309, N87, N199);
nand NAND2 (N317, N316, N170);
buf BUF1 (N318, N280);
not NOT1 (N319, N299);
xor XOR2 (N320, N311, N241);
nor NOR4 (N321, N318, N92, N274, N275);
buf BUF1 (N322, N312);
nor NOR2 (N323, N315, N110);
and AND4 (N324, N321, N115, N48, N188);
buf BUF1 (N325, N286);
not NOT1 (N326, N324);
not NOT1 (N327, N326);
or OR2 (N328, N317, N327);
nand NAND2 (N329, N277, N108);
and AND4 (N330, N322, N75, N205, N45);
nor NOR4 (N331, N319, N236, N10, N319);
not NOT1 (N332, N323);
and AND2 (N333, N332, N168);
and AND2 (N334, N306, N140);
nor NOR4 (N335, N330, N77, N71, N177);
nor NOR2 (N336, N313, N176);
xor XOR2 (N337, N295, N276);
and AND2 (N338, N331, N294);
and AND2 (N339, N328, N91);
xor XOR2 (N340, N335, N29);
buf BUF1 (N341, N333);
nor NOR2 (N342, N320, N59);
buf BUF1 (N343, N339);
buf BUF1 (N344, N337);
nand NAND2 (N345, N329, N283);
nand NAND3 (N346, N341, N104, N277);
nor NOR3 (N347, N346, N58, N224);
and AND3 (N348, N325, N7, N132);
nand NAND4 (N349, N344, N298, N86, N131);
buf BUF1 (N350, N349);
nor NOR3 (N351, N348, N75, N317);
and AND3 (N352, N343, N243, N318);
nor NOR4 (N353, N345, N343, N157, N178);
nand NAND4 (N354, N351, N210, N14, N64);
nand NAND4 (N355, N353, N300, N190, N76);
not NOT1 (N356, N347);
nor NOR2 (N357, N342, N253);
not NOT1 (N358, N352);
and AND3 (N359, N336, N19, N303);
xor XOR2 (N360, N350, N290);
or OR2 (N361, N359, N227);
xor XOR2 (N362, N340, N11);
buf BUF1 (N363, N338);
and AND2 (N364, N361, N74);
not NOT1 (N365, N363);
and AND4 (N366, N356, N280, N227, N83);
or OR3 (N367, N366, N347, N343);
or OR2 (N368, N364, N128);
nand NAND4 (N369, N367, N176, N234, N100);
xor XOR2 (N370, N355, N36);
nand NAND2 (N371, N368, N218);
or OR3 (N372, N371, N229, N214);
nand NAND3 (N373, N354, N349, N245);
or OR4 (N374, N370, N372, N172, N87);
nand NAND4 (N375, N339, N243, N360, N204);
buf BUF1 (N376, N271);
nand NAND2 (N377, N374, N312);
buf BUF1 (N378, N377);
or OR4 (N379, N334, N296, N84, N213);
xor XOR2 (N380, N373, N36);
buf BUF1 (N381, N369);
or OR3 (N382, N378, N326, N126);
buf BUF1 (N383, N357);
nor NOR4 (N384, N375, N266, N73, N116);
nand NAND3 (N385, N380, N29, N378);
nor NOR3 (N386, N362, N17, N161);
nor NOR3 (N387, N358, N348, N177);
nand NAND3 (N388, N382, N262, N20);
nand NAND4 (N389, N388, N135, N184, N316);
not NOT1 (N390, N389);
buf BUF1 (N391, N381);
nor NOR3 (N392, N384, N76, N123);
buf BUF1 (N393, N386);
xor XOR2 (N394, N383, N287);
and AND3 (N395, N385, N106, N232);
xor XOR2 (N396, N391, N200);
or OR2 (N397, N376, N118);
nor NOR3 (N398, N396, N233, N54);
or OR4 (N399, N397, N362, N155, N230);
or OR3 (N400, N390, N188, N273);
not NOT1 (N401, N395);
xor XOR2 (N402, N365, N98);
or OR2 (N403, N398, N332);
nor NOR4 (N404, N403, N39, N375, N27);
nand NAND2 (N405, N379, N150);
or OR4 (N406, N399, N13, N302, N24);
nor NOR4 (N407, N402, N162, N89, N47);
or OR3 (N408, N394, N191, N104);
and AND2 (N409, N393, N96);
buf BUF1 (N410, N405);
not NOT1 (N411, N392);
nand NAND4 (N412, N401, N278, N317, N298);
not NOT1 (N413, N387);
or OR3 (N414, N411, N348, N405);
or OR4 (N415, N404, N89, N371, N130);
nor NOR3 (N416, N400, N293, N93);
nand NAND3 (N417, N410, N215, N226);
xor XOR2 (N418, N408, N52);
nand NAND4 (N419, N413, N63, N328, N29);
and AND4 (N420, N414, N346, N92, N90);
nand NAND3 (N421, N419, N294, N179);
nor NOR2 (N422, N409, N157);
buf BUF1 (N423, N406);
xor XOR2 (N424, N421, N171);
nor NOR3 (N425, N407, N40, N109);
and AND4 (N426, N423, N32, N106, N84);
or OR3 (N427, N425, N17, N208);
nor NOR3 (N428, N416, N359, N62);
xor XOR2 (N429, N422, N227);
xor XOR2 (N430, N429, N7);
buf BUF1 (N431, N426);
not NOT1 (N432, N412);
nand NAND4 (N433, N427, N395, N276, N89);
not NOT1 (N434, N433);
not NOT1 (N435, N424);
xor XOR2 (N436, N428, N177);
and AND2 (N437, N435, N403);
xor XOR2 (N438, N436, N397);
xor XOR2 (N439, N420, N116);
xor XOR2 (N440, N439, N3);
nor NOR2 (N441, N434, N156);
or OR2 (N442, N431, N385);
buf BUF1 (N443, N417);
and AND2 (N444, N418, N185);
nand NAND3 (N445, N440, N435, N94);
buf BUF1 (N446, N437);
nand NAND2 (N447, N415, N191);
buf BUF1 (N448, N446);
or OR4 (N449, N430, N269, N393, N437);
xor XOR2 (N450, N441, N376);
or OR2 (N451, N443, N212);
nor NOR3 (N452, N447, N135, N26);
buf BUF1 (N453, N432);
and AND3 (N454, N445, N157, N239);
buf BUF1 (N455, N453);
or OR3 (N456, N452, N161, N226);
or OR2 (N457, N444, N67);
nand NAND4 (N458, N455, N440, N27, N236);
buf BUF1 (N459, N448);
xor XOR2 (N460, N442, N10);
or OR4 (N461, N458, N39, N288, N234);
and AND2 (N462, N438, N118);
nand NAND2 (N463, N451, N123);
xor XOR2 (N464, N457, N338);
not NOT1 (N465, N461);
not NOT1 (N466, N462);
nand NAND3 (N467, N456, N215, N305);
nand NAND3 (N468, N454, N38, N433);
nand NAND4 (N469, N463, N431, N252, N65);
nor NOR3 (N470, N469, N430, N212);
xor XOR2 (N471, N460, N455);
xor XOR2 (N472, N467, N200);
nand NAND4 (N473, N470, N160, N349, N424);
xor XOR2 (N474, N465, N304);
or OR3 (N475, N472, N41, N371);
xor XOR2 (N476, N449, N120);
and AND2 (N477, N474, N462);
not NOT1 (N478, N459);
nand NAND2 (N479, N450, N383);
xor XOR2 (N480, N475, N280);
nand NAND4 (N481, N476, N349, N454, N87);
not NOT1 (N482, N481);
xor XOR2 (N483, N471, N16);
and AND2 (N484, N473, N25);
nor NOR2 (N485, N484, N185);
not NOT1 (N486, N466);
and AND2 (N487, N485, N144);
buf BUF1 (N488, N483);
xor XOR2 (N489, N464, N59);
not NOT1 (N490, N488);
nor NOR3 (N491, N468, N291, N308);
and AND2 (N492, N477, N257);
and AND3 (N493, N480, N314, N286);
nand NAND4 (N494, N479, N346, N218, N486);
xor XOR2 (N495, N29, N89);
not NOT1 (N496, N478);
and AND3 (N497, N493, N150, N418);
buf BUF1 (N498, N490);
not NOT1 (N499, N491);
nor NOR4 (N500, N498, N168, N254, N29);
or OR4 (N501, N494, N62, N462, N193);
xor XOR2 (N502, N501, N429);
or OR4 (N503, N500, N390, N220, N92);
xor XOR2 (N504, N482, N481);
buf BUF1 (N505, N495);
not NOT1 (N506, N497);
or OR3 (N507, N504, N437, N230);
not NOT1 (N508, N505);
nor NOR2 (N509, N506, N178);
not NOT1 (N510, N492);
nor NOR4 (N511, N489, N100, N362, N29);
nor NOR4 (N512, N508, N172, N134, N464);
or OR2 (N513, N496, N227);
nor NOR3 (N514, N503, N268, N250);
buf BUF1 (N515, N487);
nand NAND4 (N516, N513, N400, N247, N54);
or OR2 (N517, N499, N73);
and AND2 (N518, N512, N497);
not NOT1 (N519, N511);
nor NOR2 (N520, N507, N372);
nor NOR3 (N521, N516, N132, N197);
nor NOR2 (N522, N515, N249);
and AND2 (N523, N502, N463);
buf BUF1 (N524, N523);
nor NOR4 (N525, N510, N515, N434, N139);
and AND3 (N526, N519, N54, N192);
and AND3 (N527, N514, N321, N259);
xor XOR2 (N528, N521, N164);
not NOT1 (N529, N518);
xor XOR2 (N530, N509, N59);
or OR4 (N531, N522, N446, N108, N316);
nand NAND2 (N532, N527, N143);
not NOT1 (N533, N517);
or OR4 (N534, N529, N432, N272, N419);
or OR2 (N535, N525, N411);
and AND2 (N536, N532, N225);
buf BUF1 (N537, N528);
not NOT1 (N538, N533);
not NOT1 (N539, N526);
nor NOR3 (N540, N538, N271, N143);
xor XOR2 (N541, N531, N72);
xor XOR2 (N542, N539, N441);
xor XOR2 (N543, N534, N428);
buf BUF1 (N544, N530);
nand NAND4 (N545, N524, N59, N196, N257);
nand NAND2 (N546, N536, N535);
and AND4 (N547, N360, N164, N502, N212);
xor XOR2 (N548, N541, N185);
nor NOR4 (N549, N542, N181, N101, N126);
xor XOR2 (N550, N545, N300);
or OR3 (N551, N546, N27, N52);
nand NAND2 (N552, N544, N259);
or OR3 (N553, N520, N226, N148);
or OR2 (N554, N550, N225);
xor XOR2 (N555, N554, N496);
xor XOR2 (N556, N549, N500);
buf BUF1 (N557, N555);
xor XOR2 (N558, N543, N303);
nor NOR3 (N559, N553, N203, N156);
or OR2 (N560, N537, N557);
or OR4 (N561, N34, N424, N299, N121);
nand NAND2 (N562, N548, N363);
xor XOR2 (N563, N556, N298);
buf BUF1 (N564, N563);
and AND2 (N565, N540, N137);
nand NAND2 (N566, N562, N54);
nand NAND3 (N567, N551, N88, N555);
nor NOR2 (N568, N561, N150);
nor NOR2 (N569, N565, N263);
buf BUF1 (N570, N564);
nor NOR3 (N571, N552, N260, N432);
or OR3 (N572, N570, N381, N26);
xor XOR2 (N573, N571, N178);
and AND3 (N574, N568, N541, N245);
nand NAND2 (N575, N566, N496);
not NOT1 (N576, N567);
and AND2 (N577, N569, N509);
xor XOR2 (N578, N576, N13);
or OR4 (N579, N547, N137, N190, N565);
or OR2 (N580, N558, N217);
nor NOR3 (N581, N578, N320, N346);
not NOT1 (N582, N560);
nor NOR2 (N583, N577, N436);
and AND3 (N584, N574, N373, N103);
and AND3 (N585, N583, N326, N497);
not NOT1 (N586, N573);
xor XOR2 (N587, N581, N249);
or OR4 (N588, N586, N488, N214, N141);
buf BUF1 (N589, N575);
xor XOR2 (N590, N579, N188);
or OR3 (N591, N584, N280, N359);
nor NOR4 (N592, N587, N117, N578, N282);
and AND4 (N593, N591, N265, N2, N78);
buf BUF1 (N594, N588);
or OR2 (N595, N590, N216);
not NOT1 (N596, N594);
xor XOR2 (N597, N572, N269);
xor XOR2 (N598, N580, N566);
buf BUF1 (N599, N582);
buf BUF1 (N600, N597);
buf BUF1 (N601, N596);
and AND3 (N602, N585, N399, N384);
or OR4 (N603, N589, N115, N307, N268);
xor XOR2 (N604, N599, N557);
and AND3 (N605, N603, N237, N377);
or OR4 (N606, N598, N387, N547, N138);
xor XOR2 (N607, N602, N56);
or OR3 (N608, N593, N403, N176);
and AND4 (N609, N606, N210, N194, N104);
and AND3 (N610, N595, N311, N99);
xor XOR2 (N611, N609, N490);
buf BUF1 (N612, N604);
not NOT1 (N613, N607);
not NOT1 (N614, N613);
xor XOR2 (N615, N592, N222);
or OR2 (N616, N611, N44);
nor NOR3 (N617, N559, N67, N70);
nor NOR4 (N618, N614, N502, N324, N580);
xor XOR2 (N619, N610, N617);
xor XOR2 (N620, N436, N74);
or OR2 (N621, N605, N387);
nor NOR3 (N622, N601, N27, N611);
buf BUF1 (N623, N618);
xor XOR2 (N624, N622, N256);
buf BUF1 (N625, N619);
nor NOR3 (N626, N608, N527, N157);
nor NOR2 (N627, N623, N509);
nor NOR3 (N628, N627, N311, N132);
or OR4 (N629, N600, N245, N381, N122);
xor XOR2 (N630, N628, N204);
nand NAND4 (N631, N624, N541, N521, N363);
xor XOR2 (N632, N620, N628);
nand NAND4 (N633, N616, N386, N364, N194);
xor XOR2 (N634, N629, N349);
and AND2 (N635, N615, N107);
xor XOR2 (N636, N634, N72);
not NOT1 (N637, N621);
not NOT1 (N638, N631);
and AND4 (N639, N632, N444, N577, N340);
and AND4 (N640, N630, N602, N518, N360);
or OR4 (N641, N640, N605, N106, N386);
and AND2 (N642, N637, N197);
or OR2 (N643, N635, N381);
or OR2 (N644, N641, N184);
or OR2 (N645, N612, N279);
or OR4 (N646, N626, N321, N400, N143);
xor XOR2 (N647, N645, N295);
and AND2 (N648, N636, N548);
xor XOR2 (N649, N647, N430);
not NOT1 (N650, N646);
buf BUF1 (N651, N644);
nor NOR2 (N652, N625, N450);
nor NOR4 (N653, N651, N433, N161, N167);
not NOT1 (N654, N638);
nand NAND2 (N655, N654, N587);
buf BUF1 (N656, N653);
not NOT1 (N657, N652);
not NOT1 (N658, N633);
nor NOR3 (N659, N642, N477, N179);
xor XOR2 (N660, N658, N304);
not NOT1 (N661, N639);
buf BUF1 (N662, N660);
and AND4 (N663, N655, N218, N62, N62);
xor XOR2 (N664, N662, N584);
or OR3 (N665, N650, N455, N410);
nand NAND2 (N666, N661, N417);
and AND2 (N667, N643, N660);
or OR3 (N668, N657, N370, N169);
not NOT1 (N669, N668);
nand NAND4 (N670, N659, N211, N40, N387);
and AND4 (N671, N670, N424, N465, N446);
not NOT1 (N672, N664);
nor NOR2 (N673, N663, N19);
nor NOR4 (N674, N666, N347, N355, N311);
not NOT1 (N675, N671);
and AND3 (N676, N672, N318, N334);
nand NAND4 (N677, N665, N17, N218, N18);
or OR4 (N678, N674, N206, N391, N18);
buf BUF1 (N679, N676);
xor XOR2 (N680, N679, N188);
or OR3 (N681, N680, N528, N387);
nor NOR2 (N682, N673, N563);
or OR2 (N683, N682, N315);
xor XOR2 (N684, N667, N335);
not NOT1 (N685, N649);
buf BUF1 (N686, N656);
nand NAND2 (N687, N678, N357);
nor NOR3 (N688, N681, N306, N216);
and AND4 (N689, N687, N581, N81, N477);
nand NAND2 (N690, N675, N285);
and AND3 (N691, N684, N381, N681);
xor XOR2 (N692, N691, N361);
xor XOR2 (N693, N690, N531);
not NOT1 (N694, N677);
buf BUF1 (N695, N686);
buf BUF1 (N696, N683);
or OR2 (N697, N669, N246);
buf BUF1 (N698, N697);
nand NAND4 (N699, N694, N394, N136, N391);
buf BUF1 (N700, N648);
and AND3 (N701, N698, N420, N673);
xor XOR2 (N702, N685, N364);
buf BUF1 (N703, N689);
not NOT1 (N704, N693);
and AND3 (N705, N704, N623, N378);
and AND2 (N706, N701, N584);
xor XOR2 (N707, N706, N571);
xor XOR2 (N708, N688, N547);
nand NAND2 (N709, N707, N525);
nor NOR3 (N710, N703, N636, N334);
or OR4 (N711, N705, N564, N463, N677);
buf BUF1 (N712, N709);
nand NAND2 (N713, N695, N23);
buf BUF1 (N714, N699);
or OR3 (N715, N714, N365, N393);
or OR3 (N716, N713, N124, N46);
and AND4 (N717, N711, N89, N665, N251);
nor NOR4 (N718, N708, N479, N15, N651);
xor XOR2 (N719, N696, N651);
buf BUF1 (N720, N692);
nand NAND4 (N721, N700, N202, N675, N24);
nand NAND4 (N722, N715, N297, N335, N40);
nand NAND3 (N723, N722, N235, N488);
nor NOR3 (N724, N719, N468, N653);
xor XOR2 (N725, N724, N23);
nor NOR2 (N726, N721, N560);
nand NAND2 (N727, N718, N220);
xor XOR2 (N728, N727, N325);
xor XOR2 (N729, N702, N726);
nor NOR2 (N730, N425, N63);
and AND3 (N731, N723, N372, N359);
or OR4 (N732, N728, N617, N144, N505);
nor NOR3 (N733, N729, N540, N506);
not NOT1 (N734, N710);
xor XOR2 (N735, N720, N220);
nor NOR2 (N736, N717, N151);
not NOT1 (N737, N731);
xor XOR2 (N738, N725, N500);
buf BUF1 (N739, N734);
and AND3 (N740, N733, N229, N124);
buf BUF1 (N741, N730);
or OR3 (N742, N735, N132, N658);
not NOT1 (N743, N712);
not NOT1 (N744, N740);
nor NOR4 (N745, N716, N413, N535, N720);
xor XOR2 (N746, N741, N495);
or OR2 (N747, N744, N131);
or OR3 (N748, N737, N332, N124);
not NOT1 (N749, N738);
nand NAND2 (N750, N745, N504);
nor NOR2 (N751, N747, N744);
buf BUF1 (N752, N743);
and AND4 (N753, N748, N623, N272, N645);
or OR4 (N754, N732, N697, N458, N529);
and AND3 (N755, N750, N604, N116);
buf BUF1 (N756, N749);
buf BUF1 (N757, N746);
not NOT1 (N758, N754);
nand NAND4 (N759, N742, N272, N602, N563);
nand NAND4 (N760, N739, N163, N531, N460);
buf BUF1 (N761, N756);
nor NOR4 (N762, N752, N386, N335, N275);
or OR3 (N763, N736, N131, N242);
buf BUF1 (N764, N760);
nor NOR4 (N765, N763, N294, N329, N205);
or OR2 (N766, N759, N81);
or OR4 (N767, N765, N4, N470, N487);
or OR4 (N768, N762, N583, N223, N746);
xor XOR2 (N769, N758, N298);
nand NAND3 (N770, N755, N224, N701);
nor NOR4 (N771, N769, N456, N504, N18);
and AND3 (N772, N753, N695, N332);
and AND2 (N773, N761, N629);
not NOT1 (N774, N766);
buf BUF1 (N775, N772);
and AND4 (N776, N775, N343, N130, N63);
buf BUF1 (N777, N770);
or OR4 (N778, N774, N275, N171, N35);
and AND3 (N779, N778, N281, N427);
buf BUF1 (N780, N767);
nor NOR3 (N781, N771, N120, N487);
nand NAND4 (N782, N757, N622, N650, N131);
nand NAND4 (N783, N764, N498, N309, N427);
nor NOR2 (N784, N783, N436);
nor NOR4 (N785, N779, N544, N248, N415);
or OR2 (N786, N782, N404);
nand NAND2 (N787, N768, N158);
or OR2 (N788, N780, N570);
and AND2 (N789, N786, N433);
and AND4 (N790, N789, N179, N117, N324);
xor XOR2 (N791, N788, N533);
nand NAND2 (N792, N777, N546);
nor NOR3 (N793, N785, N21, N771);
buf BUF1 (N794, N773);
and AND2 (N795, N784, N647);
xor XOR2 (N796, N792, N528);
not NOT1 (N797, N794);
not NOT1 (N798, N795);
xor XOR2 (N799, N751, N142);
nand NAND4 (N800, N796, N169, N762, N486);
not NOT1 (N801, N799);
buf BUF1 (N802, N781);
nor NOR3 (N803, N802, N309, N686);
or OR4 (N804, N803, N711, N360, N562);
or OR4 (N805, N797, N351, N84, N319);
and AND4 (N806, N793, N459, N22, N717);
and AND4 (N807, N787, N634, N611, N720);
buf BUF1 (N808, N806);
buf BUF1 (N809, N798);
not NOT1 (N810, N807);
xor XOR2 (N811, N805, N68);
xor XOR2 (N812, N804, N86);
xor XOR2 (N813, N791, N708);
buf BUF1 (N814, N813);
buf BUF1 (N815, N800);
and AND3 (N816, N815, N513, N313);
nand NAND4 (N817, N816, N653, N130, N700);
or OR4 (N818, N801, N810, N646, N804);
or OR4 (N819, N288, N795, N541, N562);
or OR4 (N820, N808, N428, N387, N350);
nand NAND4 (N821, N776, N288, N360, N258);
nor NOR4 (N822, N820, N53, N160, N47);
nor NOR4 (N823, N822, N65, N58, N776);
not NOT1 (N824, N817);
buf BUF1 (N825, N790);
buf BUF1 (N826, N812);
not NOT1 (N827, N826);
and AND3 (N828, N809, N443, N317);
or OR4 (N829, N827, N355, N168, N610);
nor NOR3 (N830, N811, N723, N338);
nand NAND3 (N831, N824, N29, N116);
or OR2 (N832, N823, N313);
or OR4 (N833, N821, N372, N239, N416);
nand NAND4 (N834, N818, N125, N123, N492);
xor XOR2 (N835, N831, N21);
not NOT1 (N836, N829);
nor NOR4 (N837, N832, N208, N650, N225);
nand NAND3 (N838, N819, N177, N265);
not NOT1 (N839, N836);
buf BUF1 (N840, N834);
nor NOR3 (N841, N839, N355, N693);
nand NAND2 (N842, N833, N582);
and AND3 (N843, N837, N179, N469);
buf BUF1 (N844, N842);
nor NOR4 (N845, N843, N39, N323, N714);
xor XOR2 (N846, N844, N604);
nor NOR2 (N847, N830, N648);
not NOT1 (N848, N841);
not NOT1 (N849, N838);
and AND3 (N850, N835, N728, N608);
nand NAND4 (N851, N850, N337, N578, N337);
or OR2 (N852, N828, N532);
xor XOR2 (N853, N847, N439);
nor NOR3 (N854, N846, N449, N743);
buf BUF1 (N855, N854);
buf BUF1 (N856, N845);
nand NAND2 (N857, N856, N518);
xor XOR2 (N858, N855, N720);
and AND3 (N859, N851, N697, N445);
xor XOR2 (N860, N853, N55);
and AND2 (N861, N859, N255);
xor XOR2 (N862, N814, N607);
or OR4 (N863, N825, N164, N712, N144);
not NOT1 (N864, N852);
and AND4 (N865, N862, N295, N593, N567);
nor NOR2 (N866, N858, N138);
not NOT1 (N867, N840);
not NOT1 (N868, N857);
buf BUF1 (N869, N863);
buf BUF1 (N870, N861);
or OR2 (N871, N867, N237);
and AND3 (N872, N849, N612, N664);
xor XOR2 (N873, N872, N103);
and AND4 (N874, N864, N641, N661, N750);
and AND2 (N875, N848, N674);
buf BUF1 (N876, N865);
buf BUF1 (N877, N873);
xor XOR2 (N878, N870, N119);
nor NOR3 (N879, N876, N814, N47);
and AND4 (N880, N866, N766, N48, N23);
xor XOR2 (N881, N871, N39);
or OR4 (N882, N878, N34, N613, N490);
nand NAND4 (N883, N874, N235, N139, N532);
nor NOR3 (N884, N880, N13, N717);
not NOT1 (N885, N868);
buf BUF1 (N886, N877);
nand NAND2 (N887, N881, N160);
and AND4 (N888, N885, N548, N884, N43);
xor XOR2 (N889, N732, N29);
buf BUF1 (N890, N889);
not NOT1 (N891, N890);
or OR2 (N892, N882, N533);
xor XOR2 (N893, N860, N443);
xor XOR2 (N894, N892, N476);
or OR4 (N895, N875, N608, N776, N161);
buf BUF1 (N896, N879);
nand NAND4 (N897, N887, N447, N455, N673);
and AND4 (N898, N897, N64, N362, N659);
buf BUF1 (N899, N886);
nor NOR3 (N900, N898, N772, N227);
nand NAND2 (N901, N894, N272);
not NOT1 (N902, N869);
and AND4 (N903, N899, N262, N873, N427);
nor NOR3 (N904, N902, N606, N600);
xor XOR2 (N905, N904, N725);
xor XOR2 (N906, N900, N81);
not NOT1 (N907, N895);
nor NOR3 (N908, N896, N501, N898);
nand NAND2 (N909, N901, N440);
nor NOR4 (N910, N906, N114, N431, N56);
or OR2 (N911, N903, N569);
not NOT1 (N912, N907);
xor XOR2 (N913, N908, N797);
not NOT1 (N914, N912);
or OR3 (N915, N914, N440, N335);
nand NAND4 (N916, N913, N82, N124, N296);
xor XOR2 (N917, N905, N348);
and AND2 (N918, N893, N114);
nand NAND3 (N919, N911, N699, N716);
xor XOR2 (N920, N916, N640);
and AND4 (N921, N883, N70, N522, N129);
and AND2 (N922, N917, N39);
not NOT1 (N923, N915);
nor NOR4 (N924, N910, N900, N608, N556);
buf BUF1 (N925, N919);
xor XOR2 (N926, N888, N284);
or OR4 (N927, N925, N746, N351, N134);
and AND3 (N928, N921, N38, N60);
and AND3 (N929, N923, N91, N401);
buf BUF1 (N930, N920);
buf BUF1 (N931, N926);
not NOT1 (N932, N930);
or OR2 (N933, N927, N887);
nor NOR3 (N934, N932, N25, N40);
nor NOR2 (N935, N922, N365);
xor XOR2 (N936, N924, N586);
nor NOR2 (N937, N909, N511);
and AND4 (N938, N935, N317, N71, N5);
or OR4 (N939, N931, N491, N482, N429);
not NOT1 (N940, N933);
not NOT1 (N941, N934);
buf BUF1 (N942, N928);
or OR2 (N943, N938, N42);
nor NOR4 (N944, N929, N286, N427, N127);
not NOT1 (N945, N939);
nand NAND4 (N946, N940, N523, N11, N402);
buf BUF1 (N947, N946);
nor NOR3 (N948, N918, N859, N423);
or OR2 (N949, N937, N311);
xor XOR2 (N950, N944, N365);
xor XOR2 (N951, N891, N490);
xor XOR2 (N952, N942, N493);
not NOT1 (N953, N948);
buf BUF1 (N954, N947);
nor NOR3 (N955, N951, N839, N69);
not NOT1 (N956, N941);
xor XOR2 (N957, N945, N665);
buf BUF1 (N958, N936);
nand NAND2 (N959, N943, N579);
nand NAND3 (N960, N952, N496, N547);
nand NAND3 (N961, N959, N882, N232);
or OR4 (N962, N949, N443, N449, N744);
nand NAND4 (N963, N955, N565, N205, N269);
buf BUF1 (N964, N954);
nor NOR4 (N965, N961, N146, N481, N639);
not NOT1 (N966, N962);
and AND4 (N967, N956, N339, N631, N902);
nor NOR4 (N968, N957, N391, N632, N246);
xor XOR2 (N969, N966, N3);
nor NOR4 (N970, N960, N564, N186, N342);
buf BUF1 (N971, N970);
buf BUF1 (N972, N967);
and AND4 (N973, N971, N946, N748, N495);
nor NOR4 (N974, N968, N454, N176, N578);
or OR3 (N975, N963, N618, N829);
xor XOR2 (N976, N969, N137);
xor XOR2 (N977, N972, N270);
nor NOR4 (N978, N973, N938, N691, N912);
nor NOR3 (N979, N978, N230, N368);
or OR2 (N980, N975, N766);
and AND2 (N981, N980, N420);
buf BUF1 (N982, N953);
buf BUF1 (N983, N976);
or OR3 (N984, N958, N182, N754);
nor NOR3 (N985, N964, N204, N139);
not NOT1 (N986, N950);
and AND4 (N987, N982, N407, N626, N187);
not NOT1 (N988, N985);
and AND3 (N989, N981, N186, N520);
and AND3 (N990, N987, N595, N215);
not NOT1 (N991, N974);
buf BUF1 (N992, N991);
xor XOR2 (N993, N977, N817);
xor XOR2 (N994, N992, N581);
nand NAND4 (N995, N965, N231, N159, N461);
nand NAND4 (N996, N986, N362, N448, N217);
not NOT1 (N997, N995);
nand NAND4 (N998, N996, N663, N364, N955);
not NOT1 (N999, N990);
xor XOR2 (N1000, N989, N951);
and AND2 (N1001, N997, N326);
or OR4 (N1002, N993, N591, N767, N635);
buf BUF1 (N1003, N1002);
and AND3 (N1004, N979, N240, N420);
nor NOR2 (N1005, N1003, N666);
nand NAND2 (N1006, N983, N329);
buf BUF1 (N1007, N1006);
buf BUF1 (N1008, N1004);
or OR4 (N1009, N988, N255, N332, N49);
nor NOR4 (N1010, N998, N102, N156, N270);
and AND2 (N1011, N1001, N846);
nand NAND4 (N1012, N1007, N113, N66, N816);
and AND3 (N1013, N1009, N94, N317);
nand NAND3 (N1014, N984, N107, N255);
xor XOR2 (N1015, N1008, N902);
nand NAND2 (N1016, N999, N190);
xor XOR2 (N1017, N1010, N378);
or OR2 (N1018, N1016, N439);
not NOT1 (N1019, N1013);
and AND2 (N1020, N1015, N104);
xor XOR2 (N1021, N1011, N134);
or OR3 (N1022, N1020, N493, N951);
and AND4 (N1023, N1019, N73, N144, N926);
nor NOR3 (N1024, N1000, N475, N943);
buf BUF1 (N1025, N1018);
nor NOR4 (N1026, N1022, N969, N769, N550);
not NOT1 (N1027, N1014);
and AND4 (N1028, N1027, N1015, N112, N151);
buf BUF1 (N1029, N1023);
nand NAND3 (N1030, N1029, N688, N706);
nand NAND3 (N1031, N994, N260, N143);
buf BUF1 (N1032, N1005);
buf BUF1 (N1033, N1012);
or OR3 (N1034, N1032, N876, N615);
nand NAND3 (N1035, N1025, N970, N116);
nor NOR3 (N1036, N1035, N722, N18);
and AND4 (N1037, N1024, N162, N569, N423);
buf BUF1 (N1038, N1033);
buf BUF1 (N1039, N1021);
or OR3 (N1040, N1031, N922, N857);
not NOT1 (N1041, N1038);
or OR3 (N1042, N1037, N354, N308);
xor XOR2 (N1043, N1030, N189);
xor XOR2 (N1044, N1039, N909);
buf BUF1 (N1045, N1041);
nor NOR4 (N1046, N1043, N633, N16, N64);
nor NOR2 (N1047, N1036, N517);
not NOT1 (N1048, N1017);
nand NAND2 (N1049, N1040, N996);
not NOT1 (N1050, N1049);
buf BUF1 (N1051, N1042);
xor XOR2 (N1052, N1044, N524);
or OR4 (N1053, N1050, N111, N369, N261);
or OR2 (N1054, N1047, N1015);
not NOT1 (N1055, N1054);
nand NAND4 (N1056, N1045, N314, N512, N878);
nor NOR3 (N1057, N1053, N1022, N802);
and AND3 (N1058, N1048, N777, N195);
not NOT1 (N1059, N1058);
not NOT1 (N1060, N1051);
buf BUF1 (N1061, N1046);
nor NOR2 (N1062, N1056, N867);
buf BUF1 (N1063, N1057);
nand NAND4 (N1064, N1061, N892, N445, N929);
or OR2 (N1065, N1052, N839);
buf BUF1 (N1066, N1063);
buf BUF1 (N1067, N1055);
not NOT1 (N1068, N1028);
buf BUF1 (N1069, N1064);
and AND2 (N1070, N1026, N881);
not NOT1 (N1071, N1059);
not NOT1 (N1072, N1071);
nor NOR2 (N1073, N1072, N142);
nand NAND3 (N1074, N1073, N1072, N465);
not NOT1 (N1075, N1069);
nor NOR3 (N1076, N1075, N486, N167);
nor NOR2 (N1077, N1070, N823);
and AND4 (N1078, N1068, N488, N741, N637);
buf BUF1 (N1079, N1034);
nand NAND3 (N1080, N1067, N165, N806);
nand NAND2 (N1081, N1060, N1078);
nand NAND2 (N1082, N234, N113);
xor XOR2 (N1083, N1082, N788);
or OR2 (N1084, N1081, N884);
nand NAND4 (N1085, N1076, N450, N986, N916);
xor XOR2 (N1086, N1079, N716);
or OR2 (N1087, N1080, N885);
not NOT1 (N1088, N1062);
and AND3 (N1089, N1083, N12, N1011);
not NOT1 (N1090, N1089);
buf BUF1 (N1091, N1090);
not NOT1 (N1092, N1087);
or OR4 (N1093, N1085, N1007, N403, N1036);
and AND2 (N1094, N1088, N48);
buf BUF1 (N1095, N1086);
nand NAND3 (N1096, N1095, N391, N774);
xor XOR2 (N1097, N1091, N98);
nor NOR3 (N1098, N1093, N591, N151);
not NOT1 (N1099, N1066);
or OR2 (N1100, N1074, N47);
and AND2 (N1101, N1084, N954);
or OR3 (N1102, N1092, N770, N900);
or OR2 (N1103, N1101, N1005);
not NOT1 (N1104, N1099);
nand NAND2 (N1105, N1094, N884);
or OR2 (N1106, N1103, N539);
nand NAND2 (N1107, N1100, N1102);
xor XOR2 (N1108, N494, N697);
xor XOR2 (N1109, N1104, N1071);
xor XOR2 (N1110, N1106, N476);
and AND2 (N1111, N1109, N219);
nand NAND4 (N1112, N1107, N345, N977, N964);
not NOT1 (N1113, N1108);
and AND3 (N1114, N1113, N1036, N342);
nor NOR4 (N1115, N1105, N473, N756, N693);
and AND4 (N1116, N1114, N233, N245, N234);
xor XOR2 (N1117, N1065, N128);
and AND3 (N1118, N1115, N120, N707);
or OR2 (N1119, N1116, N661);
buf BUF1 (N1120, N1110);
nor NOR2 (N1121, N1111, N481);
xor XOR2 (N1122, N1097, N991);
and AND2 (N1123, N1119, N31);
or OR2 (N1124, N1118, N677);
buf BUF1 (N1125, N1098);
nand NAND3 (N1126, N1096, N60, N493);
nand NAND3 (N1127, N1117, N719, N913);
nor NOR3 (N1128, N1120, N419, N191);
or OR2 (N1129, N1125, N602);
nand NAND3 (N1130, N1127, N107, N841);
xor XOR2 (N1131, N1130, N1018);
xor XOR2 (N1132, N1112, N445);
not NOT1 (N1133, N1128);
nand NAND3 (N1134, N1124, N1020, N1101);
nand NAND2 (N1135, N1121, N681);
xor XOR2 (N1136, N1129, N410);
or OR2 (N1137, N1134, N755);
nand NAND2 (N1138, N1131, N619);
and AND4 (N1139, N1133, N623, N503, N733);
nor NOR2 (N1140, N1137, N1105);
buf BUF1 (N1141, N1122);
xor XOR2 (N1142, N1138, N199);
or OR4 (N1143, N1132, N1014, N228, N1074);
not NOT1 (N1144, N1142);
xor XOR2 (N1145, N1140, N952);
or OR2 (N1146, N1145, N950);
xor XOR2 (N1147, N1126, N950);
and AND4 (N1148, N1139, N1038, N714, N1039);
xor XOR2 (N1149, N1146, N346);
and AND3 (N1150, N1135, N200, N151);
not NOT1 (N1151, N1077);
nor NOR2 (N1152, N1147, N681);
nand NAND3 (N1153, N1150, N490, N239);
nand NAND4 (N1154, N1148, N212, N576, N706);
and AND4 (N1155, N1143, N730, N1017, N571);
not NOT1 (N1156, N1141);
xor XOR2 (N1157, N1149, N119);
and AND4 (N1158, N1136, N980, N196, N413);
or OR2 (N1159, N1153, N369);
or OR4 (N1160, N1158, N862, N261, N1051);
and AND3 (N1161, N1160, N268, N844);
not NOT1 (N1162, N1144);
not NOT1 (N1163, N1154);
buf BUF1 (N1164, N1157);
buf BUF1 (N1165, N1152);
buf BUF1 (N1166, N1163);
nor NOR2 (N1167, N1161, N840);
nand NAND2 (N1168, N1166, N490);
xor XOR2 (N1169, N1165, N1071);
nor NOR3 (N1170, N1162, N754, N111);
buf BUF1 (N1171, N1164);
or OR3 (N1172, N1156, N245, N927);
and AND3 (N1173, N1123, N471, N612);
nor NOR4 (N1174, N1168, N807, N308, N79);
xor XOR2 (N1175, N1155, N56);
nand NAND4 (N1176, N1172, N256, N305, N905);
nand NAND3 (N1177, N1173, N1144, N519);
xor XOR2 (N1178, N1169, N481);
not NOT1 (N1179, N1167);
nor NOR4 (N1180, N1177, N938, N834, N829);
xor XOR2 (N1181, N1174, N94);
nand NAND4 (N1182, N1175, N1, N1006, N838);
nand NAND3 (N1183, N1159, N896, N959);
buf BUF1 (N1184, N1183);
xor XOR2 (N1185, N1184, N850);
nand NAND4 (N1186, N1176, N868, N1177, N797);
and AND4 (N1187, N1151, N559, N755, N1030);
nand NAND4 (N1188, N1182, N506, N1156, N226);
nor NOR2 (N1189, N1179, N86);
nand NAND3 (N1190, N1180, N839, N835);
and AND2 (N1191, N1188, N572);
nand NAND2 (N1192, N1186, N761);
buf BUF1 (N1193, N1181);
and AND3 (N1194, N1187, N918, N917);
or OR4 (N1195, N1191, N24, N657, N234);
or OR2 (N1196, N1195, N660);
not NOT1 (N1197, N1193);
nand NAND4 (N1198, N1192, N314, N1156, N783);
not NOT1 (N1199, N1196);
xor XOR2 (N1200, N1185, N976);
not NOT1 (N1201, N1189);
buf BUF1 (N1202, N1198);
not NOT1 (N1203, N1178);
xor XOR2 (N1204, N1194, N830);
or OR2 (N1205, N1190, N385);
buf BUF1 (N1206, N1202);
or OR2 (N1207, N1200, N978);
nand NAND3 (N1208, N1207, N1086, N862);
or OR3 (N1209, N1208, N1177, N763);
nor NOR3 (N1210, N1170, N318, N786);
and AND2 (N1211, N1201, N1141);
not NOT1 (N1212, N1197);
and AND3 (N1213, N1209, N36, N49);
nor NOR3 (N1214, N1206, N543, N974);
xor XOR2 (N1215, N1212, N742);
nand NAND2 (N1216, N1203, N935);
nor NOR3 (N1217, N1213, N813, N625);
or OR4 (N1218, N1205, N885, N938, N1214);
nand NAND3 (N1219, N95, N796, N1100);
or OR4 (N1220, N1217, N438, N977, N860);
nand NAND2 (N1221, N1220, N508);
xor XOR2 (N1222, N1221, N1105);
not NOT1 (N1223, N1216);
nand NAND2 (N1224, N1199, N872);
nand NAND4 (N1225, N1223, N201, N1152, N1104);
nor NOR3 (N1226, N1204, N101, N656);
xor XOR2 (N1227, N1226, N42);
and AND3 (N1228, N1171, N680, N335);
nand NAND3 (N1229, N1228, N1063, N360);
buf BUF1 (N1230, N1210);
xor XOR2 (N1231, N1225, N974);
and AND4 (N1232, N1224, N742, N579, N273);
and AND3 (N1233, N1211, N192, N968);
buf BUF1 (N1234, N1227);
or OR3 (N1235, N1230, N1184, N525);
buf BUF1 (N1236, N1218);
nor NOR2 (N1237, N1235, N1025);
and AND3 (N1238, N1215, N399, N1182);
nand NAND3 (N1239, N1234, N535, N516);
nor NOR2 (N1240, N1233, N230);
xor XOR2 (N1241, N1236, N217);
buf BUF1 (N1242, N1219);
or OR2 (N1243, N1238, N1120);
xor XOR2 (N1244, N1240, N1034);
or OR4 (N1245, N1231, N384, N554, N186);
not NOT1 (N1246, N1242);
or OR4 (N1247, N1237, N83, N623, N326);
nor NOR2 (N1248, N1239, N615);
not NOT1 (N1249, N1247);
and AND4 (N1250, N1244, N1162, N269, N7);
buf BUF1 (N1251, N1250);
or OR4 (N1252, N1249, N371, N122, N137);
xor XOR2 (N1253, N1248, N1071);
and AND2 (N1254, N1229, N1116);
nand NAND4 (N1255, N1251, N146, N176, N1164);
nor NOR3 (N1256, N1252, N480, N695);
not NOT1 (N1257, N1241);
not NOT1 (N1258, N1257);
nand NAND4 (N1259, N1254, N470, N601, N701);
nand NAND2 (N1260, N1256, N503);
nand NAND3 (N1261, N1253, N675, N828);
or OR3 (N1262, N1246, N635, N745);
not NOT1 (N1263, N1222);
nor NOR2 (N1264, N1262, N1132);
buf BUF1 (N1265, N1264);
and AND3 (N1266, N1265, N33, N484);
buf BUF1 (N1267, N1245);
xor XOR2 (N1268, N1263, N1165);
not NOT1 (N1269, N1258);
xor XOR2 (N1270, N1260, N365);
and AND4 (N1271, N1267, N879, N1253, N894);
and AND2 (N1272, N1255, N1063);
not NOT1 (N1273, N1270);
or OR2 (N1274, N1243, N1251);
and AND2 (N1275, N1273, N662);
nor NOR3 (N1276, N1232, N880, N304);
or OR2 (N1277, N1266, N885);
nand NAND2 (N1278, N1272, N468);
not NOT1 (N1279, N1261);
nand NAND2 (N1280, N1277, N639);
not NOT1 (N1281, N1269);
or OR4 (N1282, N1281, N843, N928, N1058);
or OR3 (N1283, N1268, N10, N1275);
nor NOR2 (N1284, N880, N997);
not NOT1 (N1285, N1278);
and AND2 (N1286, N1285, N433);
nor NOR4 (N1287, N1280, N126, N57, N835);
nor NOR2 (N1288, N1276, N529);
nand NAND2 (N1289, N1283, N1115);
nand NAND4 (N1290, N1274, N864, N1108, N177);
and AND3 (N1291, N1279, N671, N382);
nand NAND4 (N1292, N1289, N138, N217, N575);
buf BUF1 (N1293, N1292);
buf BUF1 (N1294, N1286);
or OR4 (N1295, N1290, N882, N691, N178);
nor NOR4 (N1296, N1287, N940, N1178, N204);
buf BUF1 (N1297, N1259);
nor NOR3 (N1298, N1271, N110, N673);
nand NAND2 (N1299, N1282, N548);
or OR2 (N1300, N1297, N373);
xor XOR2 (N1301, N1300, N205);
not NOT1 (N1302, N1294);
and AND4 (N1303, N1298, N1103, N889, N1203);
buf BUF1 (N1304, N1295);
not NOT1 (N1305, N1302);
and AND4 (N1306, N1299, N218, N875, N287);
xor XOR2 (N1307, N1284, N921);
or OR2 (N1308, N1307, N662);
not NOT1 (N1309, N1306);
not NOT1 (N1310, N1308);
nor NOR3 (N1311, N1288, N766, N845);
buf BUF1 (N1312, N1301);
nand NAND3 (N1313, N1293, N1099, N231);
and AND2 (N1314, N1303, N1260);
buf BUF1 (N1315, N1291);
nand NAND2 (N1316, N1313, N284);
or OR2 (N1317, N1309, N719);
and AND3 (N1318, N1296, N1099, N775);
and AND3 (N1319, N1315, N1235, N268);
nor NOR4 (N1320, N1314, N739, N207, N1165);
buf BUF1 (N1321, N1316);
nor NOR2 (N1322, N1317, N992);
xor XOR2 (N1323, N1304, N202);
and AND3 (N1324, N1305, N349, N472);
xor XOR2 (N1325, N1312, N35);
xor XOR2 (N1326, N1323, N385);
nand NAND3 (N1327, N1326, N935, N474);
buf BUF1 (N1328, N1319);
nand NAND2 (N1329, N1324, N550);
and AND2 (N1330, N1321, N29);
or OR2 (N1331, N1329, N1212);
or OR3 (N1332, N1320, N671, N65);
or OR3 (N1333, N1330, N733, N985);
buf BUF1 (N1334, N1332);
nor NOR2 (N1335, N1327, N484);
not NOT1 (N1336, N1325);
buf BUF1 (N1337, N1318);
nor NOR2 (N1338, N1328, N21);
or OR3 (N1339, N1331, N287, N1245);
not NOT1 (N1340, N1337);
xor XOR2 (N1341, N1336, N322);
nor NOR4 (N1342, N1340, N711, N255, N669);
nand NAND3 (N1343, N1334, N38, N1320);
nand NAND3 (N1344, N1311, N475, N427);
and AND2 (N1345, N1310, N1026);
nand NAND3 (N1346, N1335, N819, N171);
nor NOR3 (N1347, N1345, N437, N240);
buf BUF1 (N1348, N1344);
nand NAND4 (N1349, N1339, N1344, N364, N444);
not NOT1 (N1350, N1322);
nand NAND4 (N1351, N1343, N1019, N22, N82);
xor XOR2 (N1352, N1350, N675);
nand NAND2 (N1353, N1341, N379);
buf BUF1 (N1354, N1353);
or OR3 (N1355, N1351, N668, N526);
and AND3 (N1356, N1347, N21, N472);
or OR4 (N1357, N1333, N137, N988, N233);
not NOT1 (N1358, N1342);
nor NOR2 (N1359, N1352, N676);
not NOT1 (N1360, N1354);
nand NAND2 (N1361, N1357, N574);
not NOT1 (N1362, N1356);
nor NOR4 (N1363, N1348, N578, N558, N403);
buf BUF1 (N1364, N1359);
or OR3 (N1365, N1355, N614, N877);
or OR3 (N1366, N1364, N433, N1061);
buf BUF1 (N1367, N1346);
xor XOR2 (N1368, N1338, N1070);
nand NAND4 (N1369, N1358, N233, N962, N983);
buf BUF1 (N1370, N1365);
xor XOR2 (N1371, N1366, N179);
or OR3 (N1372, N1361, N210, N326);
nand NAND3 (N1373, N1362, N155, N152);
nand NAND2 (N1374, N1373, N247);
nor NOR3 (N1375, N1367, N891, N247);
xor XOR2 (N1376, N1374, N287);
buf BUF1 (N1377, N1375);
nand NAND2 (N1378, N1349, N332);
and AND3 (N1379, N1360, N846, N625);
nor NOR3 (N1380, N1370, N579, N1009);
nor NOR2 (N1381, N1380, N497);
not NOT1 (N1382, N1372);
nand NAND2 (N1383, N1377, N1064);
xor XOR2 (N1384, N1369, N439);
nor NOR4 (N1385, N1383, N827, N464, N910);
nand NAND4 (N1386, N1371, N1219, N338, N384);
nand NAND4 (N1387, N1382, N1059, N310, N880);
buf BUF1 (N1388, N1386);
buf BUF1 (N1389, N1378);
nand NAND4 (N1390, N1379, N546, N61, N257);
nor NOR4 (N1391, N1381, N323, N998, N847);
or OR4 (N1392, N1368, N613, N155, N1205);
nand NAND3 (N1393, N1392, N140, N313);
nand NAND2 (N1394, N1363, N899);
or OR2 (N1395, N1390, N226);
buf BUF1 (N1396, N1394);
and AND2 (N1397, N1376, N714);
buf BUF1 (N1398, N1391);
or OR2 (N1399, N1387, N528);
xor XOR2 (N1400, N1396, N936);
nor NOR2 (N1401, N1385, N96);
nor NOR4 (N1402, N1389, N961, N1231, N589);
or OR3 (N1403, N1401, N1395, N779);
xor XOR2 (N1404, N684, N793);
nand NAND4 (N1405, N1384, N715, N814, N1297);
not NOT1 (N1406, N1400);
not NOT1 (N1407, N1399);
not NOT1 (N1408, N1407);
buf BUF1 (N1409, N1408);
nor NOR4 (N1410, N1409, N144, N538, N100);
and AND4 (N1411, N1402, N848, N492, N743);
nor NOR4 (N1412, N1410, N80, N843, N683);
not NOT1 (N1413, N1406);
nand NAND4 (N1414, N1411, N205, N16, N444);
buf BUF1 (N1415, N1403);
nor NOR3 (N1416, N1415, N1060, N183);
buf BUF1 (N1417, N1413);
nor NOR3 (N1418, N1398, N789, N1173);
nand NAND4 (N1419, N1416, N116, N785, N246);
xor XOR2 (N1420, N1393, N482);
or OR2 (N1421, N1417, N419);
not NOT1 (N1422, N1418);
nand NAND4 (N1423, N1421, N1309, N936, N1327);
and AND2 (N1424, N1423, N363);
or OR3 (N1425, N1388, N1254, N712);
nand NAND4 (N1426, N1419, N1265, N764, N388);
buf BUF1 (N1427, N1420);
and AND3 (N1428, N1414, N629, N1217);
nand NAND3 (N1429, N1427, N855, N393);
buf BUF1 (N1430, N1412);
buf BUF1 (N1431, N1430);
not NOT1 (N1432, N1424);
or OR2 (N1433, N1397, N908);
buf BUF1 (N1434, N1425);
not NOT1 (N1435, N1404);
nor NOR2 (N1436, N1433, N468);
nor NOR3 (N1437, N1434, N483, N536);
not NOT1 (N1438, N1437);
xor XOR2 (N1439, N1432, N912);
nand NAND3 (N1440, N1422, N775, N1290);
or OR2 (N1441, N1439, N424);
xor XOR2 (N1442, N1405, N89);
nand NAND4 (N1443, N1440, N1418, N746, N1096);
buf BUF1 (N1444, N1442);
nand NAND2 (N1445, N1443, N289);
not NOT1 (N1446, N1429);
xor XOR2 (N1447, N1446, N760);
nor NOR3 (N1448, N1444, N764, N768);
buf BUF1 (N1449, N1447);
buf BUF1 (N1450, N1445);
and AND2 (N1451, N1428, N506);
or OR3 (N1452, N1441, N504, N340);
and AND4 (N1453, N1451, N1067, N647, N927);
nor NOR4 (N1454, N1449, N858, N1151, N178);
or OR2 (N1455, N1454, N1097);
xor XOR2 (N1456, N1452, N30);
not NOT1 (N1457, N1435);
xor XOR2 (N1458, N1436, N603);
xor XOR2 (N1459, N1456, N942);
nand NAND3 (N1460, N1455, N26, N1028);
nand NAND4 (N1461, N1448, N901, N734, N1109);
buf BUF1 (N1462, N1458);
xor XOR2 (N1463, N1450, N1325);
and AND3 (N1464, N1426, N721, N362);
not NOT1 (N1465, N1459);
nand NAND3 (N1466, N1460, N731, N971);
xor XOR2 (N1467, N1466, N343);
not NOT1 (N1468, N1438);
and AND3 (N1469, N1464, N536, N357);
nor NOR4 (N1470, N1467, N778, N1375, N84);
nor NOR4 (N1471, N1468, N422, N524, N1047);
nor NOR2 (N1472, N1465, N1363);
not NOT1 (N1473, N1472);
xor XOR2 (N1474, N1469, N848);
nor NOR2 (N1475, N1471, N1338);
buf BUF1 (N1476, N1475);
not NOT1 (N1477, N1461);
nand NAND4 (N1478, N1462, N469, N413, N1065);
nand NAND4 (N1479, N1457, N1261, N476, N992);
not NOT1 (N1480, N1431);
nor NOR2 (N1481, N1479, N1334);
or OR2 (N1482, N1473, N1025);
nand NAND2 (N1483, N1474, N475);
or OR3 (N1484, N1483, N1055, N726);
nand NAND4 (N1485, N1481, N1448, N1267, N164);
buf BUF1 (N1486, N1478);
and AND3 (N1487, N1486, N834, N430);
nor NOR3 (N1488, N1487, N922, N1436);
nor NOR2 (N1489, N1476, N1478);
buf BUF1 (N1490, N1477);
and AND4 (N1491, N1488, N1380, N323, N214);
nor NOR2 (N1492, N1484, N696);
nor NOR4 (N1493, N1480, N857, N38, N768);
nor NOR2 (N1494, N1492, N9);
or OR3 (N1495, N1485, N554, N709);
nor NOR4 (N1496, N1453, N513, N289, N601);
nand NAND4 (N1497, N1482, N1101, N516, N609);
nor NOR4 (N1498, N1491, N976, N1403, N1075);
nand NAND4 (N1499, N1470, N1087, N523, N464);
nand NAND3 (N1500, N1497, N1271, N1477);
and AND3 (N1501, N1496, N977, N100);
or OR3 (N1502, N1493, N367, N355);
nand NAND3 (N1503, N1489, N594, N1299);
not NOT1 (N1504, N1499);
xor XOR2 (N1505, N1504, N756);
nand NAND2 (N1506, N1494, N1483);
not NOT1 (N1507, N1495);
or OR4 (N1508, N1507, N904, N859, N1438);
nand NAND3 (N1509, N1505, N1258, N902);
nand NAND4 (N1510, N1490, N854, N973, N414);
xor XOR2 (N1511, N1509, N1154);
and AND2 (N1512, N1508, N543);
buf BUF1 (N1513, N1502);
not NOT1 (N1514, N1513);
nor NOR2 (N1515, N1506, N798);
nor NOR4 (N1516, N1514, N1443, N1145, N785);
and AND4 (N1517, N1516, N1202, N952, N983);
buf BUF1 (N1518, N1500);
and AND3 (N1519, N1498, N691, N1360);
buf BUF1 (N1520, N1512);
and AND2 (N1521, N1463, N78);
or OR3 (N1522, N1511, N994, N587);
not NOT1 (N1523, N1521);
or OR3 (N1524, N1520, N1489, N253);
nand NAND4 (N1525, N1524, N901, N728, N616);
nand NAND2 (N1526, N1518, N1413);
not NOT1 (N1527, N1503);
nand NAND3 (N1528, N1517, N1480, N531);
or OR2 (N1529, N1515, N642);
xor XOR2 (N1530, N1526, N824);
nand NAND2 (N1531, N1522, N686);
nand NAND4 (N1532, N1525, N455, N1306, N1088);
not NOT1 (N1533, N1528);
xor XOR2 (N1534, N1523, N586);
and AND4 (N1535, N1510, N633, N1408, N759);
nor NOR2 (N1536, N1532, N1216);
and AND4 (N1537, N1531, N143, N782, N1446);
and AND3 (N1538, N1533, N631, N1145);
nand NAND4 (N1539, N1519, N150, N1430, N1223);
not NOT1 (N1540, N1529);
not NOT1 (N1541, N1536);
not NOT1 (N1542, N1501);
buf BUF1 (N1543, N1538);
or OR2 (N1544, N1537, N1415);
not NOT1 (N1545, N1535);
not NOT1 (N1546, N1530);
nor NOR3 (N1547, N1543, N1132, N460);
nor NOR4 (N1548, N1541, N543, N1133, N468);
nand NAND2 (N1549, N1539, N1158);
xor XOR2 (N1550, N1544, N1196);
and AND2 (N1551, N1540, N144);
nand NAND4 (N1552, N1551, N347, N635, N511);
xor XOR2 (N1553, N1552, N1154);
or OR3 (N1554, N1548, N679, N223);
nor NOR3 (N1555, N1542, N789, N831);
not NOT1 (N1556, N1545);
buf BUF1 (N1557, N1547);
nor NOR4 (N1558, N1527, N426, N314, N533);
and AND2 (N1559, N1556, N779);
or OR2 (N1560, N1559, N816);
buf BUF1 (N1561, N1553);
or OR2 (N1562, N1557, N1289);
nand NAND4 (N1563, N1550, N972, N759, N379);
xor XOR2 (N1564, N1555, N723);
nor NOR3 (N1565, N1560, N1379, N1245);
buf BUF1 (N1566, N1549);
nor NOR4 (N1567, N1546, N567, N369, N921);
nand NAND3 (N1568, N1534, N780, N706);
and AND2 (N1569, N1563, N505);
nand NAND4 (N1570, N1564, N959, N1213, N263);
buf BUF1 (N1571, N1562);
or OR3 (N1572, N1566, N17, N1493);
nor NOR4 (N1573, N1572, N1439, N987, N1264);
or OR4 (N1574, N1554, N147, N847, N1155);
not NOT1 (N1575, N1567);
not NOT1 (N1576, N1568);
and AND3 (N1577, N1570, N378, N965);
and AND4 (N1578, N1558, N1414, N606, N341);
xor XOR2 (N1579, N1571, N1154);
nand NAND3 (N1580, N1575, N103, N1290);
xor XOR2 (N1581, N1577, N114);
nand NAND3 (N1582, N1580, N324, N427);
buf BUF1 (N1583, N1582);
buf BUF1 (N1584, N1573);
nor NOR2 (N1585, N1574, N330);
not NOT1 (N1586, N1585);
nor NOR3 (N1587, N1586, N1310, N476);
and AND3 (N1588, N1565, N213, N1300);
buf BUF1 (N1589, N1583);
xor XOR2 (N1590, N1578, N940);
not NOT1 (N1591, N1569);
or OR4 (N1592, N1590, N959, N497, N122);
xor XOR2 (N1593, N1591, N34);
nor NOR3 (N1594, N1584, N718, N1384);
or OR4 (N1595, N1593, N912, N1494, N1403);
nand NAND4 (N1596, N1581, N1526, N1564, N435);
and AND2 (N1597, N1576, N323);
or OR2 (N1598, N1596, N267);
nand NAND3 (N1599, N1588, N1484, N820);
buf BUF1 (N1600, N1598);
nand NAND2 (N1601, N1589, N820);
and AND4 (N1602, N1600, N124, N675, N332);
or OR4 (N1603, N1561, N1463, N351, N292);
nor NOR4 (N1604, N1597, N981, N898, N980);
nand NAND2 (N1605, N1592, N849);
nand NAND3 (N1606, N1579, N452, N345);
not NOT1 (N1607, N1594);
and AND4 (N1608, N1605, N216, N531, N617);
or OR4 (N1609, N1599, N1153, N1380, N1362);
not NOT1 (N1610, N1587);
and AND2 (N1611, N1608, N1390);
and AND2 (N1612, N1609, N161);
or OR3 (N1613, N1604, N284, N1564);
or OR2 (N1614, N1610, N483);
xor XOR2 (N1615, N1611, N1444);
xor XOR2 (N1616, N1614, N1458);
buf BUF1 (N1617, N1595);
and AND2 (N1618, N1615, N1557);
and AND4 (N1619, N1603, N112, N897, N1434);
or OR3 (N1620, N1613, N322, N274);
nor NOR4 (N1621, N1607, N574, N797, N1247);
nand NAND3 (N1622, N1621, N498, N1440);
not NOT1 (N1623, N1602);
buf BUF1 (N1624, N1617);
buf BUF1 (N1625, N1624);
nor NOR2 (N1626, N1623, N1578);
buf BUF1 (N1627, N1622);
xor XOR2 (N1628, N1616, N44);
not NOT1 (N1629, N1606);
nor NOR3 (N1630, N1618, N1605, N495);
and AND4 (N1631, N1630, N1323, N723, N1216);
buf BUF1 (N1632, N1625);
nor NOR2 (N1633, N1632, N1228);
buf BUF1 (N1634, N1620);
buf BUF1 (N1635, N1633);
nand NAND4 (N1636, N1629, N603, N332, N458);
nor NOR2 (N1637, N1634, N510);
and AND3 (N1638, N1627, N1278, N1369);
buf BUF1 (N1639, N1635);
or OR4 (N1640, N1636, N513, N904, N1256);
or OR4 (N1641, N1639, N1174, N1293, N638);
nand NAND4 (N1642, N1641, N13, N576, N827);
xor XOR2 (N1643, N1638, N46);
or OR2 (N1644, N1637, N958);
nand NAND3 (N1645, N1628, N1550, N795);
or OR3 (N1646, N1645, N1642, N681);
buf BUF1 (N1647, N982);
and AND2 (N1648, N1644, N122);
and AND4 (N1649, N1631, N660, N307, N305);
or OR4 (N1650, N1649, N1278, N346, N469);
nand NAND4 (N1651, N1646, N1314, N612, N898);
or OR2 (N1652, N1648, N1297);
buf BUF1 (N1653, N1651);
and AND3 (N1654, N1640, N1437, N729);
xor XOR2 (N1655, N1654, N430);
nand NAND2 (N1656, N1655, N53);
buf BUF1 (N1657, N1650);
buf BUF1 (N1658, N1652);
buf BUF1 (N1659, N1626);
xor XOR2 (N1660, N1643, N123);
not NOT1 (N1661, N1619);
xor XOR2 (N1662, N1601, N747);
or OR3 (N1663, N1661, N347, N1119);
nand NAND3 (N1664, N1647, N189, N891);
xor XOR2 (N1665, N1662, N607);
nand NAND2 (N1666, N1657, N663);
nor NOR4 (N1667, N1612, N1111, N1474, N1280);
nand NAND3 (N1668, N1658, N261, N356);
nand NAND3 (N1669, N1665, N31, N1048);
buf BUF1 (N1670, N1664);
nor NOR4 (N1671, N1659, N1631, N398, N853);
not NOT1 (N1672, N1653);
nand NAND4 (N1673, N1656, N620, N1291, N36);
nor NOR4 (N1674, N1673, N850, N129, N1239);
xor XOR2 (N1675, N1667, N1093);
nand NAND2 (N1676, N1670, N554);
not NOT1 (N1677, N1674);
or OR3 (N1678, N1677, N178, N363);
nor NOR2 (N1679, N1678, N1520);
nor NOR3 (N1680, N1672, N336, N399);
buf BUF1 (N1681, N1675);
nand NAND2 (N1682, N1679, N334);
and AND4 (N1683, N1671, N471, N1342, N331);
nand NAND2 (N1684, N1663, N448);
and AND4 (N1685, N1660, N52, N1671, N1102);
nor NOR4 (N1686, N1684, N16, N670, N1096);
xor XOR2 (N1687, N1685, N159);
nor NOR2 (N1688, N1668, N1035);
not NOT1 (N1689, N1681);
buf BUF1 (N1690, N1676);
nor NOR3 (N1691, N1666, N1458, N704);
or OR4 (N1692, N1691, N543, N1665, N1554);
nand NAND2 (N1693, N1687, N307);
or OR2 (N1694, N1688, N798);
or OR2 (N1695, N1689, N1547);
buf BUF1 (N1696, N1669);
or OR4 (N1697, N1682, N992, N1395, N27);
nand NAND3 (N1698, N1680, N1344, N918);
xor XOR2 (N1699, N1695, N1317);
or OR2 (N1700, N1699, N1498);
xor XOR2 (N1701, N1694, N1132);
nor NOR3 (N1702, N1698, N973, N281);
and AND2 (N1703, N1686, N907);
and AND2 (N1704, N1696, N917);
nor NOR3 (N1705, N1692, N44, N606);
buf BUF1 (N1706, N1702);
nor NOR4 (N1707, N1706, N1550, N1584, N1170);
nand NAND2 (N1708, N1704, N1549);
nor NOR2 (N1709, N1707, N601);
buf BUF1 (N1710, N1690);
nor NOR2 (N1711, N1701, N987);
nand NAND2 (N1712, N1708, N771);
and AND2 (N1713, N1710, N112);
and AND4 (N1714, N1709, N1504, N1651, N467);
xor XOR2 (N1715, N1693, N1215);
xor XOR2 (N1716, N1703, N150);
buf BUF1 (N1717, N1697);
buf BUF1 (N1718, N1714);
xor XOR2 (N1719, N1705, N317);
or OR4 (N1720, N1712, N478, N1691, N1242);
nand NAND4 (N1721, N1719, N450, N1058, N1083);
or OR3 (N1722, N1721, N1538, N1607);
nand NAND2 (N1723, N1717, N1501);
buf BUF1 (N1724, N1711);
nand NAND2 (N1725, N1700, N1580);
buf BUF1 (N1726, N1716);
nand NAND2 (N1727, N1725, N1506);
xor XOR2 (N1728, N1727, N788);
and AND3 (N1729, N1726, N38, N944);
nor NOR2 (N1730, N1718, N100);
nor NOR3 (N1731, N1729, N503, N449);
nand NAND2 (N1732, N1720, N1147);
xor XOR2 (N1733, N1730, N1335);
or OR2 (N1734, N1733, N46);
nor NOR3 (N1735, N1734, N1317, N645);
nand NAND4 (N1736, N1724, N986, N1282, N190);
nand NAND2 (N1737, N1731, N167);
and AND4 (N1738, N1737, N1203, N50, N386);
and AND3 (N1739, N1723, N1255, N1438);
buf BUF1 (N1740, N1715);
nand NAND4 (N1741, N1736, N988, N547, N699);
not NOT1 (N1742, N1735);
not NOT1 (N1743, N1722);
xor XOR2 (N1744, N1713, N1159);
nor NOR4 (N1745, N1741, N165, N545, N1069);
xor XOR2 (N1746, N1732, N41);
or OR3 (N1747, N1738, N1548, N168);
or OR4 (N1748, N1742, N938, N1126, N1571);
buf BUF1 (N1749, N1745);
nand NAND3 (N1750, N1749, N647, N1671);
or OR3 (N1751, N1744, N156, N1081);
nor NOR2 (N1752, N1748, N614);
xor XOR2 (N1753, N1747, N1746);
xor XOR2 (N1754, N835, N1254);
or OR4 (N1755, N1750, N408, N251, N1738);
nor NOR4 (N1756, N1754, N546, N676, N971);
not NOT1 (N1757, N1739);
nand NAND3 (N1758, N1752, N805, N1032);
nand NAND2 (N1759, N1740, N1387);
nor NOR4 (N1760, N1755, N404, N1081, N1410);
or OR3 (N1761, N1753, N952, N1026);
nor NOR4 (N1762, N1761, N975, N259, N721);
and AND2 (N1763, N1756, N1050);
buf BUF1 (N1764, N1751);
xor XOR2 (N1765, N1758, N1499);
nor NOR4 (N1766, N1728, N1399, N356, N1527);
not NOT1 (N1767, N1757);
not NOT1 (N1768, N1763);
buf BUF1 (N1769, N1767);
buf BUF1 (N1770, N1768);
or OR2 (N1771, N1759, N1671);
or OR2 (N1772, N1769, N1311);
nor NOR2 (N1773, N1762, N1205);
not NOT1 (N1774, N1764);
and AND4 (N1775, N1773, N393, N499, N1689);
buf BUF1 (N1776, N1760);
buf BUF1 (N1777, N1765);
and AND4 (N1778, N1770, N27, N1546, N1658);
not NOT1 (N1779, N1743);
and AND2 (N1780, N1778, N1762);
xor XOR2 (N1781, N1772, N9);
nand NAND2 (N1782, N1775, N710);
and AND3 (N1783, N1774, N1742, N1434);
nor NOR3 (N1784, N1782, N124, N1027);
buf BUF1 (N1785, N1779);
and AND2 (N1786, N1780, N456);
not NOT1 (N1787, N1766);
buf BUF1 (N1788, N1786);
not NOT1 (N1789, N1785);
xor XOR2 (N1790, N1776, N1136);
or OR2 (N1791, N1771, N1525);
or OR2 (N1792, N1790, N37);
not NOT1 (N1793, N1791);
nand NAND4 (N1794, N1788, N152, N1327, N364);
buf BUF1 (N1795, N1683);
nor NOR4 (N1796, N1794, N538, N1023, N1704);
xor XOR2 (N1797, N1781, N1281);
nor NOR2 (N1798, N1792, N1003);
nor NOR4 (N1799, N1797, N739, N775, N666);
nor NOR4 (N1800, N1787, N995, N492, N395);
not NOT1 (N1801, N1798);
or OR2 (N1802, N1800, N818);
or OR3 (N1803, N1799, N1694, N19);
not NOT1 (N1804, N1801);
nand NAND3 (N1805, N1795, N794, N209);
or OR4 (N1806, N1777, N1677, N561, N107);
nor NOR2 (N1807, N1804, N1722);
nand NAND4 (N1808, N1784, N1701, N855, N652);
and AND4 (N1809, N1807, N175, N86, N202);
nand NAND4 (N1810, N1809, N377, N1341, N1145);
buf BUF1 (N1811, N1789);
xor XOR2 (N1812, N1793, N846);
nor NOR2 (N1813, N1783, N379);
and AND4 (N1814, N1810, N1407, N4, N380);
buf BUF1 (N1815, N1813);
and AND2 (N1816, N1806, N1033);
buf BUF1 (N1817, N1803);
not NOT1 (N1818, N1805);
nand NAND2 (N1819, N1808, N697);
and AND2 (N1820, N1812, N802);
buf BUF1 (N1821, N1815);
or OR2 (N1822, N1814, N346);
xor XOR2 (N1823, N1819, N1547);
nand NAND2 (N1824, N1816, N278);
or OR4 (N1825, N1796, N1536, N836, N205);
xor XOR2 (N1826, N1802, N1141);
buf BUF1 (N1827, N1817);
nor NOR3 (N1828, N1824, N1505, N1767);
nor NOR2 (N1829, N1825, N274);
nand NAND4 (N1830, N1821, N1318, N1227, N1609);
nor NOR2 (N1831, N1818, N1655);
nand NAND2 (N1832, N1831, N617);
nor NOR4 (N1833, N1811, N1387, N213, N1166);
nor NOR4 (N1834, N1829, N1516, N1583, N574);
nand NAND3 (N1835, N1833, N1245, N1510);
not NOT1 (N1836, N1823);
buf BUF1 (N1837, N1822);
nand NAND3 (N1838, N1826, N755, N1470);
and AND3 (N1839, N1820, N618, N974);
nor NOR2 (N1840, N1828, N835);
xor XOR2 (N1841, N1835, N1485);
xor XOR2 (N1842, N1838, N1357);
not NOT1 (N1843, N1832);
not NOT1 (N1844, N1843);
nand NAND4 (N1845, N1839, N919, N1083, N1535);
not NOT1 (N1846, N1840);
not NOT1 (N1847, N1834);
nor NOR2 (N1848, N1847, N1076);
xor XOR2 (N1849, N1844, N1415);
xor XOR2 (N1850, N1827, N439);
xor XOR2 (N1851, N1830, N1314);
xor XOR2 (N1852, N1836, N922);
nor NOR3 (N1853, N1837, N337, N278);
buf BUF1 (N1854, N1850);
or OR4 (N1855, N1848, N849, N194, N604);
not NOT1 (N1856, N1846);
not NOT1 (N1857, N1856);
buf BUF1 (N1858, N1849);
and AND4 (N1859, N1852, N731, N1348, N1486);
nand NAND3 (N1860, N1855, N233, N490);
and AND3 (N1861, N1857, N1706, N1089);
nor NOR4 (N1862, N1861, N1128, N1431, N837);
xor XOR2 (N1863, N1854, N931);
buf BUF1 (N1864, N1851);
buf BUF1 (N1865, N1845);
xor XOR2 (N1866, N1862, N754);
xor XOR2 (N1867, N1860, N598);
buf BUF1 (N1868, N1866);
nor NOR3 (N1869, N1867, N1156, N899);
nand NAND4 (N1870, N1869, N1463, N4, N143);
nor NOR2 (N1871, N1853, N828);
nor NOR2 (N1872, N1842, N1064);
and AND2 (N1873, N1841, N1020);
nand NAND2 (N1874, N1872, N1826);
or OR2 (N1875, N1873, N140);
nor NOR3 (N1876, N1874, N1819, N277);
nand NAND4 (N1877, N1859, N1086, N813, N700);
nor NOR4 (N1878, N1875, N582, N919, N264);
not NOT1 (N1879, N1864);
xor XOR2 (N1880, N1877, N94);
or OR2 (N1881, N1863, N648);
nor NOR3 (N1882, N1858, N1036, N1817);
not NOT1 (N1883, N1876);
xor XOR2 (N1884, N1871, N1326);
xor XOR2 (N1885, N1878, N1423);
nand NAND3 (N1886, N1883, N75, N92);
and AND4 (N1887, N1886, N187, N865, N348);
and AND2 (N1888, N1879, N1536);
nand NAND4 (N1889, N1870, N444, N700, N912);
and AND3 (N1890, N1889, N702, N141);
not NOT1 (N1891, N1868);
or OR3 (N1892, N1884, N1488, N433);
not NOT1 (N1893, N1865);
nor NOR4 (N1894, N1881, N1103, N1829, N88);
xor XOR2 (N1895, N1894, N1059);
or OR3 (N1896, N1882, N686, N366);
or OR2 (N1897, N1887, N313);
or OR2 (N1898, N1885, N299);
and AND3 (N1899, N1880, N1703, N751);
xor XOR2 (N1900, N1895, N264);
and AND3 (N1901, N1897, N1119, N105);
buf BUF1 (N1902, N1892);
or OR2 (N1903, N1898, N1650);
or OR2 (N1904, N1901, N340);
nor NOR4 (N1905, N1891, N1128, N1721, N1432);
nor NOR3 (N1906, N1904, N506, N474);
buf BUF1 (N1907, N1903);
buf BUF1 (N1908, N1888);
nor NOR4 (N1909, N1906, N1837, N1651, N1871);
xor XOR2 (N1910, N1900, N814);
buf BUF1 (N1911, N1910);
buf BUF1 (N1912, N1893);
buf BUF1 (N1913, N1909);
buf BUF1 (N1914, N1908);
buf BUF1 (N1915, N1905);
nor NOR3 (N1916, N1914, N372, N403);
not NOT1 (N1917, N1902);
and AND3 (N1918, N1915, N1700, N1765);
and AND3 (N1919, N1907, N1639, N1164);
xor XOR2 (N1920, N1913, N1917);
nand NAND2 (N1921, N411, N1502);
nor NOR4 (N1922, N1890, N881, N1521, N1880);
buf BUF1 (N1923, N1922);
not NOT1 (N1924, N1920);
xor XOR2 (N1925, N1919, N931);
or OR2 (N1926, N1912, N1506);
nor NOR2 (N1927, N1918, N1385);
or OR3 (N1928, N1927, N976, N1127);
xor XOR2 (N1929, N1899, N1087);
not NOT1 (N1930, N1923);
nand NAND3 (N1931, N1929, N697, N1089);
not NOT1 (N1932, N1928);
or OR3 (N1933, N1916, N1792, N992);
nand NAND3 (N1934, N1926, N695, N105);
not NOT1 (N1935, N1932);
or OR2 (N1936, N1935, N1420);
nor NOR3 (N1937, N1925, N940, N1658);
nor NOR4 (N1938, N1936, N1689, N1225, N1292);
and AND4 (N1939, N1896, N705, N57, N885);
nand NAND3 (N1940, N1911, N1136, N1135);
xor XOR2 (N1941, N1933, N217);
not NOT1 (N1942, N1924);
buf BUF1 (N1943, N1921);
nor NOR4 (N1944, N1939, N1486, N909, N1372);
or OR3 (N1945, N1941, N1690, N385);
xor XOR2 (N1946, N1940, N563);
or OR2 (N1947, N1944, N1494);
buf BUF1 (N1948, N1934);
buf BUF1 (N1949, N1930);
not NOT1 (N1950, N1949);
xor XOR2 (N1951, N1946, N981);
not NOT1 (N1952, N1950);
nor NOR3 (N1953, N1948, N216, N647);
xor XOR2 (N1954, N1951, N1376);
xor XOR2 (N1955, N1942, N195);
nor NOR4 (N1956, N1952, N1810, N1763, N41);
nand NAND3 (N1957, N1945, N953, N1017);
and AND3 (N1958, N1953, N398, N1859);
or OR2 (N1959, N1955, N681);
nor NOR4 (N1960, N1958, N335, N623, N645);
buf BUF1 (N1961, N1937);
not NOT1 (N1962, N1959);
not NOT1 (N1963, N1947);
nor NOR3 (N1964, N1963, N397, N1570);
not NOT1 (N1965, N1960);
buf BUF1 (N1966, N1931);
not NOT1 (N1967, N1961);
and AND4 (N1968, N1967, N1496, N1324, N162);
buf BUF1 (N1969, N1968);
nor NOR2 (N1970, N1943, N1286);
or OR2 (N1971, N1954, N1703);
or OR3 (N1972, N1966, N503, N303);
not NOT1 (N1973, N1962);
not NOT1 (N1974, N1973);
xor XOR2 (N1975, N1956, N1162);
and AND2 (N1976, N1957, N1219);
nand NAND4 (N1977, N1976, N1326, N466, N942);
nand NAND3 (N1978, N1977, N1721, N1409);
and AND3 (N1979, N1974, N784, N1172);
nor NOR2 (N1980, N1971, N1062);
or OR3 (N1981, N1964, N451, N269);
and AND2 (N1982, N1969, N1569);
nand NAND2 (N1983, N1980, N773);
xor XOR2 (N1984, N1979, N20);
nand NAND3 (N1985, N1965, N1502, N955);
xor XOR2 (N1986, N1982, N80);
not NOT1 (N1987, N1984);
not NOT1 (N1988, N1972);
nand NAND2 (N1989, N1975, N1364);
and AND2 (N1990, N1985, N1013);
not NOT1 (N1991, N1988);
nor NOR2 (N1992, N1970, N330);
xor XOR2 (N1993, N1987, N1397);
nand NAND4 (N1994, N1993, N1666, N1153, N1286);
buf BUF1 (N1995, N1938);
buf BUF1 (N1996, N1994);
not NOT1 (N1997, N1983);
not NOT1 (N1998, N1981);
nor NOR3 (N1999, N1989, N1886, N1020);
nor NOR4 (N2000, N1999, N1882, N1537, N1562);
and AND4 (N2001, N1998, N949, N1354, N695);
and AND4 (N2002, N1986, N639, N1089, N160);
nor NOR4 (N2003, N1997, N1640, N1056, N1437);
nor NOR3 (N2004, N1992, N647, N636);
nor NOR3 (N2005, N1991, N1385, N1471);
nand NAND4 (N2006, N1978, N786, N963, N861);
and AND4 (N2007, N2000, N211, N1661, N308);
nand NAND2 (N2008, N2003, N912);
buf BUF1 (N2009, N2001);
and AND3 (N2010, N1996, N1103, N1165);
and AND3 (N2011, N2002, N58, N656);
not NOT1 (N2012, N2006);
not NOT1 (N2013, N2008);
xor XOR2 (N2014, N1995, N1607);
nand NAND2 (N2015, N2013, N301);
buf BUF1 (N2016, N2014);
nor NOR2 (N2017, N1990, N458);
and AND4 (N2018, N2005, N1907, N719, N1573);
nor NOR3 (N2019, N2009, N1658, N1402);
not NOT1 (N2020, N2007);
nor NOR2 (N2021, N2010, N686);
not NOT1 (N2022, N2012);
buf BUF1 (N2023, N2018);
xor XOR2 (N2024, N2011, N1853);
buf BUF1 (N2025, N2019);
nand NAND3 (N2026, N2004, N1320, N487);
buf BUF1 (N2027, N2022);
nor NOR3 (N2028, N2025, N321, N1604);
nand NAND3 (N2029, N2026, N2028, N705);
xor XOR2 (N2030, N1285, N1124);
nor NOR2 (N2031, N2015, N1726);
nand NAND2 (N2032, N2016, N1297);
and AND4 (N2033, N2024, N1922, N1263, N1231);
not NOT1 (N2034, N2027);
xor XOR2 (N2035, N2034, N1375);
nor NOR3 (N2036, N2021, N1901, N1184);
not NOT1 (N2037, N2023);
not NOT1 (N2038, N2030);
nor NOR4 (N2039, N2037, N597, N224, N1659);
nor NOR4 (N2040, N2035, N561, N6, N470);
xor XOR2 (N2041, N2038, N896);
buf BUF1 (N2042, N2020);
or OR2 (N2043, N2029, N1813);
nand NAND3 (N2044, N2039, N985, N607);
and AND3 (N2045, N2031, N136, N1420);
and AND4 (N2046, N2043, N70, N1470, N1181);
not NOT1 (N2047, N2046);
not NOT1 (N2048, N2036);
buf BUF1 (N2049, N2044);
and AND2 (N2050, N2045, N244);
not NOT1 (N2051, N2049);
xor XOR2 (N2052, N2040, N1971);
buf BUF1 (N2053, N2032);
and AND3 (N2054, N2050, N1983, N1134);
nor NOR3 (N2055, N2052, N1453, N1702);
nor NOR4 (N2056, N2041, N1840, N1298, N1703);
buf BUF1 (N2057, N2054);
not NOT1 (N2058, N2042);
or OR3 (N2059, N2048, N1814, N1720);
and AND2 (N2060, N2057, N1738);
buf BUF1 (N2061, N2047);
xor XOR2 (N2062, N2060, N371);
not NOT1 (N2063, N2053);
xor XOR2 (N2064, N2058, N169);
nand NAND2 (N2065, N2061, N799);
xor XOR2 (N2066, N2051, N635);
nor NOR4 (N2067, N2062, N1515, N1461, N1689);
xor XOR2 (N2068, N2017, N1180);
xor XOR2 (N2069, N2059, N1892);
not NOT1 (N2070, N2069);
nor NOR4 (N2071, N2066, N1970, N524, N298);
xor XOR2 (N2072, N2065, N1080);
and AND2 (N2073, N2071, N1477);
or OR3 (N2074, N2056, N441, N2006);
xor XOR2 (N2075, N2074, N247);
xor XOR2 (N2076, N2073, N815);
nor NOR4 (N2077, N2076, N1573, N874, N1606);
or OR4 (N2078, N2075, N1503, N232, N1630);
or OR3 (N2079, N2033, N1174, N457);
or OR2 (N2080, N2063, N727);
nor NOR4 (N2081, N2064, N561, N1007, N2049);
not NOT1 (N2082, N2055);
or OR2 (N2083, N2077, N1283);
nand NAND4 (N2084, N2080, N1874, N1759, N1258);
nor NOR2 (N2085, N2072, N1409);
or OR3 (N2086, N2067, N780, N867);
not NOT1 (N2087, N2081);
or OR2 (N2088, N2086, N1690);
not NOT1 (N2089, N2083);
or OR2 (N2090, N2078, N1965);
buf BUF1 (N2091, N2079);
buf BUF1 (N2092, N2090);
not NOT1 (N2093, N2084);
buf BUF1 (N2094, N2087);
nand NAND2 (N2095, N2091, N1471);
or OR2 (N2096, N2089, N1137);
buf BUF1 (N2097, N2092);
buf BUF1 (N2098, N2097);
and AND2 (N2099, N2082, N1244);
nor NOR4 (N2100, N2095, N1961, N542, N1801);
and AND4 (N2101, N2085, N670, N2, N2055);
nand NAND2 (N2102, N2098, N1876);
and AND2 (N2103, N2094, N501);
xor XOR2 (N2104, N2088, N116);
nor NOR4 (N2105, N2093, N1256, N1343, N147);
nor NOR2 (N2106, N2096, N688);
buf BUF1 (N2107, N2103);
nand NAND3 (N2108, N2105, N1893, N1170);
nor NOR4 (N2109, N2068, N1968, N1197, N1262);
not NOT1 (N2110, N2104);
and AND4 (N2111, N2108, N1632, N21, N1890);
not NOT1 (N2112, N2101);
buf BUF1 (N2113, N2107);
xor XOR2 (N2114, N2099, N573);
or OR3 (N2115, N2110, N748, N1697);
and AND2 (N2116, N2113, N499);
nand NAND2 (N2117, N2102, N11);
and AND2 (N2118, N2116, N1344);
nand NAND4 (N2119, N2114, N581, N1704, N1858);
nor NOR4 (N2120, N2070, N270, N1439, N1656);
and AND3 (N2121, N2119, N1992, N1832);
nand NAND3 (N2122, N2118, N1658, N2095);
and AND4 (N2123, N2115, N1097, N391, N1236);
nand NAND3 (N2124, N2112, N689, N110);
not NOT1 (N2125, N2121);
xor XOR2 (N2126, N2117, N1131);
not NOT1 (N2127, N2106);
or OR4 (N2128, N2111, N1162, N143, N456);
nor NOR4 (N2129, N2120, N788, N1929, N1814);
xor XOR2 (N2130, N2129, N385);
xor XOR2 (N2131, N2123, N389);
and AND4 (N2132, N2124, N1675, N215, N1642);
and AND4 (N2133, N2128, N975, N1091, N1689);
or OR3 (N2134, N2133, N1361, N511);
nand NAND3 (N2135, N2131, N454, N1316);
nand NAND4 (N2136, N2130, N30, N2107, N1043);
nor NOR2 (N2137, N2135, N1589);
xor XOR2 (N2138, N2132, N492);
nand NAND2 (N2139, N2127, N1301);
nand NAND2 (N2140, N2122, N1091);
and AND4 (N2141, N2100, N30, N859, N714);
xor XOR2 (N2142, N2109, N1442);
or OR2 (N2143, N2141, N1021);
or OR4 (N2144, N2136, N944, N1717, N2089);
buf BUF1 (N2145, N2139);
buf BUF1 (N2146, N2145);
nor NOR2 (N2147, N2126, N1793);
and AND3 (N2148, N2142, N1189, N910);
xor XOR2 (N2149, N2138, N1279);
buf BUF1 (N2150, N2146);
xor XOR2 (N2151, N2149, N1589);
not NOT1 (N2152, N2143);
xor XOR2 (N2153, N2137, N2090);
nor NOR2 (N2154, N2134, N1476);
not NOT1 (N2155, N2148);
and AND4 (N2156, N2150, N265, N767, N713);
or OR2 (N2157, N2147, N689);
nand NAND4 (N2158, N2156, N1618, N1710, N671);
or OR2 (N2159, N2155, N546);
xor XOR2 (N2160, N2144, N366);
nand NAND2 (N2161, N2157, N1003);
xor XOR2 (N2162, N2125, N270);
xor XOR2 (N2163, N2140, N2103);
and AND3 (N2164, N2153, N1588, N1579);
xor XOR2 (N2165, N2162, N2053);
nand NAND4 (N2166, N2152, N1397, N1092, N933);
buf BUF1 (N2167, N2151);
and AND3 (N2168, N2154, N276, N43);
xor XOR2 (N2169, N2160, N635);
buf BUF1 (N2170, N2165);
nand NAND2 (N2171, N2164, N380);
buf BUF1 (N2172, N2170);
not NOT1 (N2173, N2172);
and AND3 (N2174, N2158, N1785, N944);
buf BUF1 (N2175, N2168);
nor NOR2 (N2176, N2171, N71);
or OR3 (N2177, N2161, N1994, N1441);
and AND2 (N2178, N2176, N1013);
xor XOR2 (N2179, N2169, N1424);
and AND4 (N2180, N2166, N1742, N741, N2112);
and AND4 (N2181, N2177, N1436, N1194, N620);
nor NOR2 (N2182, N2180, N1738);
and AND3 (N2183, N2175, N772, N799);
not NOT1 (N2184, N2178);
or OR3 (N2185, N2179, N471, N1991);
nand NAND4 (N2186, N2167, N1072, N328, N193);
nor NOR3 (N2187, N2159, N914, N1297);
nand NAND3 (N2188, N2182, N1044, N122);
nor NOR2 (N2189, N2185, N232);
and AND2 (N2190, N2173, N756);
or OR2 (N2191, N2163, N1988);
nor NOR2 (N2192, N2174, N1266);
nor NOR4 (N2193, N2192, N400, N377, N38);
not NOT1 (N2194, N2187);
nor NOR2 (N2195, N2186, N398);
xor XOR2 (N2196, N2193, N886);
not NOT1 (N2197, N2188);
buf BUF1 (N2198, N2190);
and AND4 (N2199, N2196, N622, N463, N518);
xor XOR2 (N2200, N2198, N2019);
xor XOR2 (N2201, N2189, N437);
not NOT1 (N2202, N2184);
nor NOR4 (N2203, N2200, N422, N1157, N1360);
xor XOR2 (N2204, N2203, N405);
or OR2 (N2205, N2197, N338);
and AND2 (N2206, N2195, N1729);
nand NAND4 (N2207, N2181, N1661, N1401, N1341);
buf BUF1 (N2208, N2191);
and AND3 (N2209, N2199, N821, N402);
and AND4 (N2210, N2183, N235, N913, N1492);
or OR4 (N2211, N2205, N1295, N17, N463);
and AND3 (N2212, N2211, N1374, N243);
xor XOR2 (N2213, N2202, N683);
nor NOR3 (N2214, N2212, N1582, N1129);
buf BUF1 (N2215, N2208);
not NOT1 (N2216, N2207);
xor XOR2 (N2217, N2214, N1248);
and AND3 (N2218, N2209, N176, N931);
nand NAND4 (N2219, N2218, N432, N1410, N1308);
xor XOR2 (N2220, N2217, N660);
nand NAND3 (N2221, N2210, N399, N1944);
or OR4 (N2222, N2220, N996, N1206, N1625);
nand NAND2 (N2223, N2219, N1507);
or OR2 (N2224, N2194, N2051);
or OR2 (N2225, N2204, N76);
not NOT1 (N2226, N2213);
xor XOR2 (N2227, N2221, N829);
not NOT1 (N2228, N2206);
and AND3 (N2229, N2224, N229, N2223);
or OR4 (N2230, N784, N264, N851, N323);
xor XOR2 (N2231, N2229, N896);
not NOT1 (N2232, N2230);
nor NOR3 (N2233, N2226, N1727, N41);
nor NOR3 (N2234, N2233, N685, N1057);
nor NOR4 (N2235, N2225, N309, N1570, N225);
and AND2 (N2236, N2232, N1879);
not NOT1 (N2237, N2201);
nor NOR4 (N2238, N2216, N1562, N1142, N741);
buf BUF1 (N2239, N2237);
nor NOR2 (N2240, N2231, N1203);
or OR3 (N2241, N2238, N1221, N1377);
buf BUF1 (N2242, N2215);
and AND2 (N2243, N2227, N542);
nand NAND4 (N2244, N2235, N1927, N48, N2006);
not NOT1 (N2245, N2241);
nand NAND2 (N2246, N2242, N2095);
not NOT1 (N2247, N2244);
and AND2 (N2248, N2234, N564);
buf BUF1 (N2249, N2245);
buf BUF1 (N2250, N2243);
or OR3 (N2251, N2248, N286, N2042);
xor XOR2 (N2252, N2240, N183);
buf BUF1 (N2253, N2252);
buf BUF1 (N2254, N2236);
or OR2 (N2255, N2228, N1216);
or OR4 (N2256, N2254, N2130, N1864, N1358);
buf BUF1 (N2257, N2247);
nand NAND3 (N2258, N2255, N871, N863);
nor NOR2 (N2259, N2251, N1096);
not NOT1 (N2260, N2256);
nand NAND2 (N2261, N2250, N1156);
not NOT1 (N2262, N2246);
not NOT1 (N2263, N2258);
buf BUF1 (N2264, N2257);
and AND3 (N2265, N2249, N905, N592);
xor XOR2 (N2266, N2263, N937);
not NOT1 (N2267, N2262);
xor XOR2 (N2268, N2222, N1166);
and AND4 (N2269, N2261, N491, N803, N2142);
not NOT1 (N2270, N2253);
buf BUF1 (N2271, N2270);
nor NOR3 (N2272, N2266, N1437, N223);
and AND3 (N2273, N2272, N956, N686);
xor XOR2 (N2274, N2239, N977);
nand NAND2 (N2275, N2268, N1998);
or OR4 (N2276, N2259, N1434, N1125, N1970);
or OR3 (N2277, N2267, N1511, N1747);
xor XOR2 (N2278, N2265, N773);
xor XOR2 (N2279, N2276, N481);
nand NAND4 (N2280, N2275, N1887, N892, N579);
and AND3 (N2281, N2271, N2120, N587);
xor XOR2 (N2282, N2279, N735);
buf BUF1 (N2283, N2273);
nor NOR3 (N2284, N2264, N1759, N76);
nor NOR3 (N2285, N2274, N1465, N1269);
or OR3 (N2286, N2282, N891, N2186);
not NOT1 (N2287, N2269);
and AND3 (N2288, N2287, N1048, N1682);
not NOT1 (N2289, N2260);
and AND4 (N2290, N2278, N541, N750, N1101);
xor XOR2 (N2291, N2277, N1426);
nor NOR3 (N2292, N2290, N1825, N1848);
or OR2 (N2293, N2284, N724);
not NOT1 (N2294, N2283);
xor XOR2 (N2295, N2285, N1987);
not NOT1 (N2296, N2292);
not NOT1 (N2297, N2281);
or OR3 (N2298, N2293, N522, N1836);
nand NAND4 (N2299, N2289, N462, N447, N900);
and AND3 (N2300, N2296, N20, N371);
xor XOR2 (N2301, N2295, N623);
or OR3 (N2302, N2301, N1841, N832);
xor XOR2 (N2303, N2298, N809);
nand NAND4 (N2304, N2288, N2203, N841, N1888);
xor XOR2 (N2305, N2300, N782);
and AND3 (N2306, N2302, N836, N385);
buf BUF1 (N2307, N2299);
or OR3 (N2308, N2291, N1915, N175);
nor NOR4 (N2309, N2306, N2228, N752, N1497);
not NOT1 (N2310, N2307);
xor XOR2 (N2311, N2304, N43);
nor NOR2 (N2312, N2310, N434);
or OR4 (N2313, N2286, N1457, N1172, N231);
or OR4 (N2314, N2309, N2181, N1669, N940);
or OR4 (N2315, N2312, N1014, N232, N117);
and AND3 (N2316, N2297, N2291, N1633);
xor XOR2 (N2317, N2308, N1160);
and AND3 (N2318, N2305, N2268, N2110);
nor NOR2 (N2319, N2311, N2075);
nor NOR3 (N2320, N2315, N96, N1554);
nor NOR4 (N2321, N2317, N1682, N1861, N1866);
buf BUF1 (N2322, N2313);
not NOT1 (N2323, N2322);
nor NOR4 (N2324, N2314, N1519, N615, N1672);
nand NAND2 (N2325, N2318, N698);
and AND2 (N2326, N2280, N1812);
not NOT1 (N2327, N2325);
xor XOR2 (N2328, N2294, N2325);
or OR2 (N2329, N2319, N1241);
buf BUF1 (N2330, N2326);
not NOT1 (N2331, N2327);
nor NOR3 (N2332, N2320, N1215, N1443);
and AND3 (N2333, N2324, N669, N103);
and AND4 (N2334, N2316, N1822, N2307, N659);
xor XOR2 (N2335, N2321, N1834);
or OR2 (N2336, N2329, N575);
nor NOR2 (N2337, N2332, N1792);
nand NAND2 (N2338, N2303, N1302);
or OR2 (N2339, N2331, N1554);
not NOT1 (N2340, N2323);
not NOT1 (N2341, N2339);
not NOT1 (N2342, N2333);
and AND4 (N2343, N2336, N59, N197, N429);
and AND2 (N2344, N2328, N392);
or OR3 (N2345, N2340, N1130, N418);
nand NAND3 (N2346, N2335, N702, N1972);
nor NOR2 (N2347, N2344, N212);
buf BUF1 (N2348, N2337);
nand NAND4 (N2349, N2345, N51, N300, N1598);
not NOT1 (N2350, N2349);
xor XOR2 (N2351, N2347, N2173);
and AND2 (N2352, N2338, N1780);
and AND4 (N2353, N2350, N368, N899, N1372);
xor XOR2 (N2354, N2341, N2053);
nor NOR2 (N2355, N2351, N1200);
buf BUF1 (N2356, N2354);
buf BUF1 (N2357, N2346);
buf BUF1 (N2358, N2355);
and AND3 (N2359, N2330, N850, N1023);
buf BUF1 (N2360, N2358);
nand NAND2 (N2361, N2334, N1616);
nand NAND2 (N2362, N2359, N1211);
xor XOR2 (N2363, N2357, N1355);
xor XOR2 (N2364, N2353, N1321);
and AND4 (N2365, N2352, N1236, N211, N1488);
not NOT1 (N2366, N2360);
not NOT1 (N2367, N2356);
not NOT1 (N2368, N2367);
and AND3 (N2369, N2343, N1146, N2115);
buf BUF1 (N2370, N2363);
and AND2 (N2371, N2361, N1968);
buf BUF1 (N2372, N2364);
not NOT1 (N2373, N2371);
xor XOR2 (N2374, N2373, N1684);
buf BUF1 (N2375, N2374);
or OR2 (N2376, N2365, N1914);
nand NAND4 (N2377, N2362, N138, N233, N696);
nand NAND2 (N2378, N2370, N1279);
buf BUF1 (N2379, N2372);
nor NOR4 (N2380, N2342, N657, N451, N316);
xor XOR2 (N2381, N2366, N237);
nand NAND4 (N2382, N2377, N2145, N2228, N1930);
xor XOR2 (N2383, N2379, N1996);
xor XOR2 (N2384, N2368, N926);
nand NAND3 (N2385, N2369, N1729, N88);
buf BUF1 (N2386, N2375);
buf BUF1 (N2387, N2380);
xor XOR2 (N2388, N2387, N1797);
and AND3 (N2389, N2383, N1100, N1675);
nand NAND3 (N2390, N2376, N754, N712);
buf BUF1 (N2391, N2381);
xor XOR2 (N2392, N2388, N334);
not NOT1 (N2393, N2391);
xor XOR2 (N2394, N2390, N1196);
not NOT1 (N2395, N2389);
nor NOR2 (N2396, N2386, N451);
nor NOR4 (N2397, N2384, N2036, N73, N216);
nand NAND2 (N2398, N2394, N151);
nand NAND2 (N2399, N2398, N943);
nand NAND3 (N2400, N2378, N1475, N509);
xor XOR2 (N2401, N2382, N1074);
xor XOR2 (N2402, N2393, N1012);
buf BUF1 (N2403, N2400);
or OR4 (N2404, N2396, N803, N2103, N810);
and AND4 (N2405, N2402, N1256, N495, N2079);
and AND3 (N2406, N2405, N1072, N1147);
xor XOR2 (N2407, N2404, N2333);
and AND2 (N2408, N2392, N1326);
nand NAND3 (N2409, N2397, N886, N545);
not NOT1 (N2410, N2407);
nand NAND2 (N2411, N2408, N1961);
nor NOR3 (N2412, N2348, N350, N2140);
nand NAND2 (N2413, N2409, N1076);
not NOT1 (N2414, N2412);
not NOT1 (N2415, N2410);
and AND4 (N2416, N2399, N2411, N954, N65);
not NOT1 (N2417, N1796);
and AND4 (N2418, N2385, N422, N945, N1633);
and AND3 (N2419, N2414, N1769, N1321);
xor XOR2 (N2420, N2419, N587);
or OR4 (N2421, N2401, N912, N992, N1303);
nand NAND3 (N2422, N2403, N488, N1140);
nand NAND3 (N2423, N2420, N917, N1777);
xor XOR2 (N2424, N2415, N1155);
buf BUF1 (N2425, N2418);
nand NAND4 (N2426, N2416, N1908, N2387, N1440);
or OR2 (N2427, N2413, N2249);
or OR3 (N2428, N2406, N1634, N2269);
and AND4 (N2429, N2427, N2274, N96, N1135);
buf BUF1 (N2430, N2422);
buf BUF1 (N2431, N2421);
and AND4 (N2432, N2429, N41, N1421, N2394);
not NOT1 (N2433, N2426);
xor XOR2 (N2434, N2432, N968);
nand NAND2 (N2435, N2431, N467);
not NOT1 (N2436, N2417);
and AND2 (N2437, N2428, N2235);
nor NOR2 (N2438, N2424, N1228);
nor NOR2 (N2439, N2438, N1912);
nor NOR2 (N2440, N2430, N1543);
buf BUF1 (N2441, N2433);
xor XOR2 (N2442, N2395, N66);
nand NAND4 (N2443, N2442, N734, N1288, N1068);
nor NOR4 (N2444, N2434, N2112, N301, N1089);
buf BUF1 (N2445, N2423);
buf BUF1 (N2446, N2436);
nor NOR3 (N2447, N2443, N277, N962);
nand NAND2 (N2448, N2425, N1168);
nor NOR3 (N2449, N2444, N1667, N965);
nand NAND4 (N2450, N2449, N1034, N764, N2184);
buf BUF1 (N2451, N2446);
or OR4 (N2452, N2435, N2223, N1456, N1077);
nor NOR4 (N2453, N2439, N1574, N2199, N1882);
or OR2 (N2454, N2453, N869);
nor NOR4 (N2455, N2450, N1234, N638, N1051);
and AND3 (N2456, N2455, N462, N2164);
or OR4 (N2457, N2440, N482, N1791, N1097);
xor XOR2 (N2458, N2451, N1061);
nor NOR2 (N2459, N2441, N2120);
buf BUF1 (N2460, N2457);
or OR2 (N2461, N2458, N235);
and AND4 (N2462, N2447, N2276, N468, N1159);
buf BUF1 (N2463, N2448);
buf BUF1 (N2464, N2462);
xor XOR2 (N2465, N2464, N992);
or OR2 (N2466, N2454, N290);
not NOT1 (N2467, N2465);
xor XOR2 (N2468, N2437, N1914);
buf BUF1 (N2469, N2461);
xor XOR2 (N2470, N2460, N1811);
not NOT1 (N2471, N2445);
nand NAND2 (N2472, N2463, N1731);
nand NAND3 (N2473, N2471, N1933, N579);
xor XOR2 (N2474, N2467, N60);
or OR3 (N2475, N2459, N232, N294);
nand NAND3 (N2476, N2472, N770, N1826);
nand NAND2 (N2477, N2466, N2205);
not NOT1 (N2478, N2456);
and AND3 (N2479, N2469, N621, N1917);
xor XOR2 (N2480, N2478, N2046);
and AND3 (N2481, N2470, N305, N1523);
not NOT1 (N2482, N2476);
and AND4 (N2483, N2480, N826, N1712, N1756);
and AND3 (N2484, N2475, N2036, N1003);
xor XOR2 (N2485, N2452, N2087);
and AND2 (N2486, N2474, N2413);
nand NAND2 (N2487, N2486, N1342);
nand NAND4 (N2488, N2484, N1948, N477, N2068);
or OR3 (N2489, N2485, N1673, N1897);
nand NAND2 (N2490, N2487, N1070);
or OR4 (N2491, N2482, N555, N1810, N92);
xor XOR2 (N2492, N2477, N1248);
or OR4 (N2493, N2479, N2066, N2374, N622);
or OR4 (N2494, N2488, N1528, N1797, N2392);
and AND2 (N2495, N2483, N872);
nor NOR3 (N2496, N2489, N1440, N604);
nand NAND3 (N2497, N2493, N2130, N1289);
nor NOR2 (N2498, N2496, N671);
nor NOR3 (N2499, N2473, N1602, N1526);
buf BUF1 (N2500, N2499);
and AND2 (N2501, N2492, N2427);
and AND4 (N2502, N2481, N1317, N1502, N1701);
xor XOR2 (N2503, N2501, N2336);
not NOT1 (N2504, N2495);
xor XOR2 (N2505, N2494, N323);
xor XOR2 (N2506, N2500, N1055);
not NOT1 (N2507, N2502);
xor XOR2 (N2508, N2507, N1112);
xor XOR2 (N2509, N2498, N1541);
xor XOR2 (N2510, N2509, N714);
buf BUF1 (N2511, N2503);
buf BUF1 (N2512, N2497);
or OR4 (N2513, N2512, N1888, N1166, N212);
nand NAND4 (N2514, N2490, N1327, N2084, N1511);
buf BUF1 (N2515, N2504);
and AND3 (N2516, N2468, N1012, N283);
nand NAND2 (N2517, N2491, N601);
nor NOR2 (N2518, N2517, N101);
nor NOR2 (N2519, N2515, N64);
endmodule