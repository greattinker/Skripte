// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18;

output N586,N609,N613,N606,N617,N615,N616,N604,N612,N618;

nor NOR3 (N19, N14, N18, N9);
or OR3 (N20, N10, N16, N16);
nor NOR4 (N21, N15, N5, N13, N8);
buf BUF1 (N22, N11);
and AND3 (N23, N5, N11, N19);
and AND3 (N24, N22, N14, N13);
not NOT1 (N25, N5);
nor NOR2 (N26, N25, N20);
nor NOR3 (N27, N9, N23, N17);
or OR4 (N28, N8, N19, N4, N9);
or OR4 (N29, N8, N2, N2, N22);
buf BUF1 (N30, N28);
xor XOR2 (N31, N7, N24);
nand NAND4 (N32, N1, N18, N8, N17);
and AND3 (N33, N14, N25, N17);
and AND4 (N34, N3, N23, N21, N26);
nor NOR4 (N35, N18, N9, N1, N2);
and AND4 (N36, N20, N1, N23, N26);
not NOT1 (N37, N21);
buf BUF1 (N38, N33);
buf BUF1 (N39, N36);
and AND2 (N40, N27, N23);
nand NAND2 (N41, N31, N16);
nor NOR2 (N42, N41, N30);
not NOT1 (N43, N19);
buf BUF1 (N44, N32);
nand NAND4 (N45, N42, N39, N42, N3);
buf BUF1 (N46, N14);
not NOT1 (N47, N45);
xor XOR2 (N48, N44, N12);
buf BUF1 (N49, N48);
or OR2 (N50, N47, N40);
and AND2 (N51, N20, N38);
buf BUF1 (N52, N19);
not NOT1 (N53, N50);
or OR2 (N54, N49, N38);
xor XOR2 (N55, N54, N28);
nor NOR2 (N56, N37, N8);
and AND4 (N57, N46, N5, N54, N2);
not NOT1 (N58, N35);
and AND2 (N59, N29, N28);
nor NOR4 (N60, N59, N2, N25, N44);
buf BUF1 (N61, N43);
nand NAND3 (N62, N55, N36, N26);
not NOT1 (N63, N34);
and AND4 (N64, N58, N17, N10, N20);
or OR4 (N65, N56, N50, N39, N38);
nand NAND3 (N66, N62, N9, N54);
xor XOR2 (N67, N64, N49);
xor XOR2 (N68, N65, N43);
or OR2 (N69, N51, N43);
and AND4 (N70, N53, N11, N19, N21);
or OR2 (N71, N57, N47);
not NOT1 (N72, N66);
and AND2 (N73, N60, N26);
and AND2 (N74, N67, N55);
xor XOR2 (N75, N63, N17);
and AND2 (N76, N75, N59);
not NOT1 (N77, N52);
xor XOR2 (N78, N68, N59);
xor XOR2 (N79, N61, N78);
nand NAND3 (N80, N79, N16, N3);
or OR2 (N81, N8, N35);
not NOT1 (N82, N71);
nand NAND3 (N83, N69, N66, N27);
not NOT1 (N84, N82);
and AND4 (N85, N74, N46, N22, N61);
and AND2 (N86, N84, N39);
buf BUF1 (N87, N85);
xor XOR2 (N88, N72, N43);
xor XOR2 (N89, N80, N33);
buf BUF1 (N90, N86);
nor NOR2 (N91, N88, N55);
and AND3 (N92, N76, N85, N46);
nor NOR4 (N93, N81, N68, N8, N85);
not NOT1 (N94, N92);
xor XOR2 (N95, N91, N71);
or OR3 (N96, N77, N43, N39);
nor NOR3 (N97, N96, N19, N70);
not NOT1 (N98, N62);
nor NOR4 (N99, N87, N85, N5, N75);
nand NAND2 (N100, N94, N49);
buf BUF1 (N101, N98);
xor XOR2 (N102, N95, N33);
buf BUF1 (N103, N93);
or OR3 (N104, N90, N77, N59);
nand NAND4 (N105, N73, N25, N80, N58);
nor NOR3 (N106, N103, N18, N55);
xor XOR2 (N107, N101, N28);
and AND3 (N108, N89, N28, N54);
not NOT1 (N109, N97);
or OR2 (N110, N108, N92);
xor XOR2 (N111, N102, N27);
and AND4 (N112, N107, N55, N88, N111);
buf BUF1 (N113, N46);
and AND4 (N114, N99, N54, N80, N44);
and AND2 (N115, N110, N99);
not NOT1 (N116, N109);
not NOT1 (N117, N83);
buf BUF1 (N118, N105);
nor NOR2 (N119, N116, N33);
or OR2 (N120, N106, N93);
xor XOR2 (N121, N104, N55);
nand NAND4 (N122, N100, N36, N50, N4);
and AND4 (N123, N121, N65, N108, N52);
and AND2 (N124, N119, N74);
xor XOR2 (N125, N115, N49);
nand NAND2 (N126, N125, N5);
nor NOR2 (N127, N123, N125);
xor XOR2 (N128, N126, N43);
nor NOR4 (N129, N112, N94, N19, N21);
nand NAND2 (N130, N113, N122);
not NOT1 (N131, N35);
buf BUF1 (N132, N131);
buf BUF1 (N133, N114);
nor NOR3 (N134, N130, N58, N131);
xor XOR2 (N135, N118, N108);
buf BUF1 (N136, N127);
and AND3 (N137, N136, N21, N117);
not NOT1 (N138, N36);
or OR4 (N139, N137, N30, N125, N29);
and AND4 (N140, N138, N138, N104, N35);
and AND4 (N141, N132, N97, N29, N63);
xor XOR2 (N142, N141, N20);
or OR2 (N143, N124, N100);
or OR4 (N144, N135, N113, N26, N119);
or OR3 (N145, N144, N20, N102);
or OR2 (N146, N128, N90);
nor NOR3 (N147, N129, N101, N127);
xor XOR2 (N148, N120, N74);
not NOT1 (N149, N140);
or OR2 (N150, N143, N17);
and AND4 (N151, N148, N94, N54, N121);
nor NOR2 (N152, N134, N70);
or OR2 (N153, N146, N68);
nand NAND3 (N154, N152, N114, N130);
or OR4 (N155, N139, N106, N24, N59);
nand NAND4 (N156, N154, N42, N23, N105);
or OR2 (N157, N147, N54);
and AND3 (N158, N151, N18, N105);
nor NOR3 (N159, N156, N148, N16);
nand NAND3 (N160, N157, N42, N32);
and AND4 (N161, N150, N6, N142, N32);
and AND2 (N162, N5, N86);
and AND4 (N163, N162, N58, N52, N141);
xor XOR2 (N164, N158, N113);
xor XOR2 (N165, N155, N155);
xor XOR2 (N166, N160, N31);
nand NAND3 (N167, N164, N95, N32);
nand NAND2 (N168, N153, N51);
nor NOR4 (N169, N165, N88, N60, N131);
not NOT1 (N170, N167);
nand NAND2 (N171, N145, N25);
nand NAND4 (N172, N170, N150, N103, N134);
buf BUF1 (N173, N172);
nand NAND2 (N174, N169, N96);
not NOT1 (N175, N174);
nand NAND4 (N176, N163, N73, N106, N127);
xor XOR2 (N177, N161, N113);
or OR2 (N178, N159, N37);
and AND3 (N179, N173, N26, N176);
nand NAND4 (N180, N59, N178, N87, N109);
xor XOR2 (N181, N110, N10);
xor XOR2 (N182, N180, N133);
and AND4 (N183, N5, N167, N95, N119);
not NOT1 (N184, N166);
nor NOR2 (N185, N168, N132);
not NOT1 (N186, N185);
not NOT1 (N187, N183);
nor NOR2 (N188, N181, N178);
xor XOR2 (N189, N177, N150);
buf BUF1 (N190, N171);
and AND4 (N191, N187, N157, N95, N129);
nand NAND3 (N192, N175, N106, N30);
buf BUF1 (N193, N184);
buf BUF1 (N194, N190);
not NOT1 (N195, N149);
buf BUF1 (N196, N191);
and AND3 (N197, N196, N178, N67);
buf BUF1 (N198, N189);
xor XOR2 (N199, N188, N36);
nand NAND2 (N200, N194, N72);
or OR3 (N201, N179, N189, N68);
and AND4 (N202, N198, N148, N132, N101);
nor NOR4 (N203, N192, N22, N33, N87);
buf BUF1 (N204, N200);
buf BUF1 (N205, N203);
nand NAND2 (N206, N199, N19);
buf BUF1 (N207, N205);
nor NOR4 (N208, N207, N16, N31, N181);
and AND4 (N209, N193, N106, N167, N199);
buf BUF1 (N210, N186);
and AND3 (N211, N182, N11, N67);
buf BUF1 (N212, N204);
not NOT1 (N213, N209);
buf BUF1 (N214, N208);
nor NOR3 (N215, N201, N180, N104);
or OR2 (N216, N195, N156);
buf BUF1 (N217, N215);
not NOT1 (N218, N210);
buf BUF1 (N219, N218);
not NOT1 (N220, N219);
buf BUF1 (N221, N216);
and AND4 (N222, N220, N21, N12, N43);
not NOT1 (N223, N206);
nor NOR3 (N224, N222, N217, N39);
and AND4 (N225, N14, N145, N62, N216);
and AND2 (N226, N197, N2);
nor NOR3 (N227, N226, N78, N81);
buf BUF1 (N228, N223);
nor NOR2 (N229, N202, N86);
not NOT1 (N230, N227);
xor XOR2 (N231, N224, N206);
xor XOR2 (N232, N212, N148);
or OR2 (N233, N229, N168);
buf BUF1 (N234, N211);
nor NOR3 (N235, N225, N67, N45);
nand NAND3 (N236, N235, N35, N82);
not NOT1 (N237, N230);
not NOT1 (N238, N231);
and AND2 (N239, N232, N140);
xor XOR2 (N240, N214, N28);
nor NOR4 (N241, N228, N8, N84, N44);
nand NAND4 (N242, N234, N85, N21, N11);
nor NOR3 (N243, N213, N109, N195);
buf BUF1 (N244, N242);
nand NAND4 (N245, N243, N46, N166, N156);
not NOT1 (N246, N221);
buf BUF1 (N247, N245);
buf BUF1 (N248, N233);
nand NAND3 (N249, N246, N62, N231);
buf BUF1 (N250, N249);
and AND2 (N251, N239, N220);
and AND2 (N252, N236, N191);
or OR3 (N253, N240, N234, N144);
or OR4 (N254, N253, N221, N30, N201);
nor NOR4 (N255, N238, N107, N168, N182);
and AND4 (N256, N255, N77, N70, N152);
not NOT1 (N257, N248);
not NOT1 (N258, N251);
not NOT1 (N259, N258);
and AND3 (N260, N257, N172, N174);
buf BUF1 (N261, N259);
not NOT1 (N262, N254);
and AND2 (N263, N250, N148);
and AND2 (N264, N252, N57);
buf BUF1 (N265, N263);
nand NAND4 (N266, N265, N221, N184, N17);
not NOT1 (N267, N262);
or OR2 (N268, N260, N229);
buf BUF1 (N269, N237);
buf BUF1 (N270, N266);
nand NAND2 (N271, N267, N244);
nor NOR4 (N272, N96, N217, N206, N186);
xor XOR2 (N273, N272, N21);
and AND2 (N274, N256, N77);
or OR2 (N275, N247, N253);
nor NOR3 (N276, N271, N142, N1);
buf BUF1 (N277, N241);
not NOT1 (N278, N261);
nand NAND2 (N279, N278, N230);
nand NAND3 (N280, N270, N277, N214);
buf BUF1 (N281, N89);
or OR3 (N282, N269, N237, N218);
and AND3 (N283, N282, N86, N211);
nor NOR3 (N284, N273, N257, N144);
xor XOR2 (N285, N264, N215);
nand NAND4 (N286, N280, N70, N265, N178);
nand NAND3 (N287, N285, N182, N153);
and AND4 (N288, N284, N153, N255, N107);
and AND4 (N289, N281, N209, N252, N23);
nor NOR3 (N290, N287, N236, N220);
not NOT1 (N291, N275);
or OR2 (N292, N279, N242);
buf BUF1 (N293, N288);
not NOT1 (N294, N276);
nand NAND2 (N295, N294, N95);
nand NAND2 (N296, N289, N105);
or OR4 (N297, N274, N199, N106, N116);
not NOT1 (N298, N295);
nor NOR4 (N299, N291, N28, N193, N225);
buf BUF1 (N300, N268);
and AND4 (N301, N299, N258, N248, N230);
not NOT1 (N302, N293);
xor XOR2 (N303, N296, N196);
or OR3 (N304, N292, N130, N188);
not NOT1 (N305, N301);
nand NAND2 (N306, N298, N292);
nand NAND4 (N307, N302, N212, N184, N70);
not NOT1 (N308, N304);
and AND3 (N309, N306, N72, N213);
buf BUF1 (N310, N300);
buf BUF1 (N311, N290);
or OR4 (N312, N311, N215, N280, N151);
xor XOR2 (N313, N297, N286);
or OR2 (N314, N246, N200);
and AND4 (N315, N308, N114, N160, N190);
nand NAND4 (N316, N307, N40, N6, N108);
not NOT1 (N317, N283);
buf BUF1 (N318, N312);
and AND4 (N319, N309, N283, N190, N316);
or OR2 (N320, N242, N229);
and AND4 (N321, N310, N101, N283, N110);
buf BUF1 (N322, N318);
nand NAND2 (N323, N321, N174);
buf BUF1 (N324, N305);
nor NOR2 (N325, N313, N243);
and AND4 (N326, N319, N21, N131, N315);
buf BUF1 (N327, N271);
or OR3 (N328, N325, N21, N314);
or OR3 (N329, N93, N55, N89);
xor XOR2 (N330, N320, N121);
nor NOR2 (N331, N303, N165);
and AND4 (N332, N326, N327, N51, N155);
and AND2 (N333, N254, N64);
not NOT1 (N334, N328);
or OR4 (N335, N317, N317, N334, N300);
or OR2 (N336, N316, N237);
or OR3 (N337, N323, N22, N65);
nor NOR2 (N338, N333, N158);
nand NAND3 (N339, N336, N12, N141);
xor XOR2 (N340, N335, N268);
not NOT1 (N341, N331);
buf BUF1 (N342, N338);
not NOT1 (N343, N324);
xor XOR2 (N344, N322, N295);
and AND4 (N345, N340, N93, N173, N83);
xor XOR2 (N346, N337, N247);
buf BUF1 (N347, N345);
and AND2 (N348, N347, N202);
not NOT1 (N349, N329);
nand NAND3 (N350, N342, N258, N156);
buf BUF1 (N351, N346);
not NOT1 (N352, N343);
and AND4 (N353, N332, N69, N151, N223);
buf BUF1 (N354, N353);
or OR4 (N355, N349, N226, N235, N26);
and AND4 (N356, N339, N34, N212, N284);
not NOT1 (N357, N348);
xor XOR2 (N358, N350, N85);
and AND2 (N359, N358, N72);
xor XOR2 (N360, N351, N103);
not NOT1 (N361, N354);
and AND4 (N362, N341, N95, N354, N283);
buf BUF1 (N363, N360);
and AND2 (N364, N330, N328);
or OR3 (N365, N362, N43, N284);
nor NOR3 (N366, N356, N96, N31);
buf BUF1 (N367, N357);
not NOT1 (N368, N366);
buf BUF1 (N369, N352);
nand NAND4 (N370, N363, N53, N347, N318);
xor XOR2 (N371, N344, N207);
nor NOR4 (N372, N368, N219, N261, N301);
nor NOR2 (N373, N359, N84);
xor XOR2 (N374, N361, N231);
xor XOR2 (N375, N371, N66);
nor NOR4 (N376, N370, N2, N295, N260);
nor NOR4 (N377, N376, N84, N177, N171);
xor XOR2 (N378, N375, N133);
or OR4 (N379, N377, N215, N250, N205);
and AND4 (N380, N367, N233, N343, N79);
and AND2 (N381, N372, N211);
or OR4 (N382, N378, N212, N357, N266);
nand NAND4 (N383, N365, N7, N28, N340);
or OR2 (N384, N374, N250);
nor NOR2 (N385, N369, N3);
nand NAND4 (N386, N364, N235, N38, N107);
and AND3 (N387, N385, N301, N274);
nor NOR4 (N388, N373, N89, N318, N19);
buf BUF1 (N389, N387);
nor NOR2 (N390, N388, N323);
nor NOR3 (N391, N380, N148, N22);
and AND4 (N392, N384, N211, N15, N96);
and AND2 (N393, N389, N16);
nand NAND3 (N394, N379, N216, N343);
xor XOR2 (N395, N390, N165);
or OR3 (N396, N393, N146, N71);
xor XOR2 (N397, N383, N334);
not NOT1 (N398, N392);
xor XOR2 (N399, N355, N332);
xor XOR2 (N400, N382, N225);
nor NOR3 (N401, N399, N333, N384);
or OR4 (N402, N396, N399, N166, N109);
xor XOR2 (N403, N400, N374);
or OR2 (N404, N401, N344);
nand NAND2 (N405, N381, N216);
buf BUF1 (N406, N395);
buf BUF1 (N407, N386);
and AND3 (N408, N405, N336, N67);
and AND2 (N409, N391, N368);
or OR4 (N410, N402, N99, N15, N345);
or OR4 (N411, N403, N270, N296, N334);
buf BUF1 (N412, N394);
or OR2 (N413, N398, N101);
nand NAND3 (N414, N404, N320, N85);
buf BUF1 (N415, N406);
xor XOR2 (N416, N397, N353);
buf BUF1 (N417, N414);
not NOT1 (N418, N409);
and AND4 (N419, N410, N43, N90, N410);
nand NAND4 (N420, N413, N7, N163, N222);
buf BUF1 (N421, N412);
and AND4 (N422, N417, N42, N312, N207);
not NOT1 (N423, N416);
nand NAND2 (N424, N420, N44);
or OR4 (N425, N408, N319, N171, N105);
buf BUF1 (N426, N425);
not NOT1 (N427, N422);
not NOT1 (N428, N419);
and AND2 (N429, N421, N332);
and AND3 (N430, N429, N258, N363);
buf BUF1 (N431, N418);
or OR4 (N432, N407, N313, N274, N80);
nor NOR4 (N433, N431, N196, N147, N338);
buf BUF1 (N434, N427);
or OR3 (N435, N433, N39, N372);
nor NOR4 (N436, N423, N25, N54, N124);
buf BUF1 (N437, N411);
not NOT1 (N438, N430);
nand NAND3 (N439, N435, N55, N96);
xor XOR2 (N440, N437, N267);
not NOT1 (N441, N426);
and AND2 (N442, N440, N196);
buf BUF1 (N443, N436);
or OR4 (N444, N415, N431, N309, N252);
nand NAND4 (N445, N424, N247, N266, N147);
nor NOR3 (N446, N441, N78, N49);
not NOT1 (N447, N446);
or OR3 (N448, N442, N384, N100);
and AND2 (N449, N439, N360);
nand NAND2 (N450, N432, N445);
not NOT1 (N451, N131);
buf BUF1 (N452, N450);
nand NAND4 (N453, N434, N448, N258, N149);
not NOT1 (N454, N14);
buf BUF1 (N455, N454);
nand NAND3 (N456, N447, N227, N453);
nand NAND3 (N457, N54, N440, N431);
nand NAND2 (N458, N428, N31);
not NOT1 (N459, N458);
nand NAND3 (N460, N456, N167, N59);
nand NAND3 (N461, N449, N409, N325);
nand NAND2 (N462, N459, N109);
not NOT1 (N463, N457);
nand NAND2 (N464, N462, N178);
and AND3 (N465, N451, N321, N214);
nand NAND4 (N466, N444, N127, N129, N83);
nand NAND2 (N467, N460, N249);
or OR4 (N468, N463, N20, N9, N385);
nand NAND2 (N469, N443, N305);
nor NOR4 (N470, N455, N313, N62, N285);
buf BUF1 (N471, N467);
nand NAND3 (N472, N469, N443, N401);
not NOT1 (N473, N461);
nor NOR4 (N474, N473, N376, N185, N22);
nand NAND4 (N475, N452, N397, N471, N142);
buf BUF1 (N476, N467);
nor NOR2 (N477, N468, N476);
buf BUF1 (N478, N229);
nand NAND2 (N479, N475, N109);
xor XOR2 (N480, N470, N346);
buf BUF1 (N481, N478);
nor NOR4 (N482, N477, N186, N131, N403);
nand NAND4 (N483, N438, N345, N63, N399);
nand NAND4 (N484, N481, N236, N376, N349);
or OR3 (N485, N484, N254, N313);
not NOT1 (N486, N480);
not NOT1 (N487, N485);
nor NOR2 (N488, N482, N58);
nand NAND3 (N489, N472, N445, N264);
nor NOR3 (N490, N483, N211, N456);
and AND4 (N491, N466, N436, N431, N479);
nor NOR4 (N492, N264, N118, N294, N479);
not NOT1 (N493, N489);
not NOT1 (N494, N493);
and AND4 (N495, N464, N380, N372, N236);
buf BUF1 (N496, N491);
nor NOR2 (N497, N488, N377);
nor NOR4 (N498, N490, N82, N435, N204);
nor NOR3 (N499, N487, N11, N113);
not NOT1 (N500, N497);
xor XOR2 (N501, N486, N212);
and AND3 (N502, N501, N23, N322);
nor NOR4 (N503, N502, N280, N348, N185);
or OR3 (N504, N492, N308, N26);
not NOT1 (N505, N494);
nand NAND2 (N506, N495, N214);
xor XOR2 (N507, N499, N384);
buf BUF1 (N508, N498);
xor XOR2 (N509, N505, N243);
nor NOR4 (N510, N506, N472, N375, N415);
nor NOR3 (N511, N509, N131, N249);
not NOT1 (N512, N511);
and AND2 (N513, N504, N227);
xor XOR2 (N514, N496, N409);
nor NOR3 (N515, N503, N238, N396);
and AND4 (N516, N474, N184, N333, N144);
nor NOR4 (N517, N500, N224, N109, N433);
not NOT1 (N518, N507);
buf BUF1 (N519, N512);
nand NAND2 (N520, N519, N260);
xor XOR2 (N521, N514, N408);
or OR3 (N522, N510, N175, N415);
buf BUF1 (N523, N522);
and AND2 (N524, N520, N340);
nand NAND4 (N525, N521, N125, N373, N439);
buf BUF1 (N526, N465);
and AND4 (N527, N523, N83, N287, N113);
or OR2 (N528, N518, N17);
xor XOR2 (N529, N517, N471);
nand NAND4 (N530, N525, N192, N172, N31);
nand NAND2 (N531, N515, N176);
nor NOR3 (N532, N528, N411, N182);
not NOT1 (N533, N508);
nand NAND3 (N534, N524, N285, N362);
nand NAND2 (N535, N513, N422);
and AND2 (N536, N526, N365);
nand NAND2 (N537, N534, N519);
xor XOR2 (N538, N537, N288);
nand NAND4 (N539, N538, N303, N20, N420);
or OR2 (N540, N535, N226);
and AND3 (N541, N527, N14, N57);
nand NAND2 (N542, N529, N468);
not NOT1 (N543, N540);
or OR2 (N544, N536, N216);
xor XOR2 (N545, N533, N158);
xor XOR2 (N546, N531, N467);
and AND3 (N547, N542, N502, N148);
and AND2 (N548, N547, N286);
not NOT1 (N549, N546);
or OR2 (N550, N532, N80);
buf BUF1 (N551, N530);
and AND4 (N552, N539, N72, N182, N367);
buf BUF1 (N553, N550);
nor NOR2 (N554, N545, N14);
nor NOR2 (N555, N541, N61);
nand NAND3 (N556, N554, N405, N294);
and AND2 (N557, N549, N170);
and AND4 (N558, N544, N385, N491, N34);
not NOT1 (N559, N556);
buf BUF1 (N560, N543);
nor NOR2 (N561, N548, N354);
xor XOR2 (N562, N560, N184);
buf BUF1 (N563, N553);
buf BUF1 (N564, N555);
buf BUF1 (N565, N559);
buf BUF1 (N566, N564);
nand NAND4 (N567, N562, N359, N310, N215);
or OR3 (N568, N567, N131, N347);
or OR2 (N569, N557, N351);
buf BUF1 (N570, N516);
xor XOR2 (N571, N566, N478);
and AND3 (N572, N552, N92, N503);
or OR2 (N573, N568, N186);
buf BUF1 (N574, N571);
not NOT1 (N575, N563);
not NOT1 (N576, N565);
nand NAND3 (N577, N572, N444, N434);
buf BUF1 (N578, N558);
xor XOR2 (N579, N578, N128);
xor XOR2 (N580, N570, N273);
nand NAND2 (N581, N577, N316);
and AND3 (N582, N569, N581, N379);
not NOT1 (N583, N180);
nor NOR2 (N584, N582, N94);
xor XOR2 (N585, N576, N184);
not NOT1 (N586, N584);
and AND4 (N587, N583, N61, N566, N165);
and AND3 (N588, N580, N129, N362);
nand NAND3 (N589, N575, N418, N128);
and AND4 (N590, N561, N149, N276, N142);
buf BUF1 (N591, N551);
nor NOR4 (N592, N574, N263, N169, N26);
nor NOR2 (N593, N573, N115);
nand NAND4 (N594, N587, N212, N474, N444);
and AND3 (N595, N590, N286, N518);
buf BUF1 (N596, N588);
not NOT1 (N597, N579);
nor NOR2 (N598, N589, N332);
and AND3 (N599, N594, N354, N542);
not NOT1 (N600, N598);
xor XOR2 (N601, N593, N309);
or OR2 (N602, N600, N215);
buf BUF1 (N603, N595);
not NOT1 (N604, N596);
and AND2 (N605, N592, N300);
buf BUF1 (N606, N597);
and AND3 (N607, N599, N78, N90);
and AND3 (N608, N602, N74, N50);
nand NAND4 (N609, N607, N571, N265, N67);
xor XOR2 (N610, N601, N181);
xor XOR2 (N611, N591, N264);
nand NAND4 (N612, N603, N115, N513, N521);
xor XOR2 (N613, N610, N492);
xor XOR2 (N614, N585, N114);
nor NOR2 (N615, N608, N531);
buf BUF1 (N616, N614);
xor XOR2 (N617, N611, N443);
nand NAND4 (N618, N605, N553, N472, N236);
endmodule