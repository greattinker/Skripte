// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10;

output N1003,N1009,N995,N1005,N997,N1007,N1008,N991,N1001,N1010;

nor NOR2 (N11, N4, N8);
xor XOR2 (N12, N5, N2);
xor XOR2 (N13, N12, N10);
not NOT1 (N14, N4);
buf BUF1 (N15, N1);
nand NAND2 (N16, N2, N10);
xor XOR2 (N17, N2, N14);
not NOT1 (N18, N16);
nor NOR4 (N19, N3, N4, N2, N18);
or OR2 (N20, N9, N19);
and AND4 (N21, N18, N15, N4, N8);
not NOT1 (N22, N8);
buf BUF1 (N23, N17);
buf BUF1 (N24, N14);
or OR2 (N25, N6, N24);
or OR4 (N26, N17, N17, N18, N19);
or OR2 (N27, N5, N3);
or OR3 (N28, N23, N16, N26);
buf BUF1 (N29, N15);
and AND3 (N30, N29, N2, N12);
not NOT1 (N31, N4);
or OR4 (N32, N22, N25, N13, N18);
nor NOR2 (N33, N11, N4);
or OR4 (N34, N31, N14, N20, N31);
buf BUF1 (N35, N8);
not NOT1 (N36, N15);
xor XOR2 (N37, N19, N25);
nand NAND2 (N38, N32, N20);
buf BUF1 (N39, N21);
xor XOR2 (N40, N34, N23);
not NOT1 (N41, N35);
or OR4 (N42, N40, N25, N40, N13);
and AND4 (N43, N30, N8, N1, N41);
nand NAND4 (N44, N19, N8, N42, N12);
buf BUF1 (N45, N5);
xor XOR2 (N46, N39, N36);
xor XOR2 (N47, N39, N7);
buf BUF1 (N48, N27);
nand NAND3 (N49, N28, N22, N5);
nand NAND3 (N50, N47, N15, N20);
and AND4 (N51, N33, N13, N2, N11);
xor XOR2 (N52, N45, N11);
and AND2 (N53, N52, N27);
xor XOR2 (N54, N37, N23);
or OR2 (N55, N38, N2);
buf BUF1 (N56, N49);
nand NAND4 (N57, N48, N31, N22, N20);
buf BUF1 (N58, N43);
xor XOR2 (N59, N56, N51);
not NOT1 (N60, N2);
xor XOR2 (N61, N53, N2);
not NOT1 (N62, N54);
nor NOR2 (N63, N46, N61);
and AND4 (N64, N18, N46, N13, N6);
and AND3 (N65, N60, N9, N46);
or OR4 (N66, N55, N9, N44, N8);
not NOT1 (N67, N3);
and AND3 (N68, N59, N4, N9);
buf BUF1 (N69, N64);
or OR4 (N70, N66, N34, N43, N23);
buf BUF1 (N71, N67);
buf BUF1 (N72, N50);
nor NOR2 (N73, N72, N27);
nand NAND4 (N74, N73, N61, N67, N6);
nor NOR4 (N75, N71, N46, N21, N11);
nor NOR3 (N76, N57, N12, N23);
nand NAND4 (N77, N65, N40, N35, N57);
nand NAND4 (N78, N70, N12, N34, N42);
and AND2 (N79, N77, N55);
xor XOR2 (N80, N79, N17);
not NOT1 (N81, N76);
xor XOR2 (N82, N75, N19);
nand NAND2 (N83, N69, N45);
and AND4 (N84, N68, N48, N64, N27);
and AND4 (N85, N62, N61, N74, N39);
or OR3 (N86, N81, N65, N25);
nor NOR4 (N87, N4, N73, N6, N60);
buf BUF1 (N88, N82);
nand NAND4 (N89, N85, N19, N54, N63);
nor NOR4 (N90, N1, N28, N7, N79);
nor NOR3 (N91, N83, N20, N70);
buf BUF1 (N92, N88);
nand NAND2 (N93, N90, N24);
buf BUF1 (N94, N78);
nor NOR3 (N95, N86, N69, N44);
not NOT1 (N96, N80);
buf BUF1 (N97, N87);
nand NAND3 (N98, N91, N54, N56);
not NOT1 (N99, N84);
not NOT1 (N100, N58);
or OR4 (N101, N99, N96, N58, N42);
not NOT1 (N102, N86);
nor NOR3 (N103, N92, N21, N7);
or OR4 (N104, N97, N77, N81, N34);
nor NOR4 (N105, N98, N38, N31, N98);
nor NOR3 (N106, N104, N72, N18);
xor XOR2 (N107, N105, N64);
nor NOR3 (N108, N103, N19, N86);
buf BUF1 (N109, N102);
not NOT1 (N110, N108);
and AND4 (N111, N89, N17, N41, N20);
and AND4 (N112, N110, N75, N30, N93);
nor NOR3 (N113, N97, N92, N34);
and AND3 (N114, N101, N60, N34);
buf BUF1 (N115, N114);
not NOT1 (N116, N112);
xor XOR2 (N117, N100, N94);
xor XOR2 (N118, N24, N4);
nor NOR4 (N119, N111, N69, N30, N55);
nor NOR3 (N120, N109, N116, N41);
and AND2 (N121, N117, N9);
and AND2 (N122, N38, N74);
and AND3 (N123, N119, N98, N89);
nand NAND2 (N124, N106, N50);
buf BUF1 (N125, N122);
nor NOR4 (N126, N120, N95, N80, N80);
or OR3 (N127, N1, N38, N63);
xor XOR2 (N128, N118, N7);
buf BUF1 (N129, N123);
nand NAND2 (N130, N129, N18);
not NOT1 (N131, N126);
and AND4 (N132, N127, N92, N69, N66);
not NOT1 (N133, N132);
nor NOR4 (N134, N107, N32, N89, N74);
buf BUF1 (N135, N134);
and AND4 (N136, N135, N44, N113, N107);
not NOT1 (N137, N11);
buf BUF1 (N138, N131);
xor XOR2 (N139, N136, N33);
xor XOR2 (N140, N130, N19);
or OR2 (N141, N138, N96);
not NOT1 (N142, N121);
xor XOR2 (N143, N142, N83);
and AND4 (N144, N128, N66, N56, N89);
and AND3 (N145, N124, N94, N103);
nand NAND3 (N146, N115, N38, N44);
xor XOR2 (N147, N145, N109);
buf BUF1 (N148, N146);
nand NAND4 (N149, N143, N87, N53, N130);
or OR3 (N150, N133, N15, N134);
buf BUF1 (N151, N141);
xor XOR2 (N152, N144, N42);
nand NAND3 (N153, N147, N117, N42);
or OR2 (N154, N148, N105);
xor XOR2 (N155, N153, N60);
not NOT1 (N156, N154);
and AND4 (N157, N137, N81, N138, N93);
not NOT1 (N158, N150);
nand NAND2 (N159, N158, N112);
buf BUF1 (N160, N152);
nor NOR2 (N161, N151, N51);
nor NOR2 (N162, N125, N101);
or OR3 (N163, N139, N142, N55);
nand NAND2 (N164, N160, N122);
and AND2 (N165, N155, N3);
or OR2 (N166, N165, N108);
buf BUF1 (N167, N159);
buf BUF1 (N168, N140);
buf BUF1 (N169, N149);
nor NOR4 (N170, N169, N113, N161, N11);
and AND4 (N171, N54, N161, N100, N20);
xor XOR2 (N172, N162, N83);
nor NOR2 (N173, N170, N60);
buf BUF1 (N174, N156);
or OR4 (N175, N157, N58, N18, N47);
or OR4 (N176, N175, N138, N12, N102);
nor NOR3 (N177, N163, N107, N81);
nand NAND2 (N178, N164, N66);
and AND2 (N179, N178, N113);
xor XOR2 (N180, N167, N10);
not NOT1 (N181, N179);
xor XOR2 (N182, N180, N56);
not NOT1 (N183, N174);
and AND4 (N184, N181, N35, N62, N177);
xor XOR2 (N185, N159, N115);
buf BUF1 (N186, N172);
or OR4 (N187, N182, N73, N72, N150);
buf BUF1 (N188, N173);
not NOT1 (N189, N171);
or OR3 (N190, N188, N61, N34);
and AND3 (N191, N166, N140, N29);
nor NOR2 (N192, N189, N159);
buf BUF1 (N193, N176);
buf BUF1 (N194, N191);
and AND2 (N195, N168, N174);
nor NOR3 (N196, N194, N186, N79);
or OR4 (N197, N5, N18, N79, N1);
xor XOR2 (N198, N183, N190);
nand NAND4 (N199, N41, N37, N174, N67);
or OR3 (N200, N195, N194, N43);
nand NAND3 (N201, N185, N199, N39);
nand NAND3 (N202, N24, N42, N107);
xor XOR2 (N203, N202, N23);
not NOT1 (N204, N198);
and AND3 (N205, N193, N79, N201);
buf BUF1 (N206, N91);
nand NAND2 (N207, N196, N18);
nor NOR4 (N208, N200, N87, N41, N206);
nand NAND2 (N209, N75, N6);
xor XOR2 (N210, N207, N176);
not NOT1 (N211, N204);
xor XOR2 (N212, N209, N145);
not NOT1 (N213, N210);
and AND2 (N214, N213, N135);
nand NAND3 (N215, N192, N169, N152);
xor XOR2 (N216, N197, N24);
or OR4 (N217, N215, N25, N111, N47);
not NOT1 (N218, N203);
not NOT1 (N219, N217);
not NOT1 (N220, N208);
not NOT1 (N221, N220);
or OR4 (N222, N218, N88, N97, N63);
buf BUF1 (N223, N184);
nor NOR3 (N224, N187, N189, N50);
xor XOR2 (N225, N219, N130);
nor NOR4 (N226, N211, N78, N81, N140);
nand NAND4 (N227, N224, N74, N48, N178);
not NOT1 (N228, N214);
not NOT1 (N229, N225);
not NOT1 (N230, N212);
or OR3 (N231, N223, N39, N105);
not NOT1 (N232, N227);
or OR4 (N233, N228, N183, N31, N164);
nand NAND4 (N234, N216, N178, N187, N21);
buf BUF1 (N235, N205);
nor NOR3 (N236, N235, N110, N214);
not NOT1 (N237, N234);
or OR2 (N238, N230, N75);
nor NOR2 (N239, N237, N165);
or OR3 (N240, N239, N110, N43);
and AND3 (N241, N221, N59, N210);
buf BUF1 (N242, N233);
xor XOR2 (N243, N240, N10);
nand NAND2 (N244, N232, N24);
buf BUF1 (N245, N243);
not NOT1 (N246, N244);
nand NAND2 (N247, N236, N169);
nand NAND4 (N248, N229, N219, N18, N247);
buf BUF1 (N249, N124);
or OR2 (N250, N248, N174);
xor XOR2 (N251, N238, N132);
and AND3 (N252, N249, N36, N81);
nor NOR4 (N253, N250, N97, N197, N245);
and AND3 (N254, N217, N212, N52);
not NOT1 (N255, N231);
xor XOR2 (N256, N252, N63);
buf BUF1 (N257, N222);
and AND3 (N258, N257, N75, N218);
nand NAND3 (N259, N253, N50, N120);
buf BUF1 (N260, N241);
not NOT1 (N261, N255);
and AND3 (N262, N226, N172, N31);
and AND3 (N263, N256, N179, N85);
or OR2 (N264, N246, N194);
xor XOR2 (N265, N261, N90);
or OR2 (N266, N265, N185);
not NOT1 (N267, N266);
not NOT1 (N268, N251);
and AND2 (N269, N242, N98);
nand NAND4 (N270, N254, N64, N86, N173);
xor XOR2 (N271, N263, N194);
nand NAND4 (N272, N267, N182, N97, N270);
not NOT1 (N273, N93);
not NOT1 (N274, N260);
and AND4 (N275, N274, N13, N105, N101);
not NOT1 (N276, N268);
xor XOR2 (N277, N276, N85);
and AND4 (N278, N273, N106, N38, N189);
not NOT1 (N279, N259);
xor XOR2 (N280, N269, N85);
not NOT1 (N281, N277);
xor XOR2 (N282, N264, N239);
nor NOR2 (N283, N272, N67);
not NOT1 (N284, N281);
xor XOR2 (N285, N279, N8);
not NOT1 (N286, N285);
xor XOR2 (N287, N278, N207);
buf BUF1 (N288, N258);
buf BUF1 (N289, N283);
or OR3 (N290, N282, N162, N253);
and AND4 (N291, N288, N283, N264, N276);
and AND2 (N292, N291, N178);
nor NOR4 (N293, N290, N14, N290, N132);
buf BUF1 (N294, N286);
buf BUF1 (N295, N280);
nor NOR4 (N296, N293, N159, N221, N8);
nand NAND2 (N297, N294, N45);
not NOT1 (N298, N289);
nand NAND2 (N299, N298, N134);
and AND2 (N300, N296, N241);
nand NAND2 (N301, N275, N300);
xor XOR2 (N302, N177, N60);
nand NAND2 (N303, N299, N108);
xor XOR2 (N304, N302, N249);
or OR2 (N305, N262, N253);
xor XOR2 (N306, N301, N184);
not NOT1 (N307, N271);
nor NOR3 (N308, N306, N51, N238);
or OR3 (N309, N303, N73, N174);
nand NAND3 (N310, N284, N178, N55);
not NOT1 (N311, N295);
nor NOR2 (N312, N308, N7);
nand NAND2 (N313, N309, N239);
xor XOR2 (N314, N313, N273);
nor NOR3 (N315, N310, N104, N79);
nand NAND3 (N316, N304, N268, N193);
and AND2 (N317, N316, N95);
buf BUF1 (N318, N315);
not NOT1 (N319, N305);
buf BUF1 (N320, N287);
not NOT1 (N321, N311);
nand NAND4 (N322, N312, N55, N167, N164);
nor NOR2 (N323, N297, N32);
and AND2 (N324, N322, N76);
xor XOR2 (N325, N324, N52);
or OR4 (N326, N317, N200, N302, N13);
nor NOR3 (N327, N323, N251, N310);
nor NOR3 (N328, N327, N123, N218);
nand NAND2 (N329, N319, N144);
and AND4 (N330, N325, N309, N11, N68);
not NOT1 (N331, N329);
nand NAND2 (N332, N326, N214);
xor XOR2 (N333, N331, N131);
nand NAND2 (N334, N330, N293);
and AND3 (N335, N314, N24, N197);
and AND4 (N336, N328, N256, N154, N83);
buf BUF1 (N337, N318);
nand NAND3 (N338, N321, N216, N163);
nand NAND2 (N339, N307, N70);
nor NOR2 (N340, N334, N131);
xor XOR2 (N341, N333, N204);
nand NAND2 (N342, N292, N282);
nand NAND3 (N343, N342, N258, N118);
buf BUF1 (N344, N337);
or OR4 (N345, N341, N3, N1, N198);
nand NAND2 (N346, N340, N165);
nor NOR3 (N347, N344, N274, N164);
not NOT1 (N348, N346);
not NOT1 (N349, N338);
nand NAND3 (N350, N347, N164, N96);
nand NAND3 (N351, N343, N94, N120);
and AND2 (N352, N345, N91);
nand NAND3 (N353, N335, N37, N159);
xor XOR2 (N354, N352, N175);
not NOT1 (N355, N332);
or OR2 (N356, N348, N270);
and AND3 (N357, N320, N245, N95);
not NOT1 (N358, N355);
nor NOR3 (N359, N339, N53, N88);
nor NOR4 (N360, N354, N292, N266, N271);
xor XOR2 (N361, N357, N276);
nor NOR3 (N362, N336, N119, N275);
and AND3 (N363, N361, N46, N302);
or OR3 (N364, N353, N122, N238);
nand NAND3 (N365, N362, N39, N73);
nand NAND4 (N366, N360, N349, N316, N24);
buf BUF1 (N367, N289);
xor XOR2 (N368, N365, N133);
or OR4 (N369, N359, N320, N130, N131);
xor XOR2 (N370, N351, N198);
or OR2 (N371, N358, N187);
nand NAND2 (N372, N350, N207);
xor XOR2 (N373, N368, N292);
or OR4 (N374, N373, N150, N343, N262);
nor NOR4 (N375, N364, N46, N119, N5);
and AND3 (N376, N372, N164, N251);
or OR2 (N377, N371, N45);
xor XOR2 (N378, N376, N337);
nand NAND3 (N379, N363, N8, N70);
or OR3 (N380, N356, N163, N291);
xor XOR2 (N381, N375, N207);
nand NAND3 (N382, N369, N6, N274);
buf BUF1 (N383, N378);
not NOT1 (N384, N374);
not NOT1 (N385, N366);
xor XOR2 (N386, N379, N59);
nor NOR3 (N387, N367, N339, N340);
nor NOR2 (N388, N381, N203);
buf BUF1 (N389, N377);
and AND4 (N390, N383, N87, N228, N63);
nor NOR4 (N391, N387, N307, N70, N28);
not NOT1 (N392, N380);
and AND2 (N393, N386, N279);
nor NOR4 (N394, N382, N52, N312, N320);
buf BUF1 (N395, N385);
xor XOR2 (N396, N394, N67);
or OR3 (N397, N388, N97, N369);
nor NOR4 (N398, N390, N96, N93, N44);
and AND3 (N399, N392, N332, N269);
not NOT1 (N400, N384);
or OR4 (N401, N398, N112, N198, N269);
or OR2 (N402, N400, N280);
nor NOR2 (N403, N397, N170);
xor XOR2 (N404, N389, N88);
and AND3 (N405, N396, N311, N382);
not NOT1 (N406, N399);
nor NOR4 (N407, N395, N246, N97, N118);
not NOT1 (N408, N403);
or OR2 (N409, N370, N213);
nor NOR2 (N410, N405, N241);
buf BUF1 (N411, N402);
nor NOR3 (N412, N393, N224, N135);
or OR2 (N413, N406, N65);
buf BUF1 (N414, N409);
and AND3 (N415, N408, N394, N23);
or OR2 (N416, N412, N113);
buf BUF1 (N417, N391);
buf BUF1 (N418, N407);
or OR2 (N419, N410, N239);
nor NOR4 (N420, N415, N38, N223, N412);
xor XOR2 (N421, N404, N71);
and AND4 (N422, N401, N170, N414, N168);
or OR2 (N423, N374, N197);
nand NAND3 (N424, N423, N78, N120);
buf BUF1 (N425, N418);
nand NAND4 (N426, N422, N275, N36, N178);
nand NAND2 (N427, N413, N262);
not NOT1 (N428, N421);
or OR2 (N429, N427, N410);
or OR3 (N430, N424, N138, N242);
or OR4 (N431, N417, N37, N77, N393);
xor XOR2 (N432, N420, N365);
nand NAND3 (N433, N431, N3, N416);
xor XOR2 (N434, N100, N269);
and AND2 (N435, N411, N7);
xor XOR2 (N436, N429, N299);
and AND2 (N437, N432, N91);
nor NOR2 (N438, N434, N2);
nand NAND3 (N439, N419, N362, N101);
buf BUF1 (N440, N436);
nand NAND2 (N441, N426, N151);
nor NOR2 (N442, N439, N224);
nor NOR4 (N443, N440, N301, N433, N315);
nor NOR3 (N444, N141, N352, N100);
or OR4 (N445, N425, N383, N268, N410);
xor XOR2 (N446, N442, N20);
xor XOR2 (N447, N445, N98);
not NOT1 (N448, N430);
or OR3 (N449, N447, N196, N6);
nand NAND2 (N450, N428, N338);
nand NAND4 (N451, N435, N422, N60, N126);
nand NAND2 (N452, N444, N44);
nand NAND2 (N453, N449, N426);
not NOT1 (N454, N451);
not NOT1 (N455, N450);
xor XOR2 (N456, N441, N160);
nor NOR4 (N457, N453, N418, N246, N361);
buf BUF1 (N458, N457);
or OR2 (N459, N448, N44);
nor NOR2 (N460, N446, N9);
nand NAND4 (N461, N438, N163, N367, N412);
nand NAND4 (N462, N452, N382, N375, N2);
and AND3 (N463, N462, N64, N364);
or OR4 (N464, N443, N259, N204, N143);
and AND3 (N465, N454, N80, N197);
not NOT1 (N466, N459);
nor NOR3 (N467, N437, N105, N457);
or OR2 (N468, N464, N124);
nor NOR3 (N469, N465, N24, N454);
nand NAND2 (N470, N467, N384);
and AND4 (N471, N458, N259, N141, N355);
or OR2 (N472, N469, N169);
or OR3 (N473, N456, N158, N346);
and AND4 (N474, N460, N110, N375, N249);
or OR3 (N475, N470, N428, N398);
or OR2 (N476, N455, N35);
not NOT1 (N477, N463);
and AND4 (N478, N473, N49, N347, N463);
or OR3 (N479, N468, N192, N465);
nand NAND4 (N480, N471, N284, N470, N398);
and AND2 (N481, N478, N461);
not NOT1 (N482, N462);
and AND3 (N483, N472, N480, N21);
not NOT1 (N484, N477);
and AND4 (N485, N157, N306, N421, N284);
or OR4 (N486, N483, N73, N225, N387);
or OR3 (N487, N476, N243, N167);
buf BUF1 (N488, N474);
nand NAND4 (N489, N485, N433, N316, N47);
or OR2 (N490, N489, N270);
buf BUF1 (N491, N481);
buf BUF1 (N492, N487);
or OR4 (N493, N492, N361, N18, N348);
or OR3 (N494, N466, N426, N304);
xor XOR2 (N495, N484, N299);
xor XOR2 (N496, N479, N33);
xor XOR2 (N497, N494, N251);
or OR4 (N498, N490, N190, N325, N223);
nor NOR2 (N499, N486, N386);
xor XOR2 (N500, N496, N472);
xor XOR2 (N501, N500, N179);
buf BUF1 (N502, N497);
xor XOR2 (N503, N498, N117);
xor XOR2 (N504, N493, N410);
or OR3 (N505, N502, N71, N383);
xor XOR2 (N506, N503, N61);
and AND4 (N507, N505, N21, N23, N462);
not NOT1 (N508, N501);
xor XOR2 (N509, N507, N96);
not NOT1 (N510, N504);
nand NAND2 (N511, N488, N321);
and AND3 (N512, N475, N394, N51);
buf BUF1 (N513, N495);
or OR2 (N514, N509, N394);
nand NAND3 (N515, N512, N294, N118);
nand NAND2 (N516, N508, N422);
and AND3 (N517, N499, N379, N380);
nand NAND4 (N518, N491, N74, N386, N250);
buf BUF1 (N519, N506);
or OR3 (N520, N515, N214, N484);
xor XOR2 (N521, N517, N194);
and AND3 (N522, N513, N375, N18);
and AND3 (N523, N482, N306, N313);
and AND3 (N524, N514, N16, N102);
not NOT1 (N525, N522);
and AND3 (N526, N511, N271, N514);
or OR4 (N527, N524, N276, N143, N179);
buf BUF1 (N528, N525);
or OR2 (N529, N528, N96);
or OR3 (N530, N529, N37, N413);
xor XOR2 (N531, N518, N168);
nand NAND3 (N532, N526, N152, N172);
and AND4 (N533, N520, N507, N369, N299);
not NOT1 (N534, N533);
xor XOR2 (N535, N516, N269);
nor NOR4 (N536, N531, N176, N445, N174);
not NOT1 (N537, N523);
not NOT1 (N538, N534);
or OR4 (N539, N536, N281, N341, N495);
buf BUF1 (N540, N538);
and AND4 (N541, N527, N216, N128, N416);
not NOT1 (N542, N519);
not NOT1 (N543, N541);
or OR3 (N544, N537, N105, N55);
or OR2 (N545, N544, N448);
xor XOR2 (N546, N545, N15);
buf BUF1 (N547, N535);
or OR3 (N548, N542, N415, N331);
and AND2 (N549, N540, N35);
xor XOR2 (N550, N543, N14);
or OR4 (N551, N521, N546, N480, N489);
and AND2 (N552, N159, N78);
or OR3 (N553, N547, N57, N139);
nand NAND2 (N554, N551, N530);
not NOT1 (N555, N413);
or OR2 (N556, N552, N383);
nand NAND4 (N557, N556, N543, N365, N163);
nand NAND2 (N558, N550, N334);
nor NOR2 (N559, N553, N304);
or OR2 (N560, N548, N228);
or OR4 (N561, N555, N464, N526, N151);
nand NAND2 (N562, N557, N470);
xor XOR2 (N563, N549, N178);
nand NAND2 (N564, N561, N407);
or OR2 (N565, N564, N499);
xor XOR2 (N566, N558, N423);
nand NAND4 (N567, N563, N128, N328, N470);
not NOT1 (N568, N510);
buf BUF1 (N569, N554);
or OR4 (N570, N565, N248, N416, N179);
not NOT1 (N571, N560);
buf BUF1 (N572, N570);
not NOT1 (N573, N532);
and AND4 (N574, N559, N225, N86, N177);
not NOT1 (N575, N562);
and AND3 (N576, N567, N89, N112);
nor NOR4 (N577, N566, N15, N507, N324);
not NOT1 (N578, N575);
and AND3 (N579, N572, N466, N180);
nand NAND3 (N580, N539, N244, N355);
nand NAND2 (N581, N576, N365);
and AND2 (N582, N577, N111);
xor XOR2 (N583, N568, N90);
nand NAND2 (N584, N578, N419);
buf BUF1 (N585, N579);
and AND3 (N586, N569, N558, N535);
or OR3 (N587, N585, N289, N213);
not NOT1 (N588, N580);
or OR4 (N589, N571, N308, N499, N438);
not NOT1 (N590, N574);
or OR2 (N591, N587, N460);
not NOT1 (N592, N573);
xor XOR2 (N593, N584, N263);
nor NOR2 (N594, N590, N293);
xor XOR2 (N595, N592, N158);
nor NOR4 (N596, N582, N248, N224, N82);
and AND3 (N597, N591, N5, N526);
not NOT1 (N598, N583);
buf BUF1 (N599, N593);
xor XOR2 (N600, N596, N250);
and AND2 (N601, N598, N451);
and AND2 (N602, N594, N160);
nor NOR4 (N603, N588, N455, N392, N455);
nor NOR3 (N604, N589, N560, N533);
and AND3 (N605, N586, N240, N69);
or OR3 (N606, N597, N353, N223);
nor NOR2 (N607, N600, N388);
nand NAND4 (N608, N605, N292, N362, N577);
xor XOR2 (N609, N601, N237);
and AND4 (N610, N609, N160, N526, N245);
or OR2 (N611, N606, N267);
or OR4 (N612, N610, N109, N197, N55);
and AND2 (N613, N581, N424);
xor XOR2 (N614, N603, N317);
nand NAND3 (N615, N611, N305, N144);
xor XOR2 (N616, N615, N13);
or OR4 (N617, N604, N336, N9, N129);
nor NOR4 (N618, N612, N282, N190, N423);
and AND2 (N619, N607, N532);
and AND3 (N620, N608, N584, N199);
buf BUF1 (N621, N616);
buf BUF1 (N622, N619);
nand NAND2 (N623, N622, N42);
and AND4 (N624, N614, N322, N552, N90);
buf BUF1 (N625, N602);
and AND3 (N626, N595, N463, N32);
xor XOR2 (N627, N623, N106);
or OR2 (N628, N627, N473);
not NOT1 (N629, N624);
xor XOR2 (N630, N620, N612);
xor XOR2 (N631, N625, N248);
and AND2 (N632, N617, N586);
xor XOR2 (N633, N629, N531);
or OR2 (N634, N633, N513);
buf BUF1 (N635, N628);
nor NOR4 (N636, N634, N142, N565, N59);
xor XOR2 (N637, N630, N24);
nor NOR4 (N638, N613, N11, N384, N413);
not NOT1 (N639, N636);
and AND2 (N640, N637, N425);
or OR2 (N641, N639, N179);
not NOT1 (N642, N631);
nand NAND2 (N643, N621, N638);
xor XOR2 (N644, N271, N228);
and AND4 (N645, N644, N46, N243, N283);
nor NOR2 (N646, N599, N479);
and AND3 (N647, N641, N1, N81);
nand NAND3 (N648, N626, N345, N166);
nand NAND2 (N649, N632, N434);
not NOT1 (N650, N640);
nor NOR3 (N651, N643, N355, N190);
nor NOR2 (N652, N651, N588);
nand NAND2 (N653, N652, N513);
nand NAND2 (N654, N653, N220);
buf BUF1 (N655, N645);
or OR3 (N656, N649, N623, N401);
nand NAND4 (N657, N618, N378, N271, N557);
buf BUF1 (N658, N648);
buf BUF1 (N659, N642);
nor NOR2 (N660, N646, N98);
buf BUF1 (N661, N656);
or OR2 (N662, N635, N526);
or OR4 (N663, N661, N385, N473, N205);
or OR2 (N664, N647, N546);
and AND2 (N665, N658, N487);
or OR2 (N666, N659, N398);
nand NAND3 (N667, N664, N477, N493);
not NOT1 (N668, N650);
nand NAND4 (N669, N667, N307, N102, N230);
or OR2 (N670, N657, N493);
buf BUF1 (N671, N668);
and AND2 (N672, N662, N241);
not NOT1 (N673, N671);
xor XOR2 (N674, N665, N514);
nor NOR3 (N675, N663, N506, N501);
buf BUF1 (N676, N674);
nor NOR3 (N677, N655, N199, N48);
or OR4 (N678, N675, N306, N423, N186);
buf BUF1 (N679, N660);
or OR4 (N680, N670, N459, N3, N518);
or OR3 (N681, N672, N660, N667);
and AND4 (N682, N679, N172, N99, N485);
or OR4 (N683, N681, N335, N514, N144);
xor XOR2 (N684, N683, N240);
xor XOR2 (N685, N676, N600);
and AND4 (N686, N684, N389, N424, N489);
nand NAND2 (N687, N673, N501);
and AND2 (N688, N666, N524);
or OR2 (N689, N686, N172);
or OR2 (N690, N654, N631);
or OR2 (N691, N687, N597);
xor XOR2 (N692, N680, N122);
nand NAND2 (N693, N677, N453);
buf BUF1 (N694, N685);
nor NOR4 (N695, N692, N642, N39, N49);
nor NOR3 (N696, N695, N235, N75);
nor NOR3 (N697, N682, N218, N166);
nand NAND3 (N698, N688, N409, N39);
buf BUF1 (N699, N678);
or OR2 (N700, N697, N158);
or OR2 (N701, N698, N100);
not NOT1 (N702, N694);
or OR3 (N703, N701, N251, N289);
nor NOR4 (N704, N690, N268, N162, N320);
buf BUF1 (N705, N689);
not NOT1 (N706, N699);
buf BUF1 (N707, N706);
buf BUF1 (N708, N704);
nand NAND4 (N709, N702, N603, N612, N638);
nor NOR2 (N710, N700, N59);
nor NOR3 (N711, N707, N48, N651);
not NOT1 (N712, N708);
or OR2 (N713, N705, N453);
buf BUF1 (N714, N691);
nand NAND4 (N715, N696, N97, N17, N650);
xor XOR2 (N716, N713, N46);
not NOT1 (N717, N715);
buf BUF1 (N718, N710);
nor NOR2 (N719, N716, N65);
nor NOR3 (N720, N669, N279, N645);
nand NAND2 (N721, N711, N395);
xor XOR2 (N722, N717, N613);
not NOT1 (N723, N712);
and AND2 (N724, N709, N250);
nand NAND2 (N725, N720, N218);
xor XOR2 (N726, N714, N367);
and AND4 (N727, N722, N4, N158, N281);
or OR3 (N728, N726, N694, N631);
not NOT1 (N729, N725);
or OR2 (N730, N693, N628);
and AND2 (N731, N719, N173);
buf BUF1 (N732, N731);
or OR4 (N733, N718, N505, N445, N600);
nor NOR2 (N734, N703, N572);
nand NAND3 (N735, N724, N117, N123);
xor XOR2 (N736, N729, N329);
not NOT1 (N737, N736);
and AND2 (N738, N727, N376);
and AND3 (N739, N738, N507, N533);
nor NOR4 (N740, N723, N166, N401, N430);
nand NAND3 (N741, N737, N351, N485);
and AND4 (N742, N741, N278, N572, N126);
not NOT1 (N743, N733);
xor XOR2 (N744, N740, N56);
and AND4 (N745, N734, N660, N297, N70);
not NOT1 (N746, N728);
xor XOR2 (N747, N742, N234);
nor NOR3 (N748, N730, N321, N212);
nor NOR3 (N749, N739, N99, N363);
buf BUF1 (N750, N749);
nand NAND2 (N751, N746, N508);
or OR4 (N752, N735, N678, N397, N26);
xor XOR2 (N753, N743, N100);
xor XOR2 (N754, N751, N489);
nor NOR3 (N755, N745, N442, N203);
nor NOR2 (N756, N753, N435);
and AND4 (N757, N721, N203, N291, N464);
xor XOR2 (N758, N744, N665);
buf BUF1 (N759, N750);
and AND3 (N760, N732, N452, N33);
nor NOR3 (N761, N754, N12, N456);
not NOT1 (N762, N757);
buf BUF1 (N763, N752);
nor NOR4 (N764, N747, N410, N581, N120);
and AND3 (N765, N758, N536, N70);
xor XOR2 (N766, N748, N349);
buf BUF1 (N767, N764);
xor XOR2 (N768, N759, N245);
and AND4 (N769, N755, N336, N150, N331);
buf BUF1 (N770, N765);
and AND3 (N771, N762, N321, N518);
or OR2 (N772, N769, N419);
and AND4 (N773, N767, N11, N246, N126);
nand NAND2 (N774, N770, N452);
nor NOR4 (N775, N766, N574, N350, N362);
nor NOR4 (N776, N773, N589, N737, N424);
not NOT1 (N777, N763);
nand NAND2 (N778, N768, N474);
or OR4 (N779, N771, N655, N610, N334);
not NOT1 (N780, N761);
nor NOR3 (N781, N772, N192, N675);
or OR2 (N782, N780, N239);
and AND2 (N783, N775, N319);
nand NAND4 (N784, N779, N741, N144, N140);
xor XOR2 (N785, N783, N210);
nor NOR2 (N786, N776, N782);
nor NOR4 (N787, N546, N455, N759, N60);
and AND2 (N788, N785, N6);
and AND3 (N789, N784, N166, N735);
nand NAND3 (N790, N778, N736, N184);
xor XOR2 (N791, N788, N589);
and AND2 (N792, N787, N307);
nor NOR2 (N793, N789, N48);
nor NOR2 (N794, N792, N478);
not NOT1 (N795, N791);
not NOT1 (N796, N794);
and AND2 (N797, N781, N207);
nor NOR4 (N798, N760, N577, N178, N762);
not NOT1 (N799, N777);
buf BUF1 (N800, N786);
nand NAND4 (N801, N790, N245, N387, N732);
xor XOR2 (N802, N800, N712);
buf BUF1 (N803, N795);
or OR4 (N804, N803, N726, N54, N9);
xor XOR2 (N805, N804, N372);
not NOT1 (N806, N802);
nand NAND4 (N807, N797, N259, N705, N248);
nor NOR3 (N808, N806, N502, N202);
or OR2 (N809, N796, N764);
xor XOR2 (N810, N799, N618);
buf BUF1 (N811, N774);
and AND3 (N812, N801, N600, N285);
or OR3 (N813, N809, N778, N746);
xor XOR2 (N814, N810, N341);
buf BUF1 (N815, N814);
not NOT1 (N816, N812);
nand NAND3 (N817, N813, N754, N538);
xor XOR2 (N818, N807, N416);
and AND2 (N819, N818, N251);
xor XOR2 (N820, N816, N197);
nor NOR3 (N821, N808, N400, N7);
not NOT1 (N822, N819);
nand NAND3 (N823, N822, N337, N150);
xor XOR2 (N824, N815, N352);
and AND4 (N825, N805, N422, N9, N237);
not NOT1 (N826, N821);
nor NOR2 (N827, N824, N246);
and AND3 (N828, N820, N396, N519);
or OR2 (N829, N811, N159);
and AND2 (N830, N825, N739);
or OR2 (N831, N826, N200);
and AND4 (N832, N817, N10, N115, N792);
xor XOR2 (N833, N827, N15);
or OR4 (N834, N830, N235, N766, N458);
and AND3 (N835, N823, N66, N43);
xor XOR2 (N836, N798, N517);
buf BUF1 (N837, N836);
nor NOR3 (N838, N835, N251, N468);
nor NOR2 (N839, N756, N422);
not NOT1 (N840, N833);
buf BUF1 (N841, N839);
not NOT1 (N842, N828);
and AND2 (N843, N841, N246);
or OR2 (N844, N838, N687);
buf BUF1 (N845, N843);
buf BUF1 (N846, N793);
xor XOR2 (N847, N837, N317);
buf BUF1 (N848, N846);
buf BUF1 (N849, N831);
not NOT1 (N850, N849);
not NOT1 (N851, N850);
not NOT1 (N852, N845);
not NOT1 (N853, N844);
or OR4 (N854, N853, N482, N590, N418);
not NOT1 (N855, N832);
xor XOR2 (N856, N847, N68);
nor NOR3 (N857, N851, N797, N854);
nor NOR4 (N858, N378, N739, N793, N358);
buf BUF1 (N859, N829);
nor NOR4 (N860, N848, N81, N414, N244);
and AND4 (N861, N857, N120, N854, N624);
nor NOR2 (N862, N852, N634);
xor XOR2 (N863, N860, N303);
and AND3 (N864, N834, N495, N151);
nand NAND2 (N865, N842, N739);
nor NOR2 (N866, N864, N152);
nand NAND3 (N867, N862, N6, N707);
xor XOR2 (N868, N866, N660);
and AND2 (N869, N865, N767);
not NOT1 (N870, N858);
not NOT1 (N871, N870);
and AND2 (N872, N861, N287);
buf BUF1 (N873, N872);
buf BUF1 (N874, N855);
nor NOR2 (N875, N840, N316);
nand NAND2 (N876, N867, N621);
nor NOR4 (N877, N875, N482, N76, N177);
buf BUF1 (N878, N871);
nand NAND4 (N879, N874, N567, N184, N276);
xor XOR2 (N880, N859, N51);
nand NAND4 (N881, N879, N173, N851, N308);
or OR3 (N882, N877, N837, N171);
not NOT1 (N883, N876);
buf BUF1 (N884, N873);
nor NOR4 (N885, N884, N737, N163, N211);
nor NOR4 (N886, N885, N623, N170, N26);
buf BUF1 (N887, N882);
nor NOR4 (N888, N878, N661, N322, N304);
nor NOR3 (N889, N881, N853, N217);
xor XOR2 (N890, N886, N25);
buf BUF1 (N891, N868);
buf BUF1 (N892, N891);
buf BUF1 (N893, N863);
nand NAND3 (N894, N889, N123, N156);
or OR3 (N895, N887, N810, N22);
nor NOR3 (N896, N893, N408, N660);
or OR2 (N897, N894, N627);
and AND2 (N898, N888, N554);
nor NOR4 (N899, N880, N288, N681, N785);
and AND4 (N900, N883, N698, N832, N359);
nor NOR4 (N901, N892, N699, N746, N757);
buf BUF1 (N902, N897);
not NOT1 (N903, N890);
or OR3 (N904, N896, N527, N613);
nor NOR2 (N905, N895, N446);
not NOT1 (N906, N904);
nand NAND2 (N907, N905, N292);
not NOT1 (N908, N906);
not NOT1 (N909, N907);
or OR4 (N910, N898, N389, N732, N186);
nor NOR2 (N911, N856, N466);
nand NAND2 (N912, N911, N593);
or OR4 (N913, N909, N598, N539, N650);
not NOT1 (N914, N869);
not NOT1 (N915, N899);
not NOT1 (N916, N908);
buf BUF1 (N917, N901);
buf BUF1 (N918, N915);
and AND4 (N919, N912, N192, N546, N195);
nand NAND2 (N920, N902, N844);
or OR2 (N921, N919, N740);
nor NOR2 (N922, N910, N188);
xor XOR2 (N923, N914, N599);
nand NAND4 (N924, N916, N246, N882, N117);
nor NOR4 (N925, N922, N579, N297, N667);
nor NOR3 (N926, N923, N603, N459);
not NOT1 (N927, N917);
or OR4 (N928, N913, N366, N117, N876);
nor NOR4 (N929, N924, N756, N866, N734);
not NOT1 (N930, N929);
not NOT1 (N931, N926);
nand NAND3 (N932, N928, N16, N111);
xor XOR2 (N933, N900, N410);
nand NAND4 (N934, N932, N308, N804, N592);
nor NOR2 (N935, N933, N266);
nand NAND4 (N936, N920, N445, N213, N599);
or OR4 (N937, N925, N46, N370, N23);
xor XOR2 (N938, N930, N604);
not NOT1 (N939, N931);
xor XOR2 (N940, N918, N406);
buf BUF1 (N941, N935);
and AND4 (N942, N937, N91, N475, N240);
nor NOR4 (N943, N942, N750, N76, N77);
nor NOR2 (N944, N943, N194);
not NOT1 (N945, N927);
or OR2 (N946, N903, N242);
nand NAND4 (N947, N921, N893, N927, N818);
not NOT1 (N948, N936);
nor NOR4 (N949, N944, N599, N23, N130);
or OR3 (N950, N941, N33, N467);
not NOT1 (N951, N947);
or OR4 (N952, N950, N453, N372, N150);
or OR4 (N953, N940, N120, N507, N224);
not NOT1 (N954, N951);
xor XOR2 (N955, N939, N569);
or OR3 (N956, N952, N333, N69);
nor NOR4 (N957, N938, N840, N699, N893);
and AND4 (N958, N957, N178, N694, N707);
nand NAND4 (N959, N953, N516, N788, N475);
nor NOR3 (N960, N959, N248, N393);
nor NOR3 (N961, N954, N634, N907);
or OR4 (N962, N960, N788, N506, N762);
not NOT1 (N963, N955);
nand NAND2 (N964, N949, N531);
nor NOR3 (N965, N963, N291, N636);
nor NOR3 (N966, N948, N310, N906);
nand NAND2 (N967, N962, N507);
buf BUF1 (N968, N945);
and AND2 (N969, N946, N433);
nand NAND3 (N970, N965, N517, N375);
and AND2 (N971, N964, N87);
xor XOR2 (N972, N961, N490);
nor NOR3 (N973, N970, N811, N899);
nand NAND4 (N974, N934, N590, N527, N692);
not NOT1 (N975, N969);
nor NOR3 (N976, N958, N813, N237);
or OR4 (N977, N975, N291, N87, N66);
nor NOR3 (N978, N956, N753, N928);
not NOT1 (N979, N968);
and AND2 (N980, N974, N553);
and AND3 (N981, N977, N783, N164);
nand NAND2 (N982, N981, N396);
nand NAND4 (N983, N978, N703, N92, N585);
and AND3 (N984, N983, N386, N309);
xor XOR2 (N985, N979, N527);
not NOT1 (N986, N980);
or OR2 (N987, N985, N396);
nor NOR4 (N988, N971, N107, N701, N292);
and AND4 (N989, N966, N32, N59, N91);
nand NAND4 (N990, N988, N449, N39, N299);
buf BUF1 (N991, N973);
nand NAND3 (N992, N976, N407, N989);
and AND2 (N993, N789, N115);
not NOT1 (N994, N986);
not NOT1 (N995, N990);
nand NAND4 (N996, N993, N611, N230, N795);
not NOT1 (N997, N992);
nand NAND3 (N998, N987, N310, N460);
xor XOR2 (N999, N967, N130);
xor XOR2 (N1000, N984, N224);
buf BUF1 (N1001, N996);
xor XOR2 (N1002, N982, N751);
nor NOR4 (N1003, N999, N323, N662, N179);
not NOT1 (N1004, N994);
buf BUF1 (N1005, N1002);
xor XOR2 (N1006, N972, N675);
buf BUF1 (N1007, N998);
xor XOR2 (N1008, N1004, N297);
or OR2 (N1009, N1006, N562);
buf BUF1 (N1010, N1000);
endmodule