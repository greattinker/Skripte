// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20;

output N2014,N2002,N2012,N2017,N2015,N2007,N2016,N2018,N2019,N2020;

not NOT1 (N21, N18);
buf BUF1 (N22, N3);
not NOT1 (N23, N10);
not NOT1 (N24, N15);
nand NAND2 (N25, N3, N20);
and AND2 (N26, N9, N12);
nor NOR2 (N27, N20, N5);
or OR3 (N28, N16, N18, N8);
nor NOR3 (N29, N13, N28, N23);
and AND4 (N30, N11, N11, N6, N26);
nand NAND2 (N31, N28, N27);
or OR3 (N32, N12, N27, N29);
nand NAND3 (N33, N26, N20, N14);
not NOT1 (N34, N8);
not NOT1 (N35, N13);
buf BUF1 (N36, N24);
nor NOR2 (N37, N35, N27);
and AND3 (N38, N32, N16, N18);
or OR4 (N39, N30, N37, N28, N37);
xor XOR2 (N40, N22, N38);
nand NAND4 (N41, N3, N15, N40, N20);
and AND4 (N42, N22, N26, N31, N12);
nand NAND2 (N43, N13, N39);
nor NOR4 (N44, N27, N25, N3, N8);
buf BUF1 (N45, N44);
nor NOR3 (N46, N8, N25, N21);
not NOT1 (N47, N10);
xor XOR2 (N48, N34, N8);
and AND3 (N49, N39, N32, N39);
nor NOR2 (N50, N43, N16);
xor XOR2 (N51, N33, N12);
not NOT1 (N52, N46);
nand NAND3 (N53, N42, N22, N43);
or OR4 (N54, N36, N12, N13, N11);
not NOT1 (N55, N41);
xor XOR2 (N56, N52, N7);
not NOT1 (N57, N53);
and AND3 (N58, N57, N25, N25);
not NOT1 (N59, N48);
buf BUF1 (N60, N54);
xor XOR2 (N61, N51, N32);
not NOT1 (N62, N61);
nand NAND4 (N63, N47, N9, N27, N35);
buf BUF1 (N64, N63);
buf BUF1 (N65, N45);
buf BUF1 (N66, N56);
and AND3 (N67, N58, N5, N13);
nand NAND2 (N68, N60, N30);
nand NAND4 (N69, N66, N32, N18, N21);
nor NOR2 (N70, N59, N49);
buf BUF1 (N71, N63);
or OR3 (N72, N65, N49, N14);
or OR2 (N73, N71, N36);
nor NOR2 (N74, N70, N13);
xor XOR2 (N75, N50, N17);
not NOT1 (N76, N73);
and AND4 (N77, N64, N7, N71, N5);
nor NOR2 (N78, N74, N8);
buf BUF1 (N79, N69);
and AND2 (N80, N75, N34);
or OR3 (N81, N78, N6, N67);
or OR4 (N82, N46, N36, N19, N29);
xor XOR2 (N83, N80, N13);
and AND4 (N84, N62, N42, N47, N52);
nor NOR4 (N85, N68, N18, N34, N52);
and AND3 (N86, N72, N29, N58);
buf BUF1 (N87, N55);
not NOT1 (N88, N79);
or OR4 (N89, N86, N23, N39, N3);
xor XOR2 (N90, N84, N31);
not NOT1 (N91, N77);
and AND2 (N92, N89, N82);
nand NAND2 (N93, N57, N53);
xor XOR2 (N94, N92, N48);
and AND4 (N95, N88, N61, N88, N35);
nand NAND3 (N96, N91, N66, N28);
xor XOR2 (N97, N81, N28);
not NOT1 (N98, N97);
not NOT1 (N99, N96);
xor XOR2 (N100, N87, N33);
buf BUF1 (N101, N85);
nand NAND2 (N102, N99, N63);
or OR3 (N103, N102, N5, N91);
nand NAND4 (N104, N94, N40, N94, N70);
or OR3 (N105, N95, N3, N47);
nor NOR2 (N106, N90, N82);
nor NOR2 (N107, N98, N35);
buf BUF1 (N108, N93);
xor XOR2 (N109, N103, N60);
and AND3 (N110, N83, N56, N36);
xor XOR2 (N111, N107, N7);
nor NOR2 (N112, N108, N88);
nor NOR4 (N113, N101, N16, N47, N84);
nor NOR2 (N114, N106, N58);
not NOT1 (N115, N105);
nor NOR2 (N116, N109, N98);
nand NAND3 (N117, N112, N96, N32);
buf BUF1 (N118, N115);
nand NAND4 (N119, N118, N28, N9, N100);
xor XOR2 (N120, N38, N58);
nand NAND3 (N121, N110, N30, N21);
and AND3 (N122, N117, N89, N12);
and AND3 (N123, N119, N2, N91);
xor XOR2 (N124, N116, N61);
or OR3 (N125, N76, N5, N52);
xor XOR2 (N126, N104, N30);
or OR2 (N127, N124, N86);
xor XOR2 (N128, N123, N37);
nand NAND3 (N129, N127, N56, N48);
xor XOR2 (N130, N113, N61);
and AND4 (N131, N130, N104, N7, N103);
or OR4 (N132, N125, N103, N66, N16);
buf BUF1 (N133, N131);
nor NOR2 (N134, N129, N83);
buf BUF1 (N135, N134);
not NOT1 (N136, N132);
and AND4 (N137, N111, N21, N27, N53);
xor XOR2 (N138, N126, N39);
nand NAND2 (N139, N120, N43);
nand NAND3 (N140, N138, N54, N61);
and AND2 (N141, N114, N91);
nand NAND4 (N142, N135, N68, N123, N129);
and AND3 (N143, N122, N21, N127);
not NOT1 (N144, N140);
or OR3 (N145, N137, N24, N72);
and AND4 (N146, N141, N59, N3, N82);
or OR3 (N147, N146, N135, N95);
and AND4 (N148, N144, N137, N57, N24);
not NOT1 (N149, N148);
nand NAND2 (N150, N133, N6);
and AND2 (N151, N136, N36);
buf BUF1 (N152, N150);
xor XOR2 (N153, N128, N146);
buf BUF1 (N154, N142);
buf BUF1 (N155, N151);
not NOT1 (N156, N143);
and AND3 (N157, N152, N132, N135);
nor NOR3 (N158, N155, N59, N24);
buf BUF1 (N159, N121);
nor NOR4 (N160, N145, N20, N130, N42);
or OR3 (N161, N159, N40, N156);
buf BUF1 (N162, N153);
not NOT1 (N163, N132);
nand NAND4 (N164, N162, N83, N94, N135);
and AND4 (N165, N161, N146, N159, N162);
xor XOR2 (N166, N158, N159);
not NOT1 (N167, N165);
xor XOR2 (N168, N154, N124);
nand NAND3 (N169, N167, N109, N80);
or OR2 (N170, N157, N81);
not NOT1 (N171, N169);
and AND3 (N172, N163, N9, N61);
not NOT1 (N173, N170);
buf BUF1 (N174, N168);
not NOT1 (N175, N172);
nand NAND4 (N176, N174, N65, N106, N53);
and AND2 (N177, N149, N117);
not NOT1 (N178, N173);
and AND2 (N179, N164, N125);
and AND3 (N180, N177, N144, N35);
buf BUF1 (N181, N139);
not NOT1 (N182, N175);
or OR3 (N183, N147, N118, N43);
nor NOR4 (N184, N176, N146, N15, N154);
buf BUF1 (N185, N166);
nor NOR4 (N186, N184, N10, N133, N87);
or OR2 (N187, N180, N80);
not NOT1 (N188, N185);
and AND2 (N189, N179, N92);
not NOT1 (N190, N183);
buf BUF1 (N191, N171);
not NOT1 (N192, N188);
buf BUF1 (N193, N182);
and AND2 (N194, N160, N170);
nor NOR3 (N195, N193, N170, N153);
xor XOR2 (N196, N187, N98);
nand NAND4 (N197, N196, N185, N140, N196);
and AND3 (N198, N186, N79, N10);
xor XOR2 (N199, N198, N73);
not NOT1 (N200, N197);
buf BUF1 (N201, N200);
and AND4 (N202, N189, N194, N154, N145);
xor XOR2 (N203, N172, N75);
and AND2 (N204, N195, N167);
nand NAND4 (N205, N199, N164, N91, N112);
xor XOR2 (N206, N181, N33);
not NOT1 (N207, N191);
nor NOR2 (N208, N201, N91);
nand NAND4 (N209, N202, N131, N52, N155);
not NOT1 (N210, N204);
xor XOR2 (N211, N207, N37);
xor XOR2 (N212, N178, N61);
nand NAND2 (N213, N192, N130);
nor NOR2 (N214, N213, N86);
and AND3 (N215, N209, N138, N131);
nor NOR3 (N216, N214, N178, N80);
not NOT1 (N217, N206);
or OR3 (N218, N217, N108, N167);
and AND2 (N219, N218, N199);
buf BUF1 (N220, N203);
nor NOR3 (N221, N211, N142, N122);
and AND4 (N222, N219, N145, N97, N72);
or OR3 (N223, N222, N81, N106);
nand NAND2 (N224, N212, N94);
nand NAND4 (N225, N210, N176, N119, N67);
and AND4 (N226, N221, N115, N89, N80);
xor XOR2 (N227, N224, N47);
nand NAND4 (N228, N208, N213, N209, N91);
and AND2 (N229, N226, N205);
xor XOR2 (N230, N216, N116);
nor NOR2 (N231, N72, N74);
xor XOR2 (N232, N231, N198);
buf BUF1 (N233, N225);
and AND4 (N234, N223, N109, N5, N162);
or OR4 (N235, N232, N234, N139, N221);
and AND3 (N236, N48, N101, N139);
nor NOR3 (N237, N236, N96, N169);
nand NAND4 (N238, N229, N236, N193, N109);
nor NOR4 (N239, N233, N50, N177, N70);
xor XOR2 (N240, N235, N197);
buf BUF1 (N241, N238);
xor XOR2 (N242, N220, N92);
nor NOR3 (N243, N241, N214, N39);
buf BUF1 (N244, N227);
and AND3 (N245, N244, N75, N170);
not NOT1 (N246, N240);
xor XOR2 (N247, N243, N65);
xor XOR2 (N248, N237, N44);
nor NOR4 (N249, N247, N166, N148, N166);
not NOT1 (N250, N215);
buf BUF1 (N251, N242);
and AND2 (N252, N251, N156);
xor XOR2 (N253, N228, N227);
nor NOR4 (N254, N253, N193, N130, N235);
not NOT1 (N255, N230);
not NOT1 (N256, N255);
nor NOR4 (N257, N250, N228, N52, N66);
nand NAND2 (N258, N246, N236);
nor NOR2 (N259, N252, N118);
buf BUF1 (N260, N190);
buf BUF1 (N261, N239);
or OR2 (N262, N248, N37);
or OR4 (N263, N256, N205, N147, N170);
buf BUF1 (N264, N249);
xor XOR2 (N265, N264, N185);
not NOT1 (N266, N245);
nand NAND2 (N267, N257, N178);
nand NAND3 (N268, N260, N252, N246);
nor NOR3 (N269, N268, N181, N92);
not NOT1 (N270, N269);
or OR4 (N271, N270, N240, N113, N89);
or OR4 (N272, N271, N80, N183, N181);
and AND4 (N273, N258, N50, N47, N198);
nand NAND3 (N274, N267, N7, N178);
and AND3 (N275, N263, N62, N199);
xor XOR2 (N276, N272, N220);
xor XOR2 (N277, N254, N175);
xor XOR2 (N278, N262, N63);
or OR2 (N279, N259, N74);
nand NAND2 (N280, N277, N233);
nor NOR2 (N281, N273, N81);
not NOT1 (N282, N266);
nand NAND2 (N283, N265, N225);
xor XOR2 (N284, N276, N233);
xor XOR2 (N285, N278, N122);
or OR2 (N286, N281, N274);
nor NOR3 (N287, N118, N217, N111);
xor XOR2 (N288, N284, N200);
nor NOR4 (N289, N285, N22, N19, N219);
xor XOR2 (N290, N288, N261);
or OR2 (N291, N202, N157);
and AND4 (N292, N291, N33, N279, N81);
xor XOR2 (N293, N201, N172);
or OR4 (N294, N286, N39, N43, N10);
buf BUF1 (N295, N292);
nor NOR3 (N296, N283, N284, N134);
or OR2 (N297, N280, N149);
buf BUF1 (N298, N289);
nand NAND4 (N299, N294, N33, N190, N121);
or OR2 (N300, N298, N89);
xor XOR2 (N301, N275, N40);
and AND3 (N302, N299, N198, N195);
xor XOR2 (N303, N295, N13);
or OR3 (N304, N282, N101, N195);
nand NAND4 (N305, N290, N115, N294, N118);
nor NOR4 (N306, N297, N21, N229, N248);
and AND2 (N307, N287, N125);
nor NOR2 (N308, N302, N6);
nand NAND3 (N309, N304, N292, N30);
nand NAND4 (N310, N296, N129, N148, N167);
nand NAND2 (N311, N300, N180);
xor XOR2 (N312, N308, N304);
xor XOR2 (N313, N312, N306);
and AND3 (N314, N46, N126, N210);
nor NOR3 (N315, N303, N150, N166);
nor NOR4 (N316, N309, N208, N150, N306);
nand NAND2 (N317, N293, N78);
and AND3 (N318, N305, N100, N24);
nor NOR3 (N319, N314, N314, N316);
buf BUF1 (N320, N210);
not NOT1 (N321, N319);
or OR3 (N322, N318, N50, N220);
or OR3 (N323, N310, N275, N149);
nand NAND3 (N324, N301, N61, N149);
nand NAND3 (N325, N317, N247, N201);
nor NOR4 (N326, N322, N75, N223, N145);
not NOT1 (N327, N315);
and AND3 (N328, N311, N65, N166);
xor XOR2 (N329, N323, N157);
and AND4 (N330, N329, N212, N314, N68);
not NOT1 (N331, N307);
not NOT1 (N332, N327);
nor NOR3 (N333, N332, N142, N40);
nand NAND4 (N334, N325, N10, N265, N303);
nor NOR4 (N335, N313, N330, N140, N79);
buf BUF1 (N336, N224);
xor XOR2 (N337, N335, N75);
nand NAND4 (N338, N321, N305, N41, N184);
not NOT1 (N339, N326);
and AND4 (N340, N331, N270, N287, N89);
or OR2 (N341, N334, N9);
or OR2 (N342, N320, N75);
buf BUF1 (N343, N328);
buf BUF1 (N344, N343);
nand NAND3 (N345, N337, N320, N75);
and AND3 (N346, N341, N12, N341);
nand NAND3 (N347, N342, N239, N143);
or OR2 (N348, N333, N74);
nor NOR3 (N349, N336, N133, N67);
nor NOR2 (N350, N349, N183);
buf BUF1 (N351, N346);
buf BUF1 (N352, N347);
and AND2 (N353, N351, N105);
buf BUF1 (N354, N352);
and AND2 (N355, N324, N47);
not NOT1 (N356, N339);
buf BUF1 (N357, N345);
and AND4 (N358, N356, N150, N301, N32);
and AND4 (N359, N340, N106, N235, N309);
xor XOR2 (N360, N354, N13);
buf BUF1 (N361, N338);
or OR2 (N362, N357, N29);
xor XOR2 (N363, N348, N106);
and AND2 (N364, N362, N179);
not NOT1 (N365, N363);
xor XOR2 (N366, N358, N60);
not NOT1 (N367, N344);
buf BUF1 (N368, N355);
xor XOR2 (N369, N368, N170);
or OR2 (N370, N359, N181);
nor NOR4 (N371, N370, N327, N35, N256);
not NOT1 (N372, N350);
buf BUF1 (N373, N371);
nand NAND3 (N374, N367, N187, N267);
nor NOR4 (N375, N360, N166, N81, N281);
nor NOR4 (N376, N369, N315, N276, N328);
nor NOR3 (N377, N376, N213, N302);
buf BUF1 (N378, N366);
and AND4 (N379, N378, N272, N56, N105);
or OR4 (N380, N379, N61, N330, N57);
nor NOR3 (N381, N365, N133, N85);
xor XOR2 (N382, N372, N343);
or OR2 (N383, N364, N108);
xor XOR2 (N384, N373, N214);
or OR2 (N385, N384, N55);
or OR2 (N386, N374, N135);
and AND2 (N387, N386, N222);
and AND2 (N388, N383, N59);
buf BUF1 (N389, N380);
or OR2 (N390, N361, N311);
or OR2 (N391, N390, N358);
nor NOR2 (N392, N391, N132);
buf BUF1 (N393, N353);
and AND2 (N394, N387, N255);
nor NOR2 (N395, N375, N266);
buf BUF1 (N396, N392);
xor XOR2 (N397, N377, N88);
nand NAND3 (N398, N395, N53, N258);
or OR2 (N399, N388, N35);
or OR3 (N400, N381, N46, N36);
buf BUF1 (N401, N398);
xor XOR2 (N402, N400, N211);
xor XOR2 (N403, N396, N364);
nand NAND2 (N404, N385, N339);
or OR4 (N405, N382, N159, N128, N276);
nand NAND3 (N406, N403, N162, N118);
buf BUF1 (N407, N393);
xor XOR2 (N408, N406, N247);
buf BUF1 (N409, N404);
buf BUF1 (N410, N402);
xor XOR2 (N411, N399, N265);
xor XOR2 (N412, N401, N255);
buf BUF1 (N413, N389);
and AND4 (N414, N408, N277, N273, N406);
or OR3 (N415, N397, N22, N146);
buf BUF1 (N416, N410);
not NOT1 (N417, N407);
not NOT1 (N418, N417);
not NOT1 (N419, N416);
buf BUF1 (N420, N405);
or OR2 (N421, N413, N44);
and AND4 (N422, N414, N397, N151, N43);
buf BUF1 (N423, N421);
nor NOR2 (N424, N423, N422);
buf BUF1 (N425, N143);
nand NAND4 (N426, N420, N115, N177, N390);
and AND4 (N427, N424, N362, N184, N366);
or OR2 (N428, N427, N347);
and AND3 (N429, N428, N383, N406);
nor NOR3 (N430, N425, N322, N56);
or OR2 (N431, N415, N214);
or OR2 (N432, N411, N146);
or OR4 (N433, N419, N93, N351, N352);
xor XOR2 (N434, N412, N111);
nand NAND3 (N435, N418, N140, N242);
not NOT1 (N436, N426);
or OR4 (N437, N433, N275, N35, N219);
not NOT1 (N438, N429);
nand NAND2 (N439, N394, N351);
buf BUF1 (N440, N435);
buf BUF1 (N441, N432);
buf BUF1 (N442, N434);
and AND4 (N443, N431, N149, N235, N276);
and AND4 (N444, N409, N26, N243, N256);
nand NAND2 (N445, N442, N414);
not NOT1 (N446, N430);
buf BUF1 (N447, N438);
buf BUF1 (N448, N440);
not NOT1 (N449, N447);
buf BUF1 (N450, N439);
nand NAND4 (N451, N441, N445, N11, N211);
not NOT1 (N452, N372);
nand NAND3 (N453, N443, N216, N368);
xor XOR2 (N454, N453, N121);
and AND3 (N455, N454, N89, N391);
buf BUF1 (N456, N449);
xor XOR2 (N457, N451, N254);
nor NOR4 (N458, N436, N142, N219, N81);
not NOT1 (N459, N452);
nor NOR2 (N460, N455, N416);
nor NOR3 (N461, N446, N205, N160);
buf BUF1 (N462, N437);
buf BUF1 (N463, N461);
and AND2 (N464, N460, N300);
not NOT1 (N465, N444);
nor NOR2 (N466, N463, N195);
xor XOR2 (N467, N459, N67);
or OR3 (N468, N467, N420, N422);
and AND4 (N469, N465, N261, N36, N252);
xor XOR2 (N470, N450, N240);
nand NAND2 (N471, N468, N274);
not NOT1 (N472, N448);
or OR3 (N473, N470, N367, N438);
buf BUF1 (N474, N464);
xor XOR2 (N475, N457, N423);
xor XOR2 (N476, N462, N397);
xor XOR2 (N477, N475, N462);
and AND4 (N478, N473, N237, N98, N446);
or OR3 (N479, N471, N133, N178);
nor NOR4 (N480, N477, N371, N153, N380);
nand NAND3 (N481, N472, N362, N202);
not NOT1 (N482, N466);
nor NOR2 (N483, N481, N271);
xor XOR2 (N484, N476, N33);
not NOT1 (N485, N456);
buf BUF1 (N486, N483);
buf BUF1 (N487, N478);
or OR3 (N488, N474, N305, N272);
not NOT1 (N489, N480);
nand NAND3 (N490, N482, N176, N4);
xor XOR2 (N491, N484, N118);
nand NAND3 (N492, N488, N94, N236);
buf BUF1 (N493, N469);
or OR3 (N494, N493, N354, N392);
buf BUF1 (N495, N485);
and AND2 (N496, N458, N320);
xor XOR2 (N497, N492, N145);
xor XOR2 (N498, N497, N248);
and AND2 (N499, N487, N34);
buf BUF1 (N500, N486);
buf BUF1 (N501, N499);
nor NOR4 (N502, N496, N221, N249, N310);
not NOT1 (N503, N501);
nor NOR3 (N504, N500, N177, N60);
or OR2 (N505, N479, N119);
not NOT1 (N506, N494);
nor NOR2 (N507, N505, N381);
or OR4 (N508, N490, N338, N139, N367);
xor XOR2 (N509, N502, N414);
nor NOR3 (N510, N508, N503, N343);
and AND3 (N511, N199, N394, N321);
not NOT1 (N512, N511);
buf BUF1 (N513, N512);
nor NOR4 (N514, N506, N276, N496, N483);
and AND4 (N515, N498, N301, N250, N33);
and AND2 (N516, N491, N443);
not NOT1 (N517, N504);
xor XOR2 (N518, N495, N373);
nor NOR4 (N519, N509, N159, N25, N218);
xor XOR2 (N520, N514, N443);
xor XOR2 (N521, N489, N42);
nand NAND4 (N522, N521, N227, N22, N271);
buf BUF1 (N523, N516);
xor XOR2 (N524, N520, N7);
buf BUF1 (N525, N510);
or OR4 (N526, N525, N160, N392, N485);
and AND2 (N527, N524, N64);
nand NAND3 (N528, N513, N142, N193);
or OR2 (N529, N527, N88);
xor XOR2 (N530, N519, N322);
not NOT1 (N531, N522);
buf BUF1 (N532, N515);
and AND4 (N533, N530, N181, N370, N103);
not NOT1 (N534, N529);
not NOT1 (N535, N528);
nor NOR2 (N536, N517, N509);
xor XOR2 (N537, N531, N420);
nor NOR4 (N538, N523, N406, N372, N189);
and AND4 (N539, N532, N9, N17, N390);
nor NOR2 (N540, N533, N285);
xor XOR2 (N541, N536, N147);
buf BUF1 (N542, N518);
nand NAND4 (N543, N537, N210, N81, N218);
nor NOR4 (N544, N543, N423, N242, N199);
buf BUF1 (N545, N535);
nand NAND4 (N546, N526, N219, N82, N191);
or OR2 (N547, N541, N30);
or OR4 (N548, N540, N251, N448, N220);
nand NAND3 (N549, N546, N530, N34);
and AND4 (N550, N534, N50, N504, N165);
buf BUF1 (N551, N550);
buf BUF1 (N552, N544);
xor XOR2 (N553, N545, N63);
xor XOR2 (N554, N549, N196);
and AND4 (N555, N548, N290, N445, N267);
nor NOR3 (N556, N547, N421, N195);
buf BUF1 (N557, N554);
nand NAND3 (N558, N538, N281, N396);
xor XOR2 (N559, N556, N137);
not NOT1 (N560, N557);
buf BUF1 (N561, N551);
xor XOR2 (N562, N559, N396);
or OR3 (N563, N562, N100, N32);
and AND2 (N564, N539, N54);
nor NOR4 (N565, N553, N82, N362, N464);
or OR3 (N566, N560, N393, N394);
and AND3 (N567, N566, N7, N86);
or OR4 (N568, N563, N416, N29, N445);
nor NOR3 (N569, N558, N166, N125);
not NOT1 (N570, N561);
buf BUF1 (N571, N555);
and AND4 (N572, N568, N217, N114, N470);
or OR4 (N573, N565, N33, N409, N132);
nand NAND4 (N574, N572, N113, N292, N520);
and AND2 (N575, N569, N168);
or OR4 (N576, N567, N207, N114, N47);
xor XOR2 (N577, N574, N415);
xor XOR2 (N578, N576, N471);
nand NAND3 (N579, N577, N294, N436);
nor NOR4 (N580, N552, N471, N536, N310);
buf BUF1 (N581, N575);
or OR4 (N582, N579, N324, N201, N304);
or OR2 (N583, N570, N176);
or OR3 (N584, N571, N512, N324);
xor XOR2 (N585, N578, N254);
not NOT1 (N586, N582);
and AND2 (N587, N564, N194);
not NOT1 (N588, N573);
nand NAND2 (N589, N586, N408);
nand NAND4 (N590, N507, N10, N553, N513);
and AND4 (N591, N584, N283, N81, N315);
not NOT1 (N592, N589);
nor NOR2 (N593, N590, N415);
nor NOR4 (N594, N587, N61, N587, N153);
or OR2 (N595, N594, N330);
nand NAND3 (N596, N592, N379, N361);
nor NOR3 (N597, N542, N76, N494);
xor XOR2 (N598, N595, N355);
buf BUF1 (N599, N583);
xor XOR2 (N600, N593, N155);
nor NOR3 (N601, N588, N523, N129);
nand NAND3 (N602, N580, N11, N515);
or OR4 (N603, N600, N224, N542, N137);
buf BUF1 (N604, N596);
buf BUF1 (N605, N604);
not NOT1 (N606, N603);
nand NAND4 (N607, N585, N143, N311, N96);
nor NOR4 (N608, N599, N385, N155, N209);
or OR3 (N609, N605, N208, N474);
and AND2 (N610, N597, N190);
or OR4 (N611, N607, N28, N32, N356);
not NOT1 (N612, N606);
and AND4 (N613, N601, N586, N197, N299);
not NOT1 (N614, N598);
or OR2 (N615, N614, N188);
and AND2 (N616, N611, N566);
buf BUF1 (N617, N581);
nand NAND4 (N618, N617, N304, N507, N272);
buf BUF1 (N619, N616);
or OR2 (N620, N610, N208);
or OR3 (N621, N591, N496, N348);
buf BUF1 (N622, N613);
not NOT1 (N623, N612);
and AND3 (N624, N623, N38, N55);
or OR4 (N625, N621, N212, N106, N52);
buf BUF1 (N626, N620);
xor XOR2 (N627, N609, N385);
or OR2 (N628, N627, N196);
or OR2 (N629, N608, N433);
xor XOR2 (N630, N628, N321);
nor NOR4 (N631, N622, N410, N114, N522);
or OR2 (N632, N625, N119);
nor NOR2 (N633, N618, N237);
nor NOR3 (N634, N619, N85, N240);
xor XOR2 (N635, N602, N432);
or OR4 (N636, N624, N433, N249, N190);
xor XOR2 (N637, N634, N46);
buf BUF1 (N638, N637);
or OR3 (N639, N615, N18, N74);
and AND2 (N640, N633, N183);
and AND2 (N641, N638, N593);
nor NOR2 (N642, N636, N313);
xor XOR2 (N643, N641, N348);
nor NOR2 (N644, N631, N360);
xor XOR2 (N645, N643, N284);
nor NOR3 (N646, N644, N515, N362);
buf BUF1 (N647, N645);
nand NAND3 (N648, N629, N536, N103);
nand NAND3 (N649, N647, N399, N234);
xor XOR2 (N650, N642, N555);
nand NAND3 (N651, N632, N306, N80);
nand NAND2 (N652, N650, N221);
buf BUF1 (N653, N630);
not NOT1 (N654, N652);
not NOT1 (N655, N640);
and AND4 (N656, N635, N367, N520, N252);
and AND3 (N657, N626, N338, N60);
or OR2 (N658, N655, N651);
and AND3 (N659, N505, N534, N529);
nor NOR2 (N660, N639, N190);
nor NOR4 (N661, N656, N176, N432, N80);
not NOT1 (N662, N649);
nand NAND3 (N663, N662, N49, N405);
nand NAND4 (N664, N654, N538, N407, N263);
nor NOR4 (N665, N657, N646, N364, N260);
buf BUF1 (N666, N100);
or OR2 (N667, N660, N361);
or OR3 (N668, N665, N54, N403);
not NOT1 (N669, N666);
and AND3 (N670, N648, N169, N67);
nand NAND3 (N671, N669, N27, N615);
buf BUF1 (N672, N661);
nor NOR4 (N673, N668, N64, N229, N448);
nand NAND4 (N674, N667, N337, N131, N7);
not NOT1 (N675, N674);
buf BUF1 (N676, N663);
buf BUF1 (N677, N664);
buf BUF1 (N678, N671);
xor XOR2 (N679, N673, N59);
nand NAND2 (N680, N658, N645);
or OR4 (N681, N678, N399, N429, N95);
buf BUF1 (N682, N672);
nand NAND3 (N683, N679, N176, N256);
or OR4 (N684, N681, N371, N160, N461);
not NOT1 (N685, N682);
and AND4 (N686, N675, N296, N254, N317);
not NOT1 (N687, N686);
or OR4 (N688, N680, N615, N631, N99);
nand NAND3 (N689, N688, N99, N321);
and AND2 (N690, N670, N324);
nand NAND3 (N691, N677, N428, N484);
not NOT1 (N692, N685);
or OR4 (N693, N687, N277, N93, N523);
nand NAND3 (N694, N653, N661, N351);
xor XOR2 (N695, N692, N328);
xor XOR2 (N696, N659, N46);
xor XOR2 (N697, N696, N210);
buf BUF1 (N698, N683);
not NOT1 (N699, N698);
xor XOR2 (N700, N697, N490);
not NOT1 (N701, N700);
nand NAND3 (N702, N694, N45, N414);
buf BUF1 (N703, N691);
not NOT1 (N704, N676);
or OR2 (N705, N689, N650);
nor NOR4 (N706, N701, N253, N408, N286);
buf BUF1 (N707, N706);
buf BUF1 (N708, N705);
not NOT1 (N709, N704);
buf BUF1 (N710, N690);
nor NOR4 (N711, N702, N218, N633, N94);
xor XOR2 (N712, N699, N125);
not NOT1 (N713, N695);
xor XOR2 (N714, N711, N185);
not NOT1 (N715, N714);
nand NAND3 (N716, N709, N142, N73);
or OR2 (N717, N707, N534);
and AND2 (N718, N715, N66);
buf BUF1 (N719, N712);
or OR4 (N720, N693, N41, N476, N200);
and AND2 (N721, N713, N203);
or OR3 (N722, N703, N85, N82);
buf BUF1 (N723, N719);
and AND2 (N724, N720, N454);
nor NOR4 (N725, N718, N342, N116, N551);
not NOT1 (N726, N708);
not NOT1 (N727, N726);
nor NOR2 (N728, N710, N605);
nand NAND2 (N729, N723, N225);
nand NAND4 (N730, N717, N567, N504, N712);
xor XOR2 (N731, N729, N309);
nor NOR3 (N732, N684, N661, N568);
and AND4 (N733, N728, N23, N415, N676);
buf BUF1 (N734, N730);
not NOT1 (N735, N724);
and AND2 (N736, N716, N208);
or OR2 (N737, N731, N486);
not NOT1 (N738, N734);
buf BUF1 (N739, N737);
not NOT1 (N740, N732);
and AND4 (N741, N722, N192, N259, N523);
xor XOR2 (N742, N738, N673);
and AND2 (N743, N727, N702);
buf BUF1 (N744, N725);
or OR3 (N745, N743, N341, N69);
nor NOR4 (N746, N721, N490, N423, N173);
nand NAND2 (N747, N739, N649);
not NOT1 (N748, N742);
not NOT1 (N749, N735);
nor NOR3 (N750, N745, N610, N635);
and AND2 (N751, N744, N298);
or OR4 (N752, N733, N204, N238, N580);
and AND4 (N753, N748, N738, N505, N286);
and AND2 (N754, N751, N129);
and AND4 (N755, N747, N180, N651, N471);
nor NOR2 (N756, N750, N87);
buf BUF1 (N757, N755);
buf BUF1 (N758, N753);
nor NOR2 (N759, N757, N287);
xor XOR2 (N760, N741, N734);
and AND3 (N761, N736, N315, N494);
or OR3 (N762, N754, N138, N458);
not NOT1 (N763, N749);
or OR3 (N764, N740, N114, N490);
xor XOR2 (N765, N763, N760);
nor NOR3 (N766, N101, N59, N500);
nand NAND4 (N767, N756, N57, N469, N553);
not NOT1 (N768, N759);
or OR4 (N769, N746, N64, N423, N493);
or OR3 (N770, N765, N526, N78);
nor NOR2 (N771, N764, N666);
or OR2 (N772, N768, N178);
or OR2 (N773, N758, N142);
and AND2 (N774, N767, N675);
nor NOR3 (N775, N769, N204, N522);
and AND4 (N776, N770, N251, N186, N707);
and AND3 (N777, N762, N184, N86);
nand NAND2 (N778, N752, N776);
not NOT1 (N779, N233);
nor NOR4 (N780, N772, N96, N387, N235);
buf BUF1 (N781, N780);
xor XOR2 (N782, N779, N642);
not NOT1 (N783, N771);
buf BUF1 (N784, N773);
and AND2 (N785, N777, N552);
nor NOR3 (N786, N783, N557, N672);
not NOT1 (N787, N775);
buf BUF1 (N788, N761);
or OR3 (N789, N781, N379, N726);
buf BUF1 (N790, N784);
and AND4 (N791, N788, N733, N3, N473);
nand NAND4 (N792, N787, N45, N376, N113);
xor XOR2 (N793, N789, N543);
and AND4 (N794, N766, N771, N132, N550);
nor NOR3 (N795, N782, N380, N555);
or OR3 (N796, N774, N655, N269);
not NOT1 (N797, N790);
or OR3 (N798, N785, N797, N97);
not NOT1 (N799, N474);
buf BUF1 (N800, N796);
nand NAND4 (N801, N795, N248, N792, N489);
nor NOR4 (N802, N300, N632, N642, N563);
buf BUF1 (N803, N794);
buf BUF1 (N804, N791);
not NOT1 (N805, N778);
and AND3 (N806, N805, N59, N86);
xor XOR2 (N807, N786, N734);
buf BUF1 (N808, N800);
not NOT1 (N809, N804);
nand NAND2 (N810, N807, N16);
buf BUF1 (N811, N793);
not NOT1 (N812, N799);
buf BUF1 (N813, N810);
and AND4 (N814, N808, N456, N590, N792);
not NOT1 (N815, N812);
not NOT1 (N816, N802);
nor NOR4 (N817, N806, N349, N66, N468);
buf BUF1 (N818, N801);
xor XOR2 (N819, N816, N16);
nand NAND4 (N820, N818, N235, N329, N546);
buf BUF1 (N821, N817);
not NOT1 (N822, N821);
xor XOR2 (N823, N814, N502);
nand NAND3 (N824, N820, N804, N279);
not NOT1 (N825, N809);
and AND2 (N826, N819, N231);
nor NOR4 (N827, N798, N459, N297, N71);
and AND4 (N828, N825, N266, N202, N17);
nor NOR2 (N829, N824, N818);
nor NOR3 (N830, N828, N450, N117);
xor XOR2 (N831, N811, N89);
nand NAND3 (N832, N803, N566, N7);
not NOT1 (N833, N831);
buf BUF1 (N834, N826);
buf BUF1 (N835, N822);
nor NOR4 (N836, N832, N148, N732, N227);
or OR4 (N837, N835, N434, N537, N400);
xor XOR2 (N838, N823, N247);
xor XOR2 (N839, N834, N137);
nor NOR2 (N840, N837, N152);
nand NAND4 (N841, N839, N527, N341, N645);
or OR4 (N842, N841, N160, N750, N136);
or OR4 (N843, N836, N598, N327, N344);
nor NOR4 (N844, N840, N452, N588, N728);
buf BUF1 (N845, N844);
xor XOR2 (N846, N833, N306);
nand NAND3 (N847, N815, N75, N390);
or OR3 (N848, N846, N416, N627);
nand NAND2 (N849, N830, N695);
nor NOR2 (N850, N848, N186);
or OR2 (N851, N842, N774);
and AND3 (N852, N850, N528, N28);
nand NAND2 (N853, N813, N612);
buf BUF1 (N854, N849);
nand NAND4 (N855, N827, N119, N415, N624);
xor XOR2 (N856, N852, N18);
nand NAND3 (N857, N851, N458, N828);
buf BUF1 (N858, N854);
buf BUF1 (N859, N838);
nand NAND4 (N860, N853, N339, N252, N746);
not NOT1 (N861, N845);
nor NOR4 (N862, N856, N315, N510, N459);
xor XOR2 (N863, N855, N395);
nand NAND3 (N864, N857, N783, N561);
or OR4 (N865, N862, N315, N458, N244);
xor XOR2 (N866, N843, N194);
and AND2 (N867, N860, N214);
buf BUF1 (N868, N858);
and AND3 (N869, N847, N113, N164);
nand NAND4 (N870, N865, N88, N440, N660);
nor NOR4 (N871, N829, N748, N432, N664);
or OR3 (N872, N866, N660, N435);
not NOT1 (N873, N861);
buf BUF1 (N874, N873);
buf BUF1 (N875, N869);
and AND4 (N876, N863, N308, N274, N735);
not NOT1 (N877, N874);
xor XOR2 (N878, N859, N30);
not NOT1 (N879, N877);
nand NAND2 (N880, N876, N877);
not NOT1 (N881, N868);
buf BUF1 (N882, N871);
not NOT1 (N883, N867);
xor XOR2 (N884, N864, N33);
nor NOR3 (N885, N881, N722, N604);
or OR4 (N886, N884, N731, N466, N210);
and AND4 (N887, N870, N569, N729, N227);
not NOT1 (N888, N880);
not NOT1 (N889, N882);
not NOT1 (N890, N875);
nor NOR4 (N891, N886, N582, N230, N449);
buf BUF1 (N892, N890);
and AND4 (N893, N887, N71, N747, N404);
nand NAND4 (N894, N888, N799, N752, N177);
buf BUF1 (N895, N879);
nand NAND3 (N896, N892, N267, N363);
and AND3 (N897, N889, N677, N741);
and AND3 (N898, N885, N132, N99);
nor NOR3 (N899, N894, N258, N600);
and AND3 (N900, N891, N345, N384);
and AND3 (N901, N899, N441, N877);
xor XOR2 (N902, N901, N647);
xor XOR2 (N903, N872, N448);
or OR3 (N904, N897, N618, N335);
buf BUF1 (N905, N900);
not NOT1 (N906, N883);
nand NAND2 (N907, N896, N181);
and AND3 (N908, N878, N188, N577);
nand NAND2 (N909, N905, N794);
xor XOR2 (N910, N904, N892);
nor NOR2 (N911, N908, N170);
nor NOR3 (N912, N906, N305, N562);
not NOT1 (N913, N910);
nand NAND4 (N914, N913, N187, N647, N872);
nand NAND2 (N915, N914, N911);
xor XOR2 (N916, N191, N286);
nand NAND4 (N917, N893, N643, N604, N235);
and AND3 (N918, N917, N286, N837);
not NOT1 (N919, N902);
not NOT1 (N920, N903);
not NOT1 (N921, N920);
nand NAND2 (N922, N898, N492);
not NOT1 (N923, N907);
nand NAND3 (N924, N895, N71, N691);
and AND4 (N925, N921, N662, N261, N156);
nand NAND3 (N926, N916, N316, N865);
buf BUF1 (N927, N925);
nor NOR3 (N928, N922, N577, N47);
nand NAND3 (N929, N918, N379, N918);
and AND4 (N930, N926, N58, N568, N169);
xor XOR2 (N931, N929, N875);
buf BUF1 (N932, N927);
xor XOR2 (N933, N930, N51);
xor XOR2 (N934, N932, N312);
nor NOR4 (N935, N923, N272, N520, N8);
nand NAND3 (N936, N909, N599, N273);
nor NOR3 (N937, N919, N339, N258);
and AND2 (N938, N935, N892);
nor NOR2 (N939, N928, N5);
nor NOR4 (N940, N939, N438, N812, N607);
xor XOR2 (N941, N924, N107);
nor NOR4 (N942, N938, N331, N350, N206);
xor XOR2 (N943, N933, N499);
and AND2 (N944, N934, N409);
nand NAND2 (N945, N943, N187);
xor XOR2 (N946, N941, N97);
xor XOR2 (N947, N946, N131);
xor XOR2 (N948, N931, N213);
buf BUF1 (N949, N915);
and AND2 (N950, N940, N211);
or OR4 (N951, N942, N148, N773, N891);
or OR4 (N952, N945, N609, N604, N17);
or OR2 (N953, N937, N219);
or OR4 (N954, N948, N406, N626, N459);
not NOT1 (N955, N951);
xor XOR2 (N956, N912, N4);
nor NOR2 (N957, N954, N651);
and AND2 (N958, N936, N290);
xor XOR2 (N959, N958, N504);
nand NAND4 (N960, N952, N426, N178, N64);
nor NOR2 (N961, N957, N653);
nand NAND3 (N962, N960, N93, N428);
or OR4 (N963, N961, N23, N102, N507);
nor NOR3 (N964, N959, N330, N204);
or OR3 (N965, N956, N718, N569);
nand NAND4 (N966, N953, N524, N792, N207);
nor NOR2 (N967, N962, N623);
xor XOR2 (N968, N955, N231);
and AND2 (N969, N966, N595);
xor XOR2 (N970, N950, N662);
nand NAND4 (N971, N963, N569, N157, N408);
nor NOR2 (N972, N971, N407);
buf BUF1 (N973, N969);
not NOT1 (N974, N972);
xor XOR2 (N975, N974, N376);
nand NAND2 (N976, N970, N748);
nor NOR2 (N977, N975, N46);
not NOT1 (N978, N977);
nor NOR2 (N979, N976, N384);
and AND2 (N980, N944, N540);
and AND2 (N981, N980, N266);
buf BUF1 (N982, N949);
or OR4 (N983, N965, N300, N676, N580);
nor NOR3 (N984, N964, N943, N269);
nand NAND4 (N985, N947, N564, N427, N925);
and AND4 (N986, N968, N168, N307, N145);
nor NOR3 (N987, N982, N398, N513);
buf BUF1 (N988, N987);
nor NOR4 (N989, N981, N382, N960, N142);
nand NAND2 (N990, N989, N47);
buf BUF1 (N991, N990);
not NOT1 (N992, N988);
nand NAND4 (N993, N992, N981, N970, N200);
buf BUF1 (N994, N983);
or OR2 (N995, N979, N319);
buf BUF1 (N996, N984);
or OR4 (N997, N967, N176, N261, N448);
buf BUF1 (N998, N993);
buf BUF1 (N999, N996);
and AND2 (N1000, N999, N610);
xor XOR2 (N1001, N986, N272);
nor NOR3 (N1002, N998, N521, N808);
nor NOR3 (N1003, N1001, N630, N506);
and AND4 (N1004, N1003, N469, N840, N331);
not NOT1 (N1005, N973);
xor XOR2 (N1006, N1000, N433);
xor XOR2 (N1007, N1002, N765);
xor XOR2 (N1008, N991, N843);
or OR2 (N1009, N1005, N127);
nand NAND3 (N1010, N985, N315, N456);
and AND3 (N1011, N995, N392, N86);
nand NAND2 (N1012, N1008, N238);
buf BUF1 (N1013, N994);
nor NOR4 (N1014, N1011, N16, N423, N627);
buf BUF1 (N1015, N1006);
not NOT1 (N1016, N1012);
nand NAND2 (N1017, N978, N938);
buf BUF1 (N1018, N1004);
nor NOR3 (N1019, N1007, N807, N706);
and AND2 (N1020, N1016, N610);
or OR2 (N1021, N1013, N559);
nor NOR4 (N1022, N1010, N549, N704, N347);
nand NAND2 (N1023, N1020, N940);
xor XOR2 (N1024, N1014, N983);
buf BUF1 (N1025, N1024);
or OR4 (N1026, N1009, N972, N845, N1000);
xor XOR2 (N1027, N1025, N64);
and AND2 (N1028, N1018, N593);
xor XOR2 (N1029, N1019, N539);
nand NAND2 (N1030, N1017, N221);
xor XOR2 (N1031, N1026, N942);
nand NAND3 (N1032, N1030, N108, N134);
buf BUF1 (N1033, N1028);
nor NOR3 (N1034, N1027, N539, N734);
or OR3 (N1035, N1015, N115, N797);
xor XOR2 (N1036, N1034, N593);
not NOT1 (N1037, N1035);
nor NOR4 (N1038, N997, N95, N286, N792);
xor XOR2 (N1039, N1031, N98);
or OR2 (N1040, N1039, N159);
or OR3 (N1041, N1022, N983, N324);
not NOT1 (N1042, N1029);
xor XOR2 (N1043, N1042, N322);
or OR3 (N1044, N1036, N732, N250);
buf BUF1 (N1045, N1037);
buf BUF1 (N1046, N1038);
nand NAND3 (N1047, N1021, N221, N112);
nand NAND2 (N1048, N1032, N666);
not NOT1 (N1049, N1046);
xor XOR2 (N1050, N1047, N902);
or OR2 (N1051, N1033, N254);
xor XOR2 (N1052, N1045, N219);
not NOT1 (N1053, N1050);
nor NOR4 (N1054, N1051, N662, N1002, N520);
nor NOR2 (N1055, N1048, N911);
nor NOR2 (N1056, N1049, N685);
nor NOR2 (N1057, N1055, N825);
buf BUF1 (N1058, N1043);
or OR2 (N1059, N1023, N608);
and AND2 (N1060, N1053, N2);
not NOT1 (N1061, N1040);
nand NAND4 (N1062, N1056, N39, N48, N464);
buf BUF1 (N1063, N1041);
not NOT1 (N1064, N1058);
nand NAND3 (N1065, N1057, N105, N379);
and AND2 (N1066, N1060, N730);
buf BUF1 (N1067, N1064);
or OR3 (N1068, N1065, N789, N112);
nor NOR4 (N1069, N1066, N152, N195, N1);
nor NOR3 (N1070, N1063, N814, N37);
and AND3 (N1071, N1044, N850, N723);
or OR4 (N1072, N1067, N98, N605, N488);
xor XOR2 (N1073, N1052, N642);
nand NAND3 (N1074, N1070, N301, N135);
nor NOR2 (N1075, N1054, N237);
nand NAND2 (N1076, N1074, N990);
buf BUF1 (N1077, N1059);
and AND2 (N1078, N1068, N252);
nand NAND3 (N1079, N1071, N753, N168);
nand NAND4 (N1080, N1062, N341, N187, N600);
nor NOR3 (N1081, N1079, N674, N880);
nand NAND2 (N1082, N1078, N658);
or OR3 (N1083, N1080, N411, N209);
and AND4 (N1084, N1073, N126, N134, N107);
not NOT1 (N1085, N1082);
nand NAND3 (N1086, N1084, N876, N804);
xor XOR2 (N1087, N1076, N749);
nor NOR3 (N1088, N1081, N805, N48);
or OR4 (N1089, N1087, N951, N49, N824);
not NOT1 (N1090, N1086);
not NOT1 (N1091, N1085);
or OR4 (N1092, N1075, N421, N544, N968);
not NOT1 (N1093, N1061);
buf BUF1 (N1094, N1093);
not NOT1 (N1095, N1089);
not NOT1 (N1096, N1088);
nor NOR2 (N1097, N1092, N730);
nand NAND3 (N1098, N1096, N26, N1084);
nor NOR3 (N1099, N1090, N489, N438);
or OR4 (N1100, N1094, N1079, N933, N428);
nor NOR2 (N1101, N1097, N448);
and AND3 (N1102, N1083, N118, N60);
not NOT1 (N1103, N1100);
or OR3 (N1104, N1102, N660, N456);
or OR2 (N1105, N1104, N851);
xor XOR2 (N1106, N1101, N82);
and AND2 (N1107, N1095, N248);
or OR2 (N1108, N1103, N1074);
or OR2 (N1109, N1105, N778);
buf BUF1 (N1110, N1099);
or OR3 (N1111, N1109, N75, N825);
or OR4 (N1112, N1072, N530, N950, N857);
or OR3 (N1113, N1111, N495, N517);
and AND3 (N1114, N1098, N408, N39);
not NOT1 (N1115, N1108);
buf BUF1 (N1116, N1110);
buf BUF1 (N1117, N1106);
nor NOR4 (N1118, N1117, N562, N1065, N760);
buf BUF1 (N1119, N1115);
nand NAND2 (N1120, N1069, N922);
not NOT1 (N1121, N1091);
xor XOR2 (N1122, N1120, N716);
nor NOR3 (N1123, N1122, N946, N564);
not NOT1 (N1124, N1077);
nand NAND2 (N1125, N1114, N818);
or OR4 (N1126, N1119, N323, N332, N1003);
buf BUF1 (N1127, N1107);
buf BUF1 (N1128, N1118);
or OR2 (N1129, N1116, N954);
not NOT1 (N1130, N1124);
not NOT1 (N1131, N1125);
not NOT1 (N1132, N1123);
nand NAND2 (N1133, N1131, N523);
and AND4 (N1134, N1127, N1068, N326, N1017);
xor XOR2 (N1135, N1126, N739);
or OR4 (N1136, N1121, N546, N204, N130);
or OR3 (N1137, N1136, N20, N721);
buf BUF1 (N1138, N1135);
xor XOR2 (N1139, N1138, N819);
xor XOR2 (N1140, N1113, N38);
nor NOR3 (N1141, N1128, N417, N881);
nor NOR4 (N1142, N1140, N711, N661, N681);
or OR2 (N1143, N1132, N705);
nor NOR2 (N1144, N1139, N482);
not NOT1 (N1145, N1112);
not NOT1 (N1146, N1134);
and AND2 (N1147, N1145, N193);
buf BUF1 (N1148, N1144);
xor XOR2 (N1149, N1143, N620);
buf BUF1 (N1150, N1146);
and AND3 (N1151, N1129, N473, N537);
not NOT1 (N1152, N1149);
or OR2 (N1153, N1151, N57);
buf BUF1 (N1154, N1152);
buf BUF1 (N1155, N1133);
buf BUF1 (N1156, N1148);
nand NAND3 (N1157, N1142, N1018, N1130);
and AND3 (N1158, N1055, N309, N304);
or OR4 (N1159, N1157, N1032, N904, N530);
and AND4 (N1160, N1155, N963, N191, N163);
and AND2 (N1161, N1156, N388);
buf BUF1 (N1162, N1158);
not NOT1 (N1163, N1161);
nand NAND2 (N1164, N1147, N1060);
xor XOR2 (N1165, N1160, N765);
nand NAND3 (N1166, N1165, N534, N181);
and AND4 (N1167, N1164, N82, N781, N235);
nor NOR4 (N1168, N1162, N351, N1116, N515);
buf BUF1 (N1169, N1137);
nor NOR3 (N1170, N1159, N592, N273);
nor NOR2 (N1171, N1154, N1061);
not NOT1 (N1172, N1166);
and AND3 (N1173, N1171, N953, N697);
nor NOR3 (N1174, N1173, N1063, N796);
or OR4 (N1175, N1172, N1166, N457, N699);
buf BUF1 (N1176, N1170);
buf BUF1 (N1177, N1153);
or OR2 (N1178, N1175, N74);
not NOT1 (N1179, N1174);
buf BUF1 (N1180, N1176);
xor XOR2 (N1181, N1141, N844);
and AND3 (N1182, N1163, N581, N29);
buf BUF1 (N1183, N1181);
not NOT1 (N1184, N1168);
not NOT1 (N1185, N1150);
and AND2 (N1186, N1185, N706);
not NOT1 (N1187, N1177);
nor NOR4 (N1188, N1184, N1166, N858, N746);
and AND4 (N1189, N1167, N273, N1020, N764);
nor NOR3 (N1190, N1169, N223, N1042);
nand NAND4 (N1191, N1179, N1048, N1113, N932);
nor NOR4 (N1192, N1186, N463, N70, N98);
or OR4 (N1193, N1190, N30, N536, N817);
nor NOR2 (N1194, N1188, N908);
and AND2 (N1195, N1187, N1059);
xor XOR2 (N1196, N1183, N572);
nor NOR2 (N1197, N1193, N1039);
or OR4 (N1198, N1192, N205, N523, N963);
and AND4 (N1199, N1191, N1094, N208, N272);
or OR4 (N1200, N1189, N943, N868, N1195);
nand NAND3 (N1201, N145, N388, N456);
xor XOR2 (N1202, N1182, N838);
xor XOR2 (N1203, N1197, N595);
nor NOR3 (N1204, N1199, N438, N1039);
xor XOR2 (N1205, N1201, N871);
nand NAND4 (N1206, N1202, N336, N794, N699);
nor NOR3 (N1207, N1196, N638, N150);
not NOT1 (N1208, N1207);
xor XOR2 (N1209, N1178, N534);
nand NAND3 (N1210, N1209, N538, N591);
or OR3 (N1211, N1208, N938, N132);
and AND2 (N1212, N1198, N839);
buf BUF1 (N1213, N1204);
or OR4 (N1214, N1180, N336, N749, N198);
or OR2 (N1215, N1214, N269);
not NOT1 (N1216, N1210);
and AND4 (N1217, N1216, N633, N648, N816);
not NOT1 (N1218, N1205);
or OR3 (N1219, N1212, N668, N1124);
not NOT1 (N1220, N1219);
nand NAND4 (N1221, N1211, N55, N963, N33);
nor NOR3 (N1222, N1218, N800, N738);
buf BUF1 (N1223, N1206);
nand NAND2 (N1224, N1220, N853);
nand NAND4 (N1225, N1217, N460, N1150, N1089);
or OR3 (N1226, N1194, N4, N792);
xor XOR2 (N1227, N1224, N257);
nor NOR4 (N1228, N1222, N204, N973, N785);
xor XOR2 (N1229, N1226, N668);
or OR4 (N1230, N1229, N807, N242, N526);
and AND2 (N1231, N1228, N620);
or OR4 (N1232, N1221, N207, N1213, N106);
not NOT1 (N1233, N633);
nand NAND2 (N1234, N1233, N519);
nand NAND4 (N1235, N1227, N964, N296, N311);
not NOT1 (N1236, N1235);
buf BUF1 (N1237, N1236);
not NOT1 (N1238, N1230);
nor NOR3 (N1239, N1225, N1061, N1077);
nor NOR4 (N1240, N1239, N245, N1212, N520);
buf BUF1 (N1241, N1237);
nand NAND2 (N1242, N1231, N334);
xor XOR2 (N1243, N1223, N86);
buf BUF1 (N1244, N1241);
buf BUF1 (N1245, N1234);
xor XOR2 (N1246, N1232, N26);
nand NAND3 (N1247, N1203, N214, N759);
buf BUF1 (N1248, N1215);
buf BUF1 (N1249, N1247);
not NOT1 (N1250, N1238);
xor XOR2 (N1251, N1240, N1177);
nand NAND2 (N1252, N1246, N691);
not NOT1 (N1253, N1249);
and AND4 (N1254, N1200, N324, N1159, N315);
xor XOR2 (N1255, N1251, N442);
nand NAND2 (N1256, N1252, N317);
and AND4 (N1257, N1245, N153, N705, N849);
or OR2 (N1258, N1253, N552);
or OR3 (N1259, N1243, N588, N491);
xor XOR2 (N1260, N1254, N360);
not NOT1 (N1261, N1244);
and AND3 (N1262, N1255, N441, N572);
xor XOR2 (N1263, N1257, N260);
and AND2 (N1264, N1259, N229);
and AND3 (N1265, N1256, N387, N602);
and AND3 (N1266, N1262, N1213, N35);
nand NAND4 (N1267, N1265, N703, N1253, N464);
not NOT1 (N1268, N1264);
or OR3 (N1269, N1258, N231, N1152);
not NOT1 (N1270, N1268);
nor NOR3 (N1271, N1263, N796, N939);
buf BUF1 (N1272, N1271);
or OR4 (N1273, N1272, N82, N1250, N201);
and AND2 (N1274, N981, N873);
or OR4 (N1275, N1273, N867, N184, N356);
nor NOR2 (N1276, N1260, N403);
and AND4 (N1277, N1270, N812, N986, N323);
and AND2 (N1278, N1266, N734);
not NOT1 (N1279, N1242);
nand NAND2 (N1280, N1267, N206);
nand NAND2 (N1281, N1248, N1043);
xor XOR2 (N1282, N1281, N1192);
buf BUF1 (N1283, N1261);
not NOT1 (N1284, N1276);
nor NOR4 (N1285, N1279, N1145, N690, N1268);
xor XOR2 (N1286, N1274, N1203);
nand NAND2 (N1287, N1277, N229);
not NOT1 (N1288, N1275);
xor XOR2 (N1289, N1269, N1194);
and AND3 (N1290, N1278, N1022, N1028);
buf BUF1 (N1291, N1288);
not NOT1 (N1292, N1282);
xor XOR2 (N1293, N1289, N251);
nand NAND2 (N1294, N1285, N451);
nor NOR4 (N1295, N1293, N715, N653, N261);
or OR4 (N1296, N1294, N192, N899, N59);
nand NAND4 (N1297, N1287, N75, N459, N87);
buf BUF1 (N1298, N1280);
and AND2 (N1299, N1298, N1050);
buf BUF1 (N1300, N1297);
or OR2 (N1301, N1284, N267);
or OR2 (N1302, N1296, N677);
not NOT1 (N1303, N1301);
and AND2 (N1304, N1290, N278);
xor XOR2 (N1305, N1299, N889);
xor XOR2 (N1306, N1292, N754);
xor XOR2 (N1307, N1291, N693);
buf BUF1 (N1308, N1305);
not NOT1 (N1309, N1303);
nor NOR3 (N1310, N1302, N651, N1001);
and AND2 (N1311, N1310, N761);
not NOT1 (N1312, N1309);
and AND2 (N1313, N1283, N86);
xor XOR2 (N1314, N1307, N759);
buf BUF1 (N1315, N1312);
buf BUF1 (N1316, N1300);
xor XOR2 (N1317, N1315, N481);
nor NOR4 (N1318, N1304, N590, N222, N575);
or OR4 (N1319, N1306, N1162, N733, N1188);
nand NAND2 (N1320, N1319, N857);
nand NAND4 (N1321, N1313, N153, N98, N470);
and AND2 (N1322, N1317, N1171);
nand NAND4 (N1323, N1311, N959, N87, N437);
not NOT1 (N1324, N1322);
and AND4 (N1325, N1308, N980, N665, N1152);
not NOT1 (N1326, N1318);
buf BUF1 (N1327, N1320);
nor NOR4 (N1328, N1323, N254, N133, N1123);
nor NOR2 (N1329, N1324, N743);
nand NAND2 (N1330, N1326, N571);
not NOT1 (N1331, N1321);
buf BUF1 (N1332, N1314);
xor XOR2 (N1333, N1295, N1053);
not NOT1 (N1334, N1316);
not NOT1 (N1335, N1327);
or OR3 (N1336, N1334, N1172, N321);
buf BUF1 (N1337, N1329);
not NOT1 (N1338, N1332);
nand NAND2 (N1339, N1337, N420);
nand NAND3 (N1340, N1336, N541, N826);
not NOT1 (N1341, N1335);
nor NOR4 (N1342, N1325, N1069, N110, N805);
or OR2 (N1343, N1342, N295);
and AND2 (N1344, N1331, N773);
or OR2 (N1345, N1340, N1044);
xor XOR2 (N1346, N1286, N184);
not NOT1 (N1347, N1344);
buf BUF1 (N1348, N1343);
not NOT1 (N1349, N1338);
nand NAND3 (N1350, N1347, N1129, N1030);
and AND3 (N1351, N1349, N941, N1292);
nand NAND2 (N1352, N1348, N1069);
xor XOR2 (N1353, N1351, N398);
nand NAND4 (N1354, N1345, N261, N1203, N993);
not NOT1 (N1355, N1346);
or OR2 (N1356, N1353, N54);
and AND3 (N1357, N1356, N1290, N255);
and AND3 (N1358, N1339, N194, N684);
and AND4 (N1359, N1330, N860, N1031, N512);
and AND4 (N1360, N1354, N336, N60, N423);
xor XOR2 (N1361, N1360, N723);
buf BUF1 (N1362, N1352);
nand NAND3 (N1363, N1350, N1174, N1028);
nand NAND3 (N1364, N1355, N349, N402);
not NOT1 (N1365, N1333);
nand NAND3 (N1366, N1328, N504, N682);
buf BUF1 (N1367, N1361);
or OR3 (N1368, N1366, N381, N550);
nor NOR3 (N1369, N1363, N240, N955);
not NOT1 (N1370, N1359);
buf BUF1 (N1371, N1370);
and AND4 (N1372, N1364, N586, N1187, N305);
or OR2 (N1373, N1365, N1314);
or OR3 (N1374, N1341, N1152, N576);
nor NOR3 (N1375, N1371, N253, N1211);
buf BUF1 (N1376, N1369);
not NOT1 (N1377, N1373);
nand NAND3 (N1378, N1358, N152, N667);
nor NOR2 (N1379, N1368, N159);
nand NAND4 (N1380, N1362, N952, N286, N267);
and AND2 (N1381, N1378, N82);
nor NOR2 (N1382, N1367, N287);
and AND2 (N1383, N1377, N638);
nand NAND3 (N1384, N1376, N1280, N470);
buf BUF1 (N1385, N1383);
nand NAND4 (N1386, N1385, N262, N1291, N1334);
nor NOR2 (N1387, N1357, N335);
buf BUF1 (N1388, N1375);
nand NAND2 (N1389, N1388, N1153);
not NOT1 (N1390, N1379);
and AND4 (N1391, N1390, N626, N999, N1356);
xor XOR2 (N1392, N1381, N781);
nor NOR3 (N1393, N1372, N241, N544);
buf BUF1 (N1394, N1380);
buf BUF1 (N1395, N1389);
not NOT1 (N1396, N1374);
or OR4 (N1397, N1396, N952, N850, N1173);
nor NOR2 (N1398, N1386, N204);
nand NAND4 (N1399, N1391, N947, N1228, N491);
xor XOR2 (N1400, N1397, N387);
and AND2 (N1401, N1387, N547);
or OR4 (N1402, N1393, N808, N947, N527);
or OR3 (N1403, N1399, N225, N1040);
and AND3 (N1404, N1384, N415, N1077);
not NOT1 (N1405, N1392);
and AND3 (N1406, N1398, N149, N441);
xor XOR2 (N1407, N1400, N1399);
not NOT1 (N1408, N1405);
nand NAND4 (N1409, N1402, N1381, N580, N1117);
or OR2 (N1410, N1409, N155);
or OR4 (N1411, N1407, N229, N600, N1303);
nor NOR2 (N1412, N1395, N1164);
not NOT1 (N1413, N1382);
xor XOR2 (N1414, N1410, N955);
and AND2 (N1415, N1411, N1025);
nor NOR4 (N1416, N1406, N1117, N888, N570);
or OR2 (N1417, N1403, N658);
xor XOR2 (N1418, N1415, N458);
nand NAND4 (N1419, N1404, N271, N1251, N440);
nor NOR2 (N1420, N1414, N794);
nor NOR2 (N1421, N1408, N180);
nor NOR2 (N1422, N1419, N1081);
or OR4 (N1423, N1394, N110, N590, N526);
buf BUF1 (N1424, N1423);
not NOT1 (N1425, N1401);
and AND2 (N1426, N1418, N1219);
and AND2 (N1427, N1420, N1006);
nand NAND2 (N1428, N1425, N103);
not NOT1 (N1429, N1424);
and AND4 (N1430, N1422, N1065, N793, N414);
nand NAND2 (N1431, N1416, N1200);
nor NOR2 (N1432, N1412, N430);
not NOT1 (N1433, N1417);
xor XOR2 (N1434, N1431, N1093);
not NOT1 (N1435, N1428);
xor XOR2 (N1436, N1435, N93);
xor XOR2 (N1437, N1413, N682);
buf BUF1 (N1438, N1437);
or OR3 (N1439, N1421, N330, N633);
xor XOR2 (N1440, N1436, N1273);
xor XOR2 (N1441, N1440, N1100);
buf BUF1 (N1442, N1426);
nand NAND4 (N1443, N1434, N943, N406, N1247);
or OR3 (N1444, N1427, N454, N771);
nand NAND2 (N1445, N1433, N1177);
buf BUF1 (N1446, N1443);
not NOT1 (N1447, N1444);
not NOT1 (N1448, N1432);
or OR4 (N1449, N1438, N1035, N1025, N502);
nor NOR4 (N1450, N1442, N1349, N505, N1052);
buf BUF1 (N1451, N1430);
xor XOR2 (N1452, N1445, N628);
xor XOR2 (N1453, N1446, N204);
nand NAND2 (N1454, N1439, N1317);
buf BUF1 (N1455, N1448);
nand NAND4 (N1456, N1451, N870, N1190, N880);
not NOT1 (N1457, N1441);
xor XOR2 (N1458, N1429, N1101);
nor NOR2 (N1459, N1454, N606);
xor XOR2 (N1460, N1450, N1396);
xor XOR2 (N1461, N1457, N1014);
nor NOR3 (N1462, N1458, N150, N1319);
not NOT1 (N1463, N1452);
and AND4 (N1464, N1456, N386, N866, N991);
not NOT1 (N1465, N1460);
xor XOR2 (N1466, N1464, N358);
buf BUF1 (N1467, N1459);
nor NOR4 (N1468, N1455, N782, N871, N589);
nand NAND3 (N1469, N1461, N1468, N25);
not NOT1 (N1470, N1033);
xor XOR2 (N1471, N1466, N542);
buf BUF1 (N1472, N1469);
xor XOR2 (N1473, N1449, N74);
xor XOR2 (N1474, N1465, N709);
and AND4 (N1475, N1467, N610, N600, N788);
xor XOR2 (N1476, N1473, N967);
buf BUF1 (N1477, N1470);
buf BUF1 (N1478, N1462);
or OR3 (N1479, N1474, N10, N757);
nand NAND4 (N1480, N1476, N1402, N335, N1316);
nand NAND4 (N1481, N1472, N717, N678, N668);
nand NAND4 (N1482, N1481, N1464, N518, N129);
not NOT1 (N1483, N1479);
xor XOR2 (N1484, N1483, N658);
nand NAND4 (N1485, N1453, N745, N1439, N490);
buf BUF1 (N1486, N1478);
xor XOR2 (N1487, N1484, N1136);
not NOT1 (N1488, N1485);
nand NAND4 (N1489, N1477, N292, N266, N493);
xor XOR2 (N1490, N1480, N997);
not NOT1 (N1491, N1490);
buf BUF1 (N1492, N1482);
and AND3 (N1493, N1491, N791, N1366);
and AND3 (N1494, N1487, N338, N1321);
not NOT1 (N1495, N1471);
xor XOR2 (N1496, N1486, N437);
not NOT1 (N1497, N1489);
xor XOR2 (N1498, N1493, N410);
nor NOR3 (N1499, N1463, N531, N728);
buf BUF1 (N1500, N1475);
xor XOR2 (N1501, N1499, N703);
buf BUF1 (N1502, N1488);
buf BUF1 (N1503, N1498);
not NOT1 (N1504, N1496);
buf BUF1 (N1505, N1502);
or OR4 (N1506, N1492, N241, N1033, N1035);
or OR4 (N1507, N1506, N350, N1339, N219);
not NOT1 (N1508, N1497);
buf BUF1 (N1509, N1501);
not NOT1 (N1510, N1500);
nor NOR4 (N1511, N1510, N161, N661, N233);
buf BUF1 (N1512, N1511);
xor XOR2 (N1513, N1507, N856);
nand NAND2 (N1514, N1504, N293);
not NOT1 (N1515, N1494);
and AND3 (N1516, N1515, N116, N1394);
nor NOR2 (N1517, N1508, N1394);
and AND3 (N1518, N1512, N279, N1412);
buf BUF1 (N1519, N1514);
and AND2 (N1520, N1517, N112);
nor NOR2 (N1521, N1495, N294);
and AND3 (N1522, N1521, N378, N875);
xor XOR2 (N1523, N1520, N391);
not NOT1 (N1524, N1519);
not NOT1 (N1525, N1524);
buf BUF1 (N1526, N1505);
nand NAND3 (N1527, N1526, N1198, N551);
nor NOR3 (N1528, N1516, N1020, N1167);
buf BUF1 (N1529, N1447);
buf BUF1 (N1530, N1522);
nand NAND3 (N1531, N1527, N5, N1430);
or OR4 (N1532, N1528, N957, N1422, N417);
nor NOR3 (N1533, N1532, N1090, N187);
nor NOR4 (N1534, N1530, N519, N1427, N177);
or OR2 (N1535, N1523, N541);
nor NOR2 (N1536, N1518, N880);
buf BUF1 (N1537, N1536);
or OR4 (N1538, N1534, N310, N1049, N575);
xor XOR2 (N1539, N1513, N564);
nor NOR3 (N1540, N1538, N485, N859);
nor NOR3 (N1541, N1525, N143, N935);
not NOT1 (N1542, N1540);
buf BUF1 (N1543, N1503);
or OR3 (N1544, N1542, N362, N243);
xor XOR2 (N1545, N1537, N901);
not NOT1 (N1546, N1535);
buf BUF1 (N1547, N1539);
nand NAND4 (N1548, N1533, N714, N913, N1047);
buf BUF1 (N1549, N1529);
buf BUF1 (N1550, N1543);
or OR4 (N1551, N1509, N595, N888, N811);
xor XOR2 (N1552, N1544, N300);
buf BUF1 (N1553, N1547);
xor XOR2 (N1554, N1546, N660);
and AND4 (N1555, N1551, N691, N907, N1000);
nand NAND4 (N1556, N1549, N411, N4, N886);
nand NAND3 (N1557, N1554, N1364, N618);
buf BUF1 (N1558, N1555);
nor NOR4 (N1559, N1548, N1085, N1364, N1399);
or OR3 (N1560, N1559, N161, N660);
not NOT1 (N1561, N1560);
or OR2 (N1562, N1531, N621);
or OR3 (N1563, N1541, N1084, N200);
nand NAND3 (N1564, N1552, N135, N300);
xor XOR2 (N1565, N1550, N1466);
buf BUF1 (N1566, N1563);
nand NAND3 (N1567, N1566, N103, N1120);
not NOT1 (N1568, N1553);
buf BUF1 (N1569, N1557);
buf BUF1 (N1570, N1561);
nand NAND4 (N1571, N1565, N1035, N126, N1564);
not NOT1 (N1572, N870);
nor NOR2 (N1573, N1556, N229);
not NOT1 (N1574, N1570);
xor XOR2 (N1575, N1545, N44);
buf BUF1 (N1576, N1571);
nand NAND3 (N1577, N1558, N211, N1158);
nor NOR2 (N1578, N1569, N1251);
xor XOR2 (N1579, N1567, N292);
nor NOR3 (N1580, N1576, N1096, N138);
or OR2 (N1581, N1574, N1111);
not NOT1 (N1582, N1572);
and AND4 (N1583, N1568, N1411, N1329, N777);
or OR2 (N1584, N1573, N1327);
and AND4 (N1585, N1584, N1417, N1199, N489);
xor XOR2 (N1586, N1582, N1264);
buf BUF1 (N1587, N1586);
nand NAND3 (N1588, N1579, N188, N1467);
nor NOR2 (N1589, N1575, N747);
nand NAND2 (N1590, N1583, N1433);
xor XOR2 (N1591, N1589, N1475);
and AND3 (N1592, N1591, N814, N265);
and AND3 (N1593, N1585, N1410, N187);
buf BUF1 (N1594, N1590);
buf BUF1 (N1595, N1592);
not NOT1 (N1596, N1588);
xor XOR2 (N1597, N1581, N1139);
xor XOR2 (N1598, N1597, N1597);
or OR2 (N1599, N1595, N924);
xor XOR2 (N1600, N1594, N1182);
nor NOR3 (N1601, N1598, N1005, N482);
or OR2 (N1602, N1596, N640);
and AND4 (N1603, N1602, N270, N1506, N1028);
or OR4 (N1604, N1562, N839, N1415, N549);
not NOT1 (N1605, N1603);
nand NAND2 (N1606, N1604, N203);
nor NOR4 (N1607, N1605, N917, N119, N536);
xor XOR2 (N1608, N1599, N9);
xor XOR2 (N1609, N1578, N70);
xor XOR2 (N1610, N1609, N913);
xor XOR2 (N1611, N1607, N1420);
not NOT1 (N1612, N1593);
and AND4 (N1613, N1610, N482, N1037, N1116);
buf BUF1 (N1614, N1600);
or OR4 (N1615, N1601, N1056, N257, N1056);
nand NAND3 (N1616, N1614, N9, N632);
nand NAND2 (N1617, N1611, N1584);
and AND3 (N1618, N1577, N351, N1234);
not NOT1 (N1619, N1616);
or OR3 (N1620, N1580, N956, N178);
nor NOR3 (N1621, N1606, N1521, N1213);
nor NOR2 (N1622, N1618, N1575);
buf BUF1 (N1623, N1612);
or OR3 (N1624, N1621, N48, N1431);
or OR3 (N1625, N1613, N1110, N1228);
xor XOR2 (N1626, N1622, N1413);
nor NOR2 (N1627, N1587, N1384);
and AND2 (N1628, N1620, N323);
not NOT1 (N1629, N1615);
xor XOR2 (N1630, N1626, N282);
not NOT1 (N1631, N1630);
xor XOR2 (N1632, N1619, N1042);
and AND3 (N1633, N1631, N295, N1479);
or OR4 (N1634, N1608, N885, N1102, N881);
buf BUF1 (N1635, N1634);
buf BUF1 (N1636, N1627);
nor NOR2 (N1637, N1625, N71);
and AND2 (N1638, N1636, N1308);
xor XOR2 (N1639, N1624, N783);
nand NAND2 (N1640, N1628, N573);
and AND2 (N1641, N1639, N626);
nor NOR2 (N1642, N1623, N998);
or OR4 (N1643, N1641, N432, N952, N573);
nand NAND2 (N1644, N1635, N910);
and AND2 (N1645, N1640, N1582);
not NOT1 (N1646, N1644);
or OR4 (N1647, N1617, N1118, N843, N515);
buf BUF1 (N1648, N1645);
and AND3 (N1649, N1642, N550, N436);
and AND3 (N1650, N1648, N1423, N255);
and AND3 (N1651, N1646, N1566, N691);
or OR2 (N1652, N1637, N1109);
nand NAND4 (N1653, N1652, N817, N550, N57);
nand NAND4 (N1654, N1650, N1271, N1526, N737);
nand NAND4 (N1655, N1632, N1425, N1451, N930);
or OR2 (N1656, N1643, N269);
nand NAND2 (N1657, N1653, N676);
and AND3 (N1658, N1655, N259, N937);
nand NAND4 (N1659, N1629, N23, N42, N387);
not NOT1 (N1660, N1659);
buf BUF1 (N1661, N1647);
or OR2 (N1662, N1657, N1504);
nand NAND2 (N1663, N1658, N266);
and AND4 (N1664, N1638, N407, N1583, N1435);
nand NAND4 (N1665, N1633, N1411, N574, N604);
nor NOR4 (N1666, N1660, N680, N1550, N719);
buf BUF1 (N1667, N1664);
and AND4 (N1668, N1656, N218, N1227, N1340);
nand NAND3 (N1669, N1668, N1620, N279);
and AND3 (N1670, N1667, N916, N1224);
nand NAND4 (N1671, N1651, N600, N1338, N273);
or OR2 (N1672, N1670, N603);
or OR4 (N1673, N1661, N717, N449, N297);
nand NAND4 (N1674, N1649, N354, N1241, N827);
xor XOR2 (N1675, N1663, N883);
or OR2 (N1676, N1669, N624);
nand NAND2 (N1677, N1665, N730);
buf BUF1 (N1678, N1672);
xor XOR2 (N1679, N1666, N1206);
and AND2 (N1680, N1662, N197);
xor XOR2 (N1681, N1654, N635);
nor NOR4 (N1682, N1681, N771, N323, N386);
or OR3 (N1683, N1671, N117, N626);
not NOT1 (N1684, N1680);
nand NAND4 (N1685, N1679, N1391, N353, N202);
or OR3 (N1686, N1675, N145, N429);
xor XOR2 (N1687, N1683, N530);
buf BUF1 (N1688, N1676);
or OR2 (N1689, N1686, N1290);
buf BUF1 (N1690, N1674);
buf BUF1 (N1691, N1690);
xor XOR2 (N1692, N1687, N1397);
buf BUF1 (N1693, N1689);
nor NOR4 (N1694, N1685, N804, N1531, N140);
xor XOR2 (N1695, N1677, N33);
not NOT1 (N1696, N1695);
xor XOR2 (N1697, N1688, N1004);
xor XOR2 (N1698, N1692, N190);
not NOT1 (N1699, N1682);
nand NAND4 (N1700, N1699, N1185, N667, N667);
xor XOR2 (N1701, N1691, N4);
and AND4 (N1702, N1697, N549, N386, N1605);
and AND3 (N1703, N1701, N1617, N843);
buf BUF1 (N1704, N1703);
and AND2 (N1705, N1694, N502);
xor XOR2 (N1706, N1704, N308);
nand NAND4 (N1707, N1698, N1544, N1610, N1210);
buf BUF1 (N1708, N1684);
not NOT1 (N1709, N1700);
nor NOR4 (N1710, N1709, N1405, N234, N974);
or OR4 (N1711, N1702, N489, N847, N499);
buf BUF1 (N1712, N1708);
not NOT1 (N1713, N1706);
and AND4 (N1714, N1693, N1635, N412, N613);
and AND4 (N1715, N1678, N931, N1322, N1578);
buf BUF1 (N1716, N1696);
xor XOR2 (N1717, N1714, N1231);
buf BUF1 (N1718, N1711);
or OR2 (N1719, N1707, N1466);
nand NAND2 (N1720, N1705, N660);
and AND4 (N1721, N1673, N636, N1388, N75);
and AND4 (N1722, N1710, N1210, N1423, N345);
nand NAND3 (N1723, N1716, N1521, N184);
and AND3 (N1724, N1718, N1233, N326);
or OR3 (N1725, N1717, N1561, N1719);
and AND2 (N1726, N1486, N1651);
buf BUF1 (N1727, N1713);
not NOT1 (N1728, N1726);
xor XOR2 (N1729, N1720, N109);
xor XOR2 (N1730, N1721, N1496);
xor XOR2 (N1731, N1715, N1716);
not NOT1 (N1732, N1723);
or OR2 (N1733, N1727, N1458);
not NOT1 (N1734, N1733);
nor NOR2 (N1735, N1722, N314);
nand NAND4 (N1736, N1734, N1015, N470, N1687);
xor XOR2 (N1737, N1732, N116);
not NOT1 (N1738, N1725);
and AND3 (N1739, N1730, N108, N901);
or OR3 (N1740, N1736, N930, N1104);
nand NAND2 (N1741, N1739, N1678);
or OR4 (N1742, N1740, N1523, N378, N270);
and AND4 (N1743, N1735, N1364, N1584, N814);
or OR3 (N1744, N1728, N19, N1099);
not NOT1 (N1745, N1738);
xor XOR2 (N1746, N1729, N962);
nor NOR2 (N1747, N1731, N1086);
not NOT1 (N1748, N1712);
not NOT1 (N1749, N1724);
buf BUF1 (N1750, N1747);
not NOT1 (N1751, N1744);
buf BUF1 (N1752, N1737);
nand NAND4 (N1753, N1742, N850, N643, N1016);
nand NAND2 (N1754, N1751, N821);
xor XOR2 (N1755, N1745, N774);
buf BUF1 (N1756, N1746);
not NOT1 (N1757, N1741);
and AND2 (N1758, N1750, N392);
or OR4 (N1759, N1753, N580, N1232, N625);
and AND3 (N1760, N1758, N282, N1638);
xor XOR2 (N1761, N1749, N221);
buf BUF1 (N1762, N1761);
nor NOR3 (N1763, N1752, N588, N1362);
or OR4 (N1764, N1755, N728, N494, N55);
xor XOR2 (N1765, N1764, N1689);
and AND2 (N1766, N1756, N743);
nor NOR4 (N1767, N1757, N337, N582, N220);
nand NAND2 (N1768, N1765, N431);
nor NOR4 (N1769, N1762, N1585, N1628, N922);
nor NOR3 (N1770, N1759, N1466, N503);
nor NOR3 (N1771, N1763, N1466, N753);
nand NAND4 (N1772, N1770, N1116, N1073, N1003);
xor XOR2 (N1773, N1754, N1771);
buf BUF1 (N1774, N993);
nand NAND4 (N1775, N1774, N683, N1047, N609);
and AND2 (N1776, N1748, N777);
nand NAND4 (N1777, N1769, N564, N788, N727);
not NOT1 (N1778, N1743);
or OR4 (N1779, N1760, N1523, N1516, N449);
or OR4 (N1780, N1766, N1159, N1578, N809);
not NOT1 (N1781, N1773);
xor XOR2 (N1782, N1767, N1325);
or OR3 (N1783, N1777, N536, N954);
and AND3 (N1784, N1768, N1305, N1274);
not NOT1 (N1785, N1776);
or OR2 (N1786, N1784, N1035);
nor NOR3 (N1787, N1778, N1550, N535);
not NOT1 (N1788, N1781);
or OR3 (N1789, N1787, N1010, N749);
and AND4 (N1790, N1779, N515, N1520, N302);
nand NAND4 (N1791, N1790, N1441, N305, N194);
buf BUF1 (N1792, N1783);
nand NAND3 (N1793, N1792, N1001, N806);
or OR4 (N1794, N1782, N1611, N1121, N632);
nand NAND4 (N1795, N1788, N1073, N596, N287);
or OR3 (N1796, N1795, N1139, N1548);
nor NOR3 (N1797, N1780, N1235, N1792);
and AND2 (N1798, N1775, N865);
and AND2 (N1799, N1796, N276);
nand NAND2 (N1800, N1786, N538);
nand NAND4 (N1801, N1799, N1615, N1029, N1679);
xor XOR2 (N1802, N1797, N457);
not NOT1 (N1803, N1800);
and AND4 (N1804, N1798, N1559, N784, N1491);
nand NAND2 (N1805, N1794, N1611);
not NOT1 (N1806, N1804);
nand NAND2 (N1807, N1772, N1516);
and AND4 (N1808, N1785, N1399, N853, N1312);
or OR3 (N1809, N1793, N1722, N38);
buf BUF1 (N1810, N1808);
buf BUF1 (N1811, N1791);
nor NOR3 (N1812, N1802, N1585, N1172);
and AND4 (N1813, N1810, N194, N1348, N826);
xor XOR2 (N1814, N1789, N1422);
not NOT1 (N1815, N1807);
or OR3 (N1816, N1805, N1802, N1040);
not NOT1 (N1817, N1814);
not NOT1 (N1818, N1813);
or OR2 (N1819, N1809, N346);
or OR3 (N1820, N1815, N245, N895);
xor XOR2 (N1821, N1803, N250);
nand NAND2 (N1822, N1801, N691);
nand NAND2 (N1823, N1821, N1087);
nor NOR4 (N1824, N1806, N1263, N1354, N560);
not NOT1 (N1825, N1811);
nand NAND4 (N1826, N1822, N680, N1673, N1298);
nor NOR4 (N1827, N1826, N468, N536, N917);
nand NAND3 (N1828, N1827, N1176, N296);
or OR2 (N1829, N1824, N283);
or OR4 (N1830, N1812, N1793, N139, N306);
and AND3 (N1831, N1818, N1669, N1606);
xor XOR2 (N1832, N1820, N693);
not NOT1 (N1833, N1828);
and AND4 (N1834, N1831, N1628, N717, N967);
or OR2 (N1835, N1829, N713);
nand NAND2 (N1836, N1817, N1758);
or OR4 (N1837, N1816, N670, N404, N1734);
xor XOR2 (N1838, N1834, N139);
xor XOR2 (N1839, N1830, N772);
nor NOR2 (N1840, N1825, N1255);
or OR2 (N1841, N1832, N1140);
not NOT1 (N1842, N1838);
nand NAND3 (N1843, N1823, N39, N682);
not NOT1 (N1844, N1835);
buf BUF1 (N1845, N1840);
not NOT1 (N1846, N1842);
buf BUF1 (N1847, N1841);
buf BUF1 (N1848, N1843);
nand NAND2 (N1849, N1848, N50);
not NOT1 (N1850, N1847);
buf BUF1 (N1851, N1844);
or OR3 (N1852, N1851, N750, N663);
not NOT1 (N1853, N1839);
nand NAND4 (N1854, N1845, N967, N1030, N1557);
buf BUF1 (N1855, N1833);
and AND3 (N1856, N1850, N1416, N383);
nor NOR2 (N1857, N1846, N357);
xor XOR2 (N1858, N1857, N1784);
or OR3 (N1859, N1855, N213, N1358);
xor XOR2 (N1860, N1819, N211);
and AND3 (N1861, N1858, N893, N1547);
xor XOR2 (N1862, N1854, N1270);
nand NAND2 (N1863, N1860, N875);
nand NAND4 (N1864, N1849, N1646, N783, N224);
nand NAND3 (N1865, N1836, N1299, N900);
buf BUF1 (N1866, N1862);
or OR4 (N1867, N1866, N998, N1386, N263);
and AND4 (N1868, N1853, N1553, N622, N1667);
or OR2 (N1869, N1856, N1582);
xor XOR2 (N1870, N1868, N40);
and AND4 (N1871, N1865, N875, N1329, N686);
and AND4 (N1872, N1863, N1494, N283, N712);
xor XOR2 (N1873, N1837, N1543);
nand NAND2 (N1874, N1859, N746);
nor NOR4 (N1875, N1873, N841, N472, N174);
and AND3 (N1876, N1870, N572, N1776);
not NOT1 (N1877, N1871);
and AND4 (N1878, N1877, N1536, N11, N416);
and AND3 (N1879, N1878, N180, N187);
not NOT1 (N1880, N1864);
and AND3 (N1881, N1852, N408, N1100);
buf BUF1 (N1882, N1867);
nand NAND3 (N1883, N1861, N1392, N900);
not NOT1 (N1884, N1883);
not NOT1 (N1885, N1872);
buf BUF1 (N1886, N1884);
xor XOR2 (N1887, N1880, N1638);
nor NOR2 (N1888, N1876, N1884);
not NOT1 (N1889, N1882);
buf BUF1 (N1890, N1881);
buf BUF1 (N1891, N1869);
not NOT1 (N1892, N1891);
buf BUF1 (N1893, N1887);
xor XOR2 (N1894, N1888, N1071);
xor XOR2 (N1895, N1894, N1027);
or OR2 (N1896, N1889, N1110);
xor XOR2 (N1897, N1885, N1654);
not NOT1 (N1898, N1893);
not NOT1 (N1899, N1895);
not NOT1 (N1900, N1892);
xor XOR2 (N1901, N1896, N531);
xor XOR2 (N1902, N1900, N1235);
buf BUF1 (N1903, N1886);
nand NAND2 (N1904, N1890, N178);
nor NOR4 (N1905, N1902, N1715, N675, N835);
nand NAND2 (N1906, N1901, N777);
and AND4 (N1907, N1899, N274, N1349, N508);
xor XOR2 (N1908, N1879, N1401);
and AND2 (N1909, N1905, N1882);
and AND2 (N1910, N1874, N752);
or OR3 (N1911, N1906, N555, N46);
xor XOR2 (N1912, N1907, N672);
not NOT1 (N1913, N1912);
nand NAND2 (N1914, N1903, N153);
xor XOR2 (N1915, N1913, N1335);
and AND2 (N1916, N1904, N1890);
not NOT1 (N1917, N1914);
buf BUF1 (N1918, N1910);
nor NOR4 (N1919, N1875, N1547, N97, N827);
buf BUF1 (N1920, N1898);
not NOT1 (N1921, N1919);
or OR4 (N1922, N1916, N1820, N1512, N346);
not NOT1 (N1923, N1909);
not NOT1 (N1924, N1897);
buf BUF1 (N1925, N1920);
nand NAND4 (N1926, N1925, N399, N474, N1196);
and AND4 (N1927, N1908, N414, N892, N1413);
xor XOR2 (N1928, N1926, N1613);
buf BUF1 (N1929, N1911);
buf BUF1 (N1930, N1924);
nand NAND4 (N1931, N1917, N1685, N1068, N1888);
nand NAND4 (N1932, N1928, N729, N349, N1139);
xor XOR2 (N1933, N1932, N466);
buf BUF1 (N1934, N1931);
not NOT1 (N1935, N1921);
or OR2 (N1936, N1929, N304);
xor XOR2 (N1937, N1935, N1491);
or OR3 (N1938, N1937, N1048, N1402);
not NOT1 (N1939, N1922);
xor XOR2 (N1940, N1927, N1801);
xor XOR2 (N1941, N1915, N1913);
nand NAND4 (N1942, N1938, N369, N1533, N1691);
buf BUF1 (N1943, N1930);
xor XOR2 (N1944, N1939, N1892);
not NOT1 (N1945, N1934);
not NOT1 (N1946, N1936);
and AND2 (N1947, N1943, N1591);
and AND4 (N1948, N1940, N310, N235, N829);
nor NOR4 (N1949, N1945, N395, N227, N763);
or OR4 (N1950, N1949, N1531, N51, N1614);
nor NOR4 (N1951, N1933, N1500, N1528, N1816);
not NOT1 (N1952, N1942);
and AND3 (N1953, N1923, N110, N240);
nor NOR3 (N1954, N1918, N39, N504);
buf BUF1 (N1955, N1941);
buf BUF1 (N1956, N1947);
or OR3 (N1957, N1944, N1632, N1338);
buf BUF1 (N1958, N1956);
or OR4 (N1959, N1950, N393, N654, N1070);
xor XOR2 (N1960, N1946, N1213);
buf BUF1 (N1961, N1948);
nand NAND3 (N1962, N1955, N1700, N1633);
and AND3 (N1963, N1960, N1182, N90);
not NOT1 (N1964, N1951);
not NOT1 (N1965, N1957);
buf BUF1 (N1966, N1959);
and AND4 (N1967, N1962, N783, N1137, N603);
and AND3 (N1968, N1961, N1944, N338);
and AND4 (N1969, N1963, N1820, N90, N1263);
not NOT1 (N1970, N1966);
buf BUF1 (N1971, N1965);
nand NAND4 (N1972, N1952, N1601, N1334, N982);
buf BUF1 (N1973, N1953);
nand NAND3 (N1974, N1970, N703, N826);
and AND3 (N1975, N1973, N45, N632);
nor NOR3 (N1976, N1954, N1133, N765);
xor XOR2 (N1977, N1975, N504);
nand NAND2 (N1978, N1972, N1347);
or OR4 (N1979, N1974, N1542, N246, N1347);
xor XOR2 (N1980, N1964, N1585);
xor XOR2 (N1981, N1977, N1039);
or OR2 (N1982, N1978, N1938);
buf BUF1 (N1983, N1982);
xor XOR2 (N1984, N1979, N1814);
and AND3 (N1985, N1976, N1304, N1395);
xor XOR2 (N1986, N1967, N1930);
or OR3 (N1987, N1969, N1265, N1003);
buf BUF1 (N1988, N1971);
nand NAND3 (N1989, N1983, N829, N1627);
buf BUF1 (N1990, N1968);
nand NAND4 (N1991, N1984, N1783, N864, N1990);
nand NAND2 (N1992, N525, N301);
xor XOR2 (N1993, N1991, N1338);
buf BUF1 (N1994, N1981);
not NOT1 (N1995, N1993);
and AND3 (N1996, N1958, N725, N1073);
nor NOR3 (N1997, N1995, N1662, N1933);
and AND3 (N1998, N1992, N1432, N257);
nand NAND4 (N1999, N1987, N1744, N474, N1190);
buf BUF1 (N2000, N1980);
nand NAND4 (N2001, N1997, N1448, N1041, N94);
not NOT1 (N2002, N1989);
xor XOR2 (N2003, N2001, N1495);
xor XOR2 (N2004, N1994, N961);
xor XOR2 (N2005, N1985, N1199);
nand NAND2 (N2006, N1998, N243);
nand NAND4 (N2007, N2000, N982, N417, N1441);
nor NOR4 (N2008, N1986, N1536, N351, N1859);
not NOT1 (N2009, N1999);
nor NOR3 (N2010, N1996, N1454, N425);
nand NAND2 (N2011, N2006, N1632);
nand NAND3 (N2012, N2010, N781, N780);
and AND4 (N2013, N2008, N796, N725, N1574);
xor XOR2 (N2014, N2011, N347);
buf BUF1 (N2015, N2005);
or OR4 (N2016, N2009, N931, N1229, N1465);
and AND4 (N2017, N2003, N521, N1134, N1431);
or OR3 (N2018, N2013, N29, N381);
and AND2 (N2019, N1988, N1002);
nand NAND2 (N2020, N2004, N93);
endmodule