// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24;

output N1017,N1014,N1022,N1009,N1010,N1019,N1018,N1020,N1016,N1024;

xor XOR2 (N25, N8, N7);
xor XOR2 (N26, N1, N1);
nor NOR2 (N27, N3, N1);
or OR4 (N28, N2, N22, N18, N19);
and AND3 (N29, N20, N25, N16);
and AND4 (N30, N11, N29, N7, N9);
not NOT1 (N31, N5);
xor XOR2 (N32, N22, N26);
nand NAND4 (N33, N32, N29, N17, N6);
nand NAND2 (N34, N11, N6);
nor NOR2 (N35, N32, N9);
nor NOR3 (N36, N12, N20, N2);
not NOT1 (N37, N15);
and AND4 (N38, N18, N8, N6, N7);
nand NAND2 (N39, N37, N12);
not NOT1 (N40, N28);
not NOT1 (N41, N35);
nand NAND2 (N42, N33, N15);
and AND4 (N43, N34, N16, N16, N11);
not NOT1 (N44, N39);
xor XOR2 (N45, N30, N16);
or OR3 (N46, N36, N24, N5);
and AND2 (N47, N43, N28);
or OR4 (N48, N31, N4, N12, N6);
not NOT1 (N49, N46);
xor XOR2 (N50, N27, N45);
and AND2 (N51, N32, N47);
and AND3 (N52, N4, N50, N43);
buf BUF1 (N53, N1);
and AND3 (N54, N53, N40, N49);
xor XOR2 (N55, N38, N52);
nand NAND2 (N56, N35, N35);
and AND3 (N57, N9, N21, N52);
or OR4 (N58, N38, N54, N50, N28);
nor NOR4 (N59, N31, N33, N48, N7);
nor NOR3 (N60, N21, N29, N23);
buf BUF1 (N61, N44);
xor XOR2 (N62, N59, N19);
nor NOR4 (N63, N41, N61, N23, N5);
nand NAND4 (N64, N39, N20, N8, N13);
and AND2 (N65, N60, N13);
buf BUF1 (N66, N62);
nand NAND4 (N67, N64, N34, N39, N3);
not NOT1 (N68, N55);
nor NOR2 (N69, N65, N50);
and AND3 (N70, N57, N50, N11);
nand NAND2 (N71, N66, N48);
not NOT1 (N72, N51);
or OR4 (N73, N72, N42, N19, N8);
xor XOR2 (N74, N13, N40);
xor XOR2 (N75, N69, N25);
nor NOR4 (N76, N67, N50, N38, N35);
nand NAND3 (N77, N68, N51, N13);
and AND4 (N78, N73, N76, N37, N60);
and AND2 (N79, N44, N13);
nor NOR4 (N80, N75, N73, N12, N47);
nand NAND2 (N81, N78, N3);
nor NOR4 (N82, N77, N23, N35, N56);
xor XOR2 (N83, N43, N59);
nand NAND3 (N84, N70, N60, N5);
or OR2 (N85, N71, N21);
buf BUF1 (N86, N58);
or OR4 (N87, N63, N21, N2, N30);
buf BUF1 (N88, N86);
and AND2 (N89, N87, N30);
or OR2 (N90, N80, N9);
and AND4 (N91, N82, N37, N74, N41);
nor NOR2 (N92, N12, N20);
xor XOR2 (N93, N81, N20);
buf BUF1 (N94, N90);
or OR4 (N95, N93, N67, N30, N44);
nor NOR2 (N96, N92, N65);
and AND3 (N97, N79, N82, N30);
nand NAND4 (N98, N85, N9, N85, N57);
not NOT1 (N99, N84);
or OR3 (N100, N97, N25, N84);
and AND3 (N101, N95, N39, N36);
nor NOR2 (N102, N94, N66);
buf BUF1 (N103, N100);
nor NOR3 (N104, N91, N7, N70);
xor XOR2 (N105, N102, N35);
nor NOR4 (N106, N103, N99, N30, N50);
xor XOR2 (N107, N48, N50);
nor NOR3 (N108, N89, N76, N11);
buf BUF1 (N109, N104);
xor XOR2 (N110, N96, N10);
xor XOR2 (N111, N110, N81);
nor NOR2 (N112, N83, N38);
not NOT1 (N113, N101);
not NOT1 (N114, N113);
not NOT1 (N115, N108);
or OR3 (N116, N106, N42, N57);
or OR2 (N117, N115, N116);
not NOT1 (N118, N98);
nand NAND4 (N119, N23, N4, N22, N38);
or OR3 (N120, N119, N45, N59);
nor NOR4 (N121, N88, N30, N85, N63);
xor XOR2 (N122, N118, N67);
buf BUF1 (N123, N117);
xor XOR2 (N124, N109, N96);
buf BUF1 (N125, N112);
buf BUF1 (N126, N120);
nand NAND3 (N127, N107, N84, N11);
buf BUF1 (N128, N124);
and AND3 (N129, N105, N76, N24);
xor XOR2 (N130, N122, N81);
buf BUF1 (N131, N130);
xor XOR2 (N132, N123, N3);
xor XOR2 (N133, N126, N82);
buf BUF1 (N134, N125);
not NOT1 (N135, N133);
nand NAND3 (N136, N132, N34, N96);
or OR4 (N137, N135, N136, N91, N76);
nor NOR3 (N138, N40, N121, N88);
xor XOR2 (N139, N60, N97);
xor XOR2 (N140, N114, N135);
xor XOR2 (N141, N129, N130);
not NOT1 (N142, N137);
not NOT1 (N143, N134);
or OR2 (N144, N128, N60);
xor XOR2 (N145, N141, N119);
or OR2 (N146, N138, N63);
nand NAND2 (N147, N140, N82);
nor NOR2 (N148, N127, N142);
not NOT1 (N149, N11);
nor NOR2 (N150, N143, N149);
not NOT1 (N151, N9);
nor NOR3 (N152, N147, N100, N76);
or OR2 (N153, N150, N137);
nand NAND4 (N154, N152, N99, N48, N141);
buf BUF1 (N155, N153);
nor NOR2 (N156, N111, N90);
nor NOR3 (N157, N155, N80, N88);
nor NOR3 (N158, N144, N14, N4);
nand NAND4 (N159, N151, N64, N136, N101);
xor XOR2 (N160, N158, N69);
xor XOR2 (N161, N145, N9);
and AND2 (N162, N157, N39);
nor NOR3 (N163, N161, N155, N77);
and AND3 (N164, N146, N5, N156);
buf BUF1 (N165, N64);
buf BUF1 (N166, N163);
nand NAND2 (N167, N154, N7);
nor NOR3 (N168, N162, N73, N76);
xor XOR2 (N169, N166, N116);
not NOT1 (N170, N164);
not NOT1 (N171, N160);
or OR2 (N172, N159, N18);
buf BUF1 (N173, N148);
nor NOR3 (N174, N171, N35, N4);
buf BUF1 (N175, N173);
not NOT1 (N176, N168);
xor XOR2 (N177, N139, N124);
not NOT1 (N178, N170);
nand NAND4 (N179, N176, N15, N123, N148);
xor XOR2 (N180, N131, N142);
not NOT1 (N181, N165);
nand NAND3 (N182, N181, N135, N133);
nor NOR3 (N183, N179, N150, N16);
or OR3 (N184, N182, N22, N153);
not NOT1 (N185, N167);
and AND3 (N186, N172, N15, N174);
buf BUF1 (N187, N6);
or OR2 (N188, N187, N106);
or OR4 (N189, N186, N16, N127, N108);
buf BUF1 (N190, N184);
or OR4 (N191, N178, N81, N52, N132);
nand NAND3 (N192, N189, N155, N169);
nand NAND3 (N193, N44, N165, N11);
xor XOR2 (N194, N175, N182);
and AND2 (N195, N185, N164);
and AND3 (N196, N188, N34, N132);
nand NAND3 (N197, N195, N40, N187);
nand NAND3 (N198, N190, N143, N26);
nand NAND4 (N199, N177, N87, N36, N167);
not NOT1 (N200, N197);
nand NAND4 (N201, N200, N192, N82, N56);
not NOT1 (N202, N1);
xor XOR2 (N203, N193, N26);
not NOT1 (N204, N201);
nand NAND2 (N205, N199, N31);
not NOT1 (N206, N203);
buf BUF1 (N207, N183);
not NOT1 (N208, N207);
and AND3 (N209, N180, N144, N92);
not NOT1 (N210, N208);
buf BUF1 (N211, N209);
and AND4 (N212, N204, N143, N53, N95);
xor XOR2 (N213, N198, N80);
nor NOR3 (N214, N191, N126, N206);
and AND2 (N215, N192, N208);
nor NOR4 (N216, N211, N157, N184, N133);
not NOT1 (N217, N212);
nor NOR2 (N218, N210, N132);
and AND2 (N219, N194, N79);
or OR3 (N220, N219, N131, N94);
or OR4 (N221, N220, N208, N51, N46);
not NOT1 (N222, N218);
nand NAND3 (N223, N196, N187, N168);
not NOT1 (N224, N202);
not NOT1 (N225, N214);
buf BUF1 (N226, N223);
and AND3 (N227, N217, N36, N77);
xor XOR2 (N228, N227, N203);
or OR4 (N229, N224, N116, N68, N72);
nor NOR3 (N230, N213, N135, N95);
xor XOR2 (N231, N221, N198);
nand NAND3 (N232, N226, N211, N106);
nand NAND3 (N233, N231, N179, N224);
nand NAND3 (N234, N233, N36, N170);
and AND4 (N235, N205, N213, N9, N171);
buf BUF1 (N236, N228);
buf BUF1 (N237, N230);
and AND3 (N238, N225, N29, N143);
or OR3 (N239, N222, N71, N44);
or OR4 (N240, N216, N41, N51, N18);
or OR2 (N241, N237, N93);
xor XOR2 (N242, N236, N157);
nor NOR3 (N243, N229, N131, N162);
not NOT1 (N244, N242);
not NOT1 (N245, N234);
xor XOR2 (N246, N243, N168);
nor NOR2 (N247, N238, N215);
and AND3 (N248, N45, N79, N130);
nor NOR3 (N249, N247, N76, N196);
buf BUF1 (N250, N249);
not NOT1 (N251, N246);
buf BUF1 (N252, N245);
and AND3 (N253, N241, N222, N250);
or OR4 (N254, N117, N248, N80, N42);
buf BUF1 (N255, N126);
and AND2 (N256, N232, N239);
nor NOR2 (N257, N58, N104);
xor XOR2 (N258, N252, N132);
and AND2 (N259, N251, N175);
and AND4 (N260, N254, N247, N31, N236);
nand NAND4 (N261, N256, N159, N185, N158);
xor XOR2 (N262, N244, N106);
not NOT1 (N263, N261);
nand NAND4 (N264, N257, N256, N41, N242);
nor NOR2 (N265, N258, N162);
xor XOR2 (N266, N263, N130);
nor NOR3 (N267, N255, N129, N132);
and AND3 (N268, N253, N255, N102);
buf BUF1 (N269, N265);
xor XOR2 (N270, N262, N39);
xor XOR2 (N271, N270, N231);
buf BUF1 (N272, N269);
xor XOR2 (N273, N271, N80);
nand NAND3 (N274, N260, N2, N14);
not NOT1 (N275, N274);
not NOT1 (N276, N235);
buf BUF1 (N277, N266);
nand NAND2 (N278, N240, N265);
nor NOR3 (N279, N273, N145, N61);
nand NAND2 (N280, N264, N145);
nand NAND2 (N281, N278, N85);
and AND3 (N282, N267, N245, N74);
buf BUF1 (N283, N268);
buf BUF1 (N284, N276);
buf BUF1 (N285, N283);
or OR3 (N286, N280, N258, N240);
not NOT1 (N287, N281);
not NOT1 (N288, N279);
buf BUF1 (N289, N287);
nand NAND3 (N290, N259, N266, N198);
nand NAND2 (N291, N288, N90);
nor NOR2 (N292, N275, N39);
or OR2 (N293, N291, N10);
nand NAND3 (N294, N290, N74, N66);
xor XOR2 (N295, N293, N269);
buf BUF1 (N296, N286);
xor XOR2 (N297, N294, N146);
and AND4 (N298, N297, N99, N127, N227);
nor NOR3 (N299, N298, N58, N60);
xor XOR2 (N300, N299, N67);
and AND2 (N301, N300, N10);
nor NOR4 (N302, N289, N77, N223, N250);
buf BUF1 (N303, N282);
nor NOR2 (N304, N272, N201);
and AND3 (N305, N284, N217, N126);
or OR2 (N306, N295, N10);
or OR2 (N307, N301, N151);
nand NAND4 (N308, N277, N289, N178, N184);
nor NOR4 (N309, N308, N15, N227, N179);
nor NOR3 (N310, N306, N177, N157);
nor NOR2 (N311, N302, N80);
not NOT1 (N312, N303);
buf BUF1 (N313, N310);
not NOT1 (N314, N312);
or OR2 (N315, N292, N42);
nor NOR4 (N316, N313, N242, N189, N68);
nand NAND3 (N317, N316, N242, N108);
nor NOR3 (N318, N317, N151, N286);
buf BUF1 (N319, N309);
not NOT1 (N320, N296);
xor XOR2 (N321, N304, N100);
not NOT1 (N322, N320);
buf BUF1 (N323, N318);
nor NOR2 (N324, N322, N208);
or OR2 (N325, N315, N309);
and AND2 (N326, N307, N287);
buf BUF1 (N327, N325);
or OR4 (N328, N319, N169, N36, N199);
not NOT1 (N329, N328);
nand NAND4 (N330, N329, N3, N75, N58);
buf BUF1 (N331, N326);
xor XOR2 (N332, N311, N282);
xor XOR2 (N333, N285, N226);
or OR4 (N334, N331, N26, N5, N158);
or OR2 (N335, N332, N245);
nor NOR2 (N336, N333, N150);
nor NOR4 (N337, N335, N128, N143, N298);
xor XOR2 (N338, N334, N104);
and AND2 (N339, N327, N24);
buf BUF1 (N340, N338);
xor XOR2 (N341, N336, N249);
not NOT1 (N342, N341);
nor NOR2 (N343, N314, N325);
nor NOR2 (N344, N323, N135);
xor XOR2 (N345, N339, N42);
and AND4 (N346, N344, N237, N90, N208);
buf BUF1 (N347, N337);
nand NAND3 (N348, N346, N38, N168);
xor XOR2 (N349, N321, N152);
nand NAND2 (N350, N324, N349);
buf BUF1 (N351, N90);
buf BUF1 (N352, N347);
nor NOR2 (N353, N343, N169);
not NOT1 (N354, N350);
or OR2 (N355, N353, N18);
and AND2 (N356, N345, N234);
xor XOR2 (N357, N330, N19);
or OR3 (N358, N351, N58, N211);
xor XOR2 (N359, N356, N187);
not NOT1 (N360, N354);
buf BUF1 (N361, N342);
xor XOR2 (N362, N360, N332);
and AND4 (N363, N359, N287, N11, N282);
xor XOR2 (N364, N358, N165);
xor XOR2 (N365, N352, N97);
nor NOR2 (N366, N362, N29);
nand NAND4 (N367, N355, N271, N14, N330);
nor NOR3 (N368, N340, N143, N129);
buf BUF1 (N369, N363);
xor XOR2 (N370, N348, N171);
not NOT1 (N371, N305);
nor NOR3 (N372, N371, N153, N74);
nor NOR2 (N373, N372, N205);
and AND4 (N374, N369, N159, N363, N233);
nor NOR4 (N375, N368, N32, N171, N229);
buf BUF1 (N376, N361);
xor XOR2 (N377, N365, N178);
nor NOR4 (N378, N366, N269, N233, N91);
or OR2 (N379, N357, N46);
and AND4 (N380, N376, N1, N91, N219);
and AND2 (N381, N380, N298);
not NOT1 (N382, N381);
xor XOR2 (N383, N364, N181);
not NOT1 (N384, N374);
nand NAND2 (N385, N378, N108);
xor XOR2 (N386, N385, N50);
nor NOR3 (N387, N373, N316, N308);
buf BUF1 (N388, N386);
and AND3 (N389, N377, N249, N19);
and AND3 (N390, N382, N239, N284);
xor XOR2 (N391, N375, N281);
nand NAND4 (N392, N379, N301, N43, N199);
and AND3 (N393, N370, N208, N9);
nor NOR2 (N394, N383, N104);
and AND3 (N395, N392, N83, N46);
buf BUF1 (N396, N384);
and AND4 (N397, N393, N364, N146, N271);
nand NAND2 (N398, N397, N247);
nand NAND4 (N399, N390, N71, N243, N25);
buf BUF1 (N400, N394);
not NOT1 (N401, N389);
not NOT1 (N402, N399);
or OR3 (N403, N395, N248, N72);
nand NAND2 (N404, N401, N337);
nand NAND3 (N405, N391, N90, N302);
xor XOR2 (N406, N396, N361);
buf BUF1 (N407, N403);
nand NAND3 (N408, N406, N144, N77);
buf BUF1 (N409, N404);
or OR2 (N410, N367, N125);
not NOT1 (N411, N398);
not NOT1 (N412, N400);
not NOT1 (N413, N410);
or OR4 (N414, N411, N378, N367, N88);
or OR2 (N415, N412, N411);
nand NAND2 (N416, N415, N294);
nand NAND2 (N417, N416, N295);
not NOT1 (N418, N414);
or OR4 (N419, N418, N113, N72, N183);
not NOT1 (N420, N413);
not NOT1 (N421, N408);
and AND3 (N422, N405, N25, N81);
buf BUF1 (N423, N409);
or OR4 (N424, N422, N90, N246, N77);
buf BUF1 (N425, N388);
xor XOR2 (N426, N423, N328);
xor XOR2 (N427, N426, N334);
and AND4 (N428, N427, N334, N360, N13);
nand NAND4 (N429, N428, N374, N276, N20);
nor NOR2 (N430, N387, N107);
or OR4 (N431, N407, N195, N287, N152);
nand NAND3 (N432, N417, N130, N115);
xor XOR2 (N433, N421, N142);
xor XOR2 (N434, N431, N300);
xor XOR2 (N435, N430, N187);
nor NOR3 (N436, N434, N403, N198);
buf BUF1 (N437, N419);
xor XOR2 (N438, N402, N373);
xor XOR2 (N439, N424, N152);
and AND3 (N440, N435, N61, N282);
or OR2 (N441, N440, N14);
not NOT1 (N442, N433);
xor XOR2 (N443, N436, N435);
not NOT1 (N444, N441);
nor NOR4 (N445, N438, N51, N126, N83);
buf BUF1 (N446, N439);
not NOT1 (N447, N444);
xor XOR2 (N448, N446, N284);
buf BUF1 (N449, N425);
not NOT1 (N450, N448);
not NOT1 (N451, N432);
buf BUF1 (N452, N420);
xor XOR2 (N453, N442, N75);
buf BUF1 (N454, N451);
or OR3 (N455, N437, N437, N94);
nand NAND2 (N456, N443, N350);
buf BUF1 (N457, N445);
nand NAND3 (N458, N450, N36, N256);
buf BUF1 (N459, N458);
nor NOR4 (N460, N452, N98, N84, N96);
and AND3 (N461, N455, N389, N351);
nor NOR3 (N462, N454, N31, N211);
nor NOR3 (N463, N453, N428, N399);
nand NAND3 (N464, N449, N81, N255);
buf BUF1 (N465, N464);
and AND2 (N466, N429, N150);
buf BUF1 (N467, N463);
xor XOR2 (N468, N447, N267);
nor NOR4 (N469, N462, N297, N106, N360);
or OR2 (N470, N460, N312);
xor XOR2 (N471, N469, N461);
or OR4 (N472, N50, N286, N293, N260);
nand NAND4 (N473, N456, N6, N398, N157);
buf BUF1 (N474, N472);
or OR2 (N475, N457, N44);
and AND2 (N476, N468, N56);
nor NOR2 (N477, N473, N199);
nand NAND2 (N478, N476, N451);
not NOT1 (N479, N474);
nand NAND4 (N480, N467, N99, N184, N328);
not NOT1 (N481, N475);
nor NOR3 (N482, N481, N29, N451);
or OR2 (N483, N465, N93);
nand NAND3 (N484, N482, N250, N242);
nand NAND2 (N485, N477, N357);
and AND4 (N486, N483, N397, N404, N443);
nor NOR2 (N487, N478, N314);
and AND3 (N488, N485, N180, N362);
buf BUF1 (N489, N459);
or OR4 (N490, N480, N199, N422, N219);
and AND2 (N491, N489, N433);
not NOT1 (N492, N486);
not NOT1 (N493, N487);
not NOT1 (N494, N490);
and AND4 (N495, N493, N277, N139, N22);
xor XOR2 (N496, N484, N301);
xor XOR2 (N497, N491, N27);
not NOT1 (N498, N488);
not NOT1 (N499, N492);
and AND2 (N500, N494, N475);
xor XOR2 (N501, N498, N366);
xor XOR2 (N502, N471, N439);
and AND3 (N503, N470, N427, N485);
nand NAND3 (N504, N501, N486, N192);
buf BUF1 (N505, N503);
and AND4 (N506, N500, N426, N356, N327);
not NOT1 (N507, N506);
buf BUF1 (N508, N505);
not NOT1 (N509, N479);
nor NOR4 (N510, N508, N97, N156, N240);
nand NAND2 (N511, N499, N404);
and AND4 (N512, N495, N400, N234, N256);
buf BUF1 (N513, N502);
xor XOR2 (N514, N513, N491);
xor XOR2 (N515, N466, N287);
and AND4 (N516, N515, N330, N50, N59);
buf BUF1 (N517, N507);
xor XOR2 (N518, N504, N377);
nor NOR3 (N519, N516, N422, N119);
not NOT1 (N520, N518);
or OR3 (N521, N520, N327, N154);
or OR2 (N522, N497, N129);
nand NAND3 (N523, N512, N34, N138);
nor NOR2 (N524, N511, N354);
buf BUF1 (N525, N509);
not NOT1 (N526, N496);
nor NOR3 (N527, N517, N233, N491);
not NOT1 (N528, N514);
nor NOR4 (N529, N526, N465, N95, N66);
not NOT1 (N530, N521);
and AND3 (N531, N529, N40, N154);
nand NAND4 (N532, N530, N84, N521, N27);
xor XOR2 (N533, N527, N459);
not NOT1 (N534, N525);
not NOT1 (N535, N534);
xor XOR2 (N536, N531, N446);
nand NAND4 (N537, N524, N213, N285, N51);
buf BUF1 (N538, N528);
xor XOR2 (N539, N522, N130);
or OR4 (N540, N536, N28, N205, N166);
nand NAND2 (N541, N533, N165);
nor NOR2 (N542, N538, N191);
xor XOR2 (N543, N537, N449);
xor XOR2 (N544, N542, N452);
not NOT1 (N545, N523);
nand NAND4 (N546, N510, N5, N148, N44);
nand NAND4 (N547, N541, N427, N96, N512);
not NOT1 (N548, N545);
xor XOR2 (N549, N532, N342);
and AND4 (N550, N549, N168, N342, N84);
and AND4 (N551, N548, N256, N384, N350);
and AND2 (N552, N540, N187);
buf BUF1 (N553, N551);
buf BUF1 (N554, N547);
nor NOR3 (N555, N535, N308, N450);
nand NAND4 (N556, N553, N432, N409, N521);
nand NAND3 (N557, N550, N287, N46);
and AND3 (N558, N552, N480, N215);
xor XOR2 (N559, N543, N148);
and AND3 (N560, N519, N242, N536);
nand NAND3 (N561, N558, N506, N489);
buf BUF1 (N562, N556);
buf BUF1 (N563, N559);
and AND3 (N564, N539, N19, N42);
not NOT1 (N565, N557);
nor NOR3 (N566, N554, N27, N245);
nor NOR3 (N567, N562, N152, N253);
not NOT1 (N568, N560);
nor NOR3 (N569, N567, N381, N128);
or OR2 (N570, N568, N53);
nand NAND2 (N571, N569, N219);
and AND2 (N572, N563, N19);
nand NAND3 (N573, N555, N165, N447);
xor XOR2 (N574, N573, N536);
or OR2 (N575, N565, N33);
nand NAND3 (N576, N544, N469, N359);
xor XOR2 (N577, N546, N560);
nand NAND4 (N578, N564, N260, N547, N173);
nand NAND3 (N579, N561, N449, N254);
buf BUF1 (N580, N566);
and AND2 (N581, N579, N397);
nor NOR3 (N582, N577, N442, N464);
nand NAND3 (N583, N570, N289, N482);
buf BUF1 (N584, N582);
buf BUF1 (N585, N576);
buf BUF1 (N586, N581);
buf BUF1 (N587, N572);
and AND4 (N588, N587, N262, N454, N320);
not NOT1 (N589, N583);
or OR4 (N590, N589, N211, N189, N58);
xor XOR2 (N591, N571, N479);
nand NAND4 (N592, N590, N193, N66, N138);
nor NOR3 (N593, N591, N403, N354);
xor XOR2 (N594, N575, N512);
nor NOR4 (N595, N592, N196, N287, N43);
buf BUF1 (N596, N595);
not NOT1 (N597, N593);
not NOT1 (N598, N584);
and AND2 (N599, N596, N389);
xor XOR2 (N600, N588, N294);
xor XOR2 (N601, N585, N570);
nand NAND2 (N602, N578, N159);
nand NAND4 (N603, N598, N286, N17, N158);
or OR4 (N604, N574, N558, N602, N281);
nor NOR2 (N605, N529, N540);
and AND3 (N606, N597, N127, N545);
nor NOR3 (N607, N594, N144, N222);
nand NAND4 (N608, N605, N232, N25, N583);
nand NAND4 (N609, N603, N174, N461, N226);
xor XOR2 (N610, N604, N203);
buf BUF1 (N611, N599);
nor NOR3 (N612, N610, N274, N476);
or OR4 (N613, N609, N480, N167, N540);
xor XOR2 (N614, N601, N257);
and AND2 (N615, N608, N427);
not NOT1 (N616, N580);
nor NOR4 (N617, N606, N242, N49, N419);
buf BUF1 (N618, N600);
buf BUF1 (N619, N617);
not NOT1 (N620, N586);
or OR4 (N621, N620, N195, N388, N53);
nand NAND4 (N622, N614, N139, N423, N4);
or OR2 (N623, N607, N543);
xor XOR2 (N624, N618, N423);
and AND4 (N625, N612, N449, N88, N303);
nand NAND2 (N626, N624, N28);
and AND4 (N627, N619, N60, N491, N112);
and AND3 (N628, N626, N293, N448);
nand NAND4 (N629, N611, N434, N18, N235);
not NOT1 (N630, N621);
nand NAND4 (N631, N615, N312, N286, N499);
buf BUF1 (N632, N631);
and AND3 (N633, N628, N484, N407);
buf BUF1 (N634, N627);
and AND4 (N635, N633, N153, N24, N69);
and AND2 (N636, N625, N525);
or OR3 (N637, N613, N121, N431);
not NOT1 (N638, N632);
xor XOR2 (N639, N636, N134);
nor NOR3 (N640, N635, N193, N439);
and AND2 (N641, N634, N77);
nor NOR3 (N642, N641, N513, N37);
nand NAND3 (N643, N623, N100, N392);
xor XOR2 (N644, N630, N258);
buf BUF1 (N645, N638);
not NOT1 (N646, N644);
and AND4 (N647, N645, N144, N509, N44);
nor NOR4 (N648, N640, N13, N422, N83);
nor NOR2 (N649, N647, N174);
and AND2 (N650, N629, N370);
nand NAND3 (N651, N616, N206, N29);
xor XOR2 (N652, N622, N11);
xor XOR2 (N653, N649, N417);
and AND3 (N654, N643, N441, N70);
xor XOR2 (N655, N639, N396);
buf BUF1 (N656, N637);
not NOT1 (N657, N655);
and AND4 (N658, N653, N45, N477, N227);
xor XOR2 (N659, N656, N425);
or OR3 (N660, N659, N456, N527);
not NOT1 (N661, N646);
and AND3 (N662, N642, N45, N588);
buf BUF1 (N663, N657);
nand NAND4 (N664, N660, N404, N43, N442);
not NOT1 (N665, N664);
nand NAND4 (N666, N663, N443, N362, N592);
buf BUF1 (N667, N650);
and AND2 (N668, N661, N210);
nor NOR4 (N669, N668, N282, N110, N30);
nand NAND2 (N670, N651, N68);
or OR2 (N671, N652, N398);
nor NOR4 (N672, N667, N369, N612, N64);
nor NOR4 (N673, N666, N317, N589, N520);
buf BUF1 (N674, N672);
not NOT1 (N675, N674);
or OR2 (N676, N658, N412);
xor XOR2 (N677, N675, N417);
and AND4 (N678, N673, N95, N349, N392);
not NOT1 (N679, N678);
buf BUF1 (N680, N671);
not NOT1 (N681, N676);
or OR4 (N682, N670, N423, N240, N611);
nor NOR2 (N683, N677, N654);
not NOT1 (N684, N484);
not NOT1 (N685, N648);
buf BUF1 (N686, N669);
nand NAND4 (N687, N681, N474, N8, N397);
xor XOR2 (N688, N687, N417);
not NOT1 (N689, N680);
buf BUF1 (N690, N684);
xor XOR2 (N691, N665, N635);
buf BUF1 (N692, N686);
nor NOR3 (N693, N662, N416, N305);
and AND4 (N694, N690, N203, N102, N457);
and AND4 (N695, N693, N445, N294, N579);
xor XOR2 (N696, N688, N259);
buf BUF1 (N697, N691);
xor XOR2 (N698, N692, N201);
xor XOR2 (N699, N694, N543);
nor NOR2 (N700, N685, N415);
xor XOR2 (N701, N689, N108);
not NOT1 (N702, N695);
not NOT1 (N703, N696);
not NOT1 (N704, N683);
or OR4 (N705, N697, N159, N681, N400);
xor XOR2 (N706, N682, N366);
and AND3 (N707, N702, N481, N79);
not NOT1 (N708, N705);
nand NAND4 (N709, N698, N33, N412, N163);
not NOT1 (N710, N708);
nand NAND3 (N711, N703, N552, N568);
buf BUF1 (N712, N709);
not NOT1 (N713, N701);
buf BUF1 (N714, N679);
buf BUF1 (N715, N704);
nor NOR4 (N716, N710, N349, N155, N333);
nand NAND2 (N717, N707, N181);
or OR3 (N718, N715, N76, N416);
or OR2 (N719, N700, N33);
nand NAND4 (N720, N717, N257, N334, N66);
and AND2 (N721, N716, N537);
buf BUF1 (N722, N706);
nand NAND2 (N723, N712, N240);
and AND4 (N724, N713, N508, N25, N34);
and AND4 (N725, N720, N374, N478, N655);
xor XOR2 (N726, N724, N199);
nand NAND2 (N727, N719, N476);
and AND2 (N728, N718, N188);
nor NOR4 (N729, N722, N401, N633, N271);
and AND4 (N730, N711, N160, N97, N367);
xor XOR2 (N731, N723, N723);
or OR4 (N732, N699, N64, N715, N663);
not NOT1 (N733, N731);
nand NAND3 (N734, N727, N539, N673);
buf BUF1 (N735, N721);
not NOT1 (N736, N726);
nor NOR4 (N737, N725, N333, N661, N27);
xor XOR2 (N738, N734, N595);
not NOT1 (N739, N733);
buf BUF1 (N740, N738);
nor NOR3 (N741, N728, N658, N470);
not NOT1 (N742, N741);
nor NOR2 (N743, N736, N227);
nor NOR2 (N744, N743, N253);
buf BUF1 (N745, N744);
xor XOR2 (N746, N730, N420);
xor XOR2 (N747, N729, N466);
nand NAND3 (N748, N740, N537, N709);
nand NAND4 (N749, N747, N261, N465, N203);
xor XOR2 (N750, N745, N335);
and AND2 (N751, N746, N725);
nor NOR3 (N752, N748, N348, N638);
and AND2 (N753, N737, N17);
nand NAND2 (N754, N739, N204);
not NOT1 (N755, N749);
nor NOR3 (N756, N754, N590, N127);
or OR2 (N757, N750, N109);
nand NAND4 (N758, N714, N654, N43, N696);
not NOT1 (N759, N757);
nor NOR2 (N760, N732, N10);
nor NOR3 (N761, N753, N64, N219);
nor NOR4 (N762, N760, N342, N134, N449);
nor NOR3 (N763, N762, N316, N184);
nor NOR3 (N764, N756, N644, N530);
nor NOR2 (N765, N742, N537);
or OR2 (N766, N765, N439);
xor XOR2 (N767, N735, N168);
nand NAND4 (N768, N766, N5, N81, N651);
xor XOR2 (N769, N763, N95);
nand NAND2 (N770, N761, N629);
or OR3 (N771, N769, N549, N152);
nand NAND4 (N772, N755, N738, N428, N260);
buf BUF1 (N773, N770);
nor NOR4 (N774, N768, N445, N361, N550);
buf BUF1 (N775, N771);
buf BUF1 (N776, N775);
not NOT1 (N777, N751);
buf BUF1 (N778, N759);
not NOT1 (N779, N767);
nor NOR2 (N780, N752, N274);
nand NAND2 (N781, N764, N189);
not NOT1 (N782, N772);
xor XOR2 (N783, N777, N356);
nand NAND2 (N784, N779, N740);
nand NAND2 (N785, N784, N490);
buf BUF1 (N786, N774);
buf BUF1 (N787, N785);
and AND2 (N788, N776, N79);
buf BUF1 (N789, N780);
buf BUF1 (N790, N782);
buf BUF1 (N791, N758);
and AND2 (N792, N791, N118);
buf BUF1 (N793, N787);
xor XOR2 (N794, N778, N145);
buf BUF1 (N795, N794);
nor NOR4 (N796, N781, N795, N579, N191);
xor XOR2 (N797, N438, N474);
not NOT1 (N798, N783);
nand NAND3 (N799, N789, N89, N695);
nor NOR3 (N800, N798, N183, N689);
and AND2 (N801, N797, N491);
and AND4 (N802, N800, N551, N471, N104);
nor NOR2 (N803, N801, N101);
xor XOR2 (N804, N786, N578);
buf BUF1 (N805, N796);
nand NAND4 (N806, N773, N220, N275, N305);
not NOT1 (N807, N788);
and AND3 (N808, N806, N63, N556);
xor XOR2 (N809, N790, N263);
and AND4 (N810, N805, N197, N430, N138);
or OR3 (N811, N799, N220, N657);
buf BUF1 (N812, N804);
or OR2 (N813, N808, N706);
buf BUF1 (N814, N809);
xor XOR2 (N815, N793, N217);
buf BUF1 (N816, N803);
buf BUF1 (N817, N802);
nor NOR4 (N818, N807, N783, N490, N438);
not NOT1 (N819, N814);
buf BUF1 (N820, N812);
buf BUF1 (N821, N817);
and AND2 (N822, N792, N512);
buf BUF1 (N823, N811);
and AND4 (N824, N819, N73, N52, N743);
buf BUF1 (N825, N810);
xor XOR2 (N826, N824, N633);
and AND3 (N827, N813, N648, N116);
nor NOR2 (N828, N825, N352);
buf BUF1 (N829, N821);
nand NAND4 (N830, N826, N807, N398, N265);
not NOT1 (N831, N823);
or OR2 (N832, N829, N725);
nand NAND4 (N833, N820, N188, N534, N446);
not NOT1 (N834, N815);
nor NOR2 (N835, N831, N345);
or OR4 (N836, N822, N23, N509, N297);
buf BUF1 (N837, N818);
buf BUF1 (N838, N832);
not NOT1 (N839, N830);
or OR4 (N840, N828, N149, N245, N724);
buf BUF1 (N841, N827);
or OR2 (N842, N838, N819);
and AND3 (N843, N841, N655, N560);
buf BUF1 (N844, N840);
nor NOR3 (N845, N842, N538, N633);
buf BUF1 (N846, N834);
or OR4 (N847, N843, N1, N700, N485);
buf BUF1 (N848, N836);
not NOT1 (N849, N816);
buf BUF1 (N850, N835);
buf BUF1 (N851, N837);
buf BUF1 (N852, N847);
and AND2 (N853, N848, N547);
buf BUF1 (N854, N850);
and AND4 (N855, N852, N124, N642, N778);
xor XOR2 (N856, N853, N753);
buf BUF1 (N857, N845);
or OR2 (N858, N844, N46);
not NOT1 (N859, N857);
or OR4 (N860, N854, N771, N627, N76);
nand NAND2 (N861, N833, N475);
xor XOR2 (N862, N855, N67);
buf BUF1 (N863, N839);
nand NAND4 (N864, N862, N531, N353, N620);
or OR4 (N865, N849, N249, N429, N219);
nor NOR4 (N866, N861, N730, N297, N426);
and AND3 (N867, N864, N578, N160);
and AND3 (N868, N858, N44, N36);
nor NOR2 (N869, N867, N860);
or OR2 (N870, N179, N294);
and AND2 (N871, N870, N10);
or OR2 (N872, N869, N366);
not NOT1 (N873, N851);
not NOT1 (N874, N865);
or OR2 (N875, N871, N659);
nand NAND3 (N876, N859, N527, N718);
or OR2 (N877, N866, N243);
nor NOR4 (N878, N872, N801, N1, N732);
nor NOR3 (N879, N878, N393, N84);
or OR4 (N880, N877, N786, N854, N318);
nand NAND4 (N881, N863, N667, N146, N553);
nor NOR3 (N882, N846, N777, N125);
and AND4 (N883, N868, N157, N821, N328);
nor NOR4 (N884, N873, N480, N614, N332);
buf BUF1 (N885, N883);
nand NAND2 (N886, N875, N612);
xor XOR2 (N887, N879, N513);
nor NOR3 (N888, N882, N872, N625);
and AND3 (N889, N856, N610, N626);
or OR2 (N890, N876, N581);
nand NAND3 (N891, N885, N430, N721);
and AND2 (N892, N888, N111);
nor NOR4 (N893, N887, N763, N378, N408);
buf BUF1 (N894, N892);
and AND2 (N895, N891, N630);
buf BUF1 (N896, N890);
buf BUF1 (N897, N886);
buf BUF1 (N898, N881);
xor XOR2 (N899, N896, N133);
nand NAND3 (N900, N874, N372, N375);
not NOT1 (N901, N897);
xor XOR2 (N902, N898, N378);
nor NOR2 (N903, N880, N605);
nand NAND4 (N904, N884, N334, N767, N74);
nor NOR3 (N905, N894, N791, N159);
nand NAND2 (N906, N899, N488);
nor NOR4 (N907, N902, N31, N661, N379);
nor NOR3 (N908, N895, N620, N78);
not NOT1 (N909, N904);
nand NAND4 (N910, N906, N131, N100, N704);
or OR3 (N911, N909, N153, N345);
not NOT1 (N912, N910);
or OR2 (N913, N903, N389);
nand NAND2 (N914, N905, N689);
not NOT1 (N915, N893);
buf BUF1 (N916, N901);
not NOT1 (N917, N911);
not NOT1 (N918, N908);
buf BUF1 (N919, N889);
not NOT1 (N920, N915);
and AND2 (N921, N918, N423);
or OR3 (N922, N912, N320, N899);
nor NOR3 (N923, N922, N166, N714);
or OR2 (N924, N907, N554);
and AND4 (N925, N919, N355, N643, N196);
nand NAND3 (N926, N921, N849, N37);
nand NAND4 (N927, N917, N590, N349, N433);
or OR3 (N928, N913, N355, N77);
buf BUF1 (N929, N924);
not NOT1 (N930, N927);
or OR4 (N931, N914, N741, N800, N197);
not NOT1 (N932, N916);
nand NAND2 (N933, N920, N651);
nor NOR4 (N934, N931, N542, N198, N759);
and AND2 (N935, N934, N153);
and AND4 (N936, N929, N524, N55, N676);
nor NOR2 (N937, N933, N829);
nor NOR3 (N938, N930, N343, N39);
xor XOR2 (N939, N923, N35);
or OR4 (N940, N900, N606, N105, N929);
and AND2 (N941, N935, N192);
not NOT1 (N942, N925);
and AND3 (N943, N926, N312, N535);
or OR4 (N944, N932, N783, N634, N889);
nand NAND3 (N945, N943, N921, N413);
and AND4 (N946, N936, N885, N200, N489);
buf BUF1 (N947, N937);
and AND3 (N948, N944, N850, N713);
not NOT1 (N949, N928);
or OR3 (N950, N938, N239, N819);
and AND4 (N951, N939, N248, N796, N39);
nor NOR3 (N952, N945, N11, N574);
nor NOR2 (N953, N951, N571);
nor NOR3 (N954, N946, N106, N491);
and AND2 (N955, N950, N98);
buf BUF1 (N956, N948);
not NOT1 (N957, N942);
or OR4 (N958, N940, N829, N271, N268);
or OR4 (N959, N952, N693, N139, N120);
and AND2 (N960, N954, N333);
xor XOR2 (N961, N953, N718);
xor XOR2 (N962, N949, N272);
nor NOR4 (N963, N955, N487, N434, N586);
or OR3 (N964, N962, N606, N293);
buf BUF1 (N965, N964);
and AND4 (N966, N941, N173, N475, N429);
and AND3 (N967, N966, N839, N744);
or OR4 (N968, N967, N657, N394, N18);
not NOT1 (N969, N965);
and AND4 (N970, N963, N796, N922, N917);
nand NAND3 (N971, N968, N699, N508);
not NOT1 (N972, N958);
nor NOR2 (N973, N971, N138);
or OR2 (N974, N972, N651);
and AND4 (N975, N961, N840, N778, N282);
xor XOR2 (N976, N960, N525);
buf BUF1 (N977, N973);
xor XOR2 (N978, N959, N377);
or OR2 (N979, N976, N84);
nand NAND4 (N980, N957, N816, N201, N829);
buf BUF1 (N981, N974);
nor NOR3 (N982, N970, N286, N609);
not NOT1 (N983, N982);
buf BUF1 (N984, N979);
nand NAND2 (N985, N980, N528);
or OR4 (N986, N978, N950, N486, N483);
not NOT1 (N987, N977);
or OR3 (N988, N985, N779, N724);
not NOT1 (N989, N988);
not NOT1 (N990, N956);
and AND2 (N991, N983, N403);
not NOT1 (N992, N975);
or OR2 (N993, N947, N361);
and AND2 (N994, N969, N158);
and AND3 (N995, N994, N872, N221);
nand NAND3 (N996, N995, N309, N437);
not NOT1 (N997, N989);
or OR4 (N998, N981, N423, N730, N108);
xor XOR2 (N999, N984, N116);
xor XOR2 (N1000, N990, N661);
buf BUF1 (N1001, N1000);
not NOT1 (N1002, N986);
and AND4 (N1003, N1001, N516, N223, N939);
and AND3 (N1004, N999, N290, N417);
buf BUF1 (N1005, N997);
not NOT1 (N1006, N1002);
buf BUF1 (N1007, N1006);
nor NOR2 (N1008, N987, N83);
not NOT1 (N1009, N998);
or OR4 (N1010, N992, N252, N290, N368);
nor NOR3 (N1011, N991, N643, N674);
buf BUF1 (N1012, N1004);
xor XOR2 (N1013, N1003, N82);
not NOT1 (N1014, N1008);
or OR3 (N1015, N996, N374, N182);
nor NOR2 (N1016, N1011, N164);
nor NOR2 (N1017, N1012, N760);
or OR3 (N1018, N1013, N279, N840);
nor NOR2 (N1019, N1015, N643);
not NOT1 (N1020, N1007);
not NOT1 (N1021, N993);
not NOT1 (N1022, N1021);
and AND3 (N1023, N1005, N778, N828);
and AND3 (N1024, N1023, N82, N739);
endmodule