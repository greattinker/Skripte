// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20;

output N217,N219,N218,N200,N207,N216,N212,N215,N204,N220;

and AND4 (N21, N19, N19, N6, N15);
xor XOR2 (N22, N11, N2);
nand NAND4 (N23, N20, N21, N10, N10);
buf BUF1 (N24, N7);
buf BUF1 (N25, N10);
buf BUF1 (N26, N11);
nor NOR2 (N27, N20, N19);
and AND2 (N28, N12, N11);
nor NOR3 (N29, N3, N26, N6);
nor NOR3 (N30, N19, N22, N26);
xor XOR2 (N31, N5, N3);
nor NOR4 (N32, N8, N4, N29, N30);
and AND2 (N33, N31, N10);
xor XOR2 (N34, N4, N9);
or OR4 (N35, N9, N32, N22, N19);
nand NAND4 (N36, N35, N6, N23, N3);
or OR3 (N37, N17, N8, N14);
buf BUF1 (N38, N4);
xor XOR2 (N39, N29, N15);
nand NAND2 (N40, N39, N21);
nand NAND2 (N41, N27, N33);
buf BUF1 (N42, N28);
nand NAND4 (N43, N27, N35, N23, N30);
or OR3 (N44, N37, N40, N2);
xor XOR2 (N45, N8, N40);
buf BUF1 (N46, N36);
nand NAND4 (N47, N41, N27, N21, N43);
nor NOR4 (N48, N37, N36, N24, N10);
nor NOR2 (N49, N19, N11);
or OR3 (N50, N45, N14, N2);
nand NAND3 (N51, N46, N13, N50);
nor NOR4 (N52, N29, N9, N37, N13);
buf BUF1 (N53, N52);
nor NOR2 (N54, N49, N27);
not NOT1 (N55, N54);
xor XOR2 (N56, N42, N24);
or OR2 (N57, N53, N40);
xor XOR2 (N58, N47, N25);
nor NOR4 (N59, N44, N47, N23, N28);
buf BUF1 (N60, N22);
and AND3 (N61, N38, N37, N13);
buf BUF1 (N62, N59);
buf BUF1 (N63, N61);
or OR4 (N64, N63, N26, N9, N49);
not NOT1 (N65, N55);
not NOT1 (N66, N56);
nand NAND3 (N67, N62, N1, N1);
nand NAND2 (N68, N58, N22);
nor NOR3 (N69, N48, N21, N52);
and AND2 (N70, N69, N64);
xor XOR2 (N71, N36, N45);
nor NOR4 (N72, N51, N44, N28, N23);
and AND2 (N73, N71, N59);
xor XOR2 (N74, N57, N30);
xor XOR2 (N75, N34, N74);
xor XOR2 (N76, N64, N33);
buf BUF1 (N77, N67);
not NOT1 (N78, N68);
nor NOR2 (N79, N75, N34);
nand NAND3 (N80, N66, N40, N31);
nand NAND4 (N81, N73, N70, N59, N70);
buf BUF1 (N82, N81);
buf BUF1 (N83, N5);
not NOT1 (N84, N83);
not NOT1 (N85, N60);
not NOT1 (N86, N82);
and AND4 (N87, N65, N9, N2, N50);
nand NAND2 (N88, N85, N51);
not NOT1 (N89, N80);
xor XOR2 (N90, N84, N23);
or OR2 (N91, N88, N75);
xor XOR2 (N92, N89, N80);
nand NAND2 (N93, N90, N75);
or OR4 (N94, N79, N26, N13, N69);
or OR3 (N95, N93, N47, N45);
and AND2 (N96, N95, N26);
or OR4 (N97, N87, N68, N72, N92);
not NOT1 (N98, N3);
xor XOR2 (N99, N73, N83);
xor XOR2 (N100, N86, N75);
buf BUF1 (N101, N91);
not NOT1 (N102, N76);
nor NOR2 (N103, N96, N47);
buf BUF1 (N104, N77);
xor XOR2 (N105, N101, N5);
xor XOR2 (N106, N103, N57);
or OR3 (N107, N105, N50, N42);
nor NOR2 (N108, N94, N85);
nand NAND4 (N109, N107, N66, N34, N42);
or OR4 (N110, N106, N92, N19, N95);
nand NAND3 (N111, N102, N50, N27);
buf BUF1 (N112, N104);
or OR2 (N113, N112, N48);
xor XOR2 (N114, N108, N14);
or OR3 (N115, N100, N2, N74);
or OR4 (N116, N97, N56, N54, N109);
nor NOR4 (N117, N33, N4, N93, N110);
not NOT1 (N118, N39);
buf BUF1 (N119, N113);
or OR4 (N120, N98, N13, N97, N33);
nand NAND2 (N121, N115, N41);
not NOT1 (N122, N116);
xor XOR2 (N123, N118, N60);
nor NOR4 (N124, N120, N3, N83, N55);
or OR2 (N125, N119, N85);
xor XOR2 (N126, N117, N116);
xor XOR2 (N127, N124, N56);
not NOT1 (N128, N122);
xor XOR2 (N129, N127, N18);
buf BUF1 (N130, N99);
xor XOR2 (N131, N125, N14);
buf BUF1 (N132, N114);
or OR2 (N133, N132, N81);
or OR4 (N134, N129, N34, N119, N105);
not NOT1 (N135, N134);
and AND4 (N136, N135, N114, N106, N124);
xor XOR2 (N137, N111, N110);
nand NAND2 (N138, N121, N104);
xor XOR2 (N139, N128, N119);
xor XOR2 (N140, N136, N119);
not NOT1 (N141, N133);
nor NOR2 (N142, N141, N96);
nand NAND3 (N143, N140, N48, N14);
or OR4 (N144, N130, N118, N89, N112);
xor XOR2 (N145, N143, N13);
buf BUF1 (N146, N142);
nand NAND4 (N147, N126, N29, N105, N31);
nand NAND3 (N148, N139, N14, N68);
buf BUF1 (N149, N144);
buf BUF1 (N150, N78);
and AND3 (N151, N123, N42, N75);
or OR3 (N152, N151, N58, N88);
and AND4 (N153, N137, N54, N30, N47);
not NOT1 (N154, N152);
nand NAND4 (N155, N138, N36, N102, N66);
xor XOR2 (N156, N150, N114);
xor XOR2 (N157, N156, N108);
buf BUF1 (N158, N148);
nand NAND2 (N159, N147, N42);
nand NAND3 (N160, N157, N42, N24);
nand NAND2 (N161, N131, N122);
buf BUF1 (N162, N154);
xor XOR2 (N163, N158, N128);
not NOT1 (N164, N153);
or OR4 (N165, N149, N84, N15, N10);
xor XOR2 (N166, N159, N158);
xor XOR2 (N167, N155, N52);
or OR4 (N168, N160, N86, N98, N149);
not NOT1 (N169, N165);
and AND4 (N170, N166, N83, N94, N138);
and AND4 (N171, N170, N91, N135, N91);
nand NAND3 (N172, N145, N53, N125);
and AND2 (N173, N164, N72);
or OR4 (N174, N172, N164, N36, N111);
xor XOR2 (N175, N162, N169);
buf BUF1 (N176, N119);
nor NOR2 (N177, N174, N159);
not NOT1 (N178, N171);
nand NAND4 (N179, N173, N2, N110, N159);
and AND2 (N180, N146, N59);
not NOT1 (N181, N180);
xor XOR2 (N182, N178, N11);
nand NAND4 (N183, N179, N68, N52, N133);
or OR4 (N184, N168, N17, N158, N150);
not NOT1 (N185, N184);
nor NOR3 (N186, N177, N5, N157);
xor XOR2 (N187, N186, N105);
buf BUF1 (N188, N163);
or OR4 (N189, N175, N94, N183, N133);
not NOT1 (N190, N117);
and AND3 (N191, N176, N123, N24);
not NOT1 (N192, N161);
buf BUF1 (N193, N187);
or OR3 (N194, N182, N178, N6);
nor NOR3 (N195, N193, N119, N55);
and AND2 (N196, N167, N27);
nand NAND2 (N197, N194, N135);
nor NOR3 (N198, N197, N197, N37);
nand NAND4 (N199, N181, N58, N105, N103);
nor NOR3 (N200, N196, N121, N198);
or OR4 (N201, N52, N43, N69, N36);
buf BUF1 (N202, N189);
not NOT1 (N203, N199);
nand NAND4 (N204, N195, N72, N89, N164);
not NOT1 (N205, N190);
xor XOR2 (N206, N192, N29);
and AND4 (N207, N203, N197, N205, N73);
not NOT1 (N208, N185);
not NOT1 (N209, N58);
or OR4 (N210, N206, N185, N88, N165);
buf BUF1 (N211, N210);
buf BUF1 (N212, N191);
or OR2 (N213, N208, N194);
not NOT1 (N214, N202);
or OR3 (N215, N211, N154, N206);
nor NOR4 (N216, N214, N22, N93, N133);
nand NAND3 (N217, N188, N128, N63);
nor NOR4 (N218, N213, N154, N152, N68);
and AND4 (N219, N201, N14, N202, N161);
nand NAND2 (N220, N209, N91);
endmodule