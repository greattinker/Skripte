// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23;

output N8021,N8008,N8020,N8017,N8010,N8002,N8014,N7963,N8015,N8023;

nand NAND3 (N24, N1, N23, N16);
nand NAND2 (N25, N12, N19);
or OR3 (N26, N25, N5, N13);
nand NAND4 (N27, N26, N10, N2, N18);
buf BUF1 (N28, N26);
nor NOR4 (N29, N5, N28, N25, N22);
xor XOR2 (N30, N12, N2);
buf BUF1 (N31, N4);
buf BUF1 (N32, N3);
nand NAND3 (N33, N10, N17, N12);
and AND2 (N34, N26, N23);
xor XOR2 (N35, N16, N17);
not NOT1 (N36, N6);
buf BUF1 (N37, N30);
and AND3 (N38, N34, N31, N10);
or OR3 (N39, N33, N8, N30);
buf BUF1 (N40, N27);
and AND3 (N41, N10, N23, N3);
xor XOR2 (N42, N24, N6);
nand NAND3 (N43, N40, N41, N25);
xor XOR2 (N44, N26, N8);
nand NAND2 (N45, N36, N2);
buf BUF1 (N46, N35);
not NOT1 (N47, N29);
not NOT1 (N48, N32);
or OR4 (N49, N38, N1, N32, N19);
xor XOR2 (N50, N37, N40);
xor XOR2 (N51, N45, N43);
nor NOR3 (N52, N37, N34, N41);
nand NAND2 (N53, N42, N10);
xor XOR2 (N54, N48, N31);
or OR2 (N55, N54, N31);
nor NOR4 (N56, N53, N18, N34, N25);
nand NAND3 (N57, N44, N52, N47);
nand NAND2 (N58, N40, N43);
buf BUF1 (N59, N36);
nand NAND4 (N60, N46, N21, N34, N28);
not NOT1 (N61, N59);
xor XOR2 (N62, N49, N51);
xor XOR2 (N63, N45, N27);
or OR2 (N64, N55, N15);
or OR3 (N65, N60, N50, N9);
and AND2 (N66, N3, N44);
buf BUF1 (N67, N56);
buf BUF1 (N68, N66);
nor NOR4 (N69, N58, N33, N43, N57);
nand NAND3 (N70, N31, N7, N18);
nor NOR3 (N71, N65, N7, N55);
xor XOR2 (N72, N62, N62);
nor NOR2 (N73, N64, N34);
not NOT1 (N74, N72);
nand NAND3 (N75, N73, N45, N51);
or OR4 (N76, N71, N15, N47, N54);
buf BUF1 (N77, N76);
nor NOR3 (N78, N63, N28, N44);
or OR4 (N79, N74, N3, N52, N61);
nand NAND3 (N80, N22, N7, N9);
not NOT1 (N81, N75);
buf BUF1 (N82, N77);
buf BUF1 (N83, N80);
buf BUF1 (N84, N68);
or OR2 (N85, N83, N67);
nand NAND3 (N86, N35, N63, N36);
or OR3 (N87, N85, N26, N5);
not NOT1 (N88, N79);
xor XOR2 (N89, N82, N22);
buf BUF1 (N90, N89);
xor XOR2 (N91, N39, N42);
buf BUF1 (N92, N81);
not NOT1 (N93, N88);
not NOT1 (N94, N86);
buf BUF1 (N95, N70);
or OR2 (N96, N91, N44);
xor XOR2 (N97, N87, N41);
not NOT1 (N98, N90);
and AND4 (N99, N94, N50, N5, N95);
not NOT1 (N100, N17);
or OR2 (N101, N99, N6);
buf BUF1 (N102, N96);
not NOT1 (N103, N101);
xor XOR2 (N104, N100, N74);
or OR2 (N105, N93, N11);
not NOT1 (N106, N102);
or OR4 (N107, N103, N17, N1, N102);
or OR4 (N108, N107, N40, N75, N73);
nand NAND4 (N109, N92, N91, N4, N29);
nor NOR3 (N110, N109, N85, N32);
buf BUF1 (N111, N104);
or OR3 (N112, N98, N42, N62);
nor NOR4 (N113, N69, N29, N41, N27);
xor XOR2 (N114, N97, N95);
nor NOR4 (N115, N114, N95, N92, N89);
or OR2 (N116, N78, N66);
buf BUF1 (N117, N111);
xor XOR2 (N118, N115, N45);
nor NOR3 (N119, N116, N27, N18);
buf BUF1 (N120, N112);
not NOT1 (N121, N118);
nor NOR3 (N122, N121, N51, N23);
nor NOR4 (N123, N122, N100, N103, N35);
not NOT1 (N124, N110);
nand NAND4 (N125, N113, N61, N29, N35);
not NOT1 (N126, N106);
and AND2 (N127, N105, N63);
nand NAND4 (N128, N125, N70, N59, N24);
xor XOR2 (N129, N108, N69);
buf BUF1 (N130, N119);
and AND3 (N131, N120, N103, N51);
buf BUF1 (N132, N131);
and AND3 (N133, N126, N103, N92);
xor XOR2 (N134, N130, N121);
nor NOR4 (N135, N124, N75, N16, N123);
and AND3 (N136, N32, N47, N84);
nor NOR4 (N137, N135, N92, N37, N135);
or OR3 (N138, N74, N24, N56);
or OR2 (N139, N128, N44);
not NOT1 (N140, N129);
xor XOR2 (N141, N117, N138);
nor NOR3 (N142, N32, N115, N99);
nand NAND4 (N143, N140, N46, N120, N60);
xor XOR2 (N144, N133, N62);
not NOT1 (N145, N141);
or OR3 (N146, N143, N51, N125);
and AND4 (N147, N137, N101, N51, N136);
nor NOR2 (N148, N110, N111);
xor XOR2 (N149, N142, N9);
nor NOR4 (N150, N144, N39, N59, N71);
xor XOR2 (N151, N148, N7);
buf BUF1 (N152, N139);
buf BUF1 (N153, N149);
and AND4 (N154, N145, N85, N97, N92);
or OR2 (N155, N151, N67);
and AND2 (N156, N153, N102);
not NOT1 (N157, N152);
and AND3 (N158, N127, N86, N51);
nand NAND4 (N159, N154, N76, N131, N16);
nor NOR2 (N160, N159, N25);
and AND3 (N161, N158, N109, N53);
and AND2 (N162, N157, N97);
buf BUF1 (N163, N146);
buf BUF1 (N164, N160);
xor XOR2 (N165, N147, N159);
and AND2 (N166, N155, N161);
and AND2 (N167, N74, N4);
and AND3 (N168, N165, N73, N161);
xor XOR2 (N169, N150, N54);
nor NOR2 (N170, N132, N9);
nand NAND2 (N171, N169, N70);
or OR3 (N172, N162, N151, N48);
buf BUF1 (N173, N172);
nand NAND2 (N174, N156, N85);
buf BUF1 (N175, N164);
xor XOR2 (N176, N167, N146);
nor NOR3 (N177, N174, N171, N35);
and AND3 (N178, N152, N160, N60);
nand NAND3 (N179, N173, N11, N28);
not NOT1 (N180, N179);
xor XOR2 (N181, N134, N142);
and AND2 (N182, N176, N52);
nor NOR2 (N183, N170, N52);
not NOT1 (N184, N177);
or OR4 (N185, N168, N151, N175, N162);
nor NOR3 (N186, N153, N137, N15);
buf BUF1 (N187, N185);
nor NOR2 (N188, N163, N18);
or OR4 (N189, N166, N130, N30, N4);
xor XOR2 (N190, N180, N103);
nor NOR3 (N191, N184, N177, N176);
not NOT1 (N192, N187);
xor XOR2 (N193, N181, N22);
not NOT1 (N194, N186);
xor XOR2 (N195, N192, N181);
buf BUF1 (N196, N182);
not NOT1 (N197, N195);
nor NOR3 (N198, N189, N20, N64);
nor NOR4 (N199, N194, N88, N180, N65);
xor XOR2 (N200, N199, N53);
not NOT1 (N201, N200);
and AND4 (N202, N178, N79, N102, N74);
nand NAND2 (N203, N193, N148);
xor XOR2 (N204, N198, N88);
not NOT1 (N205, N191);
and AND4 (N206, N204, N144, N62, N27);
nor NOR4 (N207, N188, N89, N188, N67);
not NOT1 (N208, N201);
nor NOR3 (N209, N205, N171, N23);
nor NOR4 (N210, N190, N89, N25, N191);
and AND2 (N211, N207, N41);
and AND3 (N212, N210, N89, N208);
buf BUF1 (N213, N83);
nor NOR3 (N214, N212, N199, N99);
not NOT1 (N215, N213);
or OR2 (N216, N197, N96);
or OR4 (N217, N203, N21, N174, N74);
and AND2 (N218, N209, N203);
buf BUF1 (N219, N214);
nand NAND4 (N220, N183, N45, N29, N111);
or OR3 (N221, N211, N59, N109);
xor XOR2 (N222, N216, N108);
not NOT1 (N223, N222);
xor XOR2 (N224, N218, N125);
nor NOR3 (N225, N196, N85, N118);
and AND2 (N226, N223, N105);
buf BUF1 (N227, N221);
and AND2 (N228, N217, N10);
buf BUF1 (N229, N202);
nor NOR2 (N230, N220, N31);
not NOT1 (N231, N225);
or OR2 (N232, N224, N230);
buf BUF1 (N233, N90);
nor NOR3 (N234, N215, N78, N44);
xor XOR2 (N235, N228, N163);
and AND2 (N236, N232, N103);
nor NOR2 (N237, N235, N123);
or OR2 (N238, N237, N124);
buf BUF1 (N239, N206);
buf BUF1 (N240, N219);
and AND3 (N241, N226, N171, N115);
and AND2 (N242, N236, N67);
nor NOR4 (N243, N229, N82, N168, N34);
or OR2 (N244, N227, N165);
and AND2 (N245, N243, N37);
and AND2 (N246, N238, N9);
not NOT1 (N247, N233);
and AND4 (N248, N241, N120, N247, N142);
nor NOR4 (N249, N175, N134, N121, N63);
and AND4 (N250, N240, N177, N71, N60);
nor NOR4 (N251, N239, N190, N131, N162);
or OR4 (N252, N234, N28, N204, N87);
nand NAND4 (N253, N250, N9, N85, N16);
buf BUF1 (N254, N251);
nand NAND4 (N255, N254, N190, N106, N222);
nor NOR3 (N256, N242, N72, N149);
not NOT1 (N257, N249);
and AND3 (N258, N231, N223, N55);
nor NOR3 (N259, N258, N248, N125);
nor NOR3 (N260, N76, N8, N180);
and AND4 (N261, N257, N37, N158, N250);
nor NOR4 (N262, N253, N248, N116, N105);
nor NOR4 (N263, N255, N260, N65, N3);
not NOT1 (N264, N166);
and AND4 (N265, N245, N114, N83, N25);
buf BUF1 (N266, N262);
nand NAND3 (N267, N264, N191, N244);
or OR3 (N268, N257, N2, N238);
buf BUF1 (N269, N252);
not NOT1 (N270, N263);
not NOT1 (N271, N261);
or OR3 (N272, N271, N72, N120);
or OR3 (N273, N270, N198, N130);
buf BUF1 (N274, N273);
xor XOR2 (N275, N272, N236);
buf BUF1 (N276, N246);
or OR4 (N277, N256, N124, N147, N79);
nand NAND2 (N278, N259, N19);
nor NOR3 (N279, N268, N247, N59);
xor XOR2 (N280, N275, N75);
or OR4 (N281, N274, N112, N136, N77);
buf BUF1 (N282, N265);
nand NAND4 (N283, N279, N245, N122, N45);
buf BUF1 (N284, N280);
not NOT1 (N285, N284);
or OR2 (N286, N269, N57);
nand NAND2 (N287, N266, N272);
nand NAND2 (N288, N283, N51);
or OR4 (N289, N281, N90, N186, N259);
xor XOR2 (N290, N276, N145);
buf BUF1 (N291, N288);
nor NOR3 (N292, N287, N39, N161);
or OR3 (N293, N282, N133, N116);
not NOT1 (N294, N285);
nand NAND3 (N295, N290, N48, N202);
nand NAND3 (N296, N289, N69, N160);
buf BUF1 (N297, N278);
and AND4 (N298, N291, N129, N207, N222);
or OR2 (N299, N296, N118);
xor XOR2 (N300, N297, N127);
buf BUF1 (N301, N293);
nor NOR2 (N302, N267, N298);
nor NOR2 (N303, N106, N58);
nor NOR2 (N304, N301, N51);
nor NOR4 (N305, N300, N281, N35, N81);
xor XOR2 (N306, N277, N4);
xor XOR2 (N307, N304, N185);
buf BUF1 (N308, N295);
nor NOR2 (N309, N303, N189);
nand NAND2 (N310, N306, N137);
or OR4 (N311, N307, N84, N278, N69);
not NOT1 (N312, N309);
buf BUF1 (N313, N308);
buf BUF1 (N314, N310);
xor XOR2 (N315, N292, N97);
xor XOR2 (N316, N314, N225);
or OR2 (N317, N286, N173);
or OR2 (N318, N311, N107);
nand NAND4 (N319, N317, N264, N267, N202);
xor XOR2 (N320, N315, N261);
buf BUF1 (N321, N312);
xor XOR2 (N322, N302, N275);
buf BUF1 (N323, N321);
not NOT1 (N324, N318);
and AND3 (N325, N320, N219, N282);
nor NOR2 (N326, N319, N76);
xor XOR2 (N327, N326, N283);
nand NAND4 (N328, N305, N178, N33, N176);
nor NOR4 (N329, N324, N232, N278, N125);
not NOT1 (N330, N323);
not NOT1 (N331, N325);
and AND4 (N332, N330, N92, N8, N281);
buf BUF1 (N333, N294);
nor NOR4 (N334, N316, N275, N65, N159);
and AND2 (N335, N299, N267);
and AND4 (N336, N327, N213, N202, N281);
buf BUF1 (N337, N335);
nor NOR2 (N338, N333, N189);
not NOT1 (N339, N332);
not NOT1 (N340, N328);
xor XOR2 (N341, N322, N172);
buf BUF1 (N342, N338);
nor NOR3 (N343, N342, N225, N171);
or OR4 (N344, N336, N207, N211, N217);
nor NOR4 (N345, N339, N309, N17, N170);
buf BUF1 (N346, N341);
and AND4 (N347, N334, N61, N273, N280);
not NOT1 (N348, N347);
or OR2 (N349, N331, N68);
nor NOR3 (N350, N344, N140, N213);
not NOT1 (N351, N345);
nor NOR3 (N352, N346, N201, N23);
nor NOR3 (N353, N348, N251, N31);
or OR3 (N354, N352, N115, N4);
nand NAND2 (N355, N351, N339);
nand NAND3 (N356, N355, N194, N338);
or OR3 (N357, N356, N276, N154);
buf BUF1 (N358, N340);
nand NAND3 (N359, N337, N174, N210);
buf BUF1 (N360, N358);
or OR2 (N361, N357, N225);
buf BUF1 (N362, N360);
nor NOR3 (N363, N362, N347, N204);
nor NOR2 (N364, N361, N254);
nand NAND4 (N365, N353, N37, N168, N158);
nand NAND3 (N366, N313, N269, N138);
and AND4 (N367, N349, N90, N79, N245);
nor NOR4 (N368, N329, N25, N348, N121);
or OR3 (N369, N364, N328, N35);
not NOT1 (N370, N359);
not NOT1 (N371, N369);
and AND4 (N372, N350, N249, N138, N339);
nand NAND4 (N373, N367, N236, N124, N240);
not NOT1 (N374, N368);
and AND3 (N375, N363, N273, N21);
not NOT1 (N376, N371);
nor NOR2 (N377, N376, N113);
nand NAND3 (N378, N365, N62, N37);
buf BUF1 (N379, N354);
or OR2 (N380, N343, N229);
not NOT1 (N381, N379);
nor NOR2 (N382, N370, N184);
xor XOR2 (N383, N380, N298);
nand NAND4 (N384, N377, N81, N338, N43);
or OR3 (N385, N382, N145, N281);
nand NAND3 (N386, N366, N68, N134);
nor NOR2 (N387, N375, N379);
or OR2 (N388, N378, N31);
and AND4 (N389, N384, N24, N380, N72);
nor NOR2 (N390, N385, N82);
buf BUF1 (N391, N389);
xor XOR2 (N392, N373, N145);
xor XOR2 (N393, N388, N51);
nand NAND4 (N394, N391, N88, N378, N324);
nor NOR3 (N395, N374, N388, N267);
not NOT1 (N396, N394);
or OR2 (N397, N372, N62);
and AND4 (N398, N381, N102, N319, N241);
buf BUF1 (N399, N392);
nand NAND3 (N400, N383, N147, N338);
or OR4 (N401, N395, N270, N220, N132);
xor XOR2 (N402, N393, N194);
or OR2 (N403, N401, N134);
and AND3 (N404, N400, N263, N298);
nor NOR4 (N405, N398, N397, N28, N280);
buf BUF1 (N406, N342);
nand NAND3 (N407, N406, N92, N62);
or OR4 (N408, N390, N43, N377, N48);
nand NAND4 (N409, N403, N300, N116, N74);
nor NOR3 (N410, N396, N311, N41);
or OR3 (N411, N408, N1, N38);
xor XOR2 (N412, N405, N287);
nor NOR4 (N413, N407, N276, N150, N344);
or OR4 (N414, N410, N149, N175, N122);
and AND2 (N415, N409, N255);
and AND2 (N416, N399, N260);
nand NAND4 (N417, N413, N23, N272, N24);
nand NAND2 (N418, N415, N69);
not NOT1 (N419, N417);
xor XOR2 (N420, N387, N364);
and AND2 (N421, N414, N239);
xor XOR2 (N422, N418, N318);
nand NAND4 (N423, N412, N91, N314, N237);
or OR2 (N424, N423, N342);
buf BUF1 (N425, N386);
and AND4 (N426, N419, N81, N158, N77);
and AND3 (N427, N402, N150, N142);
nor NOR4 (N428, N420, N398, N94, N9);
or OR3 (N429, N416, N211, N121);
not NOT1 (N430, N421);
nand NAND3 (N431, N427, N411, N42);
nor NOR2 (N432, N56, N118);
not NOT1 (N433, N422);
and AND3 (N434, N430, N279, N343);
and AND2 (N435, N425, N264);
or OR2 (N436, N426, N60);
buf BUF1 (N437, N432);
nand NAND4 (N438, N424, N147, N128, N71);
or OR3 (N439, N438, N288, N237);
buf BUF1 (N440, N428);
nor NOR2 (N441, N440, N316);
xor XOR2 (N442, N436, N68);
nor NOR4 (N443, N442, N176, N321, N174);
and AND3 (N444, N439, N244, N330);
not NOT1 (N445, N435);
nand NAND3 (N446, N433, N411, N316);
not NOT1 (N447, N441);
or OR3 (N448, N404, N440, N19);
buf BUF1 (N449, N446);
not NOT1 (N450, N448);
nor NOR2 (N451, N445, N211);
and AND4 (N452, N450, N28, N357, N253);
not NOT1 (N453, N447);
xor XOR2 (N454, N449, N70);
not NOT1 (N455, N434);
xor XOR2 (N456, N454, N442);
and AND3 (N457, N444, N446, N206);
nand NAND2 (N458, N437, N323);
nand NAND2 (N459, N456, N296);
not NOT1 (N460, N443);
not NOT1 (N461, N451);
or OR2 (N462, N459, N291);
xor XOR2 (N463, N431, N145);
and AND3 (N464, N462, N377, N55);
xor XOR2 (N465, N452, N346);
nor NOR3 (N466, N460, N108, N290);
buf BUF1 (N467, N457);
and AND4 (N468, N466, N300, N54, N82);
or OR4 (N469, N458, N37, N384, N315);
and AND3 (N470, N467, N243, N337);
and AND2 (N471, N468, N293);
buf BUF1 (N472, N461);
xor XOR2 (N473, N429, N341);
xor XOR2 (N474, N465, N385);
not NOT1 (N475, N464);
and AND2 (N476, N470, N387);
or OR2 (N477, N476, N378);
xor XOR2 (N478, N455, N47);
xor XOR2 (N479, N473, N400);
nand NAND3 (N480, N471, N326, N161);
nand NAND2 (N481, N475, N148);
nor NOR2 (N482, N472, N320);
nand NAND2 (N483, N477, N437);
nor NOR4 (N484, N482, N471, N301, N457);
or OR4 (N485, N478, N117, N459, N436);
not NOT1 (N486, N469);
nor NOR3 (N487, N486, N418, N382);
and AND2 (N488, N479, N209);
nor NOR4 (N489, N453, N473, N171, N202);
buf BUF1 (N490, N488);
not NOT1 (N491, N481);
nor NOR3 (N492, N490, N360, N480);
or OR4 (N493, N453, N352, N470, N84);
or OR3 (N494, N492, N300, N412);
nand NAND3 (N495, N474, N383, N342);
nor NOR3 (N496, N495, N383, N198);
not NOT1 (N497, N463);
xor XOR2 (N498, N496, N270);
buf BUF1 (N499, N487);
and AND2 (N500, N498, N282);
xor XOR2 (N501, N493, N399);
buf BUF1 (N502, N499);
buf BUF1 (N503, N489);
nor NOR3 (N504, N502, N426, N173);
or OR2 (N505, N497, N52);
nand NAND2 (N506, N491, N71);
buf BUF1 (N507, N500);
buf BUF1 (N508, N501);
or OR2 (N509, N505, N131);
or OR3 (N510, N504, N386, N68);
xor XOR2 (N511, N485, N111);
or OR3 (N512, N507, N289, N221);
nand NAND3 (N513, N506, N498, N122);
buf BUF1 (N514, N483);
nand NAND4 (N515, N484, N332, N308, N147);
buf BUF1 (N516, N511);
xor XOR2 (N517, N510, N339);
xor XOR2 (N518, N508, N178);
not NOT1 (N519, N503);
not NOT1 (N520, N516);
or OR2 (N521, N494, N281);
nand NAND3 (N522, N518, N241, N251);
and AND3 (N523, N512, N63, N119);
nor NOR2 (N524, N517, N503);
nand NAND3 (N525, N519, N22, N316);
nor NOR3 (N526, N520, N186, N206);
buf BUF1 (N527, N524);
nor NOR3 (N528, N525, N146, N122);
not NOT1 (N529, N522);
buf BUF1 (N530, N513);
and AND3 (N531, N526, N231, N100);
and AND4 (N532, N529, N306, N306, N43);
buf BUF1 (N533, N530);
or OR2 (N534, N515, N143);
nand NAND4 (N535, N527, N5, N512, N260);
and AND2 (N536, N521, N39);
buf BUF1 (N537, N523);
nor NOR4 (N538, N536, N231, N406, N499);
or OR3 (N539, N531, N389, N447);
buf BUF1 (N540, N533);
nand NAND4 (N541, N535, N301, N391, N259);
nor NOR4 (N542, N539, N361, N250, N250);
nor NOR3 (N543, N532, N360, N166);
xor XOR2 (N544, N537, N434);
and AND3 (N545, N509, N410, N535);
and AND4 (N546, N542, N423, N347, N270);
or OR4 (N547, N528, N424, N518, N480);
xor XOR2 (N548, N543, N257);
nand NAND2 (N549, N514, N253);
and AND4 (N550, N547, N193, N64, N518);
nand NAND3 (N551, N549, N399, N306);
nand NAND3 (N552, N548, N478, N125);
nand NAND4 (N553, N540, N462, N65, N325);
nor NOR2 (N554, N544, N310);
nand NAND4 (N555, N546, N370, N94, N85);
buf BUF1 (N556, N550);
xor XOR2 (N557, N553, N299);
xor XOR2 (N558, N557, N387);
not NOT1 (N559, N545);
nand NAND2 (N560, N541, N204);
or OR2 (N561, N556, N67);
nor NOR3 (N562, N538, N556, N64);
not NOT1 (N563, N552);
nand NAND2 (N564, N554, N164);
nand NAND4 (N565, N563, N349, N493, N492);
not NOT1 (N566, N562);
xor XOR2 (N567, N565, N86);
nor NOR3 (N568, N551, N70, N200);
nor NOR3 (N569, N567, N340, N362);
buf BUF1 (N570, N566);
nor NOR3 (N571, N555, N110, N358);
and AND4 (N572, N560, N55, N43, N287);
and AND3 (N573, N561, N476, N483);
or OR3 (N574, N570, N14, N117);
and AND2 (N575, N564, N125);
buf BUF1 (N576, N573);
or OR3 (N577, N571, N433, N183);
and AND4 (N578, N559, N13, N436, N192);
or OR3 (N579, N558, N373, N79);
buf BUF1 (N580, N569);
nand NAND4 (N581, N572, N251, N272, N33);
nor NOR3 (N582, N577, N182, N251);
and AND2 (N583, N576, N208);
xor XOR2 (N584, N574, N195);
or OR3 (N585, N582, N231, N228);
not NOT1 (N586, N584);
or OR2 (N587, N575, N320);
and AND3 (N588, N579, N554, N434);
buf BUF1 (N589, N587);
nand NAND2 (N590, N578, N163);
nor NOR3 (N591, N581, N41, N515);
nand NAND3 (N592, N585, N327, N32);
nand NAND4 (N593, N592, N120, N130, N439);
or OR2 (N594, N568, N374);
buf BUF1 (N595, N586);
nand NAND2 (N596, N590, N347);
and AND4 (N597, N534, N138, N27, N563);
nand NAND2 (N598, N591, N451);
or OR3 (N599, N588, N335, N470);
or OR4 (N600, N597, N423, N522, N502);
nor NOR3 (N601, N600, N367, N440);
or OR2 (N602, N598, N298);
nand NAND2 (N603, N593, N72);
not NOT1 (N604, N589);
xor XOR2 (N605, N580, N45);
buf BUF1 (N606, N595);
xor XOR2 (N607, N594, N137);
not NOT1 (N608, N607);
and AND2 (N609, N606, N336);
buf BUF1 (N610, N605);
nand NAND3 (N611, N603, N233, N276);
or OR4 (N612, N608, N491, N455, N415);
nand NAND4 (N613, N611, N462, N206, N127);
buf BUF1 (N614, N596);
not NOT1 (N615, N610);
nor NOR2 (N616, N612, N103);
nor NOR3 (N617, N602, N380, N616);
xor XOR2 (N618, N126, N273);
and AND4 (N619, N583, N32, N401, N358);
nand NAND4 (N620, N618, N560, N239, N136);
xor XOR2 (N621, N613, N605);
and AND3 (N622, N614, N24, N209);
or OR3 (N623, N604, N105, N126);
nor NOR4 (N624, N621, N153, N298, N276);
and AND3 (N625, N624, N74, N71);
nor NOR2 (N626, N609, N326);
nor NOR2 (N627, N623, N541);
or OR3 (N628, N617, N152, N621);
buf BUF1 (N629, N599);
buf BUF1 (N630, N615);
nor NOR4 (N631, N622, N157, N527, N268);
xor XOR2 (N632, N625, N589);
nor NOR2 (N633, N632, N596);
nand NAND3 (N634, N619, N228, N548);
buf BUF1 (N635, N631);
or OR4 (N636, N626, N118, N510, N204);
nand NAND2 (N637, N635, N5);
and AND2 (N638, N630, N197);
and AND3 (N639, N629, N123, N634);
nand NAND2 (N640, N130, N96);
and AND4 (N641, N620, N416, N332, N547);
and AND4 (N642, N639, N481, N626, N290);
buf BUF1 (N643, N642);
xor XOR2 (N644, N643, N72);
nand NAND2 (N645, N636, N142);
nand NAND2 (N646, N633, N122);
xor XOR2 (N647, N640, N551);
nand NAND4 (N648, N644, N339, N485, N448);
buf BUF1 (N649, N637);
nor NOR4 (N650, N648, N501, N388, N282);
not NOT1 (N651, N646);
buf BUF1 (N652, N647);
not NOT1 (N653, N628);
xor XOR2 (N654, N641, N473);
buf BUF1 (N655, N645);
nor NOR3 (N656, N654, N422, N409);
nor NOR3 (N657, N601, N393, N184);
or OR2 (N658, N657, N284);
not NOT1 (N659, N652);
and AND4 (N660, N638, N287, N113, N260);
not NOT1 (N661, N627);
or OR2 (N662, N651, N110);
not NOT1 (N663, N656);
nand NAND3 (N664, N655, N408, N207);
nor NOR3 (N665, N664, N435, N93);
nand NAND2 (N666, N662, N274);
nand NAND2 (N667, N650, N465);
nor NOR2 (N668, N659, N615);
nor NOR2 (N669, N658, N233);
nand NAND4 (N670, N661, N360, N292, N92);
or OR3 (N671, N669, N341, N21);
not NOT1 (N672, N670);
nor NOR4 (N673, N668, N117, N570, N479);
nand NAND4 (N674, N666, N604, N260, N212);
not NOT1 (N675, N660);
nand NAND3 (N676, N673, N340, N607);
nand NAND3 (N677, N672, N346, N356);
buf BUF1 (N678, N667);
buf BUF1 (N679, N676);
or OR3 (N680, N653, N104, N252);
nor NOR2 (N681, N665, N31);
not NOT1 (N682, N671);
nor NOR4 (N683, N680, N21, N266, N660);
not NOT1 (N684, N649);
nand NAND3 (N685, N682, N489, N278);
and AND3 (N686, N678, N617, N457);
buf BUF1 (N687, N681);
buf BUF1 (N688, N683);
and AND3 (N689, N684, N221, N287);
and AND4 (N690, N689, N250, N82, N234);
buf BUF1 (N691, N679);
or OR2 (N692, N687, N235);
buf BUF1 (N693, N691);
and AND2 (N694, N677, N332);
xor XOR2 (N695, N694, N68);
buf BUF1 (N696, N695);
nor NOR2 (N697, N675, N695);
not NOT1 (N698, N696);
buf BUF1 (N699, N698);
buf BUF1 (N700, N693);
buf BUF1 (N701, N697);
xor XOR2 (N702, N699, N8);
nand NAND3 (N703, N692, N405, N25);
and AND3 (N704, N674, N515, N679);
nor NOR3 (N705, N703, N120, N190);
not NOT1 (N706, N705);
or OR2 (N707, N663, N86);
nor NOR4 (N708, N685, N629, N700, N377);
buf BUF1 (N709, N433);
nor NOR2 (N710, N709, N157);
or OR4 (N711, N688, N378, N106, N220);
nand NAND2 (N712, N686, N323);
xor XOR2 (N713, N701, N466);
or OR4 (N714, N712, N130, N555, N498);
nand NAND2 (N715, N713, N399);
not NOT1 (N716, N690);
or OR4 (N717, N715, N261, N576, N448);
or OR4 (N718, N702, N396, N216, N303);
nand NAND2 (N719, N717, N191);
not NOT1 (N720, N716);
not NOT1 (N721, N714);
nor NOR3 (N722, N711, N421, N92);
nor NOR4 (N723, N722, N179, N695, N79);
and AND3 (N724, N710, N254, N596);
nand NAND2 (N725, N718, N12);
not NOT1 (N726, N708);
xor XOR2 (N727, N725, N98);
and AND4 (N728, N723, N641, N634, N116);
or OR3 (N729, N721, N278, N212);
xor XOR2 (N730, N727, N140);
xor XOR2 (N731, N704, N72);
not NOT1 (N732, N720);
or OR4 (N733, N706, N264, N59, N180);
nor NOR4 (N734, N731, N472, N387, N431);
or OR2 (N735, N707, N350);
nor NOR3 (N736, N732, N296, N589);
not NOT1 (N737, N724);
nand NAND3 (N738, N735, N176, N405);
xor XOR2 (N739, N728, N477);
not NOT1 (N740, N734);
nand NAND2 (N741, N737, N685);
not NOT1 (N742, N730);
nand NAND4 (N743, N739, N334, N637, N464);
not NOT1 (N744, N736);
not NOT1 (N745, N719);
nand NAND4 (N746, N729, N733, N522, N731);
not NOT1 (N747, N575);
or OR3 (N748, N742, N741, N694);
or OR3 (N749, N492, N261, N582);
nor NOR4 (N750, N726, N736, N101, N100);
nor NOR4 (N751, N743, N302, N449, N84);
not NOT1 (N752, N738);
xor XOR2 (N753, N747, N731);
or OR2 (N754, N745, N322);
or OR3 (N755, N754, N748, N594);
buf BUF1 (N756, N731);
nor NOR2 (N757, N755, N575);
nor NOR2 (N758, N751, N401);
nor NOR2 (N759, N749, N464);
and AND2 (N760, N752, N414);
nand NAND2 (N761, N744, N658);
buf BUF1 (N762, N759);
buf BUF1 (N763, N756);
nand NAND4 (N764, N757, N136, N307, N53);
or OR3 (N765, N753, N172, N6);
nor NOR4 (N766, N746, N122, N480, N526);
buf BUF1 (N767, N760);
nor NOR2 (N768, N767, N722);
and AND3 (N769, N761, N542, N617);
buf BUF1 (N770, N766);
buf BUF1 (N771, N762);
not NOT1 (N772, N770);
not NOT1 (N773, N765);
buf BUF1 (N774, N768);
or OR2 (N775, N774, N682);
and AND3 (N776, N775, N179, N454);
xor XOR2 (N777, N776, N295);
or OR4 (N778, N750, N214, N234, N727);
xor XOR2 (N779, N763, N361);
buf BUF1 (N780, N779);
buf BUF1 (N781, N771);
nor NOR2 (N782, N777, N549);
not NOT1 (N783, N773);
or OR2 (N784, N772, N20);
nand NAND3 (N785, N783, N137, N367);
xor XOR2 (N786, N782, N217);
not NOT1 (N787, N784);
nand NAND3 (N788, N780, N266, N129);
or OR2 (N789, N740, N362);
not NOT1 (N790, N764);
buf BUF1 (N791, N787);
nor NOR4 (N792, N785, N116, N638, N520);
and AND3 (N793, N778, N475, N738);
buf BUF1 (N794, N793);
and AND2 (N795, N788, N608);
nand NAND3 (N796, N758, N405, N513);
nor NOR3 (N797, N769, N791, N192);
or OR3 (N798, N738, N738, N740);
nand NAND4 (N799, N789, N658, N45, N228);
not NOT1 (N800, N798);
not NOT1 (N801, N800);
buf BUF1 (N802, N781);
not NOT1 (N803, N794);
or OR3 (N804, N803, N599, N686);
nand NAND3 (N805, N802, N773, N297);
nor NOR3 (N806, N796, N271, N659);
or OR2 (N807, N797, N583);
nor NOR4 (N808, N799, N233, N493, N263);
and AND3 (N809, N790, N414, N679);
nand NAND2 (N810, N808, N291);
or OR3 (N811, N801, N536, N325);
not NOT1 (N812, N795);
nor NOR4 (N813, N806, N486, N325, N478);
nor NOR4 (N814, N812, N390, N606, N117);
xor XOR2 (N815, N810, N373);
buf BUF1 (N816, N792);
or OR2 (N817, N809, N182);
nor NOR2 (N818, N805, N210);
buf BUF1 (N819, N807);
nor NOR3 (N820, N817, N239, N392);
nand NAND2 (N821, N815, N132);
nand NAND3 (N822, N804, N751, N309);
not NOT1 (N823, N822);
nor NOR3 (N824, N786, N484, N566);
not NOT1 (N825, N813);
nor NOR2 (N826, N811, N495);
not NOT1 (N827, N816);
and AND2 (N828, N824, N240);
and AND3 (N829, N828, N672, N423);
buf BUF1 (N830, N819);
nor NOR3 (N831, N818, N736, N531);
not NOT1 (N832, N829);
xor XOR2 (N833, N827, N188);
nand NAND2 (N834, N833, N515);
buf BUF1 (N835, N823);
or OR3 (N836, N820, N460, N192);
nand NAND3 (N837, N832, N587, N348);
buf BUF1 (N838, N837);
nor NOR3 (N839, N836, N248, N576);
and AND3 (N840, N826, N561, N140);
not NOT1 (N841, N835);
xor XOR2 (N842, N834, N15);
and AND2 (N843, N831, N138);
and AND2 (N844, N830, N313);
or OR4 (N845, N825, N311, N139, N247);
nand NAND2 (N846, N841, N102);
nand NAND2 (N847, N845, N691);
nand NAND2 (N848, N814, N782);
nor NOR2 (N849, N839, N34);
or OR3 (N850, N838, N419, N840);
and AND2 (N851, N342, N186);
nor NOR4 (N852, N844, N157, N259, N252);
and AND2 (N853, N848, N229);
xor XOR2 (N854, N842, N611);
nand NAND2 (N855, N846, N424);
xor XOR2 (N856, N851, N422);
nand NAND3 (N857, N849, N336, N350);
and AND3 (N858, N847, N826, N793);
nand NAND3 (N859, N856, N530, N434);
nor NOR3 (N860, N850, N675, N238);
xor XOR2 (N861, N859, N520);
not NOT1 (N862, N857);
or OR4 (N863, N854, N527, N265, N98);
nand NAND2 (N864, N853, N35);
and AND3 (N865, N863, N13, N44);
nand NAND2 (N866, N852, N753);
or OR2 (N867, N858, N1);
buf BUF1 (N868, N862);
xor XOR2 (N869, N866, N122);
buf BUF1 (N870, N864);
xor XOR2 (N871, N821, N123);
xor XOR2 (N872, N855, N77);
xor XOR2 (N873, N868, N71);
buf BUF1 (N874, N860);
or OR4 (N875, N843, N272, N131, N842);
nand NAND4 (N876, N861, N3, N98, N336);
buf BUF1 (N877, N874);
nand NAND2 (N878, N869, N90);
buf BUF1 (N879, N873);
xor XOR2 (N880, N865, N88);
and AND2 (N881, N879, N149);
nor NOR2 (N882, N877, N121);
xor XOR2 (N883, N870, N855);
xor XOR2 (N884, N883, N88);
and AND2 (N885, N880, N40);
buf BUF1 (N886, N882);
or OR3 (N887, N878, N122, N261);
or OR3 (N888, N887, N711, N325);
not NOT1 (N889, N884);
nor NOR2 (N890, N875, N369);
not NOT1 (N891, N889);
or OR3 (N892, N867, N888, N140);
xor XOR2 (N893, N531, N563);
and AND3 (N894, N872, N173, N539);
buf BUF1 (N895, N881);
or OR2 (N896, N892, N271);
nor NOR2 (N897, N895, N580);
buf BUF1 (N898, N894);
nand NAND3 (N899, N886, N711, N645);
nor NOR4 (N900, N885, N718, N231, N813);
not NOT1 (N901, N900);
not NOT1 (N902, N871);
nor NOR4 (N903, N891, N622, N237, N397);
and AND3 (N904, N898, N388, N655);
nor NOR2 (N905, N890, N162);
nor NOR2 (N906, N903, N17);
buf BUF1 (N907, N893);
not NOT1 (N908, N876);
nand NAND4 (N909, N901, N517, N745, N163);
nor NOR2 (N910, N908, N586);
not NOT1 (N911, N906);
buf BUF1 (N912, N911);
not NOT1 (N913, N902);
and AND4 (N914, N913, N129, N638, N151);
not NOT1 (N915, N905);
and AND4 (N916, N897, N79, N795, N283);
nor NOR4 (N917, N896, N17, N387, N527);
xor XOR2 (N918, N917, N42);
nor NOR3 (N919, N915, N849, N259);
nand NAND3 (N920, N899, N558, N691);
and AND2 (N921, N904, N476);
or OR2 (N922, N912, N673);
buf BUF1 (N923, N916);
nor NOR4 (N924, N918, N330, N892, N731);
nor NOR3 (N925, N921, N463, N722);
and AND2 (N926, N914, N476);
nand NAND3 (N927, N919, N719, N446);
nand NAND4 (N928, N923, N856, N424, N247);
nand NAND4 (N929, N927, N764, N723, N103);
xor XOR2 (N930, N920, N502);
nor NOR2 (N931, N926, N670);
buf BUF1 (N932, N928);
and AND4 (N933, N922, N416, N416, N162);
xor XOR2 (N934, N907, N51);
and AND3 (N935, N929, N130, N667);
or OR4 (N936, N925, N322, N444, N456);
nand NAND4 (N937, N934, N218, N208, N889);
not NOT1 (N938, N937);
or OR3 (N939, N936, N349, N438);
nor NOR2 (N940, N938, N171);
not NOT1 (N941, N909);
buf BUF1 (N942, N932);
or OR3 (N943, N941, N487, N530);
nor NOR3 (N944, N910, N478, N893);
or OR3 (N945, N939, N726, N256);
not NOT1 (N946, N930);
nand NAND2 (N947, N946, N272);
nand NAND3 (N948, N931, N584, N552);
nand NAND2 (N949, N940, N206);
nor NOR2 (N950, N949, N836);
nor NOR3 (N951, N950, N270, N359);
and AND3 (N952, N944, N589, N223);
or OR3 (N953, N945, N322, N231);
buf BUF1 (N954, N942);
or OR2 (N955, N947, N155);
buf BUF1 (N956, N935);
and AND4 (N957, N956, N723, N802, N660);
or OR3 (N958, N957, N67, N666);
buf BUF1 (N959, N952);
and AND4 (N960, N924, N652, N391, N697);
nand NAND2 (N961, N959, N344);
or OR3 (N962, N961, N665, N385);
buf BUF1 (N963, N960);
and AND2 (N964, N943, N124);
not NOT1 (N965, N954);
buf BUF1 (N966, N964);
not NOT1 (N967, N955);
or OR4 (N968, N948, N767, N792, N928);
buf BUF1 (N969, N962);
or OR2 (N970, N966, N921);
not NOT1 (N971, N965);
nand NAND4 (N972, N951, N184, N424, N235);
not NOT1 (N973, N958);
not NOT1 (N974, N963);
xor XOR2 (N975, N953, N556);
or OR3 (N976, N968, N889, N389);
nand NAND2 (N977, N975, N856);
xor XOR2 (N978, N933, N38);
nand NAND2 (N979, N977, N68);
not NOT1 (N980, N972);
buf BUF1 (N981, N978);
or OR4 (N982, N969, N76, N611, N386);
nand NAND3 (N983, N982, N942, N684);
buf BUF1 (N984, N971);
nand NAND4 (N985, N974, N805, N522, N863);
buf BUF1 (N986, N980);
nand NAND4 (N987, N983, N508, N656, N199);
buf BUF1 (N988, N987);
not NOT1 (N989, N970);
or OR3 (N990, N981, N901, N289);
nor NOR4 (N991, N976, N330, N253, N64);
or OR2 (N992, N991, N640);
or OR3 (N993, N985, N607, N445);
nor NOR2 (N994, N992, N344);
xor XOR2 (N995, N967, N224);
and AND3 (N996, N990, N617, N926);
nor NOR3 (N997, N988, N128, N214);
or OR3 (N998, N986, N526, N71);
xor XOR2 (N999, N996, N30);
not NOT1 (N1000, N973);
buf BUF1 (N1001, N995);
buf BUF1 (N1002, N1001);
xor XOR2 (N1003, N989, N342);
and AND4 (N1004, N1002, N11, N945, N442);
nor NOR4 (N1005, N984, N522, N779, N819);
buf BUF1 (N1006, N999);
xor XOR2 (N1007, N1000, N961);
buf BUF1 (N1008, N993);
nor NOR3 (N1009, N979, N445, N666);
or OR4 (N1010, N997, N360, N320, N848);
not NOT1 (N1011, N1009);
xor XOR2 (N1012, N1006, N837);
buf BUF1 (N1013, N1007);
xor XOR2 (N1014, N994, N416);
not NOT1 (N1015, N998);
or OR2 (N1016, N1004, N78);
nand NAND2 (N1017, N1012, N681);
nor NOR3 (N1018, N1008, N590, N724);
nand NAND2 (N1019, N1011, N165);
xor XOR2 (N1020, N1010, N136);
buf BUF1 (N1021, N1013);
and AND2 (N1022, N1003, N635);
xor XOR2 (N1023, N1022, N950);
buf BUF1 (N1024, N1005);
not NOT1 (N1025, N1020);
and AND4 (N1026, N1025, N165, N591, N47);
nand NAND4 (N1027, N1026, N229, N1003, N634);
and AND4 (N1028, N1017, N414, N301, N661);
buf BUF1 (N1029, N1015);
xor XOR2 (N1030, N1024, N985);
nor NOR4 (N1031, N1018, N85, N550, N28);
buf BUF1 (N1032, N1014);
nor NOR4 (N1033, N1029, N477, N633, N377);
buf BUF1 (N1034, N1033);
not NOT1 (N1035, N1016);
nand NAND2 (N1036, N1030, N81);
or OR2 (N1037, N1021, N652);
not NOT1 (N1038, N1031);
nor NOR4 (N1039, N1038, N815, N788, N842);
not NOT1 (N1040, N1039);
not NOT1 (N1041, N1036);
or OR4 (N1042, N1019, N649, N521, N412);
buf BUF1 (N1043, N1023);
or OR3 (N1044, N1034, N194, N521);
and AND2 (N1045, N1044, N838);
or OR3 (N1046, N1041, N1042, N871);
and AND3 (N1047, N352, N34, N179);
nand NAND2 (N1048, N1032, N77);
and AND2 (N1049, N1035, N360);
and AND4 (N1050, N1028, N19, N52, N246);
and AND3 (N1051, N1027, N862, N718);
nor NOR2 (N1052, N1046, N84);
buf BUF1 (N1053, N1043);
nand NAND4 (N1054, N1052, N676, N1018, N68);
nand NAND4 (N1055, N1048, N823, N38, N44);
xor XOR2 (N1056, N1045, N644);
and AND3 (N1057, N1037, N614, N790);
xor XOR2 (N1058, N1056, N620);
not NOT1 (N1059, N1050);
not NOT1 (N1060, N1055);
xor XOR2 (N1061, N1047, N539);
buf BUF1 (N1062, N1053);
not NOT1 (N1063, N1049);
and AND3 (N1064, N1059, N655, N668);
nand NAND3 (N1065, N1060, N1030, N227);
nand NAND3 (N1066, N1058, N666, N541);
xor XOR2 (N1067, N1040, N792);
or OR2 (N1068, N1054, N638);
nor NOR2 (N1069, N1057, N615);
nand NAND3 (N1070, N1069, N131, N371);
nand NAND2 (N1071, N1070, N1040);
not NOT1 (N1072, N1071);
buf BUF1 (N1073, N1068);
and AND4 (N1074, N1065, N493, N398, N759);
nor NOR2 (N1075, N1064, N686);
nor NOR2 (N1076, N1067, N471);
and AND4 (N1077, N1076, N240, N864, N208);
nand NAND3 (N1078, N1072, N149, N289);
not NOT1 (N1079, N1077);
not NOT1 (N1080, N1079);
not NOT1 (N1081, N1080);
or OR3 (N1082, N1063, N50, N837);
not NOT1 (N1083, N1082);
and AND3 (N1084, N1075, N330, N212);
nor NOR4 (N1085, N1078, N903, N490, N807);
or OR4 (N1086, N1083, N136, N860, N148);
not NOT1 (N1087, N1051);
not NOT1 (N1088, N1085);
not NOT1 (N1089, N1074);
nor NOR3 (N1090, N1073, N249, N1016);
not NOT1 (N1091, N1089);
nand NAND2 (N1092, N1084, N96);
not NOT1 (N1093, N1086);
xor XOR2 (N1094, N1061, N502);
xor XOR2 (N1095, N1087, N291);
not NOT1 (N1096, N1062);
buf BUF1 (N1097, N1091);
nand NAND2 (N1098, N1092, N290);
buf BUF1 (N1099, N1081);
nand NAND2 (N1100, N1099, N849);
nor NOR2 (N1101, N1066, N850);
nand NAND3 (N1102, N1094, N1076, N368);
xor XOR2 (N1103, N1097, N759);
nand NAND4 (N1104, N1103, N812, N459, N150);
buf BUF1 (N1105, N1102);
nand NAND3 (N1106, N1104, N383, N327);
not NOT1 (N1107, N1106);
buf BUF1 (N1108, N1093);
not NOT1 (N1109, N1088);
buf BUF1 (N1110, N1098);
and AND3 (N1111, N1105, N446, N347);
buf BUF1 (N1112, N1090);
and AND2 (N1113, N1112, N429);
or OR3 (N1114, N1096, N717, N568);
or OR2 (N1115, N1095, N837);
nand NAND4 (N1116, N1108, N1110, N150, N385);
buf BUF1 (N1117, N894);
or OR4 (N1118, N1101, N740, N1105, N556);
buf BUF1 (N1119, N1107);
not NOT1 (N1120, N1117);
nor NOR2 (N1121, N1118, N213);
and AND4 (N1122, N1119, N154, N756, N688);
or OR3 (N1123, N1120, N598, N426);
or OR2 (N1124, N1114, N531);
not NOT1 (N1125, N1109);
buf BUF1 (N1126, N1121);
nand NAND2 (N1127, N1115, N352);
nand NAND3 (N1128, N1126, N181, N107);
buf BUF1 (N1129, N1100);
not NOT1 (N1130, N1113);
nand NAND2 (N1131, N1129, N620);
and AND4 (N1132, N1122, N893, N888, N1075);
nand NAND4 (N1133, N1127, N142, N373, N775);
nand NAND4 (N1134, N1132, N1100, N336, N824);
or OR2 (N1135, N1133, N1097);
nand NAND3 (N1136, N1128, N4, N865);
or OR2 (N1137, N1125, N61);
xor XOR2 (N1138, N1134, N277);
xor XOR2 (N1139, N1111, N629);
nor NOR2 (N1140, N1139, N587);
or OR3 (N1141, N1130, N996, N15);
xor XOR2 (N1142, N1138, N675);
xor XOR2 (N1143, N1140, N144);
and AND4 (N1144, N1124, N457, N499, N199);
nand NAND3 (N1145, N1135, N438, N911);
or OR4 (N1146, N1131, N655, N83, N469);
or OR4 (N1147, N1137, N472, N951, N816);
nor NOR2 (N1148, N1142, N429);
buf BUF1 (N1149, N1136);
nor NOR3 (N1150, N1123, N253, N777);
nand NAND4 (N1151, N1145, N967, N217, N879);
nor NOR4 (N1152, N1141, N257, N837, N1094);
nand NAND4 (N1153, N1151, N1100, N724, N893);
xor XOR2 (N1154, N1150, N1021);
or OR3 (N1155, N1152, N426, N288);
xor XOR2 (N1156, N1149, N949);
not NOT1 (N1157, N1148);
not NOT1 (N1158, N1116);
or OR2 (N1159, N1153, N452);
or OR2 (N1160, N1146, N808);
xor XOR2 (N1161, N1147, N768);
buf BUF1 (N1162, N1144);
buf BUF1 (N1163, N1156);
nor NOR2 (N1164, N1160, N819);
nor NOR2 (N1165, N1161, N940);
buf BUF1 (N1166, N1155);
or OR4 (N1167, N1157, N1160, N1021, N324);
buf BUF1 (N1168, N1162);
or OR3 (N1169, N1167, N551, N428);
xor XOR2 (N1170, N1165, N814);
not NOT1 (N1171, N1164);
nor NOR4 (N1172, N1158, N719, N1136, N1025);
nand NAND3 (N1173, N1169, N219, N1084);
buf BUF1 (N1174, N1171);
not NOT1 (N1175, N1174);
nor NOR2 (N1176, N1166, N878);
buf BUF1 (N1177, N1170);
nand NAND3 (N1178, N1168, N224, N1115);
nor NOR3 (N1179, N1177, N1153, N678);
nor NOR3 (N1180, N1159, N64, N935);
not NOT1 (N1181, N1176);
nand NAND3 (N1182, N1163, N441, N963);
buf BUF1 (N1183, N1173);
or OR2 (N1184, N1179, N373);
nand NAND4 (N1185, N1175, N256, N551, N1141);
not NOT1 (N1186, N1143);
nand NAND2 (N1187, N1178, N131);
or OR2 (N1188, N1187, N724);
nor NOR4 (N1189, N1188, N839, N767, N344);
xor XOR2 (N1190, N1181, N541);
not NOT1 (N1191, N1182);
not NOT1 (N1192, N1184);
or OR4 (N1193, N1154, N215, N554, N344);
nand NAND2 (N1194, N1186, N759);
or OR2 (N1195, N1192, N982);
not NOT1 (N1196, N1194);
not NOT1 (N1197, N1172);
nor NOR2 (N1198, N1180, N924);
or OR3 (N1199, N1195, N400, N450);
nor NOR3 (N1200, N1198, N1139, N986);
and AND3 (N1201, N1193, N1194, N866);
and AND3 (N1202, N1201, N212, N393);
not NOT1 (N1203, N1189);
xor XOR2 (N1204, N1199, N555);
nand NAND3 (N1205, N1190, N197, N831);
nand NAND2 (N1206, N1196, N173);
nand NAND3 (N1207, N1191, N1205, N944);
nand NAND3 (N1208, N519, N684, N159);
or OR2 (N1209, N1200, N938);
or OR2 (N1210, N1207, N152);
and AND2 (N1211, N1204, N185);
buf BUF1 (N1212, N1211);
xor XOR2 (N1213, N1197, N841);
or OR4 (N1214, N1210, N59, N839, N439);
nand NAND3 (N1215, N1206, N1021, N401);
and AND4 (N1216, N1213, N168, N498, N682);
and AND2 (N1217, N1208, N783);
buf BUF1 (N1218, N1214);
not NOT1 (N1219, N1183);
and AND2 (N1220, N1202, N777);
buf BUF1 (N1221, N1220);
nor NOR3 (N1222, N1209, N632, N362);
and AND4 (N1223, N1221, N632, N835, N1153);
nor NOR2 (N1224, N1218, N547);
nor NOR2 (N1225, N1215, N449);
not NOT1 (N1226, N1224);
buf BUF1 (N1227, N1226);
or OR4 (N1228, N1227, N1089, N1015, N1118);
or OR3 (N1229, N1185, N13, N596);
buf BUF1 (N1230, N1217);
and AND2 (N1231, N1228, N982);
or OR3 (N1232, N1212, N628, N91);
nand NAND3 (N1233, N1230, N186, N367);
xor XOR2 (N1234, N1231, N175);
buf BUF1 (N1235, N1232);
nor NOR2 (N1236, N1229, N159);
or OR3 (N1237, N1225, N656, N140);
nor NOR4 (N1238, N1233, N697, N826, N946);
nor NOR4 (N1239, N1219, N232, N139, N1063);
nand NAND2 (N1240, N1216, N754);
xor XOR2 (N1241, N1203, N68);
xor XOR2 (N1242, N1236, N515);
nor NOR4 (N1243, N1234, N38, N985, N632);
or OR2 (N1244, N1235, N731);
buf BUF1 (N1245, N1241);
nand NAND3 (N1246, N1239, N1219, N991);
and AND2 (N1247, N1244, N415);
nor NOR2 (N1248, N1247, N300);
and AND4 (N1249, N1238, N127, N643, N735);
or OR3 (N1250, N1246, N152, N624);
buf BUF1 (N1251, N1222);
nand NAND2 (N1252, N1242, N1088);
or OR4 (N1253, N1250, N1085, N186, N1103);
or OR4 (N1254, N1253, N339, N501, N247);
buf BUF1 (N1255, N1243);
buf BUF1 (N1256, N1254);
not NOT1 (N1257, N1255);
buf BUF1 (N1258, N1240);
not NOT1 (N1259, N1245);
nor NOR4 (N1260, N1251, N566, N605, N1090);
buf BUF1 (N1261, N1259);
xor XOR2 (N1262, N1258, N503);
and AND4 (N1263, N1252, N1182, N221, N452);
buf BUF1 (N1264, N1248);
buf BUF1 (N1265, N1256);
xor XOR2 (N1266, N1260, N917);
nand NAND3 (N1267, N1263, N1073, N703);
buf BUF1 (N1268, N1249);
nand NAND2 (N1269, N1267, N286);
buf BUF1 (N1270, N1266);
or OR4 (N1271, N1264, N745, N555, N253);
nor NOR4 (N1272, N1262, N982, N753, N133);
and AND4 (N1273, N1271, N1087, N1228, N1194);
or OR3 (N1274, N1272, N395, N1051);
not NOT1 (N1275, N1237);
buf BUF1 (N1276, N1268);
or OR3 (N1277, N1223, N309, N1239);
and AND4 (N1278, N1276, N93, N716, N1007);
xor XOR2 (N1279, N1274, N912);
nand NAND2 (N1280, N1278, N390);
not NOT1 (N1281, N1275);
nand NAND3 (N1282, N1269, N847, N588);
and AND2 (N1283, N1281, N716);
not NOT1 (N1284, N1257);
and AND3 (N1285, N1265, N606, N1172);
xor XOR2 (N1286, N1284, N73);
xor XOR2 (N1287, N1270, N505);
nand NAND2 (N1288, N1261, N14);
buf BUF1 (N1289, N1283);
xor XOR2 (N1290, N1288, N837);
and AND3 (N1291, N1287, N581, N35);
nand NAND4 (N1292, N1285, N316, N909, N630);
nor NOR3 (N1293, N1273, N281, N1239);
nor NOR3 (N1294, N1289, N137, N190);
and AND3 (N1295, N1292, N529, N79);
xor XOR2 (N1296, N1290, N438);
and AND2 (N1297, N1279, N11);
xor XOR2 (N1298, N1293, N337);
or OR3 (N1299, N1294, N846, N703);
not NOT1 (N1300, N1297);
xor XOR2 (N1301, N1296, N1089);
nand NAND4 (N1302, N1301, N142, N782, N678);
buf BUF1 (N1303, N1298);
or OR2 (N1304, N1300, N807);
xor XOR2 (N1305, N1277, N96);
xor XOR2 (N1306, N1291, N1098);
buf BUF1 (N1307, N1286);
buf BUF1 (N1308, N1305);
and AND2 (N1309, N1304, N1105);
not NOT1 (N1310, N1308);
buf BUF1 (N1311, N1303);
nand NAND3 (N1312, N1309, N512, N426);
buf BUF1 (N1313, N1307);
nor NOR4 (N1314, N1306, N845, N482, N503);
or OR2 (N1315, N1310, N215);
and AND3 (N1316, N1282, N971, N1267);
xor XOR2 (N1317, N1312, N1088);
not NOT1 (N1318, N1313);
nand NAND2 (N1319, N1317, N1167);
buf BUF1 (N1320, N1315);
or OR2 (N1321, N1318, N1175);
buf BUF1 (N1322, N1314);
nand NAND2 (N1323, N1316, N159);
or OR4 (N1324, N1323, N499, N444, N748);
nor NOR4 (N1325, N1324, N858, N35, N366);
buf BUF1 (N1326, N1311);
nor NOR3 (N1327, N1280, N28, N381);
nand NAND2 (N1328, N1299, N1068);
nand NAND3 (N1329, N1328, N391, N446);
or OR3 (N1330, N1322, N769, N1068);
or OR2 (N1331, N1295, N918);
or OR3 (N1332, N1325, N493, N551);
xor XOR2 (N1333, N1302, N317);
or OR4 (N1334, N1326, N674, N334, N19);
buf BUF1 (N1335, N1334);
or OR3 (N1336, N1329, N211, N499);
nand NAND2 (N1337, N1333, N749);
nor NOR2 (N1338, N1335, N529);
buf BUF1 (N1339, N1330);
buf BUF1 (N1340, N1319);
not NOT1 (N1341, N1336);
not NOT1 (N1342, N1337);
buf BUF1 (N1343, N1341);
not NOT1 (N1344, N1327);
xor XOR2 (N1345, N1344, N1135);
and AND3 (N1346, N1342, N1231, N1133);
xor XOR2 (N1347, N1345, N83);
xor XOR2 (N1348, N1339, N205);
or OR3 (N1349, N1338, N844, N562);
not NOT1 (N1350, N1343);
buf BUF1 (N1351, N1332);
or OR2 (N1352, N1349, N168);
and AND3 (N1353, N1346, N249, N1290);
and AND4 (N1354, N1321, N579, N155, N685);
nor NOR3 (N1355, N1354, N437, N244);
and AND4 (N1356, N1350, N184, N737, N184);
xor XOR2 (N1357, N1352, N106);
nor NOR2 (N1358, N1356, N214);
xor XOR2 (N1359, N1331, N1225);
and AND3 (N1360, N1357, N483, N1075);
nor NOR2 (N1361, N1340, N88);
and AND2 (N1362, N1355, N778);
nand NAND3 (N1363, N1351, N560, N1182);
not NOT1 (N1364, N1358);
xor XOR2 (N1365, N1347, N537);
and AND2 (N1366, N1320, N879);
nor NOR2 (N1367, N1363, N1076);
nor NOR2 (N1368, N1365, N636);
not NOT1 (N1369, N1360);
xor XOR2 (N1370, N1367, N181);
nor NOR4 (N1371, N1370, N117, N222, N279);
nand NAND2 (N1372, N1359, N924);
buf BUF1 (N1373, N1362);
nand NAND4 (N1374, N1353, N451, N626, N445);
xor XOR2 (N1375, N1374, N987);
or OR2 (N1376, N1372, N30);
xor XOR2 (N1377, N1348, N721);
buf BUF1 (N1378, N1376);
nand NAND3 (N1379, N1369, N1224, N1325);
not NOT1 (N1380, N1371);
buf BUF1 (N1381, N1378);
buf BUF1 (N1382, N1364);
buf BUF1 (N1383, N1379);
not NOT1 (N1384, N1383);
not NOT1 (N1385, N1380);
and AND3 (N1386, N1373, N867, N931);
or OR2 (N1387, N1384, N625);
nand NAND3 (N1388, N1382, N211, N158);
not NOT1 (N1389, N1385);
nor NOR2 (N1390, N1388, N321);
not NOT1 (N1391, N1390);
and AND2 (N1392, N1361, N310);
xor XOR2 (N1393, N1387, N397);
xor XOR2 (N1394, N1391, N1085);
not NOT1 (N1395, N1389);
not NOT1 (N1396, N1377);
or OR4 (N1397, N1366, N1279, N493, N1006);
or OR4 (N1398, N1397, N895, N455, N444);
nand NAND4 (N1399, N1375, N571, N599, N1354);
xor XOR2 (N1400, N1399, N989);
nor NOR4 (N1401, N1396, N518, N1010, N350);
xor XOR2 (N1402, N1368, N300);
not NOT1 (N1403, N1398);
buf BUF1 (N1404, N1381);
not NOT1 (N1405, N1403);
nand NAND4 (N1406, N1392, N15, N380, N821);
and AND3 (N1407, N1400, N196, N107);
and AND3 (N1408, N1402, N576, N1039);
xor XOR2 (N1409, N1395, N308);
not NOT1 (N1410, N1407);
nand NAND4 (N1411, N1386, N21, N55, N342);
nor NOR2 (N1412, N1406, N177);
and AND3 (N1413, N1410, N616, N1377);
nand NAND4 (N1414, N1405, N104, N279, N701);
and AND3 (N1415, N1394, N229, N83);
not NOT1 (N1416, N1415);
or OR2 (N1417, N1401, N1106);
nor NOR2 (N1418, N1393, N259);
buf BUF1 (N1419, N1414);
and AND3 (N1420, N1412, N1218, N1015);
and AND2 (N1421, N1419, N1064);
or OR3 (N1422, N1409, N1230, N1334);
xor XOR2 (N1423, N1418, N184);
buf BUF1 (N1424, N1417);
nand NAND3 (N1425, N1416, N756, N138);
nor NOR3 (N1426, N1422, N879, N1357);
nor NOR4 (N1427, N1420, N1260, N436, N1410);
not NOT1 (N1428, N1426);
xor XOR2 (N1429, N1408, N350);
nor NOR4 (N1430, N1428, N406, N121, N1088);
nand NAND2 (N1431, N1421, N313);
nand NAND4 (N1432, N1427, N878, N1307, N705);
and AND2 (N1433, N1431, N736);
nand NAND4 (N1434, N1404, N1009, N1327, N1239);
and AND3 (N1435, N1429, N127, N913);
or OR4 (N1436, N1435, N153, N649, N882);
xor XOR2 (N1437, N1423, N544);
and AND4 (N1438, N1432, N818, N742, N729);
not NOT1 (N1439, N1411);
buf BUF1 (N1440, N1430);
xor XOR2 (N1441, N1413, N143);
and AND4 (N1442, N1425, N557, N1135, N569);
and AND4 (N1443, N1439, N1322, N1087, N374);
and AND3 (N1444, N1437, N194, N1138);
and AND2 (N1445, N1440, N1313);
nand NAND3 (N1446, N1438, N973, N906);
and AND2 (N1447, N1424, N703);
nand NAND4 (N1448, N1436, N243, N1127, N2);
not NOT1 (N1449, N1443);
or OR4 (N1450, N1445, N28, N1177, N1197);
and AND2 (N1451, N1441, N668);
and AND3 (N1452, N1447, N1050, N1207);
nor NOR2 (N1453, N1442, N719);
buf BUF1 (N1454, N1452);
and AND3 (N1455, N1433, N762, N1020);
xor XOR2 (N1456, N1450, N125);
xor XOR2 (N1457, N1453, N499);
buf BUF1 (N1458, N1455);
nor NOR3 (N1459, N1444, N203, N1272);
nand NAND2 (N1460, N1458, N343);
not NOT1 (N1461, N1446);
nand NAND4 (N1462, N1451, N1192, N1384, N822);
nor NOR3 (N1463, N1462, N557, N867);
and AND4 (N1464, N1456, N231, N129, N818);
xor XOR2 (N1465, N1464, N49);
xor XOR2 (N1466, N1457, N487);
and AND2 (N1467, N1434, N1034);
nand NAND3 (N1468, N1449, N1422, N1244);
or OR3 (N1469, N1463, N822, N670);
or OR3 (N1470, N1467, N839, N1340);
or OR4 (N1471, N1448, N1102, N124, N718);
and AND4 (N1472, N1454, N511, N1470, N439);
or OR2 (N1473, N1394, N1457);
buf BUF1 (N1474, N1472);
nand NAND3 (N1475, N1461, N1344, N317);
nor NOR4 (N1476, N1469, N1023, N1262, N36);
nor NOR2 (N1477, N1466, N111);
xor XOR2 (N1478, N1477, N237);
buf BUF1 (N1479, N1460);
buf BUF1 (N1480, N1479);
xor XOR2 (N1481, N1476, N633);
nor NOR4 (N1482, N1473, N63, N323, N730);
not NOT1 (N1483, N1482);
not NOT1 (N1484, N1480);
xor XOR2 (N1485, N1475, N536);
xor XOR2 (N1486, N1468, N969);
xor XOR2 (N1487, N1481, N454);
nor NOR4 (N1488, N1485, N182, N1348, N297);
xor XOR2 (N1489, N1487, N1329);
not NOT1 (N1490, N1483);
xor XOR2 (N1491, N1484, N1313);
and AND3 (N1492, N1474, N1399, N55);
buf BUF1 (N1493, N1471);
not NOT1 (N1494, N1459);
buf BUF1 (N1495, N1478);
nor NOR4 (N1496, N1489, N1238, N36, N301);
or OR4 (N1497, N1493, N650, N721, N1081);
nand NAND2 (N1498, N1494, N1443);
nor NOR3 (N1499, N1496, N1038, N688);
buf BUF1 (N1500, N1497);
xor XOR2 (N1501, N1492, N926);
xor XOR2 (N1502, N1498, N614);
nand NAND3 (N1503, N1465, N1198, N596);
nand NAND4 (N1504, N1502, N993, N690, N243);
nand NAND2 (N1505, N1503, N201);
or OR3 (N1506, N1500, N902, N365);
not NOT1 (N1507, N1490);
nor NOR2 (N1508, N1499, N1307);
or OR3 (N1509, N1505, N1188, N971);
or OR2 (N1510, N1504, N1253);
or OR4 (N1511, N1495, N287, N818, N279);
nor NOR3 (N1512, N1510, N965, N879);
not NOT1 (N1513, N1512);
nand NAND3 (N1514, N1488, N1501, N47);
not NOT1 (N1515, N409);
and AND2 (N1516, N1514, N1332);
nand NAND4 (N1517, N1513, N595, N100, N1059);
not NOT1 (N1518, N1507);
buf BUF1 (N1519, N1508);
or OR4 (N1520, N1515, N209, N712, N840);
nand NAND3 (N1521, N1486, N1444, N1354);
or OR4 (N1522, N1520, N697, N1084, N517);
and AND4 (N1523, N1518, N1262, N1160, N293);
not NOT1 (N1524, N1516);
and AND4 (N1525, N1522, N1395, N187, N1275);
xor XOR2 (N1526, N1525, N1143);
or OR4 (N1527, N1524, N982, N791, N292);
not NOT1 (N1528, N1526);
buf BUF1 (N1529, N1506);
buf BUF1 (N1530, N1521);
xor XOR2 (N1531, N1509, N1255);
xor XOR2 (N1532, N1529, N745);
nor NOR3 (N1533, N1511, N672, N993);
buf BUF1 (N1534, N1531);
or OR4 (N1535, N1528, N1261, N950, N366);
not NOT1 (N1536, N1534);
or OR3 (N1537, N1533, N1429, N1178);
xor XOR2 (N1538, N1536, N270);
and AND2 (N1539, N1517, N88);
xor XOR2 (N1540, N1527, N1182);
or OR3 (N1541, N1519, N76, N1189);
xor XOR2 (N1542, N1541, N220);
nand NAND2 (N1543, N1532, N626);
and AND4 (N1544, N1538, N764, N831, N594);
nand NAND2 (N1545, N1539, N461);
or OR3 (N1546, N1537, N549, N320);
nor NOR4 (N1547, N1523, N713, N802, N1267);
buf BUF1 (N1548, N1547);
xor XOR2 (N1549, N1545, N360);
or OR2 (N1550, N1530, N579);
buf BUF1 (N1551, N1549);
xor XOR2 (N1552, N1535, N1392);
or OR2 (N1553, N1543, N251);
and AND4 (N1554, N1546, N530, N740, N1329);
not NOT1 (N1555, N1553);
not NOT1 (N1556, N1552);
nor NOR3 (N1557, N1548, N1268, N1343);
not NOT1 (N1558, N1556);
nor NOR2 (N1559, N1550, N322);
not NOT1 (N1560, N1540);
xor XOR2 (N1561, N1559, N937);
buf BUF1 (N1562, N1544);
xor XOR2 (N1563, N1562, N1471);
xor XOR2 (N1564, N1551, N1476);
buf BUF1 (N1565, N1564);
buf BUF1 (N1566, N1554);
xor XOR2 (N1567, N1563, N107);
not NOT1 (N1568, N1565);
or OR3 (N1569, N1491, N1289, N418);
buf BUF1 (N1570, N1569);
xor XOR2 (N1571, N1555, N1432);
and AND4 (N1572, N1560, N523, N1536, N1014);
nor NOR3 (N1573, N1570, N715, N326);
buf BUF1 (N1574, N1572);
not NOT1 (N1575, N1558);
and AND2 (N1576, N1571, N1523);
not NOT1 (N1577, N1574);
nand NAND2 (N1578, N1557, N1028);
nor NOR3 (N1579, N1578, N451, N1516);
nand NAND3 (N1580, N1561, N871, N614);
nor NOR3 (N1581, N1568, N1354, N291);
buf BUF1 (N1582, N1580);
not NOT1 (N1583, N1582);
xor XOR2 (N1584, N1579, N351);
or OR2 (N1585, N1577, N1447);
xor XOR2 (N1586, N1573, N507);
and AND2 (N1587, N1576, N1197);
not NOT1 (N1588, N1587);
and AND3 (N1589, N1566, N57, N737);
or OR3 (N1590, N1575, N882, N570);
nand NAND3 (N1591, N1584, N1176, N232);
not NOT1 (N1592, N1586);
or OR2 (N1593, N1590, N1507);
nor NOR3 (N1594, N1589, N1125, N1407);
nor NOR4 (N1595, N1581, N1470, N98, N1498);
nand NAND4 (N1596, N1593, N1176, N159, N895);
xor XOR2 (N1597, N1567, N1291);
not NOT1 (N1598, N1591);
or OR2 (N1599, N1542, N1555);
nor NOR4 (N1600, N1594, N1256, N1117, N1349);
nand NAND3 (N1601, N1597, N1381, N1451);
xor XOR2 (N1602, N1598, N134);
xor XOR2 (N1603, N1583, N826);
buf BUF1 (N1604, N1585);
xor XOR2 (N1605, N1603, N1309);
buf BUF1 (N1606, N1599);
nand NAND2 (N1607, N1602, N1572);
buf BUF1 (N1608, N1601);
not NOT1 (N1609, N1605);
or OR3 (N1610, N1604, N69, N1180);
nor NOR4 (N1611, N1607, N408, N750, N44);
buf BUF1 (N1612, N1592);
xor XOR2 (N1613, N1606, N896);
nor NOR2 (N1614, N1608, N255);
xor XOR2 (N1615, N1600, N779);
and AND3 (N1616, N1609, N509, N779);
or OR4 (N1617, N1613, N1236, N440, N1612);
nor NOR2 (N1618, N867, N1238);
or OR3 (N1619, N1596, N1331, N1375);
nand NAND3 (N1620, N1615, N287, N625);
xor XOR2 (N1621, N1614, N523);
or OR3 (N1622, N1620, N712, N201);
and AND3 (N1623, N1621, N1009, N1103);
xor XOR2 (N1624, N1623, N963);
nor NOR2 (N1625, N1618, N1265);
xor XOR2 (N1626, N1617, N1191);
xor XOR2 (N1627, N1595, N1165);
nand NAND2 (N1628, N1619, N1103);
not NOT1 (N1629, N1627);
xor XOR2 (N1630, N1625, N1180);
buf BUF1 (N1631, N1610);
nand NAND4 (N1632, N1588, N873, N60, N1536);
or OR3 (N1633, N1626, N288, N622);
xor XOR2 (N1634, N1630, N797);
not NOT1 (N1635, N1632);
nor NOR4 (N1636, N1634, N1044, N1432, N1491);
xor XOR2 (N1637, N1636, N1195);
and AND3 (N1638, N1624, N1139, N1534);
xor XOR2 (N1639, N1633, N946);
xor XOR2 (N1640, N1629, N972);
nor NOR3 (N1641, N1639, N183, N594);
or OR2 (N1642, N1638, N510);
or OR2 (N1643, N1622, N91);
xor XOR2 (N1644, N1643, N1042);
nor NOR3 (N1645, N1628, N385, N1617);
xor XOR2 (N1646, N1631, N838);
nand NAND2 (N1647, N1640, N135);
not NOT1 (N1648, N1646);
xor XOR2 (N1649, N1641, N240);
nor NOR4 (N1650, N1635, N311, N1334, N375);
not NOT1 (N1651, N1649);
or OR2 (N1652, N1611, N1558);
nor NOR4 (N1653, N1651, N1497, N476, N1287);
xor XOR2 (N1654, N1642, N1165);
not NOT1 (N1655, N1654);
and AND4 (N1656, N1655, N862, N784, N188);
nand NAND2 (N1657, N1652, N1492);
nor NOR2 (N1658, N1650, N1613);
xor XOR2 (N1659, N1648, N241);
buf BUF1 (N1660, N1645);
and AND4 (N1661, N1657, N1551, N1041, N1159);
not NOT1 (N1662, N1653);
buf BUF1 (N1663, N1644);
not NOT1 (N1664, N1660);
nand NAND4 (N1665, N1647, N55, N230, N1252);
nand NAND4 (N1666, N1663, N948, N482, N318);
not NOT1 (N1667, N1665);
xor XOR2 (N1668, N1664, N1073);
and AND2 (N1669, N1658, N733);
nand NAND2 (N1670, N1662, N292);
nand NAND3 (N1671, N1637, N857, N912);
not NOT1 (N1672, N1669);
buf BUF1 (N1673, N1671);
nor NOR2 (N1674, N1666, N370);
buf BUF1 (N1675, N1672);
nand NAND2 (N1676, N1667, N1054);
nand NAND2 (N1677, N1675, N134);
nor NOR3 (N1678, N1659, N118, N1013);
or OR2 (N1679, N1676, N622);
nor NOR2 (N1680, N1673, N1002);
nor NOR3 (N1681, N1656, N831, N1445);
xor XOR2 (N1682, N1678, N1228);
or OR4 (N1683, N1668, N879, N857, N1243);
xor XOR2 (N1684, N1661, N1060);
nor NOR2 (N1685, N1677, N1131);
nor NOR3 (N1686, N1683, N1438, N721);
nor NOR2 (N1687, N1682, N1159);
or OR3 (N1688, N1616, N480, N1409);
xor XOR2 (N1689, N1686, N210);
buf BUF1 (N1690, N1687);
buf BUF1 (N1691, N1670);
and AND2 (N1692, N1690, N1382);
xor XOR2 (N1693, N1688, N210);
or OR3 (N1694, N1691, N1666, N1148);
nor NOR4 (N1695, N1679, N624, N1201, N1503);
not NOT1 (N1696, N1693);
not NOT1 (N1697, N1695);
and AND2 (N1698, N1684, N1053);
nor NOR4 (N1699, N1697, N748, N462, N1199);
buf BUF1 (N1700, N1698);
not NOT1 (N1701, N1674);
not NOT1 (N1702, N1701);
nor NOR4 (N1703, N1689, N461, N840, N1599);
nand NAND3 (N1704, N1702, N1620, N1379);
and AND3 (N1705, N1692, N1519, N208);
buf BUF1 (N1706, N1700);
nor NOR3 (N1707, N1696, N1442, N647);
buf BUF1 (N1708, N1681);
not NOT1 (N1709, N1685);
not NOT1 (N1710, N1705);
xor XOR2 (N1711, N1703, N59);
or OR3 (N1712, N1694, N1159, N1551);
buf BUF1 (N1713, N1711);
and AND4 (N1714, N1704, N767, N478, N300);
nor NOR2 (N1715, N1708, N1085);
or OR3 (N1716, N1715, N703, N50);
not NOT1 (N1717, N1710);
and AND3 (N1718, N1709, N1203, N195);
nand NAND2 (N1719, N1699, N1655);
xor XOR2 (N1720, N1717, N425);
and AND2 (N1721, N1719, N951);
and AND4 (N1722, N1713, N997, N1462, N1122);
xor XOR2 (N1723, N1714, N849);
xor XOR2 (N1724, N1720, N1377);
xor XOR2 (N1725, N1718, N1168);
and AND3 (N1726, N1706, N1336, N930);
nand NAND3 (N1727, N1725, N14, N1607);
not NOT1 (N1728, N1724);
not NOT1 (N1729, N1728);
buf BUF1 (N1730, N1729);
not NOT1 (N1731, N1707);
buf BUF1 (N1732, N1730);
not NOT1 (N1733, N1726);
nand NAND3 (N1734, N1727, N1156, N904);
buf BUF1 (N1735, N1731);
not NOT1 (N1736, N1712);
buf BUF1 (N1737, N1732);
nor NOR4 (N1738, N1736, N1342, N286, N1428);
nor NOR2 (N1739, N1735, N207);
or OR4 (N1740, N1680, N626, N1644, N313);
not NOT1 (N1741, N1739);
and AND2 (N1742, N1734, N507);
nor NOR4 (N1743, N1738, N1369, N901, N1437);
and AND3 (N1744, N1741, N1609, N396);
nand NAND4 (N1745, N1722, N582, N1117, N688);
xor XOR2 (N1746, N1737, N1569);
or OR4 (N1747, N1723, N502, N27, N1595);
not NOT1 (N1748, N1740);
not NOT1 (N1749, N1745);
or OR2 (N1750, N1747, N582);
nand NAND4 (N1751, N1744, N1677, N1254, N1391);
nor NOR4 (N1752, N1716, N1411, N1611, N1031);
nand NAND3 (N1753, N1743, N93, N879);
xor XOR2 (N1754, N1752, N1668);
nand NAND3 (N1755, N1748, N540, N1732);
not NOT1 (N1756, N1755);
or OR2 (N1757, N1750, N588);
or OR4 (N1758, N1757, N710, N280, N865);
or OR3 (N1759, N1756, N440, N71);
and AND4 (N1760, N1742, N564, N307, N1028);
and AND3 (N1761, N1758, N251, N596);
and AND3 (N1762, N1761, N1468, N962);
nand NAND4 (N1763, N1760, N912, N1191, N1161);
not NOT1 (N1764, N1749);
nand NAND4 (N1765, N1733, N376, N824, N275);
not NOT1 (N1766, N1721);
and AND2 (N1767, N1759, N1675);
and AND4 (N1768, N1764, N368, N1531, N864);
not NOT1 (N1769, N1754);
buf BUF1 (N1770, N1746);
nor NOR2 (N1771, N1768, N1388);
not NOT1 (N1772, N1767);
nor NOR2 (N1773, N1769, N889);
xor XOR2 (N1774, N1773, N1295);
xor XOR2 (N1775, N1751, N1657);
nor NOR3 (N1776, N1774, N1524, N1452);
and AND3 (N1777, N1762, N848, N707);
nand NAND2 (N1778, N1766, N1034);
nor NOR3 (N1779, N1771, N913, N1758);
nand NAND2 (N1780, N1779, N174);
nor NOR2 (N1781, N1778, N180);
nor NOR2 (N1782, N1781, N579);
buf BUF1 (N1783, N1775);
or OR2 (N1784, N1753, N15);
nand NAND2 (N1785, N1783, N275);
not NOT1 (N1786, N1765);
nor NOR4 (N1787, N1786, N1033, N373, N1163);
buf BUF1 (N1788, N1787);
or OR2 (N1789, N1788, N195);
xor XOR2 (N1790, N1763, N552);
nor NOR2 (N1791, N1777, N1572);
or OR4 (N1792, N1791, N951, N1210, N1032);
and AND4 (N1793, N1784, N235, N1090, N354);
nand NAND4 (N1794, N1772, N426, N465, N1574);
or OR2 (N1795, N1793, N1279);
or OR2 (N1796, N1785, N1114);
nor NOR3 (N1797, N1794, N1078, N5);
not NOT1 (N1798, N1796);
buf BUF1 (N1799, N1798);
nor NOR2 (N1800, N1770, N262);
buf BUF1 (N1801, N1789);
buf BUF1 (N1802, N1790);
not NOT1 (N1803, N1780);
nor NOR4 (N1804, N1800, N1439, N1098, N882);
and AND3 (N1805, N1804, N1301, N585);
buf BUF1 (N1806, N1782);
or OR2 (N1807, N1806, N1736);
or OR4 (N1808, N1795, N1151, N517, N502);
or OR4 (N1809, N1792, N262, N765, N1016);
nand NAND4 (N1810, N1803, N1163, N858, N814);
nand NAND4 (N1811, N1807, N1188, N397, N920);
buf BUF1 (N1812, N1811);
and AND3 (N1813, N1808, N1210, N739);
nand NAND4 (N1814, N1812, N262, N1031, N75);
nor NOR4 (N1815, N1801, N1732, N610, N1537);
xor XOR2 (N1816, N1797, N241);
xor XOR2 (N1817, N1815, N821);
not NOT1 (N1818, N1799);
nand NAND3 (N1819, N1814, N281, N173);
not NOT1 (N1820, N1813);
buf BUF1 (N1821, N1805);
xor XOR2 (N1822, N1820, N1698);
nand NAND4 (N1823, N1821, N1190, N1710, N76);
nand NAND4 (N1824, N1776, N1543, N1039, N1581);
nand NAND3 (N1825, N1817, N1084, N634);
nor NOR2 (N1826, N1819, N623);
not NOT1 (N1827, N1810);
nand NAND3 (N1828, N1825, N332, N64);
buf BUF1 (N1829, N1826);
xor XOR2 (N1830, N1823, N829);
and AND3 (N1831, N1802, N531, N1205);
and AND4 (N1832, N1830, N1504, N1532, N96);
or OR3 (N1833, N1816, N1619, N221);
nand NAND4 (N1834, N1818, N678, N1373, N240);
nor NOR2 (N1835, N1832, N1065);
not NOT1 (N1836, N1828);
not NOT1 (N1837, N1835);
nor NOR3 (N1838, N1809, N1315, N825);
not NOT1 (N1839, N1837);
or OR3 (N1840, N1833, N1647, N1661);
buf BUF1 (N1841, N1834);
nor NOR2 (N1842, N1836, N308);
nand NAND3 (N1843, N1827, N399, N238);
nor NOR3 (N1844, N1843, N1418, N1336);
xor XOR2 (N1845, N1840, N550);
and AND3 (N1846, N1842, N442, N1238);
buf BUF1 (N1847, N1846);
not NOT1 (N1848, N1831);
buf BUF1 (N1849, N1824);
nand NAND3 (N1850, N1849, N1293, N36);
buf BUF1 (N1851, N1845);
nand NAND3 (N1852, N1841, N785, N1030);
buf BUF1 (N1853, N1848);
xor XOR2 (N1854, N1838, N31);
or OR3 (N1855, N1852, N1235, N1170);
or OR2 (N1856, N1850, N931);
xor XOR2 (N1857, N1839, N1032);
xor XOR2 (N1858, N1847, N1624);
and AND4 (N1859, N1844, N423, N768, N620);
or OR4 (N1860, N1856, N358, N518, N462);
and AND3 (N1861, N1857, N1403, N335);
buf BUF1 (N1862, N1861);
nand NAND2 (N1863, N1854, N1105);
or OR4 (N1864, N1855, N1181, N670, N948);
nand NAND2 (N1865, N1853, N10);
not NOT1 (N1866, N1864);
buf BUF1 (N1867, N1863);
not NOT1 (N1868, N1822);
and AND4 (N1869, N1865, N805, N12, N489);
buf BUF1 (N1870, N1866);
or OR2 (N1871, N1868, N1139);
nand NAND2 (N1872, N1870, N661);
or OR3 (N1873, N1869, N252, N489);
nand NAND3 (N1874, N1851, N1421, N1693);
or OR2 (N1875, N1860, N816);
nand NAND2 (N1876, N1829, N693);
buf BUF1 (N1877, N1858);
nand NAND3 (N1878, N1862, N836, N1233);
xor XOR2 (N1879, N1871, N38);
and AND4 (N1880, N1874, N587, N1396, N1585);
xor XOR2 (N1881, N1875, N1556);
not NOT1 (N1882, N1876);
and AND2 (N1883, N1867, N1463);
and AND2 (N1884, N1882, N505);
or OR3 (N1885, N1859, N1402, N1552);
xor XOR2 (N1886, N1881, N1558);
xor XOR2 (N1887, N1873, N1570);
not NOT1 (N1888, N1878);
buf BUF1 (N1889, N1872);
not NOT1 (N1890, N1888);
not NOT1 (N1891, N1877);
not NOT1 (N1892, N1891);
xor XOR2 (N1893, N1887, N566);
nor NOR4 (N1894, N1880, N778, N433, N1430);
and AND3 (N1895, N1883, N745, N189);
buf BUF1 (N1896, N1893);
xor XOR2 (N1897, N1896, N248);
nand NAND4 (N1898, N1894, N1200, N33, N736);
and AND2 (N1899, N1895, N1353);
buf BUF1 (N1900, N1879);
or OR3 (N1901, N1885, N870, N1177);
nand NAND2 (N1902, N1897, N824);
or OR4 (N1903, N1898, N975, N914, N1353);
buf BUF1 (N1904, N1886);
and AND3 (N1905, N1901, N225, N1884);
xor XOR2 (N1906, N1240, N1391);
and AND2 (N1907, N1889, N477);
nand NAND4 (N1908, N1907, N1052, N1149, N1152);
and AND3 (N1909, N1905, N1245, N1097);
not NOT1 (N1910, N1906);
or OR4 (N1911, N1892, N123, N644, N186);
or OR2 (N1912, N1908, N1512);
buf BUF1 (N1913, N1903);
nand NAND2 (N1914, N1913, N372);
or OR2 (N1915, N1912, N564);
nand NAND4 (N1916, N1899, N1454, N241, N1750);
or OR4 (N1917, N1911, N1622, N55, N202);
and AND3 (N1918, N1916, N695, N1715);
or OR2 (N1919, N1900, N1097);
xor XOR2 (N1920, N1918, N813);
nand NAND3 (N1921, N1904, N471, N584);
xor XOR2 (N1922, N1915, N100);
and AND3 (N1923, N1920, N1140, N331);
not NOT1 (N1924, N1914);
or OR3 (N1925, N1923, N1242, N552);
nand NAND4 (N1926, N1919, N1600, N724, N465);
buf BUF1 (N1927, N1922);
nor NOR4 (N1928, N1910, N575, N11, N574);
or OR4 (N1929, N1926, N1620, N950, N623);
nor NOR3 (N1930, N1927, N1122, N948);
xor XOR2 (N1931, N1925, N1928);
or OR3 (N1932, N1652, N916, N747);
and AND3 (N1933, N1890, N1311, N5);
buf BUF1 (N1934, N1930);
xor XOR2 (N1935, N1917, N1479);
not NOT1 (N1936, N1933);
nor NOR3 (N1937, N1902, N1804, N466);
nand NAND2 (N1938, N1924, N1350);
nor NOR2 (N1939, N1921, N1443);
buf BUF1 (N1940, N1932);
nand NAND2 (N1941, N1931, N968);
buf BUF1 (N1942, N1934);
or OR4 (N1943, N1942, N1720, N1583, N1917);
nand NAND3 (N1944, N1938, N347, N184);
nand NAND3 (N1945, N1909, N1930, N1356);
buf BUF1 (N1946, N1944);
buf BUF1 (N1947, N1945);
xor XOR2 (N1948, N1941, N676);
nor NOR3 (N1949, N1929, N753, N1258);
buf BUF1 (N1950, N1937);
buf BUF1 (N1951, N1939);
not NOT1 (N1952, N1943);
xor XOR2 (N1953, N1950, N1189);
nor NOR4 (N1954, N1949, N1120, N592, N14);
buf BUF1 (N1955, N1947);
buf BUF1 (N1956, N1935);
not NOT1 (N1957, N1956);
buf BUF1 (N1958, N1940);
nand NAND3 (N1959, N1954, N1935, N1313);
nor NOR4 (N1960, N1951, N332, N126, N1597);
xor XOR2 (N1961, N1955, N1015);
and AND3 (N1962, N1958, N409, N944);
or OR4 (N1963, N1960, N187, N1313, N1864);
and AND4 (N1964, N1936, N1568, N369, N1658);
not NOT1 (N1965, N1957);
nand NAND2 (N1966, N1959, N403);
not NOT1 (N1967, N1946);
nor NOR2 (N1968, N1948, N260);
or OR3 (N1969, N1964, N163, N257);
xor XOR2 (N1970, N1966, N126);
nand NAND3 (N1971, N1952, N653, N1711);
buf BUF1 (N1972, N1965);
and AND4 (N1973, N1962, N1828, N180, N1451);
nor NOR4 (N1974, N1968, N1825, N1066, N13);
nand NAND2 (N1975, N1972, N1450);
or OR3 (N1976, N1963, N1465, N1723);
and AND3 (N1977, N1971, N1077, N1486);
and AND2 (N1978, N1975, N1699);
not NOT1 (N1979, N1974);
and AND2 (N1980, N1977, N1712);
not NOT1 (N1981, N1980);
or OR2 (N1982, N1970, N807);
nor NOR3 (N1983, N1979, N96, N708);
nor NOR3 (N1984, N1969, N1519, N602);
and AND2 (N1985, N1976, N430);
buf BUF1 (N1986, N1982);
and AND4 (N1987, N1985, N570, N1656, N1824);
buf BUF1 (N1988, N1978);
or OR4 (N1989, N1988, N1985, N1059, N1123);
nand NAND2 (N1990, N1989, N1314);
and AND4 (N1991, N1981, N623, N1506, N1775);
xor XOR2 (N1992, N1973, N1123);
buf BUF1 (N1993, N1990);
buf BUF1 (N1994, N1967);
nand NAND4 (N1995, N1984, N407, N142, N1515);
buf BUF1 (N1996, N1987);
xor XOR2 (N1997, N1986, N1121);
xor XOR2 (N1998, N1991, N756);
or OR2 (N1999, N1995, N284);
xor XOR2 (N2000, N1994, N488);
or OR3 (N2001, N1997, N1009, N1364);
nand NAND2 (N2002, N2001, N1384);
nand NAND3 (N2003, N1999, N14, N1070);
nor NOR2 (N2004, N1992, N1652);
xor XOR2 (N2005, N1993, N891);
nand NAND3 (N2006, N2000, N1614, N45);
not NOT1 (N2007, N1996);
or OR4 (N2008, N2004, N2004, N74, N1067);
and AND2 (N2009, N2008, N898);
not NOT1 (N2010, N2003);
nor NOR4 (N2011, N2010, N1030, N1674, N1647);
and AND2 (N2012, N1983, N1166);
not NOT1 (N2013, N2002);
not NOT1 (N2014, N1998);
and AND2 (N2015, N2013, N1810);
nand NAND2 (N2016, N2005, N1053);
and AND3 (N2017, N1953, N374, N1642);
or OR4 (N2018, N2016, N1848, N1369, N1916);
nor NOR3 (N2019, N2014, N1118, N441);
buf BUF1 (N2020, N2019);
or OR2 (N2021, N1961, N593);
nand NAND2 (N2022, N2009, N584);
nor NOR3 (N2023, N2011, N1700, N1144);
buf BUF1 (N2024, N2018);
xor XOR2 (N2025, N2024, N218);
and AND2 (N2026, N2017, N1489);
or OR3 (N2027, N2007, N552, N1665);
buf BUF1 (N2028, N2012);
not NOT1 (N2029, N2023);
nand NAND2 (N2030, N2026, N1417);
or OR3 (N2031, N2027, N72, N1285);
nor NOR2 (N2032, N2030, N1338);
xor XOR2 (N2033, N2025, N23);
nand NAND4 (N2034, N2029, N638, N1976, N738);
nand NAND3 (N2035, N2015, N865, N416);
not NOT1 (N2036, N2031);
not NOT1 (N2037, N2028);
nor NOR4 (N2038, N2006, N1879, N1415, N1047);
xor XOR2 (N2039, N2022, N1888);
and AND3 (N2040, N2039, N1362, N2015);
nor NOR2 (N2041, N2035, N396);
buf BUF1 (N2042, N2036);
not NOT1 (N2043, N2038);
xor XOR2 (N2044, N2034, N514);
buf BUF1 (N2045, N2021);
buf BUF1 (N2046, N2037);
nand NAND2 (N2047, N2020, N270);
buf BUF1 (N2048, N2040);
or OR4 (N2049, N2046, N87, N312, N1882);
xor XOR2 (N2050, N2041, N1936);
nor NOR2 (N2051, N2042, N1334);
buf BUF1 (N2052, N2049);
or OR2 (N2053, N2052, N412);
and AND4 (N2054, N2053, N1155, N101, N92);
or OR2 (N2055, N2033, N1196);
buf BUF1 (N2056, N2054);
or OR4 (N2057, N2045, N673, N108, N1073);
nand NAND4 (N2058, N2057, N483, N1955, N1764);
nand NAND4 (N2059, N2050, N769, N907, N409);
buf BUF1 (N2060, N2059);
and AND3 (N2061, N2058, N46, N473);
nand NAND4 (N2062, N2047, N1383, N809, N981);
nand NAND3 (N2063, N2061, N1130, N626);
not NOT1 (N2064, N2062);
and AND4 (N2065, N2044, N426, N1177, N1360);
not NOT1 (N2066, N2055);
or OR3 (N2067, N2060, N1030, N1449);
or OR3 (N2068, N2063, N292, N558);
not NOT1 (N2069, N2048);
buf BUF1 (N2070, N2043);
and AND3 (N2071, N2065, N1279, N1928);
and AND4 (N2072, N2068, N932, N1303, N1735);
buf BUF1 (N2073, N2070);
not NOT1 (N2074, N2056);
and AND4 (N2075, N2069, N597, N1049, N1421);
or OR4 (N2076, N2067, N1430, N1036, N1846);
nand NAND4 (N2077, N2071, N1147, N37, N735);
xor XOR2 (N2078, N2066, N1354);
buf BUF1 (N2079, N2064);
not NOT1 (N2080, N2078);
xor XOR2 (N2081, N2077, N1957);
and AND3 (N2082, N2072, N330, N649);
not NOT1 (N2083, N2051);
xor XOR2 (N2084, N2074, N117);
nand NAND2 (N2085, N2073, N364);
and AND2 (N2086, N2080, N1963);
not NOT1 (N2087, N2079);
nor NOR3 (N2088, N2087, N1465, N1756);
nand NAND3 (N2089, N2088, N1634, N332);
buf BUF1 (N2090, N2086);
nand NAND3 (N2091, N2085, N328, N528);
xor XOR2 (N2092, N2089, N1949);
and AND2 (N2093, N2090, N2068);
buf BUF1 (N2094, N2032);
nor NOR4 (N2095, N2093, N795, N1313, N1319);
nand NAND2 (N2096, N2084, N668);
nand NAND4 (N2097, N2076, N360, N1501, N728);
not NOT1 (N2098, N2095);
buf BUF1 (N2099, N2094);
nand NAND2 (N2100, N2091, N382);
nor NOR2 (N2101, N2075, N638);
or OR3 (N2102, N2099, N1883, N380);
buf BUF1 (N2103, N2101);
buf BUF1 (N2104, N2097);
nand NAND2 (N2105, N2081, N476);
buf BUF1 (N2106, N2105);
not NOT1 (N2107, N2106);
xor XOR2 (N2108, N2100, N1295);
and AND3 (N2109, N2102, N153, N1962);
nand NAND4 (N2110, N2109, N281, N1617, N1266);
buf BUF1 (N2111, N2104);
nand NAND2 (N2112, N2082, N1020);
and AND2 (N2113, N2103, N1049);
nand NAND4 (N2114, N2112, N288, N97, N2105);
or OR3 (N2115, N2108, N879, N1443);
nand NAND2 (N2116, N2114, N168);
and AND4 (N2117, N2098, N1724, N670, N856);
not NOT1 (N2118, N2116);
nor NOR3 (N2119, N2117, N352, N270);
buf BUF1 (N2120, N2083);
xor XOR2 (N2121, N2107, N696);
xor XOR2 (N2122, N2110, N987);
nor NOR4 (N2123, N2115, N1242, N129, N640);
nand NAND3 (N2124, N2113, N1253, N566);
nor NOR3 (N2125, N2121, N680, N1209);
xor XOR2 (N2126, N2118, N1640);
buf BUF1 (N2127, N2126);
not NOT1 (N2128, N2119);
buf BUF1 (N2129, N2128);
not NOT1 (N2130, N2124);
and AND2 (N2131, N2092, N199);
nand NAND3 (N2132, N2130, N986, N372);
and AND2 (N2133, N2123, N1735);
or OR2 (N2134, N2131, N617);
or OR2 (N2135, N2129, N1919);
and AND2 (N2136, N2096, N1406);
and AND2 (N2137, N2135, N1820);
nand NAND4 (N2138, N2137, N273, N1, N1092);
and AND3 (N2139, N2133, N128, N1066);
xor XOR2 (N2140, N2125, N1952);
nand NAND3 (N2141, N2127, N134, N102);
not NOT1 (N2142, N2111);
nand NAND2 (N2143, N2139, N149);
or OR2 (N2144, N2132, N330);
buf BUF1 (N2145, N2138);
xor XOR2 (N2146, N2136, N1966);
nor NOR2 (N2147, N2142, N747);
xor XOR2 (N2148, N2144, N1615);
xor XOR2 (N2149, N2122, N1701);
xor XOR2 (N2150, N2149, N1488);
not NOT1 (N2151, N2143);
xor XOR2 (N2152, N2148, N1374);
or OR3 (N2153, N2140, N492, N1299);
and AND4 (N2154, N2134, N313, N1746, N1657);
nand NAND4 (N2155, N2147, N358, N1562, N532);
not NOT1 (N2156, N2153);
not NOT1 (N2157, N2156);
and AND4 (N2158, N2157, N1021, N1934, N67);
or OR4 (N2159, N2155, N1270, N498, N1470);
xor XOR2 (N2160, N2151, N1904);
buf BUF1 (N2161, N2152);
and AND3 (N2162, N2154, N1077, N1578);
buf BUF1 (N2163, N2158);
or OR3 (N2164, N2146, N455, N2010);
buf BUF1 (N2165, N2162);
nor NOR2 (N2166, N2165, N1182);
xor XOR2 (N2167, N2164, N1734);
not NOT1 (N2168, N2166);
not NOT1 (N2169, N2145);
nand NAND4 (N2170, N2150, N1243, N2100, N92);
nor NOR2 (N2171, N2168, N1948);
nor NOR4 (N2172, N2169, N1241, N529, N772);
nor NOR2 (N2173, N2170, N553);
xor XOR2 (N2174, N2160, N509);
not NOT1 (N2175, N2172);
or OR4 (N2176, N2174, N461, N137, N1630);
nand NAND4 (N2177, N2161, N599, N1522, N1519);
xor XOR2 (N2178, N2159, N1318);
buf BUF1 (N2179, N2163);
or OR2 (N2180, N2167, N735);
nand NAND2 (N2181, N2120, N509);
buf BUF1 (N2182, N2141);
and AND2 (N2183, N2177, N93);
and AND2 (N2184, N2176, N1872);
buf BUF1 (N2185, N2171);
nor NOR4 (N2186, N2175, N1103, N1320, N1746);
nand NAND3 (N2187, N2180, N1623, N1850);
buf BUF1 (N2188, N2185);
nand NAND3 (N2189, N2178, N1831, N1212);
buf BUF1 (N2190, N2173);
xor XOR2 (N2191, N2183, N1425);
nor NOR2 (N2192, N2186, N991);
or OR3 (N2193, N2184, N1246, N1544);
xor XOR2 (N2194, N2191, N1135);
and AND3 (N2195, N2188, N2024, N207);
or OR3 (N2196, N2195, N1020, N200);
not NOT1 (N2197, N2194);
and AND2 (N2198, N2187, N1626);
xor XOR2 (N2199, N2192, N421);
or OR4 (N2200, N2179, N512, N882, N631);
nand NAND3 (N2201, N2196, N1122, N803);
nand NAND4 (N2202, N2198, N1181, N518, N1759);
nor NOR4 (N2203, N2190, N164, N1537, N1102);
and AND3 (N2204, N2202, N1265, N521);
or OR4 (N2205, N2199, N735, N1311, N2176);
or OR4 (N2206, N2189, N485, N755, N666);
nor NOR4 (N2207, N2200, N1725, N1381, N74);
buf BUF1 (N2208, N2203);
xor XOR2 (N2209, N2204, N497);
or OR4 (N2210, N2206, N383, N593, N99);
and AND3 (N2211, N2207, N1205, N991);
and AND2 (N2212, N2208, N711);
nor NOR4 (N2213, N2182, N1414, N125, N399);
and AND4 (N2214, N2212, N1547, N2162, N223);
and AND2 (N2215, N2181, N1439);
not NOT1 (N2216, N2193);
nand NAND3 (N2217, N2211, N1709, N1074);
nor NOR2 (N2218, N2201, N573);
nor NOR4 (N2219, N2217, N752, N1852, N150);
or OR4 (N2220, N2197, N1671, N1437, N1518);
buf BUF1 (N2221, N2219);
xor XOR2 (N2222, N2215, N1872);
or OR4 (N2223, N2214, N129, N1278, N1539);
nor NOR4 (N2224, N2213, N67, N138, N1935);
not NOT1 (N2225, N2223);
and AND2 (N2226, N2220, N672);
and AND3 (N2227, N2226, N1871, N1509);
and AND3 (N2228, N2227, N1598, N1826);
xor XOR2 (N2229, N2218, N529);
not NOT1 (N2230, N2225);
nor NOR2 (N2231, N2221, N1591);
or OR3 (N2232, N2205, N1556, N1226);
not NOT1 (N2233, N2210);
or OR4 (N2234, N2216, N1376, N780, N85);
nand NAND3 (N2235, N2234, N1837, N2030);
nand NAND2 (N2236, N2222, N1606);
buf BUF1 (N2237, N2236);
buf BUF1 (N2238, N2229);
xor XOR2 (N2239, N2209, N536);
not NOT1 (N2240, N2230);
and AND4 (N2241, N2240, N1854, N1022, N94);
not NOT1 (N2242, N2235);
not NOT1 (N2243, N2232);
and AND2 (N2244, N2233, N1526);
xor XOR2 (N2245, N2244, N1144);
nor NOR2 (N2246, N2231, N837);
nor NOR2 (N2247, N2239, N2201);
xor XOR2 (N2248, N2242, N730);
nand NAND4 (N2249, N2247, N2221, N308, N2011);
nor NOR2 (N2250, N2249, N2113);
nor NOR4 (N2251, N2237, N284, N1568, N1667);
or OR2 (N2252, N2224, N725);
and AND2 (N2253, N2243, N1038);
not NOT1 (N2254, N2250);
not NOT1 (N2255, N2241);
buf BUF1 (N2256, N2248);
not NOT1 (N2257, N2238);
not NOT1 (N2258, N2228);
and AND4 (N2259, N2245, N593, N382, N1998);
or OR4 (N2260, N2259, N862, N988, N2111);
nor NOR3 (N2261, N2246, N1249, N2114);
buf BUF1 (N2262, N2253);
and AND2 (N2263, N2260, N769);
or OR4 (N2264, N2252, N821, N876, N381);
not NOT1 (N2265, N2258);
or OR3 (N2266, N2254, N282, N942);
not NOT1 (N2267, N2264);
nor NOR3 (N2268, N2261, N871, N818);
and AND2 (N2269, N2257, N417);
xor XOR2 (N2270, N2265, N603);
xor XOR2 (N2271, N2256, N541);
nand NAND4 (N2272, N2266, N270, N894, N179);
buf BUF1 (N2273, N2271);
and AND3 (N2274, N2269, N1314, N1944);
or OR4 (N2275, N2267, N1303, N331, N426);
and AND3 (N2276, N2275, N1374, N1685);
nand NAND4 (N2277, N2268, N1711, N73, N988);
not NOT1 (N2278, N2270);
or OR2 (N2279, N2272, N726);
or OR2 (N2280, N2277, N1416);
not NOT1 (N2281, N2279);
or OR3 (N2282, N2273, N1892, N25);
or OR4 (N2283, N2255, N1464, N271, N1305);
and AND3 (N2284, N2280, N374, N2005);
and AND4 (N2285, N2281, N1883, N1024, N1960);
and AND2 (N2286, N2274, N1260);
xor XOR2 (N2287, N2263, N1483);
buf BUF1 (N2288, N2282);
or OR3 (N2289, N2262, N79, N984);
or OR4 (N2290, N2289, N1664, N255, N1409);
or OR3 (N2291, N2278, N1838, N2047);
and AND2 (N2292, N2276, N2278);
and AND2 (N2293, N2285, N331);
not NOT1 (N2294, N2251);
nor NOR4 (N2295, N2293, N1946, N121, N1394);
not NOT1 (N2296, N2287);
buf BUF1 (N2297, N2294);
buf BUF1 (N2298, N2283);
nor NOR4 (N2299, N2286, N1218, N2145, N1479);
not NOT1 (N2300, N2298);
nor NOR4 (N2301, N2297, N685, N699, N477);
xor XOR2 (N2302, N2292, N860);
nand NAND2 (N2303, N2295, N421);
or OR4 (N2304, N2299, N1897, N2052, N37);
xor XOR2 (N2305, N2300, N520);
xor XOR2 (N2306, N2303, N922);
not NOT1 (N2307, N2302);
xor XOR2 (N2308, N2307, N1206);
and AND2 (N2309, N2304, N637);
xor XOR2 (N2310, N2284, N90);
nand NAND3 (N2311, N2291, N87, N155);
buf BUF1 (N2312, N2305);
buf BUF1 (N2313, N2301);
not NOT1 (N2314, N2311);
nand NAND3 (N2315, N2296, N1775, N1015);
or OR2 (N2316, N2308, N665);
not NOT1 (N2317, N2312);
nor NOR2 (N2318, N2316, N1983);
nor NOR4 (N2319, N2314, N2168, N55, N2286);
or OR3 (N2320, N2319, N2122, N1202);
xor XOR2 (N2321, N2318, N291);
not NOT1 (N2322, N2310);
buf BUF1 (N2323, N2306);
not NOT1 (N2324, N2315);
or OR4 (N2325, N2324, N2212, N995, N1806);
xor XOR2 (N2326, N2317, N1938);
nor NOR4 (N2327, N2290, N1379, N262, N311);
nand NAND2 (N2328, N2323, N360);
buf BUF1 (N2329, N2322);
xor XOR2 (N2330, N2320, N715);
or OR4 (N2331, N2326, N1783, N717, N815);
or OR3 (N2332, N2309, N690, N2116);
nor NOR2 (N2333, N2332, N1728);
xor XOR2 (N2334, N2329, N1439);
buf BUF1 (N2335, N2325);
buf BUF1 (N2336, N2321);
nor NOR3 (N2337, N2330, N627, N2282);
not NOT1 (N2338, N2335);
not NOT1 (N2339, N2334);
nor NOR2 (N2340, N2337, N2316);
nand NAND2 (N2341, N2333, N2113);
or OR4 (N2342, N2340, N939, N32, N1763);
buf BUF1 (N2343, N2327);
or OR2 (N2344, N2328, N1202);
nand NAND3 (N2345, N2339, N2270, N1388);
buf BUF1 (N2346, N2338);
or OR4 (N2347, N2313, N1830, N1921, N646);
nor NOR3 (N2348, N2342, N1767, N582);
and AND4 (N2349, N2343, N120, N1326, N319);
xor XOR2 (N2350, N2336, N772);
xor XOR2 (N2351, N2341, N1385);
and AND3 (N2352, N2348, N77, N677);
xor XOR2 (N2353, N2351, N241);
or OR2 (N2354, N2350, N2265);
and AND2 (N2355, N2331, N839);
not NOT1 (N2356, N2344);
or OR4 (N2357, N2352, N1033, N1757, N479);
nor NOR3 (N2358, N2356, N1721, N1617);
buf BUF1 (N2359, N2355);
buf BUF1 (N2360, N2354);
nor NOR4 (N2361, N2353, N869, N1553, N1340);
xor XOR2 (N2362, N2359, N518);
buf BUF1 (N2363, N2288);
or OR3 (N2364, N2361, N210, N65);
nor NOR2 (N2365, N2349, N109);
or OR4 (N2366, N2365, N331, N254, N1400);
and AND3 (N2367, N2366, N193, N1140);
not NOT1 (N2368, N2362);
buf BUF1 (N2369, N2368);
buf BUF1 (N2370, N2345);
or OR3 (N2371, N2363, N1550, N2062);
nand NAND3 (N2372, N2370, N847, N889);
buf BUF1 (N2373, N2346);
not NOT1 (N2374, N2373);
and AND2 (N2375, N2357, N2280);
and AND3 (N2376, N2374, N2126, N1371);
nor NOR3 (N2377, N2371, N784, N484);
or OR4 (N2378, N2360, N1839, N119, N544);
not NOT1 (N2379, N2358);
nor NOR2 (N2380, N2375, N1347);
nor NOR3 (N2381, N2378, N10, N667);
buf BUF1 (N2382, N2364);
not NOT1 (N2383, N2381);
buf BUF1 (N2384, N2383);
nand NAND4 (N2385, N2384, N1165, N1761, N1165);
xor XOR2 (N2386, N2385, N1398);
not NOT1 (N2387, N2386);
nor NOR4 (N2388, N2377, N779, N1190, N638);
and AND2 (N2389, N2372, N2241);
buf BUF1 (N2390, N2376);
and AND2 (N2391, N2369, N1983);
nand NAND4 (N2392, N2390, N593, N1822, N1835);
or OR4 (N2393, N2387, N1688, N1842, N2222);
nor NOR3 (N2394, N2393, N1834, N2028);
xor XOR2 (N2395, N2388, N2178);
not NOT1 (N2396, N2380);
buf BUF1 (N2397, N2391);
xor XOR2 (N2398, N2347, N629);
or OR4 (N2399, N2392, N1716, N1566, N1987);
and AND2 (N2400, N2399, N895);
not NOT1 (N2401, N2397);
nor NOR2 (N2402, N2379, N1646);
nand NAND3 (N2403, N2367, N515, N1189);
nor NOR3 (N2404, N2400, N755, N201);
nor NOR4 (N2405, N2401, N829, N735, N1987);
nor NOR3 (N2406, N2405, N1070, N641);
xor XOR2 (N2407, N2396, N2049);
buf BUF1 (N2408, N2404);
not NOT1 (N2409, N2389);
and AND3 (N2410, N2409, N598, N1675);
or OR3 (N2411, N2402, N318, N2010);
not NOT1 (N2412, N2408);
xor XOR2 (N2413, N2407, N2239);
xor XOR2 (N2414, N2413, N169);
nand NAND2 (N2415, N2403, N1323);
not NOT1 (N2416, N2412);
not NOT1 (N2417, N2398);
not NOT1 (N2418, N2411);
and AND3 (N2419, N2415, N588, N811);
or OR3 (N2420, N2395, N1421, N2081);
buf BUF1 (N2421, N2414);
or OR2 (N2422, N2394, N1324);
nand NAND2 (N2423, N2406, N23);
and AND3 (N2424, N2420, N2080, N128);
nand NAND3 (N2425, N2424, N1582, N1411);
xor XOR2 (N2426, N2418, N1472);
and AND4 (N2427, N2410, N1315, N270, N1871);
or OR2 (N2428, N2419, N86);
nor NOR3 (N2429, N2426, N1845, N300);
nand NAND4 (N2430, N2382, N844, N1537, N693);
and AND3 (N2431, N2425, N1405, N2186);
buf BUF1 (N2432, N2417);
not NOT1 (N2433, N2430);
nor NOR2 (N2434, N2421, N1038);
nand NAND2 (N2435, N2432, N2098);
nor NOR2 (N2436, N2433, N900);
and AND3 (N2437, N2436, N363, N505);
xor XOR2 (N2438, N2416, N1878);
xor XOR2 (N2439, N2437, N2242);
nor NOR4 (N2440, N2428, N2068, N189, N630);
xor XOR2 (N2441, N2434, N685);
buf BUF1 (N2442, N2429);
buf BUF1 (N2443, N2422);
buf BUF1 (N2444, N2427);
xor XOR2 (N2445, N2443, N2313);
nor NOR4 (N2446, N2431, N2159, N1088, N1947);
or OR4 (N2447, N2446, N1914, N2301, N2360);
nor NOR3 (N2448, N2442, N116, N2000);
xor XOR2 (N2449, N2447, N2038);
nor NOR4 (N2450, N2444, N1624, N2355, N207);
or OR2 (N2451, N2449, N2392);
and AND2 (N2452, N2441, N1722);
nor NOR4 (N2453, N2440, N1477, N2097, N2320);
or OR3 (N2454, N2445, N994, N2090);
or OR3 (N2455, N2450, N1670, N1984);
buf BUF1 (N2456, N2435);
xor XOR2 (N2457, N2438, N1964);
buf BUF1 (N2458, N2457);
nand NAND4 (N2459, N2452, N2019, N1034, N15);
and AND2 (N2460, N2454, N854);
nor NOR3 (N2461, N2455, N2029, N1217);
not NOT1 (N2462, N2460);
not NOT1 (N2463, N2462);
or OR4 (N2464, N2439, N1498, N304, N165);
or OR4 (N2465, N2458, N70, N830, N1229);
buf BUF1 (N2466, N2461);
and AND3 (N2467, N2463, N1586, N738);
not NOT1 (N2468, N2459);
xor XOR2 (N2469, N2468, N2299);
nand NAND3 (N2470, N2469, N18, N425);
not NOT1 (N2471, N2456);
or OR4 (N2472, N2423, N1866, N935, N1615);
buf BUF1 (N2473, N2448);
and AND2 (N2474, N2470, N936);
nor NOR4 (N2475, N2472, N2451, N1529, N73);
xor XOR2 (N2476, N2148, N2069);
or OR3 (N2477, N2465, N1574, N1821);
nor NOR4 (N2478, N2471, N2184, N564, N1650);
or OR3 (N2479, N2477, N217, N996);
xor XOR2 (N2480, N2473, N2004);
buf BUF1 (N2481, N2475);
or OR2 (N2482, N2481, N994);
buf BUF1 (N2483, N2482);
buf BUF1 (N2484, N2478);
xor XOR2 (N2485, N2484, N2014);
nand NAND3 (N2486, N2485, N1882, N1541);
and AND4 (N2487, N2480, N1152, N1382, N1029);
not NOT1 (N2488, N2453);
buf BUF1 (N2489, N2483);
and AND4 (N2490, N2464, N890, N1459, N2087);
buf BUF1 (N2491, N2479);
nand NAND2 (N2492, N2466, N1155);
buf BUF1 (N2493, N2486);
and AND2 (N2494, N2467, N1902);
or OR4 (N2495, N2474, N1325, N233, N380);
xor XOR2 (N2496, N2493, N2423);
nor NOR2 (N2497, N2488, N853);
xor XOR2 (N2498, N2490, N2125);
and AND3 (N2499, N2496, N397, N611);
nor NOR3 (N2500, N2495, N271, N2370);
buf BUF1 (N2501, N2489);
nand NAND3 (N2502, N2487, N2186, N1253);
or OR3 (N2503, N2476, N2473, N1334);
nor NOR3 (N2504, N2492, N1687, N438);
xor XOR2 (N2505, N2499, N1220);
xor XOR2 (N2506, N2501, N1890);
nand NAND2 (N2507, N2497, N508);
buf BUF1 (N2508, N2505);
nand NAND2 (N2509, N2491, N125);
or OR2 (N2510, N2494, N2041);
xor XOR2 (N2511, N2507, N2263);
not NOT1 (N2512, N2510);
nand NAND3 (N2513, N2509, N254, N1618);
nand NAND2 (N2514, N2508, N918);
nor NOR2 (N2515, N2500, N2293);
buf BUF1 (N2516, N2511);
nor NOR4 (N2517, N2502, N1313, N248, N1177);
not NOT1 (N2518, N2513);
or OR2 (N2519, N2504, N2079);
or OR2 (N2520, N2517, N1700);
nand NAND4 (N2521, N2515, N127, N1144, N769);
xor XOR2 (N2522, N2514, N954);
xor XOR2 (N2523, N2512, N1272);
nor NOR2 (N2524, N2516, N1777);
nor NOR3 (N2525, N2524, N1784, N258);
not NOT1 (N2526, N2521);
and AND2 (N2527, N2526, N715);
buf BUF1 (N2528, N2527);
and AND3 (N2529, N2520, N1023, N1776);
nor NOR4 (N2530, N2518, N1303, N1331, N937);
buf BUF1 (N2531, N2522);
nor NOR3 (N2532, N2498, N988, N862);
buf BUF1 (N2533, N2519);
buf BUF1 (N2534, N2530);
nor NOR4 (N2535, N2532, N1970, N1106, N1340);
xor XOR2 (N2536, N2528, N1503);
and AND4 (N2537, N2503, N1762, N1845, N468);
xor XOR2 (N2538, N2523, N1216);
nor NOR4 (N2539, N2529, N1755, N376, N2264);
or OR3 (N2540, N2506, N1879, N2230);
nor NOR4 (N2541, N2525, N1642, N2262, N248);
and AND4 (N2542, N2531, N1156, N852, N1162);
nor NOR3 (N2543, N2535, N1395, N1561);
nand NAND4 (N2544, N2540, N964, N1632, N44);
nor NOR4 (N2545, N2539, N393, N811, N381);
buf BUF1 (N2546, N2534);
buf BUF1 (N2547, N2544);
nor NOR4 (N2548, N2538, N1852, N583, N2156);
and AND2 (N2549, N2547, N82);
nand NAND2 (N2550, N2549, N1099);
or OR2 (N2551, N2536, N1496);
nand NAND3 (N2552, N2548, N2434, N116);
nor NOR2 (N2553, N2552, N669);
and AND4 (N2554, N2550, N2192, N2084, N1677);
buf BUF1 (N2555, N2553);
nor NOR4 (N2556, N2546, N728, N1091, N1473);
nand NAND2 (N2557, N2555, N676);
nand NAND4 (N2558, N2542, N2287, N1417, N792);
or OR3 (N2559, N2551, N2091, N1653);
or OR4 (N2560, N2554, N2519, N1148, N1780);
xor XOR2 (N2561, N2545, N365);
xor XOR2 (N2562, N2556, N1208);
xor XOR2 (N2563, N2562, N186);
nor NOR3 (N2564, N2559, N1625, N676);
xor XOR2 (N2565, N2564, N2400);
xor XOR2 (N2566, N2560, N653);
xor XOR2 (N2567, N2533, N1571);
nor NOR2 (N2568, N2543, N2519);
or OR3 (N2569, N2565, N843, N2388);
buf BUF1 (N2570, N2557);
or OR2 (N2571, N2567, N136);
or OR2 (N2572, N2537, N452);
and AND3 (N2573, N2572, N1212, N9);
xor XOR2 (N2574, N2561, N1731);
and AND4 (N2575, N2568, N2110, N1884, N520);
xor XOR2 (N2576, N2558, N1264);
buf BUF1 (N2577, N2575);
xor XOR2 (N2578, N2569, N2478);
xor XOR2 (N2579, N2571, N911);
nor NOR2 (N2580, N2570, N473);
nand NAND2 (N2581, N2574, N1026);
not NOT1 (N2582, N2580);
and AND4 (N2583, N2578, N2348, N419, N2505);
and AND4 (N2584, N2581, N1445, N1564, N849);
not NOT1 (N2585, N2563);
nor NOR3 (N2586, N2541, N2583, N893);
or OR4 (N2587, N507, N1175, N2504, N1747);
buf BUF1 (N2588, N2582);
not NOT1 (N2589, N2584);
nand NAND3 (N2590, N2579, N342, N1843);
buf BUF1 (N2591, N2566);
buf BUF1 (N2592, N2588);
not NOT1 (N2593, N2573);
xor XOR2 (N2594, N2585, N248);
not NOT1 (N2595, N2594);
and AND3 (N2596, N2592, N106, N2333);
buf BUF1 (N2597, N2593);
not NOT1 (N2598, N2590);
buf BUF1 (N2599, N2576);
not NOT1 (N2600, N2598);
nor NOR2 (N2601, N2587, N2468);
nand NAND4 (N2602, N2601, N569, N1186, N1256);
nor NOR2 (N2603, N2596, N57);
xor XOR2 (N2604, N2603, N887);
or OR2 (N2605, N2577, N2334);
not NOT1 (N2606, N2602);
buf BUF1 (N2607, N2589);
buf BUF1 (N2608, N2607);
not NOT1 (N2609, N2595);
or OR2 (N2610, N2600, N1191);
nor NOR4 (N2611, N2599, N1146, N1079, N2116);
not NOT1 (N2612, N2604);
nand NAND2 (N2613, N2597, N1786);
nand NAND2 (N2614, N2586, N2522);
or OR3 (N2615, N2608, N1119, N1592);
nor NOR4 (N2616, N2610, N2326, N1839, N1216);
nor NOR2 (N2617, N2606, N1938);
not NOT1 (N2618, N2613);
nand NAND3 (N2619, N2611, N267, N1579);
nor NOR3 (N2620, N2617, N1117, N755);
buf BUF1 (N2621, N2615);
or OR2 (N2622, N2621, N2469);
buf BUF1 (N2623, N2591);
or OR3 (N2624, N2614, N792, N1929);
not NOT1 (N2625, N2622);
or OR4 (N2626, N2624, N2301, N2338, N1512);
not NOT1 (N2627, N2620);
or OR2 (N2628, N2619, N854);
and AND3 (N2629, N2616, N145, N1889);
and AND4 (N2630, N2618, N1942, N941, N2022);
xor XOR2 (N2631, N2629, N1248);
nor NOR2 (N2632, N2627, N1979);
nand NAND3 (N2633, N2632, N71, N2501);
and AND3 (N2634, N2612, N1842, N2319);
xor XOR2 (N2635, N2626, N1301);
xor XOR2 (N2636, N2630, N1136);
not NOT1 (N2637, N2635);
and AND2 (N2638, N2633, N2350);
and AND2 (N2639, N2636, N2614);
nor NOR3 (N2640, N2637, N2297, N892);
buf BUF1 (N2641, N2634);
or OR3 (N2642, N2623, N1868, N1316);
or OR2 (N2643, N2639, N965);
nor NOR3 (N2644, N2609, N2425, N587);
nand NAND4 (N2645, N2631, N2457, N255, N1943);
xor XOR2 (N2646, N2643, N1965);
xor XOR2 (N2647, N2642, N2411);
not NOT1 (N2648, N2647);
nand NAND4 (N2649, N2628, N1488, N2209, N1072);
not NOT1 (N2650, N2641);
and AND4 (N2651, N2625, N1392, N1664, N585);
or OR3 (N2652, N2646, N167, N1079);
xor XOR2 (N2653, N2605, N1084);
not NOT1 (N2654, N2645);
xor XOR2 (N2655, N2650, N614);
or OR3 (N2656, N2651, N1287, N2134);
nor NOR3 (N2657, N2652, N666, N2183);
xor XOR2 (N2658, N2644, N1438);
or OR4 (N2659, N2657, N1257, N414, N2087);
or OR4 (N2660, N2640, N1350, N1381, N2596);
nor NOR3 (N2661, N2656, N2327, N432);
xor XOR2 (N2662, N2648, N1713);
buf BUF1 (N2663, N2662);
xor XOR2 (N2664, N2663, N8);
and AND4 (N2665, N2653, N859, N2150, N894);
xor XOR2 (N2666, N2664, N2616);
buf BUF1 (N2667, N2654);
not NOT1 (N2668, N2658);
not NOT1 (N2669, N2649);
nand NAND3 (N2670, N2666, N595, N1344);
buf BUF1 (N2671, N2655);
nor NOR3 (N2672, N2667, N1907, N1018);
or OR2 (N2673, N2670, N1926);
not NOT1 (N2674, N2668);
xor XOR2 (N2675, N2661, N1187);
buf BUF1 (N2676, N2638);
nor NOR4 (N2677, N2660, N1821, N524, N2210);
and AND2 (N2678, N2675, N1491);
and AND2 (N2679, N2672, N110);
and AND2 (N2680, N2679, N962);
xor XOR2 (N2681, N2674, N534);
not NOT1 (N2682, N2659);
buf BUF1 (N2683, N2682);
and AND2 (N2684, N2665, N910);
not NOT1 (N2685, N2680);
xor XOR2 (N2686, N2676, N2128);
or OR3 (N2687, N2677, N767, N1801);
and AND4 (N2688, N2684, N1773, N2459, N1666);
buf BUF1 (N2689, N2687);
nor NOR3 (N2690, N2669, N483, N2586);
xor XOR2 (N2691, N2686, N251);
not NOT1 (N2692, N2681);
xor XOR2 (N2693, N2683, N254);
or OR2 (N2694, N2671, N615);
not NOT1 (N2695, N2690);
buf BUF1 (N2696, N2689);
nor NOR3 (N2697, N2693, N765, N1605);
and AND3 (N2698, N2696, N925, N260);
buf BUF1 (N2699, N2691);
xor XOR2 (N2700, N2688, N286);
or OR3 (N2701, N2697, N2290, N92);
nor NOR2 (N2702, N2699, N701);
or OR4 (N2703, N2701, N938, N888, N205);
or OR4 (N2704, N2685, N288, N252, N2600);
nand NAND4 (N2705, N2695, N1853, N969, N1784);
nor NOR2 (N2706, N2692, N2052);
xor XOR2 (N2707, N2703, N783);
not NOT1 (N2708, N2694);
buf BUF1 (N2709, N2702);
not NOT1 (N2710, N2708);
or OR3 (N2711, N2710, N2219, N841);
nor NOR2 (N2712, N2678, N807);
buf BUF1 (N2713, N2706);
or OR4 (N2714, N2705, N2467, N472, N376);
not NOT1 (N2715, N2698);
or OR3 (N2716, N2707, N2441, N693);
xor XOR2 (N2717, N2716, N695);
or OR2 (N2718, N2713, N2280);
or OR4 (N2719, N2709, N65, N2464, N455);
or OR3 (N2720, N2719, N1587, N247);
or OR4 (N2721, N2673, N1398, N2583, N100);
and AND3 (N2722, N2711, N492, N1599);
not NOT1 (N2723, N2721);
nand NAND3 (N2724, N2715, N1006, N1152);
not NOT1 (N2725, N2718);
nand NAND2 (N2726, N2723, N1321);
nor NOR3 (N2727, N2724, N1743, N110);
buf BUF1 (N2728, N2722);
buf BUF1 (N2729, N2720);
or OR4 (N2730, N2729, N2439, N1051, N658);
and AND4 (N2731, N2725, N2706, N995, N2124);
and AND2 (N2732, N2730, N1143);
nand NAND2 (N2733, N2732, N1078);
buf BUF1 (N2734, N2714);
nor NOR2 (N2735, N2717, N1246);
buf BUF1 (N2736, N2731);
and AND2 (N2737, N2728, N857);
nor NOR4 (N2738, N2736, N1152, N44, N949);
and AND3 (N2739, N2733, N1345, N837);
nand NAND2 (N2740, N2727, N2221);
buf BUF1 (N2741, N2740);
or OR3 (N2742, N2726, N42, N14);
and AND2 (N2743, N2700, N7);
not NOT1 (N2744, N2734);
and AND2 (N2745, N2704, N1577);
not NOT1 (N2746, N2742);
not NOT1 (N2747, N2735);
and AND4 (N2748, N2712, N2017, N290, N23);
nand NAND3 (N2749, N2737, N2676, N1604);
and AND3 (N2750, N2745, N1505, N1098);
buf BUF1 (N2751, N2739);
buf BUF1 (N2752, N2749);
buf BUF1 (N2753, N2752);
nand NAND2 (N2754, N2738, N2049);
or OR3 (N2755, N2744, N29, N1053);
nor NOR2 (N2756, N2755, N458);
and AND2 (N2757, N2748, N469);
and AND2 (N2758, N2741, N418);
buf BUF1 (N2759, N2750);
nor NOR3 (N2760, N2746, N178, N2563);
buf BUF1 (N2761, N2757);
nor NOR4 (N2762, N2753, N1743, N504, N2075);
nor NOR4 (N2763, N2759, N2761, N1469, N39);
nor NOR4 (N2764, N543, N218, N963, N2737);
nor NOR2 (N2765, N2760, N2360);
xor XOR2 (N2766, N2764, N1263);
xor XOR2 (N2767, N2747, N1971);
xor XOR2 (N2768, N2763, N940);
xor XOR2 (N2769, N2766, N1542);
xor XOR2 (N2770, N2754, N2572);
xor XOR2 (N2771, N2756, N1153);
or OR4 (N2772, N2743, N894, N981, N1136);
buf BUF1 (N2773, N2765);
not NOT1 (N2774, N2772);
and AND4 (N2775, N2762, N453, N554, N1859);
or OR4 (N2776, N2769, N930, N594, N1395);
not NOT1 (N2777, N2771);
or OR2 (N2778, N2770, N1368);
and AND2 (N2779, N2775, N1726);
and AND2 (N2780, N2779, N334);
not NOT1 (N2781, N2751);
xor XOR2 (N2782, N2774, N2335);
nor NOR3 (N2783, N2768, N356, N2233);
or OR2 (N2784, N2776, N2252);
and AND4 (N2785, N2773, N990, N2593, N1775);
xor XOR2 (N2786, N2778, N618);
buf BUF1 (N2787, N2777);
and AND2 (N2788, N2787, N2085);
buf BUF1 (N2789, N2780);
xor XOR2 (N2790, N2785, N226);
buf BUF1 (N2791, N2783);
not NOT1 (N2792, N2791);
not NOT1 (N2793, N2758);
and AND3 (N2794, N2782, N2665, N824);
xor XOR2 (N2795, N2788, N403);
not NOT1 (N2796, N2792);
not NOT1 (N2797, N2767);
not NOT1 (N2798, N2790);
buf BUF1 (N2799, N2798);
not NOT1 (N2800, N2789);
and AND3 (N2801, N2800, N38, N2265);
and AND4 (N2802, N2786, N146, N1986, N2322);
nand NAND4 (N2803, N2784, N538, N528, N52);
and AND4 (N2804, N2793, N699, N1344, N2438);
nor NOR2 (N2805, N2803, N470);
nor NOR3 (N2806, N2795, N2262, N2255);
not NOT1 (N2807, N2802);
not NOT1 (N2808, N2799);
and AND4 (N2809, N2781, N2702, N2006, N2245);
and AND4 (N2810, N2801, N1187, N539, N2563);
xor XOR2 (N2811, N2809, N1354);
or OR2 (N2812, N2808, N2313);
or OR2 (N2813, N2796, N2148);
or OR4 (N2814, N2807, N2214, N1556, N1716);
not NOT1 (N2815, N2806);
buf BUF1 (N2816, N2805);
or OR4 (N2817, N2815, N2204, N163, N1124);
or OR4 (N2818, N2814, N1993, N1930, N1387);
buf BUF1 (N2819, N2794);
nand NAND3 (N2820, N2812, N2639, N13);
and AND3 (N2821, N2819, N1168, N621);
and AND4 (N2822, N2813, N1862, N1236, N630);
not NOT1 (N2823, N2811);
and AND2 (N2824, N2822, N221);
xor XOR2 (N2825, N2823, N1023);
buf BUF1 (N2826, N2816);
or OR2 (N2827, N2818, N1020);
xor XOR2 (N2828, N2825, N2370);
nand NAND2 (N2829, N2817, N144);
buf BUF1 (N2830, N2826);
and AND4 (N2831, N2829, N1611, N246, N2055);
nand NAND2 (N2832, N2821, N2362);
buf BUF1 (N2833, N2830);
xor XOR2 (N2834, N2804, N995);
nor NOR3 (N2835, N2824, N2274, N2023);
nor NOR4 (N2836, N2831, N577, N100, N2526);
or OR3 (N2837, N2834, N1910, N1810);
nand NAND2 (N2838, N2828, N1911);
nor NOR3 (N2839, N2835, N1743, N461);
nand NAND3 (N2840, N2836, N586, N764);
and AND3 (N2841, N2840, N2357, N2209);
nor NOR2 (N2842, N2832, N1244);
nand NAND4 (N2843, N2837, N1393, N1629, N2344);
buf BUF1 (N2844, N2827);
xor XOR2 (N2845, N2843, N1413);
buf BUF1 (N2846, N2844);
or OR4 (N2847, N2810, N1442, N342, N991);
and AND4 (N2848, N2838, N1185, N1890, N1236);
nor NOR4 (N2849, N2846, N848, N361, N2638);
not NOT1 (N2850, N2833);
or OR2 (N2851, N2849, N686);
nand NAND2 (N2852, N2839, N2353);
buf BUF1 (N2853, N2847);
buf BUF1 (N2854, N2851);
not NOT1 (N2855, N2848);
xor XOR2 (N2856, N2845, N2315);
xor XOR2 (N2857, N2853, N1475);
xor XOR2 (N2858, N2820, N1245);
buf BUF1 (N2859, N2857);
xor XOR2 (N2860, N2842, N2766);
buf BUF1 (N2861, N2841);
nand NAND2 (N2862, N2856, N1230);
or OR2 (N2863, N2862, N333);
buf BUF1 (N2864, N2861);
nand NAND3 (N2865, N2797, N374, N2302);
nand NAND2 (N2866, N2863, N2241);
and AND2 (N2867, N2866, N1399);
nor NOR2 (N2868, N2854, N2469);
or OR4 (N2869, N2868, N257, N653, N2412);
buf BUF1 (N2870, N2850);
and AND2 (N2871, N2858, N606);
not NOT1 (N2872, N2859);
or OR2 (N2873, N2855, N2057);
buf BUF1 (N2874, N2852);
not NOT1 (N2875, N2860);
xor XOR2 (N2876, N2872, N558);
or OR3 (N2877, N2874, N1327, N216);
and AND4 (N2878, N2869, N1544, N706, N635);
nand NAND3 (N2879, N2870, N1496, N1790);
not NOT1 (N2880, N2875);
nor NOR3 (N2881, N2877, N1925, N796);
not NOT1 (N2882, N2867);
nor NOR4 (N2883, N2871, N2592, N1345, N453);
and AND2 (N2884, N2865, N2708);
not NOT1 (N2885, N2864);
buf BUF1 (N2886, N2884);
buf BUF1 (N2887, N2879);
nand NAND2 (N2888, N2878, N1974);
not NOT1 (N2889, N2880);
and AND2 (N2890, N2881, N2870);
not NOT1 (N2891, N2873);
and AND2 (N2892, N2882, N482);
buf BUF1 (N2893, N2892);
xor XOR2 (N2894, N2889, N1330);
nand NAND3 (N2895, N2891, N1535, N2665);
and AND4 (N2896, N2895, N1819, N1477, N2388);
and AND2 (N2897, N2893, N2611);
not NOT1 (N2898, N2888);
xor XOR2 (N2899, N2890, N959);
buf BUF1 (N2900, N2899);
nand NAND4 (N2901, N2885, N2193, N2355, N1430);
and AND2 (N2902, N2900, N1742);
or OR3 (N2903, N2898, N1776, N1450);
nand NAND2 (N2904, N2902, N2340);
not NOT1 (N2905, N2904);
not NOT1 (N2906, N2897);
not NOT1 (N2907, N2887);
nor NOR4 (N2908, N2883, N1603, N1040, N2381);
and AND4 (N2909, N2896, N839, N931, N593);
or OR3 (N2910, N2907, N2634, N1904);
nand NAND2 (N2911, N2886, N1984);
nor NOR3 (N2912, N2903, N363, N2698);
xor XOR2 (N2913, N2894, N1119);
nor NOR3 (N2914, N2912, N877, N873);
nand NAND4 (N2915, N2906, N433, N1525, N1461);
buf BUF1 (N2916, N2915);
not NOT1 (N2917, N2913);
not NOT1 (N2918, N2908);
and AND2 (N2919, N2901, N870);
buf BUF1 (N2920, N2919);
xor XOR2 (N2921, N2911, N2846);
and AND4 (N2922, N2876, N2580, N843, N1056);
buf BUF1 (N2923, N2917);
and AND2 (N2924, N2923, N1148);
and AND3 (N2925, N2910, N1088, N1595);
nand NAND3 (N2926, N2918, N862, N276);
nor NOR3 (N2927, N2914, N2568, N359);
not NOT1 (N2928, N2909);
and AND4 (N2929, N2920, N2730, N1884, N1639);
not NOT1 (N2930, N2924);
xor XOR2 (N2931, N2929, N475);
xor XOR2 (N2932, N2922, N1286);
or OR3 (N2933, N2928, N907, N904);
nand NAND3 (N2934, N2933, N2712, N853);
xor XOR2 (N2935, N2905, N1970);
not NOT1 (N2936, N2935);
buf BUF1 (N2937, N2926);
nand NAND4 (N2938, N2936, N2171, N482, N1484);
buf BUF1 (N2939, N2937);
buf BUF1 (N2940, N2921);
xor XOR2 (N2941, N2932, N1443);
and AND2 (N2942, N2934, N2931);
xor XOR2 (N2943, N1863, N875);
nand NAND3 (N2944, N2930, N810, N1153);
buf BUF1 (N2945, N2943);
buf BUF1 (N2946, N2940);
buf BUF1 (N2947, N2942);
nand NAND4 (N2948, N2946, N1026, N59, N455);
nand NAND2 (N2949, N2925, N2505);
not NOT1 (N2950, N2938);
nand NAND3 (N2951, N2916, N2035, N466);
buf BUF1 (N2952, N2949);
or OR4 (N2953, N2951, N1966, N1179, N1589);
buf BUF1 (N2954, N2939);
not NOT1 (N2955, N2953);
nor NOR3 (N2956, N2945, N447, N1945);
xor XOR2 (N2957, N2956, N2107);
nor NOR2 (N2958, N2941, N1970);
xor XOR2 (N2959, N2958, N1883);
nor NOR3 (N2960, N2959, N307, N1846);
buf BUF1 (N2961, N2952);
not NOT1 (N2962, N2957);
or OR2 (N2963, N2950, N1759);
or OR4 (N2964, N2948, N751, N980, N2021);
nand NAND4 (N2965, N2947, N934, N1231, N1663);
xor XOR2 (N2966, N2962, N2393);
buf BUF1 (N2967, N2944);
xor XOR2 (N2968, N2967, N2424);
xor XOR2 (N2969, N2961, N1821);
xor XOR2 (N2970, N2963, N2091);
xor XOR2 (N2971, N2964, N7);
buf BUF1 (N2972, N2955);
nor NOR2 (N2973, N2965, N1239);
nand NAND2 (N2974, N2972, N1853);
buf BUF1 (N2975, N2971);
xor XOR2 (N2976, N2975, N2111);
buf BUF1 (N2977, N2966);
and AND4 (N2978, N2973, N2319, N2293, N2291);
xor XOR2 (N2979, N2969, N2396);
nor NOR4 (N2980, N2968, N1523, N694, N1789);
nand NAND3 (N2981, N2978, N1671, N129);
not NOT1 (N2982, N2979);
and AND3 (N2983, N2960, N1989, N14);
xor XOR2 (N2984, N2977, N2053);
nor NOR4 (N2985, N2974, N1449, N2087, N2651);
nor NOR4 (N2986, N2927, N2447, N1409, N394);
or OR3 (N2987, N2954, N2817, N250);
or OR4 (N2988, N2981, N2867, N1819, N282);
nand NAND4 (N2989, N2983, N2371, N739, N224);
nor NOR2 (N2990, N2985, N614);
not NOT1 (N2991, N2986);
nor NOR4 (N2992, N2970, N2853, N726, N502);
and AND3 (N2993, N2980, N2818, N2204);
or OR2 (N2994, N2987, N1886);
buf BUF1 (N2995, N2991);
nand NAND2 (N2996, N2990, N19);
not NOT1 (N2997, N2992);
xor XOR2 (N2998, N2989, N510);
buf BUF1 (N2999, N2984);
or OR3 (N3000, N2996, N200, N1871);
not NOT1 (N3001, N2995);
buf BUF1 (N3002, N2988);
and AND2 (N3003, N3001, N1369);
or OR4 (N3004, N2982, N2448, N1735, N929);
and AND4 (N3005, N3003, N2082, N2282, N305);
or OR2 (N3006, N3002, N1961);
nand NAND3 (N3007, N3000, N823, N2225);
and AND4 (N3008, N3007, N2080, N21, N2375);
and AND2 (N3009, N2999, N1087);
nor NOR3 (N3010, N3005, N354, N2212);
not NOT1 (N3011, N3006);
or OR4 (N3012, N3008, N2195, N571, N1432);
and AND4 (N3013, N3004, N1646, N2523, N2432);
and AND3 (N3014, N3010, N1241, N195);
nor NOR3 (N3015, N3009, N498, N464);
xor XOR2 (N3016, N3012, N50);
and AND3 (N3017, N3011, N85, N2367);
not NOT1 (N3018, N2976);
nand NAND3 (N3019, N3014, N1520, N1181);
and AND4 (N3020, N3017, N798, N2967, N908);
nand NAND4 (N3021, N3016, N1141, N123, N680);
not NOT1 (N3022, N3018);
xor XOR2 (N3023, N2994, N2151);
buf BUF1 (N3024, N3022);
nand NAND3 (N3025, N2997, N1580, N2074);
and AND4 (N3026, N2998, N2365, N1104, N729);
xor XOR2 (N3027, N3019, N465);
buf BUF1 (N3028, N3020);
nor NOR4 (N3029, N3023, N1990, N1229, N1229);
nand NAND2 (N3030, N3013, N1830);
and AND3 (N3031, N2993, N1738, N264);
xor XOR2 (N3032, N3024, N1341);
or OR4 (N3033, N3015, N2167, N2605, N1517);
not NOT1 (N3034, N3029);
buf BUF1 (N3035, N3026);
buf BUF1 (N3036, N3033);
buf BUF1 (N3037, N3032);
nand NAND4 (N3038, N3036, N594, N2934, N1029);
or OR2 (N3039, N3038, N1287);
or OR3 (N3040, N3027, N275, N1858);
or OR2 (N3041, N3021, N1598);
nand NAND4 (N3042, N3028, N2228, N315, N668);
buf BUF1 (N3043, N3042);
and AND3 (N3044, N3025, N3011, N123);
nor NOR4 (N3045, N3037, N1889, N337, N188);
xor XOR2 (N3046, N3035, N1332);
xor XOR2 (N3047, N3044, N2941);
nand NAND4 (N3048, N3043, N2047, N1033, N159);
xor XOR2 (N3049, N3045, N2536);
nand NAND2 (N3050, N3031, N2823);
or OR4 (N3051, N3041, N2854, N2295, N245);
and AND2 (N3052, N3039, N783);
not NOT1 (N3053, N3030);
not NOT1 (N3054, N3048);
and AND4 (N3055, N3046, N710, N1199, N2362);
or OR2 (N3056, N3049, N804);
not NOT1 (N3057, N3051);
or OR2 (N3058, N3040, N52);
and AND4 (N3059, N3034, N381, N1336, N2783);
nand NAND4 (N3060, N3052, N1950, N2461, N2980);
not NOT1 (N3061, N3057);
nor NOR4 (N3062, N3050, N2654, N2417, N170);
or OR2 (N3063, N3058, N2941);
or OR3 (N3064, N3060, N2474, N2489);
nor NOR4 (N3065, N3055, N2266, N671, N2273);
not NOT1 (N3066, N3053);
or OR2 (N3067, N3056, N2399);
xor XOR2 (N3068, N3054, N389);
buf BUF1 (N3069, N3061);
and AND3 (N3070, N3064, N642, N470);
xor XOR2 (N3071, N3047, N1330);
nor NOR2 (N3072, N3068, N1294);
xor XOR2 (N3073, N3063, N3003);
xor XOR2 (N3074, N3059, N1763);
or OR3 (N3075, N3074, N2197, N912);
buf BUF1 (N3076, N3072);
nor NOR4 (N3077, N3071, N2042, N1430, N1472);
nor NOR4 (N3078, N3070, N768, N2725, N688);
nand NAND3 (N3079, N3067, N2647, N479);
buf BUF1 (N3080, N3076);
and AND3 (N3081, N3073, N701, N544);
not NOT1 (N3082, N3081);
and AND4 (N3083, N3065, N2638, N354, N483);
nand NAND4 (N3084, N3075, N728, N1938, N1901);
or OR3 (N3085, N3069, N37, N702);
nand NAND4 (N3086, N3083, N120, N1047, N1049);
not NOT1 (N3087, N3086);
nand NAND3 (N3088, N3066, N2479, N517);
not NOT1 (N3089, N3078);
nand NAND3 (N3090, N3089, N1426, N2492);
or OR4 (N3091, N3077, N1899, N449, N591);
not NOT1 (N3092, N3088);
buf BUF1 (N3093, N3079);
or OR4 (N3094, N3062, N1109, N2001, N1802);
buf BUF1 (N3095, N3085);
nand NAND4 (N3096, N3092, N767, N756, N62);
and AND3 (N3097, N3091, N775, N362);
nand NAND3 (N3098, N3084, N1950, N2029);
not NOT1 (N3099, N3097);
xor XOR2 (N3100, N3080, N2158);
or OR4 (N3101, N3095, N2429, N280, N3066);
buf BUF1 (N3102, N3100);
xor XOR2 (N3103, N3096, N2787);
not NOT1 (N3104, N3101);
and AND2 (N3105, N3094, N2981);
or OR3 (N3106, N3093, N2579, N2549);
nand NAND2 (N3107, N3105, N342);
nand NAND3 (N3108, N3103, N589, N143);
nor NOR2 (N3109, N3107, N1919);
and AND4 (N3110, N3099, N2394, N2655, N1061);
nor NOR2 (N3111, N3110, N2896);
or OR2 (N3112, N3098, N2046);
or OR4 (N3113, N3106, N2321, N2008, N1506);
nor NOR4 (N3114, N3108, N2385, N1840, N1950);
and AND4 (N3115, N3102, N2443, N248, N534);
buf BUF1 (N3116, N3109);
not NOT1 (N3117, N3114);
nor NOR2 (N3118, N3090, N2416);
and AND3 (N3119, N3118, N2495, N2045);
nor NOR2 (N3120, N3113, N1184);
nand NAND2 (N3121, N3111, N2748);
xor XOR2 (N3122, N3117, N1349);
nor NOR3 (N3123, N3104, N2433, N2456);
not NOT1 (N3124, N3112);
nand NAND4 (N3125, N3122, N2246, N251, N2925);
xor XOR2 (N3126, N3120, N1426);
nand NAND3 (N3127, N3116, N92, N1201);
nand NAND2 (N3128, N3115, N2011);
and AND2 (N3129, N3124, N2348);
nand NAND3 (N3130, N3127, N2575, N2948);
or OR2 (N3131, N3126, N1050);
nor NOR3 (N3132, N3131, N1083, N2469);
not NOT1 (N3133, N3082);
nor NOR2 (N3134, N3125, N98);
not NOT1 (N3135, N3132);
and AND2 (N3136, N3119, N2024);
or OR3 (N3137, N3134, N2023, N900);
not NOT1 (N3138, N3136);
or OR4 (N3139, N3130, N114, N2263, N1751);
nand NAND2 (N3140, N3133, N655);
buf BUF1 (N3141, N3139);
xor XOR2 (N3142, N3135, N1722);
and AND4 (N3143, N3140, N2538, N900, N2052);
or OR2 (N3144, N3137, N1299);
not NOT1 (N3145, N3129);
or OR3 (N3146, N3121, N725, N3111);
not NOT1 (N3147, N3146);
not NOT1 (N3148, N3138);
and AND4 (N3149, N3145, N2393, N1635, N1726);
and AND4 (N3150, N3141, N2608, N839, N1776);
buf BUF1 (N3151, N3150);
not NOT1 (N3152, N3147);
xor XOR2 (N3153, N3152, N2313);
or OR2 (N3154, N3128, N1175);
not NOT1 (N3155, N3123);
and AND4 (N3156, N3148, N2734, N724, N2849);
not NOT1 (N3157, N3144);
and AND3 (N3158, N3149, N2576, N2491);
nor NOR4 (N3159, N3142, N410, N1796, N625);
or OR3 (N3160, N3157, N243, N2194);
nand NAND4 (N3161, N3143, N2669, N2005, N2545);
or OR3 (N3162, N3155, N2133, N1059);
and AND4 (N3163, N3158, N396, N1149, N1527);
or OR3 (N3164, N3153, N242, N3027);
and AND3 (N3165, N3087, N1968, N3035);
nand NAND2 (N3166, N3163, N110);
buf BUF1 (N3167, N3160);
buf BUF1 (N3168, N3151);
nand NAND2 (N3169, N3156, N382);
nand NAND3 (N3170, N3159, N2022, N694);
nand NAND4 (N3171, N3161, N1562, N1021, N2657);
or OR4 (N3172, N3167, N720, N651, N2335);
or OR4 (N3173, N3172, N1272, N681, N2839);
buf BUF1 (N3174, N3168);
nand NAND2 (N3175, N3162, N612);
buf BUF1 (N3176, N3175);
not NOT1 (N3177, N3176);
buf BUF1 (N3178, N3170);
xor XOR2 (N3179, N3174, N2141);
or OR3 (N3180, N3166, N3131, N31);
nor NOR4 (N3181, N3165, N1359, N1255, N85);
not NOT1 (N3182, N3180);
nand NAND3 (N3183, N3171, N49, N21);
and AND2 (N3184, N3181, N1657);
buf BUF1 (N3185, N3164);
or OR4 (N3186, N3184, N1971, N239, N428);
buf BUF1 (N3187, N3182);
xor XOR2 (N3188, N3185, N2125);
and AND3 (N3189, N3187, N3050, N1965);
xor XOR2 (N3190, N3186, N960);
buf BUF1 (N3191, N3179);
and AND4 (N3192, N3190, N1547, N2747, N2346);
nand NAND3 (N3193, N3192, N2789, N735);
nor NOR2 (N3194, N3177, N1554);
not NOT1 (N3195, N3189);
nor NOR4 (N3196, N3188, N2189, N2242, N1703);
not NOT1 (N3197, N3193);
nand NAND3 (N3198, N3178, N2820, N1111);
nor NOR2 (N3199, N3196, N2871);
nand NAND3 (N3200, N3169, N3016, N1288);
xor XOR2 (N3201, N3154, N1636);
nand NAND4 (N3202, N3173, N757, N2421, N1661);
not NOT1 (N3203, N3197);
nor NOR3 (N3204, N3201, N1458, N1017);
or OR3 (N3205, N3198, N121, N2245);
nor NOR2 (N3206, N3183, N50);
not NOT1 (N3207, N3194);
not NOT1 (N3208, N3207);
not NOT1 (N3209, N3200);
xor XOR2 (N3210, N3202, N750);
nor NOR4 (N3211, N3204, N29, N3076, N3194);
and AND2 (N3212, N3195, N909);
or OR3 (N3213, N3206, N2362, N2031);
not NOT1 (N3214, N3203);
nand NAND2 (N3215, N3205, N2864);
and AND4 (N3216, N3199, N1230, N327, N107);
buf BUF1 (N3217, N3211);
or OR4 (N3218, N3213, N280, N2111, N733);
not NOT1 (N3219, N3214);
nand NAND3 (N3220, N3218, N1212, N1825);
not NOT1 (N3221, N3215);
or OR3 (N3222, N3191, N2384, N1633);
xor XOR2 (N3223, N3216, N990);
or OR4 (N3224, N3210, N2434, N2840, N359);
or OR4 (N3225, N3212, N3049, N227, N650);
not NOT1 (N3226, N3217);
and AND4 (N3227, N3221, N489, N2699, N56);
xor XOR2 (N3228, N3219, N1590);
nor NOR3 (N3229, N3228, N3029, N1771);
and AND4 (N3230, N3225, N1932, N3160, N1905);
buf BUF1 (N3231, N3227);
buf BUF1 (N3232, N3222);
not NOT1 (N3233, N3220);
or OR4 (N3234, N3226, N762, N1868, N1111);
and AND2 (N3235, N3231, N649);
nor NOR3 (N3236, N3224, N2287, N1322);
nor NOR4 (N3237, N3236, N1866, N1865, N286);
xor XOR2 (N3238, N3208, N810);
or OR2 (N3239, N3234, N291);
xor XOR2 (N3240, N3230, N617);
nor NOR2 (N3241, N3240, N1547);
buf BUF1 (N3242, N3238);
not NOT1 (N3243, N3241);
xor XOR2 (N3244, N3233, N777);
not NOT1 (N3245, N3209);
buf BUF1 (N3246, N3244);
or OR4 (N3247, N3235, N2552, N548, N1466);
xor XOR2 (N3248, N3242, N1501);
nor NOR2 (N3249, N3229, N1246);
xor XOR2 (N3250, N3223, N2797);
xor XOR2 (N3251, N3245, N218);
not NOT1 (N3252, N3250);
nand NAND3 (N3253, N3237, N412, N1949);
nor NOR4 (N3254, N3248, N1955, N2009, N1700);
buf BUF1 (N3255, N3253);
nor NOR3 (N3256, N3255, N1094, N1758);
and AND4 (N3257, N3239, N289, N996, N1778);
not NOT1 (N3258, N3247);
not NOT1 (N3259, N3251);
not NOT1 (N3260, N3258);
nand NAND2 (N3261, N3249, N209);
nor NOR2 (N3262, N3254, N3172);
nand NAND3 (N3263, N3260, N1187, N1479);
xor XOR2 (N3264, N3252, N447);
xor XOR2 (N3265, N3232, N111);
nand NAND3 (N3266, N3264, N2501, N2344);
and AND3 (N3267, N3266, N1510, N60);
nor NOR3 (N3268, N3246, N2476, N241);
xor XOR2 (N3269, N3256, N2533);
xor XOR2 (N3270, N3261, N417);
buf BUF1 (N3271, N3243);
and AND3 (N3272, N3267, N2456, N3035);
nand NAND3 (N3273, N3271, N1988, N2488);
xor XOR2 (N3274, N3257, N592);
not NOT1 (N3275, N3262);
nor NOR2 (N3276, N3274, N86);
xor XOR2 (N3277, N3269, N2225);
nand NAND2 (N3278, N3263, N1381);
not NOT1 (N3279, N3273);
not NOT1 (N3280, N3259);
buf BUF1 (N3281, N3278);
buf BUF1 (N3282, N3280);
or OR3 (N3283, N3279, N2461, N3070);
nand NAND3 (N3284, N3275, N2160, N503);
not NOT1 (N3285, N3283);
not NOT1 (N3286, N3277);
or OR2 (N3287, N3286, N779);
nor NOR2 (N3288, N3268, N2067);
buf BUF1 (N3289, N3272);
or OR2 (N3290, N3289, N160);
and AND2 (N3291, N3281, N3071);
buf BUF1 (N3292, N3287);
nor NOR2 (N3293, N3276, N1451);
nand NAND2 (N3294, N3265, N1109);
nor NOR4 (N3295, N3284, N248, N300, N1157);
not NOT1 (N3296, N3288);
nand NAND3 (N3297, N3285, N2505, N2889);
or OR4 (N3298, N3291, N655, N2377, N839);
nand NAND4 (N3299, N3270, N3195, N2067, N182);
and AND3 (N3300, N3295, N2702, N651);
buf BUF1 (N3301, N3282);
nor NOR3 (N3302, N3292, N537, N820);
nand NAND2 (N3303, N3302, N2372);
or OR4 (N3304, N3298, N770, N3132, N1111);
and AND4 (N3305, N3300, N792, N1597, N1437);
xor XOR2 (N3306, N3296, N1859);
xor XOR2 (N3307, N3294, N2637);
nand NAND4 (N3308, N3303, N800, N3169, N710);
or OR2 (N3309, N3308, N1423);
or OR3 (N3310, N3293, N1560, N3253);
and AND2 (N3311, N3290, N1227);
and AND2 (N3312, N3306, N175);
nor NOR3 (N3313, N3304, N3291, N3071);
buf BUF1 (N3314, N3299);
xor XOR2 (N3315, N3305, N276);
nand NAND3 (N3316, N3301, N2004, N1414);
not NOT1 (N3317, N3316);
or OR3 (N3318, N3311, N1908, N3158);
not NOT1 (N3319, N3312);
or OR2 (N3320, N3318, N330);
and AND2 (N3321, N3313, N1438);
buf BUF1 (N3322, N3314);
xor XOR2 (N3323, N3320, N3132);
xor XOR2 (N3324, N3319, N698);
nor NOR4 (N3325, N3324, N2334, N3195, N872);
not NOT1 (N3326, N3321);
or OR2 (N3327, N3326, N1542);
buf BUF1 (N3328, N3315);
and AND3 (N3329, N3322, N1258, N1975);
and AND3 (N3330, N3328, N3034, N903);
not NOT1 (N3331, N3297);
xor XOR2 (N3332, N3327, N2699);
or OR2 (N3333, N3310, N2039);
and AND4 (N3334, N3307, N1082, N3135, N1123);
xor XOR2 (N3335, N3334, N1061);
not NOT1 (N3336, N3333);
or OR2 (N3337, N3332, N1714);
buf BUF1 (N3338, N3317);
not NOT1 (N3339, N3337);
or OR2 (N3340, N3336, N1687);
not NOT1 (N3341, N3331);
not NOT1 (N3342, N3309);
and AND4 (N3343, N3330, N777, N2442, N431);
buf BUF1 (N3344, N3325);
or OR2 (N3345, N3335, N2486);
nor NOR2 (N3346, N3323, N2350);
or OR3 (N3347, N3340, N1691, N966);
buf BUF1 (N3348, N3345);
nand NAND2 (N3349, N3338, N1457);
or OR3 (N3350, N3343, N850, N2247);
and AND2 (N3351, N3344, N1876);
buf BUF1 (N3352, N3346);
not NOT1 (N3353, N3329);
or OR3 (N3354, N3341, N421, N2714);
not NOT1 (N3355, N3342);
xor XOR2 (N3356, N3347, N578);
nor NOR2 (N3357, N3348, N2903);
and AND3 (N3358, N3351, N3269, N2749);
buf BUF1 (N3359, N3339);
and AND2 (N3360, N3355, N2495);
xor XOR2 (N3361, N3358, N2773);
nor NOR3 (N3362, N3353, N1744, N420);
xor XOR2 (N3363, N3354, N3335);
nand NAND3 (N3364, N3349, N1744, N2196);
xor XOR2 (N3365, N3350, N1374);
nor NOR4 (N3366, N3362, N2968, N936, N1745);
or OR2 (N3367, N3356, N756);
or OR3 (N3368, N3366, N2574, N181);
buf BUF1 (N3369, N3357);
nor NOR2 (N3370, N3361, N2873);
or OR3 (N3371, N3370, N650, N1771);
nand NAND2 (N3372, N3369, N1123);
nor NOR2 (N3373, N3371, N835);
nor NOR4 (N3374, N3359, N862, N1385, N3173);
not NOT1 (N3375, N3374);
buf BUF1 (N3376, N3372);
buf BUF1 (N3377, N3367);
xor XOR2 (N3378, N3364, N1462);
not NOT1 (N3379, N3377);
buf BUF1 (N3380, N3363);
and AND4 (N3381, N3373, N2942, N1027, N251);
nand NAND2 (N3382, N3380, N2789);
xor XOR2 (N3383, N3368, N2649);
xor XOR2 (N3384, N3378, N2525);
not NOT1 (N3385, N3381);
or OR2 (N3386, N3352, N2131);
not NOT1 (N3387, N3384);
xor XOR2 (N3388, N3365, N1789);
not NOT1 (N3389, N3387);
not NOT1 (N3390, N3375);
buf BUF1 (N3391, N3385);
nor NOR3 (N3392, N3376, N1455, N445);
buf BUF1 (N3393, N3389);
or OR3 (N3394, N3393, N2054, N3007);
or OR2 (N3395, N3388, N559);
or OR3 (N3396, N3379, N2370, N2571);
buf BUF1 (N3397, N3390);
buf BUF1 (N3398, N3383);
not NOT1 (N3399, N3394);
buf BUF1 (N3400, N3396);
and AND3 (N3401, N3399, N2363, N1076);
not NOT1 (N3402, N3382);
nand NAND2 (N3403, N3395, N3268);
nor NOR3 (N3404, N3403, N1503, N232);
not NOT1 (N3405, N3402);
xor XOR2 (N3406, N3392, N3402);
or OR4 (N3407, N3406, N3364, N615, N2826);
not NOT1 (N3408, N3397);
or OR4 (N3409, N3404, N1433, N2451, N2914);
buf BUF1 (N3410, N3386);
and AND4 (N3411, N3408, N3113, N1473, N508);
not NOT1 (N3412, N3410);
not NOT1 (N3413, N3405);
nor NOR4 (N3414, N3398, N2630, N648, N56);
or OR4 (N3415, N3391, N3412, N2445, N1393);
not NOT1 (N3416, N2927);
xor XOR2 (N3417, N3415, N1923);
xor XOR2 (N3418, N3413, N314);
xor XOR2 (N3419, N3400, N1751);
or OR4 (N3420, N3360, N604, N975, N2517);
not NOT1 (N3421, N3411);
and AND2 (N3422, N3419, N3121);
not NOT1 (N3423, N3417);
nand NAND2 (N3424, N3422, N3332);
nor NOR2 (N3425, N3418, N3332);
and AND4 (N3426, N3420, N2734, N2281, N2124);
buf BUF1 (N3427, N3424);
xor XOR2 (N3428, N3423, N2698);
or OR4 (N3429, N3409, N2041, N195, N277);
and AND3 (N3430, N3425, N2704, N337);
xor XOR2 (N3431, N3430, N3208);
or OR3 (N3432, N3428, N2326, N2550);
nor NOR4 (N3433, N3416, N2107, N2981, N1108);
buf BUF1 (N3434, N3407);
nand NAND3 (N3435, N3429, N2315, N1514);
nand NAND4 (N3436, N3421, N345, N2389, N676);
not NOT1 (N3437, N3414);
nor NOR2 (N3438, N3434, N1104);
not NOT1 (N3439, N3436);
xor XOR2 (N3440, N3438, N3323);
nor NOR2 (N3441, N3426, N774);
buf BUF1 (N3442, N3437);
nor NOR3 (N3443, N3435, N2143, N2115);
nor NOR4 (N3444, N3443, N1684, N3425, N1317);
xor XOR2 (N3445, N3444, N743);
and AND2 (N3446, N3440, N2764);
xor XOR2 (N3447, N3441, N34);
buf BUF1 (N3448, N3431);
or OR2 (N3449, N3427, N2888);
and AND2 (N3450, N3447, N840);
nor NOR4 (N3451, N3433, N2642, N2429, N1560);
xor XOR2 (N3452, N3450, N1506);
nor NOR3 (N3453, N3401, N818, N2202);
and AND3 (N3454, N3449, N2385, N631);
xor XOR2 (N3455, N3448, N137);
nand NAND3 (N3456, N3439, N804, N1506);
and AND2 (N3457, N3445, N365);
nand NAND2 (N3458, N3432, N908);
nand NAND4 (N3459, N3456, N2874, N2205, N2584);
not NOT1 (N3460, N3452);
and AND2 (N3461, N3454, N67);
xor XOR2 (N3462, N3459, N3180);
buf BUF1 (N3463, N3458);
buf BUF1 (N3464, N3446);
nor NOR2 (N3465, N3457, N2312);
nor NOR3 (N3466, N3442, N1580, N3001);
not NOT1 (N3467, N3466);
and AND2 (N3468, N3467, N1171);
and AND4 (N3469, N3468, N3137, N2550, N889);
nand NAND4 (N3470, N3465, N2336, N726, N208);
and AND4 (N3471, N3455, N1442, N2995, N1902);
xor XOR2 (N3472, N3461, N3413);
and AND3 (N3473, N3453, N1922, N235);
xor XOR2 (N3474, N3469, N135);
or OR2 (N3475, N3472, N781);
nor NOR3 (N3476, N3474, N1972, N3090);
and AND2 (N3477, N3476, N1209);
not NOT1 (N3478, N3477);
xor XOR2 (N3479, N3471, N68);
not NOT1 (N3480, N3473);
nor NOR4 (N3481, N3464, N1235, N2803, N2118);
xor XOR2 (N3482, N3470, N1954);
xor XOR2 (N3483, N3463, N2353);
buf BUF1 (N3484, N3460);
or OR2 (N3485, N3475, N2030);
and AND3 (N3486, N3480, N2145, N2877);
xor XOR2 (N3487, N3485, N2822);
nand NAND4 (N3488, N3482, N2728, N2671, N3282);
and AND3 (N3489, N3487, N2977, N662);
xor XOR2 (N3490, N3489, N317);
nand NAND2 (N3491, N3478, N1376);
or OR3 (N3492, N3483, N1300, N1499);
not NOT1 (N3493, N3451);
nor NOR2 (N3494, N3479, N2681);
nand NAND2 (N3495, N3462, N3386);
xor XOR2 (N3496, N3494, N1521);
not NOT1 (N3497, N3491);
or OR3 (N3498, N3493, N858, N2091);
buf BUF1 (N3499, N3481);
and AND2 (N3500, N3497, N2638);
xor XOR2 (N3501, N3498, N2335);
nand NAND3 (N3502, N3496, N1946, N2284);
or OR2 (N3503, N3502, N2479);
and AND4 (N3504, N3495, N1580, N381, N2452);
buf BUF1 (N3505, N3490);
buf BUF1 (N3506, N3499);
xor XOR2 (N3507, N3492, N1851);
buf BUF1 (N3508, N3488);
xor XOR2 (N3509, N3507, N2421);
nand NAND4 (N3510, N3503, N2209, N3127, N274);
and AND4 (N3511, N3500, N21, N2651, N410);
nand NAND4 (N3512, N3501, N2788, N2209, N929);
and AND4 (N3513, N3505, N3294, N2444, N1039);
buf BUF1 (N3514, N3508);
xor XOR2 (N3515, N3514, N481);
not NOT1 (N3516, N3486);
or OR3 (N3517, N3504, N2182, N1505);
buf BUF1 (N3518, N3511);
nand NAND3 (N3519, N3506, N3453, N1810);
not NOT1 (N3520, N3513);
buf BUF1 (N3521, N3512);
and AND2 (N3522, N3518, N3151);
xor XOR2 (N3523, N3519, N1718);
xor XOR2 (N3524, N3516, N2029);
and AND4 (N3525, N3523, N626, N2353, N2479);
buf BUF1 (N3526, N3517);
or OR2 (N3527, N3521, N204);
nand NAND4 (N3528, N3527, N2285, N2736, N1347);
and AND4 (N3529, N3515, N3097, N453, N2149);
nor NOR3 (N3530, N3528, N2551, N3356);
nor NOR4 (N3531, N3510, N3168, N2345, N1128);
buf BUF1 (N3532, N3530);
xor XOR2 (N3533, N3524, N595);
not NOT1 (N3534, N3522);
buf BUF1 (N3535, N3520);
or OR4 (N3536, N3534, N2344, N2154, N722);
or OR3 (N3537, N3529, N2238, N654);
buf BUF1 (N3538, N3526);
buf BUF1 (N3539, N3536);
not NOT1 (N3540, N3533);
nor NOR4 (N3541, N3531, N226, N3460, N1562);
nand NAND3 (N3542, N3539, N2831, N239);
not NOT1 (N3543, N3525);
xor XOR2 (N3544, N3542, N1539);
or OR4 (N3545, N3541, N1252, N2249, N445);
not NOT1 (N3546, N3535);
xor XOR2 (N3547, N3537, N2126);
nor NOR2 (N3548, N3540, N2212);
and AND3 (N3549, N3547, N522, N2872);
nor NOR2 (N3550, N3532, N957);
xor XOR2 (N3551, N3484, N908);
not NOT1 (N3552, N3549);
buf BUF1 (N3553, N3552);
or OR4 (N3554, N3550, N1715, N1976, N1560);
or OR4 (N3555, N3551, N2209, N3058, N1699);
or OR2 (N3556, N3545, N2047);
nand NAND3 (N3557, N3554, N911, N2357);
not NOT1 (N3558, N3555);
nand NAND2 (N3559, N3553, N1052);
xor XOR2 (N3560, N3538, N3332);
nand NAND4 (N3561, N3557, N743, N102, N1804);
buf BUF1 (N3562, N3561);
not NOT1 (N3563, N3559);
nor NOR2 (N3564, N3546, N275);
and AND2 (N3565, N3544, N1337);
xor XOR2 (N3566, N3548, N2281);
nor NOR4 (N3567, N3509, N1140, N256, N980);
nor NOR2 (N3568, N3565, N1443);
nor NOR3 (N3569, N3563, N1708, N3196);
or OR2 (N3570, N3556, N1687);
or OR4 (N3571, N3543, N2999, N1119, N1344);
or OR3 (N3572, N3570, N349, N643);
nor NOR3 (N3573, N3564, N2717, N2220);
buf BUF1 (N3574, N3560);
xor XOR2 (N3575, N3573, N814);
not NOT1 (N3576, N3572);
not NOT1 (N3577, N3568);
not NOT1 (N3578, N3558);
not NOT1 (N3579, N3567);
or OR3 (N3580, N3578, N1424, N3129);
not NOT1 (N3581, N3579);
not NOT1 (N3582, N3575);
nand NAND3 (N3583, N3569, N2843, N2864);
and AND4 (N3584, N3583, N176, N545, N118);
nor NOR4 (N3585, N3581, N2475, N811, N91);
buf BUF1 (N3586, N3584);
and AND4 (N3587, N3580, N2848, N320, N1858);
nor NOR4 (N3588, N3566, N2069, N3398, N2231);
xor XOR2 (N3589, N3585, N1937);
nor NOR4 (N3590, N3588, N2008, N1604, N578);
nor NOR4 (N3591, N3577, N2058, N2495, N391);
nand NAND4 (N3592, N3571, N187, N2779, N3063);
nor NOR3 (N3593, N3590, N2077, N3181);
nor NOR4 (N3594, N3592, N1322, N726, N3041);
or OR2 (N3595, N3591, N1858);
buf BUF1 (N3596, N3582);
and AND4 (N3597, N3596, N1471, N169, N1809);
xor XOR2 (N3598, N3595, N2386);
nand NAND4 (N3599, N3589, N1991, N1578, N490);
nand NAND3 (N3600, N3574, N1464, N2403);
and AND2 (N3601, N3586, N1585);
nand NAND4 (N3602, N3599, N1075, N2069, N564);
nor NOR3 (N3603, N3576, N1771, N2486);
nand NAND4 (N3604, N3600, N1114, N1224, N179);
nand NAND2 (N3605, N3604, N1024);
buf BUF1 (N3606, N3603);
not NOT1 (N3607, N3597);
nand NAND3 (N3608, N3587, N708, N610);
or OR4 (N3609, N3605, N2588, N525, N1414);
nor NOR3 (N3610, N3609, N3191, N2731);
and AND3 (N3611, N3601, N347, N3088);
and AND4 (N3612, N3610, N1766, N1487, N2792);
nor NOR2 (N3613, N3611, N796);
xor XOR2 (N3614, N3608, N3104);
xor XOR2 (N3615, N3562, N433);
xor XOR2 (N3616, N3615, N2849);
not NOT1 (N3617, N3602);
and AND4 (N3618, N3606, N299, N1201, N2561);
or OR2 (N3619, N3618, N3573);
nor NOR4 (N3620, N3594, N1695, N2477, N1569);
buf BUF1 (N3621, N3612);
nor NOR4 (N3622, N3617, N3073, N2993, N1391);
or OR3 (N3623, N3614, N2017, N2905);
and AND2 (N3624, N3622, N953);
and AND4 (N3625, N3621, N833, N2904, N409);
or OR4 (N3626, N3620, N1913, N1256, N343);
nand NAND2 (N3627, N3613, N2537);
and AND3 (N3628, N3624, N1563, N558);
nand NAND3 (N3629, N3626, N2216, N2965);
buf BUF1 (N3630, N3616);
or OR3 (N3631, N3619, N2659, N950);
nand NAND2 (N3632, N3631, N2245);
xor XOR2 (N3633, N3627, N1224);
buf BUF1 (N3634, N3629);
buf BUF1 (N3635, N3593);
buf BUF1 (N3636, N3623);
and AND3 (N3637, N3635, N1728, N872);
nor NOR4 (N3638, N3636, N2066, N2300, N858);
nand NAND2 (N3639, N3634, N3144);
nand NAND2 (N3640, N3632, N2254);
buf BUF1 (N3641, N3640);
nand NAND2 (N3642, N3625, N3013);
nand NAND3 (N3643, N3639, N1810, N535);
nand NAND2 (N3644, N3642, N116);
xor XOR2 (N3645, N3641, N3516);
xor XOR2 (N3646, N3633, N1658);
or OR3 (N3647, N3646, N2251, N937);
nand NAND3 (N3648, N3598, N1127, N927);
or OR4 (N3649, N3638, N1965, N251, N809);
not NOT1 (N3650, N3644);
nand NAND4 (N3651, N3643, N1281, N3117, N818);
buf BUF1 (N3652, N3648);
xor XOR2 (N3653, N3651, N520);
nor NOR2 (N3654, N3652, N1736);
buf BUF1 (N3655, N3637);
buf BUF1 (N3656, N3655);
xor XOR2 (N3657, N3628, N2418);
buf BUF1 (N3658, N3607);
xor XOR2 (N3659, N3658, N642);
not NOT1 (N3660, N3649);
xor XOR2 (N3661, N3660, N1388);
and AND3 (N3662, N3653, N1058, N3487);
buf BUF1 (N3663, N3661);
buf BUF1 (N3664, N3650);
nand NAND2 (N3665, N3645, N1460);
buf BUF1 (N3666, N3654);
xor XOR2 (N3667, N3657, N1690);
nand NAND2 (N3668, N3656, N2275);
or OR4 (N3669, N3667, N1430, N281, N1558);
not NOT1 (N3670, N3665);
nand NAND2 (N3671, N3647, N1646);
xor XOR2 (N3672, N3671, N1340);
and AND2 (N3673, N3669, N1277);
not NOT1 (N3674, N3659);
not NOT1 (N3675, N3630);
or OR3 (N3676, N3672, N636, N430);
and AND4 (N3677, N3664, N2493, N262, N369);
not NOT1 (N3678, N3675);
nor NOR2 (N3679, N3666, N1660);
and AND4 (N3680, N3670, N1189, N2960, N1404);
nor NOR4 (N3681, N3673, N1070, N921, N1048);
xor XOR2 (N3682, N3663, N1038);
xor XOR2 (N3683, N3678, N3399);
not NOT1 (N3684, N3677);
nor NOR2 (N3685, N3684, N3055);
and AND3 (N3686, N3683, N3553, N936);
xor XOR2 (N3687, N3662, N561);
or OR3 (N3688, N3676, N1724, N3583);
and AND2 (N3689, N3687, N3521);
nand NAND4 (N3690, N3681, N2406, N2905, N2889);
and AND4 (N3691, N3688, N666, N1772, N560);
not NOT1 (N3692, N3674);
or OR3 (N3693, N3690, N3131, N1779);
or OR3 (N3694, N3679, N2834, N220);
xor XOR2 (N3695, N3694, N2379);
buf BUF1 (N3696, N3668);
buf BUF1 (N3697, N3680);
and AND4 (N3698, N3693, N765, N2698, N3398);
xor XOR2 (N3699, N3695, N3229);
nand NAND3 (N3700, N3685, N3371, N2338);
and AND3 (N3701, N3692, N1545, N102);
or OR4 (N3702, N3700, N765, N1387, N102);
or OR4 (N3703, N3702, N1577, N1103, N3010);
or OR2 (N3704, N3696, N434);
or OR2 (N3705, N3682, N236);
buf BUF1 (N3706, N3691);
and AND2 (N3707, N3699, N1826);
and AND4 (N3708, N3701, N2828, N1590, N3084);
buf BUF1 (N3709, N3706);
or OR4 (N3710, N3698, N1739, N1102, N2543);
not NOT1 (N3711, N3707);
buf BUF1 (N3712, N3711);
or OR2 (N3713, N3709, N1228);
not NOT1 (N3714, N3689);
xor XOR2 (N3715, N3703, N3572);
buf BUF1 (N3716, N3708);
nor NOR3 (N3717, N3704, N1205, N2208);
buf BUF1 (N3718, N3710);
nand NAND2 (N3719, N3716, N3049);
nor NOR3 (N3720, N3713, N1187, N2845);
nand NAND2 (N3721, N3715, N818);
xor XOR2 (N3722, N3721, N1276);
buf BUF1 (N3723, N3718);
or OR4 (N3724, N3712, N333, N22, N2710);
xor XOR2 (N3725, N3723, N3155);
and AND2 (N3726, N3722, N1769);
xor XOR2 (N3727, N3724, N1330);
and AND3 (N3728, N3725, N2103, N297);
or OR4 (N3729, N3705, N1810, N3172, N2175);
not NOT1 (N3730, N3697);
xor XOR2 (N3731, N3720, N1234);
buf BUF1 (N3732, N3730);
not NOT1 (N3733, N3686);
buf BUF1 (N3734, N3732);
buf BUF1 (N3735, N3733);
not NOT1 (N3736, N3714);
nor NOR4 (N3737, N3717, N343, N95, N3223);
xor XOR2 (N3738, N3734, N176);
and AND3 (N3739, N3729, N1774, N883);
or OR3 (N3740, N3731, N1657, N1526);
nand NAND3 (N3741, N3719, N3540, N3199);
buf BUF1 (N3742, N3741);
xor XOR2 (N3743, N3727, N1456);
xor XOR2 (N3744, N3726, N2056);
or OR2 (N3745, N3743, N2489);
buf BUF1 (N3746, N3738);
nand NAND4 (N3747, N3742, N839, N698, N636);
not NOT1 (N3748, N3747);
nor NOR4 (N3749, N3737, N1001, N1723, N961);
xor XOR2 (N3750, N3745, N2889);
and AND4 (N3751, N3739, N2914, N2415, N954);
and AND4 (N3752, N3746, N2838, N2436, N95);
buf BUF1 (N3753, N3740);
not NOT1 (N3754, N3744);
and AND4 (N3755, N3752, N1862, N865, N2172);
or OR2 (N3756, N3748, N2917);
not NOT1 (N3757, N3753);
or OR3 (N3758, N3735, N3231, N65);
nor NOR2 (N3759, N3751, N2792);
xor XOR2 (N3760, N3755, N3016);
nor NOR2 (N3761, N3749, N1578);
or OR4 (N3762, N3728, N1947, N2901, N1214);
buf BUF1 (N3763, N3759);
nand NAND3 (N3764, N3757, N163, N2535);
buf BUF1 (N3765, N3761);
not NOT1 (N3766, N3754);
and AND2 (N3767, N3764, N2487);
nor NOR3 (N3768, N3756, N3416, N727);
or OR4 (N3769, N3768, N3670, N2363, N1787);
and AND4 (N3770, N3767, N2091, N317, N1850);
or OR4 (N3771, N3766, N2648, N1620, N3144);
nor NOR2 (N3772, N3758, N2329);
and AND4 (N3773, N3769, N1653, N2179, N432);
not NOT1 (N3774, N3762);
xor XOR2 (N3775, N3772, N1519);
and AND4 (N3776, N3770, N1610, N1481, N1458);
not NOT1 (N3777, N3775);
not NOT1 (N3778, N3765);
and AND4 (N3779, N3773, N2185, N455, N1225);
xor XOR2 (N3780, N3777, N417);
nor NOR3 (N3781, N3760, N328, N907);
and AND4 (N3782, N3774, N139, N2182, N3175);
not NOT1 (N3783, N3781);
and AND4 (N3784, N3750, N1193, N2011, N3089);
nor NOR4 (N3785, N3778, N1814, N3463, N2194);
buf BUF1 (N3786, N3771);
or OR4 (N3787, N3736, N1964, N2171, N3105);
and AND3 (N3788, N3787, N358, N1754);
or OR4 (N3789, N3779, N2552, N3601, N501);
and AND4 (N3790, N3784, N3423, N2402, N2310);
nor NOR3 (N3791, N3790, N3303, N202);
nor NOR2 (N3792, N3776, N3716);
nor NOR3 (N3793, N3788, N291, N2660);
buf BUF1 (N3794, N3786);
buf BUF1 (N3795, N3783);
not NOT1 (N3796, N3792);
not NOT1 (N3797, N3796);
nor NOR3 (N3798, N3780, N2544, N1357);
not NOT1 (N3799, N3791);
nand NAND3 (N3800, N3793, N2519, N2154);
nor NOR2 (N3801, N3763, N1138);
or OR2 (N3802, N3789, N1500);
not NOT1 (N3803, N3800);
not NOT1 (N3804, N3799);
nor NOR2 (N3805, N3798, N2570);
buf BUF1 (N3806, N3797);
nor NOR4 (N3807, N3803, N1835, N2699, N3291);
nor NOR2 (N3808, N3801, N3775);
and AND3 (N3809, N3808, N423, N838);
xor XOR2 (N3810, N3809, N2815);
nor NOR4 (N3811, N3782, N2927, N56, N2277);
xor XOR2 (N3812, N3806, N390);
xor XOR2 (N3813, N3785, N2676);
or OR3 (N3814, N3813, N1752, N3032);
xor XOR2 (N3815, N3810, N3241);
or OR2 (N3816, N3794, N3792);
xor XOR2 (N3817, N3814, N2367);
not NOT1 (N3818, N3815);
xor XOR2 (N3819, N3807, N2308);
not NOT1 (N3820, N3818);
nor NOR4 (N3821, N3819, N3144, N145, N1130);
xor XOR2 (N3822, N3817, N347);
not NOT1 (N3823, N3812);
not NOT1 (N3824, N3820);
or OR2 (N3825, N3816, N3224);
and AND3 (N3826, N3804, N1623, N800);
or OR4 (N3827, N3823, N1686, N3017, N1701);
or OR3 (N3828, N3821, N2389, N48);
or OR2 (N3829, N3828, N1131);
xor XOR2 (N3830, N3795, N86);
or OR2 (N3831, N3824, N523);
buf BUF1 (N3832, N3829);
and AND2 (N3833, N3827, N1874);
and AND3 (N3834, N3833, N3159, N675);
buf BUF1 (N3835, N3811);
or OR4 (N3836, N3805, N536, N285, N496);
buf BUF1 (N3837, N3822);
nor NOR2 (N3838, N3835, N2167);
buf BUF1 (N3839, N3834);
or OR2 (N3840, N3825, N2305);
and AND2 (N3841, N3839, N2511);
and AND3 (N3842, N3836, N5, N2334);
or OR4 (N3843, N3830, N2552, N3591, N1602);
nand NAND3 (N3844, N3837, N2827, N2631);
nor NOR3 (N3845, N3842, N688, N2983);
xor XOR2 (N3846, N3832, N1415);
and AND2 (N3847, N3843, N2225);
buf BUF1 (N3848, N3841);
buf BUF1 (N3849, N3848);
not NOT1 (N3850, N3840);
and AND4 (N3851, N3850, N374, N994, N351);
and AND2 (N3852, N3846, N1496);
or OR2 (N3853, N3845, N1076);
nand NAND4 (N3854, N3838, N1318, N1249, N651);
or OR3 (N3855, N3849, N2456, N1815);
buf BUF1 (N3856, N3847);
not NOT1 (N3857, N3831);
buf BUF1 (N3858, N3844);
buf BUF1 (N3859, N3856);
and AND2 (N3860, N3857, N1322);
nor NOR4 (N3861, N3852, N873, N2189, N1342);
and AND2 (N3862, N3860, N714);
nand NAND2 (N3863, N3851, N3276);
not NOT1 (N3864, N3854);
not NOT1 (N3865, N3859);
xor XOR2 (N3866, N3861, N1881);
nor NOR4 (N3867, N3858, N2012, N1899, N3772);
and AND2 (N3868, N3864, N3061);
and AND4 (N3869, N3853, N2846, N589, N3682);
or OR4 (N3870, N3865, N646, N678, N3519);
nand NAND3 (N3871, N3869, N1613, N2726);
nor NOR2 (N3872, N3870, N2823);
and AND2 (N3873, N3872, N963);
xor XOR2 (N3874, N3873, N800);
buf BUF1 (N3875, N3862);
not NOT1 (N3876, N3868);
and AND2 (N3877, N3876, N1635);
or OR3 (N3878, N3863, N802, N2834);
not NOT1 (N3879, N3826);
nor NOR2 (N3880, N3875, N2129);
or OR3 (N3881, N3866, N471, N76);
not NOT1 (N3882, N3867);
nor NOR2 (N3883, N3802, N1910);
not NOT1 (N3884, N3883);
xor XOR2 (N3885, N3880, N828);
not NOT1 (N3886, N3855);
and AND3 (N3887, N3877, N3116, N2901);
nor NOR2 (N3888, N3879, N2768);
and AND2 (N3889, N3886, N1708);
buf BUF1 (N3890, N3874);
and AND2 (N3891, N3885, N2298);
nor NOR2 (N3892, N3882, N3169);
and AND3 (N3893, N3891, N100, N3327);
or OR2 (N3894, N3881, N230);
xor XOR2 (N3895, N3888, N3035);
xor XOR2 (N3896, N3884, N580);
nor NOR4 (N3897, N3878, N3539, N1583, N840);
buf BUF1 (N3898, N3890);
nor NOR3 (N3899, N3898, N175, N1996);
nor NOR4 (N3900, N3899, N1731, N1463, N887);
nor NOR3 (N3901, N3887, N1019, N371);
nor NOR2 (N3902, N3871, N1224);
xor XOR2 (N3903, N3896, N857);
not NOT1 (N3904, N3901);
not NOT1 (N3905, N3897);
nand NAND4 (N3906, N3902, N585, N594, N2530);
xor XOR2 (N3907, N3894, N244);
not NOT1 (N3908, N3900);
not NOT1 (N3909, N3892);
nand NAND3 (N3910, N3909, N1086, N948);
nor NOR2 (N3911, N3905, N2021);
not NOT1 (N3912, N3903);
or OR3 (N3913, N3911, N3289, N998);
buf BUF1 (N3914, N3904);
nor NOR2 (N3915, N3906, N3059);
and AND3 (N3916, N3907, N909, N1283);
buf BUF1 (N3917, N3895);
nand NAND2 (N3918, N3908, N1896);
nand NAND2 (N3919, N3889, N1396);
nand NAND3 (N3920, N3917, N357, N520);
or OR4 (N3921, N3913, N2175, N2444, N171);
nand NAND2 (N3922, N3916, N3805);
nor NOR3 (N3923, N3918, N3239, N1525);
not NOT1 (N3924, N3919);
nor NOR4 (N3925, N3914, N1458, N3268, N364);
and AND4 (N3926, N3920, N1330, N3248, N3002);
buf BUF1 (N3927, N3924);
nand NAND2 (N3928, N3915, N2240);
xor XOR2 (N3929, N3927, N474);
or OR4 (N3930, N3926, N3639, N2990, N3135);
and AND4 (N3931, N3922, N1848, N2445, N560);
buf BUF1 (N3932, N3910);
or OR3 (N3933, N3930, N1030, N2227);
and AND3 (N3934, N3925, N2757, N1072);
xor XOR2 (N3935, N3921, N848);
nand NAND3 (N3936, N3934, N1993, N3485);
xor XOR2 (N3937, N3932, N3919);
not NOT1 (N3938, N3893);
xor XOR2 (N3939, N3928, N3174);
xor XOR2 (N3940, N3933, N3395);
and AND3 (N3941, N3937, N2474, N3462);
xor XOR2 (N3942, N3929, N780);
and AND2 (N3943, N3938, N3002);
buf BUF1 (N3944, N3923);
nand NAND2 (N3945, N3936, N441);
not NOT1 (N3946, N3944);
and AND2 (N3947, N3931, N485);
or OR3 (N3948, N3912, N1085, N3247);
nand NAND3 (N3949, N3947, N3432, N1372);
nand NAND4 (N3950, N3940, N2261, N3617, N725);
not NOT1 (N3951, N3946);
and AND2 (N3952, N3948, N1651);
and AND3 (N3953, N3951, N1157, N3077);
nand NAND3 (N3954, N3935, N3139, N3581);
and AND2 (N3955, N3939, N289);
or OR3 (N3956, N3942, N2428, N2573);
nand NAND4 (N3957, N3943, N3623, N849, N2098);
or OR4 (N3958, N3956, N1425, N2090, N1262);
and AND2 (N3959, N3950, N3830);
buf BUF1 (N3960, N3958);
not NOT1 (N3961, N3949);
nor NOR2 (N3962, N3941, N401);
buf BUF1 (N3963, N3945);
xor XOR2 (N3964, N3961, N3642);
and AND4 (N3965, N3963, N3375, N481, N547);
xor XOR2 (N3966, N3955, N3275);
nand NAND4 (N3967, N3954, N733, N3665, N45);
buf BUF1 (N3968, N3960);
buf BUF1 (N3969, N3962);
or OR3 (N3970, N3965, N3191, N3429);
buf BUF1 (N3971, N3953);
nand NAND3 (N3972, N3959, N2907, N844);
and AND3 (N3973, N3971, N3463, N1263);
buf BUF1 (N3974, N3972);
nand NAND3 (N3975, N3974, N3619, N355);
nor NOR2 (N3976, N3973, N967);
nor NOR4 (N3977, N3968, N2758, N352, N1296);
nor NOR2 (N3978, N3976, N2735);
and AND2 (N3979, N3964, N2343);
and AND4 (N3980, N3978, N64, N723, N1902);
and AND4 (N3981, N3966, N2081, N1964, N2271);
xor XOR2 (N3982, N3970, N1380);
xor XOR2 (N3983, N3967, N3232);
nor NOR3 (N3984, N3981, N2477, N1730);
nand NAND4 (N3985, N3969, N3632, N3439, N3821);
buf BUF1 (N3986, N3980);
and AND4 (N3987, N3957, N2873, N570, N1152);
nand NAND2 (N3988, N3985, N2154);
buf BUF1 (N3989, N3979);
nand NAND4 (N3990, N3988, N1661, N173, N198);
xor XOR2 (N3991, N3984, N564);
or OR4 (N3992, N3990, N2569, N3778, N1487);
nand NAND2 (N3993, N3991, N1934);
and AND2 (N3994, N3982, N3023);
not NOT1 (N3995, N3952);
not NOT1 (N3996, N3992);
buf BUF1 (N3997, N3996);
xor XOR2 (N3998, N3994, N747);
nor NOR4 (N3999, N3995, N3613, N1501, N1135);
xor XOR2 (N4000, N3983, N2386);
xor XOR2 (N4001, N3999, N3265);
xor XOR2 (N4002, N3977, N3593);
xor XOR2 (N4003, N3986, N901);
buf BUF1 (N4004, N3997);
or OR3 (N4005, N4004, N447, N723);
or OR4 (N4006, N3993, N2846, N3522, N2833);
or OR3 (N4007, N4003, N1277, N2765);
nand NAND3 (N4008, N3989, N1151, N1756);
and AND3 (N4009, N4001, N2775, N3462);
nand NAND3 (N4010, N4002, N961, N2754);
and AND3 (N4011, N3998, N1083, N1844);
xor XOR2 (N4012, N3987, N286);
nor NOR3 (N4013, N4008, N2325, N3692);
or OR2 (N4014, N4006, N4000);
xor XOR2 (N4015, N2712, N832);
nor NOR2 (N4016, N4014, N230);
or OR3 (N4017, N4016, N1997, N3488);
and AND2 (N4018, N4010, N1219);
or OR2 (N4019, N4009, N1865);
and AND3 (N4020, N3975, N110, N533);
or OR4 (N4021, N4018, N962, N1608, N21);
or OR4 (N4022, N4017, N3632, N3923, N1912);
nand NAND3 (N4023, N4021, N3640, N3286);
and AND2 (N4024, N4013, N1816);
xor XOR2 (N4025, N4007, N2498);
nand NAND4 (N4026, N4022, N1562, N1592, N208);
or OR2 (N4027, N4025, N1528);
nand NAND4 (N4028, N4012, N2587, N1390, N1967);
buf BUF1 (N4029, N4024);
or OR2 (N4030, N4029, N1675);
nand NAND2 (N4031, N4015, N1409);
not NOT1 (N4032, N4011);
buf BUF1 (N4033, N4026);
and AND4 (N4034, N4019, N3778, N2313, N3116);
nand NAND4 (N4035, N4028, N175, N2078, N779);
and AND4 (N4036, N4023, N1295, N2731, N2283);
nand NAND2 (N4037, N4032, N1039);
xor XOR2 (N4038, N4030, N3513);
xor XOR2 (N4039, N4038, N2877);
nand NAND3 (N4040, N4027, N1342, N2091);
nand NAND3 (N4041, N4035, N1340, N1931);
buf BUF1 (N4042, N4031);
nand NAND3 (N4043, N4033, N2117, N514);
buf BUF1 (N4044, N4039);
nor NOR3 (N4045, N4044, N3221, N2885);
xor XOR2 (N4046, N4005, N3806);
xor XOR2 (N4047, N4034, N3019);
not NOT1 (N4048, N4042);
and AND3 (N4049, N4046, N1053, N1564);
and AND3 (N4050, N4045, N1540, N131);
or OR3 (N4051, N4036, N2332, N559);
xor XOR2 (N4052, N4020, N3728);
and AND4 (N4053, N4049, N1926, N2625, N2753);
xor XOR2 (N4054, N4041, N3541);
nand NAND3 (N4055, N4052, N2806, N3127);
or OR3 (N4056, N4040, N3629, N3934);
buf BUF1 (N4057, N4051);
nand NAND3 (N4058, N4043, N2781, N3301);
buf BUF1 (N4059, N4055);
nand NAND2 (N4060, N4054, N621);
xor XOR2 (N4061, N4047, N764);
xor XOR2 (N4062, N4060, N1312);
and AND4 (N4063, N4037, N1192, N768, N560);
xor XOR2 (N4064, N4048, N1377);
xor XOR2 (N4065, N4063, N2329);
or OR3 (N4066, N4061, N2362, N2660);
and AND3 (N4067, N4066, N356, N230);
and AND4 (N4068, N4064, N4017, N892, N3045);
xor XOR2 (N4069, N4058, N560);
not NOT1 (N4070, N4068);
and AND2 (N4071, N4050, N917);
buf BUF1 (N4072, N4067);
or OR3 (N4073, N4071, N814, N3550);
buf BUF1 (N4074, N4059);
nand NAND2 (N4075, N4065, N1857);
nand NAND4 (N4076, N4072, N958, N2003, N556);
and AND2 (N4077, N4062, N838);
buf BUF1 (N4078, N4056);
buf BUF1 (N4079, N4077);
not NOT1 (N4080, N4057);
buf BUF1 (N4081, N4079);
and AND3 (N4082, N4080, N892, N1274);
or OR4 (N4083, N4076, N3772, N1103, N1602);
nor NOR2 (N4084, N4083, N2257);
and AND2 (N4085, N4081, N3617);
xor XOR2 (N4086, N4084, N1254);
nand NAND3 (N4087, N4069, N2219, N1889);
xor XOR2 (N4088, N4075, N505);
not NOT1 (N4089, N4086);
or OR2 (N4090, N4074, N938);
and AND3 (N4091, N4070, N1097, N1897);
nor NOR4 (N4092, N4053, N1330, N493, N1591);
not NOT1 (N4093, N4090);
buf BUF1 (N4094, N4088);
xor XOR2 (N4095, N4091, N3676);
nor NOR4 (N4096, N4095, N3490, N3042, N1237);
and AND3 (N4097, N4092, N3114, N1597);
nor NOR3 (N4098, N4087, N908, N3681);
or OR4 (N4099, N4085, N374, N3142, N3339);
or OR4 (N4100, N4093, N3324, N1376, N1639);
and AND2 (N4101, N4094, N141);
or OR4 (N4102, N4100, N3159, N963, N2368);
or OR2 (N4103, N4102, N1203);
nor NOR3 (N4104, N4098, N2483, N1686);
and AND4 (N4105, N4097, N1232, N3176, N2424);
xor XOR2 (N4106, N4105, N2344);
and AND4 (N4107, N4103, N1804, N1322, N1641);
and AND3 (N4108, N4096, N266, N2533);
or OR4 (N4109, N4106, N3516, N1406, N3423);
nand NAND3 (N4110, N4107, N1427, N2192);
nor NOR4 (N4111, N4104, N2795, N639, N3738);
and AND3 (N4112, N4111, N1273, N939);
or OR3 (N4113, N4110, N1560, N2494);
buf BUF1 (N4114, N4101);
not NOT1 (N4115, N4114);
nor NOR3 (N4116, N4115, N3540, N664);
xor XOR2 (N4117, N4073, N1014);
nand NAND4 (N4118, N4113, N4026, N2805, N461);
xor XOR2 (N4119, N4117, N818);
nand NAND4 (N4120, N4089, N3098, N526, N3235);
buf BUF1 (N4121, N4078);
xor XOR2 (N4122, N4121, N1161);
or OR3 (N4123, N4116, N3519, N91);
not NOT1 (N4124, N4099);
not NOT1 (N4125, N4124);
xor XOR2 (N4126, N4108, N2802);
or OR2 (N4127, N4109, N3056);
and AND2 (N4128, N4118, N2954);
and AND4 (N4129, N4127, N2160, N108, N2675);
nor NOR2 (N4130, N4126, N2904);
xor XOR2 (N4131, N4112, N873);
nor NOR3 (N4132, N4125, N1520, N1075);
xor XOR2 (N4133, N4132, N378);
not NOT1 (N4134, N4128);
and AND3 (N4135, N4082, N2958, N795);
not NOT1 (N4136, N4120);
and AND2 (N4137, N4133, N1659);
xor XOR2 (N4138, N4122, N719);
and AND3 (N4139, N4136, N2171, N786);
nor NOR4 (N4140, N4130, N2200, N2237, N1005);
xor XOR2 (N4141, N4140, N1837);
xor XOR2 (N4142, N4134, N3160);
nand NAND3 (N4143, N4129, N685, N325);
and AND2 (N4144, N4141, N1549);
buf BUF1 (N4145, N4131);
nor NOR2 (N4146, N4143, N3973);
or OR4 (N4147, N4123, N788, N877, N2484);
or OR3 (N4148, N4135, N95, N4078);
nor NOR4 (N4149, N4142, N720, N1381, N1327);
buf BUF1 (N4150, N4147);
nand NAND2 (N4151, N4137, N1945);
xor XOR2 (N4152, N4149, N4149);
not NOT1 (N4153, N4151);
nor NOR4 (N4154, N4145, N1540, N389, N2181);
nand NAND2 (N4155, N4139, N2550);
buf BUF1 (N4156, N4152);
buf BUF1 (N4157, N4119);
or OR4 (N4158, N4146, N3468, N1352, N541);
nand NAND4 (N4159, N4148, N3926, N3301, N2112);
buf BUF1 (N4160, N4150);
nand NAND4 (N4161, N4138, N249, N1826, N182);
buf BUF1 (N4162, N4144);
not NOT1 (N4163, N4156);
nand NAND2 (N4164, N4157, N1929);
and AND2 (N4165, N4154, N3322);
nor NOR3 (N4166, N4159, N979, N3426);
and AND3 (N4167, N4166, N1681, N1371);
or OR3 (N4168, N4165, N2669, N1603);
and AND4 (N4169, N4162, N3613, N1516, N3724);
or OR2 (N4170, N4161, N1095);
and AND2 (N4171, N4164, N3449);
not NOT1 (N4172, N4158);
nor NOR3 (N4173, N4167, N2390, N176);
buf BUF1 (N4174, N4170);
and AND3 (N4175, N4172, N3520, N3748);
nand NAND2 (N4176, N4171, N403);
nand NAND3 (N4177, N4153, N1594, N2839);
xor XOR2 (N4178, N4168, N3842);
nand NAND3 (N4179, N4175, N2658, N1895);
and AND4 (N4180, N4176, N78, N1093, N2933);
not NOT1 (N4181, N4155);
or OR3 (N4182, N4160, N2494, N3996);
or OR3 (N4183, N4169, N766, N346);
and AND3 (N4184, N4174, N315, N2781);
nor NOR4 (N4185, N4173, N2116, N2363, N2230);
and AND4 (N4186, N4178, N1603, N4042, N2830);
or OR3 (N4187, N4181, N871, N2310);
or OR3 (N4188, N4177, N1240, N3363);
nor NOR3 (N4189, N4163, N2357, N407);
buf BUF1 (N4190, N4184);
or OR4 (N4191, N4180, N3847, N1991, N23);
or OR3 (N4192, N4186, N3443, N1800);
and AND4 (N4193, N4179, N1250, N757, N2749);
nand NAND2 (N4194, N4191, N3959);
not NOT1 (N4195, N4185);
or OR2 (N4196, N4189, N2539);
xor XOR2 (N4197, N4195, N1043);
and AND4 (N4198, N4194, N2189, N2762, N1636);
nor NOR3 (N4199, N4182, N1761, N1371);
nor NOR3 (N4200, N4183, N691, N2503);
nor NOR4 (N4201, N4190, N3083, N681, N1810);
or OR3 (N4202, N4200, N3416, N3169);
not NOT1 (N4203, N4199);
buf BUF1 (N4204, N4197);
buf BUF1 (N4205, N4198);
buf BUF1 (N4206, N4204);
not NOT1 (N4207, N4203);
xor XOR2 (N4208, N4188, N1862);
or OR2 (N4209, N4207, N3457);
xor XOR2 (N4210, N4206, N451);
and AND3 (N4211, N4210, N2276, N1851);
buf BUF1 (N4212, N4193);
or OR3 (N4213, N4196, N3821, N2681);
nand NAND3 (N4214, N4202, N107, N401);
buf BUF1 (N4215, N4208);
nand NAND3 (N4216, N4212, N476, N3783);
not NOT1 (N4217, N4187);
and AND3 (N4218, N4216, N140, N2133);
xor XOR2 (N4219, N4209, N968);
not NOT1 (N4220, N4211);
not NOT1 (N4221, N4217);
nor NOR3 (N4222, N4192, N2099, N4218);
nor NOR3 (N4223, N2315, N3320, N1389);
and AND3 (N4224, N4215, N3448, N3955);
xor XOR2 (N4225, N4222, N1449);
and AND4 (N4226, N4220, N2611, N1386, N2093);
or OR2 (N4227, N4224, N1606);
buf BUF1 (N4228, N4201);
or OR4 (N4229, N4225, N2643, N2421, N2766);
buf BUF1 (N4230, N4226);
buf BUF1 (N4231, N4219);
nor NOR3 (N4232, N4214, N3337, N699);
buf BUF1 (N4233, N4231);
nor NOR3 (N4234, N4233, N4219, N3937);
not NOT1 (N4235, N4223);
xor XOR2 (N4236, N4227, N740);
and AND3 (N4237, N4205, N2271, N217);
buf BUF1 (N4238, N4235);
xor XOR2 (N4239, N4236, N718);
nor NOR2 (N4240, N4213, N3394);
buf BUF1 (N4241, N4228);
nand NAND3 (N4242, N4234, N3977, N1465);
xor XOR2 (N4243, N4221, N861);
nor NOR2 (N4244, N4242, N1372);
buf BUF1 (N4245, N4238);
buf BUF1 (N4246, N4239);
buf BUF1 (N4247, N4240);
not NOT1 (N4248, N4246);
buf BUF1 (N4249, N4241);
xor XOR2 (N4250, N4232, N2917);
buf BUF1 (N4251, N4229);
and AND3 (N4252, N4247, N556, N563);
and AND3 (N4253, N4249, N4060, N2327);
nand NAND3 (N4254, N4230, N3887, N1038);
not NOT1 (N4255, N4245);
nor NOR2 (N4256, N4251, N3930);
or OR4 (N4257, N4254, N3444, N2342, N831);
nor NOR4 (N4258, N4253, N1185, N88, N1091);
nand NAND4 (N4259, N4243, N1253, N2127, N4113);
buf BUF1 (N4260, N4259);
and AND3 (N4261, N4256, N2904, N103);
xor XOR2 (N4262, N4261, N3002);
or OR2 (N4263, N4250, N1002);
nor NOR4 (N4264, N4263, N3104, N345, N2825);
xor XOR2 (N4265, N4252, N1193);
and AND2 (N4266, N4255, N1618);
not NOT1 (N4267, N4262);
buf BUF1 (N4268, N4248);
xor XOR2 (N4269, N4260, N2530);
xor XOR2 (N4270, N4244, N399);
xor XOR2 (N4271, N4264, N2436);
nand NAND2 (N4272, N4237, N2987);
or OR4 (N4273, N4269, N2990, N1619, N2224);
or OR3 (N4274, N4267, N1157, N3221);
nand NAND4 (N4275, N4273, N590, N1774, N2707);
nor NOR4 (N4276, N4274, N3261, N1913, N2026);
and AND3 (N4277, N4270, N2946, N181);
nor NOR3 (N4278, N4268, N1764, N3906);
xor XOR2 (N4279, N4272, N365);
nand NAND2 (N4280, N4276, N843);
nor NOR3 (N4281, N4266, N2698, N3077);
xor XOR2 (N4282, N4275, N824);
nand NAND2 (N4283, N4281, N741);
or OR4 (N4284, N4257, N516, N2119, N2910);
nor NOR2 (N4285, N4258, N3540);
or OR2 (N4286, N4285, N678);
and AND3 (N4287, N4283, N1388, N2091);
nand NAND3 (N4288, N4282, N2454, N3901);
or OR3 (N4289, N4287, N211, N1886);
not NOT1 (N4290, N4289);
nor NOR2 (N4291, N4280, N62);
or OR3 (N4292, N4286, N1021, N985);
not NOT1 (N4293, N4279);
xor XOR2 (N4294, N4277, N596);
and AND2 (N4295, N4288, N1536);
xor XOR2 (N4296, N4293, N1945);
or OR3 (N4297, N4296, N3926, N3454);
and AND4 (N4298, N4271, N2291, N3829, N1985);
nor NOR3 (N4299, N4298, N2004, N3286);
and AND3 (N4300, N4295, N3728, N2687);
xor XOR2 (N4301, N4291, N4127);
not NOT1 (N4302, N4300);
and AND2 (N4303, N4284, N1717);
buf BUF1 (N4304, N4297);
xor XOR2 (N4305, N4278, N2556);
nand NAND3 (N4306, N4305, N255, N867);
or OR3 (N4307, N4304, N183, N539);
and AND3 (N4308, N4299, N3884, N3538);
or OR4 (N4309, N4307, N2338, N1998, N2808);
not NOT1 (N4310, N4290);
buf BUF1 (N4311, N4265);
nand NAND3 (N4312, N4306, N1988, N4287);
not NOT1 (N4313, N4301);
nand NAND2 (N4314, N4302, N3132);
not NOT1 (N4315, N4308);
not NOT1 (N4316, N4313);
nor NOR2 (N4317, N4315, N3701);
buf BUF1 (N4318, N4303);
and AND2 (N4319, N4312, N1132);
xor XOR2 (N4320, N4319, N2406);
xor XOR2 (N4321, N4309, N1404);
or OR3 (N4322, N4321, N516, N3686);
buf BUF1 (N4323, N4311);
nand NAND2 (N4324, N4322, N3631);
not NOT1 (N4325, N4310);
not NOT1 (N4326, N4316);
not NOT1 (N4327, N4324);
nand NAND3 (N4328, N4325, N3654, N2100);
and AND2 (N4329, N4314, N3805);
and AND2 (N4330, N4329, N2347);
not NOT1 (N4331, N4294);
buf BUF1 (N4332, N4320);
xor XOR2 (N4333, N4332, N1117);
buf BUF1 (N4334, N4328);
nand NAND4 (N4335, N4330, N2982, N3762, N303);
buf BUF1 (N4336, N4318);
or OR4 (N4337, N4326, N2666, N1420, N1804);
nor NOR3 (N4338, N4331, N194, N2507);
xor XOR2 (N4339, N4338, N1910);
nor NOR2 (N4340, N4292, N164);
and AND4 (N4341, N4334, N354, N3809, N2327);
nor NOR2 (N4342, N4333, N651);
xor XOR2 (N4343, N4317, N208);
nor NOR2 (N4344, N4342, N1324);
nor NOR4 (N4345, N4323, N1992, N3583, N3028);
xor XOR2 (N4346, N4336, N836);
nand NAND3 (N4347, N4339, N2763, N1204);
nand NAND4 (N4348, N4341, N1361, N4112, N2301);
not NOT1 (N4349, N4345);
not NOT1 (N4350, N4348);
xor XOR2 (N4351, N4335, N1694);
xor XOR2 (N4352, N4337, N1140);
not NOT1 (N4353, N4350);
xor XOR2 (N4354, N4349, N729);
nor NOR3 (N4355, N4351, N414, N1601);
not NOT1 (N4356, N4355);
nand NAND2 (N4357, N4347, N3594);
or OR2 (N4358, N4352, N1049);
buf BUF1 (N4359, N4343);
nor NOR3 (N4360, N4358, N1912, N1534);
buf BUF1 (N4361, N4353);
or OR4 (N4362, N4344, N2436, N3109, N2234);
and AND2 (N4363, N4360, N3753);
or OR2 (N4364, N4354, N335);
or OR4 (N4365, N4327, N200, N4161, N3040);
nand NAND4 (N4366, N4361, N2821, N1207, N3786);
or OR2 (N4367, N4357, N2760);
and AND3 (N4368, N4365, N3668, N2172);
not NOT1 (N4369, N4366);
nor NOR2 (N4370, N4340, N4216);
nor NOR2 (N4371, N4368, N1786);
or OR2 (N4372, N4359, N3975);
and AND4 (N4373, N4362, N3617, N1691, N503);
nor NOR3 (N4374, N4363, N3740, N2075);
xor XOR2 (N4375, N4374, N1103);
not NOT1 (N4376, N4375);
not NOT1 (N4377, N4372);
nand NAND3 (N4378, N4373, N3457, N805);
buf BUF1 (N4379, N4356);
buf BUF1 (N4380, N4371);
nor NOR2 (N4381, N4367, N2390);
xor XOR2 (N4382, N4377, N1041);
and AND3 (N4383, N4364, N2416, N1178);
not NOT1 (N4384, N4378);
and AND4 (N4385, N4384, N1714, N987, N436);
nor NOR2 (N4386, N4370, N1654);
buf BUF1 (N4387, N4386);
nor NOR2 (N4388, N4369, N4063);
not NOT1 (N4389, N4376);
nand NAND4 (N4390, N4380, N1411, N305, N805);
buf BUF1 (N4391, N4381);
xor XOR2 (N4392, N4346, N160);
nor NOR2 (N4393, N4385, N2174);
or OR4 (N4394, N4382, N2338, N2379, N1174);
or OR2 (N4395, N4390, N490);
xor XOR2 (N4396, N4388, N3062);
not NOT1 (N4397, N4392);
or OR3 (N4398, N4395, N2837, N4137);
xor XOR2 (N4399, N4393, N2300);
not NOT1 (N4400, N4394);
buf BUF1 (N4401, N4397);
not NOT1 (N4402, N4398);
and AND4 (N4403, N4379, N1556, N3208, N1419);
nor NOR4 (N4404, N4402, N1267, N3496, N1237);
buf BUF1 (N4405, N4403);
xor XOR2 (N4406, N4400, N2279);
and AND4 (N4407, N4391, N1178, N3956, N726);
buf BUF1 (N4408, N4407);
nand NAND4 (N4409, N4399, N1684, N2276, N2032);
nand NAND3 (N4410, N4404, N3686, N4049);
and AND2 (N4411, N4389, N3674);
nor NOR3 (N4412, N4401, N1457, N3733);
not NOT1 (N4413, N4408);
or OR4 (N4414, N4412, N3134, N2901, N2357);
not NOT1 (N4415, N4387);
and AND3 (N4416, N4410, N4187, N3033);
nand NAND2 (N4417, N4409, N44);
or OR2 (N4418, N4416, N2071);
nor NOR2 (N4419, N4413, N1799);
xor XOR2 (N4420, N4418, N4102);
nand NAND3 (N4421, N4383, N1132, N3509);
nor NOR2 (N4422, N4419, N2891);
or OR2 (N4423, N4422, N134);
or OR3 (N4424, N4405, N925, N472);
or OR3 (N4425, N4414, N2817, N418);
and AND3 (N4426, N4423, N1457, N523);
not NOT1 (N4427, N4417);
not NOT1 (N4428, N4426);
or OR3 (N4429, N4411, N798, N3768);
nand NAND4 (N4430, N4427, N3613, N1459, N446);
or OR4 (N4431, N4428, N1346, N1933, N3386);
nand NAND2 (N4432, N4431, N1388);
or OR2 (N4433, N4425, N3295);
xor XOR2 (N4434, N4415, N3081);
nand NAND3 (N4435, N4429, N1818, N2653);
xor XOR2 (N4436, N4406, N946);
or OR3 (N4437, N4424, N567, N3907);
and AND2 (N4438, N4435, N1366);
or OR2 (N4439, N4432, N4049);
nor NOR3 (N4440, N4396, N44, N4123);
or OR2 (N4441, N4434, N2224);
xor XOR2 (N4442, N4439, N3835);
and AND2 (N4443, N4440, N2482);
nor NOR4 (N4444, N4433, N1639, N117, N2609);
or OR2 (N4445, N4438, N2540);
xor XOR2 (N4446, N4420, N2540);
or OR4 (N4447, N4430, N2633, N1429, N1235);
xor XOR2 (N4448, N4446, N3299);
or OR2 (N4449, N4437, N812);
xor XOR2 (N4450, N4436, N3124);
nand NAND2 (N4451, N4445, N3521);
xor XOR2 (N4452, N4421, N1789);
not NOT1 (N4453, N4443);
and AND4 (N4454, N4447, N2662, N402, N2391);
and AND4 (N4455, N4451, N1886, N2366, N4135);
not NOT1 (N4456, N4453);
nand NAND2 (N4457, N4450, N3599);
xor XOR2 (N4458, N4448, N879);
xor XOR2 (N4459, N4441, N4448);
buf BUF1 (N4460, N4457);
or OR4 (N4461, N4459, N1432, N3336, N3058);
or OR4 (N4462, N4456, N1757, N2069, N1314);
nor NOR3 (N4463, N4442, N3055, N881);
buf BUF1 (N4464, N4461);
or OR2 (N4465, N4460, N3365);
nand NAND4 (N4466, N4444, N665, N4132, N727);
or OR4 (N4467, N4455, N1436, N4357, N3212);
buf BUF1 (N4468, N4449);
nand NAND4 (N4469, N4466, N2260, N1433, N3374);
and AND4 (N4470, N4458, N2995, N4024, N2028);
nand NAND4 (N4471, N4465, N2950, N3775, N381);
and AND2 (N4472, N4454, N282);
xor XOR2 (N4473, N4464, N1329);
xor XOR2 (N4474, N4470, N4141);
or OR4 (N4475, N4471, N2830, N3647, N2703);
not NOT1 (N4476, N4463);
not NOT1 (N4477, N4469);
buf BUF1 (N4478, N4452);
xor XOR2 (N4479, N4462, N2110);
xor XOR2 (N4480, N4474, N3519);
or OR2 (N4481, N4467, N2856);
or OR2 (N4482, N4480, N581);
buf BUF1 (N4483, N4478);
not NOT1 (N4484, N4475);
nand NAND2 (N4485, N4479, N1993);
xor XOR2 (N4486, N4484, N1261);
or OR3 (N4487, N4481, N1660, N1932);
nand NAND3 (N4488, N4473, N3321, N1687);
or OR2 (N4489, N4486, N1952);
or OR4 (N4490, N4472, N889, N1893, N2410);
nor NOR4 (N4491, N4482, N992, N2676, N2151);
nand NAND4 (N4492, N4490, N4385, N2543, N3659);
or OR4 (N4493, N4491, N3486, N2898, N995);
nor NOR2 (N4494, N4489, N4112);
nand NAND3 (N4495, N4485, N1473, N1205);
not NOT1 (N4496, N4483);
or OR4 (N4497, N4476, N2202, N1526, N914);
and AND2 (N4498, N4468, N1615);
not NOT1 (N4499, N4488);
nor NOR2 (N4500, N4497, N817);
buf BUF1 (N4501, N4500);
and AND3 (N4502, N4492, N4, N353);
or OR3 (N4503, N4493, N1324, N1712);
not NOT1 (N4504, N4501);
nor NOR4 (N4505, N4477, N2270, N3855, N2907);
nor NOR2 (N4506, N4505, N2690);
buf BUF1 (N4507, N4495);
and AND3 (N4508, N4502, N2513, N1961);
and AND3 (N4509, N4499, N3348, N3150);
buf BUF1 (N4510, N4506);
xor XOR2 (N4511, N4510, N848);
and AND2 (N4512, N4487, N2189);
and AND2 (N4513, N4512, N3549);
nand NAND3 (N4514, N4498, N1543, N3902);
and AND3 (N4515, N4509, N416, N647);
or OR2 (N4516, N4504, N4364);
nor NOR3 (N4517, N4508, N4301, N683);
and AND4 (N4518, N4507, N2424, N4111, N474);
xor XOR2 (N4519, N4503, N299);
and AND3 (N4520, N4516, N758, N2748);
nor NOR3 (N4521, N4514, N3001, N969);
nor NOR3 (N4522, N4496, N3778, N67);
nor NOR4 (N4523, N4519, N188, N664, N2431);
nand NAND3 (N4524, N4521, N2035, N2592);
buf BUF1 (N4525, N4513);
nor NOR3 (N4526, N4522, N33, N3330);
xor XOR2 (N4527, N4526, N3253);
or OR3 (N4528, N4527, N4501, N3100);
and AND2 (N4529, N4524, N426);
and AND4 (N4530, N4515, N1750, N2267, N2179);
buf BUF1 (N4531, N4517);
and AND3 (N4532, N4520, N3543, N100);
nand NAND3 (N4533, N4528, N1568, N4422);
nor NOR2 (N4534, N4511, N4533);
buf BUF1 (N4535, N430);
not NOT1 (N4536, N4535);
not NOT1 (N4537, N4536);
xor XOR2 (N4538, N4494, N2148);
not NOT1 (N4539, N4525);
nor NOR3 (N4540, N4537, N864, N1044);
nand NAND3 (N4541, N4540, N3046, N1549);
buf BUF1 (N4542, N4532);
buf BUF1 (N4543, N4539);
and AND3 (N4544, N4538, N4055, N4036);
and AND3 (N4545, N4544, N1715, N1888);
nand NAND2 (N4546, N4530, N2920);
not NOT1 (N4547, N4534);
or OR4 (N4548, N4546, N516, N4420, N2776);
nor NOR4 (N4549, N4523, N2420, N3500, N978);
or OR4 (N4550, N4548, N4402, N859, N2607);
buf BUF1 (N4551, N4550);
nor NOR4 (N4552, N4542, N4508, N1157, N4421);
or OR2 (N4553, N4543, N3128);
and AND2 (N4554, N4549, N2864);
and AND3 (N4555, N4554, N128, N2820);
and AND3 (N4556, N4551, N568, N2397);
nand NAND2 (N4557, N4545, N3421);
not NOT1 (N4558, N4555);
xor XOR2 (N4559, N4531, N1636);
nor NOR2 (N4560, N4552, N3684);
and AND4 (N4561, N4560, N2248, N1153, N2154);
or OR2 (N4562, N4558, N717);
not NOT1 (N4563, N4557);
and AND3 (N4564, N4562, N760, N417);
buf BUF1 (N4565, N4563);
and AND4 (N4566, N4565, N2052, N910, N2622);
nor NOR4 (N4567, N4547, N3385, N4094, N3537);
nand NAND4 (N4568, N4518, N987, N54, N572);
xor XOR2 (N4569, N4556, N3886);
not NOT1 (N4570, N4567);
not NOT1 (N4571, N4570);
not NOT1 (N4572, N4561);
buf BUF1 (N4573, N4571);
or OR2 (N4574, N4564, N2976);
xor XOR2 (N4575, N4541, N887);
and AND3 (N4576, N4574, N3878, N4161);
nor NOR4 (N4577, N4575, N2667, N3385, N19);
nand NAND4 (N4578, N4568, N1624, N543, N4108);
xor XOR2 (N4579, N4553, N4065);
nand NAND3 (N4580, N4566, N869, N3075);
and AND3 (N4581, N4578, N2878, N914);
nor NOR2 (N4582, N4581, N4234);
buf BUF1 (N4583, N4573);
not NOT1 (N4584, N4576);
and AND3 (N4585, N4572, N2154, N2299);
and AND3 (N4586, N4584, N3321, N1996);
xor XOR2 (N4587, N4569, N399);
not NOT1 (N4588, N4587);
nand NAND4 (N4589, N4580, N4248, N1677, N1437);
and AND4 (N4590, N4586, N1021, N4262, N1937);
or OR2 (N4591, N4529, N2805);
nand NAND4 (N4592, N4583, N1856, N2330, N258);
buf BUF1 (N4593, N4582);
and AND3 (N4594, N4577, N2126, N1026);
not NOT1 (N4595, N4591);
nor NOR4 (N4596, N4595, N2129, N1595, N1270);
and AND3 (N4597, N4589, N2460, N804);
nand NAND4 (N4598, N4596, N4484, N3067, N2795);
or OR4 (N4599, N4592, N4478, N2571, N4291);
and AND2 (N4600, N4594, N3923);
not NOT1 (N4601, N4593);
not NOT1 (N4602, N4599);
not NOT1 (N4603, N4588);
and AND4 (N4604, N4559, N548, N425, N1730);
or OR4 (N4605, N4603, N342, N2511, N796);
and AND4 (N4606, N4604, N4071, N1938, N1487);
and AND2 (N4607, N4579, N4196);
nand NAND2 (N4608, N4590, N2273);
xor XOR2 (N4609, N4585, N2270);
not NOT1 (N4610, N4605);
nor NOR4 (N4611, N4597, N2097, N899, N1174);
buf BUF1 (N4612, N4610);
or OR4 (N4613, N4601, N849, N324, N4465);
or OR2 (N4614, N4598, N4124);
buf BUF1 (N4615, N4614);
xor XOR2 (N4616, N4609, N811);
nor NOR4 (N4617, N4616, N1920, N1601, N1495);
not NOT1 (N4618, N4613);
not NOT1 (N4619, N4615);
or OR3 (N4620, N4602, N4489, N3208);
xor XOR2 (N4621, N4612, N769);
nand NAND2 (N4622, N4600, N3625);
buf BUF1 (N4623, N4618);
buf BUF1 (N4624, N4621);
nor NOR2 (N4625, N4620, N3732);
xor XOR2 (N4626, N4625, N3950);
nor NOR4 (N4627, N4623, N232, N2398, N1147);
or OR3 (N4628, N4617, N932, N4215);
buf BUF1 (N4629, N4611);
not NOT1 (N4630, N4619);
xor XOR2 (N4631, N4622, N2065);
nor NOR3 (N4632, N4606, N2834, N846);
xor XOR2 (N4633, N4627, N2090);
xor XOR2 (N4634, N4630, N3834);
not NOT1 (N4635, N4628);
nand NAND4 (N4636, N4608, N90, N2394, N2374);
buf BUF1 (N4637, N4635);
nand NAND4 (N4638, N4626, N1505, N2554, N4068);
nand NAND2 (N4639, N4607, N1287);
and AND4 (N4640, N4639, N4259, N3823, N868);
nor NOR4 (N4641, N4633, N3608, N1156, N3358);
or OR2 (N4642, N4629, N2019);
nand NAND3 (N4643, N4637, N3374, N3770);
nor NOR3 (N4644, N4624, N3258, N3638);
nand NAND4 (N4645, N4634, N1294, N2757, N2531);
or OR3 (N4646, N4643, N1472, N568);
nor NOR2 (N4647, N4641, N2014);
nor NOR3 (N4648, N4646, N1202, N1738);
or OR4 (N4649, N4636, N2530, N1459, N2363);
xor XOR2 (N4650, N4645, N3658);
buf BUF1 (N4651, N4644);
nand NAND3 (N4652, N4651, N3088, N4095);
and AND4 (N4653, N4652, N2607, N205, N654);
xor XOR2 (N4654, N4648, N2312);
nor NOR3 (N4655, N4640, N2400, N3067);
xor XOR2 (N4656, N4647, N1346);
not NOT1 (N4657, N4656);
nand NAND2 (N4658, N4653, N1456);
or OR2 (N4659, N4631, N1746);
or OR2 (N4660, N4642, N973);
nand NAND4 (N4661, N4659, N617, N1145, N1179);
and AND2 (N4662, N4649, N163);
not NOT1 (N4663, N4660);
buf BUF1 (N4664, N4632);
and AND3 (N4665, N4664, N961, N2990);
not NOT1 (N4666, N4655);
buf BUF1 (N4667, N4650);
nor NOR3 (N4668, N4661, N4555, N2045);
and AND4 (N4669, N4667, N2584, N4386, N3761);
not NOT1 (N4670, N4669);
not NOT1 (N4671, N4670);
nor NOR3 (N4672, N4668, N2568, N453);
or OR4 (N4673, N4665, N3757, N1676, N3398);
xor XOR2 (N4674, N4671, N1608);
not NOT1 (N4675, N4674);
xor XOR2 (N4676, N4662, N2688);
nor NOR2 (N4677, N4676, N4026);
nor NOR4 (N4678, N4654, N2636, N4125, N512);
not NOT1 (N4679, N4666);
xor XOR2 (N4680, N4658, N2992);
buf BUF1 (N4681, N4679);
and AND2 (N4682, N4678, N1639);
and AND4 (N4683, N4682, N2340, N3713, N4666);
buf BUF1 (N4684, N4680);
not NOT1 (N4685, N4672);
buf BUF1 (N4686, N4683);
buf BUF1 (N4687, N4686);
xor XOR2 (N4688, N4638, N4542);
or OR4 (N4689, N4685, N3998, N39, N2714);
and AND3 (N4690, N4673, N1902, N4438);
not NOT1 (N4691, N4687);
not NOT1 (N4692, N4691);
xor XOR2 (N4693, N4689, N2337);
xor XOR2 (N4694, N4675, N4305);
nand NAND2 (N4695, N4692, N359);
buf BUF1 (N4696, N4677);
nand NAND3 (N4697, N4695, N3897, N1411);
buf BUF1 (N4698, N4697);
xor XOR2 (N4699, N4693, N3175);
or OR4 (N4700, N4657, N2687, N3517, N3642);
buf BUF1 (N4701, N4700);
or OR4 (N4702, N4684, N2814, N622, N2255);
or OR2 (N4703, N4694, N3302);
buf BUF1 (N4704, N4696);
or OR2 (N4705, N4688, N732);
not NOT1 (N4706, N4704);
or OR4 (N4707, N4705, N2243, N357, N3111);
xor XOR2 (N4708, N4702, N2673);
buf BUF1 (N4709, N4663);
nor NOR4 (N4710, N4708, N1040, N3081, N1251);
or OR2 (N4711, N4709, N4654);
xor XOR2 (N4712, N4698, N1055);
not NOT1 (N4713, N4701);
xor XOR2 (N4714, N4703, N4126);
xor XOR2 (N4715, N4713, N3153);
and AND2 (N4716, N4711, N329);
nor NOR2 (N4717, N4706, N2020);
nor NOR4 (N4718, N4707, N1709, N4615, N2099);
not NOT1 (N4719, N4681);
buf BUF1 (N4720, N4714);
xor XOR2 (N4721, N4712, N3822);
and AND3 (N4722, N4699, N2175, N370);
and AND2 (N4723, N4715, N1644);
or OR4 (N4724, N4710, N158, N3103, N3668);
and AND4 (N4725, N4722, N3714, N3696, N4305);
nor NOR2 (N4726, N4716, N394);
not NOT1 (N4727, N4690);
nand NAND3 (N4728, N4726, N1145, N2023);
nor NOR2 (N4729, N4728, N4257);
buf BUF1 (N4730, N4723);
nand NAND4 (N4731, N4724, N2481, N4532, N2548);
and AND2 (N4732, N4725, N4247);
xor XOR2 (N4733, N4718, N2984);
nor NOR2 (N4734, N4717, N17);
nand NAND3 (N4735, N4720, N3159, N2396);
xor XOR2 (N4736, N4731, N2286);
xor XOR2 (N4737, N4734, N3856);
not NOT1 (N4738, N4727);
and AND3 (N4739, N4736, N3072, N2952);
or OR4 (N4740, N4733, N1125, N1459, N2302);
xor XOR2 (N4741, N4730, N3979);
nor NOR4 (N4742, N4740, N1566, N677, N1664);
nand NAND3 (N4743, N4737, N3778, N4020);
not NOT1 (N4744, N4742);
nand NAND4 (N4745, N4729, N1115, N2258, N636);
xor XOR2 (N4746, N4745, N813);
xor XOR2 (N4747, N4744, N3223);
nor NOR4 (N4748, N4741, N1720, N1187, N2436);
buf BUF1 (N4749, N4735);
nor NOR2 (N4750, N4739, N519);
or OR4 (N4751, N4750, N2435, N812, N4526);
or OR2 (N4752, N4748, N3624);
xor XOR2 (N4753, N4721, N4515);
or OR3 (N4754, N4746, N3413, N1430);
and AND4 (N4755, N4732, N3306, N4054, N484);
or OR4 (N4756, N4738, N681, N4630, N2959);
not NOT1 (N4757, N4755);
buf BUF1 (N4758, N4754);
xor XOR2 (N4759, N4749, N970);
not NOT1 (N4760, N4751);
and AND3 (N4761, N4758, N1797, N4578);
or OR2 (N4762, N4747, N1009);
not NOT1 (N4763, N4752);
nor NOR3 (N4764, N4763, N1156, N2681);
nor NOR2 (N4765, N4764, N4);
or OR3 (N4766, N4743, N1150, N864);
and AND3 (N4767, N4759, N1167, N4271);
nor NOR2 (N4768, N4757, N1674);
nand NAND4 (N4769, N4768, N2031, N3789, N3449);
xor XOR2 (N4770, N4765, N253);
nand NAND3 (N4771, N4770, N422, N246);
nand NAND3 (N4772, N4761, N1482, N1319);
or OR4 (N4773, N4769, N4453, N2475, N959);
nor NOR3 (N4774, N4773, N1313, N1821);
buf BUF1 (N4775, N4771);
buf BUF1 (N4776, N4772);
and AND3 (N4777, N4753, N3119, N2613);
nand NAND3 (N4778, N4774, N3106, N648);
nor NOR2 (N4779, N4762, N4288);
and AND4 (N4780, N4766, N3221, N1341, N2279);
nor NOR3 (N4781, N4756, N3384, N454);
not NOT1 (N4782, N4780);
xor XOR2 (N4783, N4778, N3748);
nand NAND2 (N4784, N4783, N3195);
nor NOR4 (N4785, N4760, N1266, N1538, N967);
xor XOR2 (N4786, N4776, N4369);
not NOT1 (N4787, N4779);
not NOT1 (N4788, N4786);
not NOT1 (N4789, N4784);
nand NAND2 (N4790, N4788, N1657);
nor NOR4 (N4791, N4782, N453, N4712, N4145);
nand NAND4 (N4792, N4785, N1882, N1284, N1426);
or OR2 (N4793, N4789, N329);
buf BUF1 (N4794, N4775);
buf BUF1 (N4795, N4719);
nor NOR4 (N4796, N4787, N4475, N2741, N1671);
buf BUF1 (N4797, N4795);
and AND3 (N4798, N4777, N197, N3009);
nand NAND4 (N4799, N4793, N2206, N3541, N967);
and AND2 (N4800, N4797, N790);
buf BUF1 (N4801, N4798);
buf BUF1 (N4802, N4792);
and AND2 (N4803, N4796, N3030);
buf BUF1 (N4804, N4767);
nor NOR2 (N4805, N4781, N1130);
xor XOR2 (N4806, N4801, N2918);
nand NAND2 (N4807, N4802, N1066);
buf BUF1 (N4808, N4807);
or OR2 (N4809, N4805, N364);
and AND2 (N4810, N4804, N4057);
nor NOR4 (N4811, N4810, N2998, N4060, N886);
and AND4 (N4812, N4794, N4459, N4212, N4323);
and AND3 (N4813, N4803, N3418, N4447);
buf BUF1 (N4814, N4799);
or OR3 (N4815, N4813, N2576, N4765);
xor XOR2 (N4816, N4812, N2198);
and AND2 (N4817, N4815, N4110);
nor NOR2 (N4818, N4806, N2493);
nor NOR2 (N4819, N4811, N2356);
nor NOR4 (N4820, N4818, N4344, N1707, N3307);
and AND4 (N4821, N4800, N730, N1234, N1390);
xor XOR2 (N4822, N4817, N3132);
buf BUF1 (N4823, N4822);
not NOT1 (N4824, N4821);
or OR2 (N4825, N4823, N1022);
xor XOR2 (N4826, N4808, N721);
and AND3 (N4827, N4816, N2367, N2398);
xor XOR2 (N4828, N4824, N1559);
not NOT1 (N4829, N4826);
or OR2 (N4830, N4790, N3354);
buf BUF1 (N4831, N4825);
not NOT1 (N4832, N4831);
nand NAND4 (N4833, N4814, N3782, N897, N3604);
or OR2 (N4834, N4828, N4695);
and AND2 (N4835, N4791, N3764);
nor NOR4 (N4836, N4832, N4280, N3805, N348);
nand NAND3 (N4837, N4827, N3650, N400);
not NOT1 (N4838, N4834);
nand NAND4 (N4839, N4836, N2303, N3787, N3075);
or OR2 (N4840, N4837, N4346);
nand NAND2 (N4841, N4830, N3221);
or OR4 (N4842, N4809, N1063, N3411, N2518);
and AND4 (N4843, N4838, N3369, N3511, N4069);
not NOT1 (N4844, N4835);
and AND4 (N4845, N4844, N1356, N1444, N3878);
nand NAND3 (N4846, N4819, N4780, N2018);
xor XOR2 (N4847, N4829, N2638);
xor XOR2 (N4848, N4845, N836);
and AND4 (N4849, N4843, N2873, N4532, N1302);
and AND2 (N4850, N4847, N796);
not NOT1 (N4851, N4839);
nor NOR3 (N4852, N4833, N2013, N2016);
nand NAND4 (N4853, N4852, N3295, N1619, N3697);
buf BUF1 (N4854, N4820);
xor XOR2 (N4855, N4849, N1206);
not NOT1 (N4856, N4842);
nor NOR4 (N4857, N4854, N3819, N1090, N2660);
nand NAND2 (N4858, N4841, N3670);
not NOT1 (N4859, N4857);
nor NOR2 (N4860, N4856, N3733);
buf BUF1 (N4861, N4840);
and AND3 (N4862, N4848, N559, N2795);
nor NOR4 (N4863, N4853, N4049, N4020, N1746);
nor NOR3 (N4864, N4860, N1864, N1801);
buf BUF1 (N4865, N4851);
nand NAND3 (N4866, N4846, N4407, N4090);
not NOT1 (N4867, N4866);
nor NOR4 (N4868, N4858, N3976, N4347, N2722);
or OR3 (N4869, N4861, N3498, N1248);
nor NOR2 (N4870, N4868, N4421);
nand NAND2 (N4871, N4869, N2423);
not NOT1 (N4872, N4863);
nor NOR3 (N4873, N4855, N3012, N3422);
and AND3 (N4874, N4873, N989, N2816);
or OR2 (N4875, N4850, N4501);
not NOT1 (N4876, N4871);
and AND4 (N4877, N4864, N2409, N3699, N1544);
xor XOR2 (N4878, N4874, N1870);
nand NAND2 (N4879, N4867, N181);
nand NAND2 (N4880, N4879, N3945);
nor NOR3 (N4881, N4876, N281, N553);
or OR3 (N4882, N4878, N1534, N731);
nor NOR3 (N4883, N4882, N3488, N4302);
xor XOR2 (N4884, N4870, N4217);
nor NOR3 (N4885, N4877, N4036, N2648);
nor NOR2 (N4886, N4880, N544);
buf BUF1 (N4887, N4886);
xor XOR2 (N4888, N4859, N1514);
or OR2 (N4889, N4881, N452);
xor XOR2 (N4890, N4887, N2680);
xor XOR2 (N4891, N4889, N2994);
and AND3 (N4892, N4862, N4308, N81);
buf BUF1 (N4893, N4884);
or OR4 (N4894, N4885, N4192, N3592, N2140);
nand NAND3 (N4895, N4872, N236, N4425);
and AND2 (N4896, N4890, N1923);
or OR4 (N4897, N4893, N4081, N620, N3744);
or OR2 (N4898, N4894, N2039);
nor NOR2 (N4899, N4895, N3908);
nand NAND4 (N4900, N4883, N4774, N4538, N4456);
and AND4 (N4901, N4897, N610, N387, N670);
nor NOR3 (N4902, N4899, N2958, N2962);
buf BUF1 (N4903, N4865);
xor XOR2 (N4904, N4903, N3414);
nor NOR2 (N4905, N4901, N1818);
buf BUF1 (N4906, N4904);
nand NAND4 (N4907, N4898, N4333, N2050, N536);
or OR2 (N4908, N4891, N45);
buf BUF1 (N4909, N4905);
xor XOR2 (N4910, N4896, N3719);
nor NOR3 (N4911, N4908, N1096, N3255);
buf BUF1 (N4912, N4911);
nor NOR3 (N4913, N4875, N2184, N2681);
and AND2 (N4914, N4912, N4096);
nand NAND4 (N4915, N4909, N2286, N4560, N2179);
xor XOR2 (N4916, N4888, N2601);
xor XOR2 (N4917, N4914, N2688);
buf BUF1 (N4918, N4915);
xor XOR2 (N4919, N4917, N3353);
nor NOR2 (N4920, N4913, N4783);
not NOT1 (N4921, N4920);
and AND3 (N4922, N4906, N3184, N4605);
buf BUF1 (N4923, N4900);
and AND3 (N4924, N4907, N503, N3888);
buf BUF1 (N4925, N4922);
xor XOR2 (N4926, N4902, N3843);
buf BUF1 (N4927, N4919);
xor XOR2 (N4928, N4926, N1272);
nand NAND4 (N4929, N4927, N3168, N1158, N4784);
and AND4 (N4930, N4925, N3376, N3456, N694);
nor NOR2 (N4931, N4916, N2320);
and AND3 (N4932, N4928, N537, N916);
nand NAND4 (N4933, N4910, N2975, N4895, N1101);
buf BUF1 (N4934, N4930);
or OR3 (N4935, N4923, N4674, N4817);
or OR4 (N4936, N4929, N1433, N1345, N3822);
nand NAND2 (N4937, N4918, N4327);
and AND3 (N4938, N4931, N3979, N4178);
xor XOR2 (N4939, N4935, N4551);
not NOT1 (N4940, N4932);
or OR4 (N4941, N4934, N2547, N2168, N2957);
nand NAND2 (N4942, N4940, N3462);
and AND3 (N4943, N4942, N3328, N925);
xor XOR2 (N4944, N4924, N1239);
not NOT1 (N4945, N4943);
not NOT1 (N4946, N4939);
nand NAND3 (N4947, N4945, N4529, N4017);
and AND2 (N4948, N4921, N137);
xor XOR2 (N4949, N4944, N3052);
nand NAND2 (N4950, N4936, N4470);
buf BUF1 (N4951, N4941);
or OR4 (N4952, N4950, N1731, N3068, N1559);
xor XOR2 (N4953, N4947, N2791);
or OR3 (N4954, N4952, N4558, N2935);
not NOT1 (N4955, N4933);
nand NAND3 (N4956, N4948, N2052, N49);
nor NOR4 (N4957, N4949, N2957, N3205, N1760);
nand NAND4 (N4958, N4956, N4768, N341, N516);
and AND2 (N4959, N4955, N2266);
xor XOR2 (N4960, N4938, N247);
buf BUF1 (N4961, N4937);
buf BUF1 (N4962, N4953);
xor XOR2 (N4963, N4951, N4785);
not NOT1 (N4964, N4946);
nor NOR2 (N4965, N4964, N717);
or OR2 (N4966, N4961, N4718);
or OR4 (N4967, N4966, N594, N740, N4598);
and AND4 (N4968, N4960, N3297, N3443, N2173);
buf BUF1 (N4969, N4965);
buf BUF1 (N4970, N4962);
xor XOR2 (N4971, N4970, N3403);
buf BUF1 (N4972, N4959);
nor NOR2 (N4973, N4968, N90);
xor XOR2 (N4974, N4957, N4489);
not NOT1 (N4975, N4974);
and AND3 (N4976, N4958, N3767, N4255);
not NOT1 (N4977, N4967);
not NOT1 (N4978, N4977);
xor XOR2 (N4979, N4978, N21);
and AND4 (N4980, N4975, N2063, N4948, N661);
xor XOR2 (N4981, N4971, N2345);
nand NAND2 (N4982, N4969, N160);
nand NAND2 (N4983, N4979, N2295);
or OR2 (N4984, N4981, N1812);
nor NOR4 (N4985, N4972, N476, N866, N1209);
buf BUF1 (N4986, N4976);
nor NOR2 (N4987, N4963, N2658);
nor NOR2 (N4988, N4973, N1561);
not NOT1 (N4989, N4954);
or OR4 (N4990, N4986, N678, N510, N3416);
and AND4 (N4991, N4988, N3000, N4428, N2415);
or OR2 (N4992, N4991, N498);
not NOT1 (N4993, N4987);
or OR3 (N4994, N4989, N453, N1176);
buf BUF1 (N4995, N4980);
xor XOR2 (N4996, N4994, N1995);
xor XOR2 (N4997, N4992, N601);
not NOT1 (N4998, N4892);
nor NOR2 (N4999, N4984, N3279);
nand NAND4 (N5000, N4997, N4334, N2521, N2114);
not NOT1 (N5001, N5000);
buf BUF1 (N5002, N4982);
nor NOR2 (N5003, N5002, N1052);
nor NOR4 (N5004, N5001, N4763, N2233, N2351);
xor XOR2 (N5005, N5004, N3115);
nand NAND4 (N5006, N4993, N3152, N1378, N4549);
or OR3 (N5007, N4985, N2053, N3845);
buf BUF1 (N5008, N5003);
or OR4 (N5009, N5005, N331, N404, N599);
nand NAND3 (N5010, N5008, N3912, N923);
nor NOR3 (N5011, N4998, N2250, N1979);
xor XOR2 (N5012, N4990, N1622);
or OR4 (N5013, N5007, N2706, N3554, N1176);
not NOT1 (N5014, N5010);
xor XOR2 (N5015, N4995, N162);
buf BUF1 (N5016, N5012);
and AND4 (N5017, N5009, N3198, N3434, N4850);
not NOT1 (N5018, N4983);
not NOT1 (N5019, N5018);
or OR2 (N5020, N4996, N1356);
xor XOR2 (N5021, N5014, N3906);
buf BUF1 (N5022, N5015);
and AND3 (N5023, N5020, N952, N588);
or OR4 (N5024, N5016, N3283, N4198, N512);
or OR4 (N5025, N5021, N4983, N378, N4658);
and AND4 (N5026, N4999, N1324, N441, N690);
nor NOR2 (N5027, N5019, N2648);
nor NOR2 (N5028, N5026, N1016);
or OR3 (N5029, N5028, N4564, N3288);
or OR3 (N5030, N5017, N3679, N3262);
not NOT1 (N5031, N5027);
not NOT1 (N5032, N5023);
or OR3 (N5033, N5032, N609, N3028);
buf BUF1 (N5034, N5013);
not NOT1 (N5035, N5033);
xor XOR2 (N5036, N5030, N2217);
nor NOR2 (N5037, N5031, N2430);
xor XOR2 (N5038, N5036, N556);
or OR4 (N5039, N5038, N3554, N1743, N2034);
and AND3 (N5040, N5029, N2616, N2054);
nor NOR3 (N5041, N5006, N3588, N2411);
not NOT1 (N5042, N5041);
xor XOR2 (N5043, N5022, N2673);
xor XOR2 (N5044, N5024, N3906);
or OR2 (N5045, N5011, N1285);
or OR3 (N5046, N5035, N4263, N3581);
or OR3 (N5047, N5025, N3175, N456);
nand NAND2 (N5048, N5044, N4198);
not NOT1 (N5049, N5042);
nor NOR2 (N5050, N5049, N3399);
and AND4 (N5051, N5039, N4541, N3472, N488);
or OR4 (N5052, N5046, N222, N933, N2166);
nand NAND4 (N5053, N5034, N2801, N3596, N87);
not NOT1 (N5054, N5048);
or OR2 (N5055, N5053, N3866);
not NOT1 (N5056, N5051);
nor NOR4 (N5057, N5055, N4560, N1212, N2952);
nor NOR4 (N5058, N5052, N2925, N427, N269);
not NOT1 (N5059, N5043);
buf BUF1 (N5060, N5059);
not NOT1 (N5061, N5058);
nor NOR4 (N5062, N5054, N4178, N2768, N3725);
nand NAND4 (N5063, N5057, N4227, N1125, N1052);
nand NAND4 (N5064, N5040, N225, N3961, N356);
not NOT1 (N5065, N5045);
buf BUF1 (N5066, N5065);
nor NOR3 (N5067, N5061, N2580, N2646);
xor XOR2 (N5068, N5064, N2865);
buf BUF1 (N5069, N5050);
not NOT1 (N5070, N5056);
and AND3 (N5071, N5060, N1252, N1867);
not NOT1 (N5072, N5037);
xor XOR2 (N5073, N5067, N4041);
or OR2 (N5074, N5066, N1410);
or OR3 (N5075, N5072, N4153, N4844);
buf BUF1 (N5076, N5070);
xor XOR2 (N5077, N5068, N1646);
xor XOR2 (N5078, N5076, N791);
nor NOR4 (N5079, N5063, N3159, N1349, N3930);
buf BUF1 (N5080, N5078);
buf BUF1 (N5081, N5047);
and AND3 (N5082, N5074, N2323, N3377);
nor NOR3 (N5083, N5077, N1655, N104);
nor NOR2 (N5084, N5082, N4547);
nand NAND3 (N5085, N5075, N2589, N2578);
nor NOR3 (N5086, N5069, N136, N3425);
and AND3 (N5087, N5071, N1223, N305);
buf BUF1 (N5088, N5081);
nand NAND3 (N5089, N5083, N4331, N2947);
nand NAND4 (N5090, N5062, N740, N1251, N3267);
nand NAND2 (N5091, N5085, N4134);
nor NOR4 (N5092, N5089, N2052, N1092, N3450);
nand NAND4 (N5093, N5080, N4284, N4752, N4300);
not NOT1 (N5094, N5084);
buf BUF1 (N5095, N5094);
or OR4 (N5096, N5093, N2504, N2717, N79);
or OR3 (N5097, N5091, N63, N290);
nor NOR3 (N5098, N5073, N1254, N4960);
or OR3 (N5099, N5098, N1737, N340);
xor XOR2 (N5100, N5095, N2577);
nand NAND4 (N5101, N5090, N5077, N1873, N4627);
or OR2 (N5102, N5079, N117);
or OR2 (N5103, N5088, N307);
buf BUF1 (N5104, N5102);
nand NAND4 (N5105, N5092, N612, N2759, N4151);
or OR4 (N5106, N5103, N940, N3449, N2746);
buf BUF1 (N5107, N5086);
nand NAND2 (N5108, N5087, N3927);
and AND3 (N5109, N5099, N1892, N1132);
or OR3 (N5110, N5096, N3351, N1556);
nand NAND4 (N5111, N5110, N1804, N4538, N1081);
and AND2 (N5112, N5111, N4704);
nand NAND4 (N5113, N5108, N2942, N3474, N1069);
and AND3 (N5114, N5112, N1470, N232);
nand NAND4 (N5115, N5106, N4794, N1705, N1217);
nor NOR4 (N5116, N5115, N1519, N2790, N3398);
not NOT1 (N5117, N5107);
xor XOR2 (N5118, N5109, N2049);
not NOT1 (N5119, N5114);
nand NAND3 (N5120, N5119, N1885, N51);
nor NOR3 (N5121, N5113, N4545, N4063);
or OR4 (N5122, N5104, N583, N1427, N4521);
or OR3 (N5123, N5121, N4839, N3702);
not NOT1 (N5124, N5105);
buf BUF1 (N5125, N5100);
xor XOR2 (N5126, N5123, N294);
and AND2 (N5127, N5118, N3961);
or OR3 (N5128, N5101, N2607, N979);
nor NOR2 (N5129, N5117, N4554);
or OR3 (N5130, N5116, N3827, N1926);
not NOT1 (N5131, N5129);
and AND4 (N5132, N5124, N2412, N2379, N2104);
nor NOR4 (N5133, N5097, N3246, N525, N564);
or OR4 (N5134, N5127, N679, N4330, N2840);
buf BUF1 (N5135, N5132);
buf BUF1 (N5136, N5128);
buf BUF1 (N5137, N5126);
xor XOR2 (N5138, N5125, N3968);
not NOT1 (N5139, N5131);
or OR2 (N5140, N5138, N2313);
nor NOR4 (N5141, N5134, N2223, N3138, N5045);
nor NOR2 (N5142, N5133, N2216);
not NOT1 (N5143, N5120);
nor NOR2 (N5144, N5142, N128);
nand NAND4 (N5145, N5136, N1511, N2418, N3832);
nand NAND3 (N5146, N5140, N1192, N4016);
and AND2 (N5147, N5130, N1932);
nor NOR2 (N5148, N5135, N2589);
or OR3 (N5149, N5137, N3930, N1163);
or OR4 (N5150, N5145, N1281, N1853, N2874);
not NOT1 (N5151, N5146);
not NOT1 (N5152, N5122);
and AND4 (N5153, N5152, N2783, N3235, N360);
and AND4 (N5154, N5141, N5133, N3491, N1771);
buf BUF1 (N5155, N5154);
not NOT1 (N5156, N5149);
buf BUF1 (N5157, N5150);
or OR4 (N5158, N5155, N516, N1833, N1173);
not NOT1 (N5159, N5151);
nand NAND4 (N5160, N5148, N2646, N3461, N4668);
nor NOR3 (N5161, N5139, N4951, N148);
not NOT1 (N5162, N5143);
or OR3 (N5163, N5144, N4786, N2198);
not NOT1 (N5164, N5161);
and AND2 (N5165, N5157, N2158);
xor XOR2 (N5166, N5164, N4273);
and AND3 (N5167, N5160, N4765, N2705);
or OR3 (N5168, N5166, N1369, N4682);
or OR4 (N5169, N5147, N613, N968, N2496);
nor NOR2 (N5170, N5169, N5131);
or OR4 (N5171, N5156, N4244, N45, N865);
buf BUF1 (N5172, N5162);
and AND4 (N5173, N5167, N310, N3240, N4429);
nor NOR3 (N5174, N5170, N1357, N2836);
xor XOR2 (N5175, N5158, N1291);
nand NAND4 (N5176, N5175, N2544, N4052, N4878);
and AND2 (N5177, N5172, N3929);
and AND3 (N5178, N5165, N4348, N4540);
xor XOR2 (N5179, N5153, N2103);
and AND4 (N5180, N5159, N2867, N4466, N1394);
not NOT1 (N5181, N5176);
or OR4 (N5182, N5171, N1903, N4736, N5007);
nor NOR3 (N5183, N5174, N1708, N4540);
nor NOR4 (N5184, N5163, N13, N4211, N379);
and AND4 (N5185, N5181, N338, N1332, N3060);
and AND3 (N5186, N5173, N10, N3621);
buf BUF1 (N5187, N5182);
or OR2 (N5188, N5183, N2096);
xor XOR2 (N5189, N5180, N2050);
buf BUF1 (N5190, N5179);
xor XOR2 (N5191, N5190, N3253);
and AND4 (N5192, N5188, N908, N1032, N1366);
and AND4 (N5193, N5192, N1261, N3106, N4540);
buf BUF1 (N5194, N5184);
nand NAND2 (N5195, N5185, N818);
nand NAND2 (N5196, N5187, N2219);
buf BUF1 (N5197, N5194);
or OR2 (N5198, N5177, N857);
buf BUF1 (N5199, N5168);
xor XOR2 (N5200, N5189, N164);
buf BUF1 (N5201, N5186);
or OR3 (N5202, N5197, N2563, N1600);
buf BUF1 (N5203, N5196);
nor NOR3 (N5204, N5202, N1638, N4402);
and AND3 (N5205, N5204, N3701, N3469);
buf BUF1 (N5206, N5203);
and AND3 (N5207, N5206, N3255, N3678);
nand NAND3 (N5208, N5198, N4882, N1694);
buf BUF1 (N5209, N5205);
buf BUF1 (N5210, N5209);
and AND4 (N5211, N5200, N3816, N1097, N4648);
nor NOR3 (N5212, N5193, N2135, N3866);
nor NOR2 (N5213, N5212, N49);
nor NOR3 (N5214, N5195, N1502, N3855);
nor NOR4 (N5215, N5178, N4098, N3839, N1521);
nor NOR4 (N5216, N5191, N2813, N4122, N4851);
nand NAND3 (N5217, N5211, N3750, N4174);
buf BUF1 (N5218, N5207);
and AND2 (N5219, N5216, N5207);
buf BUF1 (N5220, N5217);
nor NOR2 (N5221, N5210, N320);
nor NOR3 (N5222, N5221, N4004, N3346);
buf BUF1 (N5223, N5208);
and AND4 (N5224, N5201, N3620, N3945, N1887);
buf BUF1 (N5225, N5220);
xor XOR2 (N5226, N5225, N957);
nor NOR3 (N5227, N5213, N1214, N1357);
xor XOR2 (N5228, N5224, N1387);
not NOT1 (N5229, N5223);
or OR4 (N5230, N5228, N1164, N4215, N1730);
nand NAND3 (N5231, N5227, N127, N3410);
or OR2 (N5232, N5199, N1763);
xor XOR2 (N5233, N5231, N1197);
or OR2 (N5234, N5222, N1121);
not NOT1 (N5235, N5229);
or OR3 (N5236, N5226, N1246, N663);
or OR2 (N5237, N5234, N2685);
not NOT1 (N5238, N5230);
not NOT1 (N5239, N5236);
nor NOR3 (N5240, N5235, N3662, N4765);
xor XOR2 (N5241, N5240, N3587);
or OR3 (N5242, N5214, N900, N4239);
xor XOR2 (N5243, N5218, N1379);
buf BUF1 (N5244, N5232);
not NOT1 (N5245, N5239);
or OR3 (N5246, N5244, N666, N3725);
nor NOR2 (N5247, N5246, N402);
or OR2 (N5248, N5237, N1604);
not NOT1 (N5249, N5219);
nand NAND2 (N5250, N5248, N3716);
and AND4 (N5251, N5249, N5021, N2238, N2988);
buf BUF1 (N5252, N5215);
nor NOR3 (N5253, N5251, N1041, N2797);
xor XOR2 (N5254, N5250, N1117);
xor XOR2 (N5255, N5247, N3683);
and AND3 (N5256, N5252, N1520, N51);
or OR4 (N5257, N5238, N578, N204, N2725);
nand NAND4 (N5258, N5242, N692, N2526, N2741);
buf BUF1 (N5259, N5245);
xor XOR2 (N5260, N5255, N4422);
buf BUF1 (N5261, N5241);
nor NOR4 (N5262, N5258, N590, N2562, N218);
xor XOR2 (N5263, N5257, N1704);
or OR4 (N5264, N5256, N4217, N2820, N1517);
buf BUF1 (N5265, N5260);
nor NOR2 (N5266, N5253, N2033);
and AND4 (N5267, N5264, N3798, N4597, N1855);
not NOT1 (N5268, N5262);
nand NAND2 (N5269, N5267, N4390);
nor NOR2 (N5270, N5259, N4641);
buf BUF1 (N5271, N5268);
nand NAND3 (N5272, N5261, N1904, N3077);
buf BUF1 (N5273, N5243);
nor NOR4 (N5274, N5263, N4974, N2602, N3061);
xor XOR2 (N5275, N5254, N1504);
buf BUF1 (N5276, N5272);
and AND4 (N5277, N5269, N4624, N3114, N4725);
nor NOR2 (N5278, N5274, N3346);
buf BUF1 (N5279, N5273);
xor XOR2 (N5280, N5275, N4348);
and AND2 (N5281, N5270, N925);
or OR2 (N5282, N5279, N4839);
buf BUF1 (N5283, N5266);
buf BUF1 (N5284, N5265);
xor XOR2 (N5285, N5271, N1562);
or OR3 (N5286, N5281, N3037, N3233);
nor NOR3 (N5287, N5280, N4658, N692);
buf BUF1 (N5288, N5285);
or OR4 (N5289, N5287, N626, N4348, N208);
buf BUF1 (N5290, N5286);
or OR3 (N5291, N5284, N3019, N2127);
xor XOR2 (N5292, N5291, N4249);
or OR4 (N5293, N5277, N2085, N576, N2879);
and AND2 (N5294, N5293, N4364);
nor NOR2 (N5295, N5288, N4909);
nor NOR2 (N5296, N5292, N765);
nor NOR4 (N5297, N5290, N4397, N102, N4442);
buf BUF1 (N5298, N5278);
nor NOR4 (N5299, N5289, N376, N3251, N2926);
nand NAND2 (N5300, N5296, N3803);
xor XOR2 (N5301, N5283, N932);
not NOT1 (N5302, N5299);
nor NOR2 (N5303, N5302, N4731);
and AND2 (N5304, N5301, N4841);
and AND2 (N5305, N5294, N2026);
or OR3 (N5306, N5295, N271, N973);
nor NOR2 (N5307, N5276, N868);
or OR2 (N5308, N5297, N24);
or OR3 (N5309, N5298, N3083, N2769);
and AND4 (N5310, N5303, N228, N4550, N450);
buf BUF1 (N5311, N5307);
nor NOR2 (N5312, N5305, N2074);
xor XOR2 (N5313, N5311, N3627);
or OR3 (N5314, N5312, N442, N1128);
xor XOR2 (N5315, N5309, N1047);
not NOT1 (N5316, N5306);
not NOT1 (N5317, N5315);
buf BUF1 (N5318, N5308);
not NOT1 (N5319, N5310);
xor XOR2 (N5320, N5233, N4803);
and AND2 (N5321, N5320, N302);
or OR3 (N5322, N5314, N4045, N1398);
nand NAND2 (N5323, N5318, N1938);
xor XOR2 (N5324, N5323, N3444);
and AND3 (N5325, N5304, N1365, N3801);
not NOT1 (N5326, N5313);
xor XOR2 (N5327, N5324, N3285);
or OR3 (N5328, N5327, N3534, N207);
and AND2 (N5329, N5300, N1652);
nor NOR4 (N5330, N5321, N1455, N994, N3286);
and AND2 (N5331, N5282, N3578);
xor XOR2 (N5332, N5331, N4242);
nor NOR3 (N5333, N5325, N704, N3979);
not NOT1 (N5334, N5330);
xor XOR2 (N5335, N5329, N38);
or OR3 (N5336, N5334, N2089, N4740);
xor XOR2 (N5337, N5316, N4876);
and AND3 (N5338, N5322, N1443, N415);
or OR4 (N5339, N5333, N2694, N2635, N1195);
xor XOR2 (N5340, N5336, N2452);
buf BUF1 (N5341, N5319);
nor NOR3 (N5342, N5332, N3023, N1975);
nor NOR4 (N5343, N5341, N464, N1319, N600);
nor NOR4 (N5344, N5326, N4972, N536, N1743);
nor NOR4 (N5345, N5342, N951, N2615, N442);
not NOT1 (N5346, N5345);
not NOT1 (N5347, N5340);
not NOT1 (N5348, N5344);
or OR2 (N5349, N5337, N3861);
xor XOR2 (N5350, N5346, N5202);
buf BUF1 (N5351, N5317);
nand NAND2 (N5352, N5343, N4260);
nand NAND2 (N5353, N5350, N4148);
buf BUF1 (N5354, N5352);
nand NAND3 (N5355, N5351, N1072, N340);
buf BUF1 (N5356, N5335);
buf BUF1 (N5357, N5356);
nor NOR4 (N5358, N5328, N2899, N2619, N5275);
or OR4 (N5359, N5357, N1973, N4824, N32);
xor XOR2 (N5360, N5339, N1416);
nor NOR3 (N5361, N5358, N5247, N4351);
nand NAND2 (N5362, N5355, N3277);
and AND4 (N5363, N5348, N4754, N361, N54);
xor XOR2 (N5364, N5362, N1781);
buf BUF1 (N5365, N5360);
xor XOR2 (N5366, N5363, N109);
nor NOR3 (N5367, N5338, N4106, N2481);
or OR3 (N5368, N5354, N3250, N5187);
nand NAND3 (N5369, N5353, N3302, N3250);
and AND4 (N5370, N5365, N4994, N4977, N4771);
not NOT1 (N5371, N5349);
or OR4 (N5372, N5368, N2131, N3633, N939);
or OR2 (N5373, N5367, N3128);
xor XOR2 (N5374, N5361, N537);
not NOT1 (N5375, N5370);
buf BUF1 (N5376, N5373);
nor NOR2 (N5377, N5366, N4549);
nand NAND3 (N5378, N5364, N4420, N3210);
nor NOR2 (N5379, N5377, N1572);
or OR4 (N5380, N5372, N4722, N93, N3195);
not NOT1 (N5381, N5375);
xor XOR2 (N5382, N5369, N4649);
buf BUF1 (N5383, N5376);
xor XOR2 (N5384, N5382, N4905);
nand NAND3 (N5385, N5347, N2493, N5138);
xor XOR2 (N5386, N5381, N2462);
or OR3 (N5387, N5385, N4106, N2543);
xor XOR2 (N5388, N5374, N2784);
or OR3 (N5389, N5383, N4730, N4963);
not NOT1 (N5390, N5386);
nand NAND3 (N5391, N5380, N2706, N4515);
xor XOR2 (N5392, N5371, N1015);
or OR4 (N5393, N5359, N3291, N1736, N2286);
or OR3 (N5394, N5387, N4834, N4137);
buf BUF1 (N5395, N5378);
xor XOR2 (N5396, N5389, N1566);
or OR3 (N5397, N5391, N4444, N1094);
or OR4 (N5398, N5396, N473, N842, N2632);
buf BUF1 (N5399, N5395);
xor XOR2 (N5400, N5398, N4513);
buf BUF1 (N5401, N5388);
and AND2 (N5402, N5393, N4347);
nand NAND3 (N5403, N5384, N2448, N2931);
and AND4 (N5404, N5400, N3769, N3735, N3911);
not NOT1 (N5405, N5399);
nor NOR3 (N5406, N5403, N400, N416);
not NOT1 (N5407, N5379);
not NOT1 (N5408, N5401);
nand NAND3 (N5409, N5390, N3561, N5018);
or OR2 (N5410, N5405, N4853);
nor NOR3 (N5411, N5394, N2509, N3208);
or OR3 (N5412, N5392, N3672, N4060);
and AND2 (N5413, N5411, N3178);
nor NOR2 (N5414, N5407, N5063);
nor NOR3 (N5415, N5406, N2500, N629);
not NOT1 (N5416, N5414);
and AND3 (N5417, N5402, N4289, N1610);
not NOT1 (N5418, N5408);
and AND3 (N5419, N5417, N5076, N4270);
nand NAND4 (N5420, N5410, N3534, N4509, N3421);
xor XOR2 (N5421, N5419, N1221);
and AND2 (N5422, N5413, N1702);
or OR4 (N5423, N5422, N3668, N2352, N1880);
and AND2 (N5424, N5415, N710);
xor XOR2 (N5425, N5416, N2916);
nand NAND4 (N5426, N5404, N363, N3988, N3484);
nand NAND2 (N5427, N5409, N583);
xor XOR2 (N5428, N5420, N329);
nand NAND2 (N5429, N5423, N4149);
buf BUF1 (N5430, N5418);
or OR2 (N5431, N5412, N3926);
xor XOR2 (N5432, N5427, N2466);
buf BUF1 (N5433, N5397);
or OR4 (N5434, N5428, N260, N2000, N4960);
buf BUF1 (N5435, N5425);
buf BUF1 (N5436, N5430);
buf BUF1 (N5437, N5431);
or OR3 (N5438, N5421, N1382, N164);
and AND2 (N5439, N5424, N942);
xor XOR2 (N5440, N5429, N3197);
buf BUF1 (N5441, N5435);
buf BUF1 (N5442, N5436);
nor NOR3 (N5443, N5432, N1615, N4138);
buf BUF1 (N5444, N5442);
buf BUF1 (N5445, N5440);
or OR4 (N5446, N5441, N239, N2638, N3806);
nand NAND4 (N5447, N5445, N1365, N818, N4683);
xor XOR2 (N5448, N5446, N5420);
xor XOR2 (N5449, N5444, N1170);
nor NOR3 (N5450, N5447, N1513, N5108);
or OR2 (N5451, N5439, N4890);
xor XOR2 (N5452, N5449, N5228);
or OR2 (N5453, N5448, N4066);
buf BUF1 (N5454, N5426);
xor XOR2 (N5455, N5433, N2862);
nor NOR2 (N5456, N5434, N3320);
not NOT1 (N5457, N5453);
or OR4 (N5458, N5456, N445, N1889, N2660);
nor NOR3 (N5459, N5438, N1440, N5211);
nor NOR4 (N5460, N5450, N80, N2746, N3559);
nor NOR3 (N5461, N5437, N1605, N4155);
and AND3 (N5462, N5443, N2154, N4245);
xor XOR2 (N5463, N5452, N2440);
nor NOR3 (N5464, N5463, N1905, N2894);
not NOT1 (N5465, N5461);
nand NAND3 (N5466, N5455, N2007, N938);
nor NOR2 (N5467, N5462, N4896);
nor NOR2 (N5468, N5451, N3287);
nand NAND4 (N5469, N5459, N929, N2655, N1738);
nand NAND2 (N5470, N5467, N1611);
nor NOR4 (N5471, N5466, N4031, N1521, N3537);
nor NOR3 (N5472, N5469, N1031, N718);
buf BUF1 (N5473, N5464);
buf BUF1 (N5474, N5460);
buf BUF1 (N5475, N5473);
or OR3 (N5476, N5468, N2235, N3853);
nor NOR4 (N5477, N5475, N3449, N4397, N2706);
not NOT1 (N5478, N5477);
not NOT1 (N5479, N5458);
buf BUF1 (N5480, N5454);
and AND3 (N5481, N5478, N2696, N4124);
nor NOR4 (N5482, N5457, N750, N3480, N160);
nand NAND4 (N5483, N5480, N3653, N5068, N235);
buf BUF1 (N5484, N5481);
not NOT1 (N5485, N5474);
or OR3 (N5486, N5482, N1552, N687);
buf BUF1 (N5487, N5476);
or OR2 (N5488, N5472, N4070);
not NOT1 (N5489, N5487);
and AND3 (N5490, N5486, N974, N278);
nor NOR4 (N5491, N5490, N3633, N267, N4599);
and AND4 (N5492, N5489, N76, N5348, N4462);
or OR2 (N5493, N5470, N3861);
or OR4 (N5494, N5488, N3438, N4457, N4788);
and AND4 (N5495, N5465, N5024, N5066, N3635);
nand NAND3 (N5496, N5495, N5345, N4461);
and AND3 (N5497, N5494, N3717, N3810);
nand NAND2 (N5498, N5492, N4758);
nand NAND2 (N5499, N5491, N1123);
nand NAND2 (N5500, N5497, N2473);
nor NOR2 (N5501, N5479, N3715);
nor NOR4 (N5502, N5483, N3362, N125, N2619);
not NOT1 (N5503, N5485);
and AND4 (N5504, N5496, N1406, N4446, N5285);
or OR4 (N5505, N5493, N1771, N1294, N5171);
buf BUF1 (N5506, N5500);
xor XOR2 (N5507, N5484, N777);
buf BUF1 (N5508, N5501);
nand NAND4 (N5509, N5502, N3842, N1224, N4427);
nand NAND4 (N5510, N5498, N635, N2391, N3305);
or OR4 (N5511, N5509, N4174, N3993, N1542);
and AND4 (N5512, N5508, N2600, N804, N2428);
or OR4 (N5513, N5499, N1719, N3621, N1170);
nand NAND4 (N5514, N5503, N3496, N2060, N2935);
xor XOR2 (N5515, N5471, N620);
xor XOR2 (N5516, N5507, N3927);
xor XOR2 (N5517, N5504, N3222);
buf BUF1 (N5518, N5505);
buf BUF1 (N5519, N5510);
nand NAND2 (N5520, N5517, N1461);
not NOT1 (N5521, N5511);
or OR2 (N5522, N5518, N3725);
nand NAND2 (N5523, N5506, N4416);
xor XOR2 (N5524, N5515, N4280);
nand NAND2 (N5525, N5519, N3803);
xor XOR2 (N5526, N5524, N3304);
not NOT1 (N5527, N5513);
or OR4 (N5528, N5525, N5076, N1922, N2675);
nor NOR3 (N5529, N5528, N5516, N3669);
not NOT1 (N5530, N4250);
and AND3 (N5531, N5526, N3121, N1714);
nand NAND4 (N5532, N5512, N5348, N5373, N2539);
buf BUF1 (N5533, N5529);
not NOT1 (N5534, N5521);
and AND3 (N5535, N5523, N1668, N2189);
nor NOR2 (N5536, N5527, N4363);
xor XOR2 (N5537, N5530, N4198);
xor XOR2 (N5538, N5520, N1594);
or OR4 (N5539, N5535, N5247, N5011, N5524);
or OR4 (N5540, N5534, N2641, N3108, N2113);
not NOT1 (N5541, N5536);
or OR2 (N5542, N5537, N279);
or OR4 (N5543, N5531, N2139, N4026, N1505);
xor XOR2 (N5544, N5532, N4110);
buf BUF1 (N5545, N5538);
or OR3 (N5546, N5539, N3706, N5282);
and AND4 (N5547, N5542, N4508, N3078, N3157);
buf BUF1 (N5548, N5533);
and AND2 (N5549, N5522, N1507);
buf BUF1 (N5550, N5544);
nor NOR3 (N5551, N5549, N35, N3247);
xor XOR2 (N5552, N5550, N5527);
or OR3 (N5553, N5540, N2707, N3477);
not NOT1 (N5554, N5543);
nor NOR2 (N5555, N5547, N1702);
xor XOR2 (N5556, N5553, N423);
or OR3 (N5557, N5555, N2569, N445);
and AND4 (N5558, N5548, N3757, N732, N796);
buf BUF1 (N5559, N5514);
xor XOR2 (N5560, N5557, N1729);
and AND3 (N5561, N5554, N3267, N4550);
xor XOR2 (N5562, N5561, N260);
nand NAND4 (N5563, N5558, N997, N5230, N2402);
xor XOR2 (N5564, N5541, N880);
buf BUF1 (N5565, N5560);
or OR4 (N5566, N5546, N3261, N415, N1583);
buf BUF1 (N5567, N5559);
or OR2 (N5568, N5552, N2004);
or OR4 (N5569, N5565, N228, N3146, N3978);
nand NAND4 (N5570, N5551, N4588, N1138, N577);
or OR3 (N5571, N5564, N453, N2709);
not NOT1 (N5572, N5570);
nor NOR4 (N5573, N5556, N3310, N3256, N4064);
buf BUF1 (N5574, N5562);
nor NOR3 (N5575, N5569, N4830, N5046);
nand NAND4 (N5576, N5545, N1317, N2088, N2240);
or OR3 (N5577, N5566, N3772, N796);
or OR4 (N5578, N5568, N3741, N541, N2388);
not NOT1 (N5579, N5576);
buf BUF1 (N5580, N5575);
xor XOR2 (N5581, N5567, N3586);
and AND2 (N5582, N5572, N4336);
buf BUF1 (N5583, N5573);
xor XOR2 (N5584, N5571, N291);
xor XOR2 (N5585, N5563, N4456);
and AND2 (N5586, N5579, N607);
xor XOR2 (N5587, N5574, N2583);
nor NOR2 (N5588, N5587, N3171);
nand NAND2 (N5589, N5583, N4308);
buf BUF1 (N5590, N5580);
xor XOR2 (N5591, N5577, N22);
and AND3 (N5592, N5591, N1089, N3605);
and AND2 (N5593, N5581, N2961);
xor XOR2 (N5594, N5592, N2369);
xor XOR2 (N5595, N5578, N3743);
not NOT1 (N5596, N5582);
not NOT1 (N5597, N5585);
buf BUF1 (N5598, N5586);
not NOT1 (N5599, N5589);
xor XOR2 (N5600, N5598, N98);
buf BUF1 (N5601, N5590);
nor NOR4 (N5602, N5596, N1503, N191, N3999);
not NOT1 (N5603, N5601);
xor XOR2 (N5604, N5593, N2429);
nand NAND2 (N5605, N5588, N1317);
or OR2 (N5606, N5599, N3528);
xor XOR2 (N5607, N5597, N1512);
buf BUF1 (N5608, N5600);
and AND4 (N5609, N5594, N4132, N4367, N2866);
xor XOR2 (N5610, N5607, N3147);
not NOT1 (N5611, N5606);
not NOT1 (N5612, N5602);
nor NOR4 (N5613, N5611, N1311, N3412, N1687);
xor XOR2 (N5614, N5613, N519);
nor NOR4 (N5615, N5610, N4793, N5307, N1500);
xor XOR2 (N5616, N5608, N4005);
and AND3 (N5617, N5612, N5002, N1273);
buf BUF1 (N5618, N5615);
buf BUF1 (N5619, N5617);
not NOT1 (N5620, N5619);
buf BUF1 (N5621, N5614);
buf BUF1 (N5622, N5605);
not NOT1 (N5623, N5620);
nand NAND2 (N5624, N5584, N2587);
and AND2 (N5625, N5622, N4838);
xor XOR2 (N5626, N5595, N5564);
buf BUF1 (N5627, N5621);
nor NOR3 (N5628, N5616, N1543, N2505);
nor NOR2 (N5629, N5626, N3070);
nor NOR4 (N5630, N5618, N757, N1495, N5169);
or OR4 (N5631, N5623, N2388, N4920, N1515);
xor XOR2 (N5632, N5630, N1567);
or OR4 (N5633, N5627, N5362, N5075, N1128);
or OR2 (N5634, N5604, N40);
or OR4 (N5635, N5634, N3219, N5143, N73);
xor XOR2 (N5636, N5625, N868);
nor NOR4 (N5637, N5629, N2450, N5633, N5441);
and AND4 (N5638, N1537, N5492, N1076, N3612);
buf BUF1 (N5639, N5603);
or OR4 (N5640, N5624, N2290, N651, N3615);
xor XOR2 (N5641, N5632, N2256);
nor NOR4 (N5642, N5609, N3784, N1462, N1529);
or OR2 (N5643, N5637, N377);
buf BUF1 (N5644, N5642);
and AND2 (N5645, N5636, N416);
nand NAND3 (N5646, N5635, N5458, N3800);
or OR3 (N5647, N5641, N4095, N1174);
nand NAND3 (N5648, N5647, N3427, N2191);
not NOT1 (N5649, N5631);
or OR3 (N5650, N5644, N3056, N21);
and AND4 (N5651, N5646, N170, N3947, N3003);
or OR4 (N5652, N5640, N2516, N3777, N3769);
and AND3 (N5653, N5651, N1721, N3885);
or OR3 (N5654, N5645, N4942, N3976);
buf BUF1 (N5655, N5639);
not NOT1 (N5656, N5652);
buf BUF1 (N5657, N5648);
and AND4 (N5658, N5650, N5275, N1428, N3930);
nor NOR4 (N5659, N5656, N808, N1818, N5486);
xor XOR2 (N5660, N5653, N2981);
buf BUF1 (N5661, N5658);
and AND2 (N5662, N5655, N443);
not NOT1 (N5663, N5657);
nand NAND3 (N5664, N5659, N2078, N5540);
buf BUF1 (N5665, N5643);
buf BUF1 (N5666, N5662);
xor XOR2 (N5667, N5654, N896);
nand NAND2 (N5668, N5666, N283);
not NOT1 (N5669, N5661);
nand NAND2 (N5670, N5667, N3103);
xor XOR2 (N5671, N5664, N802);
buf BUF1 (N5672, N5665);
buf BUF1 (N5673, N5671);
not NOT1 (N5674, N5672);
not NOT1 (N5675, N5649);
nand NAND4 (N5676, N5638, N368, N1166, N5132);
nand NAND3 (N5677, N5675, N2658, N3758);
or OR2 (N5678, N5677, N3155);
and AND4 (N5679, N5663, N2290, N5135, N4529);
nand NAND4 (N5680, N5628, N1416, N3562, N2655);
nor NOR4 (N5681, N5676, N1371, N1961, N255);
xor XOR2 (N5682, N5681, N3560);
and AND4 (N5683, N5680, N3230, N3144, N732);
buf BUF1 (N5684, N5669);
buf BUF1 (N5685, N5684);
nand NAND4 (N5686, N5682, N5268, N173, N1823);
buf BUF1 (N5687, N5674);
nor NOR4 (N5688, N5683, N7, N5054, N5278);
xor XOR2 (N5689, N5678, N5098);
or OR2 (N5690, N5689, N1707);
and AND4 (N5691, N5668, N2713, N5674, N4570);
nand NAND4 (N5692, N5688, N5361, N1853, N4513);
buf BUF1 (N5693, N5670);
xor XOR2 (N5694, N5690, N711);
and AND2 (N5695, N5685, N1281);
or OR3 (N5696, N5693, N3866, N1478);
and AND4 (N5697, N5692, N438, N651, N772);
and AND4 (N5698, N5679, N32, N49, N2057);
nand NAND3 (N5699, N5697, N4172, N5030);
and AND2 (N5700, N5699, N994);
nor NOR3 (N5701, N5687, N4870, N4814);
buf BUF1 (N5702, N5695);
not NOT1 (N5703, N5702);
not NOT1 (N5704, N5691);
xor XOR2 (N5705, N5686, N5298);
nor NOR2 (N5706, N5703, N2722);
buf BUF1 (N5707, N5673);
xor XOR2 (N5708, N5698, N4972);
or OR3 (N5709, N5700, N4279, N2479);
xor XOR2 (N5710, N5708, N2019);
and AND4 (N5711, N5710, N2001, N587, N1334);
and AND3 (N5712, N5706, N2878, N4975);
and AND4 (N5713, N5704, N43, N4739, N619);
not NOT1 (N5714, N5696);
xor XOR2 (N5715, N5660, N5511);
xor XOR2 (N5716, N5694, N1613);
nor NOR3 (N5717, N5709, N141, N5265);
nand NAND4 (N5718, N5712, N2243, N610, N4509);
not NOT1 (N5719, N5715);
not NOT1 (N5720, N5719);
nand NAND3 (N5721, N5717, N4681, N1437);
not NOT1 (N5722, N5701);
nor NOR3 (N5723, N5714, N2591, N4443);
and AND2 (N5724, N5707, N4762);
buf BUF1 (N5725, N5724);
nor NOR3 (N5726, N5713, N5701, N1722);
buf BUF1 (N5727, N5726);
nand NAND2 (N5728, N5725, N1409);
or OR2 (N5729, N5705, N1570);
nor NOR3 (N5730, N5729, N1971, N3721);
not NOT1 (N5731, N5718);
nor NOR3 (N5732, N5711, N3532, N4771);
nor NOR3 (N5733, N5728, N3818, N2396);
buf BUF1 (N5734, N5716);
nor NOR4 (N5735, N5722, N4235, N5396, N1377);
not NOT1 (N5736, N5721);
not NOT1 (N5737, N5735);
not NOT1 (N5738, N5732);
xor XOR2 (N5739, N5738, N567);
buf BUF1 (N5740, N5739);
buf BUF1 (N5741, N5720);
xor XOR2 (N5742, N5731, N3035);
nand NAND2 (N5743, N5733, N4545);
nand NAND2 (N5744, N5730, N4301);
or OR2 (N5745, N5727, N659);
or OR4 (N5746, N5741, N5715, N647, N1241);
nand NAND4 (N5747, N5737, N792, N4818, N3778);
and AND4 (N5748, N5743, N4666, N1034, N320);
nor NOR2 (N5749, N5744, N4898);
nor NOR3 (N5750, N5748, N987, N385);
and AND4 (N5751, N5734, N2561, N5190, N228);
nor NOR2 (N5752, N5749, N5663);
buf BUF1 (N5753, N5723);
or OR3 (N5754, N5740, N1088, N175);
or OR3 (N5755, N5750, N5219, N891);
buf BUF1 (N5756, N5751);
or OR4 (N5757, N5747, N3945, N103, N814);
not NOT1 (N5758, N5754);
xor XOR2 (N5759, N5742, N1494);
buf BUF1 (N5760, N5757);
not NOT1 (N5761, N5752);
and AND4 (N5762, N5736, N2597, N1931, N4950);
and AND2 (N5763, N5745, N5056);
not NOT1 (N5764, N5753);
buf BUF1 (N5765, N5758);
or OR4 (N5766, N5763, N3324, N803, N1209);
nand NAND4 (N5767, N5755, N2711, N4139, N1956);
xor XOR2 (N5768, N5756, N2027);
buf BUF1 (N5769, N5746);
or OR2 (N5770, N5766, N3238);
nor NOR2 (N5771, N5768, N1409);
nor NOR2 (N5772, N5762, N950);
and AND3 (N5773, N5770, N4317, N2056);
buf BUF1 (N5774, N5765);
or OR4 (N5775, N5769, N1038, N1914, N3225);
nor NOR4 (N5776, N5775, N5688, N2253, N1365);
buf BUF1 (N5777, N5760);
nand NAND3 (N5778, N5776, N2843, N2760);
xor XOR2 (N5779, N5773, N4177);
not NOT1 (N5780, N5779);
not NOT1 (N5781, N5764);
nor NOR4 (N5782, N5781, N4928, N4514, N610);
nor NOR4 (N5783, N5780, N1907, N5200, N3519);
nor NOR3 (N5784, N5783, N1816, N357);
not NOT1 (N5785, N5782);
nor NOR4 (N5786, N5784, N1033, N3258, N2525);
and AND3 (N5787, N5772, N5258, N4404);
buf BUF1 (N5788, N5774);
xor XOR2 (N5789, N5767, N5503);
xor XOR2 (N5790, N5786, N4156);
not NOT1 (N5791, N5777);
nor NOR4 (N5792, N5789, N2448, N5086, N3511);
and AND2 (N5793, N5788, N441);
xor XOR2 (N5794, N5792, N5251);
and AND2 (N5795, N5778, N4790);
nand NAND2 (N5796, N5790, N228);
not NOT1 (N5797, N5793);
nand NAND4 (N5798, N5771, N2025, N2164, N5634);
not NOT1 (N5799, N5796);
nand NAND4 (N5800, N5785, N1108, N3099, N760);
nand NAND2 (N5801, N5798, N4955);
buf BUF1 (N5802, N5795);
and AND2 (N5803, N5799, N3453);
buf BUF1 (N5804, N5802);
nor NOR3 (N5805, N5761, N2933, N4630);
nor NOR2 (N5806, N5803, N3767);
xor XOR2 (N5807, N5804, N1536);
nand NAND2 (N5808, N5800, N3848);
not NOT1 (N5809, N5794);
xor XOR2 (N5810, N5805, N5281);
not NOT1 (N5811, N5807);
nor NOR4 (N5812, N5809, N5793, N3287, N1008);
and AND3 (N5813, N5811, N420, N5450);
xor XOR2 (N5814, N5812, N4669);
or OR2 (N5815, N5814, N1653);
nor NOR3 (N5816, N5806, N5388, N3255);
or OR3 (N5817, N5810, N4204, N1229);
nand NAND3 (N5818, N5815, N586, N3608);
buf BUF1 (N5819, N5818);
buf BUF1 (N5820, N5787);
and AND4 (N5821, N5816, N4459, N1451, N1536);
and AND4 (N5822, N5801, N894, N1475, N421);
not NOT1 (N5823, N5797);
and AND4 (N5824, N5823, N5353, N1095, N2891);
buf BUF1 (N5825, N5820);
not NOT1 (N5826, N5791);
or OR2 (N5827, N5813, N5304);
and AND2 (N5828, N5817, N701);
xor XOR2 (N5829, N5822, N1194);
or OR3 (N5830, N5826, N1017, N1691);
and AND3 (N5831, N5830, N3946, N3898);
nor NOR4 (N5832, N5759, N621, N2416, N1103);
or OR4 (N5833, N5827, N2639, N1719, N1936);
not NOT1 (N5834, N5824);
nand NAND2 (N5835, N5829, N4813);
or OR4 (N5836, N5819, N4163, N4640, N1138);
buf BUF1 (N5837, N5834);
buf BUF1 (N5838, N5835);
xor XOR2 (N5839, N5831, N2879);
and AND2 (N5840, N5828, N1911);
and AND4 (N5841, N5839, N4339, N878, N2441);
xor XOR2 (N5842, N5840, N5071);
or OR2 (N5843, N5837, N3265);
xor XOR2 (N5844, N5808, N369);
nand NAND4 (N5845, N5843, N5079, N970, N1164);
buf BUF1 (N5846, N5842);
xor XOR2 (N5847, N5844, N321);
xor XOR2 (N5848, N5845, N4937);
or OR4 (N5849, N5841, N3075, N2640, N4751);
buf BUF1 (N5850, N5846);
xor XOR2 (N5851, N5849, N2271);
nand NAND4 (N5852, N5833, N2222, N3903, N1958);
or OR3 (N5853, N5825, N5209, N1366);
nand NAND4 (N5854, N5832, N2144, N3850, N440);
nand NAND2 (N5855, N5851, N5504);
xor XOR2 (N5856, N5821, N3566);
nor NOR4 (N5857, N5856, N2155, N3862, N876);
or OR3 (N5858, N5852, N3880, N130);
not NOT1 (N5859, N5848);
or OR3 (N5860, N5859, N5659, N3884);
xor XOR2 (N5861, N5850, N2178);
buf BUF1 (N5862, N5853);
nor NOR4 (N5863, N5860, N698, N2896, N1779);
nor NOR3 (N5864, N5858, N5185, N2040);
buf BUF1 (N5865, N5862);
xor XOR2 (N5866, N5865, N1501);
or OR2 (N5867, N5854, N2662);
and AND3 (N5868, N5864, N2132, N366);
buf BUF1 (N5869, N5847);
and AND2 (N5870, N5869, N3666);
nor NOR4 (N5871, N5838, N3450, N3862, N517);
not NOT1 (N5872, N5871);
not NOT1 (N5873, N5836);
nand NAND3 (N5874, N5861, N640, N2102);
not NOT1 (N5875, N5870);
buf BUF1 (N5876, N5868);
buf BUF1 (N5877, N5866);
nor NOR2 (N5878, N5877, N4964);
buf BUF1 (N5879, N5872);
buf BUF1 (N5880, N5875);
nor NOR4 (N5881, N5867, N3021, N5128, N3189);
not NOT1 (N5882, N5879);
buf BUF1 (N5883, N5873);
buf BUF1 (N5884, N5855);
xor XOR2 (N5885, N5878, N2052);
buf BUF1 (N5886, N5882);
not NOT1 (N5887, N5880);
nor NOR3 (N5888, N5876, N4897, N3814);
and AND2 (N5889, N5881, N660);
nand NAND4 (N5890, N5857, N5140, N5703, N5509);
and AND2 (N5891, N5890, N1803);
xor XOR2 (N5892, N5891, N3382);
or OR4 (N5893, N5889, N5814, N4849, N5453);
buf BUF1 (N5894, N5886);
nand NAND3 (N5895, N5874, N5452, N1743);
buf BUF1 (N5896, N5895);
nand NAND4 (N5897, N5885, N2564, N5687, N3340);
xor XOR2 (N5898, N5892, N4236);
nor NOR4 (N5899, N5893, N405, N4585, N4300);
nor NOR4 (N5900, N5899, N5723, N1770, N368);
nand NAND2 (N5901, N5900, N1141);
buf BUF1 (N5902, N5884);
xor XOR2 (N5903, N5902, N3973);
nand NAND2 (N5904, N5887, N18);
nor NOR3 (N5905, N5883, N5538, N1827);
buf BUF1 (N5906, N5863);
not NOT1 (N5907, N5894);
and AND4 (N5908, N5888, N3589, N837, N4453);
xor XOR2 (N5909, N5897, N3178);
buf BUF1 (N5910, N5898);
not NOT1 (N5911, N5901);
and AND3 (N5912, N5907, N3760, N2943);
or OR4 (N5913, N5896, N5834, N5653, N2499);
nor NOR2 (N5914, N5912, N2808);
not NOT1 (N5915, N5911);
nor NOR3 (N5916, N5909, N3873, N4755);
not NOT1 (N5917, N5906);
nand NAND4 (N5918, N5915, N546, N86, N4250);
and AND3 (N5919, N5903, N4039, N470);
and AND3 (N5920, N5919, N1574, N3599);
xor XOR2 (N5921, N5913, N3730);
not NOT1 (N5922, N5914);
xor XOR2 (N5923, N5916, N648);
nand NAND4 (N5924, N5908, N1351, N4195, N3675);
xor XOR2 (N5925, N5923, N4468);
nor NOR2 (N5926, N5925, N5915);
nand NAND4 (N5927, N5910, N2833, N3985, N4599);
not NOT1 (N5928, N5927);
nor NOR2 (N5929, N5904, N5775);
buf BUF1 (N5930, N5929);
buf BUF1 (N5931, N5905);
nand NAND2 (N5932, N5930, N3082);
nor NOR3 (N5933, N5922, N4880, N5126);
buf BUF1 (N5934, N5918);
nor NOR4 (N5935, N5917, N4825, N3817, N3655);
not NOT1 (N5936, N5935);
and AND3 (N5937, N5924, N2250, N4922);
nor NOR4 (N5938, N5926, N1968, N5191, N2079);
buf BUF1 (N5939, N5938);
not NOT1 (N5940, N5939);
and AND4 (N5941, N5933, N4242, N1502, N4663);
and AND2 (N5942, N5940, N4040);
and AND2 (N5943, N5937, N5528);
nand NAND4 (N5944, N5941, N5717, N3503, N861);
not NOT1 (N5945, N5931);
nand NAND4 (N5946, N5934, N5731, N1950, N4400);
and AND4 (N5947, N5943, N4963, N2014, N3314);
nand NAND3 (N5948, N5945, N868, N249);
not NOT1 (N5949, N5920);
not NOT1 (N5950, N5936);
and AND4 (N5951, N5932, N4691, N3681, N5259);
and AND2 (N5952, N5950, N3520);
nand NAND2 (N5953, N5928, N4807);
not NOT1 (N5954, N5949);
buf BUF1 (N5955, N5948);
xor XOR2 (N5956, N5921, N1222);
nand NAND3 (N5957, N5953, N707, N4949);
and AND2 (N5958, N5946, N744);
nand NAND3 (N5959, N5958, N4333, N3491);
not NOT1 (N5960, N5944);
not NOT1 (N5961, N5947);
buf BUF1 (N5962, N5955);
nand NAND4 (N5963, N5962, N3450, N4497, N4327);
and AND2 (N5964, N5959, N3625);
or OR4 (N5965, N5957, N620, N3299, N109);
nand NAND4 (N5966, N5960, N3876, N1460, N841);
not NOT1 (N5967, N5952);
xor XOR2 (N5968, N5965, N2906);
nor NOR4 (N5969, N5951, N4980, N3879, N5636);
or OR4 (N5970, N5969, N2168, N2546, N718);
xor XOR2 (N5971, N5963, N3751);
and AND2 (N5972, N5970, N247);
nor NOR4 (N5973, N5942, N3548, N5271, N5945);
buf BUF1 (N5974, N5964);
xor XOR2 (N5975, N5966, N4865);
nand NAND2 (N5976, N5968, N3447);
not NOT1 (N5977, N5976);
xor XOR2 (N5978, N5974, N3073);
not NOT1 (N5979, N5972);
nor NOR4 (N5980, N5973, N1403, N2226, N4397);
buf BUF1 (N5981, N5980);
nor NOR4 (N5982, N5954, N216, N3496, N4173);
nor NOR4 (N5983, N5975, N5420, N3936, N235);
and AND3 (N5984, N5961, N2979, N4818);
nor NOR4 (N5985, N5979, N1639, N1031, N2322);
buf BUF1 (N5986, N5971);
xor XOR2 (N5987, N5977, N2974);
nand NAND3 (N5988, N5983, N3955, N4782);
buf BUF1 (N5989, N5981);
nand NAND4 (N5990, N5986, N541, N2529, N2394);
xor XOR2 (N5991, N5978, N3582);
and AND4 (N5992, N5984, N41, N244, N1210);
or OR4 (N5993, N5985, N5659, N3320, N169);
xor XOR2 (N5994, N5993, N1009);
xor XOR2 (N5995, N5991, N2939);
xor XOR2 (N5996, N5994, N3284);
not NOT1 (N5997, N5987);
buf BUF1 (N5998, N5995);
xor XOR2 (N5999, N5988, N4305);
buf BUF1 (N6000, N5982);
nor NOR4 (N6001, N6000, N3417, N2118, N757);
xor XOR2 (N6002, N5997, N4045);
not NOT1 (N6003, N5967);
or OR4 (N6004, N5956, N4613, N4517, N2301);
nor NOR4 (N6005, N6004, N2793, N2149, N230);
buf BUF1 (N6006, N6001);
nand NAND4 (N6007, N6005, N2299, N2960, N202);
buf BUF1 (N6008, N5990);
not NOT1 (N6009, N5989);
and AND2 (N6010, N6008, N1018);
nand NAND2 (N6011, N5998, N5143);
xor XOR2 (N6012, N6002, N1443);
or OR3 (N6013, N6007, N1309, N5484);
buf BUF1 (N6014, N6003);
not NOT1 (N6015, N6011);
not NOT1 (N6016, N6009);
xor XOR2 (N6017, N5992, N4528);
or OR3 (N6018, N5996, N2917, N1921);
or OR2 (N6019, N6016, N3958);
nand NAND2 (N6020, N6015, N4476);
not NOT1 (N6021, N6010);
nor NOR3 (N6022, N6006, N2430, N1458);
or OR4 (N6023, N6019, N5371, N4336, N2358);
xor XOR2 (N6024, N5999, N1510);
and AND3 (N6025, N6017, N2433, N3672);
or OR4 (N6026, N6020, N5081, N126, N1166);
buf BUF1 (N6027, N6014);
or OR4 (N6028, N6024, N210, N4483, N5774);
nor NOR3 (N6029, N6013, N3441, N1834);
nor NOR2 (N6030, N6026, N4679);
or OR3 (N6031, N6022, N5241, N6002);
not NOT1 (N6032, N6028);
buf BUF1 (N6033, N6012);
buf BUF1 (N6034, N6030);
not NOT1 (N6035, N6031);
or OR3 (N6036, N6032, N331, N537);
xor XOR2 (N6037, N6035, N2324);
xor XOR2 (N6038, N6034, N5513);
xor XOR2 (N6039, N6033, N4022);
not NOT1 (N6040, N6029);
xor XOR2 (N6041, N6027, N618);
nand NAND4 (N6042, N6023, N1184, N5181, N3252);
buf BUF1 (N6043, N6042);
or OR3 (N6044, N6041, N3313, N2027);
and AND3 (N6045, N6038, N69, N3827);
buf BUF1 (N6046, N6045);
and AND3 (N6047, N6046, N373, N4282);
or OR4 (N6048, N6021, N582, N927, N4672);
nand NAND3 (N6049, N6048, N1209, N1688);
buf BUF1 (N6050, N6049);
and AND2 (N6051, N6040, N5765);
or OR3 (N6052, N6037, N1465, N4853);
nand NAND2 (N6053, N6036, N2201);
not NOT1 (N6054, N6052);
not NOT1 (N6055, N6039);
and AND2 (N6056, N6047, N5178);
nand NAND4 (N6057, N6054, N2667, N2937, N2415);
buf BUF1 (N6058, N6018);
buf BUF1 (N6059, N6050);
or OR3 (N6060, N6043, N3491, N1194);
buf BUF1 (N6061, N6044);
buf BUF1 (N6062, N6061);
buf BUF1 (N6063, N6059);
and AND3 (N6064, N6056, N910, N5208);
and AND3 (N6065, N6060, N1592, N974);
xor XOR2 (N6066, N6062, N4900);
buf BUF1 (N6067, N6066);
nor NOR2 (N6068, N6065, N5897);
not NOT1 (N6069, N6057);
buf BUF1 (N6070, N6067);
buf BUF1 (N6071, N6069);
nor NOR2 (N6072, N6071, N3798);
and AND2 (N6073, N6063, N537);
not NOT1 (N6074, N6051);
buf BUF1 (N6075, N6074);
nor NOR4 (N6076, N6075, N5507, N925, N5797);
nor NOR2 (N6077, N6068, N295);
buf BUF1 (N6078, N6073);
nand NAND3 (N6079, N6053, N4468, N743);
nor NOR4 (N6080, N6070, N4377, N4508, N4677);
or OR3 (N6081, N6077, N3700, N1518);
nor NOR2 (N6082, N6064, N4824);
not NOT1 (N6083, N6058);
and AND2 (N6084, N6025, N1356);
not NOT1 (N6085, N6076);
xor XOR2 (N6086, N6084, N4401);
xor XOR2 (N6087, N6082, N5622);
nor NOR2 (N6088, N6079, N2471);
buf BUF1 (N6089, N6078);
nor NOR2 (N6090, N6085, N1077);
nor NOR4 (N6091, N6083, N3345, N3121, N4876);
nor NOR3 (N6092, N6055, N1620, N1654);
xor XOR2 (N6093, N6080, N5003);
xor XOR2 (N6094, N6087, N103);
nor NOR4 (N6095, N6088, N4350, N2996, N3889);
not NOT1 (N6096, N6089);
not NOT1 (N6097, N6096);
xor XOR2 (N6098, N6091, N2068);
nand NAND4 (N6099, N6093, N1037, N1650, N3283);
and AND2 (N6100, N6099, N6028);
buf BUF1 (N6101, N6100);
nor NOR2 (N6102, N6086, N603);
not NOT1 (N6103, N6097);
nand NAND4 (N6104, N6090, N4221, N1928, N5101);
not NOT1 (N6105, N6072);
nand NAND2 (N6106, N6095, N3010);
or OR4 (N6107, N6081, N1865, N1584, N3950);
or OR2 (N6108, N6104, N3340);
nand NAND4 (N6109, N6107, N4718, N826, N5331);
or OR2 (N6110, N6101, N3955);
nand NAND4 (N6111, N6105, N4288, N1654, N3130);
xor XOR2 (N6112, N6094, N5316);
nor NOR3 (N6113, N6102, N2621, N5094);
nor NOR4 (N6114, N6110, N1372, N5910, N2687);
xor XOR2 (N6115, N6109, N3518);
buf BUF1 (N6116, N6098);
and AND3 (N6117, N6106, N2221, N6003);
not NOT1 (N6118, N6117);
or OR3 (N6119, N6112, N3477, N5365);
and AND2 (N6120, N6116, N3773);
not NOT1 (N6121, N6092);
not NOT1 (N6122, N6115);
buf BUF1 (N6123, N6121);
not NOT1 (N6124, N6122);
buf BUF1 (N6125, N6108);
nand NAND3 (N6126, N6111, N1057, N2242);
nand NAND4 (N6127, N6114, N5794, N1139, N1284);
or OR4 (N6128, N6125, N4588, N2348, N4958);
xor XOR2 (N6129, N6118, N427);
buf BUF1 (N6130, N6128);
nor NOR2 (N6131, N6124, N1518);
not NOT1 (N6132, N6119);
buf BUF1 (N6133, N6113);
xor XOR2 (N6134, N6130, N2937);
not NOT1 (N6135, N6123);
nand NAND2 (N6136, N6129, N3158);
buf BUF1 (N6137, N6133);
and AND3 (N6138, N6131, N6023, N3724);
xor XOR2 (N6139, N6126, N4065);
buf BUF1 (N6140, N6136);
buf BUF1 (N6141, N6140);
nand NAND4 (N6142, N6103, N1948, N3310, N183);
nor NOR2 (N6143, N6142, N3247);
nor NOR4 (N6144, N6139, N525, N4176, N5464);
xor XOR2 (N6145, N6134, N853);
and AND2 (N6146, N6137, N157);
not NOT1 (N6147, N6146);
not NOT1 (N6148, N6145);
and AND2 (N6149, N6132, N2864);
buf BUF1 (N6150, N6143);
buf BUF1 (N6151, N6149);
or OR2 (N6152, N6120, N3125);
or OR2 (N6153, N6151, N1150);
or OR2 (N6154, N6135, N4107);
nor NOR2 (N6155, N6138, N3063);
nand NAND3 (N6156, N6147, N5280, N4516);
or OR4 (N6157, N6144, N2539, N2444, N4025);
and AND2 (N6158, N6152, N3262);
nor NOR3 (N6159, N6157, N6095, N1876);
buf BUF1 (N6160, N6159);
nor NOR3 (N6161, N6148, N4204, N289);
xor XOR2 (N6162, N6160, N2018);
and AND3 (N6163, N6154, N5721, N5930);
buf BUF1 (N6164, N6161);
nor NOR2 (N6165, N6141, N5483);
nor NOR2 (N6166, N6164, N2656);
or OR3 (N6167, N6163, N5393, N1021);
or OR3 (N6168, N6165, N5445, N1111);
and AND3 (N6169, N6127, N2560, N697);
buf BUF1 (N6170, N6162);
not NOT1 (N6171, N6169);
buf BUF1 (N6172, N6170);
and AND2 (N6173, N6167, N5569);
nor NOR4 (N6174, N6168, N3482, N3386, N3417);
not NOT1 (N6175, N6155);
xor XOR2 (N6176, N6173, N5477);
xor XOR2 (N6177, N6175, N1274);
xor XOR2 (N6178, N6177, N3840);
nand NAND4 (N6179, N6158, N3161, N482, N5703);
xor XOR2 (N6180, N6179, N614);
nor NOR4 (N6181, N6153, N303, N597, N1750);
not NOT1 (N6182, N6166);
or OR3 (N6183, N6174, N2031, N5818);
and AND3 (N6184, N6172, N4067, N1126);
buf BUF1 (N6185, N6183);
and AND4 (N6186, N6184, N2608, N2885, N3210);
nor NOR3 (N6187, N6181, N431, N4903);
nor NOR3 (N6188, N6186, N765, N1618);
nand NAND2 (N6189, N6178, N2970);
nor NOR3 (N6190, N6171, N5693, N1786);
or OR2 (N6191, N6188, N3825);
nor NOR3 (N6192, N6176, N4610, N5164);
and AND3 (N6193, N6189, N3306, N5261);
not NOT1 (N6194, N6191);
xor XOR2 (N6195, N6150, N3932);
xor XOR2 (N6196, N6182, N867);
not NOT1 (N6197, N6187);
buf BUF1 (N6198, N6156);
not NOT1 (N6199, N6190);
and AND3 (N6200, N6196, N4910, N3982);
buf BUF1 (N6201, N6199);
nor NOR3 (N6202, N6185, N4887, N2240);
and AND2 (N6203, N6200, N5553);
not NOT1 (N6204, N6197);
buf BUF1 (N6205, N6193);
not NOT1 (N6206, N6205);
nor NOR2 (N6207, N6194, N6009);
xor XOR2 (N6208, N6201, N802);
buf BUF1 (N6209, N6207);
or OR2 (N6210, N6198, N143);
nor NOR2 (N6211, N6208, N1604);
buf BUF1 (N6212, N6206);
not NOT1 (N6213, N6211);
not NOT1 (N6214, N6195);
nand NAND4 (N6215, N6204, N5375, N355, N3711);
nor NOR2 (N6216, N6215, N2307);
xor XOR2 (N6217, N6192, N4445);
xor XOR2 (N6218, N6209, N4549);
buf BUF1 (N6219, N6214);
or OR2 (N6220, N6210, N1253);
and AND2 (N6221, N6180, N156);
nand NAND4 (N6222, N6203, N2880, N1826, N4490);
and AND4 (N6223, N6217, N1314, N1186, N5993);
not NOT1 (N6224, N6218);
and AND3 (N6225, N6219, N5750, N3895);
or OR3 (N6226, N6223, N2787, N1183);
nor NOR2 (N6227, N6221, N2152);
buf BUF1 (N6228, N6212);
or OR4 (N6229, N6227, N1801, N3088, N847);
not NOT1 (N6230, N6216);
xor XOR2 (N6231, N6225, N2238);
and AND4 (N6232, N6229, N5700, N1284, N5103);
or OR3 (N6233, N6232, N5341, N1953);
nor NOR4 (N6234, N6202, N4750, N3985, N3845);
and AND4 (N6235, N6213, N2983, N5792, N2521);
and AND4 (N6236, N6231, N558, N4946, N1710);
and AND2 (N6237, N6235, N2571);
not NOT1 (N6238, N6226);
and AND4 (N6239, N6224, N1228, N4734, N4270);
and AND4 (N6240, N6220, N3045, N2967, N2300);
and AND2 (N6241, N6233, N4158);
xor XOR2 (N6242, N6240, N960);
nor NOR3 (N6243, N6234, N3798, N1362);
nor NOR4 (N6244, N6230, N3723, N4382, N582);
and AND3 (N6245, N6243, N5183, N2936);
or OR3 (N6246, N6245, N3523, N2470);
not NOT1 (N6247, N6239);
buf BUF1 (N6248, N6246);
nand NAND2 (N6249, N6236, N6164);
nand NAND2 (N6250, N6249, N5130);
nand NAND4 (N6251, N6228, N4732, N2639, N1034);
nor NOR4 (N6252, N6222, N5771, N3520, N3053);
or OR4 (N6253, N6247, N2415, N3419, N897);
and AND3 (N6254, N6242, N1534, N6211);
nand NAND3 (N6255, N6244, N1772, N5941);
and AND4 (N6256, N6253, N1182, N609, N1508);
buf BUF1 (N6257, N6255);
and AND4 (N6258, N6257, N243, N1486, N5985);
xor XOR2 (N6259, N6256, N4499);
buf BUF1 (N6260, N6238);
not NOT1 (N6261, N6241);
not NOT1 (N6262, N6261);
nand NAND4 (N6263, N6252, N737, N1561, N5230);
nand NAND3 (N6264, N6251, N2876, N3940);
buf BUF1 (N6265, N6254);
and AND4 (N6266, N6262, N2906, N4323, N5837);
nor NOR4 (N6267, N6263, N5742, N1807, N4287);
nand NAND4 (N6268, N6264, N1734, N5269, N5439);
or OR4 (N6269, N6248, N4255, N5510, N5121);
not NOT1 (N6270, N6268);
xor XOR2 (N6271, N6270, N3040);
not NOT1 (N6272, N6267);
xor XOR2 (N6273, N6259, N2105);
or OR3 (N6274, N6272, N607, N4422);
buf BUF1 (N6275, N6266);
not NOT1 (N6276, N6265);
not NOT1 (N6277, N6273);
and AND2 (N6278, N6276, N4563);
not NOT1 (N6279, N6271);
nor NOR4 (N6280, N6260, N4704, N4940, N4164);
and AND3 (N6281, N6280, N4384, N4893);
nand NAND4 (N6282, N6258, N4959, N3379, N1851);
buf BUF1 (N6283, N6250);
not NOT1 (N6284, N6282);
xor XOR2 (N6285, N6283, N1968);
or OR4 (N6286, N6269, N3939, N4824, N1501);
nor NOR3 (N6287, N6278, N1864, N6109);
and AND3 (N6288, N6284, N2514, N5270);
xor XOR2 (N6289, N6279, N3676);
nor NOR3 (N6290, N6277, N1542, N6030);
buf BUF1 (N6291, N6286);
nor NOR4 (N6292, N6285, N3201, N587, N3330);
or OR4 (N6293, N6237, N2075, N2506, N2936);
buf BUF1 (N6294, N6288);
xor XOR2 (N6295, N6281, N2573);
not NOT1 (N6296, N6294);
not NOT1 (N6297, N6293);
not NOT1 (N6298, N6275);
nand NAND4 (N6299, N6296, N5109, N2115, N1845);
or OR3 (N6300, N6297, N1127, N3909);
and AND2 (N6301, N6300, N5356);
buf BUF1 (N6302, N6299);
or OR3 (N6303, N6298, N1157, N2131);
buf BUF1 (N6304, N6289);
nor NOR2 (N6305, N6292, N4893);
not NOT1 (N6306, N6304);
nor NOR2 (N6307, N6287, N3478);
or OR3 (N6308, N6274, N4298, N2205);
xor XOR2 (N6309, N6301, N2789);
or OR4 (N6310, N6291, N3840, N2166, N2117);
not NOT1 (N6311, N6306);
nand NAND4 (N6312, N6295, N5579, N4398, N1139);
not NOT1 (N6313, N6305);
nand NAND3 (N6314, N6312, N4967, N5030);
nor NOR3 (N6315, N6302, N2700, N495);
nor NOR2 (N6316, N6290, N5606);
not NOT1 (N6317, N6307);
nand NAND3 (N6318, N6314, N5319, N452);
nor NOR4 (N6319, N6308, N4033, N5945, N794);
and AND3 (N6320, N6313, N3538, N3018);
or OR4 (N6321, N6310, N1954, N140, N5487);
buf BUF1 (N6322, N6311);
xor XOR2 (N6323, N6316, N4425);
buf BUF1 (N6324, N6319);
or OR3 (N6325, N6320, N3902, N4205);
or OR4 (N6326, N6317, N226, N1799, N5395);
nand NAND3 (N6327, N6309, N2430, N708);
not NOT1 (N6328, N6318);
nand NAND4 (N6329, N6323, N3526, N6023, N4036);
or OR2 (N6330, N6315, N2271);
nand NAND3 (N6331, N6324, N2687, N3868);
xor XOR2 (N6332, N6325, N3251);
and AND3 (N6333, N6322, N6054, N3433);
not NOT1 (N6334, N6329);
not NOT1 (N6335, N6326);
nand NAND3 (N6336, N6334, N2274, N658);
not NOT1 (N6337, N6332);
or OR4 (N6338, N6321, N3188, N4844, N268);
buf BUF1 (N6339, N6330);
not NOT1 (N6340, N6335);
buf BUF1 (N6341, N6328);
nand NAND2 (N6342, N6327, N942);
not NOT1 (N6343, N6342);
or OR2 (N6344, N6331, N5805);
buf BUF1 (N6345, N6333);
not NOT1 (N6346, N6340);
nor NOR4 (N6347, N6344, N2493, N6097, N5334);
nor NOR2 (N6348, N6346, N2645);
nor NOR4 (N6349, N6347, N4063, N3598, N1943);
nor NOR2 (N6350, N6345, N1632);
nor NOR2 (N6351, N6348, N4079);
nand NAND2 (N6352, N6303, N482);
not NOT1 (N6353, N6343);
or OR4 (N6354, N6341, N4053, N5056, N2265);
xor XOR2 (N6355, N6350, N726);
not NOT1 (N6356, N6349);
xor XOR2 (N6357, N6351, N5875);
nand NAND4 (N6358, N6357, N5027, N3617, N3758);
xor XOR2 (N6359, N6339, N270);
or OR2 (N6360, N6337, N3328);
or OR4 (N6361, N6355, N459, N1327, N443);
and AND4 (N6362, N6360, N2349, N816, N3622);
nand NAND4 (N6363, N6336, N6046, N4076, N174);
nand NAND4 (N6364, N6362, N3226, N3854, N6102);
nor NOR2 (N6365, N6338, N6029);
and AND4 (N6366, N6359, N2926, N749, N1231);
not NOT1 (N6367, N6364);
nand NAND2 (N6368, N6358, N4087);
nor NOR3 (N6369, N6366, N3402, N2407);
and AND4 (N6370, N6368, N945, N1855, N2940);
buf BUF1 (N6371, N6354);
nand NAND2 (N6372, N6371, N1686);
buf BUF1 (N6373, N6363);
not NOT1 (N6374, N6369);
and AND2 (N6375, N6373, N3425);
and AND2 (N6376, N6370, N3389);
nand NAND2 (N6377, N6353, N5629);
nor NOR4 (N6378, N6372, N2624, N5604, N836);
or OR4 (N6379, N6375, N6197, N2286, N3392);
or OR2 (N6380, N6377, N4572);
nand NAND4 (N6381, N6361, N1082, N4121, N71);
not NOT1 (N6382, N6376);
or OR4 (N6383, N6382, N4255, N4518, N1790);
xor XOR2 (N6384, N6378, N5734);
buf BUF1 (N6385, N6380);
xor XOR2 (N6386, N6367, N3363);
buf BUF1 (N6387, N6386);
and AND4 (N6388, N6365, N228, N4086, N2553);
xor XOR2 (N6389, N6374, N4366);
or OR2 (N6390, N6356, N5368);
buf BUF1 (N6391, N6389);
nor NOR4 (N6392, N6387, N5707, N5173, N577);
not NOT1 (N6393, N6392);
or OR3 (N6394, N6384, N5868, N1925);
buf BUF1 (N6395, N6393);
nand NAND2 (N6396, N6390, N1061);
not NOT1 (N6397, N6395);
and AND2 (N6398, N6352, N395);
or OR3 (N6399, N6396, N5386, N2871);
or OR3 (N6400, N6399, N4426, N5467);
not NOT1 (N6401, N6388);
nor NOR2 (N6402, N6398, N2212);
buf BUF1 (N6403, N6383);
nand NAND2 (N6404, N6397, N4195);
buf BUF1 (N6405, N6379);
or OR2 (N6406, N6401, N630);
or OR4 (N6407, N6403, N100, N360, N4334);
buf BUF1 (N6408, N6404);
or OR3 (N6409, N6406, N19, N1044);
nor NOR3 (N6410, N6405, N3151, N1745);
and AND3 (N6411, N6385, N838, N809);
not NOT1 (N6412, N6411);
nand NAND3 (N6413, N6400, N106, N5101);
and AND3 (N6414, N6394, N521, N3392);
and AND3 (N6415, N6407, N948, N4924);
or OR4 (N6416, N6402, N2357, N29, N5533);
or OR3 (N6417, N6410, N1297, N413);
xor XOR2 (N6418, N6413, N981);
nor NOR2 (N6419, N6408, N1826);
nor NOR3 (N6420, N6417, N540, N2420);
and AND3 (N6421, N6391, N233, N3002);
nand NAND4 (N6422, N6421, N4240, N2192, N6092);
and AND2 (N6423, N6414, N2522);
nand NAND4 (N6424, N6420, N1877, N2639, N5388);
or OR2 (N6425, N6418, N2817);
and AND4 (N6426, N6425, N350, N3621, N4922);
xor XOR2 (N6427, N6419, N3535);
buf BUF1 (N6428, N6416);
nand NAND4 (N6429, N6422, N4819, N3915, N4163);
xor XOR2 (N6430, N6426, N1648);
nor NOR2 (N6431, N6381, N2749);
not NOT1 (N6432, N6430);
xor XOR2 (N6433, N6424, N2906);
buf BUF1 (N6434, N6429);
and AND2 (N6435, N6423, N5282);
not NOT1 (N6436, N6434);
nand NAND4 (N6437, N6409, N113, N722, N3069);
nor NOR2 (N6438, N6436, N5186);
nand NAND2 (N6439, N6432, N6022);
nand NAND2 (N6440, N6427, N3489);
and AND4 (N6441, N6431, N1670, N310, N3249);
nor NOR2 (N6442, N6439, N1598);
or OR2 (N6443, N6415, N2354);
nor NOR4 (N6444, N6440, N158, N5292, N6227);
or OR3 (N6445, N6438, N1841, N4610);
xor XOR2 (N6446, N6442, N4839);
nand NAND3 (N6447, N6435, N119, N6014);
and AND2 (N6448, N6412, N3678);
buf BUF1 (N6449, N6437);
xor XOR2 (N6450, N6428, N766);
and AND2 (N6451, N6448, N4171);
or OR3 (N6452, N6450, N2391, N6009);
or OR3 (N6453, N6445, N2475, N5793);
and AND3 (N6454, N6449, N1581, N3953);
buf BUF1 (N6455, N6441);
nand NAND2 (N6456, N6451, N974);
and AND2 (N6457, N6444, N4978);
not NOT1 (N6458, N6452);
or OR4 (N6459, N6455, N787, N3750, N4881);
nand NAND3 (N6460, N6457, N4290, N2810);
or OR4 (N6461, N6460, N4366, N2864, N5796);
or OR3 (N6462, N6433, N4875, N1637);
or OR2 (N6463, N6447, N1394);
xor XOR2 (N6464, N6461, N2662);
and AND2 (N6465, N6463, N4325);
nor NOR4 (N6466, N6446, N2610, N2216, N2765);
buf BUF1 (N6467, N6462);
nand NAND2 (N6468, N6458, N333);
or OR3 (N6469, N6468, N5066, N3576);
and AND3 (N6470, N6456, N3927, N3076);
nand NAND2 (N6471, N6469, N2906);
buf BUF1 (N6472, N6465);
buf BUF1 (N6473, N6472);
and AND3 (N6474, N6470, N2571, N3241);
nand NAND3 (N6475, N6459, N1493, N2877);
nand NAND4 (N6476, N6473, N608, N2991, N644);
not NOT1 (N6477, N6443);
nand NAND4 (N6478, N6476, N4936, N3882, N825);
not NOT1 (N6479, N6471);
nor NOR3 (N6480, N6475, N105, N575);
or OR3 (N6481, N6477, N1743, N1505);
not NOT1 (N6482, N6453);
buf BUF1 (N6483, N6481);
or OR2 (N6484, N6454, N3619);
xor XOR2 (N6485, N6464, N5371);
not NOT1 (N6486, N6479);
or OR4 (N6487, N6484, N238, N5795, N735);
xor XOR2 (N6488, N6486, N5903);
not NOT1 (N6489, N6488);
and AND4 (N6490, N6474, N4332, N954, N3430);
buf BUF1 (N6491, N6487);
nor NOR4 (N6492, N6489, N814, N1549, N4934);
xor XOR2 (N6493, N6478, N2504);
nand NAND3 (N6494, N6493, N6468, N2706);
xor XOR2 (N6495, N6480, N1791);
nor NOR2 (N6496, N6485, N1407);
not NOT1 (N6497, N6467);
nor NOR3 (N6498, N6490, N4670, N2297);
or OR4 (N6499, N6495, N4888, N1873, N3159);
buf BUF1 (N6500, N6496);
xor XOR2 (N6501, N6494, N1639);
and AND3 (N6502, N6501, N5098, N4774);
and AND4 (N6503, N6482, N4900, N2187, N1955);
nand NAND2 (N6504, N6491, N5144);
xor XOR2 (N6505, N6492, N1786);
nand NAND3 (N6506, N6504, N475, N1142);
or OR3 (N6507, N6505, N4822, N4349);
nor NOR4 (N6508, N6499, N331, N5278, N4246);
nor NOR4 (N6509, N6498, N4102, N5723, N1437);
buf BUF1 (N6510, N6506);
or OR4 (N6511, N6497, N5829, N1730, N6251);
xor XOR2 (N6512, N6503, N1926);
not NOT1 (N6513, N6509);
or OR2 (N6514, N6502, N3916);
and AND3 (N6515, N6514, N2831, N4200);
or OR3 (N6516, N6510, N6102, N1773);
nor NOR2 (N6517, N6511, N6285);
and AND4 (N6518, N6508, N4267, N683, N4208);
not NOT1 (N6519, N6516);
buf BUF1 (N6520, N6500);
not NOT1 (N6521, N6513);
nand NAND3 (N6522, N6521, N1850, N3996);
buf BUF1 (N6523, N6515);
or OR4 (N6524, N6518, N3317, N3914, N907);
xor XOR2 (N6525, N6512, N1258);
and AND3 (N6526, N6525, N1759, N4488);
and AND2 (N6527, N6507, N5824);
not NOT1 (N6528, N6523);
or OR3 (N6529, N6517, N1982, N2052);
and AND3 (N6530, N6483, N1907, N2048);
or OR2 (N6531, N6519, N4364);
xor XOR2 (N6532, N6530, N3076);
and AND3 (N6533, N6532, N3433, N4891);
or OR4 (N6534, N6531, N4300, N2225, N3337);
nand NAND3 (N6535, N6466, N3801, N55);
or OR2 (N6536, N6533, N5888);
not NOT1 (N6537, N6522);
buf BUF1 (N6538, N6537);
nor NOR2 (N6539, N6520, N312);
and AND2 (N6540, N6528, N927);
nand NAND3 (N6541, N6538, N4523, N2715);
or OR4 (N6542, N6534, N1544, N5098, N4976);
xor XOR2 (N6543, N6524, N1329);
not NOT1 (N6544, N6541);
or OR3 (N6545, N6543, N6178, N5452);
buf BUF1 (N6546, N6542);
nor NOR4 (N6547, N6540, N822, N4143, N5241);
and AND2 (N6548, N6539, N322);
nor NOR2 (N6549, N6536, N4030);
not NOT1 (N6550, N6535);
nand NAND2 (N6551, N6526, N386);
nor NOR4 (N6552, N6545, N1304, N1066, N4334);
nor NOR4 (N6553, N6551, N1452, N2364, N1755);
nand NAND4 (N6554, N6529, N4293, N3218, N5910);
or OR2 (N6555, N6554, N6500);
buf BUF1 (N6556, N6555);
buf BUF1 (N6557, N6547);
and AND2 (N6558, N6552, N917);
and AND2 (N6559, N6557, N2421);
nor NOR4 (N6560, N6556, N5935, N5259, N766);
not NOT1 (N6561, N6548);
nor NOR2 (N6562, N6561, N603);
xor XOR2 (N6563, N6553, N4795);
xor XOR2 (N6564, N6563, N1752);
nand NAND3 (N6565, N6549, N93, N4397);
xor XOR2 (N6566, N6544, N2329);
nor NOR3 (N6567, N6566, N3408, N3873);
and AND4 (N6568, N6562, N2618, N4390, N4095);
and AND3 (N6569, N6565, N2493, N3887);
buf BUF1 (N6570, N6559);
nor NOR3 (N6571, N6564, N5986, N3083);
nand NAND3 (N6572, N6570, N337, N1836);
or OR2 (N6573, N6572, N5699);
or OR2 (N6574, N6550, N2355);
or OR2 (N6575, N6568, N2696);
nor NOR3 (N6576, N6560, N3285, N1909);
or OR3 (N6577, N6527, N1674, N2563);
not NOT1 (N6578, N6571);
buf BUF1 (N6579, N6574);
nor NOR3 (N6580, N6546, N6117, N5210);
and AND4 (N6581, N6558, N160, N93, N2047);
and AND4 (N6582, N6569, N869, N5337, N6095);
buf BUF1 (N6583, N6580);
and AND3 (N6584, N6576, N6092, N4720);
nand NAND2 (N6585, N6575, N3623);
and AND2 (N6586, N6573, N3191);
not NOT1 (N6587, N6581);
not NOT1 (N6588, N6577);
nand NAND4 (N6589, N6586, N3446, N1138, N1912);
not NOT1 (N6590, N6588);
nand NAND4 (N6591, N6579, N4120, N6293, N1676);
xor XOR2 (N6592, N6590, N4583);
nor NOR4 (N6593, N6584, N2977, N397, N3602);
nor NOR4 (N6594, N6582, N4792, N536, N1733);
or OR3 (N6595, N6594, N2858, N5381);
not NOT1 (N6596, N6567);
nand NAND2 (N6597, N6585, N1287);
or OR2 (N6598, N6578, N3817);
xor XOR2 (N6599, N6598, N1356);
nor NOR3 (N6600, N6583, N2284, N4007);
buf BUF1 (N6601, N6596);
nand NAND3 (N6602, N6601, N1973, N2595);
or OR2 (N6603, N6587, N775);
nor NOR3 (N6604, N6602, N5879, N403);
buf BUF1 (N6605, N6597);
xor XOR2 (N6606, N6591, N825);
buf BUF1 (N6607, N6606);
xor XOR2 (N6608, N6593, N5401);
not NOT1 (N6609, N6589);
nor NOR2 (N6610, N6599, N4740);
or OR2 (N6611, N6592, N3254);
and AND4 (N6612, N6611, N124, N5070, N1871);
buf BUF1 (N6613, N6609);
buf BUF1 (N6614, N6600);
or OR4 (N6615, N6613, N4174, N655, N3264);
nor NOR4 (N6616, N6608, N2541, N901, N5980);
nand NAND3 (N6617, N6612, N2564, N521);
and AND4 (N6618, N6617, N1672, N1235, N2361);
not NOT1 (N6619, N6616);
not NOT1 (N6620, N6607);
buf BUF1 (N6621, N6603);
and AND4 (N6622, N6605, N3028, N4360, N539);
or OR3 (N6623, N6614, N2034, N1106);
xor XOR2 (N6624, N6621, N1377);
and AND4 (N6625, N6620, N5013, N4167, N4070);
buf BUF1 (N6626, N6604);
or OR4 (N6627, N6619, N5953, N4085, N4468);
not NOT1 (N6628, N6626);
and AND2 (N6629, N6610, N6020);
buf BUF1 (N6630, N6595);
nor NOR4 (N6631, N6622, N3512, N3419, N5809);
nand NAND4 (N6632, N6625, N1649, N1707, N6601);
not NOT1 (N6633, N6631);
not NOT1 (N6634, N6615);
and AND4 (N6635, N6618, N3784, N2319, N5609);
buf BUF1 (N6636, N6630);
nor NOR2 (N6637, N6627, N1211);
buf BUF1 (N6638, N6633);
nand NAND2 (N6639, N6634, N4646);
nor NOR3 (N6640, N6636, N6123, N5163);
nor NOR3 (N6641, N6637, N1423, N5720);
buf BUF1 (N6642, N6640);
xor XOR2 (N6643, N6632, N3126);
buf BUF1 (N6644, N6624);
nand NAND3 (N6645, N6642, N3760, N6029);
xor XOR2 (N6646, N6645, N61);
or OR4 (N6647, N6646, N4467, N2845, N489);
buf BUF1 (N6648, N6635);
and AND3 (N6649, N6641, N6559, N1410);
nand NAND2 (N6650, N6639, N4269);
xor XOR2 (N6651, N6647, N3797);
xor XOR2 (N6652, N6628, N3841);
or OR2 (N6653, N6649, N668);
nand NAND3 (N6654, N6623, N2635, N6528);
not NOT1 (N6655, N6643);
xor XOR2 (N6656, N6638, N4916);
xor XOR2 (N6657, N6629, N3278);
not NOT1 (N6658, N6657);
nor NOR3 (N6659, N6655, N4140, N4216);
nor NOR4 (N6660, N6654, N4975, N1118, N1674);
and AND4 (N6661, N6648, N3273, N5459, N6458);
buf BUF1 (N6662, N6651);
buf BUF1 (N6663, N6658);
nand NAND3 (N6664, N6653, N4715, N2291);
and AND2 (N6665, N6664, N5901);
nand NAND4 (N6666, N6652, N3645, N554, N2497);
buf BUF1 (N6667, N6663);
and AND2 (N6668, N6650, N1136);
and AND3 (N6669, N6662, N6086, N1312);
and AND2 (N6670, N6660, N1297);
or OR2 (N6671, N6670, N2565);
buf BUF1 (N6672, N6656);
xor XOR2 (N6673, N6644, N4180);
xor XOR2 (N6674, N6668, N4213);
or OR2 (N6675, N6672, N972);
not NOT1 (N6676, N6669);
xor XOR2 (N6677, N6675, N3597);
or OR4 (N6678, N6674, N5867, N2654, N5985);
xor XOR2 (N6679, N6678, N1534);
buf BUF1 (N6680, N6671);
nor NOR4 (N6681, N6666, N4736, N2940, N346);
nor NOR3 (N6682, N6676, N2905, N3483);
or OR4 (N6683, N6679, N5633, N1245, N2808);
not NOT1 (N6684, N6680);
nor NOR4 (N6685, N6661, N5164, N6613, N4397);
nand NAND4 (N6686, N6684, N1246, N6437, N3457);
buf BUF1 (N6687, N6667);
xor XOR2 (N6688, N6683, N2348);
nand NAND4 (N6689, N6659, N4747, N1462, N6280);
xor XOR2 (N6690, N6677, N865);
nand NAND3 (N6691, N6665, N4307, N2419);
or OR4 (N6692, N6690, N66, N6182, N3293);
nand NAND4 (N6693, N6689, N5431, N5569, N2126);
nand NAND2 (N6694, N6688, N718);
nand NAND3 (N6695, N6685, N355, N6417);
nand NAND4 (N6696, N6693, N1090, N2728, N1889);
or OR4 (N6697, N6695, N2010, N4826, N3051);
xor XOR2 (N6698, N6686, N150);
not NOT1 (N6699, N6698);
buf BUF1 (N6700, N6692);
and AND3 (N6701, N6697, N6272, N3499);
or OR4 (N6702, N6682, N5979, N4137, N14);
not NOT1 (N6703, N6702);
xor XOR2 (N6704, N6681, N2043);
buf BUF1 (N6705, N6704);
not NOT1 (N6706, N6694);
not NOT1 (N6707, N6703);
buf BUF1 (N6708, N6705);
or OR4 (N6709, N6706, N6046, N1349, N625);
not NOT1 (N6710, N6709);
nor NOR4 (N6711, N6687, N5304, N530, N1039);
not NOT1 (N6712, N6711);
or OR3 (N6713, N6712, N1476, N5123);
xor XOR2 (N6714, N6713, N2298);
buf BUF1 (N6715, N6696);
nand NAND4 (N6716, N6691, N2646, N3659, N3430);
nor NOR2 (N6717, N6708, N10);
not NOT1 (N6718, N6700);
or OR4 (N6719, N6710, N3431, N1769, N3308);
and AND2 (N6720, N6701, N449);
nor NOR3 (N6721, N6718, N5794, N2087);
not NOT1 (N6722, N6721);
not NOT1 (N6723, N6673);
nor NOR4 (N6724, N6715, N1316, N1611, N5536);
not NOT1 (N6725, N6719);
nor NOR3 (N6726, N6717, N1626, N2057);
and AND4 (N6727, N6726, N6245, N1400, N6191);
and AND3 (N6728, N6725, N2838, N3251);
not NOT1 (N6729, N6724);
and AND2 (N6730, N6728, N4298);
or OR2 (N6731, N6699, N1994);
and AND4 (N6732, N6731, N1699, N2196, N3221);
not NOT1 (N6733, N6716);
or OR3 (N6734, N6707, N3075, N4125);
buf BUF1 (N6735, N6733);
and AND3 (N6736, N6730, N3164, N6238);
xor XOR2 (N6737, N6734, N5743);
or OR3 (N6738, N6732, N4783, N3299);
nand NAND3 (N6739, N6714, N3201, N2933);
nand NAND3 (N6740, N6739, N1021, N1570);
buf BUF1 (N6741, N6723);
xor XOR2 (N6742, N6722, N5806);
nand NAND4 (N6743, N6738, N2909, N4336, N2604);
xor XOR2 (N6744, N6741, N3094);
not NOT1 (N6745, N6744);
buf BUF1 (N6746, N6720);
and AND2 (N6747, N6742, N3081);
and AND4 (N6748, N6743, N4014, N5843, N4083);
buf BUF1 (N6749, N6745);
and AND3 (N6750, N6749, N1765, N1047);
or OR3 (N6751, N6740, N219, N315);
nand NAND3 (N6752, N6748, N5220, N4728);
xor XOR2 (N6753, N6747, N1658);
not NOT1 (N6754, N6753);
and AND4 (N6755, N6750, N4705, N3599, N2271);
nor NOR2 (N6756, N6755, N6665);
nand NAND3 (N6757, N6727, N3734, N3391);
or OR2 (N6758, N6751, N3333);
buf BUF1 (N6759, N6756);
not NOT1 (N6760, N6759);
and AND3 (N6761, N6735, N5441, N5055);
and AND3 (N6762, N6760, N577, N4416);
nor NOR3 (N6763, N6762, N683, N1906);
buf BUF1 (N6764, N6746);
or OR3 (N6765, N6752, N4921, N5300);
nor NOR2 (N6766, N6757, N983);
or OR2 (N6767, N6736, N6366);
or OR4 (N6768, N6758, N3570, N240, N1628);
buf BUF1 (N6769, N6729);
nor NOR4 (N6770, N6754, N5076, N6174, N65);
xor XOR2 (N6771, N6767, N214);
buf BUF1 (N6772, N6770);
and AND3 (N6773, N6766, N5235, N4516);
and AND4 (N6774, N6737, N6261, N6691, N6734);
nor NOR3 (N6775, N6769, N2620, N4210);
nor NOR3 (N6776, N6765, N1599, N4028);
buf BUF1 (N6777, N6773);
and AND3 (N6778, N6775, N3778, N6069);
nor NOR2 (N6779, N6771, N893);
and AND2 (N6780, N6761, N4432);
not NOT1 (N6781, N6774);
buf BUF1 (N6782, N6763);
buf BUF1 (N6783, N6768);
nand NAND3 (N6784, N6777, N48, N1158);
not NOT1 (N6785, N6780);
nor NOR3 (N6786, N6784, N3303, N5856);
nor NOR4 (N6787, N6778, N5357, N161, N4055);
xor XOR2 (N6788, N6783, N1632);
and AND3 (N6789, N6764, N419, N3314);
and AND4 (N6790, N6779, N598, N4614, N5052);
or OR2 (N6791, N6788, N1961);
not NOT1 (N6792, N6776);
nor NOR3 (N6793, N6781, N4285, N6554);
nor NOR2 (N6794, N6791, N1318);
and AND2 (N6795, N6787, N649);
or OR4 (N6796, N6772, N3324, N2487, N2718);
nor NOR3 (N6797, N6785, N4284, N931);
and AND3 (N6798, N6786, N3994, N1184);
not NOT1 (N6799, N6792);
and AND3 (N6800, N6790, N3557, N2197);
nor NOR4 (N6801, N6795, N2965, N3111, N782);
buf BUF1 (N6802, N6801);
buf BUF1 (N6803, N6793);
and AND4 (N6804, N6797, N1725, N5671, N2163);
nor NOR2 (N6805, N6802, N5397);
nand NAND4 (N6806, N6798, N562, N2067, N3464);
nand NAND2 (N6807, N6805, N3808);
or OR4 (N6808, N6807, N6714, N2802, N510);
not NOT1 (N6809, N6800);
not NOT1 (N6810, N6806);
xor XOR2 (N6811, N6804, N3317);
and AND3 (N6812, N6803, N6184, N168);
xor XOR2 (N6813, N6799, N1135);
nor NOR3 (N6814, N6789, N5866, N1001);
not NOT1 (N6815, N6810);
and AND4 (N6816, N6811, N6624, N4977, N3857);
xor XOR2 (N6817, N6782, N5946);
not NOT1 (N6818, N6816);
and AND2 (N6819, N6817, N2560);
buf BUF1 (N6820, N6796);
and AND2 (N6821, N6809, N85);
buf BUF1 (N6822, N6815);
and AND3 (N6823, N6813, N3006, N4950);
buf BUF1 (N6824, N6819);
xor XOR2 (N6825, N6818, N1566);
and AND3 (N6826, N6812, N828, N5280);
xor XOR2 (N6827, N6820, N2451);
nor NOR2 (N6828, N6822, N6613);
nor NOR4 (N6829, N6808, N3318, N104, N5485);
not NOT1 (N6830, N6829);
xor XOR2 (N6831, N6824, N905);
and AND2 (N6832, N6827, N2811);
xor XOR2 (N6833, N6826, N1612);
nand NAND4 (N6834, N6821, N1427, N5554, N1104);
and AND2 (N6835, N6830, N6579);
nand NAND4 (N6836, N6828, N4151, N518, N5374);
not NOT1 (N6837, N6825);
not NOT1 (N6838, N6831);
nand NAND3 (N6839, N6823, N3985, N2795);
and AND4 (N6840, N6834, N6700, N3124, N4135);
nor NOR2 (N6841, N6840, N4665);
nor NOR2 (N6842, N6841, N1336);
xor XOR2 (N6843, N6833, N778);
not NOT1 (N6844, N6794);
not NOT1 (N6845, N6814);
or OR2 (N6846, N6842, N2598);
or OR2 (N6847, N6845, N4355);
not NOT1 (N6848, N6846);
buf BUF1 (N6849, N6839);
xor XOR2 (N6850, N6836, N6350);
or OR2 (N6851, N6838, N6418);
or OR3 (N6852, N6837, N1304, N2933);
buf BUF1 (N6853, N6851);
nor NOR4 (N6854, N6852, N4416, N6081, N2196);
nand NAND3 (N6855, N6832, N5900, N2447);
or OR4 (N6856, N6835, N2618, N4054, N3918);
and AND4 (N6857, N6856, N6050, N2145, N1996);
nand NAND3 (N6858, N6854, N661, N1966);
nor NOR3 (N6859, N6849, N6260, N3486);
and AND2 (N6860, N6859, N4725);
xor XOR2 (N6861, N6860, N4030);
nand NAND3 (N6862, N6843, N3468, N2096);
nor NOR4 (N6863, N6862, N840, N6176, N4659);
xor XOR2 (N6864, N6855, N4132);
and AND2 (N6865, N6857, N5457);
and AND3 (N6866, N6850, N4861, N2531);
nor NOR2 (N6867, N6853, N4217);
buf BUF1 (N6868, N6848);
xor XOR2 (N6869, N6847, N816);
buf BUF1 (N6870, N6858);
nand NAND4 (N6871, N6861, N6706, N3424, N6049);
not NOT1 (N6872, N6867);
buf BUF1 (N6873, N6870);
xor XOR2 (N6874, N6844, N356);
or OR2 (N6875, N6874, N4923);
buf BUF1 (N6876, N6869);
not NOT1 (N6877, N6863);
buf BUF1 (N6878, N6873);
buf BUF1 (N6879, N6878);
buf BUF1 (N6880, N6868);
or OR3 (N6881, N6877, N5572, N4286);
xor XOR2 (N6882, N6876, N846);
buf BUF1 (N6883, N6866);
buf BUF1 (N6884, N6875);
nand NAND4 (N6885, N6880, N125, N4468, N3179);
nor NOR2 (N6886, N6881, N6380);
or OR3 (N6887, N6879, N6300, N4259);
xor XOR2 (N6888, N6864, N1538);
nand NAND2 (N6889, N6887, N2873);
nand NAND4 (N6890, N6882, N6349, N4518, N897);
xor XOR2 (N6891, N6884, N3812);
nand NAND3 (N6892, N6888, N343, N1168);
buf BUF1 (N6893, N6892);
nor NOR3 (N6894, N6893, N4773, N602);
and AND2 (N6895, N6894, N421);
and AND4 (N6896, N6886, N1781, N2848, N4508);
or OR2 (N6897, N6889, N3062);
nor NOR3 (N6898, N6891, N74, N4570);
nand NAND4 (N6899, N6865, N977, N6297, N4901);
nand NAND2 (N6900, N6883, N6285);
nor NOR3 (N6901, N6899, N2869, N4968);
not NOT1 (N6902, N6885);
nand NAND2 (N6903, N6871, N5506);
nand NAND4 (N6904, N6890, N6193, N6161, N5324);
nand NAND2 (N6905, N6903, N851);
nor NOR2 (N6906, N6900, N4041);
or OR3 (N6907, N6902, N4061, N3395);
xor XOR2 (N6908, N6906, N4996);
nor NOR3 (N6909, N6905, N1931, N2857);
nand NAND3 (N6910, N6909, N563, N1943);
xor XOR2 (N6911, N6896, N2316);
not NOT1 (N6912, N6897);
xor XOR2 (N6913, N6908, N3177);
nand NAND3 (N6914, N6911, N4190, N4247);
nor NOR4 (N6915, N6872, N6891, N3164, N4508);
buf BUF1 (N6916, N6910);
buf BUF1 (N6917, N6895);
and AND2 (N6918, N6913, N6109);
buf BUF1 (N6919, N6907);
not NOT1 (N6920, N6898);
nand NAND4 (N6921, N6915, N5941, N6565, N3458);
buf BUF1 (N6922, N6921);
buf BUF1 (N6923, N6904);
and AND3 (N6924, N6923, N6122, N6260);
nor NOR3 (N6925, N6917, N5159, N6467);
not NOT1 (N6926, N6901);
xor XOR2 (N6927, N6925, N6429);
buf BUF1 (N6928, N6922);
nand NAND2 (N6929, N6918, N239);
xor XOR2 (N6930, N6926, N1651);
buf BUF1 (N6931, N6914);
and AND4 (N6932, N6919, N1810, N393, N3279);
nand NAND2 (N6933, N6930, N2118);
not NOT1 (N6934, N6916);
xor XOR2 (N6935, N6929, N2882);
buf BUF1 (N6936, N6935);
buf BUF1 (N6937, N6932);
buf BUF1 (N6938, N6912);
or OR4 (N6939, N6934, N2495, N122, N5364);
not NOT1 (N6940, N6920);
xor XOR2 (N6941, N6937, N5331);
nand NAND4 (N6942, N6931, N3942, N6678, N3835);
not NOT1 (N6943, N6939);
and AND2 (N6944, N6933, N5247);
xor XOR2 (N6945, N6942, N5190);
nand NAND3 (N6946, N6936, N4857, N2810);
nor NOR2 (N6947, N6941, N2174);
not NOT1 (N6948, N6946);
or OR3 (N6949, N6927, N1091, N4006);
not NOT1 (N6950, N6949);
nand NAND4 (N6951, N6938, N794, N2622, N4695);
or OR4 (N6952, N6945, N1651, N4887, N612);
or OR2 (N6953, N6948, N686);
and AND3 (N6954, N6924, N2981, N4073);
and AND3 (N6955, N6943, N1270, N2524);
and AND2 (N6956, N6947, N2296);
nand NAND3 (N6957, N6928, N3706, N3645);
and AND3 (N6958, N6955, N5603, N738);
nand NAND3 (N6959, N6958, N2528, N835);
nor NOR3 (N6960, N6940, N423, N6108);
buf BUF1 (N6961, N6953);
xor XOR2 (N6962, N6957, N571);
nor NOR4 (N6963, N6952, N4145, N5860, N5423);
nand NAND4 (N6964, N6954, N5384, N6072, N6050);
buf BUF1 (N6965, N6956);
or OR3 (N6966, N6959, N3453, N5691);
or OR3 (N6967, N6960, N5211, N2634);
nor NOR3 (N6968, N6951, N5524, N4002);
xor XOR2 (N6969, N6968, N44);
and AND4 (N6970, N6964, N3681, N2407, N3571);
and AND3 (N6971, N6965, N3720, N2302);
buf BUF1 (N6972, N6963);
nand NAND3 (N6973, N6969, N2666, N126);
xor XOR2 (N6974, N6961, N5575);
buf BUF1 (N6975, N6967);
and AND3 (N6976, N6966, N2769, N1561);
not NOT1 (N6977, N6974);
nor NOR4 (N6978, N6962, N1737, N3316, N3707);
not NOT1 (N6979, N6971);
buf BUF1 (N6980, N6979);
nor NOR4 (N6981, N6975, N2432, N1918, N2575);
xor XOR2 (N6982, N6978, N5227);
or OR3 (N6983, N6973, N1558, N6504);
nand NAND4 (N6984, N6982, N6602, N1063, N4788);
nand NAND4 (N6985, N6980, N4999, N1438, N3970);
nand NAND2 (N6986, N6981, N5315);
not NOT1 (N6987, N6970);
nor NOR4 (N6988, N6972, N1618, N4115, N1649);
buf BUF1 (N6989, N6988);
nand NAND3 (N6990, N6984, N151, N3008);
and AND3 (N6991, N6977, N3152, N6427);
nor NOR2 (N6992, N6944, N5290);
or OR4 (N6993, N6976, N6097, N896, N3408);
nand NAND2 (N6994, N6989, N3991);
buf BUF1 (N6995, N6985);
buf BUF1 (N6996, N6991);
or OR4 (N6997, N6996, N5789, N6807, N3149);
and AND4 (N6998, N6994, N1901, N2886, N5075);
or OR4 (N6999, N6995, N1377, N1776, N5509);
not NOT1 (N7000, N6998);
not NOT1 (N7001, N6983);
and AND3 (N7002, N6993, N1028, N2965);
not NOT1 (N7003, N7001);
xor XOR2 (N7004, N6986, N395);
nand NAND3 (N7005, N6950, N1977, N5189);
nand NAND4 (N7006, N6997, N151, N2707, N4914);
nor NOR3 (N7007, N6990, N5012, N378);
xor XOR2 (N7008, N7005, N4282);
nor NOR3 (N7009, N7007, N4471, N1461);
nor NOR4 (N7010, N7004, N418, N4470, N6875);
or OR2 (N7011, N7010, N1649);
nor NOR4 (N7012, N7003, N2000, N1909, N2509);
nor NOR3 (N7013, N7006, N202, N3639);
nor NOR3 (N7014, N7011, N1020, N5461);
not NOT1 (N7015, N7012);
nand NAND3 (N7016, N7008, N1385, N3598);
not NOT1 (N7017, N7013);
xor XOR2 (N7018, N7000, N6884);
not NOT1 (N7019, N7018);
not NOT1 (N7020, N7014);
buf BUF1 (N7021, N7002);
xor XOR2 (N7022, N6999, N6857);
nand NAND3 (N7023, N7015, N6469, N350);
or OR4 (N7024, N7022, N2764, N4833, N1891);
xor XOR2 (N7025, N7020, N6777);
and AND4 (N7026, N7017, N477, N3372, N4847);
not NOT1 (N7027, N7009);
and AND2 (N7028, N7021, N982);
buf BUF1 (N7029, N7019);
xor XOR2 (N7030, N6987, N1143);
buf BUF1 (N7031, N7030);
nand NAND3 (N7032, N7016, N6626, N4718);
xor XOR2 (N7033, N6992, N6102);
buf BUF1 (N7034, N7031);
xor XOR2 (N7035, N7034, N2755);
nand NAND2 (N7036, N7026, N6490);
xor XOR2 (N7037, N7029, N5768);
nor NOR2 (N7038, N7036, N1294);
xor XOR2 (N7039, N7025, N6140);
or OR2 (N7040, N7037, N7020);
or OR4 (N7041, N7039, N800, N3728, N5250);
xor XOR2 (N7042, N7028, N6204);
not NOT1 (N7043, N7042);
buf BUF1 (N7044, N7043);
buf BUF1 (N7045, N7038);
buf BUF1 (N7046, N7027);
or OR3 (N7047, N7032, N3428, N968);
xor XOR2 (N7048, N7040, N1548);
nand NAND3 (N7049, N7041, N3790, N2614);
xor XOR2 (N7050, N7044, N3937);
nand NAND3 (N7051, N7033, N6040, N4289);
nor NOR3 (N7052, N7048, N6008, N45);
or OR2 (N7053, N7023, N3056);
nand NAND4 (N7054, N7035, N5493, N6441, N5348);
nor NOR2 (N7055, N7051, N5583);
nand NAND4 (N7056, N7052, N5969, N3729, N3336);
xor XOR2 (N7057, N7045, N3028);
nor NOR2 (N7058, N7049, N3445);
xor XOR2 (N7059, N7046, N5009);
nor NOR2 (N7060, N7057, N2167);
xor XOR2 (N7061, N7047, N2012);
and AND4 (N7062, N7059, N6059, N5344, N1236);
xor XOR2 (N7063, N7056, N3128);
buf BUF1 (N7064, N7061);
nor NOR2 (N7065, N7054, N6254);
xor XOR2 (N7066, N7058, N1748);
xor XOR2 (N7067, N7060, N346);
buf BUF1 (N7068, N7062);
buf BUF1 (N7069, N7067);
buf BUF1 (N7070, N7066);
buf BUF1 (N7071, N7064);
xor XOR2 (N7072, N7070, N5714);
nor NOR2 (N7073, N7053, N5195);
xor XOR2 (N7074, N7065, N3287);
or OR2 (N7075, N7063, N5353);
nand NAND2 (N7076, N7069, N1949);
xor XOR2 (N7077, N7071, N5966);
nor NOR2 (N7078, N7077, N1961);
nand NAND4 (N7079, N7074, N3310, N1140, N6957);
nor NOR2 (N7080, N7079, N995);
and AND4 (N7081, N7050, N4185, N6293, N1953);
nor NOR2 (N7082, N7055, N6266);
xor XOR2 (N7083, N7076, N3809);
nor NOR2 (N7084, N7081, N5061);
not NOT1 (N7085, N7083);
or OR4 (N7086, N7068, N2257, N3566, N3675);
or OR3 (N7087, N7075, N768, N2382);
buf BUF1 (N7088, N7084);
and AND3 (N7089, N7082, N1299, N413);
nand NAND2 (N7090, N7085, N1300);
xor XOR2 (N7091, N7089, N3127);
buf BUF1 (N7092, N7080);
xor XOR2 (N7093, N7078, N2746);
buf BUF1 (N7094, N7072);
xor XOR2 (N7095, N7088, N5695);
or OR2 (N7096, N7091, N3074);
or OR2 (N7097, N7093, N6402);
nor NOR2 (N7098, N7087, N3880);
nand NAND2 (N7099, N7092, N2435);
or OR4 (N7100, N7024, N5394, N440, N1813);
xor XOR2 (N7101, N7094, N6875);
not NOT1 (N7102, N7095);
not NOT1 (N7103, N7098);
xor XOR2 (N7104, N7100, N1624);
not NOT1 (N7105, N7104);
buf BUF1 (N7106, N7097);
and AND4 (N7107, N7090, N2768, N6688, N6933);
nor NOR4 (N7108, N7103, N6711, N4746, N1581);
xor XOR2 (N7109, N7106, N1495);
and AND2 (N7110, N7108, N1631);
and AND3 (N7111, N7086, N5779, N6866);
nand NAND4 (N7112, N7109, N2685, N963, N2753);
and AND4 (N7113, N7112, N28, N5145, N6188);
nand NAND4 (N7114, N7107, N6069, N1671, N5500);
nand NAND2 (N7115, N7073, N1981);
not NOT1 (N7116, N7105);
nand NAND2 (N7117, N7101, N6834);
or OR3 (N7118, N7096, N3115, N2856);
buf BUF1 (N7119, N7115);
and AND2 (N7120, N7117, N5856);
not NOT1 (N7121, N7102);
nand NAND2 (N7122, N7110, N4789);
and AND3 (N7123, N7119, N2913, N1418);
buf BUF1 (N7124, N7121);
nand NAND4 (N7125, N7118, N339, N3663, N4717);
and AND3 (N7126, N7113, N6394, N6144);
not NOT1 (N7127, N7122);
xor XOR2 (N7128, N7124, N169);
not NOT1 (N7129, N7114);
nor NOR2 (N7130, N7116, N1874);
or OR2 (N7131, N7123, N3193);
and AND4 (N7132, N7126, N3204, N1702, N6230);
nand NAND3 (N7133, N7120, N5882, N2298);
nor NOR3 (N7134, N7099, N5011, N3766);
or OR3 (N7135, N7125, N3946, N5632);
and AND2 (N7136, N7129, N4832);
buf BUF1 (N7137, N7132);
and AND4 (N7138, N7137, N4290, N5539, N2537);
nor NOR2 (N7139, N7138, N101);
nor NOR3 (N7140, N7131, N4932, N2912);
or OR2 (N7141, N7139, N5308);
nor NOR2 (N7142, N7141, N6557);
not NOT1 (N7143, N7135);
and AND2 (N7144, N7127, N2143);
nor NOR2 (N7145, N7133, N780);
or OR2 (N7146, N7140, N5602);
xor XOR2 (N7147, N7136, N1701);
not NOT1 (N7148, N7146);
buf BUF1 (N7149, N7111);
and AND2 (N7150, N7148, N2557);
not NOT1 (N7151, N7134);
nor NOR3 (N7152, N7151, N6212, N1116);
buf BUF1 (N7153, N7142);
nor NOR4 (N7154, N7147, N2341, N6850, N310);
buf BUF1 (N7155, N7128);
nor NOR4 (N7156, N7152, N287, N1914, N671);
xor XOR2 (N7157, N7149, N1196);
nand NAND4 (N7158, N7143, N6707, N2581, N346);
or OR4 (N7159, N7156, N3866, N3578, N4539);
nor NOR4 (N7160, N7155, N6475, N2336, N5372);
nand NAND3 (N7161, N7159, N1291, N4188);
xor XOR2 (N7162, N7161, N2131);
and AND4 (N7163, N7144, N4612, N3659, N3629);
nand NAND2 (N7164, N7154, N395);
not NOT1 (N7165, N7157);
buf BUF1 (N7166, N7165);
nand NAND3 (N7167, N7162, N322, N1340);
and AND4 (N7168, N7164, N2397, N3891, N405);
xor XOR2 (N7169, N7153, N7006);
or OR3 (N7170, N7168, N3020, N2801);
or OR2 (N7171, N7169, N5355);
xor XOR2 (N7172, N7170, N2799);
nand NAND4 (N7173, N7163, N968, N6547, N3538);
or OR3 (N7174, N7130, N5866, N4185);
or OR4 (N7175, N7166, N7171, N1447, N1164);
nor NOR3 (N7176, N1643, N2657, N5207);
and AND2 (N7177, N7167, N5176);
and AND3 (N7178, N7177, N5985, N333);
xor XOR2 (N7179, N7160, N353);
xor XOR2 (N7180, N7145, N6218);
and AND3 (N7181, N7174, N5299, N4723);
xor XOR2 (N7182, N7181, N3977);
and AND3 (N7183, N7173, N6608, N5847);
nand NAND4 (N7184, N7182, N4861, N5091, N4812);
nand NAND3 (N7185, N7180, N5246, N6122);
nor NOR2 (N7186, N7175, N5716);
and AND4 (N7187, N7183, N3859, N276, N449);
and AND4 (N7188, N7185, N2629, N5339, N20);
nor NOR2 (N7189, N7186, N4868);
xor XOR2 (N7190, N7176, N2888);
and AND4 (N7191, N7158, N5227, N5128, N1840);
nor NOR3 (N7192, N7189, N1395, N2329);
nand NAND2 (N7193, N7191, N2101);
buf BUF1 (N7194, N7187);
nand NAND4 (N7195, N7184, N3927, N3614, N4917);
and AND3 (N7196, N7194, N5337, N971);
xor XOR2 (N7197, N7190, N551);
or OR4 (N7198, N7196, N183, N5121, N6832);
not NOT1 (N7199, N7192);
nand NAND4 (N7200, N7198, N2275, N1829, N4079);
buf BUF1 (N7201, N7179);
not NOT1 (N7202, N7197);
or OR4 (N7203, N7193, N3891, N1127, N4191);
buf BUF1 (N7204, N7200);
nor NOR2 (N7205, N7204, N6374);
and AND3 (N7206, N7188, N3677, N5472);
not NOT1 (N7207, N7199);
nand NAND2 (N7208, N7202, N3113);
nor NOR3 (N7209, N7178, N5906, N5236);
nor NOR4 (N7210, N7206, N6139, N5486, N4717);
buf BUF1 (N7211, N7201);
not NOT1 (N7212, N7205);
buf BUF1 (N7213, N7211);
xor XOR2 (N7214, N7213, N6132);
nor NOR3 (N7215, N7214, N6144, N7045);
nand NAND4 (N7216, N7212, N2541, N1562, N3370);
buf BUF1 (N7217, N7209);
not NOT1 (N7218, N7195);
and AND3 (N7219, N7203, N4091, N3672);
buf BUF1 (N7220, N7215);
and AND4 (N7221, N7216, N3654, N1025, N2427);
buf BUF1 (N7222, N7172);
nor NOR4 (N7223, N7217, N94, N7041, N2510);
nor NOR4 (N7224, N7218, N3155, N1143, N1077);
or OR2 (N7225, N7221, N5455);
xor XOR2 (N7226, N7150, N893);
and AND2 (N7227, N7219, N5612);
or OR2 (N7228, N7220, N1356);
xor XOR2 (N7229, N7222, N3240);
nor NOR3 (N7230, N7207, N2927, N2563);
buf BUF1 (N7231, N7224);
nor NOR4 (N7232, N7210, N908, N3864, N6242);
nor NOR3 (N7233, N7231, N51, N1823);
buf BUF1 (N7234, N7227);
and AND2 (N7235, N7232, N4077);
nor NOR2 (N7236, N7234, N5116);
nor NOR4 (N7237, N7233, N510, N6243, N1444);
and AND3 (N7238, N7225, N370, N672);
buf BUF1 (N7239, N7230);
buf BUF1 (N7240, N7237);
xor XOR2 (N7241, N7236, N3018);
and AND3 (N7242, N7208, N4806, N5257);
not NOT1 (N7243, N7238);
nor NOR4 (N7244, N7240, N511, N6885, N4730);
xor XOR2 (N7245, N7229, N1833);
nand NAND3 (N7246, N7243, N1701, N6510);
not NOT1 (N7247, N7244);
and AND2 (N7248, N7239, N2685);
or OR2 (N7249, N7242, N2547);
buf BUF1 (N7250, N7241);
xor XOR2 (N7251, N7226, N2738);
buf BUF1 (N7252, N7235);
buf BUF1 (N7253, N7247);
nand NAND3 (N7254, N7250, N44, N3592);
xor XOR2 (N7255, N7223, N4383);
buf BUF1 (N7256, N7251);
nor NOR2 (N7257, N7254, N4728);
xor XOR2 (N7258, N7228, N1183);
nor NOR3 (N7259, N7255, N2030, N2744);
xor XOR2 (N7260, N7258, N3057);
nor NOR4 (N7261, N7249, N703, N3324, N3273);
xor XOR2 (N7262, N7252, N277);
nand NAND3 (N7263, N7260, N2683, N4808);
buf BUF1 (N7264, N7262);
buf BUF1 (N7265, N7259);
nand NAND4 (N7266, N7253, N5493, N2166, N5826);
or OR4 (N7267, N7245, N1887, N1573, N157);
or OR2 (N7268, N7263, N6302);
and AND2 (N7269, N7248, N2183);
or OR2 (N7270, N7269, N3116);
and AND2 (N7271, N7268, N2003);
and AND2 (N7272, N7265, N3669);
nand NAND3 (N7273, N7267, N6049, N2110);
nand NAND2 (N7274, N7246, N6304);
not NOT1 (N7275, N7271);
not NOT1 (N7276, N7257);
xor XOR2 (N7277, N7270, N2759);
nand NAND3 (N7278, N7275, N4742, N3390);
not NOT1 (N7279, N7272);
or OR2 (N7280, N7276, N7258);
or OR2 (N7281, N7256, N2279);
xor XOR2 (N7282, N7277, N3031);
and AND2 (N7283, N7266, N3047);
buf BUF1 (N7284, N7264);
or OR4 (N7285, N7278, N2444, N1243, N3291);
nand NAND3 (N7286, N7273, N1320, N3750);
buf BUF1 (N7287, N7282);
buf BUF1 (N7288, N7280);
or OR4 (N7289, N7279, N7155, N3714, N6267);
nor NOR4 (N7290, N7274, N3448, N5308, N3343);
and AND3 (N7291, N7286, N6036, N6210);
nand NAND4 (N7292, N7289, N4716, N3072, N4327);
nand NAND4 (N7293, N7285, N2735, N3022, N415);
nor NOR2 (N7294, N7284, N3830);
nand NAND2 (N7295, N7281, N6275);
or OR4 (N7296, N7287, N6239, N3568, N2490);
nor NOR3 (N7297, N7283, N2041, N6754);
nand NAND2 (N7298, N7261, N1367);
xor XOR2 (N7299, N7296, N4448);
buf BUF1 (N7300, N7294);
nand NAND2 (N7301, N7291, N4120);
and AND2 (N7302, N7298, N3054);
nor NOR4 (N7303, N7297, N306, N4779, N31);
nor NOR4 (N7304, N7299, N448, N1336, N6852);
and AND2 (N7305, N7304, N2972);
or OR2 (N7306, N7295, N1193);
nand NAND4 (N7307, N7293, N3305, N4051, N6117);
or OR2 (N7308, N7292, N6558);
nand NAND3 (N7309, N7305, N4716, N2993);
xor XOR2 (N7310, N7302, N489);
xor XOR2 (N7311, N7310, N5925);
buf BUF1 (N7312, N7300);
or OR2 (N7313, N7311, N3017);
nor NOR2 (N7314, N7306, N191);
buf BUF1 (N7315, N7301);
nand NAND4 (N7316, N7309, N3383, N410, N6598);
not NOT1 (N7317, N7307);
nand NAND2 (N7318, N7314, N190);
nand NAND3 (N7319, N7312, N5151, N715);
nand NAND4 (N7320, N7288, N1052, N3341, N6413);
not NOT1 (N7321, N7303);
xor XOR2 (N7322, N7308, N3101);
or OR4 (N7323, N7321, N6081, N5261, N7272);
nand NAND3 (N7324, N7322, N710, N4953);
xor XOR2 (N7325, N7315, N858);
xor XOR2 (N7326, N7323, N7035);
not NOT1 (N7327, N7316);
not NOT1 (N7328, N7319);
xor XOR2 (N7329, N7317, N1984);
xor XOR2 (N7330, N7325, N2135);
nand NAND4 (N7331, N7318, N2089, N3873, N3105);
or OR4 (N7332, N7290, N3599, N68, N4097);
nor NOR4 (N7333, N7313, N2531, N5348, N6787);
not NOT1 (N7334, N7333);
xor XOR2 (N7335, N7334, N3398);
nor NOR4 (N7336, N7328, N6994, N984, N2436);
and AND3 (N7337, N7326, N6225, N3934);
nor NOR4 (N7338, N7327, N4752, N2687, N4135);
and AND2 (N7339, N7336, N3124);
nor NOR4 (N7340, N7337, N2789, N5248, N1289);
not NOT1 (N7341, N7330);
nor NOR4 (N7342, N7324, N3162, N4989, N3713);
xor XOR2 (N7343, N7331, N7003);
xor XOR2 (N7344, N7341, N6327);
not NOT1 (N7345, N7320);
not NOT1 (N7346, N7335);
nor NOR3 (N7347, N7343, N5038, N5953);
not NOT1 (N7348, N7339);
xor XOR2 (N7349, N7332, N3413);
buf BUF1 (N7350, N7344);
not NOT1 (N7351, N7347);
buf BUF1 (N7352, N7342);
and AND3 (N7353, N7329, N942, N158);
buf BUF1 (N7354, N7353);
xor XOR2 (N7355, N7354, N6220);
buf BUF1 (N7356, N7340);
nand NAND4 (N7357, N7348, N4474, N729, N6204);
nor NOR4 (N7358, N7357, N6678, N4519, N1290);
and AND2 (N7359, N7349, N5295);
buf BUF1 (N7360, N7350);
nor NOR3 (N7361, N7351, N5595, N6129);
and AND4 (N7362, N7358, N214, N982, N2563);
buf BUF1 (N7363, N7346);
and AND4 (N7364, N7352, N6709, N5284, N7134);
nand NAND4 (N7365, N7338, N3585, N1944, N3877);
and AND4 (N7366, N7345, N1257, N2074, N2447);
nand NAND2 (N7367, N7361, N6699);
not NOT1 (N7368, N7367);
or OR3 (N7369, N7360, N1000, N7027);
xor XOR2 (N7370, N7362, N4406);
buf BUF1 (N7371, N7359);
nand NAND3 (N7372, N7355, N2207, N5340);
or OR4 (N7373, N7371, N5305, N4752, N2657);
nand NAND2 (N7374, N7370, N3910);
not NOT1 (N7375, N7363);
nor NOR4 (N7376, N7374, N6518, N436, N368);
xor XOR2 (N7377, N7364, N6040);
not NOT1 (N7378, N7365);
nor NOR3 (N7379, N7376, N1108, N5277);
nor NOR3 (N7380, N7368, N3373, N379);
not NOT1 (N7381, N7378);
or OR3 (N7382, N7366, N5778, N5969);
buf BUF1 (N7383, N7381);
xor XOR2 (N7384, N7375, N6976);
or OR3 (N7385, N7377, N5281, N6738);
not NOT1 (N7386, N7372);
nand NAND2 (N7387, N7369, N6414);
not NOT1 (N7388, N7373);
not NOT1 (N7389, N7356);
xor XOR2 (N7390, N7383, N6298);
buf BUF1 (N7391, N7389);
buf BUF1 (N7392, N7384);
not NOT1 (N7393, N7380);
or OR2 (N7394, N7388, N1237);
not NOT1 (N7395, N7393);
nand NAND4 (N7396, N7387, N297, N3402, N2725);
not NOT1 (N7397, N7391);
xor XOR2 (N7398, N7397, N5431);
and AND3 (N7399, N7392, N1030, N6581);
buf BUF1 (N7400, N7390);
or OR3 (N7401, N7385, N1920, N946);
not NOT1 (N7402, N7394);
xor XOR2 (N7403, N7396, N6075);
buf BUF1 (N7404, N7386);
not NOT1 (N7405, N7382);
buf BUF1 (N7406, N7395);
not NOT1 (N7407, N7401);
and AND4 (N7408, N7398, N4192, N1879, N5429);
and AND3 (N7409, N7404, N5997, N1828);
nor NOR2 (N7410, N7408, N7287);
buf BUF1 (N7411, N7399);
nor NOR2 (N7412, N7411, N3426);
buf BUF1 (N7413, N7405);
xor XOR2 (N7414, N7412, N6324);
buf BUF1 (N7415, N7414);
buf BUF1 (N7416, N7407);
nor NOR3 (N7417, N7410, N108, N1458);
nand NAND2 (N7418, N7413, N4227);
or OR3 (N7419, N7416, N6945, N2822);
nand NAND2 (N7420, N7418, N1791);
or OR4 (N7421, N7406, N2731, N3043, N6250);
nand NAND3 (N7422, N7421, N1194, N4636);
or OR2 (N7423, N7420, N3);
or OR2 (N7424, N7403, N158);
and AND2 (N7425, N7402, N2953);
and AND2 (N7426, N7422, N5659);
and AND3 (N7427, N7424, N2467, N6763);
nand NAND4 (N7428, N7379, N2661, N1407, N795);
buf BUF1 (N7429, N7415);
nand NAND4 (N7430, N7427, N4827, N2159, N220);
or OR4 (N7431, N7428, N2712, N4525, N5707);
buf BUF1 (N7432, N7426);
or OR4 (N7433, N7423, N4441, N4151, N5333);
nand NAND2 (N7434, N7419, N3051);
not NOT1 (N7435, N7432);
and AND3 (N7436, N7417, N6837, N6263);
xor XOR2 (N7437, N7429, N4299);
and AND3 (N7438, N7409, N1269, N128);
xor XOR2 (N7439, N7436, N4942);
and AND3 (N7440, N7434, N2711, N4490);
nand NAND2 (N7441, N7430, N2092);
not NOT1 (N7442, N7425);
not NOT1 (N7443, N7437);
nand NAND2 (N7444, N7400, N5864);
not NOT1 (N7445, N7444);
not NOT1 (N7446, N7441);
not NOT1 (N7447, N7431);
not NOT1 (N7448, N7446);
not NOT1 (N7449, N7435);
nand NAND3 (N7450, N7442, N29, N4530);
nand NAND4 (N7451, N7449, N6931, N7284, N1384);
nand NAND3 (N7452, N7433, N5468, N4477);
or OR3 (N7453, N7448, N1688, N1422);
buf BUF1 (N7454, N7453);
xor XOR2 (N7455, N7440, N3962);
nor NOR3 (N7456, N7438, N1018, N1432);
and AND4 (N7457, N7452, N5770, N2600, N6208);
or OR3 (N7458, N7455, N3344, N1020);
nor NOR4 (N7459, N7443, N2937, N3400, N2055);
not NOT1 (N7460, N7439);
nand NAND3 (N7461, N7459, N2892, N2589);
nor NOR4 (N7462, N7450, N5708, N378, N404);
xor XOR2 (N7463, N7461, N2644);
and AND4 (N7464, N7463, N1487, N2107, N4983);
and AND2 (N7465, N7460, N4928);
buf BUF1 (N7466, N7464);
or OR3 (N7467, N7447, N4327, N7171);
xor XOR2 (N7468, N7462, N6498);
not NOT1 (N7469, N7466);
and AND4 (N7470, N7451, N3719, N848, N3642);
buf BUF1 (N7471, N7457);
and AND2 (N7472, N7467, N6394);
not NOT1 (N7473, N7469);
nor NOR2 (N7474, N7470, N761);
or OR2 (N7475, N7458, N1422);
or OR4 (N7476, N7474, N3019, N7163, N6147);
nor NOR3 (N7477, N7475, N5259, N2419);
nand NAND3 (N7478, N7476, N6301, N5421);
buf BUF1 (N7479, N7478);
buf BUF1 (N7480, N7471);
nor NOR4 (N7481, N7454, N6635, N474, N86);
not NOT1 (N7482, N7472);
or OR4 (N7483, N7479, N5228, N4911, N1760);
xor XOR2 (N7484, N7445, N5799);
nor NOR4 (N7485, N7483, N2424, N3248, N889);
nor NOR3 (N7486, N7482, N5333, N4746);
nand NAND3 (N7487, N7473, N1258, N6201);
and AND3 (N7488, N7477, N3075, N1911);
nor NOR2 (N7489, N7456, N333);
and AND2 (N7490, N7484, N1636);
xor XOR2 (N7491, N7480, N4774);
nand NAND3 (N7492, N7468, N371, N1608);
nand NAND3 (N7493, N7488, N4895, N7151);
buf BUF1 (N7494, N7493);
xor XOR2 (N7495, N7486, N4932);
or OR4 (N7496, N7491, N1417, N7204, N7391);
and AND3 (N7497, N7465, N2630, N6425);
nor NOR3 (N7498, N7492, N872, N1086);
and AND4 (N7499, N7490, N5005, N3926, N7356);
nor NOR3 (N7500, N7489, N3554, N5437);
or OR3 (N7501, N7499, N5152, N7096);
nor NOR4 (N7502, N7485, N6992, N3191, N3697);
not NOT1 (N7503, N7487);
buf BUF1 (N7504, N7500);
or OR2 (N7505, N7494, N6911);
nand NAND3 (N7506, N7502, N5858, N613);
or OR4 (N7507, N7504, N1350, N7069, N6464);
not NOT1 (N7508, N7507);
or OR2 (N7509, N7503, N1280);
or OR4 (N7510, N7496, N7405, N75, N6262);
xor XOR2 (N7511, N7505, N4563);
or OR3 (N7512, N7511, N4109, N4881);
not NOT1 (N7513, N7510);
nor NOR3 (N7514, N7497, N7333, N4510);
xor XOR2 (N7515, N7512, N6119);
or OR2 (N7516, N7506, N1343);
or OR3 (N7517, N7513, N7434, N3934);
xor XOR2 (N7518, N7509, N3923);
and AND4 (N7519, N7501, N2992, N6820, N2525);
xor XOR2 (N7520, N7516, N497);
not NOT1 (N7521, N7520);
nor NOR3 (N7522, N7514, N1346, N3546);
and AND4 (N7523, N7517, N4697, N6465, N6568);
not NOT1 (N7524, N7495);
buf BUF1 (N7525, N7518);
not NOT1 (N7526, N7521);
xor XOR2 (N7527, N7526, N5983);
not NOT1 (N7528, N7515);
and AND2 (N7529, N7523, N1120);
nor NOR2 (N7530, N7525, N1171);
nand NAND2 (N7531, N7527, N3583);
not NOT1 (N7532, N7528);
buf BUF1 (N7533, N7519);
and AND2 (N7534, N7498, N2701);
buf BUF1 (N7535, N7532);
not NOT1 (N7536, N7534);
nor NOR3 (N7537, N7529, N6030, N4507);
buf BUF1 (N7538, N7508);
nor NOR3 (N7539, N7524, N5431, N2136);
and AND3 (N7540, N7481, N7392, N177);
nor NOR4 (N7541, N7535, N2319, N2146, N2819);
or OR2 (N7542, N7536, N596);
not NOT1 (N7543, N7540);
nand NAND4 (N7544, N7531, N4887, N1068, N1742);
not NOT1 (N7545, N7541);
or OR2 (N7546, N7537, N1740);
not NOT1 (N7547, N7542);
xor XOR2 (N7548, N7522, N1473);
buf BUF1 (N7549, N7548);
nor NOR2 (N7550, N7549, N6417);
not NOT1 (N7551, N7533);
nand NAND2 (N7552, N7545, N136);
or OR4 (N7553, N7547, N5481, N7303, N4528);
and AND4 (N7554, N7543, N4232, N3288, N3717);
not NOT1 (N7555, N7544);
not NOT1 (N7556, N7553);
buf BUF1 (N7557, N7554);
xor XOR2 (N7558, N7557, N1321);
and AND4 (N7559, N7555, N5649, N6446, N7137);
and AND3 (N7560, N7530, N4322, N1880);
nor NOR2 (N7561, N7551, N7007);
nand NAND3 (N7562, N7552, N6937, N6289);
and AND3 (N7563, N7556, N4124, N2128);
not NOT1 (N7564, N7562);
nor NOR4 (N7565, N7561, N1391, N7149, N6547);
or OR4 (N7566, N7560, N5841, N2249, N4266);
buf BUF1 (N7567, N7546);
xor XOR2 (N7568, N7559, N5964);
or OR4 (N7569, N7539, N6131, N4291, N12);
buf BUF1 (N7570, N7558);
or OR4 (N7571, N7569, N4688, N108, N6542);
or OR4 (N7572, N7566, N6483, N5601, N320);
and AND4 (N7573, N7567, N5929, N3630, N2564);
or OR4 (N7574, N7538, N5166, N40, N2141);
not NOT1 (N7575, N7564);
and AND4 (N7576, N7550, N7550, N2706, N1940);
nand NAND3 (N7577, N7570, N5294, N2568);
or OR4 (N7578, N7577, N1292, N2173, N2538);
nor NOR3 (N7579, N7572, N4536, N7384);
buf BUF1 (N7580, N7579);
and AND2 (N7581, N7563, N1863);
nor NOR3 (N7582, N7565, N7237, N3005);
nor NOR2 (N7583, N7576, N7335);
buf BUF1 (N7584, N7574);
nor NOR4 (N7585, N7571, N1734, N2632, N510);
or OR4 (N7586, N7583, N5714, N4190, N1846);
xor XOR2 (N7587, N7580, N5064);
xor XOR2 (N7588, N7575, N6366);
buf BUF1 (N7589, N7586);
and AND4 (N7590, N7587, N1379, N2832, N1780);
nor NOR2 (N7591, N7584, N5774);
xor XOR2 (N7592, N7581, N6658);
xor XOR2 (N7593, N7582, N7481);
xor XOR2 (N7594, N7590, N5485);
not NOT1 (N7595, N7589);
nand NAND4 (N7596, N7592, N56, N593, N808);
nor NOR2 (N7597, N7585, N4140);
xor XOR2 (N7598, N7595, N3519);
xor XOR2 (N7599, N7596, N4365);
and AND3 (N7600, N7578, N444, N5263);
nor NOR3 (N7601, N7568, N6508, N5344);
nor NOR3 (N7602, N7597, N1431, N7182);
buf BUF1 (N7603, N7593);
and AND3 (N7604, N7588, N4604, N419);
or OR2 (N7605, N7603, N7518);
xor XOR2 (N7606, N7599, N4727);
not NOT1 (N7607, N7598);
buf BUF1 (N7608, N7591);
not NOT1 (N7609, N7600);
buf BUF1 (N7610, N7601);
nand NAND3 (N7611, N7607, N1134, N4067);
buf BUF1 (N7612, N7610);
and AND3 (N7613, N7602, N2596, N5276);
xor XOR2 (N7614, N7613, N3156);
nand NAND3 (N7615, N7573, N3710, N5962);
nor NOR4 (N7616, N7611, N5329, N1665, N3832);
nor NOR3 (N7617, N7594, N3698, N5202);
or OR2 (N7618, N7606, N3432);
and AND4 (N7619, N7605, N1196, N6556, N3688);
nand NAND3 (N7620, N7616, N1303, N2665);
nand NAND3 (N7621, N7604, N4406, N6007);
and AND4 (N7622, N7620, N287, N1222, N5279);
buf BUF1 (N7623, N7615);
nor NOR3 (N7624, N7623, N6613, N5020);
and AND4 (N7625, N7608, N3860, N1971, N7464);
xor XOR2 (N7626, N7609, N2209);
or OR2 (N7627, N7618, N378);
buf BUF1 (N7628, N7621);
nor NOR4 (N7629, N7622, N1839, N6006, N5170);
nand NAND4 (N7630, N7614, N6165, N3025, N4353);
not NOT1 (N7631, N7612);
buf BUF1 (N7632, N7626);
buf BUF1 (N7633, N7630);
and AND2 (N7634, N7619, N2402);
nor NOR3 (N7635, N7632, N928, N7211);
nand NAND4 (N7636, N7631, N4014, N4730, N5767);
and AND4 (N7637, N7635, N7089, N2615, N3335);
nand NAND3 (N7638, N7617, N6019, N7015);
nor NOR2 (N7639, N7624, N307);
nand NAND2 (N7640, N7633, N4075);
nor NOR3 (N7641, N7627, N4652, N802);
and AND2 (N7642, N7636, N7010);
buf BUF1 (N7643, N7638);
buf BUF1 (N7644, N7641);
xor XOR2 (N7645, N7640, N2374);
nor NOR4 (N7646, N7634, N759, N1675, N2643);
nor NOR4 (N7647, N7637, N5012, N4777, N5064);
buf BUF1 (N7648, N7629);
nand NAND2 (N7649, N7639, N1461);
nand NAND2 (N7650, N7645, N830);
and AND4 (N7651, N7650, N4746, N7474, N6693);
and AND4 (N7652, N7646, N3905, N4698, N3982);
nor NOR2 (N7653, N7647, N1105);
or OR4 (N7654, N7649, N2115, N5061, N1166);
buf BUF1 (N7655, N7628);
nor NOR4 (N7656, N7642, N5268, N5656, N5197);
buf BUF1 (N7657, N7643);
nand NAND3 (N7658, N7656, N1208, N7104);
nor NOR2 (N7659, N7657, N3281);
not NOT1 (N7660, N7648);
or OR4 (N7661, N7651, N2787, N231, N3747);
and AND4 (N7662, N7644, N1107, N4347, N5675);
nand NAND2 (N7663, N7658, N3141);
nand NAND3 (N7664, N7653, N3171, N5506);
not NOT1 (N7665, N7660);
not NOT1 (N7666, N7664);
not NOT1 (N7667, N7654);
nand NAND3 (N7668, N7655, N4122, N250);
nand NAND4 (N7669, N7625, N2859, N7497, N5828);
nand NAND3 (N7670, N7661, N4765, N4020);
or OR3 (N7671, N7666, N2559, N7022);
nand NAND4 (N7672, N7652, N4124, N367, N6065);
xor XOR2 (N7673, N7669, N4347);
not NOT1 (N7674, N7670);
nand NAND3 (N7675, N7667, N383, N4119);
nor NOR2 (N7676, N7671, N1123);
or OR2 (N7677, N7675, N4171);
nand NAND3 (N7678, N7677, N6576, N1721);
nand NAND2 (N7679, N7673, N2049);
and AND4 (N7680, N7659, N654, N6796, N6057);
xor XOR2 (N7681, N7680, N4399);
xor XOR2 (N7682, N7665, N7003);
and AND3 (N7683, N7662, N3887, N2257);
xor XOR2 (N7684, N7678, N860);
and AND3 (N7685, N7681, N945, N3070);
buf BUF1 (N7686, N7682);
or OR4 (N7687, N7683, N4718, N2149, N6542);
nor NOR4 (N7688, N7676, N3682, N3014, N2996);
xor XOR2 (N7689, N7684, N1252);
nor NOR4 (N7690, N7674, N128, N5923, N6745);
buf BUF1 (N7691, N7663);
nor NOR4 (N7692, N7672, N611, N6100, N1106);
nand NAND4 (N7693, N7689, N4731, N2806, N5446);
and AND4 (N7694, N7688, N4723, N6679, N5313);
nor NOR2 (N7695, N7668, N4504);
xor XOR2 (N7696, N7693, N4730);
or OR3 (N7697, N7687, N4950, N4630);
and AND4 (N7698, N7691, N648, N7431, N1376);
nand NAND3 (N7699, N7690, N6675, N5552);
or OR3 (N7700, N7699, N7509, N2733);
xor XOR2 (N7701, N7698, N6863);
or OR3 (N7702, N7679, N7344, N5571);
not NOT1 (N7703, N7695);
nor NOR4 (N7704, N7697, N6106, N4505, N3238);
and AND2 (N7705, N7704, N5253);
and AND3 (N7706, N7685, N4047, N1108);
nand NAND3 (N7707, N7706, N4659, N1297);
and AND4 (N7708, N7703, N7124, N6870, N2337);
or OR3 (N7709, N7694, N6328, N7428);
not NOT1 (N7710, N7701);
nor NOR2 (N7711, N7692, N7240);
nor NOR4 (N7712, N7707, N1679, N2135, N5471);
xor XOR2 (N7713, N7696, N4917);
xor XOR2 (N7714, N7702, N6568);
not NOT1 (N7715, N7705);
nand NAND2 (N7716, N7700, N3909);
xor XOR2 (N7717, N7716, N2171);
not NOT1 (N7718, N7717);
and AND4 (N7719, N7715, N3031, N1534, N2034);
or OR3 (N7720, N7718, N6617, N4567);
nand NAND3 (N7721, N7686, N3805, N1229);
and AND3 (N7722, N7720, N2090, N2476);
buf BUF1 (N7723, N7722);
nor NOR2 (N7724, N7712, N3865);
not NOT1 (N7725, N7721);
not NOT1 (N7726, N7711);
nor NOR4 (N7727, N7726, N2405, N6221, N5161);
buf BUF1 (N7728, N7727);
nor NOR2 (N7729, N7709, N5298);
nand NAND4 (N7730, N7714, N3348, N5575, N5219);
nand NAND3 (N7731, N7729, N4965, N1942);
nor NOR4 (N7732, N7723, N1270, N3879, N6693);
and AND2 (N7733, N7719, N7675);
not NOT1 (N7734, N7713);
not NOT1 (N7735, N7730);
buf BUF1 (N7736, N7731);
buf BUF1 (N7737, N7736);
and AND3 (N7738, N7725, N2894, N5279);
nand NAND2 (N7739, N7710, N1287);
xor XOR2 (N7740, N7735, N6516);
and AND2 (N7741, N7738, N4295);
buf BUF1 (N7742, N7728);
not NOT1 (N7743, N7742);
and AND2 (N7744, N7739, N7690);
and AND3 (N7745, N7733, N1247, N2152);
buf BUF1 (N7746, N7732);
not NOT1 (N7747, N7724);
nor NOR3 (N7748, N7734, N3017, N5566);
xor XOR2 (N7749, N7708, N4996);
or OR2 (N7750, N7749, N7510);
nor NOR4 (N7751, N7743, N3513, N6376, N144);
or OR3 (N7752, N7751, N2813, N7535);
buf BUF1 (N7753, N7740);
buf BUF1 (N7754, N7753);
not NOT1 (N7755, N7741);
nand NAND3 (N7756, N7737, N4833, N5100);
buf BUF1 (N7757, N7755);
buf BUF1 (N7758, N7745);
and AND3 (N7759, N7746, N3759, N2863);
or OR2 (N7760, N7754, N4291);
and AND4 (N7761, N7756, N4289, N6313, N2611);
nor NOR4 (N7762, N7752, N6711, N4571, N2537);
or OR3 (N7763, N7757, N6578, N4498);
xor XOR2 (N7764, N7763, N7458);
nor NOR3 (N7765, N7748, N1331, N6376);
not NOT1 (N7766, N7764);
buf BUF1 (N7767, N7747);
not NOT1 (N7768, N7762);
xor XOR2 (N7769, N7760, N6330);
and AND2 (N7770, N7767, N2850);
nor NOR3 (N7771, N7768, N638, N6599);
buf BUF1 (N7772, N7769);
buf BUF1 (N7773, N7750);
xor XOR2 (N7774, N7759, N3409);
buf BUF1 (N7775, N7744);
or OR4 (N7776, N7765, N1859, N773, N5351);
and AND4 (N7777, N7771, N7190, N1439, N4112);
not NOT1 (N7778, N7777);
and AND2 (N7779, N7778, N1943);
nand NAND3 (N7780, N7776, N136, N5533);
xor XOR2 (N7781, N7772, N1470);
xor XOR2 (N7782, N7766, N1936);
nand NAND4 (N7783, N7774, N4136, N5235, N1503);
xor XOR2 (N7784, N7773, N6783);
nand NAND3 (N7785, N7780, N6149, N7153);
nand NAND2 (N7786, N7781, N2077);
not NOT1 (N7787, N7775);
nand NAND2 (N7788, N7785, N4991);
buf BUF1 (N7789, N7783);
or OR4 (N7790, N7770, N5995, N4886, N513);
xor XOR2 (N7791, N7782, N4269);
nor NOR2 (N7792, N7784, N7675);
or OR2 (N7793, N7761, N2032);
or OR4 (N7794, N7788, N5175, N7165, N5641);
not NOT1 (N7795, N7790);
nor NOR4 (N7796, N7786, N7539, N7794, N6992);
xor XOR2 (N7797, N5377, N5176);
xor XOR2 (N7798, N7758, N5177);
not NOT1 (N7799, N7796);
nor NOR3 (N7800, N7799, N996, N5335);
not NOT1 (N7801, N7795);
buf BUF1 (N7802, N7787);
buf BUF1 (N7803, N7789);
buf BUF1 (N7804, N7792);
or OR3 (N7805, N7802, N6705, N5579);
xor XOR2 (N7806, N7803, N6702);
and AND2 (N7807, N7805, N2841);
or OR3 (N7808, N7806, N7229, N1907);
and AND2 (N7809, N7804, N7042);
buf BUF1 (N7810, N7798);
buf BUF1 (N7811, N7808);
or OR4 (N7812, N7811, N749, N1802, N2699);
nor NOR3 (N7813, N7801, N6889, N78);
xor XOR2 (N7814, N7797, N5545);
nor NOR3 (N7815, N7809, N3838, N2753);
nor NOR4 (N7816, N7791, N5731, N2393, N368);
or OR2 (N7817, N7807, N3533);
not NOT1 (N7818, N7813);
and AND4 (N7819, N7817, N7265, N2384, N3054);
not NOT1 (N7820, N7812);
xor XOR2 (N7821, N7818, N7562);
or OR4 (N7822, N7820, N6562, N1828, N3187);
not NOT1 (N7823, N7816);
buf BUF1 (N7824, N7800);
xor XOR2 (N7825, N7814, N4266);
and AND2 (N7826, N7821, N5648);
and AND2 (N7827, N7822, N2223);
nand NAND3 (N7828, N7815, N2469, N4994);
or OR4 (N7829, N7779, N5328, N3668, N7410);
xor XOR2 (N7830, N7810, N5025);
xor XOR2 (N7831, N7828, N299);
not NOT1 (N7832, N7824);
nand NAND3 (N7833, N7830, N298, N4734);
nand NAND2 (N7834, N7823, N6174);
buf BUF1 (N7835, N7834);
and AND3 (N7836, N7832, N224, N5720);
not NOT1 (N7837, N7829);
and AND2 (N7838, N7826, N4253);
and AND4 (N7839, N7837, N4955, N5344, N6139);
nand NAND2 (N7840, N7835, N5898);
not NOT1 (N7841, N7793);
buf BUF1 (N7842, N7836);
xor XOR2 (N7843, N7841, N6401);
xor XOR2 (N7844, N7840, N664);
nand NAND4 (N7845, N7825, N2736, N4197, N7231);
and AND4 (N7846, N7839, N2792, N5089, N505);
and AND2 (N7847, N7844, N4415);
or OR2 (N7848, N7846, N5121);
and AND4 (N7849, N7847, N6421, N86, N7521);
nand NAND2 (N7850, N7848, N6451);
xor XOR2 (N7851, N7842, N4092);
or OR4 (N7852, N7819, N129, N4970, N1247);
and AND4 (N7853, N7843, N6507, N5893, N5949);
nor NOR2 (N7854, N7831, N2553);
not NOT1 (N7855, N7852);
and AND3 (N7856, N7845, N4804, N1189);
and AND3 (N7857, N7850, N3887, N3487);
buf BUF1 (N7858, N7833);
not NOT1 (N7859, N7849);
buf BUF1 (N7860, N7855);
nor NOR3 (N7861, N7853, N3878, N7809);
nor NOR2 (N7862, N7827, N4506);
xor XOR2 (N7863, N7838, N7533);
buf BUF1 (N7864, N7857);
not NOT1 (N7865, N7859);
buf BUF1 (N7866, N7864);
not NOT1 (N7867, N7866);
nor NOR3 (N7868, N7851, N3749, N2239);
not NOT1 (N7869, N7861);
and AND3 (N7870, N7863, N2328, N4069);
nor NOR3 (N7871, N7856, N5193, N4408);
or OR4 (N7872, N7868, N1597, N6190, N4310);
or OR4 (N7873, N7854, N983, N1666, N7682);
and AND2 (N7874, N7873, N1584);
nor NOR4 (N7875, N7871, N5792, N3697, N3295);
not NOT1 (N7876, N7865);
and AND4 (N7877, N7872, N7819, N4559, N4109);
buf BUF1 (N7878, N7862);
nor NOR4 (N7879, N7870, N3207, N5475, N2227);
buf BUF1 (N7880, N7860);
nor NOR3 (N7881, N7874, N3593, N5719);
and AND4 (N7882, N7875, N2055, N5768, N1152);
and AND3 (N7883, N7882, N5963, N4739);
not NOT1 (N7884, N7876);
buf BUF1 (N7885, N7878);
nand NAND3 (N7886, N7877, N4184, N6815);
nand NAND4 (N7887, N7884, N600, N1793, N3737);
nor NOR3 (N7888, N7881, N2771, N2733);
nor NOR2 (N7889, N7879, N3072);
and AND4 (N7890, N7885, N385, N2972, N296);
nand NAND2 (N7891, N7887, N4541);
nand NAND2 (N7892, N7883, N6900);
or OR4 (N7893, N7886, N2364, N860, N3163);
and AND3 (N7894, N7867, N2958, N1332);
nand NAND4 (N7895, N7893, N6825, N7078, N3726);
nor NOR3 (N7896, N7892, N3935, N4285);
nor NOR4 (N7897, N7895, N4886, N6151, N338);
xor XOR2 (N7898, N7894, N7199);
nand NAND3 (N7899, N7891, N2939, N2750);
xor XOR2 (N7900, N7888, N844);
xor XOR2 (N7901, N7869, N345);
and AND3 (N7902, N7880, N332, N3607);
xor XOR2 (N7903, N7897, N7105);
or OR3 (N7904, N7900, N3830, N6903);
and AND2 (N7905, N7889, N6507);
or OR4 (N7906, N7903, N3998, N904, N4579);
nor NOR2 (N7907, N7905, N3446);
buf BUF1 (N7908, N7904);
buf BUF1 (N7909, N7858);
xor XOR2 (N7910, N7907, N943);
buf BUF1 (N7911, N7898);
nor NOR3 (N7912, N7909, N6112, N5166);
not NOT1 (N7913, N7902);
and AND2 (N7914, N7910, N7415);
or OR4 (N7915, N7912, N4709, N6633, N2057);
or OR2 (N7916, N7906, N5969);
nand NAND4 (N7917, N7908, N4242, N5341, N7903);
nor NOR3 (N7918, N7917, N6298, N1594);
xor XOR2 (N7919, N7890, N4806);
nand NAND4 (N7920, N7918, N2678, N1452, N4096);
nand NAND2 (N7921, N7913, N3964);
xor XOR2 (N7922, N7899, N1103);
and AND4 (N7923, N7922, N1411, N6234, N7221);
not NOT1 (N7924, N7920);
xor XOR2 (N7925, N7919, N4332);
buf BUF1 (N7926, N7896);
and AND2 (N7927, N7914, N6829);
or OR3 (N7928, N7915, N5212, N6273);
xor XOR2 (N7929, N7928, N797);
xor XOR2 (N7930, N7926, N5361);
xor XOR2 (N7931, N7927, N2216);
nor NOR3 (N7932, N7901, N2777, N800);
or OR2 (N7933, N7932, N2435);
nand NAND3 (N7934, N7923, N3111, N28);
nor NOR3 (N7935, N7934, N4699, N1684);
xor XOR2 (N7936, N7921, N7379);
or OR2 (N7937, N7924, N6653);
buf BUF1 (N7938, N7937);
and AND4 (N7939, N7931, N4263, N2619, N4311);
and AND4 (N7940, N7916, N4618, N2199, N4781);
nor NOR3 (N7941, N7933, N3781, N4003);
not NOT1 (N7942, N7929);
or OR4 (N7943, N7935, N3476, N2902, N3099);
nor NOR3 (N7944, N7930, N6890, N7088);
and AND2 (N7945, N7911, N1637);
buf BUF1 (N7946, N7925);
buf BUF1 (N7947, N7945);
nand NAND4 (N7948, N7939, N1076, N538, N3562);
xor XOR2 (N7949, N7941, N6470);
or OR4 (N7950, N7948, N1087, N3680, N3124);
xor XOR2 (N7951, N7949, N1022);
nor NOR3 (N7952, N7951, N7261, N1869);
or OR3 (N7953, N7946, N6127, N4778);
buf BUF1 (N7954, N7950);
xor XOR2 (N7955, N7952, N6816);
nor NOR4 (N7956, N7942, N1331, N515, N4808);
or OR4 (N7957, N7944, N4176, N3644, N106);
nor NOR2 (N7958, N7955, N6190);
nand NAND4 (N7959, N7940, N4142, N2357, N3511);
nand NAND2 (N7960, N7936, N1754);
or OR4 (N7961, N7953, N1338, N2938, N7151);
or OR4 (N7962, N7960, N1082, N3895, N5324);
buf BUF1 (N7963, N7959);
nand NAND3 (N7964, N7938, N936, N5014);
not NOT1 (N7965, N7957);
xor XOR2 (N7966, N7943, N5855);
xor XOR2 (N7967, N7956, N4262);
nand NAND2 (N7968, N7947, N101);
xor XOR2 (N7969, N7967, N387);
buf BUF1 (N7970, N7954);
nor NOR2 (N7971, N7958, N79);
buf BUF1 (N7972, N7968);
and AND4 (N7973, N7971, N2387, N7024, N4690);
not NOT1 (N7974, N7973);
nor NOR3 (N7975, N7961, N3946, N7613);
and AND3 (N7976, N7974, N1744, N4412);
and AND3 (N7977, N7970, N2536, N6877);
nor NOR4 (N7978, N7975, N6099, N5746, N49);
nand NAND4 (N7979, N7965, N6792, N6386, N3074);
not NOT1 (N7980, N7976);
buf BUF1 (N7981, N7966);
or OR3 (N7982, N7972, N6262, N5550);
not NOT1 (N7983, N7977);
xor XOR2 (N7984, N7982, N4218);
or OR3 (N7985, N7962, N4957, N6424);
not NOT1 (N7986, N7985);
or OR2 (N7987, N7986, N279);
nand NAND2 (N7988, N7981, N314);
nor NOR4 (N7989, N7980, N1664, N186, N6743);
and AND2 (N7990, N7984, N2659);
nor NOR2 (N7991, N7983, N7759);
nand NAND3 (N7992, N7964, N4680, N6405);
buf BUF1 (N7993, N7991);
and AND3 (N7994, N7969, N7887, N4043);
or OR3 (N7995, N7979, N6209, N497);
nand NAND2 (N7996, N7992, N1424);
not NOT1 (N7997, N7987);
and AND2 (N7998, N7990, N3275);
nor NOR4 (N7999, N7988, N5331, N6909, N395);
buf BUF1 (N8000, N7998);
and AND2 (N8001, N7978, N3322);
not NOT1 (N8002, N8001);
or OR4 (N8003, N7994, N2595, N1445, N2672);
buf BUF1 (N8004, N7995);
not NOT1 (N8005, N8004);
or OR2 (N8006, N7989, N7825);
not NOT1 (N8007, N8000);
or OR3 (N8008, N7997, N6107, N4800);
or OR2 (N8009, N8003, N5965);
and AND3 (N8010, N8009, N1911, N6945);
or OR3 (N8011, N7996, N6853, N7362);
not NOT1 (N8012, N7993);
nand NAND3 (N8013, N7999, N3962, N2777);
nor NOR2 (N8014, N8006, N535);
and AND2 (N8015, N8012, N2724);
nor NOR3 (N8016, N8007, N6026, N7131);
nand NAND2 (N8017, N8011, N4333);
nor NOR2 (N8018, N8005, N4950);
nand NAND3 (N8019, N8013, N3586, N3803);
or OR2 (N8020, N8019, N624);
nor NOR3 (N8021, N8018, N705, N7001);
and AND2 (N8022, N8016, N2881);
nor NOR4 (N8023, N8022, N1200, N4912, N4516);
endmodule