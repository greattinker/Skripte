// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13;

output N15995,N15991,N16012,N16000,N16011,N16009,N16006,N15974,N16010,N16013;

buf BUF1 (N14, N3);
buf BUF1 (N15, N4);
nor NOR4 (N16, N13, N6, N5, N7);
nor NOR4 (N17, N14, N4, N15, N11);
or OR2 (N18, N7, N6);
or OR4 (N19, N9, N17, N6, N9);
nor NOR4 (N20, N10, N7, N3, N18);
and AND3 (N21, N17, N18, N20);
nand NAND4 (N22, N11, N12, N16, N20);
nor NOR4 (N23, N10, N16, N20, N12);
buf BUF1 (N24, N23);
nand NAND4 (N25, N4, N10, N6, N18);
and AND2 (N26, N6, N4);
and AND3 (N27, N19, N12, N16);
not NOT1 (N28, N3);
xor XOR2 (N29, N25, N6);
nor NOR3 (N30, N19, N9, N17);
nand NAND2 (N31, N12, N11);
nand NAND3 (N32, N3, N12, N29);
nor NOR4 (N33, N19, N21, N11, N12);
and AND2 (N34, N1, N10);
and AND4 (N35, N22, N6, N9, N9);
and AND3 (N36, N26, N10, N25);
nor NOR3 (N37, N33, N27, N28);
and AND3 (N38, N34, N30, N12);
and AND2 (N39, N29, N38);
not NOT1 (N40, N11);
buf BUF1 (N41, N30);
buf BUF1 (N42, N36);
and AND3 (N43, N7, N39, N14);
not NOT1 (N44, N13);
not NOT1 (N45, N35);
nand NAND4 (N46, N45, N5, N42, N33);
not NOT1 (N47, N8);
or OR2 (N48, N47, N3);
buf BUF1 (N49, N44);
buf BUF1 (N50, N24);
nor NOR3 (N51, N31, N7, N35);
and AND2 (N52, N41, N40);
or OR4 (N53, N17, N10, N24, N17);
and AND4 (N54, N53, N3, N17, N12);
and AND4 (N55, N43, N14, N14, N27);
or OR2 (N56, N52, N47);
not NOT1 (N57, N32);
xor XOR2 (N58, N57, N17);
xor XOR2 (N59, N50, N53);
or OR4 (N60, N54, N53, N42, N39);
nand NAND2 (N61, N37, N60);
buf BUF1 (N62, N43);
nand NAND2 (N63, N48, N21);
xor XOR2 (N64, N56, N40);
nand NAND4 (N65, N55, N7, N1, N6);
not NOT1 (N66, N61);
or OR4 (N67, N63, N57, N3, N6);
xor XOR2 (N68, N62, N11);
buf BUF1 (N69, N65);
nor NOR4 (N70, N69, N22, N15, N27);
or OR3 (N71, N49, N34, N21);
nor NOR4 (N72, N59, N45, N54, N40);
not NOT1 (N73, N71);
nor NOR2 (N74, N70, N60);
buf BUF1 (N75, N73);
and AND2 (N76, N46, N44);
not NOT1 (N77, N68);
or OR2 (N78, N67, N66);
buf BUF1 (N79, N6);
or OR4 (N80, N75, N50, N7, N10);
not NOT1 (N81, N64);
not NOT1 (N82, N74);
xor XOR2 (N83, N79, N81);
nor NOR4 (N84, N35, N63, N35, N82);
or OR4 (N85, N56, N20, N71, N54);
nor NOR4 (N86, N78, N25, N70, N25);
and AND4 (N87, N80, N75, N2, N43);
xor XOR2 (N88, N51, N57);
and AND4 (N89, N85, N43, N80, N3);
nor NOR4 (N90, N77, N89, N18, N85);
nand NAND4 (N91, N10, N11, N36, N2);
or OR2 (N92, N87, N25);
or OR2 (N93, N76, N89);
xor XOR2 (N94, N93, N71);
xor XOR2 (N95, N88, N84);
nand NAND2 (N96, N58, N18);
and AND3 (N97, N87, N91, N18);
or OR2 (N98, N47, N46);
nor NOR2 (N99, N95, N64);
or OR2 (N100, N90, N97);
nand NAND4 (N101, N77, N7, N73, N15);
nand NAND3 (N102, N83, N27, N30);
buf BUF1 (N103, N92);
xor XOR2 (N104, N102, N80);
buf BUF1 (N105, N103);
or OR3 (N106, N105, N33, N15);
or OR4 (N107, N99, N106, N67, N79);
xor XOR2 (N108, N32, N9);
nor NOR2 (N109, N86, N71);
nand NAND2 (N110, N108, N67);
and AND2 (N111, N104, N80);
nor NOR3 (N112, N96, N92, N108);
or OR2 (N113, N100, N36);
not NOT1 (N114, N72);
xor XOR2 (N115, N101, N53);
or OR3 (N116, N110, N12, N12);
and AND4 (N117, N94, N105, N71, N35);
nor NOR4 (N118, N114, N57, N81, N2);
and AND4 (N119, N115, N19, N66, N10);
not NOT1 (N120, N111);
and AND4 (N121, N117, N78, N34, N29);
or OR3 (N122, N116, N7, N10);
and AND3 (N123, N112, N7, N114);
buf BUF1 (N124, N118);
buf BUF1 (N125, N119);
not NOT1 (N126, N120);
buf BUF1 (N127, N107);
nor NOR4 (N128, N121, N111, N20, N109);
buf BUF1 (N129, N67);
nand NAND3 (N130, N98, N129, N79);
not NOT1 (N131, N28);
xor XOR2 (N132, N123, N104);
not NOT1 (N133, N113);
and AND3 (N134, N130, N44, N10);
and AND4 (N135, N127, N125, N115, N26);
not NOT1 (N136, N94);
xor XOR2 (N137, N131, N7);
buf BUF1 (N138, N126);
not NOT1 (N139, N138);
nor NOR3 (N140, N124, N90, N99);
nor NOR2 (N141, N128, N83);
xor XOR2 (N142, N134, N23);
buf BUF1 (N143, N136);
or OR2 (N144, N122, N125);
and AND4 (N145, N144, N132, N80, N111);
nand NAND3 (N146, N20, N118, N51);
and AND4 (N147, N142, N18, N19, N131);
nor NOR3 (N148, N147, N94, N140);
buf BUF1 (N149, N144);
or OR4 (N150, N143, N77, N149, N44);
or OR2 (N151, N93, N82);
not NOT1 (N152, N133);
or OR3 (N153, N151, N88, N147);
nor NOR4 (N154, N148, N81, N105, N83);
buf BUF1 (N155, N152);
or OR2 (N156, N150, N109);
buf BUF1 (N157, N146);
not NOT1 (N158, N135);
xor XOR2 (N159, N141, N89);
nand NAND3 (N160, N153, N16, N98);
not NOT1 (N161, N145);
nor NOR3 (N162, N154, N74, N37);
nor NOR4 (N163, N137, N147, N112, N67);
and AND4 (N164, N155, N25, N11, N101);
xor XOR2 (N165, N157, N145);
nor NOR4 (N166, N139, N37, N101, N38);
buf BUF1 (N167, N164);
buf BUF1 (N168, N162);
and AND3 (N169, N156, N65, N150);
or OR3 (N170, N166, N51, N55);
nor NOR4 (N171, N158, N21, N27, N94);
nor NOR2 (N172, N171, N142);
xor XOR2 (N173, N167, N6);
and AND3 (N174, N159, N57, N36);
xor XOR2 (N175, N160, N102);
buf BUF1 (N176, N175);
or OR3 (N177, N176, N31, N99);
and AND2 (N178, N161, N152);
xor XOR2 (N179, N169, N173);
nor NOR4 (N180, N62, N150, N13, N20);
xor XOR2 (N181, N163, N35);
not NOT1 (N182, N177);
buf BUF1 (N183, N178);
or OR3 (N184, N168, N118, N74);
nor NOR4 (N185, N172, N44, N153, N16);
nand NAND2 (N186, N184, N23);
or OR3 (N187, N181, N79, N9);
and AND4 (N188, N180, N169, N90, N28);
nand NAND4 (N189, N186, N51, N47, N40);
and AND2 (N190, N179, N75);
nand NAND2 (N191, N188, N147);
not NOT1 (N192, N183);
xor XOR2 (N193, N170, N53);
buf BUF1 (N194, N182);
buf BUF1 (N195, N185);
buf BUF1 (N196, N194);
buf BUF1 (N197, N165);
not NOT1 (N198, N195);
nand NAND4 (N199, N174, N127, N193, N26);
nor NOR4 (N200, N123, N165, N29, N29);
buf BUF1 (N201, N189);
and AND2 (N202, N200, N134);
not NOT1 (N203, N201);
or OR3 (N204, N191, N61, N23);
nand NAND2 (N205, N199, N15);
buf BUF1 (N206, N205);
or OR3 (N207, N192, N141, N56);
buf BUF1 (N208, N198);
xor XOR2 (N209, N197, N138);
xor XOR2 (N210, N209, N160);
nand NAND4 (N211, N208, N72, N206, N21);
or OR2 (N212, N64, N122);
nand NAND4 (N213, N196, N154, N94, N4);
nand NAND3 (N214, N211, N112, N126);
nand NAND4 (N215, N187, N134, N147, N93);
nor NOR2 (N216, N190, N186);
buf BUF1 (N217, N213);
xor XOR2 (N218, N210, N216);
and AND4 (N219, N176, N34, N38, N57);
buf BUF1 (N220, N207);
not NOT1 (N221, N220);
nor NOR4 (N222, N218, N52, N167, N202);
xor XOR2 (N223, N166, N206);
not NOT1 (N224, N203);
nor NOR2 (N225, N222, N81);
xor XOR2 (N226, N224, N124);
not NOT1 (N227, N223);
buf BUF1 (N228, N225);
nor NOR4 (N229, N228, N205, N78, N190);
xor XOR2 (N230, N204, N192);
nor NOR3 (N231, N214, N186, N80);
nand NAND3 (N232, N221, N84, N212);
xor XOR2 (N233, N98, N72);
nor NOR4 (N234, N232, N212, N192, N25);
xor XOR2 (N235, N217, N79);
nor NOR2 (N236, N230, N155);
nor NOR3 (N237, N233, N175, N205);
xor XOR2 (N238, N226, N78);
xor XOR2 (N239, N234, N115);
nor NOR3 (N240, N215, N201, N137);
buf BUF1 (N241, N236);
xor XOR2 (N242, N227, N213);
and AND2 (N243, N241, N110);
nor NOR4 (N244, N231, N136, N139, N190);
xor XOR2 (N245, N242, N183);
and AND2 (N246, N244, N174);
or OR3 (N247, N245, N3, N17);
and AND2 (N248, N238, N221);
nor NOR3 (N249, N229, N237, N120);
or OR3 (N250, N11, N146, N117);
buf BUF1 (N251, N219);
or OR4 (N252, N235, N61, N178, N90);
xor XOR2 (N253, N247, N146);
or OR3 (N254, N248, N236, N35);
or OR4 (N255, N249, N61, N236, N86);
not NOT1 (N256, N246);
nand NAND3 (N257, N252, N173, N188);
not NOT1 (N258, N240);
nand NAND3 (N259, N253, N194, N164);
and AND2 (N260, N243, N255);
not NOT1 (N261, N177);
and AND3 (N262, N254, N46, N1);
or OR4 (N263, N259, N171, N116, N133);
not NOT1 (N264, N261);
not NOT1 (N265, N260);
xor XOR2 (N266, N263, N176);
buf BUF1 (N267, N251);
and AND3 (N268, N262, N232, N119);
nor NOR4 (N269, N264, N198, N263, N217);
and AND2 (N270, N256, N142);
and AND3 (N271, N265, N126, N181);
buf BUF1 (N272, N267);
nand NAND3 (N273, N250, N171, N47);
nand NAND3 (N274, N258, N138, N45);
and AND3 (N275, N257, N259, N68);
xor XOR2 (N276, N271, N41);
or OR3 (N277, N269, N184, N152);
not NOT1 (N278, N277);
xor XOR2 (N279, N273, N121);
nor NOR2 (N280, N270, N231);
xor XOR2 (N281, N239, N27);
or OR4 (N282, N266, N115, N171, N254);
nor NOR4 (N283, N279, N281, N51, N255);
or OR4 (N284, N223, N96, N45, N137);
nor NOR2 (N285, N276, N87);
xor XOR2 (N286, N275, N52);
or OR2 (N287, N278, N284);
or OR2 (N288, N19, N175);
or OR3 (N289, N274, N7, N44);
buf BUF1 (N290, N289);
not NOT1 (N291, N282);
buf BUF1 (N292, N285);
nand NAND3 (N293, N287, N114, N223);
nand NAND3 (N294, N283, N98, N185);
or OR3 (N295, N292, N55, N50);
buf BUF1 (N296, N268);
and AND4 (N297, N296, N3, N73, N220);
not NOT1 (N298, N280);
nor NOR3 (N299, N294, N137, N280);
nand NAND4 (N300, N295, N24, N119, N28);
nor NOR4 (N301, N286, N20, N40, N72);
not NOT1 (N302, N301);
nand NAND3 (N303, N300, N190, N127);
not NOT1 (N304, N293);
buf BUF1 (N305, N291);
xor XOR2 (N306, N298, N67);
nor NOR2 (N307, N302, N270);
nor NOR4 (N308, N305, N234, N4, N207);
and AND2 (N309, N299, N230);
nand NAND2 (N310, N288, N90);
nor NOR2 (N311, N304, N31);
xor XOR2 (N312, N290, N162);
nor NOR4 (N313, N306, N158, N176, N22);
nor NOR2 (N314, N311, N244);
nand NAND3 (N315, N314, N191, N242);
buf BUF1 (N316, N297);
nor NOR2 (N317, N307, N276);
xor XOR2 (N318, N317, N1);
or OR3 (N319, N309, N270, N302);
or OR3 (N320, N308, N28, N307);
nand NAND4 (N321, N315, N87, N186, N221);
nor NOR4 (N322, N321, N203, N16, N134);
and AND4 (N323, N322, N58, N269, N49);
buf BUF1 (N324, N320);
buf BUF1 (N325, N318);
or OR3 (N326, N272, N273, N269);
nor NOR2 (N327, N325, N321);
or OR2 (N328, N310, N45);
and AND2 (N329, N327, N111);
nand NAND4 (N330, N319, N295, N205, N297);
xor XOR2 (N331, N316, N77);
not NOT1 (N332, N313);
nand NAND4 (N333, N312, N160, N243, N327);
and AND4 (N334, N328, N314, N67, N297);
nor NOR2 (N335, N331, N87);
xor XOR2 (N336, N330, N45);
xor XOR2 (N337, N333, N135);
xor XOR2 (N338, N335, N159);
and AND3 (N339, N303, N125, N159);
xor XOR2 (N340, N332, N222);
nand NAND3 (N341, N324, N53, N131);
or OR4 (N342, N336, N296, N102, N72);
nor NOR4 (N343, N323, N207, N142, N234);
or OR3 (N344, N339, N30, N246);
nand NAND2 (N345, N341, N60);
and AND4 (N346, N338, N328, N207, N315);
xor XOR2 (N347, N334, N156);
or OR2 (N348, N346, N7);
buf BUF1 (N349, N343);
and AND2 (N350, N340, N269);
nand NAND3 (N351, N342, N345, N161);
nor NOR4 (N352, N262, N94, N7, N64);
xor XOR2 (N353, N347, N292);
nor NOR2 (N354, N350, N260);
xor XOR2 (N355, N349, N91);
not NOT1 (N356, N354);
not NOT1 (N357, N348);
xor XOR2 (N358, N344, N357);
and AND3 (N359, N342, N95, N267);
buf BUF1 (N360, N337);
xor XOR2 (N361, N329, N49);
buf BUF1 (N362, N326);
xor XOR2 (N363, N356, N18);
and AND4 (N364, N361, N231, N302, N323);
nor NOR2 (N365, N358, N117);
nor NOR3 (N366, N362, N8, N165);
nor NOR4 (N367, N366, N169, N71, N348);
nor NOR4 (N368, N360, N110, N221, N194);
buf BUF1 (N369, N364);
or OR4 (N370, N351, N258, N188, N361);
buf BUF1 (N371, N359);
buf BUF1 (N372, N353);
nand NAND4 (N373, N352, N289, N247, N71);
nor NOR4 (N374, N355, N227, N30, N147);
buf BUF1 (N375, N369);
nand NAND4 (N376, N368, N137, N183, N271);
not NOT1 (N377, N370);
nor NOR3 (N378, N371, N217, N338);
not NOT1 (N379, N377);
nor NOR2 (N380, N374, N214);
nand NAND3 (N381, N375, N338, N45);
buf BUF1 (N382, N363);
nand NAND2 (N383, N372, N164);
buf BUF1 (N384, N378);
or OR3 (N385, N380, N65, N11);
xor XOR2 (N386, N383, N54);
or OR3 (N387, N373, N192, N98);
xor XOR2 (N388, N384, N301);
buf BUF1 (N389, N367);
nor NOR2 (N390, N388, N237);
xor XOR2 (N391, N389, N19);
and AND2 (N392, N376, N140);
buf BUF1 (N393, N390);
xor XOR2 (N394, N365, N33);
nor NOR3 (N395, N393, N327, N80);
or OR2 (N396, N392, N383);
nor NOR4 (N397, N396, N199, N105, N185);
or OR2 (N398, N381, N57);
and AND3 (N399, N394, N277, N47);
nor NOR4 (N400, N397, N287, N143, N181);
nand NAND4 (N401, N395, N82, N63, N180);
xor XOR2 (N402, N401, N157);
nor NOR4 (N403, N382, N299, N81, N248);
nor NOR4 (N404, N387, N228, N96, N365);
nor NOR4 (N405, N404, N320, N140, N53);
not NOT1 (N406, N399);
not NOT1 (N407, N379);
or OR4 (N408, N402, N293, N332, N37);
not NOT1 (N409, N403);
nand NAND4 (N410, N400, N84, N409, N104);
buf BUF1 (N411, N392);
nand NAND2 (N412, N398, N167);
and AND2 (N413, N412, N196);
buf BUF1 (N414, N408);
xor XOR2 (N415, N386, N115);
nand NAND3 (N416, N385, N283, N151);
nand NAND4 (N417, N405, N255, N38, N27);
not NOT1 (N418, N415);
nor NOR3 (N419, N413, N46, N242);
xor XOR2 (N420, N419, N393);
and AND2 (N421, N420, N261);
buf BUF1 (N422, N391);
not NOT1 (N423, N410);
or OR2 (N424, N417, N312);
and AND2 (N425, N414, N160);
not NOT1 (N426, N422);
not NOT1 (N427, N426);
nor NOR3 (N428, N423, N240, N318);
and AND3 (N429, N407, N170, N287);
xor XOR2 (N430, N418, N298);
nor NOR2 (N431, N427, N34);
and AND2 (N432, N428, N32);
nor NOR2 (N433, N416, N216);
nand NAND2 (N434, N431, N6);
nor NOR3 (N435, N424, N322, N135);
not NOT1 (N436, N406);
nor NOR3 (N437, N435, N271, N101);
nor NOR4 (N438, N411, N124, N102, N334);
nand NAND4 (N439, N425, N349, N296, N241);
not NOT1 (N440, N433);
buf BUF1 (N441, N429);
nor NOR3 (N442, N440, N317, N345);
or OR3 (N443, N442, N279, N356);
not NOT1 (N444, N430);
and AND3 (N445, N438, N29, N189);
buf BUF1 (N446, N444);
nand NAND4 (N447, N421, N328, N318, N167);
and AND3 (N448, N441, N128, N340);
and AND4 (N449, N445, N220, N379, N23);
or OR2 (N450, N447, N129);
or OR3 (N451, N432, N309, N284);
and AND3 (N452, N437, N46, N61);
nor NOR3 (N453, N451, N419, N395);
not NOT1 (N454, N443);
nand NAND4 (N455, N453, N283, N252, N376);
nand NAND4 (N456, N455, N116, N232, N203);
nand NAND4 (N457, N434, N447, N354, N243);
nor NOR4 (N458, N457, N190, N89, N177);
or OR2 (N459, N456, N276);
or OR4 (N460, N439, N132, N26, N435);
nand NAND4 (N461, N452, N300, N56, N275);
not NOT1 (N462, N446);
not NOT1 (N463, N448);
buf BUF1 (N464, N454);
nand NAND3 (N465, N458, N92, N380);
or OR3 (N466, N462, N219, N206);
and AND4 (N467, N460, N274, N152, N192);
xor XOR2 (N468, N467, N373);
or OR4 (N469, N463, N164, N7, N413);
and AND3 (N470, N449, N156, N194);
and AND3 (N471, N450, N98, N378);
and AND3 (N472, N471, N447, N213);
nand NAND3 (N473, N461, N22, N342);
and AND4 (N474, N469, N13, N3, N206);
nor NOR2 (N475, N464, N283);
and AND2 (N476, N473, N368);
or OR2 (N477, N468, N273);
xor XOR2 (N478, N470, N231);
nor NOR4 (N479, N459, N336, N41, N305);
xor XOR2 (N480, N478, N468);
nor NOR4 (N481, N474, N139, N274, N101);
and AND4 (N482, N466, N156, N328, N373);
not NOT1 (N483, N475);
nand NAND4 (N484, N482, N324, N469, N312);
nand NAND4 (N485, N481, N397, N266, N10);
or OR2 (N486, N479, N258);
not NOT1 (N487, N436);
and AND3 (N488, N483, N38, N319);
xor XOR2 (N489, N486, N162);
and AND2 (N490, N465, N377);
or OR3 (N491, N477, N255, N407);
xor XOR2 (N492, N484, N4);
and AND4 (N493, N490, N226, N120, N19);
not NOT1 (N494, N493);
nand NAND4 (N495, N492, N79, N237, N348);
not NOT1 (N496, N495);
nor NOR2 (N497, N489, N237);
not NOT1 (N498, N491);
and AND3 (N499, N498, N448, N492);
or OR4 (N500, N499, N179, N69, N481);
buf BUF1 (N501, N494);
and AND3 (N502, N497, N463, N478);
xor XOR2 (N503, N487, N205);
xor XOR2 (N504, N472, N365);
or OR3 (N505, N485, N374, N443);
nand NAND4 (N506, N504, N485, N259, N3);
not NOT1 (N507, N488);
and AND2 (N508, N500, N81);
nor NOR2 (N509, N480, N445);
and AND3 (N510, N502, N279, N44);
or OR4 (N511, N501, N455, N233, N108);
nand NAND2 (N512, N510, N289);
nor NOR4 (N513, N503, N129, N326, N373);
buf BUF1 (N514, N509);
and AND4 (N515, N476, N17, N239, N35);
nor NOR2 (N516, N496, N111);
not NOT1 (N517, N511);
and AND3 (N518, N514, N115, N141);
and AND4 (N519, N515, N145, N424, N56);
nor NOR3 (N520, N516, N2, N69);
not NOT1 (N521, N520);
not NOT1 (N522, N508);
and AND4 (N523, N517, N108, N329, N494);
and AND3 (N524, N523, N422, N227);
buf BUF1 (N525, N513);
not NOT1 (N526, N524);
buf BUF1 (N527, N507);
nor NOR2 (N528, N521, N241);
nor NOR3 (N529, N512, N525, N338);
not NOT1 (N530, N343);
or OR3 (N531, N527, N39, N55);
buf BUF1 (N532, N530);
nand NAND4 (N533, N519, N425, N406, N29);
not NOT1 (N534, N528);
buf BUF1 (N535, N518);
xor XOR2 (N536, N505, N264);
xor XOR2 (N537, N532, N100);
not NOT1 (N538, N536);
not NOT1 (N539, N534);
xor XOR2 (N540, N538, N264);
nand NAND4 (N541, N522, N488, N137, N435);
nor NOR2 (N542, N529, N298);
and AND3 (N543, N526, N540, N276);
or OR3 (N544, N451, N288, N412);
not NOT1 (N545, N539);
and AND3 (N546, N544, N428, N412);
buf BUF1 (N547, N542);
xor XOR2 (N548, N531, N344);
buf BUF1 (N549, N506);
xor XOR2 (N550, N533, N297);
and AND4 (N551, N549, N304, N314, N213);
nor NOR4 (N552, N551, N218, N420, N417);
nand NAND4 (N553, N541, N370, N495, N191);
buf BUF1 (N554, N548);
xor XOR2 (N555, N546, N239);
nor NOR4 (N556, N553, N431, N420, N372);
nor NOR2 (N557, N537, N166);
buf BUF1 (N558, N547);
and AND4 (N559, N554, N119, N33, N447);
and AND2 (N560, N556, N206);
not NOT1 (N561, N545);
buf BUF1 (N562, N560);
not NOT1 (N563, N535);
nand NAND2 (N564, N558, N212);
nor NOR3 (N565, N563, N361, N34);
not NOT1 (N566, N559);
nand NAND3 (N567, N562, N434, N173);
nor NOR3 (N568, N567, N337, N57);
nor NOR2 (N569, N543, N426);
not NOT1 (N570, N564);
xor XOR2 (N571, N552, N262);
not NOT1 (N572, N561);
not NOT1 (N573, N565);
or OR3 (N574, N573, N65, N23);
or OR3 (N575, N555, N146, N117);
nand NAND4 (N576, N572, N464, N402, N529);
not NOT1 (N577, N575);
nand NAND4 (N578, N568, N99, N128, N557);
not NOT1 (N579, N136);
nor NOR2 (N580, N577, N373);
nand NAND2 (N581, N571, N456);
nand NAND4 (N582, N569, N572, N235, N8);
nand NAND4 (N583, N581, N217, N273, N529);
and AND3 (N584, N576, N173, N446);
nand NAND2 (N585, N583, N325);
nand NAND4 (N586, N580, N115, N115, N161);
buf BUF1 (N587, N550);
or OR3 (N588, N570, N218, N208);
not NOT1 (N589, N582);
nor NOR2 (N590, N585, N458);
xor XOR2 (N591, N590, N310);
xor XOR2 (N592, N591, N313);
nor NOR3 (N593, N584, N392, N454);
nor NOR4 (N594, N578, N466, N577, N194);
or OR3 (N595, N589, N429, N94);
nand NAND2 (N596, N594, N63);
or OR2 (N597, N588, N334);
xor XOR2 (N598, N579, N594);
nor NOR2 (N599, N586, N560);
buf BUF1 (N600, N595);
buf BUF1 (N601, N587);
nand NAND4 (N602, N601, N517, N345, N174);
or OR3 (N603, N592, N393, N31);
nand NAND3 (N604, N599, N239, N205);
and AND2 (N605, N600, N363);
buf BUF1 (N606, N605);
and AND4 (N607, N598, N271, N587, N152);
buf BUF1 (N608, N604);
or OR4 (N609, N593, N273, N388, N573);
or OR2 (N610, N596, N349);
nand NAND4 (N611, N610, N440, N278, N262);
buf BUF1 (N612, N611);
or OR3 (N613, N607, N48, N262);
buf BUF1 (N614, N603);
buf BUF1 (N615, N614);
nor NOR3 (N616, N606, N92, N270);
nor NOR4 (N617, N566, N347, N198, N392);
nand NAND2 (N618, N615, N558);
nor NOR4 (N619, N597, N22, N478, N286);
or OR2 (N620, N617, N571);
not NOT1 (N621, N574);
not NOT1 (N622, N612);
not NOT1 (N623, N616);
nor NOR2 (N624, N609, N448);
nand NAND3 (N625, N621, N276, N577);
or OR3 (N626, N608, N435, N401);
and AND3 (N627, N624, N197, N542);
and AND2 (N628, N620, N20);
xor XOR2 (N629, N618, N120);
nand NAND3 (N630, N627, N621, N180);
nand NAND3 (N631, N622, N120, N485);
xor XOR2 (N632, N619, N267);
nor NOR2 (N633, N628, N440);
and AND3 (N634, N629, N375, N471);
and AND2 (N635, N634, N598);
nand NAND2 (N636, N632, N209);
not NOT1 (N637, N613);
and AND3 (N638, N630, N247, N91);
not NOT1 (N639, N631);
and AND3 (N640, N633, N163, N248);
xor XOR2 (N641, N623, N193);
nor NOR4 (N642, N641, N232, N81, N103);
and AND4 (N643, N640, N119, N455, N108);
or OR2 (N644, N635, N132);
xor XOR2 (N645, N602, N603);
buf BUF1 (N646, N642);
and AND2 (N647, N639, N281);
not NOT1 (N648, N625);
or OR2 (N649, N644, N179);
nor NOR3 (N650, N637, N605, N69);
or OR4 (N651, N650, N442, N46, N512);
nor NOR3 (N652, N638, N379, N373);
nor NOR3 (N653, N645, N478, N335);
or OR4 (N654, N652, N141, N533, N178);
nand NAND3 (N655, N651, N165, N643);
nor NOR3 (N656, N233, N483, N89);
nand NAND4 (N657, N647, N246, N44, N631);
nor NOR4 (N658, N646, N80, N229, N234);
nor NOR3 (N659, N656, N443, N441);
nand NAND2 (N660, N653, N194);
and AND2 (N661, N655, N638);
or OR2 (N662, N626, N637);
buf BUF1 (N663, N661);
nand NAND2 (N664, N657, N346);
or OR3 (N665, N654, N381, N567);
not NOT1 (N666, N659);
nand NAND3 (N667, N664, N523, N261);
not NOT1 (N668, N666);
nand NAND2 (N669, N663, N276);
and AND4 (N670, N658, N258, N105, N456);
xor XOR2 (N671, N649, N560);
and AND3 (N672, N662, N247, N447);
and AND2 (N673, N648, N82);
xor XOR2 (N674, N665, N157);
nor NOR2 (N675, N660, N240);
xor XOR2 (N676, N673, N371);
not NOT1 (N677, N674);
and AND2 (N678, N668, N334);
nand NAND4 (N679, N670, N118, N385, N571);
xor XOR2 (N680, N679, N339);
not NOT1 (N681, N680);
xor XOR2 (N682, N672, N98);
buf BUF1 (N683, N636);
nor NOR2 (N684, N681, N249);
xor XOR2 (N685, N669, N603);
and AND2 (N686, N685, N77);
xor XOR2 (N687, N682, N402);
xor XOR2 (N688, N684, N139);
or OR3 (N689, N676, N631, N393);
buf BUF1 (N690, N689);
xor XOR2 (N691, N690, N3);
xor XOR2 (N692, N667, N664);
xor XOR2 (N693, N677, N40);
nand NAND4 (N694, N678, N270, N531, N437);
or OR3 (N695, N675, N288, N683);
not NOT1 (N696, N88);
buf BUF1 (N697, N671);
nor NOR4 (N698, N686, N405, N625, N308);
buf BUF1 (N699, N696);
buf BUF1 (N700, N699);
buf BUF1 (N701, N697);
nand NAND3 (N702, N701, N254, N323);
xor XOR2 (N703, N698, N168);
xor XOR2 (N704, N692, N546);
xor XOR2 (N705, N688, N702);
nor NOR2 (N706, N611, N657);
not NOT1 (N707, N703);
nand NAND3 (N708, N687, N372, N520);
not NOT1 (N709, N708);
nand NAND3 (N710, N691, N274, N477);
or OR3 (N711, N693, N500, N123);
and AND3 (N712, N710, N50, N638);
not NOT1 (N713, N705);
nand NAND2 (N714, N707, N111);
buf BUF1 (N715, N706);
and AND2 (N716, N711, N576);
not NOT1 (N717, N716);
or OR4 (N718, N700, N717, N339, N97);
nor NOR3 (N719, N436, N5, N324);
buf BUF1 (N720, N695);
not NOT1 (N721, N712);
or OR3 (N722, N709, N626, N340);
not NOT1 (N723, N704);
nand NAND2 (N724, N723, N100);
not NOT1 (N725, N715);
nor NOR2 (N726, N720, N11);
nand NAND4 (N727, N719, N161, N551, N355);
not NOT1 (N728, N714);
or OR4 (N729, N713, N472, N539, N133);
nor NOR4 (N730, N728, N675, N668, N186);
buf BUF1 (N731, N722);
or OR4 (N732, N727, N46, N587, N165);
nand NAND3 (N733, N725, N133, N434);
xor XOR2 (N734, N726, N221);
buf BUF1 (N735, N733);
xor XOR2 (N736, N730, N241);
and AND4 (N737, N729, N330, N89, N186);
nor NOR2 (N738, N731, N491);
or OR4 (N739, N736, N481, N301, N152);
nand NAND2 (N740, N738, N15);
or OR4 (N741, N724, N630, N454, N243);
not NOT1 (N742, N718);
and AND2 (N743, N732, N345);
not NOT1 (N744, N694);
buf BUF1 (N745, N742);
or OR2 (N746, N737, N279);
nor NOR4 (N747, N743, N476, N163, N256);
not NOT1 (N748, N747);
nand NAND4 (N749, N741, N159, N536, N229);
nor NOR3 (N750, N744, N741, N295);
nand NAND4 (N751, N745, N53, N493, N28);
nand NAND4 (N752, N735, N222, N235, N194);
xor XOR2 (N753, N721, N702);
or OR2 (N754, N739, N23);
nor NOR3 (N755, N749, N173, N63);
or OR4 (N756, N755, N2, N389, N539);
buf BUF1 (N757, N734);
not NOT1 (N758, N756);
buf BUF1 (N759, N753);
nor NOR4 (N760, N759, N389, N640, N249);
nand NAND2 (N761, N760, N339);
or OR2 (N762, N746, N439);
buf BUF1 (N763, N762);
nand NAND2 (N764, N751, N122);
nor NOR3 (N765, N758, N298, N440);
or OR4 (N766, N761, N145, N422, N379);
buf BUF1 (N767, N748);
not NOT1 (N768, N752);
nor NOR2 (N769, N768, N394);
and AND2 (N770, N766, N750);
buf BUF1 (N771, N623);
and AND4 (N772, N770, N142, N429, N457);
nor NOR2 (N773, N772, N329);
or OR3 (N774, N764, N737, N572);
buf BUF1 (N775, N767);
nand NAND4 (N776, N774, N152, N273, N448);
nand NAND2 (N777, N740, N11);
not NOT1 (N778, N769);
nand NAND3 (N779, N757, N303, N88);
or OR3 (N780, N776, N116, N24);
nand NAND4 (N781, N775, N604, N11, N269);
not NOT1 (N782, N779);
nand NAND4 (N783, N754, N118, N30, N569);
xor XOR2 (N784, N781, N595);
and AND2 (N785, N777, N494);
xor XOR2 (N786, N765, N633);
nand NAND2 (N787, N785, N440);
not NOT1 (N788, N763);
and AND2 (N789, N787, N294);
buf BUF1 (N790, N782);
xor XOR2 (N791, N789, N730);
xor XOR2 (N792, N784, N471);
xor XOR2 (N793, N783, N410);
xor XOR2 (N794, N786, N558);
not NOT1 (N795, N791);
and AND3 (N796, N792, N432, N795);
and AND2 (N797, N284, N544);
buf BUF1 (N798, N796);
nor NOR4 (N799, N771, N608, N93, N23);
nor NOR4 (N800, N778, N644, N94, N323);
and AND2 (N801, N800, N488);
and AND2 (N802, N801, N26);
nor NOR3 (N803, N773, N406, N582);
or OR4 (N804, N798, N399, N238, N760);
or OR2 (N805, N793, N218);
not NOT1 (N806, N803);
and AND4 (N807, N788, N268, N468, N396);
nand NAND3 (N808, N780, N419, N309);
and AND3 (N809, N808, N220, N12);
buf BUF1 (N810, N809);
nor NOR3 (N811, N799, N736, N45);
and AND4 (N812, N797, N489, N26, N802);
xor XOR2 (N813, N245, N659);
or OR4 (N814, N794, N161, N100, N290);
buf BUF1 (N815, N811);
xor XOR2 (N816, N812, N157);
buf BUF1 (N817, N810);
not NOT1 (N818, N804);
buf BUF1 (N819, N807);
not NOT1 (N820, N816);
not NOT1 (N821, N818);
nand NAND4 (N822, N819, N750, N93, N156);
nor NOR4 (N823, N806, N554, N416, N81);
buf BUF1 (N824, N790);
and AND3 (N825, N824, N614, N340);
and AND4 (N826, N813, N317, N464, N177);
and AND4 (N827, N823, N332, N688, N242);
xor XOR2 (N828, N817, N185);
or OR3 (N829, N826, N663, N725);
nand NAND4 (N830, N814, N522, N388, N408);
or OR2 (N831, N815, N125);
nand NAND3 (N832, N830, N46, N767);
or OR3 (N833, N821, N806, N746);
not NOT1 (N834, N827);
buf BUF1 (N835, N805);
not NOT1 (N836, N825);
not NOT1 (N837, N835);
buf BUF1 (N838, N831);
nand NAND3 (N839, N834, N264, N777);
nand NAND4 (N840, N838, N316, N348, N403);
nor NOR3 (N841, N840, N488, N621);
not NOT1 (N842, N839);
and AND3 (N843, N833, N225, N109);
nor NOR3 (N844, N837, N731, N399);
and AND3 (N845, N836, N742, N13);
xor XOR2 (N846, N829, N415);
buf BUF1 (N847, N843);
not NOT1 (N848, N844);
nand NAND3 (N849, N848, N314, N338);
or OR2 (N850, N847, N630);
xor XOR2 (N851, N841, N588);
or OR2 (N852, N846, N321);
nor NOR2 (N853, N852, N682);
buf BUF1 (N854, N842);
and AND2 (N855, N851, N204);
or OR4 (N856, N828, N479, N847, N35);
buf BUF1 (N857, N854);
nand NAND4 (N858, N853, N131, N273, N224);
not NOT1 (N859, N850);
nor NOR3 (N860, N855, N487, N198);
nor NOR4 (N861, N820, N836, N848, N57);
or OR4 (N862, N849, N306, N278, N232);
not NOT1 (N863, N859);
and AND3 (N864, N858, N860, N732);
xor XOR2 (N865, N277, N102);
nor NOR3 (N866, N857, N721, N146);
buf BUF1 (N867, N866);
xor XOR2 (N868, N845, N613);
not NOT1 (N869, N867);
and AND2 (N870, N868, N133);
buf BUF1 (N871, N862);
xor XOR2 (N872, N864, N159);
and AND4 (N873, N832, N418, N127, N654);
xor XOR2 (N874, N861, N730);
nor NOR4 (N875, N871, N508, N334, N671);
nor NOR4 (N876, N875, N123, N443, N570);
or OR3 (N877, N872, N742, N550);
and AND3 (N878, N870, N589, N702);
or OR3 (N879, N878, N846, N406);
or OR2 (N880, N876, N251);
xor XOR2 (N881, N874, N357);
nand NAND4 (N882, N877, N548, N17, N790);
not NOT1 (N883, N882);
not NOT1 (N884, N873);
xor XOR2 (N885, N880, N140);
not NOT1 (N886, N863);
buf BUF1 (N887, N856);
buf BUF1 (N888, N885);
or OR4 (N889, N888, N341, N834, N485);
buf BUF1 (N890, N889);
and AND4 (N891, N890, N275, N361, N6);
buf BUF1 (N892, N891);
and AND2 (N893, N881, N204);
and AND2 (N894, N886, N454);
xor XOR2 (N895, N894, N156);
nor NOR2 (N896, N869, N136);
xor XOR2 (N897, N865, N687);
not NOT1 (N898, N879);
xor XOR2 (N899, N887, N301);
xor XOR2 (N900, N896, N645);
nor NOR4 (N901, N883, N520, N32, N883);
nand NAND2 (N902, N899, N717);
and AND3 (N903, N901, N501, N8);
not NOT1 (N904, N903);
not NOT1 (N905, N897);
nand NAND2 (N906, N900, N255);
buf BUF1 (N907, N906);
not NOT1 (N908, N904);
buf BUF1 (N909, N905);
or OR3 (N910, N893, N665, N721);
xor XOR2 (N911, N908, N566);
xor XOR2 (N912, N898, N744);
and AND2 (N913, N895, N711);
not NOT1 (N914, N911);
or OR4 (N915, N914, N619, N658, N642);
buf BUF1 (N916, N892);
nor NOR3 (N917, N916, N694, N378);
nor NOR3 (N918, N917, N302, N104);
nor NOR2 (N919, N884, N392);
buf BUF1 (N920, N915);
nand NAND4 (N921, N919, N574, N829, N354);
buf BUF1 (N922, N913);
not NOT1 (N923, N912);
and AND2 (N924, N923, N509);
buf BUF1 (N925, N918);
and AND2 (N926, N921, N249);
not NOT1 (N927, N926);
or OR2 (N928, N925, N494);
nor NOR2 (N929, N920, N535);
and AND4 (N930, N929, N489, N739, N921);
nor NOR4 (N931, N907, N781, N361, N882);
xor XOR2 (N932, N924, N96);
nor NOR2 (N933, N922, N125);
nand NAND3 (N934, N902, N618, N397);
and AND3 (N935, N930, N461, N670);
xor XOR2 (N936, N933, N412);
buf BUF1 (N937, N910);
buf BUF1 (N938, N928);
nand NAND3 (N939, N931, N403, N171);
xor XOR2 (N940, N936, N308);
buf BUF1 (N941, N932);
not NOT1 (N942, N934);
or OR3 (N943, N938, N643, N396);
not NOT1 (N944, N937);
nor NOR4 (N945, N941, N259, N262, N389);
nor NOR4 (N946, N939, N763, N458, N502);
buf BUF1 (N947, N945);
buf BUF1 (N948, N935);
nand NAND4 (N949, N822, N42, N596, N223);
and AND3 (N950, N947, N191, N681);
xor XOR2 (N951, N942, N699);
buf BUF1 (N952, N927);
buf BUF1 (N953, N948);
nor NOR4 (N954, N944, N881, N616, N403);
and AND4 (N955, N946, N320, N525, N139);
xor XOR2 (N956, N949, N326);
nand NAND4 (N957, N953, N815, N298, N360);
buf BUF1 (N958, N951);
not NOT1 (N959, N940);
and AND4 (N960, N955, N203, N261, N739);
xor XOR2 (N961, N943, N939);
buf BUF1 (N962, N954);
not NOT1 (N963, N956);
nor NOR3 (N964, N963, N897, N213);
or OR2 (N965, N952, N305);
and AND3 (N966, N960, N111, N354);
buf BUF1 (N967, N965);
and AND4 (N968, N950, N322, N465, N185);
not NOT1 (N969, N966);
buf BUF1 (N970, N964);
xor XOR2 (N971, N967, N194);
nor NOR4 (N972, N961, N865, N64, N464);
nor NOR4 (N973, N959, N498, N1, N332);
or OR3 (N974, N909, N401, N828);
xor XOR2 (N975, N968, N254);
buf BUF1 (N976, N958);
xor XOR2 (N977, N957, N946);
not NOT1 (N978, N972);
nor NOR2 (N979, N974, N784);
and AND3 (N980, N971, N31, N289);
nor NOR2 (N981, N979, N146);
and AND3 (N982, N978, N648, N161);
not NOT1 (N983, N973);
buf BUF1 (N984, N982);
xor XOR2 (N985, N983, N496);
buf BUF1 (N986, N980);
nand NAND2 (N987, N969, N69);
nor NOR2 (N988, N986, N113);
buf BUF1 (N989, N970);
and AND2 (N990, N989, N140);
nor NOR4 (N991, N981, N113, N414, N287);
nand NAND2 (N992, N977, N547);
nand NAND3 (N993, N984, N805, N925);
nand NAND4 (N994, N991, N40, N10, N99);
nand NAND3 (N995, N975, N71, N404);
buf BUF1 (N996, N988);
or OR2 (N997, N962, N989);
not NOT1 (N998, N996);
xor XOR2 (N999, N985, N618);
nor NOR3 (N1000, N999, N756, N788);
buf BUF1 (N1001, N976);
xor XOR2 (N1002, N992, N676);
buf BUF1 (N1003, N998);
nand NAND4 (N1004, N997, N63, N910, N86);
xor XOR2 (N1005, N993, N409);
nor NOR3 (N1006, N994, N690, N344);
xor XOR2 (N1007, N1004, N897);
buf BUF1 (N1008, N1005);
not NOT1 (N1009, N987);
or OR3 (N1010, N1000, N820, N448);
nor NOR3 (N1011, N1009, N441, N572);
nor NOR2 (N1012, N1006, N700);
not NOT1 (N1013, N1011);
buf BUF1 (N1014, N1008);
nor NOR3 (N1015, N1007, N587, N629);
xor XOR2 (N1016, N1015, N747);
not NOT1 (N1017, N1014);
and AND4 (N1018, N1016, N27, N979, N1008);
nand NAND4 (N1019, N1010, N980, N135, N827);
nand NAND3 (N1020, N995, N308, N441);
nand NAND4 (N1021, N1020, N574, N1019, N945);
nor NOR2 (N1022, N735, N755);
nor NOR2 (N1023, N1013, N100);
not NOT1 (N1024, N1018);
or OR2 (N1025, N1022, N754);
nor NOR3 (N1026, N1017, N663, N790);
and AND4 (N1027, N1025, N691, N167, N610);
or OR4 (N1028, N1027, N767, N319, N1015);
nor NOR4 (N1029, N1012, N324, N686, N762);
and AND4 (N1030, N1026, N900, N451, N656);
xor XOR2 (N1031, N1001, N374);
and AND4 (N1032, N1003, N284, N469, N921);
or OR2 (N1033, N1023, N70);
nor NOR3 (N1034, N1031, N880, N543);
nand NAND4 (N1035, N1021, N7, N735, N894);
xor XOR2 (N1036, N1034, N207);
xor XOR2 (N1037, N1002, N688);
not NOT1 (N1038, N990);
nor NOR2 (N1039, N1035, N913);
buf BUF1 (N1040, N1036);
or OR2 (N1041, N1037, N46);
xor XOR2 (N1042, N1033, N393);
nand NAND2 (N1043, N1038, N596);
nand NAND2 (N1044, N1029, N974);
buf BUF1 (N1045, N1042);
or OR4 (N1046, N1044, N827, N424, N187);
nand NAND3 (N1047, N1045, N858, N156);
nand NAND3 (N1048, N1024, N274, N911);
nor NOR4 (N1049, N1041, N995, N358, N540);
nor NOR2 (N1050, N1046, N591);
buf BUF1 (N1051, N1050);
not NOT1 (N1052, N1043);
buf BUF1 (N1053, N1048);
buf BUF1 (N1054, N1053);
or OR2 (N1055, N1047, N1012);
xor XOR2 (N1056, N1055, N30);
or OR3 (N1057, N1040, N1047, N339);
not NOT1 (N1058, N1054);
not NOT1 (N1059, N1052);
and AND4 (N1060, N1056, N956, N456, N805);
not NOT1 (N1061, N1028);
or OR3 (N1062, N1049, N277, N186);
xor XOR2 (N1063, N1060, N728);
not NOT1 (N1064, N1062);
not NOT1 (N1065, N1063);
nand NAND4 (N1066, N1032, N526, N336, N415);
nor NOR4 (N1067, N1057, N915, N631, N498);
nor NOR3 (N1068, N1051, N362, N558);
or OR3 (N1069, N1058, N900, N112);
nor NOR2 (N1070, N1066, N627);
buf BUF1 (N1071, N1064);
xor XOR2 (N1072, N1069, N430);
and AND4 (N1073, N1059, N93, N102, N269);
nor NOR4 (N1074, N1065, N542, N141, N44);
nor NOR3 (N1075, N1030, N596, N357);
nor NOR4 (N1076, N1075, N701, N817, N1046);
xor XOR2 (N1077, N1071, N64);
or OR3 (N1078, N1070, N815, N281);
not NOT1 (N1079, N1067);
buf BUF1 (N1080, N1068);
or OR3 (N1081, N1073, N284, N197);
xor XOR2 (N1082, N1061, N352);
or OR3 (N1083, N1081, N264, N766);
not NOT1 (N1084, N1074);
nor NOR2 (N1085, N1039, N611);
xor XOR2 (N1086, N1083, N556);
buf BUF1 (N1087, N1080);
xor XOR2 (N1088, N1087, N987);
nor NOR4 (N1089, N1076, N512, N6, N105);
nor NOR2 (N1090, N1078, N786);
not NOT1 (N1091, N1072);
nand NAND2 (N1092, N1079, N529);
buf BUF1 (N1093, N1092);
or OR3 (N1094, N1077, N80, N900);
and AND3 (N1095, N1093, N271, N633);
xor XOR2 (N1096, N1086, N171);
or OR2 (N1097, N1088, N1022);
buf BUF1 (N1098, N1090);
nand NAND4 (N1099, N1084, N861, N455, N7);
xor XOR2 (N1100, N1089, N14);
not NOT1 (N1101, N1082);
buf BUF1 (N1102, N1094);
nand NAND3 (N1103, N1099, N834, N750);
or OR3 (N1104, N1101, N842, N106);
not NOT1 (N1105, N1102);
nand NAND3 (N1106, N1085, N591, N579);
not NOT1 (N1107, N1103);
not NOT1 (N1108, N1107);
nor NOR4 (N1109, N1098, N28, N438, N944);
or OR2 (N1110, N1105, N454);
nor NOR2 (N1111, N1095, N375);
xor XOR2 (N1112, N1100, N659);
and AND4 (N1113, N1111, N492, N269, N487);
xor XOR2 (N1114, N1108, N873);
nand NAND3 (N1115, N1096, N195, N280);
xor XOR2 (N1116, N1091, N1028);
and AND3 (N1117, N1114, N150, N586);
xor XOR2 (N1118, N1106, N151);
buf BUF1 (N1119, N1104);
or OR3 (N1120, N1110, N458, N588);
xor XOR2 (N1121, N1097, N772);
not NOT1 (N1122, N1121);
nand NAND3 (N1123, N1115, N465, N528);
buf BUF1 (N1124, N1109);
xor XOR2 (N1125, N1116, N652);
buf BUF1 (N1126, N1120);
not NOT1 (N1127, N1126);
nand NAND2 (N1128, N1127, N264);
buf BUF1 (N1129, N1118);
nand NAND2 (N1130, N1129, N836);
not NOT1 (N1131, N1119);
nor NOR2 (N1132, N1113, N38);
and AND4 (N1133, N1123, N162, N410, N837);
or OR2 (N1134, N1117, N760);
nor NOR3 (N1135, N1128, N311, N620);
and AND2 (N1136, N1124, N1097);
not NOT1 (N1137, N1133);
buf BUF1 (N1138, N1134);
nor NOR4 (N1139, N1132, N169, N601, N483);
and AND2 (N1140, N1139, N267);
nor NOR3 (N1141, N1122, N635, N127);
xor XOR2 (N1142, N1140, N225);
nand NAND4 (N1143, N1136, N1021, N801, N1005);
nand NAND4 (N1144, N1112, N867, N432, N257);
nand NAND4 (N1145, N1144, N595, N979, N389);
not NOT1 (N1146, N1137);
xor XOR2 (N1147, N1146, N891);
nor NOR2 (N1148, N1147, N876);
and AND3 (N1149, N1148, N754, N21);
buf BUF1 (N1150, N1130);
buf BUF1 (N1151, N1145);
buf BUF1 (N1152, N1141);
or OR2 (N1153, N1135, N786);
nand NAND3 (N1154, N1138, N803, N1016);
nor NOR3 (N1155, N1143, N674, N880);
not NOT1 (N1156, N1142);
nand NAND2 (N1157, N1151, N256);
and AND2 (N1158, N1153, N738);
buf BUF1 (N1159, N1131);
xor XOR2 (N1160, N1157, N925);
and AND4 (N1161, N1159, N1068, N564, N517);
nor NOR2 (N1162, N1158, N390);
xor XOR2 (N1163, N1156, N724);
buf BUF1 (N1164, N1155);
and AND3 (N1165, N1162, N815, N395);
nand NAND4 (N1166, N1163, N433, N391, N225);
or OR4 (N1167, N1150, N538, N1066, N726);
or OR3 (N1168, N1149, N1085, N1066);
or OR2 (N1169, N1167, N251);
buf BUF1 (N1170, N1166);
buf BUF1 (N1171, N1165);
buf BUF1 (N1172, N1169);
buf BUF1 (N1173, N1164);
nor NOR3 (N1174, N1161, N274, N702);
nand NAND3 (N1175, N1170, N765, N2);
not NOT1 (N1176, N1175);
or OR3 (N1177, N1154, N887, N757);
or OR3 (N1178, N1125, N396, N1058);
nor NOR2 (N1179, N1174, N597);
or OR4 (N1180, N1178, N458, N1035, N988);
and AND3 (N1181, N1173, N855, N163);
or OR2 (N1182, N1171, N354);
xor XOR2 (N1183, N1182, N163);
nand NAND2 (N1184, N1176, N740);
not NOT1 (N1185, N1179);
nor NOR4 (N1186, N1180, N1162, N575, N1170);
buf BUF1 (N1187, N1172);
nor NOR4 (N1188, N1160, N1087, N78, N975);
and AND3 (N1189, N1181, N346, N989);
buf BUF1 (N1190, N1187);
or OR2 (N1191, N1188, N994);
nor NOR3 (N1192, N1168, N467, N1168);
not NOT1 (N1193, N1177);
nor NOR2 (N1194, N1186, N1029);
not NOT1 (N1195, N1190);
nand NAND3 (N1196, N1189, N307, N913);
or OR4 (N1197, N1184, N34, N480, N167);
not NOT1 (N1198, N1192);
xor XOR2 (N1199, N1197, N670);
nand NAND2 (N1200, N1194, N906);
xor XOR2 (N1201, N1200, N255);
nand NAND4 (N1202, N1152, N213, N6, N584);
buf BUF1 (N1203, N1195);
buf BUF1 (N1204, N1185);
nand NAND3 (N1205, N1201, N1154, N914);
buf BUF1 (N1206, N1204);
and AND2 (N1207, N1203, N20);
not NOT1 (N1208, N1206);
and AND3 (N1209, N1196, N635, N646);
buf BUF1 (N1210, N1208);
and AND3 (N1211, N1210, N475, N162);
buf BUF1 (N1212, N1198);
xor XOR2 (N1213, N1211, N758);
xor XOR2 (N1214, N1202, N1166);
nor NOR3 (N1215, N1205, N1027, N896);
or OR2 (N1216, N1183, N1157);
or OR4 (N1217, N1215, N423, N215, N715);
or OR4 (N1218, N1213, N1213, N207, N890);
or OR2 (N1219, N1209, N944);
and AND4 (N1220, N1207, N358, N596, N399);
or OR3 (N1221, N1217, N768, N969);
nor NOR4 (N1222, N1199, N872, N1215, N15);
nor NOR3 (N1223, N1222, N955, N914);
nor NOR2 (N1224, N1191, N1117);
nand NAND3 (N1225, N1219, N278, N186);
and AND3 (N1226, N1224, N739, N967);
not NOT1 (N1227, N1226);
not NOT1 (N1228, N1212);
nand NAND2 (N1229, N1193, N103);
xor XOR2 (N1230, N1214, N158);
and AND4 (N1231, N1216, N40, N664, N1020);
buf BUF1 (N1232, N1223);
buf BUF1 (N1233, N1229);
or OR3 (N1234, N1218, N703, N482);
buf BUF1 (N1235, N1234);
or OR2 (N1236, N1230, N940);
nor NOR3 (N1237, N1235, N991, N270);
nand NAND2 (N1238, N1236, N806);
nor NOR2 (N1239, N1237, N271);
and AND2 (N1240, N1220, N299);
nor NOR2 (N1241, N1233, N805);
nor NOR4 (N1242, N1240, N669, N369, N897);
nand NAND4 (N1243, N1241, N850, N87, N855);
and AND3 (N1244, N1232, N797, N1162);
and AND4 (N1245, N1225, N635, N544, N690);
nor NOR2 (N1246, N1239, N9);
or OR4 (N1247, N1238, N134, N83, N1223);
and AND3 (N1248, N1228, N415, N995);
not NOT1 (N1249, N1247);
nand NAND4 (N1250, N1244, N1161, N449, N498);
buf BUF1 (N1251, N1250);
nand NAND2 (N1252, N1242, N1202);
not NOT1 (N1253, N1246);
xor XOR2 (N1254, N1251, N644);
xor XOR2 (N1255, N1221, N908);
xor XOR2 (N1256, N1248, N495);
buf BUF1 (N1257, N1252);
nor NOR4 (N1258, N1256, N1073, N693, N1021);
or OR2 (N1259, N1257, N135);
nand NAND2 (N1260, N1227, N413);
and AND4 (N1261, N1231, N498, N727, N1183);
not NOT1 (N1262, N1249);
and AND2 (N1263, N1245, N397);
buf BUF1 (N1264, N1259);
not NOT1 (N1265, N1263);
and AND3 (N1266, N1261, N187, N526);
nand NAND2 (N1267, N1258, N991);
or OR2 (N1268, N1266, N101);
and AND4 (N1269, N1253, N123, N104, N330);
nand NAND4 (N1270, N1260, N1012, N111, N712);
xor XOR2 (N1271, N1254, N57);
and AND2 (N1272, N1269, N961);
or OR2 (N1273, N1268, N131);
nand NAND3 (N1274, N1270, N1220, N960);
buf BUF1 (N1275, N1271);
nor NOR2 (N1276, N1262, N1273);
nand NAND4 (N1277, N1016, N1154, N784, N273);
xor XOR2 (N1278, N1274, N66);
or OR4 (N1279, N1267, N955, N47, N972);
buf BUF1 (N1280, N1279);
nand NAND3 (N1281, N1275, N716, N677);
not NOT1 (N1282, N1265);
xor XOR2 (N1283, N1272, N104);
xor XOR2 (N1284, N1283, N256);
or OR3 (N1285, N1281, N1121, N1168);
not NOT1 (N1286, N1243);
not NOT1 (N1287, N1276);
nand NAND2 (N1288, N1280, N374);
nor NOR2 (N1289, N1277, N519);
or OR4 (N1290, N1288, N75, N535, N873);
nand NAND3 (N1291, N1278, N386, N1008);
nor NOR4 (N1292, N1285, N1226, N1250, N1016);
not NOT1 (N1293, N1292);
xor XOR2 (N1294, N1287, N773);
and AND3 (N1295, N1286, N147, N1258);
or OR3 (N1296, N1255, N153, N427);
xor XOR2 (N1297, N1284, N492);
or OR4 (N1298, N1293, N1206, N449, N998);
nor NOR2 (N1299, N1295, N131);
xor XOR2 (N1300, N1289, N104);
or OR4 (N1301, N1297, N261, N1117, N825);
or OR3 (N1302, N1299, N151, N402);
or OR2 (N1303, N1290, N221);
nor NOR4 (N1304, N1296, N132, N1058, N300);
xor XOR2 (N1305, N1304, N90);
not NOT1 (N1306, N1301);
nand NAND4 (N1307, N1294, N671, N1028, N476);
or OR4 (N1308, N1264, N748, N1064, N243);
nor NOR3 (N1309, N1302, N1117, N1215);
nand NAND4 (N1310, N1291, N898, N818, N1034);
nand NAND4 (N1311, N1300, N1307, N987, N735);
not NOT1 (N1312, N160);
not NOT1 (N1313, N1298);
nor NOR2 (N1314, N1306, N264);
nor NOR3 (N1315, N1313, N420, N113);
and AND4 (N1316, N1314, N705, N1053, N784);
or OR3 (N1317, N1316, N685, N759);
not NOT1 (N1318, N1311);
nor NOR2 (N1319, N1315, N197);
buf BUF1 (N1320, N1308);
and AND2 (N1321, N1282, N436);
not NOT1 (N1322, N1318);
and AND4 (N1323, N1321, N1027, N250, N216);
nor NOR2 (N1324, N1317, N1188);
and AND4 (N1325, N1323, N729, N228, N786);
xor XOR2 (N1326, N1319, N409);
buf BUF1 (N1327, N1320);
or OR4 (N1328, N1303, N892, N133, N614);
buf BUF1 (N1329, N1322);
or OR4 (N1330, N1309, N103, N1311, N753);
buf BUF1 (N1331, N1326);
nor NOR3 (N1332, N1324, N878, N188);
nand NAND4 (N1333, N1312, N1118, N479, N582);
nor NOR3 (N1334, N1333, N1141, N736);
or OR3 (N1335, N1310, N314, N1040);
and AND3 (N1336, N1334, N1314, N123);
xor XOR2 (N1337, N1325, N274);
nand NAND4 (N1338, N1331, N51, N371, N644);
and AND4 (N1339, N1329, N399, N984, N1278);
nor NOR4 (N1340, N1337, N1011, N224, N1065);
or OR4 (N1341, N1339, N1035, N259, N1236);
not NOT1 (N1342, N1327);
and AND4 (N1343, N1336, N740, N1161, N1005);
nor NOR2 (N1344, N1340, N1139);
nor NOR3 (N1345, N1330, N1138, N1314);
not NOT1 (N1346, N1338);
and AND2 (N1347, N1328, N248);
nor NOR4 (N1348, N1343, N735, N891, N547);
xor XOR2 (N1349, N1345, N925);
xor XOR2 (N1350, N1349, N390);
buf BUF1 (N1351, N1344);
nor NOR4 (N1352, N1346, N885, N64, N88);
xor XOR2 (N1353, N1305, N58);
or OR4 (N1354, N1347, N705, N192, N561);
and AND2 (N1355, N1342, N597);
nand NAND2 (N1356, N1353, N405);
and AND3 (N1357, N1352, N230, N807);
nand NAND4 (N1358, N1355, N354, N820, N641);
nor NOR3 (N1359, N1358, N312, N1229);
not NOT1 (N1360, N1332);
and AND4 (N1361, N1341, N406, N456, N264);
nor NOR4 (N1362, N1350, N675, N372, N582);
and AND4 (N1363, N1362, N1233, N335, N673);
or OR4 (N1364, N1357, N136, N351, N180);
and AND3 (N1365, N1348, N696, N1082);
xor XOR2 (N1366, N1364, N976);
nand NAND4 (N1367, N1359, N1073, N66, N552);
nor NOR3 (N1368, N1363, N754, N1354);
and AND3 (N1369, N684, N434, N566);
buf BUF1 (N1370, N1361);
not NOT1 (N1371, N1335);
xor XOR2 (N1372, N1371, N1249);
and AND4 (N1373, N1366, N272, N258, N677);
or OR4 (N1374, N1365, N855, N320, N300);
not NOT1 (N1375, N1360);
xor XOR2 (N1376, N1374, N1002);
nand NAND3 (N1377, N1376, N139, N78);
or OR2 (N1378, N1369, N858);
nor NOR4 (N1379, N1377, N1318, N947, N1063);
buf BUF1 (N1380, N1372);
xor XOR2 (N1381, N1379, N536);
or OR4 (N1382, N1380, N261, N666, N625);
not NOT1 (N1383, N1381);
not NOT1 (N1384, N1375);
nand NAND4 (N1385, N1378, N1259, N33, N1221);
xor XOR2 (N1386, N1356, N635);
xor XOR2 (N1387, N1385, N198);
buf BUF1 (N1388, N1383);
xor XOR2 (N1389, N1384, N240);
or OR4 (N1390, N1387, N1350, N982, N186);
nand NAND2 (N1391, N1370, N657);
nand NAND3 (N1392, N1367, N430, N630);
xor XOR2 (N1393, N1382, N154);
and AND3 (N1394, N1389, N709, N1381);
or OR2 (N1395, N1388, N700);
xor XOR2 (N1396, N1391, N105);
nand NAND4 (N1397, N1386, N475, N1034, N549);
and AND3 (N1398, N1396, N806, N1327);
xor XOR2 (N1399, N1397, N589);
or OR4 (N1400, N1373, N165, N641, N1);
not NOT1 (N1401, N1399);
xor XOR2 (N1402, N1394, N970);
not NOT1 (N1403, N1351);
or OR3 (N1404, N1401, N630, N176);
nor NOR2 (N1405, N1402, N1072);
nor NOR4 (N1406, N1392, N496, N276, N173);
xor XOR2 (N1407, N1395, N369);
or OR2 (N1408, N1390, N21);
nor NOR4 (N1409, N1398, N189, N247, N1220);
buf BUF1 (N1410, N1409);
buf BUF1 (N1411, N1400);
not NOT1 (N1412, N1406);
nor NOR4 (N1413, N1404, N328, N757, N688);
xor XOR2 (N1414, N1403, N1048);
or OR3 (N1415, N1412, N346, N836);
not NOT1 (N1416, N1411);
buf BUF1 (N1417, N1413);
nand NAND4 (N1418, N1405, N105, N1012, N664);
and AND2 (N1419, N1407, N876);
buf BUF1 (N1420, N1408);
or OR4 (N1421, N1418, N948, N1089, N471);
not NOT1 (N1422, N1415);
nor NOR2 (N1423, N1368, N1408);
nor NOR3 (N1424, N1421, N887, N462);
buf BUF1 (N1425, N1422);
buf BUF1 (N1426, N1424);
buf BUF1 (N1427, N1414);
or OR3 (N1428, N1423, N944, N641);
nand NAND2 (N1429, N1393, N531);
or OR2 (N1430, N1427, N278);
buf BUF1 (N1431, N1410);
and AND4 (N1432, N1429, N117, N713, N1265);
xor XOR2 (N1433, N1428, N180);
or OR4 (N1434, N1432, N1159, N137, N1);
buf BUF1 (N1435, N1431);
buf BUF1 (N1436, N1417);
or OR2 (N1437, N1436, N727);
xor XOR2 (N1438, N1435, N447);
buf BUF1 (N1439, N1438);
not NOT1 (N1440, N1434);
buf BUF1 (N1441, N1440);
xor XOR2 (N1442, N1430, N147);
or OR4 (N1443, N1416, N711, N1299, N30);
xor XOR2 (N1444, N1439, N974);
xor XOR2 (N1445, N1444, N1248);
or OR3 (N1446, N1425, N665, N270);
not NOT1 (N1447, N1442);
xor XOR2 (N1448, N1445, N325);
nand NAND4 (N1449, N1433, N1301, N1426, N927);
xor XOR2 (N1450, N1308, N1414);
not NOT1 (N1451, N1437);
not NOT1 (N1452, N1451);
nand NAND3 (N1453, N1446, N354, N365);
and AND3 (N1454, N1419, N73, N708);
or OR4 (N1455, N1420, N1010, N1419, N1001);
and AND2 (N1456, N1452, N622);
xor XOR2 (N1457, N1443, N555);
nand NAND4 (N1458, N1447, N266, N466, N116);
buf BUF1 (N1459, N1450);
nor NOR4 (N1460, N1454, N1381, N302, N288);
buf BUF1 (N1461, N1448);
nor NOR2 (N1462, N1453, N1152);
xor XOR2 (N1463, N1458, N1448);
nor NOR4 (N1464, N1462, N1187, N444, N474);
nor NOR2 (N1465, N1459, N240);
or OR3 (N1466, N1449, N826, N123);
and AND2 (N1467, N1463, N873);
not NOT1 (N1468, N1465);
nand NAND2 (N1469, N1455, N862);
or OR4 (N1470, N1456, N307, N1117, N173);
or OR4 (N1471, N1468, N855, N36, N1153);
xor XOR2 (N1472, N1441, N1285);
not NOT1 (N1473, N1461);
not NOT1 (N1474, N1473);
not NOT1 (N1475, N1457);
nand NAND2 (N1476, N1466, N519);
buf BUF1 (N1477, N1464);
nor NOR4 (N1478, N1470, N679, N1296, N1308);
nand NAND3 (N1479, N1472, N372, N1002);
not NOT1 (N1480, N1460);
not NOT1 (N1481, N1477);
xor XOR2 (N1482, N1469, N1241);
or OR4 (N1483, N1471, N863, N595, N1392);
nor NOR3 (N1484, N1482, N569, N605);
and AND3 (N1485, N1480, N320, N1396);
xor XOR2 (N1486, N1467, N961);
xor XOR2 (N1487, N1485, N1080);
nand NAND3 (N1488, N1474, N1128, N1140);
and AND2 (N1489, N1476, N340);
not NOT1 (N1490, N1475);
nor NOR2 (N1491, N1486, N1437);
or OR3 (N1492, N1490, N550, N393);
nor NOR3 (N1493, N1483, N63, N894);
and AND3 (N1494, N1488, N282, N644);
nand NAND4 (N1495, N1478, N170, N734, N173);
nor NOR4 (N1496, N1495, N507, N278, N129);
not NOT1 (N1497, N1489);
or OR3 (N1498, N1487, N811, N1348);
xor XOR2 (N1499, N1481, N1430);
buf BUF1 (N1500, N1492);
not NOT1 (N1501, N1498);
or OR3 (N1502, N1494, N650, N1228);
xor XOR2 (N1503, N1500, N1087);
not NOT1 (N1504, N1479);
nor NOR3 (N1505, N1502, N1383, N681);
xor XOR2 (N1506, N1504, N1384);
buf BUF1 (N1507, N1496);
not NOT1 (N1508, N1501);
xor XOR2 (N1509, N1508, N1239);
buf BUF1 (N1510, N1509);
xor XOR2 (N1511, N1505, N159);
xor XOR2 (N1512, N1499, N736);
nor NOR3 (N1513, N1491, N915, N782);
buf BUF1 (N1514, N1513);
nand NAND2 (N1515, N1506, N1117);
nor NOR3 (N1516, N1484, N1231, N843);
and AND3 (N1517, N1510, N398, N506);
xor XOR2 (N1518, N1507, N113);
not NOT1 (N1519, N1497);
and AND2 (N1520, N1514, N295);
or OR4 (N1521, N1493, N231, N1086, N490);
not NOT1 (N1522, N1517);
or OR3 (N1523, N1503, N478, N1486);
and AND4 (N1524, N1520, N1397, N500, N1444);
or OR2 (N1525, N1524, N1513);
buf BUF1 (N1526, N1522);
not NOT1 (N1527, N1521);
xor XOR2 (N1528, N1519, N762);
and AND2 (N1529, N1516, N403);
and AND3 (N1530, N1529, N670, N1264);
not NOT1 (N1531, N1523);
xor XOR2 (N1532, N1515, N8);
buf BUF1 (N1533, N1526);
or OR4 (N1534, N1531, N1526, N149, N529);
buf BUF1 (N1535, N1528);
buf BUF1 (N1536, N1532);
or OR2 (N1537, N1512, N1138);
or OR3 (N1538, N1511, N1113, N1168);
not NOT1 (N1539, N1534);
or OR2 (N1540, N1539, N222);
buf BUF1 (N1541, N1533);
not NOT1 (N1542, N1537);
nand NAND2 (N1543, N1530, N323);
nor NOR3 (N1544, N1538, N730, N1161);
nand NAND3 (N1545, N1525, N101, N263);
xor XOR2 (N1546, N1543, N915);
or OR3 (N1547, N1518, N1495, N317);
nor NOR4 (N1548, N1541, N354, N724, N820);
nand NAND4 (N1549, N1544, N1009, N713, N1224);
not NOT1 (N1550, N1545);
nand NAND3 (N1551, N1546, N915, N432);
not NOT1 (N1552, N1540);
and AND3 (N1553, N1548, N413, N1287);
not NOT1 (N1554, N1550);
not NOT1 (N1555, N1535);
not NOT1 (N1556, N1527);
or OR3 (N1557, N1547, N595, N1067);
buf BUF1 (N1558, N1551);
and AND3 (N1559, N1536, N382, N776);
and AND4 (N1560, N1553, N112, N112, N518);
buf BUF1 (N1561, N1557);
and AND4 (N1562, N1561, N20, N1069, N952);
not NOT1 (N1563, N1562);
nand NAND4 (N1564, N1549, N1218, N1402, N1183);
or OR3 (N1565, N1542, N1111, N336);
nand NAND2 (N1566, N1563, N1037);
not NOT1 (N1567, N1555);
xor XOR2 (N1568, N1554, N1226);
not NOT1 (N1569, N1552);
buf BUF1 (N1570, N1567);
xor XOR2 (N1571, N1564, N1088);
nand NAND2 (N1572, N1556, N1009);
nor NOR4 (N1573, N1558, N731, N60, N88);
buf BUF1 (N1574, N1559);
and AND2 (N1575, N1560, N501);
xor XOR2 (N1576, N1570, N999);
nand NAND2 (N1577, N1569, N35);
nor NOR2 (N1578, N1574, N120);
nor NOR2 (N1579, N1573, N1063);
nand NAND4 (N1580, N1579, N702, N1229, N863);
not NOT1 (N1581, N1577);
or OR3 (N1582, N1571, N1173, N469);
or OR2 (N1583, N1581, N1229);
or OR2 (N1584, N1565, N311);
nand NAND3 (N1585, N1578, N107, N275);
or OR3 (N1586, N1575, N1153, N603);
and AND3 (N1587, N1582, N138, N499);
not NOT1 (N1588, N1572);
and AND2 (N1589, N1580, N1343);
nand NAND2 (N1590, N1586, N264);
not NOT1 (N1591, N1585);
nand NAND2 (N1592, N1566, N364);
nand NAND3 (N1593, N1592, N1038, N1127);
xor XOR2 (N1594, N1589, N1048);
and AND3 (N1595, N1594, N108, N785);
nor NOR3 (N1596, N1593, N718, N305);
or OR4 (N1597, N1584, N909, N857, N450);
xor XOR2 (N1598, N1595, N359);
not NOT1 (N1599, N1597);
xor XOR2 (N1600, N1568, N1486);
and AND3 (N1601, N1600, N1283, N192);
buf BUF1 (N1602, N1590);
not NOT1 (N1603, N1576);
nand NAND2 (N1604, N1598, N1587);
not NOT1 (N1605, N309);
nand NAND3 (N1606, N1596, N546, N1040);
buf BUF1 (N1607, N1601);
and AND4 (N1608, N1604, N320, N808, N256);
or OR2 (N1609, N1606, N538);
not NOT1 (N1610, N1607);
and AND2 (N1611, N1602, N325);
nor NOR2 (N1612, N1591, N1047);
nand NAND4 (N1613, N1608, N66, N1194, N1509);
nand NAND4 (N1614, N1605, N434, N1285, N271);
or OR3 (N1615, N1610, N96, N1032);
nor NOR4 (N1616, N1609, N498, N1178, N1147);
or OR2 (N1617, N1611, N1458);
nor NOR2 (N1618, N1615, N353);
xor XOR2 (N1619, N1616, N946);
and AND3 (N1620, N1603, N653, N1425);
xor XOR2 (N1621, N1599, N1118);
xor XOR2 (N1622, N1612, N101);
nand NAND2 (N1623, N1619, N272);
buf BUF1 (N1624, N1614);
not NOT1 (N1625, N1618);
buf BUF1 (N1626, N1625);
or OR2 (N1627, N1621, N337);
buf BUF1 (N1628, N1613);
not NOT1 (N1629, N1588);
nor NOR2 (N1630, N1583, N999);
not NOT1 (N1631, N1627);
and AND2 (N1632, N1630, N666);
not NOT1 (N1633, N1632);
or OR4 (N1634, N1628, N88, N1246, N208);
buf BUF1 (N1635, N1624);
nor NOR3 (N1636, N1634, N580, N144);
xor XOR2 (N1637, N1636, N1225);
and AND3 (N1638, N1629, N974, N245);
or OR2 (N1639, N1617, N242);
nand NAND2 (N1640, N1622, N707);
nor NOR3 (N1641, N1623, N53, N353);
nor NOR3 (N1642, N1641, N1394, N461);
nor NOR2 (N1643, N1620, N494);
nand NAND2 (N1644, N1637, N1274);
nand NAND3 (N1645, N1631, N756, N1609);
buf BUF1 (N1646, N1642);
not NOT1 (N1647, N1644);
nor NOR4 (N1648, N1635, N343, N605, N329);
or OR4 (N1649, N1646, N1323, N1555, N1087);
not NOT1 (N1650, N1633);
xor XOR2 (N1651, N1639, N1552);
xor XOR2 (N1652, N1643, N535);
buf BUF1 (N1653, N1650);
nor NOR4 (N1654, N1648, N1082, N1488, N1099);
nor NOR4 (N1655, N1654, N666, N1087, N1186);
nand NAND4 (N1656, N1652, N1400, N392, N1485);
and AND2 (N1657, N1645, N62);
buf BUF1 (N1658, N1638);
nand NAND2 (N1659, N1655, N1503);
not NOT1 (N1660, N1640);
buf BUF1 (N1661, N1649);
nor NOR3 (N1662, N1659, N1236, N1202);
nand NAND3 (N1663, N1658, N638, N1103);
not NOT1 (N1664, N1653);
nor NOR2 (N1665, N1657, N882);
not NOT1 (N1666, N1651);
nand NAND4 (N1667, N1660, N239, N595, N214);
not NOT1 (N1668, N1665);
xor XOR2 (N1669, N1647, N565);
and AND3 (N1670, N1626, N919, N94);
buf BUF1 (N1671, N1656);
not NOT1 (N1672, N1668);
and AND4 (N1673, N1671, N805, N496, N677);
not NOT1 (N1674, N1661);
or OR3 (N1675, N1662, N111, N341);
or OR4 (N1676, N1673, N621, N978, N993);
nand NAND4 (N1677, N1670, N933, N1376, N1566);
buf BUF1 (N1678, N1664);
buf BUF1 (N1679, N1676);
buf BUF1 (N1680, N1663);
or OR4 (N1681, N1669, N815, N1563, N1420);
not NOT1 (N1682, N1677);
and AND4 (N1683, N1672, N208, N711, N280);
xor XOR2 (N1684, N1681, N920);
nor NOR4 (N1685, N1666, N1380, N391, N744);
or OR2 (N1686, N1674, N1161);
nor NOR4 (N1687, N1678, N507, N722, N640);
and AND3 (N1688, N1682, N230, N219);
xor XOR2 (N1689, N1684, N1272);
not NOT1 (N1690, N1688);
and AND2 (N1691, N1689, N1337);
and AND2 (N1692, N1679, N505);
buf BUF1 (N1693, N1680);
xor XOR2 (N1694, N1686, N852);
not NOT1 (N1695, N1690);
or OR2 (N1696, N1675, N477);
and AND3 (N1697, N1695, N1052, N759);
buf BUF1 (N1698, N1687);
xor XOR2 (N1699, N1692, N54);
buf BUF1 (N1700, N1693);
nand NAND3 (N1701, N1700, N993, N709);
or OR3 (N1702, N1694, N960, N322);
xor XOR2 (N1703, N1699, N1417);
or OR4 (N1704, N1683, N1261, N1053, N732);
or OR2 (N1705, N1685, N623);
nand NAND2 (N1706, N1702, N407);
buf BUF1 (N1707, N1691);
nor NOR4 (N1708, N1706, N472, N1177, N550);
buf BUF1 (N1709, N1707);
not NOT1 (N1710, N1708);
buf BUF1 (N1711, N1709);
nor NOR4 (N1712, N1698, N665, N828, N732);
not NOT1 (N1713, N1703);
xor XOR2 (N1714, N1667, N443);
buf BUF1 (N1715, N1696);
or OR2 (N1716, N1710, N914);
nor NOR2 (N1717, N1711, N1131);
nor NOR4 (N1718, N1701, N286, N510, N1212);
not NOT1 (N1719, N1704);
nand NAND4 (N1720, N1719, N1199, N58, N883);
and AND2 (N1721, N1712, N1311);
nor NOR3 (N1722, N1705, N1504, N1601);
buf BUF1 (N1723, N1715);
buf BUF1 (N1724, N1713);
and AND2 (N1725, N1721, N1601);
nor NOR3 (N1726, N1720, N808, N1318);
xor XOR2 (N1727, N1722, N1122);
not NOT1 (N1728, N1723);
xor XOR2 (N1729, N1718, N187);
and AND4 (N1730, N1724, N1642, N657, N1346);
or OR4 (N1731, N1716, N235, N97, N825);
buf BUF1 (N1732, N1717);
or OR4 (N1733, N1725, N376, N392, N1581);
or OR2 (N1734, N1733, N373);
and AND4 (N1735, N1730, N384, N1632, N47);
not NOT1 (N1736, N1727);
and AND3 (N1737, N1728, N712, N803);
not NOT1 (N1738, N1732);
nand NAND2 (N1739, N1735, N170);
xor XOR2 (N1740, N1697, N236);
or OR3 (N1741, N1740, N1634, N127);
nand NAND4 (N1742, N1741, N417, N238, N216);
nand NAND3 (N1743, N1738, N1126, N1736);
xor XOR2 (N1744, N127, N244);
xor XOR2 (N1745, N1743, N67);
nor NOR2 (N1746, N1734, N22);
or OR4 (N1747, N1744, N1584, N43, N725);
xor XOR2 (N1748, N1747, N1673);
and AND3 (N1749, N1731, N128, N8);
and AND4 (N1750, N1714, N243, N1146, N1200);
xor XOR2 (N1751, N1739, N348);
nand NAND3 (N1752, N1751, N1151, N334);
or OR3 (N1753, N1726, N1352, N1376);
or OR2 (N1754, N1742, N1398);
and AND3 (N1755, N1748, N907, N1177);
nand NAND3 (N1756, N1755, N546, N1060);
xor XOR2 (N1757, N1753, N923);
buf BUF1 (N1758, N1757);
nand NAND3 (N1759, N1745, N501, N733);
buf BUF1 (N1760, N1759);
buf BUF1 (N1761, N1758);
and AND3 (N1762, N1761, N697, N578);
xor XOR2 (N1763, N1752, N821);
nand NAND2 (N1764, N1760, N1262);
xor XOR2 (N1765, N1729, N107);
buf BUF1 (N1766, N1750);
or OR4 (N1767, N1754, N745, N1618, N889);
buf BUF1 (N1768, N1767);
xor XOR2 (N1769, N1737, N1531);
and AND2 (N1770, N1749, N310);
or OR3 (N1771, N1768, N746, N1385);
nand NAND3 (N1772, N1763, N1568, N206);
nand NAND4 (N1773, N1764, N75, N150, N1152);
or OR4 (N1774, N1773, N1465, N1213, N1643);
or OR3 (N1775, N1771, N1600, N582);
or OR2 (N1776, N1765, N1348);
not NOT1 (N1777, N1775);
nor NOR4 (N1778, N1770, N1451, N1533, N541);
nand NAND4 (N1779, N1769, N598, N751, N45);
not NOT1 (N1780, N1778);
xor XOR2 (N1781, N1766, N1182);
and AND3 (N1782, N1781, N1394, N1735);
buf BUF1 (N1783, N1756);
buf BUF1 (N1784, N1779);
nor NOR2 (N1785, N1774, N217);
not NOT1 (N1786, N1782);
nor NOR2 (N1787, N1772, N870);
not NOT1 (N1788, N1786);
not NOT1 (N1789, N1783);
nor NOR4 (N1790, N1787, N1474, N903, N1474);
not NOT1 (N1791, N1785);
not NOT1 (N1792, N1790);
buf BUF1 (N1793, N1788);
nor NOR2 (N1794, N1791, N1545);
nor NOR2 (N1795, N1789, N616);
or OR4 (N1796, N1746, N475, N809, N41);
or OR3 (N1797, N1780, N695, N991);
and AND3 (N1798, N1784, N1674, N693);
nor NOR4 (N1799, N1798, N71, N1271, N888);
nand NAND2 (N1800, N1799, N553);
nor NOR2 (N1801, N1794, N350);
buf BUF1 (N1802, N1776);
nor NOR2 (N1803, N1797, N404);
nor NOR3 (N1804, N1796, N595, N1382);
nand NAND2 (N1805, N1801, N1005);
nand NAND2 (N1806, N1793, N629);
xor XOR2 (N1807, N1762, N90);
xor XOR2 (N1808, N1792, N1119);
and AND2 (N1809, N1802, N94);
or OR2 (N1810, N1807, N508);
xor XOR2 (N1811, N1795, N483);
or OR2 (N1812, N1777, N1450);
not NOT1 (N1813, N1800);
or OR4 (N1814, N1806, N1138, N1254, N594);
nor NOR2 (N1815, N1814, N240);
nor NOR3 (N1816, N1812, N129, N1423);
xor XOR2 (N1817, N1810, N1672);
or OR2 (N1818, N1808, N192);
buf BUF1 (N1819, N1804);
or OR3 (N1820, N1811, N14, N1644);
or OR4 (N1821, N1818, N159, N213, N1809);
nor NOR2 (N1822, N1778, N1783);
nand NAND2 (N1823, N1817, N189);
xor XOR2 (N1824, N1813, N1221);
nand NAND4 (N1825, N1805, N225, N15, N1524);
xor XOR2 (N1826, N1816, N1050);
not NOT1 (N1827, N1824);
nand NAND4 (N1828, N1823, N578, N959, N851);
not NOT1 (N1829, N1827);
or OR4 (N1830, N1803, N541, N1162, N472);
xor XOR2 (N1831, N1825, N529);
not NOT1 (N1832, N1829);
buf BUF1 (N1833, N1819);
buf BUF1 (N1834, N1826);
and AND4 (N1835, N1834, N1057, N717, N183);
buf BUF1 (N1836, N1821);
nor NOR2 (N1837, N1820, N791);
nor NOR2 (N1838, N1831, N385);
nor NOR3 (N1839, N1837, N610, N1620);
not NOT1 (N1840, N1822);
xor XOR2 (N1841, N1840, N1579);
nand NAND3 (N1842, N1835, N105, N1077);
not NOT1 (N1843, N1842);
buf BUF1 (N1844, N1839);
nand NAND3 (N1845, N1843, N888, N1378);
and AND2 (N1846, N1828, N1756);
nand NAND2 (N1847, N1844, N1632);
nor NOR4 (N1848, N1847, N565, N751, N430);
nor NOR4 (N1849, N1815, N1729, N1810, N1122);
not NOT1 (N1850, N1848);
and AND4 (N1851, N1833, N971, N588, N1555);
xor XOR2 (N1852, N1830, N695);
not NOT1 (N1853, N1841);
not NOT1 (N1854, N1851);
buf BUF1 (N1855, N1832);
or OR2 (N1856, N1853, N364);
not NOT1 (N1857, N1849);
buf BUF1 (N1858, N1838);
xor XOR2 (N1859, N1855, N1757);
nor NOR2 (N1860, N1850, N473);
xor XOR2 (N1861, N1859, N1082);
and AND4 (N1862, N1854, N437, N1316, N1263);
nand NAND2 (N1863, N1862, N178);
and AND4 (N1864, N1860, N1088, N1797, N1783);
not NOT1 (N1865, N1861);
not NOT1 (N1866, N1858);
and AND4 (N1867, N1845, N915, N450, N1810);
or OR3 (N1868, N1846, N1296, N221);
not NOT1 (N1869, N1867);
or OR3 (N1870, N1864, N1100, N3);
nor NOR2 (N1871, N1856, N645);
xor XOR2 (N1872, N1857, N507);
nor NOR2 (N1873, N1872, N53);
xor XOR2 (N1874, N1852, N1794);
buf BUF1 (N1875, N1870);
buf BUF1 (N1876, N1873);
nor NOR4 (N1877, N1874, N112, N309, N1756);
nor NOR3 (N1878, N1836, N1173, N428);
nor NOR3 (N1879, N1866, N1334, N723);
buf BUF1 (N1880, N1877);
and AND2 (N1881, N1863, N1486);
and AND3 (N1882, N1875, N1119, N1234);
or OR2 (N1883, N1880, N1438);
nand NAND2 (N1884, N1881, N1854);
or OR4 (N1885, N1883, N1119, N762, N152);
not NOT1 (N1886, N1879);
and AND4 (N1887, N1885, N589, N419, N195);
and AND2 (N1888, N1865, N1659);
and AND4 (N1889, N1876, N351, N257, N886);
not NOT1 (N1890, N1887);
buf BUF1 (N1891, N1886);
nand NAND2 (N1892, N1890, N1416);
or OR2 (N1893, N1889, N1543);
or OR3 (N1894, N1882, N1243, N1883);
xor XOR2 (N1895, N1891, N1610);
xor XOR2 (N1896, N1895, N1870);
nor NOR3 (N1897, N1878, N99, N371);
or OR3 (N1898, N1888, N141, N306);
or OR3 (N1899, N1893, N1865, N1150);
xor XOR2 (N1900, N1894, N1771);
nor NOR2 (N1901, N1897, N365);
buf BUF1 (N1902, N1900);
not NOT1 (N1903, N1892);
xor XOR2 (N1904, N1901, N37);
buf BUF1 (N1905, N1884);
or OR2 (N1906, N1905, N351);
not NOT1 (N1907, N1869);
or OR4 (N1908, N1907, N520, N1101, N1091);
not NOT1 (N1909, N1906);
nand NAND2 (N1910, N1908, N1795);
or OR4 (N1911, N1868, N1478, N1397, N252);
xor XOR2 (N1912, N1896, N1380);
and AND4 (N1913, N1871, N893, N649, N1389);
xor XOR2 (N1914, N1899, N694);
and AND4 (N1915, N1902, N763, N43, N733);
or OR4 (N1916, N1912, N223, N1460, N324);
or OR4 (N1917, N1916, N557, N1626, N1049);
not NOT1 (N1918, N1915);
and AND4 (N1919, N1909, N6, N666, N1039);
nand NAND4 (N1920, N1898, N248, N890, N926);
and AND2 (N1921, N1914, N29);
xor XOR2 (N1922, N1913, N1881);
nor NOR4 (N1923, N1922, N861, N1790, N1252);
or OR3 (N1924, N1918, N985, N29);
xor XOR2 (N1925, N1904, N1629);
nor NOR3 (N1926, N1910, N1761, N179);
nor NOR3 (N1927, N1920, N1771, N553);
and AND2 (N1928, N1903, N497);
nor NOR2 (N1929, N1921, N1776);
not NOT1 (N1930, N1927);
xor XOR2 (N1931, N1924, N164);
not NOT1 (N1932, N1929);
nor NOR4 (N1933, N1911, N1876, N1577, N1326);
xor XOR2 (N1934, N1932, N1689);
buf BUF1 (N1935, N1928);
nor NOR2 (N1936, N1933, N1472);
xor XOR2 (N1937, N1925, N258);
nor NOR2 (N1938, N1931, N1229);
and AND2 (N1939, N1930, N1801);
or OR4 (N1940, N1936, N1392, N1640, N838);
nor NOR4 (N1941, N1923, N1024, N546, N1483);
nand NAND4 (N1942, N1940, N1519, N585, N1085);
nor NOR4 (N1943, N1938, N180, N185, N708);
and AND4 (N1944, N1917, N1105, N1354, N1478);
and AND3 (N1945, N1939, N574, N1023);
not NOT1 (N1946, N1941);
nand NAND4 (N1947, N1926, N226, N1838, N914);
and AND2 (N1948, N1919, N1709);
not NOT1 (N1949, N1947);
buf BUF1 (N1950, N1934);
and AND3 (N1951, N1949, N1798, N1708);
nor NOR2 (N1952, N1948, N1189);
buf BUF1 (N1953, N1952);
nand NAND3 (N1954, N1945, N1531, N1554);
buf BUF1 (N1955, N1954);
nor NOR3 (N1956, N1946, N543, N1800);
nand NAND4 (N1957, N1943, N1426, N446, N729);
nor NOR3 (N1958, N1935, N539, N67);
xor XOR2 (N1959, N1956, N662);
and AND4 (N1960, N1951, N1376, N1381, N1936);
nand NAND4 (N1961, N1937, N752, N1704, N723);
xor XOR2 (N1962, N1960, N419);
and AND2 (N1963, N1957, N349);
or OR3 (N1964, N1944, N302, N1027);
and AND4 (N1965, N1962, N1330, N1518, N693);
and AND2 (N1966, N1965, N438);
xor XOR2 (N1967, N1963, N240);
not NOT1 (N1968, N1953);
buf BUF1 (N1969, N1968);
not NOT1 (N1970, N1967);
or OR2 (N1971, N1964, N1767);
buf BUF1 (N1972, N1950);
buf BUF1 (N1973, N1969);
and AND2 (N1974, N1955, N1195);
or OR3 (N1975, N1973, N602, N1218);
buf BUF1 (N1976, N1972);
buf BUF1 (N1977, N1966);
and AND3 (N1978, N1958, N1832, N157);
not NOT1 (N1979, N1961);
nand NAND4 (N1980, N1975, N1537, N1774, N1515);
nand NAND4 (N1981, N1978, N392, N1368, N1731);
and AND2 (N1982, N1980, N985);
not NOT1 (N1983, N1976);
buf BUF1 (N1984, N1974);
not NOT1 (N1985, N1981);
and AND3 (N1986, N1982, N232, N134);
nand NAND4 (N1987, N1985, N1510, N572, N9);
nor NOR3 (N1988, N1959, N1867, N90);
xor XOR2 (N1989, N1988, N1650);
xor XOR2 (N1990, N1986, N1789);
buf BUF1 (N1991, N1970);
not NOT1 (N1992, N1991);
nand NAND2 (N1993, N1992, N1085);
nand NAND4 (N1994, N1989, N202, N884, N985);
and AND2 (N1995, N1994, N1374);
nor NOR3 (N1996, N1979, N1994, N60);
not NOT1 (N1997, N1942);
not NOT1 (N1998, N1984);
and AND3 (N1999, N1998, N1988, N1044);
nand NAND4 (N2000, N1977, N1283, N572, N1592);
and AND3 (N2001, N1997, N581, N918);
nand NAND4 (N2002, N2001, N794, N157, N1960);
xor XOR2 (N2003, N2000, N459);
buf BUF1 (N2004, N1996);
nand NAND2 (N2005, N1993, N1635);
nor NOR2 (N2006, N1983, N1770);
not NOT1 (N2007, N1995);
nor NOR2 (N2008, N1971, N1615);
or OR4 (N2009, N1990, N1255, N1799, N729);
not NOT1 (N2010, N2008);
or OR4 (N2011, N1999, N1109, N1513, N1229);
nand NAND4 (N2012, N2003, N548, N912, N225);
and AND4 (N2013, N2002, N778, N1227, N1716);
or OR4 (N2014, N1987, N1646, N1384, N1770);
xor XOR2 (N2015, N2009, N2013);
nor NOR3 (N2016, N316, N1712, N1339);
or OR4 (N2017, N2014, N334, N980, N1599);
or OR3 (N2018, N2005, N1576, N1003);
or OR3 (N2019, N2017, N1489, N291);
buf BUF1 (N2020, N2011);
buf BUF1 (N2021, N2019);
and AND3 (N2022, N2020, N1337, N1007);
nor NOR3 (N2023, N2016, N818, N1458);
not NOT1 (N2024, N2012);
and AND3 (N2025, N2023, N1163, N1220);
buf BUF1 (N2026, N2007);
xor XOR2 (N2027, N2022, N1785);
or OR4 (N2028, N2004, N1984, N889, N589);
xor XOR2 (N2029, N2024, N1828);
buf BUF1 (N2030, N2006);
xor XOR2 (N2031, N2029, N232);
and AND3 (N2032, N2025, N484, N236);
nor NOR3 (N2033, N2010, N712, N600);
and AND2 (N2034, N2028, N558);
buf BUF1 (N2035, N2015);
and AND4 (N2036, N2033, N1121, N373, N330);
or OR2 (N2037, N2018, N1070);
or OR2 (N2038, N2034, N1146);
nand NAND2 (N2039, N2038, N1273);
xor XOR2 (N2040, N2030, N767);
nor NOR2 (N2041, N2032, N301);
nor NOR2 (N2042, N2040, N1374);
and AND3 (N2043, N2042, N1837, N1197);
and AND3 (N2044, N2026, N664, N1277);
and AND3 (N2045, N2041, N1818, N885);
buf BUF1 (N2046, N2043);
not NOT1 (N2047, N2027);
nand NAND2 (N2048, N2039, N310);
and AND2 (N2049, N2035, N746);
buf BUF1 (N2050, N2046);
and AND2 (N2051, N2044, N1434);
nand NAND4 (N2052, N2031, N1927, N1887, N1005);
nand NAND2 (N2053, N2045, N1308);
nor NOR3 (N2054, N2049, N1827, N1792);
nor NOR4 (N2055, N2050, N915, N2025, N237);
buf BUF1 (N2056, N2047);
buf BUF1 (N2057, N2051);
or OR2 (N2058, N2053, N808);
or OR4 (N2059, N2052, N175, N1505, N233);
not NOT1 (N2060, N2048);
nand NAND2 (N2061, N2021, N874);
xor XOR2 (N2062, N2037, N1755);
nand NAND3 (N2063, N2057, N213, N1979);
buf BUF1 (N2064, N2063);
not NOT1 (N2065, N2054);
buf BUF1 (N2066, N2061);
buf BUF1 (N2067, N2055);
or OR2 (N2068, N2067, N1503);
and AND3 (N2069, N2064, N1191, N458);
not NOT1 (N2070, N2056);
not NOT1 (N2071, N2065);
buf BUF1 (N2072, N2070);
nand NAND3 (N2073, N2062, N494, N458);
nor NOR2 (N2074, N2069, N1369);
xor XOR2 (N2075, N2066, N1792);
xor XOR2 (N2076, N2036, N1130);
nor NOR3 (N2077, N2076, N1165, N540);
and AND4 (N2078, N2068, N228, N626, N2049);
not NOT1 (N2079, N2059);
not NOT1 (N2080, N2074);
nand NAND4 (N2081, N2075, N1175, N1814, N548);
buf BUF1 (N2082, N2072);
buf BUF1 (N2083, N2080);
xor XOR2 (N2084, N2079, N731);
or OR4 (N2085, N2071, N1749, N490, N2031);
not NOT1 (N2086, N2073);
not NOT1 (N2087, N2082);
buf BUF1 (N2088, N2087);
not NOT1 (N2089, N2083);
nand NAND2 (N2090, N2078, N149);
and AND3 (N2091, N2090, N730, N845);
or OR4 (N2092, N2091, N1955, N621, N338);
not NOT1 (N2093, N2081);
and AND4 (N2094, N2085, N1552, N390, N211);
and AND2 (N2095, N2094, N328);
and AND4 (N2096, N2077, N560, N709, N60);
xor XOR2 (N2097, N2060, N1491);
xor XOR2 (N2098, N2089, N406);
and AND3 (N2099, N2095, N1312, N1876);
nor NOR3 (N2100, N2098, N159, N1752);
nand NAND4 (N2101, N2097, N315, N1655, N1923);
nand NAND2 (N2102, N2099, N355);
nor NOR3 (N2103, N2092, N1479, N1729);
not NOT1 (N2104, N2103);
or OR2 (N2105, N2101, N116);
buf BUF1 (N2106, N2086);
xor XOR2 (N2107, N2106, N1608);
nor NOR3 (N2108, N2088, N1723, N1259);
xor XOR2 (N2109, N2058, N1568);
buf BUF1 (N2110, N2093);
or OR2 (N2111, N2084, N1193);
buf BUF1 (N2112, N2110);
nor NOR3 (N2113, N2102, N2029, N442);
nor NOR3 (N2114, N2105, N118, N1331);
buf BUF1 (N2115, N2107);
nor NOR4 (N2116, N2114, N1942, N1468, N514);
not NOT1 (N2117, N2100);
nor NOR4 (N2118, N2113, N82, N588, N1483);
nand NAND3 (N2119, N2118, N1850, N1204);
or OR2 (N2120, N2109, N1984);
not NOT1 (N2121, N2111);
or OR2 (N2122, N2096, N1938);
or OR3 (N2123, N2116, N954, N1994);
nor NOR4 (N2124, N2121, N1588, N339, N1308);
buf BUF1 (N2125, N2122);
or OR4 (N2126, N2119, N1304, N320, N1993);
or OR2 (N2127, N2125, N1994);
not NOT1 (N2128, N2126);
or OR3 (N2129, N2127, N1018, N139);
xor XOR2 (N2130, N2120, N2015);
nor NOR4 (N2131, N2130, N1397, N337, N1151);
buf BUF1 (N2132, N2123);
nor NOR2 (N2133, N2124, N84);
buf BUF1 (N2134, N2117);
and AND3 (N2135, N2108, N1675, N1756);
nor NOR4 (N2136, N2129, N2115, N1129, N1133);
not NOT1 (N2137, N275);
nor NOR2 (N2138, N2134, N1122);
not NOT1 (N2139, N2104);
nand NAND4 (N2140, N2131, N2056, N286, N1057);
or OR2 (N2141, N2138, N1296);
not NOT1 (N2142, N2137);
not NOT1 (N2143, N2128);
buf BUF1 (N2144, N2139);
xor XOR2 (N2145, N2144, N1118);
xor XOR2 (N2146, N2142, N1398);
nand NAND2 (N2147, N2143, N297);
nor NOR4 (N2148, N2112, N1102, N1342, N931);
or OR4 (N2149, N2133, N1933, N1856, N1609);
buf BUF1 (N2150, N2145);
not NOT1 (N2151, N2132);
nor NOR4 (N2152, N2146, N2088, N1222, N1974);
or OR2 (N2153, N2141, N602);
not NOT1 (N2154, N2153);
and AND2 (N2155, N2149, N1179);
nand NAND3 (N2156, N2152, N734, N1256);
nand NAND3 (N2157, N2140, N1503, N542);
nand NAND2 (N2158, N2148, N1533);
xor XOR2 (N2159, N2135, N1357);
nor NOR3 (N2160, N2151, N311, N1900);
buf BUF1 (N2161, N2147);
and AND4 (N2162, N2160, N1308, N556, N1013);
nor NOR3 (N2163, N2155, N2043, N1662);
or OR2 (N2164, N2157, N1056);
and AND4 (N2165, N2136, N936, N756, N1217);
buf BUF1 (N2166, N2165);
or OR3 (N2167, N2163, N1313, N1126);
nor NOR3 (N2168, N2150, N144, N956);
or OR4 (N2169, N2168, N2062, N1444, N1297);
or OR4 (N2170, N2159, N818, N1688, N1159);
and AND4 (N2171, N2158, N1700, N327, N1068);
not NOT1 (N2172, N2162);
nor NOR2 (N2173, N2171, N308);
or OR2 (N2174, N2172, N853);
xor XOR2 (N2175, N2161, N1497);
or OR3 (N2176, N2175, N1276, N1821);
not NOT1 (N2177, N2164);
or OR2 (N2178, N2177, N1099);
and AND3 (N2179, N2173, N1055, N450);
buf BUF1 (N2180, N2176);
xor XOR2 (N2181, N2156, N1167);
buf BUF1 (N2182, N2179);
or OR3 (N2183, N2166, N1257, N1039);
nand NAND3 (N2184, N2183, N366, N2066);
or OR3 (N2185, N2178, N265, N663);
nand NAND4 (N2186, N2154, N1442, N937, N742);
nor NOR4 (N2187, N2186, N2008, N240, N1881);
xor XOR2 (N2188, N2187, N481);
nand NAND2 (N2189, N2167, N1734);
nor NOR2 (N2190, N2170, N1347);
buf BUF1 (N2191, N2188);
nand NAND2 (N2192, N2182, N194);
nor NOR2 (N2193, N2169, N1976);
xor XOR2 (N2194, N2191, N568);
nor NOR4 (N2195, N2190, N1873, N2149, N1218);
or OR2 (N2196, N2194, N633);
buf BUF1 (N2197, N2174);
not NOT1 (N2198, N2184);
not NOT1 (N2199, N2189);
nand NAND2 (N2200, N2180, N494);
xor XOR2 (N2201, N2198, N810);
nor NOR4 (N2202, N2181, N387, N605, N328);
buf BUF1 (N2203, N2185);
buf BUF1 (N2204, N2193);
nand NAND2 (N2205, N2195, N971);
nor NOR2 (N2206, N2197, N2170);
buf BUF1 (N2207, N2200);
and AND2 (N2208, N2203, N1920);
nor NOR3 (N2209, N2207, N2114, N821);
buf BUF1 (N2210, N2205);
buf BUF1 (N2211, N2206);
and AND4 (N2212, N2204, N130, N285, N1992);
buf BUF1 (N2213, N2199);
buf BUF1 (N2214, N2209);
nor NOR3 (N2215, N2202, N370, N622);
xor XOR2 (N2216, N2214, N1419);
not NOT1 (N2217, N2216);
and AND4 (N2218, N2213, N2027, N1486, N2137);
not NOT1 (N2219, N2208);
not NOT1 (N2220, N2215);
nand NAND3 (N2221, N2220, N1670, N1514);
nor NOR4 (N2222, N2218, N1908, N470, N1360);
nand NAND3 (N2223, N2221, N1108, N1990);
buf BUF1 (N2224, N2196);
not NOT1 (N2225, N2210);
nor NOR3 (N2226, N2219, N2124, N510);
buf BUF1 (N2227, N2192);
nand NAND4 (N2228, N2224, N502, N1616, N2063);
nor NOR3 (N2229, N2226, N1949, N2071);
xor XOR2 (N2230, N2227, N1783);
xor XOR2 (N2231, N2217, N196);
nor NOR3 (N2232, N2231, N285, N1024);
and AND3 (N2233, N2223, N1335, N1115);
or OR2 (N2234, N2233, N1103);
or OR3 (N2235, N2201, N890, N867);
xor XOR2 (N2236, N2225, N1390);
nor NOR2 (N2237, N2236, N1869);
nand NAND3 (N2238, N2234, N863, N1757);
xor XOR2 (N2239, N2229, N2069);
nor NOR3 (N2240, N2228, N929, N404);
nor NOR4 (N2241, N2222, N880, N2083, N592);
xor XOR2 (N2242, N2230, N1911);
or OR3 (N2243, N2212, N607, N1042);
nand NAND3 (N2244, N2238, N40, N162);
nor NOR4 (N2245, N2237, N1648, N1706, N1972);
xor XOR2 (N2246, N2242, N1022);
nor NOR2 (N2247, N2246, N2087);
buf BUF1 (N2248, N2247);
buf BUF1 (N2249, N2241);
nor NOR2 (N2250, N2240, N1069);
nand NAND3 (N2251, N2244, N1042, N2101);
buf BUF1 (N2252, N2250);
buf BUF1 (N2253, N2239);
xor XOR2 (N2254, N2211, N1662);
buf BUF1 (N2255, N2243);
buf BUF1 (N2256, N2255);
or OR4 (N2257, N2254, N946, N1830, N1231);
nand NAND4 (N2258, N2235, N363, N1814, N194);
buf BUF1 (N2259, N2253);
or OR3 (N2260, N2249, N479, N1634);
and AND2 (N2261, N2257, N1445);
or OR2 (N2262, N2248, N1780);
and AND4 (N2263, N2261, N1335, N2262, N2070);
xor XOR2 (N2264, N1616, N1487);
nand NAND2 (N2265, N2263, N1432);
buf BUF1 (N2266, N2260);
nand NAND3 (N2267, N2259, N697, N861);
nand NAND2 (N2268, N2232, N1068);
buf BUF1 (N2269, N2245);
nand NAND4 (N2270, N2258, N27, N398, N178);
not NOT1 (N2271, N2269);
nand NAND3 (N2272, N2256, N1799, N1858);
not NOT1 (N2273, N2265);
nor NOR3 (N2274, N2270, N1412, N2269);
buf BUF1 (N2275, N2272);
buf BUF1 (N2276, N2274);
buf BUF1 (N2277, N2267);
nor NOR4 (N2278, N2271, N2230, N174, N709);
nand NAND2 (N2279, N2268, N2171);
xor XOR2 (N2280, N2273, N1872);
and AND2 (N2281, N2278, N1279);
nor NOR2 (N2282, N2280, N395);
buf BUF1 (N2283, N2279);
xor XOR2 (N2284, N2275, N925);
xor XOR2 (N2285, N2276, N1993);
nand NAND4 (N2286, N2281, N2008, N2189, N391);
and AND2 (N2287, N2286, N400);
nor NOR3 (N2288, N2285, N1592, N1851);
and AND4 (N2289, N2277, N950, N1987, N2132);
not NOT1 (N2290, N2266);
xor XOR2 (N2291, N2284, N1345);
and AND3 (N2292, N2290, N747, N2259);
buf BUF1 (N2293, N2292);
not NOT1 (N2294, N2283);
buf BUF1 (N2295, N2251);
and AND2 (N2296, N2295, N1750);
not NOT1 (N2297, N2252);
nand NAND2 (N2298, N2288, N711);
and AND4 (N2299, N2296, N1791, N2284, N694);
nor NOR4 (N2300, N2264, N599, N1495, N1528);
or OR2 (N2301, N2293, N1507);
and AND2 (N2302, N2294, N2158);
not NOT1 (N2303, N2291);
xor XOR2 (N2304, N2297, N1903);
not NOT1 (N2305, N2299);
nand NAND2 (N2306, N2302, N1587);
nor NOR4 (N2307, N2306, N1255, N690, N2278);
buf BUF1 (N2308, N2300);
xor XOR2 (N2309, N2305, N461);
buf BUF1 (N2310, N2298);
not NOT1 (N2311, N2301);
nand NAND3 (N2312, N2311, N541, N582);
not NOT1 (N2313, N2310);
buf BUF1 (N2314, N2303);
nor NOR2 (N2315, N2309, N423);
and AND2 (N2316, N2289, N1415);
buf BUF1 (N2317, N2315);
and AND2 (N2318, N2316, N1255);
buf BUF1 (N2319, N2282);
or OR2 (N2320, N2319, N751);
not NOT1 (N2321, N2304);
nor NOR2 (N2322, N2314, N1433);
nor NOR3 (N2323, N2322, N1839, N1846);
not NOT1 (N2324, N2308);
or OR3 (N2325, N2312, N57, N377);
nor NOR2 (N2326, N2321, N309);
and AND3 (N2327, N2320, N541, N429);
xor XOR2 (N2328, N2307, N998);
not NOT1 (N2329, N2317);
or OR4 (N2330, N2325, N1355, N811, N1924);
nor NOR4 (N2331, N2329, N839, N1145, N475);
nor NOR2 (N2332, N2287, N2171);
buf BUF1 (N2333, N2332);
not NOT1 (N2334, N2330);
not NOT1 (N2335, N2318);
not NOT1 (N2336, N2323);
not NOT1 (N2337, N2313);
and AND4 (N2338, N2333, N2188, N772, N1179);
xor XOR2 (N2339, N2334, N677);
xor XOR2 (N2340, N2335, N1325);
or OR2 (N2341, N2328, N1586);
and AND2 (N2342, N2340, N761);
not NOT1 (N2343, N2327);
buf BUF1 (N2344, N2324);
nor NOR2 (N2345, N2337, N1772);
xor XOR2 (N2346, N2331, N74);
not NOT1 (N2347, N2343);
xor XOR2 (N2348, N2344, N1263);
not NOT1 (N2349, N2345);
nand NAND4 (N2350, N2341, N644, N1346, N1829);
buf BUF1 (N2351, N2346);
nor NOR2 (N2352, N2339, N290);
xor XOR2 (N2353, N2350, N1148);
not NOT1 (N2354, N2352);
nand NAND3 (N2355, N2353, N1767, N1821);
or OR2 (N2356, N2348, N287);
not NOT1 (N2357, N2351);
buf BUF1 (N2358, N2342);
buf BUF1 (N2359, N2355);
xor XOR2 (N2360, N2358, N1745);
or OR4 (N2361, N2326, N624, N1317, N812);
buf BUF1 (N2362, N2336);
or OR3 (N2363, N2347, N799, N685);
nand NAND3 (N2364, N2362, N2297, N1204);
buf BUF1 (N2365, N2363);
or OR4 (N2366, N2356, N1567, N2240, N1011);
not NOT1 (N2367, N2338);
buf BUF1 (N2368, N2359);
nor NOR3 (N2369, N2354, N432, N2183);
buf BUF1 (N2370, N2365);
nor NOR3 (N2371, N2366, N562, N795);
xor XOR2 (N2372, N2369, N1160);
or OR4 (N2373, N2349, N1146, N993, N98);
xor XOR2 (N2374, N2367, N102);
not NOT1 (N2375, N2374);
nor NOR4 (N2376, N2370, N358, N324, N2005);
xor XOR2 (N2377, N2364, N336);
not NOT1 (N2378, N2375);
nor NOR2 (N2379, N2372, N1276);
buf BUF1 (N2380, N2361);
not NOT1 (N2381, N2368);
or OR4 (N2382, N2378, N287, N1104, N2143);
xor XOR2 (N2383, N2376, N1502);
not NOT1 (N2384, N2360);
xor XOR2 (N2385, N2380, N1713);
xor XOR2 (N2386, N2383, N1176);
buf BUF1 (N2387, N2377);
nor NOR2 (N2388, N2382, N511);
xor XOR2 (N2389, N2386, N2129);
buf BUF1 (N2390, N2373);
and AND3 (N2391, N2389, N1920, N88);
and AND4 (N2392, N2387, N168, N1163, N1378);
buf BUF1 (N2393, N2379);
and AND4 (N2394, N2393, N1590, N1448, N1098);
xor XOR2 (N2395, N2388, N202);
buf BUF1 (N2396, N2392);
buf BUF1 (N2397, N2371);
and AND2 (N2398, N2391, N816);
nand NAND4 (N2399, N2396, N2157, N1930, N1739);
or OR3 (N2400, N2357, N739, N1768);
xor XOR2 (N2401, N2400, N473);
and AND4 (N2402, N2390, N1665, N193, N2258);
buf BUF1 (N2403, N2398);
nor NOR4 (N2404, N2402, N453, N29, N1515);
xor XOR2 (N2405, N2384, N637);
or OR3 (N2406, N2395, N700, N624);
not NOT1 (N2407, N2381);
or OR3 (N2408, N2406, N162, N163);
nand NAND2 (N2409, N2405, N415);
buf BUF1 (N2410, N2399);
and AND4 (N2411, N2385, N863, N95, N2390);
or OR3 (N2412, N2394, N803, N2314);
not NOT1 (N2413, N2403);
or OR2 (N2414, N2408, N583);
buf BUF1 (N2415, N2412);
and AND4 (N2416, N2411, N787, N2133, N2017);
nand NAND4 (N2417, N2413, N1708, N78, N229);
not NOT1 (N2418, N2414);
buf BUF1 (N2419, N2409);
not NOT1 (N2420, N2407);
not NOT1 (N2421, N2417);
nor NOR3 (N2422, N2415, N866, N2225);
not NOT1 (N2423, N2404);
nor NOR2 (N2424, N2401, N1583);
buf BUF1 (N2425, N2424);
or OR3 (N2426, N2422, N869, N1141);
nor NOR3 (N2427, N2397, N32, N907);
nand NAND4 (N2428, N2427, N554, N2033, N107);
not NOT1 (N2429, N2418);
or OR3 (N2430, N2423, N681, N2156);
or OR3 (N2431, N2428, N1322, N2293);
or OR3 (N2432, N2429, N2302, N1251);
xor XOR2 (N2433, N2421, N2427);
and AND2 (N2434, N2419, N1533);
or OR2 (N2435, N2434, N1977);
nand NAND4 (N2436, N2430, N390, N80, N2156);
buf BUF1 (N2437, N2426);
and AND2 (N2438, N2433, N399);
or OR3 (N2439, N2420, N972, N2392);
and AND3 (N2440, N2432, N912, N991);
xor XOR2 (N2441, N2436, N503);
buf BUF1 (N2442, N2425);
or OR2 (N2443, N2416, N321);
not NOT1 (N2444, N2410);
nor NOR4 (N2445, N2437, N2390, N611, N1774);
buf BUF1 (N2446, N2442);
or OR2 (N2447, N2435, N483);
and AND2 (N2448, N2440, N686);
or OR3 (N2449, N2439, N589, N1099);
and AND3 (N2450, N2447, N481, N739);
buf BUF1 (N2451, N2441);
xor XOR2 (N2452, N2443, N566);
nand NAND4 (N2453, N2444, N1489, N1316, N1150);
nor NOR2 (N2454, N2438, N2013);
xor XOR2 (N2455, N2446, N1344);
or OR3 (N2456, N2454, N855, N109);
nand NAND4 (N2457, N2452, N1306, N49, N1053);
and AND3 (N2458, N2453, N1755, N1951);
nand NAND2 (N2459, N2451, N410);
and AND4 (N2460, N2449, N1611, N1355, N28);
xor XOR2 (N2461, N2457, N1478);
xor XOR2 (N2462, N2459, N764);
or OR2 (N2463, N2445, N566);
or OR4 (N2464, N2456, N1148, N559, N1918);
buf BUF1 (N2465, N2464);
or OR3 (N2466, N2458, N1227, N1233);
and AND4 (N2467, N2460, N877, N602, N734);
buf BUF1 (N2468, N2465);
nand NAND4 (N2469, N2448, N493, N1459, N2233);
nand NAND4 (N2470, N2469, N2427, N2325, N1305);
not NOT1 (N2471, N2455);
buf BUF1 (N2472, N2470);
not NOT1 (N2473, N2461);
nand NAND3 (N2474, N2431, N542, N1914);
xor XOR2 (N2475, N2462, N2081);
not NOT1 (N2476, N2475);
nand NAND4 (N2477, N2476, N2380, N1045, N1068);
and AND4 (N2478, N2473, N1839, N1463, N203);
xor XOR2 (N2479, N2468, N23);
not NOT1 (N2480, N2463);
or OR4 (N2481, N2480, N2153, N2304, N2305);
nand NAND3 (N2482, N2472, N1238, N2140);
nor NOR3 (N2483, N2482, N2301, N1336);
not NOT1 (N2484, N2466);
or OR4 (N2485, N2477, N1170, N1885, N48);
or OR3 (N2486, N2481, N1020, N727);
and AND2 (N2487, N2484, N711);
xor XOR2 (N2488, N2450, N190);
or OR4 (N2489, N2479, N45, N1680, N2190);
buf BUF1 (N2490, N2489);
or OR2 (N2491, N2471, N747);
nand NAND2 (N2492, N2485, N1624);
buf BUF1 (N2493, N2486);
not NOT1 (N2494, N2492);
or OR2 (N2495, N2483, N1594);
not NOT1 (N2496, N2490);
buf BUF1 (N2497, N2478);
xor XOR2 (N2498, N2491, N2382);
or OR3 (N2499, N2467, N1610, N889);
not NOT1 (N2500, N2498);
nand NAND3 (N2501, N2488, N45, N1086);
not NOT1 (N2502, N2474);
or OR4 (N2503, N2493, N1189, N2147, N90);
and AND3 (N2504, N2502, N1639, N592);
nor NOR4 (N2505, N2504, N939, N1175, N1383);
or OR4 (N2506, N2505, N1963, N1480, N1501);
nor NOR4 (N2507, N2495, N1188, N2170, N2153);
nand NAND2 (N2508, N2506, N73);
nor NOR3 (N2509, N2500, N1494, N1475);
not NOT1 (N2510, N2503);
and AND2 (N2511, N2499, N1435);
and AND4 (N2512, N2510, N965, N1225, N1791);
nand NAND4 (N2513, N2512, N1482, N1252, N586);
buf BUF1 (N2514, N2513);
and AND3 (N2515, N2497, N49, N575);
xor XOR2 (N2516, N2514, N1234);
or OR2 (N2517, N2509, N1740);
not NOT1 (N2518, N2511);
nor NOR3 (N2519, N2507, N1600, N2039);
or OR2 (N2520, N2494, N528);
nor NOR4 (N2521, N2487, N1114, N740, N1140);
xor XOR2 (N2522, N2501, N2155);
or OR3 (N2523, N2522, N2302, N2421);
nor NOR3 (N2524, N2521, N1496, N57);
nor NOR4 (N2525, N2515, N272, N1288, N1903);
not NOT1 (N2526, N2520);
and AND4 (N2527, N2516, N1035, N1528, N1214);
buf BUF1 (N2528, N2524);
xor XOR2 (N2529, N2496, N920);
not NOT1 (N2530, N2519);
nand NAND3 (N2531, N2518, N157, N1558);
and AND4 (N2532, N2530, N1477, N1014, N2111);
not NOT1 (N2533, N2508);
nor NOR2 (N2534, N2526, N446);
nor NOR3 (N2535, N2523, N935, N1350);
and AND2 (N2536, N2533, N1736);
not NOT1 (N2537, N2532);
nand NAND3 (N2538, N2535, N878, N2500);
buf BUF1 (N2539, N2528);
and AND4 (N2540, N2537, N790, N396, N1932);
xor XOR2 (N2541, N2540, N856);
xor XOR2 (N2542, N2517, N1384);
nor NOR2 (N2543, N2539, N58);
nor NOR2 (N2544, N2531, N70);
nor NOR3 (N2545, N2544, N1522, N1792);
nor NOR2 (N2546, N2534, N2243);
not NOT1 (N2547, N2545);
buf BUF1 (N2548, N2527);
nand NAND2 (N2549, N2542, N1816);
and AND3 (N2550, N2525, N1348, N1574);
xor XOR2 (N2551, N2548, N2523);
and AND2 (N2552, N2550, N1644);
or OR4 (N2553, N2529, N278, N2198, N1200);
nand NAND2 (N2554, N2549, N1551);
nor NOR4 (N2555, N2551, N533, N342, N923);
not NOT1 (N2556, N2536);
or OR3 (N2557, N2538, N1346, N2056);
nor NOR3 (N2558, N2543, N732, N88);
or OR4 (N2559, N2552, N553, N1163, N1052);
xor XOR2 (N2560, N2556, N2359);
buf BUF1 (N2561, N2558);
nor NOR3 (N2562, N2541, N767, N2135);
and AND4 (N2563, N2553, N2048, N800, N1402);
nand NAND3 (N2564, N2546, N1174, N2253);
nor NOR3 (N2565, N2563, N1413, N1766);
xor XOR2 (N2566, N2555, N1004);
buf BUF1 (N2567, N2565);
or OR2 (N2568, N2547, N701);
nand NAND2 (N2569, N2560, N1130);
or OR2 (N2570, N2567, N2364);
nor NOR2 (N2571, N2561, N971);
nand NAND2 (N2572, N2569, N368);
or OR4 (N2573, N2566, N2070, N1786, N591);
nand NAND4 (N2574, N2562, N1060, N1989, N369);
nor NOR2 (N2575, N2574, N2440);
nor NOR4 (N2576, N2572, N2107, N2554, N2518);
nor NOR3 (N2577, N2072, N1792, N1072);
buf BUF1 (N2578, N2577);
nand NAND4 (N2579, N2571, N1397, N235, N200);
xor XOR2 (N2580, N2578, N2371);
nand NAND4 (N2581, N2559, N1830, N1542, N2334);
buf BUF1 (N2582, N2575);
or OR3 (N2583, N2570, N325, N384);
and AND3 (N2584, N2576, N219, N2544);
buf BUF1 (N2585, N2557);
xor XOR2 (N2586, N2584, N2351);
nand NAND4 (N2587, N2568, N444, N826, N311);
and AND2 (N2588, N2564, N236);
buf BUF1 (N2589, N2580);
or OR4 (N2590, N2587, N182, N1594, N2040);
not NOT1 (N2591, N2581);
or OR2 (N2592, N2585, N1046);
nor NOR4 (N2593, N2589, N1991, N2248, N1609);
nand NAND2 (N2594, N2590, N584);
or OR4 (N2595, N2594, N700, N2265, N1164);
xor XOR2 (N2596, N2579, N1719);
or OR2 (N2597, N2586, N346);
or OR3 (N2598, N2591, N2427, N1975);
buf BUF1 (N2599, N2582);
buf BUF1 (N2600, N2583);
nor NOR4 (N2601, N2588, N1690, N2451, N1640);
and AND2 (N2602, N2573, N933);
xor XOR2 (N2603, N2600, N752);
nand NAND4 (N2604, N2603, N579, N426, N1172);
nand NAND3 (N2605, N2592, N1299, N2129);
buf BUF1 (N2606, N2599);
and AND2 (N2607, N2602, N1514);
nand NAND4 (N2608, N2598, N2582, N1208, N112);
and AND4 (N2609, N2607, N386, N1421, N936);
or OR3 (N2610, N2595, N1451, N551);
or OR2 (N2611, N2610, N2284);
and AND3 (N2612, N2597, N1607, N2173);
xor XOR2 (N2613, N2604, N981);
nand NAND3 (N2614, N2612, N664, N741);
nor NOR3 (N2615, N2605, N1709, N1931);
or OR3 (N2616, N2613, N1493, N999);
and AND2 (N2617, N2609, N1566);
not NOT1 (N2618, N2611);
buf BUF1 (N2619, N2593);
nand NAND4 (N2620, N2608, N1009, N2604, N1174);
xor XOR2 (N2621, N2615, N2255);
or OR4 (N2622, N2614, N521, N1455, N1065);
nor NOR4 (N2623, N2617, N36, N2316, N1924);
xor XOR2 (N2624, N2623, N1428);
buf BUF1 (N2625, N2621);
nor NOR4 (N2626, N2624, N556, N1448, N1708);
nand NAND4 (N2627, N2622, N507, N510, N1799);
buf BUF1 (N2628, N2606);
nand NAND2 (N2629, N2601, N1258);
not NOT1 (N2630, N2627);
or OR2 (N2631, N2619, N1728);
or OR4 (N2632, N2628, N597, N91, N2089);
xor XOR2 (N2633, N2632, N105);
buf BUF1 (N2634, N2629);
nand NAND2 (N2635, N2634, N576);
buf BUF1 (N2636, N2626);
not NOT1 (N2637, N2636);
xor XOR2 (N2638, N2620, N1553);
xor XOR2 (N2639, N2631, N2111);
or OR4 (N2640, N2633, N1310, N692, N1445);
buf BUF1 (N2641, N2639);
nand NAND2 (N2642, N2618, N2277);
buf BUF1 (N2643, N2616);
not NOT1 (N2644, N2641);
buf BUF1 (N2645, N2644);
or OR4 (N2646, N2637, N616, N2407, N1958);
xor XOR2 (N2647, N2643, N666);
and AND2 (N2648, N2645, N1466);
nand NAND3 (N2649, N2642, N1947, N2483);
buf BUF1 (N2650, N2596);
xor XOR2 (N2651, N2635, N1153);
not NOT1 (N2652, N2640);
or OR3 (N2653, N2648, N306, N1975);
nor NOR2 (N2654, N2653, N8);
xor XOR2 (N2655, N2646, N1681);
or OR4 (N2656, N2649, N148, N1832, N1246);
or OR3 (N2657, N2652, N1624, N184);
and AND4 (N2658, N2625, N171, N2087, N2383);
nand NAND4 (N2659, N2658, N1431, N60, N2327);
or OR4 (N2660, N2650, N2467, N1019, N1388);
not NOT1 (N2661, N2638);
nand NAND4 (N2662, N2647, N1335, N54, N1870);
and AND2 (N2663, N2656, N1741);
nor NOR2 (N2664, N2662, N2598);
buf BUF1 (N2665, N2661);
nor NOR4 (N2666, N2660, N1636, N233, N483);
nand NAND2 (N2667, N2663, N2663);
or OR2 (N2668, N2657, N2585);
or OR4 (N2669, N2665, N612, N1513, N1316);
and AND4 (N2670, N2654, N1001, N594, N909);
nor NOR2 (N2671, N2666, N634);
and AND2 (N2672, N2655, N1672);
nor NOR2 (N2673, N2667, N629);
xor XOR2 (N2674, N2670, N936);
not NOT1 (N2675, N2659);
nand NAND2 (N2676, N2673, N2009);
xor XOR2 (N2677, N2676, N1678);
xor XOR2 (N2678, N2669, N2486);
xor XOR2 (N2679, N2678, N122);
xor XOR2 (N2680, N2672, N633);
nor NOR2 (N2681, N2664, N1702);
not NOT1 (N2682, N2668);
nand NAND3 (N2683, N2630, N184, N1004);
xor XOR2 (N2684, N2679, N1368);
buf BUF1 (N2685, N2683);
not NOT1 (N2686, N2671);
and AND4 (N2687, N2677, N274, N618, N1953);
not NOT1 (N2688, N2680);
or OR2 (N2689, N2682, N1357);
and AND4 (N2690, N2684, N1279, N2013, N651);
nor NOR3 (N2691, N2675, N1792, N87);
nor NOR2 (N2692, N2688, N1554);
nand NAND3 (N2693, N2681, N2244, N234);
buf BUF1 (N2694, N2692);
not NOT1 (N2695, N2685);
nand NAND2 (N2696, N2686, N1134);
nor NOR2 (N2697, N2690, N222);
nor NOR3 (N2698, N2695, N2012, N510);
not NOT1 (N2699, N2698);
nand NAND4 (N2700, N2689, N425, N1388, N2270);
nor NOR2 (N2701, N2691, N793);
nor NOR2 (N2702, N2694, N1558);
xor XOR2 (N2703, N2702, N2248);
nor NOR4 (N2704, N2687, N2578, N723, N1600);
xor XOR2 (N2705, N2703, N1106);
nand NAND2 (N2706, N2696, N2383);
nor NOR4 (N2707, N2705, N435, N629, N1690);
nand NAND3 (N2708, N2701, N7, N2032);
and AND3 (N2709, N2651, N898, N2174);
and AND3 (N2710, N2699, N2664, N835);
buf BUF1 (N2711, N2704);
nor NOR2 (N2712, N2711, N428);
nor NOR4 (N2713, N2710, N565, N2547, N417);
nand NAND3 (N2714, N2697, N137, N2360);
xor XOR2 (N2715, N2700, N1467);
not NOT1 (N2716, N2714);
and AND4 (N2717, N2709, N2317, N2077, N662);
xor XOR2 (N2718, N2716, N1054);
or OR4 (N2719, N2707, N176, N984, N2683);
buf BUF1 (N2720, N2693);
buf BUF1 (N2721, N2708);
nor NOR2 (N2722, N2706, N1159);
xor XOR2 (N2723, N2719, N1008);
or OR4 (N2724, N2720, N990, N1469, N2272);
buf BUF1 (N2725, N2717);
not NOT1 (N2726, N2722);
or OR2 (N2727, N2721, N1006);
nand NAND2 (N2728, N2712, N2340);
not NOT1 (N2729, N2725);
xor XOR2 (N2730, N2674, N2552);
xor XOR2 (N2731, N2726, N490);
not NOT1 (N2732, N2730);
or OR3 (N2733, N2724, N1970, N1722);
nor NOR3 (N2734, N2731, N1401, N2114);
and AND4 (N2735, N2728, N2306, N321, N1390);
nand NAND4 (N2736, N2727, N2058, N380, N2094);
not NOT1 (N2737, N2732);
xor XOR2 (N2738, N2715, N2524);
buf BUF1 (N2739, N2735);
not NOT1 (N2740, N2718);
nand NAND2 (N2741, N2723, N420);
and AND2 (N2742, N2741, N2171);
nor NOR4 (N2743, N2739, N726, N1651, N1738);
nand NAND3 (N2744, N2734, N722, N2030);
not NOT1 (N2745, N2738);
buf BUF1 (N2746, N2745);
nand NAND2 (N2747, N2713, N2447);
and AND4 (N2748, N2737, N2011, N2472, N1089);
and AND3 (N2749, N2729, N1927, N1603);
buf BUF1 (N2750, N2744);
nor NOR4 (N2751, N2742, N766, N1429, N311);
buf BUF1 (N2752, N2743);
and AND3 (N2753, N2752, N1974, N1117);
xor XOR2 (N2754, N2736, N1129);
xor XOR2 (N2755, N2733, N1713);
buf BUF1 (N2756, N2749);
not NOT1 (N2757, N2753);
or OR4 (N2758, N2756, N1759, N1459, N2232);
buf BUF1 (N2759, N2746);
nand NAND4 (N2760, N2757, N767, N398, N1172);
buf BUF1 (N2761, N2751);
xor XOR2 (N2762, N2747, N1538);
xor XOR2 (N2763, N2758, N1709);
buf BUF1 (N2764, N2755);
nand NAND3 (N2765, N2748, N280, N2);
not NOT1 (N2766, N2765);
nand NAND4 (N2767, N2762, N1310, N37, N2665);
xor XOR2 (N2768, N2754, N1964);
buf BUF1 (N2769, N2766);
and AND4 (N2770, N2740, N260, N1634, N2173);
buf BUF1 (N2771, N2769);
and AND4 (N2772, N2767, N463, N1121, N788);
nand NAND3 (N2773, N2750, N2531, N1133);
nand NAND2 (N2774, N2768, N1015);
or OR4 (N2775, N2774, N1646, N2429, N2426);
nand NAND2 (N2776, N2760, N1834);
and AND4 (N2777, N2770, N2077, N442, N970);
or OR2 (N2778, N2773, N1545);
xor XOR2 (N2779, N2772, N1420);
not NOT1 (N2780, N2771);
and AND3 (N2781, N2777, N2779, N2480);
or OR2 (N2782, N630, N392);
not NOT1 (N2783, N2776);
nand NAND2 (N2784, N2778, N1935);
buf BUF1 (N2785, N2782);
and AND3 (N2786, N2764, N2608, N1732);
nor NOR3 (N2787, N2786, N1470, N2330);
nand NAND2 (N2788, N2775, N2277);
buf BUF1 (N2789, N2787);
buf BUF1 (N2790, N2759);
nor NOR2 (N2791, N2785, N1089);
xor XOR2 (N2792, N2783, N106);
nand NAND3 (N2793, N2763, N2277, N1489);
nor NOR4 (N2794, N2793, N1935, N2661, N1346);
or OR2 (N2795, N2761, N853);
or OR2 (N2796, N2784, N169);
or OR2 (N2797, N2781, N1313);
or OR2 (N2798, N2791, N2664);
buf BUF1 (N2799, N2797);
nand NAND4 (N2800, N2789, N452, N1973, N775);
nor NOR4 (N2801, N2788, N2753, N1739, N1303);
xor XOR2 (N2802, N2792, N1512);
or OR3 (N2803, N2802, N1411, N259);
xor XOR2 (N2804, N2796, N905);
nand NAND4 (N2805, N2803, N1264, N1615, N1080);
not NOT1 (N2806, N2790);
or OR2 (N2807, N2804, N2213);
or OR4 (N2808, N2801, N2193, N2622, N682);
and AND4 (N2809, N2799, N78, N1946, N1311);
nor NOR3 (N2810, N2800, N869, N2717);
and AND4 (N2811, N2794, N1790, N314, N1427);
xor XOR2 (N2812, N2780, N2352);
and AND4 (N2813, N2812, N877, N300, N2586);
not NOT1 (N2814, N2810);
not NOT1 (N2815, N2798);
xor XOR2 (N2816, N2815, N303);
buf BUF1 (N2817, N2795);
not NOT1 (N2818, N2806);
buf BUF1 (N2819, N2805);
buf BUF1 (N2820, N2817);
nand NAND2 (N2821, N2807, N1861);
nand NAND3 (N2822, N2816, N945, N1036);
xor XOR2 (N2823, N2821, N2648);
nor NOR4 (N2824, N2822, N97, N1823, N1658);
buf BUF1 (N2825, N2824);
nor NOR3 (N2826, N2809, N1056, N668);
xor XOR2 (N2827, N2823, N912);
and AND3 (N2828, N2813, N799, N45);
buf BUF1 (N2829, N2808);
not NOT1 (N2830, N2827);
xor XOR2 (N2831, N2826, N2457);
or OR3 (N2832, N2820, N2240, N2013);
and AND2 (N2833, N2832, N1667);
and AND3 (N2834, N2811, N2600, N828);
not NOT1 (N2835, N2818);
not NOT1 (N2836, N2831);
or OR3 (N2837, N2829, N2489, N2017);
xor XOR2 (N2838, N2819, N544);
and AND2 (N2839, N2828, N1794);
nor NOR2 (N2840, N2814, N165);
or OR4 (N2841, N2834, N1239, N1836, N2713);
xor XOR2 (N2842, N2837, N2230);
nor NOR4 (N2843, N2836, N1488, N458, N738);
not NOT1 (N2844, N2839);
buf BUF1 (N2845, N2843);
xor XOR2 (N2846, N2844, N1476);
and AND3 (N2847, N2842, N823, N1331);
nor NOR4 (N2848, N2835, N1547, N244, N1850);
and AND2 (N2849, N2845, N2540);
not NOT1 (N2850, N2847);
nor NOR3 (N2851, N2838, N1876, N1880);
nand NAND3 (N2852, N2846, N793, N1703);
and AND4 (N2853, N2833, N1962, N466, N1890);
or OR4 (N2854, N2850, N745, N1162, N172);
not NOT1 (N2855, N2848);
nor NOR4 (N2856, N2825, N2079, N489, N1904);
nand NAND4 (N2857, N2849, N1991, N2159, N2184);
not NOT1 (N2858, N2852);
nor NOR2 (N2859, N2851, N2755);
nand NAND4 (N2860, N2856, N1288, N1047, N129);
or OR2 (N2861, N2853, N1473);
nor NOR3 (N2862, N2840, N2807, N712);
and AND4 (N2863, N2859, N1886, N744, N2443);
not NOT1 (N2864, N2858);
nor NOR3 (N2865, N2830, N1414, N590);
xor XOR2 (N2866, N2865, N1654);
and AND3 (N2867, N2857, N1491, N1611);
or OR4 (N2868, N2864, N427, N1692, N25);
nor NOR3 (N2869, N2854, N69, N1373);
or OR4 (N2870, N2866, N1332, N1015, N1049);
buf BUF1 (N2871, N2863);
and AND3 (N2872, N2871, N2123, N1816);
not NOT1 (N2873, N2872);
or OR4 (N2874, N2861, N2411, N1483, N1270);
xor XOR2 (N2875, N2855, N1625);
not NOT1 (N2876, N2870);
or OR3 (N2877, N2873, N1105, N658);
xor XOR2 (N2878, N2876, N2787);
and AND3 (N2879, N2877, N1451, N588);
and AND4 (N2880, N2841, N815, N1381, N630);
nor NOR3 (N2881, N2860, N1246, N1119);
nand NAND4 (N2882, N2880, N1039, N1689, N1723);
nand NAND3 (N2883, N2862, N2562, N2433);
nand NAND4 (N2884, N2878, N997, N2497, N2795);
nand NAND2 (N2885, N2868, N2538);
nor NOR4 (N2886, N2885, N240, N370, N818);
buf BUF1 (N2887, N2874);
or OR2 (N2888, N2875, N2312);
or OR2 (N2889, N2888, N638);
xor XOR2 (N2890, N2884, N1729);
buf BUF1 (N2891, N2887);
nand NAND3 (N2892, N2882, N2877, N903);
buf BUF1 (N2893, N2883);
not NOT1 (N2894, N2886);
buf BUF1 (N2895, N2894);
not NOT1 (N2896, N2879);
xor XOR2 (N2897, N2891, N1398);
or OR4 (N2898, N2889, N2086, N1585, N2481);
nand NAND3 (N2899, N2890, N2356, N857);
buf BUF1 (N2900, N2892);
not NOT1 (N2901, N2900);
xor XOR2 (N2902, N2895, N789);
or OR3 (N2903, N2896, N1480, N223);
nand NAND4 (N2904, N2898, N1556, N2561, N2700);
and AND3 (N2905, N2893, N2317, N218);
not NOT1 (N2906, N2905);
and AND2 (N2907, N2902, N1640);
nor NOR4 (N2908, N2867, N1614, N381, N506);
nor NOR3 (N2909, N2899, N1995, N1508);
not NOT1 (N2910, N2907);
nor NOR4 (N2911, N2903, N2045, N954, N1820);
nor NOR2 (N2912, N2910, N1735);
not NOT1 (N2913, N2908);
nand NAND4 (N2914, N2901, N1385, N349, N2252);
and AND3 (N2915, N2914, N2154, N136);
and AND4 (N2916, N2909, N1421, N2761, N681);
buf BUF1 (N2917, N2906);
and AND2 (N2918, N2911, N513);
buf BUF1 (N2919, N2917);
not NOT1 (N2920, N2918);
or OR4 (N2921, N2919, N2117, N89, N973);
and AND4 (N2922, N2912, N2763, N2723, N1277);
xor XOR2 (N2923, N2897, N2383);
nor NOR3 (N2924, N2904, N111, N269);
not NOT1 (N2925, N2869);
and AND4 (N2926, N2881, N417, N1714, N2648);
xor XOR2 (N2927, N2924, N1933);
not NOT1 (N2928, N2915);
nor NOR2 (N2929, N2916, N1179);
not NOT1 (N2930, N2922);
buf BUF1 (N2931, N2921);
nand NAND2 (N2932, N2923, N52);
nand NAND2 (N2933, N2930, N870);
nor NOR4 (N2934, N2933, N2508, N2771, N1009);
nand NAND3 (N2935, N2920, N973, N1718);
not NOT1 (N2936, N2913);
or OR3 (N2937, N2926, N625, N2323);
and AND3 (N2938, N2927, N1922, N702);
xor XOR2 (N2939, N2931, N2032);
nand NAND2 (N2940, N2934, N2822);
and AND4 (N2941, N2940, N479, N2917, N1258);
buf BUF1 (N2942, N2935);
xor XOR2 (N2943, N2937, N327);
nor NOR4 (N2944, N2932, N2466, N501, N1688);
or OR4 (N2945, N2941, N2521, N1489, N156);
xor XOR2 (N2946, N2936, N2282);
xor XOR2 (N2947, N2925, N1080);
buf BUF1 (N2948, N2929);
or OR4 (N2949, N2945, N2518, N573, N2450);
nor NOR3 (N2950, N2942, N2646, N390);
and AND3 (N2951, N2944, N984, N2591);
or OR2 (N2952, N2946, N2457);
or OR3 (N2953, N2928, N2383, N1837);
buf BUF1 (N2954, N2948);
nor NOR4 (N2955, N2953, N1704, N1949, N2854);
not NOT1 (N2956, N2950);
nand NAND3 (N2957, N2947, N282, N1645);
nand NAND2 (N2958, N2954, N1290);
nand NAND3 (N2959, N2938, N853, N2866);
buf BUF1 (N2960, N2952);
nor NOR4 (N2961, N2957, N740, N633, N2250);
nor NOR3 (N2962, N2958, N1342, N815);
buf BUF1 (N2963, N2959);
buf BUF1 (N2964, N2955);
buf BUF1 (N2965, N2951);
nor NOR2 (N2966, N2949, N1521);
xor XOR2 (N2967, N2965, N1858);
nand NAND3 (N2968, N2961, N2060, N2378);
not NOT1 (N2969, N2960);
nor NOR2 (N2970, N2963, N1581);
nor NOR2 (N2971, N2967, N2116);
xor XOR2 (N2972, N2943, N1082);
xor XOR2 (N2973, N2970, N1213);
buf BUF1 (N2974, N2969);
buf BUF1 (N2975, N2972);
or OR4 (N2976, N2939, N777, N1610, N2862);
or OR3 (N2977, N2974, N2846, N2717);
nor NOR3 (N2978, N2962, N2433, N2942);
nand NAND2 (N2979, N2977, N1107);
or OR4 (N2980, N2964, N2338, N1642, N230);
xor XOR2 (N2981, N2971, N2440);
buf BUF1 (N2982, N2978);
and AND2 (N2983, N2979, N2322);
buf BUF1 (N2984, N2975);
buf BUF1 (N2985, N2966);
xor XOR2 (N2986, N2956, N732);
nand NAND3 (N2987, N2986, N961, N2396);
not NOT1 (N2988, N2984);
or OR2 (N2989, N2981, N1194);
xor XOR2 (N2990, N2985, N1776);
not NOT1 (N2991, N2982);
or OR2 (N2992, N2983, N2783);
or OR3 (N2993, N2992, N2695, N433);
or OR4 (N2994, N2976, N1256, N2343, N296);
and AND2 (N2995, N2990, N450);
xor XOR2 (N2996, N2973, N2579);
buf BUF1 (N2997, N2989);
nand NAND4 (N2998, N2997, N2873, N1566, N2630);
or OR2 (N2999, N2996, N766);
not NOT1 (N3000, N2993);
nor NOR4 (N3001, N2999, N1116, N1706, N1907);
and AND4 (N3002, N2987, N848, N2792, N1393);
nor NOR3 (N3003, N2998, N758, N2898);
not NOT1 (N3004, N2988);
or OR4 (N3005, N3000, N1479, N1111, N2819);
xor XOR2 (N3006, N2991, N2327);
not NOT1 (N3007, N2994);
buf BUF1 (N3008, N3001);
buf BUF1 (N3009, N3002);
nor NOR4 (N3010, N2968, N2209, N185, N1016);
nor NOR2 (N3011, N3005, N505);
not NOT1 (N3012, N3008);
and AND3 (N3013, N3010, N1308, N2359);
not NOT1 (N3014, N3004);
xor XOR2 (N3015, N2995, N2891);
and AND3 (N3016, N3012, N1955, N3011);
nor NOR2 (N3017, N2551, N1343);
nor NOR3 (N3018, N3017, N601, N1760);
and AND4 (N3019, N3018, N253, N62, N962);
or OR4 (N3020, N3014, N479, N945, N1454);
and AND3 (N3021, N3003, N1576, N1309);
xor XOR2 (N3022, N3009, N628);
not NOT1 (N3023, N2980);
and AND4 (N3024, N3020, N1143, N300, N2852);
nor NOR2 (N3025, N3016, N2101);
or OR3 (N3026, N3015, N1445, N372);
or OR3 (N3027, N3013, N530, N1315);
not NOT1 (N3028, N3022);
xor XOR2 (N3029, N3007, N2003);
buf BUF1 (N3030, N3025);
nand NAND2 (N3031, N3030, N593);
not NOT1 (N3032, N3021);
nand NAND4 (N3033, N3026, N2067, N2872, N267);
or OR2 (N3034, N3031, N1463);
or OR4 (N3035, N3024, N1801, N1437, N286);
nor NOR4 (N3036, N3023, N139, N1722, N2678);
nor NOR3 (N3037, N3027, N425, N76);
buf BUF1 (N3038, N3035);
nor NOR2 (N3039, N3034, N327);
nor NOR2 (N3040, N3039, N439);
buf BUF1 (N3041, N3038);
and AND4 (N3042, N3036, N140, N2875, N2709);
nor NOR3 (N3043, N3032, N1936, N1158);
nor NOR2 (N3044, N3019, N2097);
not NOT1 (N3045, N3006);
nand NAND3 (N3046, N3029, N1454, N2518);
buf BUF1 (N3047, N3033);
nor NOR4 (N3048, N3043, N2975, N362, N1784);
not NOT1 (N3049, N3037);
xor XOR2 (N3050, N3048, N887);
nor NOR4 (N3051, N3042, N1942, N2731, N652);
nand NAND2 (N3052, N3046, N302);
xor XOR2 (N3053, N3049, N969);
not NOT1 (N3054, N3050);
xor XOR2 (N3055, N3045, N2332);
nand NAND4 (N3056, N3054, N1751, N262, N1244);
or OR4 (N3057, N3052, N2597, N2849, N1605);
nor NOR4 (N3058, N3047, N1729, N2620, N2708);
not NOT1 (N3059, N3051);
and AND4 (N3060, N3044, N2345, N779, N2530);
not NOT1 (N3061, N3041);
xor XOR2 (N3062, N3056, N2553);
buf BUF1 (N3063, N3053);
nor NOR4 (N3064, N3028, N462, N2979, N169);
not NOT1 (N3065, N3062);
xor XOR2 (N3066, N3059, N1368);
not NOT1 (N3067, N3065);
or OR3 (N3068, N3040, N2613, N878);
buf BUF1 (N3069, N3057);
nand NAND3 (N3070, N3067, N1320, N910);
buf BUF1 (N3071, N3063);
xor XOR2 (N3072, N3070, N394);
nor NOR3 (N3073, N3055, N913, N1043);
not NOT1 (N3074, N3061);
nand NAND2 (N3075, N3071, N1346);
nand NAND3 (N3076, N3064, N1757, N1463);
not NOT1 (N3077, N3058);
xor XOR2 (N3078, N3060, N787);
nor NOR3 (N3079, N3078, N1539, N1130);
xor XOR2 (N3080, N3066, N3016);
or OR3 (N3081, N3072, N367, N770);
buf BUF1 (N3082, N3076);
buf BUF1 (N3083, N3068);
xor XOR2 (N3084, N3083, N687);
buf BUF1 (N3085, N3079);
xor XOR2 (N3086, N3082, N1444);
xor XOR2 (N3087, N3073, N625);
nand NAND2 (N3088, N3086, N1016);
buf BUF1 (N3089, N3075);
and AND2 (N3090, N3077, N3006);
not NOT1 (N3091, N3089);
nor NOR4 (N3092, N3080, N413, N1084, N341);
xor XOR2 (N3093, N3081, N2018);
nand NAND2 (N3094, N3084, N759);
xor XOR2 (N3095, N3074, N1752);
nor NOR2 (N3096, N3088, N1478);
buf BUF1 (N3097, N3096);
not NOT1 (N3098, N3097);
and AND4 (N3099, N3095, N702, N2632, N1556);
and AND2 (N3100, N3099, N1963);
nor NOR2 (N3101, N3098, N332);
buf BUF1 (N3102, N3069);
xor XOR2 (N3103, N3085, N393);
and AND3 (N3104, N3103, N2108, N1386);
or OR2 (N3105, N3087, N1520);
nor NOR3 (N3106, N3102, N1674, N2311);
nand NAND4 (N3107, N3104, N2083, N1134, N1983);
or OR2 (N3108, N3101, N1341);
and AND3 (N3109, N3092, N2060, N739);
xor XOR2 (N3110, N3091, N1850);
not NOT1 (N3111, N3106);
xor XOR2 (N3112, N3100, N1511);
and AND3 (N3113, N3109, N461, N76);
nor NOR3 (N3114, N3094, N1522, N888);
nand NAND3 (N3115, N3110, N1225, N2115);
xor XOR2 (N3116, N3111, N2058);
and AND4 (N3117, N3115, N89, N1274, N2349);
and AND2 (N3118, N3112, N151);
not NOT1 (N3119, N3105);
and AND4 (N3120, N3107, N2074, N815, N296);
not NOT1 (N3121, N3118);
and AND4 (N3122, N3121, N2293, N642, N1169);
nor NOR2 (N3123, N3117, N1680);
nor NOR2 (N3124, N3113, N2101);
nand NAND4 (N3125, N3119, N2894, N2787, N1673);
buf BUF1 (N3126, N3125);
and AND3 (N3127, N3120, N1409, N1767);
and AND3 (N3128, N3090, N3040, N2959);
xor XOR2 (N3129, N3122, N1614);
not NOT1 (N3130, N3123);
nor NOR2 (N3131, N3129, N2374);
or OR4 (N3132, N3114, N1499, N434, N1037);
buf BUF1 (N3133, N3116);
nand NAND2 (N3134, N3126, N1929);
and AND4 (N3135, N3128, N1643, N1079, N2594);
not NOT1 (N3136, N3135);
or OR2 (N3137, N3132, N777);
or OR3 (N3138, N3136, N1849, N2185);
and AND3 (N3139, N3130, N2479, N1938);
or OR3 (N3140, N3138, N2694, N3115);
nand NAND2 (N3141, N3131, N2161);
nor NOR2 (N3142, N3133, N1706);
nand NAND2 (N3143, N3093, N888);
and AND3 (N3144, N3108, N1307, N1292);
not NOT1 (N3145, N3142);
nand NAND4 (N3146, N3144, N2574, N575, N1685);
buf BUF1 (N3147, N3127);
xor XOR2 (N3148, N3146, N1372);
nand NAND4 (N3149, N3137, N2610, N2825, N84);
nand NAND4 (N3150, N3140, N1323, N2996, N810);
and AND2 (N3151, N3145, N2694);
nand NAND3 (N3152, N3150, N2402, N412);
and AND2 (N3153, N3139, N2977);
not NOT1 (N3154, N3148);
buf BUF1 (N3155, N3141);
nand NAND2 (N3156, N3147, N2863);
nand NAND4 (N3157, N3149, N1538, N633, N2146);
nand NAND2 (N3158, N3157, N2021);
xor XOR2 (N3159, N3158, N3087);
not NOT1 (N3160, N3156);
nand NAND4 (N3161, N3153, N1513, N2597, N922);
buf BUF1 (N3162, N3161);
or OR3 (N3163, N3151, N1575, N360);
xor XOR2 (N3164, N3163, N1695);
not NOT1 (N3165, N3154);
not NOT1 (N3166, N3159);
or OR3 (N3167, N3143, N137, N501);
nor NOR2 (N3168, N3166, N1273);
and AND3 (N3169, N3164, N1155, N2556);
xor XOR2 (N3170, N3165, N1338);
not NOT1 (N3171, N3160);
and AND3 (N3172, N3170, N2070, N2723);
and AND2 (N3173, N3167, N520);
nor NOR2 (N3174, N3169, N1834);
xor XOR2 (N3175, N3172, N2410);
nand NAND4 (N3176, N3152, N2487, N2814, N2970);
and AND4 (N3177, N3176, N223, N2718, N919);
nand NAND4 (N3178, N3134, N2818, N390, N1373);
buf BUF1 (N3179, N3155);
xor XOR2 (N3180, N3179, N2393);
xor XOR2 (N3181, N3177, N1409);
buf BUF1 (N3182, N3175);
xor XOR2 (N3183, N3171, N269);
and AND3 (N3184, N3162, N1249, N1265);
or OR3 (N3185, N3178, N1668, N850);
not NOT1 (N3186, N3174);
nand NAND3 (N3187, N3185, N3085, N1299);
not NOT1 (N3188, N3124);
xor XOR2 (N3189, N3181, N4);
and AND4 (N3190, N3189, N2973, N535, N112);
xor XOR2 (N3191, N3186, N2696);
nor NOR4 (N3192, N3168, N812, N3173, N2661);
xor XOR2 (N3193, N238, N537);
xor XOR2 (N3194, N3182, N1076);
not NOT1 (N3195, N3183);
or OR4 (N3196, N3192, N2456, N2909, N1901);
nand NAND2 (N3197, N3191, N1407);
and AND4 (N3198, N3197, N321, N3140, N3119);
nor NOR4 (N3199, N3180, N1015, N1228, N1759);
and AND2 (N3200, N3199, N1841);
nand NAND4 (N3201, N3198, N441, N1765, N2251);
buf BUF1 (N3202, N3187);
or OR2 (N3203, N3193, N59);
and AND4 (N3204, N3202, N1597, N1797, N2842);
and AND3 (N3205, N3196, N2769, N3149);
or OR4 (N3206, N3200, N72, N2816, N1500);
and AND2 (N3207, N3195, N836);
nand NAND4 (N3208, N3206, N1952, N1035, N2677);
xor XOR2 (N3209, N3208, N617);
not NOT1 (N3210, N3194);
or OR4 (N3211, N3201, N2548, N968, N1244);
or OR2 (N3212, N3184, N574);
nand NAND2 (N3213, N3203, N284);
nor NOR2 (N3214, N3211, N2554);
buf BUF1 (N3215, N3213);
nor NOR4 (N3216, N3207, N2537, N492, N1914);
and AND2 (N3217, N3216, N1744);
xor XOR2 (N3218, N3204, N1330);
buf BUF1 (N3219, N3205);
nand NAND3 (N3220, N3188, N2243, N3072);
buf BUF1 (N3221, N3219);
nor NOR3 (N3222, N3210, N1018, N2191);
or OR3 (N3223, N3215, N2783, N2138);
or OR2 (N3224, N3218, N405);
nor NOR2 (N3225, N3217, N970);
xor XOR2 (N3226, N3212, N145);
nand NAND2 (N3227, N3226, N2180);
xor XOR2 (N3228, N3209, N3160);
buf BUF1 (N3229, N3228);
and AND2 (N3230, N3214, N1299);
buf BUF1 (N3231, N3220);
and AND4 (N3232, N3231, N1819, N265, N1571);
buf BUF1 (N3233, N3227);
or OR4 (N3234, N3190, N2148, N1736, N1085);
or OR3 (N3235, N3233, N726, N925);
not NOT1 (N3236, N3225);
xor XOR2 (N3237, N3224, N573);
nand NAND4 (N3238, N3223, N355, N15, N533);
nor NOR4 (N3239, N3237, N28, N879, N225);
buf BUF1 (N3240, N3230);
xor XOR2 (N3241, N3232, N1565);
or OR3 (N3242, N3222, N16, N2260);
buf BUF1 (N3243, N3240);
nand NAND2 (N3244, N3221, N394);
nor NOR2 (N3245, N3238, N884);
xor XOR2 (N3246, N3245, N2552);
not NOT1 (N3247, N3234);
buf BUF1 (N3248, N3229);
buf BUF1 (N3249, N3235);
not NOT1 (N3250, N3249);
nand NAND3 (N3251, N3248, N2075, N2084);
buf BUF1 (N3252, N3239);
nand NAND3 (N3253, N3247, N609, N1549);
not NOT1 (N3254, N3244);
or OR3 (N3255, N3243, N1893, N91);
or OR3 (N3256, N3251, N2250, N990);
nand NAND2 (N3257, N3236, N2660);
and AND2 (N3258, N3255, N1831);
or OR3 (N3259, N3242, N1287, N246);
or OR2 (N3260, N3250, N1600);
xor XOR2 (N3261, N3254, N2069);
or OR3 (N3262, N3241, N1617, N392);
xor XOR2 (N3263, N3256, N1035);
not NOT1 (N3264, N3262);
nor NOR4 (N3265, N3253, N2016, N3074, N653);
buf BUF1 (N3266, N3258);
not NOT1 (N3267, N3266);
nor NOR4 (N3268, N3265, N1536, N1834, N3148);
not NOT1 (N3269, N3260);
nor NOR2 (N3270, N3269, N2670);
buf BUF1 (N3271, N3261);
nor NOR2 (N3272, N3259, N2366);
not NOT1 (N3273, N3252);
not NOT1 (N3274, N3271);
nand NAND2 (N3275, N3264, N752);
or OR3 (N3276, N3267, N656, N895);
not NOT1 (N3277, N3273);
nor NOR4 (N3278, N3272, N307, N1262, N2826);
or OR4 (N3279, N3268, N2258, N2306, N2959);
nand NAND3 (N3280, N3270, N2244, N1757);
nand NAND3 (N3281, N3246, N1777, N3006);
nor NOR2 (N3282, N3280, N2626);
xor XOR2 (N3283, N3276, N2326);
and AND3 (N3284, N3281, N1722, N121);
nor NOR2 (N3285, N3275, N2196);
nand NAND4 (N3286, N3279, N27, N124, N387);
nand NAND3 (N3287, N3257, N982, N1186);
nor NOR2 (N3288, N3286, N12);
nand NAND4 (N3289, N3285, N20, N2493, N300);
or OR2 (N3290, N3289, N224);
xor XOR2 (N3291, N3277, N1805);
buf BUF1 (N3292, N3291);
nor NOR3 (N3293, N3292, N1029, N930);
buf BUF1 (N3294, N3263);
nand NAND3 (N3295, N3274, N2291, N299);
not NOT1 (N3296, N3282);
buf BUF1 (N3297, N3283);
not NOT1 (N3298, N3290);
nor NOR3 (N3299, N3298, N1307, N1719);
nand NAND4 (N3300, N3294, N348, N215, N2314);
and AND2 (N3301, N3284, N3061);
nand NAND2 (N3302, N3278, N2396);
not NOT1 (N3303, N3287);
nand NAND3 (N3304, N3299, N2808, N255);
and AND4 (N3305, N3303, N3162, N677, N1902);
or OR2 (N3306, N3295, N2309);
not NOT1 (N3307, N3304);
or OR2 (N3308, N3306, N347);
not NOT1 (N3309, N3307);
xor XOR2 (N3310, N3300, N3182);
xor XOR2 (N3311, N3309, N1081);
not NOT1 (N3312, N3302);
or OR3 (N3313, N3308, N922, N2461);
nor NOR3 (N3314, N3305, N2440, N25);
xor XOR2 (N3315, N3311, N1517);
nor NOR4 (N3316, N3310, N1138, N2234, N129);
nor NOR3 (N3317, N3293, N2286, N3053);
nor NOR4 (N3318, N3301, N2720, N2545, N3152);
xor XOR2 (N3319, N3317, N602);
buf BUF1 (N3320, N3296);
xor XOR2 (N3321, N3288, N2624);
nand NAND2 (N3322, N3319, N1161);
nor NOR4 (N3323, N3315, N1262, N784, N2953);
and AND3 (N3324, N3320, N1030, N3124);
buf BUF1 (N3325, N3321);
and AND3 (N3326, N3318, N1831, N616);
and AND3 (N3327, N3323, N111, N818);
nor NOR2 (N3328, N3322, N82);
xor XOR2 (N3329, N3327, N857);
and AND4 (N3330, N3325, N620, N428, N2127);
buf BUF1 (N3331, N3297);
or OR2 (N3332, N3326, N2606);
nand NAND4 (N3333, N3316, N3137, N2548, N896);
not NOT1 (N3334, N3313);
xor XOR2 (N3335, N3330, N307);
nor NOR4 (N3336, N3332, N1002, N533, N1130);
nand NAND3 (N3337, N3331, N2021, N1640);
xor XOR2 (N3338, N3337, N2132);
nand NAND3 (N3339, N3333, N2084, N121);
xor XOR2 (N3340, N3329, N3250);
not NOT1 (N3341, N3312);
buf BUF1 (N3342, N3328);
buf BUF1 (N3343, N3341);
or OR4 (N3344, N3334, N444, N1196, N1031);
xor XOR2 (N3345, N3338, N2145);
and AND2 (N3346, N3324, N1613);
xor XOR2 (N3347, N3342, N1931);
nor NOR4 (N3348, N3340, N1715, N1801, N1318);
and AND4 (N3349, N3346, N1047, N981, N3239);
not NOT1 (N3350, N3345);
or OR4 (N3351, N3339, N81, N2279, N3073);
xor XOR2 (N3352, N3343, N1613);
nand NAND3 (N3353, N3349, N2529, N3334);
xor XOR2 (N3354, N3335, N2658);
nor NOR4 (N3355, N3352, N924, N735, N2260);
nand NAND3 (N3356, N3336, N318, N1576);
xor XOR2 (N3357, N3347, N550);
not NOT1 (N3358, N3354);
xor XOR2 (N3359, N3356, N1620);
not NOT1 (N3360, N3314);
not NOT1 (N3361, N3353);
nand NAND3 (N3362, N3351, N3356, N1949);
xor XOR2 (N3363, N3361, N2945);
buf BUF1 (N3364, N3357);
not NOT1 (N3365, N3344);
xor XOR2 (N3366, N3364, N411);
nor NOR2 (N3367, N3358, N1915);
or OR4 (N3368, N3348, N578, N1188, N3130);
nand NAND3 (N3369, N3367, N3325, N3299);
nor NOR3 (N3370, N3359, N2576, N1428);
nor NOR3 (N3371, N3362, N422, N2062);
buf BUF1 (N3372, N3368);
not NOT1 (N3373, N3363);
buf BUF1 (N3374, N3373);
nand NAND3 (N3375, N3371, N1816, N1261);
nand NAND2 (N3376, N3365, N2719);
xor XOR2 (N3377, N3360, N331);
nor NOR2 (N3378, N3375, N424);
nand NAND2 (N3379, N3378, N1661);
not NOT1 (N3380, N3374);
nor NOR4 (N3381, N3376, N3117, N1815, N1801);
and AND3 (N3382, N3372, N1965, N2796);
nand NAND3 (N3383, N3380, N2983, N920);
and AND2 (N3384, N3370, N345);
and AND3 (N3385, N3366, N2999, N272);
nand NAND2 (N3386, N3382, N2272);
buf BUF1 (N3387, N3386);
or OR3 (N3388, N3355, N1769, N792);
or OR3 (N3389, N3388, N2823, N1947);
or OR2 (N3390, N3369, N578);
and AND3 (N3391, N3387, N3363, N2716);
buf BUF1 (N3392, N3377);
nand NAND2 (N3393, N3384, N669);
and AND4 (N3394, N3390, N1261, N2693, N1969);
or OR3 (N3395, N3391, N3251, N113);
nand NAND4 (N3396, N3389, N1975, N1714, N1014);
and AND2 (N3397, N3381, N3130);
not NOT1 (N3398, N3396);
nand NAND2 (N3399, N3392, N1328);
xor XOR2 (N3400, N3397, N1904);
buf BUF1 (N3401, N3393);
nor NOR3 (N3402, N3395, N415, N1812);
and AND4 (N3403, N3402, N1083, N2438, N2101);
xor XOR2 (N3404, N3383, N2369);
xor XOR2 (N3405, N3401, N2954);
not NOT1 (N3406, N3405);
and AND2 (N3407, N3406, N2707);
nand NAND2 (N3408, N3403, N2745);
nor NOR4 (N3409, N3379, N2475, N805, N915);
nor NOR2 (N3410, N3409, N481);
xor XOR2 (N3411, N3350, N186);
not NOT1 (N3412, N3398);
or OR2 (N3413, N3394, N3026);
nand NAND3 (N3414, N3407, N80, N3102);
buf BUF1 (N3415, N3413);
xor XOR2 (N3416, N3385, N2949);
or OR3 (N3417, N3415, N658, N2550);
and AND3 (N3418, N3404, N2848, N2316);
nor NOR2 (N3419, N3411, N298);
not NOT1 (N3420, N3412);
xor XOR2 (N3421, N3414, N1029);
and AND4 (N3422, N3399, N985, N3099, N3111);
not NOT1 (N3423, N3422);
or OR3 (N3424, N3421, N2191, N2586);
or OR2 (N3425, N3400, N1605);
nand NAND4 (N3426, N3417, N2640, N1592, N1506);
or OR3 (N3427, N3418, N3303, N722);
nor NOR4 (N3428, N3416, N1813, N1661, N2705);
or OR3 (N3429, N3419, N1061, N2490);
and AND2 (N3430, N3420, N535);
nor NOR2 (N3431, N3426, N489);
nor NOR3 (N3432, N3425, N1449, N1621);
not NOT1 (N3433, N3430);
nor NOR4 (N3434, N3427, N1607, N2657, N1017);
buf BUF1 (N3435, N3410);
not NOT1 (N3436, N3435);
xor XOR2 (N3437, N3424, N593);
not NOT1 (N3438, N3434);
xor XOR2 (N3439, N3423, N2880);
nand NAND4 (N3440, N3436, N1747, N1942, N1255);
buf BUF1 (N3441, N3440);
nor NOR4 (N3442, N3437, N2532, N2658, N694);
or OR3 (N3443, N3441, N2214, N469);
nand NAND3 (N3444, N3443, N2165, N506);
buf BUF1 (N3445, N3432);
or OR4 (N3446, N3439, N2287, N1596, N1909);
nand NAND2 (N3447, N3438, N505);
nor NOR4 (N3448, N3429, N3100, N581, N3047);
xor XOR2 (N3449, N3448, N1719);
and AND4 (N3450, N3449, N138, N1304, N1495);
or OR2 (N3451, N3447, N3239);
nor NOR4 (N3452, N3442, N1933, N1501, N3161);
xor XOR2 (N3453, N3433, N1443);
nand NAND2 (N3454, N3452, N2573);
xor XOR2 (N3455, N3451, N1282);
or OR3 (N3456, N3446, N1286, N954);
nand NAND4 (N3457, N3428, N572, N797, N1046);
nand NAND2 (N3458, N3456, N3241);
or OR3 (N3459, N3453, N1842, N2100);
nand NAND2 (N3460, N3457, N1591);
or OR2 (N3461, N3408, N3257);
or OR4 (N3462, N3455, N1513, N403, N608);
and AND4 (N3463, N3458, N3082, N1406, N2304);
nand NAND4 (N3464, N3431, N3114, N1522, N3433);
and AND4 (N3465, N3462, N1198, N1773, N2201);
and AND4 (N3466, N3445, N2212, N9, N127);
or OR3 (N3467, N3465, N2432, N1020);
and AND3 (N3468, N3450, N941, N3380);
buf BUF1 (N3469, N3460);
or OR4 (N3470, N3464, N3319, N2083, N239);
and AND2 (N3471, N3466, N3059);
nand NAND3 (N3472, N3470, N2035, N847);
nor NOR4 (N3473, N3459, N2049, N1721, N634);
xor XOR2 (N3474, N3467, N221);
or OR2 (N3475, N3472, N630);
and AND3 (N3476, N3468, N267, N1209);
nand NAND4 (N3477, N3473, N452, N2324, N364);
not NOT1 (N3478, N3463);
or OR4 (N3479, N3469, N9, N3400, N1542);
and AND2 (N3480, N3477, N3062);
not NOT1 (N3481, N3454);
and AND2 (N3482, N3476, N2622);
and AND4 (N3483, N3478, N76, N2507, N1321);
buf BUF1 (N3484, N3471);
or OR2 (N3485, N3474, N2107);
nor NOR2 (N3486, N3479, N2655);
not NOT1 (N3487, N3481);
nor NOR4 (N3488, N3480, N1064, N722, N1292);
or OR2 (N3489, N3487, N2169);
and AND2 (N3490, N3488, N2786);
nor NOR2 (N3491, N3482, N2633);
nor NOR3 (N3492, N3490, N1294, N3466);
or OR4 (N3493, N3489, N3004, N1155, N209);
and AND4 (N3494, N3491, N994, N2855, N433);
nor NOR3 (N3495, N3484, N779, N107);
nor NOR4 (N3496, N3475, N2550, N1516, N818);
nand NAND4 (N3497, N3494, N1989, N1199, N3157);
not NOT1 (N3498, N3486);
not NOT1 (N3499, N3497);
not NOT1 (N3500, N3498);
nand NAND4 (N3501, N3444, N180, N147, N1520);
nor NOR4 (N3502, N3499, N725, N543, N1896);
buf BUF1 (N3503, N3485);
nand NAND2 (N3504, N3502, N2290);
and AND4 (N3505, N3461, N791, N3168, N953);
or OR3 (N3506, N3501, N298, N2882);
or OR4 (N3507, N3492, N3474, N3503, N2297);
nand NAND3 (N3508, N3395, N3102, N1991);
nor NOR3 (N3509, N3508, N2415, N1678);
not NOT1 (N3510, N3493);
buf BUF1 (N3511, N3507);
or OR2 (N3512, N3500, N488);
and AND2 (N3513, N3504, N2224);
xor XOR2 (N3514, N3509, N1349);
and AND4 (N3515, N3511, N2299, N1200, N1294);
or OR4 (N3516, N3515, N2109, N207, N1199);
or OR3 (N3517, N3505, N2530, N3422);
xor XOR2 (N3518, N3514, N750);
buf BUF1 (N3519, N3517);
nand NAND3 (N3520, N3513, N1507, N2832);
or OR4 (N3521, N3512, N2522, N3370, N1672);
xor XOR2 (N3522, N3506, N141);
buf BUF1 (N3523, N3495);
xor XOR2 (N3524, N3483, N3045);
nor NOR4 (N3525, N3518, N176, N1008, N128);
buf BUF1 (N3526, N3516);
buf BUF1 (N3527, N3526);
and AND4 (N3528, N3527, N982, N1688, N1243);
xor XOR2 (N3529, N3524, N227);
xor XOR2 (N3530, N3496, N1316);
xor XOR2 (N3531, N3523, N2213);
nor NOR3 (N3532, N3529, N3453, N3296);
xor XOR2 (N3533, N3520, N2722);
xor XOR2 (N3534, N3531, N1907);
nor NOR2 (N3535, N3522, N2778);
or OR3 (N3536, N3528, N2914, N256);
not NOT1 (N3537, N3510);
or OR4 (N3538, N3519, N2480, N593, N3107);
and AND4 (N3539, N3537, N2833, N1124, N2130);
buf BUF1 (N3540, N3530);
not NOT1 (N3541, N3533);
nor NOR4 (N3542, N3532, N1773, N2950, N1352);
and AND2 (N3543, N3541, N2496);
xor XOR2 (N3544, N3543, N42);
nand NAND4 (N3545, N3539, N1836, N1780, N3539);
and AND4 (N3546, N3540, N3196, N1479, N2407);
nor NOR2 (N3547, N3536, N3417);
or OR3 (N3548, N3546, N1066, N1238);
buf BUF1 (N3549, N3545);
nand NAND3 (N3550, N3544, N900, N3289);
not NOT1 (N3551, N3521);
buf BUF1 (N3552, N3551);
not NOT1 (N3553, N3550);
nor NOR2 (N3554, N3525, N3457);
or OR3 (N3555, N3538, N252, N3448);
nand NAND2 (N3556, N3552, N1971);
not NOT1 (N3557, N3542);
and AND3 (N3558, N3549, N1156, N2458);
or OR4 (N3559, N3555, N2477, N3161, N1249);
xor XOR2 (N3560, N3534, N663);
or OR3 (N3561, N3548, N176, N1405);
nand NAND4 (N3562, N3558, N2548, N132, N1540);
and AND3 (N3563, N3535, N627, N1146);
xor XOR2 (N3564, N3553, N2243);
xor XOR2 (N3565, N3560, N1756);
and AND4 (N3566, N3563, N3172, N2913, N1275);
nor NOR2 (N3567, N3557, N1608);
not NOT1 (N3568, N3567);
nand NAND3 (N3569, N3562, N3116, N2837);
not NOT1 (N3570, N3564);
and AND3 (N3571, N3570, N1269, N1060);
and AND3 (N3572, N3559, N2389, N1683);
not NOT1 (N3573, N3547);
not NOT1 (N3574, N3566);
nor NOR2 (N3575, N3569, N404);
and AND2 (N3576, N3573, N1158);
or OR2 (N3577, N3576, N1189);
and AND3 (N3578, N3571, N3049, N1294);
xor XOR2 (N3579, N3556, N2511);
buf BUF1 (N3580, N3568);
nor NOR2 (N3581, N3565, N1587);
nand NAND4 (N3582, N3572, N1202, N3160, N2548);
nor NOR3 (N3583, N3579, N2458, N1577);
xor XOR2 (N3584, N3554, N2088);
buf BUF1 (N3585, N3582);
nand NAND2 (N3586, N3583, N222);
and AND2 (N3587, N3580, N896);
not NOT1 (N3588, N3578);
nand NAND4 (N3589, N3586, N1403, N1946, N1954);
or OR3 (N3590, N3575, N585, N646);
xor XOR2 (N3591, N3584, N2899);
or OR3 (N3592, N3589, N2807, N816);
nor NOR3 (N3593, N3587, N2688, N1084);
nand NAND3 (N3594, N3561, N654, N2592);
or OR4 (N3595, N3594, N2768, N2885, N2532);
nor NOR2 (N3596, N3593, N2207);
or OR3 (N3597, N3585, N2532, N724);
or OR3 (N3598, N3581, N491, N2030);
xor XOR2 (N3599, N3590, N2481);
nor NOR2 (N3600, N3597, N927);
buf BUF1 (N3601, N3588);
not NOT1 (N3602, N3601);
nor NOR3 (N3603, N3577, N1016, N2222);
and AND2 (N3604, N3602, N1408);
nand NAND2 (N3605, N3603, N2944);
buf BUF1 (N3606, N3574);
and AND3 (N3607, N3598, N3554, N2650);
nand NAND4 (N3608, N3592, N3580, N2048, N2483);
or OR3 (N3609, N3608, N1567, N2332);
or OR2 (N3610, N3604, N3109);
buf BUF1 (N3611, N3596);
and AND3 (N3612, N3606, N3048, N1556);
xor XOR2 (N3613, N3599, N1367);
or OR2 (N3614, N3591, N3198);
buf BUF1 (N3615, N3613);
buf BUF1 (N3616, N3612);
and AND3 (N3617, N3605, N2378, N1575);
buf BUF1 (N3618, N3607);
nand NAND2 (N3619, N3615, N2563);
nor NOR2 (N3620, N3618, N536);
buf BUF1 (N3621, N3616);
and AND3 (N3622, N3617, N2506, N1019);
and AND3 (N3623, N3611, N2883, N286);
buf BUF1 (N3624, N3622);
buf BUF1 (N3625, N3610);
buf BUF1 (N3626, N3595);
and AND3 (N3627, N3624, N536, N1057);
not NOT1 (N3628, N3600);
and AND4 (N3629, N3620, N1825, N379, N2870);
nand NAND2 (N3630, N3614, N3057);
nand NAND2 (N3631, N3623, N1747);
buf BUF1 (N3632, N3630);
nand NAND2 (N3633, N3627, N870);
and AND4 (N3634, N3629, N3104, N3240, N3062);
not NOT1 (N3635, N3632);
and AND4 (N3636, N3633, N3303, N1048, N1538);
or OR3 (N3637, N3609, N3235, N2945);
xor XOR2 (N3638, N3635, N3382);
not NOT1 (N3639, N3634);
not NOT1 (N3640, N3636);
nor NOR4 (N3641, N3637, N1971, N1446, N2964);
not NOT1 (N3642, N3639);
and AND2 (N3643, N3642, N71);
buf BUF1 (N3644, N3628);
xor XOR2 (N3645, N3641, N3049);
and AND3 (N3646, N3625, N2379, N181);
not NOT1 (N3647, N3646);
not NOT1 (N3648, N3619);
nor NOR2 (N3649, N3640, N2905);
buf BUF1 (N3650, N3643);
not NOT1 (N3651, N3647);
xor XOR2 (N3652, N3638, N3388);
nor NOR2 (N3653, N3650, N1144);
or OR2 (N3654, N3651, N1311);
or OR3 (N3655, N3652, N2805, N1848);
nand NAND4 (N3656, N3654, N666, N2356, N3602);
nand NAND4 (N3657, N3621, N2255, N1328, N2385);
xor XOR2 (N3658, N3656, N1394);
nor NOR3 (N3659, N3626, N2472, N1294);
not NOT1 (N3660, N3657);
nor NOR3 (N3661, N3631, N3357, N1708);
nor NOR3 (N3662, N3649, N1211, N2571);
xor XOR2 (N3663, N3661, N2007);
or OR2 (N3664, N3663, N625);
nor NOR3 (N3665, N3645, N724, N3533);
not NOT1 (N3666, N3659);
nor NOR4 (N3667, N3655, N1286, N862, N3273);
xor XOR2 (N3668, N3653, N2746);
xor XOR2 (N3669, N3644, N1024);
nand NAND4 (N3670, N3668, N40, N1074, N96);
nand NAND3 (N3671, N3665, N1015, N1667);
or OR3 (N3672, N3662, N1200, N1643);
not NOT1 (N3673, N3658);
nand NAND3 (N3674, N3671, N3260, N619);
xor XOR2 (N3675, N3660, N3459);
nand NAND2 (N3676, N3670, N3572);
nand NAND2 (N3677, N3669, N886);
not NOT1 (N3678, N3667);
nor NOR4 (N3679, N3666, N638, N3388, N3502);
and AND2 (N3680, N3648, N3301);
and AND2 (N3681, N3678, N1883);
xor XOR2 (N3682, N3674, N2181);
or OR2 (N3683, N3680, N1109);
and AND3 (N3684, N3676, N3431, N3427);
or OR4 (N3685, N3683, N2556, N2026, N962);
not NOT1 (N3686, N3682);
or OR3 (N3687, N3672, N388, N3498);
xor XOR2 (N3688, N3681, N171);
not NOT1 (N3689, N3685);
or OR3 (N3690, N3675, N2766, N54);
and AND4 (N3691, N3684, N2663, N1623, N2373);
and AND2 (N3692, N3691, N1943);
nand NAND3 (N3693, N3689, N2679, N2889);
buf BUF1 (N3694, N3677);
buf BUF1 (N3695, N3694);
xor XOR2 (N3696, N3687, N863);
and AND4 (N3697, N3664, N3520, N3536, N2744);
xor XOR2 (N3698, N3697, N1930);
xor XOR2 (N3699, N3688, N1044);
nand NAND3 (N3700, N3698, N616, N1270);
or OR2 (N3701, N3679, N3662);
nor NOR2 (N3702, N3673, N2170);
and AND2 (N3703, N3692, N375);
and AND3 (N3704, N3695, N3413, N1261);
and AND3 (N3705, N3696, N2828, N3559);
and AND3 (N3706, N3693, N2245, N2400);
buf BUF1 (N3707, N3701);
buf BUF1 (N3708, N3704);
xor XOR2 (N3709, N3705, N94);
and AND4 (N3710, N3708, N3183, N2177, N408);
or OR3 (N3711, N3686, N3475, N1962);
and AND3 (N3712, N3707, N87, N680);
or OR4 (N3713, N3702, N3244, N3675, N3447);
buf BUF1 (N3714, N3699);
not NOT1 (N3715, N3706);
buf BUF1 (N3716, N3713);
and AND2 (N3717, N3710, N3032);
nor NOR4 (N3718, N3716, N3334, N1101, N3653);
not NOT1 (N3719, N3715);
buf BUF1 (N3720, N3703);
nand NAND2 (N3721, N3690, N3007);
nor NOR2 (N3722, N3719, N455);
and AND2 (N3723, N3718, N187);
buf BUF1 (N3724, N3722);
buf BUF1 (N3725, N3724);
not NOT1 (N3726, N3714);
xor XOR2 (N3727, N3700, N3055);
not NOT1 (N3728, N3727);
xor XOR2 (N3729, N3721, N527);
buf BUF1 (N3730, N3717);
nand NAND2 (N3731, N3728, N352);
nor NOR2 (N3732, N3711, N1195);
and AND3 (N3733, N3729, N3663, N637);
xor XOR2 (N3734, N3709, N1363);
xor XOR2 (N3735, N3731, N934);
nand NAND2 (N3736, N3735, N2676);
and AND4 (N3737, N3736, N1462, N3191, N3721);
xor XOR2 (N3738, N3733, N1355);
not NOT1 (N3739, N3738);
or OR3 (N3740, N3739, N3072, N1389);
nor NOR2 (N3741, N3726, N3090);
and AND3 (N3742, N3737, N870, N211);
buf BUF1 (N3743, N3712);
buf BUF1 (N3744, N3740);
xor XOR2 (N3745, N3743, N22);
or OR2 (N3746, N3744, N1947);
nor NOR3 (N3747, N3741, N3145, N2981);
xor XOR2 (N3748, N3742, N999);
xor XOR2 (N3749, N3723, N2604);
or OR3 (N3750, N3725, N713, N2744);
nor NOR2 (N3751, N3732, N189);
buf BUF1 (N3752, N3734);
buf BUF1 (N3753, N3750);
or OR3 (N3754, N3746, N2483, N109);
not NOT1 (N3755, N3748);
or OR2 (N3756, N3753, N3443);
buf BUF1 (N3757, N3730);
nor NOR2 (N3758, N3749, N3042);
or OR2 (N3759, N3755, N3083);
not NOT1 (N3760, N3720);
buf BUF1 (N3761, N3760);
not NOT1 (N3762, N3754);
nand NAND2 (N3763, N3758, N1894);
not NOT1 (N3764, N3763);
and AND3 (N3765, N3762, N1859, N1511);
and AND3 (N3766, N3751, N38, N3571);
or OR3 (N3767, N3752, N3423, N362);
xor XOR2 (N3768, N3757, N1999);
not NOT1 (N3769, N3761);
buf BUF1 (N3770, N3767);
nand NAND4 (N3771, N3756, N1485, N3346, N2330);
nand NAND2 (N3772, N3765, N1429);
xor XOR2 (N3773, N3759, N1265);
or OR3 (N3774, N3766, N1377, N3016);
nand NAND2 (N3775, N3771, N802);
buf BUF1 (N3776, N3764);
nand NAND2 (N3777, N3768, N3426);
nand NAND2 (N3778, N3769, N3146);
buf BUF1 (N3779, N3778);
or OR2 (N3780, N3745, N2499);
nand NAND2 (N3781, N3777, N551);
nor NOR2 (N3782, N3773, N1468);
nand NAND4 (N3783, N3770, N3633, N2321, N947);
nor NOR3 (N3784, N3779, N314, N2015);
not NOT1 (N3785, N3747);
or OR2 (N3786, N3775, N572);
xor XOR2 (N3787, N3784, N751);
nor NOR3 (N3788, N3774, N198, N3619);
and AND3 (N3789, N3783, N2908, N392);
or OR4 (N3790, N3789, N1199, N607, N2195);
or OR3 (N3791, N3772, N2205, N3704);
or OR3 (N3792, N3781, N1132, N2343);
and AND2 (N3793, N3782, N3108);
xor XOR2 (N3794, N3788, N2868);
or OR3 (N3795, N3785, N3439, N717);
xor XOR2 (N3796, N3791, N2411);
buf BUF1 (N3797, N3792);
xor XOR2 (N3798, N3797, N2180);
buf BUF1 (N3799, N3780);
or OR3 (N3800, N3796, N1872, N2388);
xor XOR2 (N3801, N3799, N497);
or OR2 (N3802, N3793, N2591);
nand NAND3 (N3803, N3787, N718, N1667);
not NOT1 (N3804, N3786);
nor NOR4 (N3805, N3801, N1872, N1583, N2440);
nand NAND4 (N3806, N3804, N2085, N132, N422);
nand NAND3 (N3807, N3795, N3694, N2458);
buf BUF1 (N3808, N3807);
nor NOR2 (N3809, N3802, N1058);
or OR4 (N3810, N3809, N3353, N659, N1655);
buf BUF1 (N3811, N3810);
and AND4 (N3812, N3794, N1427, N1234, N2494);
nand NAND4 (N3813, N3805, N1692, N3773, N832);
or OR2 (N3814, N3808, N754);
nor NOR2 (N3815, N3803, N2884);
buf BUF1 (N3816, N3790);
not NOT1 (N3817, N3816);
or OR3 (N3818, N3776, N2463, N3002);
xor XOR2 (N3819, N3818, N1206);
xor XOR2 (N3820, N3813, N13);
nor NOR3 (N3821, N3798, N1333, N1807);
and AND2 (N3822, N3815, N679);
or OR4 (N3823, N3800, N2692, N1123, N2627);
buf BUF1 (N3824, N3812);
buf BUF1 (N3825, N3811);
nor NOR2 (N3826, N3806, N3741);
or OR2 (N3827, N3826, N137);
and AND4 (N3828, N3824, N1787, N1460, N2390);
buf BUF1 (N3829, N3827);
and AND2 (N3830, N3814, N3066);
nand NAND2 (N3831, N3819, N1018);
nor NOR4 (N3832, N3823, N2838, N3318, N814);
and AND3 (N3833, N3829, N2077, N513);
not NOT1 (N3834, N3830);
xor XOR2 (N3835, N3822, N1846);
nor NOR4 (N3836, N3835, N3176, N3325, N3186);
xor XOR2 (N3837, N3833, N2545);
and AND2 (N3838, N3834, N276);
nor NOR3 (N3839, N3837, N613, N444);
or OR3 (N3840, N3820, N3674, N1721);
not NOT1 (N3841, N3817);
and AND3 (N3842, N3821, N211, N3030);
nand NAND2 (N3843, N3838, N2872);
and AND2 (N3844, N3832, N1074);
nor NOR3 (N3845, N3844, N1410, N628);
buf BUF1 (N3846, N3843);
or OR4 (N3847, N3845, N2982, N3140, N2159);
or OR4 (N3848, N3842, N16, N1821, N3806);
xor XOR2 (N3849, N3831, N1273);
nor NOR4 (N3850, N3847, N298, N3755, N2869);
nand NAND4 (N3851, N3850, N574, N3757, N263);
or OR2 (N3852, N3836, N1103);
and AND3 (N3853, N3851, N1327, N1923);
nor NOR3 (N3854, N3828, N717, N3405);
buf BUF1 (N3855, N3839);
nand NAND3 (N3856, N3855, N972, N1504);
or OR4 (N3857, N3846, N832, N715, N3531);
buf BUF1 (N3858, N3854);
or OR4 (N3859, N3852, N3455, N1674, N2346);
nand NAND3 (N3860, N3848, N593, N654);
xor XOR2 (N3861, N3857, N510);
not NOT1 (N3862, N3849);
buf BUF1 (N3863, N3841);
nor NOR3 (N3864, N3859, N3246, N1214);
nor NOR4 (N3865, N3863, N3021, N1346, N200);
and AND4 (N3866, N3860, N12, N1941, N1747);
and AND3 (N3867, N3861, N1444, N2104);
buf BUF1 (N3868, N3840);
or OR2 (N3869, N3825, N3454);
or OR4 (N3870, N3865, N1105, N1796, N3747);
nand NAND4 (N3871, N3856, N1112, N1159, N221);
nand NAND4 (N3872, N3868, N748, N1086, N23);
nor NOR3 (N3873, N3872, N2830, N227);
not NOT1 (N3874, N3873);
not NOT1 (N3875, N3870);
nor NOR3 (N3876, N3866, N2105, N2945);
not NOT1 (N3877, N3876);
and AND4 (N3878, N3867, N639, N3282, N1694);
not NOT1 (N3879, N3877);
xor XOR2 (N3880, N3878, N2276);
not NOT1 (N3881, N3853);
or OR3 (N3882, N3858, N2638, N3147);
or OR2 (N3883, N3874, N3492);
and AND4 (N3884, N3881, N3134, N3603, N2879);
and AND2 (N3885, N3862, N148);
nor NOR2 (N3886, N3882, N1671);
not NOT1 (N3887, N3884);
or OR3 (N3888, N3879, N2118, N679);
nor NOR4 (N3889, N3883, N3303, N380, N2228);
buf BUF1 (N3890, N3880);
not NOT1 (N3891, N3871);
or OR3 (N3892, N3890, N2802, N2201);
and AND3 (N3893, N3891, N2789, N1037);
buf BUF1 (N3894, N3869);
xor XOR2 (N3895, N3887, N1689);
xor XOR2 (N3896, N3889, N1608);
xor XOR2 (N3897, N3864, N3747);
buf BUF1 (N3898, N3875);
not NOT1 (N3899, N3893);
nand NAND3 (N3900, N3898, N845, N549);
xor XOR2 (N3901, N3886, N402);
xor XOR2 (N3902, N3888, N3193);
nand NAND2 (N3903, N3894, N155);
buf BUF1 (N3904, N3895);
nor NOR2 (N3905, N3902, N742);
or OR2 (N3906, N3885, N3079);
nand NAND2 (N3907, N3901, N3288);
or OR2 (N3908, N3899, N389);
or OR3 (N3909, N3908, N389, N1445);
buf BUF1 (N3910, N3906);
not NOT1 (N3911, N3909);
buf BUF1 (N3912, N3896);
not NOT1 (N3913, N3907);
and AND2 (N3914, N3905, N1916);
and AND4 (N3915, N3904, N2135, N289, N2577);
nand NAND2 (N3916, N3892, N2536);
and AND4 (N3917, N3913, N2648, N3240, N2990);
and AND4 (N3918, N3903, N2758, N1065, N3484);
not NOT1 (N3919, N3900);
or OR2 (N3920, N3897, N2164);
not NOT1 (N3921, N3911);
nand NAND2 (N3922, N3915, N1158);
and AND2 (N3923, N3912, N659);
not NOT1 (N3924, N3916);
or OR3 (N3925, N3920, N1109, N810);
nor NOR3 (N3926, N3923, N1902, N2552);
or OR3 (N3927, N3921, N745, N3063);
nand NAND4 (N3928, N3918, N1781, N2821, N1591);
not NOT1 (N3929, N3917);
buf BUF1 (N3930, N3919);
nor NOR3 (N3931, N3924, N811, N3747);
nand NAND3 (N3932, N3926, N1370, N560);
nor NOR3 (N3933, N3930, N144, N2767);
or OR4 (N3934, N3932, N3192, N1086, N160);
or OR3 (N3935, N3910, N3193, N2913);
and AND2 (N3936, N3922, N2671);
xor XOR2 (N3937, N3935, N3852);
or OR4 (N3938, N3936, N2606, N3107, N2475);
not NOT1 (N3939, N3929);
buf BUF1 (N3940, N3931);
buf BUF1 (N3941, N3933);
nor NOR2 (N3942, N3941, N464);
and AND3 (N3943, N3937, N1895, N1219);
nand NAND2 (N3944, N3934, N1849);
or OR4 (N3945, N3942, N2013, N527, N154);
or OR4 (N3946, N3925, N2761, N2323, N133);
and AND2 (N3947, N3927, N1425);
not NOT1 (N3948, N3943);
xor XOR2 (N3949, N3948, N1311);
nor NOR3 (N3950, N3939, N1606, N2650);
and AND2 (N3951, N3950, N3713);
nor NOR2 (N3952, N3938, N2182);
or OR2 (N3953, N3947, N1239);
buf BUF1 (N3954, N3946);
and AND2 (N3955, N3949, N1275);
not NOT1 (N3956, N3945);
nand NAND4 (N3957, N3955, N2745, N688, N2641);
xor XOR2 (N3958, N3914, N1121);
or OR2 (N3959, N3928, N3174);
buf BUF1 (N3960, N3957);
nor NOR2 (N3961, N3954, N591);
buf BUF1 (N3962, N3960);
nand NAND3 (N3963, N3944, N67, N310);
nor NOR3 (N3964, N3940, N1819, N2643);
nand NAND4 (N3965, N3964, N2128, N1886, N1390);
nor NOR3 (N3966, N3959, N761, N1214);
not NOT1 (N3967, N3952);
nand NAND4 (N3968, N3966, N1806, N1494, N764);
nor NOR2 (N3969, N3968, N3900);
nand NAND2 (N3970, N3965, N2906);
not NOT1 (N3971, N3956);
and AND2 (N3972, N3969, N1773);
xor XOR2 (N3973, N3958, N1067);
not NOT1 (N3974, N3970);
and AND3 (N3975, N3972, N2279, N2390);
nor NOR4 (N3976, N3967, N760, N2458, N2469);
not NOT1 (N3977, N3962);
not NOT1 (N3978, N3953);
not NOT1 (N3979, N3977);
nor NOR2 (N3980, N3973, N2140);
xor XOR2 (N3981, N3961, N1279);
nand NAND4 (N3982, N3951, N3475, N696, N2235);
not NOT1 (N3983, N3979);
nand NAND3 (N3984, N3982, N2848, N3312);
xor XOR2 (N3985, N3981, N1528);
buf BUF1 (N3986, N3974);
not NOT1 (N3987, N3963);
nor NOR2 (N3988, N3983, N703);
buf BUF1 (N3989, N3980);
not NOT1 (N3990, N3976);
buf BUF1 (N3991, N3986);
buf BUF1 (N3992, N3990);
or OR3 (N3993, N3971, N2092, N3810);
nand NAND3 (N3994, N3987, N163, N767);
nand NAND3 (N3995, N3994, N291, N3554);
xor XOR2 (N3996, N3995, N192);
nand NAND4 (N3997, N3989, N3464, N1612, N3623);
nor NOR3 (N3998, N3975, N811, N1599);
nor NOR4 (N3999, N3996, N2371, N2485, N2622);
nand NAND3 (N4000, N3992, N726, N1690);
or OR2 (N4001, N3993, N1687);
nor NOR3 (N4002, N3988, N263, N2156);
and AND3 (N4003, N4000, N1353, N886);
nor NOR3 (N4004, N3991, N2976, N3311);
nand NAND2 (N4005, N3985, N225);
or OR4 (N4006, N4001, N831, N1664, N2335);
buf BUF1 (N4007, N3999);
not NOT1 (N4008, N4005);
nor NOR3 (N4009, N4002, N1399, N3449);
buf BUF1 (N4010, N4004);
xor XOR2 (N4011, N3997, N1123);
nor NOR3 (N4012, N3998, N3979, N2262);
or OR4 (N4013, N4011, N3132, N1424, N2651);
nor NOR4 (N4014, N3978, N2430, N534, N3797);
or OR3 (N4015, N4006, N2175, N690);
buf BUF1 (N4016, N4010);
nand NAND2 (N4017, N4013, N3786);
not NOT1 (N4018, N4016);
nand NAND4 (N4019, N4018, N1153, N3210, N1623);
or OR3 (N4020, N3984, N3030, N3567);
or OR3 (N4021, N4009, N2008, N1894);
nor NOR3 (N4022, N4021, N1265, N63);
nand NAND4 (N4023, N4007, N3058, N794, N208);
xor XOR2 (N4024, N4012, N612);
xor XOR2 (N4025, N4019, N3356);
nand NAND4 (N4026, N4025, N2768, N1138, N1116);
nor NOR2 (N4027, N4024, N743);
nor NOR3 (N4028, N4020, N182, N3095);
xor XOR2 (N4029, N4015, N1418);
buf BUF1 (N4030, N4003);
nor NOR2 (N4031, N4026, N133);
xor XOR2 (N4032, N4008, N3704);
xor XOR2 (N4033, N4017, N2559);
buf BUF1 (N4034, N4022);
or OR3 (N4035, N4029, N1612, N2047);
and AND3 (N4036, N4014, N1013, N527);
buf BUF1 (N4037, N4023);
or OR4 (N4038, N4032, N561, N59, N1274);
nor NOR4 (N4039, N4031, N1644, N3288, N1523);
xor XOR2 (N4040, N4039, N2779);
or OR4 (N4041, N4037, N2711, N505, N3102);
or OR4 (N4042, N4028, N360, N228, N966);
or OR2 (N4043, N4035, N1787);
nand NAND3 (N4044, N4040, N3185, N3177);
nand NAND4 (N4045, N4043, N2511, N89, N445);
and AND3 (N4046, N4042, N1947, N3922);
and AND4 (N4047, N4045, N3052, N483, N864);
buf BUF1 (N4048, N4036);
nand NAND4 (N4049, N4030, N99, N3955, N347);
xor XOR2 (N4050, N4044, N2447);
or OR3 (N4051, N4050, N370, N3230);
or OR3 (N4052, N4046, N24, N873);
and AND3 (N4053, N4052, N510, N399);
and AND3 (N4054, N4027, N537, N3583);
nor NOR4 (N4055, N4041, N3761, N1886, N3316);
nor NOR2 (N4056, N4055, N447);
nor NOR2 (N4057, N4054, N3239);
not NOT1 (N4058, N4034);
buf BUF1 (N4059, N4047);
nor NOR2 (N4060, N4048, N3815);
nand NAND3 (N4061, N4038, N1070, N165);
buf BUF1 (N4062, N4060);
and AND4 (N4063, N4058, N1522, N2784, N3088);
nor NOR2 (N4064, N4056, N3623);
nand NAND3 (N4065, N4064, N1848, N92);
not NOT1 (N4066, N4051);
not NOT1 (N4067, N4066);
not NOT1 (N4068, N4059);
nand NAND4 (N4069, N4062, N2364, N3658, N3409);
buf BUF1 (N4070, N4068);
buf BUF1 (N4071, N4070);
nand NAND4 (N4072, N4065, N1477, N3194, N2872);
buf BUF1 (N4073, N4061);
not NOT1 (N4074, N4071);
xor XOR2 (N4075, N4057, N917);
buf BUF1 (N4076, N4053);
and AND3 (N4077, N4074, N3166, N2385);
or OR2 (N4078, N4033, N1670);
or OR3 (N4079, N4077, N2181, N1669);
buf BUF1 (N4080, N4076);
nor NOR3 (N4081, N4049, N1986, N3522);
not NOT1 (N4082, N4078);
nand NAND2 (N4083, N4079, N1897);
buf BUF1 (N4084, N4083);
not NOT1 (N4085, N4075);
buf BUF1 (N4086, N4067);
nand NAND4 (N4087, N4084, N3628, N3570, N792);
and AND3 (N4088, N4087, N2337, N690);
or OR4 (N4089, N4072, N1766, N866, N3449);
and AND4 (N4090, N4063, N1422, N1446, N2416);
xor XOR2 (N4091, N4086, N3300);
xor XOR2 (N4092, N4085, N2260);
xor XOR2 (N4093, N4073, N2637);
not NOT1 (N4094, N4069);
not NOT1 (N4095, N4088);
or OR2 (N4096, N4082, N2672);
and AND3 (N4097, N4081, N3819, N3172);
not NOT1 (N4098, N4096);
or OR4 (N4099, N4093, N3191, N2951, N1887);
or OR3 (N4100, N4092, N3140, N166);
buf BUF1 (N4101, N4094);
nor NOR2 (N4102, N4091, N169);
nor NOR2 (N4103, N4099, N2262);
nand NAND4 (N4104, N4090, N1528, N1193, N3698);
and AND3 (N4105, N4101, N4041, N2629);
nor NOR3 (N4106, N4105, N1067, N3453);
nand NAND4 (N4107, N4100, N2067, N1574, N1796);
buf BUF1 (N4108, N4097);
nand NAND4 (N4109, N4080, N447, N2718, N1450);
nand NAND3 (N4110, N4108, N3547, N2304);
or OR2 (N4111, N4104, N849);
or OR3 (N4112, N4095, N1657, N887);
not NOT1 (N4113, N4102);
not NOT1 (N4114, N4089);
nor NOR4 (N4115, N4114, N2330, N1137, N1924);
nor NOR2 (N4116, N4107, N1035);
nand NAND4 (N4117, N4115, N1679, N9, N2876);
xor XOR2 (N4118, N4098, N25);
nor NOR3 (N4119, N4112, N85, N3040);
nor NOR3 (N4120, N4111, N339, N2802);
buf BUF1 (N4121, N4120);
nor NOR2 (N4122, N4103, N1580);
and AND4 (N4123, N4109, N1749, N1037, N3832);
buf BUF1 (N4124, N4110);
not NOT1 (N4125, N4122);
or OR4 (N4126, N4123, N1621, N1531, N623);
nand NAND3 (N4127, N4121, N143, N835);
not NOT1 (N4128, N4117);
or OR4 (N4129, N4119, N3322, N1313, N2373);
not NOT1 (N4130, N4124);
buf BUF1 (N4131, N4127);
not NOT1 (N4132, N4125);
buf BUF1 (N4133, N4118);
xor XOR2 (N4134, N4130, N2773);
nand NAND3 (N4135, N4131, N1039, N1922);
nand NAND3 (N4136, N4129, N2443, N2037);
not NOT1 (N4137, N4113);
xor XOR2 (N4138, N4128, N1266);
or OR3 (N4139, N4137, N1952, N1895);
not NOT1 (N4140, N4139);
not NOT1 (N4141, N4140);
or OR3 (N4142, N4136, N2562, N3318);
nand NAND2 (N4143, N4141, N2243);
not NOT1 (N4144, N4132);
and AND2 (N4145, N4142, N100);
buf BUF1 (N4146, N4116);
nand NAND2 (N4147, N4138, N1547);
not NOT1 (N4148, N4147);
and AND3 (N4149, N4134, N3899, N1319);
not NOT1 (N4150, N4149);
nor NOR4 (N4151, N4146, N3353, N3917, N3775);
or OR2 (N4152, N4151, N1633);
buf BUF1 (N4153, N4145);
xor XOR2 (N4154, N4135, N2143);
not NOT1 (N4155, N4143);
nand NAND3 (N4156, N4126, N183, N2516);
and AND2 (N4157, N4148, N481);
and AND3 (N4158, N4152, N1378, N690);
not NOT1 (N4159, N4154);
xor XOR2 (N4160, N4144, N1640);
nand NAND2 (N4161, N4153, N3818);
nor NOR4 (N4162, N4133, N3208, N1565, N4050);
nand NAND4 (N4163, N4106, N3971, N3701, N563);
xor XOR2 (N4164, N4150, N2820);
xor XOR2 (N4165, N4159, N2749);
not NOT1 (N4166, N4155);
not NOT1 (N4167, N4160);
not NOT1 (N4168, N4162);
nand NAND4 (N4169, N4165, N2022, N2934, N1211);
nand NAND2 (N4170, N4163, N1309);
or OR4 (N4171, N4161, N3087, N544, N1550);
nand NAND4 (N4172, N4156, N290, N2880, N444);
xor XOR2 (N4173, N4157, N1254);
buf BUF1 (N4174, N4170);
xor XOR2 (N4175, N4174, N2673);
nor NOR4 (N4176, N4169, N1327, N3016, N1174);
nor NOR3 (N4177, N4158, N846, N2739);
nand NAND3 (N4178, N4171, N3275, N2626);
nor NOR2 (N4179, N4168, N3089);
nor NOR3 (N4180, N4178, N3434, N2416);
and AND4 (N4181, N4175, N2744, N3048, N3861);
nor NOR2 (N4182, N4164, N4164);
and AND2 (N4183, N4172, N1638);
nor NOR2 (N4184, N4182, N2979);
xor XOR2 (N4185, N4180, N1176);
or OR2 (N4186, N4177, N1915);
buf BUF1 (N4187, N4176);
xor XOR2 (N4188, N4185, N626);
and AND3 (N4189, N4186, N2694, N3711);
and AND3 (N4190, N4167, N2776, N2470);
xor XOR2 (N4191, N4166, N2167);
xor XOR2 (N4192, N4187, N3257);
or OR4 (N4193, N4173, N1774, N3116, N3588);
or OR3 (N4194, N4179, N213, N778);
not NOT1 (N4195, N4184);
nor NOR3 (N4196, N4189, N158, N3774);
and AND2 (N4197, N4193, N1327);
nor NOR3 (N4198, N4181, N846, N891);
nand NAND2 (N4199, N4197, N3213);
xor XOR2 (N4200, N4192, N4152);
or OR4 (N4201, N4198, N3734, N2945, N916);
or OR3 (N4202, N4201, N3462, N2836);
xor XOR2 (N4203, N4199, N2327);
and AND3 (N4204, N4203, N2995, N837);
xor XOR2 (N4205, N4202, N875);
buf BUF1 (N4206, N4194);
nor NOR4 (N4207, N4204, N3412, N3131, N2484);
and AND2 (N4208, N4205, N1275);
not NOT1 (N4209, N4188);
nand NAND4 (N4210, N4206, N3285, N980, N2023);
xor XOR2 (N4211, N4190, N3558);
or OR2 (N4212, N4210, N1746);
and AND3 (N4213, N4212, N3151, N1390);
nor NOR4 (N4214, N4207, N2076, N3102, N601);
and AND2 (N4215, N4213, N712);
and AND2 (N4216, N4215, N1647);
not NOT1 (N4217, N4209);
not NOT1 (N4218, N4214);
buf BUF1 (N4219, N4183);
and AND4 (N4220, N4211, N4092, N2331, N3128);
nand NAND2 (N4221, N4195, N1551);
nor NOR3 (N4222, N4200, N4017, N1349);
buf BUF1 (N4223, N4222);
and AND3 (N4224, N4217, N4118, N2545);
or OR2 (N4225, N4223, N1133);
nor NOR3 (N4226, N4221, N670, N808);
or OR2 (N4227, N4226, N3501);
nor NOR4 (N4228, N4196, N3950, N3162, N3778);
buf BUF1 (N4229, N4224);
buf BUF1 (N4230, N4220);
buf BUF1 (N4231, N4219);
nand NAND3 (N4232, N4227, N3889, N1614);
and AND3 (N4233, N4232, N2871, N2419);
and AND3 (N4234, N4216, N3375, N3213);
nand NAND2 (N4235, N4229, N1898);
and AND4 (N4236, N4228, N2261, N4155, N156);
and AND3 (N4237, N4191, N3887, N1537);
buf BUF1 (N4238, N4225);
nor NOR4 (N4239, N4237, N3521, N3550, N3405);
buf BUF1 (N4240, N4239);
buf BUF1 (N4241, N4218);
and AND4 (N4242, N4208, N1343, N639, N1409);
or OR4 (N4243, N4241, N1458, N2224, N4021);
buf BUF1 (N4244, N4235);
xor XOR2 (N4245, N4233, N2344);
and AND3 (N4246, N4234, N3635, N935);
not NOT1 (N4247, N4238);
nand NAND3 (N4248, N4231, N663, N2526);
nand NAND2 (N4249, N4245, N1990);
nand NAND3 (N4250, N4247, N832, N1833);
or OR4 (N4251, N4249, N717, N267, N1260);
buf BUF1 (N4252, N4240);
or OR3 (N4253, N4246, N2791, N2952);
xor XOR2 (N4254, N4236, N385);
nand NAND3 (N4255, N4243, N2452, N321);
and AND3 (N4256, N4253, N1082, N3904);
nor NOR4 (N4257, N4242, N3388, N3603, N4252);
xor XOR2 (N4258, N3470, N1309);
nand NAND4 (N4259, N4256, N173, N2946, N1075);
buf BUF1 (N4260, N4258);
not NOT1 (N4261, N4250);
not NOT1 (N4262, N4257);
or OR4 (N4263, N4254, N1302, N3896, N2841);
xor XOR2 (N4264, N4255, N3892);
nand NAND4 (N4265, N4230, N3341, N2175, N1972);
or OR3 (N4266, N4244, N1523, N3615);
not NOT1 (N4267, N4264);
xor XOR2 (N4268, N4262, N3198);
nor NOR2 (N4269, N4267, N1675);
not NOT1 (N4270, N4248);
not NOT1 (N4271, N4269);
not NOT1 (N4272, N4270);
buf BUF1 (N4273, N4261);
or OR4 (N4274, N4268, N1583, N2331, N349);
buf BUF1 (N4275, N4274);
not NOT1 (N4276, N4263);
and AND2 (N4277, N4272, N3053);
or OR2 (N4278, N4275, N3517);
xor XOR2 (N4279, N4251, N2775);
nand NAND4 (N4280, N4273, N1773, N392, N2746);
or OR4 (N4281, N4279, N1572, N4161, N2496);
xor XOR2 (N4282, N4266, N89);
or OR3 (N4283, N4280, N2699, N21);
nand NAND3 (N4284, N4265, N2407, N48);
nor NOR3 (N4285, N4281, N74, N2822);
and AND2 (N4286, N4260, N1003);
or OR2 (N4287, N4278, N2212);
xor XOR2 (N4288, N4285, N730);
and AND3 (N4289, N4277, N3213, N1737);
nor NOR3 (N4290, N4286, N657, N1099);
nor NOR4 (N4291, N4282, N1044, N395, N1952);
buf BUF1 (N4292, N4271);
or OR3 (N4293, N4288, N3497, N1520);
nor NOR3 (N4294, N4290, N1703, N1820);
xor XOR2 (N4295, N4292, N249);
and AND3 (N4296, N4295, N1917, N2042);
nor NOR2 (N4297, N4283, N875);
buf BUF1 (N4298, N4296);
and AND2 (N4299, N4287, N3356);
nor NOR3 (N4300, N4289, N3792, N451);
not NOT1 (N4301, N4300);
nand NAND4 (N4302, N4299, N1978, N3911, N629);
not NOT1 (N4303, N4294);
or OR2 (N4304, N4303, N2016);
nor NOR4 (N4305, N4304, N3156, N301, N3227);
nor NOR4 (N4306, N4305, N4110, N101, N1131);
and AND2 (N4307, N4297, N1128);
nand NAND2 (N4308, N4293, N3963);
buf BUF1 (N4309, N4307);
not NOT1 (N4310, N4309);
or OR3 (N4311, N4284, N1012, N2192);
and AND3 (N4312, N4276, N773, N594);
xor XOR2 (N4313, N4298, N2745);
and AND3 (N4314, N4313, N1983, N3225);
and AND2 (N4315, N4308, N3806);
or OR3 (N4316, N4310, N401, N3309);
nand NAND4 (N4317, N4314, N1598, N3920, N3723);
xor XOR2 (N4318, N4306, N301);
and AND2 (N4319, N4259, N3800);
not NOT1 (N4320, N4302);
and AND3 (N4321, N4291, N883, N1771);
nand NAND4 (N4322, N4312, N1061, N245, N3559);
or OR3 (N4323, N4322, N3527, N2904);
and AND3 (N4324, N4315, N2338, N2466);
buf BUF1 (N4325, N4319);
buf BUF1 (N4326, N4317);
xor XOR2 (N4327, N4321, N1408);
and AND2 (N4328, N4324, N1474);
nor NOR4 (N4329, N4328, N3913, N3411, N161);
not NOT1 (N4330, N4311);
xor XOR2 (N4331, N4320, N1616);
and AND3 (N4332, N4329, N3815, N150);
or OR4 (N4333, N4301, N3528, N3871, N75);
xor XOR2 (N4334, N4330, N3534);
buf BUF1 (N4335, N4316);
and AND4 (N4336, N4331, N240, N1524, N4097);
nor NOR4 (N4337, N4332, N716, N4009, N626);
nor NOR2 (N4338, N4326, N3500);
nand NAND3 (N4339, N4335, N1563, N2096);
and AND3 (N4340, N4333, N2009, N350);
and AND4 (N4341, N4340, N2404, N519, N2790);
nand NAND2 (N4342, N4323, N4238);
nand NAND4 (N4343, N4318, N1175, N2991, N3992);
and AND3 (N4344, N4327, N2464, N3638);
nand NAND3 (N4345, N4325, N4096, N1417);
or OR3 (N4346, N4336, N1806, N1037);
nand NAND4 (N4347, N4342, N892, N1719, N2803);
not NOT1 (N4348, N4334);
nand NAND3 (N4349, N4348, N2429, N2305);
not NOT1 (N4350, N4344);
buf BUF1 (N4351, N4345);
not NOT1 (N4352, N4339);
not NOT1 (N4353, N4347);
or OR2 (N4354, N4338, N4319);
nand NAND2 (N4355, N4341, N3955);
nand NAND2 (N4356, N4351, N3853);
xor XOR2 (N4357, N4352, N820);
xor XOR2 (N4358, N4343, N3788);
buf BUF1 (N4359, N4346);
nand NAND3 (N4360, N4357, N1883, N3396);
nor NOR2 (N4361, N4356, N158);
and AND4 (N4362, N4354, N275, N1866, N4264);
and AND2 (N4363, N4358, N912);
not NOT1 (N4364, N4349);
nand NAND4 (N4365, N4363, N1354, N1232, N4363);
and AND3 (N4366, N4362, N306, N178);
nor NOR4 (N4367, N4350, N1211, N2895, N3941);
nor NOR2 (N4368, N4360, N3062);
nor NOR2 (N4369, N4359, N2406);
and AND2 (N4370, N4367, N3855);
buf BUF1 (N4371, N4353);
and AND3 (N4372, N4355, N3518, N2635);
nand NAND3 (N4373, N4372, N2364, N1487);
buf BUF1 (N4374, N4368);
and AND2 (N4375, N4366, N1077);
and AND3 (N4376, N4370, N820, N481);
xor XOR2 (N4377, N4373, N2571);
not NOT1 (N4378, N4375);
xor XOR2 (N4379, N4337, N2574);
nand NAND2 (N4380, N4365, N64);
xor XOR2 (N4381, N4371, N1932);
nor NOR4 (N4382, N4374, N2400, N1318, N246);
xor XOR2 (N4383, N4379, N452);
xor XOR2 (N4384, N4376, N1830);
xor XOR2 (N4385, N4377, N1633);
nor NOR2 (N4386, N4381, N2279);
nand NAND2 (N4387, N4382, N1032);
nor NOR4 (N4388, N4387, N1338, N2544, N3299);
nand NAND2 (N4389, N4385, N2193);
not NOT1 (N4390, N4383);
xor XOR2 (N4391, N4384, N2596);
not NOT1 (N4392, N4364);
and AND4 (N4393, N4386, N3830, N3380, N187);
and AND2 (N4394, N4388, N3127);
xor XOR2 (N4395, N4389, N2784);
buf BUF1 (N4396, N4380);
xor XOR2 (N4397, N4396, N1187);
or OR3 (N4398, N4394, N2356, N1108);
buf BUF1 (N4399, N4397);
or OR3 (N4400, N4399, N2597, N854);
xor XOR2 (N4401, N4400, N3908);
xor XOR2 (N4402, N4369, N2507);
not NOT1 (N4403, N4401);
xor XOR2 (N4404, N4403, N3292);
buf BUF1 (N4405, N4378);
or OR3 (N4406, N4361, N1941, N2508);
or OR3 (N4407, N4402, N1565, N1528);
or OR4 (N4408, N4393, N1404, N2658, N3253);
not NOT1 (N4409, N4408);
nand NAND3 (N4410, N4392, N2579, N900);
nand NAND2 (N4411, N4398, N4090);
nand NAND4 (N4412, N4395, N4066, N1658, N16);
and AND2 (N4413, N4407, N66);
or OR3 (N4414, N4409, N1786, N2199);
and AND4 (N4415, N4391, N887, N3027, N2777);
nand NAND4 (N4416, N4412, N3721, N1942, N1560);
buf BUF1 (N4417, N4416);
or OR4 (N4418, N4406, N2487, N1929, N1202);
buf BUF1 (N4419, N4410);
nor NOR4 (N4420, N4405, N3371, N1608, N2764);
nand NAND3 (N4421, N4419, N4348, N3151);
not NOT1 (N4422, N4413);
xor XOR2 (N4423, N4418, N2124);
nor NOR2 (N4424, N4422, N124);
nand NAND4 (N4425, N4424, N2739, N4089, N3678);
nand NAND4 (N4426, N4411, N2044, N743, N702);
xor XOR2 (N4427, N4417, N1354);
not NOT1 (N4428, N4425);
xor XOR2 (N4429, N4415, N2510);
nand NAND4 (N4430, N4423, N516, N833, N1010);
nor NOR4 (N4431, N4426, N2820, N3324, N3745);
and AND4 (N4432, N4421, N299, N2797, N1444);
not NOT1 (N4433, N4428);
and AND4 (N4434, N4433, N540, N1416, N2144);
nor NOR4 (N4435, N4434, N1513, N3536, N241);
nand NAND2 (N4436, N4420, N2179);
or OR3 (N4437, N4404, N3770, N2110);
nor NOR2 (N4438, N4435, N340);
or OR2 (N4439, N4437, N926);
not NOT1 (N4440, N4439);
or OR4 (N4441, N4438, N385, N91, N2454);
or OR2 (N4442, N4427, N1447);
nand NAND2 (N4443, N4441, N3235);
and AND3 (N4444, N4432, N782, N2998);
xor XOR2 (N4445, N4436, N3593);
nor NOR3 (N4446, N4429, N2958, N13);
and AND4 (N4447, N4442, N768, N3311, N3959);
nand NAND3 (N4448, N4447, N650, N3783);
not NOT1 (N4449, N4445);
not NOT1 (N4450, N4443);
and AND4 (N4451, N4450, N1663, N4448, N1440);
not NOT1 (N4452, N56);
or OR4 (N4453, N4430, N3502, N2162, N3734);
and AND2 (N4454, N4444, N802);
buf BUF1 (N4455, N4449);
buf BUF1 (N4456, N4446);
not NOT1 (N4457, N4455);
xor XOR2 (N4458, N4457, N3061);
nor NOR2 (N4459, N4454, N3406);
and AND4 (N4460, N4390, N656, N962, N435);
not NOT1 (N4461, N4453);
or OR2 (N4462, N4456, N633);
xor XOR2 (N4463, N4462, N2295);
or OR3 (N4464, N4463, N1658, N3966);
buf BUF1 (N4465, N4431);
xor XOR2 (N4466, N4461, N223);
buf BUF1 (N4467, N4466);
nor NOR4 (N4468, N4459, N1293, N4183, N1817);
and AND3 (N4469, N4460, N563, N4159);
or OR4 (N4470, N4452, N3963, N3393, N768);
nor NOR2 (N4471, N4468, N3066);
nand NAND3 (N4472, N4414, N2817, N1905);
xor XOR2 (N4473, N4472, N4257);
nand NAND2 (N4474, N4470, N4279);
nor NOR3 (N4475, N4464, N47, N2545);
xor XOR2 (N4476, N4475, N4012);
nand NAND4 (N4477, N4469, N2181, N3335, N2205);
not NOT1 (N4478, N4467);
or OR2 (N4479, N4440, N1376);
nor NOR2 (N4480, N4476, N4436);
buf BUF1 (N4481, N4478);
nand NAND3 (N4482, N4481, N1983, N2347);
nand NAND3 (N4483, N4458, N509, N3311);
not NOT1 (N4484, N4451);
buf BUF1 (N4485, N4484);
nor NOR3 (N4486, N4474, N3661, N2683);
and AND4 (N4487, N4471, N1447, N2394, N115);
buf BUF1 (N4488, N4483);
and AND4 (N4489, N4487, N952, N3357, N2759);
nor NOR2 (N4490, N4473, N1101);
not NOT1 (N4491, N4477);
not NOT1 (N4492, N4490);
or OR3 (N4493, N4488, N3751, N279);
xor XOR2 (N4494, N4492, N541);
not NOT1 (N4495, N4465);
or OR2 (N4496, N4495, N1860);
nand NAND2 (N4497, N4493, N3242);
nand NAND4 (N4498, N4482, N3283, N407, N352);
nor NOR3 (N4499, N4497, N3444, N585);
xor XOR2 (N4500, N4494, N283);
not NOT1 (N4501, N4499);
nand NAND3 (N4502, N4491, N3776, N2694);
nand NAND4 (N4503, N4500, N2001, N3409, N3761);
or OR2 (N4504, N4496, N2998);
not NOT1 (N4505, N4501);
nand NAND3 (N4506, N4485, N3740, N3827);
buf BUF1 (N4507, N4505);
xor XOR2 (N4508, N4486, N1707);
nand NAND2 (N4509, N4506, N4390);
nor NOR3 (N4510, N4479, N3093, N2402);
or OR2 (N4511, N4508, N52);
xor XOR2 (N4512, N4509, N8);
not NOT1 (N4513, N4511);
and AND3 (N4514, N4503, N3102, N816);
or OR4 (N4515, N4512, N3749, N1562, N1828);
and AND4 (N4516, N4480, N1909, N1075, N898);
and AND2 (N4517, N4514, N2022);
nor NOR4 (N4518, N4513, N2449, N3767, N2523);
and AND4 (N4519, N4502, N101, N1388, N572);
and AND3 (N4520, N4516, N1299, N880);
or OR4 (N4521, N4498, N706, N3276, N2944);
nor NOR3 (N4522, N4515, N1010, N1543);
xor XOR2 (N4523, N4489, N2212);
nand NAND2 (N4524, N4507, N1086);
buf BUF1 (N4525, N4524);
not NOT1 (N4526, N4521);
nor NOR4 (N4527, N4510, N3155, N4129, N840);
nand NAND4 (N4528, N4526, N2280, N3723, N1227);
and AND2 (N4529, N4519, N4086);
xor XOR2 (N4530, N4523, N2033);
nor NOR3 (N4531, N4528, N1986, N894);
or OR3 (N4532, N4525, N4051, N3635);
buf BUF1 (N4533, N4532);
not NOT1 (N4534, N4531);
nand NAND2 (N4535, N4504, N3638);
nand NAND3 (N4536, N4529, N3961, N2134);
xor XOR2 (N4537, N4527, N1343);
nor NOR4 (N4538, N4517, N1871, N2742, N2108);
or OR3 (N4539, N4518, N4114, N3344);
xor XOR2 (N4540, N4536, N4143);
xor XOR2 (N4541, N4538, N2213);
or OR2 (N4542, N4537, N1123);
buf BUF1 (N4543, N4522);
and AND2 (N4544, N4539, N2803);
xor XOR2 (N4545, N4544, N2633);
not NOT1 (N4546, N4530);
and AND4 (N4547, N4546, N2618, N2518, N2777);
nand NAND3 (N4548, N4520, N891, N3672);
nand NAND3 (N4549, N4543, N2720, N3911);
not NOT1 (N4550, N4535);
nor NOR2 (N4551, N4545, N1541);
not NOT1 (N4552, N4533);
xor XOR2 (N4553, N4547, N1814);
not NOT1 (N4554, N4540);
nand NAND2 (N4555, N4548, N175);
and AND4 (N4556, N4550, N2647, N1630, N879);
buf BUF1 (N4557, N4541);
buf BUF1 (N4558, N4549);
nand NAND2 (N4559, N4552, N3861);
nand NAND3 (N4560, N4554, N1955, N3974);
nor NOR4 (N4561, N4557, N3158, N4298, N1160);
nand NAND4 (N4562, N4559, N3970, N3438, N1213);
or OR3 (N4563, N4551, N1601, N485);
not NOT1 (N4564, N4553);
nor NOR3 (N4565, N4560, N879, N2395);
not NOT1 (N4566, N4556);
nand NAND3 (N4567, N4566, N4032, N3944);
nand NAND2 (N4568, N4564, N789);
nor NOR3 (N4569, N4567, N1517, N1130);
buf BUF1 (N4570, N4563);
buf BUF1 (N4571, N4568);
buf BUF1 (N4572, N4534);
nor NOR4 (N4573, N4565, N876, N3388, N4342);
nor NOR3 (N4574, N4562, N3118, N3459);
buf BUF1 (N4575, N4569);
not NOT1 (N4576, N4561);
xor XOR2 (N4577, N4542, N1003);
buf BUF1 (N4578, N4555);
nand NAND2 (N4579, N4575, N381);
buf BUF1 (N4580, N4579);
buf BUF1 (N4581, N4570);
nor NOR2 (N4582, N4577, N1783);
nand NAND4 (N4583, N4574, N4076, N2716, N1263);
xor XOR2 (N4584, N4558, N2151);
not NOT1 (N4585, N4572);
or OR4 (N4586, N4581, N4310, N1617, N2920);
xor XOR2 (N4587, N4585, N2589);
xor XOR2 (N4588, N4576, N33);
xor XOR2 (N4589, N4586, N1464);
or OR4 (N4590, N4582, N3400, N2, N1172);
buf BUF1 (N4591, N4588);
or OR3 (N4592, N4578, N3927, N1477);
or OR4 (N4593, N4584, N2321, N4278, N2136);
xor XOR2 (N4594, N4571, N859);
buf BUF1 (N4595, N4589);
buf BUF1 (N4596, N4580);
and AND3 (N4597, N4593, N4152, N2432);
and AND4 (N4598, N4583, N3678, N1179, N1508);
nand NAND3 (N4599, N4592, N4244, N2745);
or OR3 (N4600, N4599, N3946, N2472);
xor XOR2 (N4601, N4595, N1089);
nand NAND2 (N4602, N4573, N1353);
nand NAND4 (N4603, N4598, N1398, N4192, N1389);
and AND4 (N4604, N4602, N2594, N3865, N558);
nand NAND4 (N4605, N4596, N2212, N1496, N2457);
xor XOR2 (N4606, N4590, N3375);
and AND3 (N4607, N4600, N1208, N2798);
and AND3 (N4608, N4606, N926, N3310);
not NOT1 (N4609, N4605);
or OR2 (N4610, N4591, N2852);
not NOT1 (N4611, N4608);
nor NOR4 (N4612, N4610, N2269, N1651, N3582);
and AND2 (N4613, N4611, N488);
and AND3 (N4614, N4609, N748, N3835);
or OR2 (N4615, N4597, N1420);
nand NAND2 (N4616, N4614, N749);
xor XOR2 (N4617, N4603, N4204);
nand NAND3 (N4618, N4607, N3665, N328);
nor NOR4 (N4619, N4618, N2821, N503, N657);
or OR2 (N4620, N4601, N1352);
xor XOR2 (N4621, N4604, N1253);
and AND2 (N4622, N4619, N4046);
buf BUF1 (N4623, N4612);
not NOT1 (N4624, N4615);
xor XOR2 (N4625, N4622, N175);
or OR2 (N4626, N4594, N2017);
nand NAND4 (N4627, N4616, N3615, N4538, N170);
xor XOR2 (N4628, N4617, N993);
or OR3 (N4629, N4624, N1613, N4502);
not NOT1 (N4630, N4623);
not NOT1 (N4631, N4628);
and AND3 (N4632, N4621, N3728, N2779);
xor XOR2 (N4633, N4613, N3476);
nand NAND3 (N4634, N4620, N3066, N3593);
xor XOR2 (N4635, N4634, N444);
nand NAND4 (N4636, N4626, N2522, N2487, N2728);
or OR2 (N4637, N4633, N3440);
xor XOR2 (N4638, N4632, N3603);
buf BUF1 (N4639, N4638);
and AND2 (N4640, N4625, N2612);
or OR3 (N4641, N4636, N1923, N243);
xor XOR2 (N4642, N4637, N1944);
nand NAND2 (N4643, N4640, N2151);
or OR4 (N4644, N4631, N3126, N3855, N4384);
nor NOR4 (N4645, N4643, N961, N49, N476);
buf BUF1 (N4646, N4627);
or OR4 (N4647, N4642, N1414, N767, N1699);
or OR4 (N4648, N4644, N1361, N3343, N2936);
nand NAND4 (N4649, N4645, N1553, N576, N1774);
and AND2 (N4650, N4646, N569);
and AND3 (N4651, N4630, N3341, N2947);
and AND2 (N4652, N4648, N2412);
nand NAND3 (N4653, N4635, N442, N3761);
and AND2 (N4654, N4647, N4229);
buf BUF1 (N4655, N4653);
xor XOR2 (N4656, N4649, N2705);
xor XOR2 (N4657, N4650, N3124);
or OR3 (N4658, N4639, N1187, N1269);
xor XOR2 (N4659, N4657, N1703);
nand NAND4 (N4660, N4654, N3869, N2616, N1890);
and AND3 (N4661, N4660, N1334, N327);
and AND2 (N4662, N4641, N2778);
xor XOR2 (N4663, N4629, N2532);
not NOT1 (N4664, N4661);
buf BUF1 (N4665, N4655);
buf BUF1 (N4666, N4656);
not NOT1 (N4667, N4666);
or OR4 (N4668, N4658, N3815, N3690, N1215);
buf BUF1 (N4669, N4667);
nor NOR3 (N4670, N4665, N2710, N2198);
nor NOR4 (N4671, N4587, N4335, N4508, N1526);
buf BUF1 (N4672, N4671);
xor XOR2 (N4673, N4652, N3583);
buf BUF1 (N4674, N4659);
nor NOR2 (N4675, N4663, N2757);
not NOT1 (N4676, N4669);
nand NAND2 (N4677, N4675, N4256);
and AND4 (N4678, N4670, N1963, N2198, N1396);
not NOT1 (N4679, N4673);
nor NOR4 (N4680, N4664, N236, N586, N3395);
xor XOR2 (N4681, N4662, N457);
nor NOR3 (N4682, N4680, N1782, N483);
and AND4 (N4683, N4676, N1749, N1958, N3610);
buf BUF1 (N4684, N4683);
buf BUF1 (N4685, N4672);
xor XOR2 (N4686, N4651, N1026);
or OR4 (N4687, N4686, N396, N2511, N3352);
not NOT1 (N4688, N4668);
xor XOR2 (N4689, N4677, N513);
not NOT1 (N4690, N4674);
or OR4 (N4691, N4689, N2828, N4681, N3815);
nor NOR2 (N4692, N627, N2858);
xor XOR2 (N4693, N4691, N1221);
xor XOR2 (N4694, N4690, N323);
not NOT1 (N4695, N4687);
xor XOR2 (N4696, N4688, N161);
not NOT1 (N4697, N4695);
nand NAND2 (N4698, N4694, N338);
nand NAND4 (N4699, N4698, N2685, N1186, N4029);
nand NAND3 (N4700, N4693, N356, N2883);
not NOT1 (N4701, N4678);
nor NOR4 (N4702, N4684, N2069, N1239, N3464);
buf BUF1 (N4703, N4701);
nor NOR2 (N4704, N4699, N3727);
buf BUF1 (N4705, N4703);
nor NOR3 (N4706, N4679, N2574, N659);
and AND2 (N4707, N4700, N649);
and AND4 (N4708, N4696, N2553, N3188, N310);
and AND2 (N4709, N4707, N504);
or OR4 (N4710, N4682, N1153, N3628, N2145);
nand NAND2 (N4711, N4705, N2024);
xor XOR2 (N4712, N4711, N322);
or OR4 (N4713, N4692, N4556, N952, N3907);
buf BUF1 (N4714, N4685);
and AND4 (N4715, N4712, N2404, N4537, N1408);
or OR3 (N4716, N4710, N886, N3144);
and AND2 (N4717, N4714, N1954);
or OR3 (N4718, N4715, N1338, N1707);
or OR3 (N4719, N4717, N3816, N473);
and AND4 (N4720, N4709, N319, N1538, N4154);
nor NOR2 (N4721, N4718, N1709);
nand NAND3 (N4722, N4708, N3462, N4444);
nor NOR3 (N4723, N4722, N2284, N1908);
xor XOR2 (N4724, N4720, N3547);
nand NAND4 (N4725, N4724, N2478, N4648, N3377);
xor XOR2 (N4726, N4719, N4231);
not NOT1 (N4727, N4713);
nand NAND4 (N4728, N4716, N4074, N3030, N4697);
not NOT1 (N4729, N708);
and AND4 (N4730, N4704, N2755, N30, N1003);
or OR2 (N4731, N4725, N2928);
or OR4 (N4732, N4731, N1726, N172, N2427);
xor XOR2 (N4733, N4732, N3625);
and AND3 (N4734, N4702, N3516, N2494);
and AND3 (N4735, N4730, N1686, N653);
nand NAND2 (N4736, N4728, N1823);
not NOT1 (N4737, N4727);
not NOT1 (N4738, N4726);
not NOT1 (N4739, N4738);
or OR2 (N4740, N4706, N3056);
buf BUF1 (N4741, N4739);
nand NAND3 (N4742, N4721, N421, N1625);
xor XOR2 (N4743, N4735, N2666);
xor XOR2 (N4744, N4736, N3800);
xor XOR2 (N4745, N4742, N4029);
nor NOR2 (N4746, N4734, N4040);
nand NAND2 (N4747, N4741, N3427);
or OR2 (N4748, N4729, N2514);
xor XOR2 (N4749, N4745, N2109);
not NOT1 (N4750, N4746);
buf BUF1 (N4751, N4737);
buf BUF1 (N4752, N4740);
buf BUF1 (N4753, N4749);
nand NAND4 (N4754, N4750, N406, N4180, N2638);
not NOT1 (N4755, N4754);
or OR3 (N4756, N4753, N2446, N791);
nand NAND3 (N4757, N4744, N3792, N1983);
or OR4 (N4758, N4756, N690, N1605, N2940);
not NOT1 (N4759, N4751);
nor NOR3 (N4760, N4759, N397, N755);
or OR2 (N4761, N4748, N2119);
not NOT1 (N4762, N4761);
nor NOR2 (N4763, N4762, N3157);
nand NAND2 (N4764, N4760, N1346);
or OR3 (N4765, N4747, N3016, N3293);
and AND4 (N4766, N4755, N3740, N1406, N2865);
not NOT1 (N4767, N4743);
nand NAND3 (N4768, N4752, N1207, N1824);
or OR4 (N4769, N4765, N2675, N4710, N2852);
and AND2 (N4770, N4766, N4323);
nor NOR3 (N4771, N4733, N1641, N4280);
xor XOR2 (N4772, N4768, N4354);
nand NAND3 (N4773, N4770, N4651, N1795);
buf BUF1 (N4774, N4773);
or OR3 (N4775, N4769, N296, N1981);
nand NAND3 (N4776, N4774, N1525, N668);
xor XOR2 (N4777, N4758, N4252);
nor NOR3 (N4778, N4771, N2781, N4759);
not NOT1 (N4779, N4775);
nand NAND2 (N4780, N4772, N547);
buf BUF1 (N4781, N4757);
buf BUF1 (N4782, N4778);
nor NOR2 (N4783, N4781, N3675);
or OR2 (N4784, N4780, N2436);
buf BUF1 (N4785, N4782);
xor XOR2 (N4786, N4784, N2036);
or OR2 (N4787, N4785, N638);
buf BUF1 (N4788, N4764);
or OR4 (N4789, N4776, N3215, N2565, N897);
not NOT1 (N4790, N4789);
not NOT1 (N4791, N4723);
nand NAND3 (N4792, N4791, N4733, N2167);
nand NAND2 (N4793, N4767, N1679);
nor NOR4 (N4794, N4786, N364, N3061, N4681);
buf BUF1 (N4795, N4783);
and AND4 (N4796, N4777, N2870, N157, N701);
nand NAND4 (N4797, N4793, N1877, N4776, N3453);
not NOT1 (N4798, N4779);
nand NAND4 (N4799, N4763, N1687, N2032, N4572);
or OR4 (N4800, N4796, N3570, N220, N731);
xor XOR2 (N4801, N4797, N2925);
buf BUF1 (N4802, N4787);
buf BUF1 (N4803, N4802);
buf BUF1 (N4804, N4798);
xor XOR2 (N4805, N4801, N1147);
xor XOR2 (N4806, N4804, N3201);
buf BUF1 (N4807, N4792);
nand NAND3 (N4808, N4805, N3932, N3119);
not NOT1 (N4809, N4795);
buf BUF1 (N4810, N4799);
buf BUF1 (N4811, N4803);
or OR4 (N4812, N4800, N4236, N444, N3368);
xor XOR2 (N4813, N4806, N4228);
nor NOR3 (N4814, N4794, N386, N3737);
not NOT1 (N4815, N4810);
nand NAND3 (N4816, N4788, N2396, N958);
buf BUF1 (N4817, N4790);
nand NAND2 (N4818, N4814, N776);
buf BUF1 (N4819, N4807);
xor XOR2 (N4820, N4811, N1451);
nor NOR2 (N4821, N4815, N1775);
and AND4 (N4822, N4809, N2240, N1262, N3644);
and AND3 (N4823, N4808, N2376, N864);
nor NOR3 (N4824, N4819, N918, N779);
nand NAND3 (N4825, N4817, N3349, N4424);
not NOT1 (N4826, N4821);
nor NOR4 (N4827, N4818, N4293, N4727, N4126);
nand NAND2 (N4828, N4816, N1662);
nand NAND3 (N4829, N4812, N1013, N3123);
xor XOR2 (N4830, N4829, N2644);
nand NAND2 (N4831, N4826, N3598);
not NOT1 (N4832, N4823);
and AND4 (N4833, N4822, N1080, N3264, N1753);
xor XOR2 (N4834, N4820, N3449);
buf BUF1 (N4835, N4827);
and AND3 (N4836, N4813, N200, N211);
buf BUF1 (N4837, N4824);
buf BUF1 (N4838, N4832);
or OR4 (N4839, N4828, N4500, N2180, N3598);
nand NAND2 (N4840, N4825, N3556);
or OR4 (N4841, N4838, N261, N1972, N1731);
nand NAND3 (N4842, N4837, N593, N1535);
or OR2 (N4843, N4834, N1358);
xor XOR2 (N4844, N4836, N622);
xor XOR2 (N4845, N4841, N666);
and AND4 (N4846, N4844, N3328, N1941, N4357);
nor NOR2 (N4847, N4835, N320);
nand NAND4 (N4848, N4843, N101, N4070, N3943);
not NOT1 (N4849, N4848);
xor XOR2 (N4850, N4831, N3407);
buf BUF1 (N4851, N4845);
xor XOR2 (N4852, N4850, N4146);
not NOT1 (N4853, N4852);
buf BUF1 (N4854, N4839);
or OR2 (N4855, N4847, N1452);
or OR3 (N4856, N4854, N1749, N1543);
nand NAND4 (N4857, N4853, N2493, N1912, N4502);
not NOT1 (N4858, N4840);
or OR4 (N4859, N4849, N4857, N1992, N3398);
nand NAND2 (N4860, N1277, N3805);
nand NAND2 (N4861, N4830, N3179);
xor XOR2 (N4862, N4856, N3675);
nor NOR4 (N4863, N4859, N2851, N1052, N2994);
and AND3 (N4864, N4855, N1660, N4637);
buf BUF1 (N4865, N4861);
xor XOR2 (N4866, N4833, N4672);
nand NAND4 (N4867, N4864, N4208, N2663, N4665);
and AND2 (N4868, N4863, N399);
not NOT1 (N4869, N4860);
and AND2 (N4870, N4866, N4708);
xor XOR2 (N4871, N4868, N831);
nor NOR3 (N4872, N4851, N4791, N2987);
nand NAND2 (N4873, N4858, N193);
xor XOR2 (N4874, N4869, N4722);
nand NAND3 (N4875, N4871, N2308, N4385);
xor XOR2 (N4876, N4842, N2067);
or OR4 (N4877, N4874, N4144, N1918, N628);
or OR3 (N4878, N4876, N657, N540);
nor NOR2 (N4879, N4878, N803);
and AND2 (N4880, N4879, N1222);
or OR2 (N4881, N4865, N204);
nor NOR4 (N4882, N4870, N2328, N4121, N3703);
or OR3 (N4883, N4877, N3720, N1);
nor NOR3 (N4884, N4867, N4636, N4855);
and AND4 (N4885, N4883, N4175, N131, N2298);
or OR3 (N4886, N4875, N3733, N1030);
or OR2 (N4887, N4882, N1152);
xor XOR2 (N4888, N4886, N2419);
or OR4 (N4889, N4873, N623, N4652, N1368);
nand NAND4 (N4890, N4889, N1280, N826, N2103);
buf BUF1 (N4891, N4890);
buf BUF1 (N4892, N4872);
or OR3 (N4893, N4888, N4695, N2676);
xor XOR2 (N4894, N4891, N397);
or OR2 (N4895, N4893, N74);
and AND2 (N4896, N4887, N2961);
nand NAND4 (N4897, N4894, N4605, N1044, N3504);
and AND2 (N4898, N4895, N3489);
and AND2 (N4899, N4897, N3803);
not NOT1 (N4900, N4899);
buf BUF1 (N4901, N4846);
xor XOR2 (N4902, N4896, N3644);
not NOT1 (N4903, N4881);
and AND3 (N4904, N4892, N4794, N3495);
xor XOR2 (N4905, N4862, N2808);
and AND2 (N4906, N4898, N1023);
xor XOR2 (N4907, N4906, N3456);
and AND4 (N4908, N4907, N1773, N2664, N4247);
or OR3 (N4909, N4908, N2557, N4654);
xor XOR2 (N4910, N4902, N3516);
and AND4 (N4911, N4904, N480, N4060, N252);
and AND3 (N4912, N4909, N178, N4411);
and AND4 (N4913, N4912, N2832, N3769, N4566);
or OR3 (N4914, N4905, N3670, N2492);
nor NOR2 (N4915, N4900, N4175);
not NOT1 (N4916, N4910);
xor XOR2 (N4917, N4915, N123);
buf BUF1 (N4918, N4914);
nor NOR4 (N4919, N4901, N2090, N2246, N1803);
nor NOR4 (N4920, N4880, N1233, N3462, N1402);
not NOT1 (N4921, N4920);
nand NAND2 (N4922, N4921, N4683);
buf BUF1 (N4923, N4884);
xor XOR2 (N4924, N4903, N3397);
nand NAND4 (N4925, N4917, N711, N1707, N461);
not NOT1 (N4926, N4918);
not NOT1 (N4927, N4916);
xor XOR2 (N4928, N4913, N1910);
not NOT1 (N4929, N4922);
not NOT1 (N4930, N4885);
nand NAND3 (N4931, N4911, N1225, N761);
buf BUF1 (N4932, N4927);
not NOT1 (N4933, N4923);
xor XOR2 (N4934, N4928, N1537);
not NOT1 (N4935, N4930);
xor XOR2 (N4936, N4919, N4241);
xor XOR2 (N4937, N4935, N2540);
not NOT1 (N4938, N4936);
buf BUF1 (N4939, N4933);
and AND4 (N4940, N4924, N4396, N114, N1242);
not NOT1 (N4941, N4931);
not NOT1 (N4942, N4932);
or OR3 (N4943, N4939, N4880, N3489);
xor XOR2 (N4944, N4937, N3041);
buf BUF1 (N4945, N4941);
or OR3 (N4946, N4944, N441, N4801);
and AND3 (N4947, N4926, N1213, N1211);
nor NOR3 (N4948, N4940, N835, N4428);
buf BUF1 (N4949, N4942);
nand NAND2 (N4950, N4925, N71);
buf BUF1 (N4951, N4943);
nor NOR2 (N4952, N4945, N2124);
and AND4 (N4953, N4949, N1013, N3380, N4629);
nor NOR3 (N4954, N4938, N139, N1384);
nor NOR3 (N4955, N4952, N2438, N512);
or OR3 (N4956, N4929, N3092, N951);
not NOT1 (N4957, N4948);
not NOT1 (N4958, N4951);
or OR4 (N4959, N4957, N2005, N4590, N4691);
nor NOR4 (N4960, N4955, N1222, N947, N2353);
nand NAND2 (N4961, N4947, N2847);
not NOT1 (N4962, N4954);
nor NOR2 (N4963, N4958, N659);
or OR2 (N4964, N4959, N3169);
nor NOR2 (N4965, N4964, N4562);
nand NAND2 (N4966, N4950, N255);
nand NAND4 (N4967, N4962, N529, N1462, N2060);
xor XOR2 (N4968, N4946, N4779);
not NOT1 (N4969, N4961);
nand NAND3 (N4970, N4965, N2874, N2474);
nand NAND4 (N4971, N4953, N1603, N733, N2804);
or OR3 (N4972, N4970, N4068, N716);
and AND4 (N4973, N4967, N4667, N416, N4458);
nor NOR4 (N4974, N4973, N843, N2025, N995);
xor XOR2 (N4975, N4969, N111);
buf BUF1 (N4976, N4972);
or OR4 (N4977, N4976, N406, N2540, N1189);
buf BUF1 (N4978, N4960);
and AND2 (N4979, N4956, N1298);
nor NOR3 (N4980, N4977, N459, N4664);
xor XOR2 (N4981, N4978, N3633);
nor NOR4 (N4982, N4966, N2672, N3311, N416);
xor XOR2 (N4983, N4963, N3113);
buf BUF1 (N4984, N4981);
xor XOR2 (N4985, N4968, N3289);
xor XOR2 (N4986, N4975, N1996);
xor XOR2 (N4987, N4986, N810);
nor NOR3 (N4988, N4934, N2128, N4352);
buf BUF1 (N4989, N4979);
or OR2 (N4990, N4985, N1366);
nor NOR3 (N4991, N4984, N3340, N4283);
or OR2 (N4992, N4991, N2161);
buf BUF1 (N4993, N4982);
nor NOR2 (N4994, N4988, N4957);
xor XOR2 (N4995, N4994, N4961);
and AND2 (N4996, N4993, N2721);
not NOT1 (N4997, N4971);
buf BUF1 (N4998, N4983);
or OR4 (N4999, N4995, N4788, N2865, N801);
buf BUF1 (N5000, N4998);
or OR3 (N5001, N4990, N4745, N2599);
and AND4 (N5002, N4997, N4951, N2167, N3292);
nor NOR4 (N5003, N4987, N1907, N2923, N939);
nor NOR2 (N5004, N5000, N321);
xor XOR2 (N5005, N4992, N1071);
nand NAND2 (N5006, N5003, N1491);
nor NOR3 (N5007, N5004, N4776, N4011);
and AND4 (N5008, N5002, N2536, N3904, N4842);
and AND4 (N5009, N4974, N3147, N3361, N1529);
or OR3 (N5010, N4999, N3435, N1221);
buf BUF1 (N5011, N5001);
not NOT1 (N5012, N5009);
and AND3 (N5013, N5007, N204, N1708);
or OR3 (N5014, N5012, N2583, N2501);
or OR4 (N5015, N5010, N375, N4478, N4785);
nand NAND4 (N5016, N4996, N2054, N30, N4390);
and AND2 (N5017, N5013, N2339);
nor NOR2 (N5018, N5016, N3388);
buf BUF1 (N5019, N5018);
not NOT1 (N5020, N4980);
or OR2 (N5021, N5005, N2978);
nor NOR4 (N5022, N4989, N2879, N210, N4434);
not NOT1 (N5023, N5011);
nand NAND3 (N5024, N5014, N3861, N2813);
nand NAND4 (N5025, N5015, N842, N3537, N1002);
not NOT1 (N5026, N5008);
xor XOR2 (N5027, N5017, N1984);
not NOT1 (N5028, N5021);
xor XOR2 (N5029, N5026, N4998);
buf BUF1 (N5030, N5022);
or OR2 (N5031, N5027, N444);
xor XOR2 (N5032, N5025, N3074);
xor XOR2 (N5033, N5023, N1255);
not NOT1 (N5034, N5006);
not NOT1 (N5035, N5030);
xor XOR2 (N5036, N5034, N4629);
not NOT1 (N5037, N5028);
or OR4 (N5038, N5033, N4562, N4382, N3032);
nand NAND4 (N5039, N5038, N2229, N655, N2079);
nand NAND4 (N5040, N5036, N2117, N245, N1327);
buf BUF1 (N5041, N5019);
nand NAND3 (N5042, N5020, N4980, N3662);
not NOT1 (N5043, N5042);
buf BUF1 (N5044, N5031);
not NOT1 (N5045, N5029);
or OR3 (N5046, N5039, N963, N4101);
not NOT1 (N5047, N5032);
not NOT1 (N5048, N5041);
nor NOR3 (N5049, N5047, N1950, N4994);
xor XOR2 (N5050, N5035, N1654);
buf BUF1 (N5051, N5046);
buf BUF1 (N5052, N5024);
and AND4 (N5053, N5044, N1628, N537, N4343);
or OR3 (N5054, N5048, N1028, N1943);
not NOT1 (N5055, N5054);
or OR4 (N5056, N5052, N4371, N3243, N4498);
nand NAND2 (N5057, N5056, N3364);
and AND2 (N5058, N5040, N4106);
and AND4 (N5059, N5037, N2672, N4685, N417);
buf BUF1 (N5060, N5058);
xor XOR2 (N5061, N5045, N4661);
buf BUF1 (N5062, N5049);
nor NOR3 (N5063, N5055, N1450, N2345);
nor NOR3 (N5064, N5051, N3146, N4703);
and AND4 (N5065, N5057, N3221, N4168, N2290);
nor NOR3 (N5066, N5050, N4518, N656);
xor XOR2 (N5067, N5053, N4341);
xor XOR2 (N5068, N5066, N3914);
and AND4 (N5069, N5061, N1171, N988, N1104);
and AND3 (N5070, N5064, N3536, N689);
and AND3 (N5071, N5059, N4489, N3192);
or OR3 (N5072, N5065, N569, N3299);
or OR4 (N5073, N5069, N2760, N969, N3340);
and AND2 (N5074, N5043, N2807);
and AND3 (N5075, N5062, N1722, N2105);
and AND2 (N5076, N5075, N4420);
nor NOR2 (N5077, N5072, N3851);
or OR2 (N5078, N5074, N3814);
nand NAND2 (N5079, N5078, N947);
not NOT1 (N5080, N5060);
or OR4 (N5081, N5080, N4567, N2111, N14);
or OR3 (N5082, N5063, N3179, N4848);
nor NOR4 (N5083, N5079, N4944, N4297, N1590);
nand NAND4 (N5084, N5070, N243, N3055, N3327);
not NOT1 (N5085, N5071);
or OR2 (N5086, N5081, N4145);
buf BUF1 (N5087, N5077);
nand NAND2 (N5088, N5087, N2390);
not NOT1 (N5089, N5083);
nand NAND4 (N5090, N5088, N842, N58, N4871);
and AND4 (N5091, N5086, N1002, N3191, N1046);
nand NAND4 (N5092, N5073, N382, N2606, N1609);
nand NAND2 (N5093, N5092, N3858);
not NOT1 (N5094, N5090);
nand NAND2 (N5095, N5082, N2844);
buf BUF1 (N5096, N5091);
nor NOR2 (N5097, N5094, N47);
nor NOR4 (N5098, N5068, N4964, N704, N3426);
not NOT1 (N5099, N5089);
xor XOR2 (N5100, N5084, N4834);
xor XOR2 (N5101, N5096, N2717);
not NOT1 (N5102, N5101);
not NOT1 (N5103, N5067);
buf BUF1 (N5104, N5095);
and AND3 (N5105, N5098, N1214, N640);
nand NAND2 (N5106, N5099, N2333);
nor NOR2 (N5107, N5085, N3506);
and AND2 (N5108, N5076, N1111);
xor XOR2 (N5109, N5107, N865);
buf BUF1 (N5110, N5109);
xor XOR2 (N5111, N5100, N4054);
nand NAND3 (N5112, N5102, N4643, N3537);
not NOT1 (N5113, N5108);
not NOT1 (N5114, N5093);
and AND3 (N5115, N5106, N90, N4726);
nand NAND2 (N5116, N5114, N109);
not NOT1 (N5117, N5103);
nand NAND2 (N5118, N5111, N1902);
buf BUF1 (N5119, N5116);
buf BUF1 (N5120, N5097);
buf BUF1 (N5121, N5112);
and AND2 (N5122, N5104, N4339);
and AND4 (N5123, N5121, N1449, N2775, N1396);
nor NOR4 (N5124, N5113, N5122, N444, N3338);
or OR2 (N5125, N4321, N3536);
or OR2 (N5126, N5119, N478);
nor NOR3 (N5127, N5115, N1910, N528);
nor NOR3 (N5128, N5110, N2246, N1255);
and AND4 (N5129, N5118, N506, N4893, N4392);
or OR4 (N5130, N5129, N579, N2118, N2817);
buf BUF1 (N5131, N5117);
not NOT1 (N5132, N5125);
nor NOR4 (N5133, N5131, N70, N2098, N4370);
buf BUF1 (N5134, N5120);
not NOT1 (N5135, N5124);
xor XOR2 (N5136, N5130, N1104);
nor NOR4 (N5137, N5136, N3640, N4349, N3168);
nand NAND2 (N5138, N5128, N513);
not NOT1 (N5139, N5135);
not NOT1 (N5140, N5127);
xor XOR2 (N5141, N5138, N3881);
not NOT1 (N5142, N5137);
not NOT1 (N5143, N5105);
nor NOR4 (N5144, N5139, N423, N3784, N3092);
nand NAND2 (N5145, N5134, N846);
and AND2 (N5146, N5133, N1497);
not NOT1 (N5147, N5142);
and AND3 (N5148, N5126, N3923, N621);
or OR2 (N5149, N5140, N4030);
not NOT1 (N5150, N5132);
or OR3 (N5151, N5148, N3170, N662);
not NOT1 (N5152, N5144);
nor NOR2 (N5153, N5143, N2173);
xor XOR2 (N5154, N5145, N1415);
buf BUF1 (N5155, N5141);
and AND4 (N5156, N5123, N3489, N5064, N4276);
xor XOR2 (N5157, N5154, N4419);
buf BUF1 (N5158, N5147);
not NOT1 (N5159, N5152);
xor XOR2 (N5160, N5146, N265);
or OR2 (N5161, N5150, N2009);
or OR3 (N5162, N5149, N2524, N752);
not NOT1 (N5163, N5162);
xor XOR2 (N5164, N5159, N3306);
nand NAND2 (N5165, N5164, N5058);
xor XOR2 (N5166, N5161, N3701);
or OR3 (N5167, N5160, N2492, N3428);
nor NOR3 (N5168, N5151, N2181, N4302);
or OR2 (N5169, N5157, N2929);
buf BUF1 (N5170, N5167);
and AND3 (N5171, N5168, N2768, N4880);
or OR2 (N5172, N5171, N3655);
not NOT1 (N5173, N5155);
and AND3 (N5174, N5156, N1866, N756);
xor XOR2 (N5175, N5172, N1630);
nor NOR3 (N5176, N5175, N1072, N5073);
nand NAND2 (N5177, N5173, N2213);
not NOT1 (N5178, N5163);
xor XOR2 (N5179, N5166, N336);
nand NAND2 (N5180, N5177, N807);
or OR4 (N5181, N5169, N4611, N5133, N387);
buf BUF1 (N5182, N5165);
not NOT1 (N5183, N5178);
or OR4 (N5184, N5174, N437, N4282, N3125);
and AND3 (N5185, N5183, N2592, N4530);
nor NOR2 (N5186, N5185, N1869);
and AND3 (N5187, N5176, N373, N4812);
and AND3 (N5188, N5153, N128, N3374);
or OR3 (N5189, N5188, N4272, N3332);
and AND2 (N5190, N5181, N2594);
nand NAND2 (N5191, N5180, N4510);
nand NAND3 (N5192, N5190, N142, N675);
buf BUF1 (N5193, N5192);
nand NAND3 (N5194, N5158, N4282, N3550);
xor XOR2 (N5195, N5187, N2122);
nor NOR4 (N5196, N5193, N4740, N243, N345);
nor NOR3 (N5197, N5184, N2766, N1465);
not NOT1 (N5198, N5197);
and AND3 (N5199, N5189, N5080, N4453);
not NOT1 (N5200, N5198);
and AND2 (N5201, N5170, N710);
or OR2 (N5202, N5182, N4660);
nor NOR3 (N5203, N5196, N561, N2701);
not NOT1 (N5204, N5186);
xor XOR2 (N5205, N5194, N426);
buf BUF1 (N5206, N5203);
nand NAND4 (N5207, N5201, N438, N5165, N2950);
not NOT1 (N5208, N5199);
nor NOR4 (N5209, N5191, N4457, N4003, N1954);
not NOT1 (N5210, N5179);
buf BUF1 (N5211, N5208);
nand NAND3 (N5212, N5207, N2546, N5039);
buf BUF1 (N5213, N5195);
nand NAND2 (N5214, N5213, N3332);
not NOT1 (N5215, N5205);
and AND4 (N5216, N5209, N318, N1824, N3579);
or OR3 (N5217, N5214, N4119, N1382);
and AND2 (N5218, N5212, N2731);
nor NOR2 (N5219, N5211, N3900);
nor NOR4 (N5220, N5219, N4199, N4262, N2116);
not NOT1 (N5221, N5216);
xor XOR2 (N5222, N5217, N3067);
not NOT1 (N5223, N5221);
buf BUF1 (N5224, N5204);
xor XOR2 (N5225, N5218, N2700);
or OR2 (N5226, N5222, N2169);
buf BUF1 (N5227, N5200);
nand NAND4 (N5228, N5226, N4916, N4486, N4289);
not NOT1 (N5229, N5228);
or OR2 (N5230, N5229, N3533);
or OR4 (N5231, N5206, N548, N4552, N4014);
or OR2 (N5232, N5227, N4040);
xor XOR2 (N5233, N5225, N4972);
nor NOR4 (N5234, N5223, N4291, N227, N3944);
not NOT1 (N5235, N5231);
nor NOR3 (N5236, N5232, N3579, N1005);
nand NAND4 (N5237, N5202, N1608, N816, N1640);
nand NAND4 (N5238, N5235, N405, N3643, N418);
nor NOR2 (N5239, N5233, N147);
xor XOR2 (N5240, N5237, N2984);
not NOT1 (N5241, N5236);
xor XOR2 (N5242, N5239, N1655);
nand NAND2 (N5243, N5234, N4652);
and AND2 (N5244, N5238, N766);
xor XOR2 (N5245, N5241, N296);
xor XOR2 (N5246, N5244, N4383);
or OR4 (N5247, N5240, N1165, N4274, N3106);
and AND2 (N5248, N5220, N2543);
or OR3 (N5249, N5248, N1803, N1216);
not NOT1 (N5250, N5247);
buf BUF1 (N5251, N5243);
xor XOR2 (N5252, N5250, N75);
xor XOR2 (N5253, N5230, N2818);
not NOT1 (N5254, N5249);
nand NAND2 (N5255, N5210, N5169);
not NOT1 (N5256, N5246);
and AND2 (N5257, N5256, N3947);
nand NAND4 (N5258, N5215, N1290, N1424, N1172);
not NOT1 (N5259, N5255);
nor NOR4 (N5260, N5251, N4983, N4352, N2979);
buf BUF1 (N5261, N5252);
buf BUF1 (N5262, N5254);
nor NOR3 (N5263, N5261, N4586, N1578);
or OR2 (N5264, N5258, N3860);
xor XOR2 (N5265, N5263, N1780);
or OR4 (N5266, N5253, N2981, N2387, N5102);
not NOT1 (N5267, N5245);
nand NAND4 (N5268, N5259, N2349, N4325, N2080);
and AND4 (N5269, N5267, N4357, N3664, N2995);
and AND3 (N5270, N5265, N977, N3640);
buf BUF1 (N5271, N5257);
and AND2 (N5272, N5270, N2017);
xor XOR2 (N5273, N5242, N4513);
nor NOR4 (N5274, N5224, N2214, N3148, N809);
or OR3 (N5275, N5260, N4426, N3194);
buf BUF1 (N5276, N5271);
and AND3 (N5277, N5268, N5276, N572);
xor XOR2 (N5278, N4059, N2634);
or OR4 (N5279, N5275, N3599, N2382, N537);
or OR3 (N5280, N5279, N1074, N4439);
buf BUF1 (N5281, N5274);
or OR2 (N5282, N5273, N5226);
or OR2 (N5283, N5262, N3219);
xor XOR2 (N5284, N5282, N3067);
buf BUF1 (N5285, N5278);
nand NAND3 (N5286, N5266, N4880, N5011);
not NOT1 (N5287, N5264);
buf BUF1 (N5288, N5287);
not NOT1 (N5289, N5281);
nand NAND2 (N5290, N5272, N423);
nor NOR3 (N5291, N5280, N4915, N2056);
xor XOR2 (N5292, N5269, N2481);
and AND4 (N5293, N5291, N3359, N786, N1980);
nand NAND4 (N5294, N5286, N698, N4626, N3618);
nor NOR4 (N5295, N5294, N1483, N3752, N4868);
buf BUF1 (N5296, N5288);
nand NAND2 (N5297, N5295, N1806);
nor NOR3 (N5298, N5292, N16, N3793);
not NOT1 (N5299, N5289);
and AND2 (N5300, N5290, N5042);
not NOT1 (N5301, N5285);
xor XOR2 (N5302, N5296, N719);
not NOT1 (N5303, N5293);
or OR2 (N5304, N5297, N1350);
xor XOR2 (N5305, N5298, N73);
and AND4 (N5306, N5284, N2246, N4509, N3650);
buf BUF1 (N5307, N5301);
not NOT1 (N5308, N5306);
buf BUF1 (N5309, N5299);
or OR3 (N5310, N5309, N4225, N2456);
xor XOR2 (N5311, N5303, N1738);
nor NOR2 (N5312, N5308, N1824);
xor XOR2 (N5313, N5310, N4898);
nor NOR3 (N5314, N5312, N3135, N2330);
and AND2 (N5315, N5300, N5086);
xor XOR2 (N5316, N5305, N3541);
buf BUF1 (N5317, N5302);
xor XOR2 (N5318, N5283, N437);
buf BUF1 (N5319, N5307);
and AND2 (N5320, N5313, N5024);
buf BUF1 (N5321, N5319);
and AND2 (N5322, N5277, N1785);
nor NOR2 (N5323, N5314, N395);
nor NOR4 (N5324, N5317, N471, N4195, N2968);
nand NAND3 (N5325, N5320, N2748, N4425);
xor XOR2 (N5326, N5325, N2486);
xor XOR2 (N5327, N5324, N3441);
nand NAND3 (N5328, N5318, N474, N3258);
or OR4 (N5329, N5315, N2270, N4738, N4762);
nand NAND2 (N5330, N5316, N2051);
xor XOR2 (N5331, N5330, N4773);
and AND3 (N5332, N5304, N3902, N1328);
nand NAND4 (N5333, N5332, N4223, N3037, N5019);
or OR2 (N5334, N5311, N4639);
nor NOR2 (N5335, N5323, N4560);
buf BUF1 (N5336, N5327);
and AND4 (N5337, N5328, N2368, N2305, N280);
buf BUF1 (N5338, N5335);
nor NOR3 (N5339, N5337, N351, N4654);
and AND3 (N5340, N5334, N1231, N625);
not NOT1 (N5341, N5321);
buf BUF1 (N5342, N5336);
and AND3 (N5343, N5338, N1589, N2573);
and AND3 (N5344, N5331, N4827, N1257);
xor XOR2 (N5345, N5342, N3938);
xor XOR2 (N5346, N5344, N3108);
nand NAND2 (N5347, N5341, N668);
or OR3 (N5348, N5346, N3606, N2026);
nand NAND4 (N5349, N5347, N93, N1703, N2333);
buf BUF1 (N5350, N5340);
and AND3 (N5351, N5345, N4915, N3724);
xor XOR2 (N5352, N5343, N2074);
or OR3 (N5353, N5333, N5036, N5255);
not NOT1 (N5354, N5350);
buf BUF1 (N5355, N5326);
not NOT1 (N5356, N5353);
and AND4 (N5357, N5354, N1134, N1242, N1835);
not NOT1 (N5358, N5352);
nand NAND4 (N5359, N5339, N4261, N1340, N556);
or OR4 (N5360, N5358, N1844, N2850, N5253);
buf BUF1 (N5361, N5349);
not NOT1 (N5362, N5360);
buf BUF1 (N5363, N5348);
and AND2 (N5364, N5361, N2722);
nand NAND4 (N5365, N5322, N3165, N4765, N793);
buf BUF1 (N5366, N5351);
and AND4 (N5367, N5365, N972, N1750, N2161);
not NOT1 (N5368, N5329);
or OR2 (N5369, N5368, N786);
xor XOR2 (N5370, N5369, N3255);
and AND4 (N5371, N5367, N3587, N341, N3094);
and AND3 (N5372, N5357, N3857, N2978);
xor XOR2 (N5373, N5355, N3930);
and AND2 (N5374, N5371, N5320);
nand NAND2 (N5375, N5372, N1633);
not NOT1 (N5376, N5366);
nand NAND3 (N5377, N5374, N215, N865);
and AND3 (N5378, N5356, N291, N5293);
nor NOR3 (N5379, N5378, N1532, N2395);
buf BUF1 (N5380, N5363);
nand NAND2 (N5381, N5375, N2072);
not NOT1 (N5382, N5362);
nor NOR2 (N5383, N5364, N3051);
not NOT1 (N5384, N5377);
nand NAND2 (N5385, N5376, N3092);
nor NOR2 (N5386, N5384, N4264);
xor XOR2 (N5387, N5386, N3733);
nor NOR2 (N5388, N5359, N2476);
nand NAND3 (N5389, N5388, N3148, N3903);
and AND2 (N5390, N5389, N4902);
buf BUF1 (N5391, N5380);
nand NAND2 (N5392, N5382, N2652);
buf BUF1 (N5393, N5383);
not NOT1 (N5394, N5379);
and AND3 (N5395, N5393, N4063, N1803);
xor XOR2 (N5396, N5385, N1994);
and AND2 (N5397, N5381, N4191);
xor XOR2 (N5398, N5370, N4160);
buf BUF1 (N5399, N5396);
and AND3 (N5400, N5387, N2588, N642);
nor NOR2 (N5401, N5400, N4930);
buf BUF1 (N5402, N5392);
not NOT1 (N5403, N5399);
and AND3 (N5404, N5397, N5331, N1270);
xor XOR2 (N5405, N5398, N2581);
or OR2 (N5406, N5391, N3075);
not NOT1 (N5407, N5401);
not NOT1 (N5408, N5394);
and AND2 (N5409, N5395, N4552);
not NOT1 (N5410, N5390);
xor XOR2 (N5411, N5408, N2563);
and AND2 (N5412, N5406, N2765);
and AND3 (N5413, N5407, N2340, N1985);
xor XOR2 (N5414, N5412, N3768);
not NOT1 (N5415, N5402);
buf BUF1 (N5416, N5415);
and AND2 (N5417, N5403, N3670);
and AND2 (N5418, N5405, N1059);
nor NOR3 (N5419, N5418, N2800, N4524);
buf BUF1 (N5420, N5373);
buf BUF1 (N5421, N5416);
nor NOR4 (N5422, N5417, N2258, N3312, N529);
xor XOR2 (N5423, N5409, N2423);
xor XOR2 (N5424, N5413, N3961);
xor XOR2 (N5425, N5424, N3884);
or OR2 (N5426, N5419, N346);
nand NAND3 (N5427, N5404, N3159, N2332);
buf BUF1 (N5428, N5421);
nand NAND4 (N5429, N5411, N5010, N4712, N2057);
or OR3 (N5430, N5423, N3850, N2933);
not NOT1 (N5431, N5425);
not NOT1 (N5432, N5426);
nand NAND2 (N5433, N5420, N3136);
not NOT1 (N5434, N5433);
not NOT1 (N5435, N5410);
xor XOR2 (N5436, N5430, N982);
nor NOR2 (N5437, N5435, N4721);
buf BUF1 (N5438, N5431);
buf BUF1 (N5439, N5432);
nand NAND4 (N5440, N5428, N2040, N586, N4762);
buf BUF1 (N5441, N5427);
not NOT1 (N5442, N5440);
buf BUF1 (N5443, N5442);
not NOT1 (N5444, N5441);
nand NAND4 (N5445, N5434, N5422, N5138, N2052);
nand NAND3 (N5446, N2633, N84, N2806);
not NOT1 (N5447, N5438);
xor XOR2 (N5448, N5439, N4752);
buf BUF1 (N5449, N5414);
xor XOR2 (N5450, N5436, N466);
nand NAND3 (N5451, N5449, N2177, N5286);
nor NOR4 (N5452, N5448, N4870, N334, N3460);
or OR4 (N5453, N5451, N4981, N853, N5206);
nand NAND2 (N5454, N5447, N607);
buf BUF1 (N5455, N5454);
or OR3 (N5456, N5429, N2054, N695);
nor NOR4 (N5457, N5444, N5432, N3009, N3866);
or OR2 (N5458, N5452, N5096);
nor NOR3 (N5459, N5450, N1973, N3066);
buf BUF1 (N5460, N5445);
nand NAND3 (N5461, N5446, N5404, N4688);
nor NOR3 (N5462, N5458, N1282, N3943);
xor XOR2 (N5463, N5456, N5178);
nor NOR2 (N5464, N5455, N2494);
or OR2 (N5465, N5462, N3207);
nand NAND3 (N5466, N5465, N4109, N2130);
nor NOR3 (N5467, N5463, N5207, N931);
buf BUF1 (N5468, N5461);
or OR4 (N5469, N5464, N950, N1580, N1974);
and AND2 (N5470, N5443, N1818);
nand NAND2 (N5471, N5459, N1779);
and AND3 (N5472, N5437, N246, N3868);
xor XOR2 (N5473, N5472, N4404);
nor NOR4 (N5474, N5473, N531, N2064, N4040);
or OR4 (N5475, N5460, N227, N2485, N36);
and AND3 (N5476, N5457, N4238, N3056);
or OR2 (N5477, N5470, N2119);
buf BUF1 (N5478, N5453);
or OR3 (N5479, N5466, N2200, N3385);
nor NOR4 (N5480, N5469, N3244, N3061, N3345);
nand NAND2 (N5481, N5480, N2362);
nor NOR4 (N5482, N5479, N3573, N2663, N4934);
buf BUF1 (N5483, N5474);
nor NOR3 (N5484, N5478, N1141, N4618);
not NOT1 (N5485, N5481);
and AND4 (N5486, N5471, N5337, N1629, N842);
and AND4 (N5487, N5468, N3849, N2676, N652);
or OR2 (N5488, N5483, N5066);
nor NOR3 (N5489, N5488, N1105, N5285);
nor NOR4 (N5490, N5475, N3582, N687, N4146);
buf BUF1 (N5491, N5467);
and AND3 (N5492, N5487, N1556, N1968);
xor XOR2 (N5493, N5485, N1711);
nor NOR3 (N5494, N5476, N4770, N1233);
or OR4 (N5495, N5491, N4201, N4184, N3837);
not NOT1 (N5496, N5489);
or OR2 (N5497, N5484, N2883);
nand NAND3 (N5498, N5493, N4170, N3431);
or OR3 (N5499, N5496, N381, N1865);
xor XOR2 (N5500, N5490, N126);
or OR2 (N5501, N5494, N2631);
nor NOR4 (N5502, N5492, N3020, N746, N136);
nor NOR2 (N5503, N5500, N4406);
and AND4 (N5504, N5482, N490, N5143, N3474);
xor XOR2 (N5505, N5502, N4505);
and AND2 (N5506, N5505, N5083);
nand NAND2 (N5507, N5501, N4932);
or OR4 (N5508, N5507, N2383, N1838, N912);
xor XOR2 (N5509, N5499, N3822);
or OR2 (N5510, N5509, N1637);
or OR3 (N5511, N5504, N968, N583);
and AND4 (N5512, N5511, N2751, N4178, N2516);
xor XOR2 (N5513, N5503, N978);
nor NOR2 (N5514, N5495, N3743);
not NOT1 (N5515, N5477);
not NOT1 (N5516, N5506);
and AND3 (N5517, N5498, N3126, N755);
xor XOR2 (N5518, N5510, N3931);
not NOT1 (N5519, N5514);
nor NOR3 (N5520, N5512, N4191, N3050);
or OR4 (N5521, N5497, N1013, N3842, N995);
nor NOR4 (N5522, N5519, N4089, N745, N2782);
or OR2 (N5523, N5508, N1287);
nand NAND2 (N5524, N5516, N3686);
nand NAND3 (N5525, N5517, N128, N929);
xor XOR2 (N5526, N5513, N3599);
nor NOR2 (N5527, N5486, N4679);
nor NOR3 (N5528, N5515, N3598, N1619);
and AND3 (N5529, N5524, N794, N481);
buf BUF1 (N5530, N5529);
xor XOR2 (N5531, N5518, N1696);
nor NOR2 (N5532, N5527, N110);
nor NOR2 (N5533, N5532, N4369);
xor XOR2 (N5534, N5533, N3800);
nand NAND3 (N5535, N5530, N136, N4281);
nor NOR3 (N5536, N5526, N1337, N2771);
xor XOR2 (N5537, N5531, N490);
buf BUF1 (N5538, N5520);
xor XOR2 (N5539, N5523, N937);
not NOT1 (N5540, N5521);
and AND4 (N5541, N5522, N4668, N3356, N1953);
buf BUF1 (N5542, N5534);
and AND3 (N5543, N5540, N1314, N27);
not NOT1 (N5544, N5542);
and AND3 (N5545, N5525, N4010, N3330);
buf BUF1 (N5546, N5528);
and AND2 (N5547, N5544, N4192);
or OR3 (N5548, N5537, N4682, N1990);
nor NOR2 (N5549, N5548, N4829);
nand NAND3 (N5550, N5543, N3806, N2894);
nand NAND2 (N5551, N5547, N4129);
or OR2 (N5552, N5539, N4090);
or OR4 (N5553, N5546, N3031, N2347, N3759);
not NOT1 (N5554, N5551);
nand NAND3 (N5555, N5541, N660, N1331);
or OR3 (N5556, N5553, N2989, N4179);
or OR4 (N5557, N5549, N2519, N5224, N5015);
not NOT1 (N5558, N5550);
nand NAND2 (N5559, N5552, N329);
xor XOR2 (N5560, N5558, N1387);
nand NAND3 (N5561, N5557, N2801, N5483);
xor XOR2 (N5562, N5561, N1930);
and AND2 (N5563, N5538, N3558);
nand NAND2 (N5564, N5555, N1992);
buf BUF1 (N5565, N5535);
buf BUF1 (N5566, N5536);
nor NOR4 (N5567, N5565, N3478, N5166, N5337);
and AND4 (N5568, N5566, N452, N3088, N5039);
not NOT1 (N5569, N5556);
buf BUF1 (N5570, N5554);
or OR2 (N5571, N5563, N3305);
xor XOR2 (N5572, N5568, N34);
nand NAND2 (N5573, N5567, N4054);
or OR2 (N5574, N5562, N881);
or OR2 (N5575, N5570, N2833);
or OR4 (N5576, N5560, N988, N1318, N3325);
not NOT1 (N5577, N5569);
or OR2 (N5578, N5574, N4836);
buf BUF1 (N5579, N5545);
or OR2 (N5580, N5575, N3351);
nand NAND3 (N5581, N5564, N4844, N4991);
nand NAND4 (N5582, N5578, N122, N2234, N5080);
not NOT1 (N5583, N5576);
xor XOR2 (N5584, N5571, N3514);
not NOT1 (N5585, N5579);
xor XOR2 (N5586, N5572, N294);
nand NAND2 (N5587, N5586, N1883);
nor NOR2 (N5588, N5587, N319);
xor XOR2 (N5589, N5580, N1583);
and AND3 (N5590, N5585, N3422, N1818);
nand NAND3 (N5591, N5590, N3610, N1387);
xor XOR2 (N5592, N5581, N1210);
xor XOR2 (N5593, N5573, N1771);
or OR2 (N5594, N5589, N1024);
not NOT1 (N5595, N5593);
and AND2 (N5596, N5584, N2787);
and AND3 (N5597, N5594, N5398, N4930);
not NOT1 (N5598, N5595);
and AND3 (N5599, N5577, N2116, N684);
nand NAND3 (N5600, N5599, N1162, N2381);
xor XOR2 (N5601, N5596, N1199);
and AND3 (N5602, N5598, N2336, N5457);
xor XOR2 (N5603, N5601, N1076);
nor NOR3 (N5604, N5582, N2233, N2608);
and AND3 (N5605, N5591, N310, N1707);
xor XOR2 (N5606, N5603, N4921);
buf BUF1 (N5607, N5600);
nor NOR2 (N5608, N5583, N2458);
buf BUF1 (N5609, N5604);
not NOT1 (N5610, N5559);
xor XOR2 (N5611, N5609, N1098);
nor NOR3 (N5612, N5597, N719, N4010);
nor NOR3 (N5613, N5605, N1672, N2376);
xor XOR2 (N5614, N5613, N163);
nand NAND4 (N5615, N5602, N3112, N297, N2628);
not NOT1 (N5616, N5612);
nand NAND3 (N5617, N5610, N813, N2550);
nor NOR3 (N5618, N5614, N811, N2193);
nor NOR3 (N5619, N5616, N4826, N5369);
or OR3 (N5620, N5588, N1011, N4761);
nand NAND3 (N5621, N5608, N3100, N2991);
and AND3 (N5622, N5611, N1671, N2705);
buf BUF1 (N5623, N5617);
xor XOR2 (N5624, N5620, N1143);
nand NAND2 (N5625, N5621, N4733);
xor XOR2 (N5626, N5618, N3339);
xor XOR2 (N5627, N5592, N2950);
xor XOR2 (N5628, N5615, N187);
and AND4 (N5629, N5624, N723, N104, N2344);
not NOT1 (N5630, N5607);
nand NAND4 (N5631, N5619, N3723, N3717, N2437);
buf BUF1 (N5632, N5628);
not NOT1 (N5633, N5623);
nand NAND4 (N5634, N5630, N142, N3685, N2131);
buf BUF1 (N5635, N5632);
or OR2 (N5636, N5631, N5360);
nor NOR2 (N5637, N5625, N4325);
or OR4 (N5638, N5622, N5620, N1101, N3661);
nor NOR2 (N5639, N5638, N4019);
or OR4 (N5640, N5626, N796, N1105, N4671);
nand NAND2 (N5641, N5629, N2952);
nor NOR2 (N5642, N5627, N3959);
or OR2 (N5643, N5640, N144);
nand NAND4 (N5644, N5633, N1184, N2779, N2033);
buf BUF1 (N5645, N5643);
or OR4 (N5646, N5606, N2009, N4673, N5458);
buf BUF1 (N5647, N5641);
buf BUF1 (N5648, N5634);
nor NOR4 (N5649, N5644, N4149, N1432, N788);
not NOT1 (N5650, N5639);
nor NOR3 (N5651, N5635, N5324, N4764);
nand NAND4 (N5652, N5646, N4732, N81, N1699);
nor NOR4 (N5653, N5637, N5115, N996, N1812);
nor NOR2 (N5654, N5651, N4563);
or OR3 (N5655, N5649, N4782, N5341);
and AND4 (N5656, N5653, N502, N4061, N31);
or OR2 (N5657, N5636, N1943);
nand NAND4 (N5658, N5656, N1837, N1183, N1744);
not NOT1 (N5659, N5647);
buf BUF1 (N5660, N5657);
buf BUF1 (N5661, N5652);
nor NOR3 (N5662, N5659, N2611, N4304);
not NOT1 (N5663, N5658);
buf BUF1 (N5664, N5642);
buf BUF1 (N5665, N5660);
nand NAND4 (N5666, N5663, N4308, N1767, N5626);
not NOT1 (N5667, N5655);
or OR3 (N5668, N5664, N2180, N1791);
or OR3 (N5669, N5665, N3384, N131);
nand NAND3 (N5670, N5661, N1845, N3869);
xor XOR2 (N5671, N5650, N3078);
and AND4 (N5672, N5645, N4689, N5290, N4050);
xor XOR2 (N5673, N5666, N4243);
or OR3 (N5674, N5669, N4629, N3246);
nor NOR3 (N5675, N5672, N3042, N3521);
xor XOR2 (N5676, N5667, N2326);
xor XOR2 (N5677, N5675, N1034);
nand NAND3 (N5678, N5668, N2579, N1641);
buf BUF1 (N5679, N5673);
or OR4 (N5680, N5648, N591, N1038, N2269);
or OR2 (N5681, N5680, N2426);
nor NOR3 (N5682, N5677, N5620, N3656);
buf BUF1 (N5683, N5662);
xor XOR2 (N5684, N5683, N3145);
nand NAND4 (N5685, N5674, N904, N4773, N933);
xor XOR2 (N5686, N5678, N1187);
or OR2 (N5687, N5686, N4023);
buf BUF1 (N5688, N5681);
or OR3 (N5689, N5685, N3865, N1964);
nand NAND3 (N5690, N5676, N4962, N1346);
buf BUF1 (N5691, N5689);
xor XOR2 (N5692, N5688, N1577);
not NOT1 (N5693, N5679);
and AND3 (N5694, N5692, N2647, N5238);
and AND4 (N5695, N5691, N3033, N3011, N5442);
not NOT1 (N5696, N5682);
not NOT1 (N5697, N5694);
not NOT1 (N5698, N5696);
not NOT1 (N5699, N5687);
buf BUF1 (N5700, N5690);
xor XOR2 (N5701, N5698, N3272);
and AND2 (N5702, N5693, N532);
nand NAND4 (N5703, N5695, N1312, N5272, N4118);
nand NAND3 (N5704, N5670, N4062, N4523);
buf BUF1 (N5705, N5704);
and AND2 (N5706, N5701, N4458);
and AND4 (N5707, N5703, N4943, N1646, N96);
xor XOR2 (N5708, N5697, N768);
nand NAND3 (N5709, N5707, N3992, N3735);
nand NAND3 (N5710, N5700, N2786, N3694);
xor XOR2 (N5711, N5654, N1304);
nor NOR2 (N5712, N5706, N3507);
or OR4 (N5713, N5702, N4990, N3255, N5609);
not NOT1 (N5714, N5712);
xor XOR2 (N5715, N5684, N4614);
buf BUF1 (N5716, N5699);
buf BUF1 (N5717, N5705);
buf BUF1 (N5718, N5717);
xor XOR2 (N5719, N5715, N472);
nand NAND4 (N5720, N5671, N3976, N4478, N4385);
buf BUF1 (N5721, N5711);
or OR3 (N5722, N5719, N926, N581);
nor NOR2 (N5723, N5722, N5620);
nand NAND3 (N5724, N5714, N2352, N1804);
buf BUF1 (N5725, N5723);
xor XOR2 (N5726, N5710, N1181);
nand NAND3 (N5727, N5708, N2992, N4162);
nor NOR2 (N5728, N5716, N2572);
buf BUF1 (N5729, N5721);
nor NOR2 (N5730, N5729, N1931);
or OR4 (N5731, N5713, N276, N2822, N2349);
xor XOR2 (N5732, N5720, N5329);
nor NOR2 (N5733, N5730, N167);
nor NOR2 (N5734, N5718, N5647);
or OR4 (N5735, N5731, N2574, N1585, N5516);
buf BUF1 (N5736, N5728);
or OR4 (N5737, N5724, N4719, N4926, N2667);
nand NAND4 (N5738, N5725, N1302, N869, N812);
or OR3 (N5739, N5736, N4310, N1246);
and AND4 (N5740, N5727, N2941, N4983, N705);
not NOT1 (N5741, N5735);
nor NOR2 (N5742, N5738, N2327);
not NOT1 (N5743, N5740);
xor XOR2 (N5744, N5741, N3651);
not NOT1 (N5745, N5734);
buf BUF1 (N5746, N5709);
not NOT1 (N5747, N5733);
nor NOR2 (N5748, N5726, N3151);
nand NAND4 (N5749, N5745, N3001, N1303, N1972);
and AND3 (N5750, N5744, N3409, N937);
nor NOR3 (N5751, N5732, N3326, N5037);
xor XOR2 (N5752, N5742, N573);
buf BUF1 (N5753, N5737);
xor XOR2 (N5754, N5739, N3044);
buf BUF1 (N5755, N5754);
or OR3 (N5756, N5752, N4436, N4454);
buf BUF1 (N5757, N5743);
nand NAND4 (N5758, N5753, N5556, N1436, N2319);
buf BUF1 (N5759, N5751);
or OR3 (N5760, N5748, N693, N118);
or OR4 (N5761, N5747, N3809, N607, N2816);
nor NOR2 (N5762, N5749, N1510);
buf BUF1 (N5763, N5757);
or OR4 (N5764, N5758, N5595, N2105, N5065);
and AND2 (N5765, N5759, N1242);
not NOT1 (N5766, N5755);
nor NOR3 (N5767, N5756, N4359, N429);
nor NOR4 (N5768, N5746, N5600, N625, N2153);
buf BUF1 (N5769, N5762);
or OR2 (N5770, N5769, N1315);
or OR3 (N5771, N5768, N642, N5490);
nand NAND3 (N5772, N5764, N707, N632);
or OR4 (N5773, N5760, N3066, N5691, N2062);
and AND3 (N5774, N5765, N2195, N342);
xor XOR2 (N5775, N5766, N4570);
nand NAND2 (N5776, N5772, N1322);
and AND4 (N5777, N5761, N2950, N5560, N1104);
not NOT1 (N5778, N5776);
or OR4 (N5779, N5778, N726, N4332, N3318);
and AND4 (N5780, N5779, N3606, N3669, N5506);
nand NAND2 (N5781, N5770, N4891);
or OR3 (N5782, N5780, N5163, N2731);
nand NAND4 (N5783, N5774, N3789, N3892, N107);
or OR2 (N5784, N5763, N1068);
buf BUF1 (N5785, N5777);
nand NAND4 (N5786, N5775, N2308, N1222, N3221);
xor XOR2 (N5787, N5783, N2515);
or OR2 (N5788, N5781, N5136);
buf BUF1 (N5789, N5786);
buf BUF1 (N5790, N5787);
nor NOR3 (N5791, N5788, N4955, N4785);
xor XOR2 (N5792, N5784, N2903);
nand NAND3 (N5793, N5785, N1808, N420);
buf BUF1 (N5794, N5782);
not NOT1 (N5795, N5793);
xor XOR2 (N5796, N5795, N4511);
xor XOR2 (N5797, N5773, N1902);
and AND4 (N5798, N5750, N2062, N4998, N4340);
buf BUF1 (N5799, N5797);
nor NOR2 (N5800, N5798, N5053);
nor NOR4 (N5801, N5799, N889, N3209, N891);
or OR2 (N5802, N5789, N3061);
not NOT1 (N5803, N5790);
or OR2 (N5804, N5800, N1412);
xor XOR2 (N5805, N5804, N5302);
not NOT1 (N5806, N5792);
not NOT1 (N5807, N5806);
nand NAND3 (N5808, N5771, N1106, N4785);
nor NOR4 (N5809, N5808, N4312, N1176, N564);
or OR4 (N5810, N5801, N4608, N4266, N34);
not NOT1 (N5811, N5802);
and AND2 (N5812, N5810, N2284);
xor XOR2 (N5813, N5794, N4943);
nand NAND4 (N5814, N5767, N4174, N413, N3522);
or OR2 (N5815, N5811, N3540);
xor XOR2 (N5816, N5803, N5118);
not NOT1 (N5817, N5815);
nand NAND2 (N5818, N5809, N3924);
buf BUF1 (N5819, N5805);
not NOT1 (N5820, N5818);
xor XOR2 (N5821, N5791, N2630);
and AND3 (N5822, N5817, N2909, N424);
not NOT1 (N5823, N5814);
nand NAND4 (N5824, N5821, N4171, N4522, N4725);
and AND2 (N5825, N5822, N1155);
not NOT1 (N5826, N5819);
buf BUF1 (N5827, N5824);
or OR3 (N5828, N5827, N5494, N5127);
and AND2 (N5829, N5825, N2416);
buf BUF1 (N5830, N5828);
and AND2 (N5831, N5829, N785);
xor XOR2 (N5832, N5820, N2032);
nand NAND4 (N5833, N5796, N5002, N4473, N1429);
xor XOR2 (N5834, N5826, N705);
or OR2 (N5835, N5812, N4889);
not NOT1 (N5836, N5816);
nand NAND4 (N5837, N5807, N2848, N641, N4433);
buf BUF1 (N5838, N5833);
or OR4 (N5839, N5835, N5256, N4785, N1803);
buf BUF1 (N5840, N5832);
nor NOR2 (N5841, N5836, N4681);
xor XOR2 (N5842, N5839, N2012);
and AND2 (N5843, N5837, N2923);
or OR2 (N5844, N5841, N3315);
buf BUF1 (N5845, N5842);
nand NAND3 (N5846, N5831, N3791, N3296);
xor XOR2 (N5847, N5844, N426);
buf BUF1 (N5848, N5840);
nor NOR3 (N5849, N5843, N5495, N610);
nand NAND3 (N5850, N5849, N1583, N3300);
or OR2 (N5851, N5850, N5409);
nand NAND3 (N5852, N5851, N1059, N2704);
not NOT1 (N5853, N5823);
nand NAND3 (N5854, N5848, N1184, N3291);
xor XOR2 (N5855, N5845, N4372);
or OR3 (N5856, N5838, N106, N2042);
or OR2 (N5857, N5813, N2583);
not NOT1 (N5858, N5830);
nor NOR4 (N5859, N5855, N1144, N454, N3126);
nand NAND3 (N5860, N5856, N1036, N486);
and AND2 (N5861, N5857, N647);
nor NOR4 (N5862, N5858, N3576, N2824, N196);
not NOT1 (N5863, N5861);
xor XOR2 (N5864, N5862, N5487);
not NOT1 (N5865, N5853);
xor XOR2 (N5866, N5847, N1773);
nor NOR3 (N5867, N5863, N4494, N969);
buf BUF1 (N5868, N5854);
buf BUF1 (N5869, N5864);
not NOT1 (N5870, N5859);
nor NOR4 (N5871, N5869, N2249, N1673, N2431);
buf BUF1 (N5872, N5868);
buf BUF1 (N5873, N5865);
nor NOR2 (N5874, N5846, N2402);
nor NOR3 (N5875, N5871, N3498, N2127);
and AND2 (N5876, N5874, N4481);
and AND2 (N5877, N5866, N3861);
or OR2 (N5878, N5852, N3058);
not NOT1 (N5879, N5870);
nor NOR3 (N5880, N5877, N5262, N3468);
or OR2 (N5881, N5879, N4061);
xor XOR2 (N5882, N5876, N4673);
xor XOR2 (N5883, N5860, N4108);
and AND2 (N5884, N5834, N4604);
buf BUF1 (N5885, N5872);
xor XOR2 (N5886, N5875, N4450);
or OR3 (N5887, N5867, N1496, N3091);
nand NAND3 (N5888, N5882, N1054, N5525);
nand NAND3 (N5889, N5878, N2644, N1196);
or OR3 (N5890, N5889, N3002, N1702);
or OR3 (N5891, N5885, N3147, N5877);
nand NAND3 (N5892, N5883, N3783, N102);
and AND3 (N5893, N5881, N1826, N3112);
nor NOR4 (N5894, N5891, N698, N5862, N5871);
buf BUF1 (N5895, N5884);
and AND4 (N5896, N5893, N3293, N247, N4750);
or OR2 (N5897, N5888, N3435);
buf BUF1 (N5898, N5880);
not NOT1 (N5899, N5886);
not NOT1 (N5900, N5898);
not NOT1 (N5901, N5887);
and AND3 (N5902, N5895, N2249, N4240);
nand NAND4 (N5903, N5899, N2004, N3036, N4719);
nand NAND2 (N5904, N5900, N4649);
nand NAND3 (N5905, N5873, N658, N314);
buf BUF1 (N5906, N5905);
nor NOR4 (N5907, N5906, N3409, N2110, N2559);
buf BUF1 (N5908, N5904);
or OR3 (N5909, N5894, N4117, N1226);
or OR4 (N5910, N5902, N3740, N2452, N267);
not NOT1 (N5911, N5909);
buf BUF1 (N5912, N5890);
nor NOR3 (N5913, N5910, N1964, N4063);
xor XOR2 (N5914, N5908, N4069);
or OR2 (N5915, N5901, N5572);
and AND4 (N5916, N5914, N864, N121, N5859);
buf BUF1 (N5917, N5896);
or OR4 (N5918, N5913, N1534, N2077, N117);
nand NAND3 (N5919, N5907, N4707, N3116);
not NOT1 (N5920, N5897);
xor XOR2 (N5921, N5917, N2814);
nor NOR3 (N5922, N5915, N5351, N5287);
xor XOR2 (N5923, N5911, N3471);
or OR3 (N5924, N5916, N4366, N5545);
nor NOR2 (N5925, N5921, N2461);
not NOT1 (N5926, N5912);
buf BUF1 (N5927, N5923);
not NOT1 (N5928, N5903);
nor NOR2 (N5929, N5927, N2181);
buf BUF1 (N5930, N5892);
buf BUF1 (N5931, N5928);
or OR3 (N5932, N5929, N1530, N4481);
nor NOR2 (N5933, N5919, N3133);
or OR2 (N5934, N5933, N4147);
and AND3 (N5935, N5926, N1038, N718);
and AND3 (N5936, N5922, N3824, N4359);
not NOT1 (N5937, N5925);
not NOT1 (N5938, N5936);
not NOT1 (N5939, N5931);
not NOT1 (N5940, N5934);
or OR2 (N5941, N5940, N2196);
or OR4 (N5942, N5924, N244, N4620, N3070);
nand NAND3 (N5943, N5930, N2348, N1455);
buf BUF1 (N5944, N5937);
buf BUF1 (N5945, N5944);
and AND3 (N5946, N5918, N56, N1601);
nor NOR4 (N5947, N5942, N4774, N2295, N1615);
nand NAND4 (N5948, N5938, N4511, N4129, N1377);
or OR2 (N5949, N5943, N5224);
xor XOR2 (N5950, N5932, N3692);
not NOT1 (N5951, N5948);
or OR4 (N5952, N5951, N5798, N369, N4854);
buf BUF1 (N5953, N5945);
not NOT1 (N5954, N5920);
not NOT1 (N5955, N5939);
nand NAND3 (N5956, N5947, N3870, N1307);
and AND4 (N5957, N5953, N802, N1366, N1582);
nand NAND4 (N5958, N5941, N685, N602, N5240);
or OR3 (N5959, N5958, N762, N3877);
buf BUF1 (N5960, N5957);
buf BUF1 (N5961, N5950);
not NOT1 (N5962, N5946);
nand NAND2 (N5963, N5961, N36);
xor XOR2 (N5964, N5956, N2186);
not NOT1 (N5965, N5959);
or OR2 (N5966, N5965, N27);
and AND4 (N5967, N5966, N5129, N2662, N5061);
xor XOR2 (N5968, N5967, N3948);
xor XOR2 (N5969, N5963, N1609);
not NOT1 (N5970, N5968);
nor NOR2 (N5971, N5960, N5612);
xor XOR2 (N5972, N5954, N981);
and AND2 (N5973, N5952, N4836);
buf BUF1 (N5974, N5962);
buf BUF1 (N5975, N5964);
nand NAND3 (N5976, N5955, N2521, N1935);
nand NAND2 (N5977, N5974, N4980);
buf BUF1 (N5978, N5949);
or OR3 (N5979, N5973, N4983, N5240);
buf BUF1 (N5980, N5935);
xor XOR2 (N5981, N5970, N5691);
nor NOR2 (N5982, N5979, N3557);
nand NAND2 (N5983, N5978, N3173);
not NOT1 (N5984, N5975);
nor NOR3 (N5985, N5982, N5243, N4814);
buf BUF1 (N5986, N5983);
not NOT1 (N5987, N5986);
nand NAND4 (N5988, N5984, N3164, N1985, N1426);
xor XOR2 (N5989, N5981, N3988);
nor NOR2 (N5990, N5972, N335);
not NOT1 (N5991, N5977);
xor XOR2 (N5992, N5971, N2247);
and AND3 (N5993, N5991, N5926, N4075);
nor NOR4 (N5994, N5985, N467, N4879, N5663);
buf BUF1 (N5995, N5987);
nand NAND2 (N5996, N5976, N1832);
buf BUF1 (N5997, N5996);
or OR4 (N5998, N5980, N687, N4044, N282);
xor XOR2 (N5999, N5993, N1825);
nor NOR4 (N6000, N5998, N5953, N65, N558);
buf BUF1 (N6001, N5994);
not NOT1 (N6002, N5992);
or OR2 (N6003, N5997, N5317);
xor XOR2 (N6004, N5989, N3768);
xor XOR2 (N6005, N6001, N2852);
nor NOR3 (N6006, N6004, N969, N1102);
not NOT1 (N6007, N6006);
buf BUF1 (N6008, N6002);
buf BUF1 (N6009, N5999);
and AND4 (N6010, N6008, N3536, N4314, N3661);
nand NAND2 (N6011, N5990, N2199);
nand NAND2 (N6012, N6007, N4);
xor XOR2 (N6013, N5995, N4646);
xor XOR2 (N6014, N5988, N3489);
not NOT1 (N6015, N6003);
nand NAND2 (N6016, N6011, N2261);
xor XOR2 (N6017, N6012, N5925);
not NOT1 (N6018, N6009);
buf BUF1 (N6019, N6005);
nand NAND2 (N6020, N6014, N2863);
xor XOR2 (N6021, N6019, N2343);
nor NOR3 (N6022, N6015, N3927, N238);
and AND3 (N6023, N6016, N5396, N2614);
and AND4 (N6024, N6010, N5942, N1600, N5195);
nor NOR2 (N6025, N6013, N2054);
buf BUF1 (N6026, N6017);
or OR2 (N6027, N6018, N1681);
or OR2 (N6028, N6022, N3031);
or OR4 (N6029, N6026, N246, N2949, N1379);
or OR4 (N6030, N6021, N2854, N5324, N4091);
nand NAND3 (N6031, N6029, N4933, N4756);
or OR4 (N6032, N6025, N5803, N1400, N1873);
xor XOR2 (N6033, N6000, N3791);
and AND3 (N6034, N6023, N1659, N4715);
not NOT1 (N6035, N6030);
xor XOR2 (N6036, N6027, N1931);
and AND4 (N6037, N5969, N953, N99, N1269);
nand NAND3 (N6038, N6020, N231, N413);
buf BUF1 (N6039, N6036);
nor NOR3 (N6040, N6038, N1069, N474);
or OR3 (N6041, N6031, N2975, N5511);
not NOT1 (N6042, N6033);
or OR4 (N6043, N6028, N806, N4954, N1617);
and AND4 (N6044, N6034, N5335, N703, N449);
xor XOR2 (N6045, N6044, N511);
nor NOR2 (N6046, N6042, N1477);
xor XOR2 (N6047, N6046, N1655);
nor NOR4 (N6048, N6039, N5521, N627, N3569);
and AND4 (N6049, N6024, N4753, N468, N3770);
buf BUF1 (N6050, N6048);
and AND3 (N6051, N6032, N1797, N2144);
and AND4 (N6052, N6043, N3462, N1571, N3304);
or OR4 (N6053, N6051, N1895, N4224, N2989);
xor XOR2 (N6054, N6037, N4420);
nand NAND4 (N6055, N6040, N877, N3777, N3404);
and AND3 (N6056, N6041, N5154, N1967);
xor XOR2 (N6057, N6054, N5883);
nor NOR3 (N6058, N6055, N2076, N4606);
buf BUF1 (N6059, N6058);
or OR3 (N6060, N6047, N4518, N1132);
nor NOR3 (N6061, N6052, N2950, N4281);
not NOT1 (N6062, N6045);
and AND3 (N6063, N6049, N819, N2616);
nand NAND4 (N6064, N6060, N3294, N1817, N4699);
not NOT1 (N6065, N6064);
or OR3 (N6066, N6059, N1078, N5783);
nor NOR3 (N6067, N6053, N4814, N980);
nor NOR3 (N6068, N6056, N1200, N2029);
nor NOR3 (N6069, N6068, N3952, N2864);
or OR3 (N6070, N6061, N379, N5388);
xor XOR2 (N6071, N6065, N63);
xor XOR2 (N6072, N6066, N4996);
not NOT1 (N6073, N6070);
nor NOR2 (N6074, N6035, N4399);
or OR4 (N6075, N6069, N3383, N3741, N5524);
xor XOR2 (N6076, N6057, N1780);
nor NOR3 (N6077, N6072, N5445, N4526);
or OR3 (N6078, N6073, N4864, N1469);
not NOT1 (N6079, N6062);
buf BUF1 (N6080, N6079);
nand NAND3 (N6081, N6067, N4883, N337);
buf BUF1 (N6082, N6063);
not NOT1 (N6083, N6071);
nor NOR4 (N6084, N6075, N4365, N2830, N2629);
not NOT1 (N6085, N6080);
buf BUF1 (N6086, N6076);
nor NOR4 (N6087, N6082, N3987, N4683, N4516);
xor XOR2 (N6088, N6086, N3743);
or OR3 (N6089, N6074, N3353, N5608);
or OR2 (N6090, N6050, N2171);
or OR2 (N6091, N6090, N5530);
not NOT1 (N6092, N6088);
xor XOR2 (N6093, N6077, N857);
and AND2 (N6094, N6084, N2637);
and AND3 (N6095, N6093, N399, N229);
and AND3 (N6096, N6094, N865, N3946);
or OR3 (N6097, N6081, N3232, N3109);
buf BUF1 (N6098, N6085);
nand NAND4 (N6099, N6092, N6059, N4500, N5736);
xor XOR2 (N6100, N6096, N3521);
buf BUF1 (N6101, N6083);
nand NAND3 (N6102, N6089, N4380, N2887);
and AND3 (N6103, N6091, N4223, N1059);
and AND3 (N6104, N6099, N2303, N5245);
and AND4 (N6105, N6097, N2923, N1694, N2670);
and AND2 (N6106, N6105, N2662);
xor XOR2 (N6107, N6087, N3461);
or OR4 (N6108, N6101, N3106, N2266, N3709);
or OR3 (N6109, N6102, N2908, N128);
nand NAND3 (N6110, N6078, N4347, N3843);
buf BUF1 (N6111, N6110);
nand NAND4 (N6112, N6095, N547, N1650, N1712);
or OR2 (N6113, N6111, N4314);
buf BUF1 (N6114, N6098);
buf BUF1 (N6115, N6109);
nand NAND2 (N6116, N6112, N4613);
buf BUF1 (N6117, N6107);
nor NOR4 (N6118, N6100, N5844, N4229, N2204);
not NOT1 (N6119, N6104);
buf BUF1 (N6120, N6106);
nand NAND2 (N6121, N6120, N3797);
buf BUF1 (N6122, N6119);
and AND4 (N6123, N6108, N5930, N4752, N3615);
buf BUF1 (N6124, N6116);
buf BUF1 (N6125, N6114);
nor NOR2 (N6126, N6124, N1552);
and AND4 (N6127, N6117, N1522, N5232, N3779);
and AND3 (N6128, N6123, N2689, N3547);
nand NAND3 (N6129, N6128, N442, N3331);
nand NAND3 (N6130, N6113, N2961, N5524);
buf BUF1 (N6131, N6129);
buf BUF1 (N6132, N6121);
buf BUF1 (N6133, N6115);
not NOT1 (N6134, N6127);
buf BUF1 (N6135, N6122);
nand NAND2 (N6136, N6103, N3481);
nand NAND2 (N6137, N6133, N4834);
xor XOR2 (N6138, N6135, N2370);
buf BUF1 (N6139, N6126);
not NOT1 (N6140, N6139);
or OR3 (N6141, N6130, N2553, N2233);
or OR3 (N6142, N6140, N4083, N3441);
not NOT1 (N6143, N6134);
nor NOR4 (N6144, N6131, N579, N4119, N5944);
not NOT1 (N6145, N6141);
and AND4 (N6146, N6132, N2308, N3794, N4086);
xor XOR2 (N6147, N6136, N5855);
not NOT1 (N6148, N6143);
nand NAND3 (N6149, N6147, N2145, N5658);
nand NAND4 (N6150, N6144, N4714, N2746, N5815);
or OR3 (N6151, N6149, N748, N2649);
nor NOR3 (N6152, N6118, N333, N1537);
nand NAND2 (N6153, N6145, N56);
xor XOR2 (N6154, N6142, N5089);
buf BUF1 (N6155, N6146);
nor NOR3 (N6156, N6151, N813, N1959);
and AND2 (N6157, N6125, N2296);
nand NAND3 (N6158, N6157, N1810, N5670);
not NOT1 (N6159, N6148);
or OR2 (N6160, N6137, N2653);
not NOT1 (N6161, N6158);
not NOT1 (N6162, N6160);
buf BUF1 (N6163, N6162);
and AND2 (N6164, N6152, N1517);
buf BUF1 (N6165, N6159);
not NOT1 (N6166, N6164);
xor XOR2 (N6167, N6154, N2827);
buf BUF1 (N6168, N6153);
xor XOR2 (N6169, N6155, N4965);
or OR2 (N6170, N6165, N4147);
not NOT1 (N6171, N6163);
not NOT1 (N6172, N6169);
nor NOR3 (N6173, N6161, N676, N4822);
not NOT1 (N6174, N6150);
buf BUF1 (N6175, N6173);
and AND4 (N6176, N6138, N3076, N1877, N1936);
xor XOR2 (N6177, N6167, N6164);
xor XOR2 (N6178, N6177, N1745);
nor NOR4 (N6179, N6176, N1680, N1467, N4297);
nor NOR2 (N6180, N6174, N5361);
nor NOR2 (N6181, N6175, N4199);
buf BUF1 (N6182, N6170);
or OR2 (N6183, N6180, N1572);
xor XOR2 (N6184, N6156, N5099);
nand NAND3 (N6185, N6178, N4835, N2652);
not NOT1 (N6186, N6181);
nor NOR4 (N6187, N6171, N3254, N1570, N5091);
xor XOR2 (N6188, N6182, N3996);
nand NAND3 (N6189, N6185, N5288, N242);
and AND3 (N6190, N6187, N689, N191);
or OR3 (N6191, N6172, N978, N1504);
or OR4 (N6192, N6190, N2608, N200, N120);
and AND2 (N6193, N6179, N3014);
xor XOR2 (N6194, N6189, N2968);
xor XOR2 (N6195, N6194, N764);
buf BUF1 (N6196, N6192);
not NOT1 (N6197, N6195);
or OR2 (N6198, N6184, N2475);
nand NAND2 (N6199, N6191, N4809);
xor XOR2 (N6200, N6183, N2556);
xor XOR2 (N6201, N6197, N955);
xor XOR2 (N6202, N6196, N593);
nand NAND3 (N6203, N6166, N6162, N5168);
xor XOR2 (N6204, N6203, N1734);
nor NOR2 (N6205, N6168, N4978);
buf BUF1 (N6206, N6198);
not NOT1 (N6207, N6188);
nor NOR4 (N6208, N6206, N4093, N5416, N3844);
nand NAND4 (N6209, N6200, N383, N3739, N4138);
buf BUF1 (N6210, N6208);
nand NAND2 (N6211, N6210, N2242);
nor NOR3 (N6212, N6201, N2408, N1150);
xor XOR2 (N6213, N6209, N178);
nor NOR2 (N6214, N6205, N4416);
and AND3 (N6215, N6186, N82, N600);
nand NAND3 (N6216, N6193, N5092, N1952);
buf BUF1 (N6217, N6216);
buf BUF1 (N6218, N6204);
xor XOR2 (N6219, N6211, N4069);
nand NAND2 (N6220, N6212, N2082);
buf BUF1 (N6221, N6215);
nor NOR3 (N6222, N6220, N5817, N3311);
not NOT1 (N6223, N6222);
buf BUF1 (N6224, N6219);
xor XOR2 (N6225, N6202, N3044);
xor XOR2 (N6226, N6221, N5270);
or OR4 (N6227, N6213, N2410, N4252, N4583);
and AND3 (N6228, N6207, N142, N4737);
nor NOR4 (N6229, N6226, N3530, N2338, N3123);
nand NAND2 (N6230, N6199, N1776);
nand NAND2 (N6231, N6224, N1922);
and AND4 (N6232, N6217, N2812, N5714, N2229);
nor NOR4 (N6233, N6218, N4998, N619, N914);
nand NAND4 (N6234, N6223, N5491, N31, N2484);
nand NAND4 (N6235, N6233, N2529, N1711, N2825);
and AND2 (N6236, N6227, N1135);
and AND3 (N6237, N6225, N1386, N3704);
buf BUF1 (N6238, N6230);
xor XOR2 (N6239, N6232, N2889);
xor XOR2 (N6240, N6214, N683);
buf BUF1 (N6241, N6237);
xor XOR2 (N6242, N6241, N4629);
buf BUF1 (N6243, N6238);
nor NOR2 (N6244, N6236, N123);
xor XOR2 (N6245, N6244, N3927);
nand NAND2 (N6246, N6231, N5017);
nor NOR2 (N6247, N6228, N4679);
and AND4 (N6248, N6245, N5371, N1333, N4816);
buf BUF1 (N6249, N6234);
xor XOR2 (N6250, N6239, N4525);
nor NOR3 (N6251, N6242, N6163, N2756);
xor XOR2 (N6252, N6247, N1612);
nor NOR3 (N6253, N6248, N2722, N3753);
buf BUF1 (N6254, N6243);
not NOT1 (N6255, N6240);
not NOT1 (N6256, N6250);
not NOT1 (N6257, N6249);
not NOT1 (N6258, N6235);
buf BUF1 (N6259, N6229);
xor XOR2 (N6260, N6256, N6085);
and AND2 (N6261, N6257, N476);
nor NOR4 (N6262, N6246, N4037, N3751, N4272);
buf BUF1 (N6263, N6254);
xor XOR2 (N6264, N6261, N1462);
and AND4 (N6265, N6255, N1617, N1760, N5074);
nand NAND2 (N6266, N6260, N1913);
nor NOR3 (N6267, N6263, N4285, N5742);
buf BUF1 (N6268, N6266);
nor NOR3 (N6269, N6262, N912, N4530);
nor NOR2 (N6270, N6268, N3881);
or OR4 (N6271, N6253, N4126, N5167, N2185);
xor XOR2 (N6272, N6269, N6196);
and AND4 (N6273, N6251, N4955, N4916, N4984);
or OR3 (N6274, N6259, N5391, N3459);
nand NAND4 (N6275, N6264, N2423, N5261, N3576);
nor NOR2 (N6276, N6265, N5280);
not NOT1 (N6277, N6258);
nand NAND4 (N6278, N6275, N2816, N2287, N1541);
nand NAND4 (N6279, N6277, N5736, N2776, N1080);
buf BUF1 (N6280, N6267);
and AND2 (N6281, N6273, N5025);
buf BUF1 (N6282, N6281);
nor NOR2 (N6283, N6274, N705);
buf BUF1 (N6284, N6280);
and AND3 (N6285, N6252, N2919, N2379);
not NOT1 (N6286, N6283);
and AND3 (N6287, N6278, N469, N1015);
or OR2 (N6288, N6271, N3327);
or OR4 (N6289, N6270, N3449, N1486, N3898);
not NOT1 (N6290, N6286);
nand NAND4 (N6291, N6285, N5127, N4200, N1197);
nor NOR3 (N6292, N6290, N4163, N2855);
xor XOR2 (N6293, N6276, N4875);
and AND4 (N6294, N6282, N1567, N3322, N2161);
nand NAND2 (N6295, N6294, N3835);
and AND4 (N6296, N6293, N5425, N4168, N4584);
buf BUF1 (N6297, N6288);
not NOT1 (N6298, N6292);
and AND2 (N6299, N6289, N3332);
xor XOR2 (N6300, N6295, N4510);
or OR4 (N6301, N6297, N1607, N428, N2435);
xor XOR2 (N6302, N6296, N1558);
buf BUF1 (N6303, N6302);
and AND4 (N6304, N6298, N1291, N929, N471);
not NOT1 (N6305, N6272);
xor XOR2 (N6306, N6299, N4335);
xor XOR2 (N6307, N6303, N2598);
nor NOR4 (N6308, N6301, N176, N4245, N32);
nor NOR3 (N6309, N6284, N2388, N2770);
nor NOR3 (N6310, N6306, N2909, N1142);
not NOT1 (N6311, N6309);
nand NAND3 (N6312, N6305, N3509, N5353);
xor XOR2 (N6313, N6310, N997);
buf BUF1 (N6314, N6308);
nor NOR4 (N6315, N6307, N1192, N717, N4119);
xor XOR2 (N6316, N6312, N5698);
or OR3 (N6317, N6300, N213, N4962);
xor XOR2 (N6318, N6287, N4);
or OR2 (N6319, N6291, N1545);
not NOT1 (N6320, N6315);
nand NAND2 (N6321, N6313, N800);
nand NAND3 (N6322, N6320, N275, N3809);
xor XOR2 (N6323, N6311, N438);
or OR3 (N6324, N6323, N5569, N4458);
and AND2 (N6325, N6317, N2268);
xor XOR2 (N6326, N6304, N5487);
or OR3 (N6327, N6316, N5057, N4226);
buf BUF1 (N6328, N6321);
buf BUF1 (N6329, N6328);
or OR4 (N6330, N6325, N1744, N4926, N3231);
nand NAND4 (N6331, N6318, N1068, N5051, N5135);
nand NAND2 (N6332, N6326, N803);
or OR2 (N6333, N6322, N3261);
buf BUF1 (N6334, N6327);
nor NOR4 (N6335, N6279, N1010, N5897, N3347);
nand NAND3 (N6336, N6319, N3068, N3689);
or OR3 (N6337, N6329, N6323, N4902);
xor XOR2 (N6338, N6337, N2241);
and AND4 (N6339, N6333, N2774, N3401, N3291);
xor XOR2 (N6340, N6339, N80);
xor XOR2 (N6341, N6331, N5039);
and AND4 (N6342, N6340, N2105, N5558, N1623);
or OR3 (N6343, N6324, N1849, N5143);
not NOT1 (N6344, N6342);
not NOT1 (N6345, N6334);
nand NAND4 (N6346, N6336, N738, N1693, N2347);
and AND4 (N6347, N6346, N1410, N1151, N4167);
nor NOR4 (N6348, N6345, N4652, N5400, N230);
not NOT1 (N6349, N6348);
not NOT1 (N6350, N6314);
nand NAND3 (N6351, N6344, N1173, N754);
xor XOR2 (N6352, N6341, N786);
nand NAND4 (N6353, N6338, N299, N1407, N3001);
nor NOR3 (N6354, N6351, N3735, N513);
nand NAND3 (N6355, N6349, N1824, N1021);
and AND3 (N6356, N6355, N4623, N2260);
or OR4 (N6357, N6330, N145, N4368, N3844);
nor NOR2 (N6358, N6353, N2610);
nand NAND2 (N6359, N6332, N308);
or OR3 (N6360, N6354, N1557, N1901);
or OR3 (N6361, N6358, N16, N5375);
or OR2 (N6362, N6335, N5061);
not NOT1 (N6363, N6362);
or OR2 (N6364, N6356, N4120);
or OR4 (N6365, N6352, N400, N5795, N5281);
buf BUF1 (N6366, N6360);
and AND2 (N6367, N6347, N4016);
and AND4 (N6368, N6364, N6180, N4477, N2715);
xor XOR2 (N6369, N6368, N6174);
or OR4 (N6370, N6357, N3947, N5573, N661);
or OR3 (N6371, N6343, N4837, N5221);
not NOT1 (N6372, N6350);
not NOT1 (N6373, N6367);
or OR2 (N6374, N6372, N5823);
nand NAND3 (N6375, N6363, N3531, N5250);
not NOT1 (N6376, N6359);
nand NAND2 (N6377, N6361, N3383);
or OR3 (N6378, N6374, N5675, N508);
buf BUF1 (N6379, N6378);
nand NAND2 (N6380, N6370, N3565);
nand NAND2 (N6381, N6375, N6180);
xor XOR2 (N6382, N6376, N1886);
nor NOR2 (N6383, N6373, N5595);
buf BUF1 (N6384, N6365);
nor NOR2 (N6385, N6366, N1952);
xor XOR2 (N6386, N6377, N6159);
buf BUF1 (N6387, N6369);
not NOT1 (N6388, N6380);
not NOT1 (N6389, N6383);
xor XOR2 (N6390, N6388, N1445);
or OR3 (N6391, N6385, N4555, N2100);
not NOT1 (N6392, N6384);
buf BUF1 (N6393, N6387);
and AND3 (N6394, N6393, N2354, N2687);
xor XOR2 (N6395, N6392, N3303);
or OR4 (N6396, N6379, N4442, N5323, N2877);
nor NOR2 (N6397, N6382, N4900);
buf BUF1 (N6398, N6371);
nand NAND2 (N6399, N6398, N3950);
not NOT1 (N6400, N6391);
nor NOR2 (N6401, N6396, N2200);
xor XOR2 (N6402, N6389, N4303);
or OR3 (N6403, N6401, N3595, N3106);
xor XOR2 (N6404, N6397, N6193);
nor NOR4 (N6405, N6404, N6007, N6005, N1538);
and AND2 (N6406, N6405, N4602);
or OR3 (N6407, N6406, N6225, N5597);
xor XOR2 (N6408, N6400, N2683);
nand NAND4 (N6409, N6386, N54, N630, N3314);
or OR4 (N6410, N6394, N2276, N5917, N4166);
nand NAND2 (N6411, N6408, N4570);
xor XOR2 (N6412, N6390, N2219);
and AND4 (N6413, N6402, N3612, N5040, N4150);
or OR3 (N6414, N6407, N1618, N6344);
nor NOR4 (N6415, N6414, N3639, N3439, N2705);
xor XOR2 (N6416, N6403, N5514);
xor XOR2 (N6417, N6381, N4757);
or OR2 (N6418, N6412, N1209);
buf BUF1 (N6419, N6410);
not NOT1 (N6420, N6416);
or OR4 (N6421, N6417, N1091, N2050, N3560);
not NOT1 (N6422, N6413);
nor NOR2 (N6423, N6411, N4538);
xor XOR2 (N6424, N6423, N5510);
nor NOR2 (N6425, N6395, N684);
xor XOR2 (N6426, N6418, N2389);
xor XOR2 (N6427, N6409, N2112);
and AND2 (N6428, N6427, N1047);
not NOT1 (N6429, N6421);
nand NAND4 (N6430, N6429, N5533, N1335, N3048);
xor XOR2 (N6431, N6425, N4229);
buf BUF1 (N6432, N6422);
nand NAND4 (N6433, N6424, N5699, N6310, N819);
xor XOR2 (N6434, N6431, N5582);
buf BUF1 (N6435, N6430);
and AND3 (N6436, N6432, N4863, N517);
or OR3 (N6437, N6399, N5731, N5602);
nand NAND3 (N6438, N6433, N84, N2953);
buf BUF1 (N6439, N6420);
nand NAND4 (N6440, N6435, N1730, N2981, N1866);
not NOT1 (N6441, N6437);
or OR2 (N6442, N6440, N18);
xor XOR2 (N6443, N6415, N5762);
or OR3 (N6444, N6428, N3020, N2881);
or OR2 (N6445, N6438, N521);
or OR4 (N6446, N6444, N4576, N2714, N2177);
buf BUF1 (N6447, N6443);
nand NAND3 (N6448, N6445, N52, N2445);
xor XOR2 (N6449, N6446, N5379);
nor NOR2 (N6450, N6447, N416);
not NOT1 (N6451, N6434);
buf BUF1 (N6452, N6419);
or OR3 (N6453, N6448, N2622, N5928);
or OR3 (N6454, N6449, N446, N3606);
xor XOR2 (N6455, N6441, N3289);
not NOT1 (N6456, N6426);
nand NAND4 (N6457, N6456, N874, N1476, N1941);
or OR3 (N6458, N6439, N1794, N466);
nand NAND3 (N6459, N6450, N2839, N4321);
nor NOR4 (N6460, N6457, N370, N4348, N5119);
and AND2 (N6461, N6453, N3919);
not NOT1 (N6462, N6436);
nor NOR2 (N6463, N6442, N4372);
nand NAND4 (N6464, N6458, N2783, N5037, N2588);
and AND3 (N6465, N6454, N6087, N1058);
or OR3 (N6466, N6459, N6184, N268);
and AND2 (N6467, N6451, N2762);
nor NOR4 (N6468, N6455, N1369, N1864, N1249);
not NOT1 (N6469, N6461);
buf BUF1 (N6470, N6467);
nand NAND2 (N6471, N6469, N5625);
buf BUF1 (N6472, N6460);
not NOT1 (N6473, N6470);
not NOT1 (N6474, N6468);
or OR2 (N6475, N6462, N1761);
or OR3 (N6476, N6463, N2211, N648);
or OR2 (N6477, N6471, N6163);
xor XOR2 (N6478, N6452, N2856);
and AND4 (N6479, N6477, N2840, N4946, N5987);
buf BUF1 (N6480, N6466);
nor NOR2 (N6481, N6480, N4404);
nand NAND4 (N6482, N6479, N5675, N3710, N4092);
not NOT1 (N6483, N6474);
buf BUF1 (N6484, N6464);
not NOT1 (N6485, N6472);
or OR4 (N6486, N6482, N6162, N1450, N5960);
nand NAND4 (N6487, N6481, N2303, N4236, N1506);
xor XOR2 (N6488, N6483, N3345);
xor XOR2 (N6489, N6485, N1230);
not NOT1 (N6490, N6473);
or OR4 (N6491, N6484, N2028, N4100, N2281);
not NOT1 (N6492, N6476);
not NOT1 (N6493, N6487);
xor XOR2 (N6494, N6486, N6357);
xor XOR2 (N6495, N6489, N3518);
xor XOR2 (N6496, N6491, N3288);
xor XOR2 (N6497, N6478, N6183);
nor NOR3 (N6498, N6495, N4833, N1031);
nor NOR2 (N6499, N6465, N5495);
xor XOR2 (N6500, N6496, N4926);
nand NAND3 (N6501, N6500, N3034, N5358);
xor XOR2 (N6502, N6492, N934);
nand NAND3 (N6503, N6493, N6251, N2337);
buf BUF1 (N6504, N6498);
nand NAND2 (N6505, N6488, N2403);
nor NOR4 (N6506, N6497, N3428, N1687, N3192);
xor XOR2 (N6507, N6501, N5668);
and AND2 (N6508, N6507, N5678);
and AND4 (N6509, N6505, N4924, N2648, N5938);
xor XOR2 (N6510, N6503, N3294);
nand NAND2 (N6511, N6504, N4119);
not NOT1 (N6512, N6511);
xor XOR2 (N6513, N6499, N4629);
not NOT1 (N6514, N6512);
nor NOR2 (N6515, N6506, N1298);
nor NOR4 (N6516, N6475, N5950, N2250, N5757);
not NOT1 (N6517, N6490);
not NOT1 (N6518, N6502);
xor XOR2 (N6519, N6510, N4929);
buf BUF1 (N6520, N6517);
or OR4 (N6521, N6509, N5873, N5807, N246);
and AND3 (N6522, N6521, N5103, N1685);
xor XOR2 (N6523, N6520, N4248);
not NOT1 (N6524, N6519);
and AND4 (N6525, N6523, N1756, N4775, N5470);
nand NAND4 (N6526, N6522, N2007, N5092, N5936);
nand NAND4 (N6527, N6518, N5756, N2116, N398);
not NOT1 (N6528, N6516);
buf BUF1 (N6529, N6525);
buf BUF1 (N6530, N6527);
and AND2 (N6531, N6530, N2838);
not NOT1 (N6532, N6494);
or OR3 (N6533, N6529, N629, N2004);
and AND3 (N6534, N6528, N1453, N735);
nor NOR2 (N6535, N6534, N4440);
and AND4 (N6536, N6508, N1983, N6179, N3459);
nand NAND2 (N6537, N6524, N2808);
nor NOR4 (N6538, N6532, N831, N2258, N2601);
and AND4 (N6539, N6513, N3555, N2760, N4149);
nor NOR4 (N6540, N6514, N3305, N3994, N1454);
not NOT1 (N6541, N6536);
buf BUF1 (N6542, N6515);
not NOT1 (N6543, N6539);
buf BUF1 (N6544, N6531);
or OR3 (N6545, N6538, N2563, N1656);
or OR3 (N6546, N6541, N5425, N3126);
nand NAND2 (N6547, N6533, N5983);
and AND4 (N6548, N6545, N3198, N3067, N1620);
not NOT1 (N6549, N6540);
not NOT1 (N6550, N6549);
xor XOR2 (N6551, N6535, N5865);
and AND3 (N6552, N6546, N3504, N2490);
or OR3 (N6553, N6547, N2548, N3049);
nand NAND4 (N6554, N6551, N4113, N3290, N3536);
nand NAND3 (N6555, N6554, N5516, N3061);
buf BUF1 (N6556, N6552);
buf BUF1 (N6557, N6544);
not NOT1 (N6558, N6557);
nand NAND3 (N6559, N6526, N6043, N3742);
nor NOR3 (N6560, N6542, N203, N3483);
nor NOR4 (N6561, N6537, N2097, N2505, N5076);
nand NAND4 (N6562, N6561, N5473, N3590, N3677);
and AND2 (N6563, N6555, N4270);
nand NAND4 (N6564, N6558, N6045, N3724, N4108);
and AND4 (N6565, N6562, N2898, N5134, N2641);
and AND4 (N6566, N6559, N5745, N5241, N6383);
nand NAND3 (N6567, N6564, N2797, N4646);
and AND3 (N6568, N6560, N4062, N2930);
not NOT1 (N6569, N6556);
xor XOR2 (N6570, N6548, N2937);
or OR2 (N6571, N6568, N616);
not NOT1 (N6572, N6569);
or OR4 (N6573, N6572, N6124, N1650, N1577);
and AND4 (N6574, N6553, N5217, N5003, N475);
or OR2 (N6575, N6566, N1429);
nor NOR4 (N6576, N6575, N727, N966, N5492);
not NOT1 (N6577, N6571);
nor NOR2 (N6578, N6550, N1534);
xor XOR2 (N6579, N6565, N3485);
xor XOR2 (N6580, N6577, N2627);
nand NAND3 (N6581, N6579, N749, N2452);
nor NOR2 (N6582, N6576, N2605);
nor NOR2 (N6583, N6581, N621);
xor XOR2 (N6584, N6573, N691);
xor XOR2 (N6585, N6570, N6406);
and AND2 (N6586, N6580, N4818);
and AND3 (N6587, N6586, N3190, N5954);
buf BUF1 (N6588, N6585);
xor XOR2 (N6589, N6563, N2251);
buf BUF1 (N6590, N6574);
or OR4 (N6591, N6578, N1448, N5811, N3537);
and AND4 (N6592, N6587, N959, N2321, N160);
nor NOR4 (N6593, N6592, N4395, N9, N6569);
and AND4 (N6594, N6543, N3341, N1062, N6549);
not NOT1 (N6595, N6591);
xor XOR2 (N6596, N6588, N2433);
and AND4 (N6597, N6593, N4492, N3528, N3814);
not NOT1 (N6598, N6584);
buf BUF1 (N6599, N6567);
nor NOR3 (N6600, N6590, N6225, N3875);
nand NAND4 (N6601, N6597, N4022, N5083, N3738);
xor XOR2 (N6602, N6601, N2451);
not NOT1 (N6603, N6594);
xor XOR2 (N6604, N6596, N1101);
not NOT1 (N6605, N6583);
nand NAND4 (N6606, N6589, N792, N6200, N3588);
or OR3 (N6607, N6602, N3398, N1063);
nand NAND4 (N6608, N6599, N2961, N1949, N5558);
or OR2 (N6609, N6606, N369);
nor NOR4 (N6610, N6609, N4204, N762, N5135);
nand NAND2 (N6611, N6600, N4338);
buf BUF1 (N6612, N6582);
nor NOR2 (N6613, N6607, N1463);
not NOT1 (N6614, N6611);
nand NAND3 (N6615, N6603, N1288, N1957);
xor XOR2 (N6616, N6614, N5215);
buf BUF1 (N6617, N6598);
buf BUF1 (N6618, N6613);
buf BUF1 (N6619, N6617);
or OR3 (N6620, N6615, N1173, N4266);
nand NAND4 (N6621, N6608, N5342, N1129, N2109);
not NOT1 (N6622, N6618);
not NOT1 (N6623, N6616);
and AND3 (N6624, N6623, N5964, N2653);
or OR2 (N6625, N6595, N1762);
not NOT1 (N6626, N6619);
xor XOR2 (N6627, N6605, N1369);
and AND4 (N6628, N6627, N4574, N2161, N208);
not NOT1 (N6629, N6620);
not NOT1 (N6630, N6629);
nor NOR2 (N6631, N6624, N448);
and AND4 (N6632, N6622, N1533, N1265, N687);
and AND3 (N6633, N6621, N4593, N4461);
not NOT1 (N6634, N6631);
or OR2 (N6635, N6604, N1890);
not NOT1 (N6636, N6630);
not NOT1 (N6637, N6635);
not NOT1 (N6638, N6634);
nor NOR2 (N6639, N6610, N2076);
nor NOR2 (N6640, N6612, N2338);
buf BUF1 (N6641, N6625);
buf BUF1 (N6642, N6633);
and AND2 (N6643, N6632, N4220);
buf BUF1 (N6644, N6636);
nand NAND2 (N6645, N6639, N3558);
xor XOR2 (N6646, N6642, N1918);
nand NAND2 (N6647, N6626, N6145);
and AND4 (N6648, N6645, N5952, N5295, N2638);
and AND3 (N6649, N6644, N2777, N5250);
buf BUF1 (N6650, N6641);
not NOT1 (N6651, N6650);
buf BUF1 (N6652, N6637);
not NOT1 (N6653, N6640);
and AND4 (N6654, N6653, N2663, N5246, N4304);
or OR3 (N6655, N6628, N6097, N2254);
nor NOR4 (N6656, N6649, N4044, N1570, N3972);
not NOT1 (N6657, N6656);
xor XOR2 (N6658, N6647, N1872);
xor XOR2 (N6659, N6651, N4314);
nor NOR4 (N6660, N6652, N1590, N142, N3414);
nor NOR3 (N6661, N6646, N757, N923);
not NOT1 (N6662, N6657);
not NOT1 (N6663, N6648);
buf BUF1 (N6664, N6654);
xor XOR2 (N6665, N6659, N947);
not NOT1 (N6666, N6643);
or OR2 (N6667, N6638, N2486);
not NOT1 (N6668, N6662);
or OR2 (N6669, N6664, N6394);
and AND3 (N6670, N6667, N1973, N3981);
not NOT1 (N6671, N6661);
nand NAND2 (N6672, N6668, N1835);
nor NOR4 (N6673, N6671, N149, N5464, N676);
xor XOR2 (N6674, N6670, N5872);
or OR3 (N6675, N6674, N1641, N2886);
nor NOR2 (N6676, N6660, N4936);
buf BUF1 (N6677, N6676);
and AND2 (N6678, N6675, N983);
nand NAND3 (N6679, N6663, N2014, N1939);
nor NOR2 (N6680, N6658, N2431);
xor XOR2 (N6681, N6669, N6670);
nand NAND3 (N6682, N6666, N2144, N3412);
nor NOR4 (N6683, N6680, N3637, N1861, N5839);
or OR4 (N6684, N6681, N5100, N3451, N2690);
not NOT1 (N6685, N6684);
not NOT1 (N6686, N6672);
xor XOR2 (N6687, N6683, N5242);
not NOT1 (N6688, N6673);
xor XOR2 (N6689, N6679, N2990);
xor XOR2 (N6690, N6678, N3585);
nand NAND2 (N6691, N6689, N5423);
not NOT1 (N6692, N6677);
nor NOR3 (N6693, N6692, N6298, N2738);
buf BUF1 (N6694, N6688);
buf BUF1 (N6695, N6686);
nand NAND3 (N6696, N6655, N506, N3440);
buf BUF1 (N6697, N6685);
nand NAND4 (N6698, N6697, N6498, N562, N4619);
not NOT1 (N6699, N6698);
nand NAND4 (N6700, N6690, N3528, N1347, N3181);
and AND2 (N6701, N6694, N2572);
nand NAND2 (N6702, N6687, N1279);
not NOT1 (N6703, N6682);
not NOT1 (N6704, N6701);
and AND3 (N6705, N6696, N5786, N4953);
buf BUF1 (N6706, N6665);
nand NAND3 (N6707, N6703, N1927, N4120);
buf BUF1 (N6708, N6691);
and AND3 (N6709, N6706, N2967, N3067);
nor NOR4 (N6710, N6709, N3566, N2498, N5419);
or OR2 (N6711, N6705, N2565);
and AND3 (N6712, N6695, N2680, N6627);
xor XOR2 (N6713, N6700, N298);
not NOT1 (N6714, N6712);
nor NOR4 (N6715, N6693, N207, N3011, N4605);
xor XOR2 (N6716, N6707, N1387);
buf BUF1 (N6717, N6708);
not NOT1 (N6718, N6713);
and AND4 (N6719, N6711, N1746, N4186, N136);
xor XOR2 (N6720, N6718, N1870);
nand NAND2 (N6721, N6720, N6563);
not NOT1 (N6722, N6721);
and AND4 (N6723, N6716, N2592, N118, N2954);
buf BUF1 (N6724, N6702);
and AND3 (N6725, N6724, N1627, N4187);
nor NOR3 (N6726, N6725, N666, N1907);
not NOT1 (N6727, N6715);
or OR2 (N6728, N6717, N3385);
buf BUF1 (N6729, N6714);
xor XOR2 (N6730, N6728, N5148);
xor XOR2 (N6731, N6726, N6361);
xor XOR2 (N6732, N6722, N5242);
nor NOR4 (N6733, N6729, N6684, N3935, N4006);
nand NAND3 (N6734, N6710, N4262, N4004);
nor NOR3 (N6735, N6732, N1664, N3437);
nand NAND2 (N6736, N6723, N1578);
buf BUF1 (N6737, N6727);
buf BUF1 (N6738, N6734);
not NOT1 (N6739, N6738);
or OR2 (N6740, N6735, N3830);
xor XOR2 (N6741, N6719, N1360);
and AND2 (N6742, N6737, N1290);
and AND2 (N6743, N6731, N4803);
xor XOR2 (N6744, N6730, N3832);
and AND3 (N6745, N6739, N1908, N403);
not NOT1 (N6746, N6741);
nor NOR3 (N6747, N6740, N877, N4407);
nor NOR4 (N6748, N6743, N4441, N2268, N896);
xor XOR2 (N6749, N6745, N1197);
not NOT1 (N6750, N6746);
nand NAND3 (N6751, N6736, N4800, N1823);
not NOT1 (N6752, N6747);
buf BUF1 (N6753, N6748);
and AND3 (N6754, N6733, N960, N4487);
nor NOR3 (N6755, N6752, N6503, N5478);
not NOT1 (N6756, N6742);
nor NOR2 (N6757, N6750, N2839);
nor NOR3 (N6758, N6753, N3518, N3614);
not NOT1 (N6759, N6704);
not NOT1 (N6760, N6756);
buf BUF1 (N6761, N6759);
or OR4 (N6762, N6754, N346, N1357, N6564);
nor NOR4 (N6763, N6760, N2502, N4318, N2970);
and AND2 (N6764, N6744, N6034);
buf BUF1 (N6765, N6758);
nor NOR2 (N6766, N6764, N4993);
or OR2 (N6767, N6766, N3642);
and AND3 (N6768, N6755, N949, N2056);
not NOT1 (N6769, N6763);
xor XOR2 (N6770, N6757, N1813);
or OR2 (N6771, N6769, N3560);
nor NOR4 (N6772, N6761, N6752, N2547, N806);
nor NOR2 (N6773, N6771, N5804);
not NOT1 (N6774, N6772);
nor NOR3 (N6775, N6762, N5363, N4891);
or OR3 (N6776, N6699, N2706, N434);
xor XOR2 (N6777, N6770, N5002);
or OR3 (N6778, N6749, N6284, N2523);
nand NAND3 (N6779, N6775, N3930, N2475);
buf BUF1 (N6780, N6773);
xor XOR2 (N6781, N6778, N3738);
not NOT1 (N6782, N6780);
nand NAND2 (N6783, N6777, N545);
xor XOR2 (N6784, N6774, N6450);
and AND3 (N6785, N6765, N1482, N81);
nor NOR2 (N6786, N6783, N1746);
not NOT1 (N6787, N6768);
nand NAND2 (N6788, N6781, N5221);
nor NOR2 (N6789, N6786, N3289);
and AND2 (N6790, N6789, N3189);
not NOT1 (N6791, N6776);
xor XOR2 (N6792, N6779, N2554);
not NOT1 (N6793, N6787);
not NOT1 (N6794, N6790);
xor XOR2 (N6795, N6794, N3136);
nor NOR2 (N6796, N6793, N1049);
nand NAND3 (N6797, N6785, N5405, N4024);
nand NAND4 (N6798, N6782, N5596, N5665, N2594);
xor XOR2 (N6799, N6797, N3857);
or OR2 (N6800, N6784, N3130);
buf BUF1 (N6801, N6800);
not NOT1 (N6802, N6791);
nor NOR3 (N6803, N6795, N5888, N4967);
buf BUF1 (N6804, N6802);
nor NOR4 (N6805, N6788, N2327, N3397, N4563);
nand NAND2 (N6806, N6804, N6392);
not NOT1 (N6807, N6803);
buf BUF1 (N6808, N6806);
nor NOR2 (N6809, N6796, N3581);
nand NAND2 (N6810, N6809, N2862);
xor XOR2 (N6811, N6807, N4435);
not NOT1 (N6812, N6767);
xor XOR2 (N6813, N6792, N2758);
xor XOR2 (N6814, N6811, N1175);
and AND2 (N6815, N6751, N3596);
xor XOR2 (N6816, N6798, N1904);
buf BUF1 (N6817, N6812);
nor NOR2 (N6818, N6817, N3128);
not NOT1 (N6819, N6810);
nor NOR2 (N6820, N6801, N4943);
and AND3 (N6821, N6820, N6530, N5557);
nor NOR3 (N6822, N6819, N4510, N4356);
not NOT1 (N6823, N6808);
buf BUF1 (N6824, N6821);
nand NAND4 (N6825, N6813, N5312, N2992, N3245);
nand NAND3 (N6826, N6824, N5056, N3441);
and AND3 (N6827, N6815, N4321, N924);
nand NAND2 (N6828, N6805, N2611);
or OR4 (N6829, N6828, N2741, N2724, N5843);
xor XOR2 (N6830, N6818, N711);
xor XOR2 (N6831, N6799, N3838);
or OR3 (N6832, N6825, N37, N4193);
nor NOR4 (N6833, N6822, N182, N4628, N608);
buf BUF1 (N6834, N6829);
buf BUF1 (N6835, N6833);
not NOT1 (N6836, N6823);
or OR3 (N6837, N6827, N4529, N808);
nor NOR3 (N6838, N6835, N2825, N1738);
xor XOR2 (N6839, N6826, N245);
buf BUF1 (N6840, N6816);
nor NOR2 (N6841, N6839, N3590);
nor NOR2 (N6842, N6836, N2143);
or OR2 (N6843, N6841, N6828);
or OR3 (N6844, N6837, N4987, N6658);
xor XOR2 (N6845, N6843, N4572);
xor XOR2 (N6846, N6834, N4006);
and AND3 (N6847, N6842, N3370, N5730);
xor XOR2 (N6848, N6831, N1148);
and AND2 (N6849, N6830, N6716);
not NOT1 (N6850, N6844);
nor NOR2 (N6851, N6850, N4471);
or OR2 (N6852, N6832, N1317);
buf BUF1 (N6853, N6840);
xor XOR2 (N6854, N6846, N4456);
nand NAND3 (N6855, N6838, N3521, N5552);
nand NAND4 (N6856, N6849, N2636, N3176, N3093);
nor NOR4 (N6857, N6853, N6086, N2505, N230);
and AND4 (N6858, N6852, N3286, N6678, N4931);
nand NAND2 (N6859, N6847, N6288);
or OR3 (N6860, N6856, N5494, N4301);
nand NAND3 (N6861, N6854, N3386, N5039);
xor XOR2 (N6862, N6855, N5662);
and AND3 (N6863, N6857, N5060, N3171);
buf BUF1 (N6864, N6859);
nand NAND2 (N6865, N6860, N3546);
nor NOR4 (N6866, N6864, N5731, N5218, N3929);
buf BUF1 (N6867, N6851);
or OR3 (N6868, N6863, N6685, N5421);
nor NOR3 (N6869, N6848, N3453, N4861);
xor XOR2 (N6870, N6814, N5463);
xor XOR2 (N6871, N6858, N6137);
nand NAND4 (N6872, N6869, N2674, N4442, N1101);
nand NAND4 (N6873, N6866, N1764, N1234, N1324);
or OR4 (N6874, N6865, N854, N425, N2355);
nor NOR4 (N6875, N6862, N4264, N1859, N5439);
or OR4 (N6876, N6871, N637, N953, N4296);
and AND4 (N6877, N6868, N2740, N579, N5513);
or OR3 (N6878, N6872, N2589, N1541);
and AND3 (N6879, N6867, N5644, N5817);
xor XOR2 (N6880, N6876, N3697);
nand NAND2 (N6881, N6879, N210);
buf BUF1 (N6882, N6875);
buf BUF1 (N6883, N6870);
xor XOR2 (N6884, N6883, N5867);
or OR4 (N6885, N6873, N6795, N5247, N6483);
nor NOR4 (N6886, N6884, N3174, N788, N3236);
nand NAND3 (N6887, N6845, N1286, N6042);
or OR4 (N6888, N6882, N4541, N1181, N5767);
xor XOR2 (N6889, N6886, N2258);
buf BUF1 (N6890, N6878);
nand NAND4 (N6891, N6881, N5183, N4739, N3969);
buf BUF1 (N6892, N6890);
nor NOR3 (N6893, N6887, N6214, N4099);
or OR4 (N6894, N6874, N3803, N320, N19);
nor NOR2 (N6895, N6885, N2589);
nand NAND2 (N6896, N6889, N232);
buf BUF1 (N6897, N6895);
nand NAND2 (N6898, N6880, N1198);
buf BUF1 (N6899, N6896);
or OR4 (N6900, N6877, N2459, N5207, N4881);
xor XOR2 (N6901, N6892, N239);
or OR4 (N6902, N6899, N4777, N3209, N2633);
buf BUF1 (N6903, N6888);
not NOT1 (N6904, N6861);
and AND4 (N6905, N6902, N2646, N685, N3252);
and AND4 (N6906, N6897, N2394, N1800, N2175);
not NOT1 (N6907, N6898);
and AND4 (N6908, N6894, N6888, N537, N6427);
and AND3 (N6909, N6908, N678, N2038);
xor XOR2 (N6910, N6907, N5751);
nand NAND3 (N6911, N6909, N2917, N407);
or OR3 (N6912, N6891, N6398, N1702);
nor NOR2 (N6913, N6900, N731);
and AND2 (N6914, N6904, N957);
nor NOR2 (N6915, N6903, N1238);
not NOT1 (N6916, N6893);
buf BUF1 (N6917, N6912);
not NOT1 (N6918, N6915);
buf BUF1 (N6919, N6901);
not NOT1 (N6920, N6906);
or OR3 (N6921, N6913, N850, N730);
nand NAND2 (N6922, N6918, N4172);
buf BUF1 (N6923, N6917);
nor NOR4 (N6924, N6921, N2818, N551, N964);
nor NOR3 (N6925, N6919, N5142, N5047);
not NOT1 (N6926, N6914);
not NOT1 (N6927, N6923);
not NOT1 (N6928, N6910);
nand NAND4 (N6929, N6916, N837, N542, N4398);
not NOT1 (N6930, N6925);
and AND2 (N6931, N6905, N5559);
and AND3 (N6932, N6911, N5049, N5113);
and AND3 (N6933, N6932, N6797, N4295);
xor XOR2 (N6934, N6930, N638);
not NOT1 (N6935, N6922);
not NOT1 (N6936, N6920);
nand NAND3 (N6937, N6929, N1227, N5379);
buf BUF1 (N6938, N6936);
not NOT1 (N6939, N6927);
nand NAND3 (N6940, N6931, N972, N2923);
nand NAND2 (N6941, N6933, N6375);
buf BUF1 (N6942, N6940);
nand NAND3 (N6943, N6935, N5790, N3365);
buf BUF1 (N6944, N6941);
nand NAND3 (N6945, N6943, N6511, N2211);
or OR2 (N6946, N6942, N2455);
not NOT1 (N6947, N6926);
xor XOR2 (N6948, N6946, N3469);
buf BUF1 (N6949, N6947);
nand NAND2 (N6950, N6924, N6530);
nand NAND3 (N6951, N6950, N53, N3333);
nand NAND2 (N6952, N6949, N1008);
not NOT1 (N6953, N6951);
xor XOR2 (N6954, N6952, N5845);
buf BUF1 (N6955, N6945);
nand NAND4 (N6956, N6937, N4276, N2484, N3756);
or OR4 (N6957, N6956, N6208, N1592, N1913);
xor XOR2 (N6958, N6939, N888);
and AND4 (N6959, N6938, N1857, N2514, N4108);
nand NAND3 (N6960, N6948, N1706, N3248);
not NOT1 (N6961, N6959);
and AND4 (N6962, N6934, N917, N2572, N289);
not NOT1 (N6963, N6955);
nand NAND2 (N6964, N6928, N1957);
not NOT1 (N6965, N6953);
nand NAND2 (N6966, N6964, N6344);
xor XOR2 (N6967, N6962, N5603);
nor NOR3 (N6968, N6958, N5977, N5754);
xor XOR2 (N6969, N6957, N753);
xor XOR2 (N6970, N6968, N2397);
xor XOR2 (N6971, N6960, N3815);
or OR2 (N6972, N6970, N2126);
nor NOR3 (N6973, N6969, N1382, N943);
nand NAND4 (N6974, N6965, N2105, N1174, N5904);
or OR3 (N6975, N6963, N514, N3425);
buf BUF1 (N6976, N6967);
nand NAND3 (N6977, N6972, N1132, N6390);
nor NOR3 (N6978, N6973, N833, N4168);
nor NOR2 (N6979, N6976, N4457);
nor NOR3 (N6980, N6978, N4775, N5981);
or OR2 (N6981, N6966, N3784);
xor XOR2 (N6982, N6944, N6585);
not NOT1 (N6983, N6979);
buf BUF1 (N6984, N6974);
and AND3 (N6985, N6954, N3916, N4748);
xor XOR2 (N6986, N6984, N5007);
nor NOR4 (N6987, N6985, N4748, N2803, N3764);
nand NAND2 (N6988, N6981, N5756);
buf BUF1 (N6989, N6975);
xor XOR2 (N6990, N6987, N3084);
nand NAND4 (N6991, N6983, N6787, N1360, N3144);
not NOT1 (N6992, N6988);
not NOT1 (N6993, N6982);
nor NOR2 (N6994, N6993, N2527);
not NOT1 (N6995, N6990);
nand NAND2 (N6996, N6980, N1645);
and AND4 (N6997, N6989, N6360, N3172, N6949);
buf BUF1 (N6998, N6977);
not NOT1 (N6999, N6961);
or OR4 (N7000, N6994, N1307, N4113, N260);
nand NAND4 (N7001, N7000, N3788, N6465, N2318);
and AND3 (N7002, N7001, N1783, N4523);
buf BUF1 (N7003, N6986);
nand NAND4 (N7004, N6991, N4340, N4214, N6057);
not NOT1 (N7005, N6995);
xor XOR2 (N7006, N6971, N343);
not NOT1 (N7007, N7003);
not NOT1 (N7008, N6999);
not NOT1 (N7009, N7006);
not NOT1 (N7010, N6996);
nor NOR2 (N7011, N7008, N2257);
nor NOR2 (N7012, N6998, N3025);
nor NOR2 (N7013, N7010, N4816);
or OR4 (N7014, N7002, N3190, N2598, N78);
and AND3 (N7015, N7013, N2535, N716);
nor NOR3 (N7016, N7007, N5289, N5885);
nor NOR4 (N7017, N7004, N6372, N5535, N3137);
nor NOR3 (N7018, N7017, N4154, N5483);
and AND3 (N7019, N7016, N5730, N1851);
xor XOR2 (N7020, N7015, N2815);
buf BUF1 (N7021, N7014);
buf BUF1 (N7022, N7021);
and AND3 (N7023, N7019, N3938, N6705);
not NOT1 (N7024, N6997);
nor NOR2 (N7025, N7009, N1644);
nand NAND2 (N7026, N6992, N2715);
or OR2 (N7027, N7012, N5759);
nand NAND4 (N7028, N7018, N4556, N1071, N427);
xor XOR2 (N7029, N7005, N4708);
nand NAND2 (N7030, N7020, N999);
nand NAND3 (N7031, N7025, N6388, N3544);
xor XOR2 (N7032, N7026, N4964);
xor XOR2 (N7033, N7027, N6736);
and AND3 (N7034, N7031, N6355, N2162);
and AND4 (N7035, N7034, N2133, N5291, N325);
not NOT1 (N7036, N7011);
nand NAND3 (N7037, N7023, N2715, N469);
nor NOR4 (N7038, N7028, N2614, N3180, N5562);
and AND3 (N7039, N7030, N2787, N4386);
nor NOR4 (N7040, N7035, N3974, N5311, N1754);
buf BUF1 (N7041, N7033);
or OR4 (N7042, N7022, N566, N563, N4742);
nor NOR4 (N7043, N7038, N6141, N3841, N5391);
xor XOR2 (N7044, N7039, N3066);
and AND4 (N7045, N7042, N1902, N2097, N4613);
xor XOR2 (N7046, N7036, N497);
xor XOR2 (N7047, N7045, N2894);
or OR2 (N7048, N7029, N44);
and AND4 (N7049, N7037, N1755, N1875, N1672);
and AND2 (N7050, N7024, N5669);
nand NAND3 (N7051, N7050, N3874, N558);
or OR3 (N7052, N7032, N1480, N4490);
not NOT1 (N7053, N7051);
and AND4 (N7054, N7052, N532, N2163, N4518);
xor XOR2 (N7055, N7054, N5071);
and AND3 (N7056, N7055, N1564, N6785);
or OR4 (N7057, N7053, N2816, N6500, N5865);
not NOT1 (N7058, N7041);
nand NAND4 (N7059, N7043, N6741, N5563, N5683);
and AND4 (N7060, N7056, N2716, N2154, N5196);
or OR2 (N7061, N7040, N4892);
or OR4 (N7062, N7048, N1291, N1542, N1102);
buf BUF1 (N7063, N7059);
nor NOR2 (N7064, N7062, N1621);
nor NOR4 (N7065, N7049, N4821, N4611, N76);
buf BUF1 (N7066, N7044);
buf BUF1 (N7067, N7058);
not NOT1 (N7068, N7063);
or OR3 (N7069, N7047, N3428, N4737);
or OR4 (N7070, N7061, N6863, N4064, N3827);
nand NAND4 (N7071, N7065, N6112, N5613, N3317);
or OR2 (N7072, N7069, N6725);
buf BUF1 (N7073, N7060);
and AND4 (N7074, N7068, N5979, N4139, N392);
xor XOR2 (N7075, N7057, N6136);
buf BUF1 (N7076, N7072);
not NOT1 (N7077, N7075);
not NOT1 (N7078, N7073);
buf BUF1 (N7079, N7064);
not NOT1 (N7080, N7071);
nor NOR4 (N7081, N7079, N2985, N5381, N527);
not NOT1 (N7082, N7070);
nand NAND3 (N7083, N7078, N1738, N7015);
nor NOR2 (N7084, N7066, N3215);
nor NOR4 (N7085, N7084, N4979, N2727, N550);
nor NOR2 (N7086, N7082, N539);
nand NAND2 (N7087, N7046, N1677);
or OR4 (N7088, N7085, N6565, N1910, N4888);
nor NOR2 (N7089, N7086, N5500);
not NOT1 (N7090, N7081);
nand NAND2 (N7091, N7089, N6524);
or OR2 (N7092, N7067, N3190);
buf BUF1 (N7093, N7083);
buf BUF1 (N7094, N7076);
nand NAND3 (N7095, N7080, N7071, N966);
and AND3 (N7096, N7094, N3644, N2381);
or OR2 (N7097, N7093, N3438);
nor NOR4 (N7098, N7095, N5131, N3170, N3253);
nor NOR2 (N7099, N7092, N5958);
buf BUF1 (N7100, N7096);
and AND3 (N7101, N7099, N4106, N1792);
not NOT1 (N7102, N7098);
nand NAND4 (N7103, N7087, N684, N6277, N4740);
or OR4 (N7104, N7103, N693, N3867, N3771);
or OR3 (N7105, N7090, N148, N661);
buf BUF1 (N7106, N7097);
nor NOR4 (N7107, N7105, N5359, N1181, N914);
and AND4 (N7108, N7102, N6943, N5501, N2529);
xor XOR2 (N7109, N7108, N5049);
nand NAND4 (N7110, N7109, N582, N2444, N604);
nand NAND4 (N7111, N7091, N4618, N5614, N1930);
nor NOR2 (N7112, N7104, N2676);
nand NAND2 (N7113, N7112, N4396);
and AND4 (N7114, N7088, N6644, N2338, N1226);
buf BUF1 (N7115, N7101);
nor NOR2 (N7116, N7113, N6786);
xor XOR2 (N7117, N7100, N5376);
or OR2 (N7118, N7074, N302);
nor NOR2 (N7119, N7117, N3628);
nand NAND2 (N7120, N7116, N2473);
nand NAND2 (N7121, N7106, N2244);
nand NAND3 (N7122, N7121, N4895, N3299);
and AND3 (N7123, N7110, N4284, N3612);
nand NAND3 (N7124, N7118, N3961, N2990);
nand NAND2 (N7125, N7119, N3275);
and AND3 (N7126, N7122, N6719, N2074);
and AND3 (N7127, N7077, N904, N4420);
buf BUF1 (N7128, N7123);
and AND4 (N7129, N7126, N6891, N5859, N3001);
or OR2 (N7130, N7127, N3905);
xor XOR2 (N7131, N7129, N5226);
nand NAND2 (N7132, N7124, N4253);
nor NOR3 (N7133, N7111, N6878, N6950);
not NOT1 (N7134, N7120);
xor XOR2 (N7135, N7125, N5280);
not NOT1 (N7136, N7131);
buf BUF1 (N7137, N7135);
and AND2 (N7138, N7133, N1791);
or OR3 (N7139, N7132, N2626, N3757);
nand NAND4 (N7140, N7114, N4205, N4890, N3676);
xor XOR2 (N7141, N7139, N3699);
or OR2 (N7142, N7115, N4259);
nand NAND4 (N7143, N7142, N4545, N5109, N6770);
buf BUF1 (N7144, N7138);
not NOT1 (N7145, N7140);
nor NOR3 (N7146, N7144, N3159, N5228);
buf BUF1 (N7147, N7134);
or OR4 (N7148, N7128, N2453, N6864, N5230);
nor NOR3 (N7149, N7148, N1121, N27);
xor XOR2 (N7150, N7145, N1907);
xor XOR2 (N7151, N7147, N5102);
not NOT1 (N7152, N7151);
or OR3 (N7153, N7107, N4409, N1879);
buf BUF1 (N7154, N7149);
and AND3 (N7155, N7150, N6829, N2616);
nor NOR3 (N7156, N7136, N5707, N5613);
buf BUF1 (N7157, N7146);
buf BUF1 (N7158, N7153);
nor NOR4 (N7159, N7137, N6508, N1930, N2438);
and AND2 (N7160, N7159, N346);
not NOT1 (N7161, N7143);
xor XOR2 (N7162, N7156, N6053);
xor XOR2 (N7163, N7141, N2014);
nand NAND4 (N7164, N7161, N5833, N3777, N508);
buf BUF1 (N7165, N7163);
xor XOR2 (N7166, N7130, N3825);
nand NAND3 (N7167, N7162, N2010, N2400);
not NOT1 (N7168, N7165);
nand NAND2 (N7169, N7158, N1671);
nand NAND3 (N7170, N7160, N4581, N6945);
and AND3 (N7171, N7157, N3452, N4194);
nor NOR3 (N7172, N7166, N3387, N1264);
not NOT1 (N7173, N7170);
or OR3 (N7174, N7173, N228, N5438);
and AND3 (N7175, N7171, N1086, N6674);
nor NOR2 (N7176, N7169, N5558);
not NOT1 (N7177, N7176);
buf BUF1 (N7178, N7164);
and AND4 (N7179, N7177, N2659, N3269, N6870);
buf BUF1 (N7180, N7175);
xor XOR2 (N7181, N7152, N3276);
and AND4 (N7182, N7155, N352, N5465, N4809);
or OR4 (N7183, N7182, N1452, N3506, N5503);
xor XOR2 (N7184, N7178, N3972);
nand NAND4 (N7185, N7154, N3301, N2530, N511);
nor NOR2 (N7186, N7181, N2082);
xor XOR2 (N7187, N7179, N126);
not NOT1 (N7188, N7174);
nand NAND4 (N7189, N7168, N6370, N73, N5977);
buf BUF1 (N7190, N7184);
buf BUF1 (N7191, N7189);
buf BUF1 (N7192, N7190);
nor NOR2 (N7193, N7183, N3010);
xor XOR2 (N7194, N7185, N2518);
xor XOR2 (N7195, N7167, N1389);
nor NOR2 (N7196, N7187, N4172);
xor XOR2 (N7197, N7193, N4539);
not NOT1 (N7198, N7186);
or OR2 (N7199, N7194, N4897);
nand NAND2 (N7200, N7199, N2063);
not NOT1 (N7201, N7196);
xor XOR2 (N7202, N7195, N3383);
or OR4 (N7203, N7180, N189, N3208, N6116);
nand NAND3 (N7204, N7188, N5042, N547);
not NOT1 (N7205, N7198);
nor NOR3 (N7206, N7172, N3353, N6482);
or OR3 (N7207, N7201, N3819, N2625);
buf BUF1 (N7208, N7192);
or OR2 (N7209, N7203, N133);
or OR2 (N7210, N7207, N4142);
xor XOR2 (N7211, N7206, N6562);
nor NOR2 (N7212, N7202, N6916);
or OR4 (N7213, N7205, N3636, N3532, N3565);
not NOT1 (N7214, N7212);
buf BUF1 (N7215, N7209);
xor XOR2 (N7216, N7214, N5086);
xor XOR2 (N7217, N7213, N3270);
nand NAND3 (N7218, N7197, N2702, N1715);
and AND4 (N7219, N7200, N5729, N3152, N2447);
and AND2 (N7220, N7208, N3801);
or OR4 (N7221, N7191, N1319, N6087, N82);
not NOT1 (N7222, N7204);
nand NAND4 (N7223, N7210, N3279, N1391, N5684);
nor NOR2 (N7224, N7219, N1863);
nor NOR3 (N7225, N7221, N3776, N1509);
nand NAND2 (N7226, N7225, N6933);
xor XOR2 (N7227, N7217, N4392);
nand NAND4 (N7228, N7215, N3710, N1023, N6205);
nand NAND2 (N7229, N7218, N3712);
or OR3 (N7230, N7211, N2525, N3259);
or OR2 (N7231, N7229, N6040);
nand NAND4 (N7232, N7220, N977, N2108, N3555);
nor NOR2 (N7233, N7232, N7016);
or OR3 (N7234, N7216, N1109, N5648);
not NOT1 (N7235, N7226);
nor NOR3 (N7236, N7230, N3265, N5603);
or OR4 (N7237, N7227, N4387, N3960, N7011);
or OR4 (N7238, N7224, N6573, N882, N6741);
nor NOR4 (N7239, N7234, N6846, N5671, N4538);
not NOT1 (N7240, N7235);
and AND4 (N7241, N7231, N6942, N3467, N5184);
nor NOR4 (N7242, N7238, N5882, N4833, N6704);
and AND3 (N7243, N7222, N2319, N3030);
and AND3 (N7244, N7228, N886, N4000);
buf BUF1 (N7245, N7244);
or OR4 (N7246, N7242, N214, N4121, N4103);
nand NAND4 (N7247, N7236, N4632, N5329, N3030);
nand NAND3 (N7248, N7239, N5422, N5713);
nor NOR2 (N7249, N7247, N3188);
nand NAND2 (N7250, N7243, N6782);
and AND2 (N7251, N7223, N7207);
not NOT1 (N7252, N7245);
and AND2 (N7253, N7249, N3464);
nand NAND2 (N7254, N7248, N5194);
xor XOR2 (N7255, N7241, N6338);
and AND2 (N7256, N7240, N6721);
buf BUF1 (N7257, N7256);
and AND2 (N7258, N7257, N2038);
not NOT1 (N7259, N7233);
or OR3 (N7260, N7253, N3977, N4633);
or OR3 (N7261, N7251, N3572, N2374);
nor NOR2 (N7262, N7261, N647);
not NOT1 (N7263, N7252);
and AND3 (N7264, N7250, N6094, N2619);
nand NAND3 (N7265, N7259, N488, N2576);
nor NOR4 (N7266, N7254, N7016, N3856, N59);
nor NOR4 (N7267, N7258, N2107, N2682, N1685);
and AND4 (N7268, N7260, N6653, N3252, N4770);
nor NOR3 (N7269, N7246, N2065, N2757);
not NOT1 (N7270, N7263);
nor NOR2 (N7271, N7267, N744);
xor XOR2 (N7272, N7264, N6863);
nand NAND4 (N7273, N7271, N4543, N4937, N5537);
not NOT1 (N7274, N7237);
not NOT1 (N7275, N7272);
buf BUF1 (N7276, N7262);
nor NOR2 (N7277, N7255, N5027);
xor XOR2 (N7278, N7276, N1399);
and AND4 (N7279, N7275, N3433, N3334, N5718);
xor XOR2 (N7280, N7274, N856);
or OR2 (N7281, N7280, N1302);
nor NOR2 (N7282, N7265, N5015);
nand NAND4 (N7283, N7270, N2472, N838, N5556);
and AND4 (N7284, N7282, N6205, N2842, N3141);
or OR2 (N7285, N7269, N3854);
nand NAND4 (N7286, N7281, N4482, N4892, N1445);
xor XOR2 (N7287, N7284, N2513);
and AND2 (N7288, N7278, N3207);
nor NOR3 (N7289, N7279, N3661, N2805);
and AND3 (N7290, N7266, N4403, N4416);
and AND3 (N7291, N7273, N6573, N2841);
xor XOR2 (N7292, N7288, N254);
and AND3 (N7293, N7285, N5120, N2476);
and AND2 (N7294, N7290, N6640);
nor NOR4 (N7295, N7287, N179, N2017, N3315);
buf BUF1 (N7296, N7286);
and AND2 (N7297, N7283, N6929);
and AND2 (N7298, N7291, N2269);
or OR2 (N7299, N7289, N7118);
nor NOR3 (N7300, N7299, N1823, N257);
xor XOR2 (N7301, N7296, N4612);
and AND2 (N7302, N7292, N485);
xor XOR2 (N7303, N7300, N3056);
nor NOR2 (N7304, N7293, N1927);
nor NOR3 (N7305, N7301, N956, N5339);
and AND3 (N7306, N7277, N3078, N4079);
xor XOR2 (N7307, N7302, N4886);
nor NOR3 (N7308, N7294, N2845, N6912);
nor NOR2 (N7309, N7308, N5088);
buf BUF1 (N7310, N7306);
buf BUF1 (N7311, N7304);
and AND2 (N7312, N7297, N7219);
not NOT1 (N7313, N7310);
xor XOR2 (N7314, N7311, N2289);
and AND2 (N7315, N7268, N4845);
or OR4 (N7316, N7313, N2173, N6076, N1814);
not NOT1 (N7317, N7305);
or OR3 (N7318, N7309, N5284, N6461);
nand NAND2 (N7319, N7316, N1465);
buf BUF1 (N7320, N7314);
or OR2 (N7321, N7317, N2627);
and AND3 (N7322, N7320, N6039, N2627);
and AND3 (N7323, N7318, N3340, N5012);
xor XOR2 (N7324, N7315, N6331);
not NOT1 (N7325, N7295);
or OR3 (N7326, N7298, N3503, N4658);
not NOT1 (N7327, N7321);
buf BUF1 (N7328, N7323);
not NOT1 (N7329, N7326);
buf BUF1 (N7330, N7307);
or OR4 (N7331, N7329, N2335, N4687, N6085);
nor NOR4 (N7332, N7327, N3965, N2630, N6696);
nor NOR2 (N7333, N7331, N5300);
or OR4 (N7334, N7330, N1555, N5488, N162);
buf BUF1 (N7335, N7334);
xor XOR2 (N7336, N7312, N2677);
buf BUF1 (N7337, N7328);
nor NOR3 (N7338, N7319, N4045, N6170);
or OR2 (N7339, N7322, N859);
or OR2 (N7340, N7324, N3755);
nor NOR3 (N7341, N7339, N5760, N5071);
not NOT1 (N7342, N7333);
not NOT1 (N7343, N7337);
nand NAND3 (N7344, N7335, N988, N7019);
nand NAND4 (N7345, N7344, N2890, N3285, N1132);
and AND2 (N7346, N7341, N5965);
buf BUF1 (N7347, N7338);
and AND2 (N7348, N7303, N2012);
nand NAND4 (N7349, N7325, N7204, N2006, N4173);
xor XOR2 (N7350, N7332, N6819);
not NOT1 (N7351, N7342);
or OR2 (N7352, N7347, N1575);
and AND4 (N7353, N7343, N6870, N802, N6836);
or OR3 (N7354, N7348, N2444, N6504);
xor XOR2 (N7355, N7353, N2879);
not NOT1 (N7356, N7346);
not NOT1 (N7357, N7349);
or OR4 (N7358, N7350, N1748, N7106, N5854);
and AND3 (N7359, N7356, N2252, N3934);
and AND2 (N7360, N7352, N4659);
and AND4 (N7361, N7355, N566, N4623, N871);
nor NOR3 (N7362, N7360, N4256, N4389);
nor NOR3 (N7363, N7345, N7144, N3870);
nor NOR2 (N7364, N7357, N3038);
nor NOR3 (N7365, N7351, N3374, N2819);
nor NOR4 (N7366, N7336, N7098, N2175, N307);
nor NOR2 (N7367, N7359, N3361);
or OR2 (N7368, N7363, N1515);
or OR4 (N7369, N7340, N3603, N6578, N5126);
not NOT1 (N7370, N7366);
buf BUF1 (N7371, N7367);
xor XOR2 (N7372, N7369, N2285);
not NOT1 (N7373, N7368);
buf BUF1 (N7374, N7362);
and AND4 (N7375, N7370, N1869, N4240, N3789);
or OR4 (N7376, N7354, N1660, N3465, N6422);
buf BUF1 (N7377, N7373);
xor XOR2 (N7378, N7372, N2116);
and AND4 (N7379, N7358, N462, N3125, N1289);
buf BUF1 (N7380, N7377);
buf BUF1 (N7381, N7374);
and AND3 (N7382, N7365, N4789, N5544);
not NOT1 (N7383, N7379);
buf BUF1 (N7384, N7364);
nor NOR4 (N7385, N7378, N4715, N2433, N7180);
and AND4 (N7386, N7375, N4725, N5372, N5277);
and AND2 (N7387, N7386, N353);
or OR2 (N7388, N7383, N5995);
nand NAND3 (N7389, N7376, N4055, N5892);
buf BUF1 (N7390, N7371);
buf BUF1 (N7391, N7361);
and AND4 (N7392, N7384, N2415, N7112, N4448);
or OR4 (N7393, N7381, N5095, N1140, N6113);
buf BUF1 (N7394, N7391);
not NOT1 (N7395, N7393);
not NOT1 (N7396, N7395);
xor XOR2 (N7397, N7394, N1417);
not NOT1 (N7398, N7390);
nand NAND2 (N7399, N7385, N1430);
or OR2 (N7400, N7399, N1037);
and AND2 (N7401, N7388, N1035);
nand NAND4 (N7402, N7397, N4547, N3807, N4645);
or OR2 (N7403, N7389, N95);
xor XOR2 (N7404, N7396, N1728);
or OR3 (N7405, N7382, N6968, N6765);
nand NAND3 (N7406, N7402, N108, N2226);
or OR2 (N7407, N7387, N2029);
and AND3 (N7408, N7406, N1409, N4449);
and AND2 (N7409, N7403, N3070);
nand NAND2 (N7410, N7392, N3632);
buf BUF1 (N7411, N7407);
and AND2 (N7412, N7410, N892);
buf BUF1 (N7413, N7398);
nand NAND4 (N7414, N7411, N5073, N6501, N7267);
or OR3 (N7415, N7405, N6971, N860);
nor NOR4 (N7416, N7415, N3333, N1946, N718);
buf BUF1 (N7417, N7400);
and AND4 (N7418, N7409, N5613, N5980, N3000);
nor NOR2 (N7419, N7412, N5493);
or OR2 (N7420, N7404, N6205);
and AND4 (N7421, N7401, N6642, N7205, N6001);
not NOT1 (N7422, N7414);
buf BUF1 (N7423, N7408);
not NOT1 (N7424, N7416);
and AND4 (N7425, N7380, N4954, N3669, N2458);
not NOT1 (N7426, N7422);
and AND2 (N7427, N7418, N4957);
buf BUF1 (N7428, N7419);
xor XOR2 (N7429, N7423, N6251);
nand NAND2 (N7430, N7417, N5600);
or OR4 (N7431, N7430, N4477, N1459, N6453);
and AND3 (N7432, N7429, N4993, N2690);
nor NOR2 (N7433, N7431, N5586);
buf BUF1 (N7434, N7413);
nor NOR2 (N7435, N7434, N101);
xor XOR2 (N7436, N7433, N411);
not NOT1 (N7437, N7426);
not NOT1 (N7438, N7425);
and AND2 (N7439, N7420, N6758);
nor NOR2 (N7440, N7439, N3469);
or OR4 (N7441, N7421, N1215, N868, N6952);
nand NAND4 (N7442, N7428, N1198, N7420, N6204);
xor XOR2 (N7443, N7440, N2009);
nor NOR3 (N7444, N7437, N5414, N7331);
xor XOR2 (N7445, N7442, N1369);
xor XOR2 (N7446, N7445, N6628);
xor XOR2 (N7447, N7444, N4207);
buf BUF1 (N7448, N7435);
xor XOR2 (N7449, N7424, N1299);
or OR4 (N7450, N7443, N4135, N3753, N974);
nor NOR3 (N7451, N7446, N6726, N6283);
and AND3 (N7452, N7441, N942, N716);
and AND4 (N7453, N7450, N5886, N524, N6261);
and AND2 (N7454, N7447, N6528);
nand NAND2 (N7455, N7453, N6767);
and AND2 (N7456, N7436, N5921);
nand NAND4 (N7457, N7451, N2531, N1833, N2057);
buf BUF1 (N7458, N7432);
or OR4 (N7459, N7458, N2160, N6892, N5222);
buf BUF1 (N7460, N7457);
nor NOR4 (N7461, N7460, N7438, N4680, N2668);
nand NAND4 (N7462, N3587, N2572, N1866, N6405);
nor NOR2 (N7463, N7456, N7441);
nor NOR3 (N7464, N7449, N5502, N3286);
or OR2 (N7465, N7427, N1615);
buf BUF1 (N7466, N7464);
and AND4 (N7467, N7448, N206, N2809, N620);
or OR4 (N7468, N7467, N3869, N1986, N1055);
nand NAND2 (N7469, N7466, N1215);
and AND3 (N7470, N7459, N5649, N1903);
or OR2 (N7471, N7465, N7);
nor NOR3 (N7472, N7461, N6950, N7040);
nand NAND3 (N7473, N7452, N7328, N5140);
or OR2 (N7474, N7468, N3992);
nor NOR3 (N7475, N7463, N3077, N7284);
not NOT1 (N7476, N7473);
and AND2 (N7477, N7469, N7263);
not NOT1 (N7478, N7470);
xor XOR2 (N7479, N7478, N4231);
nor NOR4 (N7480, N7477, N862, N6572, N3767);
buf BUF1 (N7481, N7462);
buf BUF1 (N7482, N7480);
xor XOR2 (N7483, N7481, N4746);
nor NOR3 (N7484, N7479, N5856, N140);
and AND3 (N7485, N7475, N3402, N792);
nor NOR2 (N7486, N7484, N721);
or OR3 (N7487, N7472, N1426, N13);
not NOT1 (N7488, N7476);
xor XOR2 (N7489, N7454, N2789);
or OR3 (N7490, N7487, N490, N2867);
nor NOR3 (N7491, N7488, N583, N2755);
or OR3 (N7492, N7486, N3155, N735);
buf BUF1 (N7493, N7491);
buf BUF1 (N7494, N7489);
not NOT1 (N7495, N7471);
nand NAND4 (N7496, N7455, N7276, N4525, N7492);
and AND3 (N7497, N5784, N2125, N3035);
xor XOR2 (N7498, N7496, N3352);
nand NAND3 (N7499, N7485, N6134, N3992);
nor NOR2 (N7500, N7494, N1214);
buf BUF1 (N7501, N7500);
buf BUF1 (N7502, N7493);
nand NAND3 (N7503, N7474, N6646, N6587);
buf BUF1 (N7504, N7490);
or OR2 (N7505, N7495, N5461);
nor NOR4 (N7506, N7497, N5308, N1493, N5589);
xor XOR2 (N7507, N7505, N7017);
or OR2 (N7508, N7483, N3710);
and AND2 (N7509, N7508, N714);
nor NOR2 (N7510, N7509, N6151);
xor XOR2 (N7511, N7501, N6269);
and AND4 (N7512, N7504, N5326, N2847, N5742);
nor NOR3 (N7513, N7482, N4939, N6009);
not NOT1 (N7514, N7507);
and AND2 (N7515, N7499, N5826);
buf BUF1 (N7516, N7515);
buf BUF1 (N7517, N7503);
nor NOR2 (N7518, N7506, N4583);
nand NAND3 (N7519, N7512, N5914, N2530);
nor NOR2 (N7520, N7516, N2386);
not NOT1 (N7521, N7498);
and AND2 (N7522, N7514, N68);
and AND3 (N7523, N7521, N2105, N195);
nand NAND4 (N7524, N7502, N6037, N6209, N4268);
nor NOR2 (N7525, N7520, N5170);
not NOT1 (N7526, N7519);
not NOT1 (N7527, N7517);
not NOT1 (N7528, N7518);
nand NAND3 (N7529, N7523, N5553, N1450);
not NOT1 (N7530, N7526);
and AND2 (N7531, N7525, N4127);
not NOT1 (N7532, N7531);
and AND2 (N7533, N7511, N6261);
nand NAND3 (N7534, N7533, N4854, N4408);
and AND2 (N7535, N7532, N1944);
and AND4 (N7536, N7510, N5441, N3506, N1028);
nand NAND4 (N7537, N7527, N2000, N782, N708);
nor NOR4 (N7538, N7513, N2902, N6723, N474);
xor XOR2 (N7539, N7529, N2958);
buf BUF1 (N7540, N7538);
and AND2 (N7541, N7534, N5038);
xor XOR2 (N7542, N7522, N4472);
and AND2 (N7543, N7535, N6553);
and AND4 (N7544, N7530, N3018, N2041, N5762);
xor XOR2 (N7545, N7541, N2090);
or OR2 (N7546, N7543, N2300);
xor XOR2 (N7547, N7545, N5847);
xor XOR2 (N7548, N7524, N4137);
buf BUF1 (N7549, N7547);
buf BUF1 (N7550, N7549);
xor XOR2 (N7551, N7528, N6477);
not NOT1 (N7552, N7550);
and AND3 (N7553, N7542, N497, N2881);
buf BUF1 (N7554, N7544);
and AND2 (N7555, N7537, N5559);
nand NAND3 (N7556, N7546, N6831, N5042);
xor XOR2 (N7557, N7556, N5439);
nor NOR2 (N7558, N7554, N1973);
or OR3 (N7559, N7536, N6501, N154);
and AND2 (N7560, N7551, N1563);
not NOT1 (N7561, N7555);
buf BUF1 (N7562, N7560);
xor XOR2 (N7563, N7548, N1663);
nand NAND2 (N7564, N7562, N2119);
xor XOR2 (N7565, N7539, N450);
or OR3 (N7566, N7565, N4907, N711);
nor NOR3 (N7567, N7558, N6272, N1378);
buf BUF1 (N7568, N7561);
nor NOR4 (N7569, N7552, N7217, N5720, N4265);
nand NAND2 (N7570, N7540, N4510);
nor NOR4 (N7571, N7566, N4962, N4436, N853);
nand NAND2 (N7572, N7557, N7457);
and AND4 (N7573, N7564, N3207, N18, N606);
not NOT1 (N7574, N7573);
xor XOR2 (N7575, N7568, N6159);
and AND3 (N7576, N7563, N4195, N1140);
or OR4 (N7577, N7569, N6782, N2326, N82);
and AND3 (N7578, N7570, N421, N4200);
buf BUF1 (N7579, N7567);
nor NOR3 (N7580, N7559, N6955, N2287);
not NOT1 (N7581, N7571);
buf BUF1 (N7582, N7553);
buf BUF1 (N7583, N7578);
or OR4 (N7584, N7580, N5250, N511, N6812);
nand NAND2 (N7585, N7579, N1638);
or OR4 (N7586, N7582, N4398, N5594, N2636);
buf BUF1 (N7587, N7583);
nor NOR3 (N7588, N7585, N1035, N4744);
nor NOR4 (N7589, N7575, N2714, N7312, N7565);
nand NAND3 (N7590, N7574, N1344, N1570);
not NOT1 (N7591, N7584);
not NOT1 (N7592, N7588);
xor XOR2 (N7593, N7576, N218);
not NOT1 (N7594, N7577);
nor NOR2 (N7595, N7586, N5430);
buf BUF1 (N7596, N7593);
xor XOR2 (N7597, N7587, N2891);
nor NOR2 (N7598, N7591, N4786);
buf BUF1 (N7599, N7597);
or OR2 (N7600, N7596, N6056);
or OR2 (N7601, N7600, N3127);
not NOT1 (N7602, N7594);
not NOT1 (N7603, N7589);
nor NOR2 (N7604, N7590, N4187);
xor XOR2 (N7605, N7598, N7256);
or OR3 (N7606, N7599, N640, N4761);
and AND3 (N7607, N7592, N279, N6264);
nor NOR3 (N7608, N7581, N5273, N5318);
or OR2 (N7609, N7608, N5151);
or OR3 (N7610, N7605, N5003, N2024);
or OR3 (N7611, N7595, N3659, N621);
and AND2 (N7612, N7606, N3445);
and AND4 (N7613, N7610, N665, N931, N1482);
xor XOR2 (N7614, N7572, N1190);
not NOT1 (N7615, N7614);
xor XOR2 (N7616, N7603, N616);
xor XOR2 (N7617, N7604, N1749);
nand NAND2 (N7618, N7609, N2642);
buf BUF1 (N7619, N7612);
nand NAND2 (N7620, N7613, N5701);
buf BUF1 (N7621, N7601);
nand NAND4 (N7622, N7617, N2833, N6949, N1765);
not NOT1 (N7623, N7602);
or OR4 (N7624, N7607, N4393, N2431, N5194);
not NOT1 (N7625, N7622);
not NOT1 (N7626, N7611);
nor NOR3 (N7627, N7615, N2202, N747);
nand NAND4 (N7628, N7621, N5087, N6285, N457);
nor NOR3 (N7629, N7623, N2702, N764);
buf BUF1 (N7630, N7627);
or OR4 (N7631, N7625, N3520, N540, N3848);
xor XOR2 (N7632, N7620, N4184);
nor NOR3 (N7633, N7618, N6375, N4536);
nor NOR4 (N7634, N7626, N3810, N1818, N3470);
buf BUF1 (N7635, N7619);
and AND3 (N7636, N7628, N5628, N1693);
xor XOR2 (N7637, N7629, N1916);
xor XOR2 (N7638, N7631, N2504);
and AND2 (N7639, N7616, N2959);
not NOT1 (N7640, N7637);
or OR4 (N7641, N7639, N5476, N631, N777);
nor NOR3 (N7642, N7630, N747, N3871);
nor NOR2 (N7643, N7632, N2903);
or OR2 (N7644, N7641, N5631);
buf BUF1 (N7645, N7638);
or OR3 (N7646, N7640, N4678, N3417);
nand NAND3 (N7647, N7634, N3099, N6836);
buf BUF1 (N7648, N7647);
xor XOR2 (N7649, N7643, N5599);
xor XOR2 (N7650, N7648, N2404);
and AND2 (N7651, N7649, N2579);
nor NOR2 (N7652, N7642, N2766);
nand NAND3 (N7653, N7646, N3402, N7523);
buf BUF1 (N7654, N7651);
xor XOR2 (N7655, N7636, N6775);
nor NOR2 (N7656, N7635, N531);
not NOT1 (N7657, N7656);
and AND2 (N7658, N7653, N790);
xor XOR2 (N7659, N7633, N5147);
nand NAND2 (N7660, N7657, N4278);
not NOT1 (N7661, N7655);
buf BUF1 (N7662, N7654);
not NOT1 (N7663, N7661);
or OR3 (N7664, N7645, N41, N5615);
nand NAND2 (N7665, N7664, N4952);
xor XOR2 (N7666, N7624, N6227);
not NOT1 (N7667, N7663);
or OR2 (N7668, N7665, N2125);
xor XOR2 (N7669, N7658, N3405);
not NOT1 (N7670, N7662);
xor XOR2 (N7671, N7666, N3793);
nor NOR4 (N7672, N7660, N5963, N2916, N5921);
not NOT1 (N7673, N7659);
xor XOR2 (N7674, N7668, N5235);
and AND4 (N7675, N7652, N6461, N4251, N731);
and AND4 (N7676, N7673, N5635, N4921, N1907);
nand NAND2 (N7677, N7669, N4962);
nor NOR4 (N7678, N7677, N314, N3366, N2711);
and AND4 (N7679, N7672, N4469, N4150, N681);
nand NAND3 (N7680, N7644, N3046, N1686);
not NOT1 (N7681, N7676);
and AND4 (N7682, N7680, N1804, N4788, N713);
xor XOR2 (N7683, N7682, N603);
not NOT1 (N7684, N7674);
not NOT1 (N7685, N7667);
not NOT1 (N7686, N7681);
nor NOR2 (N7687, N7675, N4710);
or OR2 (N7688, N7683, N1955);
not NOT1 (N7689, N7687);
nand NAND3 (N7690, N7650, N679, N301);
xor XOR2 (N7691, N7671, N2019);
and AND4 (N7692, N7688, N5265, N6842, N3419);
nand NAND2 (N7693, N7685, N893);
nor NOR4 (N7694, N7689, N4889, N5911, N5862);
buf BUF1 (N7695, N7693);
not NOT1 (N7696, N7691);
xor XOR2 (N7697, N7694, N1148);
buf BUF1 (N7698, N7695);
and AND2 (N7699, N7679, N6559);
nand NAND3 (N7700, N7697, N2113, N606);
and AND3 (N7701, N7684, N6849, N311);
xor XOR2 (N7702, N7698, N3184);
buf BUF1 (N7703, N7678);
not NOT1 (N7704, N7702);
buf BUF1 (N7705, N7700);
not NOT1 (N7706, N7686);
not NOT1 (N7707, N7692);
not NOT1 (N7708, N7701);
not NOT1 (N7709, N7696);
not NOT1 (N7710, N7699);
or OR3 (N7711, N7705, N1082, N5521);
xor XOR2 (N7712, N7709, N3358);
buf BUF1 (N7713, N7670);
and AND4 (N7714, N7706, N686, N748, N3130);
or OR4 (N7715, N7703, N6427, N6178, N6860);
and AND4 (N7716, N7704, N1787, N4919, N1148);
not NOT1 (N7717, N7712);
nand NAND4 (N7718, N7708, N3050, N4812, N4278);
xor XOR2 (N7719, N7711, N408);
nand NAND4 (N7720, N7710, N636, N4972, N4636);
nand NAND4 (N7721, N7717, N7659, N6718, N3920);
buf BUF1 (N7722, N7716);
or OR4 (N7723, N7713, N2444, N5757, N7638);
not NOT1 (N7724, N7715);
or OR3 (N7725, N7720, N6296, N5803);
not NOT1 (N7726, N7725);
nand NAND2 (N7727, N7726, N6016);
and AND4 (N7728, N7719, N4575, N6255, N4291);
nor NOR2 (N7729, N7728, N1390);
xor XOR2 (N7730, N7727, N5233);
xor XOR2 (N7731, N7730, N3702);
buf BUF1 (N7732, N7718);
nand NAND4 (N7733, N7724, N7292, N5546, N1534);
buf BUF1 (N7734, N7731);
nor NOR2 (N7735, N7722, N4523);
buf BUF1 (N7736, N7734);
and AND4 (N7737, N7733, N6159, N2932, N881);
and AND3 (N7738, N7732, N5499, N1180);
xor XOR2 (N7739, N7735, N5357);
nand NAND2 (N7740, N7707, N181);
xor XOR2 (N7741, N7740, N3889);
or OR2 (N7742, N7737, N3055);
nor NOR3 (N7743, N7739, N4085, N119);
or OR2 (N7744, N7741, N338);
nand NAND3 (N7745, N7729, N5510, N2050);
not NOT1 (N7746, N7721);
and AND4 (N7747, N7746, N7388, N345, N4782);
or OR3 (N7748, N7742, N1148, N4297);
buf BUF1 (N7749, N7736);
nor NOR4 (N7750, N7738, N1163, N634, N6366);
not NOT1 (N7751, N7690);
buf BUF1 (N7752, N7749);
or OR3 (N7753, N7747, N4743, N7067);
nand NAND3 (N7754, N7743, N6380, N2912);
nor NOR4 (N7755, N7753, N2401, N5470, N899);
and AND3 (N7756, N7714, N174, N5926);
and AND2 (N7757, N7748, N7699);
xor XOR2 (N7758, N7756, N401);
or OR3 (N7759, N7754, N103, N6027);
or OR3 (N7760, N7759, N3288, N3423);
nand NAND3 (N7761, N7751, N2310, N5984);
nor NOR3 (N7762, N7760, N6248, N4710);
buf BUF1 (N7763, N7758);
buf BUF1 (N7764, N7763);
and AND3 (N7765, N7755, N1620, N6821);
and AND3 (N7766, N7765, N1939, N1969);
and AND2 (N7767, N7764, N3952);
not NOT1 (N7768, N7752);
nand NAND2 (N7769, N7723, N6218);
and AND2 (N7770, N7757, N4645);
and AND3 (N7771, N7761, N461, N855);
nor NOR2 (N7772, N7750, N7446);
nor NOR3 (N7773, N7744, N2560, N2975);
or OR2 (N7774, N7766, N3524);
not NOT1 (N7775, N7774);
nand NAND4 (N7776, N7769, N5233, N4652, N5583);
nand NAND4 (N7777, N7772, N112, N4376, N478);
or OR3 (N7778, N7773, N566, N963);
and AND3 (N7779, N7776, N2552, N851);
xor XOR2 (N7780, N7745, N925);
buf BUF1 (N7781, N7780);
or OR3 (N7782, N7779, N1197, N2021);
not NOT1 (N7783, N7762);
nor NOR2 (N7784, N7767, N5670);
nor NOR4 (N7785, N7771, N2075, N2253, N3716);
buf BUF1 (N7786, N7782);
buf BUF1 (N7787, N7770);
nand NAND4 (N7788, N7775, N4572, N2549, N216);
not NOT1 (N7789, N7777);
or OR2 (N7790, N7787, N1308);
not NOT1 (N7791, N7790);
nand NAND3 (N7792, N7791, N2995, N4329);
buf BUF1 (N7793, N7784);
nand NAND2 (N7794, N7788, N2779);
buf BUF1 (N7795, N7783);
and AND4 (N7796, N7785, N761, N581, N763);
nor NOR2 (N7797, N7794, N6067);
nand NAND4 (N7798, N7795, N6262, N6729, N4666);
xor XOR2 (N7799, N7781, N1337);
or OR2 (N7800, N7793, N3792);
nand NAND2 (N7801, N7792, N1035);
or OR3 (N7802, N7800, N6154, N5371);
nor NOR3 (N7803, N7797, N7261, N6701);
not NOT1 (N7804, N7789);
not NOT1 (N7805, N7799);
not NOT1 (N7806, N7804);
nor NOR4 (N7807, N7778, N2428, N4545, N1320);
xor XOR2 (N7808, N7805, N1229);
nand NAND3 (N7809, N7803, N860, N6867);
buf BUF1 (N7810, N7768);
buf BUF1 (N7811, N7807);
or OR3 (N7812, N7798, N3118, N6440);
not NOT1 (N7813, N7796);
or OR4 (N7814, N7813, N391, N5271, N949);
xor XOR2 (N7815, N7810, N6869);
nor NOR3 (N7816, N7786, N6702, N87);
xor XOR2 (N7817, N7814, N2838);
or OR2 (N7818, N7809, N251);
not NOT1 (N7819, N7808);
nor NOR2 (N7820, N7811, N5052);
and AND3 (N7821, N7801, N5667, N1511);
xor XOR2 (N7822, N7815, N3735);
not NOT1 (N7823, N7816);
nor NOR4 (N7824, N7818, N2341, N3238, N3050);
xor XOR2 (N7825, N7806, N3073);
nor NOR4 (N7826, N7802, N981, N96, N3879);
and AND2 (N7827, N7812, N4819);
and AND4 (N7828, N7827, N7686, N2613, N3632);
not NOT1 (N7829, N7820);
xor XOR2 (N7830, N7823, N2703);
nand NAND2 (N7831, N7819, N5079);
nand NAND2 (N7832, N7828, N7198);
nor NOR2 (N7833, N7825, N3439);
nor NOR2 (N7834, N7824, N5610);
xor XOR2 (N7835, N7826, N2105);
not NOT1 (N7836, N7830);
not NOT1 (N7837, N7817);
xor XOR2 (N7838, N7833, N858);
xor XOR2 (N7839, N7838, N40);
nand NAND2 (N7840, N7837, N6561);
nor NOR3 (N7841, N7839, N581, N2397);
or OR2 (N7842, N7829, N1398);
buf BUF1 (N7843, N7821);
nand NAND3 (N7844, N7822, N5678, N7039);
buf BUF1 (N7845, N7835);
not NOT1 (N7846, N7834);
nor NOR2 (N7847, N7840, N6354);
xor XOR2 (N7848, N7843, N688);
nand NAND4 (N7849, N7831, N1147, N3104, N3059);
not NOT1 (N7850, N7845);
nand NAND4 (N7851, N7849, N5117, N3486, N1794);
buf BUF1 (N7852, N7848);
nor NOR3 (N7853, N7847, N5284, N1727);
and AND2 (N7854, N7850, N3413);
not NOT1 (N7855, N7836);
xor XOR2 (N7856, N7853, N2686);
or OR2 (N7857, N7854, N4909);
or OR2 (N7858, N7856, N5019);
nand NAND2 (N7859, N7852, N3587);
xor XOR2 (N7860, N7855, N3698);
and AND2 (N7861, N7858, N1019);
nand NAND3 (N7862, N7842, N7290, N5548);
not NOT1 (N7863, N7859);
buf BUF1 (N7864, N7844);
nand NAND2 (N7865, N7861, N1915);
and AND3 (N7866, N7863, N5000, N7817);
or OR2 (N7867, N7866, N5186);
or OR3 (N7868, N7864, N7302, N2681);
xor XOR2 (N7869, N7867, N3069);
and AND4 (N7870, N7841, N908, N2208, N1730);
or OR3 (N7871, N7870, N3999, N5617);
buf BUF1 (N7872, N7851);
xor XOR2 (N7873, N7860, N6968);
and AND3 (N7874, N7857, N6702, N3193);
or OR2 (N7875, N7872, N6944);
not NOT1 (N7876, N7869);
nand NAND4 (N7877, N7874, N2377, N987, N2223);
and AND4 (N7878, N7873, N3115, N4708, N4706);
nor NOR3 (N7879, N7862, N3812, N3223);
nand NAND3 (N7880, N7878, N6902, N3949);
not NOT1 (N7881, N7876);
nand NAND4 (N7882, N7881, N9, N5993, N7125);
not NOT1 (N7883, N7875);
and AND4 (N7884, N7879, N3256, N3251, N1836);
buf BUF1 (N7885, N7846);
xor XOR2 (N7886, N7880, N2780);
or OR2 (N7887, N7877, N865);
xor XOR2 (N7888, N7884, N4924);
buf BUF1 (N7889, N7832);
not NOT1 (N7890, N7887);
nor NOR4 (N7891, N7868, N4066, N565, N3628);
buf BUF1 (N7892, N7882);
nand NAND3 (N7893, N7883, N6465, N2353);
not NOT1 (N7894, N7891);
nand NAND2 (N7895, N7871, N4947);
and AND2 (N7896, N7893, N55);
not NOT1 (N7897, N7896);
or OR3 (N7898, N7885, N3912, N3252);
or OR2 (N7899, N7886, N1824);
nor NOR3 (N7900, N7889, N456, N2722);
nor NOR2 (N7901, N7892, N169);
not NOT1 (N7902, N7901);
nor NOR4 (N7903, N7894, N7881, N7760, N3396);
buf BUF1 (N7904, N7897);
xor XOR2 (N7905, N7902, N5251);
nor NOR4 (N7906, N7899, N6929, N1377, N7905);
nor NOR3 (N7907, N2955, N5276, N5922);
or OR3 (N7908, N7888, N5732, N226);
nor NOR2 (N7909, N7907, N7212);
buf BUF1 (N7910, N7909);
not NOT1 (N7911, N7908);
or OR4 (N7912, N7895, N2897, N3411, N5230);
buf BUF1 (N7913, N7865);
nor NOR3 (N7914, N7898, N2345, N4105);
or OR2 (N7915, N7904, N4492);
nor NOR3 (N7916, N7915, N4564, N2876);
xor XOR2 (N7917, N7913, N4787);
and AND4 (N7918, N7917, N3267, N5859, N7015);
nor NOR2 (N7919, N7910, N2790);
xor XOR2 (N7920, N7911, N3173);
not NOT1 (N7921, N7918);
nor NOR3 (N7922, N7906, N5183, N5077);
or OR2 (N7923, N7916, N6214);
nor NOR2 (N7924, N7920, N587);
nor NOR4 (N7925, N7923, N7652, N4643, N7487);
not NOT1 (N7926, N7924);
buf BUF1 (N7927, N7914);
nand NAND4 (N7928, N7890, N2222, N6776, N7275);
not NOT1 (N7929, N7926);
and AND2 (N7930, N7929, N4740);
not NOT1 (N7931, N7928);
xor XOR2 (N7932, N7903, N6293);
xor XOR2 (N7933, N7925, N6135);
buf BUF1 (N7934, N7931);
buf BUF1 (N7935, N7900);
and AND2 (N7936, N7912, N3508);
nand NAND3 (N7937, N7933, N7145, N3859);
nor NOR2 (N7938, N7936, N5963);
xor XOR2 (N7939, N7930, N1142);
or OR3 (N7940, N7939, N392, N7329);
nand NAND4 (N7941, N7934, N4371, N337, N3348);
or OR4 (N7942, N7932, N4748, N6647, N524);
not NOT1 (N7943, N7935);
and AND4 (N7944, N7927, N6442, N1982, N3669);
and AND2 (N7945, N7922, N589);
nand NAND4 (N7946, N7938, N4278, N8, N3289);
nand NAND3 (N7947, N7937, N6656, N6849);
not NOT1 (N7948, N7921);
and AND2 (N7949, N7942, N3004);
or OR4 (N7950, N7941, N5300, N6353, N3447);
buf BUF1 (N7951, N7943);
not NOT1 (N7952, N7948);
not NOT1 (N7953, N7950);
nand NAND2 (N7954, N7949, N1470);
and AND2 (N7955, N7919, N1097);
nor NOR2 (N7956, N7945, N4373);
nand NAND3 (N7957, N7955, N6212, N4941);
nor NOR4 (N7958, N7944, N445, N3180, N3786);
not NOT1 (N7959, N7951);
or OR3 (N7960, N7957, N3355, N5357);
and AND2 (N7961, N7947, N2548);
or OR3 (N7962, N7960, N1766, N5151);
or OR3 (N7963, N7954, N4132, N6199);
buf BUF1 (N7964, N7958);
xor XOR2 (N7965, N7946, N2795);
and AND2 (N7966, N7956, N6077);
nor NOR3 (N7967, N7953, N4387, N3154);
nor NOR4 (N7968, N7961, N7708, N2957, N4465);
not NOT1 (N7969, N7963);
and AND2 (N7970, N7965, N6760);
nor NOR3 (N7971, N7968, N5256, N4453);
not NOT1 (N7972, N7967);
or OR4 (N7973, N7964, N1893, N7675, N4886);
nor NOR3 (N7974, N7971, N7799, N4173);
not NOT1 (N7975, N7972);
and AND3 (N7976, N7973, N2884, N4362);
buf BUF1 (N7977, N7975);
nand NAND2 (N7978, N7977, N6584);
not NOT1 (N7979, N7976);
buf BUF1 (N7980, N7959);
and AND3 (N7981, N7974, N7654, N5143);
buf BUF1 (N7982, N7979);
nor NOR2 (N7983, N7982, N1436);
nand NAND2 (N7984, N7981, N6831);
nand NAND2 (N7985, N7952, N1752);
and AND3 (N7986, N7983, N4760, N1878);
or OR3 (N7987, N7966, N5723, N884);
not NOT1 (N7988, N7984);
and AND2 (N7989, N7978, N6140);
nand NAND2 (N7990, N7986, N6010);
buf BUF1 (N7991, N7962);
and AND3 (N7992, N7987, N3321, N5339);
nand NAND2 (N7993, N7992, N475);
and AND4 (N7994, N7970, N5004, N5827, N202);
nand NAND3 (N7995, N7940, N6150, N1899);
xor XOR2 (N7996, N7990, N1575);
nor NOR4 (N7997, N7989, N5587, N7861, N668);
xor XOR2 (N7998, N7993, N5146);
and AND4 (N7999, N7991, N4652, N5414, N3465);
buf BUF1 (N8000, N7980);
buf BUF1 (N8001, N7996);
and AND4 (N8002, N7995, N5014, N2404, N2009);
nor NOR2 (N8003, N7998, N4354);
and AND4 (N8004, N7999, N7679, N4928, N6993);
nor NOR3 (N8005, N8004, N7765, N5085);
nand NAND3 (N8006, N8000, N2741, N7974);
buf BUF1 (N8007, N8006);
nor NOR3 (N8008, N8003, N3870, N4727);
not NOT1 (N8009, N8008);
not NOT1 (N8010, N7985);
nand NAND4 (N8011, N8007, N659, N6729, N5958);
or OR2 (N8012, N8002, N3991);
nand NAND3 (N8013, N7969, N4660, N3777);
and AND4 (N8014, N8013, N3256, N7278, N5888);
and AND3 (N8015, N7997, N4759, N6597);
nor NOR2 (N8016, N8015, N2389);
or OR4 (N8017, N8001, N6413, N167, N848);
and AND2 (N8018, N8005, N1790);
buf BUF1 (N8019, N8011);
or OR3 (N8020, N8016, N7844, N1242);
or OR4 (N8021, N8009, N4522, N4069, N7381);
nand NAND3 (N8022, N8010, N626, N7352);
nand NAND4 (N8023, N8018, N7910, N2633, N4878);
nor NOR3 (N8024, N7988, N6876, N2578);
and AND2 (N8025, N8017, N753);
or OR2 (N8026, N8022, N1058);
or OR4 (N8027, N8023, N3520, N3072, N84);
and AND3 (N8028, N8025, N6233, N3210);
or OR4 (N8029, N8014, N5657, N1169, N3390);
buf BUF1 (N8030, N8027);
buf BUF1 (N8031, N8029);
xor XOR2 (N8032, N8020, N2726);
and AND3 (N8033, N8026, N7652, N6065);
xor XOR2 (N8034, N8028, N3814);
buf BUF1 (N8035, N8019);
xor XOR2 (N8036, N8035, N3518);
not NOT1 (N8037, N8030);
xor XOR2 (N8038, N8034, N2919);
and AND4 (N8039, N8024, N6892, N7883, N3034);
buf BUF1 (N8040, N7994);
or OR4 (N8041, N8012, N1862, N5809, N1850);
nor NOR2 (N8042, N8041, N7369);
buf BUF1 (N8043, N8036);
xor XOR2 (N8044, N8038, N2270);
buf BUF1 (N8045, N8037);
and AND4 (N8046, N8032, N5297, N490, N4235);
xor XOR2 (N8047, N8046, N398);
nor NOR3 (N8048, N8043, N373, N4044);
buf BUF1 (N8049, N8031);
buf BUF1 (N8050, N8021);
buf BUF1 (N8051, N8042);
not NOT1 (N8052, N8044);
nor NOR4 (N8053, N8040, N5109, N3686, N6312);
nand NAND2 (N8054, N8049, N2967);
or OR2 (N8055, N8052, N4787);
or OR3 (N8056, N8048, N1539, N6073);
buf BUF1 (N8057, N8050);
nor NOR2 (N8058, N8047, N7217);
xor XOR2 (N8059, N8039, N2179);
not NOT1 (N8060, N8054);
nor NOR2 (N8061, N8059, N7362);
or OR4 (N8062, N8055, N3631, N7981, N1652);
buf BUF1 (N8063, N8061);
buf BUF1 (N8064, N8051);
nor NOR3 (N8065, N8045, N394, N5479);
not NOT1 (N8066, N8053);
not NOT1 (N8067, N8063);
xor XOR2 (N8068, N8067, N4482);
and AND4 (N8069, N8066, N7979, N4763, N1173);
nor NOR3 (N8070, N8068, N4918, N5974);
nor NOR2 (N8071, N8033, N337);
nor NOR2 (N8072, N8064, N6700);
buf BUF1 (N8073, N8071);
buf BUF1 (N8074, N8060);
xor XOR2 (N8075, N8062, N2682);
nand NAND3 (N8076, N8070, N4627, N1355);
or OR2 (N8077, N8058, N632);
xor XOR2 (N8078, N8077, N7679);
and AND2 (N8079, N8074, N4406);
nand NAND4 (N8080, N8069, N2880, N3861, N651);
not NOT1 (N8081, N8078);
nor NOR2 (N8082, N8076, N7033);
nor NOR2 (N8083, N8073, N3758);
xor XOR2 (N8084, N8082, N5981);
buf BUF1 (N8085, N8079);
not NOT1 (N8086, N8075);
xor XOR2 (N8087, N8056, N523);
nand NAND3 (N8088, N8083, N4965, N4288);
or OR2 (N8089, N8057, N7384);
xor XOR2 (N8090, N8065, N7251);
xor XOR2 (N8091, N8085, N7125);
nand NAND2 (N8092, N8088, N5176);
buf BUF1 (N8093, N8080);
or OR2 (N8094, N8086, N221);
not NOT1 (N8095, N8091);
and AND3 (N8096, N8089, N4982, N4661);
xor XOR2 (N8097, N8096, N622);
xor XOR2 (N8098, N8084, N2617);
and AND2 (N8099, N8095, N2050);
xor XOR2 (N8100, N8093, N1090);
not NOT1 (N8101, N8087);
buf BUF1 (N8102, N8081);
xor XOR2 (N8103, N8092, N5990);
nand NAND4 (N8104, N8102, N939, N6715, N5968);
or OR3 (N8105, N8103, N4769, N4478);
xor XOR2 (N8106, N8072, N5619);
and AND2 (N8107, N8099, N1315);
or OR3 (N8108, N8105, N7902, N6890);
or OR4 (N8109, N8106, N2859, N5214, N4813);
nand NAND3 (N8110, N8109, N193, N5397);
nand NAND2 (N8111, N8104, N280);
nand NAND3 (N8112, N8107, N2050, N3487);
not NOT1 (N8113, N8098);
and AND2 (N8114, N8108, N3191);
nor NOR4 (N8115, N8111, N4649, N7538, N3804);
or OR3 (N8116, N8112, N918, N7571);
xor XOR2 (N8117, N8114, N7676);
and AND4 (N8118, N8100, N2244, N3971, N7854);
and AND3 (N8119, N8118, N1937, N3598);
buf BUF1 (N8120, N8101);
xor XOR2 (N8121, N8117, N3724);
not NOT1 (N8122, N8094);
nor NOR3 (N8123, N8116, N6193, N5127);
nor NOR2 (N8124, N8120, N4556);
not NOT1 (N8125, N8090);
xor XOR2 (N8126, N8121, N4537);
nor NOR2 (N8127, N8113, N6868);
xor XOR2 (N8128, N8119, N653);
not NOT1 (N8129, N8097);
nor NOR3 (N8130, N8122, N1901, N3153);
buf BUF1 (N8131, N8129);
nor NOR3 (N8132, N8131, N5793, N3935);
buf BUF1 (N8133, N8126);
not NOT1 (N8134, N8128);
or OR4 (N8135, N8125, N1229, N6606, N6180);
and AND2 (N8136, N8115, N3657);
xor XOR2 (N8137, N8135, N4458);
nor NOR2 (N8138, N8132, N895);
or OR4 (N8139, N8110, N5106, N7036, N5006);
nand NAND2 (N8140, N8138, N1730);
nor NOR4 (N8141, N8136, N4785, N3192, N657);
buf BUF1 (N8142, N8139);
and AND3 (N8143, N8141, N1535, N7460);
and AND3 (N8144, N8143, N779, N6764);
nor NOR2 (N8145, N8140, N5660);
and AND4 (N8146, N8145, N1954, N6168, N55);
or OR3 (N8147, N8142, N1967, N6559);
not NOT1 (N8148, N8146);
or OR2 (N8149, N8124, N5702);
nor NOR2 (N8150, N8127, N7527);
or OR2 (N8151, N8133, N5288);
not NOT1 (N8152, N8149);
nand NAND3 (N8153, N8123, N6939, N7857);
nor NOR4 (N8154, N8153, N2344, N7138, N6999);
and AND4 (N8155, N8130, N97, N1232, N2429);
buf BUF1 (N8156, N8154);
buf BUF1 (N8157, N8151);
nand NAND4 (N8158, N8144, N4171, N7822, N788);
nor NOR2 (N8159, N8156, N6445);
nor NOR2 (N8160, N8157, N487);
nor NOR2 (N8161, N8160, N7206);
nor NOR4 (N8162, N8150, N3019, N5589, N2289);
nand NAND2 (N8163, N8137, N5735);
and AND3 (N8164, N8152, N2474, N162);
xor XOR2 (N8165, N8155, N7143);
or OR2 (N8166, N8134, N604);
or OR3 (N8167, N8159, N4713, N409);
not NOT1 (N8168, N8161);
and AND4 (N8169, N8147, N4080, N3567, N1286);
buf BUF1 (N8170, N8163);
not NOT1 (N8171, N8169);
not NOT1 (N8172, N8167);
xor XOR2 (N8173, N8170, N1307);
or OR3 (N8174, N8168, N42, N6797);
xor XOR2 (N8175, N8171, N6147);
nor NOR3 (N8176, N8158, N4568, N2675);
nor NOR3 (N8177, N8176, N795, N2426);
nor NOR4 (N8178, N8165, N3909, N1752, N5917);
buf BUF1 (N8179, N8164);
or OR3 (N8180, N8166, N995, N3525);
not NOT1 (N8181, N8178);
not NOT1 (N8182, N8177);
nor NOR2 (N8183, N8173, N6088);
or OR2 (N8184, N8175, N3066);
or OR3 (N8185, N8174, N260, N5275);
nand NAND2 (N8186, N8182, N7832);
nor NOR3 (N8187, N8172, N5995, N2506);
buf BUF1 (N8188, N8181);
nor NOR4 (N8189, N8187, N4597, N6804, N8001);
buf BUF1 (N8190, N8189);
not NOT1 (N8191, N8186);
not NOT1 (N8192, N8179);
or OR4 (N8193, N8192, N3638, N3490, N6376);
buf BUF1 (N8194, N8190);
xor XOR2 (N8195, N8188, N7012);
xor XOR2 (N8196, N8180, N903);
nand NAND3 (N8197, N8194, N1694, N7092);
not NOT1 (N8198, N8185);
and AND2 (N8199, N8191, N6619);
or OR3 (N8200, N8199, N7005, N3401);
xor XOR2 (N8201, N8195, N3603);
nor NOR3 (N8202, N8201, N940, N3968);
buf BUF1 (N8203, N8148);
not NOT1 (N8204, N8183);
xor XOR2 (N8205, N8198, N1477);
buf BUF1 (N8206, N8196);
buf BUF1 (N8207, N8202);
buf BUF1 (N8208, N8197);
xor XOR2 (N8209, N8208, N693);
not NOT1 (N8210, N8193);
and AND3 (N8211, N8205, N6485, N5431);
buf BUF1 (N8212, N8211);
or OR2 (N8213, N8184, N2239);
or OR3 (N8214, N8209, N1647, N6927);
and AND2 (N8215, N8213, N308);
not NOT1 (N8216, N8203);
and AND4 (N8217, N8210, N5405, N3977, N5897);
xor XOR2 (N8218, N8216, N5166);
buf BUF1 (N8219, N8218);
not NOT1 (N8220, N8206);
not NOT1 (N8221, N8212);
nor NOR3 (N8222, N8200, N3593, N2363);
buf BUF1 (N8223, N8222);
nor NOR2 (N8224, N8221, N7719);
and AND4 (N8225, N8220, N2261, N5728, N5699);
not NOT1 (N8226, N8215);
not NOT1 (N8227, N8223);
buf BUF1 (N8228, N8207);
buf BUF1 (N8229, N8217);
nand NAND3 (N8230, N8229, N5054, N4694);
not NOT1 (N8231, N8162);
and AND4 (N8232, N8225, N7955, N3380, N6538);
nand NAND4 (N8233, N8214, N2514, N7414, N4429);
not NOT1 (N8234, N8227);
xor XOR2 (N8235, N8233, N3852);
nand NAND4 (N8236, N8228, N1824, N1464, N4476);
nand NAND3 (N8237, N8226, N2331, N3577);
nand NAND3 (N8238, N8230, N8175, N5640);
or OR3 (N8239, N8219, N6369, N368);
buf BUF1 (N8240, N8231);
nand NAND3 (N8241, N8234, N7068, N2582);
and AND3 (N8242, N8236, N803, N123);
not NOT1 (N8243, N8204);
or OR2 (N8244, N8243, N6212);
not NOT1 (N8245, N8232);
xor XOR2 (N8246, N8241, N1008);
buf BUF1 (N8247, N8242);
xor XOR2 (N8248, N8239, N417);
or OR3 (N8249, N8248, N524, N1702);
not NOT1 (N8250, N8249);
xor XOR2 (N8251, N8235, N7812);
xor XOR2 (N8252, N8240, N8250);
and AND4 (N8253, N4913, N6648, N3607, N3080);
not NOT1 (N8254, N8244);
nor NOR4 (N8255, N8254, N1336, N8079, N6252);
nand NAND3 (N8256, N8237, N5843, N5755);
not NOT1 (N8257, N8238);
and AND2 (N8258, N8224, N4104);
and AND2 (N8259, N8251, N2337);
xor XOR2 (N8260, N8258, N1355);
nand NAND4 (N8261, N8252, N3025, N2253, N15);
buf BUF1 (N8262, N8259);
and AND4 (N8263, N8260, N6377, N3064, N6688);
nand NAND4 (N8264, N8247, N7111, N3564, N3626);
buf BUF1 (N8265, N8255);
nand NAND2 (N8266, N8263, N3283);
or OR3 (N8267, N8261, N4298, N886);
not NOT1 (N8268, N8267);
nand NAND4 (N8269, N8245, N1228, N1176, N792);
and AND4 (N8270, N8256, N5045, N225, N2407);
not NOT1 (N8271, N8253);
or OR3 (N8272, N8262, N6989, N4810);
nand NAND4 (N8273, N8246, N5415, N3357, N4746);
xor XOR2 (N8274, N8272, N6191);
or OR3 (N8275, N8257, N7623, N6099);
xor XOR2 (N8276, N8264, N5154);
or OR3 (N8277, N8269, N4307, N2968);
nor NOR4 (N8278, N8265, N3164, N6142, N5548);
buf BUF1 (N8279, N8271);
or OR2 (N8280, N8278, N3615);
buf BUF1 (N8281, N8276);
and AND3 (N8282, N8277, N4529, N2670);
xor XOR2 (N8283, N8280, N7472);
buf BUF1 (N8284, N8283);
or OR4 (N8285, N8284, N7986, N3212, N7886);
nor NOR3 (N8286, N8275, N7753, N4858);
or OR3 (N8287, N8279, N3981, N3301);
not NOT1 (N8288, N8281);
xor XOR2 (N8289, N8268, N7339);
xor XOR2 (N8290, N8282, N8039);
or OR3 (N8291, N8285, N5105, N5367);
buf BUF1 (N8292, N8289);
buf BUF1 (N8293, N8287);
and AND2 (N8294, N8270, N4086);
not NOT1 (N8295, N8273);
and AND3 (N8296, N8288, N5832, N7678);
not NOT1 (N8297, N8290);
xor XOR2 (N8298, N8292, N5733);
buf BUF1 (N8299, N8291);
nand NAND2 (N8300, N8296, N7337);
nand NAND4 (N8301, N8298, N4086, N7238, N1868);
nor NOR2 (N8302, N8266, N3260);
buf BUF1 (N8303, N8302);
not NOT1 (N8304, N8300);
and AND4 (N8305, N8301, N1054, N1642, N7547);
buf BUF1 (N8306, N8299);
nand NAND2 (N8307, N8306, N793);
or OR4 (N8308, N8297, N3284, N5980, N5672);
nand NAND3 (N8309, N8294, N5783, N6247);
or OR4 (N8310, N8293, N2968, N1226, N3131);
and AND3 (N8311, N8303, N3057, N4780);
buf BUF1 (N8312, N8305);
buf BUF1 (N8313, N8311);
not NOT1 (N8314, N8274);
or OR3 (N8315, N8309, N2907, N5132);
xor XOR2 (N8316, N8314, N7523);
and AND2 (N8317, N8307, N3136);
xor XOR2 (N8318, N8310, N3808);
xor XOR2 (N8319, N8316, N4522);
and AND2 (N8320, N8317, N1899);
nor NOR4 (N8321, N8319, N7297, N4114, N5218);
buf BUF1 (N8322, N8286);
buf BUF1 (N8323, N8321);
buf BUF1 (N8324, N8323);
buf BUF1 (N8325, N8295);
xor XOR2 (N8326, N8320, N3778);
xor XOR2 (N8327, N8304, N6559);
buf BUF1 (N8328, N8313);
nand NAND3 (N8329, N8322, N4925, N652);
nand NAND3 (N8330, N8327, N3372, N1941);
xor XOR2 (N8331, N8312, N4712);
or OR2 (N8332, N8308, N5390);
nor NOR4 (N8333, N8318, N41, N994, N938);
or OR3 (N8334, N8325, N8047, N1829);
buf BUF1 (N8335, N8328);
nor NOR2 (N8336, N8335, N3362);
buf BUF1 (N8337, N8333);
nor NOR4 (N8338, N8324, N3374, N6310, N5135);
buf BUF1 (N8339, N8336);
not NOT1 (N8340, N8329);
and AND3 (N8341, N8339, N4926, N7720);
and AND3 (N8342, N8315, N8146, N2693);
not NOT1 (N8343, N8340);
xor XOR2 (N8344, N8343, N7556);
xor XOR2 (N8345, N8330, N5858);
nor NOR4 (N8346, N8342, N4858, N5034, N1754);
nand NAND4 (N8347, N8344, N1357, N1763, N2556);
and AND4 (N8348, N8345, N4853, N3672, N603);
xor XOR2 (N8349, N8337, N5318);
nand NAND3 (N8350, N8341, N4509, N1491);
and AND3 (N8351, N8348, N3223, N6035);
and AND4 (N8352, N8350, N7330, N126, N1297);
xor XOR2 (N8353, N8349, N6346);
or OR4 (N8354, N8351, N7867, N1147, N7950);
and AND4 (N8355, N8353, N4868, N2222, N2221);
nor NOR3 (N8356, N8326, N1076, N4317);
nor NOR2 (N8357, N8331, N6528);
and AND4 (N8358, N8352, N5278, N1136, N8091);
or OR4 (N8359, N8356, N4116, N5382, N5644);
nand NAND3 (N8360, N8359, N7172, N2469);
xor XOR2 (N8361, N8355, N6937);
xor XOR2 (N8362, N8361, N2307);
xor XOR2 (N8363, N8347, N5644);
xor XOR2 (N8364, N8357, N4475);
not NOT1 (N8365, N8362);
xor XOR2 (N8366, N8354, N3582);
or OR2 (N8367, N8360, N3438);
not NOT1 (N8368, N8346);
xor XOR2 (N8369, N8364, N4107);
buf BUF1 (N8370, N8367);
buf BUF1 (N8371, N8370);
not NOT1 (N8372, N8365);
buf BUF1 (N8373, N8371);
not NOT1 (N8374, N8334);
nor NOR4 (N8375, N8366, N3877, N5430, N296);
and AND3 (N8376, N8375, N3538, N3677);
or OR4 (N8377, N8338, N6211, N2109, N3663);
not NOT1 (N8378, N8372);
or OR2 (N8379, N8373, N4305);
buf BUF1 (N8380, N8378);
nand NAND2 (N8381, N8374, N2666);
or OR4 (N8382, N8376, N3789, N2890, N4644);
nor NOR3 (N8383, N8369, N3833, N793);
nand NAND2 (N8384, N8382, N7529);
xor XOR2 (N8385, N8384, N3);
not NOT1 (N8386, N8358);
or OR3 (N8387, N8385, N3880, N4772);
nor NOR3 (N8388, N8379, N3595, N8079);
or OR2 (N8389, N8388, N7663);
xor XOR2 (N8390, N8368, N6900);
buf BUF1 (N8391, N8377);
nand NAND3 (N8392, N8389, N2807, N2456);
nand NAND3 (N8393, N8383, N402, N1943);
xor XOR2 (N8394, N8381, N7192);
nand NAND2 (N8395, N8392, N2608);
nand NAND4 (N8396, N8387, N2336, N2394, N6267);
buf BUF1 (N8397, N8390);
nand NAND4 (N8398, N8394, N3334, N4802, N5173);
not NOT1 (N8399, N8386);
xor XOR2 (N8400, N8397, N7703);
buf BUF1 (N8401, N8332);
and AND4 (N8402, N8380, N7698, N6059, N2258);
xor XOR2 (N8403, N8363, N1577);
nand NAND4 (N8404, N8395, N7746, N6061, N5637);
or OR3 (N8405, N8403, N3782, N18);
and AND2 (N8406, N8393, N3171);
xor XOR2 (N8407, N8391, N6673);
not NOT1 (N8408, N8406);
or OR4 (N8409, N8399, N1913, N3347, N5402);
nor NOR2 (N8410, N8402, N8088);
nor NOR4 (N8411, N8400, N8149, N3887, N1656);
xor XOR2 (N8412, N8404, N1688);
or OR3 (N8413, N8401, N4999, N7556);
and AND4 (N8414, N8408, N6395, N1126, N1329);
buf BUF1 (N8415, N8411);
and AND3 (N8416, N8415, N3809, N3889);
and AND4 (N8417, N8416, N1724, N1656, N257);
or OR3 (N8418, N8417, N8106, N5967);
xor XOR2 (N8419, N8409, N4341);
or OR4 (N8420, N8418, N489, N3880, N7066);
not NOT1 (N8421, N8413);
nor NOR4 (N8422, N8405, N7730, N6522, N5266);
or OR2 (N8423, N8407, N3485);
not NOT1 (N8424, N8419);
nand NAND4 (N8425, N8396, N5692, N265, N2789);
nand NAND4 (N8426, N8423, N7702, N5370, N1952);
not NOT1 (N8427, N8414);
not NOT1 (N8428, N8422);
or OR2 (N8429, N8410, N5079);
nor NOR3 (N8430, N8412, N4118, N1319);
or OR2 (N8431, N8424, N3289);
xor XOR2 (N8432, N8420, N5949);
buf BUF1 (N8433, N8427);
not NOT1 (N8434, N8433);
not NOT1 (N8435, N8398);
nand NAND4 (N8436, N8432, N106, N5125, N7524);
nor NOR2 (N8437, N8435, N5901);
buf BUF1 (N8438, N8430);
nor NOR4 (N8439, N8437, N1207, N970, N2554);
or OR3 (N8440, N8429, N6240, N7244);
not NOT1 (N8441, N8431);
buf BUF1 (N8442, N8436);
xor XOR2 (N8443, N8425, N3208);
not NOT1 (N8444, N8438);
nor NOR3 (N8445, N8428, N4448, N6250);
and AND4 (N8446, N8443, N1115, N6645, N6925);
xor XOR2 (N8447, N8444, N341);
not NOT1 (N8448, N8441);
xor XOR2 (N8449, N8439, N3062);
not NOT1 (N8450, N8445);
xor XOR2 (N8451, N8442, N1904);
nand NAND3 (N8452, N8447, N7945, N2699);
and AND4 (N8453, N8440, N1740, N4986, N1912);
not NOT1 (N8454, N8450);
or OR2 (N8455, N8453, N1165);
nor NOR3 (N8456, N8426, N7421, N529);
xor XOR2 (N8457, N8451, N1210);
nor NOR2 (N8458, N8449, N7581);
and AND4 (N8459, N8434, N343, N2108, N5893);
not NOT1 (N8460, N8454);
and AND2 (N8461, N8448, N3743);
nor NOR3 (N8462, N8455, N7232, N8074);
nand NAND2 (N8463, N8460, N8185);
nor NOR3 (N8464, N8446, N1752, N7860);
not NOT1 (N8465, N8452);
buf BUF1 (N8466, N8457);
nand NAND3 (N8467, N8462, N6714, N1861);
not NOT1 (N8468, N8459);
nor NOR4 (N8469, N8458, N199, N4254, N7456);
xor XOR2 (N8470, N8464, N3645);
nand NAND2 (N8471, N8467, N7347);
nand NAND3 (N8472, N8465, N2285, N6917);
and AND4 (N8473, N8461, N7558, N3156, N4580);
buf BUF1 (N8474, N8421);
nand NAND4 (N8475, N8470, N6212, N5781, N3117);
not NOT1 (N8476, N8471);
nor NOR4 (N8477, N8469, N5447, N6676, N7413);
buf BUF1 (N8478, N8456);
or OR4 (N8479, N8476, N5328, N8281, N6306);
or OR2 (N8480, N8475, N5926);
xor XOR2 (N8481, N8474, N7074);
nand NAND2 (N8482, N8468, N2215);
nand NAND3 (N8483, N8463, N1427, N3766);
xor XOR2 (N8484, N8472, N2760);
or OR2 (N8485, N8483, N4341);
nor NOR4 (N8486, N8482, N7324, N4951, N1091);
and AND2 (N8487, N8479, N4109);
not NOT1 (N8488, N8486);
nor NOR4 (N8489, N8485, N7354, N5503, N8241);
xor XOR2 (N8490, N8473, N7555);
buf BUF1 (N8491, N8488);
not NOT1 (N8492, N8487);
or OR2 (N8493, N8490, N2470);
nand NAND4 (N8494, N8489, N7437, N4448, N4779);
buf BUF1 (N8495, N8493);
nor NOR2 (N8496, N8492, N3330);
nand NAND2 (N8497, N8466, N4414);
or OR2 (N8498, N8491, N1452);
and AND2 (N8499, N8497, N2021);
nand NAND4 (N8500, N8477, N4323, N6373, N6227);
nand NAND4 (N8501, N8496, N4267, N4329, N2179);
or OR2 (N8502, N8498, N1529);
nand NAND3 (N8503, N8499, N2925, N4740);
not NOT1 (N8504, N8478);
xor XOR2 (N8505, N8503, N2317);
and AND4 (N8506, N8502, N8144, N2183, N7275);
and AND3 (N8507, N8501, N1061, N761);
nand NAND2 (N8508, N8506, N6130);
xor XOR2 (N8509, N8508, N3246);
nand NAND4 (N8510, N8480, N4714, N3850, N1853);
or OR4 (N8511, N8510, N4554, N1803, N6016);
not NOT1 (N8512, N8507);
and AND4 (N8513, N8481, N7018, N7607, N3751);
and AND3 (N8514, N8509, N8222, N3336);
buf BUF1 (N8515, N8494);
not NOT1 (N8516, N8511);
and AND3 (N8517, N8495, N6614, N3382);
nor NOR4 (N8518, N8504, N5496, N3266, N1973);
or OR2 (N8519, N8513, N5729);
or OR2 (N8520, N8517, N1450);
nand NAND3 (N8521, N8514, N3893, N4571);
nor NOR4 (N8522, N8520, N8042, N2328, N497);
xor XOR2 (N8523, N8518, N5988);
and AND4 (N8524, N8515, N6608, N1442, N7966);
and AND3 (N8525, N8522, N8353, N7643);
not NOT1 (N8526, N8500);
nand NAND4 (N8527, N8505, N7844, N8058, N5325);
xor XOR2 (N8528, N8516, N4574);
nor NOR4 (N8529, N8519, N6538, N4191, N487);
not NOT1 (N8530, N8525);
nand NAND2 (N8531, N8512, N1002);
xor XOR2 (N8532, N8523, N8276);
or OR3 (N8533, N8526, N7519, N4295);
not NOT1 (N8534, N8527);
nor NOR4 (N8535, N8528, N5435, N2739, N892);
or OR3 (N8536, N8524, N7652, N3094);
and AND2 (N8537, N8535, N3120);
nand NAND2 (N8538, N8529, N7067);
or OR2 (N8539, N8532, N4714);
xor XOR2 (N8540, N8539, N3031);
buf BUF1 (N8541, N8534);
nand NAND2 (N8542, N8521, N4088);
and AND2 (N8543, N8533, N4569);
buf BUF1 (N8544, N8536);
buf BUF1 (N8545, N8540);
nand NAND4 (N8546, N8545, N7530, N4909, N1876);
buf BUF1 (N8547, N8541);
nor NOR3 (N8548, N8547, N7722, N8098);
xor XOR2 (N8549, N8546, N3375);
buf BUF1 (N8550, N8538);
not NOT1 (N8551, N8537);
and AND2 (N8552, N8484, N6678);
buf BUF1 (N8553, N8543);
and AND4 (N8554, N8544, N7075, N6327, N6243);
nor NOR4 (N8555, N8530, N285, N2027, N482);
xor XOR2 (N8556, N8550, N7473);
or OR4 (N8557, N8553, N8115, N7650, N7007);
nor NOR4 (N8558, N8554, N344, N2235, N1019);
nand NAND3 (N8559, N8558, N7695, N2430);
buf BUF1 (N8560, N8542);
not NOT1 (N8561, N8555);
not NOT1 (N8562, N8561);
not NOT1 (N8563, N8551);
nor NOR3 (N8564, N8548, N1702, N2306);
xor XOR2 (N8565, N8560, N5075);
buf BUF1 (N8566, N8562);
buf BUF1 (N8567, N8564);
xor XOR2 (N8568, N8552, N2712);
or OR4 (N8569, N8531, N7536, N2529, N3164);
or OR2 (N8570, N8549, N3086);
nand NAND3 (N8571, N8559, N493, N5443);
xor XOR2 (N8572, N8566, N452);
and AND2 (N8573, N8565, N5585);
nor NOR4 (N8574, N8571, N3578, N8088, N5656);
or OR2 (N8575, N8567, N4897);
buf BUF1 (N8576, N8569);
not NOT1 (N8577, N8556);
not NOT1 (N8578, N8570);
and AND4 (N8579, N8576, N3375, N4814, N1967);
or OR4 (N8580, N8572, N5911, N8250, N2899);
or OR3 (N8581, N8557, N3911, N777);
nand NAND3 (N8582, N8563, N4810, N5444);
nand NAND4 (N8583, N8579, N6835, N4702, N6139);
and AND3 (N8584, N8573, N1753, N7058);
xor XOR2 (N8585, N8581, N445);
or OR3 (N8586, N8568, N2258, N6008);
buf BUF1 (N8587, N8575);
not NOT1 (N8588, N8578);
and AND3 (N8589, N8584, N5335, N2454);
and AND4 (N8590, N8583, N2169, N6081, N3164);
not NOT1 (N8591, N8586);
nand NAND3 (N8592, N8577, N1298, N148);
nor NOR4 (N8593, N8589, N1979, N1592, N7108);
xor XOR2 (N8594, N8587, N7476);
xor XOR2 (N8595, N8574, N635);
or OR2 (N8596, N8590, N6866);
and AND3 (N8597, N8594, N5857, N8146);
and AND3 (N8598, N8582, N3172, N2596);
nand NAND2 (N8599, N8592, N5202);
not NOT1 (N8600, N8593);
buf BUF1 (N8601, N8591);
and AND4 (N8602, N8599, N7122, N3032, N6747);
not NOT1 (N8603, N8600);
xor XOR2 (N8604, N8597, N7991);
and AND2 (N8605, N8595, N6430);
and AND4 (N8606, N8604, N1464, N5467, N7761);
or OR4 (N8607, N8596, N5895, N7135, N929);
not NOT1 (N8608, N8603);
nand NAND3 (N8609, N8598, N2831, N2283);
nand NAND3 (N8610, N8588, N1119, N5164);
not NOT1 (N8611, N8601);
nand NAND3 (N8612, N8580, N2493, N3570);
or OR3 (N8613, N8606, N2992, N5110);
buf BUF1 (N8614, N8613);
buf BUF1 (N8615, N8608);
not NOT1 (N8616, N8585);
xor XOR2 (N8617, N8616, N5991);
nor NOR4 (N8618, N8611, N1363, N3237, N152);
buf BUF1 (N8619, N8602);
and AND4 (N8620, N8612, N4080, N1698, N6132);
nor NOR4 (N8621, N8605, N174, N4975, N5022);
or OR4 (N8622, N8620, N6048, N4853, N2358);
buf BUF1 (N8623, N8610);
not NOT1 (N8624, N8622);
nand NAND3 (N8625, N8621, N4545, N8175);
buf BUF1 (N8626, N8614);
not NOT1 (N8627, N8623);
not NOT1 (N8628, N8627);
or OR3 (N8629, N8609, N4822, N7756);
nand NAND3 (N8630, N8625, N8473, N3631);
buf BUF1 (N8631, N8618);
nand NAND4 (N8632, N8615, N7228, N7836, N2872);
xor XOR2 (N8633, N8631, N8292);
xor XOR2 (N8634, N8624, N3632);
xor XOR2 (N8635, N8607, N1142);
nand NAND4 (N8636, N8633, N5165, N2072, N1575);
xor XOR2 (N8637, N8632, N1492);
buf BUF1 (N8638, N8619);
nand NAND3 (N8639, N8628, N6916, N7127);
nor NOR4 (N8640, N8630, N5804, N7868, N3502);
and AND3 (N8641, N8637, N8640, N6433);
nand NAND3 (N8642, N4674, N8487, N7545);
or OR3 (N8643, N8641, N3442, N5526);
and AND4 (N8644, N8617, N7341, N6883, N8507);
not NOT1 (N8645, N8629);
xor XOR2 (N8646, N8642, N3558);
not NOT1 (N8647, N8646);
nor NOR2 (N8648, N8645, N5154);
xor XOR2 (N8649, N8636, N2606);
or OR2 (N8650, N8643, N4641);
nand NAND2 (N8651, N8634, N4892);
buf BUF1 (N8652, N8649);
not NOT1 (N8653, N8652);
and AND4 (N8654, N8638, N6475, N3066, N5439);
buf BUF1 (N8655, N8653);
xor XOR2 (N8656, N8635, N1251);
not NOT1 (N8657, N8655);
nand NAND3 (N8658, N8651, N5169, N7172);
or OR4 (N8659, N8639, N7627, N7672, N950);
xor XOR2 (N8660, N8650, N4058);
buf BUF1 (N8661, N8656);
nor NOR2 (N8662, N8647, N4936);
or OR3 (N8663, N8658, N7233, N6523);
not NOT1 (N8664, N8659);
nand NAND3 (N8665, N8660, N7307, N4378);
and AND4 (N8666, N8661, N140, N1439, N1797);
or OR3 (N8667, N8657, N8180, N1071);
nor NOR2 (N8668, N8665, N2583);
and AND3 (N8669, N8662, N7369, N963);
not NOT1 (N8670, N8664);
nor NOR3 (N8671, N8654, N5765, N7286);
not NOT1 (N8672, N8668);
or OR4 (N8673, N8626, N2653, N3263, N3305);
or OR2 (N8674, N8673, N1317);
nor NOR4 (N8675, N8663, N8141, N3223, N8305);
nand NAND3 (N8676, N8672, N6192, N1972);
buf BUF1 (N8677, N8676);
or OR3 (N8678, N8677, N5222, N941);
or OR2 (N8679, N8670, N5038);
not NOT1 (N8680, N8678);
not NOT1 (N8681, N8680);
nand NAND2 (N8682, N8667, N3506);
nor NOR4 (N8683, N8671, N6848, N8117, N997);
or OR3 (N8684, N8648, N8661, N3535);
not NOT1 (N8685, N8674);
not NOT1 (N8686, N8679);
nor NOR3 (N8687, N8685, N8363, N3030);
nor NOR3 (N8688, N8666, N2441, N4466);
nor NOR3 (N8689, N8682, N669, N5442);
and AND3 (N8690, N8688, N4351, N3862);
nand NAND3 (N8691, N8675, N4398, N2503);
xor XOR2 (N8692, N8684, N4057);
nand NAND2 (N8693, N8690, N4513);
and AND2 (N8694, N8681, N1226);
xor XOR2 (N8695, N8691, N6202);
not NOT1 (N8696, N8692);
xor XOR2 (N8697, N8686, N8257);
buf BUF1 (N8698, N8697);
not NOT1 (N8699, N8696);
xor XOR2 (N8700, N8669, N2845);
and AND3 (N8701, N8693, N8397, N2952);
nand NAND3 (N8702, N8698, N2935, N8451);
or OR3 (N8703, N8687, N5234, N4379);
or OR4 (N8704, N8699, N6036, N8011, N365);
buf BUF1 (N8705, N8689);
or OR3 (N8706, N8683, N6723, N7906);
nor NOR3 (N8707, N8702, N7639, N7027);
nor NOR2 (N8708, N8705, N2884);
buf BUF1 (N8709, N8701);
nand NAND3 (N8710, N8703, N2816, N7070);
not NOT1 (N8711, N8644);
and AND4 (N8712, N8711, N1370, N511, N284);
xor XOR2 (N8713, N8704, N1168);
nor NOR4 (N8714, N8713, N5003, N5841, N6321);
buf BUF1 (N8715, N8700);
not NOT1 (N8716, N8712);
or OR4 (N8717, N8695, N3118, N560, N5727);
buf BUF1 (N8718, N8715);
and AND3 (N8719, N8717, N5775, N1652);
buf BUF1 (N8720, N8719);
and AND4 (N8721, N8716, N6914, N1019, N3444);
buf BUF1 (N8722, N8721);
and AND4 (N8723, N8722, N3983, N5061, N4542);
nand NAND2 (N8724, N8714, N5579);
nand NAND2 (N8725, N8720, N7849);
nand NAND4 (N8726, N8725, N7012, N8135, N2272);
buf BUF1 (N8727, N8726);
nand NAND3 (N8728, N8707, N5431, N3304);
or OR2 (N8729, N8727, N2658);
and AND3 (N8730, N8718, N3792, N4671);
or OR2 (N8731, N8706, N280);
xor XOR2 (N8732, N8723, N6412);
xor XOR2 (N8733, N8729, N8199);
not NOT1 (N8734, N8708);
nor NOR4 (N8735, N8710, N4754, N772, N1963);
nand NAND4 (N8736, N8730, N502, N1453, N7351);
buf BUF1 (N8737, N8735);
xor XOR2 (N8738, N8733, N7086);
buf BUF1 (N8739, N8738);
or OR2 (N8740, N8734, N4949);
nor NOR4 (N8741, N8737, N7431, N5230, N3204);
nand NAND3 (N8742, N8741, N1768, N1652);
or OR3 (N8743, N8709, N1961, N4052);
xor XOR2 (N8744, N8739, N6219);
not NOT1 (N8745, N8728);
nor NOR3 (N8746, N8694, N5349, N7844);
not NOT1 (N8747, N8736);
and AND2 (N8748, N8744, N5797);
not NOT1 (N8749, N8747);
not NOT1 (N8750, N8732);
and AND4 (N8751, N8742, N5366, N1891, N4447);
and AND3 (N8752, N8750, N440, N874);
and AND4 (N8753, N8752, N1207, N7193, N872);
not NOT1 (N8754, N8740);
and AND4 (N8755, N8754, N2960, N5386, N5178);
nor NOR2 (N8756, N8755, N617);
or OR3 (N8757, N8751, N5700, N6996);
or OR2 (N8758, N8745, N3334);
and AND3 (N8759, N8746, N2751, N1168);
not NOT1 (N8760, N8724);
xor XOR2 (N8761, N8758, N1615);
or OR4 (N8762, N8759, N3577, N771, N1216);
not NOT1 (N8763, N8753);
buf BUF1 (N8764, N8748);
not NOT1 (N8765, N8731);
and AND2 (N8766, N8762, N6774);
not NOT1 (N8767, N8764);
xor XOR2 (N8768, N8760, N5949);
or OR4 (N8769, N8756, N5484, N4906, N4010);
nand NAND3 (N8770, N8749, N6512, N5598);
nand NAND3 (N8771, N8769, N3545, N8659);
nor NOR2 (N8772, N8770, N4809);
xor XOR2 (N8773, N8772, N1670);
not NOT1 (N8774, N8766);
nor NOR4 (N8775, N8765, N2743, N2621, N4868);
nand NAND3 (N8776, N8774, N8732, N6910);
or OR2 (N8777, N8775, N2573);
nor NOR4 (N8778, N8773, N3857, N1087, N5522);
nor NOR3 (N8779, N8768, N5915, N8410);
buf BUF1 (N8780, N8743);
not NOT1 (N8781, N8763);
or OR3 (N8782, N8777, N7591, N4200);
nor NOR3 (N8783, N8757, N8664, N4124);
and AND4 (N8784, N8780, N2216, N518, N4930);
xor XOR2 (N8785, N8771, N4875);
xor XOR2 (N8786, N8776, N402);
nor NOR3 (N8787, N8784, N8062, N6805);
nand NAND2 (N8788, N8782, N1085);
nor NOR4 (N8789, N8783, N3505, N3060, N3187);
or OR2 (N8790, N8785, N4080);
buf BUF1 (N8791, N8781);
nand NAND2 (N8792, N8767, N1043);
nor NOR2 (N8793, N8787, N7034);
or OR2 (N8794, N8788, N2440);
buf BUF1 (N8795, N8791);
buf BUF1 (N8796, N8792);
or OR2 (N8797, N8761, N224);
and AND2 (N8798, N8789, N7063);
nor NOR3 (N8799, N8790, N685, N6581);
and AND3 (N8800, N8799, N3429, N3689);
nand NAND3 (N8801, N8800, N7544, N2385);
and AND3 (N8802, N8795, N2815, N511);
xor XOR2 (N8803, N8779, N1574);
and AND2 (N8804, N8794, N506);
xor XOR2 (N8805, N8798, N5409);
nor NOR3 (N8806, N8778, N2981, N5512);
or OR2 (N8807, N8804, N5616);
not NOT1 (N8808, N8797);
nor NOR4 (N8809, N8807, N7336, N8796, N8715);
not NOT1 (N8810, N5566);
nor NOR4 (N8811, N8805, N3993, N5361, N2977);
buf BUF1 (N8812, N8806);
or OR4 (N8813, N8793, N6331, N8451, N6815);
nand NAND4 (N8814, N8810, N3033, N5288, N2547);
buf BUF1 (N8815, N8803);
and AND3 (N8816, N8812, N3200, N5936);
not NOT1 (N8817, N8802);
nor NOR2 (N8818, N8811, N6618);
not NOT1 (N8819, N8816);
or OR2 (N8820, N8818, N7643);
or OR3 (N8821, N8815, N394, N152);
xor XOR2 (N8822, N8809, N4095);
xor XOR2 (N8823, N8821, N2159);
buf BUF1 (N8824, N8801);
buf BUF1 (N8825, N8813);
nor NOR3 (N8826, N8817, N7850, N1928);
nand NAND4 (N8827, N8819, N4539, N3509, N6326);
and AND3 (N8828, N8814, N1198, N4107);
and AND4 (N8829, N8826, N3599, N1432, N2824);
nand NAND3 (N8830, N8828, N6643, N6861);
nor NOR3 (N8831, N8829, N3617, N4358);
buf BUF1 (N8832, N8824);
or OR3 (N8833, N8822, N3145, N4953);
xor XOR2 (N8834, N8823, N2479);
buf BUF1 (N8835, N8832);
buf BUF1 (N8836, N8833);
xor XOR2 (N8837, N8834, N5323);
nand NAND3 (N8838, N8825, N8373, N887);
not NOT1 (N8839, N8838);
or OR3 (N8840, N8820, N5812, N2466);
nand NAND4 (N8841, N8831, N3825, N6285, N1473);
nor NOR2 (N8842, N8840, N6753);
or OR4 (N8843, N8837, N2821, N2086, N529);
or OR4 (N8844, N8835, N4645, N5319, N6279);
not NOT1 (N8845, N8844);
nand NAND4 (N8846, N8827, N3045, N5744, N2371);
not NOT1 (N8847, N8845);
or OR3 (N8848, N8846, N6428, N1029);
not NOT1 (N8849, N8808);
nand NAND3 (N8850, N8836, N1154, N1855);
or OR2 (N8851, N8847, N8306);
nand NAND3 (N8852, N8851, N410, N7113);
not NOT1 (N8853, N8786);
buf BUF1 (N8854, N8853);
or OR3 (N8855, N8848, N6173, N3238);
buf BUF1 (N8856, N8855);
or OR4 (N8857, N8843, N5155, N4186, N7478);
nor NOR4 (N8858, N8852, N5491, N8558, N7185);
nor NOR2 (N8859, N8858, N5133);
and AND3 (N8860, N8857, N8818, N7297);
nor NOR2 (N8861, N8842, N668);
not NOT1 (N8862, N8856);
or OR2 (N8863, N8850, N1906);
nand NAND4 (N8864, N8860, N8478, N8271, N5337);
not NOT1 (N8865, N8830);
not NOT1 (N8866, N8865);
nor NOR3 (N8867, N8864, N6323, N1404);
nand NAND2 (N8868, N8849, N6079);
not NOT1 (N8869, N8861);
buf BUF1 (N8870, N8862);
or OR4 (N8871, N8859, N1529, N1349, N6818);
nor NOR2 (N8872, N8869, N8721);
buf BUF1 (N8873, N8871);
buf BUF1 (N8874, N8873);
nand NAND3 (N8875, N8839, N6371, N2689);
and AND2 (N8876, N8875, N1204);
and AND2 (N8877, N8876, N4035);
nor NOR3 (N8878, N8877, N8338, N7311);
nor NOR3 (N8879, N8866, N1951, N3802);
nor NOR4 (N8880, N8863, N6707, N110, N6561);
buf BUF1 (N8881, N8872);
nand NAND4 (N8882, N8878, N7891, N1179, N4680);
xor XOR2 (N8883, N8881, N1611);
buf BUF1 (N8884, N8867);
nor NOR2 (N8885, N8884, N8766);
buf BUF1 (N8886, N8880);
and AND4 (N8887, N8870, N5833, N1420, N1954);
buf BUF1 (N8888, N8885);
nand NAND3 (N8889, N8868, N8801, N7573);
and AND4 (N8890, N8887, N5391, N1345, N6853);
or OR4 (N8891, N8854, N6674, N2583, N4265);
or OR3 (N8892, N8841, N4501, N8491);
and AND4 (N8893, N8879, N6841, N5407, N4294);
nand NAND2 (N8894, N8891, N8245);
xor XOR2 (N8895, N8882, N209);
not NOT1 (N8896, N8892);
or OR4 (N8897, N8895, N2396, N1889, N6775);
xor XOR2 (N8898, N8893, N1683);
and AND2 (N8899, N8894, N8667);
or OR4 (N8900, N8890, N2924, N3751, N2635);
not NOT1 (N8901, N8874);
nor NOR2 (N8902, N8896, N6105);
or OR3 (N8903, N8886, N2451, N505);
and AND2 (N8904, N8897, N1639);
or OR4 (N8905, N8883, N3891, N2330, N2750);
and AND2 (N8906, N8901, N7555);
or OR2 (N8907, N8888, N514);
or OR4 (N8908, N8905, N7471, N1052, N5542);
nor NOR4 (N8909, N8908, N55, N4391, N4006);
xor XOR2 (N8910, N8889, N5426);
buf BUF1 (N8911, N8902);
not NOT1 (N8912, N8900);
nand NAND3 (N8913, N8899, N6366, N2600);
nand NAND4 (N8914, N8907, N1827, N5948, N71);
or OR2 (N8915, N8903, N2796);
not NOT1 (N8916, N8913);
nor NOR3 (N8917, N8904, N1802, N8272);
nor NOR2 (N8918, N8911, N2830);
nand NAND4 (N8919, N8912, N2030, N1791, N5087);
buf BUF1 (N8920, N8906);
nand NAND3 (N8921, N8914, N6199, N1308);
nand NAND2 (N8922, N8921, N5035);
and AND3 (N8923, N8920, N463, N7019);
not NOT1 (N8924, N8917);
buf BUF1 (N8925, N8915);
nand NAND3 (N8926, N8922, N7819, N8414);
not NOT1 (N8927, N8909);
or OR3 (N8928, N8916, N5533, N2481);
xor XOR2 (N8929, N8919, N5985);
xor XOR2 (N8930, N8898, N1837);
and AND2 (N8931, N8928, N4937);
not NOT1 (N8932, N8918);
or OR3 (N8933, N8932, N501, N6680);
nand NAND2 (N8934, N8927, N7639);
buf BUF1 (N8935, N8910);
xor XOR2 (N8936, N8925, N1577);
or OR2 (N8937, N8934, N1834);
xor XOR2 (N8938, N8936, N2843);
or OR2 (N8939, N8935, N2225);
and AND2 (N8940, N8939, N5975);
nand NAND2 (N8941, N8931, N1137);
xor XOR2 (N8942, N8937, N5296);
not NOT1 (N8943, N8941);
and AND2 (N8944, N8929, N8275);
not NOT1 (N8945, N8938);
and AND2 (N8946, N8943, N174);
buf BUF1 (N8947, N8945);
nor NOR4 (N8948, N8947, N6134, N7707, N907);
buf BUF1 (N8949, N8944);
or OR2 (N8950, N8949, N1352);
xor XOR2 (N8951, N8923, N2134);
xor XOR2 (N8952, N8926, N2486);
nand NAND4 (N8953, N8940, N6742, N6304, N2318);
not NOT1 (N8954, N8946);
not NOT1 (N8955, N8930);
nor NOR2 (N8956, N8924, N2780);
buf BUF1 (N8957, N8933);
or OR4 (N8958, N8955, N3383, N2526, N6314);
nand NAND3 (N8959, N8953, N3345, N4518);
not NOT1 (N8960, N8957);
and AND2 (N8961, N8950, N1717);
nand NAND3 (N8962, N8956, N7776, N8028);
and AND3 (N8963, N8942, N7925, N3081);
and AND2 (N8964, N8952, N2258);
xor XOR2 (N8965, N8960, N1670);
buf BUF1 (N8966, N8959);
or OR4 (N8967, N8962, N8459, N6626, N3753);
not NOT1 (N8968, N8954);
or OR4 (N8969, N8948, N7987, N2854, N5999);
or OR4 (N8970, N8968, N749, N6077, N2820);
not NOT1 (N8971, N8965);
xor XOR2 (N8972, N8966, N7457);
or OR4 (N8973, N8958, N1230, N6318, N7310);
or OR2 (N8974, N8964, N4451);
or OR2 (N8975, N8967, N8500);
nor NOR2 (N8976, N8970, N3969);
nand NAND2 (N8977, N8971, N7875);
buf BUF1 (N8978, N8969);
or OR4 (N8979, N8974, N2715, N7133, N1093);
not NOT1 (N8980, N8951);
or OR4 (N8981, N8977, N5925, N8866, N7357);
buf BUF1 (N8982, N8961);
nor NOR3 (N8983, N8976, N7895, N157);
buf BUF1 (N8984, N8963);
nand NAND2 (N8985, N8983, N4338);
xor XOR2 (N8986, N8985, N4474);
or OR3 (N8987, N8986, N4524, N8857);
nor NOR3 (N8988, N8987, N3489, N50);
buf BUF1 (N8989, N8984);
nor NOR4 (N8990, N8988, N6148, N89, N632);
not NOT1 (N8991, N8989);
or OR3 (N8992, N8990, N8542, N3737);
nor NOR3 (N8993, N8975, N7607, N3193);
nor NOR2 (N8994, N8978, N3423);
buf BUF1 (N8995, N8993);
or OR2 (N8996, N8995, N7754);
not NOT1 (N8997, N8973);
or OR2 (N8998, N8994, N8375);
or OR2 (N8999, N8991, N3983);
not NOT1 (N9000, N8992);
and AND4 (N9001, N8980, N8117, N1998, N6504);
buf BUF1 (N9002, N8982);
not NOT1 (N9003, N8998);
nand NAND4 (N9004, N8972, N7343, N8214, N8948);
buf BUF1 (N9005, N8981);
or OR4 (N9006, N8996, N2205, N4288, N7833);
nor NOR4 (N9007, N9004, N7884, N5106, N877);
nand NAND2 (N9008, N9007, N8983);
xor XOR2 (N9009, N9005, N2304);
xor XOR2 (N9010, N9001, N7835);
or OR3 (N9011, N9010, N2205, N139);
xor XOR2 (N9012, N9003, N2726);
nor NOR4 (N9013, N9011, N7925, N7936, N7012);
not NOT1 (N9014, N9008);
buf BUF1 (N9015, N9006);
or OR3 (N9016, N8979, N4957, N4155);
and AND4 (N9017, N9009, N6475, N4636, N5311);
and AND3 (N9018, N9012, N5526, N6300);
or OR2 (N9019, N9017, N8367);
nand NAND3 (N9020, N8999, N8324, N565);
nor NOR3 (N9021, N9019, N8017, N560);
and AND3 (N9022, N9018, N1414, N4147);
and AND4 (N9023, N9000, N1301, N1431, N1702);
buf BUF1 (N9024, N8997);
xor XOR2 (N9025, N9022, N5757);
nand NAND3 (N9026, N9015, N8095, N3914);
buf BUF1 (N9027, N9002);
nor NOR3 (N9028, N9013, N5001, N309);
not NOT1 (N9029, N9021);
nand NAND4 (N9030, N9029, N344, N6121, N1300);
or OR2 (N9031, N9028, N6538);
and AND2 (N9032, N9023, N4577);
nand NAND4 (N9033, N9024, N8421, N2129, N4495);
nor NOR4 (N9034, N9027, N8038, N2203, N5250);
xor XOR2 (N9035, N9031, N8366);
xor XOR2 (N9036, N9034, N8366);
nor NOR3 (N9037, N9025, N8331, N7352);
and AND3 (N9038, N9016, N6682, N8966);
or OR3 (N9039, N9014, N4760, N2676);
nor NOR2 (N9040, N9035, N8886);
or OR3 (N9041, N9030, N4134, N8368);
not NOT1 (N9042, N9037);
and AND2 (N9043, N9033, N1913);
buf BUF1 (N9044, N9038);
buf BUF1 (N9045, N9026);
and AND4 (N9046, N9020, N2588, N7919, N5256);
nand NAND4 (N9047, N9041, N522, N416, N7214);
buf BUF1 (N9048, N9042);
or OR4 (N9049, N9039, N2236, N5615, N8761);
nand NAND4 (N9050, N9044, N1253, N7879, N462);
xor XOR2 (N9051, N9046, N1234);
buf BUF1 (N9052, N9047);
and AND2 (N9053, N9036, N4876);
nand NAND2 (N9054, N9040, N6613);
nand NAND4 (N9055, N9049, N2121, N2804, N5077);
and AND4 (N9056, N9051, N8857, N4527, N6162);
buf BUF1 (N9057, N9045);
nand NAND4 (N9058, N9050, N8378, N6742, N6467);
nand NAND3 (N9059, N9057, N1079, N5717);
nand NAND4 (N9060, N9056, N166, N1361, N4920);
xor XOR2 (N9061, N9054, N5181);
xor XOR2 (N9062, N9061, N5590);
or OR4 (N9063, N9055, N8377, N4580, N8736);
not NOT1 (N9064, N9048);
and AND4 (N9065, N9059, N917, N2716, N4859);
buf BUF1 (N9066, N9062);
or OR3 (N9067, N9043, N1937, N5654);
nor NOR2 (N9068, N9052, N5239);
xor XOR2 (N9069, N9032, N6289);
and AND4 (N9070, N9069, N2090, N2884, N187);
buf BUF1 (N9071, N9065);
xor XOR2 (N9072, N9053, N696);
nand NAND2 (N9073, N9060, N2112);
or OR4 (N9074, N9071, N2921, N8678, N5873);
nor NOR4 (N9075, N9074, N6381, N4919, N1128);
or OR2 (N9076, N9063, N3241);
not NOT1 (N9077, N9072);
nor NOR3 (N9078, N9075, N5461, N662);
xor XOR2 (N9079, N9078, N6940);
or OR4 (N9080, N9064, N1397, N2471, N7703);
not NOT1 (N9081, N9076);
and AND3 (N9082, N9081, N6148, N3424);
xor XOR2 (N9083, N9073, N6191);
nand NAND3 (N9084, N9083, N6989, N4444);
nand NAND4 (N9085, N9067, N5225, N1363, N2834);
nor NOR2 (N9086, N9085, N1060);
xor XOR2 (N9087, N9080, N1739);
nor NOR4 (N9088, N9058, N4292, N4165, N5626);
xor XOR2 (N9089, N9068, N6114);
buf BUF1 (N9090, N9079);
xor XOR2 (N9091, N9086, N4499);
buf BUF1 (N9092, N9084);
or OR2 (N9093, N9087, N7146);
not NOT1 (N9094, N9090);
and AND4 (N9095, N9089, N4251, N1396, N1433);
nor NOR2 (N9096, N9095, N2599);
xor XOR2 (N9097, N9096, N5977);
buf BUF1 (N9098, N9094);
nor NOR2 (N9099, N9093, N4821);
or OR3 (N9100, N9091, N2980, N522);
nand NAND3 (N9101, N9099, N5179, N2456);
xor XOR2 (N9102, N9092, N8390);
buf BUF1 (N9103, N9088);
nor NOR4 (N9104, N9082, N3775, N4309, N8907);
not NOT1 (N9105, N9066);
buf BUF1 (N9106, N9105);
nand NAND4 (N9107, N9070, N3970, N631, N3168);
nand NAND2 (N9108, N9106, N5462);
buf BUF1 (N9109, N9102);
nand NAND3 (N9110, N9100, N492, N2265);
nand NAND4 (N9111, N9077, N3205, N2094, N7258);
buf BUF1 (N9112, N9101);
buf BUF1 (N9113, N9112);
or OR3 (N9114, N9109, N8986, N5366);
buf BUF1 (N9115, N9108);
nor NOR2 (N9116, N9103, N3934);
and AND2 (N9117, N9104, N7145);
and AND4 (N9118, N9116, N6894, N1195, N2787);
nor NOR3 (N9119, N9098, N5292, N6925);
nand NAND4 (N9120, N9111, N8796, N8208, N4816);
or OR2 (N9121, N9114, N9035);
nor NOR3 (N9122, N9120, N2527, N344);
xor XOR2 (N9123, N9113, N7445);
xor XOR2 (N9124, N9123, N3789);
not NOT1 (N9125, N9122);
and AND2 (N9126, N9118, N4343);
or OR4 (N9127, N9121, N8231, N4101, N1658);
nor NOR2 (N9128, N9127, N4530);
not NOT1 (N9129, N9117);
not NOT1 (N9130, N9107);
nor NOR4 (N9131, N9110, N4830, N2521, N2247);
nand NAND2 (N9132, N9126, N8902);
or OR3 (N9133, N9119, N980, N6523);
or OR3 (N9134, N9115, N3301, N2430);
buf BUF1 (N9135, N9132);
nor NOR2 (N9136, N9097, N4193);
not NOT1 (N9137, N9136);
not NOT1 (N9138, N9125);
nand NAND3 (N9139, N9128, N1380, N8379);
nor NOR2 (N9140, N9124, N7701);
and AND2 (N9141, N9130, N2913);
buf BUF1 (N9142, N9129);
and AND3 (N9143, N9138, N5925, N5023);
buf BUF1 (N9144, N9137);
xor XOR2 (N9145, N9140, N4744);
xor XOR2 (N9146, N9142, N9046);
nand NAND3 (N9147, N9135, N7232, N8997);
and AND3 (N9148, N9145, N3668, N375);
nor NOR2 (N9149, N9143, N5591);
buf BUF1 (N9150, N9131);
and AND4 (N9151, N9146, N2774, N1929, N1530);
buf BUF1 (N9152, N9149);
not NOT1 (N9153, N9134);
nand NAND4 (N9154, N9133, N3006, N6771, N8553);
nand NAND2 (N9155, N9148, N180);
buf BUF1 (N9156, N9152);
xor XOR2 (N9157, N9147, N8162);
and AND4 (N9158, N9157, N2859, N4487, N6036);
nand NAND3 (N9159, N9150, N7844, N5409);
xor XOR2 (N9160, N9158, N9058);
nand NAND2 (N9161, N9154, N4575);
or OR4 (N9162, N9159, N6628, N6370, N6138);
not NOT1 (N9163, N9162);
nand NAND2 (N9164, N9139, N7000);
buf BUF1 (N9165, N9156);
nor NOR2 (N9166, N9163, N1704);
buf BUF1 (N9167, N9166);
nor NOR2 (N9168, N9153, N6081);
not NOT1 (N9169, N9141);
nor NOR2 (N9170, N9169, N4860);
not NOT1 (N9171, N9167);
buf BUF1 (N9172, N9144);
and AND3 (N9173, N9172, N9059, N3295);
and AND4 (N9174, N9155, N4915, N7323, N1210);
or OR4 (N9175, N9173, N6734, N341, N7604);
not NOT1 (N9176, N9151);
nor NOR3 (N9177, N9164, N7331, N5124);
and AND3 (N9178, N9165, N2183, N3090);
buf BUF1 (N9179, N9177);
xor XOR2 (N9180, N9170, N4950);
nand NAND4 (N9181, N9176, N6721, N3180, N7095);
buf BUF1 (N9182, N9178);
nand NAND3 (N9183, N9180, N6608, N2515);
or OR4 (N9184, N9181, N5737, N8507, N2127);
nor NOR2 (N9185, N9160, N7362);
xor XOR2 (N9186, N9175, N9126);
nor NOR2 (N9187, N9186, N873);
nor NOR2 (N9188, N9182, N855);
and AND3 (N9189, N9171, N7981, N5584);
buf BUF1 (N9190, N9185);
and AND4 (N9191, N9188, N2067, N2089, N122);
nand NAND2 (N9192, N9168, N8349);
buf BUF1 (N9193, N9192);
nor NOR4 (N9194, N9193, N7720, N506, N6498);
nand NAND4 (N9195, N9179, N7433, N4124, N1951);
nand NAND3 (N9196, N9190, N2378, N5140);
and AND4 (N9197, N9196, N6612, N8022, N1461);
and AND4 (N9198, N9161, N8438, N3105, N7270);
xor XOR2 (N9199, N9189, N7630);
and AND3 (N9200, N9194, N8563, N6478);
not NOT1 (N9201, N9197);
buf BUF1 (N9202, N9187);
nand NAND3 (N9203, N9200, N7693, N544);
nor NOR2 (N9204, N9198, N6487);
buf BUF1 (N9205, N9183);
or OR3 (N9206, N9195, N7856, N744);
nand NAND4 (N9207, N9202, N2267, N3153, N3218);
nand NAND4 (N9208, N9203, N3040, N8328, N2602);
nand NAND4 (N9209, N9201, N7868, N7716, N8680);
nand NAND3 (N9210, N9184, N2331, N1519);
buf BUF1 (N9211, N9199);
and AND4 (N9212, N9174, N1567, N6105, N1548);
or OR3 (N9213, N9209, N795, N4074);
nand NAND3 (N9214, N9213, N7510, N5917);
not NOT1 (N9215, N9208);
xor XOR2 (N9216, N9215, N2209);
buf BUF1 (N9217, N9210);
nor NOR2 (N9218, N9205, N298);
buf BUF1 (N9219, N9204);
xor XOR2 (N9220, N9191, N7448);
not NOT1 (N9221, N9214);
or OR2 (N9222, N9207, N7802);
nand NAND3 (N9223, N9218, N6220, N3184);
nand NAND4 (N9224, N9206, N1110, N3944, N9029);
or OR2 (N9225, N9223, N7321);
buf BUF1 (N9226, N9211);
and AND2 (N9227, N9220, N5771);
not NOT1 (N9228, N9225);
or OR3 (N9229, N9226, N8656, N806);
or OR4 (N9230, N9228, N7645, N9187, N7890);
and AND2 (N9231, N9224, N5719);
nor NOR3 (N9232, N9212, N4947, N5540);
or OR3 (N9233, N9216, N9192, N7289);
nor NOR3 (N9234, N9233, N5979, N2134);
not NOT1 (N9235, N9234);
and AND2 (N9236, N9235, N2010);
xor XOR2 (N9237, N9230, N7779);
and AND4 (N9238, N9217, N8454, N8634, N2999);
not NOT1 (N9239, N9237);
nand NAND2 (N9240, N9229, N3868);
buf BUF1 (N9241, N9239);
buf BUF1 (N9242, N9227);
not NOT1 (N9243, N9219);
xor XOR2 (N9244, N9232, N1765);
and AND4 (N9245, N9236, N7816, N8864, N818);
not NOT1 (N9246, N9231);
nand NAND4 (N9247, N9244, N3451, N8590, N4222);
xor XOR2 (N9248, N9246, N2087);
and AND2 (N9249, N9247, N3954);
nand NAND4 (N9250, N9222, N603, N7678, N5231);
and AND4 (N9251, N9240, N361, N4379, N8488);
and AND4 (N9252, N9221, N1750, N6823, N8477);
not NOT1 (N9253, N9248);
nor NOR3 (N9254, N9241, N7682, N1127);
buf BUF1 (N9255, N9254);
nand NAND4 (N9256, N9250, N6776, N9041, N7312);
xor XOR2 (N9257, N9251, N3423);
xor XOR2 (N9258, N9257, N7133);
or OR2 (N9259, N9238, N189);
xor XOR2 (N9260, N9245, N2184);
xor XOR2 (N9261, N9259, N947);
or OR3 (N9262, N9261, N1996, N6508);
and AND3 (N9263, N9255, N3456, N5413);
or OR3 (N9264, N9258, N6338, N3636);
and AND2 (N9265, N9249, N8204);
nor NOR4 (N9266, N9262, N7133, N7141, N1279);
buf BUF1 (N9267, N9260);
buf BUF1 (N9268, N9266);
nand NAND2 (N9269, N9264, N1317);
and AND2 (N9270, N9252, N4819);
or OR4 (N9271, N9256, N8956, N2405, N1952);
nor NOR3 (N9272, N9271, N8074, N1305);
not NOT1 (N9273, N9270);
nand NAND4 (N9274, N9267, N3591, N7296, N6000);
buf BUF1 (N9275, N9242);
xor XOR2 (N9276, N9243, N241);
not NOT1 (N9277, N9263);
and AND3 (N9278, N9277, N6129, N5366);
nor NOR2 (N9279, N9275, N4903);
not NOT1 (N9280, N9278);
and AND4 (N9281, N9272, N4343, N8350, N3737);
not NOT1 (N9282, N9269);
or OR2 (N9283, N9273, N5253);
not NOT1 (N9284, N9276);
nor NOR3 (N9285, N9280, N1975, N5156);
xor XOR2 (N9286, N9265, N3815);
or OR3 (N9287, N9253, N4221, N375);
or OR3 (N9288, N9274, N5155, N7681);
nand NAND3 (N9289, N9288, N5422, N4517);
and AND2 (N9290, N9279, N4088);
nor NOR4 (N9291, N9286, N2221, N5423, N6408);
not NOT1 (N9292, N9290);
not NOT1 (N9293, N9283);
nor NOR2 (N9294, N9292, N421);
not NOT1 (N9295, N9282);
xor XOR2 (N9296, N9284, N5114);
and AND4 (N9297, N9287, N7065, N7391, N4920);
xor XOR2 (N9298, N9285, N2305);
and AND4 (N9299, N9295, N6276, N7755, N2331);
or OR4 (N9300, N9281, N8635, N164, N7054);
xor XOR2 (N9301, N9300, N2883);
nor NOR4 (N9302, N9301, N1633, N3182, N1215);
nand NAND2 (N9303, N9299, N9051);
buf BUF1 (N9304, N9296);
xor XOR2 (N9305, N9304, N3589);
nand NAND4 (N9306, N9291, N8119, N9229, N6611);
or OR2 (N9307, N9306, N1259);
nand NAND2 (N9308, N9302, N3836);
buf BUF1 (N9309, N9289);
nand NAND3 (N9310, N9307, N2916, N6186);
and AND3 (N9311, N9310, N6404, N5447);
xor XOR2 (N9312, N9293, N5905);
xor XOR2 (N9313, N9298, N7599);
buf BUF1 (N9314, N9312);
nand NAND3 (N9315, N9297, N8994, N2585);
not NOT1 (N9316, N9294);
not NOT1 (N9317, N9314);
xor XOR2 (N9318, N9309, N7703);
or OR2 (N9319, N9318, N677);
nand NAND4 (N9320, N9319, N9155, N7610, N3376);
nor NOR3 (N9321, N9308, N5975, N7742);
xor XOR2 (N9322, N9303, N1351);
or OR3 (N9323, N9321, N5945, N7789);
or OR3 (N9324, N9317, N1479, N91);
nand NAND4 (N9325, N9323, N4887, N4485, N5321);
nor NOR3 (N9326, N9324, N7594, N1598);
not NOT1 (N9327, N9315);
and AND3 (N9328, N9268, N7702, N7604);
nand NAND4 (N9329, N9313, N1964, N220, N567);
nor NOR2 (N9330, N9328, N2798);
buf BUF1 (N9331, N9327);
not NOT1 (N9332, N9325);
or OR2 (N9333, N9326, N8516);
nand NAND3 (N9334, N9305, N9013, N8432);
nor NOR4 (N9335, N9334, N38, N982, N419);
nor NOR3 (N9336, N9320, N5378, N3503);
buf BUF1 (N9337, N9332);
buf BUF1 (N9338, N9316);
and AND2 (N9339, N9338, N1218);
and AND4 (N9340, N9336, N5687, N7361, N1230);
and AND2 (N9341, N9311, N9047);
or OR3 (N9342, N9330, N4135, N5172);
nand NAND3 (N9343, N9333, N1211, N306);
not NOT1 (N9344, N9342);
xor XOR2 (N9345, N9322, N1079);
xor XOR2 (N9346, N9345, N4602);
nand NAND4 (N9347, N9329, N5145, N5801, N8237);
buf BUF1 (N9348, N9337);
nand NAND2 (N9349, N9343, N1055);
nand NAND2 (N9350, N9348, N2645);
nor NOR2 (N9351, N9335, N7252);
and AND2 (N9352, N9346, N7971);
and AND4 (N9353, N9340, N7946, N6519, N4719);
nand NAND3 (N9354, N9339, N154, N2516);
and AND3 (N9355, N9344, N4756, N4327);
buf BUF1 (N9356, N9352);
and AND2 (N9357, N9347, N3310);
buf BUF1 (N9358, N9341);
and AND3 (N9359, N9354, N2084, N3326);
nand NAND4 (N9360, N9331, N5234, N3510, N3089);
and AND3 (N9361, N9350, N3638, N1743);
or OR4 (N9362, N9358, N7294, N2674, N8663);
or OR3 (N9363, N9359, N7587, N2013);
xor XOR2 (N9364, N9349, N3920);
not NOT1 (N9365, N9362);
nor NOR3 (N9366, N9355, N1444, N658);
xor XOR2 (N9367, N9361, N8046);
xor XOR2 (N9368, N9365, N7517);
buf BUF1 (N9369, N9353);
nand NAND4 (N9370, N9366, N5625, N8660, N6698);
buf BUF1 (N9371, N9360);
xor XOR2 (N9372, N9370, N1190);
and AND2 (N9373, N9351, N5105);
or OR4 (N9374, N9357, N6487, N629, N6283);
not NOT1 (N9375, N9356);
nand NAND2 (N9376, N9373, N2840);
nor NOR3 (N9377, N9363, N2341, N2517);
and AND3 (N9378, N9372, N3498, N5969);
xor XOR2 (N9379, N9369, N2519);
nand NAND4 (N9380, N9378, N1912, N323, N6961);
buf BUF1 (N9381, N9368);
xor XOR2 (N9382, N9379, N959);
or OR2 (N9383, N9375, N2419);
nand NAND3 (N9384, N9374, N9218, N6113);
or OR3 (N9385, N9380, N8622, N1590);
buf BUF1 (N9386, N9377);
nor NOR4 (N9387, N9382, N892, N3208, N4046);
not NOT1 (N9388, N9364);
nand NAND2 (N9389, N9383, N2943);
nor NOR4 (N9390, N9386, N2049, N4762, N7457);
not NOT1 (N9391, N9388);
or OR3 (N9392, N9376, N6341, N3516);
buf BUF1 (N9393, N9390);
nand NAND2 (N9394, N9392, N4703);
nor NOR3 (N9395, N9394, N9135, N3272);
nand NAND2 (N9396, N9391, N3929);
or OR4 (N9397, N9367, N4238, N4248, N2601);
or OR2 (N9398, N9384, N1609);
and AND4 (N9399, N9381, N4524, N8405, N6983);
buf BUF1 (N9400, N9387);
or OR2 (N9401, N9385, N2926);
xor XOR2 (N9402, N9393, N8176);
xor XOR2 (N9403, N9396, N2829);
buf BUF1 (N9404, N9401);
or OR3 (N9405, N9402, N7068, N8040);
buf BUF1 (N9406, N9371);
xor XOR2 (N9407, N9403, N4485);
not NOT1 (N9408, N9395);
and AND2 (N9409, N9397, N8489);
nor NOR3 (N9410, N9406, N3238, N8257);
and AND4 (N9411, N9399, N2763, N7502, N6383);
not NOT1 (N9412, N9389);
not NOT1 (N9413, N9410);
xor XOR2 (N9414, N9411, N1919);
nand NAND4 (N9415, N9412, N6637, N4692, N4353);
nor NOR3 (N9416, N9408, N4586, N3528);
and AND4 (N9417, N9404, N7429, N507, N4970);
or OR4 (N9418, N9405, N4552, N3434, N4022);
nor NOR2 (N9419, N9409, N5937);
nor NOR4 (N9420, N9417, N6435, N6160, N6200);
buf BUF1 (N9421, N9400);
or OR2 (N9422, N9420, N3184);
not NOT1 (N9423, N9414);
and AND2 (N9424, N9421, N7305);
or OR4 (N9425, N9419, N417, N6791, N5498);
nand NAND4 (N9426, N9407, N1296, N1265, N7124);
and AND4 (N9427, N9425, N2207, N5224, N8336);
or OR4 (N9428, N9422, N1249, N608, N4027);
not NOT1 (N9429, N9415);
not NOT1 (N9430, N9423);
and AND3 (N9431, N9416, N7349, N3896);
nor NOR3 (N9432, N9429, N2240, N7303);
buf BUF1 (N9433, N9418);
nor NOR2 (N9434, N9433, N2168);
not NOT1 (N9435, N9427);
not NOT1 (N9436, N9432);
not NOT1 (N9437, N9434);
nor NOR3 (N9438, N9437, N1666, N524);
nand NAND3 (N9439, N9428, N1171, N2203);
nor NOR3 (N9440, N9438, N815, N1965);
not NOT1 (N9441, N9430);
nor NOR2 (N9442, N9436, N762);
nor NOR4 (N9443, N9441, N2242, N9263, N7300);
buf BUF1 (N9444, N9435);
buf BUF1 (N9445, N9424);
buf BUF1 (N9446, N9431);
nor NOR4 (N9447, N9413, N7924, N5611, N1140);
buf BUF1 (N9448, N9446);
nor NOR3 (N9449, N9443, N2074, N3826);
nor NOR3 (N9450, N9445, N6125, N5174);
xor XOR2 (N9451, N9447, N1541);
xor XOR2 (N9452, N9451, N3849);
xor XOR2 (N9453, N9448, N2116);
and AND3 (N9454, N9398, N3976, N3668);
nor NOR3 (N9455, N9449, N4198, N5797);
nand NAND3 (N9456, N9444, N7779, N3801);
or OR3 (N9457, N9456, N9047, N468);
and AND2 (N9458, N9439, N140);
nand NAND3 (N9459, N9458, N7031, N8640);
xor XOR2 (N9460, N9453, N9046);
xor XOR2 (N9461, N9450, N986);
buf BUF1 (N9462, N9461);
nand NAND4 (N9463, N9457, N2201, N4132, N2663);
and AND2 (N9464, N9460, N3355);
and AND4 (N9465, N9464, N2660, N4248, N3744);
buf BUF1 (N9466, N9452);
and AND4 (N9467, N9465, N4393, N378, N3013);
nand NAND3 (N9468, N9466, N8105, N3676);
nor NOR2 (N9469, N9462, N1572);
buf BUF1 (N9470, N9442);
buf BUF1 (N9471, N9454);
buf BUF1 (N9472, N9468);
or OR4 (N9473, N9440, N5193, N2523, N4758);
nor NOR4 (N9474, N9455, N3189, N6620, N2315);
or OR2 (N9475, N9469, N5816);
and AND3 (N9476, N9459, N5437, N749);
or OR2 (N9477, N9476, N1792);
and AND4 (N9478, N9473, N1378, N1852, N5982);
and AND3 (N9479, N9463, N108, N1932);
nand NAND2 (N9480, N9478, N1036);
xor XOR2 (N9481, N9479, N4469);
nand NAND3 (N9482, N9472, N1837, N9460);
buf BUF1 (N9483, N9426);
buf BUF1 (N9484, N9481);
and AND3 (N9485, N9480, N3722, N843);
and AND3 (N9486, N9467, N984, N1964);
not NOT1 (N9487, N9471);
not NOT1 (N9488, N9477);
nor NOR4 (N9489, N9483, N2445, N2461, N6541);
not NOT1 (N9490, N9488);
xor XOR2 (N9491, N9490, N2188);
buf BUF1 (N9492, N9491);
not NOT1 (N9493, N9489);
buf BUF1 (N9494, N9493);
nor NOR2 (N9495, N9484, N6611);
and AND4 (N9496, N9485, N5619, N9097, N5068);
nand NAND3 (N9497, N9495, N7746, N1839);
and AND3 (N9498, N9492, N1104, N7775);
nand NAND2 (N9499, N9486, N2568);
nor NOR4 (N9500, N9498, N3137, N1266, N4519);
nor NOR3 (N9501, N9475, N7792, N7286);
xor XOR2 (N9502, N9470, N4805);
and AND3 (N9503, N9487, N7142, N4469);
and AND4 (N9504, N9496, N1719, N3803, N3845);
buf BUF1 (N9505, N9499);
nor NOR4 (N9506, N9494, N8255, N327, N6626);
nand NAND4 (N9507, N9503, N5326, N1218, N6850);
nor NOR3 (N9508, N9500, N5458, N4627);
xor XOR2 (N9509, N9508, N4738);
or OR2 (N9510, N9474, N7443);
nor NOR4 (N9511, N9497, N3966, N1060, N3842);
not NOT1 (N9512, N9509);
nor NOR2 (N9513, N9510, N7546);
xor XOR2 (N9514, N9505, N5446);
not NOT1 (N9515, N9501);
nor NOR2 (N9516, N9506, N6321);
and AND2 (N9517, N9516, N9494);
and AND2 (N9518, N9513, N2539);
nand NAND3 (N9519, N9514, N5561, N9330);
or OR3 (N9520, N9502, N1090, N7824);
nand NAND2 (N9521, N9519, N8463);
xor XOR2 (N9522, N9504, N1775);
buf BUF1 (N9523, N9511);
buf BUF1 (N9524, N9523);
xor XOR2 (N9525, N9524, N7012);
buf BUF1 (N9526, N9515);
xor XOR2 (N9527, N9525, N1082);
not NOT1 (N9528, N9526);
and AND4 (N9529, N9518, N2657, N4671, N4660);
nor NOR2 (N9530, N9520, N4415);
nand NAND2 (N9531, N9521, N6492);
not NOT1 (N9532, N9529);
nor NOR2 (N9533, N9527, N7857);
buf BUF1 (N9534, N9522);
nor NOR4 (N9535, N9528, N773, N5843, N1981);
and AND3 (N9536, N9535, N7574, N2527);
xor XOR2 (N9537, N9517, N3842);
or OR4 (N9538, N9482, N1396, N7105, N8375);
xor XOR2 (N9539, N9538, N2849);
or OR2 (N9540, N9536, N211);
not NOT1 (N9541, N9507);
nand NAND2 (N9542, N9530, N4970);
buf BUF1 (N9543, N9533);
or OR4 (N9544, N9531, N3108, N8958, N5583);
not NOT1 (N9545, N9512);
not NOT1 (N9546, N9541);
nor NOR3 (N9547, N9542, N864, N1434);
xor XOR2 (N9548, N9544, N9196);
nand NAND4 (N9549, N9545, N1782, N7484, N1466);
and AND3 (N9550, N9537, N3912, N9213);
or OR3 (N9551, N9543, N52, N3616);
buf BUF1 (N9552, N9539);
buf BUF1 (N9553, N9551);
xor XOR2 (N9554, N9550, N5989);
xor XOR2 (N9555, N9553, N5464);
nor NOR3 (N9556, N9555, N1465, N2146);
or OR4 (N9557, N9532, N6662, N1570, N9186);
xor XOR2 (N9558, N9540, N5674);
nor NOR3 (N9559, N9552, N4535, N4749);
buf BUF1 (N9560, N9556);
xor XOR2 (N9561, N9547, N9201);
buf BUF1 (N9562, N9534);
and AND2 (N9563, N9560, N453);
not NOT1 (N9564, N9554);
xor XOR2 (N9565, N9549, N1303);
and AND3 (N9566, N9559, N7652, N7376);
nand NAND4 (N9567, N9561, N5455, N1217, N9544);
or OR2 (N9568, N9557, N5586);
not NOT1 (N9569, N9558);
and AND2 (N9570, N9564, N4524);
buf BUF1 (N9571, N9569);
not NOT1 (N9572, N9567);
nor NOR3 (N9573, N9566, N8672, N608);
not NOT1 (N9574, N9572);
not NOT1 (N9575, N9563);
xor XOR2 (N9576, N9565, N4871);
xor XOR2 (N9577, N9546, N6934);
buf BUF1 (N9578, N9570);
nand NAND4 (N9579, N9562, N6163, N6600, N9272);
and AND4 (N9580, N9577, N602, N9120, N2622);
nor NOR4 (N9581, N9576, N5593, N4674, N4535);
not NOT1 (N9582, N9580);
not NOT1 (N9583, N9575);
not NOT1 (N9584, N9571);
buf BUF1 (N9585, N9573);
and AND3 (N9586, N9584, N8727, N7592);
and AND4 (N9587, N9582, N4261, N5008, N3129);
nor NOR2 (N9588, N9568, N9010);
and AND3 (N9589, N9588, N3541, N7820);
not NOT1 (N9590, N9579);
nand NAND3 (N9591, N9581, N7986, N5950);
xor XOR2 (N9592, N9591, N7255);
nand NAND2 (N9593, N9586, N2648);
buf BUF1 (N9594, N9592);
nand NAND2 (N9595, N9574, N6911);
nor NOR2 (N9596, N9585, N4754);
nor NOR4 (N9597, N9590, N8383, N8474, N9166);
and AND3 (N9598, N9548, N5033, N4176);
or OR4 (N9599, N9596, N6956, N7734, N5874);
buf BUF1 (N9600, N9589);
buf BUF1 (N9601, N9583);
buf BUF1 (N9602, N9597);
and AND2 (N9603, N9595, N6559);
nor NOR3 (N9604, N9601, N7932, N6204);
xor XOR2 (N9605, N9604, N7576);
not NOT1 (N9606, N9602);
and AND2 (N9607, N9603, N4064);
or OR2 (N9608, N9600, N6357);
nor NOR2 (N9609, N9608, N2549);
nand NAND4 (N9610, N9587, N4152, N8054, N1745);
xor XOR2 (N9611, N9606, N379);
xor XOR2 (N9612, N9594, N1730);
and AND2 (N9613, N9605, N1341);
not NOT1 (N9614, N9612);
nor NOR3 (N9615, N9614, N6729, N523);
buf BUF1 (N9616, N9609);
buf BUF1 (N9617, N9615);
or OR3 (N9618, N9616, N8819, N398);
nand NAND4 (N9619, N9598, N4007, N7573, N8863);
and AND4 (N9620, N9599, N4089, N1402, N3967);
nand NAND4 (N9621, N9613, N3095, N3657, N5965);
or OR2 (N9622, N9618, N2868);
xor XOR2 (N9623, N9619, N3967);
xor XOR2 (N9624, N9611, N3531);
buf BUF1 (N9625, N9622);
buf BUF1 (N9626, N9617);
nor NOR3 (N9627, N9621, N7528, N1375);
buf BUF1 (N9628, N9578);
not NOT1 (N9629, N9624);
and AND3 (N9630, N9626, N16, N2504);
not NOT1 (N9631, N9629);
nand NAND2 (N9632, N9623, N8407);
nand NAND2 (N9633, N9630, N2404);
xor XOR2 (N9634, N9620, N9019);
not NOT1 (N9635, N9625);
not NOT1 (N9636, N9607);
nand NAND4 (N9637, N9633, N8967, N8168, N2834);
buf BUF1 (N9638, N9632);
xor XOR2 (N9639, N9628, N8708);
nor NOR2 (N9640, N9610, N5535);
nor NOR4 (N9641, N9636, N625, N101, N793);
nor NOR3 (N9642, N9641, N8550, N2486);
or OR2 (N9643, N9642, N3123);
not NOT1 (N9644, N9637);
and AND4 (N9645, N9634, N9128, N3409, N104);
xor XOR2 (N9646, N9643, N8262);
xor XOR2 (N9647, N9639, N6587);
nand NAND2 (N9648, N9638, N8134);
nor NOR2 (N9649, N9645, N4921);
or OR4 (N9650, N9631, N1900, N6610, N4301);
xor XOR2 (N9651, N9646, N1612);
nand NAND4 (N9652, N9649, N2541, N8925, N7258);
and AND4 (N9653, N9627, N9405, N326, N1860);
nand NAND3 (N9654, N9648, N6162, N6508);
nand NAND4 (N9655, N9653, N1452, N2954, N863);
nor NOR3 (N9656, N9635, N7705, N893);
and AND3 (N9657, N9651, N4383, N2798);
buf BUF1 (N9658, N9652);
buf BUF1 (N9659, N9647);
buf BUF1 (N9660, N9658);
or OR3 (N9661, N9654, N2550, N9063);
not NOT1 (N9662, N9660);
buf BUF1 (N9663, N9593);
not NOT1 (N9664, N9655);
not NOT1 (N9665, N9663);
and AND2 (N9666, N9664, N9129);
buf BUF1 (N9667, N9640);
not NOT1 (N9668, N9662);
buf BUF1 (N9669, N9668);
buf BUF1 (N9670, N9644);
nor NOR4 (N9671, N9665, N8134, N7895, N8102);
or OR3 (N9672, N9650, N6932, N2910);
xor XOR2 (N9673, N9672, N6600);
nor NOR3 (N9674, N9670, N4958, N3876);
or OR3 (N9675, N9669, N9377, N4516);
and AND2 (N9676, N9667, N7308);
or OR3 (N9677, N9666, N9240, N5317);
nand NAND4 (N9678, N9656, N2833, N2039, N9381);
and AND2 (N9679, N9678, N8394);
nor NOR3 (N9680, N9657, N2947, N9340);
not NOT1 (N9681, N9659);
and AND3 (N9682, N9681, N6036, N2831);
and AND4 (N9683, N9676, N8016, N7467, N6167);
not NOT1 (N9684, N9682);
buf BUF1 (N9685, N9675);
buf BUF1 (N9686, N9679);
and AND4 (N9687, N9685, N6689, N932, N4698);
and AND4 (N9688, N9687, N4779, N8624, N7394);
nand NAND4 (N9689, N9686, N8896, N3307, N2985);
not NOT1 (N9690, N9671);
xor XOR2 (N9691, N9661, N7410);
buf BUF1 (N9692, N9680);
nor NOR2 (N9693, N9684, N9493);
nor NOR2 (N9694, N9693, N7076);
xor XOR2 (N9695, N9688, N6381);
xor XOR2 (N9696, N9673, N1488);
nand NAND4 (N9697, N9674, N1377, N5209, N3334);
buf BUF1 (N9698, N9697);
and AND4 (N9699, N9698, N5369, N4487, N1607);
nor NOR4 (N9700, N9691, N9394, N4022, N7124);
nor NOR3 (N9701, N9696, N7779, N4591);
and AND3 (N9702, N9690, N3378, N8043);
and AND2 (N9703, N9683, N4453);
xor XOR2 (N9704, N9689, N1147);
nand NAND3 (N9705, N9695, N4916, N280);
nand NAND4 (N9706, N9699, N3898, N6206, N3029);
nand NAND3 (N9707, N9692, N1214, N3101);
and AND2 (N9708, N9694, N8885);
nor NOR4 (N9709, N9702, N3421, N3425, N8252);
nand NAND4 (N9710, N9707, N265, N6653, N9698);
xor XOR2 (N9711, N9708, N8474);
not NOT1 (N9712, N9677);
or OR3 (N9713, N9706, N2440, N2237);
not NOT1 (N9714, N9709);
nand NAND4 (N9715, N9701, N3556, N1553, N698);
not NOT1 (N9716, N9712);
nand NAND3 (N9717, N9711, N2883, N898);
nor NOR2 (N9718, N9710, N4783);
not NOT1 (N9719, N9714);
buf BUF1 (N9720, N9718);
nand NAND2 (N9721, N9703, N3760);
nand NAND2 (N9722, N9713, N7717);
not NOT1 (N9723, N9721);
xor XOR2 (N9724, N9719, N8402);
nor NOR2 (N9725, N9716, N3682);
buf BUF1 (N9726, N9717);
nor NOR4 (N9727, N9704, N6769, N4393, N3307);
and AND3 (N9728, N9727, N163, N6897);
nand NAND3 (N9729, N9724, N5182, N6353);
or OR2 (N9730, N9728, N250);
and AND2 (N9731, N9705, N4216);
nor NOR4 (N9732, N9722, N1711, N7165, N9052);
buf BUF1 (N9733, N9729);
nand NAND4 (N9734, N9715, N6349, N58, N6901);
buf BUF1 (N9735, N9730);
buf BUF1 (N9736, N9732);
nor NOR4 (N9737, N9700, N8446, N190, N6177);
xor XOR2 (N9738, N9725, N4256);
xor XOR2 (N9739, N9726, N3090);
or OR3 (N9740, N9739, N5465, N3013);
xor XOR2 (N9741, N9736, N5620);
nor NOR4 (N9742, N9735, N1936, N6595, N3640);
nand NAND2 (N9743, N9742, N1781);
or OR3 (N9744, N9720, N6139, N586);
not NOT1 (N9745, N9738);
buf BUF1 (N9746, N9723);
and AND4 (N9747, N9743, N6831, N6971, N1303);
buf BUF1 (N9748, N9747);
and AND4 (N9749, N9737, N8516, N1571, N3386);
xor XOR2 (N9750, N9744, N2571);
or OR2 (N9751, N9734, N4935);
or OR3 (N9752, N9733, N8219, N8351);
and AND4 (N9753, N9745, N692, N3778, N8645);
and AND4 (N9754, N9749, N1720, N6008, N3915);
xor XOR2 (N9755, N9731, N7462);
nand NAND3 (N9756, N9752, N1833, N9124);
not NOT1 (N9757, N9753);
nand NAND2 (N9758, N9754, N1100);
xor XOR2 (N9759, N9758, N2996);
not NOT1 (N9760, N9756);
nor NOR2 (N9761, N9748, N319);
and AND4 (N9762, N9760, N2261, N2447, N9071);
nand NAND2 (N9763, N9746, N5315);
or OR2 (N9764, N9763, N1475);
xor XOR2 (N9765, N9759, N2258);
or OR2 (N9766, N9740, N7774);
xor XOR2 (N9767, N9766, N9053);
nor NOR2 (N9768, N9741, N1164);
and AND3 (N9769, N9761, N9463, N9600);
buf BUF1 (N9770, N9768);
or OR4 (N9771, N9767, N1545, N5873, N7076);
and AND3 (N9772, N9770, N3336, N2223);
nand NAND3 (N9773, N9765, N7800, N3971);
not NOT1 (N9774, N9769);
not NOT1 (N9775, N9774);
xor XOR2 (N9776, N9751, N93);
xor XOR2 (N9777, N9764, N3772);
or OR2 (N9778, N9777, N5650);
buf BUF1 (N9779, N9775);
or OR3 (N9780, N9776, N7337, N20);
buf BUF1 (N9781, N9773);
or OR3 (N9782, N9762, N1704, N2298);
nand NAND3 (N9783, N9782, N2586, N8434);
nor NOR2 (N9784, N9780, N1505);
nor NOR4 (N9785, N9771, N4516, N666, N2312);
buf BUF1 (N9786, N9781);
and AND4 (N9787, N9783, N6012, N4806, N6017);
xor XOR2 (N9788, N9772, N2892);
not NOT1 (N9789, N9750);
xor XOR2 (N9790, N9788, N7388);
xor XOR2 (N9791, N9755, N3383);
and AND4 (N9792, N9779, N9548, N9226, N2340);
or OR2 (N9793, N9785, N2819);
nor NOR4 (N9794, N9791, N6431, N6190, N5354);
nand NAND4 (N9795, N9787, N5602, N154, N4304);
xor XOR2 (N9796, N9794, N9786);
or OR2 (N9797, N8160, N6400);
buf BUF1 (N9798, N9792);
nor NOR3 (N9799, N9798, N7899, N4827);
or OR4 (N9800, N9797, N7732, N6717, N9152);
and AND2 (N9801, N9784, N6138);
nor NOR4 (N9802, N9801, N7334, N767, N9017);
not NOT1 (N9803, N9795);
xor XOR2 (N9804, N9789, N447);
nand NAND2 (N9805, N9790, N4794);
nand NAND2 (N9806, N9805, N2083);
nand NAND2 (N9807, N9793, N2406);
or OR4 (N9808, N9778, N621, N4585, N8020);
buf BUF1 (N9809, N9802);
nand NAND2 (N9810, N9799, N6792);
xor XOR2 (N9811, N9800, N2433);
buf BUF1 (N9812, N9809);
xor XOR2 (N9813, N9804, N7844);
and AND4 (N9814, N9803, N6574, N6123, N5646);
xor XOR2 (N9815, N9808, N2478);
buf BUF1 (N9816, N9812);
nand NAND2 (N9817, N9796, N7869);
xor XOR2 (N9818, N9816, N1892);
nand NAND3 (N9819, N9811, N32, N5850);
and AND3 (N9820, N9813, N8867, N4327);
or OR2 (N9821, N9757, N4059);
and AND2 (N9822, N9821, N8713);
nor NOR4 (N9823, N9817, N832, N6112, N7596);
not NOT1 (N9824, N9819);
and AND3 (N9825, N9822, N559, N692);
xor XOR2 (N9826, N9815, N9278);
buf BUF1 (N9827, N9826);
xor XOR2 (N9828, N9825, N9710);
buf BUF1 (N9829, N9814);
xor XOR2 (N9830, N9818, N1317);
nand NAND4 (N9831, N9820, N8093, N3736, N8465);
not NOT1 (N9832, N9806);
nor NOR3 (N9833, N9827, N8822, N9714);
or OR3 (N9834, N9810, N345, N2385);
nor NOR3 (N9835, N9834, N1122, N8185);
nor NOR4 (N9836, N9807, N1993, N8578, N5502);
buf BUF1 (N9837, N9832);
xor XOR2 (N9838, N9836, N4778);
nand NAND2 (N9839, N9835, N1315);
or OR4 (N9840, N9823, N2312, N2612, N3234);
xor XOR2 (N9841, N9833, N4555);
not NOT1 (N9842, N9837);
buf BUF1 (N9843, N9831);
and AND4 (N9844, N9829, N2021, N9016, N9271);
nand NAND2 (N9845, N9844, N6827);
not NOT1 (N9846, N9843);
not NOT1 (N9847, N9839);
not NOT1 (N9848, N9842);
not NOT1 (N9849, N9848);
nand NAND4 (N9850, N9828, N3266, N5123, N1290);
xor XOR2 (N9851, N9840, N6970);
nor NOR3 (N9852, N9851, N9262, N7596);
nand NAND2 (N9853, N9841, N9115);
not NOT1 (N9854, N9845);
or OR4 (N9855, N9850, N2457, N7434, N3588);
nand NAND3 (N9856, N9855, N9292, N7624);
buf BUF1 (N9857, N9852);
buf BUF1 (N9858, N9830);
or OR2 (N9859, N9856, N8479);
xor XOR2 (N9860, N9838, N2563);
buf BUF1 (N9861, N9860);
and AND4 (N9862, N9859, N5050, N3293, N2552);
nand NAND2 (N9863, N9857, N2327);
buf BUF1 (N9864, N9846);
not NOT1 (N9865, N9861);
xor XOR2 (N9866, N9854, N6980);
not NOT1 (N9867, N9849);
and AND2 (N9868, N9866, N5350);
nand NAND4 (N9869, N9853, N5737, N5991, N5534);
not NOT1 (N9870, N9824);
buf BUF1 (N9871, N9867);
buf BUF1 (N9872, N9847);
not NOT1 (N9873, N9870);
or OR2 (N9874, N9868, N5566);
and AND3 (N9875, N9863, N5060, N6394);
xor XOR2 (N9876, N9858, N6592);
xor XOR2 (N9877, N9871, N5835);
buf BUF1 (N9878, N9864);
buf BUF1 (N9879, N9869);
nor NOR3 (N9880, N9876, N6890, N1656);
nand NAND2 (N9881, N9878, N2230);
nor NOR4 (N9882, N9873, N82, N5218, N7066);
buf BUF1 (N9883, N9874);
nand NAND2 (N9884, N9881, N7167);
not NOT1 (N9885, N9877);
nand NAND4 (N9886, N9882, N4127, N3975, N1499);
nand NAND3 (N9887, N9879, N989, N9842);
not NOT1 (N9888, N9872);
xor XOR2 (N9889, N9875, N5009);
nor NOR2 (N9890, N9883, N5668);
xor XOR2 (N9891, N9890, N9888);
or OR2 (N9892, N2509, N1649);
not NOT1 (N9893, N9885);
xor XOR2 (N9894, N9892, N1920);
nor NOR4 (N9895, N9887, N6206, N2532, N2806);
or OR2 (N9896, N9893, N368);
nor NOR2 (N9897, N9884, N5848);
buf BUF1 (N9898, N9886);
nand NAND3 (N9899, N9880, N3662, N4329);
nand NAND2 (N9900, N9865, N5961);
or OR3 (N9901, N9894, N6645, N6128);
and AND3 (N9902, N9895, N7654, N500);
buf BUF1 (N9903, N9891);
nand NAND4 (N9904, N9902, N2447, N4926, N2010);
nand NAND3 (N9905, N9901, N6508, N8652);
or OR4 (N9906, N9896, N5542, N9627, N4051);
or OR4 (N9907, N9889, N5761, N3159, N7264);
not NOT1 (N9908, N9900);
nand NAND3 (N9909, N9897, N5805, N3566);
nand NAND3 (N9910, N9907, N190, N6488);
nand NAND3 (N9911, N9903, N2448, N9022);
not NOT1 (N9912, N9908);
and AND3 (N9913, N9899, N7109, N4414);
nor NOR3 (N9914, N9906, N6204, N6415);
or OR2 (N9915, N9904, N2648);
nand NAND4 (N9916, N9915, N4224, N5508, N2100);
not NOT1 (N9917, N9912);
nand NAND4 (N9918, N9913, N4707, N7917, N5495);
nand NAND4 (N9919, N9914, N6771, N2608, N7230);
buf BUF1 (N9920, N9905);
or OR3 (N9921, N9918, N3487, N8178);
buf BUF1 (N9922, N9910);
and AND3 (N9923, N9917, N8756, N4116);
nand NAND2 (N9924, N9916, N2929);
or OR3 (N9925, N9920, N5306, N6087);
and AND2 (N9926, N9898, N4264);
xor XOR2 (N9927, N9911, N3698);
and AND4 (N9928, N9923, N3723, N3604, N3547);
nand NAND2 (N9929, N9862, N9760);
not NOT1 (N9930, N9925);
not NOT1 (N9931, N9924);
or OR4 (N9932, N9921, N5122, N6741, N5778);
and AND3 (N9933, N9932, N7189, N3076);
nor NOR2 (N9934, N9926, N4828);
and AND2 (N9935, N9922, N5997);
nor NOR2 (N9936, N9933, N7296);
and AND3 (N9937, N9930, N7415, N3866);
nor NOR3 (N9938, N9928, N8078, N6415);
or OR4 (N9939, N9929, N833, N4034, N5805);
nor NOR3 (N9940, N9936, N1750, N736);
and AND2 (N9941, N9938, N1244);
not NOT1 (N9942, N9931);
not NOT1 (N9943, N9939);
nand NAND4 (N9944, N9919, N9500, N3472, N1602);
buf BUF1 (N9945, N9940);
xor XOR2 (N9946, N9935, N5449);
nand NAND3 (N9947, N9909, N9159, N3401);
or OR2 (N9948, N9937, N8756);
and AND2 (N9949, N9927, N6235);
not NOT1 (N9950, N9947);
or OR4 (N9951, N9943, N597, N5688, N87);
and AND3 (N9952, N9945, N9220, N5125);
or OR3 (N9953, N9946, N37, N9811);
and AND4 (N9954, N9944, N8922, N3149, N1418);
xor XOR2 (N9955, N9952, N912);
or OR3 (N9956, N9953, N4125, N9066);
and AND3 (N9957, N9954, N7091, N9777);
nand NAND2 (N9958, N9950, N3250);
xor XOR2 (N9959, N9958, N1255);
buf BUF1 (N9960, N9959);
not NOT1 (N9961, N9948);
buf BUF1 (N9962, N9941);
and AND2 (N9963, N9960, N7789);
nor NOR2 (N9964, N9957, N8859);
or OR3 (N9965, N9949, N1365, N9503);
nor NOR2 (N9966, N9963, N6031);
or OR2 (N9967, N9956, N8259);
xor XOR2 (N9968, N9967, N8245);
nor NOR3 (N9969, N9951, N8771, N786);
nor NOR2 (N9970, N9934, N4003);
not NOT1 (N9971, N9965);
or OR2 (N9972, N9961, N3563);
xor XOR2 (N9973, N9964, N7692);
buf BUF1 (N9974, N9962);
buf BUF1 (N9975, N9966);
and AND4 (N9976, N9975, N395, N3978, N4228);
xor XOR2 (N9977, N9970, N393);
not NOT1 (N9978, N9977);
xor XOR2 (N9979, N9976, N9523);
nand NAND3 (N9980, N9971, N2103, N8952);
or OR3 (N9981, N9978, N2379, N3767);
nor NOR4 (N9982, N9955, N1056, N3391, N9139);
nand NAND3 (N9983, N9942, N9367, N7917);
or OR4 (N9984, N9980, N221, N4435, N9885);
or OR4 (N9985, N9981, N3881, N4034, N304);
nor NOR2 (N9986, N9984, N9600);
or OR3 (N9987, N9973, N9653, N4911);
not NOT1 (N9988, N9986);
and AND4 (N9989, N9969, N9540, N1606, N3938);
and AND4 (N9990, N9983, N1244, N3561, N3403);
nor NOR3 (N9991, N9968, N4106, N4831);
and AND4 (N9992, N9972, N5384, N5498, N6223);
buf BUF1 (N9993, N9985);
not NOT1 (N9994, N9979);
nand NAND3 (N9995, N9992, N3960, N5618);
and AND4 (N9996, N9974, N3505, N8483, N859);
nand NAND2 (N9997, N9989, N9859);
buf BUF1 (N9998, N9996);
and AND4 (N9999, N9994, N3428, N1177, N3446);
nor NOR4 (N10000, N9999, N1534, N3821, N5241);
nand NAND3 (N10001, N9993, N3857, N7217);
buf BUF1 (N10002, N9997);
or OR3 (N10003, N9995, N4676, N6780);
nor NOR3 (N10004, N9990, N7964, N1363);
nor NOR2 (N10005, N9982, N5663);
nand NAND4 (N10006, N10003, N9673, N7637, N937);
not NOT1 (N10007, N10005);
nor NOR4 (N10008, N9991, N9327, N2579, N9161);
not NOT1 (N10009, N9987);
not NOT1 (N10010, N10002);
xor XOR2 (N10011, N10006, N1793);
nor NOR2 (N10012, N10009, N1657);
not NOT1 (N10013, N10011);
buf BUF1 (N10014, N10012);
buf BUF1 (N10015, N10014);
not NOT1 (N10016, N10013);
nand NAND2 (N10017, N9988, N3518);
nand NAND4 (N10018, N10001, N1407, N1014, N9326);
xor XOR2 (N10019, N9998, N4568);
xor XOR2 (N10020, N10000, N5815);
or OR4 (N10021, N10018, N2614, N8457, N6656);
buf BUF1 (N10022, N10021);
and AND2 (N10023, N10015, N7313);
nand NAND2 (N10024, N10007, N6351);
and AND4 (N10025, N10024, N2214, N3220, N8417);
nand NAND2 (N10026, N10008, N5198);
buf BUF1 (N10027, N10023);
or OR2 (N10028, N10004, N1851);
xor XOR2 (N10029, N10010, N7073);
xor XOR2 (N10030, N10029, N356);
xor XOR2 (N10031, N10026, N5466);
or OR4 (N10032, N10025, N3069, N9322, N7885);
nand NAND3 (N10033, N10030, N918, N8155);
buf BUF1 (N10034, N10019);
and AND4 (N10035, N10020, N7747, N6301, N7684);
xor XOR2 (N10036, N10034, N8180);
xor XOR2 (N10037, N10032, N9784);
not NOT1 (N10038, N10016);
and AND3 (N10039, N10022, N7399, N4116);
buf BUF1 (N10040, N10038);
buf BUF1 (N10041, N10033);
buf BUF1 (N10042, N10035);
not NOT1 (N10043, N10017);
nor NOR2 (N10044, N10042, N3184);
xor XOR2 (N10045, N10044, N3504);
nor NOR3 (N10046, N10040, N5728, N4004);
nand NAND4 (N10047, N10028, N8862, N8661, N1509);
buf BUF1 (N10048, N10047);
not NOT1 (N10049, N10046);
nand NAND3 (N10050, N10037, N3405, N9783);
not NOT1 (N10051, N10048);
buf BUF1 (N10052, N10036);
nor NOR2 (N10053, N10049, N49);
xor XOR2 (N10054, N10045, N9983);
nand NAND4 (N10055, N10051, N9904, N9076, N3497);
buf BUF1 (N10056, N10054);
or OR2 (N10057, N10056, N290);
xor XOR2 (N10058, N10039, N2991);
and AND2 (N10059, N10055, N2914);
and AND3 (N10060, N10041, N5596, N6373);
buf BUF1 (N10061, N10027);
and AND2 (N10062, N10057, N8522);
not NOT1 (N10063, N10031);
not NOT1 (N10064, N10061);
nor NOR3 (N10065, N10064, N955, N2290);
nor NOR4 (N10066, N10065, N6610, N6320, N4798);
and AND3 (N10067, N10050, N3412, N4107);
buf BUF1 (N10068, N10060);
and AND4 (N10069, N10058, N325, N2230, N6156);
nor NOR2 (N10070, N10063, N9601);
nand NAND2 (N10071, N10070, N3344);
nor NOR2 (N10072, N10069, N649);
or OR4 (N10073, N10043, N7455, N41, N7137);
or OR2 (N10074, N10073, N2736);
or OR2 (N10075, N10068, N6162);
and AND3 (N10076, N10074, N868, N8621);
xor XOR2 (N10077, N10076, N3475);
and AND3 (N10078, N10072, N8518, N6978);
xor XOR2 (N10079, N10071, N2121);
and AND2 (N10080, N10079, N271);
nor NOR4 (N10081, N10077, N8628, N2328, N4626);
or OR2 (N10082, N10078, N7492);
nand NAND3 (N10083, N10062, N1235, N5379);
not NOT1 (N10084, N10066);
and AND2 (N10085, N10084, N5483);
not NOT1 (N10086, N10085);
not NOT1 (N10087, N10067);
xor XOR2 (N10088, N10059, N2083);
buf BUF1 (N10089, N10081);
not NOT1 (N10090, N10080);
or OR2 (N10091, N10083, N7013);
buf BUF1 (N10092, N10087);
and AND2 (N10093, N10082, N1844);
or OR3 (N10094, N10092, N15, N3806);
or OR2 (N10095, N10091, N9541);
or OR3 (N10096, N10094, N9419, N6848);
or OR2 (N10097, N10088, N6238);
xor XOR2 (N10098, N10075, N7735);
not NOT1 (N10099, N10098);
nand NAND3 (N10100, N10097, N6540, N3775);
xor XOR2 (N10101, N10089, N9823);
or OR2 (N10102, N10090, N6207);
nor NOR4 (N10103, N10096, N5856, N3839, N7273);
nand NAND4 (N10104, N10103, N7958, N4190, N8365);
buf BUF1 (N10105, N10099);
buf BUF1 (N10106, N10102);
nand NAND4 (N10107, N10105, N7916, N677, N6557);
nor NOR3 (N10108, N10053, N985, N721);
and AND4 (N10109, N10100, N8400, N9638, N227);
buf BUF1 (N10110, N10109);
xor XOR2 (N10111, N10107, N6791);
xor XOR2 (N10112, N10110, N263);
and AND4 (N10113, N10101, N3114, N7312, N5641);
not NOT1 (N10114, N10113);
not NOT1 (N10115, N10108);
and AND4 (N10116, N10104, N1265, N7484, N2924);
and AND3 (N10117, N10111, N2643, N3);
not NOT1 (N10118, N10052);
or OR2 (N10119, N10117, N4033);
buf BUF1 (N10120, N10114);
and AND4 (N10121, N10115, N2804, N2701, N9540);
nor NOR2 (N10122, N10121, N2424);
and AND4 (N10123, N10116, N8310, N3249, N2709);
and AND3 (N10124, N10120, N3607, N1492);
not NOT1 (N10125, N10119);
and AND3 (N10126, N10112, N6020, N2874);
or OR4 (N10127, N10122, N9097, N2504, N4892);
buf BUF1 (N10128, N10126);
nor NOR3 (N10129, N10093, N8964, N7876);
or OR2 (N10130, N10106, N1398);
buf BUF1 (N10131, N10129);
nand NAND4 (N10132, N10124, N1135, N3585, N5575);
and AND4 (N10133, N10132, N8934, N6341, N5614);
nor NOR3 (N10134, N10130, N2126, N4652);
xor XOR2 (N10135, N10095, N4902);
buf BUF1 (N10136, N10127);
not NOT1 (N10137, N10086);
nand NAND2 (N10138, N10123, N4226);
nand NAND4 (N10139, N10118, N6702, N1086, N8463);
nand NAND2 (N10140, N10137, N6908);
xor XOR2 (N10141, N10136, N3630);
or OR2 (N10142, N10133, N8394);
not NOT1 (N10143, N10135);
nor NOR2 (N10144, N10139, N7355);
not NOT1 (N10145, N10125);
and AND4 (N10146, N10138, N6095, N4034, N4883);
or OR3 (N10147, N10146, N8081, N3290);
nand NAND4 (N10148, N10142, N5620, N5503, N9736);
buf BUF1 (N10149, N10145);
and AND4 (N10150, N10144, N1929, N2303, N5337);
buf BUF1 (N10151, N10134);
and AND3 (N10152, N10141, N2236, N6767);
xor XOR2 (N10153, N10149, N5655);
nor NOR2 (N10154, N10151, N9314);
nand NAND2 (N10155, N10143, N5012);
buf BUF1 (N10156, N10147);
nor NOR2 (N10157, N10150, N4727);
buf BUF1 (N10158, N10154);
xor XOR2 (N10159, N10153, N469);
and AND3 (N10160, N10128, N7, N407);
buf BUF1 (N10161, N10148);
or OR2 (N10162, N10161, N5868);
not NOT1 (N10163, N10160);
or OR4 (N10164, N10152, N10024, N5618, N9679);
not NOT1 (N10165, N10162);
nor NOR4 (N10166, N10131, N1941, N8993, N4825);
not NOT1 (N10167, N10156);
not NOT1 (N10168, N10155);
buf BUF1 (N10169, N10140);
xor XOR2 (N10170, N10163, N5898);
buf BUF1 (N10171, N10166);
buf BUF1 (N10172, N10167);
nand NAND2 (N10173, N10172, N3803);
xor XOR2 (N10174, N10173, N4124);
nand NAND3 (N10175, N10164, N5912, N6192);
buf BUF1 (N10176, N10171);
and AND2 (N10177, N10175, N1470);
nor NOR4 (N10178, N10176, N9852, N4130, N8128);
buf BUF1 (N10179, N10177);
nor NOR4 (N10180, N10179, N4794, N6093, N3024);
nor NOR4 (N10181, N10158, N9709, N2546, N2434);
buf BUF1 (N10182, N10168);
nand NAND2 (N10183, N10157, N7524);
buf BUF1 (N10184, N10180);
xor XOR2 (N10185, N10181, N7493);
not NOT1 (N10186, N10184);
nor NOR3 (N10187, N10182, N1491, N7085);
nand NAND4 (N10188, N10187, N199, N5805, N496);
and AND2 (N10189, N10165, N4066);
nor NOR3 (N10190, N10188, N1005, N2855);
nand NAND2 (N10191, N10186, N8971);
xor XOR2 (N10192, N10183, N7969);
buf BUF1 (N10193, N10185);
or OR3 (N10194, N10193, N4290, N2001);
xor XOR2 (N10195, N10170, N791);
or OR2 (N10196, N10195, N8161);
xor XOR2 (N10197, N10191, N6234);
not NOT1 (N10198, N10197);
buf BUF1 (N10199, N10159);
or OR3 (N10200, N10178, N7248, N7006);
xor XOR2 (N10201, N10169, N7288);
or OR2 (N10202, N10199, N5467);
nand NAND4 (N10203, N10198, N5316, N2207, N5128);
not NOT1 (N10204, N10190);
not NOT1 (N10205, N10204);
buf BUF1 (N10206, N10200);
xor XOR2 (N10207, N10174, N9209);
and AND2 (N10208, N10192, N1627);
or OR2 (N10209, N10189, N4431);
or OR2 (N10210, N10208, N9380);
and AND2 (N10211, N10194, N8934);
buf BUF1 (N10212, N10211);
or OR4 (N10213, N10203, N1119, N6159, N8931);
or OR2 (N10214, N10209, N1738);
not NOT1 (N10215, N10213);
not NOT1 (N10216, N10206);
nand NAND4 (N10217, N10196, N9920, N4655, N6453);
not NOT1 (N10218, N10215);
nor NOR4 (N10219, N10202, N5945, N9507, N7146);
or OR3 (N10220, N10214, N5358, N4538);
and AND3 (N10221, N10218, N5992, N9722);
buf BUF1 (N10222, N10201);
or OR2 (N10223, N10207, N4751);
not NOT1 (N10224, N10217);
nand NAND4 (N10225, N10220, N8073, N9452, N5965);
xor XOR2 (N10226, N10224, N479);
not NOT1 (N10227, N10210);
nand NAND3 (N10228, N10219, N9799, N8367);
nand NAND4 (N10229, N10227, N8434, N680, N1466);
buf BUF1 (N10230, N10212);
nor NOR4 (N10231, N10228, N4033, N483, N4602);
xor XOR2 (N10232, N10223, N4698);
not NOT1 (N10233, N10230);
buf BUF1 (N10234, N10232);
not NOT1 (N10235, N10233);
not NOT1 (N10236, N10231);
nor NOR2 (N10237, N10225, N6734);
nand NAND4 (N10238, N10205, N6296, N4716, N5080);
buf BUF1 (N10239, N10216);
nor NOR2 (N10240, N10229, N2379);
buf BUF1 (N10241, N10240);
xor XOR2 (N10242, N10234, N2820);
buf BUF1 (N10243, N10241);
or OR2 (N10244, N10239, N4003);
nand NAND4 (N10245, N10226, N8378, N7760, N3445);
and AND2 (N10246, N10243, N6336);
nor NOR3 (N10247, N10222, N2432, N7730);
nor NOR4 (N10248, N10244, N2061, N7245, N8954);
buf BUF1 (N10249, N10246);
and AND2 (N10250, N10235, N8256);
nand NAND2 (N10251, N10245, N4681);
nand NAND3 (N10252, N10242, N8206, N1397);
or OR4 (N10253, N10237, N7893, N3177, N8128);
not NOT1 (N10254, N10238);
or OR2 (N10255, N10252, N4902);
and AND4 (N10256, N10221, N7012, N1060, N5224);
nand NAND4 (N10257, N10255, N1193, N3277, N903);
nor NOR4 (N10258, N10248, N2910, N3378, N1665);
buf BUF1 (N10259, N10247);
not NOT1 (N10260, N10253);
xor XOR2 (N10261, N10250, N3896);
buf BUF1 (N10262, N10256);
not NOT1 (N10263, N10251);
and AND2 (N10264, N10263, N49);
xor XOR2 (N10265, N10259, N4742);
not NOT1 (N10266, N10249);
xor XOR2 (N10267, N10262, N545);
xor XOR2 (N10268, N10258, N8765);
buf BUF1 (N10269, N10260);
nor NOR3 (N10270, N10268, N9268, N9440);
nand NAND3 (N10271, N10270, N9192, N3573);
and AND3 (N10272, N10271, N2447, N8236);
nand NAND2 (N10273, N10261, N1383);
nand NAND3 (N10274, N10269, N3120, N4644);
not NOT1 (N10275, N10257);
xor XOR2 (N10276, N10254, N3586);
buf BUF1 (N10277, N10266);
and AND2 (N10278, N10277, N2799);
nand NAND4 (N10279, N10275, N4419, N7583, N9015);
or OR2 (N10280, N10236, N7260);
nor NOR2 (N10281, N10265, N7127);
not NOT1 (N10282, N10273);
or OR2 (N10283, N10282, N6013);
not NOT1 (N10284, N10283);
nor NOR3 (N10285, N10284, N5742, N3177);
or OR4 (N10286, N10267, N8882, N4466, N1010);
not NOT1 (N10287, N10272);
xor XOR2 (N10288, N10286, N2829);
buf BUF1 (N10289, N10280);
and AND4 (N10290, N10289, N8989, N3882, N8746);
buf BUF1 (N10291, N10288);
not NOT1 (N10292, N10264);
or OR2 (N10293, N10291, N2338);
buf BUF1 (N10294, N10293);
nand NAND2 (N10295, N10276, N4769);
xor XOR2 (N10296, N10295, N4590);
xor XOR2 (N10297, N10281, N7392);
buf BUF1 (N10298, N10274);
and AND2 (N10299, N10297, N1473);
and AND2 (N10300, N10279, N8747);
and AND4 (N10301, N10299, N8289, N6350, N4388);
xor XOR2 (N10302, N10296, N5575);
xor XOR2 (N10303, N10301, N961);
nand NAND3 (N10304, N10290, N3657, N6981);
and AND4 (N10305, N10304, N9240, N3324, N1622);
nand NAND2 (N10306, N10305, N1781);
buf BUF1 (N10307, N10278);
not NOT1 (N10308, N10302);
not NOT1 (N10309, N10306);
nand NAND4 (N10310, N10285, N4102, N3177, N2366);
buf BUF1 (N10311, N10308);
and AND3 (N10312, N10292, N1383, N441);
or OR3 (N10313, N10307, N4577, N8832);
nor NOR3 (N10314, N10294, N56, N715);
or OR2 (N10315, N10313, N2643);
buf BUF1 (N10316, N10287);
nand NAND2 (N10317, N10303, N3111);
buf BUF1 (N10318, N10309);
xor XOR2 (N10319, N10318, N1639);
or OR2 (N10320, N10300, N4514);
not NOT1 (N10321, N10312);
and AND2 (N10322, N10310, N8105);
buf BUF1 (N10323, N10311);
buf BUF1 (N10324, N10322);
and AND2 (N10325, N10317, N3752);
nand NAND3 (N10326, N10323, N1935, N5964);
or OR2 (N10327, N10321, N2744);
and AND3 (N10328, N10320, N5134, N1604);
or OR4 (N10329, N10326, N7248, N365, N8204);
xor XOR2 (N10330, N10327, N7808);
and AND4 (N10331, N10325, N9655, N2039, N7347);
xor XOR2 (N10332, N10328, N4316);
not NOT1 (N10333, N10316);
or OR3 (N10334, N10324, N1071, N9757);
nor NOR4 (N10335, N10332, N7191, N6502, N9170);
or OR4 (N10336, N10314, N6955, N8150, N4251);
nand NAND2 (N10337, N10319, N4047);
or OR2 (N10338, N10335, N9483);
not NOT1 (N10339, N10333);
not NOT1 (N10340, N10331);
buf BUF1 (N10341, N10334);
or OR3 (N10342, N10329, N2506, N2099);
buf BUF1 (N10343, N10339);
nand NAND4 (N10344, N10315, N1944, N9838, N5957);
or OR4 (N10345, N10330, N1315, N7432, N3725);
buf BUF1 (N10346, N10338);
or OR4 (N10347, N10298, N10321, N3513, N82);
nand NAND4 (N10348, N10342, N9603, N3340, N8192);
and AND2 (N10349, N10344, N5242);
buf BUF1 (N10350, N10336);
xor XOR2 (N10351, N10340, N2272);
buf BUF1 (N10352, N10349);
nor NOR2 (N10353, N10347, N5769);
not NOT1 (N10354, N10337);
buf BUF1 (N10355, N10353);
or OR4 (N10356, N10350, N7740, N6185, N9445);
buf BUF1 (N10357, N10351);
xor XOR2 (N10358, N10343, N1430);
and AND3 (N10359, N10358, N1414, N6257);
nand NAND3 (N10360, N10356, N5989, N7);
nand NAND2 (N10361, N10354, N5674);
buf BUF1 (N10362, N10361);
not NOT1 (N10363, N10355);
and AND4 (N10364, N10357, N5586, N1922, N8337);
nor NOR2 (N10365, N10352, N8396);
not NOT1 (N10366, N10360);
not NOT1 (N10367, N10366);
buf BUF1 (N10368, N10365);
xor XOR2 (N10369, N10341, N3264);
and AND2 (N10370, N10368, N3227);
and AND4 (N10371, N10367, N2129, N3824, N1879);
buf BUF1 (N10372, N10364);
xor XOR2 (N10373, N10362, N293);
or OR2 (N10374, N10348, N8002);
or OR2 (N10375, N10359, N4317);
buf BUF1 (N10376, N10374);
nand NAND2 (N10377, N10372, N7696);
nor NOR3 (N10378, N10377, N7765, N795);
buf BUF1 (N10379, N10371);
or OR4 (N10380, N10373, N5801, N6617, N8935);
and AND4 (N10381, N10345, N3493, N6432, N3203);
and AND2 (N10382, N10370, N3133);
not NOT1 (N10383, N10369);
xor XOR2 (N10384, N10380, N9386);
buf BUF1 (N10385, N10375);
or OR4 (N10386, N10378, N1915, N985, N9358);
xor XOR2 (N10387, N10382, N6499);
nor NOR2 (N10388, N10346, N394);
or OR2 (N10389, N10376, N4096);
and AND3 (N10390, N10388, N8424, N1847);
or OR4 (N10391, N10379, N6652, N1380, N3689);
buf BUF1 (N10392, N10381);
xor XOR2 (N10393, N10392, N7915);
nand NAND4 (N10394, N10391, N6456, N7572, N2494);
or OR2 (N10395, N10393, N4866);
or OR3 (N10396, N10363, N8799, N4696);
and AND3 (N10397, N10390, N678, N8788);
and AND3 (N10398, N10389, N1124, N1168);
xor XOR2 (N10399, N10398, N8205);
and AND4 (N10400, N10395, N4380, N5492, N2072);
nand NAND3 (N10401, N10383, N9345, N4674);
nand NAND2 (N10402, N10400, N2917);
or OR2 (N10403, N10385, N7424);
buf BUF1 (N10404, N10394);
not NOT1 (N10405, N10399);
or OR4 (N10406, N10404, N3212, N7602, N9162);
nand NAND4 (N10407, N10396, N8192, N6217, N9975);
xor XOR2 (N10408, N10402, N5624);
buf BUF1 (N10409, N10387);
buf BUF1 (N10410, N10408);
not NOT1 (N10411, N10405);
xor XOR2 (N10412, N10406, N5536);
not NOT1 (N10413, N10409);
not NOT1 (N10414, N10397);
nor NOR4 (N10415, N10407, N10165, N6691, N2546);
xor XOR2 (N10416, N10384, N6652);
or OR2 (N10417, N10411, N4355);
or OR4 (N10418, N10410, N3064, N9475, N10034);
nand NAND2 (N10419, N10403, N7613);
buf BUF1 (N10420, N10414);
nand NAND2 (N10421, N10420, N2082);
or OR3 (N10422, N10415, N10153, N672);
and AND4 (N10423, N10419, N942, N9703, N7108);
not NOT1 (N10424, N10416);
buf BUF1 (N10425, N10423);
not NOT1 (N10426, N10417);
and AND2 (N10427, N10422, N6014);
not NOT1 (N10428, N10425);
and AND3 (N10429, N10426, N3269, N4378);
nor NOR3 (N10430, N10424, N2730, N4021);
nor NOR4 (N10431, N10421, N3997, N3723, N6989);
nand NAND4 (N10432, N10418, N1942, N3791, N1825);
nand NAND4 (N10433, N10431, N3055, N3302, N7154);
buf BUF1 (N10434, N10412);
nor NOR3 (N10435, N10401, N6003, N4260);
and AND4 (N10436, N10413, N545, N3794, N6979);
and AND2 (N10437, N10433, N2066);
xor XOR2 (N10438, N10430, N380);
nor NOR2 (N10439, N10386, N5299);
or OR3 (N10440, N10434, N4760, N6359);
and AND3 (N10441, N10432, N6616, N8057);
and AND4 (N10442, N10438, N10034, N2808, N4870);
xor XOR2 (N10443, N10442, N2406);
or OR3 (N10444, N10436, N8177, N5237);
not NOT1 (N10445, N10439);
and AND4 (N10446, N10435, N2982, N10160, N7631);
not NOT1 (N10447, N10437);
and AND2 (N10448, N10441, N5358);
buf BUF1 (N10449, N10428);
buf BUF1 (N10450, N10445);
nor NOR4 (N10451, N10444, N2723, N119, N5441);
buf BUF1 (N10452, N10443);
nand NAND3 (N10453, N10447, N434, N10377);
nand NAND3 (N10454, N10449, N3356, N3613);
or OR4 (N10455, N10427, N10006, N3115, N9047);
not NOT1 (N10456, N10446);
and AND2 (N10457, N10456, N5569);
nor NOR2 (N10458, N10454, N7755);
buf BUF1 (N10459, N10458);
and AND3 (N10460, N10448, N1838, N6209);
buf BUF1 (N10461, N10457);
nor NOR4 (N10462, N10459, N4141, N4146, N5144);
not NOT1 (N10463, N10461);
or OR2 (N10464, N10451, N9277);
and AND3 (N10465, N10463, N383, N9691);
xor XOR2 (N10466, N10460, N9260);
and AND3 (N10467, N10462, N2770, N10330);
nand NAND4 (N10468, N10453, N5082, N9409, N2083);
buf BUF1 (N10469, N10464);
nor NOR3 (N10470, N10452, N1902, N7733);
or OR4 (N10471, N10455, N10361, N4953, N3236);
buf BUF1 (N10472, N10450);
nor NOR2 (N10473, N10472, N7414);
or OR2 (N10474, N10468, N7888);
buf BUF1 (N10475, N10466);
xor XOR2 (N10476, N10429, N8900);
nand NAND3 (N10477, N10474, N8634, N6836);
or OR2 (N10478, N10440, N5913);
nor NOR3 (N10479, N10470, N3041, N7167);
not NOT1 (N10480, N10467);
nand NAND3 (N10481, N10476, N9568, N6626);
nand NAND2 (N10482, N10480, N7411);
nor NOR2 (N10483, N10481, N5574);
nor NOR2 (N10484, N10477, N8733);
or OR3 (N10485, N10478, N2433, N8762);
buf BUF1 (N10486, N10484);
not NOT1 (N10487, N10479);
nor NOR3 (N10488, N10465, N2425, N9327);
xor XOR2 (N10489, N10487, N9191);
nor NOR2 (N10490, N10485, N1570);
and AND4 (N10491, N10488, N4988, N5652, N6758);
not NOT1 (N10492, N10473);
buf BUF1 (N10493, N10471);
buf BUF1 (N10494, N10491);
not NOT1 (N10495, N10492);
or OR4 (N10496, N10475, N10020, N9413, N1577);
not NOT1 (N10497, N10469);
not NOT1 (N10498, N10489);
not NOT1 (N10499, N10495);
not NOT1 (N10500, N10490);
not NOT1 (N10501, N10493);
xor XOR2 (N10502, N10499, N7346);
not NOT1 (N10503, N10496);
nand NAND2 (N10504, N10482, N1197);
not NOT1 (N10505, N10497);
nand NAND4 (N10506, N10503, N6216, N9744, N4100);
buf BUF1 (N10507, N10494);
xor XOR2 (N10508, N10505, N4588);
buf BUF1 (N10509, N10486);
nand NAND3 (N10510, N10501, N5727, N8702);
nand NAND3 (N10511, N10508, N7632, N3568);
nand NAND3 (N10512, N10498, N7053, N8838);
nand NAND3 (N10513, N10511, N6526, N7892);
xor XOR2 (N10514, N10510, N10367);
not NOT1 (N10515, N10506);
buf BUF1 (N10516, N10512);
or OR3 (N10517, N10509, N585, N9728);
not NOT1 (N10518, N10504);
or OR3 (N10519, N10483, N9317, N3987);
and AND2 (N10520, N10502, N5734);
buf BUF1 (N10521, N10517);
xor XOR2 (N10522, N10514, N9694);
not NOT1 (N10523, N10519);
xor XOR2 (N10524, N10516, N7358);
not NOT1 (N10525, N10520);
or OR2 (N10526, N10522, N9456);
not NOT1 (N10527, N10521);
buf BUF1 (N10528, N10526);
or OR4 (N10529, N10525, N7412, N272, N7790);
buf BUF1 (N10530, N10529);
xor XOR2 (N10531, N10507, N4668);
nor NOR3 (N10532, N10515, N1865, N9607);
buf BUF1 (N10533, N10518);
and AND3 (N10534, N10524, N6909, N5658);
or OR2 (N10535, N10532, N9137);
nand NAND4 (N10536, N10533, N2739, N578, N9308);
xor XOR2 (N10537, N10530, N6319);
nand NAND4 (N10538, N10531, N10294, N966, N1168);
and AND2 (N10539, N10528, N3516);
not NOT1 (N10540, N10537);
and AND2 (N10541, N10534, N2720);
buf BUF1 (N10542, N10540);
buf BUF1 (N10543, N10513);
not NOT1 (N10544, N10538);
xor XOR2 (N10545, N10543, N10046);
or OR4 (N10546, N10539, N2760, N8657, N9150);
xor XOR2 (N10547, N10523, N2828);
nor NOR2 (N10548, N10536, N8549);
not NOT1 (N10549, N10500);
not NOT1 (N10550, N10548);
nand NAND2 (N10551, N10546, N9135);
not NOT1 (N10552, N10551);
and AND2 (N10553, N10541, N7276);
nor NOR4 (N10554, N10544, N4821, N2221, N8092);
buf BUF1 (N10555, N10554);
not NOT1 (N10556, N10555);
or OR2 (N10557, N10535, N5358);
and AND3 (N10558, N10542, N4429, N1852);
nand NAND3 (N10559, N10527, N9439, N7814);
or OR2 (N10560, N10556, N8906);
and AND2 (N10561, N10557, N7603);
or OR3 (N10562, N10547, N6819, N7544);
or OR2 (N10563, N10559, N152);
nand NAND3 (N10564, N10563, N10038, N3728);
xor XOR2 (N10565, N10561, N6245);
not NOT1 (N10566, N10553);
xor XOR2 (N10567, N10562, N9947);
nand NAND3 (N10568, N10565, N1578, N10531);
xor XOR2 (N10569, N10567, N3018);
or OR4 (N10570, N10552, N3356, N8687, N3211);
xor XOR2 (N10571, N10564, N10420);
and AND2 (N10572, N10558, N5249);
xor XOR2 (N10573, N10569, N8111);
nor NOR3 (N10574, N10550, N7674, N2071);
buf BUF1 (N10575, N10572);
buf BUF1 (N10576, N10568);
not NOT1 (N10577, N10549);
xor XOR2 (N10578, N10574, N273);
nand NAND2 (N10579, N10566, N3906);
not NOT1 (N10580, N10575);
or OR4 (N10581, N10576, N6750, N8718, N6796);
nor NOR3 (N10582, N10577, N309, N4706);
or OR4 (N10583, N10582, N4270, N6254, N5576);
not NOT1 (N10584, N10583);
and AND3 (N10585, N10579, N1820, N2366);
nor NOR2 (N10586, N10578, N10501);
or OR2 (N10587, N10580, N122);
or OR4 (N10588, N10585, N7915, N4808, N9827);
or OR3 (N10589, N10573, N103, N2867);
and AND4 (N10590, N10588, N6535, N8387, N1908);
nand NAND2 (N10591, N10571, N4917);
or OR4 (N10592, N10545, N693, N668, N2692);
or OR2 (N10593, N10584, N2171);
nand NAND3 (N10594, N10592, N3317, N6197);
and AND4 (N10595, N10587, N8003, N5265, N2723);
and AND3 (N10596, N10591, N1417, N6124);
nor NOR2 (N10597, N10586, N5738);
or OR3 (N10598, N10594, N9425, N5312);
and AND2 (N10599, N10570, N6322);
and AND3 (N10600, N10597, N5959, N10025);
or OR2 (N10601, N10593, N2495);
buf BUF1 (N10602, N10596);
buf BUF1 (N10603, N10599);
and AND2 (N10604, N10590, N8800);
buf BUF1 (N10605, N10604);
nor NOR2 (N10606, N10560, N668);
or OR2 (N10607, N10598, N2525);
nor NOR3 (N10608, N10607, N8375, N2080);
buf BUF1 (N10609, N10595);
xor XOR2 (N10610, N10606, N8769);
not NOT1 (N10611, N10581);
xor XOR2 (N10612, N10589, N6089);
xor XOR2 (N10613, N10601, N2460);
buf BUF1 (N10614, N10608);
not NOT1 (N10615, N10603);
buf BUF1 (N10616, N10614);
nor NOR4 (N10617, N10605, N4138, N3565, N2914);
buf BUF1 (N10618, N10613);
or OR3 (N10619, N10602, N7300, N89);
and AND2 (N10620, N10615, N9041);
and AND3 (N10621, N10609, N66, N553);
nor NOR2 (N10622, N10620, N6569);
nor NOR3 (N10623, N10622, N8729, N8411);
or OR2 (N10624, N10619, N2795);
xor XOR2 (N10625, N10611, N9554);
nor NOR2 (N10626, N10610, N6158);
nand NAND4 (N10627, N10616, N6542, N373, N3910);
or OR3 (N10628, N10625, N4857, N8613);
nand NAND3 (N10629, N10618, N7304, N352);
and AND3 (N10630, N10626, N3476, N10196);
buf BUF1 (N10631, N10630);
and AND4 (N10632, N10612, N10008, N8152, N1283);
or OR4 (N10633, N10623, N8447, N3392, N9866);
and AND2 (N10634, N10627, N835);
nand NAND2 (N10635, N10629, N3762);
buf BUF1 (N10636, N10633);
not NOT1 (N10637, N10636);
not NOT1 (N10638, N10624);
xor XOR2 (N10639, N10634, N7281);
and AND3 (N10640, N10637, N10268, N3349);
and AND3 (N10641, N10638, N2050, N119);
xor XOR2 (N10642, N10600, N4413);
nor NOR4 (N10643, N10632, N952, N5095, N10044);
not NOT1 (N10644, N10640);
or OR3 (N10645, N10642, N9269, N8051);
not NOT1 (N10646, N10641);
nor NOR2 (N10647, N10628, N3109);
or OR2 (N10648, N10621, N2649);
xor XOR2 (N10649, N10617, N3526);
not NOT1 (N10650, N10644);
not NOT1 (N10651, N10639);
or OR2 (N10652, N10650, N5807);
or OR3 (N10653, N10646, N3951, N2377);
or OR3 (N10654, N10652, N4087, N9498);
and AND2 (N10655, N10645, N917);
xor XOR2 (N10656, N10654, N7343);
nor NOR2 (N10657, N10653, N4147);
nand NAND3 (N10658, N10651, N7110, N7343);
and AND2 (N10659, N10647, N3312);
nor NOR4 (N10660, N10631, N4816, N2902, N10313);
buf BUF1 (N10661, N10655);
or OR2 (N10662, N10643, N372);
nor NOR4 (N10663, N10660, N6404, N9236, N237);
nor NOR3 (N10664, N10635, N8309, N3475);
or OR3 (N10665, N10648, N3363, N2502);
xor XOR2 (N10666, N10663, N1042);
nand NAND2 (N10667, N10662, N8858);
nand NAND4 (N10668, N10665, N5313, N4790, N5249);
and AND3 (N10669, N10664, N4721, N4900);
and AND3 (N10670, N10649, N656, N4142);
xor XOR2 (N10671, N10669, N3712);
xor XOR2 (N10672, N10667, N8361);
nor NOR2 (N10673, N10661, N9907);
not NOT1 (N10674, N10672);
and AND2 (N10675, N10659, N5249);
not NOT1 (N10676, N10674);
nor NOR4 (N10677, N10657, N2304, N7079, N1750);
buf BUF1 (N10678, N10676);
or OR2 (N10679, N10675, N6411);
nand NAND2 (N10680, N10673, N5431);
nand NAND3 (N10681, N10658, N8268, N6011);
xor XOR2 (N10682, N10677, N7833);
xor XOR2 (N10683, N10678, N8142);
nor NOR4 (N10684, N10668, N1194, N1434, N4294);
nor NOR2 (N10685, N10682, N2334);
buf BUF1 (N10686, N10680);
nand NAND3 (N10687, N10656, N6483, N1111);
nor NOR4 (N10688, N10666, N399, N8868, N5149);
not NOT1 (N10689, N10670);
not NOT1 (N10690, N10689);
nor NOR2 (N10691, N10683, N2249);
or OR2 (N10692, N10684, N4610);
and AND2 (N10693, N10671, N674);
nor NOR3 (N10694, N10685, N9530, N4437);
nand NAND3 (N10695, N10679, N294, N9868);
or OR4 (N10696, N10695, N3124, N5324, N9661);
or OR4 (N10697, N10687, N338, N2250, N6187);
nor NOR4 (N10698, N10697, N4088, N7134, N9542);
xor XOR2 (N10699, N10681, N709);
nand NAND4 (N10700, N10699, N6298, N2483, N8228);
nand NAND2 (N10701, N10693, N3694);
nor NOR2 (N10702, N10700, N1993);
and AND3 (N10703, N10701, N2274, N5644);
not NOT1 (N10704, N10698);
and AND3 (N10705, N10704, N6309, N7338);
not NOT1 (N10706, N10696);
and AND2 (N10707, N10690, N4091);
nand NAND2 (N10708, N10707, N5734);
xor XOR2 (N10709, N10702, N4253);
nor NOR3 (N10710, N10703, N1158, N9242);
buf BUF1 (N10711, N10691);
buf BUF1 (N10712, N10694);
not NOT1 (N10713, N10706);
and AND4 (N10714, N10686, N9818, N1105, N1895);
and AND3 (N10715, N10709, N3338, N4989);
not NOT1 (N10716, N10712);
buf BUF1 (N10717, N10692);
nand NAND2 (N10718, N10705, N1765);
or OR3 (N10719, N10710, N4984, N222);
not NOT1 (N10720, N10716);
buf BUF1 (N10721, N10708);
and AND2 (N10722, N10718, N6217);
or OR2 (N10723, N10717, N5143);
xor XOR2 (N10724, N10711, N8718);
and AND2 (N10725, N10688, N4510);
nand NAND2 (N10726, N10722, N9986);
or OR4 (N10727, N10713, N545, N9332, N9686);
nor NOR4 (N10728, N10714, N5273, N6124, N6960);
and AND4 (N10729, N10715, N5911, N2806, N5950);
nand NAND2 (N10730, N10723, N5197);
and AND2 (N10731, N10720, N8218);
nand NAND4 (N10732, N10729, N8034, N8924, N1838);
xor XOR2 (N10733, N10725, N8193);
buf BUF1 (N10734, N10726);
buf BUF1 (N10735, N10721);
buf BUF1 (N10736, N10734);
xor XOR2 (N10737, N10731, N4068);
nand NAND4 (N10738, N10735, N10374, N62, N9704);
nor NOR4 (N10739, N10733, N9200, N10015, N10539);
or OR3 (N10740, N10739, N10446, N9699);
xor XOR2 (N10741, N10727, N3227);
nor NOR4 (N10742, N10741, N2697, N4064, N3700);
buf BUF1 (N10743, N10738);
nor NOR4 (N10744, N10737, N8402, N8084, N8070);
nand NAND4 (N10745, N10719, N8426, N1426, N463);
or OR2 (N10746, N10732, N6070);
xor XOR2 (N10747, N10740, N9976);
or OR3 (N10748, N10747, N8376, N5774);
or OR2 (N10749, N10743, N2584);
and AND3 (N10750, N10728, N8823, N4058);
and AND2 (N10751, N10744, N5757);
nand NAND3 (N10752, N10746, N5010, N10462);
and AND2 (N10753, N10750, N9612);
nand NAND3 (N10754, N10724, N9557, N7688);
xor XOR2 (N10755, N10745, N5996);
and AND3 (N10756, N10753, N9489, N2006);
buf BUF1 (N10757, N10754);
buf BUF1 (N10758, N10730);
xor XOR2 (N10759, N10755, N5674);
nand NAND4 (N10760, N10758, N5224, N8271, N2206);
nand NAND4 (N10761, N10760, N1502, N2685, N6382);
buf BUF1 (N10762, N10748);
or OR2 (N10763, N10759, N1615);
buf BUF1 (N10764, N10761);
and AND3 (N10765, N10764, N9226, N10673);
and AND2 (N10766, N10765, N8972);
and AND4 (N10767, N10762, N2287, N2327, N1376);
nor NOR4 (N10768, N10767, N7683, N5439, N721);
buf BUF1 (N10769, N10756);
xor XOR2 (N10770, N10749, N10450);
and AND4 (N10771, N10742, N1928, N6231, N8038);
buf BUF1 (N10772, N10763);
buf BUF1 (N10773, N10757);
not NOT1 (N10774, N10769);
xor XOR2 (N10775, N10770, N5829);
xor XOR2 (N10776, N10752, N7298);
xor XOR2 (N10777, N10775, N602);
xor XOR2 (N10778, N10736, N7182);
nand NAND4 (N10779, N10774, N8516, N2541, N845);
nand NAND3 (N10780, N10771, N5425, N3269);
buf BUF1 (N10781, N10777);
nor NOR3 (N10782, N10779, N9474, N853);
not NOT1 (N10783, N10781);
nand NAND4 (N10784, N10783, N769, N410, N9968);
xor XOR2 (N10785, N10776, N8839);
xor XOR2 (N10786, N10751, N3546);
and AND3 (N10787, N10768, N6599, N6647);
not NOT1 (N10788, N10784);
not NOT1 (N10789, N10782);
nand NAND2 (N10790, N10772, N6344);
and AND2 (N10791, N10787, N536);
nand NAND3 (N10792, N10766, N9299, N9763);
not NOT1 (N10793, N10786);
and AND2 (N10794, N10785, N8765);
or OR2 (N10795, N10794, N5824);
nand NAND2 (N10796, N10778, N4690);
nand NAND2 (N10797, N10780, N5681);
not NOT1 (N10798, N10797);
buf BUF1 (N10799, N10773);
and AND3 (N10800, N10789, N1037, N7993);
buf BUF1 (N10801, N10800);
or OR3 (N10802, N10788, N10104, N2188);
xor XOR2 (N10803, N10801, N469);
or OR4 (N10804, N10803, N9917, N6616, N7362);
xor XOR2 (N10805, N10790, N8402);
xor XOR2 (N10806, N10796, N2094);
nor NOR4 (N10807, N10806, N5666, N2943, N2867);
buf BUF1 (N10808, N10793);
nor NOR3 (N10809, N10795, N9421, N2329);
buf BUF1 (N10810, N10791);
buf BUF1 (N10811, N10810);
nand NAND3 (N10812, N10809, N1633, N1604);
or OR3 (N10813, N10792, N6655, N5184);
xor XOR2 (N10814, N10813, N10623);
nand NAND4 (N10815, N10812, N10433, N9950, N135);
and AND3 (N10816, N10802, N1977, N5693);
and AND2 (N10817, N10814, N8004);
nand NAND2 (N10818, N10816, N3765);
xor XOR2 (N10819, N10807, N9327);
nor NOR2 (N10820, N10818, N5869);
buf BUF1 (N10821, N10798);
nor NOR2 (N10822, N10817, N2835);
nand NAND4 (N10823, N10819, N4148, N2483, N10496);
nor NOR3 (N10824, N10823, N5394, N327);
buf BUF1 (N10825, N10804);
and AND2 (N10826, N10825, N1427);
nand NAND4 (N10827, N10811, N8683, N9068, N9842);
buf BUF1 (N10828, N10821);
or OR2 (N10829, N10826, N1479);
xor XOR2 (N10830, N10822, N9145);
not NOT1 (N10831, N10824);
buf BUF1 (N10832, N10828);
nand NAND3 (N10833, N10805, N4143, N10200);
xor XOR2 (N10834, N10827, N2566);
xor XOR2 (N10835, N10831, N4719);
not NOT1 (N10836, N10830);
and AND2 (N10837, N10832, N8697);
not NOT1 (N10838, N10829);
buf BUF1 (N10839, N10838);
xor XOR2 (N10840, N10835, N9797);
not NOT1 (N10841, N10836);
nand NAND3 (N10842, N10840, N10057, N2099);
nand NAND3 (N10843, N10815, N7262, N6018);
not NOT1 (N10844, N10834);
buf BUF1 (N10845, N10820);
nor NOR3 (N10846, N10842, N3796, N815);
xor XOR2 (N10847, N10837, N3676);
nand NAND3 (N10848, N10841, N7453, N2402);
and AND2 (N10849, N10846, N8981);
not NOT1 (N10850, N10843);
nand NAND4 (N10851, N10839, N5404, N8831, N321);
not NOT1 (N10852, N10847);
xor XOR2 (N10853, N10852, N9612);
or OR3 (N10854, N10808, N7140, N7721);
buf BUF1 (N10855, N10849);
and AND3 (N10856, N10854, N7959, N5889);
or OR2 (N10857, N10848, N9373);
nor NOR3 (N10858, N10833, N10336, N8679);
not NOT1 (N10859, N10857);
or OR4 (N10860, N10859, N4475, N10372, N3726);
not NOT1 (N10861, N10844);
and AND4 (N10862, N10855, N5225, N678, N9701);
not NOT1 (N10863, N10860);
buf BUF1 (N10864, N10799);
or OR4 (N10865, N10850, N1893, N290, N4634);
nor NOR2 (N10866, N10853, N10861);
xor XOR2 (N10867, N8422, N2311);
nand NAND4 (N10868, N10865, N10434, N2707, N6237);
buf BUF1 (N10869, N10856);
not NOT1 (N10870, N10866);
and AND2 (N10871, N10863, N8311);
not NOT1 (N10872, N10845);
nand NAND3 (N10873, N10858, N1050, N3773);
not NOT1 (N10874, N10872);
and AND3 (N10875, N10873, N3719, N8760);
not NOT1 (N10876, N10862);
not NOT1 (N10877, N10868);
buf BUF1 (N10878, N10870);
and AND3 (N10879, N10864, N9934, N2138);
or OR3 (N10880, N10851, N1713, N1490);
and AND4 (N10881, N10876, N10671, N10880, N8503);
buf BUF1 (N10882, N3955);
and AND3 (N10883, N10874, N1523, N1387);
xor XOR2 (N10884, N10877, N6292);
buf BUF1 (N10885, N10875);
not NOT1 (N10886, N10884);
or OR2 (N10887, N10878, N9669);
not NOT1 (N10888, N10885);
xor XOR2 (N10889, N10867, N5558);
or OR4 (N10890, N10886, N2840, N2761, N10410);
and AND2 (N10891, N10883, N4962);
or OR4 (N10892, N10879, N6034, N7041, N8979);
nor NOR3 (N10893, N10891, N5799, N9305);
buf BUF1 (N10894, N10881);
not NOT1 (N10895, N10894);
xor XOR2 (N10896, N10893, N2992);
not NOT1 (N10897, N10889);
xor XOR2 (N10898, N10871, N2934);
nor NOR2 (N10899, N10869, N6016);
or OR4 (N10900, N10895, N2456, N10567, N5855);
nand NAND3 (N10901, N10899, N8521, N2130);
not NOT1 (N10902, N10882);
xor XOR2 (N10903, N10888, N3951);
nor NOR2 (N10904, N10903, N5737);
and AND2 (N10905, N10897, N6121);
buf BUF1 (N10906, N10902);
not NOT1 (N10907, N10896);
or OR3 (N10908, N10905, N8882, N2574);
xor XOR2 (N10909, N10892, N78);
not NOT1 (N10910, N10904);
buf BUF1 (N10911, N10906);
nand NAND2 (N10912, N10890, N9953);
or OR2 (N10913, N10909, N2040);
buf BUF1 (N10914, N10913);
and AND3 (N10915, N10887, N7179, N1293);
nand NAND4 (N10916, N10898, N7792, N4893, N7971);
or OR2 (N10917, N10912, N3502);
nand NAND2 (N10918, N10901, N1578);
buf BUF1 (N10919, N10910);
nand NAND2 (N10920, N10914, N8293);
buf BUF1 (N10921, N10917);
buf BUF1 (N10922, N10916);
xor XOR2 (N10923, N10918, N2782);
not NOT1 (N10924, N10907);
xor XOR2 (N10925, N10915, N486);
and AND3 (N10926, N10925, N4326, N9902);
not NOT1 (N10927, N10926);
or OR2 (N10928, N10911, N9025);
or OR2 (N10929, N10922, N2221);
and AND3 (N10930, N10921, N5778, N7975);
xor XOR2 (N10931, N10929, N5700);
xor XOR2 (N10932, N10927, N6182);
nor NOR4 (N10933, N10908, N22, N5997, N3544);
and AND3 (N10934, N10930, N9452, N2316);
nor NOR4 (N10935, N10924, N2156, N4113, N4999);
xor XOR2 (N10936, N10932, N4328);
not NOT1 (N10937, N10936);
buf BUF1 (N10938, N10931);
or OR4 (N10939, N10900, N9324, N7061, N9144);
or OR4 (N10940, N10937, N2250, N9729, N8202);
and AND4 (N10941, N10923, N6405, N7346, N3076);
xor XOR2 (N10942, N10939, N1283);
xor XOR2 (N10943, N10935, N1093);
not NOT1 (N10944, N10933);
buf BUF1 (N10945, N10920);
not NOT1 (N10946, N10938);
nand NAND2 (N10947, N10941, N6508);
xor XOR2 (N10948, N10947, N6021);
buf BUF1 (N10949, N10928);
nor NOR4 (N10950, N10949, N7931, N885, N6580);
or OR4 (N10951, N10945, N5039, N2582, N10740);
and AND4 (N10952, N10919, N2231, N668, N1726);
and AND3 (N10953, N10951, N8005, N9293);
nand NAND4 (N10954, N10952, N9062, N3938, N2109);
buf BUF1 (N10955, N10950);
or OR2 (N10956, N10943, N3405);
nor NOR3 (N10957, N10954, N7100, N10174);
buf BUF1 (N10958, N10956);
or OR2 (N10959, N10957, N8618);
xor XOR2 (N10960, N10948, N4943);
and AND2 (N10961, N10946, N3150);
nor NOR2 (N10962, N10942, N1520);
nor NOR3 (N10963, N10944, N7818, N10576);
xor XOR2 (N10964, N10962, N9084);
xor XOR2 (N10965, N10953, N10129);
or OR4 (N10966, N10934, N6420, N7399, N436);
or OR2 (N10967, N10963, N9317);
nand NAND3 (N10968, N10967, N1084, N1896);
or OR4 (N10969, N10958, N8444, N4253, N6745);
xor XOR2 (N10970, N10968, N4647);
buf BUF1 (N10971, N10966);
not NOT1 (N10972, N10969);
buf BUF1 (N10973, N10940);
nand NAND2 (N10974, N10961, N4589);
xor XOR2 (N10975, N10955, N7950);
xor XOR2 (N10976, N10965, N1834);
nor NOR2 (N10977, N10970, N4803);
and AND2 (N10978, N10973, N8084);
not NOT1 (N10979, N10964);
and AND4 (N10980, N10971, N3644, N5517, N5900);
not NOT1 (N10981, N10979);
xor XOR2 (N10982, N10976, N256);
nand NAND2 (N10983, N10981, N9345);
and AND4 (N10984, N10959, N7317, N5215, N1140);
xor XOR2 (N10985, N10974, N6261);
xor XOR2 (N10986, N10975, N7073);
buf BUF1 (N10987, N10986);
not NOT1 (N10988, N10960);
not NOT1 (N10989, N10987);
not NOT1 (N10990, N10983);
buf BUF1 (N10991, N10990);
buf BUF1 (N10992, N10988);
and AND4 (N10993, N10985, N8306, N10162, N2323);
not NOT1 (N10994, N10977);
buf BUF1 (N10995, N10984);
and AND3 (N10996, N10978, N8405, N4137);
nor NOR2 (N10997, N10982, N3341);
or OR4 (N10998, N10996, N2334, N4190, N2680);
buf BUF1 (N10999, N10997);
buf BUF1 (N11000, N10993);
not NOT1 (N11001, N10992);
nand NAND3 (N11002, N10995, N10269, N6306);
nor NOR4 (N11003, N10999, N2225, N9915, N1677);
and AND2 (N11004, N10998, N8493);
not NOT1 (N11005, N10972);
nor NOR2 (N11006, N10991, N9356);
buf BUF1 (N11007, N11004);
or OR3 (N11008, N11001, N2721, N10479);
nor NOR4 (N11009, N10989, N7979, N10233, N7776);
and AND2 (N11010, N10980, N6323);
or OR4 (N11011, N11009, N7102, N5536, N9799);
buf BUF1 (N11012, N11000);
nand NAND4 (N11013, N11008, N6738, N1276, N5795);
and AND4 (N11014, N11011, N6107, N3597, N8254);
xor XOR2 (N11015, N11005, N3962);
nor NOR3 (N11016, N11003, N2780, N9356);
nor NOR4 (N11017, N11012, N5129, N5567, N3313);
or OR3 (N11018, N11017, N2054, N6600);
not NOT1 (N11019, N11018);
buf BUF1 (N11020, N11019);
xor XOR2 (N11021, N11002, N5736);
buf BUF1 (N11022, N10994);
not NOT1 (N11023, N11020);
nor NOR2 (N11024, N11021, N3063);
buf BUF1 (N11025, N11010);
nand NAND2 (N11026, N11006, N1787);
and AND4 (N11027, N11023, N8014, N428, N5238);
and AND2 (N11028, N11016, N3245);
not NOT1 (N11029, N11027);
not NOT1 (N11030, N11013);
nand NAND2 (N11031, N11030, N10800);
and AND2 (N11032, N11015, N8720);
or OR2 (N11033, N11029, N8837);
not NOT1 (N11034, N11032);
and AND3 (N11035, N11007, N2310, N6101);
nor NOR2 (N11036, N11031, N513);
nand NAND2 (N11037, N11025, N637);
nor NOR3 (N11038, N11037, N8424, N4751);
or OR2 (N11039, N11024, N9787);
buf BUF1 (N11040, N11039);
not NOT1 (N11041, N11040);
xor XOR2 (N11042, N11028, N8075);
or OR4 (N11043, N11026, N3232, N15, N9677);
not NOT1 (N11044, N11043);
not NOT1 (N11045, N11033);
and AND2 (N11046, N11036, N300);
nand NAND2 (N11047, N11044, N2534);
buf BUF1 (N11048, N11038);
or OR2 (N11049, N11014, N4481);
buf BUF1 (N11050, N11022);
xor XOR2 (N11051, N11047, N9326);
not NOT1 (N11052, N11041);
or OR2 (N11053, N11046, N6365);
nand NAND3 (N11054, N11045, N3702, N3984);
nand NAND3 (N11055, N11048, N5075, N2534);
or OR3 (N11056, N11051, N97, N7646);
nand NAND3 (N11057, N11055, N4414, N1298);
or OR2 (N11058, N11056, N9880);
xor XOR2 (N11059, N11053, N9698);
nor NOR4 (N11060, N11042, N9043, N7151, N1513);
or OR2 (N11061, N11035, N1430);
xor XOR2 (N11062, N11049, N10403);
and AND2 (N11063, N11054, N8658);
and AND3 (N11064, N11059, N6120, N9372);
nand NAND3 (N11065, N11034, N5330, N4309);
buf BUF1 (N11066, N11058);
or OR2 (N11067, N11052, N3983);
xor XOR2 (N11068, N11063, N7959);
and AND3 (N11069, N11061, N543, N3675);
nand NAND4 (N11070, N11062, N3002, N9995, N10925);
buf BUF1 (N11071, N11050);
not NOT1 (N11072, N11070);
nand NAND3 (N11073, N11068, N9531, N5565);
buf BUF1 (N11074, N11065);
nand NAND3 (N11075, N11060, N8925, N8962);
or OR2 (N11076, N11057, N3763);
nor NOR4 (N11077, N11072, N1615, N5304, N6610);
nor NOR4 (N11078, N11071, N7329, N10784, N7184);
not NOT1 (N11079, N11069);
nand NAND4 (N11080, N11076, N7115, N4522, N4935);
nor NOR2 (N11081, N11078, N8704);
nand NAND3 (N11082, N11080, N2130, N5962);
xor XOR2 (N11083, N11073, N9469);
not NOT1 (N11084, N11074);
buf BUF1 (N11085, N11066);
xor XOR2 (N11086, N11082, N4869);
and AND2 (N11087, N11064, N242);
buf BUF1 (N11088, N11086);
and AND4 (N11089, N11085, N6102, N1558, N6674);
not NOT1 (N11090, N11075);
xor XOR2 (N11091, N11084, N2879);
or OR3 (N11092, N11083, N5031, N2614);
buf BUF1 (N11093, N11090);
buf BUF1 (N11094, N11092);
and AND3 (N11095, N11077, N7416, N6877);
and AND4 (N11096, N11091, N8787, N10039, N4581);
buf BUF1 (N11097, N11089);
nand NAND2 (N11098, N11094, N1114);
and AND4 (N11099, N11087, N5559, N10463, N8919);
not NOT1 (N11100, N11067);
nor NOR3 (N11101, N11081, N1724, N7337);
nor NOR2 (N11102, N11097, N10326);
or OR3 (N11103, N11096, N5276, N9352);
not NOT1 (N11104, N11079);
nand NAND2 (N11105, N11099, N938);
not NOT1 (N11106, N11100);
or OR3 (N11107, N11101, N9510, N6843);
not NOT1 (N11108, N11107);
nor NOR3 (N11109, N11088, N5084, N6712);
or OR2 (N11110, N11105, N5969);
nand NAND4 (N11111, N11106, N1854, N5727, N2854);
or OR2 (N11112, N11110, N1516);
and AND3 (N11113, N11103, N4148, N3114);
buf BUF1 (N11114, N11108);
and AND3 (N11115, N11112, N4317, N1243);
or OR4 (N11116, N11115, N8757, N9471, N10240);
nor NOR3 (N11117, N11095, N1115, N8681);
nand NAND2 (N11118, N11098, N8986);
nand NAND4 (N11119, N11109, N2228, N9987, N2855);
or OR3 (N11120, N11102, N6159, N2454);
not NOT1 (N11121, N11117);
xor XOR2 (N11122, N11118, N4392);
buf BUF1 (N11123, N11111);
nand NAND2 (N11124, N11093, N7034);
nand NAND4 (N11125, N11121, N1831, N935, N7721);
not NOT1 (N11126, N11122);
nor NOR4 (N11127, N11125, N21, N7467, N10510);
not NOT1 (N11128, N11127);
and AND3 (N11129, N11119, N11073, N9267);
and AND3 (N11130, N11104, N7703, N9107);
not NOT1 (N11131, N11114);
nand NAND2 (N11132, N11129, N7323);
nand NAND3 (N11133, N11128, N5828, N10022);
and AND4 (N11134, N11133, N1769, N10658, N7998);
buf BUF1 (N11135, N11120);
or OR3 (N11136, N11116, N2777, N2684);
xor XOR2 (N11137, N11123, N7065);
buf BUF1 (N11138, N11135);
not NOT1 (N11139, N11132);
nor NOR3 (N11140, N11136, N4252, N10964);
buf BUF1 (N11141, N11139);
nor NOR2 (N11142, N11140, N8632);
and AND2 (N11143, N11124, N10149);
nand NAND4 (N11144, N11141, N3727, N1569, N5254);
xor XOR2 (N11145, N11143, N3113);
not NOT1 (N11146, N11138);
nor NOR3 (N11147, N11131, N4618, N10417);
buf BUF1 (N11148, N11146);
and AND2 (N11149, N11144, N2412);
not NOT1 (N11150, N11145);
xor XOR2 (N11151, N11147, N3320);
not NOT1 (N11152, N11151);
xor XOR2 (N11153, N11150, N7705);
not NOT1 (N11154, N11148);
or OR3 (N11155, N11154, N9788, N1435);
nor NOR3 (N11156, N11155, N9785, N1380);
buf BUF1 (N11157, N11134);
buf BUF1 (N11158, N11149);
and AND2 (N11159, N11137, N3477);
nor NOR3 (N11160, N11158, N6164, N5006);
buf BUF1 (N11161, N11126);
or OR2 (N11162, N11156, N1021);
nand NAND2 (N11163, N11130, N5031);
not NOT1 (N11164, N11152);
nor NOR3 (N11165, N11142, N4887, N701);
nor NOR4 (N11166, N11162, N10589, N2419, N2096);
xor XOR2 (N11167, N11113, N2270);
buf BUF1 (N11168, N11153);
xor XOR2 (N11169, N11157, N3192);
not NOT1 (N11170, N11161);
buf BUF1 (N11171, N11164);
nor NOR3 (N11172, N11160, N8182, N1904);
nand NAND3 (N11173, N11169, N7672, N997);
and AND4 (N11174, N11168, N1277, N1530, N4783);
nand NAND2 (N11175, N11163, N10625);
nand NAND2 (N11176, N11159, N8761);
buf BUF1 (N11177, N11166);
xor XOR2 (N11178, N11173, N10766);
or OR3 (N11179, N11165, N3870, N9266);
not NOT1 (N11180, N11174);
xor XOR2 (N11181, N11178, N10274);
not NOT1 (N11182, N11179);
nand NAND4 (N11183, N11171, N3024, N1680, N5334);
nand NAND2 (N11184, N11176, N9828);
nor NOR3 (N11185, N11180, N10796, N2393);
not NOT1 (N11186, N11184);
and AND4 (N11187, N11172, N4224, N2228, N2186);
and AND3 (N11188, N11170, N9742, N10490);
and AND4 (N11189, N11175, N11014, N9910, N10586);
not NOT1 (N11190, N11189);
nor NOR3 (N11191, N11186, N10757, N8336);
nor NOR3 (N11192, N11177, N10246, N10023);
nand NAND3 (N11193, N11191, N4879, N3883);
and AND4 (N11194, N11185, N3292, N4414, N6587);
xor XOR2 (N11195, N11183, N2947);
nor NOR2 (N11196, N11190, N7686);
and AND4 (N11197, N11167, N3568, N8143, N1056);
nor NOR4 (N11198, N11196, N8150, N10573, N5771);
nand NAND2 (N11199, N11192, N2365);
not NOT1 (N11200, N11187);
nor NOR2 (N11201, N11200, N10432);
and AND2 (N11202, N11194, N764);
nand NAND2 (N11203, N11195, N8361);
buf BUF1 (N11204, N11181);
and AND4 (N11205, N11193, N9467, N8341, N356);
not NOT1 (N11206, N11204);
xor XOR2 (N11207, N11202, N8315);
nand NAND4 (N11208, N11201, N8239, N7045, N7294);
nand NAND2 (N11209, N11203, N5614);
or OR4 (N11210, N11199, N3550, N2055, N10808);
not NOT1 (N11211, N11208);
not NOT1 (N11212, N11188);
nor NOR3 (N11213, N11209, N581, N1366);
nand NAND2 (N11214, N11198, N5911);
not NOT1 (N11215, N11197);
nor NOR4 (N11216, N11207, N4134, N6311, N7700);
buf BUF1 (N11217, N11214);
not NOT1 (N11218, N11210);
and AND2 (N11219, N11182, N3495);
or OR3 (N11220, N11215, N2067, N2102);
or OR4 (N11221, N11212, N2873, N1013, N4726);
and AND4 (N11222, N11206, N8140, N363, N249);
nand NAND4 (N11223, N11205, N5246, N5623, N5243);
and AND4 (N11224, N11216, N9250, N9331, N9219);
nor NOR2 (N11225, N11220, N10274);
not NOT1 (N11226, N11224);
or OR2 (N11227, N11222, N3302);
and AND3 (N11228, N11218, N5755, N7320);
xor XOR2 (N11229, N11213, N10318);
nor NOR3 (N11230, N11226, N5364, N3786);
buf BUF1 (N11231, N11217);
xor XOR2 (N11232, N11211, N675);
buf BUF1 (N11233, N11219);
xor XOR2 (N11234, N11230, N8000);
buf BUF1 (N11235, N11229);
and AND4 (N11236, N11235, N10113, N7155, N5154);
buf BUF1 (N11237, N11232);
buf BUF1 (N11238, N11228);
and AND4 (N11239, N11231, N5713, N3925, N5879);
xor XOR2 (N11240, N11238, N7968);
xor XOR2 (N11241, N11221, N5835);
nand NAND2 (N11242, N11223, N9693);
xor XOR2 (N11243, N11236, N490);
not NOT1 (N11244, N11239);
nand NAND4 (N11245, N11241, N2549, N7082, N3902);
and AND4 (N11246, N11225, N2245, N9663, N11117);
and AND2 (N11247, N11227, N8836);
xor XOR2 (N11248, N11233, N10442);
buf BUF1 (N11249, N11240);
or OR3 (N11250, N11237, N8579, N6034);
not NOT1 (N11251, N11248);
not NOT1 (N11252, N11234);
xor XOR2 (N11253, N11252, N5411);
nand NAND2 (N11254, N11246, N9065);
buf BUF1 (N11255, N11251);
buf BUF1 (N11256, N11255);
and AND3 (N11257, N11247, N236, N3502);
xor XOR2 (N11258, N11250, N6667);
nand NAND2 (N11259, N11245, N2412);
buf BUF1 (N11260, N11253);
nor NOR4 (N11261, N11244, N8095, N4640, N6861);
buf BUF1 (N11262, N11249);
not NOT1 (N11263, N11256);
and AND4 (N11264, N11254, N8617, N8857, N5871);
nand NAND4 (N11265, N11260, N8130, N3602, N10429);
or OR4 (N11266, N11261, N802, N831, N239);
xor XOR2 (N11267, N11257, N7223);
not NOT1 (N11268, N11243);
nor NOR2 (N11269, N11263, N4504);
or OR4 (N11270, N11266, N7645, N9416, N3270);
or OR2 (N11271, N11258, N7659);
buf BUF1 (N11272, N11270);
buf BUF1 (N11273, N11242);
not NOT1 (N11274, N11262);
xor XOR2 (N11275, N11271, N9501);
and AND2 (N11276, N11269, N86);
and AND2 (N11277, N11276, N900);
or OR2 (N11278, N11272, N8824);
not NOT1 (N11279, N11277);
xor XOR2 (N11280, N11278, N1701);
buf BUF1 (N11281, N11265);
and AND2 (N11282, N11281, N1330);
and AND2 (N11283, N11280, N9194);
not NOT1 (N11284, N11273);
not NOT1 (N11285, N11283);
and AND2 (N11286, N11268, N10708);
xor XOR2 (N11287, N11279, N7577);
buf BUF1 (N11288, N11284);
not NOT1 (N11289, N11286);
nand NAND3 (N11290, N11285, N1856, N3423);
or OR2 (N11291, N11274, N9845);
not NOT1 (N11292, N11264);
not NOT1 (N11293, N11259);
nand NAND4 (N11294, N11288, N1343, N448, N3760);
nand NAND3 (N11295, N11291, N2068, N3174);
buf BUF1 (N11296, N11292);
xor XOR2 (N11297, N11275, N2280);
nor NOR2 (N11298, N11282, N875);
nand NAND3 (N11299, N11294, N5558, N8011);
nand NAND4 (N11300, N11297, N2931, N10132, N9905);
nor NOR4 (N11301, N11296, N245, N9886, N7283);
buf BUF1 (N11302, N11298);
xor XOR2 (N11303, N11287, N10948);
xor XOR2 (N11304, N11289, N4302);
nand NAND3 (N11305, N11267, N10668, N6781);
nand NAND2 (N11306, N11300, N9606);
buf BUF1 (N11307, N11303);
nor NOR2 (N11308, N11293, N6421);
and AND4 (N11309, N11299, N9111, N10604, N4099);
not NOT1 (N11310, N11309);
nand NAND3 (N11311, N11295, N7627, N10811);
xor XOR2 (N11312, N11302, N2614);
or OR2 (N11313, N11308, N8435);
and AND3 (N11314, N11290, N4015, N5194);
not NOT1 (N11315, N11305);
buf BUF1 (N11316, N11304);
not NOT1 (N11317, N11311);
nor NOR2 (N11318, N11312, N9606);
xor XOR2 (N11319, N11316, N489);
not NOT1 (N11320, N11317);
xor XOR2 (N11321, N11314, N7000);
nand NAND3 (N11322, N11307, N3409, N11279);
xor XOR2 (N11323, N11301, N11278);
not NOT1 (N11324, N11313);
and AND2 (N11325, N11324, N9518);
buf BUF1 (N11326, N11323);
buf BUF1 (N11327, N11319);
buf BUF1 (N11328, N11321);
or OR4 (N11329, N11325, N9459, N2811, N2068);
and AND3 (N11330, N11327, N4559, N2634);
xor XOR2 (N11331, N11328, N5351);
nor NOR2 (N11332, N11310, N1407);
nor NOR4 (N11333, N11322, N4388, N1203, N8557);
nand NAND4 (N11334, N11326, N2149, N1454, N75);
and AND3 (N11335, N11333, N7767, N2194);
and AND3 (N11336, N11315, N5164, N567);
nor NOR3 (N11337, N11332, N4110, N4934);
or OR2 (N11338, N11306, N11225);
not NOT1 (N11339, N11330);
not NOT1 (N11340, N11336);
xor XOR2 (N11341, N11320, N9735);
not NOT1 (N11342, N11341);
not NOT1 (N11343, N11331);
or OR3 (N11344, N11334, N6946, N676);
and AND2 (N11345, N11343, N6863);
buf BUF1 (N11346, N11335);
not NOT1 (N11347, N11338);
and AND2 (N11348, N11347, N782);
nand NAND2 (N11349, N11318, N6577);
buf BUF1 (N11350, N11340);
or OR4 (N11351, N11346, N4402, N5863, N8333);
not NOT1 (N11352, N11351);
not NOT1 (N11353, N11329);
or OR4 (N11354, N11353, N6644, N9064, N6272);
and AND3 (N11355, N11348, N10505, N7252);
xor XOR2 (N11356, N11354, N3976);
xor XOR2 (N11357, N11344, N4013);
buf BUF1 (N11358, N11350);
xor XOR2 (N11359, N11355, N465);
nand NAND3 (N11360, N11349, N10200, N11084);
nor NOR2 (N11361, N11342, N10216);
or OR4 (N11362, N11361, N8227, N11204, N8603);
not NOT1 (N11363, N11352);
nand NAND4 (N11364, N11358, N7165, N1627, N2002);
or OR3 (N11365, N11364, N11335, N5699);
not NOT1 (N11366, N11345);
buf BUF1 (N11367, N11359);
nor NOR2 (N11368, N11360, N8992);
and AND4 (N11369, N11368, N4379, N3073, N3768);
or OR4 (N11370, N11369, N4397, N6785, N1995);
buf BUF1 (N11371, N11357);
nor NOR3 (N11372, N11370, N2891, N2417);
buf BUF1 (N11373, N11339);
not NOT1 (N11374, N11337);
buf BUF1 (N11375, N11373);
xor XOR2 (N11376, N11371, N6701);
and AND4 (N11377, N11365, N4549, N8204, N10963);
xor XOR2 (N11378, N11362, N2076);
nand NAND4 (N11379, N11367, N6275, N5173, N11306);
nand NAND2 (N11380, N11378, N1707);
nor NOR2 (N11381, N11380, N2367);
xor XOR2 (N11382, N11379, N5595);
not NOT1 (N11383, N11377);
or OR3 (N11384, N11372, N8531, N479);
or OR2 (N11385, N11382, N32);
nor NOR2 (N11386, N11375, N9420);
nand NAND4 (N11387, N11384, N3623, N459, N8607);
not NOT1 (N11388, N11374);
xor XOR2 (N11389, N11386, N11366);
buf BUF1 (N11390, N7617);
buf BUF1 (N11391, N11376);
nor NOR2 (N11392, N11390, N2001);
nor NOR3 (N11393, N11387, N2674, N5064);
nor NOR2 (N11394, N11356, N7013);
buf BUF1 (N11395, N11388);
nand NAND2 (N11396, N11392, N10579);
nand NAND2 (N11397, N11393, N828);
and AND2 (N11398, N11385, N8069);
xor XOR2 (N11399, N11363, N8748);
not NOT1 (N11400, N11394);
xor XOR2 (N11401, N11381, N4677);
buf BUF1 (N11402, N11397);
and AND2 (N11403, N11396, N2691);
not NOT1 (N11404, N11399);
nand NAND4 (N11405, N11400, N3914, N6989, N7777);
or OR2 (N11406, N11389, N6622);
xor XOR2 (N11407, N11405, N5570);
nand NAND4 (N11408, N11383, N3479, N5187, N8621);
and AND2 (N11409, N11398, N1749);
buf BUF1 (N11410, N11403);
buf BUF1 (N11411, N11391);
buf BUF1 (N11412, N11411);
and AND2 (N11413, N11410, N2378);
nor NOR2 (N11414, N11409, N4282);
or OR2 (N11415, N11402, N167);
and AND3 (N11416, N11413, N7638, N466);
xor XOR2 (N11417, N11412, N1898);
nand NAND4 (N11418, N11415, N377, N9586, N1170);
nand NAND2 (N11419, N11418, N760);
or OR4 (N11420, N11419, N9222, N8981, N4876);
buf BUF1 (N11421, N11401);
nor NOR4 (N11422, N11408, N3280, N10117, N7351);
buf BUF1 (N11423, N11422);
xor XOR2 (N11424, N11423, N8813);
not NOT1 (N11425, N11421);
xor XOR2 (N11426, N11414, N8073);
nand NAND3 (N11427, N11404, N7532, N9212);
xor XOR2 (N11428, N11407, N4553);
not NOT1 (N11429, N11426);
and AND4 (N11430, N11420, N1415, N2251, N5395);
or OR3 (N11431, N11424, N9292, N6610);
or OR3 (N11432, N11427, N8282, N4394);
nor NOR2 (N11433, N11406, N7724);
or OR2 (N11434, N11416, N9347);
nor NOR2 (N11435, N11434, N1241);
nor NOR3 (N11436, N11429, N10914, N601);
xor XOR2 (N11437, N11430, N8024);
or OR2 (N11438, N11395, N158);
and AND3 (N11439, N11435, N6419, N2716);
not NOT1 (N11440, N11432);
nand NAND2 (N11441, N11436, N1970);
or OR2 (N11442, N11441, N2903);
nor NOR4 (N11443, N11439, N3177, N5778, N2458);
nor NOR4 (N11444, N11437, N1075, N7331, N6510);
and AND2 (N11445, N11431, N2586);
xor XOR2 (N11446, N11433, N1596);
and AND2 (N11447, N11425, N10369);
nand NAND3 (N11448, N11438, N8493, N7054);
buf BUF1 (N11449, N11445);
nor NOR3 (N11450, N11417, N2324, N5222);
or OR2 (N11451, N11448, N6474);
xor XOR2 (N11452, N11449, N3642);
nand NAND3 (N11453, N11450, N1059, N11083);
or OR4 (N11454, N11443, N192, N6995, N4535);
nor NOR3 (N11455, N11452, N5566, N8335);
nand NAND4 (N11456, N11440, N7438, N10399, N10686);
nor NOR4 (N11457, N11444, N1724, N8280, N10734);
buf BUF1 (N11458, N11456);
buf BUF1 (N11459, N11428);
buf BUF1 (N11460, N11459);
buf BUF1 (N11461, N11447);
and AND2 (N11462, N11460, N6365);
xor XOR2 (N11463, N11455, N11285);
buf BUF1 (N11464, N11463);
nor NOR4 (N11465, N11457, N10584, N10905, N5435);
nor NOR2 (N11466, N11462, N2552);
not NOT1 (N11467, N11466);
nor NOR4 (N11468, N11454, N3500, N1060, N610);
or OR2 (N11469, N11467, N3091);
or OR4 (N11470, N11442, N8290, N742, N3938);
not NOT1 (N11471, N11451);
xor XOR2 (N11472, N11468, N4163);
not NOT1 (N11473, N11461);
buf BUF1 (N11474, N11446);
or OR4 (N11475, N11458, N6698, N11307, N1128);
buf BUF1 (N11476, N11475);
not NOT1 (N11477, N11473);
nor NOR2 (N11478, N11465, N9473);
nor NOR2 (N11479, N11469, N2552);
or OR3 (N11480, N11453, N3134, N3455);
buf BUF1 (N11481, N11478);
and AND2 (N11482, N11474, N460);
or OR4 (N11483, N11470, N3817, N6947, N7832);
nand NAND4 (N11484, N11476, N68, N1730, N10964);
buf BUF1 (N11485, N11472);
xor XOR2 (N11486, N11477, N4630);
and AND4 (N11487, N11484, N2581, N6417, N9575);
or OR3 (N11488, N11479, N10775, N3894);
nand NAND3 (N11489, N11471, N6194, N10385);
buf BUF1 (N11490, N11487);
nand NAND2 (N11491, N11490, N4529);
nand NAND3 (N11492, N11481, N10484, N11182);
buf BUF1 (N11493, N11485);
or OR2 (N11494, N11493, N10537);
not NOT1 (N11495, N11486);
nand NAND4 (N11496, N11464, N884, N2457, N10686);
or OR4 (N11497, N11482, N8316, N5345, N3382);
xor XOR2 (N11498, N11497, N10187);
buf BUF1 (N11499, N11483);
not NOT1 (N11500, N11491);
buf BUF1 (N11501, N11500);
nor NOR3 (N11502, N11495, N3411, N4134);
and AND3 (N11503, N11494, N8825, N3203);
not NOT1 (N11504, N11502);
not NOT1 (N11505, N11492);
and AND2 (N11506, N11498, N1173);
or OR3 (N11507, N11480, N9680, N6129);
and AND4 (N11508, N11499, N8789, N277, N5763);
buf BUF1 (N11509, N11503);
nand NAND3 (N11510, N11505, N11112, N10679);
xor XOR2 (N11511, N11509, N5587);
nor NOR4 (N11512, N11507, N10731, N3568, N3462);
not NOT1 (N11513, N11510);
buf BUF1 (N11514, N11513);
or OR4 (N11515, N11514, N10203, N7078, N156);
nand NAND2 (N11516, N11496, N9208);
and AND2 (N11517, N11516, N7264);
xor XOR2 (N11518, N11515, N247);
and AND2 (N11519, N11508, N4208);
and AND3 (N11520, N11519, N5284, N2355);
xor XOR2 (N11521, N11511, N10258);
nor NOR4 (N11522, N11489, N1987, N6842, N10432);
not NOT1 (N11523, N11521);
nor NOR4 (N11524, N11517, N423, N2891, N7224);
nor NOR4 (N11525, N11524, N687, N3086, N241);
and AND3 (N11526, N11525, N2378, N4135);
not NOT1 (N11527, N11501);
and AND2 (N11528, N11527, N7274);
xor XOR2 (N11529, N11526, N138);
nor NOR2 (N11530, N11528, N10460);
nand NAND2 (N11531, N11530, N7907);
xor XOR2 (N11532, N11522, N6149);
nor NOR3 (N11533, N11504, N8708, N3388);
buf BUF1 (N11534, N11488);
nand NAND2 (N11535, N11523, N11418);
buf BUF1 (N11536, N11520);
not NOT1 (N11537, N11518);
buf BUF1 (N11538, N11536);
not NOT1 (N11539, N11512);
buf BUF1 (N11540, N11534);
buf BUF1 (N11541, N11533);
xor XOR2 (N11542, N11506, N6154);
and AND3 (N11543, N11538, N6788, N10405);
not NOT1 (N11544, N11539);
not NOT1 (N11545, N11540);
xor XOR2 (N11546, N11543, N6868);
buf BUF1 (N11547, N11535);
or OR2 (N11548, N11547, N1672);
nand NAND2 (N11549, N11542, N9399);
and AND4 (N11550, N11537, N10217, N657, N362);
or OR2 (N11551, N11541, N9378);
or OR4 (N11552, N11550, N1026, N5533, N9011);
xor XOR2 (N11553, N11548, N1971);
buf BUF1 (N11554, N11553);
nand NAND4 (N11555, N11552, N9763, N8341, N6298);
nand NAND4 (N11556, N11546, N729, N2529, N3474);
and AND4 (N11557, N11544, N2034, N4446, N1000);
buf BUF1 (N11558, N11557);
not NOT1 (N11559, N11531);
or OR3 (N11560, N11545, N640, N823);
or OR3 (N11561, N11555, N1456, N1148);
and AND2 (N11562, N11556, N1155);
buf BUF1 (N11563, N11558);
buf BUF1 (N11564, N11551);
nor NOR2 (N11565, N11564, N10415);
xor XOR2 (N11566, N11561, N898);
buf BUF1 (N11567, N11563);
not NOT1 (N11568, N11566);
or OR2 (N11569, N11568, N10380);
nor NOR3 (N11570, N11554, N1078, N36);
nand NAND2 (N11571, N11529, N9766);
and AND3 (N11572, N11571, N6618, N255);
and AND3 (N11573, N11572, N8244, N2579);
buf BUF1 (N11574, N11562);
or OR3 (N11575, N11549, N4425, N4331);
not NOT1 (N11576, N11532);
and AND3 (N11577, N11567, N6967, N4651);
and AND2 (N11578, N11565, N10540);
xor XOR2 (N11579, N11578, N10433);
nor NOR4 (N11580, N11570, N3985, N7054, N6045);
or OR2 (N11581, N11573, N4637);
buf BUF1 (N11582, N11569);
and AND4 (N11583, N11559, N7385, N2957, N3022);
or OR2 (N11584, N11574, N10546);
xor XOR2 (N11585, N11584, N9214);
not NOT1 (N11586, N11582);
or OR4 (N11587, N11586, N6691, N7483, N5034);
and AND3 (N11588, N11575, N10933, N10346);
xor XOR2 (N11589, N11560, N8618);
nor NOR2 (N11590, N11580, N673);
not NOT1 (N11591, N11587);
xor XOR2 (N11592, N11576, N6026);
xor XOR2 (N11593, N11589, N8831);
not NOT1 (N11594, N11581);
xor XOR2 (N11595, N11590, N9157);
nor NOR4 (N11596, N11577, N10067, N7279, N3997);
and AND2 (N11597, N11591, N5726);
nor NOR4 (N11598, N11596, N5742, N2349, N578);
nand NAND3 (N11599, N11583, N5585, N6448);
nor NOR4 (N11600, N11599, N532, N4604, N3918);
or OR3 (N11601, N11597, N11145, N10580);
xor XOR2 (N11602, N11601, N7365);
xor XOR2 (N11603, N11592, N10088);
nor NOR4 (N11604, N11585, N5921, N9100, N10485);
or OR2 (N11605, N11594, N1326);
or OR4 (N11606, N11605, N4661, N1298, N10561);
or OR4 (N11607, N11598, N3354, N2697, N3333);
buf BUF1 (N11608, N11602);
xor XOR2 (N11609, N11607, N10463);
nand NAND4 (N11610, N11608, N324, N2166, N739);
buf BUF1 (N11611, N11595);
and AND4 (N11612, N11600, N5084, N4769, N1432);
buf BUF1 (N11613, N11604);
xor XOR2 (N11614, N11579, N5914);
nand NAND4 (N11615, N11612, N3180, N6463, N6082);
and AND4 (N11616, N11614, N6296, N6349, N8424);
or OR2 (N11617, N11609, N9064);
nand NAND3 (N11618, N11606, N9143, N5479);
not NOT1 (N11619, N11610);
not NOT1 (N11620, N11619);
nor NOR4 (N11621, N11620, N9557, N4531, N9345);
not NOT1 (N11622, N11611);
not NOT1 (N11623, N11603);
not NOT1 (N11624, N11613);
nor NOR3 (N11625, N11623, N789, N4029);
buf BUF1 (N11626, N11617);
nand NAND4 (N11627, N11626, N8854, N1388, N6061);
xor XOR2 (N11628, N11588, N1670);
nor NOR4 (N11629, N11625, N7578, N10471, N9872);
buf BUF1 (N11630, N11593);
or OR2 (N11631, N11628, N8244);
and AND2 (N11632, N11621, N2495);
buf BUF1 (N11633, N11622);
and AND3 (N11634, N11627, N9588, N6158);
not NOT1 (N11635, N11632);
nor NOR3 (N11636, N11631, N7221, N10529);
and AND3 (N11637, N11633, N11424, N5703);
not NOT1 (N11638, N11618);
xor XOR2 (N11639, N11616, N4677);
nor NOR2 (N11640, N11629, N8865);
not NOT1 (N11641, N11630);
not NOT1 (N11642, N11636);
and AND2 (N11643, N11641, N5070);
xor XOR2 (N11644, N11624, N11573);
xor XOR2 (N11645, N11615, N8774);
buf BUF1 (N11646, N11644);
buf BUF1 (N11647, N11635);
xor XOR2 (N11648, N11643, N11204);
or OR4 (N11649, N11648, N1280, N1843, N1481);
nor NOR4 (N11650, N11639, N2239, N10767, N2550);
xor XOR2 (N11651, N11634, N8426);
xor XOR2 (N11652, N11650, N8527);
buf BUF1 (N11653, N11649);
xor XOR2 (N11654, N11638, N6238);
nand NAND2 (N11655, N11652, N11406);
buf BUF1 (N11656, N11651);
or OR2 (N11657, N11646, N11091);
not NOT1 (N11658, N11657);
and AND4 (N11659, N11656, N2278, N9198, N2379);
and AND3 (N11660, N11655, N2500, N722);
xor XOR2 (N11661, N11645, N5370);
and AND2 (N11662, N11647, N3585);
nand NAND4 (N11663, N11654, N9543, N8107, N5663);
xor XOR2 (N11664, N11662, N4331);
buf BUF1 (N11665, N11653);
xor XOR2 (N11666, N11664, N10548);
and AND3 (N11667, N11661, N2781, N3444);
buf BUF1 (N11668, N11637);
buf BUF1 (N11669, N11666);
and AND3 (N11670, N11668, N5784, N2684);
buf BUF1 (N11671, N11640);
buf BUF1 (N11672, N11659);
nand NAND4 (N11673, N11642, N6535, N9379, N8606);
buf BUF1 (N11674, N11672);
or OR2 (N11675, N11663, N7394);
not NOT1 (N11676, N11673);
nor NOR4 (N11677, N11658, N6479, N6476, N4294);
and AND4 (N11678, N11674, N9006, N713, N10670);
nand NAND3 (N11679, N11667, N9859, N4048);
or OR2 (N11680, N11660, N5229);
xor XOR2 (N11681, N11670, N7048);
buf BUF1 (N11682, N11669);
nor NOR3 (N11683, N11676, N8742, N488);
nor NOR2 (N11684, N11678, N26);
buf BUF1 (N11685, N11679);
nand NAND4 (N11686, N11683, N6967, N1118, N2721);
not NOT1 (N11687, N11665);
nor NOR3 (N11688, N11687, N6576, N5564);
nor NOR3 (N11689, N11680, N9675, N2935);
nand NAND4 (N11690, N11685, N7200, N10194, N7405);
nand NAND2 (N11691, N11690, N4912);
nand NAND3 (N11692, N11691, N6014, N3909);
and AND3 (N11693, N11677, N10887, N3744);
nor NOR2 (N11694, N11682, N4811);
nand NAND4 (N11695, N11686, N1846, N465, N9219);
nor NOR2 (N11696, N11671, N4854);
not NOT1 (N11697, N11681);
xor XOR2 (N11698, N11675, N2701);
or OR4 (N11699, N11697, N6987, N4927, N660);
and AND4 (N11700, N11696, N5862, N3040, N11337);
and AND2 (N11701, N11694, N7104);
nor NOR2 (N11702, N11698, N8795);
or OR2 (N11703, N11693, N9452);
xor XOR2 (N11704, N11699, N3400);
nand NAND3 (N11705, N11695, N2490, N1887);
nor NOR3 (N11706, N11701, N9386, N3936);
xor XOR2 (N11707, N11702, N9605);
nor NOR2 (N11708, N11684, N6990);
not NOT1 (N11709, N11703);
and AND4 (N11710, N11700, N7226, N6700, N3679);
buf BUF1 (N11711, N11710);
not NOT1 (N11712, N11689);
xor XOR2 (N11713, N11712, N980);
xor XOR2 (N11714, N11704, N9699);
not NOT1 (N11715, N11706);
xor XOR2 (N11716, N11713, N939);
nor NOR3 (N11717, N11707, N440, N7333);
buf BUF1 (N11718, N11705);
nor NOR4 (N11719, N11716, N1886, N7085, N10960);
nand NAND3 (N11720, N11708, N10421, N7323);
or OR3 (N11721, N11718, N2950, N11027);
nor NOR3 (N11722, N11688, N5044, N11619);
not NOT1 (N11723, N11719);
xor XOR2 (N11724, N11717, N8828);
xor XOR2 (N11725, N11722, N1884);
buf BUF1 (N11726, N11714);
nand NAND3 (N11727, N11723, N4116, N8347);
xor XOR2 (N11728, N11721, N11006);
and AND3 (N11729, N11724, N1823, N7286);
nor NOR2 (N11730, N11728, N6867);
nor NOR2 (N11731, N11715, N4481);
and AND4 (N11732, N11720, N1796, N5828, N9724);
nand NAND4 (N11733, N11692, N2587, N8301, N1276);
and AND4 (N11734, N11732, N3402, N9908, N7507);
xor XOR2 (N11735, N11733, N7875);
nand NAND3 (N11736, N11727, N11413, N8233);
buf BUF1 (N11737, N11709);
not NOT1 (N11738, N11734);
not NOT1 (N11739, N11726);
nor NOR3 (N11740, N11737, N10605, N1146);
buf BUF1 (N11741, N11711);
nor NOR3 (N11742, N11731, N10176, N5649);
or OR2 (N11743, N11740, N11282);
xor XOR2 (N11744, N11729, N11041);
and AND4 (N11745, N11741, N10365, N10466, N3160);
and AND3 (N11746, N11743, N3715, N8535);
or OR4 (N11747, N11736, N6042, N5032, N9514);
xor XOR2 (N11748, N11739, N5302);
nor NOR4 (N11749, N11744, N9330, N2698, N10783);
buf BUF1 (N11750, N11747);
xor XOR2 (N11751, N11735, N11464);
nor NOR2 (N11752, N11748, N969);
and AND2 (N11753, N11730, N6114);
buf BUF1 (N11754, N11725);
and AND4 (N11755, N11742, N3048, N3549, N7378);
nor NOR3 (N11756, N11750, N4618, N3832);
xor XOR2 (N11757, N11754, N8319);
nor NOR4 (N11758, N11746, N5448, N9926, N6032);
and AND4 (N11759, N11751, N1480, N2970, N2555);
buf BUF1 (N11760, N11749);
and AND2 (N11761, N11758, N4802);
nand NAND4 (N11762, N11755, N1546, N4983, N11695);
not NOT1 (N11763, N11753);
or OR3 (N11764, N11762, N7427, N2011);
or OR4 (N11765, N11756, N928, N7350, N6468);
nor NOR2 (N11766, N11760, N11165);
or OR3 (N11767, N11757, N1404, N1071);
nand NAND4 (N11768, N11761, N7110, N11541, N4851);
and AND2 (N11769, N11759, N7879);
nor NOR2 (N11770, N11745, N1287);
or OR4 (N11771, N11763, N4590, N8344, N837);
not NOT1 (N11772, N11765);
buf BUF1 (N11773, N11771);
xor XOR2 (N11774, N11770, N5824);
xor XOR2 (N11775, N11764, N5112);
not NOT1 (N11776, N11769);
xor XOR2 (N11777, N11776, N1196);
xor XOR2 (N11778, N11766, N9592);
and AND4 (N11779, N11778, N8810, N2905, N8424);
nor NOR2 (N11780, N11768, N8190);
nand NAND4 (N11781, N11774, N4380, N1763, N6357);
nand NAND4 (N11782, N11781, N6959, N6301, N9353);
nor NOR4 (N11783, N11779, N2914, N1489, N10221);
xor XOR2 (N11784, N11772, N620);
and AND2 (N11785, N11767, N4876);
and AND4 (N11786, N11780, N9524, N7456, N6957);
and AND2 (N11787, N11786, N10458);
nand NAND3 (N11788, N11787, N1115, N11321);
buf BUF1 (N11789, N11788);
nand NAND4 (N11790, N11785, N5857, N7852, N5511);
xor XOR2 (N11791, N11790, N8872);
or OR4 (N11792, N11777, N10289, N10281, N4328);
and AND2 (N11793, N11738, N2336);
xor XOR2 (N11794, N11752, N7843);
and AND4 (N11795, N11791, N7610, N4400, N6665);
nand NAND4 (N11796, N11783, N1187, N8581, N3841);
not NOT1 (N11797, N11789);
or OR3 (N11798, N11782, N6604, N9124);
nor NOR3 (N11799, N11773, N1050, N7236);
buf BUF1 (N11800, N11799);
nand NAND2 (N11801, N11792, N1099);
xor XOR2 (N11802, N11798, N6923);
xor XOR2 (N11803, N11795, N6441);
xor XOR2 (N11804, N11801, N9628);
buf BUF1 (N11805, N11802);
or OR3 (N11806, N11796, N9796, N2057);
xor XOR2 (N11807, N11794, N2981);
or OR3 (N11808, N11803, N3915, N4295);
not NOT1 (N11809, N11800);
nand NAND3 (N11810, N11804, N8663, N8984);
or OR4 (N11811, N11793, N11554, N7531, N104);
nor NOR2 (N11812, N11808, N4112);
or OR3 (N11813, N11806, N4125, N3915);
and AND2 (N11814, N11810, N10040);
buf BUF1 (N11815, N11811);
nor NOR3 (N11816, N11805, N11157, N10081);
buf BUF1 (N11817, N11797);
or OR3 (N11818, N11812, N9856, N9866);
nor NOR3 (N11819, N11818, N10732, N6469);
and AND2 (N11820, N11817, N4697);
and AND2 (N11821, N11775, N496);
nand NAND3 (N11822, N11814, N7648, N814);
nor NOR4 (N11823, N11809, N11558, N8071, N9092);
xor XOR2 (N11824, N11822, N2915);
nor NOR3 (N11825, N11807, N6615, N831);
or OR4 (N11826, N11819, N7111, N7506, N11067);
or OR3 (N11827, N11823, N8227, N7463);
buf BUF1 (N11828, N11827);
not NOT1 (N11829, N11828);
not NOT1 (N11830, N11820);
buf BUF1 (N11831, N11825);
xor XOR2 (N11832, N11829, N5885);
nand NAND2 (N11833, N11832, N11793);
nor NOR3 (N11834, N11833, N3284, N6575);
not NOT1 (N11835, N11830);
and AND3 (N11836, N11835, N8882, N10446);
xor XOR2 (N11837, N11826, N7491);
buf BUF1 (N11838, N11813);
xor XOR2 (N11839, N11838, N3271);
and AND2 (N11840, N11836, N7134);
or OR3 (N11841, N11816, N6885, N1933);
nor NOR3 (N11842, N11821, N3442, N3078);
and AND4 (N11843, N11824, N9793, N11300, N2816);
nand NAND3 (N11844, N11840, N7462, N8169);
nor NOR3 (N11845, N11842, N8888, N4284);
xor XOR2 (N11846, N11815, N8663);
nor NOR4 (N11847, N11841, N4268, N7340, N11171);
and AND4 (N11848, N11843, N8786, N5508, N11527);
not NOT1 (N11849, N11844);
or OR2 (N11850, N11839, N5961);
and AND2 (N11851, N11831, N8340);
nor NOR4 (N11852, N11848, N10611, N8442, N4122);
nand NAND4 (N11853, N11847, N10365, N10404, N7065);
xor XOR2 (N11854, N11834, N8401);
and AND2 (N11855, N11846, N7933);
and AND4 (N11856, N11837, N4000, N7647, N11033);
not NOT1 (N11857, N11851);
nand NAND3 (N11858, N11853, N2006, N4949);
nor NOR2 (N11859, N11850, N72);
or OR2 (N11860, N11856, N1224);
and AND4 (N11861, N11854, N11207, N11413, N10416);
or OR3 (N11862, N11849, N858, N7148);
xor XOR2 (N11863, N11845, N6765);
and AND2 (N11864, N11858, N8805);
buf BUF1 (N11865, N11852);
not NOT1 (N11866, N11862);
and AND2 (N11867, N11860, N4791);
xor XOR2 (N11868, N11859, N3450);
and AND4 (N11869, N11857, N11003, N7937, N632);
xor XOR2 (N11870, N11869, N10370);
xor XOR2 (N11871, N11870, N5619);
nor NOR3 (N11872, N11855, N486, N5430);
buf BUF1 (N11873, N11866);
nand NAND2 (N11874, N11873, N4187);
and AND4 (N11875, N11872, N8164, N5460, N333);
or OR2 (N11876, N11863, N4292);
or OR4 (N11877, N11871, N9441, N7192, N9096);
xor XOR2 (N11878, N11874, N4348);
xor XOR2 (N11879, N11875, N11724);
or OR3 (N11880, N11879, N10486, N3856);
xor XOR2 (N11881, N11867, N9723);
not NOT1 (N11882, N11878);
nand NAND2 (N11883, N11864, N4998);
buf BUF1 (N11884, N11876);
nand NAND3 (N11885, N11861, N7127, N8867);
nor NOR4 (N11886, N11880, N11273, N7041, N10435);
nand NAND4 (N11887, N11885, N3582, N2207, N1315);
nand NAND3 (N11888, N11886, N4686, N9187);
and AND2 (N11889, N11865, N190);
xor XOR2 (N11890, N11883, N2149);
or OR4 (N11891, N11784, N2837, N4701, N1775);
or OR4 (N11892, N11868, N4150, N9570, N2299);
buf BUF1 (N11893, N11887);
or OR4 (N11894, N11881, N10408, N10874, N8509);
not NOT1 (N11895, N11884);
xor XOR2 (N11896, N11894, N4684);
and AND2 (N11897, N11882, N7460);
buf BUF1 (N11898, N11893);
nand NAND4 (N11899, N11888, N10573, N4496, N2684);
xor XOR2 (N11900, N11877, N9556);
nand NAND3 (N11901, N11900, N4114, N4659);
buf BUF1 (N11902, N11892);
not NOT1 (N11903, N11889);
xor XOR2 (N11904, N11902, N3208);
or OR3 (N11905, N11901, N2455, N6450);
xor XOR2 (N11906, N11896, N8701);
and AND3 (N11907, N11891, N8122, N9783);
or OR4 (N11908, N11890, N1026, N359, N10254);
buf BUF1 (N11909, N11908);
xor XOR2 (N11910, N11909, N2178);
and AND3 (N11911, N11905, N10037, N2253);
nand NAND3 (N11912, N11903, N7502, N5991);
or OR2 (N11913, N11898, N6625);
or OR4 (N11914, N11906, N6270, N6477, N8615);
nand NAND4 (N11915, N11912, N6032, N11812, N103);
nor NOR3 (N11916, N11914, N11569, N8911);
buf BUF1 (N11917, N11897);
and AND4 (N11918, N11907, N9517, N8184, N6813);
not NOT1 (N11919, N11904);
nor NOR2 (N11920, N11899, N4642);
or OR3 (N11921, N11910, N11666, N9568);
buf BUF1 (N11922, N11918);
nand NAND2 (N11923, N11919, N6248);
and AND2 (N11924, N11917, N5594);
nor NOR3 (N11925, N11895, N1208, N4720);
nand NAND4 (N11926, N11920, N8814, N10167, N9329);
and AND4 (N11927, N11926, N6559, N4369, N6347);
xor XOR2 (N11928, N11927, N11253);
not NOT1 (N11929, N11925);
buf BUF1 (N11930, N11923);
buf BUF1 (N11931, N11929);
buf BUF1 (N11932, N11915);
xor XOR2 (N11933, N11922, N9519);
nand NAND4 (N11934, N11933, N1188, N5208, N7180);
buf BUF1 (N11935, N11916);
buf BUF1 (N11936, N11934);
xor XOR2 (N11937, N11931, N4913);
not NOT1 (N11938, N11921);
and AND2 (N11939, N11911, N5270);
or OR2 (N11940, N11935, N6715);
nor NOR3 (N11941, N11937, N10827, N10741);
and AND3 (N11942, N11930, N11597, N1492);
or OR3 (N11943, N11938, N8125, N6051);
and AND3 (N11944, N11940, N9325, N2307);
nor NOR2 (N11945, N11936, N8635);
xor XOR2 (N11946, N11939, N9447);
buf BUF1 (N11947, N11924);
and AND3 (N11948, N11947, N6192, N10130);
and AND4 (N11949, N11932, N9522, N3716, N5753);
not NOT1 (N11950, N11913);
nor NOR3 (N11951, N11943, N1529, N884);
xor XOR2 (N11952, N11950, N473);
and AND3 (N11953, N11948, N8822, N11766);
nor NOR4 (N11954, N11953, N5738, N11223, N10916);
or OR2 (N11955, N11944, N9469);
or OR2 (N11956, N11946, N7162);
nand NAND4 (N11957, N11952, N8817, N11534, N10396);
buf BUF1 (N11958, N11954);
nand NAND3 (N11959, N11957, N6952, N7501);
buf BUF1 (N11960, N11958);
nor NOR3 (N11961, N11960, N6433, N7266);
buf BUF1 (N11962, N11942);
or OR2 (N11963, N11962, N2928);
nand NAND3 (N11964, N11945, N1855, N4956);
not NOT1 (N11965, N11963);
buf BUF1 (N11966, N11949);
not NOT1 (N11967, N11961);
not NOT1 (N11968, N11967);
xor XOR2 (N11969, N11928, N1477);
and AND2 (N11970, N11955, N6460);
or OR4 (N11971, N11965, N10144, N516, N8645);
xor XOR2 (N11972, N11951, N4204);
buf BUF1 (N11973, N11966);
nand NAND4 (N11974, N11970, N4361, N6152, N8303);
or OR3 (N11975, N11973, N9911, N11646);
not NOT1 (N11976, N11956);
and AND4 (N11977, N11971, N7469, N8352, N11716);
xor XOR2 (N11978, N11941, N6314);
not NOT1 (N11979, N11959);
not NOT1 (N11980, N11976);
not NOT1 (N11981, N11964);
buf BUF1 (N11982, N11974);
nor NOR3 (N11983, N11972, N4631, N7302);
buf BUF1 (N11984, N11980);
nand NAND2 (N11985, N11982, N5961);
xor XOR2 (N11986, N11969, N6615);
nand NAND4 (N11987, N11979, N11832, N6394, N8819);
or OR2 (N11988, N11984, N6591);
nand NAND3 (N11989, N11987, N10351, N4742);
not NOT1 (N11990, N11989);
or OR4 (N11991, N11988, N11267, N8725, N4471);
or OR3 (N11992, N11983, N2241, N3903);
xor XOR2 (N11993, N11975, N1697);
and AND3 (N11994, N11978, N6056, N1830);
not NOT1 (N11995, N11991);
buf BUF1 (N11996, N11977);
buf BUF1 (N11997, N11986);
nand NAND4 (N11998, N11993, N8325, N7628, N2235);
or OR3 (N11999, N11996, N4942, N2860);
and AND2 (N12000, N11994, N4905);
nand NAND3 (N12001, N11981, N8296, N9251);
nor NOR3 (N12002, N11997, N8718, N9567);
or OR2 (N12003, N11995, N3090);
buf BUF1 (N12004, N12002);
buf BUF1 (N12005, N11999);
not NOT1 (N12006, N12005);
and AND4 (N12007, N12003, N11658, N10305, N2800);
and AND3 (N12008, N11992, N4285, N7388);
nor NOR3 (N12009, N11998, N6734, N9607);
xor XOR2 (N12010, N12006, N6066);
or OR4 (N12011, N12007, N2582, N3534, N161);
not NOT1 (N12012, N11968);
and AND4 (N12013, N11985, N4052, N6878, N10671);
buf BUF1 (N12014, N11990);
or OR2 (N12015, N12008, N8702);
or OR4 (N12016, N12010, N11640, N12012, N3355);
buf BUF1 (N12017, N6721);
not NOT1 (N12018, N12014);
or OR3 (N12019, N12000, N4050, N7575);
not NOT1 (N12020, N12013);
or OR2 (N12021, N12011, N2092);
nor NOR2 (N12022, N12004, N4235);
and AND2 (N12023, N12017, N9104);
or OR2 (N12024, N12022, N8513);
and AND3 (N12025, N12024, N4727, N7336);
or OR3 (N12026, N12001, N2933, N5227);
xor XOR2 (N12027, N12023, N10387);
not NOT1 (N12028, N12021);
nor NOR4 (N12029, N12019, N962, N7494, N8743);
xor XOR2 (N12030, N12025, N764);
or OR3 (N12031, N12029, N7718, N6868);
and AND2 (N12032, N12027, N10225);
not NOT1 (N12033, N12009);
nand NAND4 (N12034, N12018, N9677, N1780, N10672);
xor XOR2 (N12035, N12026, N6448);
and AND2 (N12036, N12020, N3741);
nor NOR4 (N12037, N12016, N2674, N3389, N9497);
not NOT1 (N12038, N12031);
xor XOR2 (N12039, N12036, N10197);
buf BUF1 (N12040, N12039);
or OR4 (N12041, N12032, N3261, N8028, N4915);
and AND3 (N12042, N12040, N4895, N4739);
nor NOR4 (N12043, N12028, N11193, N5107, N6611);
and AND3 (N12044, N12030, N6403, N615);
or OR3 (N12045, N12038, N7858, N1542);
not NOT1 (N12046, N12041);
or OR3 (N12047, N12045, N3225, N1904);
nor NOR2 (N12048, N12037, N3187);
and AND2 (N12049, N12015, N8948);
and AND4 (N12050, N12049, N5233, N781, N1594);
not NOT1 (N12051, N12033);
xor XOR2 (N12052, N12047, N3805);
nor NOR2 (N12053, N12052, N1800);
nor NOR2 (N12054, N12051, N6228);
buf BUF1 (N12055, N12050);
nor NOR3 (N12056, N12034, N2909, N7246);
xor XOR2 (N12057, N12044, N3613);
xor XOR2 (N12058, N12042, N9971);
buf BUF1 (N12059, N12048);
and AND4 (N12060, N12035, N6938, N10056, N1057);
xor XOR2 (N12061, N12058, N3657);
or OR3 (N12062, N12061, N5229, N9275);
and AND2 (N12063, N12053, N7463);
xor XOR2 (N12064, N12043, N8920);
or OR4 (N12065, N12046, N3067, N11692, N12055);
xor XOR2 (N12066, N5995, N5);
xor XOR2 (N12067, N12063, N6324);
and AND3 (N12068, N12060, N5206, N5441);
nand NAND4 (N12069, N12068, N699, N1469, N97);
nand NAND4 (N12070, N12054, N5187, N7450, N6820);
xor XOR2 (N12071, N12069, N7621);
nor NOR2 (N12072, N12067, N9194);
and AND2 (N12073, N12066, N4464);
xor XOR2 (N12074, N12072, N7460);
nor NOR2 (N12075, N12059, N9211);
and AND4 (N12076, N12065, N2203, N5993, N3971);
not NOT1 (N12077, N12056);
not NOT1 (N12078, N12071);
buf BUF1 (N12079, N12074);
nand NAND3 (N12080, N12079, N2361, N5845);
nand NAND4 (N12081, N12073, N7712, N3680, N9856);
buf BUF1 (N12082, N12076);
nand NAND3 (N12083, N12082, N6679, N1802);
xor XOR2 (N12084, N12081, N1659);
or OR4 (N12085, N12070, N10850, N3488, N4556);
and AND3 (N12086, N12078, N7528, N5592);
not NOT1 (N12087, N12085);
xor XOR2 (N12088, N12083, N1047);
nand NAND4 (N12089, N12064, N4117, N3092, N6603);
and AND3 (N12090, N12086, N5580, N7837);
and AND4 (N12091, N12075, N9044, N3525, N5106);
nor NOR3 (N12092, N12088, N7200, N8722);
xor XOR2 (N12093, N12090, N8310);
buf BUF1 (N12094, N12077);
nand NAND2 (N12095, N12087, N1972);
xor XOR2 (N12096, N12089, N174);
nor NOR4 (N12097, N12094, N1555, N3257, N2699);
and AND3 (N12098, N12080, N9002, N10522);
nor NOR4 (N12099, N12098, N3133, N5482, N9823);
not NOT1 (N12100, N12084);
xor XOR2 (N12101, N12092, N11221);
or OR2 (N12102, N12062, N11711);
nor NOR4 (N12103, N12101, N1790, N5585, N6175);
or OR3 (N12104, N12102, N10671, N4230);
buf BUF1 (N12105, N12057);
and AND4 (N12106, N12091, N4235, N9354, N8396);
nor NOR2 (N12107, N12095, N1026);
and AND2 (N12108, N12103, N5259);
or OR3 (N12109, N12093, N4955, N7621);
buf BUF1 (N12110, N12106);
nor NOR2 (N12111, N12110, N534);
and AND2 (N12112, N12108, N5139);
nor NOR2 (N12113, N12099, N2710);
not NOT1 (N12114, N12096);
buf BUF1 (N12115, N12114);
nor NOR3 (N12116, N12111, N6731, N6925);
nor NOR3 (N12117, N12105, N8346, N377);
not NOT1 (N12118, N12107);
nand NAND2 (N12119, N12112, N11097);
and AND4 (N12120, N12109, N9096, N10951, N10483);
not NOT1 (N12121, N12100);
not NOT1 (N12122, N12118);
xor XOR2 (N12123, N12120, N4837);
xor XOR2 (N12124, N12123, N688);
or OR4 (N12125, N12121, N9588, N7565, N5938);
nand NAND3 (N12126, N12124, N10715, N4693);
not NOT1 (N12127, N12117);
buf BUF1 (N12128, N12104);
xor XOR2 (N12129, N12128, N11077);
buf BUF1 (N12130, N12115);
or OR2 (N12131, N12116, N7130);
xor XOR2 (N12132, N12122, N1194);
or OR2 (N12133, N12119, N6591);
and AND2 (N12134, N12129, N6701);
not NOT1 (N12135, N12113);
xor XOR2 (N12136, N12133, N1054);
nand NAND3 (N12137, N12097, N9076, N8376);
not NOT1 (N12138, N12125);
or OR4 (N12139, N12127, N8231, N1176, N10431);
and AND3 (N12140, N12126, N7016, N4624);
nor NOR4 (N12141, N12140, N11452, N5927, N1963);
and AND4 (N12142, N12130, N1129, N9813, N1864);
buf BUF1 (N12143, N12136);
xor XOR2 (N12144, N12142, N1618);
or OR2 (N12145, N12138, N1130);
and AND2 (N12146, N12135, N11344);
nor NOR4 (N12147, N12131, N10625, N6972, N1780);
or OR4 (N12148, N12143, N10010, N4889, N5417);
and AND4 (N12149, N12147, N8260, N9914, N7652);
or OR4 (N12150, N12144, N3423, N2160, N7142);
and AND4 (N12151, N12145, N1331, N866, N6240);
xor XOR2 (N12152, N12151, N10092);
or OR2 (N12153, N12137, N1359);
not NOT1 (N12154, N12148);
and AND4 (N12155, N12150, N2440, N1760, N10227);
nand NAND4 (N12156, N12141, N1799, N8099, N11554);
nor NOR3 (N12157, N12149, N9244, N11827);
buf BUF1 (N12158, N12154);
nor NOR4 (N12159, N12153, N7353, N1111, N3531);
nand NAND2 (N12160, N12157, N8881);
xor XOR2 (N12161, N12139, N9658);
and AND2 (N12162, N12146, N10813);
nor NOR4 (N12163, N12158, N4283, N4682, N6402);
xor XOR2 (N12164, N12162, N2122);
nand NAND2 (N12165, N12156, N5016);
buf BUF1 (N12166, N12132);
or OR2 (N12167, N12165, N2410);
buf BUF1 (N12168, N12166);
xor XOR2 (N12169, N12163, N2204);
nor NOR3 (N12170, N12152, N11559, N10389);
not NOT1 (N12171, N12155);
and AND3 (N12172, N12134, N3316, N8533);
nand NAND2 (N12173, N12167, N5204);
nor NOR2 (N12174, N12169, N1819);
nand NAND4 (N12175, N12174, N1098, N6578, N4688);
nor NOR2 (N12176, N12171, N8651);
not NOT1 (N12177, N12160);
or OR3 (N12178, N12176, N8415, N9564);
buf BUF1 (N12179, N12172);
buf BUF1 (N12180, N12178);
xor XOR2 (N12181, N12179, N6141);
and AND2 (N12182, N12180, N7331);
buf BUF1 (N12183, N12159);
not NOT1 (N12184, N12164);
buf BUF1 (N12185, N12161);
xor XOR2 (N12186, N12170, N8267);
not NOT1 (N12187, N12168);
buf BUF1 (N12188, N12181);
nand NAND2 (N12189, N12183, N941);
xor XOR2 (N12190, N12173, N2080);
buf BUF1 (N12191, N12189);
nand NAND2 (N12192, N12184, N1973);
xor XOR2 (N12193, N12185, N2938);
and AND2 (N12194, N12190, N3713);
not NOT1 (N12195, N12193);
nand NAND4 (N12196, N12187, N10849, N8563, N9416);
or OR3 (N12197, N12194, N10710, N1746);
or OR4 (N12198, N12196, N2363, N5482, N5802);
nor NOR3 (N12199, N12197, N11469, N3611);
buf BUF1 (N12200, N12186);
or OR4 (N12201, N12200, N1305, N8093, N11348);
not NOT1 (N12202, N12191);
not NOT1 (N12203, N12177);
buf BUF1 (N12204, N12201);
and AND3 (N12205, N12204, N222, N11309);
nor NOR4 (N12206, N12188, N12019, N1893, N6595);
buf BUF1 (N12207, N12205);
nor NOR3 (N12208, N12198, N3507, N8188);
buf BUF1 (N12209, N12208);
and AND4 (N12210, N12206, N3461, N676, N9262);
not NOT1 (N12211, N12182);
not NOT1 (N12212, N12192);
xor XOR2 (N12213, N12211, N3984);
xor XOR2 (N12214, N12209, N696);
or OR4 (N12215, N12213, N6576, N7169, N1626);
not NOT1 (N12216, N12210);
nand NAND2 (N12217, N12212, N10963);
nor NOR4 (N12218, N12216, N21, N12105, N11543);
and AND2 (N12219, N12202, N11625);
and AND3 (N12220, N12175, N6506, N1952);
and AND4 (N12221, N12195, N5714, N8714, N9608);
or OR4 (N12222, N12203, N2195, N9200, N8159);
or OR2 (N12223, N12214, N1536);
nand NAND3 (N12224, N12215, N4870, N12080);
and AND4 (N12225, N12220, N1031, N6749, N1789);
and AND2 (N12226, N12219, N816);
nor NOR2 (N12227, N12223, N12196);
or OR2 (N12228, N12224, N5268);
and AND4 (N12229, N12222, N7132, N3793, N7639);
and AND2 (N12230, N12218, N8454);
nand NAND4 (N12231, N12227, N2694, N7823, N11049);
nand NAND3 (N12232, N12229, N8155, N5120);
or OR4 (N12233, N12199, N7193, N85, N11714);
buf BUF1 (N12234, N12207);
buf BUF1 (N12235, N12230);
or OR2 (N12236, N12225, N409);
nor NOR2 (N12237, N12233, N2353);
and AND2 (N12238, N12236, N4426);
or OR2 (N12239, N12232, N6547);
and AND4 (N12240, N12234, N8954, N10513, N8487);
buf BUF1 (N12241, N12235);
or OR4 (N12242, N12241, N6178, N10817, N105);
buf BUF1 (N12243, N12217);
not NOT1 (N12244, N12228);
or OR2 (N12245, N12231, N3915);
not NOT1 (N12246, N12243);
xor XOR2 (N12247, N12245, N5703);
or OR2 (N12248, N12246, N8696);
buf BUF1 (N12249, N12242);
xor XOR2 (N12250, N12238, N6703);
or OR2 (N12251, N12239, N10463);
nand NAND3 (N12252, N12249, N11394, N11511);
buf BUF1 (N12253, N12248);
nor NOR3 (N12254, N12226, N12066, N8687);
nand NAND3 (N12255, N12221, N9457, N4374);
not NOT1 (N12256, N12253);
nand NAND4 (N12257, N12240, N7295, N1452, N5095);
xor XOR2 (N12258, N12256, N2687);
and AND2 (N12259, N12252, N4046);
buf BUF1 (N12260, N12259);
not NOT1 (N12261, N12260);
xor XOR2 (N12262, N12244, N3183);
not NOT1 (N12263, N12255);
not NOT1 (N12264, N12254);
not NOT1 (N12265, N12261);
nand NAND4 (N12266, N12237, N1728, N7242, N3291);
xor XOR2 (N12267, N12263, N2730);
or OR4 (N12268, N12258, N2787, N5593, N9945);
not NOT1 (N12269, N12257);
not NOT1 (N12270, N12262);
not NOT1 (N12271, N12265);
and AND2 (N12272, N12266, N1684);
or OR4 (N12273, N12269, N8591, N9369, N6306);
buf BUF1 (N12274, N12267);
not NOT1 (N12275, N12274);
nand NAND3 (N12276, N12250, N10429, N10850);
and AND2 (N12277, N12275, N5901);
nor NOR3 (N12278, N12251, N10950, N6422);
not NOT1 (N12279, N12278);
nand NAND3 (N12280, N12277, N11776, N6066);
and AND4 (N12281, N12273, N3824, N8082, N9520);
or OR4 (N12282, N12247, N11306, N1013, N1648);
or OR4 (N12283, N12272, N8429, N5668, N5152);
buf BUF1 (N12284, N12281);
nor NOR4 (N12285, N12283, N777, N11709, N3791);
and AND4 (N12286, N12264, N3671, N6115, N5964);
or OR2 (N12287, N12282, N5183);
xor XOR2 (N12288, N12286, N11062);
nand NAND4 (N12289, N12284, N2075, N918, N8361);
and AND3 (N12290, N12276, N401, N4843);
nor NOR3 (N12291, N12288, N7864, N8743);
xor XOR2 (N12292, N12268, N4697);
nor NOR3 (N12293, N12289, N617, N8612);
and AND3 (N12294, N12280, N322, N11291);
xor XOR2 (N12295, N12287, N2722);
and AND2 (N12296, N12295, N5257);
buf BUF1 (N12297, N12293);
nor NOR3 (N12298, N12292, N1948, N498);
buf BUF1 (N12299, N12296);
or OR4 (N12300, N12271, N7708, N8115, N5509);
xor XOR2 (N12301, N12297, N7805);
not NOT1 (N12302, N12294);
not NOT1 (N12303, N12300);
nand NAND2 (N12304, N12301, N10617);
or OR4 (N12305, N12302, N4256, N3494, N7484);
buf BUF1 (N12306, N12304);
buf BUF1 (N12307, N12270);
nand NAND2 (N12308, N12305, N1481);
nor NOR4 (N12309, N12299, N2270, N8032, N10796);
not NOT1 (N12310, N12298);
and AND3 (N12311, N12308, N7322, N524);
nor NOR2 (N12312, N12291, N2270);
xor XOR2 (N12313, N12306, N474);
buf BUF1 (N12314, N12303);
and AND3 (N12315, N12307, N6200, N8860);
nand NAND3 (N12316, N12285, N3464, N3177);
or OR2 (N12317, N12290, N2957);
nor NOR4 (N12318, N12310, N975, N7692, N337);
not NOT1 (N12319, N12313);
xor XOR2 (N12320, N12317, N7866);
nand NAND2 (N12321, N12318, N7182);
not NOT1 (N12322, N12311);
buf BUF1 (N12323, N12312);
and AND4 (N12324, N12321, N3259, N7079, N2457);
buf BUF1 (N12325, N12320);
not NOT1 (N12326, N12279);
nand NAND4 (N12327, N12314, N12180, N1432, N11800);
or OR4 (N12328, N12316, N6884, N48, N7184);
not NOT1 (N12329, N12325);
buf BUF1 (N12330, N12328);
and AND2 (N12331, N12324, N5810);
not NOT1 (N12332, N12330);
not NOT1 (N12333, N12322);
or OR4 (N12334, N12315, N11770, N5251, N6847);
nor NOR3 (N12335, N12329, N5033, N9929);
xor XOR2 (N12336, N12309, N9087);
xor XOR2 (N12337, N12319, N2182);
not NOT1 (N12338, N12323);
xor XOR2 (N12339, N12326, N8307);
not NOT1 (N12340, N12335);
not NOT1 (N12341, N12333);
and AND4 (N12342, N12331, N1185, N6873, N7260);
nand NAND2 (N12343, N12342, N4434);
or OR2 (N12344, N12341, N2447);
not NOT1 (N12345, N12334);
nor NOR4 (N12346, N12345, N8990, N742, N5484);
nor NOR2 (N12347, N12344, N11384);
or OR4 (N12348, N12337, N11224, N10676, N6738);
not NOT1 (N12349, N12336);
or OR4 (N12350, N12338, N8017, N3930, N6879);
nor NOR4 (N12351, N12346, N8035, N297, N3891);
or OR4 (N12352, N12340, N1392, N8677, N21);
nor NOR2 (N12353, N12343, N2701);
and AND3 (N12354, N12348, N8394, N214);
nor NOR3 (N12355, N12350, N7400, N257);
buf BUF1 (N12356, N12347);
xor XOR2 (N12357, N12356, N1612);
or OR4 (N12358, N12354, N5078, N9982, N10991);
buf BUF1 (N12359, N12355);
xor XOR2 (N12360, N12349, N7739);
buf BUF1 (N12361, N12352);
nor NOR4 (N12362, N12353, N11070, N1988, N1844);
nor NOR4 (N12363, N12360, N1413, N11132, N9730);
nor NOR4 (N12364, N12361, N3073, N7691, N5957);
and AND2 (N12365, N12357, N521);
nand NAND2 (N12366, N12363, N1712);
or OR2 (N12367, N12365, N4083);
xor XOR2 (N12368, N12364, N10664);
xor XOR2 (N12369, N12359, N11114);
buf BUF1 (N12370, N12327);
nand NAND3 (N12371, N12368, N3936, N9746);
and AND3 (N12372, N12367, N9905, N11623);
nand NAND3 (N12373, N12362, N11140, N3416);
buf BUF1 (N12374, N12371);
nor NOR2 (N12375, N12369, N1087);
buf BUF1 (N12376, N12332);
or OR4 (N12377, N12339, N8869, N7829, N6001);
and AND4 (N12378, N12370, N1567, N8367, N2923);
and AND2 (N12379, N12372, N11968);
nor NOR2 (N12380, N12377, N2574);
nand NAND3 (N12381, N12351, N9607, N8586);
nor NOR4 (N12382, N12374, N76, N7443, N9380);
nor NOR3 (N12383, N12375, N5540, N4866);
buf BUF1 (N12384, N12383);
not NOT1 (N12385, N12376);
xor XOR2 (N12386, N12366, N2164);
xor XOR2 (N12387, N12373, N10581);
buf BUF1 (N12388, N12385);
and AND3 (N12389, N12381, N4006, N10696);
nor NOR3 (N12390, N12388, N4274, N2047);
and AND3 (N12391, N12378, N10202, N204);
nor NOR4 (N12392, N12379, N3365, N9805, N8807);
nand NAND3 (N12393, N12380, N3652, N9542);
buf BUF1 (N12394, N12389);
and AND3 (N12395, N12394, N3233, N562);
xor XOR2 (N12396, N12393, N1781);
and AND2 (N12397, N12387, N7947);
nand NAND3 (N12398, N12384, N1388, N7768);
or OR4 (N12399, N12390, N2253, N11223, N7932);
or OR3 (N12400, N12386, N285, N9006);
or OR4 (N12401, N12400, N4933, N3898, N5115);
buf BUF1 (N12402, N12398);
not NOT1 (N12403, N12391);
nand NAND2 (N12404, N12402, N7379);
nor NOR4 (N12405, N12404, N3719, N9417, N279);
nor NOR3 (N12406, N12358, N2137, N11375);
not NOT1 (N12407, N12405);
and AND2 (N12408, N12403, N3000);
or OR3 (N12409, N12392, N7640, N1753);
xor XOR2 (N12410, N12409, N6985);
xor XOR2 (N12411, N12397, N3935);
buf BUF1 (N12412, N12395);
or OR3 (N12413, N12401, N3059, N83);
nand NAND3 (N12414, N12410, N9536, N12093);
nand NAND2 (N12415, N12407, N6452);
or OR2 (N12416, N12414, N9283);
or OR3 (N12417, N12406, N8163, N3261);
and AND4 (N12418, N12412, N2687, N4966, N11495);
xor XOR2 (N12419, N12382, N1089);
xor XOR2 (N12420, N12411, N4708);
xor XOR2 (N12421, N12396, N6069);
xor XOR2 (N12422, N12420, N9784);
or OR2 (N12423, N12408, N133);
or OR3 (N12424, N12413, N8567, N11581);
nand NAND2 (N12425, N12421, N938);
not NOT1 (N12426, N12399);
or OR4 (N12427, N12419, N8287, N8161, N8652);
nand NAND2 (N12428, N12417, N1026);
buf BUF1 (N12429, N12428);
nand NAND3 (N12430, N12425, N11888, N6367);
nand NAND3 (N12431, N12416, N10131, N12175);
or OR3 (N12432, N12422, N8393, N7846);
and AND2 (N12433, N12415, N8463);
xor XOR2 (N12434, N12433, N15);
not NOT1 (N12435, N12430);
and AND3 (N12436, N12418, N4988, N1367);
or OR4 (N12437, N12424, N11241, N12055, N5238);
buf BUF1 (N12438, N12423);
nand NAND3 (N12439, N12434, N6616, N9026);
buf BUF1 (N12440, N12437);
or OR3 (N12441, N12438, N7358, N4445);
not NOT1 (N12442, N12440);
or OR2 (N12443, N12429, N3280);
not NOT1 (N12444, N12427);
or OR2 (N12445, N12426, N557);
or OR4 (N12446, N12441, N11668, N12022, N639);
not NOT1 (N12447, N12439);
nor NOR3 (N12448, N12442, N11934, N7662);
not NOT1 (N12449, N12435);
or OR3 (N12450, N12449, N3244, N6883);
not NOT1 (N12451, N12448);
and AND4 (N12452, N12444, N10199, N9211, N2059);
xor XOR2 (N12453, N12431, N1836);
and AND4 (N12454, N12447, N2022, N1511, N3140);
nand NAND3 (N12455, N12446, N1250, N6172);
or OR4 (N12456, N12454, N3157, N5316, N7810);
and AND2 (N12457, N12452, N4928);
nor NOR2 (N12458, N12450, N5656);
xor XOR2 (N12459, N12458, N7239);
buf BUF1 (N12460, N12445);
not NOT1 (N12461, N12453);
buf BUF1 (N12462, N12456);
or OR3 (N12463, N12459, N1580, N11639);
buf BUF1 (N12464, N12443);
or OR3 (N12465, N12462, N11834, N11530);
nor NOR2 (N12466, N12457, N10773);
or OR4 (N12467, N12436, N5242, N1884, N1379);
buf BUF1 (N12468, N12455);
and AND2 (N12469, N12464, N3203);
buf BUF1 (N12470, N12460);
nand NAND3 (N12471, N12466, N9377, N1978);
or OR3 (N12472, N12470, N5213, N7362);
and AND2 (N12473, N12451, N2933);
xor XOR2 (N12474, N12472, N10656);
buf BUF1 (N12475, N12463);
or OR3 (N12476, N12467, N4523, N7826);
buf BUF1 (N12477, N12473);
or OR3 (N12478, N12469, N9145, N3653);
nand NAND4 (N12479, N12461, N5751, N1598, N4831);
or OR2 (N12480, N12471, N3123);
nor NOR3 (N12481, N12468, N2300, N9905);
not NOT1 (N12482, N12481);
or OR2 (N12483, N12465, N4382);
not NOT1 (N12484, N12432);
not NOT1 (N12485, N12479);
buf BUF1 (N12486, N12475);
buf BUF1 (N12487, N12486);
nand NAND3 (N12488, N12483, N3948, N4963);
xor XOR2 (N12489, N12482, N5215);
not NOT1 (N12490, N12485);
or OR3 (N12491, N12487, N2161, N3839);
not NOT1 (N12492, N12484);
and AND3 (N12493, N12488, N1702, N11748);
nor NOR3 (N12494, N12492, N2576, N4231);
not NOT1 (N12495, N12491);
or OR2 (N12496, N12474, N2318);
or OR2 (N12497, N12480, N7687);
nor NOR3 (N12498, N12495, N5901, N4241);
not NOT1 (N12499, N12478);
nand NAND4 (N12500, N12494, N500, N7309, N10401);
buf BUF1 (N12501, N12498);
not NOT1 (N12502, N12497);
nor NOR2 (N12503, N12493, N7396);
xor XOR2 (N12504, N12477, N2815);
or OR2 (N12505, N12501, N1221);
xor XOR2 (N12506, N12502, N11526);
and AND2 (N12507, N12496, N10778);
buf BUF1 (N12508, N12505);
or OR4 (N12509, N12507, N2823, N5331, N8232);
and AND2 (N12510, N12500, N6699);
or OR2 (N12511, N12509, N12154);
xor XOR2 (N12512, N12489, N5220);
not NOT1 (N12513, N12511);
nor NOR4 (N12514, N12499, N6256, N11049, N11030);
buf BUF1 (N12515, N12513);
nand NAND3 (N12516, N12514, N10925, N3695);
not NOT1 (N12517, N12504);
and AND2 (N12518, N12476, N10070);
nand NAND3 (N12519, N12490, N9644, N1951);
buf BUF1 (N12520, N12519);
nor NOR3 (N12521, N12508, N3289, N1463);
buf BUF1 (N12522, N12521);
and AND2 (N12523, N12517, N2639);
buf BUF1 (N12524, N12510);
buf BUF1 (N12525, N12516);
nand NAND3 (N12526, N12524, N8813, N2799);
or OR2 (N12527, N12518, N1255);
and AND2 (N12528, N12506, N10820);
nand NAND4 (N12529, N12527, N7292, N11572, N4136);
nor NOR2 (N12530, N12520, N169);
not NOT1 (N12531, N12526);
buf BUF1 (N12532, N12531);
nand NAND3 (N12533, N12523, N11378, N860);
or OR4 (N12534, N12529, N1485, N12505, N9120);
and AND4 (N12535, N12528, N4250, N2269, N8007);
and AND3 (N12536, N12522, N8023, N3229);
nand NAND3 (N12537, N12515, N7092, N8799);
or OR3 (N12538, N12530, N9543, N2359);
nor NOR3 (N12539, N12534, N6167, N295);
or OR2 (N12540, N12503, N6096);
and AND2 (N12541, N12539, N531);
nor NOR2 (N12542, N12533, N4085);
xor XOR2 (N12543, N12537, N3949);
nor NOR4 (N12544, N12542, N6314, N3260, N9091);
and AND2 (N12545, N12536, N7698);
nand NAND4 (N12546, N12512, N1678, N7632, N6686);
or OR2 (N12547, N12545, N10665);
xor XOR2 (N12548, N12538, N11204);
nand NAND4 (N12549, N12546, N10305, N5628, N3759);
nor NOR3 (N12550, N12535, N1111, N1010);
not NOT1 (N12551, N12540);
and AND3 (N12552, N12549, N4081, N886);
not NOT1 (N12553, N12547);
nor NOR3 (N12554, N12551, N3425, N8816);
not NOT1 (N12555, N12554);
nor NOR2 (N12556, N12552, N8280);
xor XOR2 (N12557, N12548, N3779);
nand NAND4 (N12558, N12557, N11978, N3844, N9676);
and AND4 (N12559, N12553, N9356, N7718, N12168);
and AND2 (N12560, N12532, N7175);
buf BUF1 (N12561, N12559);
nand NAND3 (N12562, N12556, N1611, N11986);
xor XOR2 (N12563, N12525, N6261);
or OR2 (N12564, N12543, N2349);
or OR4 (N12565, N12564, N2559, N3051, N3502);
and AND3 (N12566, N12544, N7574, N2746);
not NOT1 (N12567, N12561);
nand NAND4 (N12568, N12558, N3139, N7659, N3782);
and AND3 (N12569, N12563, N1814, N8649);
xor XOR2 (N12570, N12568, N8733);
or OR3 (N12571, N12560, N9001, N4524);
and AND2 (N12572, N12566, N2422);
not NOT1 (N12573, N12570);
xor XOR2 (N12574, N12571, N2896);
or OR4 (N12575, N12541, N8001, N11526, N11280);
and AND4 (N12576, N12573, N4378, N5351, N160);
and AND4 (N12577, N12550, N7205, N300, N5190);
xor XOR2 (N12578, N12577, N9505);
xor XOR2 (N12579, N12574, N7775);
not NOT1 (N12580, N12578);
nand NAND2 (N12581, N12565, N8200);
xor XOR2 (N12582, N12572, N5917);
xor XOR2 (N12583, N12569, N10607);
xor XOR2 (N12584, N12582, N6324);
or OR4 (N12585, N12584, N9177, N157, N2376);
nor NOR3 (N12586, N12562, N7151, N8910);
and AND4 (N12587, N12579, N7574, N10451, N11571);
nor NOR3 (N12588, N12587, N9809, N12541);
xor XOR2 (N12589, N12583, N570);
buf BUF1 (N12590, N12567);
and AND3 (N12591, N12588, N10251, N3476);
xor XOR2 (N12592, N12591, N9941);
and AND3 (N12593, N12581, N11060, N798);
and AND3 (N12594, N12575, N10445, N5522);
nand NAND2 (N12595, N12580, N3333);
not NOT1 (N12596, N12592);
xor XOR2 (N12597, N12593, N11864);
buf BUF1 (N12598, N12596);
nand NAND2 (N12599, N12576, N5039);
not NOT1 (N12600, N12555);
and AND3 (N12601, N12597, N12298, N3616);
or OR3 (N12602, N12601, N10757, N1813);
nor NOR4 (N12603, N12589, N1952, N5173, N5469);
or OR3 (N12604, N12598, N11204, N5717);
nand NAND2 (N12605, N12585, N8437);
and AND4 (N12606, N12605, N5082, N10736, N6531);
and AND2 (N12607, N12602, N11961);
nor NOR4 (N12608, N12604, N10905, N8988, N9529);
or OR4 (N12609, N12594, N1982, N5834, N5758);
nor NOR4 (N12610, N12595, N2378, N620, N10526);
and AND4 (N12611, N12606, N215, N11162, N1043);
buf BUF1 (N12612, N12599);
nand NAND4 (N12613, N12608, N965, N8995, N2505);
nor NOR2 (N12614, N12610, N6906);
and AND2 (N12615, N12600, N824);
and AND2 (N12616, N12611, N937);
not NOT1 (N12617, N12612);
not NOT1 (N12618, N12590);
not NOT1 (N12619, N12617);
nand NAND2 (N12620, N12586, N10449);
or OR3 (N12621, N12619, N9277, N12044);
xor XOR2 (N12622, N12616, N10531);
nor NOR3 (N12623, N12603, N7209, N8566);
nor NOR2 (N12624, N12613, N500);
nor NOR2 (N12625, N12614, N7756);
and AND3 (N12626, N12624, N4736, N2014);
or OR4 (N12627, N12625, N4974, N10345, N4558);
and AND2 (N12628, N12615, N255);
and AND4 (N12629, N12627, N6590, N5473, N8589);
buf BUF1 (N12630, N12609);
not NOT1 (N12631, N12622);
buf BUF1 (N12632, N12618);
xor XOR2 (N12633, N12623, N8989);
nand NAND3 (N12634, N12626, N11904, N7148);
not NOT1 (N12635, N12628);
and AND4 (N12636, N12634, N11626, N5255, N11309);
or OR3 (N12637, N12621, N1064, N2395);
and AND4 (N12638, N12635, N4160, N9944, N3848);
not NOT1 (N12639, N12636);
or OR3 (N12640, N12637, N6385, N12281);
nor NOR3 (N12641, N12632, N499, N10409);
not NOT1 (N12642, N12633);
nor NOR4 (N12643, N12630, N7294, N10995, N11490);
not NOT1 (N12644, N12607);
not NOT1 (N12645, N12640);
xor XOR2 (N12646, N12638, N2740);
xor XOR2 (N12647, N12641, N576);
not NOT1 (N12648, N12643);
and AND2 (N12649, N12644, N3803);
nand NAND2 (N12650, N12631, N9850);
xor XOR2 (N12651, N12648, N158);
not NOT1 (N12652, N12650);
buf BUF1 (N12653, N12652);
xor XOR2 (N12654, N12651, N12302);
and AND2 (N12655, N12654, N8208);
buf BUF1 (N12656, N12649);
buf BUF1 (N12657, N12642);
xor XOR2 (N12658, N12646, N7836);
not NOT1 (N12659, N12645);
not NOT1 (N12660, N12657);
nor NOR4 (N12661, N12655, N3433, N9466, N1308);
nor NOR4 (N12662, N12659, N4165, N8926, N10678);
xor XOR2 (N12663, N12647, N8010);
nand NAND2 (N12664, N12658, N2570);
or OR3 (N12665, N12629, N9619, N10836);
nor NOR3 (N12666, N12620, N78, N9837);
not NOT1 (N12667, N12653);
nand NAND3 (N12668, N12664, N7235, N5357);
or OR2 (N12669, N12662, N578);
not NOT1 (N12670, N12660);
not NOT1 (N12671, N12656);
xor XOR2 (N12672, N12670, N12440);
and AND2 (N12673, N12665, N7161);
xor XOR2 (N12674, N12661, N2383);
nand NAND3 (N12675, N12639, N9106, N4150);
nor NOR3 (N12676, N12673, N12597, N9587);
buf BUF1 (N12677, N12669);
nor NOR4 (N12678, N12668, N1439, N12370, N12666);
or OR2 (N12679, N6127, N2735);
not NOT1 (N12680, N12679);
buf BUF1 (N12681, N12677);
or OR4 (N12682, N12663, N1442, N11512, N4791);
and AND3 (N12683, N12671, N12310, N8985);
not NOT1 (N12684, N12674);
nand NAND3 (N12685, N12667, N4581, N106);
or OR2 (N12686, N12685, N4075);
nand NAND3 (N12687, N12683, N3083, N10719);
nand NAND2 (N12688, N12684, N7381);
buf BUF1 (N12689, N12687);
or OR2 (N12690, N12675, N10012);
buf BUF1 (N12691, N12676);
nor NOR2 (N12692, N12681, N2732);
buf BUF1 (N12693, N12672);
or OR3 (N12694, N12691, N10689, N2026);
or OR4 (N12695, N12688, N9594, N3466, N11720);
or OR2 (N12696, N12678, N11875);
not NOT1 (N12697, N12693);
or OR3 (N12698, N12689, N1936, N816);
nand NAND2 (N12699, N12695, N3527);
not NOT1 (N12700, N12697);
xor XOR2 (N12701, N12694, N7487);
buf BUF1 (N12702, N12701);
or OR3 (N12703, N12698, N1566, N10658);
nor NOR2 (N12704, N12700, N2070);
buf BUF1 (N12705, N12692);
or OR3 (N12706, N12699, N856, N6105);
not NOT1 (N12707, N12704);
xor XOR2 (N12708, N12705, N5651);
xor XOR2 (N12709, N12690, N11248);
nor NOR4 (N12710, N12708, N8167, N5144, N6537);
and AND4 (N12711, N12709, N6289, N5929, N3687);
nand NAND4 (N12712, N12686, N3427, N1241, N12283);
buf BUF1 (N12713, N12696);
buf BUF1 (N12714, N12680);
nand NAND2 (N12715, N12711, N229);
nor NOR4 (N12716, N12706, N4344, N1721, N2217);
or OR3 (N12717, N12703, N7232, N893);
or OR3 (N12718, N12712, N6855, N296);
not NOT1 (N12719, N12715);
or OR3 (N12720, N12717, N6836, N7391);
buf BUF1 (N12721, N12716);
xor XOR2 (N12722, N12721, N9096);
not NOT1 (N12723, N12710);
nor NOR2 (N12724, N12720, N2347);
xor XOR2 (N12725, N12713, N7216);
and AND4 (N12726, N12707, N2043, N2269, N10652);
nand NAND4 (N12727, N12723, N7346, N7113, N8456);
or OR4 (N12728, N12718, N5941, N134, N11680);
buf BUF1 (N12729, N12702);
buf BUF1 (N12730, N12724);
and AND4 (N12731, N12729, N8564, N3545, N10309);
nand NAND4 (N12732, N12725, N4513, N9098, N5632);
nor NOR4 (N12733, N12719, N4635, N9024, N2782);
or OR4 (N12734, N12714, N5129, N3400, N1110);
not NOT1 (N12735, N12727);
not NOT1 (N12736, N12682);
and AND4 (N12737, N12728, N6459, N3538, N1386);
nand NAND3 (N12738, N12737, N7508, N419);
not NOT1 (N12739, N12722);
nand NAND3 (N12740, N12735, N3826, N10721);
and AND4 (N12741, N12739, N703, N10528, N6402);
or OR4 (N12742, N12736, N10951, N8907, N6298);
or OR4 (N12743, N12741, N2165, N7035, N1656);
xor XOR2 (N12744, N12742, N481);
buf BUF1 (N12745, N12726);
nand NAND3 (N12746, N12730, N5360, N4400);
not NOT1 (N12747, N12738);
buf BUF1 (N12748, N12733);
or OR4 (N12749, N12746, N199, N4208, N11113);
or OR3 (N12750, N12749, N7258, N1755);
and AND2 (N12751, N12750, N3847);
not NOT1 (N12752, N12740);
and AND3 (N12753, N12747, N7962, N2678);
not NOT1 (N12754, N12751);
xor XOR2 (N12755, N12753, N8696);
nand NAND2 (N12756, N12743, N8536);
not NOT1 (N12757, N12744);
not NOT1 (N12758, N12748);
or OR2 (N12759, N12731, N9689);
nand NAND4 (N12760, N12732, N9579, N7760, N8218);
xor XOR2 (N12761, N12754, N3874);
or OR2 (N12762, N12752, N2502);
nor NOR3 (N12763, N12762, N8555, N5368);
and AND4 (N12764, N12759, N11733, N2847, N141);
nand NAND4 (N12765, N12761, N9984, N3626, N3732);
nand NAND4 (N12766, N12755, N8267, N1684, N7172);
or OR3 (N12767, N12758, N7544, N11760);
nand NAND2 (N12768, N12760, N11882);
nor NOR3 (N12769, N12734, N3388, N9395);
or OR3 (N12770, N12764, N4383, N2396);
and AND2 (N12771, N12769, N6316);
not NOT1 (N12772, N12763);
or OR3 (N12773, N12768, N2253, N11164);
and AND2 (N12774, N12757, N7194);
nand NAND2 (N12775, N12745, N8892);
not NOT1 (N12776, N12756);
nand NAND4 (N12777, N12773, N3898, N7895, N2735);
buf BUF1 (N12778, N12777);
not NOT1 (N12779, N12771);
or OR4 (N12780, N12776, N7245, N5906, N6868);
or OR3 (N12781, N12767, N839, N5341);
not NOT1 (N12782, N12781);
or OR2 (N12783, N12766, N4595);
or OR3 (N12784, N12778, N4793, N9153);
buf BUF1 (N12785, N12774);
xor XOR2 (N12786, N12783, N7442);
nand NAND2 (N12787, N12780, N6226);
xor XOR2 (N12788, N12782, N1132);
or OR3 (N12789, N12786, N8891, N413);
nor NOR2 (N12790, N12775, N1181);
buf BUF1 (N12791, N12790);
not NOT1 (N12792, N12770);
nor NOR3 (N12793, N12788, N10503, N4424);
or OR4 (N12794, N12779, N6084, N10423, N3495);
and AND4 (N12795, N12791, N6172, N11672, N8915);
nand NAND3 (N12796, N12789, N8490, N12016);
xor XOR2 (N12797, N12784, N9544);
xor XOR2 (N12798, N12796, N1876);
or OR4 (N12799, N12765, N10442, N5761, N10066);
nor NOR4 (N12800, N12787, N5086, N11248, N12144);
or OR3 (N12801, N12795, N9523, N10893);
nand NAND4 (N12802, N12798, N3107, N5775, N1422);
and AND4 (N12803, N12772, N9321, N1912, N11601);
buf BUF1 (N12804, N12794);
and AND3 (N12805, N12804, N3981, N2802);
not NOT1 (N12806, N12793);
and AND4 (N12807, N12797, N952, N1212, N5427);
buf BUF1 (N12808, N12806);
xor XOR2 (N12809, N12800, N7939);
nand NAND2 (N12810, N12802, N12736);
or OR2 (N12811, N12803, N1938);
not NOT1 (N12812, N12807);
and AND3 (N12813, N12805, N2649, N3563);
buf BUF1 (N12814, N12813);
buf BUF1 (N12815, N12801);
not NOT1 (N12816, N12809);
xor XOR2 (N12817, N12811, N9928);
not NOT1 (N12818, N12817);
xor XOR2 (N12819, N12818, N4240);
nor NOR4 (N12820, N12799, N8179, N1195, N3834);
nor NOR3 (N12821, N12792, N7821, N7069);
not NOT1 (N12822, N12808);
xor XOR2 (N12823, N12816, N7358);
and AND2 (N12824, N12823, N9494);
or OR3 (N12825, N12812, N12778, N3697);
nor NOR3 (N12826, N12815, N1802, N3885);
or OR2 (N12827, N12810, N572);
not NOT1 (N12828, N12821);
buf BUF1 (N12829, N12820);
nor NOR2 (N12830, N12829, N6338);
buf BUF1 (N12831, N12785);
or OR3 (N12832, N12827, N10138, N10112);
nand NAND2 (N12833, N12824, N2569);
not NOT1 (N12834, N12826);
nand NAND4 (N12835, N12825, N3258, N6928, N5311);
not NOT1 (N12836, N12835);
and AND3 (N12837, N12830, N8431, N9110);
not NOT1 (N12838, N12834);
or OR4 (N12839, N12819, N401, N103, N4954);
xor XOR2 (N12840, N12831, N5332);
and AND2 (N12841, N12833, N11068);
nand NAND4 (N12842, N12836, N11206, N211, N1937);
not NOT1 (N12843, N12832);
and AND4 (N12844, N12828, N12126, N2353, N1467);
nand NAND2 (N12845, N12839, N9226);
and AND4 (N12846, N12838, N5233, N6302, N6904);
not NOT1 (N12847, N12822);
and AND3 (N12848, N12845, N9850, N8601);
and AND2 (N12849, N12842, N970);
nor NOR2 (N12850, N12843, N5396);
buf BUF1 (N12851, N12837);
xor XOR2 (N12852, N12844, N11045);
xor XOR2 (N12853, N12814, N9006);
or OR2 (N12854, N12852, N8549);
not NOT1 (N12855, N12854);
nand NAND3 (N12856, N12841, N7580, N368);
not NOT1 (N12857, N12848);
nand NAND4 (N12858, N12855, N4160, N2870, N5721);
xor XOR2 (N12859, N12858, N2594);
buf BUF1 (N12860, N12840);
and AND4 (N12861, N12849, N12409, N530, N6247);
buf BUF1 (N12862, N12859);
nand NAND2 (N12863, N12860, N7142);
and AND3 (N12864, N12846, N7318, N11);
xor XOR2 (N12865, N12850, N7485);
xor XOR2 (N12866, N12847, N11052);
or OR4 (N12867, N12864, N6219, N12165, N10491);
not NOT1 (N12868, N12853);
and AND2 (N12869, N12857, N12144);
buf BUF1 (N12870, N12869);
or OR3 (N12871, N12863, N5887, N7454);
nor NOR4 (N12872, N12867, N8398, N8029, N601);
xor XOR2 (N12873, N12868, N7935);
and AND4 (N12874, N12862, N11456, N4668, N10158);
not NOT1 (N12875, N12874);
nor NOR2 (N12876, N12873, N5373);
nand NAND2 (N12877, N12876, N4557);
not NOT1 (N12878, N12875);
buf BUF1 (N12879, N12865);
and AND4 (N12880, N12872, N2058, N469, N8057);
not NOT1 (N12881, N12851);
nand NAND3 (N12882, N12870, N11196, N8172);
buf BUF1 (N12883, N12861);
nand NAND3 (N12884, N12856, N10838, N11491);
nor NOR4 (N12885, N12871, N2023, N4170, N4227);
and AND4 (N12886, N12882, N6434, N7438, N8025);
xor XOR2 (N12887, N12884, N8283);
buf BUF1 (N12888, N12885);
nor NOR2 (N12889, N12866, N7965);
or OR3 (N12890, N12880, N505, N193);
nand NAND3 (N12891, N12890, N5942, N6532);
or OR4 (N12892, N12888, N1016, N8578, N6403);
nor NOR3 (N12893, N12886, N9683, N10881);
buf BUF1 (N12894, N12887);
and AND4 (N12895, N12891, N1209, N12475, N694);
or OR2 (N12896, N12883, N11761);
or OR3 (N12897, N12889, N7537, N7707);
xor XOR2 (N12898, N12879, N1279);
xor XOR2 (N12899, N12892, N10969);
and AND4 (N12900, N12878, N154, N6490, N10107);
nand NAND3 (N12901, N12896, N6767, N1395);
nand NAND3 (N12902, N12899, N2556, N1295);
or OR3 (N12903, N12877, N9845, N8695);
not NOT1 (N12904, N12881);
and AND3 (N12905, N12902, N6183, N8694);
xor XOR2 (N12906, N12894, N4495);
buf BUF1 (N12907, N12900);
and AND4 (N12908, N12907, N11104, N4560, N10226);
buf BUF1 (N12909, N12908);
buf BUF1 (N12910, N12906);
nand NAND3 (N12911, N12897, N2259, N12579);
or OR2 (N12912, N12895, N11091);
xor XOR2 (N12913, N12898, N3401);
nor NOR3 (N12914, N12910, N5213, N10630);
nor NOR2 (N12915, N12904, N7508);
not NOT1 (N12916, N12893);
or OR2 (N12917, N12913, N12747);
or OR2 (N12918, N12901, N787);
buf BUF1 (N12919, N12917);
xor XOR2 (N12920, N12919, N5192);
buf BUF1 (N12921, N12920);
or OR4 (N12922, N12914, N10286, N10648, N1677);
not NOT1 (N12923, N12909);
nand NAND4 (N12924, N12905, N1629, N12394, N11190);
or OR3 (N12925, N12921, N12860, N10863);
and AND4 (N12926, N12925, N1569, N6260, N12219);
and AND4 (N12927, N12915, N973, N99, N2128);
not NOT1 (N12928, N12903);
buf BUF1 (N12929, N12924);
nand NAND3 (N12930, N12922, N12536, N9891);
xor XOR2 (N12931, N12916, N12725);
nand NAND3 (N12932, N12930, N8819, N10671);
buf BUF1 (N12933, N12918);
not NOT1 (N12934, N12911);
or OR4 (N12935, N12934, N526, N12145, N900);
xor XOR2 (N12936, N12928, N9386);
not NOT1 (N12937, N12927);
buf BUF1 (N12938, N12923);
xor XOR2 (N12939, N12933, N10254);
xor XOR2 (N12940, N12938, N1614);
nor NOR4 (N12941, N12935, N5354, N1837, N10826);
nand NAND2 (N12942, N12940, N10595);
nand NAND2 (N12943, N12929, N5339);
not NOT1 (N12944, N12937);
or OR2 (N12945, N12944, N530);
nand NAND3 (N12946, N12931, N12213, N6386);
not NOT1 (N12947, N12946);
buf BUF1 (N12948, N12947);
buf BUF1 (N12949, N12948);
nand NAND4 (N12950, N12932, N6328, N3300, N4443);
buf BUF1 (N12951, N12942);
nor NOR4 (N12952, N12945, N7432, N3867, N1647);
or OR3 (N12953, N12941, N7990, N7424);
buf BUF1 (N12954, N12912);
buf BUF1 (N12955, N12954);
nor NOR4 (N12956, N12949, N11993, N6476, N12139);
or OR4 (N12957, N12956, N11241, N1378, N5053);
xor XOR2 (N12958, N12939, N11062);
buf BUF1 (N12959, N12950);
nand NAND3 (N12960, N12926, N1416, N2667);
not NOT1 (N12961, N12959);
or OR3 (N12962, N12957, N4409, N1050);
buf BUF1 (N12963, N12952);
nor NOR3 (N12964, N12960, N1059, N9219);
or OR2 (N12965, N12964, N10692);
nor NOR2 (N12966, N12951, N2236);
and AND2 (N12967, N12963, N6187);
nand NAND4 (N12968, N12966, N4008, N7117, N10456);
buf BUF1 (N12969, N12962);
xor XOR2 (N12970, N12953, N5329);
nand NAND2 (N12971, N12958, N2945);
nand NAND2 (N12972, N12971, N6394);
nor NOR2 (N12973, N12972, N8468);
not NOT1 (N12974, N12967);
buf BUF1 (N12975, N12936);
not NOT1 (N12976, N12969);
nand NAND4 (N12977, N12973, N2840, N6910, N1722);
not NOT1 (N12978, N12961);
and AND3 (N12979, N12965, N3891, N8689);
and AND3 (N12980, N12979, N8960, N7795);
not NOT1 (N12981, N12975);
nand NAND2 (N12982, N12980, N3999);
buf BUF1 (N12983, N12976);
or OR4 (N12984, N12977, N117, N4163, N7727);
nor NOR2 (N12985, N12955, N2663);
nand NAND3 (N12986, N12943, N8753, N12637);
and AND3 (N12987, N12986, N1993, N6647);
and AND4 (N12988, N12968, N2792, N9776, N4522);
and AND3 (N12989, N12983, N5683, N11521);
nand NAND2 (N12990, N12982, N7794);
nor NOR3 (N12991, N12981, N7694, N2252);
buf BUF1 (N12992, N12984);
buf BUF1 (N12993, N12987);
nand NAND3 (N12994, N12990, N9109, N2818);
and AND2 (N12995, N12993, N11122);
and AND4 (N12996, N12995, N5656, N7339, N9449);
nor NOR4 (N12997, N12996, N3229, N9553, N2432);
buf BUF1 (N12998, N12985);
xor XOR2 (N12999, N12991, N12789);
not NOT1 (N13000, N12997);
nor NOR3 (N13001, N12978, N10626, N9099);
or OR2 (N13002, N12974, N3794);
or OR4 (N13003, N12992, N1945, N12934, N12989);
and AND4 (N13004, N1406, N8075, N4649, N1828);
or OR2 (N13005, N12994, N11602);
nor NOR2 (N13006, N13002, N12938);
and AND3 (N13007, N13005, N3595, N5853);
not NOT1 (N13008, N12988);
and AND2 (N13009, N13007, N9694);
and AND3 (N13010, N12999, N5068, N11839);
nor NOR2 (N13011, N13003, N7656);
nand NAND2 (N13012, N13004, N8142);
xor XOR2 (N13013, N13008, N8753);
not NOT1 (N13014, N13013);
and AND2 (N13015, N13012, N7062);
or OR4 (N13016, N13010, N9504, N8027, N7078);
xor XOR2 (N13017, N12970, N10363);
buf BUF1 (N13018, N13017);
nand NAND3 (N13019, N13000, N7735, N4430);
nor NOR2 (N13020, N13006, N4206);
buf BUF1 (N13021, N13011);
not NOT1 (N13022, N13009);
buf BUF1 (N13023, N13001);
xor XOR2 (N13024, N13015, N5819);
nor NOR2 (N13025, N13023, N431);
not NOT1 (N13026, N13025);
or OR3 (N13027, N13018, N844, N11450);
not NOT1 (N13028, N12998);
not NOT1 (N13029, N13019);
nor NOR4 (N13030, N13024, N6983, N7312, N924);
buf BUF1 (N13031, N13029);
not NOT1 (N13032, N13020);
nand NAND4 (N13033, N13030, N4658, N4403, N9382);
or OR2 (N13034, N13022, N2437);
nor NOR2 (N13035, N13033, N7804);
nor NOR4 (N13036, N13021, N891, N7554, N1768);
nor NOR4 (N13037, N13026, N8847, N11031, N12100);
or OR2 (N13038, N13016, N8183);
and AND2 (N13039, N13035, N5228);
and AND4 (N13040, N13039, N9661, N1310, N11733);
buf BUF1 (N13041, N13031);
or OR2 (N13042, N13038, N8408);
buf BUF1 (N13043, N13040);
xor XOR2 (N13044, N13043, N6463);
xor XOR2 (N13045, N13032, N6450);
xor XOR2 (N13046, N13045, N5796);
buf BUF1 (N13047, N13034);
and AND3 (N13048, N13042, N1344, N4787);
nor NOR3 (N13049, N13041, N9701, N3619);
nand NAND4 (N13050, N13044, N8414, N2151, N8569);
not NOT1 (N13051, N13048);
not NOT1 (N13052, N13014);
nand NAND2 (N13053, N13036, N11854);
nand NAND2 (N13054, N13051, N1915);
xor XOR2 (N13055, N13053, N9432);
or OR4 (N13056, N13046, N2862, N7177, N553);
buf BUF1 (N13057, N13050);
xor XOR2 (N13058, N13037, N11264);
nand NAND4 (N13059, N13056, N2159, N13032, N9);
nand NAND4 (N13060, N13049, N5205, N10799, N11316);
or OR2 (N13061, N13054, N2802);
not NOT1 (N13062, N13060);
nor NOR3 (N13063, N13058, N12474, N10618);
not NOT1 (N13064, N13057);
nand NAND4 (N13065, N13062, N8924, N8900, N8984);
and AND4 (N13066, N13055, N12813, N4796, N10811);
not NOT1 (N13067, N13047);
and AND3 (N13068, N13061, N4869, N737);
and AND4 (N13069, N13052, N9368, N171, N3993);
buf BUF1 (N13070, N13066);
buf BUF1 (N13071, N13064);
or OR3 (N13072, N13063, N5535, N10401);
nor NOR4 (N13073, N13070, N3961, N9278, N12040);
not NOT1 (N13074, N13027);
nor NOR2 (N13075, N13068, N12203);
and AND2 (N13076, N13059, N3351);
nand NAND3 (N13077, N13071, N70, N1514);
and AND2 (N13078, N13076, N1259);
nand NAND4 (N13079, N13067, N4915, N3581, N9675);
xor XOR2 (N13080, N13074, N9941);
nor NOR2 (N13081, N13069, N5396);
not NOT1 (N13082, N13080);
and AND3 (N13083, N13078, N12748, N5451);
or OR2 (N13084, N13081, N5641);
nand NAND4 (N13085, N13028, N3101, N6767, N11467);
xor XOR2 (N13086, N13079, N8783);
or OR3 (N13087, N13086, N11032, N11724);
and AND3 (N13088, N13084, N1325, N2957);
xor XOR2 (N13089, N13072, N8275);
nor NOR3 (N13090, N13082, N6655, N10481);
not NOT1 (N13091, N13088);
nand NAND3 (N13092, N13089, N11695, N5233);
nand NAND2 (N13093, N13092, N6943);
nor NOR3 (N13094, N13073, N11489, N9717);
nor NOR2 (N13095, N13093, N10917);
buf BUF1 (N13096, N13090);
and AND2 (N13097, N13095, N4356);
nor NOR2 (N13098, N13065, N10744);
nor NOR4 (N13099, N13097, N10059, N6954, N7101);
nand NAND3 (N13100, N13091, N405, N4035);
or OR4 (N13101, N13075, N63, N1085, N3283);
and AND2 (N13102, N13100, N915);
nand NAND2 (N13103, N13102, N10966);
buf BUF1 (N13104, N13094);
xor XOR2 (N13105, N13103, N8199);
buf BUF1 (N13106, N13096);
xor XOR2 (N13107, N13085, N348);
nand NAND2 (N13108, N13101, N4772);
or OR4 (N13109, N13108, N68, N2857, N3867);
and AND4 (N13110, N13105, N4198, N1581, N6989);
nor NOR4 (N13111, N13099, N2625, N6043, N4263);
nand NAND4 (N13112, N13077, N3614, N252, N1872);
nor NOR3 (N13113, N13110, N3167, N807);
buf BUF1 (N13114, N13113);
not NOT1 (N13115, N13104);
xor XOR2 (N13116, N13114, N12958);
xor XOR2 (N13117, N13116, N882);
or OR2 (N13118, N13115, N6750);
xor XOR2 (N13119, N13098, N7582);
or OR4 (N13120, N13119, N11873, N9074, N10777);
and AND2 (N13121, N13111, N6348);
nor NOR3 (N13122, N13107, N1823, N4684);
buf BUF1 (N13123, N13118);
or OR3 (N13124, N13120, N6204, N3788);
and AND4 (N13125, N13121, N12513, N4050, N8740);
not NOT1 (N13126, N13122);
nand NAND3 (N13127, N13112, N1003, N2611);
not NOT1 (N13128, N13083);
and AND3 (N13129, N13124, N7732, N5858);
xor XOR2 (N13130, N13106, N7987);
and AND2 (N13131, N13128, N8935);
and AND3 (N13132, N13117, N9905, N8732);
xor XOR2 (N13133, N13132, N11758);
xor XOR2 (N13134, N13125, N5820);
nand NAND4 (N13135, N13127, N13110, N1121, N2434);
buf BUF1 (N13136, N13087);
not NOT1 (N13137, N13131);
nand NAND3 (N13138, N13137, N1612, N11484);
not NOT1 (N13139, N13133);
buf BUF1 (N13140, N13130);
or OR4 (N13141, N13129, N7321, N10586, N4006);
nor NOR2 (N13142, N13135, N4513);
or OR2 (N13143, N13134, N10308);
or OR2 (N13144, N13139, N12038);
and AND3 (N13145, N13136, N832, N779);
nand NAND4 (N13146, N13109, N5862, N2585, N7584);
not NOT1 (N13147, N13123);
nor NOR2 (N13148, N13146, N640);
or OR2 (N13149, N13147, N788);
xor XOR2 (N13150, N13142, N10427);
buf BUF1 (N13151, N13126);
not NOT1 (N13152, N13148);
xor XOR2 (N13153, N13141, N2987);
xor XOR2 (N13154, N13151, N8430);
nor NOR2 (N13155, N13152, N1674);
or OR3 (N13156, N13154, N863, N12920);
nand NAND2 (N13157, N13144, N11763);
nand NAND3 (N13158, N13138, N6182, N9023);
and AND4 (N13159, N13149, N4955, N3973, N7605);
nand NAND4 (N13160, N13143, N9467, N3680, N10193);
and AND2 (N13161, N13160, N11411);
not NOT1 (N13162, N13153);
buf BUF1 (N13163, N13145);
nand NAND3 (N13164, N13162, N8280, N9792);
nand NAND3 (N13165, N13161, N11638, N1303);
not NOT1 (N13166, N13155);
or OR4 (N13167, N13158, N2283, N5402, N2560);
not NOT1 (N13168, N13156);
buf BUF1 (N13169, N13164);
nor NOR4 (N13170, N13157, N1836, N7490, N845);
and AND3 (N13171, N13159, N10101, N270);
buf BUF1 (N13172, N13170);
xor XOR2 (N13173, N13166, N1336);
nand NAND2 (N13174, N13172, N5501);
or OR2 (N13175, N13171, N4471);
xor XOR2 (N13176, N13167, N6391);
not NOT1 (N13177, N13173);
or OR2 (N13178, N13174, N3295);
not NOT1 (N13179, N13165);
nand NAND3 (N13180, N13177, N5415, N13066);
nand NAND3 (N13181, N13178, N9377, N8922);
buf BUF1 (N13182, N13179);
nand NAND3 (N13183, N13150, N9015, N6332);
buf BUF1 (N13184, N13169);
not NOT1 (N13185, N13175);
or OR4 (N13186, N13184, N2595, N10016, N2182);
and AND4 (N13187, N13180, N5944, N7137, N8916);
nand NAND2 (N13188, N13181, N13105);
buf BUF1 (N13189, N13187);
buf BUF1 (N13190, N13186);
not NOT1 (N13191, N13190);
nor NOR4 (N13192, N13168, N3589, N13099, N2450);
nor NOR2 (N13193, N13189, N11845);
xor XOR2 (N13194, N13188, N6681);
not NOT1 (N13195, N13191);
not NOT1 (N13196, N13140);
or OR4 (N13197, N13183, N8526, N4320, N9372);
buf BUF1 (N13198, N13176);
xor XOR2 (N13199, N13193, N371);
not NOT1 (N13200, N13197);
xor XOR2 (N13201, N13192, N10386);
or OR2 (N13202, N13199, N9994);
and AND2 (N13203, N13195, N1055);
buf BUF1 (N13204, N13201);
or OR2 (N13205, N13163, N7941);
nand NAND3 (N13206, N13203, N1443, N6258);
nor NOR4 (N13207, N13206, N2439, N12736, N12749);
and AND4 (N13208, N13200, N11288, N5516, N1180);
buf BUF1 (N13209, N13196);
or OR3 (N13210, N13182, N13018, N525);
nand NAND3 (N13211, N13194, N9182, N1043);
xor XOR2 (N13212, N13185, N6920);
nand NAND4 (N13213, N13208, N11548, N5030, N12026);
buf BUF1 (N13214, N13205);
nand NAND2 (N13215, N13207, N11994);
not NOT1 (N13216, N13204);
xor XOR2 (N13217, N13213, N10862);
or OR4 (N13218, N13217, N11898, N10861, N9191);
xor XOR2 (N13219, N13214, N2873);
nand NAND3 (N13220, N13209, N2457, N5078);
or OR2 (N13221, N13202, N1753);
and AND4 (N13222, N13221, N9871, N1218, N10299);
nand NAND2 (N13223, N13212, N3890);
nand NAND3 (N13224, N13215, N4393, N9720);
xor XOR2 (N13225, N13210, N7636);
buf BUF1 (N13226, N13222);
nand NAND3 (N13227, N13223, N1435, N10626);
or OR3 (N13228, N13211, N171, N7562);
buf BUF1 (N13229, N13226);
buf BUF1 (N13230, N13219);
or OR2 (N13231, N13224, N219);
and AND3 (N13232, N13225, N3311, N7557);
or OR3 (N13233, N13230, N1657, N8459);
or OR4 (N13234, N13233, N7587, N7312, N757);
or OR3 (N13235, N13228, N2250, N486);
buf BUF1 (N13236, N13229);
or OR2 (N13237, N13227, N994);
or OR2 (N13238, N13216, N6321);
not NOT1 (N13239, N13231);
nand NAND4 (N13240, N13239, N11006, N6622, N9175);
buf BUF1 (N13241, N13237);
not NOT1 (N13242, N13198);
not NOT1 (N13243, N13236);
nand NAND4 (N13244, N13220, N7438, N5240, N3097);
xor XOR2 (N13245, N13241, N8767);
and AND4 (N13246, N13242, N9168, N11070, N9126);
or OR2 (N13247, N13244, N6813);
xor XOR2 (N13248, N13238, N3844);
nand NAND3 (N13249, N13232, N1070, N9482);
nor NOR4 (N13250, N13234, N11632, N362, N1857);
nor NOR3 (N13251, N13218, N12463, N10367);
nor NOR2 (N13252, N13235, N5443);
buf BUF1 (N13253, N13240);
or OR4 (N13254, N13249, N1746, N9329, N2623);
and AND3 (N13255, N13243, N4175, N3392);
nand NAND2 (N13256, N13250, N6377);
nand NAND2 (N13257, N13254, N10994);
not NOT1 (N13258, N13253);
not NOT1 (N13259, N13251);
nor NOR4 (N13260, N13257, N13031, N3576, N11731);
not NOT1 (N13261, N13256);
xor XOR2 (N13262, N13247, N12999);
and AND2 (N13263, N13258, N1464);
not NOT1 (N13264, N13263);
not NOT1 (N13265, N13262);
not NOT1 (N13266, N13245);
nand NAND2 (N13267, N13252, N9833);
and AND3 (N13268, N13266, N6770, N1621);
nor NOR4 (N13269, N13246, N421, N6094, N8567);
buf BUF1 (N13270, N13261);
or OR2 (N13271, N13267, N2747);
and AND2 (N13272, N13265, N5382);
nor NOR3 (N13273, N13272, N2751, N7457);
nand NAND2 (N13274, N13248, N5827);
buf BUF1 (N13275, N13269);
not NOT1 (N13276, N13270);
and AND2 (N13277, N13264, N11019);
nand NAND4 (N13278, N13273, N2754, N1134, N6366);
or OR2 (N13279, N13278, N7827);
not NOT1 (N13280, N13275);
nand NAND2 (N13281, N13279, N3230);
xor XOR2 (N13282, N13271, N1198);
nand NAND2 (N13283, N13268, N8379);
not NOT1 (N13284, N13274);
buf BUF1 (N13285, N13255);
buf BUF1 (N13286, N13260);
or OR3 (N13287, N13281, N10494, N13113);
or OR2 (N13288, N13284, N10637);
buf BUF1 (N13289, N13285);
not NOT1 (N13290, N13286);
buf BUF1 (N13291, N13288);
buf BUF1 (N13292, N13283);
not NOT1 (N13293, N13259);
and AND3 (N13294, N13292, N13206, N12711);
not NOT1 (N13295, N13277);
nor NOR2 (N13296, N13294, N11981);
or OR3 (N13297, N13293, N13102, N10796);
buf BUF1 (N13298, N13296);
nor NOR3 (N13299, N13290, N12268, N3779);
buf BUF1 (N13300, N13295);
and AND2 (N13301, N13299, N3411);
nand NAND2 (N13302, N13300, N1048);
and AND2 (N13303, N13302, N4623);
xor XOR2 (N13304, N13298, N6282);
nor NOR4 (N13305, N13276, N7318, N10452, N9664);
and AND3 (N13306, N13282, N2986, N12646);
xor XOR2 (N13307, N13291, N11021);
and AND4 (N13308, N13303, N12564, N9097, N6921);
buf BUF1 (N13309, N13287);
nor NOR3 (N13310, N13297, N9556, N395);
buf BUF1 (N13311, N13310);
xor XOR2 (N13312, N13311, N2785);
xor XOR2 (N13313, N13312, N912);
or OR4 (N13314, N13309, N4294, N12739, N5172);
xor XOR2 (N13315, N13289, N7535);
and AND2 (N13316, N13307, N4989);
buf BUF1 (N13317, N13316);
buf BUF1 (N13318, N13314);
and AND4 (N13319, N13304, N1752, N5878, N4153);
nor NOR4 (N13320, N13319, N5248, N10764, N4233);
nand NAND2 (N13321, N13313, N5854);
and AND2 (N13322, N13320, N10214);
buf BUF1 (N13323, N13317);
and AND2 (N13324, N13308, N5795);
and AND4 (N13325, N13306, N506, N4908, N11415);
or OR4 (N13326, N13323, N5342, N2007, N7937);
nor NOR4 (N13327, N13315, N9746, N607, N13318);
not NOT1 (N13328, N1799);
buf BUF1 (N13329, N13301);
and AND4 (N13330, N13321, N9302, N3548, N1847);
or OR4 (N13331, N13322, N1591, N799, N1845);
not NOT1 (N13332, N13324);
not NOT1 (N13333, N13326);
not NOT1 (N13334, N13331);
xor XOR2 (N13335, N13329, N11515);
and AND2 (N13336, N13280, N7874);
xor XOR2 (N13337, N13327, N2883);
or OR4 (N13338, N13330, N1923, N10358, N8505);
xor XOR2 (N13339, N13337, N11626);
nand NAND4 (N13340, N13325, N10466, N4576, N13299);
buf BUF1 (N13341, N13333);
not NOT1 (N13342, N13338);
nand NAND3 (N13343, N13340, N3642, N12678);
not NOT1 (N13344, N13305);
and AND2 (N13345, N13335, N10431);
buf BUF1 (N13346, N13344);
nand NAND3 (N13347, N13341, N10822, N3583);
xor XOR2 (N13348, N13328, N5632);
nor NOR3 (N13349, N13345, N3072, N11855);
buf BUF1 (N13350, N13332);
nand NAND2 (N13351, N13346, N4908);
and AND2 (N13352, N13343, N8326);
and AND3 (N13353, N13342, N11257, N3579);
or OR4 (N13354, N13353, N7835, N1872, N2403);
nor NOR3 (N13355, N13352, N5665, N3269);
or OR2 (N13356, N13347, N9623);
nand NAND3 (N13357, N13356, N121, N7520);
or OR3 (N13358, N13348, N10760, N12074);
nand NAND2 (N13359, N13355, N2290);
and AND2 (N13360, N13357, N4408);
not NOT1 (N13361, N13351);
or OR2 (N13362, N13358, N9173);
not NOT1 (N13363, N13334);
or OR2 (N13364, N13359, N5219);
not NOT1 (N13365, N13361);
nand NAND2 (N13366, N13336, N9609);
nand NAND4 (N13367, N13354, N3206, N12473, N10169);
and AND4 (N13368, N13366, N2053, N12747, N9692);
nand NAND4 (N13369, N13367, N6901, N5719, N7087);
and AND2 (N13370, N13369, N6314);
nand NAND4 (N13371, N13349, N7431, N1502, N6089);
xor XOR2 (N13372, N13362, N8443);
not NOT1 (N13373, N13363);
xor XOR2 (N13374, N13350, N8653);
xor XOR2 (N13375, N13370, N7830);
nor NOR2 (N13376, N13364, N2520);
nand NAND2 (N13377, N13368, N10243);
nor NOR4 (N13378, N13371, N8309, N407, N12496);
and AND2 (N13379, N13376, N3336);
and AND4 (N13380, N13374, N10720, N1647, N10948);
nand NAND2 (N13381, N13377, N10000);
xor XOR2 (N13382, N13365, N10139);
not NOT1 (N13383, N13382);
xor XOR2 (N13384, N13380, N10730);
nand NAND4 (N13385, N13339, N3054, N2586, N5947);
not NOT1 (N13386, N13378);
not NOT1 (N13387, N13373);
buf BUF1 (N13388, N13379);
and AND4 (N13389, N13372, N8243, N268, N8082);
or OR2 (N13390, N13386, N5440);
buf BUF1 (N13391, N13390);
xor XOR2 (N13392, N13385, N2971);
buf BUF1 (N13393, N13383);
nor NOR2 (N13394, N13384, N8112);
not NOT1 (N13395, N13389);
xor XOR2 (N13396, N13392, N5770);
xor XOR2 (N13397, N13360, N4472);
xor XOR2 (N13398, N13375, N8207);
xor XOR2 (N13399, N13393, N7391);
buf BUF1 (N13400, N13394);
nand NAND2 (N13401, N13381, N5883);
nor NOR2 (N13402, N13398, N3450);
nand NAND2 (N13403, N13391, N8521);
not NOT1 (N13404, N13396);
nor NOR2 (N13405, N13399, N3575);
or OR4 (N13406, N13400, N10170, N8579, N1835);
buf BUF1 (N13407, N13402);
or OR4 (N13408, N13407, N1054, N7236, N1455);
nand NAND3 (N13409, N13403, N5740, N8891);
nor NOR3 (N13410, N13395, N2375, N8296);
not NOT1 (N13411, N13401);
nand NAND4 (N13412, N13404, N10843, N8986, N2959);
and AND2 (N13413, N13409, N10295);
nand NAND3 (N13414, N13405, N10252, N2222);
xor XOR2 (N13415, N13408, N3868);
and AND2 (N13416, N13410, N12780);
nand NAND2 (N13417, N13414, N2544);
xor XOR2 (N13418, N13416, N6192);
buf BUF1 (N13419, N13417);
or OR3 (N13420, N13388, N12020, N11556);
or OR3 (N13421, N13406, N8121, N5895);
buf BUF1 (N13422, N13387);
not NOT1 (N13423, N13415);
xor XOR2 (N13424, N13423, N11616);
nor NOR2 (N13425, N13424, N370);
xor XOR2 (N13426, N13418, N3056);
not NOT1 (N13427, N13411);
buf BUF1 (N13428, N13413);
buf BUF1 (N13429, N13420);
nand NAND4 (N13430, N13419, N9127, N4064, N9440);
xor XOR2 (N13431, N13397, N7474);
or OR3 (N13432, N13429, N617, N10730);
nand NAND3 (N13433, N13428, N10297, N3362);
buf BUF1 (N13434, N13425);
not NOT1 (N13435, N13427);
and AND4 (N13436, N13435, N3141, N1829, N6953);
or OR4 (N13437, N13422, N7376, N2876, N8588);
and AND4 (N13438, N13431, N8204, N4836, N3926);
not NOT1 (N13439, N13434);
or OR2 (N13440, N13426, N6905);
nand NAND2 (N13441, N13412, N3024);
and AND3 (N13442, N13433, N5825, N8083);
xor XOR2 (N13443, N13421, N4396);
nand NAND4 (N13444, N13443, N6059, N8901, N8410);
and AND4 (N13445, N13438, N9061, N2688, N7197);
or OR4 (N13446, N13430, N4160, N1902, N11481);
nor NOR2 (N13447, N13440, N7495);
or OR4 (N13448, N13445, N1689, N6487, N4045);
nor NOR4 (N13449, N13439, N10153, N6420, N45);
or OR3 (N13450, N13449, N3572, N8148);
xor XOR2 (N13451, N13448, N5728);
xor XOR2 (N13452, N13441, N12693);
xor XOR2 (N13453, N13436, N5701);
and AND2 (N13454, N13453, N3743);
and AND4 (N13455, N13446, N7768, N2087, N5065);
or OR3 (N13456, N13455, N6956, N4622);
buf BUF1 (N13457, N13437);
nand NAND4 (N13458, N13432, N12465, N5869, N11119);
nor NOR2 (N13459, N13447, N5753);
xor XOR2 (N13460, N13454, N2231);
or OR4 (N13461, N13442, N3762, N4390, N8745);
and AND2 (N13462, N13444, N10776);
not NOT1 (N13463, N13462);
and AND4 (N13464, N13459, N5539, N13050, N2903);
not NOT1 (N13465, N13457);
xor XOR2 (N13466, N13451, N4286);
buf BUF1 (N13467, N13456);
not NOT1 (N13468, N13467);
buf BUF1 (N13469, N13466);
buf BUF1 (N13470, N13461);
nand NAND4 (N13471, N13458, N1610, N7504, N8959);
nor NOR2 (N13472, N13450, N9410);
nor NOR4 (N13473, N13452, N7436, N3739, N9362);
and AND2 (N13474, N13460, N2306);
not NOT1 (N13475, N13464);
buf BUF1 (N13476, N13465);
or OR4 (N13477, N13476, N13160, N8645, N10863);
not NOT1 (N13478, N13474);
and AND2 (N13479, N13463, N7233);
nand NAND3 (N13480, N13478, N8858, N12756);
xor XOR2 (N13481, N13480, N6081);
xor XOR2 (N13482, N13471, N8319);
xor XOR2 (N13483, N13469, N11261);
buf BUF1 (N13484, N13481);
or OR2 (N13485, N13468, N650);
or OR2 (N13486, N13484, N13130);
or OR4 (N13487, N13483, N3153, N9784, N2503);
xor XOR2 (N13488, N13475, N12813);
not NOT1 (N13489, N13477);
and AND4 (N13490, N13488, N10955, N3750, N12869);
and AND4 (N13491, N13479, N9325, N4464, N5087);
nor NOR3 (N13492, N13491, N705, N8458);
nor NOR4 (N13493, N13482, N9045, N2004, N10198);
nand NAND4 (N13494, N13489, N10034, N8926, N1649);
xor XOR2 (N13495, N13494, N7843);
nand NAND2 (N13496, N13490, N10509);
xor XOR2 (N13497, N13472, N6416);
buf BUF1 (N13498, N13470);
buf BUF1 (N13499, N13496);
xor XOR2 (N13500, N13493, N6530);
buf BUF1 (N13501, N13495);
not NOT1 (N13502, N13492);
xor XOR2 (N13503, N13486, N2312);
buf BUF1 (N13504, N13503);
xor XOR2 (N13505, N13473, N6569);
not NOT1 (N13506, N13500);
buf BUF1 (N13507, N13498);
and AND4 (N13508, N13497, N10950, N5546, N8447);
or OR4 (N13509, N13501, N5031, N8228, N5872);
xor XOR2 (N13510, N13499, N5839);
not NOT1 (N13511, N13510);
xor XOR2 (N13512, N13509, N7211);
or OR2 (N13513, N13506, N5405);
nor NOR2 (N13514, N13508, N13149);
not NOT1 (N13515, N13513);
nor NOR2 (N13516, N13487, N5268);
xor XOR2 (N13517, N13504, N10238);
not NOT1 (N13518, N13517);
or OR4 (N13519, N13507, N2696, N13042, N23);
nand NAND3 (N13520, N13514, N9181, N13310);
not NOT1 (N13521, N13502);
nor NOR2 (N13522, N13505, N12274);
buf BUF1 (N13523, N13516);
nand NAND4 (N13524, N13519, N9403, N10360, N1231);
nand NAND2 (N13525, N13518, N12065);
nor NOR4 (N13526, N13521, N5725, N10168, N396);
nor NOR2 (N13527, N13526, N539);
not NOT1 (N13528, N13527);
and AND3 (N13529, N13485, N12751, N5593);
and AND3 (N13530, N13515, N8847, N4856);
not NOT1 (N13531, N13530);
or OR2 (N13532, N13531, N3799);
not NOT1 (N13533, N13524);
xor XOR2 (N13534, N13523, N10750);
or OR2 (N13535, N13529, N3830);
or OR2 (N13536, N13522, N6774);
buf BUF1 (N13537, N13536);
and AND2 (N13538, N13511, N8161);
xor XOR2 (N13539, N13534, N13283);
xor XOR2 (N13540, N13525, N2832);
nor NOR4 (N13541, N13535, N9897, N1277, N12785);
xor XOR2 (N13542, N13528, N290);
xor XOR2 (N13543, N13541, N6251);
nand NAND2 (N13544, N13539, N11073);
buf BUF1 (N13545, N13533);
xor XOR2 (N13546, N13520, N483);
or OR3 (N13547, N13546, N8457, N954);
and AND4 (N13548, N13543, N6974, N2349, N8623);
nor NOR3 (N13549, N13532, N11173, N3963);
buf BUF1 (N13550, N13540);
not NOT1 (N13551, N13548);
nor NOR2 (N13552, N13512, N8528);
nor NOR3 (N13553, N13544, N1819, N4821);
buf BUF1 (N13554, N13551);
buf BUF1 (N13555, N13545);
or OR3 (N13556, N13554, N2348, N10931);
nand NAND4 (N13557, N13553, N11845, N3055, N1467);
nand NAND2 (N13558, N13555, N7484);
xor XOR2 (N13559, N13542, N5575);
not NOT1 (N13560, N13557);
and AND4 (N13561, N13560, N7329, N10711, N4365);
nand NAND4 (N13562, N13547, N8738, N2515, N12952);
not NOT1 (N13563, N13559);
not NOT1 (N13564, N13552);
or OR2 (N13565, N13563, N1948);
or OR3 (N13566, N13550, N8041, N7899);
not NOT1 (N13567, N13566);
and AND2 (N13568, N13565, N7871);
and AND3 (N13569, N13558, N12265, N8420);
xor XOR2 (N13570, N13537, N11298);
and AND4 (N13571, N13570, N10793, N8185, N12394);
nor NOR3 (N13572, N13567, N4947, N725);
xor XOR2 (N13573, N13556, N5442);
buf BUF1 (N13574, N13549);
or OR3 (N13575, N13573, N9912, N4444);
nor NOR3 (N13576, N13571, N3841, N13064);
buf BUF1 (N13577, N13538);
nor NOR4 (N13578, N13576, N5865, N12354, N9040);
nor NOR4 (N13579, N13561, N2576, N769, N13260);
and AND2 (N13580, N13572, N343);
not NOT1 (N13581, N13579);
nand NAND2 (N13582, N13575, N9769);
not NOT1 (N13583, N13578);
not NOT1 (N13584, N13574);
and AND3 (N13585, N13582, N5305, N9909);
not NOT1 (N13586, N13583);
nand NAND2 (N13587, N13568, N101);
and AND2 (N13588, N13580, N12199);
xor XOR2 (N13589, N13585, N1659);
xor XOR2 (N13590, N13587, N4166);
or OR3 (N13591, N13562, N6275, N3081);
xor XOR2 (N13592, N13581, N13027);
nand NAND2 (N13593, N13564, N8333);
and AND2 (N13594, N13589, N6772);
or OR4 (N13595, N13592, N9565, N7429, N2563);
nand NAND4 (N13596, N13586, N3293, N2942, N10018);
or OR3 (N13597, N13584, N7214, N8949);
and AND3 (N13598, N13593, N6150, N114);
nand NAND3 (N13599, N13594, N6775, N385);
nor NOR4 (N13600, N13598, N5778, N3309, N13567);
not NOT1 (N13601, N13599);
nand NAND2 (N13602, N13601, N1425);
not NOT1 (N13603, N13597);
and AND2 (N13604, N13588, N5333);
xor XOR2 (N13605, N13595, N357);
nand NAND2 (N13606, N13605, N1360);
and AND3 (N13607, N13577, N10763, N9188);
nand NAND4 (N13608, N13590, N7250, N3041, N2026);
nor NOR4 (N13609, N13591, N4119, N706, N11662);
xor XOR2 (N13610, N13607, N8188);
not NOT1 (N13611, N13569);
and AND3 (N13612, N13600, N7170, N6927);
or OR4 (N13613, N13602, N3803, N1981, N777);
nor NOR2 (N13614, N13608, N6363);
or OR3 (N13615, N13604, N2147, N12990);
nor NOR3 (N13616, N13596, N897, N4322);
nand NAND2 (N13617, N13610, N8624);
not NOT1 (N13618, N13609);
or OR2 (N13619, N13611, N2563);
not NOT1 (N13620, N13618);
and AND4 (N13621, N13620, N1122, N8989, N4353);
buf BUF1 (N13622, N13621);
or OR2 (N13623, N13619, N10944);
or OR2 (N13624, N13623, N9643);
or OR4 (N13625, N13614, N11623, N1553, N11536);
and AND2 (N13626, N13615, N12732);
not NOT1 (N13627, N13612);
or OR3 (N13628, N13613, N4123, N12100);
xor XOR2 (N13629, N13625, N11478);
nor NOR3 (N13630, N13629, N948, N6458);
nand NAND4 (N13631, N13627, N8727, N7071, N8607);
nand NAND4 (N13632, N13616, N1089, N7567, N1547);
buf BUF1 (N13633, N13606);
not NOT1 (N13634, N13622);
and AND4 (N13635, N13634, N10670, N660, N9329);
and AND3 (N13636, N13626, N7793, N4689);
buf BUF1 (N13637, N13635);
nor NOR3 (N13638, N13631, N9229, N5243);
buf BUF1 (N13639, N13632);
and AND2 (N13640, N13636, N1033);
nor NOR3 (N13641, N13617, N8035, N378);
nand NAND3 (N13642, N13603, N10395, N9155);
not NOT1 (N13643, N13641);
nor NOR4 (N13644, N13638, N10360, N2905, N4973);
nand NAND2 (N13645, N13640, N11638);
nand NAND4 (N13646, N13637, N5699, N3543, N2093);
xor XOR2 (N13647, N13643, N2596);
nor NOR2 (N13648, N13646, N2848);
buf BUF1 (N13649, N13628);
or OR3 (N13650, N13642, N8095, N12294);
nand NAND2 (N13651, N13644, N3530);
xor XOR2 (N13652, N13630, N1751);
or OR4 (N13653, N13651, N396, N7850, N1215);
and AND2 (N13654, N13647, N9560);
and AND2 (N13655, N13639, N8886);
nor NOR2 (N13656, N13645, N1629);
nor NOR3 (N13657, N13653, N4064, N3204);
nor NOR2 (N13658, N13654, N5449);
and AND3 (N13659, N13655, N9780, N6829);
nand NAND3 (N13660, N13652, N4976, N4782);
and AND4 (N13661, N13624, N1843, N6609, N8788);
not NOT1 (N13662, N13660);
xor XOR2 (N13663, N13650, N4118);
nor NOR4 (N13664, N13633, N5634, N3978, N3392);
not NOT1 (N13665, N13663);
nor NOR3 (N13666, N13661, N9881, N10613);
buf BUF1 (N13667, N13664);
nor NOR4 (N13668, N13648, N10069, N2407, N3295);
nor NOR4 (N13669, N13662, N722, N9760, N4350);
and AND4 (N13670, N13649, N3366, N8851, N4080);
and AND2 (N13671, N13665, N8172);
and AND4 (N13672, N13659, N4065, N2788, N10686);
buf BUF1 (N13673, N13656);
nand NAND2 (N13674, N13668, N5534);
and AND3 (N13675, N13671, N4434, N4146);
buf BUF1 (N13676, N13658);
nand NAND3 (N13677, N13675, N9226, N8589);
buf BUF1 (N13678, N13677);
or OR4 (N13679, N13670, N4271, N2542, N2940);
and AND3 (N13680, N13673, N7407, N10063);
not NOT1 (N13681, N13657);
nor NOR3 (N13682, N13669, N10799, N11097);
not NOT1 (N13683, N13667);
nand NAND4 (N13684, N13672, N8558, N4937, N2710);
buf BUF1 (N13685, N13681);
nor NOR3 (N13686, N13674, N3042, N13639);
or OR4 (N13687, N13666, N10301, N4184, N3455);
buf BUF1 (N13688, N13687);
and AND3 (N13689, N13682, N7605, N122);
and AND4 (N13690, N13689, N9323, N4627, N1793);
or OR3 (N13691, N13678, N5086, N5580);
nor NOR2 (N13692, N13683, N12937);
xor XOR2 (N13693, N13684, N421);
buf BUF1 (N13694, N13688);
and AND2 (N13695, N13692, N8007);
and AND3 (N13696, N13693, N10717, N8357);
buf BUF1 (N13697, N13690);
nand NAND4 (N13698, N13695, N6922, N4274, N6029);
not NOT1 (N13699, N13680);
nor NOR4 (N13700, N13696, N1339, N11708, N8465);
xor XOR2 (N13701, N13685, N11875);
nand NAND4 (N13702, N13698, N7800, N10013, N12886);
xor XOR2 (N13703, N13694, N5310);
nor NOR2 (N13704, N13686, N11034);
and AND2 (N13705, N13702, N9202);
xor XOR2 (N13706, N13700, N1504);
buf BUF1 (N13707, N13697);
xor XOR2 (N13708, N13679, N10473);
and AND2 (N13709, N13676, N2709);
nor NOR2 (N13710, N13699, N2003);
not NOT1 (N13711, N13710);
nand NAND3 (N13712, N13707, N5932, N8657);
nor NOR3 (N13713, N13711, N5176, N8402);
and AND4 (N13714, N13713, N11071, N684, N3054);
xor XOR2 (N13715, N13701, N6119);
nand NAND3 (N13716, N13691, N5660, N6978);
xor XOR2 (N13717, N13716, N10114);
or OR4 (N13718, N13706, N8261, N3716, N2019);
or OR3 (N13719, N13715, N6958, N2871);
nand NAND4 (N13720, N13719, N11516, N9827, N6087);
xor XOR2 (N13721, N13709, N5950);
nand NAND2 (N13722, N13704, N6023);
and AND2 (N13723, N13720, N2927);
and AND2 (N13724, N13718, N2746);
nor NOR4 (N13725, N13717, N7800, N11803, N666);
or OR4 (N13726, N13703, N2142, N12221, N13491);
xor XOR2 (N13727, N13712, N9898);
nand NAND4 (N13728, N13721, N10619, N12641, N13148);
xor XOR2 (N13729, N13722, N2746);
nand NAND4 (N13730, N13708, N8609, N8546, N8449);
and AND2 (N13731, N13705, N6791);
not NOT1 (N13732, N13731);
nor NOR2 (N13733, N13732, N150);
not NOT1 (N13734, N13727);
not NOT1 (N13735, N13724);
not NOT1 (N13736, N13730);
nand NAND3 (N13737, N13729, N1823, N1542);
xor XOR2 (N13738, N13728, N898);
nor NOR2 (N13739, N13736, N4548);
buf BUF1 (N13740, N13737);
or OR3 (N13741, N13725, N775, N4809);
nor NOR2 (N13742, N13739, N13715);
buf BUF1 (N13743, N13741);
nand NAND2 (N13744, N13742, N7466);
xor XOR2 (N13745, N13734, N1871);
nand NAND3 (N13746, N13738, N10751, N7718);
not NOT1 (N13747, N13726);
and AND4 (N13748, N13745, N6608, N7336, N98);
not NOT1 (N13749, N13743);
xor XOR2 (N13750, N13746, N8241);
xor XOR2 (N13751, N13749, N10671);
nand NAND2 (N13752, N13750, N7482);
buf BUF1 (N13753, N13752);
or OR3 (N13754, N13723, N12955, N3248);
xor XOR2 (N13755, N13744, N740);
nand NAND3 (N13756, N13751, N13627, N3226);
xor XOR2 (N13757, N13740, N5273);
or OR3 (N13758, N13754, N12930, N12685);
buf BUF1 (N13759, N13747);
and AND4 (N13760, N13755, N13530, N4142, N2476);
nor NOR2 (N13761, N13757, N4137);
or OR4 (N13762, N13735, N6792, N81, N10155);
not NOT1 (N13763, N13714);
nand NAND4 (N13764, N13748, N2373, N11480, N3946);
not NOT1 (N13765, N13753);
xor XOR2 (N13766, N13758, N8743);
nor NOR2 (N13767, N13760, N4931);
not NOT1 (N13768, N13756);
buf BUF1 (N13769, N13766);
xor XOR2 (N13770, N13763, N12902);
not NOT1 (N13771, N13733);
buf BUF1 (N13772, N13770);
xor XOR2 (N13773, N13761, N9360);
or OR2 (N13774, N13759, N4901);
nand NAND3 (N13775, N13772, N12725, N11376);
and AND2 (N13776, N13765, N57);
buf BUF1 (N13777, N13773);
nor NOR3 (N13778, N13768, N11601, N1020);
not NOT1 (N13779, N13774);
nand NAND4 (N13780, N13775, N11760, N701, N4185);
nor NOR3 (N13781, N13769, N4696, N13242);
nor NOR3 (N13782, N13778, N11426, N680);
or OR3 (N13783, N13782, N8908, N11883);
or OR4 (N13784, N13783, N4546, N11172, N8071);
and AND3 (N13785, N13767, N5575, N5211);
xor XOR2 (N13786, N13771, N13467);
or OR4 (N13787, N13785, N9324, N5994, N3202);
and AND3 (N13788, N13787, N7848, N10822);
nand NAND3 (N13789, N13780, N7179, N9566);
and AND3 (N13790, N13784, N3052, N2276);
buf BUF1 (N13791, N13786);
not NOT1 (N13792, N13762);
nand NAND3 (N13793, N13779, N2140, N9155);
xor XOR2 (N13794, N13791, N413);
nor NOR3 (N13795, N13792, N6367, N528);
not NOT1 (N13796, N13795);
nand NAND4 (N13797, N13781, N12976, N12087, N962);
nor NOR2 (N13798, N13777, N288);
buf BUF1 (N13799, N13790);
not NOT1 (N13800, N13788);
and AND3 (N13801, N13764, N8737, N1895);
or OR2 (N13802, N13796, N12035);
and AND3 (N13803, N13797, N4500, N10458);
nand NAND2 (N13804, N13789, N4062);
buf BUF1 (N13805, N13803);
nor NOR3 (N13806, N13804, N3178, N13023);
nor NOR2 (N13807, N13799, N2317);
nor NOR3 (N13808, N13807, N11506, N2259);
buf BUF1 (N13809, N13808);
nor NOR4 (N13810, N13776, N11478, N3848, N12529);
not NOT1 (N13811, N13793);
nor NOR4 (N13812, N13800, N9952, N6492, N1416);
xor XOR2 (N13813, N13798, N12483);
and AND3 (N13814, N13809, N5250, N1690);
nor NOR3 (N13815, N13801, N1536, N4985);
nor NOR3 (N13816, N13802, N2896, N10064);
and AND3 (N13817, N13816, N4130, N9898);
buf BUF1 (N13818, N13811);
and AND4 (N13819, N13794, N9929, N10332, N833);
buf BUF1 (N13820, N13819);
nor NOR4 (N13821, N13817, N11570, N5016, N4530);
nand NAND2 (N13822, N13818, N11302);
nand NAND3 (N13823, N13812, N13469, N13648);
xor XOR2 (N13824, N13806, N7532);
or OR4 (N13825, N13824, N5830, N7785, N4741);
or OR3 (N13826, N13815, N9035, N8028);
not NOT1 (N13827, N13822);
nor NOR3 (N13828, N13814, N9737, N10917);
not NOT1 (N13829, N13825);
buf BUF1 (N13830, N13820);
or OR4 (N13831, N13813, N11294, N7165, N4904);
not NOT1 (N13832, N13829);
buf BUF1 (N13833, N13826);
or OR4 (N13834, N13833, N10415, N2703, N10056);
buf BUF1 (N13835, N13832);
xor XOR2 (N13836, N13835, N2528);
not NOT1 (N13837, N13810);
and AND2 (N13838, N13827, N1871);
and AND3 (N13839, N13805, N3638, N11153);
xor XOR2 (N13840, N13823, N3454);
nand NAND3 (N13841, N13831, N178, N10432);
buf BUF1 (N13842, N13839);
and AND4 (N13843, N13821, N1670, N2394, N57);
or OR4 (N13844, N13834, N4632, N1184, N5463);
nor NOR4 (N13845, N13837, N1844, N220, N4255);
not NOT1 (N13846, N13840);
nor NOR2 (N13847, N13845, N6739);
not NOT1 (N13848, N13843);
and AND4 (N13849, N13830, N11045, N7973, N3998);
nand NAND4 (N13850, N13846, N11774, N7159, N13156);
nor NOR2 (N13851, N13828, N9393);
and AND2 (N13852, N13841, N13851);
or OR4 (N13853, N13378, N8798, N5284, N10824);
nor NOR4 (N13854, N13844, N10607, N672, N13651);
or OR3 (N13855, N13852, N3573, N3861);
nand NAND4 (N13856, N13838, N12094, N12738, N1740);
xor XOR2 (N13857, N13847, N11416);
nand NAND4 (N13858, N13848, N6279, N5339, N5614);
buf BUF1 (N13859, N13855);
buf BUF1 (N13860, N13842);
nand NAND2 (N13861, N13853, N6557);
not NOT1 (N13862, N13849);
buf BUF1 (N13863, N13850);
nand NAND4 (N13864, N13836, N6713, N11321, N7597);
xor XOR2 (N13865, N13859, N8663);
buf BUF1 (N13866, N13862);
not NOT1 (N13867, N13858);
nor NOR4 (N13868, N13864, N7903, N11444, N1352);
nand NAND4 (N13869, N13854, N12927, N12883, N5350);
nand NAND3 (N13870, N13865, N12023, N4082);
nand NAND4 (N13871, N13870, N2646, N4676, N4603);
nor NOR3 (N13872, N13861, N9139, N5399);
not NOT1 (N13873, N13857);
nand NAND2 (N13874, N13868, N709);
and AND4 (N13875, N13863, N4061, N5185, N2186);
not NOT1 (N13876, N13866);
or OR4 (N13877, N13872, N4834, N12411, N4);
or OR3 (N13878, N13874, N445, N8649);
buf BUF1 (N13879, N13875);
buf BUF1 (N13880, N13867);
or OR4 (N13881, N13871, N9440, N1142, N902);
and AND4 (N13882, N13877, N6906, N11765, N4563);
nor NOR3 (N13883, N13873, N5186, N1059);
and AND4 (N13884, N13879, N4331, N12371, N4956);
and AND2 (N13885, N13860, N6060);
nor NOR3 (N13886, N13884, N3067, N1162);
not NOT1 (N13887, N13883);
or OR2 (N13888, N13887, N1470);
xor XOR2 (N13889, N13878, N10617);
buf BUF1 (N13890, N13889);
not NOT1 (N13891, N13876);
buf BUF1 (N13892, N13882);
buf BUF1 (N13893, N13869);
xor XOR2 (N13894, N13888, N1293);
or OR2 (N13895, N13881, N1322);
nand NAND2 (N13896, N13895, N5111);
or OR4 (N13897, N13856, N4048, N8736, N4676);
buf BUF1 (N13898, N13890);
nand NAND4 (N13899, N13880, N6731, N1580, N71);
or OR2 (N13900, N13892, N4251);
not NOT1 (N13901, N13900);
or OR3 (N13902, N13898, N13232, N5044);
or OR3 (N13903, N13886, N3391, N10103);
and AND3 (N13904, N13893, N3977, N2222);
xor XOR2 (N13905, N13902, N9932);
buf BUF1 (N13906, N13894);
nor NOR4 (N13907, N13897, N6256, N4630, N10406);
and AND3 (N13908, N13907, N11072, N13558);
xor XOR2 (N13909, N13908, N10795);
buf BUF1 (N13910, N13903);
and AND4 (N13911, N13906, N9447, N11305, N3622);
nand NAND3 (N13912, N13899, N11868, N2373);
buf BUF1 (N13913, N13896);
buf BUF1 (N13914, N13910);
not NOT1 (N13915, N13904);
buf BUF1 (N13916, N13915);
not NOT1 (N13917, N13891);
buf BUF1 (N13918, N13913);
xor XOR2 (N13919, N13916, N12444);
buf BUF1 (N13920, N13914);
nand NAND3 (N13921, N13919, N3422, N12681);
not NOT1 (N13922, N13901);
nand NAND4 (N13923, N13905, N281, N932, N11539);
buf BUF1 (N13924, N13911);
nor NOR4 (N13925, N13917, N1744, N9390, N2379);
nand NAND2 (N13926, N13922, N9643);
not NOT1 (N13927, N13926);
and AND4 (N13928, N13925, N11520, N10310, N2477);
or OR2 (N13929, N13918, N10553);
or OR2 (N13930, N13920, N13474);
or OR4 (N13931, N13885, N13479, N13203, N12916);
and AND2 (N13932, N13924, N7825);
buf BUF1 (N13933, N13927);
xor XOR2 (N13934, N13930, N6450);
and AND3 (N13935, N13933, N3569, N870);
nand NAND3 (N13936, N13934, N9801, N1902);
xor XOR2 (N13937, N13923, N12773);
nor NOR4 (N13938, N13929, N9407, N2918, N4665);
xor XOR2 (N13939, N13937, N4150);
or OR4 (N13940, N13936, N4407, N6914, N8503);
xor XOR2 (N13941, N13935, N872);
xor XOR2 (N13942, N13928, N9825);
xor XOR2 (N13943, N13931, N2083);
not NOT1 (N13944, N13938);
xor XOR2 (N13945, N13921, N6890);
not NOT1 (N13946, N13943);
xor XOR2 (N13947, N13942, N7067);
xor XOR2 (N13948, N13939, N8991);
nand NAND3 (N13949, N13944, N5667, N12044);
nand NAND4 (N13950, N13940, N13651, N1184, N10029);
buf BUF1 (N13951, N13946);
nor NOR3 (N13952, N13909, N10836, N2061);
nor NOR4 (N13953, N13941, N9860, N11083, N12257);
nand NAND2 (N13954, N13932, N13154);
buf BUF1 (N13955, N13948);
and AND4 (N13956, N13953, N5319, N4044, N625);
buf BUF1 (N13957, N13949);
not NOT1 (N13958, N13951);
nor NOR2 (N13959, N13947, N9597);
not NOT1 (N13960, N13958);
not NOT1 (N13961, N13912);
buf BUF1 (N13962, N13959);
buf BUF1 (N13963, N13952);
buf BUF1 (N13964, N13945);
not NOT1 (N13965, N13956);
and AND2 (N13966, N13965, N5503);
xor XOR2 (N13967, N13964, N5518);
nor NOR2 (N13968, N13954, N4148);
or OR3 (N13969, N13966, N10563, N12755);
xor XOR2 (N13970, N13960, N9289);
and AND2 (N13971, N13961, N12045);
and AND3 (N13972, N13967, N12987, N1445);
buf BUF1 (N13973, N13962);
not NOT1 (N13974, N13950);
nor NOR3 (N13975, N13969, N404, N3280);
and AND4 (N13976, N13971, N4807, N13591, N12842);
buf BUF1 (N13977, N13970);
nor NOR3 (N13978, N13974, N11887, N3178);
or OR4 (N13979, N13977, N79, N10927, N11298);
buf BUF1 (N13980, N13972);
buf BUF1 (N13981, N13973);
buf BUF1 (N13982, N13975);
nor NOR3 (N13983, N13955, N8025, N12695);
nor NOR4 (N13984, N13957, N12715, N5010, N2194);
nand NAND3 (N13985, N13976, N10387, N176);
and AND4 (N13986, N13984, N4103, N13705, N5109);
or OR2 (N13987, N13985, N5244);
not NOT1 (N13988, N13978);
and AND2 (N13989, N13968, N13415);
nor NOR3 (N13990, N13989, N5937, N3744);
xor XOR2 (N13991, N13979, N12834);
buf BUF1 (N13992, N13987);
nor NOR4 (N13993, N13980, N2121, N5224, N7133);
nand NAND2 (N13994, N13983, N7563);
xor XOR2 (N13995, N13988, N12190);
nand NAND4 (N13996, N13992, N7933, N13876, N4025);
xor XOR2 (N13997, N13991, N5846);
or OR2 (N13998, N13995, N4651);
or OR3 (N13999, N13981, N10522, N11040);
nor NOR2 (N14000, N13990, N13785);
nand NAND3 (N14001, N13993, N9907, N6615);
and AND3 (N14002, N13994, N5877, N923);
nand NAND4 (N14003, N14001, N10711, N3124, N7719);
nor NOR2 (N14004, N14000, N2328);
or OR2 (N14005, N13986, N1358);
nand NAND3 (N14006, N13963, N9637, N7292);
nand NAND2 (N14007, N13998, N2563);
not NOT1 (N14008, N13982);
and AND4 (N14009, N14002, N7065, N11232, N1633);
or OR2 (N14010, N14003, N9886);
buf BUF1 (N14011, N14006);
xor XOR2 (N14012, N14010, N5302);
or OR3 (N14013, N13996, N7671, N8606);
nand NAND4 (N14014, N14012, N2236, N124, N6112);
not NOT1 (N14015, N14008);
and AND2 (N14016, N14007, N3865);
not NOT1 (N14017, N13997);
nor NOR3 (N14018, N14017, N6408, N13533);
xor XOR2 (N14019, N14013, N812);
xor XOR2 (N14020, N14015, N3956);
or OR4 (N14021, N14018, N10040, N2841, N10436);
xor XOR2 (N14022, N14020, N350);
buf BUF1 (N14023, N14005);
nor NOR3 (N14024, N14021, N3597, N7991);
nand NAND4 (N14025, N14022, N12942, N10610, N13492);
nand NAND2 (N14026, N14004, N13754);
and AND2 (N14027, N14011, N11209);
nand NAND3 (N14028, N14009, N6605, N9385);
and AND3 (N14029, N14024, N1539, N4205);
xor XOR2 (N14030, N14029, N6549);
or OR4 (N14031, N14026, N12948, N13397, N3214);
or OR2 (N14032, N14023, N12542);
buf BUF1 (N14033, N14019);
nor NOR2 (N14034, N14033, N2408);
buf BUF1 (N14035, N13999);
or OR2 (N14036, N14028, N2493);
buf BUF1 (N14037, N14036);
buf BUF1 (N14038, N14035);
buf BUF1 (N14039, N14016);
buf BUF1 (N14040, N14039);
and AND2 (N14041, N14014, N3600);
and AND3 (N14042, N14041, N774, N6559);
and AND2 (N14043, N14030, N3414);
and AND2 (N14044, N14040, N10238);
nand NAND2 (N14045, N14042, N5674);
not NOT1 (N14046, N14045);
xor XOR2 (N14047, N14046, N10798);
not NOT1 (N14048, N14043);
and AND4 (N14049, N14047, N12885, N2843, N5013);
or OR3 (N14050, N14049, N6513, N731);
nor NOR2 (N14051, N14038, N2598);
and AND4 (N14052, N14048, N10665, N5804, N9253);
not NOT1 (N14053, N14027);
nor NOR2 (N14054, N14034, N7506);
and AND2 (N14055, N14053, N7377);
buf BUF1 (N14056, N14032);
and AND3 (N14057, N14050, N7178, N13631);
nand NAND3 (N14058, N14051, N9149, N7086);
nor NOR3 (N14059, N14052, N854, N974);
buf BUF1 (N14060, N14058);
and AND2 (N14061, N14055, N8166);
and AND2 (N14062, N14037, N12637);
buf BUF1 (N14063, N14025);
xor XOR2 (N14064, N14031, N12819);
and AND4 (N14065, N14062, N5995, N13194, N5123);
or OR2 (N14066, N14060, N563);
and AND4 (N14067, N14064, N7159, N13740, N2902);
xor XOR2 (N14068, N14066, N2913);
xor XOR2 (N14069, N14065, N3511);
or OR3 (N14070, N14063, N4627, N1085);
and AND2 (N14071, N14061, N5449);
nand NAND3 (N14072, N14069, N7219, N5492);
nand NAND3 (N14073, N14057, N2024, N11948);
buf BUF1 (N14074, N14056);
and AND4 (N14075, N14071, N11219, N3663, N10032);
xor XOR2 (N14076, N14068, N7816);
nand NAND4 (N14077, N14075, N6013, N1004, N3377);
nor NOR2 (N14078, N14059, N10078);
nand NAND4 (N14079, N14078, N1199, N1546, N6779);
xor XOR2 (N14080, N14067, N1772);
buf BUF1 (N14081, N14072);
and AND4 (N14082, N14077, N11808, N6772, N6518);
and AND2 (N14083, N14054, N9250);
xor XOR2 (N14084, N14082, N10944);
not NOT1 (N14085, N14076);
buf BUF1 (N14086, N14084);
xor XOR2 (N14087, N14044, N12353);
xor XOR2 (N14088, N14070, N3377);
nor NOR4 (N14089, N14086, N5583, N4249, N5628);
or OR4 (N14090, N14074, N13252, N10880, N10633);
nor NOR3 (N14091, N14085, N6258, N10912);
and AND4 (N14092, N14089, N8766, N2825, N1637);
and AND2 (N14093, N14091, N12129);
nor NOR2 (N14094, N14088, N4502);
nand NAND4 (N14095, N14087, N11085, N402, N6540);
and AND3 (N14096, N14093, N13304, N1126);
or OR4 (N14097, N14094, N12458, N1054, N3568);
not NOT1 (N14098, N14083);
buf BUF1 (N14099, N14080);
and AND3 (N14100, N14099, N2896, N10663);
not NOT1 (N14101, N14073);
buf BUF1 (N14102, N14079);
nand NAND4 (N14103, N14097, N1200, N8919, N3919);
or OR2 (N14104, N14090, N13365);
buf BUF1 (N14105, N14103);
or OR4 (N14106, N14102, N4014, N8104, N691);
not NOT1 (N14107, N14100);
nand NAND4 (N14108, N14107, N6303, N9840, N6734);
and AND2 (N14109, N14092, N12507);
or OR2 (N14110, N14095, N10933);
buf BUF1 (N14111, N14105);
buf BUF1 (N14112, N14096);
nor NOR2 (N14113, N14106, N4293);
nand NAND3 (N14114, N14108, N5406, N13614);
buf BUF1 (N14115, N14111);
xor XOR2 (N14116, N14113, N2852);
nor NOR4 (N14117, N14115, N11102, N4155, N12377);
buf BUF1 (N14118, N14104);
or OR4 (N14119, N14114, N10186, N3048, N11780);
or OR4 (N14120, N14109, N7780, N12371, N10390);
and AND4 (N14121, N14117, N9765, N7630, N680);
buf BUF1 (N14122, N14120);
nor NOR2 (N14123, N14119, N464);
or OR4 (N14124, N14122, N7667, N7464, N4824);
or OR2 (N14125, N14101, N5507);
or OR3 (N14126, N14123, N11578, N8589);
nand NAND3 (N14127, N14121, N1602, N9090);
or OR3 (N14128, N14126, N7072, N4641);
nand NAND4 (N14129, N14125, N9012, N3787, N13584);
or OR2 (N14130, N14110, N9430);
nand NAND3 (N14131, N14128, N6845, N7969);
and AND3 (N14132, N14098, N12305, N7721);
buf BUF1 (N14133, N14130);
nor NOR4 (N14134, N14116, N6122, N7466, N12261);
xor XOR2 (N14135, N14127, N11709);
and AND2 (N14136, N14131, N6484);
or OR2 (N14137, N14129, N3312);
and AND4 (N14138, N14112, N1269, N9515, N3558);
nand NAND2 (N14139, N14138, N2923);
xor XOR2 (N14140, N14081, N6047);
not NOT1 (N14141, N14139);
or OR2 (N14142, N14135, N4649);
or OR4 (N14143, N14142, N401, N3476, N14007);
and AND2 (N14144, N14141, N5529);
nand NAND2 (N14145, N14136, N6585);
not NOT1 (N14146, N14145);
nor NOR2 (N14147, N14137, N2164);
nor NOR4 (N14148, N14143, N680, N7622, N7585);
nand NAND4 (N14149, N14133, N12918, N6193, N1392);
or OR4 (N14150, N14147, N2652, N5125, N10662);
buf BUF1 (N14151, N14118);
not NOT1 (N14152, N14148);
nor NOR2 (N14153, N14124, N12945);
nor NOR2 (N14154, N14150, N6285);
xor XOR2 (N14155, N14153, N518);
not NOT1 (N14156, N14140);
or OR2 (N14157, N14155, N5199);
buf BUF1 (N14158, N14146);
nor NOR3 (N14159, N14151, N5872, N11750);
xor XOR2 (N14160, N14132, N1032);
buf BUF1 (N14161, N14144);
or OR2 (N14162, N14152, N6280);
or OR2 (N14163, N14154, N2745);
and AND4 (N14164, N14156, N11597, N13975, N7449);
xor XOR2 (N14165, N14162, N12255);
xor XOR2 (N14166, N14134, N10416);
not NOT1 (N14167, N14149);
or OR4 (N14168, N14159, N2198, N14046, N2817);
nand NAND2 (N14169, N14161, N4852);
and AND3 (N14170, N14167, N11599, N10139);
and AND2 (N14171, N14164, N1250);
or OR3 (N14172, N14168, N7098, N6907);
or OR2 (N14173, N14171, N13024);
not NOT1 (N14174, N14165);
nor NOR3 (N14175, N14158, N12027, N5493);
buf BUF1 (N14176, N14172);
xor XOR2 (N14177, N14160, N630);
xor XOR2 (N14178, N14170, N11310);
not NOT1 (N14179, N14178);
nand NAND4 (N14180, N14174, N8282, N3879, N3254);
xor XOR2 (N14181, N14177, N8749);
and AND2 (N14182, N14181, N11608);
nor NOR2 (N14183, N14166, N4889);
nor NOR4 (N14184, N14176, N14064, N11496, N1234);
nand NAND3 (N14185, N14163, N13709, N10117);
buf BUF1 (N14186, N14169);
xor XOR2 (N14187, N14183, N8796);
nand NAND3 (N14188, N14175, N1509, N9305);
and AND3 (N14189, N14187, N8501, N2473);
and AND4 (N14190, N14182, N10185, N3168, N10751);
nand NAND2 (N14191, N14185, N11391);
xor XOR2 (N14192, N14190, N6218);
not NOT1 (N14193, N14173);
and AND4 (N14194, N14192, N12569, N931, N12552);
nor NOR4 (N14195, N14188, N12875, N7240, N7984);
and AND2 (N14196, N14194, N817);
buf BUF1 (N14197, N14180);
or OR2 (N14198, N14184, N9541);
not NOT1 (N14199, N14197);
or OR3 (N14200, N14199, N6760, N3210);
and AND2 (N14201, N14189, N765);
nand NAND4 (N14202, N14200, N8194, N2384, N9290);
not NOT1 (N14203, N14186);
nor NOR4 (N14204, N14198, N2340, N5892, N1287);
not NOT1 (N14205, N14179);
nor NOR3 (N14206, N14203, N9621, N13041);
buf BUF1 (N14207, N14204);
nand NAND4 (N14208, N14202, N3304, N13967, N13497);
nor NOR2 (N14209, N14196, N11699);
not NOT1 (N14210, N14206);
or OR3 (N14211, N14207, N4067, N13717);
buf BUF1 (N14212, N14208);
nor NOR3 (N14213, N14157, N573, N12943);
buf BUF1 (N14214, N14205);
nand NAND3 (N14215, N14210, N11011, N9633);
buf BUF1 (N14216, N14214);
or OR3 (N14217, N14212, N5957, N4876);
nor NOR2 (N14218, N14215, N4493);
not NOT1 (N14219, N14201);
and AND2 (N14220, N14191, N11800);
xor XOR2 (N14221, N14195, N11125);
and AND3 (N14222, N14221, N11721, N1544);
nor NOR3 (N14223, N14222, N10553, N6171);
buf BUF1 (N14224, N14211);
buf BUF1 (N14225, N14193);
xor XOR2 (N14226, N14218, N13780);
not NOT1 (N14227, N14220);
nor NOR4 (N14228, N14226, N13324, N7999, N12938);
or OR2 (N14229, N14224, N5332);
or OR2 (N14230, N14229, N13913);
or OR2 (N14231, N14213, N93);
and AND2 (N14232, N14216, N13105);
buf BUF1 (N14233, N14217);
or OR2 (N14234, N14225, N13199);
and AND3 (N14235, N14232, N11450, N6606);
or OR4 (N14236, N14230, N11727, N11394, N12753);
or OR3 (N14237, N14236, N4244, N903);
and AND4 (N14238, N14235, N11627, N12408, N4632);
or OR3 (N14239, N14234, N174, N13493);
xor XOR2 (N14240, N14231, N7473);
or OR3 (N14241, N14228, N2594, N14188);
xor XOR2 (N14242, N14238, N6923);
buf BUF1 (N14243, N14219);
or OR3 (N14244, N14237, N14111, N9922);
nor NOR4 (N14245, N14244, N12267, N5963, N5938);
nor NOR2 (N14246, N14209, N931);
and AND3 (N14247, N14233, N2891, N11905);
or OR3 (N14248, N14243, N9255, N9014);
and AND3 (N14249, N14242, N10492, N5136);
xor XOR2 (N14250, N14227, N8501);
xor XOR2 (N14251, N14239, N7751);
not NOT1 (N14252, N14247);
and AND2 (N14253, N14245, N1483);
nor NOR2 (N14254, N14250, N3153);
nand NAND3 (N14255, N14246, N3039, N9035);
xor XOR2 (N14256, N14241, N3681);
buf BUF1 (N14257, N14255);
nor NOR3 (N14258, N14240, N6150, N1737);
nor NOR4 (N14259, N14254, N403, N14250, N9955);
nor NOR4 (N14260, N14253, N159, N1606, N6907);
xor XOR2 (N14261, N14251, N2167);
not NOT1 (N14262, N14252);
nor NOR3 (N14263, N14261, N6650, N9340);
or OR3 (N14264, N14259, N10713, N3746);
or OR2 (N14265, N14262, N11951);
or OR4 (N14266, N14258, N3557, N7598, N3276);
or OR4 (N14267, N14256, N4104, N2849, N1971);
not NOT1 (N14268, N14223);
nor NOR2 (N14269, N14267, N2517);
buf BUF1 (N14270, N14266);
nand NAND3 (N14271, N14257, N1715, N5449);
xor XOR2 (N14272, N14265, N171);
buf BUF1 (N14273, N14249);
or OR4 (N14274, N14269, N12840, N7712, N1000);
buf BUF1 (N14275, N14260);
not NOT1 (N14276, N14248);
and AND4 (N14277, N14276, N11016, N3722, N3048);
or OR4 (N14278, N14263, N5511, N7914, N7958);
nand NAND3 (N14279, N14272, N4452, N10774);
nand NAND2 (N14280, N14264, N11621);
xor XOR2 (N14281, N14271, N11850);
xor XOR2 (N14282, N14281, N8101);
nand NAND2 (N14283, N14279, N13637);
or OR4 (N14284, N14277, N4208, N1987, N11922);
buf BUF1 (N14285, N14274);
or OR4 (N14286, N14273, N5938, N2224, N3156);
or OR3 (N14287, N14286, N4559, N13818);
nor NOR2 (N14288, N14283, N8580);
and AND3 (N14289, N14288, N3508, N407);
and AND3 (N14290, N14287, N1130, N7930);
and AND2 (N14291, N14280, N11216);
nand NAND4 (N14292, N14290, N2878, N6852, N4143);
buf BUF1 (N14293, N14284);
and AND3 (N14294, N14291, N12999, N11645);
nor NOR2 (N14295, N14289, N2895);
nand NAND3 (N14296, N14293, N12054, N4637);
not NOT1 (N14297, N14282);
buf BUF1 (N14298, N14296);
buf BUF1 (N14299, N14270);
and AND2 (N14300, N14285, N9941);
not NOT1 (N14301, N14294);
xor XOR2 (N14302, N14268, N13818);
not NOT1 (N14303, N14295);
or OR2 (N14304, N14302, N10217);
buf BUF1 (N14305, N14300);
buf BUF1 (N14306, N14299);
not NOT1 (N14307, N14298);
not NOT1 (N14308, N14292);
and AND4 (N14309, N14275, N799, N3259, N10549);
nand NAND3 (N14310, N14297, N11731, N2646);
buf BUF1 (N14311, N14301);
or OR4 (N14312, N14303, N438, N8282, N8555);
and AND2 (N14313, N14304, N11409);
xor XOR2 (N14314, N14309, N7959);
nand NAND3 (N14315, N14311, N13775, N12589);
nand NAND3 (N14316, N14314, N3935, N13760);
xor XOR2 (N14317, N14305, N4496);
and AND4 (N14318, N14313, N6403, N9393, N11392);
buf BUF1 (N14319, N14315);
nand NAND3 (N14320, N14306, N9493, N5218);
or OR3 (N14321, N14317, N3715, N13765);
and AND4 (N14322, N14278, N13538, N162, N9448);
buf BUF1 (N14323, N14312);
or OR3 (N14324, N14321, N14201, N11124);
nor NOR4 (N14325, N14310, N11136, N3998, N6975);
nand NAND3 (N14326, N14323, N5997, N3132);
buf BUF1 (N14327, N14319);
buf BUF1 (N14328, N14308);
buf BUF1 (N14329, N14324);
nor NOR4 (N14330, N14326, N13915, N12310, N8013);
or OR3 (N14331, N14325, N763, N2208);
and AND2 (N14332, N14320, N6704);
nand NAND4 (N14333, N14328, N5503, N8176, N13247);
nor NOR4 (N14334, N14327, N10048, N13646, N14087);
and AND3 (N14335, N14316, N6045, N6898);
nand NAND4 (N14336, N14307, N10714, N10457, N3909);
xor XOR2 (N14337, N14333, N5693);
buf BUF1 (N14338, N14332);
and AND2 (N14339, N14336, N5984);
or OR3 (N14340, N14338, N11680, N11163);
and AND4 (N14341, N14335, N11101, N2933, N10690);
and AND3 (N14342, N14322, N12059, N10294);
and AND4 (N14343, N14337, N13446, N12512, N1563);
and AND3 (N14344, N14339, N5164, N6287);
not NOT1 (N14345, N14329);
nor NOR4 (N14346, N14334, N2868, N12432, N8023);
buf BUF1 (N14347, N14342);
buf BUF1 (N14348, N14344);
xor XOR2 (N14349, N14340, N1865);
or OR4 (N14350, N14343, N8768, N634, N4585);
and AND4 (N14351, N14348, N13738, N11178, N6984);
xor XOR2 (N14352, N14349, N814);
not NOT1 (N14353, N14345);
not NOT1 (N14354, N14346);
or OR3 (N14355, N14341, N10824, N87);
not NOT1 (N14356, N14355);
or OR4 (N14357, N14356, N506, N9918, N3607);
buf BUF1 (N14358, N14347);
buf BUF1 (N14359, N14350);
xor XOR2 (N14360, N14351, N13473);
buf BUF1 (N14361, N14357);
not NOT1 (N14362, N14359);
nand NAND3 (N14363, N14354, N2761, N6117);
buf BUF1 (N14364, N14360);
nand NAND2 (N14365, N14318, N11592);
and AND4 (N14366, N14365, N10179, N3667, N2283);
or OR2 (N14367, N14366, N12353);
buf BUF1 (N14368, N14353);
xor XOR2 (N14369, N14361, N8757);
xor XOR2 (N14370, N14330, N3194);
and AND4 (N14371, N14358, N4280, N1015, N9143);
and AND3 (N14372, N14364, N4586, N12000);
nand NAND2 (N14373, N14367, N75);
nand NAND3 (N14374, N14370, N9624, N3906);
not NOT1 (N14375, N14369);
nor NOR2 (N14376, N14371, N734);
and AND2 (N14377, N14352, N1906);
or OR4 (N14378, N14363, N3165, N3741, N5249);
xor XOR2 (N14379, N14374, N5030);
nand NAND2 (N14380, N14368, N13885);
xor XOR2 (N14381, N14380, N1896);
or OR4 (N14382, N14377, N3295, N9716, N2770);
or OR3 (N14383, N14331, N2445, N6263);
and AND2 (N14384, N14362, N13958);
nand NAND2 (N14385, N14382, N7118);
and AND3 (N14386, N14381, N11433, N1380);
not NOT1 (N14387, N14386);
not NOT1 (N14388, N14375);
xor XOR2 (N14389, N14384, N4445);
buf BUF1 (N14390, N14378);
or OR2 (N14391, N14388, N12866);
nor NOR2 (N14392, N14387, N4682);
and AND4 (N14393, N14379, N5860, N12261, N7055);
or OR2 (N14394, N14373, N14200);
and AND3 (N14395, N14393, N13873, N6205);
buf BUF1 (N14396, N14376);
not NOT1 (N14397, N14395);
nand NAND3 (N14398, N14397, N11195, N13663);
and AND3 (N14399, N14396, N892, N4088);
and AND3 (N14400, N14392, N4301, N1001);
and AND2 (N14401, N14390, N6329);
not NOT1 (N14402, N14372);
or OR2 (N14403, N14383, N4009);
not NOT1 (N14404, N14398);
not NOT1 (N14405, N14399);
nand NAND3 (N14406, N14400, N5279, N4902);
or OR2 (N14407, N14403, N2915);
xor XOR2 (N14408, N14407, N4039);
xor XOR2 (N14409, N14408, N14019);
xor XOR2 (N14410, N14405, N6032);
not NOT1 (N14411, N14409);
xor XOR2 (N14412, N14394, N9339);
buf BUF1 (N14413, N14404);
buf BUF1 (N14414, N14402);
buf BUF1 (N14415, N14412);
or OR4 (N14416, N14401, N591, N3974, N13251);
and AND4 (N14417, N14389, N13675, N10197, N395);
not NOT1 (N14418, N14410);
not NOT1 (N14419, N14414);
xor XOR2 (N14420, N14411, N8638);
buf BUF1 (N14421, N14420);
and AND3 (N14422, N14418, N13732, N11122);
not NOT1 (N14423, N14421);
buf BUF1 (N14424, N14413);
or OR2 (N14425, N14417, N9909);
nand NAND2 (N14426, N14391, N11332);
nor NOR3 (N14427, N14385, N8582, N4101);
nand NAND3 (N14428, N14415, N2534, N10882);
nor NOR2 (N14429, N14426, N13364);
not NOT1 (N14430, N14424);
not NOT1 (N14431, N14406);
nand NAND2 (N14432, N14428, N8578);
or OR4 (N14433, N14423, N8886, N6038, N2652);
xor XOR2 (N14434, N14419, N3173);
xor XOR2 (N14435, N14430, N517);
xor XOR2 (N14436, N14427, N275);
nor NOR2 (N14437, N14416, N2541);
and AND3 (N14438, N14433, N13274, N5048);
nor NOR4 (N14439, N14425, N1159, N4974, N9974);
and AND3 (N14440, N14435, N13197, N782);
nand NAND3 (N14441, N14437, N7702, N14432);
and AND2 (N14442, N4479, N13824);
and AND2 (N14443, N14438, N14395);
buf BUF1 (N14444, N14429);
or OR4 (N14445, N14439, N12428, N10711, N13282);
buf BUF1 (N14446, N14443);
nand NAND4 (N14447, N14422, N13157, N9708, N2773);
or OR2 (N14448, N14431, N13104);
and AND3 (N14449, N14445, N2407, N14283);
or OR2 (N14450, N14434, N12811);
and AND4 (N14451, N14440, N8347, N424, N6024);
or OR2 (N14452, N14442, N13996);
buf BUF1 (N14453, N14447);
not NOT1 (N14454, N14451);
buf BUF1 (N14455, N14453);
xor XOR2 (N14456, N14452, N12774);
not NOT1 (N14457, N14449);
not NOT1 (N14458, N14457);
not NOT1 (N14459, N14436);
buf BUF1 (N14460, N14441);
nor NOR3 (N14461, N14444, N2777, N8459);
nor NOR2 (N14462, N14456, N11114);
not NOT1 (N14463, N14446);
nor NOR2 (N14464, N14462, N14270);
or OR4 (N14465, N14460, N11406, N1958, N13368);
xor XOR2 (N14466, N14448, N13652);
not NOT1 (N14467, N14466);
buf BUF1 (N14468, N14454);
buf BUF1 (N14469, N14450);
not NOT1 (N14470, N14465);
and AND2 (N14471, N14461, N7820);
xor XOR2 (N14472, N14469, N1764);
buf BUF1 (N14473, N14455);
and AND2 (N14474, N14463, N8560);
and AND2 (N14475, N14470, N14465);
and AND4 (N14476, N14471, N7724, N4197, N6753);
and AND2 (N14477, N14473, N10698);
and AND2 (N14478, N14477, N1657);
nand NAND2 (N14479, N14459, N1511);
nor NOR2 (N14480, N14474, N990);
and AND4 (N14481, N14479, N10092, N11519, N12355);
or OR2 (N14482, N14478, N5240);
and AND2 (N14483, N14482, N2777);
and AND2 (N14484, N14483, N12360);
buf BUF1 (N14485, N14480);
and AND3 (N14486, N14472, N10358, N12083);
nor NOR2 (N14487, N14485, N13795);
or OR4 (N14488, N14481, N8396, N2010, N5964);
or OR4 (N14489, N14488, N643, N2744, N5353);
buf BUF1 (N14490, N14464);
xor XOR2 (N14491, N14486, N13544);
nand NAND4 (N14492, N14487, N3909, N7349, N11947);
not NOT1 (N14493, N14489);
xor XOR2 (N14494, N14492, N2803);
buf BUF1 (N14495, N14458);
and AND4 (N14496, N14475, N12114, N4722, N5720);
or OR4 (N14497, N14495, N5979, N11630, N1766);
and AND4 (N14498, N14494, N7456, N9176, N14441);
nor NOR4 (N14499, N14467, N5749, N11396, N13200);
and AND3 (N14500, N14491, N14202, N1154);
not NOT1 (N14501, N14498);
nor NOR2 (N14502, N14499, N2254);
and AND4 (N14503, N14468, N5112, N3893, N2123);
and AND2 (N14504, N14496, N10474);
buf BUF1 (N14505, N14502);
and AND2 (N14506, N14503, N8024);
nor NOR2 (N14507, N14506, N11096);
nor NOR2 (N14508, N14505, N2241);
not NOT1 (N14509, N14493);
and AND4 (N14510, N14501, N11596, N2242, N1896);
and AND4 (N14511, N14484, N1935, N11677, N5599);
and AND4 (N14512, N14511, N10583, N4186, N5526);
nand NAND3 (N14513, N14508, N5546, N401);
nor NOR2 (N14514, N14500, N2949);
nand NAND2 (N14515, N14512, N9842);
xor XOR2 (N14516, N14514, N10012);
buf BUF1 (N14517, N14504);
buf BUF1 (N14518, N14517);
xor XOR2 (N14519, N14513, N2507);
and AND2 (N14520, N14509, N13479);
xor XOR2 (N14521, N14519, N153);
nor NOR3 (N14522, N14510, N13634, N3768);
nand NAND4 (N14523, N14497, N10066, N6380, N11503);
nand NAND2 (N14524, N14476, N2170);
buf BUF1 (N14525, N14524);
nor NOR3 (N14526, N14525, N11516, N8275);
nor NOR4 (N14527, N14490, N6459, N12005, N4133);
or OR2 (N14528, N14523, N6590);
or OR3 (N14529, N14527, N9514, N5384);
or OR3 (N14530, N14529, N6387, N3016);
nor NOR4 (N14531, N14520, N12853, N10691, N1826);
and AND4 (N14532, N14515, N13003, N10535, N7942);
xor XOR2 (N14533, N14522, N10623);
and AND3 (N14534, N14516, N12392, N7721);
and AND4 (N14535, N14528, N13726, N7770, N9550);
buf BUF1 (N14536, N14532);
not NOT1 (N14537, N14531);
buf BUF1 (N14538, N14507);
and AND3 (N14539, N14536, N2031, N5915);
or OR2 (N14540, N14535, N5920);
buf BUF1 (N14541, N14526);
xor XOR2 (N14542, N14539, N10848);
buf BUF1 (N14543, N14542);
not NOT1 (N14544, N14538);
nand NAND2 (N14545, N14541, N8039);
not NOT1 (N14546, N14540);
or OR4 (N14547, N14546, N6538, N8843, N6902);
and AND2 (N14548, N14521, N10260);
xor XOR2 (N14549, N14534, N3961);
and AND4 (N14550, N14545, N8735, N3929, N5330);
xor XOR2 (N14551, N14518, N5279);
nor NOR3 (N14552, N14530, N2944, N8750);
buf BUF1 (N14553, N14550);
xor XOR2 (N14554, N14552, N13155);
and AND2 (N14555, N14549, N5046);
or OR3 (N14556, N14537, N13972, N6238);
nand NAND2 (N14557, N14556, N11559);
and AND4 (N14558, N14544, N5299, N12073, N11415);
nor NOR2 (N14559, N14555, N7954);
nor NOR2 (N14560, N14548, N14056);
and AND2 (N14561, N14533, N5756);
xor XOR2 (N14562, N14554, N9317);
nor NOR4 (N14563, N14543, N6846, N13161, N11162);
buf BUF1 (N14564, N14559);
not NOT1 (N14565, N14563);
nand NAND3 (N14566, N14562, N10122, N3525);
not NOT1 (N14567, N14560);
and AND3 (N14568, N14558, N11068, N6027);
or OR4 (N14569, N14557, N11574, N12282, N6346);
xor XOR2 (N14570, N14566, N3559);
nand NAND2 (N14571, N14565, N12808);
xor XOR2 (N14572, N14568, N12534);
buf BUF1 (N14573, N14572);
and AND4 (N14574, N14570, N10536, N7264, N8680);
or OR4 (N14575, N14564, N10761, N11562, N1899);
and AND3 (N14576, N14569, N140, N12178);
nor NOR3 (N14577, N14576, N376, N11123);
not NOT1 (N14578, N14561);
or OR4 (N14579, N14573, N4689, N8018, N10852);
buf BUF1 (N14580, N14575);
xor XOR2 (N14581, N14551, N9107);
buf BUF1 (N14582, N14579);
xor XOR2 (N14583, N14547, N9762);
xor XOR2 (N14584, N14553, N11537);
nand NAND2 (N14585, N14580, N9025);
and AND4 (N14586, N14585, N5379, N5381, N11085);
and AND4 (N14587, N14571, N13752, N10513, N9773);
or OR4 (N14588, N14584, N13141, N11891, N6486);
or OR3 (N14589, N14588, N12635, N8360);
nand NAND4 (N14590, N14589, N4018, N4256, N623);
not NOT1 (N14591, N14577);
not NOT1 (N14592, N14567);
not NOT1 (N14593, N14574);
or OR2 (N14594, N14593, N6095);
buf BUF1 (N14595, N14592);
buf BUF1 (N14596, N14590);
buf BUF1 (N14597, N14582);
or OR3 (N14598, N14578, N4071, N9384);
xor XOR2 (N14599, N14595, N7845);
nor NOR2 (N14600, N14597, N6195);
or OR3 (N14601, N14600, N1488, N2947);
nand NAND2 (N14602, N14598, N2258);
buf BUF1 (N14603, N14596);
nand NAND4 (N14604, N14599, N8605, N11688, N10746);
buf BUF1 (N14605, N14586);
nor NOR4 (N14606, N14602, N11049, N2751, N3478);
buf BUF1 (N14607, N14594);
or OR2 (N14608, N14603, N12382);
xor XOR2 (N14609, N14581, N4169);
and AND4 (N14610, N14606, N4058, N7061, N11609);
xor XOR2 (N14611, N14604, N1198);
not NOT1 (N14612, N14608);
or OR2 (N14613, N14609, N12216);
and AND3 (N14614, N14583, N11194, N7997);
xor XOR2 (N14615, N14587, N12246);
and AND4 (N14616, N14591, N8998, N6389, N2315);
nor NOR3 (N14617, N14605, N1336, N8224);
buf BUF1 (N14618, N14616);
nor NOR3 (N14619, N14610, N6433, N10375);
xor XOR2 (N14620, N14615, N3425);
or OR2 (N14621, N14617, N1008);
xor XOR2 (N14622, N14618, N1000);
not NOT1 (N14623, N14612);
buf BUF1 (N14624, N14607);
and AND3 (N14625, N14614, N14619, N2124);
and AND2 (N14626, N3924, N8987);
or OR4 (N14627, N14624, N9726, N358, N11434);
nor NOR2 (N14628, N14621, N6499);
xor XOR2 (N14629, N14620, N513);
or OR3 (N14630, N14626, N14579, N7633);
nand NAND4 (N14631, N14627, N11304, N5077, N1712);
buf BUF1 (N14632, N14628);
not NOT1 (N14633, N14601);
not NOT1 (N14634, N14629);
or OR2 (N14635, N14611, N13219);
or OR2 (N14636, N14623, N4032);
nand NAND3 (N14637, N14635, N14140, N767);
or OR4 (N14638, N14632, N7979, N703, N10537);
xor XOR2 (N14639, N14634, N7730);
xor XOR2 (N14640, N14638, N457);
and AND2 (N14641, N14622, N7785);
xor XOR2 (N14642, N14640, N4896);
buf BUF1 (N14643, N14633);
nor NOR3 (N14644, N14637, N476, N7761);
nand NAND3 (N14645, N14631, N7516, N1040);
and AND4 (N14646, N14630, N6357, N12897, N12717);
not NOT1 (N14647, N14643);
not NOT1 (N14648, N14644);
not NOT1 (N14649, N14636);
nor NOR4 (N14650, N14642, N1077, N9118, N1858);
buf BUF1 (N14651, N14641);
or OR4 (N14652, N14639, N7579, N8929, N9308);
nor NOR4 (N14653, N14650, N12029, N6710, N11754);
nor NOR2 (N14654, N14651, N11747);
nand NAND2 (N14655, N14654, N11133);
not NOT1 (N14656, N14647);
or OR3 (N14657, N14625, N2751, N6201);
nor NOR3 (N14658, N14648, N11711, N426);
xor XOR2 (N14659, N14658, N11278);
nand NAND4 (N14660, N14656, N11418, N4898, N7706);
not NOT1 (N14661, N14613);
or OR4 (N14662, N14652, N3416, N2047, N6390);
nand NAND3 (N14663, N14655, N9602, N11073);
buf BUF1 (N14664, N14663);
xor XOR2 (N14665, N14662, N14501);
nand NAND2 (N14666, N14657, N12380);
buf BUF1 (N14667, N14653);
buf BUF1 (N14668, N14660);
xor XOR2 (N14669, N14661, N4459);
nand NAND2 (N14670, N14668, N2922);
xor XOR2 (N14671, N14649, N2476);
not NOT1 (N14672, N14646);
xor XOR2 (N14673, N14667, N12403);
or OR3 (N14674, N14659, N5097, N13582);
xor XOR2 (N14675, N14669, N11487);
xor XOR2 (N14676, N14664, N10772);
xor XOR2 (N14677, N14674, N5913);
not NOT1 (N14678, N14676);
buf BUF1 (N14679, N14675);
and AND4 (N14680, N14673, N8788, N12368, N10931);
nor NOR4 (N14681, N14680, N9830, N6070, N1643);
xor XOR2 (N14682, N14678, N976);
and AND3 (N14683, N14666, N13109, N3844);
and AND3 (N14684, N14670, N797, N3183);
and AND4 (N14685, N14683, N2525, N10069, N7655);
nor NOR2 (N14686, N14679, N11090);
xor XOR2 (N14687, N14645, N1651);
nand NAND3 (N14688, N14682, N4529, N4808);
nand NAND4 (N14689, N14685, N11003, N6557, N11548);
or OR4 (N14690, N14686, N11469, N9047, N7123);
nor NOR2 (N14691, N14688, N9075);
nand NAND4 (N14692, N14681, N11741, N199, N8838);
nor NOR4 (N14693, N14684, N8193, N3992, N4741);
nand NAND3 (N14694, N14692, N11464, N10766);
and AND4 (N14695, N14691, N11604, N1142, N6101);
nand NAND4 (N14696, N14689, N9071, N417, N1437);
not NOT1 (N14697, N14693);
and AND3 (N14698, N14697, N10804, N5448);
or OR2 (N14699, N14690, N556);
nor NOR2 (N14700, N14672, N2274);
or OR2 (N14701, N14699, N6376);
not NOT1 (N14702, N14696);
buf BUF1 (N14703, N14694);
not NOT1 (N14704, N14701);
or OR3 (N14705, N14665, N10367, N10634);
nand NAND3 (N14706, N14677, N2363, N10060);
xor XOR2 (N14707, N14671, N12162);
and AND4 (N14708, N14700, N12489, N293, N8126);
buf BUF1 (N14709, N14698);
buf BUF1 (N14710, N14705);
nor NOR4 (N14711, N14704, N13616, N11702, N3055);
and AND3 (N14712, N14707, N451, N14202);
nor NOR3 (N14713, N14710, N7114, N11687);
nor NOR4 (N14714, N14703, N12468, N12765, N9437);
buf BUF1 (N14715, N14713);
xor XOR2 (N14716, N14708, N657);
and AND3 (N14717, N14714, N8416, N2950);
not NOT1 (N14718, N14702);
and AND4 (N14719, N14712, N12233, N1158, N12195);
nand NAND4 (N14720, N14687, N8359, N3370, N4149);
nand NAND4 (N14721, N14716, N3587, N14261, N11700);
not NOT1 (N14722, N14695);
xor XOR2 (N14723, N14717, N4206);
buf BUF1 (N14724, N14721);
or OR2 (N14725, N14718, N11796);
nand NAND2 (N14726, N14722, N4307);
nor NOR3 (N14727, N14719, N4679, N6908);
not NOT1 (N14728, N14723);
nand NAND3 (N14729, N14728, N5636, N10425);
nand NAND3 (N14730, N14727, N11544, N10993);
buf BUF1 (N14731, N14715);
not NOT1 (N14732, N14706);
xor XOR2 (N14733, N14729, N6744);
buf BUF1 (N14734, N14732);
xor XOR2 (N14735, N14726, N1646);
not NOT1 (N14736, N14733);
nor NOR2 (N14737, N14711, N5142);
not NOT1 (N14738, N14730);
xor XOR2 (N14739, N14725, N12314);
or OR4 (N14740, N14734, N6272, N10990, N4131);
nor NOR4 (N14741, N14737, N4252, N4935, N7135);
or OR2 (N14742, N14739, N8698);
or OR3 (N14743, N14720, N8613, N12346);
buf BUF1 (N14744, N14724);
not NOT1 (N14745, N14709);
nor NOR2 (N14746, N14738, N8051);
buf BUF1 (N14747, N14743);
or OR4 (N14748, N14744, N8582, N14004, N7884);
not NOT1 (N14749, N14741);
or OR2 (N14750, N14746, N9957);
and AND4 (N14751, N14745, N12743, N11977, N8219);
nand NAND3 (N14752, N14742, N4860, N771);
buf BUF1 (N14753, N14740);
not NOT1 (N14754, N14736);
xor XOR2 (N14755, N14748, N5692);
or OR4 (N14756, N14752, N9735, N7906, N646);
or OR4 (N14757, N14735, N8402, N6787, N4689);
xor XOR2 (N14758, N14754, N10738);
nor NOR3 (N14759, N14751, N383, N5280);
buf BUF1 (N14760, N14731);
not NOT1 (N14761, N14758);
nor NOR2 (N14762, N14760, N1139);
nor NOR3 (N14763, N14756, N13872, N1131);
nor NOR2 (N14764, N14749, N7109);
and AND2 (N14765, N14753, N9365);
nand NAND3 (N14766, N14762, N11359, N732);
or OR2 (N14767, N14755, N7844);
xor XOR2 (N14768, N14750, N12008);
xor XOR2 (N14769, N14765, N8267);
nand NAND2 (N14770, N14768, N7287);
or OR3 (N14771, N14770, N2590, N7611);
not NOT1 (N14772, N14757);
nand NAND3 (N14773, N14747, N12600, N7326);
or OR4 (N14774, N14773, N3767, N8346, N8100);
xor XOR2 (N14775, N14761, N12348);
and AND2 (N14776, N14774, N9628);
and AND2 (N14777, N14759, N2904);
nand NAND4 (N14778, N14767, N4746, N5785, N5917);
or OR3 (N14779, N14775, N6154, N11967);
xor XOR2 (N14780, N14769, N986);
not NOT1 (N14781, N14776);
xor XOR2 (N14782, N14772, N11567);
xor XOR2 (N14783, N14778, N9834);
xor XOR2 (N14784, N14779, N5227);
nor NOR3 (N14785, N14777, N4839, N1069);
or OR2 (N14786, N14780, N6888);
nor NOR3 (N14787, N14781, N2413, N10794);
buf BUF1 (N14788, N14766);
nand NAND2 (N14789, N14785, N12198);
nor NOR3 (N14790, N14782, N5705, N13068);
and AND2 (N14791, N14763, N11299);
nor NOR2 (N14792, N14789, N5726);
xor XOR2 (N14793, N14764, N3881);
or OR4 (N14794, N14783, N7403, N12501, N69);
buf BUF1 (N14795, N14786);
or OR2 (N14796, N14784, N9380);
nor NOR2 (N14797, N14795, N12261);
nand NAND2 (N14798, N14787, N13482);
nand NAND3 (N14799, N14771, N360, N9363);
or OR3 (N14800, N14790, N2730, N10898);
xor XOR2 (N14801, N14799, N3739);
nor NOR3 (N14802, N14793, N9536, N13027);
or OR2 (N14803, N14797, N4294);
nand NAND2 (N14804, N14798, N2248);
buf BUF1 (N14805, N14800);
buf BUF1 (N14806, N14794);
nor NOR3 (N14807, N14805, N6549, N12929);
or OR4 (N14808, N14806, N10538, N13803, N6569);
buf BUF1 (N14809, N14788);
and AND4 (N14810, N14803, N6867, N11173, N10856);
nor NOR4 (N14811, N14791, N8175, N2261, N10384);
nand NAND4 (N14812, N14796, N580, N12078, N11633);
not NOT1 (N14813, N14808);
nand NAND3 (N14814, N14804, N5854, N4212);
not NOT1 (N14815, N14802);
not NOT1 (N14816, N14792);
not NOT1 (N14817, N14813);
and AND3 (N14818, N14812, N14164, N3361);
buf BUF1 (N14819, N14809);
nand NAND3 (N14820, N14816, N9, N3235);
not NOT1 (N14821, N14820);
xor XOR2 (N14822, N14821, N644);
and AND3 (N14823, N14817, N1999, N14787);
xor XOR2 (N14824, N14807, N9072);
not NOT1 (N14825, N14824);
and AND2 (N14826, N14822, N489);
and AND2 (N14827, N14825, N8820);
and AND2 (N14828, N14811, N14575);
not NOT1 (N14829, N14827);
buf BUF1 (N14830, N14815);
and AND2 (N14831, N14826, N7174);
xor XOR2 (N14832, N14829, N4348);
nor NOR4 (N14833, N14823, N1835, N7866, N2619);
nand NAND4 (N14834, N14831, N5639, N14367, N6950);
not NOT1 (N14835, N14834);
and AND4 (N14836, N14835, N633, N7405, N12996);
not NOT1 (N14837, N14818);
and AND2 (N14838, N14836, N10467);
xor XOR2 (N14839, N14810, N4127);
and AND2 (N14840, N14828, N717);
buf BUF1 (N14841, N14840);
and AND3 (N14842, N14838, N8263, N14574);
and AND4 (N14843, N14819, N7233, N697, N10192);
xor XOR2 (N14844, N14841, N9656);
nor NOR3 (N14845, N14814, N8659, N4391);
xor XOR2 (N14846, N14844, N10017);
nor NOR2 (N14847, N14845, N11778);
xor XOR2 (N14848, N14801, N12515);
not NOT1 (N14849, N14837);
buf BUF1 (N14850, N14830);
not NOT1 (N14851, N14839);
xor XOR2 (N14852, N14851, N14627);
not NOT1 (N14853, N14833);
buf BUF1 (N14854, N14832);
buf BUF1 (N14855, N14843);
not NOT1 (N14856, N14850);
or OR4 (N14857, N14848, N6606, N8866, N2926);
and AND3 (N14858, N14853, N14362, N7036);
xor XOR2 (N14859, N14849, N4038);
xor XOR2 (N14860, N14859, N12827);
not NOT1 (N14861, N14842);
and AND2 (N14862, N14854, N1861);
or OR2 (N14863, N14862, N10640);
not NOT1 (N14864, N14856);
buf BUF1 (N14865, N14861);
xor XOR2 (N14866, N14858, N8160);
and AND4 (N14867, N14864, N11132, N3071, N11364);
not NOT1 (N14868, N14846);
buf BUF1 (N14869, N14857);
or OR3 (N14870, N14852, N508, N9660);
and AND2 (N14871, N14855, N12439);
and AND2 (N14872, N14869, N14052);
nand NAND4 (N14873, N14865, N14060, N4177, N6351);
and AND3 (N14874, N14873, N8730, N2531);
not NOT1 (N14875, N14860);
buf BUF1 (N14876, N14872);
or OR3 (N14877, N14875, N9988, N9237);
or OR3 (N14878, N14874, N3315, N1938);
xor XOR2 (N14879, N14878, N10914);
xor XOR2 (N14880, N14868, N2288);
xor XOR2 (N14881, N14876, N496);
not NOT1 (N14882, N14881);
xor XOR2 (N14883, N14870, N5195);
xor XOR2 (N14884, N14877, N9714);
buf BUF1 (N14885, N14883);
nand NAND3 (N14886, N14884, N2371, N7702);
and AND4 (N14887, N14882, N6776, N12794, N3174);
nor NOR3 (N14888, N14880, N8756, N8166);
nand NAND3 (N14889, N14863, N9016, N4941);
and AND3 (N14890, N14866, N9254, N12175);
or OR3 (N14891, N14887, N14880, N9907);
not NOT1 (N14892, N14889);
nor NOR3 (N14893, N14891, N10954, N3698);
not NOT1 (N14894, N14892);
nand NAND4 (N14895, N14888, N12828, N2734, N9218);
and AND4 (N14896, N14867, N2172, N14322, N3260);
not NOT1 (N14897, N14890);
buf BUF1 (N14898, N14896);
buf BUF1 (N14899, N14847);
buf BUF1 (N14900, N14879);
xor XOR2 (N14901, N14893, N14539);
and AND4 (N14902, N14886, N7684, N7113, N4153);
buf BUF1 (N14903, N14899);
or OR2 (N14904, N14894, N8333);
xor XOR2 (N14905, N14902, N13147);
nand NAND2 (N14906, N14901, N5962);
nor NOR4 (N14907, N14897, N1756, N8593, N10934);
not NOT1 (N14908, N14900);
or OR4 (N14909, N14907, N5018, N543, N5585);
and AND3 (N14910, N14885, N9393, N14129);
xor XOR2 (N14911, N14898, N1161);
and AND3 (N14912, N14905, N12937, N8310);
xor XOR2 (N14913, N14908, N12702);
and AND2 (N14914, N14909, N10507);
not NOT1 (N14915, N14914);
nand NAND2 (N14916, N14910, N10496);
not NOT1 (N14917, N14915);
or OR2 (N14918, N14904, N10013);
nand NAND4 (N14919, N14903, N13951, N225, N3279);
xor XOR2 (N14920, N14918, N578);
nand NAND4 (N14921, N14912, N11534, N14437, N10487);
buf BUF1 (N14922, N14921);
or OR2 (N14923, N14917, N9670);
and AND2 (N14924, N14871, N4729);
nor NOR4 (N14925, N14924, N1767, N7404, N12974);
buf BUF1 (N14926, N14922);
buf BUF1 (N14927, N14895);
or OR2 (N14928, N14906, N3053);
and AND3 (N14929, N14911, N4210, N13268);
buf BUF1 (N14930, N14929);
nand NAND4 (N14931, N14923, N12507, N10351, N3349);
and AND4 (N14932, N14925, N6876, N4594, N3101);
buf BUF1 (N14933, N14927);
or OR2 (N14934, N14930, N4375);
or OR4 (N14935, N14928, N232, N9521, N4509);
nand NAND2 (N14936, N14919, N5033);
nor NOR2 (N14937, N14920, N7951);
nor NOR4 (N14938, N14933, N12246, N13324, N606);
or OR2 (N14939, N14916, N9886);
xor XOR2 (N14940, N14931, N3850);
nand NAND2 (N14941, N14935, N13204);
not NOT1 (N14942, N14937);
or OR2 (N14943, N14926, N12412);
not NOT1 (N14944, N14913);
buf BUF1 (N14945, N14939);
xor XOR2 (N14946, N14941, N10000);
or OR2 (N14947, N14938, N3197);
or OR2 (N14948, N14943, N10321);
and AND4 (N14949, N14946, N4745, N9330, N14196);
nor NOR3 (N14950, N14944, N11398, N4336);
nor NOR4 (N14951, N14949, N6774, N9002, N3554);
and AND3 (N14952, N14951, N11534, N1641);
buf BUF1 (N14953, N14948);
or OR2 (N14954, N14953, N7678);
xor XOR2 (N14955, N14942, N3790);
nand NAND2 (N14956, N14936, N5573);
nor NOR2 (N14957, N14956, N2988);
buf BUF1 (N14958, N14934);
and AND3 (N14959, N14947, N13234, N7775);
or OR3 (N14960, N14959, N5114, N8196);
buf BUF1 (N14961, N14952);
and AND3 (N14962, N14960, N13658, N4699);
or OR2 (N14963, N14955, N11744);
and AND3 (N14964, N14945, N14160, N14441);
and AND4 (N14965, N14963, N4260, N4049, N12890);
nor NOR3 (N14966, N14932, N8001, N3246);
nand NAND4 (N14967, N14962, N12359, N7637, N8317);
or OR2 (N14968, N14954, N14904);
xor XOR2 (N14969, N14968, N9829);
xor XOR2 (N14970, N14967, N14083);
xor XOR2 (N14971, N14940, N12229);
nand NAND2 (N14972, N14957, N1910);
nand NAND3 (N14973, N14970, N11783, N14555);
xor XOR2 (N14974, N14971, N6388);
xor XOR2 (N14975, N14973, N7752);
xor XOR2 (N14976, N14965, N9210);
not NOT1 (N14977, N14958);
nand NAND4 (N14978, N14964, N9042, N4703, N5335);
nand NAND4 (N14979, N14978, N11191, N4129, N3272);
buf BUF1 (N14980, N14974);
nand NAND4 (N14981, N14950, N2312, N6582, N4815);
not NOT1 (N14982, N14969);
not NOT1 (N14983, N14972);
buf BUF1 (N14984, N14966);
xor XOR2 (N14985, N14976, N9940);
or OR2 (N14986, N14961, N2060);
buf BUF1 (N14987, N14984);
nor NOR3 (N14988, N14979, N1294, N10088);
and AND4 (N14989, N14985, N14486, N12274, N394);
not NOT1 (N14990, N14987);
nor NOR2 (N14991, N14990, N1776);
nor NOR3 (N14992, N14981, N9966, N477);
nand NAND3 (N14993, N14988, N5758, N4566);
buf BUF1 (N14994, N14975);
and AND2 (N14995, N14993, N5621);
and AND4 (N14996, N14991, N11600, N14169, N7941);
buf BUF1 (N14997, N14992);
nor NOR2 (N14998, N14982, N2851);
and AND4 (N14999, N14998, N10704, N6072, N4051);
nand NAND2 (N15000, N14997, N11483);
not NOT1 (N15001, N14986);
not NOT1 (N15002, N14996);
xor XOR2 (N15003, N14999, N1376);
and AND4 (N15004, N15000, N6963, N438, N10829);
nor NOR2 (N15005, N14995, N1384);
xor XOR2 (N15006, N15004, N10477);
and AND4 (N15007, N15005, N11825, N12193, N12053);
nand NAND2 (N15008, N14977, N13935);
xor XOR2 (N15009, N14994, N13234);
or OR3 (N15010, N15003, N12608, N3456);
xor XOR2 (N15011, N15001, N13716);
xor XOR2 (N15012, N15010, N7893);
nand NAND3 (N15013, N14980, N14204, N4299);
nor NOR3 (N15014, N15013, N10710, N13834);
buf BUF1 (N15015, N15007);
buf BUF1 (N15016, N15011);
and AND2 (N15017, N15008, N2258);
nand NAND4 (N15018, N15002, N842, N1577, N5876);
xor XOR2 (N15019, N14983, N5231);
buf BUF1 (N15020, N15009);
xor XOR2 (N15021, N15012, N12490);
not NOT1 (N15022, N15020);
xor XOR2 (N15023, N15018, N14327);
buf BUF1 (N15024, N14989);
or OR2 (N15025, N15015, N7505);
and AND4 (N15026, N15024, N7851, N1296, N4478);
buf BUF1 (N15027, N15026);
nor NOR2 (N15028, N15014, N2576);
nand NAND2 (N15029, N15022, N1983);
or OR2 (N15030, N15016, N12011);
not NOT1 (N15031, N15023);
nor NOR2 (N15032, N15031, N4166);
nand NAND4 (N15033, N15029, N2399, N6324, N10833);
and AND4 (N15034, N15027, N4295, N8582, N11853);
buf BUF1 (N15035, N15030);
buf BUF1 (N15036, N15028);
buf BUF1 (N15037, N15019);
xor XOR2 (N15038, N15035, N7130);
buf BUF1 (N15039, N15037);
xor XOR2 (N15040, N15038, N8397);
nand NAND2 (N15041, N15021, N2053);
buf BUF1 (N15042, N15039);
or OR4 (N15043, N15034, N11873, N7957, N3619);
not NOT1 (N15044, N15032);
and AND3 (N15045, N15042, N13124, N10133);
or OR2 (N15046, N15044, N6310);
xor XOR2 (N15047, N15025, N4499);
and AND2 (N15048, N15040, N14700);
nor NOR2 (N15049, N15033, N8684);
and AND4 (N15050, N15049, N2588, N293, N10571);
nor NOR4 (N15051, N15045, N4806, N10481, N10146);
or OR3 (N15052, N15036, N12427, N7230);
or OR2 (N15053, N15006, N796);
xor XOR2 (N15054, N15047, N3005);
and AND2 (N15055, N15050, N7326);
or OR3 (N15056, N15052, N187, N4356);
or OR2 (N15057, N15043, N2462);
nand NAND4 (N15058, N15048, N6321, N2622, N3087);
nor NOR3 (N15059, N15054, N10904, N9540);
not NOT1 (N15060, N15059);
and AND4 (N15061, N15055, N11444, N12222, N8406);
or OR2 (N15062, N15058, N14421);
and AND3 (N15063, N15053, N13368, N2756);
or OR4 (N15064, N15046, N1818, N13692, N3359);
not NOT1 (N15065, N15063);
nand NAND4 (N15066, N15061, N13750, N8327, N3404);
not NOT1 (N15067, N15060);
and AND3 (N15068, N15065, N10637, N11897);
and AND2 (N15069, N15064, N4014);
or OR4 (N15070, N15062, N6312, N4353, N7645);
buf BUF1 (N15071, N15069);
and AND2 (N15072, N15041, N14762);
and AND3 (N15073, N15067, N9147, N5291);
not NOT1 (N15074, N15051);
not NOT1 (N15075, N15072);
buf BUF1 (N15076, N15017);
or OR3 (N15077, N15073, N4072, N14493);
and AND2 (N15078, N15077, N1097);
nor NOR4 (N15079, N15071, N11844, N3148, N502);
buf BUF1 (N15080, N15068);
not NOT1 (N15081, N15080);
buf BUF1 (N15082, N15056);
xor XOR2 (N15083, N15082, N8429);
not NOT1 (N15084, N15070);
not NOT1 (N15085, N15079);
xor XOR2 (N15086, N15075, N7957);
nor NOR4 (N15087, N15057, N6556, N6681, N5103);
not NOT1 (N15088, N15078);
nand NAND3 (N15089, N15066, N11811, N13363);
xor XOR2 (N15090, N15074, N10885);
or OR2 (N15091, N15083, N4792);
buf BUF1 (N15092, N15086);
and AND3 (N15093, N15089, N8746, N9569);
nand NAND3 (N15094, N15084, N9918, N12718);
xor XOR2 (N15095, N15093, N267);
buf BUF1 (N15096, N15094);
xor XOR2 (N15097, N15087, N606);
and AND2 (N15098, N15097, N5927);
and AND2 (N15099, N15088, N3680);
or OR4 (N15100, N15098, N3730, N10072, N7946);
xor XOR2 (N15101, N15081, N9344);
and AND3 (N15102, N15099, N8101, N1066);
nand NAND3 (N15103, N15085, N34, N10315);
or OR4 (N15104, N15091, N11632, N91, N14692);
nor NOR3 (N15105, N15100, N12658, N1616);
nor NOR2 (N15106, N15105, N10996);
not NOT1 (N15107, N15090);
or OR2 (N15108, N15092, N2182);
buf BUF1 (N15109, N15102);
buf BUF1 (N15110, N15109);
buf BUF1 (N15111, N15108);
buf BUF1 (N15112, N15101);
not NOT1 (N15113, N15096);
nand NAND4 (N15114, N15111, N7078, N1886, N2746);
nor NOR3 (N15115, N15106, N8091, N13524);
buf BUF1 (N15116, N15107);
buf BUF1 (N15117, N15112);
nand NAND3 (N15118, N15115, N4824, N10994);
nor NOR2 (N15119, N15076, N7061);
nand NAND2 (N15120, N15118, N2916);
and AND3 (N15121, N15110, N7423, N5072);
xor XOR2 (N15122, N15116, N6343);
buf BUF1 (N15123, N15104);
nor NOR4 (N15124, N15103, N13590, N5409, N12136);
xor XOR2 (N15125, N15114, N12300);
xor XOR2 (N15126, N15095, N1179);
and AND4 (N15127, N15122, N5466, N8723, N11662);
nand NAND3 (N15128, N15117, N12271, N14942);
nor NOR4 (N15129, N15123, N2946, N12085, N11366);
or OR2 (N15130, N15125, N1871);
or OR2 (N15131, N15128, N14673);
and AND2 (N15132, N15119, N14550);
buf BUF1 (N15133, N15129);
or OR4 (N15134, N15133, N2001, N2986, N4098);
or OR2 (N15135, N15132, N9052);
not NOT1 (N15136, N15121);
nor NOR2 (N15137, N15130, N1836);
xor XOR2 (N15138, N15137, N10912);
not NOT1 (N15139, N15126);
nand NAND2 (N15140, N15134, N5450);
not NOT1 (N15141, N15136);
or OR2 (N15142, N15135, N13854);
or OR4 (N15143, N15131, N6544, N7841, N13927);
or OR3 (N15144, N15120, N735, N15074);
not NOT1 (N15145, N15140);
not NOT1 (N15146, N15145);
xor XOR2 (N15147, N15141, N15065);
nand NAND2 (N15148, N15143, N10403);
xor XOR2 (N15149, N15147, N4298);
and AND3 (N15150, N15144, N11197, N4690);
nor NOR4 (N15151, N15113, N8085, N785, N7036);
nor NOR4 (N15152, N15146, N12216, N8360, N6480);
or OR4 (N15153, N15149, N3885, N1281, N5611);
nor NOR4 (N15154, N15139, N1335, N3090, N2111);
buf BUF1 (N15155, N15150);
nand NAND2 (N15156, N15142, N14695);
buf BUF1 (N15157, N15127);
nor NOR3 (N15158, N15148, N7784, N570);
nor NOR4 (N15159, N15154, N6305, N12646, N2394);
buf BUF1 (N15160, N15159);
or OR3 (N15161, N15157, N2156, N3105);
nand NAND2 (N15162, N15158, N1386);
and AND3 (N15163, N15160, N12527, N12481);
nand NAND3 (N15164, N15161, N9765, N13452);
not NOT1 (N15165, N15162);
not NOT1 (N15166, N15156);
xor XOR2 (N15167, N15165, N7156);
not NOT1 (N15168, N15153);
not NOT1 (N15169, N15152);
buf BUF1 (N15170, N15164);
nand NAND4 (N15171, N15151, N7621, N7794, N3667);
buf BUF1 (N15172, N15124);
nor NOR2 (N15173, N15163, N4084);
buf BUF1 (N15174, N15138);
not NOT1 (N15175, N15173);
nand NAND3 (N15176, N15166, N6081, N12932);
and AND4 (N15177, N15172, N5444, N12595, N191);
not NOT1 (N15178, N15176);
not NOT1 (N15179, N15177);
xor XOR2 (N15180, N15168, N1742);
xor XOR2 (N15181, N15171, N1751);
not NOT1 (N15182, N15179);
buf BUF1 (N15183, N15180);
nor NOR3 (N15184, N15167, N3195, N14104);
not NOT1 (N15185, N15175);
and AND3 (N15186, N15174, N13390, N3656);
not NOT1 (N15187, N15155);
or OR3 (N15188, N15185, N11650, N3237);
not NOT1 (N15189, N15187);
xor XOR2 (N15190, N15170, N5666);
not NOT1 (N15191, N15169);
or OR4 (N15192, N15181, N2254, N10630, N6004);
and AND4 (N15193, N15191, N10999, N87, N2054);
xor XOR2 (N15194, N15184, N2480);
and AND3 (N15195, N15189, N9310, N5757);
not NOT1 (N15196, N15182);
nor NOR3 (N15197, N15194, N8430, N6744);
xor XOR2 (N15198, N15195, N748);
not NOT1 (N15199, N15178);
nand NAND2 (N15200, N15196, N10708);
or OR4 (N15201, N15188, N4811, N9353, N11420);
not NOT1 (N15202, N15192);
xor XOR2 (N15203, N15186, N9644);
and AND3 (N15204, N15183, N3594, N10352);
and AND4 (N15205, N15203, N13994, N10326, N199);
and AND4 (N15206, N15205, N12277, N1102, N11348);
and AND2 (N15207, N15204, N1173);
or OR3 (N15208, N15202, N13633, N15127);
and AND4 (N15209, N15198, N14087, N12228, N7884);
nand NAND4 (N15210, N15209, N12767, N12334, N1902);
nand NAND4 (N15211, N15199, N9326, N1787, N2252);
xor XOR2 (N15212, N15200, N14418);
not NOT1 (N15213, N15210);
buf BUF1 (N15214, N15193);
nand NAND4 (N15215, N15213, N14173, N6356, N11573);
and AND3 (N15216, N15206, N8543, N3569);
or OR3 (N15217, N15216, N3411, N5100);
and AND2 (N15218, N15211, N11838);
or OR3 (N15219, N15218, N7564, N3076);
nand NAND4 (N15220, N15197, N6775, N14246, N10522);
nor NOR4 (N15221, N15207, N1754, N6110, N336);
not NOT1 (N15222, N15220);
nor NOR2 (N15223, N15212, N8816);
buf BUF1 (N15224, N15208);
nand NAND3 (N15225, N15217, N5095, N11888);
buf BUF1 (N15226, N15214);
xor XOR2 (N15227, N15225, N13192);
not NOT1 (N15228, N15226);
nand NAND3 (N15229, N15219, N9339, N10306);
and AND2 (N15230, N15229, N3605);
or OR3 (N15231, N15190, N387, N13102);
and AND4 (N15232, N15215, N148, N11791, N6104);
nor NOR2 (N15233, N15201, N12926);
not NOT1 (N15234, N15231);
nor NOR4 (N15235, N15230, N11745, N9079, N2383);
not NOT1 (N15236, N15221);
buf BUF1 (N15237, N15232);
nor NOR4 (N15238, N15222, N498, N4012, N1697);
xor XOR2 (N15239, N15223, N11924);
nand NAND3 (N15240, N15233, N8032, N12425);
and AND3 (N15241, N15236, N1393, N3405);
xor XOR2 (N15242, N15239, N3969);
or OR2 (N15243, N15227, N11939);
not NOT1 (N15244, N15238);
nor NOR2 (N15245, N15241, N1570);
nand NAND3 (N15246, N15245, N775, N12037);
and AND4 (N15247, N15240, N12615, N13073, N8843);
not NOT1 (N15248, N15237);
and AND4 (N15249, N15243, N10762, N8798, N5688);
xor XOR2 (N15250, N15248, N14609);
xor XOR2 (N15251, N15228, N14518);
not NOT1 (N15252, N15224);
nor NOR2 (N15253, N15242, N6904);
or OR4 (N15254, N15244, N10541, N2371, N5941);
not NOT1 (N15255, N15235);
not NOT1 (N15256, N15254);
and AND2 (N15257, N15247, N688);
buf BUF1 (N15258, N15250);
and AND2 (N15259, N15234, N10718);
xor XOR2 (N15260, N15251, N5713);
or OR2 (N15261, N15258, N2869);
and AND2 (N15262, N15259, N1570);
nand NAND3 (N15263, N15260, N13376, N31);
nor NOR2 (N15264, N15249, N3725);
buf BUF1 (N15265, N15253);
nor NOR2 (N15266, N15261, N351);
not NOT1 (N15267, N15255);
xor XOR2 (N15268, N15265, N4498);
and AND2 (N15269, N15262, N14106);
and AND3 (N15270, N15263, N8038, N3849);
not NOT1 (N15271, N15252);
not NOT1 (N15272, N15267);
buf BUF1 (N15273, N15269);
buf BUF1 (N15274, N15266);
nand NAND4 (N15275, N15272, N13129, N1913, N10223);
not NOT1 (N15276, N15275);
not NOT1 (N15277, N15274);
nor NOR4 (N15278, N15246, N43, N735, N1986);
xor XOR2 (N15279, N15271, N9037);
xor XOR2 (N15280, N15268, N1332);
or OR3 (N15281, N15270, N3677, N4938);
and AND2 (N15282, N15279, N9732);
nand NAND2 (N15283, N15277, N8990);
not NOT1 (N15284, N15257);
buf BUF1 (N15285, N15284);
nand NAND3 (N15286, N15282, N2056, N4518);
xor XOR2 (N15287, N15276, N4841);
nor NOR3 (N15288, N15286, N7395, N11995);
and AND2 (N15289, N15273, N13112);
buf BUF1 (N15290, N15283);
buf BUF1 (N15291, N15285);
and AND2 (N15292, N15289, N1786);
nand NAND3 (N15293, N15292, N3212, N7683);
and AND3 (N15294, N15280, N13457, N5244);
and AND2 (N15295, N15287, N3742);
xor XOR2 (N15296, N15278, N12253);
or OR2 (N15297, N15256, N10965);
nor NOR3 (N15298, N15290, N9661, N7543);
nand NAND2 (N15299, N15298, N9734);
not NOT1 (N15300, N15291);
not NOT1 (N15301, N15294);
xor XOR2 (N15302, N15264, N6298);
xor XOR2 (N15303, N15301, N9778);
not NOT1 (N15304, N15296);
buf BUF1 (N15305, N15293);
not NOT1 (N15306, N15304);
or OR2 (N15307, N15306, N4211);
nand NAND4 (N15308, N15281, N2956, N533, N10189);
not NOT1 (N15309, N15295);
and AND4 (N15310, N15308, N10965, N9251, N2438);
xor XOR2 (N15311, N15288, N542);
nor NOR4 (N15312, N15307, N12463, N1262, N4608);
buf BUF1 (N15313, N15300);
and AND2 (N15314, N15303, N6595);
nand NAND2 (N15315, N15297, N3028);
buf BUF1 (N15316, N15312);
and AND4 (N15317, N15299, N873, N11127, N4792);
nand NAND4 (N15318, N15313, N4077, N5228, N10816);
or OR4 (N15319, N15305, N13327, N2530, N6045);
nand NAND4 (N15320, N15316, N7305, N9853, N6443);
or OR4 (N15321, N15319, N7309, N10124, N2278);
xor XOR2 (N15322, N15302, N1894);
nand NAND3 (N15323, N15321, N3819, N11093);
xor XOR2 (N15324, N15317, N10660);
xor XOR2 (N15325, N15314, N13374);
xor XOR2 (N15326, N15311, N6722);
and AND2 (N15327, N15320, N11002);
not NOT1 (N15328, N15324);
not NOT1 (N15329, N15322);
not NOT1 (N15330, N15326);
xor XOR2 (N15331, N15310, N4248);
buf BUF1 (N15332, N15331);
nor NOR2 (N15333, N15329, N6157);
not NOT1 (N15334, N15309);
and AND2 (N15335, N15318, N6472);
nand NAND4 (N15336, N15327, N2681, N3728, N14741);
buf BUF1 (N15337, N15334);
nor NOR4 (N15338, N15325, N8335, N6925, N10595);
nand NAND3 (N15339, N15330, N1246, N9221);
nor NOR4 (N15340, N15338, N5487, N1134, N7041);
and AND4 (N15341, N15323, N5086, N3283, N14767);
buf BUF1 (N15342, N15337);
not NOT1 (N15343, N15328);
xor XOR2 (N15344, N15340, N6830);
and AND3 (N15345, N15333, N14747, N8543);
nand NAND4 (N15346, N15336, N11458, N3738, N13632);
not NOT1 (N15347, N15344);
nand NAND4 (N15348, N15332, N15024, N2511, N8352);
nand NAND2 (N15349, N15341, N3376);
xor XOR2 (N15350, N15335, N7034);
nor NOR3 (N15351, N15343, N7146, N69);
xor XOR2 (N15352, N15315, N5583);
xor XOR2 (N15353, N15352, N4513);
and AND3 (N15354, N15348, N4544, N3138);
xor XOR2 (N15355, N15349, N13116);
xor XOR2 (N15356, N15346, N14581);
buf BUF1 (N15357, N15350);
buf BUF1 (N15358, N15356);
not NOT1 (N15359, N15357);
or OR4 (N15360, N15359, N2785, N9226, N7936);
and AND3 (N15361, N15353, N2655, N11568);
or OR3 (N15362, N15351, N9171, N1598);
nor NOR3 (N15363, N15345, N1736, N8382);
nor NOR2 (N15364, N15347, N13662);
not NOT1 (N15365, N15361);
not NOT1 (N15366, N15360);
nand NAND2 (N15367, N15362, N5543);
or OR3 (N15368, N15367, N5048, N11268);
and AND3 (N15369, N15358, N9774, N13318);
or OR2 (N15370, N15363, N13960);
and AND3 (N15371, N15366, N1331, N10602);
and AND4 (N15372, N15342, N6654, N2049, N399);
nand NAND3 (N15373, N15372, N4319, N7182);
not NOT1 (N15374, N15370);
and AND4 (N15375, N15354, N7213, N14248, N1426);
or OR4 (N15376, N15339, N1054, N1438, N141);
xor XOR2 (N15377, N15376, N8172);
or OR2 (N15378, N15364, N4564);
or OR4 (N15379, N15373, N3750, N5436, N11350);
nand NAND3 (N15380, N15377, N2585, N2235);
not NOT1 (N15381, N15355);
not NOT1 (N15382, N15368);
nand NAND3 (N15383, N15369, N10944, N4410);
or OR4 (N15384, N15365, N11052, N13356, N10383);
or OR4 (N15385, N15375, N9937, N1591, N2964);
nor NOR2 (N15386, N15380, N4831);
nor NOR4 (N15387, N15384, N10448, N5375, N5109);
xor XOR2 (N15388, N15382, N10312);
buf BUF1 (N15389, N15378);
not NOT1 (N15390, N15385);
nand NAND3 (N15391, N15379, N832, N4287);
nor NOR4 (N15392, N15374, N12087, N5161, N3335);
nand NAND2 (N15393, N15389, N5815);
nor NOR2 (N15394, N15386, N6834);
and AND2 (N15395, N15383, N7482);
and AND3 (N15396, N15394, N14652, N3814);
and AND3 (N15397, N15371, N11919, N7647);
not NOT1 (N15398, N15388);
nand NAND2 (N15399, N15396, N7672);
buf BUF1 (N15400, N15395);
buf BUF1 (N15401, N15398);
or OR4 (N15402, N15387, N15035, N10705, N6273);
buf BUF1 (N15403, N15397);
nand NAND3 (N15404, N15403, N15244, N14113);
nand NAND3 (N15405, N15402, N3574, N772);
not NOT1 (N15406, N15401);
buf BUF1 (N15407, N15405);
and AND4 (N15408, N15404, N15180, N3921, N3244);
xor XOR2 (N15409, N15408, N7343);
buf BUF1 (N15410, N15392);
nand NAND2 (N15411, N15391, N12148);
and AND3 (N15412, N15399, N9769, N6669);
and AND4 (N15413, N15411, N4630, N12813, N11890);
buf BUF1 (N15414, N15407);
or OR4 (N15415, N15393, N4883, N4478, N685);
or OR4 (N15416, N15414, N2283, N12287, N222);
buf BUF1 (N15417, N15400);
not NOT1 (N15418, N15410);
xor XOR2 (N15419, N15409, N11018);
not NOT1 (N15420, N15417);
nor NOR4 (N15421, N15420, N4624, N12817, N2724);
or OR4 (N15422, N15418, N12220, N3935, N9308);
or OR2 (N15423, N15422, N3538);
buf BUF1 (N15424, N15421);
not NOT1 (N15425, N15381);
nor NOR3 (N15426, N15406, N2770, N11074);
xor XOR2 (N15427, N15413, N13387);
nor NOR3 (N15428, N15424, N9838, N7694);
nor NOR4 (N15429, N15419, N4780, N3297, N12013);
not NOT1 (N15430, N15416);
nand NAND4 (N15431, N15429, N4872, N6536, N2986);
not NOT1 (N15432, N15431);
and AND4 (N15433, N15415, N7369, N13571, N5862);
not NOT1 (N15434, N15390);
xor XOR2 (N15435, N15430, N2666);
xor XOR2 (N15436, N15412, N12651);
nand NAND4 (N15437, N15427, N5019, N4403, N11966);
nor NOR4 (N15438, N15425, N4737, N11489, N13784);
and AND3 (N15439, N15435, N6967, N10171);
not NOT1 (N15440, N15438);
xor XOR2 (N15441, N15434, N6416);
and AND2 (N15442, N15426, N8081);
or OR3 (N15443, N15428, N2127, N12872);
nor NOR2 (N15444, N15439, N4194);
nor NOR2 (N15445, N15443, N10155);
or OR3 (N15446, N15442, N10452, N6615);
nor NOR4 (N15447, N15436, N2982, N5926, N2894);
nor NOR4 (N15448, N15444, N3083, N9159, N13872);
buf BUF1 (N15449, N15433);
buf BUF1 (N15450, N15449);
nor NOR2 (N15451, N15450, N13793);
and AND2 (N15452, N15440, N10575);
and AND2 (N15453, N15441, N1696);
nor NOR3 (N15454, N15452, N11171, N2395);
nor NOR2 (N15455, N15437, N3425);
xor XOR2 (N15456, N15451, N9414);
buf BUF1 (N15457, N15454);
and AND2 (N15458, N15448, N8020);
xor XOR2 (N15459, N15455, N8506);
xor XOR2 (N15460, N15445, N6234);
or OR4 (N15461, N15447, N10778, N4737, N6105);
and AND2 (N15462, N15459, N11570);
xor XOR2 (N15463, N15462, N369);
nor NOR4 (N15464, N15446, N14537, N3084, N1996);
or OR4 (N15465, N15463, N3780, N12074, N10686);
buf BUF1 (N15466, N15465);
xor XOR2 (N15467, N15461, N7670);
nand NAND2 (N15468, N15456, N7006);
or OR4 (N15469, N15466, N3984, N5710, N14700);
and AND3 (N15470, N15432, N10653, N14296);
and AND3 (N15471, N15470, N11450, N3041);
buf BUF1 (N15472, N15453);
nor NOR2 (N15473, N15457, N13227);
nor NOR3 (N15474, N15423, N13515, N10833);
nor NOR4 (N15475, N15468, N3612, N5516, N5750);
and AND3 (N15476, N15469, N888, N4942);
and AND2 (N15477, N15471, N5931);
nor NOR4 (N15478, N15476, N5292, N6028, N3910);
not NOT1 (N15479, N15477);
buf BUF1 (N15480, N15458);
not NOT1 (N15481, N15474);
xor XOR2 (N15482, N15460, N15141);
buf BUF1 (N15483, N15467);
xor XOR2 (N15484, N15482, N9144);
buf BUF1 (N15485, N15473);
or OR2 (N15486, N15479, N8685);
buf BUF1 (N15487, N15481);
not NOT1 (N15488, N15478);
nand NAND4 (N15489, N15475, N15292, N4111, N9469);
buf BUF1 (N15490, N15483);
or OR3 (N15491, N15480, N5149, N6438);
or OR3 (N15492, N15489, N9581, N14378);
or OR3 (N15493, N15491, N7171, N2906);
or OR4 (N15494, N15490, N1444, N6358, N349);
not NOT1 (N15495, N15487);
xor XOR2 (N15496, N15464, N6721);
not NOT1 (N15497, N15472);
and AND2 (N15498, N15485, N1080);
nand NAND2 (N15499, N15493, N7170);
buf BUF1 (N15500, N15494);
nand NAND2 (N15501, N15488, N1252);
buf BUF1 (N15502, N15496);
buf BUF1 (N15503, N15492);
not NOT1 (N15504, N15499);
or OR3 (N15505, N15503, N1196, N5422);
xor XOR2 (N15506, N15500, N6625);
and AND2 (N15507, N15484, N6684);
nand NAND2 (N15508, N15502, N13874);
nand NAND4 (N15509, N15504, N4309, N9913, N5646);
not NOT1 (N15510, N15507);
xor XOR2 (N15511, N15501, N5155);
xor XOR2 (N15512, N15511, N456);
not NOT1 (N15513, N15505);
nor NOR3 (N15514, N15498, N5671, N2099);
or OR2 (N15515, N15497, N8455);
nor NOR3 (N15516, N15513, N1140, N131);
xor XOR2 (N15517, N15486, N12257);
or OR2 (N15518, N15515, N9984);
buf BUF1 (N15519, N15518);
nor NOR3 (N15520, N15514, N9656, N2610);
or OR2 (N15521, N15517, N14065);
nor NOR2 (N15522, N15510, N4346);
nor NOR2 (N15523, N15509, N1244);
not NOT1 (N15524, N15506);
nand NAND2 (N15525, N15523, N1746);
or OR2 (N15526, N15495, N10093);
not NOT1 (N15527, N15508);
xor XOR2 (N15528, N15519, N4551);
buf BUF1 (N15529, N15522);
or OR3 (N15530, N15526, N1662, N11439);
xor XOR2 (N15531, N15528, N7647);
not NOT1 (N15532, N15524);
buf BUF1 (N15533, N15531);
xor XOR2 (N15534, N15525, N1101);
nand NAND4 (N15535, N15533, N470, N13451, N12909);
or OR4 (N15536, N15529, N2697, N8191, N66);
nor NOR3 (N15537, N15536, N14234, N12963);
and AND4 (N15538, N15537, N4952, N10183, N6561);
not NOT1 (N15539, N15527);
nor NOR4 (N15540, N15534, N4989, N1710, N1903);
nand NAND2 (N15541, N15538, N9264);
and AND4 (N15542, N15541, N13223, N10161, N6293);
nand NAND2 (N15543, N15540, N2950);
or OR4 (N15544, N15512, N14546, N14624, N8186);
or OR4 (N15545, N15539, N8191, N5635, N4365);
nand NAND4 (N15546, N15521, N6262, N10798, N8566);
or OR4 (N15547, N15516, N3687, N14853, N189);
buf BUF1 (N15548, N15535);
and AND4 (N15549, N15548, N7067, N3964, N12529);
nor NOR4 (N15550, N15545, N4439, N9937, N1794);
and AND4 (N15551, N15520, N15202, N6139, N278);
and AND2 (N15552, N15546, N1999);
buf BUF1 (N15553, N15532);
or OR2 (N15554, N15553, N10213);
not NOT1 (N15555, N15530);
nand NAND4 (N15556, N15552, N12652, N14538, N335);
nor NOR4 (N15557, N15551, N8739, N4682, N5172);
nor NOR4 (N15558, N15549, N9575, N10397, N13626);
and AND4 (N15559, N15557, N12601, N8630, N15555);
not NOT1 (N15560, N8047);
nand NAND3 (N15561, N15544, N7095, N8266);
xor XOR2 (N15562, N15543, N4800);
or OR2 (N15563, N15550, N15009);
nor NOR3 (N15564, N15559, N115, N8820);
xor XOR2 (N15565, N15560, N6694);
buf BUF1 (N15566, N15542);
nor NOR3 (N15567, N15562, N14328, N375);
not NOT1 (N15568, N15556);
or OR3 (N15569, N15563, N6472, N5759);
xor XOR2 (N15570, N15567, N1659);
or OR3 (N15571, N15561, N7069, N3578);
nand NAND4 (N15572, N15558, N1496, N13432, N13645);
nand NAND4 (N15573, N15566, N12530, N12814, N10454);
or OR4 (N15574, N15569, N10400, N10969, N5002);
nor NOR2 (N15575, N15568, N2470);
nor NOR4 (N15576, N15564, N13264, N15041, N9002);
not NOT1 (N15577, N15575);
or OR4 (N15578, N15576, N13226, N9437, N15457);
and AND2 (N15579, N15547, N1030);
xor XOR2 (N15580, N15571, N13521);
not NOT1 (N15581, N15554);
buf BUF1 (N15582, N15578);
nand NAND3 (N15583, N15581, N3430, N2681);
buf BUF1 (N15584, N15579);
nand NAND2 (N15585, N15570, N11412);
nor NOR3 (N15586, N15582, N15199, N1723);
nand NAND4 (N15587, N15583, N6311, N327, N15424);
xor XOR2 (N15588, N15572, N15130);
nor NOR4 (N15589, N15565, N4462, N15022, N6910);
nor NOR4 (N15590, N15580, N10713, N5856, N11269);
and AND2 (N15591, N15587, N14161);
nand NAND3 (N15592, N15585, N10024, N9331);
nor NOR4 (N15593, N15591, N7937, N15547, N11942);
not NOT1 (N15594, N15584);
nand NAND2 (N15595, N15590, N13234);
xor XOR2 (N15596, N15586, N13929);
nor NOR4 (N15597, N15577, N11417, N5017, N2656);
nor NOR2 (N15598, N15596, N11537);
nand NAND3 (N15599, N15592, N8154, N8587);
nor NOR3 (N15600, N15588, N12810, N5423);
xor XOR2 (N15601, N15574, N9069);
and AND2 (N15602, N15600, N4859);
nand NAND3 (N15603, N15573, N2120, N6976);
buf BUF1 (N15604, N15603);
and AND2 (N15605, N15589, N11661);
not NOT1 (N15606, N15594);
buf BUF1 (N15607, N15598);
not NOT1 (N15608, N15602);
or OR2 (N15609, N15597, N5874);
and AND3 (N15610, N15608, N2101, N10240);
xor XOR2 (N15611, N15610, N12540);
xor XOR2 (N15612, N15593, N2349);
and AND4 (N15613, N15612, N13453, N6743, N2582);
nand NAND4 (N15614, N15611, N5752, N11069, N2049);
or OR3 (N15615, N15614, N7078, N2020);
buf BUF1 (N15616, N15607);
nor NOR4 (N15617, N15606, N8335, N9085, N12022);
nor NOR2 (N15618, N15595, N6658);
xor XOR2 (N15619, N15613, N4498);
not NOT1 (N15620, N15601);
nor NOR2 (N15621, N15617, N2531);
buf BUF1 (N15622, N15604);
buf BUF1 (N15623, N15620);
and AND4 (N15624, N15616, N804, N8616, N11963);
buf BUF1 (N15625, N15619);
not NOT1 (N15626, N15618);
xor XOR2 (N15627, N15621, N13272);
not NOT1 (N15628, N15624);
buf BUF1 (N15629, N15625);
nand NAND2 (N15630, N15609, N3510);
nor NOR3 (N15631, N15628, N7378, N13689);
nand NAND2 (N15632, N15630, N7241);
nand NAND2 (N15633, N15626, N259);
not NOT1 (N15634, N15622);
buf BUF1 (N15635, N15605);
buf BUF1 (N15636, N15635);
and AND4 (N15637, N15599, N5992, N10280, N4386);
not NOT1 (N15638, N15627);
not NOT1 (N15639, N15636);
xor XOR2 (N15640, N15637, N14757);
buf BUF1 (N15641, N15640);
buf BUF1 (N15642, N15638);
and AND3 (N15643, N15631, N890, N10812);
xor XOR2 (N15644, N15629, N9024);
nor NOR2 (N15645, N15615, N2387);
or OR4 (N15646, N15639, N5066, N12420, N2760);
and AND2 (N15647, N15633, N3122);
nor NOR2 (N15648, N15646, N7829);
nand NAND3 (N15649, N15641, N3395, N11248);
xor XOR2 (N15650, N15623, N5603);
buf BUF1 (N15651, N15634);
xor XOR2 (N15652, N15650, N9311);
and AND2 (N15653, N15644, N3941);
nand NAND3 (N15654, N15651, N10729, N387);
not NOT1 (N15655, N15645);
xor XOR2 (N15656, N15653, N9657);
nor NOR3 (N15657, N15643, N5030, N7301);
buf BUF1 (N15658, N15649);
and AND3 (N15659, N15648, N11464, N13817);
nand NAND2 (N15660, N15632, N859);
or OR3 (N15661, N15655, N9734, N2844);
xor XOR2 (N15662, N15659, N11063);
xor XOR2 (N15663, N15661, N5428);
and AND2 (N15664, N15652, N2685);
not NOT1 (N15665, N15656);
and AND4 (N15666, N15658, N3936, N11911, N8026);
and AND2 (N15667, N15642, N7133);
not NOT1 (N15668, N15664);
or OR4 (N15669, N15662, N6978, N15132, N5308);
buf BUF1 (N15670, N15666);
nand NAND4 (N15671, N15663, N13386, N11267, N15400);
buf BUF1 (N15672, N15667);
not NOT1 (N15673, N15657);
and AND4 (N15674, N15654, N8456, N7456, N6913);
not NOT1 (N15675, N15647);
xor XOR2 (N15676, N15672, N7419);
and AND4 (N15677, N15665, N9293, N14041, N12363);
or OR4 (N15678, N15673, N7751, N10242, N4389);
not NOT1 (N15679, N15678);
nand NAND2 (N15680, N15674, N14951);
nor NOR2 (N15681, N15668, N8323);
buf BUF1 (N15682, N15670);
xor XOR2 (N15683, N15660, N6839);
nand NAND3 (N15684, N15671, N14761, N10219);
nand NAND4 (N15685, N15682, N5975, N11942, N5759);
nand NAND3 (N15686, N15677, N7810, N14981);
and AND3 (N15687, N15684, N5918, N8847);
buf BUF1 (N15688, N15685);
xor XOR2 (N15689, N15686, N1857);
or OR2 (N15690, N15675, N466);
buf BUF1 (N15691, N15687);
nor NOR3 (N15692, N15683, N11464, N5121);
nor NOR2 (N15693, N15691, N191);
buf BUF1 (N15694, N15669);
buf BUF1 (N15695, N15676);
nor NOR2 (N15696, N15695, N1076);
buf BUF1 (N15697, N15690);
nand NAND2 (N15698, N15696, N6344);
or OR2 (N15699, N15697, N14849);
or OR4 (N15700, N15679, N8670, N14648, N13054);
and AND4 (N15701, N15693, N2382, N15409, N2249);
or OR4 (N15702, N15701, N907, N13653, N8421);
xor XOR2 (N15703, N15689, N12303);
or OR2 (N15704, N15692, N3978);
nor NOR2 (N15705, N15699, N3988);
nand NAND3 (N15706, N15698, N15133, N96);
or OR2 (N15707, N15704, N7704);
nor NOR3 (N15708, N15707, N1861, N14313);
nor NOR3 (N15709, N15705, N15589, N5934);
or OR3 (N15710, N15700, N10816, N9920);
or OR3 (N15711, N15702, N4288, N515);
nand NAND2 (N15712, N15710, N6316);
or OR4 (N15713, N15706, N10539, N11500, N4072);
or OR4 (N15714, N15688, N10340, N5465, N7524);
and AND4 (N15715, N15708, N8487, N4649, N6859);
nand NAND3 (N15716, N15709, N4193, N14167);
buf BUF1 (N15717, N15681);
or OR2 (N15718, N15694, N11761);
not NOT1 (N15719, N15680);
xor XOR2 (N15720, N15711, N416);
nor NOR2 (N15721, N15717, N8255);
buf BUF1 (N15722, N15719);
not NOT1 (N15723, N15722);
nor NOR3 (N15724, N15718, N5460, N2726);
xor XOR2 (N15725, N15715, N6798);
or OR3 (N15726, N15720, N1650, N227);
or OR4 (N15727, N15713, N7300, N1119, N4598);
not NOT1 (N15728, N15723);
not NOT1 (N15729, N15728);
nand NAND2 (N15730, N15724, N12813);
xor XOR2 (N15731, N15703, N11987);
nand NAND4 (N15732, N15726, N9920, N10869, N4912);
nor NOR4 (N15733, N15727, N11149, N8571, N12048);
nand NAND3 (N15734, N15730, N1461, N4054);
xor XOR2 (N15735, N15734, N9679);
nand NAND4 (N15736, N15716, N7575, N7804, N14877);
nor NOR4 (N15737, N15729, N4198, N4036, N5601);
buf BUF1 (N15738, N15732);
not NOT1 (N15739, N15731);
xor XOR2 (N15740, N15733, N10141);
nand NAND4 (N15741, N15714, N3620, N2153, N6935);
not NOT1 (N15742, N15737);
buf BUF1 (N15743, N15735);
buf BUF1 (N15744, N15741);
and AND3 (N15745, N15725, N9090, N11955);
not NOT1 (N15746, N15738);
nor NOR2 (N15747, N15721, N2942);
nand NAND4 (N15748, N15739, N38, N994, N9664);
buf BUF1 (N15749, N15745);
and AND2 (N15750, N15736, N4376);
nor NOR2 (N15751, N15747, N6040);
buf BUF1 (N15752, N15748);
buf BUF1 (N15753, N15742);
and AND3 (N15754, N15743, N6741, N2143);
xor XOR2 (N15755, N15744, N7494);
not NOT1 (N15756, N15746);
xor XOR2 (N15757, N15754, N13211);
nor NOR3 (N15758, N15740, N12689, N15033);
nand NAND2 (N15759, N15755, N13394);
not NOT1 (N15760, N15752);
not NOT1 (N15761, N15760);
not NOT1 (N15762, N15750);
nor NOR4 (N15763, N15759, N12187, N15364, N11585);
buf BUF1 (N15764, N15757);
not NOT1 (N15765, N15749);
not NOT1 (N15766, N15762);
xor XOR2 (N15767, N15766, N9809);
nor NOR2 (N15768, N15751, N4606);
nor NOR2 (N15769, N15767, N8077);
and AND2 (N15770, N15712, N9235);
or OR4 (N15771, N15763, N3520, N2710, N9212);
nor NOR4 (N15772, N15770, N9953, N7598, N3169);
nor NOR3 (N15773, N15761, N7344, N1828);
nand NAND3 (N15774, N15772, N9193, N2138);
and AND2 (N15775, N15769, N4687);
buf BUF1 (N15776, N15775);
and AND3 (N15777, N15768, N9722, N1734);
buf BUF1 (N15778, N15777);
buf BUF1 (N15779, N15758);
not NOT1 (N15780, N15756);
xor XOR2 (N15781, N15771, N7385);
buf BUF1 (N15782, N15776);
or OR2 (N15783, N15781, N1377);
nor NOR2 (N15784, N15773, N10021);
or OR3 (N15785, N15778, N1419, N2896);
xor XOR2 (N15786, N15780, N13122);
or OR3 (N15787, N15765, N9715, N10266);
or OR3 (N15788, N15753, N14552, N5304);
nand NAND2 (N15789, N15774, N12443);
nor NOR2 (N15790, N15782, N11871);
nor NOR2 (N15791, N15785, N8010);
buf BUF1 (N15792, N15789);
or OR3 (N15793, N15783, N15022, N2891);
nand NAND2 (N15794, N15787, N1918);
buf BUF1 (N15795, N15788);
nand NAND4 (N15796, N15793, N11726, N11958, N15489);
and AND3 (N15797, N15791, N4032, N15263);
and AND2 (N15798, N15792, N3645);
nand NAND4 (N15799, N15784, N12254, N13210, N15107);
or OR4 (N15800, N15797, N6708, N11825, N5847);
and AND3 (N15801, N15795, N7276, N15399);
or OR4 (N15802, N15800, N959, N1298, N12305);
not NOT1 (N15803, N15798);
nand NAND4 (N15804, N15764, N11502, N12958, N10276);
buf BUF1 (N15805, N15801);
nor NOR2 (N15806, N15786, N13803);
nor NOR2 (N15807, N15804, N13611);
and AND4 (N15808, N15806, N12740, N1936, N500);
xor XOR2 (N15809, N15807, N7672);
buf BUF1 (N15810, N15790);
nor NOR2 (N15811, N15809, N10537);
xor XOR2 (N15812, N15779, N11666);
nor NOR4 (N15813, N15799, N6979, N13190, N15597);
and AND4 (N15814, N15794, N12322, N4352, N12388);
xor XOR2 (N15815, N15805, N7400);
nand NAND4 (N15816, N15815, N3103, N628, N6602);
nor NOR2 (N15817, N15808, N9788);
xor XOR2 (N15818, N15817, N546);
or OR4 (N15819, N15803, N12342, N2030, N3969);
and AND4 (N15820, N15818, N5664, N8332, N6366);
nor NOR3 (N15821, N15820, N7786, N14597);
xor XOR2 (N15822, N15816, N1531);
or OR3 (N15823, N15814, N11241, N12949);
nand NAND3 (N15824, N15812, N15179, N10027);
and AND3 (N15825, N15821, N6752, N4046);
not NOT1 (N15826, N15823);
not NOT1 (N15827, N15822);
xor XOR2 (N15828, N15826, N4813);
nand NAND2 (N15829, N15811, N8742);
and AND4 (N15830, N15813, N12585, N10707, N10061);
nand NAND3 (N15831, N15810, N5076, N15353);
buf BUF1 (N15832, N15827);
or OR4 (N15833, N15796, N11710, N8045, N2792);
or OR4 (N15834, N15833, N12221, N4978, N10226);
nand NAND3 (N15835, N15830, N3543, N5363);
not NOT1 (N15836, N15832);
and AND2 (N15837, N15829, N13524);
xor XOR2 (N15838, N15819, N2257);
buf BUF1 (N15839, N15835);
nand NAND4 (N15840, N15837, N13860, N1458, N9752);
nand NAND4 (N15841, N15824, N4112, N12637, N3144);
nor NOR2 (N15842, N15825, N8200);
not NOT1 (N15843, N15836);
xor XOR2 (N15844, N15841, N6268);
and AND2 (N15845, N15802, N4722);
nand NAND4 (N15846, N15842, N13931, N13153, N2949);
nand NAND3 (N15847, N15831, N14992, N6159);
and AND4 (N15848, N15834, N15060, N3695, N3335);
nand NAND4 (N15849, N15845, N5006, N13646, N5231);
nor NOR3 (N15850, N15844, N11423, N7574);
or OR2 (N15851, N15838, N13434);
xor XOR2 (N15852, N15843, N13977);
xor XOR2 (N15853, N15846, N9667);
not NOT1 (N15854, N15849);
and AND2 (N15855, N15854, N11925);
buf BUF1 (N15856, N15828);
xor XOR2 (N15857, N15840, N14838);
nand NAND2 (N15858, N15857, N8943);
buf BUF1 (N15859, N15851);
or OR4 (N15860, N15848, N10290, N2328, N5748);
or OR3 (N15861, N15847, N9539, N3791);
not NOT1 (N15862, N15856);
not NOT1 (N15863, N15858);
nand NAND2 (N15864, N15860, N15421);
not NOT1 (N15865, N15839);
nand NAND3 (N15866, N15850, N4336, N458);
nand NAND2 (N15867, N15866, N11901);
not NOT1 (N15868, N15863);
xor XOR2 (N15869, N15852, N13743);
nand NAND2 (N15870, N15855, N6268);
nor NOR4 (N15871, N15861, N1206, N4089, N3178);
nand NAND2 (N15872, N15871, N8998);
buf BUF1 (N15873, N15872);
nand NAND4 (N15874, N15873, N9307, N8117, N13035);
xor XOR2 (N15875, N15868, N5920);
xor XOR2 (N15876, N15864, N9538);
not NOT1 (N15877, N15853);
nor NOR2 (N15878, N15870, N6308);
xor XOR2 (N15879, N15878, N5671);
nand NAND4 (N15880, N15877, N13896, N4670, N10716);
or OR4 (N15881, N15869, N9947, N5913, N12463);
not NOT1 (N15882, N15876);
nand NAND4 (N15883, N15875, N2549, N10233, N2364);
nor NOR3 (N15884, N15881, N10259, N8014);
and AND4 (N15885, N15883, N9425, N10098, N11342);
nand NAND2 (N15886, N15865, N6929);
not NOT1 (N15887, N15879);
or OR2 (N15888, N15874, N14738);
nor NOR2 (N15889, N15867, N12810);
or OR4 (N15890, N15889, N5223, N10817, N11617);
not NOT1 (N15891, N15886);
nor NOR4 (N15892, N15885, N10562, N8123, N6767);
not NOT1 (N15893, N15887);
not NOT1 (N15894, N15880);
xor XOR2 (N15895, N15894, N8275);
xor XOR2 (N15896, N15882, N2924);
buf BUF1 (N15897, N15892);
not NOT1 (N15898, N15897);
not NOT1 (N15899, N15898);
buf BUF1 (N15900, N15890);
nand NAND3 (N15901, N15862, N11072, N10482);
xor XOR2 (N15902, N15900, N6183);
and AND4 (N15903, N15895, N10891, N7798, N10909);
or OR4 (N15904, N15902, N3602, N11494, N5054);
not NOT1 (N15905, N15884);
nand NAND3 (N15906, N15896, N5565, N1221);
not NOT1 (N15907, N15899);
or OR2 (N15908, N15903, N8613);
not NOT1 (N15909, N15859);
nor NOR4 (N15910, N15904, N12266, N5047, N3359);
nand NAND2 (N15911, N15901, N2463);
xor XOR2 (N15912, N15905, N3175);
nor NOR2 (N15913, N15891, N4616);
xor XOR2 (N15914, N15909, N12154);
not NOT1 (N15915, N15911);
nand NAND3 (N15916, N15888, N10360, N14626);
and AND3 (N15917, N15910, N14209, N14498);
not NOT1 (N15918, N15912);
nand NAND4 (N15919, N15918, N5261, N10482, N6036);
not NOT1 (N15920, N15914);
nand NAND3 (N15921, N15906, N12164, N7427);
nand NAND4 (N15922, N15920, N6668, N9037, N9275);
nand NAND2 (N15923, N15919, N3151);
xor XOR2 (N15924, N15913, N6065);
nor NOR3 (N15925, N15907, N4137, N8875);
nor NOR3 (N15926, N15921, N15143, N4656);
not NOT1 (N15927, N15917);
not NOT1 (N15928, N15925);
buf BUF1 (N15929, N15893);
or OR4 (N15930, N15908, N6497, N14030, N12950);
nand NAND3 (N15931, N15930, N6294, N6878);
xor XOR2 (N15932, N15931, N2209);
and AND4 (N15933, N15915, N7211, N6747, N11971);
not NOT1 (N15934, N15928);
xor XOR2 (N15935, N15929, N3571);
and AND4 (N15936, N15932, N6358, N11023, N6932);
or OR2 (N15937, N15924, N1379);
not NOT1 (N15938, N15937);
xor XOR2 (N15939, N15935, N6646);
or OR2 (N15940, N15916, N1492);
not NOT1 (N15941, N15922);
nand NAND2 (N15942, N15933, N8333);
and AND2 (N15943, N15942, N5332);
nand NAND4 (N15944, N15941, N12394, N787, N11959);
and AND4 (N15945, N15927, N4579, N13203, N15769);
not NOT1 (N15946, N15936);
buf BUF1 (N15947, N15938);
nand NAND3 (N15948, N15934, N3194, N2469);
not NOT1 (N15949, N15926);
and AND3 (N15950, N15949, N10371, N5892);
nor NOR3 (N15951, N15943, N6576, N6707);
or OR3 (N15952, N15940, N8918, N10304);
buf BUF1 (N15953, N15939);
and AND3 (N15954, N15947, N3493, N15621);
and AND3 (N15955, N15945, N5629, N2839);
not NOT1 (N15956, N15948);
nand NAND4 (N15957, N15923, N13149, N14317, N12959);
nor NOR4 (N15958, N15953, N13288, N4621, N15153);
nand NAND3 (N15959, N15946, N9916, N15818);
buf BUF1 (N15960, N15957);
and AND4 (N15961, N15944, N10320, N1666, N848);
or OR2 (N15962, N15951, N13548);
and AND3 (N15963, N15956, N49, N14773);
nand NAND3 (N15964, N15959, N13337, N1163);
xor XOR2 (N15965, N15955, N8793);
or OR3 (N15966, N15961, N11629, N6634);
not NOT1 (N15967, N15966);
not NOT1 (N15968, N15950);
buf BUF1 (N15969, N15968);
not NOT1 (N15970, N15967);
or OR2 (N15971, N15954, N5250);
or OR3 (N15972, N15958, N10866, N10095);
nand NAND2 (N15973, N15971, N7857);
buf BUF1 (N15974, N15952);
or OR4 (N15975, N15960, N228, N1079, N2061);
xor XOR2 (N15976, N15964, N14293);
xor XOR2 (N15977, N15963, N5937);
nor NOR4 (N15978, N15976, N9773, N673, N4083);
and AND3 (N15979, N15962, N13050, N6665);
buf BUF1 (N15980, N15970);
or OR3 (N15981, N15978, N5975, N4686);
or OR2 (N15982, N15973, N15839);
nand NAND4 (N15983, N15977, N3410, N2542, N11185);
nand NAND3 (N15984, N15981, N11581, N7120);
not NOT1 (N15985, N15975);
not NOT1 (N15986, N15984);
buf BUF1 (N15987, N15986);
nand NAND2 (N15988, N15965, N10807);
nand NAND3 (N15989, N15980, N9338, N8086);
nor NOR2 (N15990, N15982, N7443);
or OR4 (N15991, N15988, N11183, N12709, N12468);
nor NOR2 (N15992, N15983, N3105);
buf BUF1 (N15993, N15972);
and AND3 (N15994, N15979, N6425, N4967);
nor NOR4 (N15995, N15985, N8484, N14089, N5683);
nand NAND3 (N15996, N15989, N8107, N12107);
and AND4 (N15997, N15990, N6703, N15727, N10977);
buf BUF1 (N15998, N15987);
and AND2 (N15999, N15998, N6292);
and AND2 (N16000, N15999, N15747);
xor XOR2 (N16001, N15996, N1699);
buf BUF1 (N16002, N15992);
nand NAND2 (N16003, N16001, N10365);
not NOT1 (N16004, N15993);
nand NAND3 (N16005, N16004, N470, N12872);
buf BUF1 (N16006, N15969);
or OR3 (N16007, N15994, N1749, N12201);
xor XOR2 (N16008, N16007, N14291);
and AND4 (N16009, N16003, N12418, N7111, N11823);
nor NOR3 (N16010, N16005, N12618, N2275);
nor NOR2 (N16011, N16002, N11653);
not NOT1 (N16012, N16008);
nand NAND4 (N16013, N15997, N7178, N6866, N7970);
endmodule