// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20;

output N512,N507,N510,N494,N491,N519,N518,N502,N517,N520;

buf BUF1 (N21, N1);
buf BUF1 (N22, N3);
or OR3 (N23, N19, N19, N14);
or OR2 (N24, N11, N2);
xor XOR2 (N25, N5, N1);
or OR3 (N26, N17, N21, N20);
buf BUF1 (N27, N1);
xor XOR2 (N28, N8, N3);
and AND4 (N29, N11, N1, N27, N12);
and AND4 (N30, N9, N26, N8, N3);
not NOT1 (N31, N18);
nor NOR2 (N32, N21, N31);
xor XOR2 (N33, N15, N9);
not NOT1 (N34, N18);
xor XOR2 (N35, N34, N11);
buf BUF1 (N36, N25);
xor XOR2 (N37, N23, N32);
buf BUF1 (N38, N9);
buf BUF1 (N39, N33);
not NOT1 (N40, N38);
and AND4 (N41, N36, N16, N32, N28);
buf BUF1 (N42, N27);
nand NAND3 (N43, N29, N39, N22);
and AND3 (N44, N11, N21, N18);
buf BUF1 (N45, N27);
buf BUF1 (N46, N41);
or OR3 (N47, N46, N18, N41);
not NOT1 (N48, N40);
nand NAND3 (N49, N48, N15, N22);
nand NAND2 (N50, N24, N36);
xor XOR2 (N51, N44, N37);
buf BUF1 (N52, N51);
xor XOR2 (N53, N9, N28);
buf BUF1 (N54, N49);
buf BUF1 (N55, N35);
not NOT1 (N56, N53);
xor XOR2 (N57, N42, N22);
nand NAND3 (N58, N57, N5, N47);
and AND4 (N59, N2, N14, N27, N30);
nor NOR2 (N60, N28, N51);
xor XOR2 (N61, N50, N10);
buf BUF1 (N62, N59);
not NOT1 (N63, N60);
and AND3 (N64, N63, N61, N5);
or OR3 (N65, N25, N23, N15);
nor NOR3 (N66, N43, N41, N20);
nand NAND2 (N67, N58, N32);
and AND2 (N68, N54, N52);
not NOT1 (N69, N57);
not NOT1 (N70, N55);
nor NOR4 (N71, N64, N41, N54, N42);
xor XOR2 (N72, N45, N47);
buf BUF1 (N73, N56);
not NOT1 (N74, N66);
xor XOR2 (N75, N62, N2);
not NOT1 (N76, N68);
and AND4 (N77, N65, N49, N70, N48);
and AND2 (N78, N34, N6);
and AND2 (N79, N75, N23);
xor XOR2 (N80, N72, N10);
or OR4 (N81, N74, N6, N9, N31);
xor XOR2 (N82, N81, N60);
nand NAND3 (N83, N69, N29, N74);
not NOT1 (N84, N79);
xor XOR2 (N85, N67, N7);
nor NOR4 (N86, N85, N75, N49, N50);
and AND3 (N87, N73, N9, N7);
buf BUF1 (N88, N87);
buf BUF1 (N89, N83);
xor XOR2 (N90, N84, N46);
buf BUF1 (N91, N77);
buf BUF1 (N92, N78);
and AND4 (N93, N88, N23, N8, N76);
not NOT1 (N94, N31);
nand NAND4 (N95, N92, N82, N28, N81);
xor XOR2 (N96, N90, N29);
and AND3 (N97, N30, N43, N34);
and AND4 (N98, N89, N58, N32, N15);
nor NOR2 (N99, N93, N47);
buf BUF1 (N100, N80);
xor XOR2 (N101, N96, N70);
nand NAND2 (N102, N101, N59);
and AND4 (N103, N86, N82, N69, N97);
or OR4 (N104, N32, N63, N97, N41);
nor NOR2 (N105, N71, N76);
xor XOR2 (N106, N94, N55);
not NOT1 (N107, N104);
buf BUF1 (N108, N106);
or OR3 (N109, N100, N106, N58);
not NOT1 (N110, N103);
not NOT1 (N111, N99);
and AND2 (N112, N105, N82);
nand NAND4 (N113, N98, N104, N88, N92);
buf BUF1 (N114, N112);
not NOT1 (N115, N107);
and AND3 (N116, N102, N8, N106);
not NOT1 (N117, N111);
not NOT1 (N118, N116);
or OR4 (N119, N115, N7, N44, N75);
and AND3 (N120, N95, N39, N94);
not NOT1 (N121, N110);
nand NAND2 (N122, N120, N33);
not NOT1 (N123, N117);
nor NOR2 (N124, N122, N75);
buf BUF1 (N125, N118);
nor NOR2 (N126, N124, N50);
xor XOR2 (N127, N108, N94);
xor XOR2 (N128, N125, N23);
nor NOR3 (N129, N121, N22, N43);
buf BUF1 (N130, N109);
nand NAND3 (N131, N129, N69, N95);
buf BUF1 (N132, N113);
buf BUF1 (N133, N126);
nor NOR3 (N134, N127, N37, N91);
nor NOR4 (N135, N113, N45, N75, N37);
xor XOR2 (N136, N132, N132);
nor NOR2 (N137, N119, N112);
buf BUF1 (N138, N134);
nor NOR3 (N139, N135, N108, N10);
or OR3 (N140, N114, N84, N88);
nand NAND3 (N141, N137, N123, N133);
nor NOR2 (N142, N19, N106);
not NOT1 (N143, N79);
nand NAND4 (N144, N128, N98, N69, N90);
or OR3 (N145, N130, N143, N100);
xor XOR2 (N146, N61, N94);
buf BUF1 (N147, N140);
xor XOR2 (N148, N142, N122);
nor NOR4 (N149, N139, N68, N10, N44);
or OR3 (N150, N138, N145, N126);
or OR3 (N151, N54, N35, N81);
buf BUF1 (N152, N146);
nand NAND3 (N153, N149, N126, N138);
nor NOR4 (N154, N144, N28, N146, N53);
and AND4 (N155, N141, N81, N108, N118);
buf BUF1 (N156, N151);
nor NOR2 (N157, N156, N147);
xor XOR2 (N158, N42, N148);
or OR2 (N159, N30, N80);
nand NAND4 (N160, N131, N140, N9, N17);
nand NAND2 (N161, N155, N94);
nand NAND3 (N162, N157, N7, N123);
xor XOR2 (N163, N154, N43);
not NOT1 (N164, N163);
not NOT1 (N165, N160);
xor XOR2 (N166, N152, N108);
nor NOR2 (N167, N162, N135);
buf BUF1 (N168, N136);
and AND4 (N169, N150, N121, N52, N116);
buf BUF1 (N170, N164);
and AND4 (N171, N165, N59, N116, N129);
and AND4 (N172, N153, N106, N162, N18);
xor XOR2 (N173, N166, N52);
and AND4 (N174, N161, N105, N38, N93);
or OR3 (N175, N158, N9, N3);
nor NOR3 (N176, N169, N47, N152);
or OR4 (N177, N168, N13, N64, N36);
buf BUF1 (N178, N167);
or OR3 (N179, N159, N83, N127);
xor XOR2 (N180, N173, N76);
nand NAND3 (N181, N178, N6, N35);
buf BUF1 (N182, N177);
nand NAND3 (N183, N175, N56, N133);
buf BUF1 (N184, N179);
not NOT1 (N185, N174);
and AND2 (N186, N185, N167);
nand NAND2 (N187, N183, N11);
not NOT1 (N188, N180);
nor NOR3 (N189, N181, N166, N166);
nand NAND3 (N190, N184, N68, N101);
and AND3 (N191, N186, N186, N18);
xor XOR2 (N192, N190, N28);
and AND2 (N193, N170, N25);
and AND2 (N194, N187, N34);
and AND3 (N195, N192, N78, N69);
nor NOR2 (N196, N176, N191);
and AND4 (N197, N96, N154, N38, N71);
xor XOR2 (N198, N171, N112);
not NOT1 (N199, N197);
and AND2 (N200, N195, N115);
not NOT1 (N201, N188);
not NOT1 (N202, N194);
nor NOR2 (N203, N198, N120);
or OR3 (N204, N200, N166, N120);
buf BUF1 (N205, N202);
xor XOR2 (N206, N205, N61);
and AND3 (N207, N204, N62, N152);
nand NAND3 (N208, N199, N38, N104);
xor XOR2 (N209, N172, N198);
nand NAND2 (N210, N207, N27);
buf BUF1 (N211, N206);
nand NAND4 (N212, N201, N66, N137, N161);
xor XOR2 (N213, N209, N128);
or OR2 (N214, N208, N184);
buf BUF1 (N215, N210);
nor NOR3 (N216, N203, N142, N39);
or OR2 (N217, N193, N128);
not NOT1 (N218, N214);
xor XOR2 (N219, N213, N188);
xor XOR2 (N220, N215, N119);
nor NOR2 (N221, N219, N24);
or OR3 (N222, N216, N27, N90);
nor NOR4 (N223, N220, N132, N94, N149);
or OR2 (N224, N211, N100);
not NOT1 (N225, N196);
or OR2 (N226, N212, N209);
xor XOR2 (N227, N224, N82);
and AND4 (N228, N222, N92, N107, N129);
nor NOR3 (N229, N226, N209, N167);
or OR2 (N230, N189, N83);
xor XOR2 (N231, N229, N36);
buf BUF1 (N232, N221);
and AND3 (N233, N218, N32, N144);
buf BUF1 (N234, N230);
and AND3 (N235, N223, N161, N47);
nor NOR4 (N236, N182, N16, N222, N211);
or OR2 (N237, N233, N204);
and AND4 (N238, N235, N184, N149, N29);
not NOT1 (N239, N231);
not NOT1 (N240, N234);
nand NAND2 (N241, N236, N135);
not NOT1 (N242, N238);
not NOT1 (N243, N225);
or OR3 (N244, N237, N52, N131);
nand NAND2 (N245, N232, N54);
or OR3 (N246, N239, N230, N8);
or OR4 (N247, N246, N192, N105, N126);
nor NOR3 (N248, N244, N122, N186);
or OR4 (N249, N245, N168, N38, N223);
nand NAND4 (N250, N249, N150, N177, N130);
xor XOR2 (N251, N240, N11);
or OR4 (N252, N217, N63, N104, N94);
nor NOR4 (N253, N241, N114, N230, N54);
and AND2 (N254, N242, N29);
not NOT1 (N255, N250);
xor XOR2 (N256, N228, N197);
and AND4 (N257, N227, N171, N42, N51);
not NOT1 (N258, N252);
and AND2 (N259, N255, N192);
nand NAND4 (N260, N247, N54, N212, N105);
not NOT1 (N261, N253);
nand NAND2 (N262, N248, N26);
and AND2 (N263, N257, N256);
and AND2 (N264, N258, N152);
buf BUF1 (N265, N150);
xor XOR2 (N266, N259, N191);
xor XOR2 (N267, N265, N257);
not NOT1 (N268, N266);
nand NAND4 (N269, N254, N106, N16, N134);
not NOT1 (N270, N251);
or OR2 (N271, N264, N181);
xor XOR2 (N272, N269, N138);
nand NAND4 (N273, N268, N265, N25, N172);
nor NOR2 (N274, N263, N196);
and AND4 (N275, N261, N103, N37, N68);
nor NOR2 (N276, N274, N221);
buf BUF1 (N277, N276);
nand NAND4 (N278, N262, N104, N232, N156);
and AND4 (N279, N267, N15, N176, N129);
and AND3 (N280, N273, N127, N233);
nand NAND3 (N281, N270, N17, N67);
buf BUF1 (N282, N272);
buf BUF1 (N283, N281);
nor NOR2 (N284, N275, N218);
and AND4 (N285, N260, N77, N41, N261);
nor NOR2 (N286, N278, N109);
not NOT1 (N287, N279);
and AND3 (N288, N284, N248, N64);
xor XOR2 (N289, N288, N131);
nand NAND2 (N290, N287, N104);
buf BUF1 (N291, N282);
or OR3 (N292, N291, N141, N58);
and AND3 (N293, N286, N289, N62);
nand NAND3 (N294, N139, N202, N260);
nor NOR4 (N295, N283, N165, N90, N104);
nor NOR2 (N296, N271, N81);
xor XOR2 (N297, N280, N280);
xor XOR2 (N298, N243, N226);
nor NOR3 (N299, N296, N189, N277);
xor XOR2 (N300, N36, N99);
nand NAND4 (N301, N285, N140, N149, N46);
not NOT1 (N302, N297);
buf BUF1 (N303, N302);
nor NOR3 (N304, N295, N159, N158);
buf BUF1 (N305, N299);
not NOT1 (N306, N293);
nor NOR3 (N307, N303, N128, N93);
or OR3 (N308, N301, N65, N265);
not NOT1 (N309, N305);
buf BUF1 (N310, N300);
or OR4 (N311, N290, N214, N308, N128);
nor NOR4 (N312, N163, N184, N131, N154);
nor NOR2 (N313, N312, N269);
not NOT1 (N314, N292);
not NOT1 (N315, N298);
or OR4 (N316, N306, N204, N86, N276);
nor NOR3 (N317, N309, N59, N217);
nor NOR2 (N318, N315, N34);
or OR2 (N319, N313, N227);
and AND4 (N320, N310, N4, N217, N252);
nand NAND2 (N321, N307, N300);
and AND4 (N322, N294, N11, N232, N159);
nand NAND2 (N323, N321, N144);
or OR3 (N324, N320, N241, N108);
not NOT1 (N325, N318);
or OR2 (N326, N319, N104);
nand NAND4 (N327, N316, N161, N322, N86);
or OR4 (N328, N248, N199, N158, N52);
and AND3 (N329, N323, N180, N104);
xor XOR2 (N330, N328, N58);
nand NAND4 (N331, N324, N157, N25, N46);
nor NOR3 (N332, N325, N22, N84);
or OR2 (N333, N326, N153);
nor NOR3 (N334, N329, N124, N214);
buf BUF1 (N335, N314);
nor NOR2 (N336, N335, N230);
nor NOR3 (N337, N331, N41, N76);
not NOT1 (N338, N327);
nand NAND2 (N339, N332, N21);
buf BUF1 (N340, N339);
or OR3 (N341, N340, N16, N20);
or OR2 (N342, N341, N196);
or OR4 (N343, N337, N94, N33, N5);
xor XOR2 (N344, N330, N223);
buf BUF1 (N345, N338);
not NOT1 (N346, N333);
nor NOR4 (N347, N336, N306, N251, N215);
or OR2 (N348, N304, N341);
buf BUF1 (N349, N317);
nor NOR3 (N350, N342, N299, N184);
or OR3 (N351, N346, N325, N39);
or OR2 (N352, N349, N150);
nand NAND3 (N353, N347, N324, N56);
or OR2 (N354, N351, N220);
or OR2 (N355, N311, N302);
nor NOR3 (N356, N352, N317, N146);
buf BUF1 (N357, N355);
xor XOR2 (N358, N353, N1);
buf BUF1 (N359, N357);
nand NAND4 (N360, N343, N205, N182, N3);
and AND4 (N361, N348, N103, N51, N242);
buf BUF1 (N362, N360);
and AND4 (N363, N345, N94, N124, N206);
nor NOR3 (N364, N350, N121, N80);
or OR2 (N365, N354, N114);
xor XOR2 (N366, N365, N359);
buf BUF1 (N367, N118);
or OR4 (N368, N344, N285, N116, N357);
nand NAND4 (N369, N358, N126, N144, N32);
nand NAND2 (N370, N334, N287);
xor XOR2 (N371, N356, N237);
not NOT1 (N372, N362);
and AND3 (N373, N369, N163, N105);
and AND2 (N374, N366, N94);
and AND2 (N375, N373, N297);
nand NAND2 (N376, N363, N185);
not NOT1 (N377, N367);
nand NAND2 (N378, N376, N178);
buf BUF1 (N379, N372);
nand NAND2 (N380, N379, N256);
and AND4 (N381, N371, N140, N302, N317);
nor NOR3 (N382, N374, N106, N72);
not NOT1 (N383, N381);
and AND3 (N384, N377, N81, N95);
xor XOR2 (N385, N383, N87);
nor NOR2 (N386, N364, N317);
and AND4 (N387, N382, N249, N5, N169);
xor XOR2 (N388, N386, N120);
and AND2 (N389, N370, N268);
xor XOR2 (N390, N375, N295);
not NOT1 (N391, N387);
nor NOR2 (N392, N368, N350);
and AND3 (N393, N378, N83, N42);
not NOT1 (N394, N393);
nand NAND2 (N395, N390, N354);
xor XOR2 (N396, N380, N91);
nand NAND2 (N397, N396, N51);
xor XOR2 (N398, N361, N255);
nand NAND2 (N399, N388, N62);
nor NOR4 (N400, N398, N16, N182, N159);
and AND4 (N401, N400, N140, N84, N355);
not NOT1 (N402, N391);
xor XOR2 (N403, N384, N125);
nand NAND4 (N404, N402, N188, N242, N319);
nor NOR3 (N405, N392, N395, N47);
and AND3 (N406, N63, N88, N196);
buf BUF1 (N407, N404);
and AND3 (N408, N385, N117, N283);
xor XOR2 (N409, N389, N340);
buf BUF1 (N410, N399);
buf BUF1 (N411, N403);
not NOT1 (N412, N401);
nand NAND2 (N413, N405, N148);
buf BUF1 (N414, N410);
and AND4 (N415, N413, N61, N137, N402);
xor XOR2 (N416, N411, N371);
and AND2 (N417, N407, N153);
or OR2 (N418, N417, N161);
nand NAND4 (N419, N394, N85, N243, N415);
buf BUF1 (N420, N137);
and AND2 (N421, N409, N381);
buf BUF1 (N422, N397);
nor NOR4 (N423, N420, N326, N266, N280);
or OR2 (N424, N423, N214);
nor NOR2 (N425, N416, N67);
buf BUF1 (N426, N424);
and AND3 (N427, N418, N342, N54);
buf BUF1 (N428, N426);
buf BUF1 (N429, N406);
nand NAND2 (N430, N408, N160);
nand NAND3 (N431, N425, N394, N4);
or OR3 (N432, N428, N83, N240);
not NOT1 (N433, N419);
nand NAND3 (N434, N432, N193, N382);
nand NAND4 (N435, N431, N189, N111, N274);
or OR4 (N436, N429, N113, N12, N318);
not NOT1 (N437, N421);
nor NOR3 (N438, N414, N374, N53);
nand NAND4 (N439, N438, N1, N280, N407);
or OR4 (N440, N439, N398, N400, N344);
or OR2 (N441, N412, N372);
or OR3 (N442, N430, N167, N405);
or OR2 (N443, N427, N140);
not NOT1 (N444, N433);
nor NOR4 (N445, N435, N315, N70, N428);
xor XOR2 (N446, N442, N325);
nor NOR4 (N447, N436, N169, N124, N348);
or OR4 (N448, N446, N224, N301, N371);
buf BUF1 (N449, N441);
buf BUF1 (N450, N445);
and AND2 (N451, N440, N256);
xor XOR2 (N452, N448, N425);
and AND3 (N453, N451, N210, N85);
not NOT1 (N454, N422);
xor XOR2 (N455, N447, N2);
xor XOR2 (N456, N450, N202);
nand NAND3 (N457, N454, N227, N444);
buf BUF1 (N458, N46);
not NOT1 (N459, N443);
or OR4 (N460, N459, N324, N446, N114);
or OR2 (N461, N434, N198);
not NOT1 (N462, N437);
buf BUF1 (N463, N453);
and AND4 (N464, N458, N98, N1, N4);
or OR3 (N465, N452, N423, N132);
and AND2 (N466, N464, N361);
buf BUF1 (N467, N465);
nand NAND3 (N468, N460, N89, N404);
and AND4 (N469, N463, N413, N455, N384);
nand NAND3 (N470, N416, N89, N57);
not NOT1 (N471, N461);
nor NOR2 (N472, N466, N244);
and AND4 (N473, N449, N122, N109, N156);
nand NAND3 (N474, N472, N403, N227);
nand NAND3 (N475, N467, N160, N134);
buf BUF1 (N476, N462);
xor XOR2 (N477, N468, N52);
xor XOR2 (N478, N474, N346);
not NOT1 (N479, N475);
xor XOR2 (N480, N478, N303);
and AND3 (N481, N471, N472, N84);
xor XOR2 (N482, N456, N347);
nand NAND3 (N483, N470, N180, N456);
nor NOR3 (N484, N483, N251, N449);
or OR4 (N485, N484, N145, N279, N338);
buf BUF1 (N486, N485);
xor XOR2 (N487, N476, N428);
not NOT1 (N488, N487);
buf BUF1 (N489, N457);
buf BUF1 (N490, N480);
or OR2 (N491, N490, N353);
nand NAND4 (N492, N469, N367, N481, N477);
nand NAND3 (N493, N339, N60, N366);
nor NOR4 (N494, N22, N312, N398, N400);
not NOT1 (N495, N482);
not NOT1 (N496, N489);
not NOT1 (N497, N488);
or OR3 (N498, N495, N218, N287);
nand NAND3 (N499, N493, N293, N206);
xor XOR2 (N500, N498, N68);
not NOT1 (N501, N486);
buf BUF1 (N502, N499);
nor NOR3 (N503, N492, N12, N360);
not NOT1 (N504, N503);
and AND3 (N505, N479, N349, N58);
xor XOR2 (N506, N504, N19);
not NOT1 (N507, N497);
nand NAND4 (N508, N505, N34, N337, N341);
and AND3 (N509, N506, N336, N3);
not NOT1 (N510, N508);
and AND4 (N511, N473, N420, N269, N35);
nand NAND2 (N512, N496, N324);
buf BUF1 (N513, N500);
xor XOR2 (N514, N511, N18);
buf BUF1 (N515, N509);
or OR4 (N516, N514, N460, N389, N100);
buf BUF1 (N517, N513);
or OR3 (N518, N515, N393, N41);
nand NAND4 (N519, N516, N439, N312, N342);
xor XOR2 (N520, N501, N298);
endmodule