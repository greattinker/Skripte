// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23;

output N313,N311,N317,N315,N301,N318,N321,N322,N319,N323;

nand NAND4 (N24, N11, N22, N16, N16);
xor XOR2 (N25, N7, N24);
nor NOR2 (N26, N24, N23);
or OR3 (N27, N18, N13, N16);
or OR4 (N28, N12, N1, N14, N10);
buf BUF1 (N29, N17);
xor XOR2 (N30, N19, N16);
xor XOR2 (N31, N16, N4);
or OR2 (N32, N16, N15);
nand NAND3 (N33, N8, N30, N11);
or OR2 (N34, N28, N22);
xor XOR2 (N35, N4, N21);
nand NAND4 (N36, N22, N9, N4, N2);
buf BUF1 (N37, N27);
not NOT1 (N38, N34);
buf BUF1 (N39, N26);
and AND4 (N40, N33, N29, N22, N2);
xor XOR2 (N41, N21, N6);
and AND2 (N42, N35, N17);
and AND3 (N43, N41, N3, N6);
buf BUF1 (N44, N40);
nand NAND4 (N45, N31, N6, N17, N4);
nand NAND4 (N46, N32, N17, N11, N38);
or OR2 (N47, N39, N3);
not NOT1 (N48, N38);
xor XOR2 (N49, N25, N31);
nand NAND3 (N50, N36, N46, N21);
and AND2 (N51, N18, N16);
not NOT1 (N52, N43);
and AND3 (N53, N47, N42, N39);
or OR3 (N54, N20, N12, N18);
nand NAND2 (N55, N52, N48);
and AND4 (N56, N12, N32, N2, N39);
not NOT1 (N57, N37);
and AND4 (N58, N55, N2, N46, N14);
not NOT1 (N59, N57);
or OR3 (N60, N54, N8, N54);
nand NAND2 (N61, N58, N25);
and AND4 (N62, N56, N29, N33, N20);
nand NAND4 (N63, N51, N3, N17, N27);
nor NOR3 (N64, N61, N27, N15);
or OR3 (N65, N50, N20, N35);
and AND2 (N66, N65, N10);
nand NAND3 (N67, N63, N36, N40);
nand NAND2 (N68, N62, N29);
buf BUF1 (N69, N60);
nor NOR3 (N70, N45, N12, N55);
and AND2 (N71, N70, N36);
buf BUF1 (N72, N53);
not NOT1 (N73, N68);
nand NAND4 (N74, N49, N24, N30, N6);
not NOT1 (N75, N44);
buf BUF1 (N76, N64);
xor XOR2 (N77, N73, N49);
not NOT1 (N78, N76);
and AND2 (N79, N78, N49);
and AND4 (N80, N69, N29, N28, N46);
buf BUF1 (N81, N71);
nand NAND2 (N82, N72, N27);
xor XOR2 (N83, N59, N47);
or OR2 (N84, N67, N38);
and AND4 (N85, N74, N82, N62, N17);
and AND3 (N86, N34, N7, N58);
and AND3 (N87, N79, N75, N15);
and AND3 (N88, N43, N24, N36);
buf BUF1 (N89, N66);
nand NAND4 (N90, N84, N65, N39, N26);
nand NAND2 (N91, N83, N75);
not NOT1 (N92, N81);
buf BUF1 (N93, N77);
xor XOR2 (N94, N90, N14);
buf BUF1 (N95, N80);
and AND4 (N96, N95, N81, N72, N63);
not NOT1 (N97, N85);
not NOT1 (N98, N86);
xor XOR2 (N99, N91, N49);
buf BUF1 (N100, N92);
nor NOR3 (N101, N88, N23, N60);
and AND2 (N102, N100, N35);
xor XOR2 (N103, N97, N45);
and AND2 (N104, N98, N2);
buf BUF1 (N105, N102);
nand NAND4 (N106, N89, N4, N69, N54);
xor XOR2 (N107, N104, N38);
and AND4 (N108, N107, N80, N83, N77);
nor NOR2 (N109, N96, N60);
or OR4 (N110, N93, N6, N61, N7);
buf BUF1 (N111, N101);
xor XOR2 (N112, N99, N58);
nand NAND4 (N113, N87, N31, N98, N67);
and AND2 (N114, N108, N6);
not NOT1 (N115, N109);
nor NOR4 (N116, N110, N23, N81, N16);
and AND3 (N117, N114, N100, N76);
buf BUF1 (N118, N113);
buf BUF1 (N119, N112);
nand NAND3 (N120, N119, N117, N48);
and AND2 (N121, N85, N68);
xor XOR2 (N122, N105, N90);
and AND4 (N123, N106, N83, N82, N41);
or OR3 (N124, N121, N8, N56);
not NOT1 (N125, N94);
not NOT1 (N126, N116);
and AND3 (N127, N118, N69, N22);
not NOT1 (N128, N111);
or OR2 (N129, N125, N113);
xor XOR2 (N130, N115, N42);
xor XOR2 (N131, N103, N51);
nor NOR4 (N132, N129, N80, N8, N18);
or OR4 (N133, N132, N13, N121, N70);
nor NOR2 (N134, N122, N93);
nand NAND2 (N135, N130, N112);
nand NAND4 (N136, N123, N121, N129, N14);
and AND2 (N137, N124, N69);
xor XOR2 (N138, N127, N96);
nand NAND3 (N139, N126, N60, N72);
or OR2 (N140, N139, N38);
nand NAND4 (N141, N137, N35, N75, N37);
nand NAND2 (N142, N133, N107);
nand NAND3 (N143, N135, N4, N28);
nor NOR3 (N144, N141, N109, N126);
and AND2 (N145, N136, N37);
xor XOR2 (N146, N144, N64);
and AND4 (N147, N134, N133, N50, N26);
and AND2 (N148, N128, N96);
or OR3 (N149, N140, N7, N70);
or OR3 (N150, N142, N48, N77);
xor XOR2 (N151, N148, N72);
not NOT1 (N152, N120);
nand NAND3 (N153, N150, N99, N43);
xor XOR2 (N154, N151, N146);
and AND3 (N155, N8, N88, N17);
nand NAND2 (N156, N145, N86);
and AND4 (N157, N152, N143, N41, N56);
nand NAND2 (N158, N76, N28);
nand NAND4 (N159, N155, N108, N109, N56);
not NOT1 (N160, N156);
nand NAND2 (N161, N154, N25);
not NOT1 (N162, N158);
xor XOR2 (N163, N149, N17);
xor XOR2 (N164, N131, N156);
xor XOR2 (N165, N153, N24);
xor XOR2 (N166, N163, N51);
or OR2 (N167, N161, N44);
and AND4 (N168, N165, N69, N156, N47);
not NOT1 (N169, N138);
not NOT1 (N170, N166);
nor NOR4 (N171, N159, N145, N83, N111);
not NOT1 (N172, N170);
nand NAND4 (N173, N164, N113, N143, N95);
or OR3 (N174, N169, N30, N22);
or OR4 (N175, N160, N7, N174, N49);
xor XOR2 (N176, N15, N109);
buf BUF1 (N177, N157);
or OR2 (N178, N171, N35);
nor NOR4 (N179, N168, N29, N57, N136);
buf BUF1 (N180, N178);
xor XOR2 (N181, N167, N21);
nor NOR4 (N182, N173, N7, N53, N167);
buf BUF1 (N183, N177);
nor NOR2 (N184, N179, N81);
and AND2 (N185, N172, N62);
buf BUF1 (N186, N147);
xor XOR2 (N187, N176, N163);
nor NOR3 (N188, N182, N50, N181);
nand NAND3 (N189, N8, N16, N13);
not NOT1 (N190, N186);
xor XOR2 (N191, N183, N57);
buf BUF1 (N192, N175);
nand NAND3 (N193, N190, N160, N135);
nor NOR4 (N194, N188, N189, N102, N184);
buf BUF1 (N195, N30);
not NOT1 (N196, N160);
nand NAND4 (N197, N191, N165, N82, N189);
and AND2 (N198, N197, N124);
not NOT1 (N199, N192);
nor NOR3 (N200, N199, N25, N184);
nor NOR2 (N201, N198, N187);
nand NAND3 (N202, N50, N159, N175);
nand NAND2 (N203, N193, N137);
nand NAND2 (N204, N200, N144);
nor NOR4 (N205, N204, N59, N105, N85);
and AND2 (N206, N196, N95);
nand NAND3 (N207, N202, N156, N36);
or OR3 (N208, N162, N17, N115);
nor NOR2 (N209, N208, N138);
not NOT1 (N210, N195);
not NOT1 (N211, N205);
nor NOR3 (N212, N211, N66, N150);
not NOT1 (N213, N210);
or OR4 (N214, N203, N182, N176, N112);
nor NOR3 (N215, N194, N69, N175);
or OR3 (N216, N213, N24, N208);
buf BUF1 (N217, N209);
or OR3 (N218, N215, N26, N129);
nor NOR3 (N219, N217, N151, N63);
and AND4 (N220, N216, N52, N76, N187);
nand NAND3 (N221, N218, N177, N41);
nor NOR4 (N222, N219, N155, N36, N5);
and AND4 (N223, N220, N56, N66, N193);
or OR2 (N224, N206, N46);
and AND3 (N225, N212, N79, N40);
and AND4 (N226, N214, N35, N67, N186);
and AND2 (N227, N222, N131);
nand NAND2 (N228, N185, N54);
buf BUF1 (N229, N226);
nand NAND2 (N230, N224, N91);
nand NAND2 (N231, N225, N204);
or OR4 (N232, N228, N156, N34, N156);
and AND3 (N233, N223, N44, N107);
or OR3 (N234, N207, N112, N134);
nor NOR4 (N235, N229, N26, N225, N77);
nor NOR3 (N236, N233, N189, N168);
buf BUF1 (N237, N234);
or OR4 (N238, N237, N103, N209, N6);
nor NOR3 (N239, N180, N112, N27);
or OR2 (N240, N201, N51);
nand NAND2 (N241, N240, N227);
or OR4 (N242, N232, N17, N104, N232);
xor XOR2 (N243, N219, N95);
buf BUF1 (N244, N221);
and AND4 (N245, N231, N120, N33, N60);
or OR4 (N246, N245, N113, N119, N109);
nand NAND2 (N247, N244, N91);
buf BUF1 (N248, N247);
xor XOR2 (N249, N242, N49);
xor XOR2 (N250, N241, N96);
and AND2 (N251, N249, N182);
and AND2 (N252, N239, N178);
not NOT1 (N253, N243);
xor XOR2 (N254, N236, N195);
and AND4 (N255, N238, N198, N212, N192);
nor NOR2 (N256, N250, N174);
nor NOR3 (N257, N253, N171, N139);
buf BUF1 (N258, N256);
nand NAND2 (N259, N255, N221);
nand NAND3 (N260, N248, N37, N14);
nor NOR2 (N261, N257, N25);
and AND3 (N262, N259, N33, N81);
nor NOR2 (N263, N258, N193);
not NOT1 (N264, N251);
not NOT1 (N265, N261);
xor XOR2 (N266, N263, N166);
nor NOR3 (N267, N246, N26, N60);
buf BUF1 (N268, N265);
and AND2 (N269, N268, N14);
nand NAND3 (N270, N254, N156, N48);
nor NOR2 (N271, N262, N94);
or OR3 (N272, N267, N55, N250);
not NOT1 (N273, N271);
nor NOR2 (N274, N269, N239);
xor XOR2 (N275, N264, N235);
nand NAND2 (N276, N31, N168);
nand NAND2 (N277, N270, N56);
or OR2 (N278, N273, N74);
xor XOR2 (N279, N230, N41);
nand NAND2 (N280, N278, N165);
nand NAND3 (N281, N272, N128, N97);
or OR3 (N282, N280, N209, N161);
not NOT1 (N283, N281);
or OR3 (N284, N266, N265, N238);
and AND3 (N285, N277, N121, N272);
or OR4 (N286, N282, N89, N271, N119);
nor NOR3 (N287, N274, N117, N196);
nand NAND3 (N288, N260, N264, N184);
buf BUF1 (N289, N286);
buf BUF1 (N290, N288);
nor NOR2 (N291, N275, N286);
and AND3 (N292, N287, N20, N92);
not NOT1 (N293, N285);
xor XOR2 (N294, N252, N221);
not NOT1 (N295, N291);
not NOT1 (N296, N284);
nand NAND2 (N297, N296, N186);
not NOT1 (N298, N293);
nor NOR2 (N299, N289, N66);
xor XOR2 (N300, N292, N77);
or OR2 (N301, N299, N274);
nand NAND4 (N302, N294, N140, N182, N115);
nor NOR4 (N303, N302, N77, N276, N32);
xor XOR2 (N304, N43, N78);
xor XOR2 (N305, N298, N63);
or OR4 (N306, N305, N91, N128, N151);
xor XOR2 (N307, N283, N203);
nand NAND2 (N308, N295, N133);
nor NOR4 (N309, N279, N273, N202, N12);
nand NAND3 (N310, N290, N115, N249);
nor NOR3 (N311, N307, N53, N201);
nor NOR2 (N312, N303, N216);
or OR2 (N313, N308, N198);
nor NOR2 (N314, N309, N157);
nand NAND4 (N315, N297, N24, N295, N203);
xor XOR2 (N316, N304, N116);
or OR3 (N317, N314, N184, N223);
buf BUF1 (N318, N306);
buf BUF1 (N319, N310);
and AND2 (N320, N312, N151);
or OR2 (N321, N320, N217);
nor NOR3 (N322, N316, N167, N214);
buf BUF1 (N323, N300);
endmodule