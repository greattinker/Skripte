// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16;

output N16014,N16005,N16012,N16009,N15981,N16011,N16013,N16006,N16015,N16016;

nor NOR2 (N17, N7, N16);
xor XOR2 (N18, N10, N7);
buf BUF1 (N19, N16);
and AND2 (N20, N13, N6);
nor NOR2 (N21, N1, N7);
nor NOR2 (N22, N8, N9);
and AND4 (N23, N19, N5, N9, N19);
and AND2 (N24, N18, N4);
xor XOR2 (N25, N5, N8);
and AND4 (N26, N19, N22, N24, N15);
not NOT1 (N27, N6);
nor NOR4 (N28, N8, N12, N20, N20);
nor NOR3 (N29, N4, N22, N25);
and AND4 (N30, N25, N11, N20, N13);
nor NOR3 (N31, N24, N26, N6);
xor XOR2 (N32, N15, N18);
nor NOR2 (N33, N23, N10);
buf BUF1 (N34, N13);
not NOT1 (N35, N30);
xor XOR2 (N36, N33, N21);
buf BUF1 (N37, N10);
or OR3 (N38, N31, N23, N6);
nor NOR2 (N39, N35, N3);
and AND4 (N40, N27, N5, N16, N35);
and AND4 (N41, N39, N7, N39, N17);
not NOT1 (N42, N24);
not NOT1 (N43, N41);
xor XOR2 (N44, N37, N31);
or OR3 (N45, N43, N34, N39);
not NOT1 (N46, N7);
or OR4 (N47, N45, N28, N13, N46);
and AND3 (N48, N39, N5, N25);
nor NOR2 (N49, N24, N33);
or OR4 (N50, N44, N46, N1, N35);
nand NAND3 (N51, N38, N26, N38);
and AND4 (N52, N42, N35, N23, N26);
nor NOR3 (N53, N29, N35, N38);
not NOT1 (N54, N49);
and AND3 (N55, N32, N46, N38);
xor XOR2 (N56, N47, N2);
and AND2 (N57, N52, N1);
xor XOR2 (N58, N50, N5);
and AND2 (N59, N58, N51);
xor XOR2 (N60, N13, N20);
buf BUF1 (N61, N60);
not NOT1 (N62, N40);
nor NOR2 (N63, N48, N33);
not NOT1 (N64, N57);
not NOT1 (N65, N56);
and AND3 (N66, N62, N33, N31);
buf BUF1 (N67, N64);
not NOT1 (N68, N63);
buf BUF1 (N69, N54);
nand NAND2 (N70, N65, N61);
not NOT1 (N71, N16);
nor NOR2 (N72, N66, N26);
nor NOR4 (N73, N36, N9, N37, N42);
not NOT1 (N74, N73);
not NOT1 (N75, N70);
nand NAND2 (N76, N72, N72);
xor XOR2 (N77, N53, N9);
or OR2 (N78, N77, N64);
nand NAND4 (N79, N59, N54, N29, N10);
nor NOR4 (N80, N75, N10, N31, N69);
and AND2 (N81, N32, N21);
nand NAND3 (N82, N67, N19, N64);
buf BUF1 (N83, N81);
nor NOR2 (N84, N71, N1);
xor XOR2 (N85, N78, N25);
nand NAND2 (N86, N79, N11);
not NOT1 (N87, N83);
and AND3 (N88, N87, N76, N22);
and AND3 (N89, N9, N51, N44);
nand NAND2 (N90, N88, N3);
nand NAND3 (N91, N90, N19, N64);
buf BUF1 (N92, N86);
xor XOR2 (N93, N74, N7);
and AND4 (N94, N84, N54, N81, N47);
or OR2 (N95, N92, N59);
not NOT1 (N96, N85);
not NOT1 (N97, N80);
nand NAND2 (N98, N68, N95);
or OR4 (N99, N88, N61, N77, N2);
or OR3 (N100, N99, N20, N63);
not NOT1 (N101, N93);
and AND2 (N102, N101, N57);
nand NAND3 (N103, N98, N65, N36);
and AND4 (N104, N103, N90, N32, N38);
not NOT1 (N105, N104);
not NOT1 (N106, N94);
nand NAND2 (N107, N55, N63);
xor XOR2 (N108, N102, N65);
and AND4 (N109, N82, N53, N10, N7);
buf BUF1 (N110, N107);
nand NAND3 (N111, N108, N67, N28);
and AND4 (N112, N96, N6, N26, N67);
or OR3 (N113, N89, N43, N34);
and AND3 (N114, N113, N72, N89);
not NOT1 (N115, N110);
nand NAND3 (N116, N112, N86, N109);
nand NAND2 (N117, N13, N28);
or OR4 (N118, N111, N18, N82, N5);
not NOT1 (N119, N116);
buf BUF1 (N120, N105);
not NOT1 (N121, N117);
nor NOR2 (N122, N114, N115);
not NOT1 (N123, N19);
xor XOR2 (N124, N91, N88);
and AND3 (N125, N119, N65, N111);
or OR2 (N126, N120, N15);
nand NAND2 (N127, N125, N82);
xor XOR2 (N128, N106, N29);
and AND3 (N129, N126, N99, N88);
buf BUF1 (N130, N121);
or OR4 (N131, N127, N80, N20, N43);
and AND2 (N132, N131, N12);
buf BUF1 (N133, N100);
and AND4 (N134, N124, N116, N39, N34);
xor XOR2 (N135, N129, N74);
or OR2 (N136, N135, N58);
and AND2 (N137, N118, N131);
nor NOR4 (N138, N137, N33, N23, N93);
xor XOR2 (N139, N138, N120);
nor NOR3 (N140, N139, N73, N96);
buf BUF1 (N141, N130);
buf BUF1 (N142, N133);
not NOT1 (N143, N142);
not NOT1 (N144, N141);
nor NOR2 (N145, N128, N122);
nor NOR2 (N146, N73, N86);
and AND4 (N147, N143, N121, N16, N121);
not NOT1 (N148, N145);
not NOT1 (N149, N140);
buf BUF1 (N150, N134);
nand NAND4 (N151, N144, N46, N110, N17);
or OR4 (N152, N146, N20, N23, N118);
nand NAND3 (N153, N97, N56, N8);
and AND3 (N154, N151, N57, N136);
and AND3 (N155, N106, N25, N2);
or OR3 (N156, N149, N48, N87);
xor XOR2 (N157, N123, N21);
or OR2 (N158, N152, N59);
buf BUF1 (N159, N153);
not NOT1 (N160, N155);
and AND4 (N161, N132, N24, N55, N59);
xor XOR2 (N162, N156, N17);
not NOT1 (N163, N154);
or OR2 (N164, N150, N75);
nor NOR2 (N165, N148, N94);
and AND2 (N166, N157, N8);
buf BUF1 (N167, N165);
not NOT1 (N168, N161);
and AND4 (N169, N160, N116, N43, N68);
buf BUF1 (N170, N163);
buf BUF1 (N171, N168);
not NOT1 (N172, N147);
or OR4 (N173, N162, N29, N149, N17);
nor NOR4 (N174, N171, N12, N104, N153);
not NOT1 (N175, N172);
xor XOR2 (N176, N159, N126);
and AND4 (N177, N166, N14, N126, N133);
not NOT1 (N178, N164);
nand NAND2 (N179, N178, N166);
or OR2 (N180, N175, N177);
not NOT1 (N181, N44);
buf BUF1 (N182, N176);
not NOT1 (N183, N179);
and AND3 (N184, N158, N99, N155);
or OR2 (N185, N183, N108);
not NOT1 (N186, N169);
and AND4 (N187, N167, N29, N13, N35);
nand NAND3 (N188, N181, N25, N71);
and AND2 (N189, N185, N24);
not NOT1 (N190, N189);
not NOT1 (N191, N182);
nand NAND4 (N192, N187, N21, N26, N106);
or OR4 (N193, N191, N148, N64, N24);
and AND2 (N194, N180, N43);
xor XOR2 (N195, N186, N36);
nand NAND3 (N196, N184, N74, N85);
and AND2 (N197, N174, N2);
nor NOR2 (N198, N170, N42);
buf BUF1 (N199, N198);
xor XOR2 (N200, N196, N160);
buf BUF1 (N201, N193);
or OR4 (N202, N192, N42, N164, N196);
and AND4 (N203, N201, N14, N4, N134);
nand NAND2 (N204, N200, N124);
nor NOR2 (N205, N188, N148);
nand NAND3 (N206, N202, N36, N15);
nor NOR4 (N207, N197, N183, N178, N125);
buf BUF1 (N208, N206);
or OR2 (N209, N194, N79);
buf BUF1 (N210, N195);
buf BUF1 (N211, N173);
not NOT1 (N212, N207);
nor NOR4 (N213, N190, N192, N80, N106);
and AND3 (N214, N209, N49, N80);
nand NAND4 (N215, N203, N157, N81, N160);
or OR3 (N216, N205, N187, N156);
and AND2 (N217, N204, N99);
or OR4 (N218, N211, N123, N9, N141);
nand NAND4 (N219, N216, N23, N172, N122);
not NOT1 (N220, N219);
and AND2 (N221, N210, N101);
buf BUF1 (N222, N220);
nand NAND3 (N223, N217, N79, N17);
not NOT1 (N224, N199);
and AND3 (N225, N212, N197, N157);
not NOT1 (N226, N223);
and AND2 (N227, N214, N136);
xor XOR2 (N228, N225, N44);
not NOT1 (N229, N218);
buf BUF1 (N230, N221);
and AND3 (N231, N213, N173, N38);
nor NOR3 (N232, N227, N105, N23);
not NOT1 (N233, N224);
nand NAND4 (N234, N228, N109, N76, N127);
nand NAND2 (N235, N232, N65);
or OR4 (N236, N235, N79, N231, N37);
not NOT1 (N237, N142);
or OR3 (N238, N236, N230, N108);
not NOT1 (N239, N194);
and AND2 (N240, N215, N58);
nand NAND3 (N241, N233, N39, N34);
buf BUF1 (N242, N226);
nor NOR3 (N243, N208, N209, N145);
or OR3 (N244, N237, N132, N47);
or OR4 (N245, N240, N85, N155, N122);
buf BUF1 (N246, N242);
buf BUF1 (N247, N246);
not NOT1 (N248, N243);
xor XOR2 (N249, N229, N134);
buf BUF1 (N250, N241);
not NOT1 (N251, N245);
or OR3 (N252, N249, N222, N141);
and AND3 (N253, N123, N182, N206);
nand NAND3 (N254, N238, N53, N72);
not NOT1 (N255, N253);
nor NOR3 (N256, N254, N125, N170);
and AND3 (N257, N248, N18, N45);
or OR4 (N258, N256, N132, N157, N224);
or OR2 (N259, N252, N21);
not NOT1 (N260, N255);
nor NOR2 (N261, N251, N41);
not NOT1 (N262, N239);
nand NAND4 (N263, N261, N235, N124, N250);
and AND2 (N264, N146, N134);
not NOT1 (N265, N262);
buf BUF1 (N266, N265);
nand NAND3 (N267, N258, N64, N187);
buf BUF1 (N268, N264);
nand NAND4 (N269, N267, N130, N204, N205);
buf BUF1 (N270, N259);
and AND4 (N271, N234, N16, N264, N135);
xor XOR2 (N272, N270, N204);
nor NOR4 (N273, N263, N69, N75, N162);
not NOT1 (N274, N272);
or OR3 (N275, N244, N250, N177);
and AND3 (N276, N274, N259, N264);
buf BUF1 (N277, N268);
buf BUF1 (N278, N276);
and AND3 (N279, N271, N157, N131);
nor NOR4 (N280, N278, N5, N194, N223);
not NOT1 (N281, N280);
xor XOR2 (N282, N279, N53);
nor NOR3 (N283, N247, N107, N60);
nand NAND3 (N284, N282, N58, N268);
and AND2 (N285, N281, N146);
not NOT1 (N286, N260);
buf BUF1 (N287, N275);
xor XOR2 (N288, N269, N180);
and AND2 (N289, N283, N124);
xor XOR2 (N290, N273, N114);
xor XOR2 (N291, N284, N83);
nand NAND2 (N292, N285, N176);
nand NAND2 (N293, N287, N73);
nor NOR3 (N294, N292, N291, N78);
not NOT1 (N295, N54);
buf BUF1 (N296, N266);
nor NOR3 (N297, N293, N235, N289);
xor XOR2 (N298, N24, N268);
and AND3 (N299, N288, N261, N207);
not NOT1 (N300, N257);
and AND3 (N301, N297, N107, N137);
xor XOR2 (N302, N299, N210);
not NOT1 (N303, N294);
buf BUF1 (N304, N296);
and AND2 (N305, N300, N51);
nor NOR3 (N306, N303, N204, N199);
and AND4 (N307, N304, N222, N7, N195);
nor NOR4 (N308, N298, N293, N54, N24);
nand NAND4 (N309, N301, N40, N230, N252);
nor NOR4 (N310, N309, N269, N72, N98);
nand NAND2 (N311, N307, N271);
or OR4 (N312, N306, N173, N300, N120);
buf BUF1 (N313, N286);
not NOT1 (N314, N295);
not NOT1 (N315, N277);
nor NOR3 (N316, N315, N304, N9);
nor NOR4 (N317, N310, N177, N312, N182);
not NOT1 (N318, N108);
buf BUF1 (N319, N302);
nor NOR2 (N320, N317, N43);
or OR4 (N321, N314, N102, N33, N174);
and AND2 (N322, N319, N261);
xor XOR2 (N323, N290, N138);
nor NOR4 (N324, N305, N5, N27, N135);
nor NOR4 (N325, N318, N224, N4, N243);
nand NAND4 (N326, N311, N298, N259, N208);
nor NOR3 (N327, N313, N152, N264);
or OR3 (N328, N326, N122, N211);
buf BUF1 (N329, N323);
and AND3 (N330, N325, N284, N66);
xor XOR2 (N331, N316, N320);
nor NOR3 (N332, N275, N200, N129);
nand NAND2 (N333, N331, N317);
and AND4 (N334, N332, N96, N272, N14);
nor NOR3 (N335, N329, N32, N24);
or OR4 (N336, N328, N74, N82, N68);
nand NAND4 (N337, N334, N296, N280, N309);
and AND4 (N338, N324, N289, N247, N306);
not NOT1 (N339, N327);
nor NOR3 (N340, N333, N334, N169);
nor NOR3 (N341, N322, N335, N10);
or OR3 (N342, N293, N158, N58);
or OR2 (N343, N339, N159);
or OR3 (N344, N336, N168, N240);
nor NOR3 (N345, N308, N91, N189);
or OR3 (N346, N338, N160, N268);
nand NAND2 (N347, N321, N262);
or OR2 (N348, N343, N269);
or OR2 (N349, N348, N188);
nor NOR3 (N350, N337, N319, N38);
and AND3 (N351, N347, N30, N320);
nand NAND3 (N352, N341, N9, N17);
or OR4 (N353, N344, N234, N140, N122);
not NOT1 (N354, N342);
nand NAND3 (N355, N345, N7, N131);
and AND4 (N356, N354, N52, N178, N246);
xor XOR2 (N357, N350, N219);
buf BUF1 (N358, N351);
not NOT1 (N359, N330);
or OR4 (N360, N355, N212, N175, N54);
buf BUF1 (N361, N346);
xor XOR2 (N362, N361, N294);
or OR3 (N363, N349, N71, N164);
and AND3 (N364, N356, N90, N262);
nand NAND4 (N365, N364, N75, N360, N57);
nand NAND4 (N366, N225, N331, N355, N227);
nand NAND3 (N367, N359, N126, N138);
xor XOR2 (N368, N367, N91);
or OR3 (N369, N357, N358, N37);
not NOT1 (N370, N95);
xor XOR2 (N371, N362, N210);
nor NOR2 (N372, N353, N156);
or OR3 (N373, N371, N273, N335);
nor NOR2 (N374, N370, N73);
buf BUF1 (N375, N365);
nor NOR4 (N376, N363, N160, N145, N205);
xor XOR2 (N377, N352, N56);
and AND3 (N378, N368, N133, N53);
and AND4 (N379, N374, N228, N177, N51);
xor XOR2 (N380, N378, N160);
or OR2 (N381, N366, N136);
nand NAND2 (N382, N376, N62);
or OR2 (N383, N372, N356);
or OR2 (N384, N383, N204);
nor NOR3 (N385, N382, N111, N81);
buf BUF1 (N386, N373);
buf BUF1 (N387, N385);
nand NAND3 (N388, N377, N19, N370);
nand NAND4 (N389, N379, N68, N80, N57);
buf BUF1 (N390, N380);
buf BUF1 (N391, N369);
nand NAND4 (N392, N390, N88, N261, N266);
nor NOR3 (N393, N387, N52, N285);
buf BUF1 (N394, N381);
buf BUF1 (N395, N389);
nand NAND3 (N396, N375, N94, N209);
xor XOR2 (N397, N388, N143);
not NOT1 (N398, N394);
buf BUF1 (N399, N386);
nor NOR3 (N400, N384, N34, N65);
not NOT1 (N401, N392);
buf BUF1 (N402, N391);
nor NOR2 (N403, N340, N206);
nand NAND3 (N404, N399, N223, N274);
nor NOR4 (N405, N398, N200, N194, N300);
not NOT1 (N406, N404);
xor XOR2 (N407, N397, N101);
xor XOR2 (N408, N406, N96);
not NOT1 (N409, N396);
nor NOR2 (N410, N400, N344);
xor XOR2 (N411, N393, N189);
buf BUF1 (N412, N409);
buf BUF1 (N413, N412);
xor XOR2 (N414, N403, N310);
nor NOR3 (N415, N410, N96, N238);
and AND2 (N416, N408, N343);
not NOT1 (N417, N415);
and AND4 (N418, N407, N386, N417, N167);
and AND3 (N419, N184, N76, N400);
or OR4 (N420, N411, N115, N369, N175);
not NOT1 (N421, N418);
xor XOR2 (N422, N401, N84);
xor XOR2 (N423, N416, N250);
not NOT1 (N424, N423);
xor XOR2 (N425, N419, N2);
xor XOR2 (N426, N414, N119);
nand NAND4 (N427, N421, N297, N65, N109);
nor NOR4 (N428, N425, N419, N381, N97);
nor NOR4 (N429, N405, N370, N127, N51);
not NOT1 (N430, N427);
xor XOR2 (N431, N429, N342);
nor NOR3 (N432, N395, N160, N342);
or OR3 (N433, N432, N349, N308);
not NOT1 (N434, N413);
xor XOR2 (N435, N426, N306);
and AND3 (N436, N430, N408, N151);
or OR3 (N437, N431, N224, N368);
xor XOR2 (N438, N402, N255);
nand NAND3 (N439, N424, N105, N132);
nor NOR4 (N440, N420, N184, N415, N310);
or OR3 (N441, N436, N175, N288);
buf BUF1 (N442, N433);
nor NOR2 (N443, N422, N207);
nand NAND4 (N444, N439, N156, N264, N51);
xor XOR2 (N445, N444, N249);
or OR3 (N446, N445, N285, N22);
nor NOR2 (N447, N434, N71);
nand NAND4 (N448, N442, N251, N105, N4);
xor XOR2 (N449, N446, N7);
and AND4 (N450, N441, N188, N49, N198);
nor NOR4 (N451, N428, N402, N239, N248);
buf BUF1 (N452, N450);
nand NAND3 (N453, N447, N229, N397);
nor NOR4 (N454, N438, N302, N114, N391);
nand NAND3 (N455, N453, N437, N311);
nor NOR3 (N456, N290, N138, N305);
nand NAND2 (N457, N448, N75);
or OR2 (N458, N435, N5);
xor XOR2 (N459, N456, N54);
nand NAND2 (N460, N440, N66);
nor NOR2 (N461, N443, N127);
and AND3 (N462, N452, N334, N21);
xor XOR2 (N463, N460, N223);
nor NOR2 (N464, N455, N415);
and AND4 (N465, N459, N318, N162, N359);
and AND2 (N466, N457, N170);
nor NOR3 (N467, N465, N255, N20);
xor XOR2 (N468, N454, N317);
and AND2 (N469, N466, N165);
and AND3 (N470, N469, N52, N431);
nand NAND3 (N471, N467, N449, N343);
and AND4 (N472, N270, N168, N429, N159);
or OR3 (N473, N464, N102, N114);
nand NAND4 (N474, N458, N129, N427, N245);
or OR3 (N475, N473, N216, N404);
xor XOR2 (N476, N461, N246);
nand NAND3 (N477, N475, N456, N141);
not NOT1 (N478, N472);
not NOT1 (N479, N476);
or OR2 (N480, N462, N217);
and AND3 (N481, N478, N352, N444);
and AND2 (N482, N481, N356);
nand NAND4 (N483, N451, N196, N264, N160);
or OR2 (N484, N474, N234);
buf BUF1 (N485, N468);
nor NOR3 (N486, N470, N158, N483);
and AND3 (N487, N106, N326, N433);
xor XOR2 (N488, N484, N267);
xor XOR2 (N489, N471, N302);
xor XOR2 (N490, N482, N250);
nor NOR4 (N491, N487, N332, N33, N235);
not NOT1 (N492, N490);
not NOT1 (N493, N492);
nand NAND3 (N494, N485, N328, N251);
and AND2 (N495, N463, N203);
and AND2 (N496, N488, N63);
nand NAND3 (N497, N480, N349, N244);
not NOT1 (N498, N477);
nand NAND2 (N499, N497, N419);
or OR4 (N500, N498, N268, N353, N147);
buf BUF1 (N501, N491);
and AND3 (N502, N500, N342, N357);
buf BUF1 (N503, N493);
nand NAND4 (N504, N479, N35, N338, N231);
xor XOR2 (N505, N501, N400);
or OR3 (N506, N502, N381, N343);
buf BUF1 (N507, N486);
not NOT1 (N508, N489);
nor NOR4 (N509, N506, N345, N335, N434);
xor XOR2 (N510, N496, N24);
xor XOR2 (N511, N508, N176);
or OR4 (N512, N509, N382, N498, N280);
or OR2 (N513, N510, N45);
xor XOR2 (N514, N504, N267);
buf BUF1 (N515, N494);
nor NOR3 (N516, N507, N155, N210);
buf BUF1 (N517, N505);
nand NAND3 (N518, N503, N242, N490);
xor XOR2 (N519, N499, N308);
or OR4 (N520, N512, N250, N161, N295);
or OR2 (N521, N511, N414);
buf BUF1 (N522, N513);
not NOT1 (N523, N518);
nor NOR3 (N524, N520, N444, N169);
not NOT1 (N525, N519);
nand NAND4 (N526, N516, N414, N514, N344);
not NOT1 (N527, N162);
buf BUF1 (N528, N521);
nand NAND2 (N529, N517, N374);
not NOT1 (N530, N495);
or OR3 (N531, N528, N30, N507);
nor NOR2 (N532, N527, N331);
nor NOR2 (N533, N524, N303);
nor NOR2 (N534, N525, N70);
and AND2 (N535, N530, N530);
xor XOR2 (N536, N515, N495);
nand NAND2 (N537, N522, N91);
or OR3 (N538, N526, N524, N119);
not NOT1 (N539, N529);
or OR3 (N540, N539, N253, N522);
nand NAND4 (N541, N532, N43, N539, N117);
not NOT1 (N542, N531);
and AND3 (N543, N537, N168, N13);
nand NAND2 (N544, N535, N155);
nor NOR2 (N545, N538, N528);
xor XOR2 (N546, N533, N144);
and AND4 (N547, N534, N84, N116, N360);
xor XOR2 (N548, N544, N10);
nor NOR2 (N549, N547, N51);
and AND3 (N550, N543, N204, N28);
nor NOR4 (N551, N549, N132, N203, N235);
or OR2 (N552, N546, N40);
xor XOR2 (N553, N541, N495);
xor XOR2 (N554, N548, N516);
and AND2 (N555, N542, N471);
and AND3 (N556, N540, N235, N141);
nand NAND4 (N557, N550, N439, N405, N528);
nor NOR4 (N558, N555, N154, N482, N282);
nor NOR2 (N559, N553, N458);
buf BUF1 (N560, N554);
or OR4 (N561, N559, N221, N204, N496);
xor XOR2 (N562, N557, N343);
xor XOR2 (N563, N561, N32);
nand NAND2 (N564, N562, N488);
nand NAND4 (N565, N563, N450, N463, N120);
nand NAND2 (N566, N558, N94);
or OR3 (N567, N545, N352, N302);
or OR3 (N568, N523, N491, N216);
buf BUF1 (N569, N566);
or OR4 (N570, N560, N226, N121, N93);
nor NOR3 (N571, N565, N502, N43);
and AND2 (N572, N568, N231);
or OR3 (N573, N536, N192, N49);
buf BUF1 (N574, N571);
nand NAND2 (N575, N572, N124);
not NOT1 (N576, N574);
and AND2 (N577, N575, N89);
not NOT1 (N578, N564);
buf BUF1 (N579, N556);
and AND3 (N580, N578, N226, N397);
and AND2 (N581, N573, N315);
buf BUF1 (N582, N577);
not NOT1 (N583, N581);
xor XOR2 (N584, N579, N377);
not NOT1 (N585, N569);
nor NOR2 (N586, N570, N44);
xor XOR2 (N587, N567, N422);
not NOT1 (N588, N580);
not NOT1 (N589, N587);
or OR2 (N590, N552, N587);
nor NOR4 (N591, N585, N364, N436, N36);
nor NOR3 (N592, N576, N74, N557);
buf BUF1 (N593, N592);
xor XOR2 (N594, N551, N455);
not NOT1 (N595, N594);
nor NOR4 (N596, N589, N252, N467, N129);
and AND2 (N597, N588, N283);
or OR3 (N598, N596, N443, N87);
xor XOR2 (N599, N583, N259);
nand NAND2 (N600, N591, N480);
buf BUF1 (N601, N600);
buf BUF1 (N602, N586);
xor XOR2 (N603, N584, N175);
nor NOR4 (N604, N603, N101, N271, N35);
buf BUF1 (N605, N598);
xor XOR2 (N606, N595, N472);
buf BUF1 (N607, N604);
or OR4 (N608, N582, N236, N350, N602);
or OR4 (N609, N221, N102, N229, N421);
nor NOR4 (N610, N599, N252, N176, N148);
buf BUF1 (N611, N601);
buf BUF1 (N612, N608);
buf BUF1 (N613, N606);
or OR2 (N614, N612, N119);
and AND2 (N615, N609, N240);
not NOT1 (N616, N590);
and AND2 (N617, N616, N332);
and AND2 (N618, N605, N388);
nor NOR3 (N619, N593, N297, N566);
and AND4 (N620, N607, N517, N284, N416);
and AND2 (N621, N617, N348);
xor XOR2 (N622, N621, N115);
nor NOR2 (N623, N611, N587);
buf BUF1 (N624, N623);
or OR4 (N625, N614, N219, N474, N27);
not NOT1 (N626, N597);
nor NOR3 (N627, N620, N400, N294);
xor XOR2 (N628, N619, N81);
xor XOR2 (N629, N622, N327);
or OR2 (N630, N618, N514);
nand NAND3 (N631, N627, N121, N446);
nand NAND2 (N632, N624, N482);
buf BUF1 (N633, N631);
nand NAND4 (N634, N626, N101, N192, N328);
nor NOR3 (N635, N634, N579, N17);
and AND4 (N636, N635, N207, N246, N614);
not NOT1 (N637, N615);
nor NOR2 (N638, N636, N417);
buf BUF1 (N639, N628);
not NOT1 (N640, N629);
nor NOR2 (N641, N613, N42);
and AND4 (N642, N637, N381, N42, N190);
buf BUF1 (N643, N639);
xor XOR2 (N644, N630, N447);
and AND3 (N645, N640, N127, N307);
or OR4 (N646, N644, N410, N309, N62);
and AND3 (N647, N645, N453, N519);
not NOT1 (N648, N642);
not NOT1 (N649, N633);
nand NAND2 (N650, N646, N207);
buf BUF1 (N651, N647);
and AND3 (N652, N650, N295, N179);
or OR2 (N653, N649, N623);
not NOT1 (N654, N648);
nor NOR2 (N655, N652, N642);
nand NAND2 (N656, N643, N603);
xor XOR2 (N657, N655, N136);
nand NAND3 (N658, N653, N23, N159);
or OR3 (N659, N658, N460, N132);
xor XOR2 (N660, N657, N217);
nand NAND3 (N661, N625, N356, N175);
nor NOR4 (N662, N610, N99, N51, N56);
xor XOR2 (N663, N659, N641);
nor NOR2 (N664, N411, N657);
nand NAND4 (N665, N638, N387, N108, N178);
nand NAND3 (N666, N662, N639, N131);
buf BUF1 (N667, N661);
buf BUF1 (N668, N667);
not NOT1 (N669, N668);
xor XOR2 (N670, N666, N38);
nand NAND4 (N671, N656, N437, N131, N233);
nor NOR4 (N672, N664, N647, N602, N561);
nor NOR3 (N673, N660, N47, N282);
not NOT1 (N674, N654);
and AND4 (N675, N674, N496, N392, N652);
or OR2 (N676, N671, N228);
xor XOR2 (N677, N632, N672);
buf BUF1 (N678, N357);
not NOT1 (N679, N676);
and AND3 (N680, N665, N377, N101);
and AND2 (N681, N677, N29);
not NOT1 (N682, N651);
buf BUF1 (N683, N681);
or OR4 (N684, N682, N495, N457, N617);
nand NAND3 (N685, N679, N440, N203);
xor XOR2 (N686, N670, N413);
xor XOR2 (N687, N669, N415);
xor XOR2 (N688, N683, N315);
or OR3 (N689, N688, N592, N284);
and AND4 (N690, N675, N403, N235, N518);
buf BUF1 (N691, N684);
not NOT1 (N692, N678);
buf BUF1 (N693, N673);
xor XOR2 (N694, N690, N27);
nor NOR4 (N695, N692, N129, N263, N153);
not NOT1 (N696, N691);
nor NOR2 (N697, N693, N272);
buf BUF1 (N698, N689);
nand NAND3 (N699, N686, N595, N615);
nand NAND4 (N700, N698, N190, N451, N63);
not NOT1 (N701, N696);
nor NOR4 (N702, N701, N477, N627, N135);
not NOT1 (N703, N700);
and AND2 (N704, N680, N411);
not NOT1 (N705, N703);
buf BUF1 (N706, N695);
nand NAND4 (N707, N685, N215, N666, N637);
and AND2 (N708, N697, N299);
xor XOR2 (N709, N706, N674);
or OR2 (N710, N708, N273);
not NOT1 (N711, N705);
nor NOR2 (N712, N687, N56);
not NOT1 (N713, N694);
nand NAND2 (N714, N702, N280);
nand NAND4 (N715, N707, N427, N174, N107);
and AND3 (N716, N712, N642, N426);
not NOT1 (N717, N713);
nand NAND3 (N718, N716, N300, N17);
or OR3 (N719, N714, N546, N375);
or OR2 (N720, N711, N618);
and AND4 (N721, N710, N158, N55, N125);
not NOT1 (N722, N699);
and AND4 (N723, N709, N291, N589, N217);
xor XOR2 (N724, N704, N403);
nor NOR2 (N725, N721, N592);
xor XOR2 (N726, N717, N138);
and AND2 (N727, N719, N51);
nand NAND4 (N728, N663, N525, N571, N606);
nand NAND3 (N729, N727, N680, N213);
or OR2 (N730, N729, N370);
nor NOR4 (N731, N722, N101, N662, N119);
buf BUF1 (N732, N730);
or OR3 (N733, N731, N142, N444);
xor XOR2 (N734, N724, N708);
not NOT1 (N735, N720);
xor XOR2 (N736, N734, N665);
buf BUF1 (N737, N733);
buf BUF1 (N738, N732);
nor NOR3 (N739, N735, N313, N249);
or OR4 (N740, N723, N591, N79, N59);
nand NAND3 (N741, N736, N341, N710);
or OR4 (N742, N726, N37, N125, N144);
nor NOR3 (N743, N742, N437, N607);
buf BUF1 (N744, N740);
or OR3 (N745, N715, N253, N21);
xor XOR2 (N746, N745, N651);
buf BUF1 (N747, N744);
or OR2 (N748, N737, N242);
xor XOR2 (N749, N747, N410);
nor NOR4 (N750, N746, N114, N365, N731);
nor NOR3 (N751, N738, N455, N183);
nor NOR4 (N752, N725, N120, N80, N597);
buf BUF1 (N753, N748);
and AND2 (N754, N743, N630);
and AND4 (N755, N753, N210, N190, N195);
and AND4 (N756, N718, N234, N202, N292);
not NOT1 (N757, N756);
or OR3 (N758, N741, N313, N497);
buf BUF1 (N759, N728);
or OR2 (N760, N754, N660);
buf BUF1 (N761, N739);
xor XOR2 (N762, N759, N163);
or OR3 (N763, N752, N473, N550);
nand NAND3 (N764, N760, N366, N464);
nor NOR2 (N765, N757, N407);
buf BUF1 (N766, N751);
xor XOR2 (N767, N763, N358);
nor NOR2 (N768, N762, N291);
not NOT1 (N769, N761);
xor XOR2 (N770, N765, N174);
nor NOR2 (N771, N750, N581);
buf BUF1 (N772, N771);
and AND4 (N773, N768, N685, N537, N380);
nor NOR4 (N774, N770, N121, N652, N497);
or OR4 (N775, N769, N696, N74, N291);
buf BUF1 (N776, N775);
xor XOR2 (N777, N767, N584);
buf BUF1 (N778, N773);
not NOT1 (N779, N774);
or OR2 (N780, N749, N42);
xor XOR2 (N781, N766, N185);
buf BUF1 (N782, N755);
nor NOR4 (N783, N776, N660, N163, N466);
buf BUF1 (N784, N779);
nand NAND2 (N785, N783, N335);
or OR4 (N786, N782, N491, N55, N57);
and AND2 (N787, N764, N516);
not NOT1 (N788, N778);
and AND2 (N789, N786, N609);
nor NOR2 (N790, N789, N715);
xor XOR2 (N791, N785, N113);
or OR3 (N792, N791, N131, N573);
nor NOR3 (N793, N777, N22, N563);
nand NAND4 (N794, N780, N696, N346, N297);
nor NOR3 (N795, N788, N718, N670);
nand NAND4 (N796, N784, N241, N234, N496);
not NOT1 (N797, N795);
or OR3 (N798, N796, N200, N254);
or OR2 (N799, N781, N753);
xor XOR2 (N800, N799, N259);
not NOT1 (N801, N772);
nor NOR2 (N802, N787, N184);
not NOT1 (N803, N792);
nand NAND3 (N804, N797, N222, N479);
or OR4 (N805, N793, N349, N716, N510);
nand NAND3 (N806, N794, N550, N28);
and AND4 (N807, N806, N128, N165, N722);
not NOT1 (N808, N800);
xor XOR2 (N809, N802, N602);
xor XOR2 (N810, N807, N94);
buf BUF1 (N811, N805);
not NOT1 (N812, N809);
xor XOR2 (N813, N812, N60);
buf BUF1 (N814, N803);
or OR3 (N815, N758, N137, N212);
or OR3 (N816, N798, N397, N297);
not NOT1 (N817, N811);
or OR4 (N818, N810, N155, N78, N236);
buf BUF1 (N819, N816);
nand NAND2 (N820, N804, N726);
buf BUF1 (N821, N790);
or OR2 (N822, N801, N662);
xor XOR2 (N823, N814, N96);
buf BUF1 (N824, N817);
or OR3 (N825, N819, N218, N415);
xor XOR2 (N826, N822, N210);
and AND3 (N827, N821, N120, N228);
nor NOR3 (N828, N827, N385, N424);
nand NAND2 (N829, N825, N181);
xor XOR2 (N830, N826, N441);
xor XOR2 (N831, N820, N318);
nand NAND4 (N832, N830, N123, N592, N830);
nand NAND3 (N833, N831, N514, N290);
nand NAND2 (N834, N833, N43);
buf BUF1 (N835, N824);
nand NAND3 (N836, N813, N507, N151);
xor XOR2 (N837, N828, N745);
xor XOR2 (N838, N808, N595);
buf BUF1 (N839, N818);
nor NOR3 (N840, N834, N602, N30);
or OR2 (N841, N815, N494);
and AND3 (N842, N832, N750, N182);
not NOT1 (N843, N836);
nand NAND3 (N844, N842, N764, N632);
nand NAND3 (N845, N838, N66, N779);
xor XOR2 (N846, N823, N289);
xor XOR2 (N847, N837, N753);
or OR2 (N848, N843, N165);
or OR2 (N849, N840, N268);
xor XOR2 (N850, N829, N212);
and AND4 (N851, N835, N415, N544, N530);
not NOT1 (N852, N849);
or OR3 (N853, N846, N410, N485);
and AND3 (N854, N851, N360, N389);
or OR4 (N855, N848, N475, N623, N463);
or OR2 (N856, N855, N128);
not NOT1 (N857, N844);
and AND3 (N858, N847, N612, N579);
buf BUF1 (N859, N850);
xor XOR2 (N860, N841, N739);
not NOT1 (N861, N859);
buf BUF1 (N862, N852);
not NOT1 (N863, N857);
or OR3 (N864, N862, N88, N671);
or OR2 (N865, N864, N741);
not NOT1 (N866, N865);
buf BUF1 (N867, N853);
xor XOR2 (N868, N845, N481);
buf BUF1 (N869, N860);
nand NAND4 (N870, N868, N440, N734, N498);
buf BUF1 (N871, N856);
or OR4 (N872, N861, N133, N692, N661);
xor XOR2 (N873, N870, N451);
or OR4 (N874, N863, N616, N687, N299);
nor NOR3 (N875, N866, N200, N670);
buf BUF1 (N876, N874);
buf BUF1 (N877, N876);
not NOT1 (N878, N871);
buf BUF1 (N879, N872);
xor XOR2 (N880, N873, N731);
xor XOR2 (N881, N879, N819);
nand NAND4 (N882, N854, N340, N178, N517);
not NOT1 (N883, N878);
nand NAND4 (N884, N883, N322, N446, N138);
buf BUF1 (N885, N858);
buf BUF1 (N886, N867);
or OR2 (N887, N839, N258);
or OR2 (N888, N875, N65);
nand NAND4 (N889, N886, N537, N348, N51);
xor XOR2 (N890, N885, N120);
buf BUF1 (N891, N889);
nand NAND2 (N892, N881, N881);
xor XOR2 (N893, N887, N414);
buf BUF1 (N894, N888);
buf BUF1 (N895, N884);
and AND3 (N896, N895, N669, N400);
nand NAND2 (N897, N869, N769);
buf BUF1 (N898, N896);
nand NAND3 (N899, N880, N378, N582);
not NOT1 (N900, N877);
nor NOR2 (N901, N893, N886);
nand NAND4 (N902, N901, N851, N455, N318);
not NOT1 (N903, N882);
and AND2 (N904, N891, N671);
nor NOR3 (N905, N902, N628, N180);
buf BUF1 (N906, N897);
nand NAND3 (N907, N903, N614, N768);
or OR2 (N908, N894, N121);
or OR4 (N909, N904, N735, N530, N489);
not NOT1 (N910, N908);
nand NAND4 (N911, N906, N5, N181, N266);
buf BUF1 (N912, N892);
or OR4 (N913, N900, N515, N600, N490);
not NOT1 (N914, N898);
nand NAND2 (N915, N909, N95);
or OR3 (N916, N905, N700, N125);
or OR2 (N917, N907, N254);
buf BUF1 (N918, N916);
buf BUF1 (N919, N910);
nand NAND3 (N920, N915, N248, N506);
buf BUF1 (N921, N917);
and AND2 (N922, N918, N465);
nand NAND4 (N923, N913, N817, N787, N570);
not NOT1 (N924, N921);
nand NAND3 (N925, N911, N679, N213);
and AND2 (N926, N899, N400);
xor XOR2 (N927, N922, N454);
nor NOR2 (N928, N926, N56);
not NOT1 (N929, N927);
buf BUF1 (N930, N928);
not NOT1 (N931, N930);
nand NAND4 (N932, N923, N249, N274, N806);
nand NAND4 (N933, N929, N427, N594, N593);
and AND2 (N934, N890, N877);
xor XOR2 (N935, N919, N584);
and AND4 (N936, N912, N711, N679, N849);
buf BUF1 (N937, N920);
xor XOR2 (N938, N937, N841);
and AND2 (N939, N931, N832);
not NOT1 (N940, N925);
xor XOR2 (N941, N939, N214);
or OR3 (N942, N941, N753, N45);
not NOT1 (N943, N933);
or OR3 (N944, N935, N618, N206);
nand NAND4 (N945, N940, N330, N151, N695);
or OR2 (N946, N945, N274);
xor XOR2 (N947, N924, N527);
or OR3 (N948, N938, N432, N707);
or OR3 (N949, N914, N390, N782);
nand NAND2 (N950, N936, N409);
nor NOR3 (N951, N944, N424, N117);
xor XOR2 (N952, N946, N656);
and AND4 (N953, N943, N636, N627, N494);
buf BUF1 (N954, N949);
not NOT1 (N955, N947);
and AND3 (N956, N955, N19, N503);
buf BUF1 (N957, N950);
nor NOR2 (N958, N952, N733);
buf BUF1 (N959, N951);
or OR2 (N960, N942, N694);
xor XOR2 (N961, N954, N423);
nor NOR3 (N962, N957, N466, N642);
not NOT1 (N963, N958);
and AND2 (N964, N963, N67);
nor NOR3 (N965, N961, N660, N317);
xor XOR2 (N966, N953, N68);
or OR4 (N967, N962, N47, N534, N794);
buf BUF1 (N968, N967);
xor XOR2 (N969, N959, N654);
xor XOR2 (N970, N956, N700);
buf BUF1 (N971, N966);
and AND3 (N972, N968, N716, N159);
nor NOR4 (N973, N964, N790, N889, N250);
or OR3 (N974, N965, N127, N553);
or OR3 (N975, N973, N431, N228);
not NOT1 (N976, N971);
or OR2 (N977, N975, N194);
and AND2 (N978, N948, N905);
not NOT1 (N979, N974);
and AND3 (N980, N934, N257, N191);
and AND4 (N981, N976, N682, N761, N182);
or OR2 (N982, N979, N685);
nand NAND4 (N983, N981, N256, N158, N395);
not NOT1 (N984, N983);
and AND3 (N985, N982, N233, N651);
not NOT1 (N986, N984);
nand NAND2 (N987, N969, N477);
not NOT1 (N988, N978);
and AND4 (N989, N986, N65, N221, N22);
or OR2 (N990, N977, N721);
xor XOR2 (N991, N932, N868);
and AND3 (N992, N987, N846, N91);
buf BUF1 (N993, N970);
and AND4 (N994, N992, N103, N600, N151);
not NOT1 (N995, N994);
buf BUF1 (N996, N960);
buf BUF1 (N997, N989);
not NOT1 (N998, N990);
and AND3 (N999, N995, N618, N609);
not NOT1 (N1000, N980);
and AND4 (N1001, N993, N37, N169, N682);
buf BUF1 (N1002, N999);
not NOT1 (N1003, N1000);
and AND2 (N1004, N985, N395);
and AND4 (N1005, N1001, N122, N447, N816);
xor XOR2 (N1006, N997, N844);
xor XOR2 (N1007, N972, N370);
nor NOR4 (N1008, N1004, N514, N886, N492);
not NOT1 (N1009, N1007);
not NOT1 (N1010, N1003);
and AND4 (N1011, N1008, N535, N460, N855);
xor XOR2 (N1012, N1009, N994);
and AND4 (N1013, N988, N516, N661, N632);
nand NAND3 (N1014, N1006, N1002, N191);
nand NAND3 (N1015, N515, N461, N242);
and AND2 (N1016, N996, N961);
and AND2 (N1017, N1015, N19);
and AND4 (N1018, N1012, N906, N284, N775);
or OR2 (N1019, N991, N971);
xor XOR2 (N1020, N1010, N374);
buf BUF1 (N1021, N1011);
xor XOR2 (N1022, N1014, N681);
not NOT1 (N1023, N1005);
nor NOR4 (N1024, N1022, N927, N188, N579);
or OR3 (N1025, N1024, N305, N862);
xor XOR2 (N1026, N1019, N875);
nand NAND3 (N1027, N998, N896, N921);
nand NAND3 (N1028, N1013, N683, N134);
nor NOR3 (N1029, N1028, N820, N597);
xor XOR2 (N1030, N1018, N403);
not NOT1 (N1031, N1029);
or OR4 (N1032, N1026, N809, N865, N718);
nand NAND2 (N1033, N1032, N851);
xor XOR2 (N1034, N1033, N667);
and AND3 (N1035, N1030, N153, N392);
nand NAND3 (N1036, N1020, N415, N796);
nor NOR3 (N1037, N1027, N476, N410);
not NOT1 (N1038, N1025);
not NOT1 (N1039, N1023);
not NOT1 (N1040, N1016);
nor NOR3 (N1041, N1034, N396, N491);
not NOT1 (N1042, N1041);
nand NAND4 (N1043, N1035, N92, N466, N542);
buf BUF1 (N1044, N1037);
or OR2 (N1045, N1021, N83);
not NOT1 (N1046, N1042);
not NOT1 (N1047, N1038);
nor NOR4 (N1048, N1036, N423, N779, N614);
not NOT1 (N1049, N1047);
and AND4 (N1050, N1044, N378, N282, N146);
not NOT1 (N1051, N1039);
nor NOR3 (N1052, N1048, N402, N417);
nand NAND4 (N1053, N1043, N408, N940, N223);
xor XOR2 (N1054, N1050, N583);
nor NOR4 (N1055, N1031, N1029, N277, N938);
nand NAND4 (N1056, N1055, N462, N185, N188);
nand NAND4 (N1057, N1017, N917, N509, N760);
buf BUF1 (N1058, N1053);
buf BUF1 (N1059, N1052);
or OR4 (N1060, N1059, N800, N299, N355);
and AND4 (N1061, N1056, N488, N943, N355);
buf BUF1 (N1062, N1045);
or OR3 (N1063, N1046, N158, N234);
and AND3 (N1064, N1049, N111, N355);
nand NAND4 (N1065, N1054, N262, N651, N412);
or OR4 (N1066, N1058, N1010, N214, N123);
nand NAND3 (N1067, N1057, N856, N573);
or OR4 (N1068, N1064, N764, N987, N26);
xor XOR2 (N1069, N1067, N94);
or OR4 (N1070, N1063, N393, N821, N7);
nor NOR2 (N1071, N1068, N113);
or OR3 (N1072, N1062, N777, N251);
buf BUF1 (N1073, N1071);
nor NOR3 (N1074, N1073, N507, N103);
buf BUF1 (N1075, N1066);
and AND3 (N1076, N1069, N496, N866);
nor NOR3 (N1077, N1065, N311, N95);
not NOT1 (N1078, N1060);
not NOT1 (N1079, N1076);
buf BUF1 (N1080, N1077);
xor XOR2 (N1081, N1074, N542);
xor XOR2 (N1082, N1070, N600);
or OR2 (N1083, N1075, N826);
buf BUF1 (N1084, N1081);
and AND3 (N1085, N1078, N677, N143);
and AND2 (N1086, N1085, N88);
or OR3 (N1087, N1082, N784, N462);
nand NAND3 (N1088, N1072, N169, N280);
xor XOR2 (N1089, N1080, N292);
or OR4 (N1090, N1084, N340, N411, N645);
not NOT1 (N1091, N1089);
and AND4 (N1092, N1086, N749, N86, N79);
nand NAND3 (N1093, N1092, N982, N963);
and AND4 (N1094, N1087, N256, N651, N818);
nand NAND3 (N1095, N1040, N1005, N941);
or OR3 (N1096, N1083, N86, N889);
or OR4 (N1097, N1088, N921, N781, N475);
nand NAND2 (N1098, N1097, N36);
xor XOR2 (N1099, N1093, N416);
xor XOR2 (N1100, N1099, N884);
xor XOR2 (N1101, N1100, N739);
nand NAND3 (N1102, N1095, N984, N233);
or OR4 (N1103, N1098, N155, N139, N941);
and AND3 (N1104, N1103, N317, N623);
nand NAND2 (N1105, N1096, N624);
not NOT1 (N1106, N1102);
buf BUF1 (N1107, N1106);
not NOT1 (N1108, N1107);
xor XOR2 (N1109, N1101, N682);
not NOT1 (N1110, N1090);
xor XOR2 (N1111, N1061, N341);
or OR2 (N1112, N1110, N584);
buf BUF1 (N1113, N1105);
buf BUF1 (N1114, N1094);
nand NAND3 (N1115, N1113, N21, N559);
and AND3 (N1116, N1079, N260, N378);
and AND3 (N1117, N1112, N531, N189);
xor XOR2 (N1118, N1116, N778);
and AND3 (N1119, N1115, N634, N835);
nand NAND4 (N1120, N1109, N11, N310, N792);
and AND3 (N1121, N1117, N644, N437);
xor XOR2 (N1122, N1121, N193);
and AND3 (N1123, N1119, N278, N994);
xor XOR2 (N1124, N1114, N206);
xor XOR2 (N1125, N1108, N524);
and AND3 (N1126, N1091, N584, N420);
and AND2 (N1127, N1120, N239);
xor XOR2 (N1128, N1122, N925);
not NOT1 (N1129, N1118);
xor XOR2 (N1130, N1124, N543);
not NOT1 (N1131, N1130);
xor XOR2 (N1132, N1123, N1071);
nor NOR3 (N1133, N1129, N276, N415);
buf BUF1 (N1134, N1126);
buf BUF1 (N1135, N1131);
or OR2 (N1136, N1104, N538);
buf BUF1 (N1137, N1125);
nor NOR2 (N1138, N1111, N167);
and AND2 (N1139, N1135, N439);
xor XOR2 (N1140, N1051, N315);
xor XOR2 (N1141, N1137, N456);
nor NOR2 (N1142, N1136, N311);
buf BUF1 (N1143, N1133);
not NOT1 (N1144, N1128);
nand NAND2 (N1145, N1134, N1081);
nand NAND2 (N1146, N1143, N363);
and AND4 (N1147, N1138, N255, N449, N148);
nand NAND2 (N1148, N1144, N391);
nor NOR2 (N1149, N1147, N301);
not NOT1 (N1150, N1146);
and AND4 (N1151, N1149, N1070, N921, N601);
not NOT1 (N1152, N1150);
xor XOR2 (N1153, N1152, N633);
nor NOR2 (N1154, N1127, N358);
or OR3 (N1155, N1140, N207, N714);
nor NOR2 (N1156, N1148, N241);
or OR4 (N1157, N1155, N653, N940, N1053);
xor XOR2 (N1158, N1157, N444);
xor XOR2 (N1159, N1154, N1105);
nand NAND4 (N1160, N1158, N223, N720, N1051);
and AND3 (N1161, N1160, N1062, N259);
buf BUF1 (N1162, N1161);
and AND4 (N1163, N1156, N755, N556, N1162);
and AND3 (N1164, N332, N383, N1093);
buf BUF1 (N1165, N1153);
and AND3 (N1166, N1164, N149, N336);
xor XOR2 (N1167, N1151, N600);
not NOT1 (N1168, N1163);
nor NOR3 (N1169, N1139, N806, N352);
or OR4 (N1170, N1141, N377, N84, N190);
nor NOR2 (N1171, N1166, N694);
xor XOR2 (N1172, N1171, N1027);
and AND4 (N1173, N1170, N442, N1093, N73);
and AND3 (N1174, N1145, N326, N865);
and AND3 (N1175, N1142, N555, N832);
not NOT1 (N1176, N1169);
xor XOR2 (N1177, N1172, N1074);
buf BUF1 (N1178, N1177);
and AND4 (N1179, N1168, N308, N946, N661);
or OR3 (N1180, N1167, N764, N767);
or OR2 (N1181, N1165, N145);
nor NOR4 (N1182, N1180, N807, N458, N373);
and AND3 (N1183, N1182, N827, N555);
not NOT1 (N1184, N1181);
nand NAND3 (N1185, N1132, N530, N1033);
not NOT1 (N1186, N1179);
nand NAND4 (N1187, N1186, N813, N91, N10);
nand NAND3 (N1188, N1176, N974, N1068);
nand NAND3 (N1189, N1174, N1069, N1121);
and AND3 (N1190, N1183, N228, N730);
and AND2 (N1191, N1187, N876);
or OR3 (N1192, N1191, N624, N605);
nand NAND2 (N1193, N1192, N217);
nor NOR3 (N1194, N1159, N587, N714);
xor XOR2 (N1195, N1189, N636);
nand NAND3 (N1196, N1190, N946, N1131);
or OR3 (N1197, N1193, N1117, N216);
xor XOR2 (N1198, N1196, N658);
buf BUF1 (N1199, N1188);
not NOT1 (N1200, N1173);
or OR2 (N1201, N1195, N956);
not NOT1 (N1202, N1198);
or OR3 (N1203, N1200, N15, N280);
nand NAND3 (N1204, N1185, N587, N161);
nor NOR3 (N1205, N1199, N827, N216);
buf BUF1 (N1206, N1203);
and AND3 (N1207, N1204, N957, N566);
xor XOR2 (N1208, N1178, N483);
xor XOR2 (N1209, N1208, N667);
buf BUF1 (N1210, N1197);
nor NOR3 (N1211, N1194, N953, N41);
and AND2 (N1212, N1175, N1181);
nor NOR2 (N1213, N1211, N92);
not NOT1 (N1214, N1213);
nor NOR2 (N1215, N1210, N107);
nor NOR4 (N1216, N1202, N337, N851, N195);
nor NOR2 (N1217, N1207, N264);
xor XOR2 (N1218, N1205, N895);
and AND3 (N1219, N1209, N171, N525);
not NOT1 (N1220, N1201);
not NOT1 (N1221, N1216);
or OR2 (N1222, N1219, N292);
not NOT1 (N1223, N1215);
buf BUF1 (N1224, N1220);
xor XOR2 (N1225, N1221, N899);
not NOT1 (N1226, N1218);
xor XOR2 (N1227, N1212, N909);
nor NOR3 (N1228, N1225, N652, N583);
and AND2 (N1229, N1214, N611);
nor NOR4 (N1230, N1224, N347, N758, N1000);
xor XOR2 (N1231, N1228, N536);
nor NOR4 (N1232, N1226, N167, N55, N1107);
xor XOR2 (N1233, N1222, N765);
nand NAND4 (N1234, N1184, N544, N682, N893);
buf BUF1 (N1235, N1206);
nor NOR3 (N1236, N1234, N298, N392);
xor XOR2 (N1237, N1232, N1148);
buf BUF1 (N1238, N1227);
or OR2 (N1239, N1217, N1131);
xor XOR2 (N1240, N1236, N661);
and AND3 (N1241, N1239, N748, N655);
nand NAND4 (N1242, N1240, N251, N1077, N446);
buf BUF1 (N1243, N1229);
nor NOR3 (N1244, N1243, N33, N1029);
nand NAND4 (N1245, N1238, N993, N1197, N89);
nand NAND3 (N1246, N1235, N600, N939);
nor NOR3 (N1247, N1244, N6, N289);
or OR3 (N1248, N1237, N619, N702);
buf BUF1 (N1249, N1242);
not NOT1 (N1250, N1241);
xor XOR2 (N1251, N1248, N714);
not NOT1 (N1252, N1247);
xor XOR2 (N1253, N1249, N1247);
nor NOR2 (N1254, N1245, N150);
xor XOR2 (N1255, N1230, N607);
not NOT1 (N1256, N1231);
buf BUF1 (N1257, N1233);
buf BUF1 (N1258, N1223);
nand NAND2 (N1259, N1258, N1022);
nor NOR2 (N1260, N1250, N381);
nor NOR3 (N1261, N1252, N784, N159);
and AND3 (N1262, N1254, N237, N729);
and AND4 (N1263, N1251, N1251, N166, N393);
and AND3 (N1264, N1255, N1102, N651);
or OR2 (N1265, N1263, N99);
or OR2 (N1266, N1262, N315);
nor NOR3 (N1267, N1246, N954, N52);
or OR3 (N1268, N1265, N1191, N103);
buf BUF1 (N1269, N1257);
buf BUF1 (N1270, N1264);
nand NAND2 (N1271, N1267, N1198);
and AND2 (N1272, N1269, N116);
and AND3 (N1273, N1261, N261, N584);
or OR3 (N1274, N1270, N201, N1141);
nand NAND3 (N1275, N1271, N772, N964);
nor NOR2 (N1276, N1259, N558);
not NOT1 (N1277, N1256);
not NOT1 (N1278, N1274);
not NOT1 (N1279, N1266);
buf BUF1 (N1280, N1273);
buf BUF1 (N1281, N1277);
and AND3 (N1282, N1275, N72, N748);
not NOT1 (N1283, N1280);
or OR2 (N1284, N1281, N1075);
xor XOR2 (N1285, N1279, N39);
nand NAND4 (N1286, N1278, N213, N547, N1105);
and AND3 (N1287, N1253, N1167, N1016);
not NOT1 (N1288, N1284);
nor NOR3 (N1289, N1286, N551, N23);
buf BUF1 (N1290, N1276);
or OR2 (N1291, N1272, N963);
and AND2 (N1292, N1287, N848);
nand NAND4 (N1293, N1292, N741, N19, N1289);
xor XOR2 (N1294, N111, N480);
nor NOR3 (N1295, N1294, N1278, N992);
not NOT1 (N1296, N1283);
not NOT1 (N1297, N1268);
nand NAND3 (N1298, N1288, N269, N1009);
buf BUF1 (N1299, N1290);
buf BUF1 (N1300, N1260);
or OR2 (N1301, N1291, N427);
and AND4 (N1302, N1298, N316, N921, N394);
and AND3 (N1303, N1282, N511, N1188);
not NOT1 (N1304, N1293);
xor XOR2 (N1305, N1304, N1063);
and AND3 (N1306, N1301, N433, N78);
or OR4 (N1307, N1306, N1287, N568, N822);
not NOT1 (N1308, N1299);
buf BUF1 (N1309, N1307);
not NOT1 (N1310, N1295);
or OR2 (N1311, N1297, N231);
not NOT1 (N1312, N1308);
nor NOR4 (N1313, N1285, N67, N725, N1051);
not NOT1 (N1314, N1305);
buf BUF1 (N1315, N1300);
buf BUF1 (N1316, N1312);
not NOT1 (N1317, N1315);
xor XOR2 (N1318, N1310, N117);
nor NOR3 (N1319, N1318, N1260, N1044);
buf BUF1 (N1320, N1303);
xor XOR2 (N1321, N1313, N578);
or OR3 (N1322, N1311, N641, N450);
nand NAND2 (N1323, N1320, N968);
not NOT1 (N1324, N1317);
or OR4 (N1325, N1316, N1181, N784, N834);
nor NOR2 (N1326, N1322, N1231);
nor NOR2 (N1327, N1321, N228);
and AND3 (N1328, N1319, N1263, N1095);
xor XOR2 (N1329, N1325, N210);
xor XOR2 (N1330, N1327, N795);
not NOT1 (N1331, N1302);
and AND3 (N1332, N1328, N336, N1259);
nor NOR4 (N1333, N1324, N1086, N287, N372);
nor NOR4 (N1334, N1296, N544, N278, N608);
xor XOR2 (N1335, N1333, N1221);
buf BUF1 (N1336, N1334);
not NOT1 (N1337, N1314);
or OR3 (N1338, N1326, N901, N1117);
and AND4 (N1339, N1309, N380, N150, N110);
nor NOR2 (N1340, N1332, N1246);
or OR4 (N1341, N1335, N1239, N1319, N295);
not NOT1 (N1342, N1338);
not NOT1 (N1343, N1329);
nor NOR4 (N1344, N1330, N370, N473, N556);
or OR2 (N1345, N1337, N1239);
xor XOR2 (N1346, N1342, N1265);
xor XOR2 (N1347, N1340, N744);
not NOT1 (N1348, N1331);
or OR4 (N1349, N1346, N1038, N1213, N577);
and AND4 (N1350, N1345, N841, N318, N1029);
nand NAND3 (N1351, N1343, N295, N167);
and AND3 (N1352, N1347, N1223, N105);
not NOT1 (N1353, N1339);
buf BUF1 (N1354, N1348);
and AND2 (N1355, N1350, N1100);
nor NOR3 (N1356, N1344, N1185, N1060);
nand NAND3 (N1357, N1355, N511, N593);
not NOT1 (N1358, N1357);
or OR4 (N1359, N1323, N854, N169, N689);
not NOT1 (N1360, N1349);
xor XOR2 (N1361, N1353, N1076);
xor XOR2 (N1362, N1356, N671);
nand NAND2 (N1363, N1351, N774);
xor XOR2 (N1364, N1363, N339);
not NOT1 (N1365, N1354);
buf BUF1 (N1366, N1361);
buf BUF1 (N1367, N1360);
nor NOR2 (N1368, N1365, N942);
buf BUF1 (N1369, N1341);
xor XOR2 (N1370, N1336, N388);
buf BUF1 (N1371, N1352);
buf BUF1 (N1372, N1371);
nor NOR2 (N1373, N1367, N304);
and AND4 (N1374, N1372, N586, N455, N145);
not NOT1 (N1375, N1366);
or OR4 (N1376, N1370, N21, N18, N1334);
or OR2 (N1377, N1368, N1012);
nand NAND3 (N1378, N1364, N964, N990);
xor XOR2 (N1379, N1378, N991);
not NOT1 (N1380, N1359);
nand NAND2 (N1381, N1373, N1234);
xor XOR2 (N1382, N1381, N33);
nand NAND2 (N1383, N1374, N208);
or OR4 (N1384, N1375, N433, N1030, N339);
or OR3 (N1385, N1376, N1048, N586);
xor XOR2 (N1386, N1362, N1156);
buf BUF1 (N1387, N1369);
nand NAND2 (N1388, N1377, N561);
nor NOR2 (N1389, N1387, N65);
or OR4 (N1390, N1388, N418, N1101, N923);
not NOT1 (N1391, N1386);
not NOT1 (N1392, N1391);
buf BUF1 (N1393, N1380);
not NOT1 (N1394, N1358);
buf BUF1 (N1395, N1382);
nand NAND2 (N1396, N1393, N951);
and AND3 (N1397, N1395, N1381, N1387);
and AND2 (N1398, N1379, N20);
xor XOR2 (N1399, N1394, N668);
and AND4 (N1400, N1396, N253, N1275, N878);
nand NAND4 (N1401, N1399, N704, N909, N102);
buf BUF1 (N1402, N1400);
and AND3 (N1403, N1401, N542, N8);
or OR4 (N1404, N1403, N1118, N313, N335);
and AND4 (N1405, N1390, N1297, N997, N1237);
or OR4 (N1406, N1405, N922, N1056, N23);
xor XOR2 (N1407, N1402, N1226);
buf BUF1 (N1408, N1404);
or OR4 (N1409, N1392, N819, N1106, N1324);
xor XOR2 (N1410, N1397, N1013);
buf BUF1 (N1411, N1406);
or OR2 (N1412, N1411, N1074);
xor XOR2 (N1413, N1383, N599);
and AND2 (N1414, N1385, N18);
nand NAND3 (N1415, N1413, N368, N1293);
and AND3 (N1416, N1412, N727, N475);
or OR3 (N1417, N1409, N371, N1309);
buf BUF1 (N1418, N1417);
not NOT1 (N1419, N1408);
or OR4 (N1420, N1419, N706, N16, N1279);
buf BUF1 (N1421, N1384);
nor NOR4 (N1422, N1420, N277, N663, N869);
nor NOR3 (N1423, N1418, N547, N1364);
buf BUF1 (N1424, N1423);
or OR2 (N1425, N1414, N401);
xor XOR2 (N1426, N1422, N335);
not NOT1 (N1427, N1424);
buf BUF1 (N1428, N1398);
not NOT1 (N1429, N1427);
xor XOR2 (N1430, N1415, N43);
nand NAND4 (N1431, N1421, N436, N511, N1208);
and AND2 (N1432, N1410, N826);
xor XOR2 (N1433, N1428, N134);
nand NAND4 (N1434, N1433, N769, N1088, N764);
buf BUF1 (N1435, N1425);
xor XOR2 (N1436, N1430, N525);
xor XOR2 (N1437, N1431, N623);
or OR2 (N1438, N1416, N719);
not NOT1 (N1439, N1426);
not NOT1 (N1440, N1435);
buf BUF1 (N1441, N1438);
nand NAND3 (N1442, N1441, N630, N321);
and AND2 (N1443, N1439, N489);
buf BUF1 (N1444, N1389);
nor NOR3 (N1445, N1432, N168, N174);
nor NOR2 (N1446, N1445, N1237);
nor NOR3 (N1447, N1434, N58, N658);
buf BUF1 (N1448, N1436);
not NOT1 (N1449, N1446);
buf BUF1 (N1450, N1442);
buf BUF1 (N1451, N1440);
not NOT1 (N1452, N1444);
buf BUF1 (N1453, N1429);
xor XOR2 (N1454, N1437, N1432);
buf BUF1 (N1455, N1450);
nand NAND2 (N1456, N1443, N1313);
not NOT1 (N1457, N1448);
not NOT1 (N1458, N1447);
xor XOR2 (N1459, N1458, N1404);
or OR3 (N1460, N1455, N114, N500);
not NOT1 (N1461, N1456);
and AND2 (N1462, N1451, N850);
buf BUF1 (N1463, N1453);
nor NOR3 (N1464, N1452, N196, N574);
xor XOR2 (N1465, N1462, N1452);
nand NAND4 (N1466, N1465, N1343, N126, N299);
nand NAND3 (N1467, N1463, N240, N382);
xor XOR2 (N1468, N1459, N1451);
buf BUF1 (N1469, N1449);
or OR4 (N1470, N1460, N1156, N14, N1102);
xor XOR2 (N1471, N1469, N116);
xor XOR2 (N1472, N1468, N605);
not NOT1 (N1473, N1457);
or OR2 (N1474, N1467, N540);
nor NOR4 (N1475, N1461, N749, N1264, N199);
not NOT1 (N1476, N1475);
or OR2 (N1477, N1472, N1325);
nand NAND2 (N1478, N1470, N1267);
or OR2 (N1479, N1473, N834);
not NOT1 (N1480, N1466);
xor XOR2 (N1481, N1407, N1108);
and AND4 (N1482, N1478, N379, N271, N11);
not NOT1 (N1483, N1479);
or OR2 (N1484, N1483, N959);
and AND4 (N1485, N1474, N1083, N894, N1432);
xor XOR2 (N1486, N1480, N632);
nor NOR4 (N1487, N1454, N18, N835, N1395);
xor XOR2 (N1488, N1481, N858);
or OR3 (N1489, N1487, N318, N1308);
and AND2 (N1490, N1484, N1234);
not NOT1 (N1491, N1488);
xor XOR2 (N1492, N1490, N699);
xor XOR2 (N1493, N1485, N839);
xor XOR2 (N1494, N1471, N745);
not NOT1 (N1495, N1486);
not NOT1 (N1496, N1476);
not NOT1 (N1497, N1493);
xor XOR2 (N1498, N1489, N452);
buf BUF1 (N1499, N1491);
and AND2 (N1500, N1499, N1145);
nand NAND4 (N1501, N1497, N1051, N340, N535);
or OR3 (N1502, N1496, N511, N341);
not NOT1 (N1503, N1492);
xor XOR2 (N1504, N1502, N20);
not NOT1 (N1505, N1504);
nand NAND2 (N1506, N1477, N1398);
buf BUF1 (N1507, N1498);
buf BUF1 (N1508, N1506);
nand NAND2 (N1509, N1482, N140);
not NOT1 (N1510, N1508);
and AND4 (N1511, N1510, N969, N207, N1179);
or OR2 (N1512, N1500, N346);
xor XOR2 (N1513, N1501, N626);
nor NOR2 (N1514, N1507, N1141);
and AND2 (N1515, N1514, N362);
xor XOR2 (N1516, N1511, N495);
nand NAND2 (N1517, N1464, N347);
nand NAND2 (N1518, N1495, N1256);
or OR3 (N1519, N1509, N1333, N719);
or OR2 (N1520, N1513, N144);
and AND4 (N1521, N1494, N377, N113, N409);
xor XOR2 (N1522, N1519, N867);
xor XOR2 (N1523, N1503, N390);
not NOT1 (N1524, N1515);
not NOT1 (N1525, N1517);
buf BUF1 (N1526, N1505);
nand NAND3 (N1527, N1518, N902, N397);
buf BUF1 (N1528, N1525);
xor XOR2 (N1529, N1516, N1133);
not NOT1 (N1530, N1523);
and AND4 (N1531, N1526, N534, N1382, N1219);
nor NOR4 (N1532, N1527, N1088, N363, N1001);
and AND2 (N1533, N1529, N1382);
xor XOR2 (N1534, N1531, N150);
xor XOR2 (N1535, N1533, N671);
buf BUF1 (N1536, N1512);
not NOT1 (N1537, N1521);
nand NAND2 (N1538, N1530, N1263);
buf BUF1 (N1539, N1536);
nand NAND2 (N1540, N1537, N1378);
xor XOR2 (N1541, N1539, N66);
or OR2 (N1542, N1528, N911);
or OR4 (N1543, N1532, N33, N1308, N821);
not NOT1 (N1544, N1538);
or OR2 (N1545, N1534, N1345);
nand NAND2 (N1546, N1522, N1150);
nand NAND4 (N1547, N1543, N1042, N1016, N871);
nor NOR4 (N1548, N1546, N820, N403, N1060);
nor NOR3 (N1549, N1540, N219, N856);
xor XOR2 (N1550, N1520, N982);
nand NAND4 (N1551, N1550, N1447, N667, N1114);
nor NOR2 (N1552, N1524, N760);
nand NAND3 (N1553, N1544, N552, N1214);
nor NOR3 (N1554, N1553, N1187, N876);
nand NAND3 (N1555, N1552, N26, N771);
not NOT1 (N1556, N1545);
not NOT1 (N1557, N1549);
and AND4 (N1558, N1547, N230, N449, N775);
nor NOR3 (N1559, N1548, N1242, N1319);
or OR2 (N1560, N1555, N1280);
not NOT1 (N1561, N1556);
nor NOR4 (N1562, N1559, N113, N492, N661);
not NOT1 (N1563, N1562);
or OR2 (N1564, N1551, N595);
or OR3 (N1565, N1563, N1258, N627);
xor XOR2 (N1566, N1561, N1550);
and AND3 (N1567, N1564, N560, N518);
buf BUF1 (N1568, N1565);
or OR4 (N1569, N1541, N610, N230, N156);
buf BUF1 (N1570, N1554);
nand NAND2 (N1571, N1567, N1348);
xor XOR2 (N1572, N1535, N1269);
or OR2 (N1573, N1557, N1018);
xor XOR2 (N1574, N1542, N1036);
and AND4 (N1575, N1570, N520, N848, N507);
or OR2 (N1576, N1573, N568);
not NOT1 (N1577, N1560);
not NOT1 (N1578, N1569);
nor NOR3 (N1579, N1568, N59, N812);
and AND2 (N1580, N1558, N1562);
not NOT1 (N1581, N1566);
and AND2 (N1582, N1574, N1063);
not NOT1 (N1583, N1582);
nand NAND2 (N1584, N1581, N986);
xor XOR2 (N1585, N1576, N212);
buf BUF1 (N1586, N1580);
or OR2 (N1587, N1586, N418);
not NOT1 (N1588, N1579);
or OR2 (N1589, N1583, N1418);
not NOT1 (N1590, N1571);
or OR3 (N1591, N1572, N22, N331);
xor XOR2 (N1592, N1584, N974);
buf BUF1 (N1593, N1592);
buf BUF1 (N1594, N1591);
xor XOR2 (N1595, N1588, N1573);
xor XOR2 (N1596, N1595, N1105);
xor XOR2 (N1597, N1585, N1374);
not NOT1 (N1598, N1593);
xor XOR2 (N1599, N1589, N198);
and AND3 (N1600, N1596, N436, N1102);
and AND2 (N1601, N1597, N1022);
buf BUF1 (N1602, N1577);
xor XOR2 (N1603, N1601, N625);
nand NAND2 (N1604, N1600, N288);
not NOT1 (N1605, N1599);
nor NOR2 (N1606, N1578, N307);
or OR4 (N1607, N1602, N737, N37, N995);
and AND2 (N1608, N1590, N1275);
nand NAND4 (N1609, N1604, N928, N697, N1311);
xor XOR2 (N1610, N1594, N49);
or OR2 (N1611, N1607, N1503);
nand NAND3 (N1612, N1611, N1070, N1275);
and AND2 (N1613, N1608, N1383);
and AND4 (N1614, N1598, N1285, N1462, N635);
nor NOR3 (N1615, N1606, N1197, N455);
nor NOR4 (N1616, N1610, N1433, N581, N1250);
nand NAND3 (N1617, N1603, N1157, N551);
not NOT1 (N1618, N1587);
nand NAND4 (N1619, N1613, N135, N21, N1172);
nand NAND2 (N1620, N1619, N621);
or OR3 (N1621, N1609, N1529, N1384);
and AND2 (N1622, N1605, N1460);
xor XOR2 (N1623, N1622, N1130);
nand NAND4 (N1624, N1615, N1372, N306, N543);
xor XOR2 (N1625, N1624, N116);
xor XOR2 (N1626, N1621, N1359);
not NOT1 (N1627, N1614);
and AND4 (N1628, N1623, N654, N299, N358);
nand NAND2 (N1629, N1575, N1264);
nand NAND3 (N1630, N1618, N1482, N533);
xor XOR2 (N1631, N1626, N599);
nand NAND4 (N1632, N1616, N1595, N942, N1101);
not NOT1 (N1633, N1627);
xor XOR2 (N1634, N1629, N1343);
not NOT1 (N1635, N1617);
nand NAND2 (N1636, N1630, N1013);
buf BUF1 (N1637, N1636);
xor XOR2 (N1638, N1635, N600);
buf BUF1 (N1639, N1631);
or OR4 (N1640, N1625, N1007, N789, N460);
nor NOR3 (N1641, N1640, N463, N628);
or OR3 (N1642, N1637, N7, N1277);
xor XOR2 (N1643, N1620, N659);
nand NAND3 (N1644, N1639, N814, N550);
and AND2 (N1645, N1628, N1534);
and AND4 (N1646, N1633, N103, N1332, N1065);
and AND3 (N1647, N1646, N1137, N72);
xor XOR2 (N1648, N1642, N113);
not NOT1 (N1649, N1644);
not NOT1 (N1650, N1643);
buf BUF1 (N1651, N1632);
and AND4 (N1652, N1651, N1495, N162, N483);
xor XOR2 (N1653, N1634, N17);
nand NAND4 (N1654, N1645, N562, N1334, N249);
not NOT1 (N1655, N1653);
nand NAND2 (N1656, N1641, N831);
and AND3 (N1657, N1612, N1190, N353);
nor NOR2 (N1658, N1647, N804);
xor XOR2 (N1659, N1656, N1477);
or OR2 (N1660, N1655, N210);
xor XOR2 (N1661, N1649, N1653);
nor NOR2 (N1662, N1657, N921);
or OR2 (N1663, N1654, N569);
not NOT1 (N1664, N1648);
not NOT1 (N1665, N1660);
buf BUF1 (N1666, N1638);
nor NOR2 (N1667, N1664, N1190);
or OR3 (N1668, N1662, N1017, N1060);
not NOT1 (N1669, N1650);
buf BUF1 (N1670, N1668);
buf BUF1 (N1671, N1661);
or OR3 (N1672, N1665, N276, N1152);
or OR4 (N1673, N1652, N488, N508, N926);
nand NAND4 (N1674, N1663, N771, N699, N742);
nand NAND3 (N1675, N1670, N1114, N196);
nand NAND3 (N1676, N1671, N1086, N1482);
buf BUF1 (N1677, N1669);
not NOT1 (N1678, N1666);
buf BUF1 (N1679, N1677);
not NOT1 (N1680, N1675);
and AND4 (N1681, N1667, N508, N376, N1628);
nand NAND2 (N1682, N1659, N454);
xor XOR2 (N1683, N1673, N1583);
or OR2 (N1684, N1658, N1319);
or OR4 (N1685, N1683, N845, N679, N1043);
buf BUF1 (N1686, N1685);
nor NOR3 (N1687, N1678, N1120, N1661);
nor NOR4 (N1688, N1686, N582, N1082, N1477);
and AND4 (N1689, N1682, N1472, N1643, N1333);
or OR2 (N1690, N1688, N919);
xor XOR2 (N1691, N1690, N994);
not NOT1 (N1692, N1672);
not NOT1 (N1693, N1689);
nor NOR2 (N1694, N1684, N182);
nor NOR3 (N1695, N1681, N1223, N944);
nor NOR4 (N1696, N1687, N365, N670, N143);
not NOT1 (N1697, N1674);
nor NOR2 (N1698, N1695, N442);
or OR2 (N1699, N1679, N1619);
and AND2 (N1700, N1692, N302);
or OR4 (N1701, N1676, N1373, N1323, N88);
and AND3 (N1702, N1699, N548, N16);
buf BUF1 (N1703, N1691);
and AND3 (N1704, N1697, N1031, N1626);
nand NAND4 (N1705, N1696, N1055, N1462, N316);
and AND4 (N1706, N1703, N1486, N891, N826);
or OR2 (N1707, N1680, N337);
xor XOR2 (N1708, N1705, N776);
buf BUF1 (N1709, N1701);
not NOT1 (N1710, N1709);
not NOT1 (N1711, N1708);
and AND3 (N1712, N1700, N913, N949);
not NOT1 (N1713, N1694);
not NOT1 (N1714, N1698);
xor XOR2 (N1715, N1706, N791);
and AND2 (N1716, N1702, N145);
nor NOR2 (N1717, N1715, N1148);
nand NAND4 (N1718, N1712, N1487, N994, N475);
and AND3 (N1719, N1710, N1612, N1702);
nand NAND3 (N1720, N1713, N708, N121);
buf BUF1 (N1721, N1693);
xor XOR2 (N1722, N1719, N1547);
or OR2 (N1723, N1720, N790);
buf BUF1 (N1724, N1718);
xor XOR2 (N1725, N1711, N890);
xor XOR2 (N1726, N1725, N1551);
nor NOR2 (N1727, N1704, N1503);
and AND4 (N1728, N1721, N1055, N1586, N1123);
buf BUF1 (N1729, N1726);
buf BUF1 (N1730, N1714);
or OR2 (N1731, N1730, N246);
and AND3 (N1732, N1729, N640, N126);
buf BUF1 (N1733, N1716);
nor NOR4 (N1734, N1724, N1132, N968, N498);
or OR2 (N1735, N1732, N429);
and AND2 (N1736, N1733, N312);
nand NAND2 (N1737, N1723, N629);
not NOT1 (N1738, N1736);
nand NAND3 (N1739, N1728, N1101, N47);
buf BUF1 (N1740, N1707);
or OR4 (N1741, N1727, N814, N1131, N514);
and AND4 (N1742, N1739, N508, N307, N793);
nand NAND2 (N1743, N1740, N1080);
and AND3 (N1744, N1734, N1438, N85);
nor NOR2 (N1745, N1738, N929);
not NOT1 (N1746, N1722);
buf BUF1 (N1747, N1745);
and AND4 (N1748, N1742, N1682, N1241, N664);
or OR2 (N1749, N1744, N290);
not NOT1 (N1750, N1731);
nor NOR3 (N1751, N1737, N278, N394);
or OR4 (N1752, N1717, N825, N1522, N1147);
or OR3 (N1753, N1750, N731, N1387);
and AND2 (N1754, N1743, N727);
xor XOR2 (N1755, N1746, N498);
xor XOR2 (N1756, N1735, N1264);
nor NOR4 (N1757, N1753, N1352, N1476, N1687);
buf BUF1 (N1758, N1751);
buf BUF1 (N1759, N1741);
xor XOR2 (N1760, N1755, N661);
not NOT1 (N1761, N1748);
nor NOR3 (N1762, N1757, N1392, N321);
nor NOR2 (N1763, N1752, N1393);
xor XOR2 (N1764, N1756, N1750);
buf BUF1 (N1765, N1763);
xor XOR2 (N1766, N1760, N476);
xor XOR2 (N1767, N1762, N25);
nor NOR4 (N1768, N1754, N781, N430, N1081);
and AND3 (N1769, N1766, N1493, N596);
nand NAND4 (N1770, N1747, N357, N1511, N1065);
nor NOR2 (N1771, N1770, N772);
not NOT1 (N1772, N1759);
nand NAND3 (N1773, N1771, N1591, N431);
nand NAND3 (N1774, N1749, N92, N1602);
not NOT1 (N1775, N1774);
not NOT1 (N1776, N1767);
nor NOR3 (N1777, N1758, N668, N1436);
and AND4 (N1778, N1776, N604, N424, N544);
nor NOR3 (N1779, N1772, N180, N38);
xor XOR2 (N1780, N1779, N128);
or OR3 (N1781, N1778, N821, N717);
buf BUF1 (N1782, N1765);
or OR4 (N1783, N1780, N856, N833, N799);
xor XOR2 (N1784, N1777, N360);
xor XOR2 (N1785, N1761, N1112);
or OR2 (N1786, N1785, N299);
buf BUF1 (N1787, N1783);
not NOT1 (N1788, N1773);
xor XOR2 (N1789, N1764, N1661);
or OR3 (N1790, N1789, N1359, N1677);
and AND2 (N1791, N1784, N567);
nand NAND3 (N1792, N1788, N949, N1351);
nand NAND3 (N1793, N1769, N1107, N686);
buf BUF1 (N1794, N1787);
or OR4 (N1795, N1790, N966, N637, N1411);
and AND2 (N1796, N1786, N1719);
nor NOR3 (N1797, N1775, N1060, N380);
or OR4 (N1798, N1791, N906, N852, N1666);
nor NOR4 (N1799, N1768, N612, N1439, N575);
xor XOR2 (N1800, N1798, N1481);
nand NAND4 (N1801, N1796, N1181, N110, N1628);
nor NOR4 (N1802, N1801, N558, N468, N1623);
nand NAND3 (N1803, N1781, N1378, N1372);
and AND3 (N1804, N1800, N260, N729);
not NOT1 (N1805, N1795);
nand NAND2 (N1806, N1805, N373);
buf BUF1 (N1807, N1793);
buf BUF1 (N1808, N1803);
nor NOR4 (N1809, N1804, N1505, N1636, N417);
nor NOR3 (N1810, N1794, N219, N1527);
xor XOR2 (N1811, N1792, N1639);
nand NAND2 (N1812, N1799, N289);
or OR4 (N1813, N1808, N1032, N91, N319);
xor XOR2 (N1814, N1782, N338);
buf BUF1 (N1815, N1810);
nand NAND2 (N1816, N1814, N835);
nor NOR2 (N1817, N1811, N1143);
buf BUF1 (N1818, N1807);
and AND2 (N1819, N1816, N632);
buf BUF1 (N1820, N1818);
xor XOR2 (N1821, N1817, N1182);
buf BUF1 (N1822, N1821);
nand NAND4 (N1823, N1820, N1591, N1653, N607);
or OR3 (N1824, N1822, N965, N97);
xor XOR2 (N1825, N1815, N1077);
and AND3 (N1826, N1806, N1704, N728);
not NOT1 (N1827, N1823);
nand NAND3 (N1828, N1797, N211, N1532);
nand NAND2 (N1829, N1828, N178);
xor XOR2 (N1830, N1819, N374);
xor XOR2 (N1831, N1802, N1581);
or OR4 (N1832, N1826, N920, N1019, N22);
not NOT1 (N1833, N1831);
xor XOR2 (N1834, N1827, N458);
not NOT1 (N1835, N1812);
not NOT1 (N1836, N1832);
not NOT1 (N1837, N1824);
nand NAND2 (N1838, N1829, N1763);
or OR4 (N1839, N1838, N399, N337, N1151);
buf BUF1 (N1840, N1833);
nor NOR2 (N1841, N1834, N1073);
nand NAND3 (N1842, N1837, N1078, N883);
nand NAND3 (N1843, N1841, N897, N1496);
nand NAND3 (N1844, N1835, N1290, N455);
xor XOR2 (N1845, N1839, N1683);
buf BUF1 (N1846, N1825);
buf BUF1 (N1847, N1830);
buf BUF1 (N1848, N1843);
not NOT1 (N1849, N1847);
and AND4 (N1850, N1809, N1006, N1366, N1504);
and AND3 (N1851, N1836, N998, N558);
or OR4 (N1852, N1840, N1655, N1101, N1193);
nor NOR4 (N1853, N1848, N1565, N1749, N1509);
and AND3 (N1854, N1813, N1593, N1676);
and AND3 (N1855, N1845, N69, N738);
buf BUF1 (N1856, N1849);
xor XOR2 (N1857, N1846, N910);
or OR3 (N1858, N1857, N1231, N1494);
buf BUF1 (N1859, N1855);
xor XOR2 (N1860, N1856, N1150);
xor XOR2 (N1861, N1854, N1400);
or OR2 (N1862, N1858, N1267);
xor XOR2 (N1863, N1860, N1204);
not NOT1 (N1864, N1853);
and AND3 (N1865, N1844, N1559, N1190);
xor XOR2 (N1866, N1863, N1804);
nor NOR2 (N1867, N1864, N697);
and AND2 (N1868, N1862, N1173);
buf BUF1 (N1869, N1867);
xor XOR2 (N1870, N1842, N173);
buf BUF1 (N1871, N1850);
xor XOR2 (N1872, N1852, N1088);
or OR3 (N1873, N1872, N367, N471);
nor NOR3 (N1874, N1866, N1465, N1105);
and AND2 (N1875, N1859, N293);
nand NAND3 (N1876, N1871, N1043, N1000);
nand NAND2 (N1877, N1865, N713);
xor XOR2 (N1878, N1876, N975);
nand NAND4 (N1879, N1870, N990, N500, N1252);
nor NOR3 (N1880, N1861, N814, N811);
not NOT1 (N1881, N1875);
nand NAND4 (N1882, N1877, N1018, N1794, N474);
xor XOR2 (N1883, N1874, N1019);
not NOT1 (N1884, N1883);
nor NOR2 (N1885, N1881, N541);
not NOT1 (N1886, N1885);
buf BUF1 (N1887, N1868);
or OR4 (N1888, N1869, N930, N1475, N1845);
and AND3 (N1889, N1851, N1826, N668);
xor XOR2 (N1890, N1884, N1092);
and AND4 (N1891, N1886, N439, N1359, N475);
buf BUF1 (N1892, N1891);
or OR3 (N1893, N1890, N1006, N80);
or OR4 (N1894, N1889, N723, N995, N186);
buf BUF1 (N1895, N1878);
and AND2 (N1896, N1893, N1136);
or OR4 (N1897, N1894, N1645, N1499, N1610);
xor XOR2 (N1898, N1879, N490);
or OR2 (N1899, N1888, N735);
not NOT1 (N1900, N1892);
nor NOR3 (N1901, N1896, N1675, N210);
and AND3 (N1902, N1895, N677, N915);
not NOT1 (N1903, N1899);
nand NAND4 (N1904, N1882, N71, N316, N1467);
xor XOR2 (N1905, N1903, N912);
nand NAND3 (N1906, N1905, N1822, N463);
nor NOR3 (N1907, N1897, N739, N1467);
not NOT1 (N1908, N1880);
and AND4 (N1909, N1906, N1188, N1843, N1200);
or OR3 (N1910, N1900, N3, N1140);
nand NAND4 (N1911, N1907, N1108, N1195, N655);
not NOT1 (N1912, N1910);
buf BUF1 (N1913, N1912);
buf BUF1 (N1914, N1911);
not NOT1 (N1915, N1898);
buf BUF1 (N1916, N1902);
and AND4 (N1917, N1914, N1625, N1849, N269);
not NOT1 (N1918, N1916);
nor NOR2 (N1919, N1918, N1390);
or OR2 (N1920, N1915, N1145);
buf BUF1 (N1921, N1873);
or OR4 (N1922, N1904, N1130, N765, N1318);
or OR3 (N1923, N1887, N833, N1127);
or OR3 (N1924, N1909, N535, N244);
xor XOR2 (N1925, N1922, N1409);
or OR4 (N1926, N1923, N32, N1516, N1652);
buf BUF1 (N1927, N1919);
not NOT1 (N1928, N1926);
nand NAND4 (N1929, N1920, N1432, N989, N726);
buf BUF1 (N1930, N1908);
buf BUF1 (N1931, N1921);
and AND4 (N1932, N1927, N454, N19, N1729);
buf BUF1 (N1933, N1932);
not NOT1 (N1934, N1913);
nor NOR4 (N1935, N1931, N1336, N1858, N1621);
nor NOR2 (N1936, N1924, N613);
nor NOR3 (N1937, N1901, N327, N518);
or OR2 (N1938, N1934, N1721);
nor NOR4 (N1939, N1930, N446, N1733, N758);
not NOT1 (N1940, N1929);
or OR2 (N1941, N1935, N952);
nor NOR2 (N1942, N1940, N925);
buf BUF1 (N1943, N1938);
nor NOR3 (N1944, N1937, N713, N445);
nand NAND2 (N1945, N1944, N1639);
and AND3 (N1946, N1941, N503, N522);
or OR3 (N1947, N1925, N885, N1674);
buf BUF1 (N1948, N1928);
nand NAND4 (N1949, N1936, N318, N981, N1004);
not NOT1 (N1950, N1945);
and AND4 (N1951, N1942, N488, N1869, N535);
or OR3 (N1952, N1939, N1339, N970);
xor XOR2 (N1953, N1950, N1696);
or OR2 (N1954, N1946, N1278);
nand NAND4 (N1955, N1952, N1504, N1198, N118);
xor XOR2 (N1956, N1953, N1042);
nand NAND3 (N1957, N1943, N116, N1190);
nor NOR3 (N1958, N1917, N1363, N466);
nand NAND3 (N1959, N1956, N1389, N4);
nor NOR4 (N1960, N1947, N1287, N224, N1618);
buf BUF1 (N1961, N1933);
not NOT1 (N1962, N1955);
not NOT1 (N1963, N1962);
and AND3 (N1964, N1957, N1485, N246);
or OR3 (N1965, N1964, N18, N1197);
not NOT1 (N1966, N1958);
nand NAND4 (N1967, N1959, N879, N1397, N1488);
xor XOR2 (N1968, N1965, N751);
nor NOR2 (N1969, N1948, N1090);
nor NOR3 (N1970, N1966, N650, N847);
buf BUF1 (N1971, N1963);
nor NOR2 (N1972, N1967, N1892);
nor NOR2 (N1973, N1960, N1884);
or OR2 (N1974, N1971, N1693);
or OR2 (N1975, N1961, N1706);
and AND3 (N1976, N1951, N1704, N530);
buf BUF1 (N1977, N1949);
nand NAND4 (N1978, N1976, N1013, N100, N1323);
nand NAND2 (N1979, N1973, N294);
not NOT1 (N1980, N1969);
buf BUF1 (N1981, N1980);
buf BUF1 (N1982, N1968);
or OR4 (N1983, N1974, N1136, N659, N947);
not NOT1 (N1984, N1983);
xor XOR2 (N1985, N1975, N310);
xor XOR2 (N1986, N1982, N597);
buf BUF1 (N1987, N1985);
or OR3 (N1988, N1977, N1778, N1180);
not NOT1 (N1989, N1972);
not NOT1 (N1990, N1989);
buf BUF1 (N1991, N1981);
nand NAND3 (N1992, N1988, N1439, N706);
buf BUF1 (N1993, N1990);
xor XOR2 (N1994, N1970, N426);
and AND4 (N1995, N1992, N1167, N11, N1232);
nand NAND2 (N1996, N1993, N500);
nand NAND4 (N1997, N1979, N142, N1212, N477);
not NOT1 (N1998, N1984);
or OR4 (N1999, N1978, N139, N1872, N933);
and AND4 (N2000, N1987, N1694, N955, N1107);
nor NOR3 (N2001, N1995, N1682, N1487);
xor XOR2 (N2002, N1999, N522);
or OR3 (N2003, N1954, N1760, N1262);
nor NOR3 (N2004, N1996, N1109, N64);
and AND2 (N2005, N2001, N760);
or OR3 (N2006, N1997, N911, N1072);
xor XOR2 (N2007, N2002, N900);
nand NAND2 (N2008, N2004, N633);
buf BUF1 (N2009, N2008);
or OR4 (N2010, N2007, N499, N1011, N1367);
nand NAND3 (N2011, N1991, N1620, N1973);
nand NAND4 (N2012, N2003, N1704, N1475, N441);
and AND3 (N2013, N2000, N957, N1563);
nor NOR3 (N2014, N1998, N1881, N1450);
nor NOR3 (N2015, N2012, N1182, N1673);
xor XOR2 (N2016, N1994, N257);
buf BUF1 (N2017, N1986);
nand NAND2 (N2018, N2015, N197);
or OR2 (N2019, N2013, N750);
xor XOR2 (N2020, N2014, N284);
buf BUF1 (N2021, N2019);
buf BUF1 (N2022, N2005);
not NOT1 (N2023, N2020);
not NOT1 (N2024, N2006);
xor XOR2 (N2025, N2018, N535);
and AND4 (N2026, N2023, N555, N130, N805);
buf BUF1 (N2027, N2021);
not NOT1 (N2028, N2026);
nand NAND4 (N2029, N2024, N1955, N1016, N1701);
nand NAND3 (N2030, N2010, N1598, N901);
not NOT1 (N2031, N2017);
or OR2 (N2032, N2031, N1693);
nand NAND4 (N2033, N2030, N1121, N802, N938);
not NOT1 (N2034, N2028);
nor NOR2 (N2035, N2027, N1227);
nand NAND3 (N2036, N2009, N906, N1449);
not NOT1 (N2037, N2032);
not NOT1 (N2038, N2011);
nand NAND3 (N2039, N2033, N1364, N2004);
xor XOR2 (N2040, N2029, N233);
nor NOR2 (N2041, N2035, N1841);
or OR2 (N2042, N2040, N169);
xor XOR2 (N2043, N2034, N306);
xor XOR2 (N2044, N2042, N618);
xor XOR2 (N2045, N2039, N673);
nand NAND2 (N2046, N2025, N785);
buf BUF1 (N2047, N2022);
not NOT1 (N2048, N2037);
or OR4 (N2049, N2048, N595, N855, N531);
nand NAND2 (N2050, N2041, N1346);
buf BUF1 (N2051, N2016);
xor XOR2 (N2052, N2036, N605);
nor NOR4 (N2053, N2038, N366, N1027, N1829);
nand NAND2 (N2054, N2047, N352);
nand NAND2 (N2055, N2052, N161);
or OR3 (N2056, N2055, N9, N965);
and AND2 (N2057, N2046, N1506);
and AND3 (N2058, N2044, N1273, N1805);
not NOT1 (N2059, N2056);
not NOT1 (N2060, N2057);
xor XOR2 (N2061, N2043, N236);
not NOT1 (N2062, N2050);
not NOT1 (N2063, N2060);
nor NOR4 (N2064, N2053, N1854, N1490, N1656);
not NOT1 (N2065, N2063);
buf BUF1 (N2066, N2062);
buf BUF1 (N2067, N2066);
and AND4 (N2068, N2051, N234, N1889, N1846);
or OR3 (N2069, N2058, N1277, N404);
buf BUF1 (N2070, N2064);
nand NAND3 (N2071, N2069, N2058, N128);
and AND3 (N2072, N2070, N1722, N786);
or OR4 (N2073, N2065, N826, N765, N716);
xor XOR2 (N2074, N2071, N1814);
nor NOR2 (N2075, N2061, N682);
nand NAND2 (N2076, N2068, N1809);
buf BUF1 (N2077, N2045);
nor NOR3 (N2078, N2049, N1132, N122);
buf BUF1 (N2079, N2059);
nand NAND4 (N2080, N2078, N415, N1534, N348);
and AND4 (N2081, N2076, N623, N1075, N268);
buf BUF1 (N2082, N2067);
not NOT1 (N2083, N2073);
nand NAND4 (N2084, N2077, N533, N999, N2014);
buf BUF1 (N2085, N2083);
nor NOR3 (N2086, N2074, N1490, N1229);
buf BUF1 (N2087, N2085);
nand NAND2 (N2088, N2075, N323);
or OR2 (N2089, N2082, N687);
nand NAND3 (N2090, N2079, N1638, N1405);
and AND2 (N2091, N2072, N1469);
nand NAND3 (N2092, N2054, N30, N931);
nand NAND4 (N2093, N2090, N779, N1078, N1633);
buf BUF1 (N2094, N2087);
buf BUF1 (N2095, N2094);
xor XOR2 (N2096, N2089, N496);
buf BUF1 (N2097, N2092);
not NOT1 (N2098, N2095);
nor NOR3 (N2099, N2098, N1187, N511);
and AND2 (N2100, N2081, N1285);
nor NOR3 (N2101, N2100, N821, N243);
nor NOR2 (N2102, N2093, N696);
and AND3 (N2103, N2088, N593, N77);
or OR2 (N2104, N2084, N34);
xor XOR2 (N2105, N2104, N2007);
nor NOR3 (N2106, N2103, N1774, N310);
buf BUF1 (N2107, N2101);
not NOT1 (N2108, N2102);
nor NOR4 (N2109, N2099, N1448, N1439, N717);
xor XOR2 (N2110, N2108, N1544);
or OR2 (N2111, N2109, N415);
or OR4 (N2112, N2097, N650, N1690, N750);
buf BUF1 (N2113, N2112);
nor NOR4 (N2114, N2113, N415, N713, N2078);
not NOT1 (N2115, N2106);
nand NAND2 (N2116, N2086, N934);
and AND4 (N2117, N2096, N493, N1250, N1355);
xor XOR2 (N2118, N2105, N927);
buf BUF1 (N2119, N2110);
xor XOR2 (N2120, N2107, N1825);
or OR3 (N2121, N2119, N1796, N857);
and AND4 (N2122, N2117, N1115, N1093, N2100);
not NOT1 (N2123, N2111);
or OR3 (N2124, N2114, N1235, N1084);
nor NOR3 (N2125, N2091, N1905, N914);
not NOT1 (N2126, N2125);
not NOT1 (N2127, N2120);
xor XOR2 (N2128, N2127, N605);
buf BUF1 (N2129, N2080);
nand NAND3 (N2130, N2118, N763, N1247);
not NOT1 (N2131, N2129);
not NOT1 (N2132, N2116);
buf BUF1 (N2133, N2122);
or OR4 (N2134, N2133, N1902, N625, N497);
or OR3 (N2135, N2115, N1894, N214);
and AND2 (N2136, N2124, N700);
xor XOR2 (N2137, N2132, N1228);
nor NOR2 (N2138, N2131, N347);
nor NOR4 (N2139, N2136, N1706, N382, N1042);
and AND2 (N2140, N2128, N305);
and AND4 (N2141, N2126, N233, N517, N1378);
xor XOR2 (N2142, N2135, N1779);
and AND2 (N2143, N2121, N311);
and AND2 (N2144, N2123, N2083);
not NOT1 (N2145, N2141);
nor NOR2 (N2146, N2143, N1860);
buf BUF1 (N2147, N2146);
buf BUF1 (N2148, N2145);
xor XOR2 (N2149, N2147, N1689);
nor NOR2 (N2150, N2139, N331);
or OR2 (N2151, N2149, N1934);
not NOT1 (N2152, N2144);
nand NAND4 (N2153, N2151, N325, N1587, N1076);
or OR4 (N2154, N2130, N2104, N813, N1277);
nor NOR2 (N2155, N2150, N653);
or OR4 (N2156, N2134, N2051, N667, N1964);
and AND2 (N2157, N2148, N93);
or OR2 (N2158, N2154, N811);
and AND4 (N2159, N2155, N558, N607, N1973);
not NOT1 (N2160, N2138);
nand NAND3 (N2161, N2140, N2064, N30);
or OR2 (N2162, N2160, N770);
or OR3 (N2163, N2159, N1520, N1451);
nor NOR4 (N2164, N2153, N784, N1426, N1790);
and AND4 (N2165, N2162, N765, N1571, N685);
xor XOR2 (N2166, N2165, N1675);
nand NAND4 (N2167, N2161, N292, N1938, N719);
not NOT1 (N2168, N2158);
xor XOR2 (N2169, N2167, N23);
nand NAND4 (N2170, N2157, N1338, N1108, N101);
not NOT1 (N2171, N2170);
buf BUF1 (N2172, N2152);
nand NAND2 (N2173, N2156, N167);
or OR3 (N2174, N2137, N1692, N33);
nand NAND4 (N2175, N2172, N1779, N989, N1813);
or OR3 (N2176, N2142, N1130, N1170);
nand NAND4 (N2177, N2171, N1938, N2094, N1202);
and AND4 (N2178, N2164, N461, N2014, N1851);
not NOT1 (N2179, N2175);
xor XOR2 (N2180, N2173, N1532);
nor NOR4 (N2181, N2169, N1074, N2074, N1168);
not NOT1 (N2182, N2176);
and AND4 (N2183, N2181, N998, N749, N1229);
xor XOR2 (N2184, N2166, N2182);
not NOT1 (N2185, N1628);
nor NOR3 (N2186, N2178, N1561, N593);
xor XOR2 (N2187, N2177, N2022);
xor XOR2 (N2188, N2163, N765);
not NOT1 (N2189, N2180);
and AND4 (N2190, N2189, N1932, N2094, N723);
not NOT1 (N2191, N2168);
nor NOR4 (N2192, N2186, N230, N1576, N1838);
xor XOR2 (N2193, N2183, N1093);
and AND3 (N2194, N2190, N1612, N1881);
not NOT1 (N2195, N2184);
nor NOR3 (N2196, N2191, N785, N593);
nand NAND4 (N2197, N2174, N969, N36, N1946);
nand NAND2 (N2198, N2195, N1449);
nor NOR4 (N2199, N2197, N1541, N422, N2011);
or OR2 (N2200, N2199, N1468);
and AND2 (N2201, N2194, N1875);
or OR4 (N2202, N2200, N1812, N281, N788);
nor NOR3 (N2203, N2192, N601, N861);
and AND2 (N2204, N2188, N169);
xor XOR2 (N2205, N2185, N27);
not NOT1 (N2206, N2204);
xor XOR2 (N2207, N2179, N1162);
not NOT1 (N2208, N2198);
buf BUF1 (N2209, N2206);
buf BUF1 (N2210, N2205);
nor NOR2 (N2211, N2187, N234);
or OR3 (N2212, N2208, N2074, N826);
buf BUF1 (N2213, N2196);
nor NOR2 (N2214, N2209, N447);
buf BUF1 (N2215, N2211);
or OR4 (N2216, N2210, N571, N776, N502);
xor XOR2 (N2217, N2212, N334);
and AND3 (N2218, N2203, N1657, N418);
or OR4 (N2219, N2216, N1408, N1732, N1727);
xor XOR2 (N2220, N2218, N609);
or OR4 (N2221, N2214, N261, N1599, N618);
nand NAND4 (N2222, N2220, N1923, N1140, N247);
nand NAND3 (N2223, N2193, N1273, N1536);
buf BUF1 (N2224, N2213);
xor XOR2 (N2225, N2221, N1072);
buf BUF1 (N2226, N2223);
nand NAND4 (N2227, N2219, N783, N973, N1399);
or OR3 (N2228, N2217, N2076, N33);
nor NOR3 (N2229, N2222, N151, N1370);
nand NAND2 (N2230, N2228, N739);
not NOT1 (N2231, N2201);
and AND2 (N2232, N2225, N1524);
nand NAND4 (N2233, N2231, N1604, N128, N1415);
nor NOR2 (N2234, N2229, N13);
not NOT1 (N2235, N2227);
and AND3 (N2236, N2207, N333, N2213);
not NOT1 (N2237, N2236);
nand NAND3 (N2238, N2226, N1335, N1230);
buf BUF1 (N2239, N2215);
nand NAND3 (N2240, N2224, N1849, N379);
not NOT1 (N2241, N2232);
buf BUF1 (N2242, N2240);
not NOT1 (N2243, N2242);
and AND4 (N2244, N2233, N252, N1273, N2118);
not NOT1 (N2245, N2239);
nand NAND4 (N2246, N2243, N252, N160, N1140);
not NOT1 (N2247, N2238);
buf BUF1 (N2248, N2235);
nand NAND3 (N2249, N2246, N2207, N950);
or OR4 (N2250, N2202, N531, N378, N1256);
xor XOR2 (N2251, N2234, N765);
not NOT1 (N2252, N2245);
nand NAND4 (N2253, N2241, N877, N126, N184);
buf BUF1 (N2254, N2253);
and AND2 (N2255, N2249, N2127);
not NOT1 (N2256, N2237);
and AND4 (N2257, N2256, N1200, N1436, N1924);
xor XOR2 (N2258, N2252, N1214);
buf BUF1 (N2259, N2230);
buf BUF1 (N2260, N2244);
not NOT1 (N2261, N2260);
nand NAND4 (N2262, N2261, N1933, N1828, N378);
nand NAND2 (N2263, N2258, N2027);
buf BUF1 (N2264, N2254);
not NOT1 (N2265, N2251);
nor NOR4 (N2266, N2265, N943, N444, N994);
xor XOR2 (N2267, N2255, N1610);
not NOT1 (N2268, N2247);
xor XOR2 (N2269, N2267, N560);
nor NOR2 (N2270, N2266, N973);
nor NOR4 (N2271, N2270, N249, N398, N103);
xor XOR2 (N2272, N2271, N1612);
xor XOR2 (N2273, N2259, N1920);
nand NAND3 (N2274, N2269, N2191, N329);
and AND2 (N2275, N2248, N1849);
buf BUF1 (N2276, N2263);
and AND4 (N2277, N2268, N865, N591, N1630);
or OR2 (N2278, N2257, N1960);
and AND4 (N2279, N2277, N1991, N724, N1183);
and AND3 (N2280, N2250, N18, N1979);
xor XOR2 (N2281, N2264, N1647);
or OR3 (N2282, N2276, N1966, N1337);
nor NOR4 (N2283, N2275, N1003, N780, N281);
not NOT1 (N2284, N2272);
nand NAND4 (N2285, N2278, N1709, N1588, N1495);
buf BUF1 (N2286, N2282);
nor NOR4 (N2287, N2284, N294, N1780, N2096);
not NOT1 (N2288, N2287);
nor NOR3 (N2289, N2281, N363, N867);
nand NAND3 (N2290, N2279, N2036, N2239);
not NOT1 (N2291, N2280);
not NOT1 (N2292, N2283);
xor XOR2 (N2293, N2273, N730);
and AND3 (N2294, N2293, N728, N898);
xor XOR2 (N2295, N2286, N735);
buf BUF1 (N2296, N2292);
nand NAND2 (N2297, N2291, N1485);
or OR2 (N2298, N2262, N365);
nor NOR2 (N2299, N2274, N2151);
not NOT1 (N2300, N2285);
nand NAND3 (N2301, N2296, N238, N444);
not NOT1 (N2302, N2297);
nor NOR3 (N2303, N2294, N2210, N567);
nor NOR3 (N2304, N2302, N1314, N323);
and AND2 (N2305, N2289, N7);
xor XOR2 (N2306, N2303, N1342);
or OR3 (N2307, N2305, N1047, N271);
and AND2 (N2308, N2300, N2292);
nor NOR3 (N2309, N2301, N1870, N1136);
not NOT1 (N2310, N2308);
and AND2 (N2311, N2304, N1924);
nand NAND4 (N2312, N2290, N2187, N2267, N2173);
buf BUF1 (N2313, N2306);
buf BUF1 (N2314, N2312);
nand NAND4 (N2315, N2295, N488, N321, N2061);
buf BUF1 (N2316, N2307);
nor NOR4 (N2317, N2309, N429, N1870, N604);
buf BUF1 (N2318, N2299);
and AND2 (N2319, N2311, N586);
xor XOR2 (N2320, N2315, N550);
buf BUF1 (N2321, N2320);
or OR4 (N2322, N2314, N1136, N869, N610);
nor NOR2 (N2323, N2310, N880);
nand NAND4 (N2324, N2298, N76, N997, N1247);
nor NOR2 (N2325, N2321, N842);
not NOT1 (N2326, N2323);
nor NOR2 (N2327, N2317, N567);
not NOT1 (N2328, N2316);
buf BUF1 (N2329, N2324);
not NOT1 (N2330, N2326);
nor NOR4 (N2331, N2319, N458, N1445, N89);
not NOT1 (N2332, N2331);
buf BUF1 (N2333, N2332);
not NOT1 (N2334, N2313);
nor NOR4 (N2335, N2334, N708, N1093, N272);
nand NAND3 (N2336, N2330, N45, N887);
buf BUF1 (N2337, N2318);
not NOT1 (N2338, N2322);
xor XOR2 (N2339, N2329, N2089);
and AND4 (N2340, N2325, N155, N768, N1510);
buf BUF1 (N2341, N2340);
or OR2 (N2342, N2337, N1856);
and AND3 (N2343, N2339, N765, N2105);
nor NOR2 (N2344, N2335, N1377);
nor NOR3 (N2345, N2344, N1795, N186);
buf BUF1 (N2346, N2343);
or OR4 (N2347, N2288, N462, N220, N1205);
xor XOR2 (N2348, N2327, N2006);
buf BUF1 (N2349, N2338);
or OR4 (N2350, N2349, N738, N1889, N2045);
nor NOR4 (N2351, N2350, N158, N241, N1877);
and AND4 (N2352, N2347, N1116, N1088, N267);
nor NOR2 (N2353, N2328, N1575);
not NOT1 (N2354, N2353);
and AND2 (N2355, N2333, N54);
xor XOR2 (N2356, N2351, N834);
xor XOR2 (N2357, N2348, N118);
nor NOR2 (N2358, N2341, N2073);
nand NAND3 (N2359, N2336, N70, N1131);
xor XOR2 (N2360, N2346, N262);
buf BUF1 (N2361, N2358);
nand NAND4 (N2362, N2357, N445, N263, N1766);
not NOT1 (N2363, N2345);
xor XOR2 (N2364, N2362, N40);
nor NOR4 (N2365, N2359, N1511, N131, N173);
not NOT1 (N2366, N2342);
buf BUF1 (N2367, N2361);
nand NAND2 (N2368, N2360, N1417);
nor NOR2 (N2369, N2367, N1308);
and AND3 (N2370, N2364, N1806, N1443);
or OR3 (N2371, N2369, N135, N408);
and AND4 (N2372, N2365, N144, N116, N2323);
not NOT1 (N2373, N2355);
and AND2 (N2374, N2366, N1362);
and AND2 (N2375, N2368, N1393);
nand NAND3 (N2376, N2352, N971, N868);
nand NAND2 (N2377, N2373, N157);
and AND3 (N2378, N2374, N349, N2311);
buf BUF1 (N2379, N2370);
not NOT1 (N2380, N2356);
and AND3 (N2381, N2371, N1283, N116);
not NOT1 (N2382, N2379);
and AND4 (N2383, N2375, N447, N550, N2004);
xor XOR2 (N2384, N2383, N880);
and AND3 (N2385, N2372, N1103, N258);
nand NAND2 (N2386, N2354, N708);
nand NAND2 (N2387, N2380, N127);
nand NAND2 (N2388, N2377, N43);
nand NAND4 (N2389, N2386, N1898, N771, N618);
xor XOR2 (N2390, N2388, N1053);
nor NOR2 (N2391, N2387, N513);
nor NOR3 (N2392, N2384, N2301, N1395);
buf BUF1 (N2393, N2363);
nor NOR2 (N2394, N2391, N168);
not NOT1 (N2395, N2382);
nand NAND3 (N2396, N2392, N299, N805);
nand NAND2 (N2397, N2376, N659);
or OR3 (N2398, N2397, N2223, N1260);
nand NAND4 (N2399, N2398, N1415, N1389, N1381);
or OR2 (N2400, N2381, N836);
and AND2 (N2401, N2393, N1652);
not NOT1 (N2402, N2395);
nor NOR4 (N2403, N2402, N2053, N967, N45);
xor XOR2 (N2404, N2390, N212);
nand NAND2 (N2405, N2396, N634);
nand NAND3 (N2406, N2385, N32, N35);
nor NOR4 (N2407, N2401, N795, N1056, N1062);
not NOT1 (N2408, N2389);
nor NOR4 (N2409, N2394, N736, N1295, N1254);
nor NOR2 (N2410, N2405, N431);
not NOT1 (N2411, N2409);
buf BUF1 (N2412, N2410);
or OR2 (N2413, N2407, N2018);
buf BUF1 (N2414, N2404);
and AND4 (N2415, N2414, N769, N2198, N1320);
or OR3 (N2416, N2411, N2398, N1831);
buf BUF1 (N2417, N2400);
nand NAND3 (N2418, N2399, N1477, N1615);
and AND2 (N2419, N2415, N530);
and AND3 (N2420, N2418, N2259, N2291);
not NOT1 (N2421, N2406);
buf BUF1 (N2422, N2417);
buf BUF1 (N2423, N2421);
or OR4 (N2424, N2403, N892, N330, N849);
nor NOR2 (N2425, N2419, N1863);
and AND3 (N2426, N2420, N769, N963);
or OR4 (N2427, N2413, N213, N1206, N649);
nor NOR3 (N2428, N2378, N641, N1941);
nor NOR2 (N2429, N2423, N952);
nand NAND2 (N2430, N2416, N92);
and AND2 (N2431, N2422, N173);
nor NOR4 (N2432, N2426, N1211, N1228, N463);
nor NOR3 (N2433, N2430, N955, N1243);
nor NOR2 (N2434, N2425, N286);
or OR3 (N2435, N2428, N545, N480);
xor XOR2 (N2436, N2424, N792);
nand NAND4 (N2437, N2412, N1964, N1672, N1452);
xor XOR2 (N2438, N2427, N1586);
not NOT1 (N2439, N2435);
xor XOR2 (N2440, N2432, N2354);
and AND4 (N2441, N2440, N733, N2261, N793);
nor NOR2 (N2442, N2434, N1255);
or OR3 (N2443, N2439, N427, N1129);
and AND2 (N2444, N2443, N22);
nor NOR3 (N2445, N2429, N1916, N1153);
nor NOR4 (N2446, N2445, N1961, N554, N2239);
and AND3 (N2447, N2438, N750, N668);
nand NAND2 (N2448, N2431, N1583);
and AND4 (N2449, N2436, N992, N2333, N2442);
buf BUF1 (N2450, N484);
buf BUF1 (N2451, N2433);
nand NAND3 (N2452, N2446, N318, N399);
or OR3 (N2453, N2450, N1964, N908);
nand NAND3 (N2454, N2451, N92, N1419);
buf BUF1 (N2455, N2447);
or OR4 (N2456, N2449, N1858, N1848, N1871);
nand NAND4 (N2457, N2453, N174, N2166, N1382);
nor NOR3 (N2458, N2437, N54, N637);
or OR2 (N2459, N2408, N582);
xor XOR2 (N2460, N2452, N1737);
xor XOR2 (N2461, N2458, N2213);
nand NAND4 (N2462, N2461, N1565, N1164, N2291);
nand NAND2 (N2463, N2462, N1942);
xor XOR2 (N2464, N2459, N621);
not NOT1 (N2465, N2463);
buf BUF1 (N2466, N2465);
and AND2 (N2467, N2448, N1908);
nor NOR3 (N2468, N2460, N1174, N1974);
and AND3 (N2469, N2468, N1176, N353);
buf BUF1 (N2470, N2466);
and AND3 (N2471, N2467, N2159, N1142);
xor XOR2 (N2472, N2444, N1051);
not NOT1 (N2473, N2470);
buf BUF1 (N2474, N2457);
nor NOR4 (N2475, N2464, N723, N1206, N229);
buf BUF1 (N2476, N2475);
xor XOR2 (N2477, N2474, N843);
nand NAND3 (N2478, N2472, N1439, N1507);
and AND2 (N2479, N2473, N1139);
nand NAND2 (N2480, N2469, N1536);
not NOT1 (N2481, N2476);
and AND4 (N2482, N2481, N1455, N1414, N1000);
buf BUF1 (N2483, N2441);
or OR4 (N2484, N2477, N1851, N1266, N2450);
nand NAND2 (N2485, N2480, N2445);
nand NAND3 (N2486, N2483, N2048, N1819);
nand NAND4 (N2487, N2482, N428, N435, N536);
and AND4 (N2488, N2456, N1527, N1502, N418);
and AND3 (N2489, N2487, N7, N1939);
nor NOR4 (N2490, N2454, N2343, N591, N1142);
nor NOR3 (N2491, N2484, N1480, N886);
nor NOR2 (N2492, N2489, N716);
and AND3 (N2493, N2485, N2215, N1731);
nor NOR4 (N2494, N2490, N354, N54, N1539);
not NOT1 (N2495, N2488);
nand NAND2 (N2496, N2478, N1504);
not NOT1 (N2497, N2496);
and AND4 (N2498, N2497, N1289, N1496, N1984);
or OR3 (N2499, N2493, N2282, N165);
xor XOR2 (N2500, N2486, N550);
xor XOR2 (N2501, N2498, N1536);
or OR3 (N2502, N2494, N519, N1657);
nor NOR2 (N2503, N2471, N902);
buf BUF1 (N2504, N2500);
not NOT1 (N2505, N2502);
and AND4 (N2506, N2495, N1236, N1076, N1250);
nor NOR2 (N2507, N2504, N2459);
or OR4 (N2508, N2503, N1222, N360, N37);
nor NOR2 (N2509, N2491, N1061);
and AND2 (N2510, N2501, N2263);
nor NOR4 (N2511, N2506, N2071, N3, N1506);
nand NAND3 (N2512, N2510, N803, N1654);
nor NOR2 (N2513, N2499, N1323);
xor XOR2 (N2514, N2455, N1578);
buf BUF1 (N2515, N2511);
nand NAND2 (N2516, N2492, N1723);
nor NOR2 (N2517, N2516, N647);
not NOT1 (N2518, N2514);
or OR4 (N2519, N2509, N1076, N1885, N741);
buf BUF1 (N2520, N2505);
nand NAND2 (N2521, N2508, N169);
or OR2 (N2522, N2519, N2332);
not NOT1 (N2523, N2520);
buf BUF1 (N2524, N2517);
nor NOR2 (N2525, N2524, N2101);
not NOT1 (N2526, N2512);
buf BUF1 (N2527, N2518);
and AND4 (N2528, N2479, N1920, N948, N1783);
nand NAND2 (N2529, N2528, N2358);
or OR4 (N2530, N2515, N572, N2209, N486);
and AND2 (N2531, N2513, N760);
not NOT1 (N2532, N2525);
xor XOR2 (N2533, N2527, N1562);
nor NOR3 (N2534, N2531, N727, N643);
buf BUF1 (N2535, N2530);
not NOT1 (N2536, N2523);
nor NOR3 (N2537, N2522, N1642, N2483);
not NOT1 (N2538, N2536);
nor NOR3 (N2539, N2538, N2400, N1950);
not NOT1 (N2540, N2521);
nand NAND4 (N2541, N2532, N790, N2458, N2428);
nor NOR3 (N2542, N2534, N522, N398);
buf BUF1 (N2543, N2537);
nor NOR3 (N2544, N2535, N1640, N1125);
not NOT1 (N2545, N2526);
nand NAND3 (N2546, N2539, N1266, N2227);
not NOT1 (N2547, N2544);
and AND3 (N2548, N2542, N265, N2408);
xor XOR2 (N2549, N2546, N561);
or OR4 (N2550, N2543, N1792, N1346, N1850);
xor XOR2 (N2551, N2540, N1607);
not NOT1 (N2552, N2507);
nand NAND4 (N2553, N2533, N2361, N870, N701);
or OR2 (N2554, N2548, N47);
or OR4 (N2555, N2551, N931, N1922, N1004);
xor XOR2 (N2556, N2529, N1959);
nand NAND2 (N2557, N2545, N1819);
not NOT1 (N2558, N2557);
and AND3 (N2559, N2541, N141, N631);
or OR3 (N2560, N2555, N199, N599);
nand NAND4 (N2561, N2556, N1657, N2379, N2090);
and AND2 (N2562, N2561, N368);
xor XOR2 (N2563, N2553, N1670);
not NOT1 (N2564, N2560);
xor XOR2 (N2565, N2559, N460);
nor NOR4 (N2566, N2562, N2070, N1995, N2056);
or OR3 (N2567, N2565, N1265, N2271);
xor XOR2 (N2568, N2558, N399);
nor NOR4 (N2569, N2549, N2285, N461, N2035);
nor NOR4 (N2570, N2567, N2133, N938, N993);
or OR3 (N2571, N2550, N1131, N1595);
not NOT1 (N2572, N2566);
nand NAND4 (N2573, N2572, N109, N2078, N1435);
or OR4 (N2574, N2554, N2435, N794, N891);
buf BUF1 (N2575, N2570);
xor XOR2 (N2576, N2569, N320);
nand NAND4 (N2577, N2547, N1888, N1832, N2549);
xor XOR2 (N2578, N2568, N1530);
nor NOR3 (N2579, N2576, N2238, N782);
buf BUF1 (N2580, N2577);
nand NAND2 (N2581, N2574, N2238);
buf BUF1 (N2582, N2563);
nand NAND4 (N2583, N2579, N1203, N2267, N1837);
not NOT1 (N2584, N2580);
xor XOR2 (N2585, N2573, N253);
xor XOR2 (N2586, N2552, N2584);
or OR4 (N2587, N2234, N1971, N523, N1769);
not NOT1 (N2588, N2587);
or OR4 (N2589, N2582, N1628, N2459, N1747);
and AND3 (N2590, N2585, N1717, N71);
or OR4 (N2591, N2581, N2525, N198, N86);
or OR3 (N2592, N2586, N1210, N51);
not NOT1 (N2593, N2578);
not NOT1 (N2594, N2564);
and AND2 (N2595, N2592, N2243);
and AND4 (N2596, N2593, N2380, N1571, N470);
xor XOR2 (N2597, N2594, N1155);
and AND2 (N2598, N2571, N963);
not NOT1 (N2599, N2589);
or OR2 (N2600, N2591, N2467);
nand NAND4 (N2601, N2596, N262, N1793, N2135);
buf BUF1 (N2602, N2598);
buf BUF1 (N2603, N2588);
nand NAND4 (N2604, N2583, N506, N1241, N823);
buf BUF1 (N2605, N2603);
nor NOR2 (N2606, N2602, N2142);
not NOT1 (N2607, N2600);
and AND3 (N2608, N2606, N850, N2470);
xor XOR2 (N2609, N2604, N1118);
nor NOR4 (N2610, N2575, N2349, N1427, N844);
nor NOR3 (N2611, N2601, N1414, N1631);
nor NOR2 (N2612, N2599, N484);
xor XOR2 (N2613, N2605, N656);
nand NAND3 (N2614, N2607, N709, N1208);
buf BUF1 (N2615, N2597);
nor NOR2 (N2616, N2590, N2613);
not NOT1 (N2617, N2578);
nor NOR3 (N2618, N2611, N2474, N515);
nor NOR3 (N2619, N2612, N2128, N2532);
and AND2 (N2620, N2595, N80);
buf BUF1 (N2621, N2616);
not NOT1 (N2622, N2609);
and AND2 (N2623, N2614, N1365);
nand NAND3 (N2624, N2621, N2145, N458);
or OR4 (N2625, N2622, N1201, N2525, N186);
xor XOR2 (N2626, N2608, N407);
xor XOR2 (N2627, N2617, N1994);
nand NAND4 (N2628, N2623, N1336, N1840, N903);
xor XOR2 (N2629, N2628, N2400);
and AND3 (N2630, N2625, N373, N630);
nor NOR4 (N2631, N2615, N1101, N634, N1871);
or OR4 (N2632, N2624, N567, N1861, N1730);
nand NAND2 (N2633, N2631, N1010);
not NOT1 (N2634, N2629);
not NOT1 (N2635, N2610);
nand NAND3 (N2636, N2634, N2158, N1155);
xor XOR2 (N2637, N2633, N909);
xor XOR2 (N2638, N2627, N1973);
or OR4 (N2639, N2618, N1263, N820, N102);
or OR4 (N2640, N2632, N988, N807, N2639);
xor XOR2 (N2641, N2360, N853);
nand NAND3 (N2642, N2626, N1389, N473);
and AND4 (N2643, N2642, N1745, N883, N2543);
nor NOR4 (N2644, N2637, N2013, N1240, N1351);
nor NOR2 (N2645, N2619, N1452);
nand NAND4 (N2646, N2645, N451, N1875, N1908);
nor NOR4 (N2647, N2646, N739, N1209, N1513);
or OR4 (N2648, N2640, N1332, N2132, N1992);
nand NAND4 (N2649, N2635, N328, N634, N393);
nor NOR4 (N2650, N2620, N1173, N366, N601);
xor XOR2 (N2651, N2638, N2056);
buf BUF1 (N2652, N2651);
not NOT1 (N2653, N2648);
and AND4 (N2654, N2636, N1462, N66, N2235);
nand NAND2 (N2655, N2652, N1976);
nor NOR4 (N2656, N2630, N834, N2238, N1553);
and AND3 (N2657, N2647, N196, N793);
not NOT1 (N2658, N2654);
or OR2 (N2659, N2649, N1442);
xor XOR2 (N2660, N2658, N1891);
nand NAND2 (N2661, N2644, N2227);
xor XOR2 (N2662, N2650, N239);
and AND2 (N2663, N2641, N2494);
nand NAND2 (N2664, N2655, N1710);
or OR2 (N2665, N2660, N1507);
nor NOR2 (N2666, N2653, N1095);
xor XOR2 (N2667, N2664, N2570);
buf BUF1 (N2668, N2657);
and AND2 (N2669, N2667, N277);
and AND2 (N2670, N2668, N2526);
nor NOR4 (N2671, N2661, N977, N916, N1868);
xor XOR2 (N2672, N2671, N1251);
and AND3 (N2673, N2670, N1409, N1840);
or OR3 (N2674, N2672, N20, N1312);
not NOT1 (N2675, N2669);
not NOT1 (N2676, N2674);
nand NAND2 (N2677, N2663, N2406);
or OR3 (N2678, N2676, N330, N1865);
nand NAND2 (N2679, N2643, N1553);
nand NAND3 (N2680, N2666, N1308, N2027);
or OR3 (N2681, N2677, N17, N136);
nor NOR2 (N2682, N2678, N807);
and AND3 (N2683, N2659, N2628, N2097);
or OR4 (N2684, N2673, N2467, N1400, N2484);
nand NAND3 (N2685, N2682, N2642, N1890);
nor NOR4 (N2686, N2685, N2001, N2107, N2509);
not NOT1 (N2687, N2675);
nand NAND2 (N2688, N2656, N2132);
or OR4 (N2689, N2681, N1075, N1453, N109);
nor NOR2 (N2690, N2665, N300);
and AND3 (N2691, N2686, N1952, N1008);
xor XOR2 (N2692, N2680, N349);
xor XOR2 (N2693, N2689, N1663);
not NOT1 (N2694, N2683);
nand NAND2 (N2695, N2691, N1415);
not NOT1 (N2696, N2688);
or OR2 (N2697, N2692, N2424);
or OR3 (N2698, N2684, N623, N423);
buf BUF1 (N2699, N2696);
or OR4 (N2700, N2693, N1680, N2465, N2690);
or OR3 (N2701, N954, N2687, N1998);
and AND2 (N2702, N1506, N488);
xor XOR2 (N2703, N2694, N2093);
nand NAND4 (N2704, N2700, N109, N1829, N463);
nand NAND2 (N2705, N2703, N2452);
xor XOR2 (N2706, N2699, N1530);
buf BUF1 (N2707, N2679);
buf BUF1 (N2708, N2662);
xor XOR2 (N2709, N2708, N1006);
and AND4 (N2710, N2705, N788, N344, N1602);
xor XOR2 (N2711, N2701, N701);
xor XOR2 (N2712, N2709, N493);
buf BUF1 (N2713, N2697);
nor NOR3 (N2714, N2710, N1135, N205);
not NOT1 (N2715, N2698);
nand NAND3 (N2716, N2712, N646, N1225);
xor XOR2 (N2717, N2713, N1220);
and AND2 (N2718, N2706, N2717);
and AND3 (N2719, N1040, N1606, N67);
buf BUF1 (N2720, N2704);
and AND3 (N2721, N2720, N907, N1001);
nand NAND4 (N2722, N2702, N1, N2713, N1794);
or OR4 (N2723, N2711, N491, N2053, N549);
nor NOR2 (N2724, N2721, N229);
and AND2 (N2725, N2718, N1898);
nand NAND4 (N2726, N2707, N1317, N1911, N2144);
or OR3 (N2727, N2716, N1904, N2185);
not NOT1 (N2728, N2714);
nand NAND3 (N2729, N2719, N2569, N2239);
and AND4 (N2730, N2725, N2376, N2151, N1529);
not NOT1 (N2731, N2723);
xor XOR2 (N2732, N2731, N282);
and AND2 (N2733, N2728, N981);
not NOT1 (N2734, N2715);
xor XOR2 (N2735, N2730, N1101);
nor NOR4 (N2736, N2727, N1501, N1958, N1126);
not NOT1 (N2737, N2722);
buf BUF1 (N2738, N2733);
nand NAND4 (N2739, N2732, N2165, N1110, N1553);
nor NOR3 (N2740, N2734, N2241, N2016);
buf BUF1 (N2741, N2729);
nor NOR3 (N2742, N2736, N1008, N1016);
nor NOR2 (N2743, N2695, N2047);
nand NAND3 (N2744, N2740, N474, N538);
not NOT1 (N2745, N2744);
not NOT1 (N2746, N2742);
nand NAND4 (N2747, N2746, N898, N2261, N1470);
not NOT1 (N2748, N2747);
buf BUF1 (N2749, N2738);
nor NOR2 (N2750, N2735, N1689);
and AND2 (N2751, N2739, N441);
and AND4 (N2752, N2750, N2398, N1437, N1681);
buf BUF1 (N2753, N2749);
and AND2 (N2754, N2753, N624);
and AND3 (N2755, N2743, N441, N2730);
xor XOR2 (N2756, N2755, N340);
and AND4 (N2757, N2741, N2307, N1126, N1279);
buf BUF1 (N2758, N2748);
or OR2 (N2759, N2758, N1769);
or OR3 (N2760, N2754, N2385, N599);
not NOT1 (N2761, N2760);
nand NAND3 (N2762, N2751, N1460, N577);
not NOT1 (N2763, N2761);
not NOT1 (N2764, N2745);
xor XOR2 (N2765, N2726, N730);
not NOT1 (N2766, N2737);
not NOT1 (N2767, N2766);
nor NOR2 (N2768, N2767, N1441);
and AND3 (N2769, N2724, N1997, N1395);
buf BUF1 (N2770, N2769);
and AND2 (N2771, N2763, N2322);
nor NOR4 (N2772, N2771, N1756, N2379, N2421);
nor NOR2 (N2773, N2759, N2687);
or OR4 (N2774, N2764, N910, N1150, N2687);
xor XOR2 (N2775, N2757, N2586);
nor NOR3 (N2776, N2768, N2768, N1767);
and AND3 (N2777, N2770, N1584, N1179);
xor XOR2 (N2778, N2775, N971);
and AND4 (N2779, N2776, N2000, N1350, N741);
not NOT1 (N2780, N2777);
buf BUF1 (N2781, N2762);
buf BUF1 (N2782, N2778);
nand NAND2 (N2783, N2779, N2249);
buf BUF1 (N2784, N2781);
not NOT1 (N2785, N2780);
not NOT1 (N2786, N2756);
nor NOR4 (N2787, N2782, N1347, N1408, N2600);
xor XOR2 (N2788, N2773, N5);
nand NAND3 (N2789, N2765, N635, N1207);
xor XOR2 (N2790, N2785, N2067);
nor NOR4 (N2791, N2790, N696, N2087, N1690);
nor NOR4 (N2792, N2774, N1862, N1831, N991);
buf BUF1 (N2793, N2791);
nor NOR2 (N2794, N2783, N2682);
not NOT1 (N2795, N2786);
nand NAND3 (N2796, N2788, N2498, N180);
xor XOR2 (N2797, N2795, N2592);
and AND4 (N2798, N2787, N987, N268, N804);
xor XOR2 (N2799, N2793, N2277);
not NOT1 (N2800, N2784);
and AND4 (N2801, N2800, N1740, N532, N1294);
nand NAND3 (N2802, N2752, N998, N2795);
nand NAND2 (N2803, N2801, N775);
buf BUF1 (N2804, N2798);
not NOT1 (N2805, N2792);
nand NAND4 (N2806, N2799, N2419, N699, N2233);
buf BUF1 (N2807, N2806);
xor XOR2 (N2808, N2789, N372);
not NOT1 (N2809, N2796);
not NOT1 (N2810, N2803);
xor XOR2 (N2811, N2809, N282);
nor NOR2 (N2812, N2805, N2115);
xor XOR2 (N2813, N2772, N1995);
or OR2 (N2814, N2794, N282);
nor NOR3 (N2815, N2810, N1445, N768);
xor XOR2 (N2816, N2802, N607);
or OR4 (N2817, N2807, N2441, N643, N2725);
nand NAND3 (N2818, N2812, N491, N1758);
or OR2 (N2819, N2808, N2755);
xor XOR2 (N2820, N2815, N1316);
buf BUF1 (N2821, N2819);
not NOT1 (N2822, N2804);
nand NAND2 (N2823, N2822, N870);
or OR3 (N2824, N2811, N600, N835);
buf BUF1 (N2825, N2824);
nand NAND4 (N2826, N2818, N918, N65, N2300);
buf BUF1 (N2827, N2826);
nor NOR3 (N2828, N2823, N536, N114);
nand NAND3 (N2829, N2797, N2261, N1442);
or OR2 (N2830, N2828, N828);
xor XOR2 (N2831, N2814, N296);
nand NAND2 (N2832, N2816, N62);
nor NOR4 (N2833, N2830, N790, N1464, N1498);
or OR4 (N2834, N2833, N1510, N2017, N1000);
not NOT1 (N2835, N2821);
not NOT1 (N2836, N2825);
xor XOR2 (N2837, N2831, N1357);
and AND4 (N2838, N2813, N2170, N434, N1172);
nand NAND3 (N2839, N2832, N2107, N895);
xor XOR2 (N2840, N2835, N2497);
not NOT1 (N2841, N2839);
nand NAND3 (N2842, N2817, N2454, N2233);
or OR3 (N2843, N2827, N814, N101);
not NOT1 (N2844, N2841);
and AND3 (N2845, N2842, N2392, N611);
buf BUF1 (N2846, N2843);
and AND3 (N2847, N2840, N271, N1870);
nor NOR4 (N2848, N2834, N557, N1349, N452);
or OR3 (N2849, N2845, N2216, N853);
and AND4 (N2850, N2820, N1916, N1025, N2336);
or OR3 (N2851, N2844, N2003, N2823);
nor NOR3 (N2852, N2847, N519, N1855);
buf BUF1 (N2853, N2851);
and AND3 (N2854, N2848, N2677, N237);
nor NOR4 (N2855, N2853, N1436, N337, N1183);
not NOT1 (N2856, N2854);
buf BUF1 (N2857, N2856);
or OR3 (N2858, N2855, N1496, N2141);
buf BUF1 (N2859, N2849);
or OR3 (N2860, N2857, N1980, N1533);
and AND2 (N2861, N2829, N1336);
nor NOR3 (N2862, N2860, N1793, N986);
xor XOR2 (N2863, N2862, N1044);
not NOT1 (N2864, N2858);
nand NAND2 (N2865, N2863, N1265);
buf BUF1 (N2866, N2861);
buf BUF1 (N2867, N2864);
buf BUF1 (N2868, N2859);
or OR4 (N2869, N2836, N55, N780, N1470);
or OR4 (N2870, N2868, N2269, N2230, N249);
and AND3 (N2871, N2846, N645, N572);
not NOT1 (N2872, N2866);
not NOT1 (N2873, N2871);
and AND3 (N2874, N2850, N706, N402);
buf BUF1 (N2875, N2874);
buf BUF1 (N2876, N2872);
not NOT1 (N2877, N2867);
buf BUF1 (N2878, N2852);
not NOT1 (N2879, N2875);
xor XOR2 (N2880, N2869, N370);
nor NOR2 (N2881, N2865, N1912);
not NOT1 (N2882, N2837);
nor NOR4 (N2883, N2877, N2322, N1831, N1461);
nand NAND2 (N2884, N2873, N2656);
and AND4 (N2885, N2882, N1963, N159, N1159);
xor XOR2 (N2886, N2838, N2426);
or OR3 (N2887, N2885, N1378, N1309);
nor NOR3 (N2888, N2883, N512, N1107);
xor XOR2 (N2889, N2870, N1247);
xor XOR2 (N2890, N2880, N1187);
or OR3 (N2891, N2889, N2217, N1868);
buf BUF1 (N2892, N2890);
nor NOR3 (N2893, N2876, N1051, N2770);
and AND3 (N2894, N2891, N2259, N2496);
and AND3 (N2895, N2893, N2554, N1801);
nor NOR4 (N2896, N2894, N2372, N2400, N1741);
and AND3 (N2897, N2896, N667, N1713);
or OR2 (N2898, N2892, N2422);
xor XOR2 (N2899, N2898, N289);
xor XOR2 (N2900, N2897, N2292);
buf BUF1 (N2901, N2899);
xor XOR2 (N2902, N2886, N2254);
nand NAND4 (N2903, N2884, N961, N2282, N2484);
nand NAND2 (N2904, N2888, N1420);
buf BUF1 (N2905, N2902);
nand NAND2 (N2906, N2878, N613);
and AND2 (N2907, N2903, N227);
not NOT1 (N2908, N2905);
nor NOR3 (N2909, N2895, N2042, N1861);
nand NAND4 (N2910, N2901, N2873, N982, N2117);
xor XOR2 (N2911, N2879, N1461);
and AND4 (N2912, N2906, N199, N259, N1537);
nor NOR3 (N2913, N2881, N2662, N723);
nand NAND4 (N2914, N2904, N1901, N1771, N2265);
buf BUF1 (N2915, N2909);
nand NAND2 (N2916, N2887, N2785);
and AND3 (N2917, N2916, N2449, N1472);
not NOT1 (N2918, N2900);
xor XOR2 (N2919, N2917, N2524);
buf BUF1 (N2920, N2914);
buf BUF1 (N2921, N2911);
and AND2 (N2922, N2912, N930);
not NOT1 (N2923, N2907);
nor NOR3 (N2924, N2908, N2792, N239);
nand NAND4 (N2925, N2913, N1174, N750, N823);
and AND4 (N2926, N2922, N2345, N2782, N1451);
not NOT1 (N2927, N2921);
not NOT1 (N2928, N2924);
and AND3 (N2929, N2918, N2756, N573);
nand NAND2 (N2930, N2926, N705);
nor NOR2 (N2931, N2910, N675);
buf BUF1 (N2932, N2927);
or OR4 (N2933, N2919, N2793, N1303, N1164);
xor XOR2 (N2934, N2923, N1352);
nand NAND4 (N2935, N2920, N300, N2801, N1914);
or OR4 (N2936, N2915, N1631, N1525, N850);
nand NAND2 (N2937, N2935, N1799);
buf BUF1 (N2938, N2936);
xor XOR2 (N2939, N2932, N2495);
nor NOR2 (N2940, N2931, N133);
and AND2 (N2941, N2925, N2261);
nor NOR3 (N2942, N2937, N2348, N1547);
nor NOR3 (N2943, N2941, N1003, N2708);
nand NAND4 (N2944, N2939, N1211, N2239, N1676);
buf BUF1 (N2945, N2938);
or OR3 (N2946, N2944, N2008, N2685);
or OR2 (N2947, N2942, N549);
or OR3 (N2948, N2945, N2005, N616);
or OR4 (N2949, N2940, N622, N1658, N1394);
or OR3 (N2950, N2934, N277, N803);
xor XOR2 (N2951, N2949, N627);
xor XOR2 (N2952, N2943, N653);
xor XOR2 (N2953, N2948, N873);
buf BUF1 (N2954, N2929);
buf BUF1 (N2955, N2951);
nand NAND2 (N2956, N2950, N2394);
buf BUF1 (N2957, N2954);
and AND2 (N2958, N2955, N942);
xor XOR2 (N2959, N2956, N2466);
nor NOR4 (N2960, N2953, N1526, N2135, N815);
nand NAND2 (N2961, N2947, N390);
xor XOR2 (N2962, N2952, N544);
not NOT1 (N2963, N2933);
nor NOR2 (N2964, N2946, N113);
not NOT1 (N2965, N2962);
not NOT1 (N2966, N2961);
nor NOR4 (N2967, N2963, N197, N1175, N1806);
nand NAND3 (N2968, N2957, N248, N1389);
and AND4 (N2969, N2958, N1411, N487, N1958);
and AND3 (N2970, N2969, N542, N1639);
or OR4 (N2971, N2964, N877, N1241, N1821);
or OR4 (N2972, N2971, N123, N2669, N2176);
and AND4 (N2973, N2967, N723, N204, N1939);
xor XOR2 (N2974, N2968, N765);
nor NOR4 (N2975, N2959, N2954, N1398, N2021);
nor NOR3 (N2976, N2972, N1711, N2698);
or OR4 (N2977, N2973, N1776, N383, N1747);
and AND4 (N2978, N2960, N1603, N1187, N1378);
not NOT1 (N2979, N2928);
or OR4 (N2980, N2970, N328, N2120, N2167);
nand NAND3 (N2981, N2965, N632, N372);
xor XOR2 (N2982, N2977, N2520);
xor XOR2 (N2983, N2980, N511);
and AND4 (N2984, N2981, N904, N1842, N2467);
not NOT1 (N2985, N2983);
and AND4 (N2986, N2982, N1705, N690, N1026);
nor NOR2 (N2987, N2986, N2113);
not NOT1 (N2988, N2987);
and AND3 (N2989, N2930, N334, N1083);
nand NAND4 (N2990, N2976, N1961, N1598, N1880);
nand NAND3 (N2991, N2989, N2209, N2490);
or OR2 (N2992, N2988, N1573);
buf BUF1 (N2993, N2984);
or OR3 (N2994, N2990, N2794, N2719);
nand NAND3 (N2995, N2979, N458, N2584);
nand NAND4 (N2996, N2994, N592, N2573, N2373);
not NOT1 (N2997, N2995);
or OR4 (N2998, N2975, N1764, N1066, N1820);
nand NAND3 (N2999, N2992, N1714, N2527);
nor NOR4 (N3000, N2997, N1594, N1724, N1075);
buf BUF1 (N3001, N2974);
and AND4 (N3002, N2966, N2489, N2599, N2487);
xor XOR2 (N3003, N3000, N1461);
xor XOR2 (N3004, N2985, N604);
nand NAND4 (N3005, N2996, N1652, N1296, N2364);
not NOT1 (N3006, N3001);
nand NAND2 (N3007, N3006, N1916);
xor XOR2 (N3008, N3005, N833);
nor NOR4 (N3009, N3008, N527, N1647, N2752);
and AND4 (N3010, N2993, N1739, N1029, N654);
xor XOR2 (N3011, N2991, N218);
xor XOR2 (N3012, N2998, N1119);
not NOT1 (N3013, N3007);
and AND3 (N3014, N3010, N2761, N54);
xor XOR2 (N3015, N3002, N2313);
or OR4 (N3016, N3011, N1008, N1741, N1946);
or OR3 (N3017, N3014, N1846, N484);
and AND2 (N3018, N3004, N2803);
not NOT1 (N3019, N2999);
nor NOR3 (N3020, N3012, N304, N1265);
not NOT1 (N3021, N3009);
nand NAND2 (N3022, N3020, N198);
nor NOR2 (N3023, N3003, N2788);
buf BUF1 (N3024, N3015);
and AND4 (N3025, N3023, N120, N1611, N254);
nand NAND4 (N3026, N3024, N332, N3023, N2764);
not NOT1 (N3027, N3016);
nor NOR2 (N3028, N3021, N2141);
or OR2 (N3029, N2978, N2109);
nor NOR4 (N3030, N3017, N1296, N2775, N2371);
not NOT1 (N3031, N3022);
or OR4 (N3032, N3029, N39, N2531, N1563);
nand NAND4 (N3033, N3028, N2836, N2562, N2431);
and AND2 (N3034, N3025, N2706);
nand NAND3 (N3035, N3013, N1197, N1298);
nand NAND3 (N3036, N3031, N361, N501);
buf BUF1 (N3037, N3035);
nor NOR2 (N3038, N3034, N1118);
nand NAND4 (N3039, N3033, N2349, N379, N2955);
buf BUF1 (N3040, N3030);
nand NAND3 (N3041, N3040, N2938, N394);
not NOT1 (N3042, N3019);
and AND3 (N3043, N3041, N2140, N694);
and AND2 (N3044, N3018, N98);
nand NAND3 (N3045, N3036, N618, N3008);
buf BUF1 (N3046, N3042);
nor NOR3 (N3047, N3045, N300, N1015);
nand NAND2 (N3048, N3046, N622);
not NOT1 (N3049, N3027);
or OR3 (N3050, N3049, N630, N3006);
nor NOR3 (N3051, N3039, N1325, N617);
not NOT1 (N3052, N3043);
or OR2 (N3053, N3038, N2020);
not NOT1 (N3054, N3026);
or OR3 (N3055, N3047, N2805, N83);
nand NAND4 (N3056, N3053, N1641, N2224, N625);
not NOT1 (N3057, N3044);
buf BUF1 (N3058, N3037);
buf BUF1 (N3059, N3050);
buf BUF1 (N3060, N3054);
buf BUF1 (N3061, N3057);
and AND4 (N3062, N3059, N426, N748, N1090);
nor NOR3 (N3063, N3055, N692, N2095);
not NOT1 (N3064, N3051);
and AND4 (N3065, N3058, N2097, N1028, N22);
nand NAND2 (N3066, N3048, N2713);
and AND3 (N3067, N3062, N2373, N555);
not NOT1 (N3068, N3065);
and AND2 (N3069, N3066, N2817);
and AND2 (N3070, N3067, N37);
xor XOR2 (N3071, N3068, N909);
buf BUF1 (N3072, N3064);
xor XOR2 (N3073, N3072, N1365);
buf BUF1 (N3074, N3070);
nor NOR4 (N3075, N3074, N1113, N413, N508);
not NOT1 (N3076, N3063);
not NOT1 (N3077, N3075);
buf BUF1 (N3078, N3032);
nand NAND3 (N3079, N3073, N1786, N2249);
nor NOR3 (N3080, N3077, N3073, N1914);
buf BUF1 (N3081, N3071);
and AND4 (N3082, N3076, N2598, N1612, N2081);
or OR2 (N3083, N3060, N1527);
and AND2 (N3084, N3061, N1863);
xor XOR2 (N3085, N3082, N1322);
or OR4 (N3086, N3085, N1427, N1524, N2618);
xor XOR2 (N3087, N3083, N2786);
nor NOR2 (N3088, N3052, N800);
buf BUF1 (N3089, N3088);
and AND4 (N3090, N3069, N1148, N152, N1453);
nor NOR4 (N3091, N3080, N3034, N602, N1956);
xor XOR2 (N3092, N3081, N1885);
not NOT1 (N3093, N3079);
or OR4 (N3094, N3078, N529, N1648, N2759);
nand NAND2 (N3095, N3094, N3080);
not NOT1 (N3096, N3086);
nor NOR2 (N3097, N3093, N2551);
xor XOR2 (N3098, N3087, N1283);
and AND2 (N3099, N3097, N2721);
nor NOR4 (N3100, N3098, N1839, N2792, N766);
and AND3 (N3101, N3091, N2725, N1063);
or OR2 (N3102, N3056, N1587);
or OR4 (N3103, N3092, N2104, N552, N2747);
nor NOR2 (N3104, N3096, N180);
xor XOR2 (N3105, N3084, N2880);
nor NOR2 (N3106, N3089, N745);
xor XOR2 (N3107, N3104, N290);
buf BUF1 (N3108, N3095);
buf BUF1 (N3109, N3105);
xor XOR2 (N3110, N3107, N2416);
or OR4 (N3111, N3108, N609, N2737, N428);
and AND3 (N3112, N3090, N1471, N219);
buf BUF1 (N3113, N3102);
nand NAND4 (N3114, N3110, N342, N1444, N2982);
not NOT1 (N3115, N3114);
and AND3 (N3116, N3103, N667, N1983);
buf BUF1 (N3117, N3112);
buf BUF1 (N3118, N3111);
xor XOR2 (N3119, N3101, N2329);
nor NOR4 (N3120, N3119, N1894, N1367, N20);
buf BUF1 (N3121, N3109);
buf BUF1 (N3122, N3099);
buf BUF1 (N3123, N3100);
not NOT1 (N3124, N3120);
nor NOR4 (N3125, N3115, N992, N1562, N1816);
and AND2 (N3126, N3125, N912);
and AND3 (N3127, N3106, N2928, N1697);
or OR2 (N3128, N3118, N59);
nand NAND3 (N3129, N3127, N2327, N2003);
or OR3 (N3130, N3117, N2817, N935);
or OR2 (N3131, N3116, N2186);
xor XOR2 (N3132, N3128, N1146);
nand NAND4 (N3133, N3113, N1698, N2058, N867);
or OR2 (N3134, N3129, N3044);
xor XOR2 (N3135, N3134, N934);
or OR4 (N3136, N3122, N1955, N1853, N2363);
and AND3 (N3137, N3126, N2080, N2317);
or OR2 (N3138, N3132, N2703);
nor NOR3 (N3139, N3135, N353, N2304);
not NOT1 (N3140, N3130);
xor XOR2 (N3141, N3136, N2748);
and AND3 (N3142, N3140, N2636, N601);
or OR3 (N3143, N3139, N693, N377);
and AND2 (N3144, N3143, N337);
xor XOR2 (N3145, N3133, N2573);
nand NAND2 (N3146, N3123, N766);
or OR4 (N3147, N3144, N577, N1568, N2093);
xor XOR2 (N3148, N3131, N641);
buf BUF1 (N3149, N3145);
nor NOR2 (N3150, N3138, N1690);
buf BUF1 (N3151, N3148);
buf BUF1 (N3152, N3121);
or OR2 (N3153, N3141, N160);
and AND4 (N3154, N3147, N851, N2281, N2089);
and AND4 (N3155, N3152, N3140, N1591, N1);
not NOT1 (N3156, N3142);
not NOT1 (N3157, N3124);
buf BUF1 (N3158, N3137);
nor NOR2 (N3159, N3150, N533);
or OR2 (N3160, N3149, N2139);
nand NAND4 (N3161, N3151, N638, N2795, N501);
buf BUF1 (N3162, N3154);
and AND4 (N3163, N3157, N992, N2836, N1191);
or OR4 (N3164, N3155, N1654, N2791, N2670);
buf BUF1 (N3165, N3161);
buf BUF1 (N3166, N3163);
nand NAND3 (N3167, N3165, N2011, N1249);
buf BUF1 (N3168, N3166);
and AND2 (N3169, N3167, N1340);
and AND4 (N3170, N3146, N737, N853, N223);
and AND4 (N3171, N3153, N2331, N323, N1039);
nor NOR2 (N3172, N3168, N2160);
nand NAND2 (N3173, N3162, N2896);
not NOT1 (N3174, N3158);
or OR3 (N3175, N3156, N1667, N2202);
nand NAND4 (N3176, N3170, N3160, N2484, N1570);
and AND2 (N3177, N1959, N104);
buf BUF1 (N3178, N3164);
nor NOR4 (N3179, N3177, N2107, N1641, N300);
xor XOR2 (N3180, N3169, N408);
and AND2 (N3181, N3176, N107);
and AND3 (N3182, N3181, N141, N963);
not NOT1 (N3183, N3178);
not NOT1 (N3184, N3171);
not NOT1 (N3185, N3183);
nand NAND4 (N3186, N3185, N1364, N808, N353);
not NOT1 (N3187, N3179);
or OR4 (N3188, N3159, N803, N1262, N2878);
and AND3 (N3189, N3172, N1044, N461);
not NOT1 (N3190, N3173);
xor XOR2 (N3191, N3190, N2520);
nand NAND4 (N3192, N3184, N636, N2984, N1109);
nand NAND2 (N3193, N3182, N510);
xor XOR2 (N3194, N3189, N1082);
not NOT1 (N3195, N3188);
buf BUF1 (N3196, N3192);
or OR4 (N3197, N3195, N2466, N1338, N247);
or OR2 (N3198, N3196, N3170);
buf BUF1 (N3199, N3180);
nand NAND2 (N3200, N3174, N2076);
not NOT1 (N3201, N3187);
nor NOR2 (N3202, N3201, N2024);
and AND3 (N3203, N3175, N791, N630);
or OR3 (N3204, N3198, N1545, N2646);
buf BUF1 (N3205, N3191);
nand NAND3 (N3206, N3199, N1158, N2775);
not NOT1 (N3207, N3203);
and AND4 (N3208, N3186, N496, N73, N2205);
buf BUF1 (N3209, N3193);
not NOT1 (N3210, N3194);
nand NAND4 (N3211, N3200, N925, N2973, N1769);
nor NOR4 (N3212, N3202, N1914, N527, N1355);
nand NAND3 (N3213, N3206, N1635, N236);
buf BUF1 (N3214, N3205);
nand NAND3 (N3215, N3204, N723, N2052);
nor NOR4 (N3216, N3213, N1352, N1712, N176);
xor XOR2 (N3217, N3212, N2141);
xor XOR2 (N3218, N3215, N2046);
nand NAND4 (N3219, N3216, N1173, N2619, N1537);
buf BUF1 (N3220, N3209);
nor NOR3 (N3221, N3220, N3183, N1777);
nand NAND2 (N3222, N3217, N1840);
buf BUF1 (N3223, N3221);
and AND4 (N3224, N3223, N3190, N1019, N1744);
nor NOR4 (N3225, N3219, N3222, N2459, N2832);
nor NOR3 (N3226, N705, N2432, N2749);
nor NOR4 (N3227, N3224, N2811, N1128, N2729);
buf BUF1 (N3228, N3227);
or OR3 (N3229, N3210, N586, N136);
or OR3 (N3230, N3228, N499, N2963);
not NOT1 (N3231, N3229);
nor NOR4 (N3232, N3231, N1211, N1784, N1885);
or OR3 (N3233, N3232, N3070, N2472);
nand NAND4 (N3234, N3218, N1209, N1934, N308);
not NOT1 (N3235, N3225);
nand NAND4 (N3236, N3211, N1583, N1719, N2514);
or OR2 (N3237, N3235, N455);
and AND3 (N3238, N3208, N414, N2263);
buf BUF1 (N3239, N3238);
nor NOR2 (N3240, N3230, N2614);
buf BUF1 (N3241, N3207);
not NOT1 (N3242, N3214);
not NOT1 (N3243, N3241);
buf BUF1 (N3244, N3236);
buf BUF1 (N3245, N3240);
buf BUF1 (N3246, N3226);
not NOT1 (N3247, N3239);
nand NAND3 (N3248, N3233, N2091, N3091);
nand NAND2 (N3249, N3234, N2473);
not NOT1 (N3250, N3244);
nor NOR4 (N3251, N3237, N836, N2290, N2948);
nand NAND3 (N3252, N3242, N3147, N711);
not NOT1 (N3253, N3248);
not NOT1 (N3254, N3246);
nor NOR2 (N3255, N3251, N1207);
not NOT1 (N3256, N3253);
not NOT1 (N3257, N3252);
or OR2 (N3258, N3254, N2992);
xor XOR2 (N3259, N3256, N308);
nor NOR4 (N3260, N3243, N2997, N2902, N1724);
or OR4 (N3261, N3260, N1122, N1610, N1300);
and AND4 (N3262, N3259, N1144, N911, N661);
and AND3 (N3263, N3255, N2159, N3192);
not NOT1 (N3264, N3245);
nand NAND4 (N3265, N3250, N3226, N563, N1257);
or OR4 (N3266, N3264, N2741, N233, N559);
not NOT1 (N3267, N3262);
not NOT1 (N3268, N3258);
nand NAND2 (N3269, N3261, N455);
xor XOR2 (N3270, N3266, N506);
xor XOR2 (N3271, N3270, N1488);
nand NAND4 (N3272, N3197, N2241, N3051, N883);
nor NOR2 (N3273, N3247, N119);
and AND3 (N3274, N3272, N2687, N1355);
xor XOR2 (N3275, N3274, N2643);
not NOT1 (N3276, N3275);
xor XOR2 (N3277, N3249, N1564);
or OR2 (N3278, N3257, N3122);
or OR3 (N3279, N3278, N1366, N447);
nor NOR4 (N3280, N3277, N1746, N5, N2829);
not NOT1 (N3281, N3279);
xor XOR2 (N3282, N3281, N2724);
xor XOR2 (N3283, N3269, N987);
and AND4 (N3284, N3283, N1500, N1702, N2543);
and AND4 (N3285, N3273, N2467, N322, N968);
nor NOR3 (N3286, N3282, N911, N1291);
and AND4 (N3287, N3284, N2033, N2478, N2868);
nor NOR4 (N3288, N3268, N283, N3093, N2376);
buf BUF1 (N3289, N3280);
and AND2 (N3290, N3286, N1954);
nand NAND4 (N3291, N3288, N1026, N33, N980);
nand NAND3 (N3292, N3267, N769, N2077);
and AND2 (N3293, N3290, N2042);
nor NOR4 (N3294, N3265, N1584, N1944, N1950);
nor NOR3 (N3295, N3287, N1078, N1795);
nand NAND4 (N3296, N3292, N626, N756, N3095);
or OR2 (N3297, N3276, N1232);
xor XOR2 (N3298, N3285, N2504);
nor NOR3 (N3299, N3271, N2532, N1402);
xor XOR2 (N3300, N3289, N1369);
xor XOR2 (N3301, N3293, N1255);
nand NAND4 (N3302, N3299, N1134, N2814, N2200);
not NOT1 (N3303, N3302);
or OR3 (N3304, N3301, N1858, N52);
xor XOR2 (N3305, N3263, N821);
or OR3 (N3306, N3296, N1447, N361);
buf BUF1 (N3307, N3305);
and AND3 (N3308, N3295, N3248, N534);
and AND2 (N3309, N3291, N598);
buf BUF1 (N3310, N3308);
nand NAND2 (N3311, N3297, N215);
nor NOR3 (N3312, N3306, N139, N1004);
not NOT1 (N3313, N3307);
not NOT1 (N3314, N3294);
or OR3 (N3315, N3304, N1191, N1431);
nand NAND2 (N3316, N3300, N2887);
nand NAND2 (N3317, N3303, N844);
nand NAND3 (N3318, N3309, N301, N2900);
or OR4 (N3319, N3310, N2962, N1571, N2512);
and AND4 (N3320, N3313, N2938, N104, N2960);
or OR3 (N3321, N3312, N927, N2041);
buf BUF1 (N3322, N3314);
and AND3 (N3323, N3320, N2054, N2954);
nand NAND2 (N3324, N3319, N2155);
nand NAND2 (N3325, N3324, N977);
nor NOR2 (N3326, N3323, N736);
and AND2 (N3327, N3316, N2345);
nor NOR4 (N3328, N3321, N2612, N360, N2534);
and AND4 (N3329, N3327, N670, N473, N2500);
not NOT1 (N3330, N3317);
xor XOR2 (N3331, N3325, N2202);
nor NOR2 (N3332, N3322, N765);
nor NOR4 (N3333, N3318, N2483, N554, N2432);
nand NAND2 (N3334, N3333, N1198);
nor NOR2 (N3335, N3328, N2148);
and AND3 (N3336, N3315, N2750, N2287);
or OR3 (N3337, N3311, N2818, N818);
nand NAND3 (N3338, N3330, N3337, N812);
not NOT1 (N3339, N1559);
nor NOR4 (N3340, N3338, N3329, N2139, N36);
buf BUF1 (N3341, N2264);
nand NAND2 (N3342, N3331, N899);
and AND3 (N3343, N3298, N2379, N1052);
or OR3 (N3344, N3339, N1305, N264);
and AND4 (N3345, N3343, N1601, N2244, N1207);
buf BUF1 (N3346, N3342);
xor XOR2 (N3347, N3341, N2123);
nor NOR4 (N3348, N3340, N2348, N2166, N2460);
and AND2 (N3349, N3335, N2223);
nor NOR2 (N3350, N3349, N1148);
xor XOR2 (N3351, N3348, N794);
nor NOR2 (N3352, N3326, N1894);
buf BUF1 (N3353, N3346);
or OR3 (N3354, N3332, N314, N51);
xor XOR2 (N3355, N3350, N2548);
and AND2 (N3356, N3354, N30);
nor NOR2 (N3357, N3356, N1537);
xor XOR2 (N3358, N3355, N1946);
or OR3 (N3359, N3353, N1803, N2045);
or OR4 (N3360, N3351, N1980, N2284, N2067);
not NOT1 (N3361, N3357);
buf BUF1 (N3362, N3360);
and AND4 (N3363, N3344, N120, N728, N2863);
nor NOR2 (N3364, N3352, N258);
not NOT1 (N3365, N3363);
nor NOR4 (N3366, N3358, N267, N3133, N3319);
buf BUF1 (N3367, N3366);
buf BUF1 (N3368, N3336);
buf BUF1 (N3369, N3362);
not NOT1 (N3370, N3334);
xor XOR2 (N3371, N3361, N1110);
or OR2 (N3372, N3365, N1718);
or OR4 (N3373, N3359, N47, N2417, N2512);
nor NOR4 (N3374, N3370, N1511, N2755, N584);
not NOT1 (N3375, N3369);
nor NOR3 (N3376, N3373, N2051, N2530);
or OR2 (N3377, N3375, N739);
nor NOR2 (N3378, N3364, N247);
xor XOR2 (N3379, N3376, N60);
buf BUF1 (N3380, N3368);
xor XOR2 (N3381, N3374, N1693);
and AND4 (N3382, N3381, N2028, N2935, N2058);
and AND3 (N3383, N3347, N2252, N2060);
buf BUF1 (N3384, N3345);
nand NAND2 (N3385, N3384, N2569);
xor XOR2 (N3386, N3378, N1592);
and AND3 (N3387, N3372, N1766, N1438);
or OR2 (N3388, N3371, N2831);
not NOT1 (N3389, N3367);
or OR2 (N3390, N3388, N386);
buf BUF1 (N3391, N3380);
or OR2 (N3392, N3383, N838);
or OR2 (N3393, N3392, N400);
buf BUF1 (N3394, N3377);
nor NOR4 (N3395, N3391, N2139, N2822, N1674);
xor XOR2 (N3396, N3394, N1601);
or OR4 (N3397, N3385, N1316, N299, N644);
not NOT1 (N3398, N3395);
not NOT1 (N3399, N3398);
or OR4 (N3400, N3399, N2313, N685, N3047);
and AND4 (N3401, N3386, N654, N2919, N3316);
buf BUF1 (N3402, N3389);
buf BUF1 (N3403, N3382);
nor NOR3 (N3404, N3379, N3187, N2861);
and AND2 (N3405, N3396, N2065);
xor XOR2 (N3406, N3401, N3056);
buf BUF1 (N3407, N3404);
nor NOR3 (N3408, N3406, N1305, N1047);
nand NAND3 (N3409, N3403, N1783, N1759);
or OR4 (N3410, N3409, N3362, N1490, N3001);
or OR4 (N3411, N3407, N709, N2055, N1347);
and AND3 (N3412, N3393, N2676, N259);
nand NAND3 (N3413, N3390, N730, N1418);
nand NAND4 (N3414, N3408, N103, N1543, N2712);
or OR4 (N3415, N3410, N444, N868, N790);
not NOT1 (N3416, N3412);
nor NOR3 (N3417, N3415, N1382, N2549);
nand NAND2 (N3418, N3411, N107);
buf BUF1 (N3419, N3405);
and AND2 (N3420, N3397, N1681);
nor NOR3 (N3421, N3420, N3413, N396);
buf BUF1 (N3422, N3049);
and AND4 (N3423, N3418, N2605, N222, N2667);
nand NAND3 (N3424, N3422, N566, N163);
xor XOR2 (N3425, N3419, N911);
and AND4 (N3426, N3421, N1756, N2834, N2004);
nor NOR2 (N3427, N3414, N841);
nand NAND3 (N3428, N3427, N1679, N2742);
nand NAND4 (N3429, N3387, N3033, N473, N3260);
and AND2 (N3430, N3428, N332);
buf BUF1 (N3431, N3400);
nand NAND4 (N3432, N3424, N402, N1940, N2915);
nand NAND2 (N3433, N3426, N1178);
nand NAND2 (N3434, N3432, N251);
or OR3 (N3435, N3433, N2723, N2149);
buf BUF1 (N3436, N3429);
nand NAND4 (N3437, N3423, N2744, N1617, N3230);
buf BUF1 (N3438, N3437);
not NOT1 (N3439, N3402);
xor XOR2 (N3440, N3438, N10);
nand NAND2 (N3441, N3435, N1127);
nand NAND3 (N3442, N3434, N2215, N1391);
buf BUF1 (N3443, N3431);
and AND3 (N3444, N3443, N160, N1019);
buf BUF1 (N3445, N3430);
not NOT1 (N3446, N3445);
and AND3 (N3447, N3436, N875, N1132);
nand NAND4 (N3448, N3417, N1868, N2503, N1645);
buf BUF1 (N3449, N3416);
buf BUF1 (N3450, N3446);
and AND3 (N3451, N3447, N3094, N935);
buf BUF1 (N3452, N3449);
not NOT1 (N3453, N3440);
and AND3 (N3454, N3444, N3327, N1362);
nor NOR4 (N3455, N3450, N2199, N2601, N1591);
nor NOR3 (N3456, N3454, N1463, N2078);
nand NAND3 (N3457, N3441, N2824, N1490);
or OR4 (N3458, N3455, N73, N753, N2727);
nor NOR3 (N3459, N3456, N1765, N1850);
or OR3 (N3460, N3459, N3364, N3117);
or OR2 (N3461, N3457, N1645);
nor NOR2 (N3462, N3461, N362);
or OR3 (N3463, N3453, N920, N1974);
and AND2 (N3464, N3439, N2175);
or OR4 (N3465, N3463, N3005, N1837, N3025);
not NOT1 (N3466, N3465);
and AND4 (N3467, N3458, N2445, N1843, N1322);
and AND2 (N3468, N3452, N268);
and AND2 (N3469, N3468, N1224);
nor NOR2 (N3470, N3462, N2664);
not NOT1 (N3471, N3442);
not NOT1 (N3472, N3469);
xor XOR2 (N3473, N3451, N2080);
nand NAND2 (N3474, N3471, N2080);
and AND3 (N3475, N3472, N354, N2501);
nand NAND4 (N3476, N3466, N1153, N1697, N73);
not NOT1 (N3477, N3475);
nand NAND3 (N3478, N3464, N3089, N502);
nand NAND4 (N3479, N3467, N394, N1197, N1979);
buf BUF1 (N3480, N3478);
or OR4 (N3481, N3479, N3154, N1570, N1568);
xor XOR2 (N3482, N3480, N1146);
and AND3 (N3483, N3482, N2746, N751);
nor NOR4 (N3484, N3483, N2458, N959, N519);
or OR4 (N3485, N3425, N1050, N2996, N216);
and AND2 (N3486, N3476, N670);
or OR2 (N3487, N3460, N3329);
not NOT1 (N3488, N3487);
and AND2 (N3489, N3486, N2201);
and AND4 (N3490, N3477, N935, N318, N105);
and AND3 (N3491, N3474, N3004, N2587);
xor XOR2 (N3492, N3448, N738);
and AND3 (N3493, N3489, N1104, N2508);
not NOT1 (N3494, N3488);
or OR2 (N3495, N3485, N1125);
buf BUF1 (N3496, N3494);
not NOT1 (N3497, N3493);
or OR3 (N3498, N3492, N2519, N1646);
nand NAND2 (N3499, N3491, N2339);
buf BUF1 (N3500, N3470);
xor XOR2 (N3501, N3495, N274);
xor XOR2 (N3502, N3499, N604);
xor XOR2 (N3503, N3490, N2529);
buf BUF1 (N3504, N3498);
and AND2 (N3505, N3503, N2502);
or OR3 (N3506, N3473, N3168, N1798);
buf BUF1 (N3507, N3506);
xor XOR2 (N3508, N3505, N1571);
and AND3 (N3509, N3496, N3187, N1612);
and AND4 (N3510, N3501, N1957, N2318, N1616);
buf BUF1 (N3511, N3510);
nor NOR2 (N3512, N3504, N3326);
or OR2 (N3513, N3511, N3003);
or OR2 (N3514, N3481, N2615);
not NOT1 (N3515, N3507);
xor XOR2 (N3516, N3515, N1033);
or OR2 (N3517, N3512, N2405);
or OR3 (N3518, N3514, N2494, N72);
buf BUF1 (N3519, N3500);
nor NOR3 (N3520, N3509, N796, N72);
and AND2 (N3521, N3518, N921);
nand NAND3 (N3522, N3497, N2611, N3370);
nor NOR4 (N3523, N3519, N479, N1473, N1425);
not NOT1 (N3524, N3523);
xor XOR2 (N3525, N3517, N3288);
xor XOR2 (N3526, N3513, N3051);
nand NAND4 (N3527, N3520, N347, N308, N2144);
buf BUF1 (N3528, N3526);
nand NAND3 (N3529, N3525, N417, N3055);
nor NOR3 (N3530, N3527, N1666, N2398);
xor XOR2 (N3531, N3508, N2145);
and AND3 (N3532, N3516, N1923, N651);
not NOT1 (N3533, N3524);
or OR3 (N3534, N3502, N562, N1423);
nand NAND3 (N3535, N3528, N797, N721);
xor XOR2 (N3536, N3522, N802);
nand NAND3 (N3537, N3531, N1038, N1731);
xor XOR2 (N3538, N3537, N3508);
or OR3 (N3539, N3534, N313, N1152);
buf BUF1 (N3540, N3533);
nor NOR3 (N3541, N3484, N2022, N1506);
or OR2 (N3542, N3532, N3227);
or OR4 (N3543, N3542, N2254, N2895, N2083);
nand NAND2 (N3544, N3543, N2678);
or OR2 (N3545, N3540, N37);
nor NOR4 (N3546, N3530, N1599, N597, N2756);
xor XOR2 (N3547, N3529, N1790);
buf BUF1 (N3548, N3541);
nand NAND4 (N3549, N3538, N2681, N2289, N87);
or OR3 (N3550, N3539, N3267, N1967);
nor NOR4 (N3551, N3547, N1543, N105, N1916);
not NOT1 (N3552, N3548);
xor XOR2 (N3553, N3536, N66);
or OR2 (N3554, N3549, N2633);
xor XOR2 (N3555, N3553, N3253);
nor NOR3 (N3556, N3550, N2556, N2650);
and AND2 (N3557, N3544, N1826);
or OR3 (N3558, N3545, N2052, N2387);
nor NOR4 (N3559, N3535, N1731, N3339, N1054);
xor XOR2 (N3560, N3552, N572);
not NOT1 (N3561, N3554);
nor NOR2 (N3562, N3557, N1886);
nor NOR2 (N3563, N3562, N2297);
xor XOR2 (N3564, N3561, N3328);
xor XOR2 (N3565, N3551, N808);
nand NAND3 (N3566, N3563, N2778, N2709);
nor NOR3 (N3567, N3555, N2594, N254);
nor NOR4 (N3568, N3566, N290, N2271, N2393);
and AND4 (N3569, N3556, N348, N280, N2871);
nand NAND3 (N3570, N3559, N3019, N163);
not NOT1 (N3571, N3521);
and AND3 (N3572, N3571, N1897, N795);
and AND4 (N3573, N3564, N118, N2873, N369);
buf BUF1 (N3574, N3565);
and AND2 (N3575, N3570, N1368);
or OR2 (N3576, N3560, N1122);
xor XOR2 (N3577, N3572, N2424);
not NOT1 (N3578, N3569);
and AND4 (N3579, N3577, N40, N2290, N285);
or OR2 (N3580, N3579, N757);
and AND2 (N3581, N3558, N3186);
nand NAND3 (N3582, N3578, N2734, N854);
buf BUF1 (N3583, N3575);
or OR4 (N3584, N3576, N389, N2600, N2989);
xor XOR2 (N3585, N3580, N2450);
nor NOR3 (N3586, N3567, N1100, N2239);
nor NOR2 (N3587, N3568, N3139);
xor XOR2 (N3588, N3573, N3161);
and AND2 (N3589, N3574, N343);
not NOT1 (N3590, N3586);
nor NOR2 (N3591, N3585, N559);
nor NOR2 (N3592, N3591, N1350);
nand NAND3 (N3593, N3587, N3248, N2858);
buf BUF1 (N3594, N3593);
nand NAND2 (N3595, N3594, N1857);
not NOT1 (N3596, N3589);
not NOT1 (N3597, N3582);
buf BUF1 (N3598, N3592);
nor NOR4 (N3599, N3588, N1691, N2202, N574);
or OR4 (N3600, N3546, N1605, N1822, N91);
not NOT1 (N3601, N3599);
nor NOR2 (N3602, N3598, N2342);
nor NOR2 (N3603, N3590, N885);
nand NAND4 (N3604, N3583, N2352, N34, N1232);
not NOT1 (N3605, N3604);
or OR2 (N3606, N3605, N683);
and AND4 (N3607, N3597, N2788, N3419, N2203);
not NOT1 (N3608, N3584);
and AND3 (N3609, N3595, N319, N2831);
or OR4 (N3610, N3607, N604, N204, N1698);
xor XOR2 (N3611, N3600, N848);
xor XOR2 (N3612, N3581, N225);
and AND4 (N3613, N3611, N2836, N2169, N2297);
xor XOR2 (N3614, N3602, N1551);
xor XOR2 (N3615, N3613, N1148);
nand NAND4 (N3616, N3615, N1882, N3533, N1124);
xor XOR2 (N3617, N3610, N485);
buf BUF1 (N3618, N3614);
or OR3 (N3619, N3608, N3419, N2910);
and AND3 (N3620, N3601, N2633, N2579);
buf BUF1 (N3621, N3609);
xor XOR2 (N3622, N3621, N1887);
nand NAND2 (N3623, N3617, N36);
nor NOR2 (N3624, N3618, N1483);
not NOT1 (N3625, N3624);
nor NOR3 (N3626, N3619, N229, N630);
nor NOR3 (N3627, N3612, N2090, N135);
nand NAND2 (N3628, N3622, N3373);
not NOT1 (N3629, N3620);
nor NOR2 (N3630, N3626, N2810);
not NOT1 (N3631, N3629);
not NOT1 (N3632, N3596);
not NOT1 (N3633, N3627);
or OR3 (N3634, N3633, N159, N1109);
xor XOR2 (N3635, N3606, N3457);
or OR4 (N3636, N3623, N852, N509, N2963);
xor XOR2 (N3637, N3603, N1785);
and AND2 (N3638, N3632, N2268);
and AND4 (N3639, N3637, N298, N188, N3463);
nor NOR4 (N3640, N3628, N181, N3023, N2315);
nand NAND2 (N3641, N3636, N1287);
or OR2 (N3642, N3640, N1621);
nor NOR4 (N3643, N3641, N3620, N587, N1427);
buf BUF1 (N3644, N3634);
or OR2 (N3645, N3638, N2592);
nand NAND3 (N3646, N3643, N3295, N297);
and AND2 (N3647, N3639, N2628);
buf BUF1 (N3648, N3642);
nor NOR3 (N3649, N3630, N2233, N274);
buf BUF1 (N3650, N3644);
or OR4 (N3651, N3625, N1543, N2841, N215);
or OR4 (N3652, N3648, N1425, N841, N1983);
and AND2 (N3653, N3652, N1308);
buf BUF1 (N3654, N3649);
and AND2 (N3655, N3616, N3164);
and AND4 (N3656, N3635, N1495, N2021, N1905);
nand NAND2 (N3657, N3651, N2089);
not NOT1 (N3658, N3657);
not NOT1 (N3659, N3656);
and AND4 (N3660, N3659, N1672, N2121, N2535);
not NOT1 (N3661, N3631);
xor XOR2 (N3662, N3650, N3285);
not NOT1 (N3663, N3660);
not NOT1 (N3664, N3647);
nand NAND2 (N3665, N3663, N2056);
xor XOR2 (N3666, N3653, N403);
nor NOR3 (N3667, N3665, N353, N3540);
nor NOR3 (N3668, N3645, N3487, N2509);
xor XOR2 (N3669, N3654, N2512);
nor NOR3 (N3670, N3662, N369, N1095);
or OR4 (N3671, N3666, N1823, N2887, N1880);
buf BUF1 (N3672, N3661);
not NOT1 (N3673, N3669);
not NOT1 (N3674, N3670);
buf BUF1 (N3675, N3664);
or OR3 (N3676, N3658, N1797, N1004);
nand NAND2 (N3677, N3675, N1617);
buf BUF1 (N3678, N3646);
xor XOR2 (N3679, N3668, N327);
and AND4 (N3680, N3671, N3245, N3471, N127);
nand NAND2 (N3681, N3678, N396);
not NOT1 (N3682, N3679);
or OR4 (N3683, N3673, N2665, N685, N1141);
not NOT1 (N3684, N3682);
and AND4 (N3685, N3667, N1070, N1748, N1219);
buf BUF1 (N3686, N3684);
nor NOR4 (N3687, N3677, N79, N2812, N2411);
nor NOR2 (N3688, N3674, N1886);
buf BUF1 (N3689, N3686);
and AND4 (N3690, N3676, N89, N656, N2962);
or OR3 (N3691, N3690, N502, N534);
not NOT1 (N3692, N3683);
xor XOR2 (N3693, N3681, N2765);
nand NAND3 (N3694, N3655, N824, N2313);
and AND4 (N3695, N3680, N812, N696, N884);
or OR3 (N3696, N3695, N2578, N1000);
nor NOR2 (N3697, N3688, N1984);
nand NAND3 (N3698, N3691, N3219, N197);
or OR2 (N3699, N3685, N3681);
or OR4 (N3700, N3698, N3676, N2194, N2555);
buf BUF1 (N3701, N3692);
buf BUF1 (N3702, N3672);
or OR2 (N3703, N3697, N2704);
buf BUF1 (N3704, N3699);
buf BUF1 (N3705, N3696);
or OR4 (N3706, N3702, N2223, N1661, N1653);
not NOT1 (N3707, N3689);
nand NAND4 (N3708, N3703, N3184, N391, N3705);
xor XOR2 (N3709, N1679, N2690);
buf BUF1 (N3710, N3706);
not NOT1 (N3711, N3709);
or OR4 (N3712, N3694, N1851, N1278, N1122);
xor XOR2 (N3713, N3710, N2178);
not NOT1 (N3714, N3711);
or OR4 (N3715, N3700, N1542, N3317, N1778);
not NOT1 (N3716, N3713);
buf BUF1 (N3717, N3716);
and AND2 (N3718, N3714, N831);
and AND4 (N3719, N3715, N2355, N2571, N1487);
nand NAND2 (N3720, N3712, N3512);
nor NOR2 (N3721, N3720, N834);
xor XOR2 (N3722, N3687, N1152);
and AND4 (N3723, N3708, N23, N1652, N75);
nand NAND4 (N3724, N3719, N51, N718, N406);
nand NAND3 (N3725, N3717, N3310, N330);
and AND3 (N3726, N3701, N1837, N2427);
not NOT1 (N3727, N3723);
nor NOR3 (N3728, N3693, N126, N2145);
nor NOR4 (N3729, N3718, N1480, N853, N761);
or OR2 (N3730, N3726, N2926);
or OR3 (N3731, N3730, N3682, N2773);
nand NAND3 (N3732, N3721, N1408, N2890);
or OR2 (N3733, N3707, N605);
buf BUF1 (N3734, N3728);
or OR3 (N3735, N3724, N3399, N429);
buf BUF1 (N3736, N3729);
nor NOR2 (N3737, N3722, N2722);
buf BUF1 (N3738, N3735);
nor NOR4 (N3739, N3734, N648, N2315, N253);
not NOT1 (N3740, N3727);
not NOT1 (N3741, N3738);
nor NOR2 (N3742, N3737, N2524);
or OR2 (N3743, N3740, N57);
xor XOR2 (N3744, N3731, N1846);
nand NAND4 (N3745, N3742, N1022, N3182, N1136);
not NOT1 (N3746, N3736);
xor XOR2 (N3747, N3746, N2582);
nor NOR4 (N3748, N3741, N592, N2064, N2224);
xor XOR2 (N3749, N3733, N2864);
buf BUF1 (N3750, N3743);
and AND3 (N3751, N3732, N3664, N3544);
xor XOR2 (N3752, N3739, N1743);
or OR3 (N3753, N3749, N3358, N3664);
buf BUF1 (N3754, N3704);
and AND4 (N3755, N3750, N1608, N3512, N3561);
not NOT1 (N3756, N3744);
nor NOR2 (N3757, N3745, N2811);
nor NOR2 (N3758, N3757, N3560);
nand NAND4 (N3759, N3756, N2542, N92, N1670);
nor NOR3 (N3760, N3753, N2030, N2792);
nand NAND4 (N3761, N3759, N1023, N2531, N3592);
nand NAND4 (N3762, N3751, N1221, N2809, N3740);
or OR2 (N3763, N3725, N1654);
xor XOR2 (N3764, N3747, N703);
not NOT1 (N3765, N3758);
not NOT1 (N3766, N3761);
nor NOR4 (N3767, N3763, N2542, N3466, N3559);
not NOT1 (N3768, N3760);
and AND2 (N3769, N3755, N2500);
and AND3 (N3770, N3769, N590, N1705);
not NOT1 (N3771, N3752);
nor NOR3 (N3772, N3771, N1173, N2413);
or OR2 (N3773, N3762, N2032);
not NOT1 (N3774, N3766);
and AND3 (N3775, N3774, N2000, N2517);
nand NAND2 (N3776, N3748, N1841);
and AND3 (N3777, N3754, N2318, N866);
or OR4 (N3778, N3772, N906, N3682, N3523);
xor XOR2 (N3779, N3767, N85);
or OR4 (N3780, N3768, N3133, N848, N3473);
not NOT1 (N3781, N3765);
buf BUF1 (N3782, N3777);
nor NOR4 (N3783, N3782, N223, N2066, N3031);
and AND3 (N3784, N3773, N96, N257);
buf BUF1 (N3785, N3775);
and AND3 (N3786, N3779, N3620, N619);
nor NOR4 (N3787, N3776, N1095, N3103, N327);
nand NAND2 (N3788, N3781, N190);
and AND4 (N3789, N3783, N15, N802, N626);
not NOT1 (N3790, N3786);
or OR2 (N3791, N3788, N566);
buf BUF1 (N3792, N3784);
not NOT1 (N3793, N3792);
nand NAND3 (N3794, N3791, N2130, N3530);
not NOT1 (N3795, N3780);
nand NAND3 (N3796, N3790, N1984, N1421);
not NOT1 (N3797, N3796);
and AND4 (N3798, N3794, N3273, N3052, N2985);
not NOT1 (N3799, N3770);
buf BUF1 (N3800, N3793);
nor NOR4 (N3801, N3785, N2037, N1440, N1847);
nand NAND3 (N3802, N3800, N2335, N3145);
or OR2 (N3803, N3795, N1407);
xor XOR2 (N3804, N3799, N577);
nand NAND4 (N3805, N3802, N1582, N2150, N1790);
or OR2 (N3806, N3789, N2190);
nand NAND2 (N3807, N3787, N745);
not NOT1 (N3808, N3797);
xor XOR2 (N3809, N3798, N3040);
or OR2 (N3810, N3805, N1912);
buf BUF1 (N3811, N3807);
nor NOR2 (N3812, N3811, N805);
xor XOR2 (N3813, N3803, N1594);
and AND2 (N3814, N3809, N3163);
not NOT1 (N3815, N3813);
or OR4 (N3816, N3814, N738, N242, N2057);
and AND2 (N3817, N3815, N588);
nand NAND4 (N3818, N3816, N120, N1384, N3165);
nand NAND3 (N3819, N3817, N970, N74);
buf BUF1 (N3820, N3804);
buf BUF1 (N3821, N3808);
buf BUF1 (N3822, N3801);
nor NOR3 (N3823, N3821, N3480, N3492);
nor NOR4 (N3824, N3778, N1431, N434, N2706);
not NOT1 (N3825, N3824);
nand NAND3 (N3826, N3812, N80, N3089);
not NOT1 (N3827, N3819);
or OR2 (N3828, N3810, N3732);
buf BUF1 (N3829, N3820);
buf BUF1 (N3830, N3818);
nand NAND4 (N3831, N3764, N836, N2172, N493);
nor NOR3 (N3832, N3825, N40, N766);
nor NOR4 (N3833, N3822, N1999, N1591, N53);
nor NOR2 (N3834, N3833, N701);
or OR3 (N3835, N3806, N504, N446);
or OR4 (N3836, N3827, N3035, N3242, N1017);
not NOT1 (N3837, N3826);
xor XOR2 (N3838, N3836, N406);
and AND3 (N3839, N3837, N2469, N1830);
buf BUF1 (N3840, N3831);
xor XOR2 (N3841, N3838, N1616);
or OR2 (N3842, N3828, N929);
nor NOR4 (N3843, N3839, N1528, N919, N1095);
nand NAND2 (N3844, N3843, N1797);
nand NAND4 (N3845, N3834, N3785, N581, N2870);
not NOT1 (N3846, N3842);
and AND3 (N3847, N3841, N522, N966);
or OR3 (N3848, N3845, N3800, N2196);
and AND3 (N3849, N3847, N423, N1351);
buf BUF1 (N3850, N3844);
buf BUF1 (N3851, N3823);
not NOT1 (N3852, N3851);
nor NOR2 (N3853, N3829, N2063);
xor XOR2 (N3854, N3840, N1628);
or OR2 (N3855, N3852, N3736);
buf BUF1 (N3856, N3835);
not NOT1 (N3857, N3848);
nor NOR4 (N3858, N3830, N3382, N2052, N3388);
not NOT1 (N3859, N3855);
and AND2 (N3860, N3849, N1032);
or OR4 (N3861, N3859, N728, N2999, N3382);
or OR2 (N3862, N3832, N467);
xor XOR2 (N3863, N3862, N1725);
xor XOR2 (N3864, N3857, N582);
not NOT1 (N3865, N3853);
buf BUF1 (N3866, N3865);
not NOT1 (N3867, N3866);
nand NAND3 (N3868, N3850, N175, N2272);
nand NAND4 (N3869, N3863, N3080, N3396, N2553);
nand NAND4 (N3870, N3861, N2537, N302, N608);
nand NAND2 (N3871, N3864, N2497);
xor XOR2 (N3872, N3868, N1277);
nand NAND4 (N3873, N3872, N1090, N267, N1588);
or OR3 (N3874, N3846, N3103, N2584);
not NOT1 (N3875, N3854);
not NOT1 (N3876, N3858);
not NOT1 (N3877, N3876);
or OR3 (N3878, N3856, N3552, N3029);
nand NAND3 (N3879, N3873, N29, N2426);
and AND4 (N3880, N3860, N2441, N1140, N2432);
and AND3 (N3881, N3879, N2707, N3741);
nand NAND4 (N3882, N3877, N1965, N3200, N2088);
not NOT1 (N3883, N3871);
nor NOR2 (N3884, N3883, N1512);
not NOT1 (N3885, N3884);
and AND2 (N3886, N3882, N633);
not NOT1 (N3887, N3885);
not NOT1 (N3888, N3870);
and AND4 (N3889, N3880, N1530, N3275, N3884);
and AND2 (N3890, N3888, N2889);
nand NAND3 (N3891, N3881, N1216, N2754);
nor NOR2 (N3892, N3889, N2752);
nor NOR2 (N3893, N3891, N782);
nor NOR4 (N3894, N3874, N2433, N830, N2599);
xor XOR2 (N3895, N3887, N1122);
nor NOR4 (N3896, N3875, N109, N2490, N2291);
nand NAND2 (N3897, N3890, N1736);
nor NOR2 (N3898, N3869, N3276);
xor XOR2 (N3899, N3892, N3691);
xor XOR2 (N3900, N3878, N801);
and AND2 (N3901, N3899, N3010);
buf BUF1 (N3902, N3894);
not NOT1 (N3903, N3896);
xor XOR2 (N3904, N3898, N3430);
xor XOR2 (N3905, N3897, N2814);
or OR2 (N3906, N3867, N2430);
nand NAND2 (N3907, N3895, N2432);
nor NOR4 (N3908, N3886, N1339, N2294, N1338);
buf BUF1 (N3909, N3901);
not NOT1 (N3910, N3900);
not NOT1 (N3911, N3910);
or OR2 (N3912, N3893, N640);
nand NAND3 (N3913, N3911, N1271, N2261);
buf BUF1 (N3914, N3909);
and AND4 (N3915, N3906, N1471, N548, N2538);
and AND2 (N3916, N3902, N1567);
xor XOR2 (N3917, N3915, N3768);
nand NAND3 (N3918, N3905, N2611, N1642);
nand NAND2 (N3919, N3917, N132);
nand NAND4 (N3920, N3919, N2628, N3354, N1812);
nand NAND3 (N3921, N3904, N34, N1613);
nor NOR3 (N3922, N3918, N2644, N387);
xor XOR2 (N3923, N3913, N3459);
nand NAND4 (N3924, N3908, N3254, N63, N2531);
nand NAND2 (N3925, N3903, N2549);
xor XOR2 (N3926, N3922, N3336);
and AND4 (N3927, N3920, N2713, N3746, N2347);
not NOT1 (N3928, N3916);
xor XOR2 (N3929, N3928, N130);
nand NAND2 (N3930, N3924, N3871);
or OR2 (N3931, N3929, N786);
not NOT1 (N3932, N3927);
buf BUF1 (N3933, N3930);
xor XOR2 (N3934, N3926, N3002);
buf BUF1 (N3935, N3932);
nor NOR2 (N3936, N3931, N3669);
and AND2 (N3937, N3921, N2326);
xor XOR2 (N3938, N3925, N2252);
not NOT1 (N3939, N3933);
nor NOR3 (N3940, N3935, N2633, N2737);
xor XOR2 (N3941, N3907, N3465);
xor XOR2 (N3942, N3937, N1021);
nor NOR4 (N3943, N3914, N742, N3857, N68);
nand NAND3 (N3944, N3939, N1385, N3099);
xor XOR2 (N3945, N3912, N2448);
or OR3 (N3946, N3938, N2253, N2160);
nor NOR4 (N3947, N3946, N2354, N1929, N3041);
or OR3 (N3948, N3943, N632, N909);
nand NAND3 (N3949, N3948, N1641, N2406);
nand NAND3 (N3950, N3934, N2294, N270);
not NOT1 (N3951, N3944);
nand NAND2 (N3952, N3936, N1584);
or OR4 (N3953, N3947, N2846, N2265, N1940);
and AND3 (N3954, N3951, N646, N879);
and AND3 (N3955, N3942, N1070, N3471);
or OR2 (N3956, N3923, N651);
not NOT1 (N3957, N3950);
nand NAND2 (N3958, N3957, N2147);
or OR3 (N3959, N3953, N3015, N484);
not NOT1 (N3960, N3958);
nor NOR3 (N3961, N3960, N1159, N3281);
or OR3 (N3962, N3940, N3528, N3676);
xor XOR2 (N3963, N3954, N780);
and AND3 (N3964, N3941, N1431, N3770);
or OR3 (N3965, N3959, N2540, N69);
not NOT1 (N3966, N3962);
nor NOR2 (N3967, N3964, N18);
xor XOR2 (N3968, N3967, N58);
and AND3 (N3969, N3966, N1145, N1631);
not NOT1 (N3970, N3955);
and AND3 (N3971, N3965, N2603, N1602);
not NOT1 (N3972, N3949);
xor XOR2 (N3973, N3969, N2636);
xor XOR2 (N3974, N3956, N1829);
buf BUF1 (N3975, N3974);
and AND3 (N3976, N3975, N1761, N2950);
buf BUF1 (N3977, N3971);
nand NAND2 (N3978, N3970, N1241);
not NOT1 (N3979, N3973);
nor NOR3 (N3980, N3961, N3201, N1289);
nor NOR2 (N3981, N3979, N664);
and AND4 (N3982, N3945, N66, N3401, N1926);
xor XOR2 (N3983, N3972, N310);
not NOT1 (N3984, N3977);
and AND4 (N3985, N3984, N2774, N2662, N3691);
or OR4 (N3986, N3983, N3185, N483, N1814);
xor XOR2 (N3987, N3980, N2520);
xor XOR2 (N3988, N3981, N2317);
buf BUF1 (N3989, N3986);
or OR4 (N3990, N3952, N3234, N683, N3647);
or OR4 (N3991, N3989, N2469, N3477, N3692);
nor NOR4 (N3992, N3985, N2261, N2015, N2892);
nor NOR3 (N3993, N3988, N3796, N3527);
buf BUF1 (N3994, N3982);
buf BUF1 (N3995, N3991);
or OR3 (N3996, N3995, N1768, N2183);
and AND3 (N3997, N3963, N666, N1665);
not NOT1 (N3998, N3997);
xor XOR2 (N3999, N3976, N263);
buf BUF1 (N4000, N3987);
xor XOR2 (N4001, N3968, N2497);
or OR2 (N4002, N3990, N1399);
buf BUF1 (N4003, N3998);
nand NAND2 (N4004, N4002, N2398);
buf BUF1 (N4005, N3996);
not NOT1 (N4006, N3999);
nor NOR2 (N4007, N4006, N3739);
and AND3 (N4008, N3978, N894, N1855);
and AND2 (N4009, N4003, N2243);
buf BUF1 (N4010, N4009);
and AND3 (N4011, N4001, N3227, N1879);
xor XOR2 (N4012, N4011, N2725);
buf BUF1 (N4013, N4010);
or OR3 (N4014, N3994, N2464, N3028);
buf BUF1 (N4015, N4004);
xor XOR2 (N4016, N4012, N2110);
nor NOR4 (N4017, N4016, N3609, N351, N204);
and AND4 (N4018, N3993, N3044, N558, N867);
buf BUF1 (N4019, N3992);
not NOT1 (N4020, N4008);
nor NOR2 (N4021, N4005, N3906);
nor NOR2 (N4022, N4019, N26);
buf BUF1 (N4023, N4007);
nor NOR2 (N4024, N4018, N155);
not NOT1 (N4025, N4017);
and AND4 (N4026, N4000, N2158, N466, N339);
and AND4 (N4027, N4013, N1310, N2135, N2608);
buf BUF1 (N4028, N4023);
not NOT1 (N4029, N4024);
nor NOR4 (N4030, N4029, N819, N2661, N78);
buf BUF1 (N4031, N4020);
nand NAND2 (N4032, N4030, N2911);
and AND4 (N4033, N4014, N2253, N1779, N1983);
xor XOR2 (N4034, N4025, N1566);
nor NOR3 (N4035, N4031, N3681, N161);
nor NOR3 (N4036, N4022, N1138, N2274);
nand NAND2 (N4037, N4032, N3120);
nor NOR3 (N4038, N4028, N2344, N737);
and AND2 (N4039, N4038, N3982);
not NOT1 (N4040, N4033);
nor NOR4 (N4041, N4026, N3910, N3394, N3078);
or OR2 (N4042, N4041, N3437);
nor NOR3 (N4043, N4042, N3752, N3930);
xor XOR2 (N4044, N4040, N2947);
or OR2 (N4045, N4021, N2608);
nor NOR2 (N4046, N4027, N293);
and AND3 (N4047, N4015, N2141, N853);
or OR3 (N4048, N4035, N3288, N3987);
and AND4 (N4049, N4048, N984, N2759, N3162);
xor XOR2 (N4050, N4039, N2273);
nor NOR3 (N4051, N4050, N3834, N683);
nand NAND3 (N4052, N4047, N1820, N2562);
and AND3 (N4053, N4044, N72, N3073);
nand NAND2 (N4054, N4049, N1046);
buf BUF1 (N4055, N4053);
nor NOR3 (N4056, N4055, N4025, N1267);
not NOT1 (N4057, N4043);
nand NAND4 (N4058, N4054, N3778, N68, N1384);
not NOT1 (N4059, N4034);
buf BUF1 (N4060, N4045);
nor NOR2 (N4061, N4046, N3605);
nor NOR4 (N4062, N4057, N3937, N2145, N2787);
and AND2 (N4063, N4058, N570);
buf BUF1 (N4064, N4061);
buf BUF1 (N4065, N4056);
buf BUF1 (N4066, N4062);
xor XOR2 (N4067, N4060, N733);
and AND4 (N4068, N4064, N1853, N2679, N373);
nand NAND4 (N4069, N4063, N3135, N2902, N3818);
buf BUF1 (N4070, N4069);
not NOT1 (N4071, N4052);
buf BUF1 (N4072, N4036);
xor XOR2 (N4073, N4072, N1996);
and AND4 (N4074, N4051, N1148, N2107, N1861);
buf BUF1 (N4075, N4067);
xor XOR2 (N4076, N4071, N1099);
not NOT1 (N4077, N4070);
not NOT1 (N4078, N4066);
not NOT1 (N4079, N4078);
xor XOR2 (N4080, N4059, N953);
nand NAND3 (N4081, N4076, N1423, N820);
and AND4 (N4082, N4080, N1927, N1454, N3196);
or OR2 (N4083, N4068, N3222);
nor NOR2 (N4084, N4075, N192);
nand NAND3 (N4085, N4084, N1890, N725);
buf BUF1 (N4086, N4079);
or OR3 (N4087, N4037, N283, N3474);
not NOT1 (N4088, N4074);
buf BUF1 (N4089, N4086);
not NOT1 (N4090, N4065);
nor NOR2 (N4091, N4085, N1236);
or OR4 (N4092, N4081, N2758, N4011, N1457);
buf BUF1 (N4093, N4090);
nor NOR4 (N4094, N4082, N3340, N1016, N2925);
not NOT1 (N4095, N4083);
buf BUF1 (N4096, N4087);
xor XOR2 (N4097, N4094, N592);
not NOT1 (N4098, N4095);
not NOT1 (N4099, N4077);
or OR2 (N4100, N4098, N2231);
and AND2 (N4101, N4092, N1707);
or OR2 (N4102, N4089, N2496);
buf BUF1 (N4103, N4097);
not NOT1 (N4104, N4088);
or OR4 (N4105, N4093, N1701, N867, N2056);
buf BUF1 (N4106, N4101);
and AND4 (N4107, N4091, N2099, N1787, N2294);
or OR2 (N4108, N4105, N922);
xor XOR2 (N4109, N4103, N837);
or OR3 (N4110, N4106, N3811, N2745);
buf BUF1 (N4111, N4100);
or OR3 (N4112, N4111, N1879, N493);
and AND3 (N4113, N4109, N2005, N572);
and AND4 (N4114, N4073, N2137, N3371, N2450);
xor XOR2 (N4115, N4104, N3398);
nand NAND2 (N4116, N4114, N2903);
or OR2 (N4117, N4112, N2913);
and AND3 (N4118, N4115, N279, N1321);
buf BUF1 (N4119, N4118);
nor NOR4 (N4120, N4102, N680, N463, N793);
xor XOR2 (N4121, N4120, N279);
buf BUF1 (N4122, N4121);
nand NAND3 (N4123, N4107, N1281, N2963);
and AND4 (N4124, N4119, N138, N3684, N2806);
nand NAND2 (N4125, N4113, N3867);
or OR2 (N4126, N4099, N1146);
not NOT1 (N4127, N4096);
not NOT1 (N4128, N4125);
buf BUF1 (N4129, N4127);
and AND2 (N4130, N4116, N1825);
nor NOR4 (N4131, N4126, N1870, N3534, N160);
buf BUF1 (N4132, N4130);
xor XOR2 (N4133, N4131, N2579);
buf BUF1 (N4134, N4128);
or OR2 (N4135, N4123, N1950);
nand NAND4 (N4136, N4135, N3401, N2072, N2335);
nand NAND4 (N4137, N4132, N2735, N1080, N1769);
and AND2 (N4138, N4122, N3592);
nand NAND3 (N4139, N4108, N843, N1312);
or OR3 (N4140, N4117, N3353, N3443);
buf BUF1 (N4141, N4110);
or OR3 (N4142, N4139, N2281, N3606);
buf BUF1 (N4143, N4142);
xor XOR2 (N4144, N4124, N1878);
xor XOR2 (N4145, N4136, N3515);
nor NOR2 (N4146, N4140, N2067);
nand NAND3 (N4147, N4129, N3872, N3371);
nand NAND3 (N4148, N4145, N174, N1912);
nor NOR3 (N4149, N4148, N1286, N2941);
and AND2 (N4150, N4144, N1714);
xor XOR2 (N4151, N4138, N3039);
xor XOR2 (N4152, N4141, N3691);
and AND2 (N4153, N4152, N3290);
not NOT1 (N4154, N4150);
not NOT1 (N4155, N4143);
nor NOR4 (N4156, N4153, N1881, N2454, N3375);
buf BUF1 (N4157, N4133);
nor NOR4 (N4158, N4155, N696, N633, N371);
nand NAND3 (N4159, N4157, N366, N1936);
nand NAND4 (N4160, N4156, N1302, N3200, N1429);
buf BUF1 (N4161, N4149);
nand NAND3 (N4162, N4134, N802, N1739);
and AND2 (N4163, N4162, N4);
nor NOR3 (N4164, N4163, N1351, N4052);
and AND3 (N4165, N4164, N854, N1438);
nor NOR2 (N4166, N4158, N861);
or OR4 (N4167, N4146, N138, N2687, N2309);
buf BUF1 (N4168, N4165);
or OR2 (N4169, N4147, N790);
xor XOR2 (N4170, N4166, N991);
and AND4 (N4171, N4151, N1407, N4071, N1098);
xor XOR2 (N4172, N4168, N1342);
or OR4 (N4173, N4172, N2827, N3567, N3949);
buf BUF1 (N4174, N4159);
nor NOR2 (N4175, N4174, N3193);
or OR2 (N4176, N4160, N1975);
or OR3 (N4177, N4175, N2420, N500);
and AND3 (N4178, N4137, N552, N491);
and AND4 (N4179, N4173, N2936, N343, N537);
and AND4 (N4180, N4177, N1125, N2375, N3108);
not NOT1 (N4181, N4171);
xor XOR2 (N4182, N4178, N1690);
nand NAND3 (N4183, N4167, N630, N2026);
buf BUF1 (N4184, N4179);
buf BUF1 (N4185, N4184);
or OR3 (N4186, N4170, N2473, N3585);
and AND4 (N4187, N4180, N1722, N343, N2062);
or OR2 (N4188, N4161, N3910);
nand NAND4 (N4189, N4186, N1259, N3796, N2027);
nor NOR3 (N4190, N4182, N2669, N874);
nor NOR2 (N4191, N4181, N433);
not NOT1 (N4192, N4176);
buf BUF1 (N4193, N4154);
buf BUF1 (N4194, N4192);
nor NOR3 (N4195, N4194, N1818, N613);
and AND3 (N4196, N4191, N3172, N91);
not NOT1 (N4197, N4188);
buf BUF1 (N4198, N4189);
not NOT1 (N4199, N4193);
and AND4 (N4200, N4187, N402, N3728, N644);
nand NAND4 (N4201, N4200, N3553, N3939, N2654);
or OR3 (N4202, N4199, N3508, N3927);
and AND2 (N4203, N4183, N2469);
nor NOR4 (N4204, N4203, N2285, N1199, N2634);
and AND3 (N4205, N4169, N1529, N3564);
nand NAND4 (N4206, N4202, N1339, N1727, N2715);
nand NAND3 (N4207, N4205, N1582, N289);
buf BUF1 (N4208, N4195);
not NOT1 (N4209, N4204);
and AND4 (N4210, N4207, N3408, N1142, N4156);
nor NOR4 (N4211, N4201, N4046, N1607, N1582);
buf BUF1 (N4212, N4196);
not NOT1 (N4213, N4206);
buf BUF1 (N4214, N4210);
or OR2 (N4215, N4190, N3281);
nor NOR3 (N4216, N4209, N2985, N923);
not NOT1 (N4217, N4215);
buf BUF1 (N4218, N4214);
nor NOR2 (N4219, N4185, N2946);
nor NOR2 (N4220, N4211, N3519);
or OR4 (N4221, N4197, N1294, N272, N1895);
or OR3 (N4222, N4198, N1841, N3009);
or OR4 (N4223, N4216, N3837, N413, N3973);
nand NAND2 (N4224, N4213, N2954);
not NOT1 (N4225, N4222);
xor XOR2 (N4226, N4217, N745);
nor NOR2 (N4227, N4220, N3315);
nand NAND4 (N4228, N4208, N1532, N2910, N383);
or OR3 (N4229, N4224, N2325, N3341);
nand NAND4 (N4230, N4225, N198, N2146, N668);
nand NAND4 (N4231, N4227, N961, N856, N308);
and AND4 (N4232, N4223, N1651, N3659, N1893);
or OR4 (N4233, N4212, N1631, N490, N3623);
buf BUF1 (N4234, N4232);
buf BUF1 (N4235, N4228);
xor XOR2 (N4236, N4221, N3530);
or OR4 (N4237, N4235, N174, N3134, N3789);
nand NAND2 (N4238, N4237, N761);
xor XOR2 (N4239, N4234, N3694);
buf BUF1 (N4240, N4230);
nor NOR4 (N4241, N4218, N910, N1807, N1802);
buf BUF1 (N4242, N4229);
or OR2 (N4243, N4238, N2792);
nand NAND3 (N4244, N4242, N2204, N4086);
or OR3 (N4245, N4231, N2468, N1225);
not NOT1 (N4246, N4240);
or OR3 (N4247, N4226, N3906, N1085);
nand NAND2 (N4248, N4236, N1065);
not NOT1 (N4249, N4244);
or OR3 (N4250, N4243, N256, N3026);
buf BUF1 (N4251, N4239);
nor NOR3 (N4252, N4245, N1047, N3759);
nor NOR2 (N4253, N4241, N1292);
buf BUF1 (N4254, N4249);
nor NOR3 (N4255, N4254, N2400, N841);
nand NAND2 (N4256, N4252, N61);
nor NOR3 (N4257, N4248, N2276, N53);
or OR4 (N4258, N4253, N3109, N1274, N3477);
nor NOR3 (N4259, N4247, N2895, N90);
buf BUF1 (N4260, N4233);
nand NAND3 (N4261, N4256, N2324, N4180);
buf BUF1 (N4262, N4259);
buf BUF1 (N4263, N4251);
not NOT1 (N4264, N4219);
xor XOR2 (N4265, N4261, N1454);
or OR2 (N4266, N4257, N624);
or OR3 (N4267, N4262, N15, N2928);
or OR3 (N4268, N4267, N2736, N1504);
and AND3 (N4269, N4255, N3954, N2909);
buf BUF1 (N4270, N4264);
and AND2 (N4271, N4258, N2262);
and AND4 (N4272, N4269, N2865, N381, N1220);
or OR2 (N4273, N4270, N1768);
or OR2 (N4274, N4266, N3233);
and AND4 (N4275, N4265, N3132, N2076, N3858);
nor NOR3 (N4276, N4268, N1755, N1579);
buf BUF1 (N4277, N4260);
xor XOR2 (N4278, N4273, N1047);
and AND4 (N4279, N4272, N2537, N2380, N2857);
xor XOR2 (N4280, N4276, N1631);
and AND2 (N4281, N4274, N2048);
not NOT1 (N4282, N4250);
nand NAND2 (N4283, N4271, N3509);
nand NAND3 (N4284, N4279, N1913, N1778);
nand NAND4 (N4285, N4280, N3650, N3504, N695);
or OR4 (N4286, N4277, N3202, N2664, N605);
nand NAND2 (N4287, N4278, N2811);
not NOT1 (N4288, N4285);
nand NAND2 (N4289, N4275, N1959);
or OR4 (N4290, N4289, N2881, N1357, N1354);
xor XOR2 (N4291, N4283, N1133);
nor NOR3 (N4292, N4286, N3715, N1627);
buf BUF1 (N4293, N4282);
nor NOR3 (N4294, N4246, N1927, N2919);
and AND3 (N4295, N4281, N1280, N1373);
xor XOR2 (N4296, N4294, N2043);
xor XOR2 (N4297, N4293, N3157);
nand NAND3 (N4298, N4297, N1542, N3820);
buf BUF1 (N4299, N4263);
and AND3 (N4300, N4295, N71, N2070);
buf BUF1 (N4301, N4299);
nor NOR4 (N4302, N4292, N557, N658, N3380);
nor NOR4 (N4303, N4296, N1665, N1585, N864);
or OR3 (N4304, N4300, N3464, N3710);
nand NAND3 (N4305, N4303, N3533, N3839);
nand NAND3 (N4306, N4305, N2505, N1671);
buf BUF1 (N4307, N4306);
or OR3 (N4308, N4284, N2159, N490);
or OR3 (N4309, N4304, N1531, N1727);
buf BUF1 (N4310, N4298);
nand NAND4 (N4311, N4291, N3285, N3642, N3206);
xor XOR2 (N4312, N4302, N1726);
nand NAND4 (N4313, N4290, N3902, N3416, N3409);
nand NAND2 (N4314, N4287, N3458);
nor NOR4 (N4315, N4313, N3005, N3520, N3811);
or OR3 (N4316, N4312, N370, N2313);
nand NAND2 (N4317, N4316, N319);
nand NAND4 (N4318, N4315, N534, N2066, N799);
nand NAND4 (N4319, N4307, N3682, N3084, N1083);
and AND2 (N4320, N4319, N3142);
buf BUF1 (N4321, N4310);
xor XOR2 (N4322, N4320, N2257);
buf BUF1 (N4323, N4311);
not NOT1 (N4324, N4309);
not NOT1 (N4325, N4308);
and AND2 (N4326, N4322, N555);
and AND2 (N4327, N4318, N3148);
nor NOR4 (N4328, N4327, N921, N336, N2569);
or OR4 (N4329, N4326, N2980, N3246, N87);
nor NOR2 (N4330, N4301, N949);
not NOT1 (N4331, N4330);
or OR2 (N4332, N4331, N3961);
nor NOR3 (N4333, N4332, N416, N3476);
not NOT1 (N4334, N4324);
xor XOR2 (N4335, N4314, N2388);
not NOT1 (N4336, N4288);
xor XOR2 (N4337, N4317, N1851);
nor NOR4 (N4338, N4335, N3305, N294, N3476);
not NOT1 (N4339, N4325);
or OR2 (N4340, N4334, N3121);
nand NAND4 (N4341, N4338, N3466, N173, N431);
buf BUF1 (N4342, N4321);
buf BUF1 (N4343, N4333);
nand NAND4 (N4344, N4323, N518, N1094, N2757);
and AND4 (N4345, N4339, N682, N1857, N3092);
and AND4 (N4346, N4328, N3467, N1271, N632);
not NOT1 (N4347, N4345);
or OR3 (N4348, N4340, N3927, N2705);
nor NOR2 (N4349, N4337, N254);
buf BUF1 (N4350, N4347);
xor XOR2 (N4351, N4342, N2511);
not NOT1 (N4352, N4343);
or OR4 (N4353, N4336, N1427, N1009, N581);
nand NAND3 (N4354, N4351, N3635, N3738);
not NOT1 (N4355, N4329);
or OR2 (N4356, N4353, N3716);
and AND4 (N4357, N4346, N416, N3228, N3028);
or OR3 (N4358, N4355, N3360, N3190);
and AND3 (N4359, N4349, N2140, N3544);
xor XOR2 (N4360, N4357, N1170);
nor NOR2 (N4361, N4359, N1235);
xor XOR2 (N4362, N4348, N1157);
xor XOR2 (N4363, N4361, N4071);
nand NAND3 (N4364, N4341, N4204, N1828);
xor XOR2 (N4365, N4362, N1793);
nand NAND3 (N4366, N4365, N4000, N1963);
not NOT1 (N4367, N4352);
xor XOR2 (N4368, N4344, N3448);
and AND2 (N4369, N4368, N1662);
or OR3 (N4370, N4354, N180, N4364);
or OR2 (N4371, N4098, N1457);
not NOT1 (N4372, N4350);
or OR4 (N4373, N4367, N32, N3882, N902);
xor XOR2 (N4374, N4363, N600);
or OR3 (N4375, N4370, N475, N123);
not NOT1 (N4376, N4369);
buf BUF1 (N4377, N4371);
not NOT1 (N4378, N4376);
or OR2 (N4379, N4356, N1269);
xor XOR2 (N4380, N4366, N1970);
buf BUF1 (N4381, N4358);
buf BUF1 (N4382, N4373);
or OR4 (N4383, N4374, N1416, N3991, N1579);
nand NAND4 (N4384, N4377, N2933, N3969, N1164);
buf BUF1 (N4385, N4360);
xor XOR2 (N4386, N4384, N3228);
nor NOR4 (N4387, N4385, N565, N4107, N1361);
not NOT1 (N4388, N4375);
buf BUF1 (N4389, N4386);
nor NOR2 (N4390, N4388, N3927);
buf BUF1 (N4391, N4382);
not NOT1 (N4392, N4387);
nor NOR3 (N4393, N4390, N2193, N1803);
buf BUF1 (N4394, N4389);
or OR4 (N4395, N4381, N1710, N4112, N2991);
nor NOR3 (N4396, N4395, N1779, N2995);
and AND4 (N4397, N4391, N3618, N2867, N1252);
and AND3 (N4398, N4397, N3118, N2757);
not NOT1 (N4399, N4379);
nor NOR2 (N4400, N4399, N2436);
xor XOR2 (N4401, N4394, N3151);
not NOT1 (N4402, N4383);
xor XOR2 (N4403, N4372, N503);
buf BUF1 (N4404, N4378);
buf BUF1 (N4405, N4404);
buf BUF1 (N4406, N4393);
not NOT1 (N4407, N4401);
xor XOR2 (N4408, N4400, N889);
nor NOR3 (N4409, N4406, N781, N1460);
not NOT1 (N4410, N4402);
or OR2 (N4411, N4407, N2252);
nand NAND4 (N4412, N4398, N3160, N3621, N3927);
or OR4 (N4413, N4380, N1148, N2222, N3359);
nor NOR2 (N4414, N4396, N3170);
nor NOR4 (N4415, N4403, N485, N1386, N1596);
or OR3 (N4416, N4412, N3070, N2053);
or OR4 (N4417, N4408, N3643, N2794, N43);
xor XOR2 (N4418, N4405, N14);
and AND2 (N4419, N4415, N1943);
nand NAND3 (N4420, N4410, N2362, N1462);
and AND4 (N4421, N4418, N2637, N3931, N3813);
not NOT1 (N4422, N4409);
nor NOR4 (N4423, N4420, N3502, N3023, N1896);
not NOT1 (N4424, N4423);
nor NOR4 (N4425, N4422, N2014, N1313, N2899);
and AND4 (N4426, N4416, N1083, N4338, N2703);
buf BUF1 (N4427, N4424);
buf BUF1 (N4428, N4392);
xor XOR2 (N4429, N4425, N2463);
and AND3 (N4430, N4417, N1847, N2121);
and AND3 (N4431, N4428, N157, N384);
xor XOR2 (N4432, N4414, N1109);
and AND4 (N4433, N4429, N57, N2104, N3479);
not NOT1 (N4434, N4411);
buf BUF1 (N4435, N4413);
not NOT1 (N4436, N4434);
buf BUF1 (N4437, N4433);
and AND4 (N4438, N4432, N1252, N1306, N2741);
and AND3 (N4439, N4421, N3486, N3642);
not NOT1 (N4440, N4437);
xor XOR2 (N4441, N4427, N33);
nand NAND3 (N4442, N4431, N609, N191);
and AND3 (N4443, N4430, N2313, N3297);
not NOT1 (N4444, N4439);
nor NOR3 (N4445, N4438, N580, N1644);
or OR4 (N4446, N4441, N531, N3473, N2401);
nor NOR4 (N4447, N4443, N25, N600, N635);
buf BUF1 (N4448, N4436);
not NOT1 (N4449, N4445);
and AND2 (N4450, N4448, N342);
nor NOR2 (N4451, N4447, N1631);
buf BUF1 (N4452, N4446);
nor NOR3 (N4453, N4449, N3188, N2518);
xor XOR2 (N4454, N4419, N4350);
nor NOR3 (N4455, N4451, N1184, N3991);
nor NOR3 (N4456, N4444, N3164, N2540);
and AND4 (N4457, N4435, N3227, N987, N1127);
and AND3 (N4458, N4457, N3722, N4242);
xor XOR2 (N4459, N4453, N4258);
or OR4 (N4460, N4459, N2813, N1318, N4227);
buf BUF1 (N4461, N4455);
nor NOR4 (N4462, N4460, N1606, N1817, N2727);
xor XOR2 (N4463, N4440, N1126);
not NOT1 (N4464, N4462);
buf BUF1 (N4465, N4426);
nand NAND2 (N4466, N4458, N1966);
not NOT1 (N4467, N4442);
nand NAND4 (N4468, N4454, N1508, N47, N4082);
nor NOR2 (N4469, N4463, N1742);
not NOT1 (N4470, N4464);
not NOT1 (N4471, N4461);
and AND3 (N4472, N4466, N2930, N3342);
nor NOR2 (N4473, N4467, N3112);
buf BUF1 (N4474, N4452);
or OR2 (N4475, N4472, N4241);
xor XOR2 (N4476, N4471, N144);
not NOT1 (N4477, N4465);
and AND4 (N4478, N4474, N2057, N159, N680);
nand NAND3 (N4479, N4470, N730, N2882);
and AND2 (N4480, N4456, N1900);
xor XOR2 (N4481, N4476, N727);
xor XOR2 (N4482, N4477, N1446);
and AND2 (N4483, N4475, N503);
nand NAND4 (N4484, N4483, N2770, N1651, N2443);
or OR4 (N4485, N4473, N41, N553, N1939);
or OR2 (N4486, N4482, N273);
nor NOR3 (N4487, N4469, N314, N4143);
nor NOR2 (N4488, N4486, N378);
and AND2 (N4489, N4479, N1586);
not NOT1 (N4490, N4468);
and AND2 (N4491, N4480, N2502);
buf BUF1 (N4492, N4481);
or OR2 (N4493, N4485, N1394);
not NOT1 (N4494, N4491);
nor NOR3 (N4495, N4488, N3595, N2552);
buf BUF1 (N4496, N4489);
nand NAND3 (N4497, N4493, N4014, N2980);
xor XOR2 (N4498, N4496, N2331);
nor NOR4 (N4499, N4497, N1162, N2741, N2051);
nor NOR3 (N4500, N4495, N1659, N3701);
xor XOR2 (N4501, N4490, N3237);
and AND3 (N4502, N4492, N3300, N4001);
nand NAND2 (N4503, N4484, N2887);
and AND3 (N4504, N4501, N231, N2385);
and AND4 (N4505, N4502, N4387, N3336, N752);
and AND2 (N4506, N4505, N179);
xor XOR2 (N4507, N4499, N3345);
buf BUF1 (N4508, N4504);
nor NOR4 (N4509, N4508, N2, N266, N1617);
nand NAND2 (N4510, N4503, N2044);
buf BUF1 (N4511, N4498);
xor XOR2 (N4512, N4494, N1945);
buf BUF1 (N4513, N4478);
xor XOR2 (N4514, N4487, N1326);
or OR3 (N4515, N4509, N1899, N567);
xor XOR2 (N4516, N4513, N1755);
xor XOR2 (N4517, N4511, N1014);
nor NOR2 (N4518, N4450, N404);
and AND3 (N4519, N4500, N3259, N3029);
nand NAND4 (N4520, N4518, N3028, N33, N1768);
and AND3 (N4521, N4510, N2696, N4097);
not NOT1 (N4522, N4515);
or OR4 (N4523, N4520, N2003, N2514, N505);
xor XOR2 (N4524, N4516, N3519);
nand NAND3 (N4525, N4517, N2164, N1911);
not NOT1 (N4526, N4519);
and AND2 (N4527, N4524, N3303);
and AND2 (N4528, N4527, N190);
xor XOR2 (N4529, N4523, N1629);
nand NAND4 (N4530, N4506, N798, N1148, N1376);
nand NAND3 (N4531, N4514, N3682, N581);
and AND4 (N4532, N4526, N1003, N738, N3357);
xor XOR2 (N4533, N4522, N4399);
nand NAND4 (N4534, N4507, N3477, N1635, N2675);
nor NOR4 (N4535, N4531, N3595, N4354, N150);
or OR2 (N4536, N4528, N4233);
not NOT1 (N4537, N4535);
and AND4 (N4538, N4512, N4409, N869, N619);
nor NOR3 (N4539, N4534, N1863, N1327);
or OR3 (N4540, N4525, N2617, N2505);
nor NOR4 (N4541, N4532, N2544, N2660, N1293);
nand NAND4 (N4542, N4537, N517, N1182, N1297);
xor XOR2 (N4543, N4536, N1962);
or OR4 (N4544, N4538, N2982, N4215, N2944);
xor XOR2 (N4545, N4529, N57);
and AND4 (N4546, N4543, N738, N1414, N2362);
and AND4 (N4547, N4530, N958, N1747, N2692);
nor NOR4 (N4548, N4545, N1055, N4052, N1494);
buf BUF1 (N4549, N4540);
nor NOR2 (N4550, N4547, N3379);
nor NOR2 (N4551, N4550, N262);
not NOT1 (N4552, N4546);
or OR3 (N4553, N4548, N1754, N4514);
not NOT1 (N4554, N4552);
nor NOR3 (N4555, N4551, N4128, N2345);
or OR2 (N4556, N4541, N2560);
buf BUF1 (N4557, N4521);
nor NOR4 (N4558, N4539, N4143, N4254, N1364);
xor XOR2 (N4559, N4554, N3995);
and AND4 (N4560, N4555, N1432, N4448, N383);
buf BUF1 (N4561, N4553);
nor NOR3 (N4562, N4549, N51, N3461);
or OR2 (N4563, N4557, N3166);
nand NAND3 (N4564, N4544, N4338, N2798);
nand NAND4 (N4565, N4561, N1404, N2867, N3011);
and AND2 (N4566, N4556, N3074);
not NOT1 (N4567, N4565);
not NOT1 (N4568, N4564);
xor XOR2 (N4569, N4542, N3346);
or OR4 (N4570, N4563, N4061, N2029, N4513);
not NOT1 (N4571, N4558);
nand NAND4 (N4572, N4568, N181, N1805, N3383);
not NOT1 (N4573, N4567);
nor NOR2 (N4574, N4570, N3738);
not NOT1 (N4575, N4562);
nor NOR4 (N4576, N4559, N4506, N1666, N2937);
buf BUF1 (N4577, N4576);
xor XOR2 (N4578, N4566, N4250);
xor XOR2 (N4579, N4577, N499);
nand NAND4 (N4580, N4571, N1926, N1594, N2261);
and AND4 (N4581, N4573, N895, N4405, N3126);
and AND3 (N4582, N4579, N3916, N4346);
xor XOR2 (N4583, N4582, N1381);
nor NOR4 (N4584, N4533, N3611, N2120, N3830);
xor XOR2 (N4585, N4578, N916);
xor XOR2 (N4586, N4574, N463);
nor NOR3 (N4587, N4584, N3436, N2692);
nor NOR4 (N4588, N4560, N3841, N1124, N555);
nand NAND3 (N4589, N4572, N1734, N2849);
and AND2 (N4590, N4575, N2359);
and AND4 (N4591, N4590, N4049, N1658, N1378);
and AND2 (N4592, N4569, N2921);
not NOT1 (N4593, N4585);
or OR4 (N4594, N4592, N4518, N2685, N2997);
and AND4 (N4595, N4587, N4410, N4215, N225);
or OR4 (N4596, N4593, N2956, N3139, N4468);
nor NOR3 (N4597, N4594, N4379, N4435);
nand NAND3 (N4598, N4591, N2792, N808);
nor NOR3 (N4599, N4595, N102, N3070);
nor NOR4 (N4600, N4598, N1780, N2797, N4344);
or OR2 (N4601, N4596, N1326);
or OR2 (N4602, N4580, N643);
nand NAND3 (N4603, N4581, N1213, N1287);
and AND2 (N4604, N4603, N846);
xor XOR2 (N4605, N4588, N369);
or OR4 (N4606, N4605, N2471, N4583, N76);
buf BUF1 (N4607, N233);
nor NOR2 (N4608, N4607, N601);
not NOT1 (N4609, N4606);
buf BUF1 (N4610, N4609);
xor XOR2 (N4611, N4610, N479);
or OR4 (N4612, N4589, N2523, N4480, N3220);
and AND3 (N4613, N4611, N239, N3778);
nor NOR4 (N4614, N4604, N2867, N2645, N3643);
nand NAND4 (N4615, N4599, N4374, N2119, N1844);
xor XOR2 (N4616, N4601, N291);
or OR4 (N4617, N4615, N4004, N705, N4051);
or OR2 (N4618, N4613, N3480);
buf BUF1 (N4619, N4616);
or OR2 (N4620, N4614, N286);
and AND3 (N4621, N4602, N3629, N115);
or OR3 (N4622, N4600, N256, N1226);
nor NOR3 (N4623, N4586, N2431, N4192);
or OR4 (N4624, N4622, N2439, N572, N3694);
and AND3 (N4625, N4623, N1396, N166);
and AND3 (N4626, N4612, N1092, N1360);
nand NAND2 (N4627, N4608, N2734);
nor NOR3 (N4628, N4625, N2700, N3702);
nand NAND4 (N4629, N4619, N2117, N2583, N1945);
buf BUF1 (N4630, N4620);
xor XOR2 (N4631, N4627, N3902);
not NOT1 (N4632, N4621);
and AND2 (N4633, N4618, N38);
and AND4 (N4634, N4630, N4606, N4330, N4582);
buf BUF1 (N4635, N4634);
nand NAND2 (N4636, N4633, N2934);
nand NAND2 (N4637, N4628, N3918);
buf BUF1 (N4638, N4636);
not NOT1 (N4639, N4638);
xor XOR2 (N4640, N4635, N1291);
buf BUF1 (N4641, N4637);
xor XOR2 (N4642, N4597, N4477);
or OR2 (N4643, N4629, N2454);
and AND3 (N4644, N4640, N317, N2440);
or OR4 (N4645, N4643, N2428, N555, N2621);
and AND2 (N4646, N4642, N1288);
nand NAND3 (N4647, N4646, N444, N4297);
and AND4 (N4648, N4624, N3279, N4251, N3232);
not NOT1 (N4649, N4648);
xor XOR2 (N4650, N4626, N4434);
buf BUF1 (N4651, N4650);
not NOT1 (N4652, N4645);
and AND4 (N4653, N4651, N2493, N2946, N3970);
nand NAND2 (N4654, N4639, N1080);
nor NOR2 (N4655, N4654, N4584);
nand NAND4 (N4656, N4649, N410, N4051, N1073);
and AND4 (N4657, N4631, N1278, N422, N3435);
buf BUF1 (N4658, N4656);
or OR2 (N4659, N4655, N4355);
or OR4 (N4660, N4617, N2152, N1511, N3903);
nor NOR4 (N4661, N4659, N1606, N3556, N368);
and AND3 (N4662, N4658, N1445, N1908);
and AND2 (N4663, N4662, N3062);
xor XOR2 (N4664, N4644, N2108);
not NOT1 (N4665, N4664);
and AND3 (N4666, N4663, N3712, N6);
xor XOR2 (N4667, N4665, N2024);
and AND3 (N4668, N4652, N1432, N2164);
nor NOR4 (N4669, N4667, N3112, N1525, N2131);
xor XOR2 (N4670, N4660, N93);
xor XOR2 (N4671, N4647, N1114);
nor NOR4 (N4672, N4666, N2279, N824, N2640);
nand NAND2 (N4673, N4672, N1694);
xor XOR2 (N4674, N4657, N2683);
nor NOR2 (N4675, N4641, N2312);
buf BUF1 (N4676, N4653);
xor XOR2 (N4677, N4676, N4458);
nor NOR4 (N4678, N4671, N4501, N4393, N856);
or OR4 (N4679, N4673, N765, N1662, N2993);
not NOT1 (N4680, N4669);
and AND3 (N4681, N4678, N2791, N2754);
nor NOR4 (N4682, N4681, N2656, N3462, N2253);
xor XOR2 (N4683, N4680, N3267);
xor XOR2 (N4684, N4675, N3454);
or OR4 (N4685, N4677, N2229, N2959, N2162);
not NOT1 (N4686, N4668);
and AND2 (N4687, N4661, N4608);
nand NAND3 (N4688, N4685, N3712, N775);
and AND4 (N4689, N4632, N1160, N1179, N2757);
and AND4 (N4690, N4686, N2909, N3289, N969);
and AND4 (N4691, N4679, N123, N1346, N3556);
buf BUF1 (N4692, N4689);
nor NOR3 (N4693, N4683, N3631, N2505);
nand NAND4 (N4694, N4684, N767, N4205, N431);
not NOT1 (N4695, N4690);
nand NAND2 (N4696, N4674, N4376);
nor NOR3 (N4697, N4670, N2592, N1417);
and AND4 (N4698, N4687, N2015, N4538, N3492);
not NOT1 (N4699, N4696);
and AND4 (N4700, N4692, N2042, N4575, N4595);
buf BUF1 (N4701, N4688);
nand NAND3 (N4702, N4700, N4338, N2964);
not NOT1 (N4703, N4698);
and AND3 (N4704, N4691, N649, N1011);
and AND4 (N4705, N4701, N4072, N965, N3760);
not NOT1 (N4706, N4705);
not NOT1 (N4707, N4706);
or OR4 (N4708, N4704, N2147, N1927, N2089);
nor NOR2 (N4709, N4694, N4654);
or OR2 (N4710, N4699, N1617);
xor XOR2 (N4711, N4709, N1034);
buf BUF1 (N4712, N4703);
nor NOR3 (N4713, N4711, N3617, N949);
nor NOR4 (N4714, N4710, N3255, N872, N1680);
or OR3 (N4715, N4682, N2402, N3835);
xor XOR2 (N4716, N4713, N2928);
nor NOR2 (N4717, N4715, N4387);
or OR2 (N4718, N4693, N3137);
and AND2 (N4719, N4702, N4685);
not NOT1 (N4720, N4719);
and AND4 (N4721, N4708, N3944, N4115, N1685);
and AND3 (N4722, N4707, N2761, N4301);
nand NAND4 (N4723, N4712, N4081, N2436, N2605);
buf BUF1 (N4724, N4722);
nor NOR3 (N4725, N4721, N2779, N270);
buf BUF1 (N4726, N4724);
nand NAND2 (N4727, N4725, N3041);
not NOT1 (N4728, N4716);
xor XOR2 (N4729, N4697, N1464);
xor XOR2 (N4730, N4695, N4355);
and AND2 (N4731, N4723, N1369);
nor NOR4 (N4732, N4727, N4156, N3848, N2146);
xor XOR2 (N4733, N4720, N3218);
or OR3 (N4734, N4728, N3369, N4179);
xor XOR2 (N4735, N4731, N2167);
not NOT1 (N4736, N4729);
and AND3 (N4737, N4732, N1383, N3891);
or OR2 (N4738, N4717, N3076);
and AND2 (N4739, N4736, N4104);
not NOT1 (N4740, N4734);
and AND4 (N4741, N4730, N3303, N3994, N3668);
nor NOR2 (N4742, N4737, N1173);
and AND3 (N4743, N4733, N1452, N797);
buf BUF1 (N4744, N4718);
buf BUF1 (N4745, N4739);
or OR2 (N4746, N4738, N2556);
buf BUF1 (N4747, N4744);
and AND3 (N4748, N4743, N2368, N1254);
not NOT1 (N4749, N4741);
nor NOR3 (N4750, N4726, N4360, N1120);
xor XOR2 (N4751, N4714, N1049);
buf BUF1 (N4752, N4750);
not NOT1 (N4753, N4752);
nor NOR4 (N4754, N4747, N792, N839, N4673);
or OR4 (N4755, N4754, N3315, N1700, N975);
buf BUF1 (N4756, N4742);
nor NOR2 (N4757, N4735, N1638);
xor XOR2 (N4758, N4755, N2776);
buf BUF1 (N4759, N4746);
not NOT1 (N4760, N4745);
nor NOR3 (N4761, N4748, N3822, N2052);
buf BUF1 (N4762, N4757);
and AND4 (N4763, N4759, N3462, N591, N3347);
not NOT1 (N4764, N4740);
and AND2 (N4765, N4761, N143);
buf BUF1 (N4766, N4760);
xor XOR2 (N4767, N4751, N2979);
xor XOR2 (N4768, N4756, N729);
or OR4 (N4769, N4765, N4193, N3954, N4569);
nand NAND3 (N4770, N4763, N3295, N2362);
not NOT1 (N4771, N4769);
not NOT1 (N4772, N4767);
not NOT1 (N4773, N4762);
and AND3 (N4774, N4772, N4555, N80);
xor XOR2 (N4775, N4753, N4065);
not NOT1 (N4776, N4768);
not NOT1 (N4777, N4758);
or OR4 (N4778, N4766, N1523, N4001, N407);
xor XOR2 (N4779, N4770, N2386);
or OR2 (N4780, N4778, N3793);
nor NOR2 (N4781, N4777, N1299);
not NOT1 (N4782, N4749);
and AND3 (N4783, N4773, N1785, N1173);
not NOT1 (N4784, N4781);
not NOT1 (N4785, N4783);
buf BUF1 (N4786, N4771);
buf BUF1 (N4787, N4774);
xor XOR2 (N4788, N4780, N4444);
xor XOR2 (N4789, N4764, N1958);
nor NOR2 (N4790, N4786, N212);
and AND4 (N4791, N4776, N1822, N2258, N2076);
buf BUF1 (N4792, N4789);
nand NAND3 (N4793, N4784, N265, N4311);
or OR3 (N4794, N4793, N732, N4717);
nor NOR3 (N4795, N4775, N3273, N2560);
nor NOR2 (N4796, N4788, N2842);
and AND4 (N4797, N4791, N3246, N3401, N4411);
nor NOR2 (N4798, N4792, N4325);
nor NOR4 (N4799, N4790, N4618, N148, N3250);
xor XOR2 (N4800, N4779, N531);
nand NAND4 (N4801, N4799, N2178, N1729, N1903);
nor NOR4 (N4802, N4795, N952, N4271, N604);
not NOT1 (N4803, N4797);
not NOT1 (N4804, N4798);
and AND3 (N4805, N4796, N3829, N3621);
nand NAND3 (N4806, N4803, N3009, N3161);
not NOT1 (N4807, N4805);
nand NAND2 (N4808, N4807, N1233);
xor XOR2 (N4809, N4787, N4535);
xor XOR2 (N4810, N4809, N161);
nand NAND2 (N4811, N4806, N317);
xor XOR2 (N4812, N4810, N2978);
xor XOR2 (N4813, N4794, N1102);
nand NAND3 (N4814, N4782, N2184, N2589);
or OR2 (N4815, N4801, N3753);
and AND4 (N4816, N4800, N2202, N3118, N1833);
nor NOR2 (N4817, N4812, N2573);
and AND2 (N4818, N4817, N1384);
nor NOR3 (N4819, N4785, N2613, N760);
nor NOR2 (N4820, N4819, N3138);
buf BUF1 (N4821, N4802);
nand NAND3 (N4822, N4811, N1231, N3205);
nor NOR4 (N4823, N4814, N3250, N3376, N1439);
nand NAND4 (N4824, N4820, N4244, N2125, N3076);
or OR4 (N4825, N4821, N1445, N2965, N2813);
buf BUF1 (N4826, N4822);
nor NOR3 (N4827, N4825, N4172, N1986);
and AND4 (N4828, N4818, N4211, N1392, N3497);
and AND3 (N4829, N4808, N3065, N148);
not NOT1 (N4830, N4823);
or OR2 (N4831, N4816, N3754);
not NOT1 (N4832, N4829);
buf BUF1 (N4833, N4826);
xor XOR2 (N4834, N4832, N2120);
and AND4 (N4835, N4833, N3973, N375, N223);
and AND3 (N4836, N4815, N1486, N4377);
and AND2 (N4837, N4824, N2353);
xor XOR2 (N4838, N4836, N865);
or OR3 (N4839, N4838, N4069, N4430);
buf BUF1 (N4840, N4834);
xor XOR2 (N4841, N4837, N4688);
xor XOR2 (N4842, N4840, N3152);
buf BUF1 (N4843, N4827);
nand NAND2 (N4844, N4830, N757);
nand NAND4 (N4845, N4828, N1790, N1451, N1036);
nor NOR3 (N4846, N4804, N2887, N4378);
nand NAND2 (N4847, N4831, N2365);
nand NAND4 (N4848, N4839, N3871, N401, N538);
buf BUF1 (N4849, N4844);
buf BUF1 (N4850, N4835);
nand NAND2 (N4851, N4850, N387);
nor NOR2 (N4852, N4845, N4446);
not NOT1 (N4853, N4847);
or OR2 (N4854, N4843, N1483);
xor XOR2 (N4855, N4853, N1106);
not NOT1 (N4856, N4813);
nor NOR3 (N4857, N4856, N588, N1657);
not NOT1 (N4858, N4841);
or OR2 (N4859, N4851, N1417);
xor XOR2 (N4860, N4852, N3153);
nand NAND2 (N4861, N4858, N363);
not NOT1 (N4862, N4859);
buf BUF1 (N4863, N4848);
nand NAND3 (N4864, N4860, N3007, N1809);
not NOT1 (N4865, N4857);
and AND3 (N4866, N4864, N10, N1891);
nand NAND3 (N4867, N4846, N280, N2164);
xor XOR2 (N4868, N4849, N3349);
nand NAND4 (N4869, N4863, N2922, N3818, N2984);
nor NOR2 (N4870, N4854, N3188);
buf BUF1 (N4871, N4865);
nor NOR4 (N4872, N4855, N2137, N4794, N4766);
buf BUF1 (N4873, N4870);
nand NAND2 (N4874, N4873, N4558);
nor NOR4 (N4875, N4861, N4395, N1844, N3403);
and AND3 (N4876, N4866, N4426, N4332);
buf BUF1 (N4877, N4869);
and AND3 (N4878, N4867, N512, N824);
buf BUF1 (N4879, N4868);
buf BUF1 (N4880, N4876);
not NOT1 (N4881, N4878);
buf BUF1 (N4882, N4871);
buf BUF1 (N4883, N4882);
buf BUF1 (N4884, N4879);
buf BUF1 (N4885, N4883);
nor NOR3 (N4886, N4881, N991, N1655);
and AND3 (N4887, N4872, N2033, N3800);
and AND4 (N4888, N4877, N1530, N1101, N1015);
or OR3 (N4889, N4888, N3124, N4445);
xor XOR2 (N4890, N4880, N1687);
nand NAND4 (N4891, N4889, N3406, N575, N3022);
not NOT1 (N4892, N4891);
nand NAND2 (N4893, N4884, N4299);
not NOT1 (N4894, N4886);
and AND3 (N4895, N4875, N4233, N4051);
and AND4 (N4896, N4893, N4360, N2498, N1226);
nand NAND4 (N4897, N4894, N469, N4497, N486);
and AND4 (N4898, N4890, N1402, N214, N4084);
nand NAND4 (N4899, N4842, N4759, N2278, N3784);
buf BUF1 (N4900, N4885);
and AND2 (N4901, N4892, N2788);
nand NAND2 (N4902, N4897, N2280);
nand NAND4 (N4903, N4900, N2276, N369, N4652);
or OR3 (N4904, N4887, N1691, N2936);
nor NOR2 (N4905, N4903, N3694);
buf BUF1 (N4906, N4874);
or OR4 (N4907, N4905, N3118, N4070, N4145);
and AND4 (N4908, N4904, N4101, N4817, N3340);
buf BUF1 (N4909, N4898);
buf BUF1 (N4910, N4895);
not NOT1 (N4911, N4899);
and AND4 (N4912, N4910, N4493, N809, N3744);
and AND3 (N4913, N4908, N2409, N4441);
buf BUF1 (N4914, N4902);
not NOT1 (N4915, N4914);
xor XOR2 (N4916, N4896, N4860);
buf BUF1 (N4917, N4862);
or OR4 (N4918, N4915, N3231, N1586, N471);
not NOT1 (N4919, N4909);
buf BUF1 (N4920, N4901);
xor XOR2 (N4921, N4906, N2303);
buf BUF1 (N4922, N4920);
nand NAND4 (N4923, N4912, N3872, N3117, N1427);
buf BUF1 (N4924, N4913);
nor NOR4 (N4925, N4923, N1180, N3, N1315);
buf BUF1 (N4926, N4917);
and AND4 (N4927, N4911, N359, N224, N4284);
nor NOR4 (N4928, N4919, N3615, N4772, N130);
buf BUF1 (N4929, N4924);
buf BUF1 (N4930, N4929);
or OR2 (N4931, N4927, N3972);
nor NOR4 (N4932, N4921, N3341, N4174, N3223);
and AND4 (N4933, N4932, N1460, N1862, N3855);
nor NOR4 (N4934, N4933, N3345, N2574, N768);
not NOT1 (N4935, N4934);
buf BUF1 (N4936, N4916);
nor NOR2 (N4937, N4907, N1242);
nor NOR2 (N4938, N4931, N2913);
and AND3 (N4939, N4937, N1814, N1866);
not NOT1 (N4940, N4918);
xor XOR2 (N4941, N4930, N3031);
nand NAND3 (N4942, N4936, N2706, N1760);
not NOT1 (N4943, N4942);
nor NOR3 (N4944, N4941, N4107, N3677);
or OR4 (N4945, N4928, N1155, N3496, N64);
buf BUF1 (N4946, N4939);
nor NOR2 (N4947, N4940, N4328);
buf BUF1 (N4948, N4946);
not NOT1 (N4949, N4944);
nor NOR4 (N4950, N4949, N3256, N242, N3605);
nand NAND3 (N4951, N4926, N3466, N3353);
or OR4 (N4952, N4922, N4231, N2211, N3587);
not NOT1 (N4953, N4951);
xor XOR2 (N4954, N4950, N695);
xor XOR2 (N4955, N4925, N2162);
and AND2 (N4956, N4935, N584);
buf BUF1 (N4957, N4953);
not NOT1 (N4958, N4945);
or OR2 (N4959, N4954, N4693);
nand NAND2 (N4960, N4947, N2556);
not NOT1 (N4961, N4959);
and AND3 (N4962, N4938, N38, N4408);
xor XOR2 (N4963, N4952, N366);
and AND3 (N4964, N4955, N2445, N1809);
or OR2 (N4965, N4948, N2931);
or OR2 (N4966, N4963, N3495);
and AND3 (N4967, N4964, N839, N1527);
and AND2 (N4968, N4966, N4781);
xor XOR2 (N4969, N4957, N1810);
nand NAND3 (N4970, N4967, N1329, N2993);
nand NAND4 (N4971, N4943, N1509, N1828, N4545);
buf BUF1 (N4972, N4969);
xor XOR2 (N4973, N4961, N582);
nor NOR2 (N4974, N4971, N4266);
nand NAND2 (N4975, N4974, N1870);
nand NAND4 (N4976, N4968, N717, N3713, N994);
and AND4 (N4977, N4960, N3704, N1050, N3990);
and AND2 (N4978, N4956, N3864);
buf BUF1 (N4979, N4958);
nor NOR4 (N4980, N4973, N3922, N1807, N4147);
and AND4 (N4981, N4976, N2915, N661, N1977);
buf BUF1 (N4982, N4972);
nand NAND3 (N4983, N4980, N3695, N981);
or OR3 (N4984, N4982, N3166, N2518);
nor NOR3 (N4985, N4978, N2203, N50);
buf BUF1 (N4986, N4983);
nor NOR2 (N4987, N4975, N913);
xor XOR2 (N4988, N4962, N1210);
or OR4 (N4989, N4988, N1230, N2673, N4401);
and AND3 (N4990, N4979, N2297, N619);
and AND3 (N4991, N4990, N4284, N2579);
or OR4 (N4992, N4981, N2053, N1954, N36);
and AND3 (N4993, N4970, N3268, N1155);
or OR4 (N4994, N4986, N3193, N4297, N2230);
and AND4 (N4995, N4977, N941, N1484, N4101);
not NOT1 (N4996, N4989);
and AND4 (N4997, N4984, N4906, N59, N119);
not NOT1 (N4998, N4965);
nor NOR3 (N4999, N4995, N3544, N1955);
buf BUF1 (N5000, N4998);
nor NOR3 (N5001, N4996, N4476, N3085);
nor NOR3 (N5002, N4994, N3995, N3209);
not NOT1 (N5003, N5000);
xor XOR2 (N5004, N4993, N4928);
nand NAND3 (N5005, N5002, N4755, N3708);
not NOT1 (N5006, N4987);
not NOT1 (N5007, N5006);
or OR3 (N5008, N4991, N1043, N3280);
buf BUF1 (N5009, N5007);
xor XOR2 (N5010, N4985, N4742);
nor NOR4 (N5011, N4999, N1938, N2635, N2639);
nand NAND2 (N5012, N4997, N2730);
buf BUF1 (N5013, N5011);
buf BUF1 (N5014, N5003);
and AND2 (N5015, N5013, N1410);
nand NAND3 (N5016, N5012, N1009, N2287);
xor XOR2 (N5017, N5010, N3422);
nor NOR3 (N5018, N5017, N3691, N511);
or OR2 (N5019, N5015, N1057);
xor XOR2 (N5020, N5004, N4202);
not NOT1 (N5021, N5001);
nor NOR3 (N5022, N5019, N1261, N820);
nor NOR3 (N5023, N5008, N1448, N2662);
xor XOR2 (N5024, N5018, N4377);
nor NOR3 (N5025, N5009, N3604, N2895);
or OR2 (N5026, N4992, N4345);
buf BUF1 (N5027, N5020);
not NOT1 (N5028, N5026);
nand NAND4 (N5029, N5028, N2963, N2415, N710);
buf BUF1 (N5030, N5016);
not NOT1 (N5031, N5021);
xor XOR2 (N5032, N5027, N3619);
nor NOR2 (N5033, N5029, N3847);
not NOT1 (N5034, N5033);
not NOT1 (N5035, N5032);
nor NOR4 (N5036, N5030, N3640, N1928, N706);
and AND2 (N5037, N5034, N333);
nand NAND4 (N5038, N5023, N2108, N1765, N2299);
not NOT1 (N5039, N5024);
xor XOR2 (N5040, N5014, N3403);
nor NOR3 (N5041, N5005, N1884, N4490);
buf BUF1 (N5042, N5036);
or OR4 (N5043, N5035, N532, N1847, N4058);
buf BUF1 (N5044, N5043);
nor NOR2 (N5045, N5037, N3995);
and AND3 (N5046, N5025, N2580, N4375);
xor XOR2 (N5047, N5031, N3047);
xor XOR2 (N5048, N5038, N1776);
xor XOR2 (N5049, N5039, N2058);
not NOT1 (N5050, N5042);
xor XOR2 (N5051, N5050, N1063);
and AND3 (N5052, N5044, N2468, N2656);
nand NAND2 (N5053, N5048, N1779);
nor NOR3 (N5054, N5040, N2811, N2285);
or OR3 (N5055, N5052, N2020, N2285);
buf BUF1 (N5056, N5045);
nor NOR4 (N5057, N5046, N4667, N4535, N1131);
buf BUF1 (N5058, N5051);
nand NAND2 (N5059, N5056, N1616);
not NOT1 (N5060, N5022);
not NOT1 (N5061, N5053);
and AND2 (N5062, N5059, N3995);
not NOT1 (N5063, N5055);
nor NOR4 (N5064, N5041, N3791, N3344, N1918);
nor NOR3 (N5065, N5058, N1799, N2518);
not NOT1 (N5066, N5062);
and AND4 (N5067, N5060, N2576, N1571, N3087);
not NOT1 (N5068, N5067);
buf BUF1 (N5069, N5065);
buf BUF1 (N5070, N5057);
xor XOR2 (N5071, N5069, N1195);
nand NAND2 (N5072, N5068, N1816);
buf BUF1 (N5073, N5072);
xor XOR2 (N5074, N5061, N3313);
and AND4 (N5075, N5073, N3937, N2296, N907);
buf BUF1 (N5076, N5075);
buf BUF1 (N5077, N5074);
nor NOR4 (N5078, N5071, N3532, N4332, N37);
xor XOR2 (N5079, N5070, N2411);
nand NAND4 (N5080, N5076, N1723, N5026, N756);
buf BUF1 (N5081, N5079);
and AND2 (N5082, N5047, N3356);
buf BUF1 (N5083, N5049);
not NOT1 (N5084, N5054);
xor XOR2 (N5085, N5084, N1146);
not NOT1 (N5086, N5082);
and AND3 (N5087, N5086, N201, N1303);
and AND3 (N5088, N5085, N187, N882);
buf BUF1 (N5089, N5066);
nand NAND2 (N5090, N5089, N4559);
or OR2 (N5091, N5078, N4078);
nor NOR3 (N5092, N5083, N2432, N4819);
not NOT1 (N5093, N5080);
nor NOR4 (N5094, N5081, N2522, N4570, N3812);
not NOT1 (N5095, N5064);
not NOT1 (N5096, N5093);
xor XOR2 (N5097, N5094, N4500);
nor NOR4 (N5098, N5091, N2975, N3094, N636);
nor NOR3 (N5099, N5063, N3182, N4576);
and AND2 (N5100, N5095, N1302);
buf BUF1 (N5101, N5100);
nand NAND4 (N5102, N5090, N2363, N1958, N2776);
xor XOR2 (N5103, N5092, N2177);
nor NOR3 (N5104, N5101, N3279, N1383);
nand NAND2 (N5105, N5102, N584);
nor NOR4 (N5106, N5077, N4904, N3365, N207);
nand NAND3 (N5107, N5087, N315, N1948);
buf BUF1 (N5108, N5107);
or OR4 (N5109, N5098, N3541, N3187, N2651);
buf BUF1 (N5110, N5109);
not NOT1 (N5111, N5096);
nor NOR3 (N5112, N5097, N4996, N1747);
or OR2 (N5113, N5099, N5008);
not NOT1 (N5114, N5110);
nand NAND2 (N5115, N5088, N2304);
buf BUF1 (N5116, N5106);
not NOT1 (N5117, N5113);
and AND2 (N5118, N5103, N2094);
nor NOR3 (N5119, N5116, N376, N1525);
buf BUF1 (N5120, N5118);
or OR4 (N5121, N5114, N405, N2592, N647);
buf BUF1 (N5122, N5108);
or OR4 (N5123, N5122, N2862, N882, N523);
not NOT1 (N5124, N5105);
nand NAND3 (N5125, N5115, N4868, N1455);
and AND3 (N5126, N5117, N1744, N3127);
buf BUF1 (N5127, N5119);
not NOT1 (N5128, N5120);
xor XOR2 (N5129, N5126, N1);
buf BUF1 (N5130, N5127);
nand NAND2 (N5131, N5130, N3556);
xor XOR2 (N5132, N5125, N4464);
nor NOR4 (N5133, N5121, N2317, N3261, N3726);
not NOT1 (N5134, N5124);
not NOT1 (N5135, N5104);
not NOT1 (N5136, N5128);
and AND4 (N5137, N5135, N4604, N1750, N2188);
buf BUF1 (N5138, N5131);
and AND2 (N5139, N5111, N1720);
nand NAND3 (N5140, N5133, N5067, N2724);
or OR3 (N5141, N5132, N2722, N4515);
nor NOR4 (N5142, N5141, N4962, N2067, N1822);
and AND2 (N5143, N5136, N3418);
buf BUF1 (N5144, N5138);
and AND4 (N5145, N5123, N4663, N3479, N3922);
nor NOR2 (N5146, N5137, N1585);
xor XOR2 (N5147, N5144, N18);
not NOT1 (N5148, N5112);
buf BUF1 (N5149, N5148);
and AND2 (N5150, N5149, N3699);
and AND3 (N5151, N5143, N3630, N2152);
nor NOR2 (N5152, N5147, N1106);
nand NAND2 (N5153, N5142, N603);
nand NAND3 (N5154, N5129, N1920, N1390);
nand NAND3 (N5155, N5139, N2143, N1288);
buf BUF1 (N5156, N5152);
buf BUF1 (N5157, N5140);
buf BUF1 (N5158, N5156);
and AND3 (N5159, N5155, N4768, N3426);
xor XOR2 (N5160, N5157, N482);
xor XOR2 (N5161, N5150, N3128);
not NOT1 (N5162, N5134);
or OR4 (N5163, N5162, N3747, N1050, N1936);
nand NAND2 (N5164, N5161, N4437);
xor XOR2 (N5165, N5160, N2629);
nand NAND2 (N5166, N5164, N3553);
and AND4 (N5167, N5153, N3415, N2422, N2638);
nor NOR3 (N5168, N5159, N1411, N1504);
nand NAND2 (N5169, N5163, N2295);
not NOT1 (N5170, N5146);
buf BUF1 (N5171, N5145);
buf BUF1 (N5172, N5166);
or OR3 (N5173, N5169, N3509, N82);
and AND4 (N5174, N5172, N4510, N4596, N2828);
nand NAND4 (N5175, N5173, N1348, N1886, N3254);
xor XOR2 (N5176, N5175, N318);
nor NOR3 (N5177, N5158, N1490, N3854);
not NOT1 (N5178, N5151);
nand NAND4 (N5179, N5168, N4716, N554, N4083);
or OR3 (N5180, N5170, N3820, N2621);
not NOT1 (N5181, N5165);
nor NOR4 (N5182, N5174, N4007, N4547, N4549);
or OR4 (N5183, N5181, N4673, N2070, N4058);
nor NOR3 (N5184, N5182, N5087, N2090);
buf BUF1 (N5185, N5184);
or OR2 (N5186, N5178, N3036);
nand NAND4 (N5187, N5179, N4886, N465, N5145);
nor NOR2 (N5188, N5154, N2802);
nor NOR3 (N5189, N5180, N1907, N4475);
and AND2 (N5190, N5187, N4643);
and AND2 (N5191, N5177, N4043);
and AND4 (N5192, N5183, N1198, N3835, N1295);
nor NOR4 (N5193, N5192, N621, N4681, N5087);
buf BUF1 (N5194, N5189);
or OR2 (N5195, N5193, N4069);
and AND3 (N5196, N5195, N2088, N792);
or OR2 (N5197, N5186, N1611);
nor NOR3 (N5198, N5196, N2151, N3755);
xor XOR2 (N5199, N5194, N2457);
buf BUF1 (N5200, N5188);
not NOT1 (N5201, N5198);
buf BUF1 (N5202, N5199);
buf BUF1 (N5203, N5201);
not NOT1 (N5204, N5176);
not NOT1 (N5205, N5204);
xor XOR2 (N5206, N5190, N3665);
not NOT1 (N5207, N5200);
and AND4 (N5208, N5191, N2883, N4873, N2403);
not NOT1 (N5209, N5203);
nand NAND3 (N5210, N5167, N2164, N4130);
not NOT1 (N5211, N5209);
not NOT1 (N5212, N5171);
not NOT1 (N5213, N5211);
nor NOR4 (N5214, N5213, N4299, N3759, N4995);
nor NOR2 (N5215, N5185, N3748);
or OR3 (N5216, N5206, N2387, N2574);
buf BUF1 (N5217, N5214);
xor XOR2 (N5218, N5208, N4249);
or OR2 (N5219, N5217, N288);
or OR2 (N5220, N5218, N243);
or OR4 (N5221, N5207, N1470, N2912, N1211);
and AND2 (N5222, N5216, N4885);
xor XOR2 (N5223, N5219, N180);
or OR2 (N5224, N5212, N2731);
or OR3 (N5225, N5220, N4622, N1991);
or OR4 (N5226, N5222, N1515, N3966, N5125);
nand NAND3 (N5227, N5197, N1759, N3959);
nand NAND2 (N5228, N5215, N2055);
and AND3 (N5229, N5223, N3434, N3067);
or OR3 (N5230, N5221, N288, N380);
nor NOR2 (N5231, N5202, N3255);
and AND2 (N5232, N5210, N1342);
or OR3 (N5233, N5231, N4709, N2602);
and AND2 (N5234, N5229, N1673);
not NOT1 (N5235, N5232);
nand NAND3 (N5236, N5226, N3173, N4066);
nor NOR4 (N5237, N5234, N4544, N1449, N1534);
or OR2 (N5238, N5233, N474);
not NOT1 (N5239, N5205);
buf BUF1 (N5240, N5238);
nand NAND3 (N5241, N5236, N872, N1016);
or OR3 (N5242, N5227, N3995, N3081);
nand NAND4 (N5243, N5228, N1179, N1994, N2978);
not NOT1 (N5244, N5224);
nand NAND4 (N5245, N5244, N3080, N1115, N2265);
or OR3 (N5246, N5242, N4367, N3957);
buf BUF1 (N5247, N5225);
or OR4 (N5248, N5237, N3295, N3308, N1342);
buf BUF1 (N5249, N5245);
buf BUF1 (N5250, N5248);
buf BUF1 (N5251, N5239);
nor NOR4 (N5252, N5243, N296, N3820, N3050);
and AND2 (N5253, N5230, N936);
and AND4 (N5254, N5235, N2514, N4929, N2820);
nor NOR3 (N5255, N5254, N547, N2160);
and AND3 (N5256, N5246, N2930, N1537);
buf BUF1 (N5257, N5252);
and AND3 (N5258, N5256, N2171, N204);
buf BUF1 (N5259, N5255);
buf BUF1 (N5260, N5257);
and AND2 (N5261, N5249, N303);
xor XOR2 (N5262, N5260, N4711);
and AND2 (N5263, N5259, N2519);
buf BUF1 (N5264, N5263);
buf BUF1 (N5265, N5240);
or OR2 (N5266, N5265, N2013);
xor XOR2 (N5267, N5266, N2974);
nand NAND2 (N5268, N5267, N1632);
or OR4 (N5269, N5251, N630, N595, N3830);
nor NOR2 (N5270, N5268, N4761);
and AND3 (N5271, N5250, N422, N1117);
and AND2 (N5272, N5247, N2730);
not NOT1 (N5273, N5258);
nand NAND2 (N5274, N5270, N1571);
nand NAND4 (N5275, N5274, N2262, N859, N2530);
xor XOR2 (N5276, N5261, N4212);
not NOT1 (N5277, N5241);
or OR4 (N5278, N5277, N3607, N1912, N4009);
nand NAND2 (N5279, N5271, N2180);
and AND4 (N5280, N5272, N23, N544, N1804);
xor XOR2 (N5281, N5276, N4197);
xor XOR2 (N5282, N5278, N4439);
nand NAND3 (N5283, N5282, N4496, N3681);
or OR3 (N5284, N5275, N5253, N4546);
and AND3 (N5285, N3420, N3641, N2334);
xor XOR2 (N5286, N5280, N3562);
or OR3 (N5287, N5273, N2865, N4158);
buf BUF1 (N5288, N5285);
nand NAND2 (N5289, N5283, N3308);
nor NOR2 (N5290, N5262, N120);
buf BUF1 (N5291, N5284);
xor XOR2 (N5292, N5264, N342);
nand NAND4 (N5293, N5287, N3126, N5113, N4342);
and AND3 (N5294, N5293, N1156, N4434);
not NOT1 (N5295, N5294);
xor XOR2 (N5296, N5286, N3064);
not NOT1 (N5297, N5288);
and AND3 (N5298, N5269, N1635, N431);
nand NAND4 (N5299, N5295, N1437, N1189, N917);
or OR3 (N5300, N5299, N12, N886);
nand NAND4 (N5301, N5279, N2905, N2500, N3970);
not NOT1 (N5302, N5289);
and AND4 (N5303, N5296, N1108, N2646, N3364);
nor NOR2 (N5304, N5290, N3476);
buf BUF1 (N5305, N5301);
and AND3 (N5306, N5297, N5182, N3684);
nor NOR3 (N5307, N5300, N1027, N2858);
or OR2 (N5308, N5281, N1563);
xor XOR2 (N5309, N5306, N3773);
or OR2 (N5310, N5304, N4381);
and AND2 (N5311, N5303, N5090);
nor NOR3 (N5312, N5311, N1042, N539);
and AND2 (N5313, N5310, N3639);
and AND2 (N5314, N5298, N3947);
or OR4 (N5315, N5292, N2454, N5144, N3439);
or OR3 (N5316, N5314, N2709, N2431);
nand NAND4 (N5317, N5302, N480, N3646, N3908);
buf BUF1 (N5318, N5317);
not NOT1 (N5319, N5315);
nor NOR2 (N5320, N5313, N1034);
or OR4 (N5321, N5291, N259, N2859, N4537);
nor NOR3 (N5322, N5305, N4461, N4699);
not NOT1 (N5323, N5312);
and AND3 (N5324, N5309, N1966, N2753);
and AND2 (N5325, N5307, N4654);
and AND4 (N5326, N5321, N2307, N5088, N3282);
or OR4 (N5327, N5326, N4607, N2125, N4572);
xor XOR2 (N5328, N5325, N1630);
nor NOR2 (N5329, N5327, N3241);
nor NOR2 (N5330, N5319, N878);
buf BUF1 (N5331, N5320);
xor XOR2 (N5332, N5316, N2080);
buf BUF1 (N5333, N5329);
or OR3 (N5334, N5318, N4305, N705);
or OR2 (N5335, N5324, N3824);
and AND3 (N5336, N5323, N1130, N729);
xor XOR2 (N5337, N5334, N2786);
nor NOR2 (N5338, N5337, N3937);
and AND4 (N5339, N5328, N980, N3391, N1915);
nor NOR4 (N5340, N5322, N2791, N522, N4604);
not NOT1 (N5341, N5333);
nand NAND4 (N5342, N5308, N710, N3854, N196);
or OR2 (N5343, N5330, N1619);
not NOT1 (N5344, N5336);
nor NOR2 (N5345, N5344, N4118);
or OR2 (N5346, N5342, N1553);
not NOT1 (N5347, N5343);
and AND4 (N5348, N5335, N2535, N183, N3409);
or OR4 (N5349, N5339, N1882, N2552, N512);
nor NOR2 (N5350, N5332, N2335);
buf BUF1 (N5351, N5348);
xor XOR2 (N5352, N5340, N4813);
xor XOR2 (N5353, N5350, N478);
not NOT1 (N5354, N5338);
nand NAND2 (N5355, N5346, N3055);
xor XOR2 (N5356, N5352, N3914);
xor XOR2 (N5357, N5341, N4219);
or OR3 (N5358, N5331, N3893, N4484);
buf BUF1 (N5359, N5357);
and AND3 (N5360, N5358, N5102, N236);
nand NAND3 (N5361, N5349, N162, N1992);
and AND3 (N5362, N5360, N853, N3839);
xor XOR2 (N5363, N5362, N3169);
nand NAND3 (N5364, N5361, N4017, N2794);
not NOT1 (N5365, N5351);
not NOT1 (N5366, N5359);
not NOT1 (N5367, N5364);
nand NAND2 (N5368, N5363, N3507);
and AND3 (N5369, N5353, N1629, N1355);
xor XOR2 (N5370, N5367, N2682);
or OR2 (N5371, N5345, N4183);
not NOT1 (N5372, N5365);
and AND4 (N5373, N5371, N281, N833, N5143);
and AND4 (N5374, N5370, N2430, N3681, N3212);
xor XOR2 (N5375, N5369, N3902);
and AND2 (N5376, N5373, N3447);
xor XOR2 (N5377, N5347, N3123);
and AND2 (N5378, N5376, N5003);
or OR2 (N5379, N5368, N2438);
buf BUF1 (N5380, N5366);
nor NOR2 (N5381, N5354, N1662);
nand NAND3 (N5382, N5379, N722, N4672);
nor NOR3 (N5383, N5374, N2109, N3064);
nand NAND3 (N5384, N5378, N60, N3994);
buf BUF1 (N5385, N5356);
buf BUF1 (N5386, N5382);
and AND2 (N5387, N5386, N492);
xor XOR2 (N5388, N5384, N4436);
buf BUF1 (N5389, N5381);
xor XOR2 (N5390, N5372, N1870);
nand NAND2 (N5391, N5389, N3722);
not NOT1 (N5392, N5380);
or OR3 (N5393, N5383, N2877, N4349);
not NOT1 (N5394, N5393);
nor NOR2 (N5395, N5394, N5348);
and AND3 (N5396, N5387, N5019, N462);
xor XOR2 (N5397, N5390, N3081);
and AND2 (N5398, N5375, N723);
buf BUF1 (N5399, N5392);
buf BUF1 (N5400, N5397);
nor NOR4 (N5401, N5388, N1803, N1657, N4637);
or OR3 (N5402, N5396, N3110, N1400);
nor NOR3 (N5403, N5385, N3690, N289);
buf BUF1 (N5404, N5355);
and AND3 (N5405, N5391, N3849, N300);
or OR3 (N5406, N5377, N2265, N1339);
buf BUF1 (N5407, N5400);
buf BUF1 (N5408, N5399);
or OR2 (N5409, N5407, N1190);
xor XOR2 (N5410, N5395, N5406);
buf BUF1 (N5411, N39);
not NOT1 (N5412, N5409);
not NOT1 (N5413, N5412);
nand NAND2 (N5414, N5410, N2177);
or OR4 (N5415, N5398, N5053, N1642, N3144);
and AND2 (N5416, N5408, N135);
xor XOR2 (N5417, N5401, N2770);
or OR4 (N5418, N5404, N608, N39, N674);
nand NAND3 (N5419, N5413, N4263, N2905);
nor NOR2 (N5420, N5414, N2504);
nor NOR4 (N5421, N5418, N1231, N1258, N2382);
not NOT1 (N5422, N5421);
buf BUF1 (N5423, N5420);
or OR4 (N5424, N5402, N3008, N87, N3153);
not NOT1 (N5425, N5422);
buf BUF1 (N5426, N5425);
not NOT1 (N5427, N5424);
xor XOR2 (N5428, N5426, N2654);
or OR4 (N5429, N5415, N5344, N3528, N137);
or OR2 (N5430, N5427, N799);
and AND2 (N5431, N5428, N4835);
not NOT1 (N5432, N5430);
and AND2 (N5433, N5411, N2474);
nor NOR3 (N5434, N5416, N3538, N250);
xor XOR2 (N5435, N5434, N1834);
nor NOR2 (N5436, N5429, N1960);
xor XOR2 (N5437, N5417, N2605);
nand NAND3 (N5438, N5432, N2298, N802);
not NOT1 (N5439, N5431);
and AND3 (N5440, N5438, N1824, N2477);
nor NOR3 (N5441, N5423, N5332, N2153);
buf BUF1 (N5442, N5435);
nor NOR4 (N5443, N5405, N3814, N1109, N5054);
nor NOR3 (N5444, N5433, N1459, N2892);
nand NAND4 (N5445, N5441, N1416, N106, N3553);
or OR2 (N5446, N5445, N1057);
xor XOR2 (N5447, N5440, N2332);
and AND4 (N5448, N5442, N4845, N1627, N5022);
and AND2 (N5449, N5446, N4220);
or OR4 (N5450, N5419, N2748, N75, N4624);
buf BUF1 (N5451, N5449);
not NOT1 (N5452, N5444);
and AND2 (N5453, N5452, N3863);
not NOT1 (N5454, N5403);
and AND2 (N5455, N5451, N1721);
or OR2 (N5456, N5453, N3380);
not NOT1 (N5457, N5437);
nor NOR2 (N5458, N5447, N4147);
and AND4 (N5459, N5443, N4994, N2304, N2896);
not NOT1 (N5460, N5459);
nor NOR3 (N5461, N5436, N3562, N5431);
buf BUF1 (N5462, N5458);
nand NAND4 (N5463, N5461, N3470, N3180, N998);
nand NAND3 (N5464, N5456, N3615, N5361);
or OR2 (N5465, N5439, N2768);
xor XOR2 (N5466, N5465, N1674);
not NOT1 (N5467, N5450);
nor NOR3 (N5468, N5463, N772, N5453);
nand NAND3 (N5469, N5468, N3306, N224);
buf BUF1 (N5470, N5462);
not NOT1 (N5471, N5448);
not NOT1 (N5472, N5464);
buf BUF1 (N5473, N5460);
or OR3 (N5474, N5473, N257, N4205);
or OR3 (N5475, N5455, N4331, N2714);
nand NAND4 (N5476, N5470, N2115, N1995, N523);
and AND3 (N5477, N5474, N3485, N2222);
nand NAND4 (N5478, N5467, N4483, N4210, N2200);
and AND2 (N5479, N5454, N4124);
nand NAND4 (N5480, N5469, N1363, N5004, N4438);
and AND4 (N5481, N5478, N192, N4838, N3483);
or OR4 (N5482, N5471, N1803, N4822, N4590);
buf BUF1 (N5483, N5479);
nor NOR3 (N5484, N5466, N255, N669);
and AND2 (N5485, N5482, N1105);
xor XOR2 (N5486, N5484, N4718);
or OR2 (N5487, N5475, N4022);
and AND2 (N5488, N5483, N4292);
xor XOR2 (N5489, N5487, N2129);
and AND4 (N5490, N5472, N1712, N1937, N2353);
nand NAND2 (N5491, N5481, N3052);
buf BUF1 (N5492, N5486);
buf BUF1 (N5493, N5488);
buf BUF1 (N5494, N5490);
nor NOR3 (N5495, N5494, N3899, N461);
xor XOR2 (N5496, N5457, N59);
not NOT1 (N5497, N5492);
or OR3 (N5498, N5497, N2068, N4199);
and AND4 (N5499, N5493, N53, N5442, N240);
buf BUF1 (N5500, N5495);
nor NOR2 (N5501, N5480, N3563);
nand NAND2 (N5502, N5501, N3463);
not NOT1 (N5503, N5491);
nand NAND2 (N5504, N5502, N1055);
xor XOR2 (N5505, N5476, N3853);
and AND2 (N5506, N5503, N3197);
and AND4 (N5507, N5505, N2640, N111, N441);
nor NOR3 (N5508, N5507, N3335, N3720);
or OR4 (N5509, N5506, N2999, N66, N5260);
and AND4 (N5510, N5509, N2928, N2433, N404);
or OR4 (N5511, N5499, N1217, N2976, N4786);
buf BUF1 (N5512, N5477);
nand NAND3 (N5513, N5496, N1748, N2697);
not NOT1 (N5514, N5504);
nor NOR3 (N5515, N5508, N3423, N2812);
buf BUF1 (N5516, N5514);
xor XOR2 (N5517, N5511, N2070);
or OR4 (N5518, N5516, N2752, N5292, N4637);
nor NOR4 (N5519, N5510, N3516, N2530, N1894);
nor NOR3 (N5520, N5519, N4983, N919);
buf BUF1 (N5521, N5485);
buf BUF1 (N5522, N5518);
buf BUF1 (N5523, N5512);
nor NOR2 (N5524, N5489, N4613);
nor NOR3 (N5525, N5521, N5131, N1744);
and AND3 (N5526, N5500, N3831, N413);
nand NAND3 (N5527, N5513, N5276, N203);
xor XOR2 (N5528, N5523, N5445);
not NOT1 (N5529, N5524);
not NOT1 (N5530, N5528);
not NOT1 (N5531, N5517);
and AND2 (N5532, N5526, N138);
buf BUF1 (N5533, N5520);
not NOT1 (N5534, N5522);
and AND2 (N5535, N5529, N3129);
nand NAND2 (N5536, N5530, N4258);
xor XOR2 (N5537, N5534, N3267);
and AND2 (N5538, N5532, N1298);
xor XOR2 (N5539, N5533, N3446);
nand NAND4 (N5540, N5537, N4395, N484, N173);
buf BUF1 (N5541, N5531);
xor XOR2 (N5542, N5538, N267);
nand NAND3 (N5543, N5535, N5260, N106);
or OR4 (N5544, N5543, N3532, N2411, N661);
xor XOR2 (N5545, N5498, N2535);
nand NAND2 (N5546, N5527, N3467);
not NOT1 (N5547, N5541);
and AND3 (N5548, N5540, N1228, N5494);
xor XOR2 (N5549, N5548, N5454);
or OR2 (N5550, N5547, N345);
not NOT1 (N5551, N5536);
xor XOR2 (N5552, N5546, N3747);
xor XOR2 (N5553, N5552, N3685);
buf BUF1 (N5554, N5549);
nor NOR3 (N5555, N5553, N4128, N3381);
nand NAND4 (N5556, N5555, N4216, N5466, N5076);
nor NOR2 (N5557, N5545, N4975);
nand NAND3 (N5558, N5556, N4316, N4308);
xor XOR2 (N5559, N5515, N2723);
nor NOR4 (N5560, N5542, N162, N829, N1891);
nor NOR3 (N5561, N5557, N5237, N4601);
or OR2 (N5562, N5554, N1118);
not NOT1 (N5563, N5539);
not NOT1 (N5564, N5563);
and AND2 (N5565, N5550, N3390);
buf BUF1 (N5566, N5558);
or OR2 (N5567, N5564, N3406);
and AND4 (N5568, N5567, N1493, N4607, N3661);
nand NAND3 (N5569, N5544, N1263, N330);
nor NOR3 (N5570, N5562, N5367, N919);
buf BUF1 (N5571, N5561);
nor NOR2 (N5572, N5551, N4194);
buf BUF1 (N5573, N5565);
and AND3 (N5574, N5573, N3447, N1190);
buf BUF1 (N5575, N5569);
xor XOR2 (N5576, N5568, N4073);
not NOT1 (N5577, N5574);
xor XOR2 (N5578, N5560, N642);
xor XOR2 (N5579, N5559, N5404);
not NOT1 (N5580, N5571);
or OR4 (N5581, N5579, N827, N5355, N1263);
nand NAND2 (N5582, N5572, N2703);
buf BUF1 (N5583, N5570);
xor XOR2 (N5584, N5566, N4649);
not NOT1 (N5585, N5581);
or OR3 (N5586, N5577, N2870, N3819);
and AND2 (N5587, N5584, N1397);
not NOT1 (N5588, N5586);
nor NOR3 (N5589, N5587, N804, N5201);
or OR2 (N5590, N5525, N3408);
buf BUF1 (N5591, N5590);
nor NOR4 (N5592, N5585, N1917, N2286, N1645);
xor XOR2 (N5593, N5588, N1327);
not NOT1 (N5594, N5575);
and AND4 (N5595, N5594, N3132, N491, N5321);
and AND2 (N5596, N5589, N1122);
nor NOR2 (N5597, N5593, N4878);
not NOT1 (N5598, N5591);
nor NOR2 (N5599, N5582, N2671);
nor NOR4 (N5600, N5599, N4435, N2040, N1956);
xor XOR2 (N5601, N5598, N5315);
and AND2 (N5602, N5592, N2792);
and AND3 (N5603, N5595, N1453, N5123);
buf BUF1 (N5604, N5596);
buf BUF1 (N5605, N5578);
and AND3 (N5606, N5603, N972, N1441);
nand NAND4 (N5607, N5600, N1706, N4711, N5506);
nand NAND3 (N5608, N5576, N1426, N1127);
buf BUF1 (N5609, N5606);
xor XOR2 (N5610, N5607, N5056);
nand NAND2 (N5611, N5609, N431);
xor XOR2 (N5612, N5583, N2943);
or OR4 (N5613, N5608, N2756, N5490, N612);
and AND3 (N5614, N5602, N305, N847);
buf BUF1 (N5615, N5604);
nand NAND2 (N5616, N5614, N3635);
or OR2 (N5617, N5611, N719);
nand NAND4 (N5618, N5601, N2969, N2365, N4798);
or OR4 (N5619, N5605, N3357, N2155, N4073);
xor XOR2 (N5620, N5615, N4809);
and AND3 (N5621, N5620, N1064, N1638);
not NOT1 (N5622, N5612);
buf BUF1 (N5623, N5617);
buf BUF1 (N5624, N5622);
nand NAND2 (N5625, N5597, N1064);
xor XOR2 (N5626, N5610, N3155);
nor NOR3 (N5627, N5580, N249, N3418);
or OR3 (N5628, N5616, N2463, N3494);
nand NAND3 (N5629, N5625, N1432, N3066);
not NOT1 (N5630, N5626);
nand NAND2 (N5631, N5630, N5194);
buf BUF1 (N5632, N5623);
and AND4 (N5633, N5613, N2438, N1511, N2695);
xor XOR2 (N5634, N5629, N3354);
buf BUF1 (N5635, N5627);
xor XOR2 (N5636, N5631, N5072);
or OR3 (N5637, N5635, N1712, N4470);
and AND3 (N5638, N5628, N5239, N734);
xor XOR2 (N5639, N5638, N5521);
xor XOR2 (N5640, N5633, N1622);
not NOT1 (N5641, N5624);
nand NAND3 (N5642, N5641, N2804, N841);
and AND2 (N5643, N5632, N1978);
nand NAND2 (N5644, N5639, N1136);
or OR2 (N5645, N5642, N4036);
not NOT1 (N5646, N5618);
xor XOR2 (N5647, N5636, N5140);
buf BUF1 (N5648, N5619);
nor NOR3 (N5649, N5637, N4385, N1840);
and AND3 (N5650, N5634, N4984, N1089);
and AND4 (N5651, N5645, N3707, N1227, N1376);
or OR2 (N5652, N5640, N1529);
nand NAND2 (N5653, N5646, N3638);
nand NAND4 (N5654, N5651, N4717, N4328, N3783);
not NOT1 (N5655, N5647);
buf BUF1 (N5656, N5644);
or OR3 (N5657, N5652, N1116, N958);
not NOT1 (N5658, N5656);
nor NOR2 (N5659, N5643, N255);
not NOT1 (N5660, N5659);
nor NOR2 (N5661, N5649, N1154);
xor XOR2 (N5662, N5650, N5392);
or OR3 (N5663, N5655, N3766, N4095);
buf BUF1 (N5664, N5663);
nor NOR4 (N5665, N5664, N4884, N4805, N2416);
and AND3 (N5666, N5653, N2759, N5063);
buf BUF1 (N5667, N5660);
and AND4 (N5668, N5665, N4824, N5455, N535);
buf BUF1 (N5669, N5648);
and AND3 (N5670, N5661, N3217, N2273);
nor NOR3 (N5671, N5654, N1810, N5329);
or OR3 (N5672, N5621, N1187, N2697);
xor XOR2 (N5673, N5662, N138);
xor XOR2 (N5674, N5667, N4493);
nor NOR2 (N5675, N5666, N4765);
nand NAND3 (N5676, N5657, N1482, N2723);
nor NOR3 (N5677, N5673, N3365, N495);
or OR2 (N5678, N5668, N412);
and AND3 (N5679, N5658, N2025, N1490);
and AND4 (N5680, N5672, N68, N1662, N4223);
or OR4 (N5681, N5671, N4552, N2562, N4734);
xor XOR2 (N5682, N5669, N3416);
or OR2 (N5683, N5680, N2915);
buf BUF1 (N5684, N5677);
xor XOR2 (N5685, N5670, N4580);
or OR3 (N5686, N5682, N4426, N3594);
xor XOR2 (N5687, N5681, N4898);
xor XOR2 (N5688, N5675, N3950);
buf BUF1 (N5689, N5684);
buf BUF1 (N5690, N5679);
xor XOR2 (N5691, N5687, N2557);
or OR3 (N5692, N5690, N2774, N1122);
nand NAND3 (N5693, N5689, N919, N2758);
nor NOR2 (N5694, N5686, N1128);
or OR2 (N5695, N5674, N3629);
or OR3 (N5696, N5693, N1661, N1636);
nand NAND2 (N5697, N5685, N5594);
or OR2 (N5698, N5696, N2213);
nor NOR4 (N5699, N5688, N2869, N2759, N3904);
or OR2 (N5700, N5678, N4743);
xor XOR2 (N5701, N5695, N4290);
and AND3 (N5702, N5699, N4885, N1713);
and AND3 (N5703, N5698, N782, N3431);
nor NOR2 (N5704, N5676, N4575);
xor XOR2 (N5705, N5704, N5168);
and AND2 (N5706, N5692, N401);
and AND4 (N5707, N5701, N4480, N765, N2083);
and AND2 (N5708, N5691, N2696);
nor NOR2 (N5709, N5705, N5467);
not NOT1 (N5710, N5703);
nand NAND3 (N5711, N5709, N74, N60);
not NOT1 (N5712, N5697);
nand NAND4 (N5713, N5706, N4425, N2270, N442);
nand NAND2 (N5714, N5707, N1930);
not NOT1 (N5715, N5710);
nor NOR2 (N5716, N5702, N2715);
and AND4 (N5717, N5700, N2721, N20, N2183);
or OR2 (N5718, N5717, N2314);
buf BUF1 (N5719, N5715);
buf BUF1 (N5720, N5718);
not NOT1 (N5721, N5714);
and AND2 (N5722, N5720, N2550);
nand NAND4 (N5723, N5722, N4762, N352, N1943);
xor XOR2 (N5724, N5694, N3572);
buf BUF1 (N5725, N5716);
nand NAND3 (N5726, N5713, N59, N5337);
buf BUF1 (N5727, N5721);
nand NAND3 (N5728, N5725, N2269, N5052);
and AND2 (N5729, N5711, N3338);
xor XOR2 (N5730, N5708, N3371);
not NOT1 (N5731, N5719);
not NOT1 (N5732, N5727);
xor XOR2 (N5733, N5732, N352);
buf BUF1 (N5734, N5728);
and AND2 (N5735, N5729, N5536);
not NOT1 (N5736, N5683);
nand NAND2 (N5737, N5712, N1349);
xor XOR2 (N5738, N5724, N2936);
nor NOR2 (N5739, N5730, N5313);
buf BUF1 (N5740, N5731);
buf BUF1 (N5741, N5726);
and AND2 (N5742, N5736, N3258);
nor NOR4 (N5743, N5737, N5181, N4488, N3236);
nand NAND2 (N5744, N5742, N4275);
and AND3 (N5745, N5735, N168, N5733);
nor NOR4 (N5746, N2756, N232, N2219, N392);
xor XOR2 (N5747, N5738, N1669);
nor NOR2 (N5748, N5743, N2281);
nor NOR2 (N5749, N5746, N3041);
nor NOR2 (N5750, N5741, N3864);
and AND2 (N5751, N5734, N5027);
xor XOR2 (N5752, N5739, N4554);
and AND2 (N5753, N5747, N5299);
or OR3 (N5754, N5752, N2899, N801);
and AND3 (N5755, N5750, N3369, N2574);
nand NAND3 (N5756, N5745, N2598, N5642);
xor XOR2 (N5757, N5753, N4608);
not NOT1 (N5758, N5723);
and AND2 (N5759, N5755, N1503);
not NOT1 (N5760, N5749);
and AND4 (N5761, N5744, N2752, N5727, N2853);
or OR3 (N5762, N5751, N1430, N5418);
nand NAND3 (N5763, N5761, N4072, N5759);
buf BUF1 (N5764, N3256);
nor NOR3 (N5765, N5748, N3101, N5690);
nor NOR4 (N5766, N5754, N2334, N2005, N5472);
and AND2 (N5767, N5763, N337);
nand NAND4 (N5768, N5764, N3779, N2738, N3490);
or OR3 (N5769, N5766, N3949, N5541);
nor NOR4 (N5770, N5757, N1696, N5528, N3336);
buf BUF1 (N5771, N5760);
nor NOR3 (N5772, N5765, N3915, N481);
not NOT1 (N5773, N5756);
and AND3 (N5774, N5771, N945, N36);
not NOT1 (N5775, N5758);
or OR2 (N5776, N5772, N3607);
buf BUF1 (N5777, N5740);
not NOT1 (N5778, N5770);
and AND4 (N5779, N5767, N577, N1920, N2567);
xor XOR2 (N5780, N5779, N2053);
nand NAND4 (N5781, N5768, N4533, N5686, N1203);
or OR3 (N5782, N5780, N5033, N349);
and AND2 (N5783, N5777, N1981);
nand NAND4 (N5784, N5776, N3582, N1436, N2421);
buf BUF1 (N5785, N5781);
not NOT1 (N5786, N5775);
and AND4 (N5787, N5769, N2065, N2985, N234);
and AND3 (N5788, N5783, N2347, N1778);
nand NAND4 (N5789, N5787, N2305, N2117, N4737);
not NOT1 (N5790, N5788);
or OR3 (N5791, N5778, N2780, N650);
nand NAND2 (N5792, N5762, N2243);
or OR3 (N5793, N5782, N3678, N3478);
nand NAND3 (N5794, N5789, N3187, N2755);
or OR2 (N5795, N5793, N1092);
nand NAND2 (N5796, N5794, N2560);
nor NOR4 (N5797, N5795, N3670, N4907, N2812);
nor NOR4 (N5798, N5773, N5796, N5683, N5168);
not NOT1 (N5799, N4002);
not NOT1 (N5800, N5785);
and AND2 (N5801, N5797, N1051);
or OR2 (N5802, N5786, N3924);
buf BUF1 (N5803, N5802);
nor NOR4 (N5804, N5798, N3916, N3221, N4986);
and AND2 (N5805, N5774, N141);
or OR3 (N5806, N5799, N3801, N603);
and AND3 (N5807, N5800, N1755, N1430);
buf BUF1 (N5808, N5801);
xor XOR2 (N5809, N5804, N3321);
buf BUF1 (N5810, N5784);
buf BUF1 (N5811, N5806);
or OR4 (N5812, N5790, N4186, N3947, N3871);
not NOT1 (N5813, N5811);
nor NOR2 (N5814, N5810, N4265);
or OR4 (N5815, N5805, N1366, N2739, N99);
or OR3 (N5816, N5807, N168, N2718);
not NOT1 (N5817, N5816);
not NOT1 (N5818, N5792);
buf BUF1 (N5819, N5815);
nor NOR2 (N5820, N5803, N4410);
or OR3 (N5821, N5819, N1494, N3166);
and AND4 (N5822, N5812, N4195, N700, N1497);
or OR4 (N5823, N5821, N319, N3303, N5157);
xor XOR2 (N5824, N5791, N1575);
nor NOR4 (N5825, N5813, N1836, N2931, N3179);
and AND4 (N5826, N5814, N2080, N3740, N3059);
nor NOR3 (N5827, N5826, N403, N2118);
not NOT1 (N5828, N5825);
not NOT1 (N5829, N5828);
xor XOR2 (N5830, N5822, N3876);
xor XOR2 (N5831, N5829, N3705);
not NOT1 (N5832, N5818);
xor XOR2 (N5833, N5827, N4827);
buf BUF1 (N5834, N5820);
and AND3 (N5835, N5809, N2573, N1019);
and AND3 (N5836, N5834, N3598, N4183);
or OR4 (N5837, N5830, N2005, N582, N1400);
buf BUF1 (N5838, N5836);
and AND3 (N5839, N5808, N1488, N2802);
buf BUF1 (N5840, N5831);
and AND2 (N5841, N5837, N3730);
xor XOR2 (N5842, N5832, N1772);
nand NAND3 (N5843, N5839, N2857, N2772);
or OR3 (N5844, N5835, N291, N3868);
nand NAND3 (N5845, N5843, N2883, N2109);
xor XOR2 (N5846, N5838, N1226);
not NOT1 (N5847, N5845);
and AND3 (N5848, N5824, N1163, N4344);
xor XOR2 (N5849, N5841, N2725);
not NOT1 (N5850, N5840);
buf BUF1 (N5851, N5842);
or OR2 (N5852, N5844, N5410);
not NOT1 (N5853, N5833);
xor XOR2 (N5854, N5817, N1465);
nor NOR3 (N5855, N5823, N4557, N2784);
nor NOR3 (N5856, N5853, N415, N5248);
xor XOR2 (N5857, N5856, N1758);
buf BUF1 (N5858, N5854);
xor XOR2 (N5859, N5851, N1512);
buf BUF1 (N5860, N5859);
and AND4 (N5861, N5855, N2362, N240, N4801);
nand NAND2 (N5862, N5847, N2618);
not NOT1 (N5863, N5849);
buf BUF1 (N5864, N5850);
nand NAND4 (N5865, N5857, N4323, N2480, N5396);
not NOT1 (N5866, N5862);
xor XOR2 (N5867, N5846, N4452);
not NOT1 (N5868, N5866);
not NOT1 (N5869, N5863);
and AND2 (N5870, N5864, N374);
buf BUF1 (N5871, N5860);
nor NOR4 (N5872, N5871, N3133, N1881, N1273);
and AND2 (N5873, N5872, N2061);
and AND4 (N5874, N5858, N1672, N3738, N2762);
or OR2 (N5875, N5861, N732);
buf BUF1 (N5876, N5865);
buf BUF1 (N5877, N5876);
buf BUF1 (N5878, N5875);
nand NAND3 (N5879, N5869, N5086, N4685);
nor NOR3 (N5880, N5870, N5664, N445);
nand NAND2 (N5881, N5867, N5860);
or OR2 (N5882, N5879, N4832);
not NOT1 (N5883, N5874);
nand NAND4 (N5884, N5878, N2134, N2620, N2223);
or OR2 (N5885, N5880, N5168);
and AND4 (N5886, N5852, N370, N5502, N3224);
or OR3 (N5887, N5868, N2506, N3077);
or OR4 (N5888, N5877, N2495, N2854, N2220);
and AND2 (N5889, N5888, N4649);
or OR2 (N5890, N5885, N46);
nor NOR3 (N5891, N5873, N1321, N3156);
and AND4 (N5892, N5886, N2740, N5558, N3872);
buf BUF1 (N5893, N5884);
or OR2 (N5894, N5881, N4139);
nor NOR4 (N5895, N5894, N4232, N5000, N3435);
nand NAND2 (N5896, N5883, N1442);
and AND3 (N5897, N5889, N3655, N3992);
xor XOR2 (N5898, N5891, N4341);
nor NOR2 (N5899, N5882, N3230);
nand NAND3 (N5900, N5892, N168, N4657);
not NOT1 (N5901, N5848);
xor XOR2 (N5902, N5897, N4290);
and AND4 (N5903, N5890, N1274, N3329, N2353);
nand NAND4 (N5904, N5895, N2164, N2590, N3504);
nand NAND2 (N5905, N5899, N1219);
nor NOR4 (N5906, N5903, N1231, N5350, N1098);
buf BUF1 (N5907, N5904);
nor NOR3 (N5908, N5906, N2246, N1258);
xor XOR2 (N5909, N5900, N1937);
nand NAND2 (N5910, N5902, N1252);
not NOT1 (N5911, N5905);
or OR3 (N5912, N5896, N1845, N917);
not NOT1 (N5913, N5911);
xor XOR2 (N5914, N5912, N3454);
nand NAND3 (N5915, N5907, N221, N4712);
not NOT1 (N5916, N5908);
buf BUF1 (N5917, N5887);
nor NOR3 (N5918, N5909, N6, N572);
buf BUF1 (N5919, N5914);
xor XOR2 (N5920, N5913, N3553);
xor XOR2 (N5921, N5917, N1531);
nand NAND3 (N5922, N5898, N3693, N5390);
not NOT1 (N5923, N5920);
nor NOR3 (N5924, N5919, N3615, N1605);
not NOT1 (N5925, N5901);
not NOT1 (N5926, N5916);
xor XOR2 (N5927, N5923, N3425);
nor NOR2 (N5928, N5915, N2615);
nor NOR3 (N5929, N5926, N3486, N2564);
not NOT1 (N5930, N5893);
xor XOR2 (N5931, N5925, N4945);
buf BUF1 (N5932, N5910);
and AND4 (N5933, N5927, N2416, N3583, N5031);
nor NOR3 (N5934, N5933, N78, N4452);
and AND3 (N5935, N5929, N2968, N948);
and AND3 (N5936, N5921, N203, N2299);
or OR4 (N5937, N5934, N2208, N242, N5486);
or OR3 (N5938, N5937, N4354, N1697);
or OR4 (N5939, N5935, N5764, N3792, N1190);
nor NOR3 (N5940, N5928, N4279, N3937);
and AND3 (N5941, N5930, N1166, N5921);
xor XOR2 (N5942, N5938, N3057);
and AND2 (N5943, N5918, N3387);
or OR2 (N5944, N5931, N1571);
nor NOR3 (N5945, N5936, N3281, N3723);
xor XOR2 (N5946, N5939, N4171);
nor NOR2 (N5947, N5944, N5792);
nand NAND3 (N5948, N5943, N3310, N2443);
nand NAND3 (N5949, N5922, N1803, N5769);
buf BUF1 (N5950, N5941);
nand NAND4 (N5951, N5932, N2529, N432, N3914);
xor XOR2 (N5952, N5940, N3708);
and AND4 (N5953, N5949, N3119, N5886, N1136);
buf BUF1 (N5954, N5942);
nor NOR2 (N5955, N5953, N1079);
not NOT1 (N5956, N5954);
not NOT1 (N5957, N5924);
nor NOR4 (N5958, N5947, N2643, N2854, N4785);
nand NAND2 (N5959, N5951, N2270);
not NOT1 (N5960, N5957);
xor XOR2 (N5961, N5959, N205);
nor NOR4 (N5962, N5945, N1181, N2132, N539);
nand NAND2 (N5963, N5956, N3195);
buf BUF1 (N5964, N5962);
not NOT1 (N5965, N5948);
buf BUF1 (N5966, N5952);
or OR3 (N5967, N5955, N5446, N4983);
not NOT1 (N5968, N5946);
nor NOR3 (N5969, N5965, N4330, N335);
nor NOR4 (N5970, N5961, N2477, N1596, N3544);
and AND4 (N5971, N5964, N3040, N2728, N4128);
not NOT1 (N5972, N5966);
or OR3 (N5973, N5971, N2185, N2403);
xor XOR2 (N5974, N5950, N3849);
or OR4 (N5975, N5970, N3117, N2392, N2855);
and AND3 (N5976, N5967, N4907, N3083);
and AND3 (N5977, N5972, N1385, N2371);
not NOT1 (N5978, N5973);
xor XOR2 (N5979, N5958, N4259);
nand NAND4 (N5980, N5963, N3776, N1353, N5029);
buf BUF1 (N5981, N5975);
nand NAND2 (N5982, N5977, N1193);
xor XOR2 (N5983, N5978, N2239);
or OR4 (N5984, N5968, N3356, N3532, N4151);
not NOT1 (N5985, N5969);
and AND3 (N5986, N5983, N2321, N2752);
or OR3 (N5987, N5985, N1654, N1066);
nor NOR3 (N5988, N5981, N4871, N5982);
and AND4 (N5989, N1976, N2971, N1131, N5776);
and AND2 (N5990, N5987, N5256);
buf BUF1 (N5991, N5984);
not NOT1 (N5992, N5989);
or OR2 (N5993, N5990, N2306);
or OR4 (N5994, N5979, N10, N1413, N590);
buf BUF1 (N5995, N5991);
or OR4 (N5996, N5995, N783, N5052, N4042);
and AND4 (N5997, N5974, N895, N1879, N2042);
or OR2 (N5998, N5994, N5967);
or OR2 (N5999, N5980, N1933);
xor XOR2 (N6000, N5997, N5261);
nor NOR4 (N6001, N5976, N4724, N4441, N5869);
and AND2 (N6002, N5999, N3240);
xor XOR2 (N6003, N6000, N4805);
nand NAND2 (N6004, N5998, N914);
xor XOR2 (N6005, N5986, N1468);
buf BUF1 (N6006, N6001);
or OR3 (N6007, N5960, N430, N4008);
buf BUF1 (N6008, N6007);
or OR4 (N6009, N5996, N4007, N375, N5288);
buf BUF1 (N6010, N5988);
xor XOR2 (N6011, N6003, N3472);
and AND4 (N6012, N6004, N306, N2656, N3046);
not NOT1 (N6013, N5992);
nand NAND4 (N6014, N6012, N3362, N4630, N4176);
or OR4 (N6015, N6008, N4421, N3214, N5565);
not NOT1 (N6016, N6009);
and AND3 (N6017, N6002, N5608, N602);
not NOT1 (N6018, N6011);
and AND2 (N6019, N6006, N4757);
nand NAND3 (N6020, N6005, N418, N3932);
nor NOR4 (N6021, N6015, N1052, N3820, N3071);
nor NOR2 (N6022, N6017, N5946);
not NOT1 (N6023, N6019);
or OR4 (N6024, N6014, N2373, N690, N1217);
and AND4 (N6025, N6021, N5485, N784, N891);
and AND4 (N6026, N6024, N2116, N3306, N1079);
not NOT1 (N6027, N6018);
xor XOR2 (N6028, N6016, N3671);
nor NOR2 (N6029, N6025, N294);
nor NOR4 (N6030, N5993, N6016, N18, N868);
or OR3 (N6031, N6029, N4922, N922);
nand NAND3 (N6032, N6028, N2074, N2067);
not NOT1 (N6033, N6026);
nor NOR4 (N6034, N6032, N5017, N4814, N5316);
xor XOR2 (N6035, N6027, N1605);
nand NAND3 (N6036, N6031, N2373, N3150);
or OR4 (N6037, N6036, N4350, N288, N380);
or OR2 (N6038, N6035, N1517);
and AND2 (N6039, N6034, N1504);
not NOT1 (N6040, N6022);
or OR3 (N6041, N6023, N4825, N1671);
and AND2 (N6042, N6041, N4843);
nor NOR4 (N6043, N6010, N559, N5756, N4117);
or OR4 (N6044, N6020, N3809, N2716, N2823);
xor XOR2 (N6045, N6033, N3525);
buf BUF1 (N6046, N6042);
xor XOR2 (N6047, N6038, N5537);
xor XOR2 (N6048, N6046, N4171);
nand NAND2 (N6049, N6047, N1657);
buf BUF1 (N6050, N6037);
not NOT1 (N6051, N6045);
buf BUF1 (N6052, N6048);
or OR4 (N6053, N6050, N2666, N1946, N233);
and AND3 (N6054, N6043, N3378, N4584);
not NOT1 (N6055, N6052);
buf BUF1 (N6056, N6039);
nor NOR2 (N6057, N6054, N5749);
or OR3 (N6058, N6053, N871, N2078);
nor NOR4 (N6059, N6057, N3950, N580, N3469);
xor XOR2 (N6060, N6049, N3970);
and AND3 (N6061, N6060, N5862, N1219);
or OR4 (N6062, N6061, N6058, N6010, N1262);
buf BUF1 (N6063, N5804);
not NOT1 (N6064, N6063);
or OR2 (N6065, N6062, N1347);
or OR4 (N6066, N6030, N55, N207, N265);
nor NOR4 (N6067, N6044, N4458, N4277, N5835);
or OR2 (N6068, N6055, N2957);
buf BUF1 (N6069, N6040);
not NOT1 (N6070, N6065);
or OR2 (N6071, N6013, N3483);
nor NOR4 (N6072, N6051, N5189, N2523, N4852);
or OR2 (N6073, N6066, N1918);
or OR2 (N6074, N6067, N1653);
xor XOR2 (N6075, N6068, N3277);
or OR4 (N6076, N6064, N5352, N2969, N4037);
and AND2 (N6077, N6070, N253);
buf BUF1 (N6078, N6076);
or OR4 (N6079, N6077, N5206, N5874, N2357);
xor XOR2 (N6080, N6078, N1612);
and AND3 (N6081, N6059, N2978, N5787);
buf BUF1 (N6082, N6073);
nand NAND4 (N6083, N6080, N10, N119, N5184);
nor NOR2 (N6084, N6079, N1428);
buf BUF1 (N6085, N6084);
or OR2 (N6086, N6083, N5384);
or OR4 (N6087, N6056, N1466, N2965, N3469);
xor XOR2 (N6088, N6081, N1570);
or OR3 (N6089, N6072, N3851, N5877);
nand NAND3 (N6090, N6086, N2, N2374);
or OR4 (N6091, N6075, N5400, N1744, N1622);
and AND2 (N6092, N6090, N5401);
and AND4 (N6093, N6089, N4881, N4323, N4190);
not NOT1 (N6094, N6088);
xor XOR2 (N6095, N6071, N4806);
buf BUF1 (N6096, N6091);
and AND3 (N6097, N6069, N1528, N4763);
nand NAND3 (N6098, N6094, N1873, N1359);
xor XOR2 (N6099, N6085, N2801);
xor XOR2 (N6100, N6099, N3961);
or OR3 (N6101, N6074, N3990, N3155);
xor XOR2 (N6102, N6092, N5751);
xor XOR2 (N6103, N6102, N1631);
or OR2 (N6104, N6082, N723);
or OR3 (N6105, N6087, N5472, N624);
nor NOR4 (N6106, N6103, N4056, N1574, N4815);
nand NAND3 (N6107, N6093, N4360, N4972);
or OR3 (N6108, N6107, N4473, N4140);
not NOT1 (N6109, N6104);
xor XOR2 (N6110, N6106, N2027);
nor NOR4 (N6111, N6110, N528, N4295, N4446);
nand NAND3 (N6112, N6111, N4325, N604);
and AND2 (N6113, N6100, N2151);
and AND3 (N6114, N6113, N1999, N4357);
xor XOR2 (N6115, N6096, N723);
not NOT1 (N6116, N6105);
buf BUF1 (N6117, N6115);
or OR4 (N6118, N6097, N3097, N2414, N407);
nor NOR3 (N6119, N6101, N5543, N534);
and AND3 (N6120, N6108, N5678, N2399);
nand NAND2 (N6121, N6120, N5998);
not NOT1 (N6122, N6116);
not NOT1 (N6123, N6112);
and AND4 (N6124, N6098, N5756, N929, N119);
xor XOR2 (N6125, N6123, N1071);
nor NOR4 (N6126, N6095, N1050, N4282, N2627);
and AND2 (N6127, N6126, N743);
not NOT1 (N6128, N6114);
or OR4 (N6129, N6128, N2458, N4974, N1591);
buf BUF1 (N6130, N6129);
or OR2 (N6131, N6117, N3790);
and AND3 (N6132, N6109, N4115, N5576);
nand NAND4 (N6133, N6125, N5221, N5295, N3164);
not NOT1 (N6134, N6124);
nor NOR3 (N6135, N6132, N5901, N494);
buf BUF1 (N6136, N6131);
nor NOR3 (N6137, N6133, N1309, N136);
nand NAND3 (N6138, N6130, N3278, N497);
or OR3 (N6139, N6135, N1846, N973);
nor NOR3 (N6140, N6137, N3680, N3725);
nand NAND4 (N6141, N6140, N2478, N3568, N489);
or OR4 (N6142, N6118, N2378, N4624, N1522);
xor XOR2 (N6143, N6119, N578);
xor XOR2 (N6144, N6141, N3941);
xor XOR2 (N6145, N6122, N3535);
not NOT1 (N6146, N6138);
nor NOR3 (N6147, N6127, N5327, N206);
and AND2 (N6148, N6145, N4199);
nor NOR3 (N6149, N6148, N2497, N5206);
xor XOR2 (N6150, N6146, N2535);
and AND4 (N6151, N6139, N4799, N1604, N5175);
buf BUF1 (N6152, N6143);
and AND3 (N6153, N6150, N3131, N3060);
buf BUF1 (N6154, N6121);
not NOT1 (N6155, N6142);
buf BUF1 (N6156, N6153);
nand NAND4 (N6157, N6154, N1215, N2092, N3432);
nand NAND2 (N6158, N6156, N3013);
xor XOR2 (N6159, N6144, N538);
nor NOR3 (N6160, N6155, N3213, N524);
or OR4 (N6161, N6151, N3763, N5885, N2573);
not NOT1 (N6162, N6136);
nor NOR4 (N6163, N6152, N3635, N4206, N5920);
xor XOR2 (N6164, N6163, N5625);
nor NOR4 (N6165, N6147, N113, N3273, N5187);
and AND2 (N6166, N6158, N4333);
buf BUF1 (N6167, N6149);
buf BUF1 (N6168, N6134);
nand NAND3 (N6169, N6168, N1955, N4022);
and AND4 (N6170, N6169, N2733, N2950, N2639);
and AND3 (N6171, N6161, N5505, N4517);
not NOT1 (N6172, N6162);
nand NAND2 (N6173, N6160, N673);
nor NOR2 (N6174, N6171, N4906);
nand NAND4 (N6175, N6172, N3052, N2700, N388);
buf BUF1 (N6176, N6174);
and AND3 (N6177, N6176, N984, N3710);
or OR4 (N6178, N6165, N4395, N2184, N203);
or OR2 (N6179, N6177, N477);
and AND4 (N6180, N6159, N3450, N100, N6046);
not NOT1 (N6181, N6179);
xor XOR2 (N6182, N6181, N4624);
or OR2 (N6183, N6164, N5523);
nand NAND2 (N6184, N6166, N5917);
buf BUF1 (N6185, N6182);
nand NAND3 (N6186, N6170, N1108, N1889);
buf BUF1 (N6187, N6184);
buf BUF1 (N6188, N6185);
nor NOR2 (N6189, N6157, N4967);
nor NOR2 (N6190, N6186, N178);
nor NOR4 (N6191, N6190, N349, N643, N5278);
buf BUF1 (N6192, N6188);
nor NOR2 (N6193, N6187, N4280);
buf BUF1 (N6194, N6183);
nand NAND2 (N6195, N6175, N4394);
or OR3 (N6196, N6193, N4095, N6129);
nor NOR3 (N6197, N6194, N4301, N5292);
nor NOR4 (N6198, N6167, N3237, N5694, N5140);
nor NOR3 (N6199, N6173, N5339, N291);
not NOT1 (N6200, N6192);
nor NOR4 (N6201, N6189, N6086, N102, N3734);
xor XOR2 (N6202, N6200, N1238);
buf BUF1 (N6203, N6178);
and AND3 (N6204, N6180, N964, N110);
buf BUF1 (N6205, N6197);
buf BUF1 (N6206, N6199);
xor XOR2 (N6207, N6202, N1371);
or OR4 (N6208, N6205, N2733, N1982, N670);
nand NAND2 (N6209, N6207, N1146);
buf BUF1 (N6210, N6208);
nand NAND3 (N6211, N6195, N2734, N2840);
xor XOR2 (N6212, N6206, N5198);
buf BUF1 (N6213, N6211);
and AND2 (N6214, N6196, N4821);
nand NAND3 (N6215, N6198, N726, N3963);
nand NAND2 (N6216, N6213, N4875);
buf BUF1 (N6217, N6216);
xor XOR2 (N6218, N6215, N1031);
buf BUF1 (N6219, N6191);
buf BUF1 (N6220, N6217);
nor NOR2 (N6221, N6204, N228);
or OR2 (N6222, N6221, N1249);
nor NOR2 (N6223, N6203, N2253);
nor NOR3 (N6224, N6212, N1615, N3320);
nand NAND4 (N6225, N6220, N685, N4933, N578);
xor XOR2 (N6226, N6218, N1097);
and AND2 (N6227, N6223, N5618);
xor XOR2 (N6228, N6219, N1698);
and AND2 (N6229, N6227, N2028);
nor NOR4 (N6230, N6201, N219, N5233, N4025);
xor XOR2 (N6231, N6225, N4124);
not NOT1 (N6232, N6210);
nand NAND3 (N6233, N6226, N2974, N2942);
or OR3 (N6234, N6230, N2959, N1831);
or OR3 (N6235, N6231, N5690, N4962);
xor XOR2 (N6236, N6234, N18);
and AND4 (N6237, N6214, N1789, N1813, N1259);
nand NAND4 (N6238, N6237, N276, N2468, N2771);
not NOT1 (N6239, N6238);
not NOT1 (N6240, N6229);
or OR3 (N6241, N6235, N6177, N5819);
buf BUF1 (N6242, N6239);
not NOT1 (N6243, N6209);
xor XOR2 (N6244, N6233, N1500);
nand NAND3 (N6245, N6232, N1616, N1940);
buf BUF1 (N6246, N6243);
buf BUF1 (N6247, N6246);
or OR2 (N6248, N6236, N1295);
buf BUF1 (N6249, N6241);
and AND4 (N6250, N6240, N2055, N4115, N276);
nor NOR2 (N6251, N6249, N4895);
buf BUF1 (N6252, N6248);
xor XOR2 (N6253, N6224, N4907);
and AND3 (N6254, N6247, N2659, N1391);
nand NAND3 (N6255, N6228, N1635, N4469);
and AND3 (N6256, N6245, N4437, N101);
nor NOR2 (N6257, N6252, N5392);
and AND2 (N6258, N6253, N5629);
not NOT1 (N6259, N6257);
and AND2 (N6260, N6222, N2971);
not NOT1 (N6261, N6251);
nor NOR4 (N6262, N6254, N788, N5606, N4883);
or OR4 (N6263, N6260, N2648, N3376, N2026);
or OR3 (N6264, N6242, N5866, N3643);
not NOT1 (N6265, N6258);
xor XOR2 (N6266, N6255, N1135);
not NOT1 (N6267, N6259);
not NOT1 (N6268, N6263);
or OR2 (N6269, N6266, N3903);
and AND2 (N6270, N6265, N4726);
and AND3 (N6271, N6250, N682, N974);
nor NOR3 (N6272, N6267, N5326, N2428);
not NOT1 (N6273, N6272);
buf BUF1 (N6274, N6261);
or OR2 (N6275, N6256, N2126);
buf BUF1 (N6276, N6262);
and AND4 (N6277, N6268, N3024, N3491, N4009);
xor XOR2 (N6278, N6244, N4938);
xor XOR2 (N6279, N6269, N5517);
nor NOR4 (N6280, N6277, N549, N5347, N4472);
xor XOR2 (N6281, N6276, N550);
and AND4 (N6282, N6273, N5984, N1462, N3627);
or OR2 (N6283, N6275, N6058);
buf BUF1 (N6284, N6278);
buf BUF1 (N6285, N6282);
and AND4 (N6286, N6285, N1195, N5341, N2051);
nor NOR4 (N6287, N6264, N3835, N91, N3966);
not NOT1 (N6288, N6287);
not NOT1 (N6289, N6288);
and AND3 (N6290, N6284, N3694, N3710);
buf BUF1 (N6291, N6283);
buf BUF1 (N6292, N6270);
not NOT1 (N6293, N6291);
nand NAND3 (N6294, N6271, N4952, N1022);
nand NAND2 (N6295, N6293, N1175);
buf BUF1 (N6296, N6281);
nor NOR3 (N6297, N6292, N6094, N2354);
nand NAND3 (N6298, N6280, N4162, N1134);
nor NOR4 (N6299, N6286, N1075, N844, N5922);
or OR2 (N6300, N6299, N3404);
or OR4 (N6301, N6300, N3695, N4391, N3317);
not NOT1 (N6302, N6298);
xor XOR2 (N6303, N6274, N1534);
not NOT1 (N6304, N6296);
nor NOR3 (N6305, N6290, N3056, N262);
nand NAND4 (N6306, N6303, N4709, N1654, N3237);
nand NAND3 (N6307, N6302, N4122, N6180);
nand NAND4 (N6308, N6294, N4365, N1930, N815);
and AND2 (N6309, N6306, N4211);
not NOT1 (N6310, N6279);
and AND3 (N6311, N6305, N2681, N2683);
nor NOR4 (N6312, N6304, N3199, N3666, N5178);
buf BUF1 (N6313, N6289);
or OR4 (N6314, N6307, N3088, N2594, N563);
not NOT1 (N6315, N6311);
and AND2 (N6316, N6313, N434);
and AND2 (N6317, N6316, N4647);
or OR2 (N6318, N6317, N4147);
buf BUF1 (N6319, N6310);
or OR4 (N6320, N6319, N5303, N1534, N4194);
not NOT1 (N6321, N6308);
and AND3 (N6322, N6297, N318, N5278);
nand NAND2 (N6323, N6320, N4849);
buf BUF1 (N6324, N6309);
and AND4 (N6325, N6312, N5684, N1271, N3071);
nand NAND3 (N6326, N6325, N5113, N1014);
or OR3 (N6327, N6324, N291, N4301);
and AND3 (N6328, N6295, N3493, N1799);
xor XOR2 (N6329, N6318, N4549);
or OR3 (N6330, N6327, N3703, N3597);
buf BUF1 (N6331, N6314);
not NOT1 (N6332, N6330);
xor XOR2 (N6333, N6322, N3548);
not NOT1 (N6334, N6301);
buf BUF1 (N6335, N6331);
nand NAND4 (N6336, N6333, N4463, N4165, N1669);
buf BUF1 (N6337, N6321);
and AND4 (N6338, N6337, N2184, N58, N6280);
or OR2 (N6339, N6326, N4042);
nor NOR3 (N6340, N6323, N4476, N2363);
nand NAND2 (N6341, N6338, N281);
nor NOR2 (N6342, N6335, N6056);
or OR4 (N6343, N6336, N3519, N3858, N2453);
buf BUF1 (N6344, N6328);
nand NAND2 (N6345, N6315, N1400);
or OR3 (N6346, N6334, N317, N3913);
nand NAND4 (N6347, N6340, N1374, N2094, N3298);
buf BUF1 (N6348, N6347);
buf BUF1 (N6349, N6332);
nor NOR2 (N6350, N6344, N2532);
xor XOR2 (N6351, N6329, N2937);
and AND4 (N6352, N6342, N6162, N728, N3364);
nor NOR3 (N6353, N6341, N6002, N2776);
xor XOR2 (N6354, N6350, N4420);
and AND4 (N6355, N6345, N2505, N4452, N806);
nand NAND2 (N6356, N6348, N1643);
or OR2 (N6357, N6351, N2693);
nor NOR2 (N6358, N6339, N4496);
and AND3 (N6359, N6343, N937, N6150);
xor XOR2 (N6360, N6355, N6299);
nor NOR4 (N6361, N6352, N3261, N6196, N1618);
xor XOR2 (N6362, N6354, N4413);
or OR3 (N6363, N6362, N600, N1759);
and AND4 (N6364, N6356, N880, N2523, N446);
and AND4 (N6365, N6346, N1835, N4895, N3666);
or OR2 (N6366, N6349, N1803);
nand NAND3 (N6367, N6353, N1161, N3132);
nor NOR2 (N6368, N6358, N1159);
or OR2 (N6369, N6364, N6191);
buf BUF1 (N6370, N6369);
nor NOR2 (N6371, N6367, N552);
nor NOR3 (N6372, N6360, N5476, N5754);
and AND2 (N6373, N6357, N6287);
xor XOR2 (N6374, N6370, N282);
nand NAND3 (N6375, N6363, N2933, N5292);
and AND3 (N6376, N6361, N3058, N592);
xor XOR2 (N6377, N6366, N228);
or OR4 (N6378, N6375, N212, N4739, N4601);
nor NOR2 (N6379, N6359, N3528);
buf BUF1 (N6380, N6372);
nor NOR2 (N6381, N6368, N2177);
nand NAND4 (N6382, N6377, N4718, N2808, N3593);
buf BUF1 (N6383, N6379);
xor XOR2 (N6384, N6378, N3933);
nor NOR2 (N6385, N6373, N1264);
buf BUF1 (N6386, N6385);
buf BUF1 (N6387, N6376);
buf BUF1 (N6388, N6383);
nand NAND2 (N6389, N6386, N5721);
and AND2 (N6390, N6365, N3167);
xor XOR2 (N6391, N6388, N4053);
xor XOR2 (N6392, N6374, N3978);
not NOT1 (N6393, N6382);
buf BUF1 (N6394, N6387);
and AND4 (N6395, N6394, N4841, N1005, N143);
xor XOR2 (N6396, N6390, N4457);
or OR2 (N6397, N6371, N188);
nor NOR2 (N6398, N6393, N905);
and AND3 (N6399, N6395, N4428, N236);
and AND3 (N6400, N6398, N5385, N4931);
xor XOR2 (N6401, N6381, N3075);
or OR2 (N6402, N6380, N2692);
and AND2 (N6403, N6391, N2426);
nand NAND2 (N6404, N6403, N2419);
not NOT1 (N6405, N6396);
not NOT1 (N6406, N6405);
not NOT1 (N6407, N6399);
buf BUF1 (N6408, N6402);
not NOT1 (N6409, N6406);
nor NOR3 (N6410, N6389, N3097, N5312);
or OR3 (N6411, N6400, N3792, N31);
nand NAND2 (N6412, N6410, N3687);
buf BUF1 (N6413, N6392);
nand NAND4 (N6414, N6413, N6141, N5661, N2721);
xor XOR2 (N6415, N6409, N1982);
nor NOR4 (N6416, N6408, N2852, N5625, N411);
not NOT1 (N6417, N6401);
nor NOR2 (N6418, N6416, N1670);
nand NAND2 (N6419, N6412, N5970);
nor NOR3 (N6420, N6407, N2036, N537);
or OR3 (N6421, N6417, N3877, N1599);
nor NOR4 (N6422, N6404, N4955, N4912, N4806);
not NOT1 (N6423, N6422);
nand NAND4 (N6424, N6423, N5781, N809, N5526);
nand NAND3 (N6425, N6419, N705, N5201);
buf BUF1 (N6426, N6415);
buf BUF1 (N6427, N6425);
buf BUF1 (N6428, N6414);
or OR2 (N6429, N6397, N6038);
or OR4 (N6430, N6424, N5721, N1125, N2239);
xor XOR2 (N6431, N6418, N4963);
nor NOR4 (N6432, N6384, N2303, N2724, N3839);
not NOT1 (N6433, N6431);
and AND3 (N6434, N6432, N2702, N2876);
or OR2 (N6435, N6433, N3452);
nand NAND2 (N6436, N6427, N2337);
or OR2 (N6437, N6411, N3872);
nor NOR2 (N6438, N6434, N4953);
buf BUF1 (N6439, N6429);
nand NAND2 (N6440, N6437, N5935);
xor XOR2 (N6441, N6438, N471);
buf BUF1 (N6442, N6441);
and AND4 (N6443, N6420, N2726, N1737, N2862);
not NOT1 (N6444, N6435);
or OR2 (N6445, N6436, N40);
or OR3 (N6446, N6439, N4743, N2624);
buf BUF1 (N6447, N6442);
xor XOR2 (N6448, N6447, N5231);
or OR4 (N6449, N6421, N3734, N2708, N4549);
buf BUF1 (N6450, N6443);
xor XOR2 (N6451, N6446, N232);
buf BUF1 (N6452, N6426);
and AND3 (N6453, N6445, N5799, N5547);
xor XOR2 (N6454, N6444, N1577);
nand NAND2 (N6455, N6454, N6205);
buf BUF1 (N6456, N6448);
nand NAND3 (N6457, N6428, N793, N5496);
not NOT1 (N6458, N6450);
xor XOR2 (N6459, N6453, N795);
buf BUF1 (N6460, N6458);
not NOT1 (N6461, N6455);
not NOT1 (N6462, N6457);
or OR3 (N6463, N6461, N5583, N5317);
xor XOR2 (N6464, N6463, N1477);
or OR4 (N6465, N6464, N4552, N3229, N2398);
or OR4 (N6466, N6462, N5817, N5616, N1901);
xor XOR2 (N6467, N6465, N1309);
or OR3 (N6468, N6467, N4523, N1626);
nand NAND3 (N6469, N6460, N1377, N5146);
xor XOR2 (N6470, N6452, N2520);
or OR4 (N6471, N6451, N4000, N3970, N154);
xor XOR2 (N6472, N6440, N67);
nand NAND4 (N6473, N6430, N5176, N3192, N5781);
or OR2 (N6474, N6469, N346);
nand NAND4 (N6475, N6472, N4807, N5060, N1095);
xor XOR2 (N6476, N6459, N4379);
nand NAND4 (N6477, N6473, N5143, N6253, N4193);
or OR4 (N6478, N6456, N5723, N3270, N1172);
nand NAND2 (N6479, N6476, N2137);
nor NOR3 (N6480, N6479, N5638, N2992);
or OR4 (N6481, N6466, N3157, N2389, N749);
xor XOR2 (N6482, N6474, N701);
nand NAND2 (N6483, N6481, N6052);
nand NAND3 (N6484, N6482, N978, N196);
nor NOR3 (N6485, N6449, N2786, N4659);
buf BUF1 (N6486, N6485);
buf BUF1 (N6487, N6486);
xor XOR2 (N6488, N6468, N2806);
buf BUF1 (N6489, N6475);
xor XOR2 (N6490, N6483, N1237);
nand NAND2 (N6491, N6488, N1067);
or OR3 (N6492, N6480, N2603, N750);
nor NOR4 (N6493, N6470, N3949, N1870, N1234);
xor XOR2 (N6494, N6493, N5622);
not NOT1 (N6495, N6471);
and AND2 (N6496, N6492, N5738);
nor NOR3 (N6497, N6478, N1422, N4604);
nand NAND4 (N6498, N6484, N6168, N3712, N5925);
and AND4 (N6499, N6487, N1469, N5128, N5171);
buf BUF1 (N6500, N6490);
not NOT1 (N6501, N6499);
and AND4 (N6502, N6489, N5489, N4507, N1958);
nor NOR3 (N6503, N6497, N576, N2751);
or OR2 (N6504, N6503, N2794);
and AND4 (N6505, N6477, N4257, N931, N3630);
nand NAND4 (N6506, N6491, N13, N3113, N3472);
buf BUF1 (N6507, N6496);
not NOT1 (N6508, N6495);
xor XOR2 (N6509, N6506, N2003);
xor XOR2 (N6510, N6509, N461);
and AND3 (N6511, N6510, N5250, N922);
or OR3 (N6512, N6511, N5138, N2685);
nand NAND4 (N6513, N6501, N1800, N3374, N2463);
nor NOR4 (N6514, N6505, N6374, N3746, N1732);
nand NAND2 (N6515, N6504, N4933);
or OR3 (N6516, N6507, N1908, N3225);
not NOT1 (N6517, N6498);
or OR2 (N6518, N6514, N2343);
and AND3 (N6519, N6508, N6245, N3499);
nor NOR3 (N6520, N6494, N1950, N2070);
not NOT1 (N6521, N6518);
buf BUF1 (N6522, N6512);
or OR2 (N6523, N6519, N1098);
nand NAND2 (N6524, N6502, N3339);
nand NAND3 (N6525, N6523, N1654, N5549);
not NOT1 (N6526, N6521);
nor NOR2 (N6527, N6526, N2124);
nand NAND2 (N6528, N6527, N3504);
and AND3 (N6529, N6524, N4729, N2611);
or OR3 (N6530, N6515, N2237, N1359);
or OR3 (N6531, N6516, N2609, N1263);
buf BUF1 (N6532, N6517);
or OR4 (N6533, N6513, N1628, N5674, N1671);
nor NOR4 (N6534, N6520, N6010, N896, N4003);
buf BUF1 (N6535, N6525);
and AND4 (N6536, N6535, N5813, N6269, N1439);
nand NAND4 (N6537, N6528, N3033, N1344, N3386);
nor NOR4 (N6538, N6532, N3741, N5154, N6268);
buf BUF1 (N6539, N6538);
not NOT1 (N6540, N6522);
nand NAND3 (N6541, N6536, N4323, N6185);
not NOT1 (N6542, N6533);
and AND2 (N6543, N6537, N4658);
nand NAND4 (N6544, N6541, N3799, N6010, N4593);
or OR4 (N6545, N6529, N1172, N2034, N2381);
or OR3 (N6546, N6539, N5992, N440);
buf BUF1 (N6547, N6540);
xor XOR2 (N6548, N6542, N3353);
and AND3 (N6549, N6548, N6279, N1412);
and AND2 (N6550, N6531, N4953);
xor XOR2 (N6551, N6550, N693);
nor NOR3 (N6552, N6547, N3427, N3701);
xor XOR2 (N6553, N6546, N3785);
buf BUF1 (N6554, N6545);
or OR3 (N6555, N6554, N5436, N4868);
or OR2 (N6556, N6543, N5875);
nor NOR4 (N6557, N6534, N2343, N307, N4157);
nand NAND2 (N6558, N6549, N299);
or OR2 (N6559, N6555, N2461);
or OR3 (N6560, N6553, N298, N60);
nand NAND2 (N6561, N6530, N5370);
not NOT1 (N6562, N6500);
not NOT1 (N6563, N6561);
or OR4 (N6564, N6563, N3617, N5385, N5415);
nand NAND4 (N6565, N6560, N4082, N6430, N5565);
nor NOR2 (N6566, N6558, N4705);
nand NAND3 (N6567, N6556, N5057, N5800);
not NOT1 (N6568, N6562);
or OR4 (N6569, N6568, N1378, N662, N1587);
not NOT1 (N6570, N6567);
and AND3 (N6571, N6557, N4092, N2702);
and AND4 (N6572, N6564, N2708, N533, N6090);
buf BUF1 (N6573, N6544);
or OR4 (N6574, N6573, N162, N2910, N6502);
buf BUF1 (N6575, N6574);
or OR3 (N6576, N6572, N31, N4105);
not NOT1 (N6577, N6571);
or OR2 (N6578, N6575, N926);
and AND2 (N6579, N6551, N6403);
nor NOR4 (N6580, N6578, N98, N158, N4005);
nor NOR4 (N6581, N6579, N5523, N3173, N888);
nand NAND2 (N6582, N6559, N6498);
or OR3 (N6583, N6582, N4571, N216);
buf BUF1 (N6584, N6581);
xor XOR2 (N6585, N6552, N2263);
buf BUF1 (N6586, N6569);
or OR4 (N6587, N6585, N6403, N1917, N889);
not NOT1 (N6588, N6587);
nor NOR3 (N6589, N6584, N2172, N1243);
xor XOR2 (N6590, N6586, N5227);
buf BUF1 (N6591, N6588);
or OR3 (N6592, N6570, N3949, N5931);
or OR2 (N6593, N6576, N635);
not NOT1 (N6594, N6580);
nand NAND3 (N6595, N6589, N4282, N1213);
nand NAND3 (N6596, N6594, N2548, N1477);
nor NOR2 (N6597, N6592, N5057);
not NOT1 (N6598, N6597);
not NOT1 (N6599, N6598);
nand NAND2 (N6600, N6565, N2353);
and AND2 (N6601, N6593, N4870);
nor NOR3 (N6602, N6599, N2510, N5847);
xor XOR2 (N6603, N6583, N1012);
nand NAND4 (N6604, N6600, N2636, N2070, N4841);
buf BUF1 (N6605, N6591);
xor XOR2 (N6606, N6605, N1873);
xor XOR2 (N6607, N6602, N1052);
xor XOR2 (N6608, N6596, N4946);
not NOT1 (N6609, N6566);
not NOT1 (N6610, N6604);
xor XOR2 (N6611, N6609, N4112);
xor XOR2 (N6612, N6577, N2389);
or OR3 (N6613, N6606, N5490, N3276);
nor NOR3 (N6614, N6613, N3485, N1632);
nand NAND2 (N6615, N6611, N3994);
or OR4 (N6616, N6612, N4092, N3890, N1564);
buf BUF1 (N6617, N6595);
nand NAND3 (N6618, N6607, N3416, N6532);
or OR3 (N6619, N6616, N3224, N2181);
buf BUF1 (N6620, N6608);
xor XOR2 (N6621, N6618, N3113);
and AND4 (N6622, N6619, N2810, N5452, N1324);
not NOT1 (N6623, N6601);
nand NAND3 (N6624, N6614, N3324, N1629);
and AND3 (N6625, N6603, N793, N2192);
nand NAND4 (N6626, N6617, N6588, N6390, N6457);
not NOT1 (N6627, N6624);
and AND3 (N6628, N6610, N4562, N1323);
and AND2 (N6629, N6621, N2826);
not NOT1 (N6630, N6628);
or OR3 (N6631, N6629, N4361, N805);
xor XOR2 (N6632, N6625, N1049);
not NOT1 (N6633, N6627);
buf BUF1 (N6634, N6626);
nor NOR4 (N6635, N6632, N6554, N4741, N3480);
nor NOR2 (N6636, N6622, N3107);
or OR2 (N6637, N6623, N2030);
not NOT1 (N6638, N6635);
xor XOR2 (N6639, N6590, N3189);
nor NOR3 (N6640, N6615, N2769, N6290);
not NOT1 (N6641, N6640);
and AND4 (N6642, N6641, N106, N1439, N2176);
and AND3 (N6643, N6638, N6079, N6608);
nor NOR2 (N6644, N6639, N2514);
nor NOR2 (N6645, N6634, N897);
and AND3 (N6646, N6633, N5882, N3526);
nor NOR3 (N6647, N6643, N3150, N4110);
nor NOR2 (N6648, N6637, N4283);
buf BUF1 (N6649, N6648);
not NOT1 (N6650, N6630);
and AND2 (N6651, N6644, N6420);
xor XOR2 (N6652, N6651, N4664);
or OR2 (N6653, N6620, N6160);
not NOT1 (N6654, N6650);
or OR4 (N6655, N6647, N3573, N1136, N5772);
buf BUF1 (N6656, N6655);
or OR4 (N6657, N6645, N282, N1652, N5098);
nand NAND2 (N6658, N6646, N5749);
nor NOR3 (N6659, N6642, N385, N2791);
buf BUF1 (N6660, N6636);
nand NAND4 (N6661, N6631, N910, N999, N1276);
and AND3 (N6662, N6656, N4449, N5683);
nor NOR3 (N6663, N6654, N3325, N4457);
or OR2 (N6664, N6653, N3908);
nand NAND4 (N6665, N6660, N3258, N3966, N4725);
nor NOR2 (N6666, N6663, N4270);
buf BUF1 (N6667, N6652);
not NOT1 (N6668, N6649);
nor NOR3 (N6669, N6665, N6565, N5086);
and AND4 (N6670, N6668, N90, N4725, N1951);
not NOT1 (N6671, N6657);
nor NOR3 (N6672, N6658, N5649, N5098);
and AND3 (N6673, N6662, N1218, N2535);
nand NAND4 (N6674, N6672, N2683, N1944, N6627);
nor NOR4 (N6675, N6669, N5075, N3739, N1418);
or OR2 (N6676, N6674, N1642);
buf BUF1 (N6677, N6673);
xor XOR2 (N6678, N6664, N5135);
or OR2 (N6679, N6675, N5411);
not NOT1 (N6680, N6667);
or OR3 (N6681, N6678, N4869, N2312);
nand NAND2 (N6682, N6676, N5163);
buf BUF1 (N6683, N6679);
nor NOR3 (N6684, N6680, N6058, N6099);
xor XOR2 (N6685, N6681, N5146);
nand NAND4 (N6686, N6684, N1440, N1396, N1523);
nand NAND2 (N6687, N6671, N4904);
buf BUF1 (N6688, N6686);
and AND2 (N6689, N6687, N1387);
nor NOR3 (N6690, N6661, N5405, N3996);
nor NOR3 (N6691, N6659, N4353, N3992);
not NOT1 (N6692, N6690);
nand NAND4 (N6693, N6683, N2040, N2443, N4412);
xor XOR2 (N6694, N6688, N1649);
or OR2 (N6695, N6691, N34);
not NOT1 (N6696, N6692);
and AND4 (N6697, N6689, N3043, N211, N5846);
xor XOR2 (N6698, N6696, N3378);
buf BUF1 (N6699, N6695);
nand NAND4 (N6700, N6677, N3695, N1202, N5418);
xor XOR2 (N6701, N6693, N881);
buf BUF1 (N6702, N6698);
nand NAND2 (N6703, N6700, N6532);
and AND3 (N6704, N6702, N2149, N4927);
not NOT1 (N6705, N6682);
buf BUF1 (N6706, N6694);
nor NOR3 (N6707, N6706, N1313, N5036);
xor XOR2 (N6708, N6666, N1318);
not NOT1 (N6709, N6705);
nand NAND3 (N6710, N6703, N5857, N1088);
nand NAND3 (N6711, N6685, N507, N2227);
or OR2 (N6712, N6710, N3505);
or OR3 (N6713, N6707, N4483, N6089);
and AND4 (N6714, N6701, N6633, N5245, N4001);
buf BUF1 (N6715, N6713);
not NOT1 (N6716, N6714);
and AND3 (N6717, N6670, N6041, N4397);
not NOT1 (N6718, N6708);
not NOT1 (N6719, N6699);
or OR2 (N6720, N6716, N1732);
buf BUF1 (N6721, N6718);
nand NAND4 (N6722, N6704, N3924, N3155, N227);
not NOT1 (N6723, N6697);
or OR2 (N6724, N6711, N1200);
nor NOR2 (N6725, N6720, N4387);
or OR4 (N6726, N6725, N3179, N3185, N5925);
nand NAND4 (N6727, N6709, N819, N5764, N1330);
or OR4 (N6728, N6724, N4595, N4131, N1362);
xor XOR2 (N6729, N6726, N2110);
not NOT1 (N6730, N6712);
buf BUF1 (N6731, N6729);
or OR3 (N6732, N6730, N2696, N2458);
buf BUF1 (N6733, N6728);
xor XOR2 (N6734, N6715, N1233);
and AND2 (N6735, N6733, N4413);
and AND2 (N6736, N6722, N564);
not NOT1 (N6737, N6717);
xor XOR2 (N6738, N6721, N3691);
nand NAND4 (N6739, N6727, N4998, N3010, N1573);
nand NAND4 (N6740, N6732, N508, N3911, N6052);
nor NOR4 (N6741, N6734, N6016, N1832, N5166);
or OR3 (N6742, N6731, N43, N5005);
xor XOR2 (N6743, N6736, N4813);
nor NOR2 (N6744, N6737, N3205);
buf BUF1 (N6745, N6741);
xor XOR2 (N6746, N6744, N3144);
nor NOR4 (N6747, N6735, N4335, N1089, N4836);
not NOT1 (N6748, N6742);
nand NAND2 (N6749, N6745, N1239);
nand NAND4 (N6750, N6740, N1113, N4194, N2858);
and AND3 (N6751, N6723, N3041, N4884);
nand NAND3 (N6752, N6719, N5582, N2733);
nand NAND2 (N6753, N6748, N536);
nand NAND2 (N6754, N6739, N662);
xor XOR2 (N6755, N6751, N1757);
nand NAND4 (N6756, N6747, N5336, N1970, N156);
buf BUF1 (N6757, N6755);
xor XOR2 (N6758, N6750, N2332);
buf BUF1 (N6759, N6743);
xor XOR2 (N6760, N6746, N6220);
and AND4 (N6761, N6757, N1761, N6532, N6679);
buf BUF1 (N6762, N6738);
not NOT1 (N6763, N6758);
xor XOR2 (N6764, N6761, N2772);
not NOT1 (N6765, N6759);
not NOT1 (N6766, N6760);
and AND3 (N6767, N6754, N2774, N3040);
xor XOR2 (N6768, N6767, N3949);
buf BUF1 (N6769, N6756);
nor NOR2 (N6770, N6753, N5624);
xor XOR2 (N6771, N6768, N2269);
and AND2 (N6772, N6763, N5238);
nor NOR4 (N6773, N6764, N4246, N436, N351);
not NOT1 (N6774, N6769);
nor NOR4 (N6775, N6766, N3839, N5848, N173);
buf BUF1 (N6776, N6762);
xor XOR2 (N6777, N6772, N3037);
buf BUF1 (N6778, N6773);
nand NAND2 (N6779, N6777, N4009);
or OR3 (N6780, N6765, N1644, N2846);
or OR2 (N6781, N6778, N5015);
not NOT1 (N6782, N6779);
xor XOR2 (N6783, N6774, N937);
xor XOR2 (N6784, N6781, N2792);
nor NOR2 (N6785, N6775, N2610);
or OR2 (N6786, N6776, N6090);
and AND4 (N6787, N6785, N6279, N365, N4469);
nor NOR4 (N6788, N6752, N4779, N1199, N5358);
not NOT1 (N6789, N6787);
nor NOR2 (N6790, N6784, N3047);
buf BUF1 (N6791, N6790);
buf BUF1 (N6792, N6749);
nand NAND4 (N6793, N6771, N1575, N35, N753);
not NOT1 (N6794, N6783);
not NOT1 (N6795, N6794);
and AND2 (N6796, N6792, N4384);
or OR4 (N6797, N6793, N3917, N4005, N2072);
and AND4 (N6798, N6789, N3698, N2239, N167);
not NOT1 (N6799, N6795);
xor XOR2 (N6800, N6799, N2195);
or OR4 (N6801, N6791, N2645, N2400, N1814);
or OR2 (N6802, N6800, N3232);
not NOT1 (N6803, N6788);
buf BUF1 (N6804, N6786);
and AND4 (N6805, N6804, N2574, N6724, N704);
not NOT1 (N6806, N6770);
nor NOR4 (N6807, N6797, N1277, N5399, N3427);
and AND3 (N6808, N6807, N6622, N727);
or OR3 (N6809, N6798, N3377, N2358);
or OR3 (N6810, N6806, N557, N4459);
xor XOR2 (N6811, N6803, N573);
nor NOR3 (N6812, N6805, N4793, N5951);
not NOT1 (N6813, N6808);
nor NOR3 (N6814, N6796, N3362, N1799);
nand NAND4 (N6815, N6810, N845, N39, N36);
xor XOR2 (N6816, N6801, N1748);
buf BUF1 (N6817, N6809);
nand NAND3 (N6818, N6815, N538, N5368);
and AND4 (N6819, N6811, N2931, N635, N6265);
and AND3 (N6820, N6816, N5387, N4950);
or OR3 (N6821, N6782, N4735, N1629);
nand NAND2 (N6822, N6813, N6051);
and AND3 (N6823, N6817, N1491, N6530);
buf BUF1 (N6824, N6823);
nand NAND3 (N6825, N6820, N5641, N6157);
or OR3 (N6826, N6825, N5137, N621);
buf BUF1 (N6827, N6821);
not NOT1 (N6828, N6827);
buf BUF1 (N6829, N6824);
or OR4 (N6830, N6818, N1259, N4042, N3420);
not NOT1 (N6831, N6830);
nor NOR2 (N6832, N6802, N2221);
or OR4 (N6833, N6826, N1416, N1511, N4935);
nor NOR2 (N6834, N6829, N6693);
and AND3 (N6835, N6812, N1840, N2699);
nor NOR3 (N6836, N6834, N1760, N3374);
and AND2 (N6837, N6828, N452);
not NOT1 (N6838, N6833);
not NOT1 (N6839, N6835);
nor NOR2 (N6840, N6838, N5022);
xor XOR2 (N6841, N6839, N1400);
nor NOR3 (N6842, N6819, N1484, N6724);
and AND4 (N6843, N6842, N4634, N2431, N5595);
or OR2 (N6844, N6836, N5588);
nor NOR2 (N6845, N6780, N6373);
nand NAND3 (N6846, N6831, N3862, N5240);
nand NAND2 (N6847, N6841, N1769);
nor NOR4 (N6848, N6847, N2673, N1367, N4305);
xor XOR2 (N6849, N6848, N3660);
xor XOR2 (N6850, N6849, N4395);
nand NAND2 (N6851, N6840, N3238);
and AND3 (N6852, N6814, N616, N56);
nor NOR3 (N6853, N6846, N5436, N3311);
not NOT1 (N6854, N6852);
and AND4 (N6855, N6845, N1731, N4589, N2564);
buf BUF1 (N6856, N6851);
and AND3 (N6857, N6856, N3452, N268);
xor XOR2 (N6858, N6855, N778);
not NOT1 (N6859, N6858);
nor NOR2 (N6860, N6854, N5015);
nor NOR2 (N6861, N6859, N748);
or OR4 (N6862, N6832, N5991, N6456, N5851);
or OR2 (N6863, N6860, N3804);
or OR3 (N6864, N6850, N1437, N6062);
and AND4 (N6865, N6864, N2350, N1050, N1398);
nand NAND4 (N6866, N6837, N1688, N1747, N3407);
nor NOR4 (N6867, N6861, N3185, N2740, N1975);
buf BUF1 (N6868, N6866);
or OR2 (N6869, N6868, N6119);
nor NOR3 (N6870, N6857, N1717, N812);
or OR3 (N6871, N6862, N4408, N5345);
xor XOR2 (N6872, N6869, N6425);
not NOT1 (N6873, N6843);
not NOT1 (N6874, N6870);
and AND4 (N6875, N6867, N3689, N5425, N4603);
buf BUF1 (N6876, N6872);
and AND4 (N6877, N6874, N2756, N1239, N3619);
nor NOR4 (N6878, N6844, N561, N212, N3654);
nand NAND3 (N6879, N6871, N1130, N1683);
buf BUF1 (N6880, N6873);
and AND2 (N6881, N6880, N4777);
and AND3 (N6882, N6863, N500, N4757);
nand NAND4 (N6883, N6853, N5479, N349, N3533);
nor NOR4 (N6884, N6883, N596, N6065, N2183);
xor XOR2 (N6885, N6879, N971);
xor XOR2 (N6886, N6884, N4351);
not NOT1 (N6887, N6877);
and AND2 (N6888, N6878, N1402);
and AND3 (N6889, N6881, N6512, N6183);
buf BUF1 (N6890, N6865);
not NOT1 (N6891, N6888);
and AND3 (N6892, N6876, N4725, N554);
nor NOR2 (N6893, N6887, N6507);
nand NAND3 (N6894, N6875, N254, N6159);
nand NAND2 (N6895, N6886, N5210);
or OR2 (N6896, N6822, N5729);
and AND4 (N6897, N6885, N5826, N2489, N2218);
nand NAND4 (N6898, N6890, N6868, N1793, N4915);
nor NOR3 (N6899, N6894, N3018, N6503);
not NOT1 (N6900, N6895);
xor XOR2 (N6901, N6892, N3037);
xor XOR2 (N6902, N6891, N3980);
and AND4 (N6903, N6896, N2874, N1464, N2532);
and AND2 (N6904, N6901, N3623);
or OR3 (N6905, N6893, N5592, N4975);
nor NOR3 (N6906, N6900, N2123, N5438);
xor XOR2 (N6907, N6899, N5717);
nand NAND2 (N6908, N6882, N4949);
and AND4 (N6909, N6905, N5170, N4457, N4813);
nand NAND3 (N6910, N6908, N2294, N4128);
and AND2 (N6911, N6906, N3864);
xor XOR2 (N6912, N6898, N3903);
not NOT1 (N6913, N6902);
nand NAND2 (N6914, N6909, N1540);
not NOT1 (N6915, N6911);
or OR4 (N6916, N6897, N2879, N532, N6412);
nand NAND4 (N6917, N6912, N2188, N5551, N6169);
and AND2 (N6918, N6910, N403);
xor XOR2 (N6919, N6914, N2145);
nand NAND3 (N6920, N6907, N1886, N502);
or OR4 (N6921, N6919, N3884, N991, N1385);
buf BUF1 (N6922, N6904);
nand NAND3 (N6923, N6921, N1197, N4991);
and AND2 (N6924, N6913, N4243);
nand NAND4 (N6925, N6922, N6913, N3810, N5208);
buf BUF1 (N6926, N6915);
or OR2 (N6927, N6903, N5665);
not NOT1 (N6928, N6920);
xor XOR2 (N6929, N6926, N2255);
nor NOR4 (N6930, N6923, N476, N6801, N6564);
buf BUF1 (N6931, N6930);
buf BUF1 (N6932, N6924);
nor NOR4 (N6933, N6928, N874, N975, N4111);
and AND3 (N6934, N6929, N878, N806);
not NOT1 (N6935, N6934);
xor XOR2 (N6936, N6925, N4975);
not NOT1 (N6937, N6935);
xor XOR2 (N6938, N6933, N5686);
or OR3 (N6939, N6918, N462, N6514);
or OR4 (N6940, N6916, N5839, N1911, N2484);
xor XOR2 (N6941, N6927, N159);
xor XOR2 (N6942, N6941, N5701);
nor NOR4 (N6943, N6936, N2498, N5938, N6751);
nor NOR4 (N6944, N6940, N3801, N3997, N3272);
not NOT1 (N6945, N6931);
and AND3 (N6946, N6889, N3294, N4422);
and AND2 (N6947, N6943, N6595);
nand NAND4 (N6948, N6938, N462, N5563, N2292);
nand NAND2 (N6949, N6939, N6921);
and AND4 (N6950, N6947, N5968, N1429, N4694);
or OR4 (N6951, N6937, N3853, N2847, N4203);
not NOT1 (N6952, N6944);
nand NAND2 (N6953, N6942, N6650);
not NOT1 (N6954, N6946);
nand NAND3 (N6955, N6948, N4375, N5275);
nand NAND2 (N6956, N6917, N5514);
nor NOR4 (N6957, N6952, N3167, N6744, N3935);
nand NAND2 (N6958, N6951, N1327);
nand NAND3 (N6959, N6957, N3055, N1319);
not NOT1 (N6960, N6949);
buf BUF1 (N6961, N6953);
xor XOR2 (N6962, N6954, N2186);
nand NAND4 (N6963, N6961, N5860, N4298, N4835);
and AND4 (N6964, N6932, N6064, N5289, N622);
nand NAND4 (N6965, N6960, N5375, N403, N830);
nor NOR3 (N6966, N6962, N6862, N1699);
not NOT1 (N6967, N6956);
or OR3 (N6968, N6955, N2455, N1347);
nor NOR2 (N6969, N6950, N2693);
not NOT1 (N6970, N6959);
not NOT1 (N6971, N6967);
or OR4 (N6972, N6969, N4065, N1292, N279);
not NOT1 (N6973, N6971);
xor XOR2 (N6974, N6965, N2425);
nand NAND4 (N6975, N6963, N4491, N849, N5594);
buf BUF1 (N6976, N6968);
nand NAND2 (N6977, N6976, N5369);
not NOT1 (N6978, N6974);
nand NAND4 (N6979, N6973, N5645, N1788, N1259);
nor NOR3 (N6980, N6958, N2721, N347);
nor NOR3 (N6981, N6945, N6263, N6485);
nand NAND2 (N6982, N6981, N4278);
nand NAND4 (N6983, N6966, N3143, N5923, N5577);
nor NOR2 (N6984, N6982, N4430);
xor XOR2 (N6985, N6980, N5960);
nor NOR2 (N6986, N6970, N441);
not NOT1 (N6987, N6985);
or OR2 (N6988, N6964, N1146);
nand NAND3 (N6989, N6977, N3255, N2537);
buf BUF1 (N6990, N6972);
or OR4 (N6991, N6990, N249, N2472, N6683);
xor XOR2 (N6992, N6983, N2350);
xor XOR2 (N6993, N6979, N1256);
or OR3 (N6994, N6993, N6315, N6090);
nor NOR3 (N6995, N6989, N6455, N699);
or OR2 (N6996, N6991, N1999);
xor XOR2 (N6997, N6984, N4554);
not NOT1 (N6998, N6994);
not NOT1 (N6999, N6998);
not NOT1 (N7000, N6988);
and AND4 (N7001, N6996, N2593, N3089, N4905);
or OR3 (N7002, N6995, N2174, N5618);
nor NOR3 (N7003, N7001, N5232, N4320);
or OR3 (N7004, N6978, N6579, N2857);
nand NAND3 (N7005, N7002, N6971, N6970);
and AND3 (N7006, N6999, N2395, N828);
not NOT1 (N7007, N7005);
not NOT1 (N7008, N7007);
nand NAND2 (N7009, N7006, N5827);
buf BUF1 (N7010, N6986);
buf BUF1 (N7011, N6987);
not NOT1 (N7012, N7000);
buf BUF1 (N7013, N7004);
buf BUF1 (N7014, N7012);
xor XOR2 (N7015, N6975, N5224);
or OR2 (N7016, N7014, N3374);
or OR4 (N7017, N6992, N3053, N1186, N494);
buf BUF1 (N7018, N7015);
and AND4 (N7019, N7017, N5305, N593, N1546);
nor NOR2 (N7020, N7010, N3791);
not NOT1 (N7021, N7019);
nor NOR3 (N7022, N7018, N5382, N3618);
and AND3 (N7023, N7021, N2921, N1147);
and AND2 (N7024, N7009, N2537);
buf BUF1 (N7025, N7013);
xor XOR2 (N7026, N7023, N7);
nor NOR2 (N7027, N7016, N5139);
and AND4 (N7028, N6997, N3830, N1898, N1016);
not NOT1 (N7029, N7026);
nor NOR3 (N7030, N7022, N3900, N5525);
or OR4 (N7031, N7008, N520, N6192, N2121);
or OR3 (N7032, N7003, N1280, N5704);
buf BUF1 (N7033, N7025);
or OR3 (N7034, N7020, N6082, N6846);
buf BUF1 (N7035, N7032);
nand NAND2 (N7036, N7031, N6823);
and AND2 (N7037, N7036, N5188);
xor XOR2 (N7038, N7030, N871);
nor NOR3 (N7039, N7028, N3791, N5631);
buf BUF1 (N7040, N7029);
nor NOR3 (N7041, N7038, N4858, N5576);
nor NOR2 (N7042, N7041, N4670);
or OR2 (N7043, N7037, N1930);
and AND2 (N7044, N7011, N1534);
buf BUF1 (N7045, N7027);
not NOT1 (N7046, N7044);
buf BUF1 (N7047, N7033);
nor NOR4 (N7048, N7024, N303, N3414, N1148);
or OR3 (N7049, N7047, N989, N4100);
buf BUF1 (N7050, N7042);
xor XOR2 (N7051, N7043, N6171);
not NOT1 (N7052, N7045);
nor NOR3 (N7053, N7048, N1615, N6041);
buf BUF1 (N7054, N7050);
not NOT1 (N7055, N7049);
buf BUF1 (N7056, N7046);
nand NAND3 (N7057, N7053, N2429, N311);
nand NAND3 (N7058, N7057, N1804, N4997);
not NOT1 (N7059, N7051);
not NOT1 (N7060, N7058);
and AND4 (N7061, N7034, N2979, N5898, N5066);
nand NAND4 (N7062, N7060, N3225, N3511, N2109);
nor NOR3 (N7063, N7056, N2867, N4203);
xor XOR2 (N7064, N7039, N6398);
buf BUF1 (N7065, N7055);
not NOT1 (N7066, N7059);
buf BUF1 (N7067, N7065);
not NOT1 (N7068, N7066);
buf BUF1 (N7069, N7035);
buf BUF1 (N7070, N7052);
or OR2 (N7071, N7054, N2473);
not NOT1 (N7072, N7062);
xor XOR2 (N7073, N7071, N1571);
not NOT1 (N7074, N7068);
or OR2 (N7075, N7069, N4141);
not NOT1 (N7076, N7061);
not NOT1 (N7077, N7063);
nand NAND4 (N7078, N7072, N6691, N2775, N4637);
or OR2 (N7079, N7074, N2667);
xor XOR2 (N7080, N7073, N4069);
nand NAND2 (N7081, N7064, N3182);
nand NAND4 (N7082, N7078, N4547, N6463, N4440);
or OR4 (N7083, N7080, N2479, N236, N5872);
not NOT1 (N7084, N7075);
buf BUF1 (N7085, N7067);
buf BUF1 (N7086, N7085);
nand NAND2 (N7087, N7086, N6287);
and AND2 (N7088, N7076, N2198);
xor XOR2 (N7089, N7082, N6988);
nand NAND3 (N7090, N7088, N6851, N6732);
buf BUF1 (N7091, N7077);
or OR4 (N7092, N7079, N3382, N3802, N3846);
buf BUF1 (N7093, N7081);
and AND3 (N7094, N7083, N289, N1359);
buf BUF1 (N7095, N7070);
nor NOR4 (N7096, N7087, N3066, N2641, N5207);
buf BUF1 (N7097, N7093);
and AND4 (N7098, N7040, N1570, N3212, N2555);
not NOT1 (N7099, N7090);
nor NOR3 (N7100, N7094, N2816, N3215);
xor XOR2 (N7101, N7091, N2572);
nor NOR3 (N7102, N7092, N1409, N3255);
and AND3 (N7103, N7084, N2714, N567);
xor XOR2 (N7104, N7102, N557);
xor XOR2 (N7105, N7100, N6315);
or OR2 (N7106, N7095, N5396);
buf BUF1 (N7107, N7101);
and AND2 (N7108, N7096, N6190);
and AND2 (N7109, N7104, N5393);
nand NAND4 (N7110, N7097, N3737, N3863, N2571);
not NOT1 (N7111, N7089);
xor XOR2 (N7112, N7106, N5629);
and AND3 (N7113, N7098, N3739, N4236);
xor XOR2 (N7114, N7111, N4464);
or OR3 (N7115, N7114, N596, N501);
not NOT1 (N7116, N7107);
nor NOR4 (N7117, N7116, N2543, N6591, N268);
nor NOR3 (N7118, N7117, N2013, N504);
or OR4 (N7119, N7099, N3091, N5167, N5738);
nand NAND2 (N7120, N7115, N1633);
xor XOR2 (N7121, N7103, N3929);
or OR3 (N7122, N7121, N5854, N5750);
buf BUF1 (N7123, N7119);
and AND4 (N7124, N7113, N2500, N4836, N5405);
nor NOR2 (N7125, N7120, N5378);
nand NAND2 (N7126, N7124, N683);
xor XOR2 (N7127, N7118, N2176);
or OR2 (N7128, N7105, N899);
or OR3 (N7129, N7122, N2479, N615);
xor XOR2 (N7130, N7110, N5090);
buf BUF1 (N7131, N7128);
and AND3 (N7132, N7126, N2944, N2102);
or OR3 (N7133, N7123, N4500, N1646);
or OR3 (N7134, N7112, N3625, N5432);
nor NOR3 (N7135, N7127, N6455, N1936);
nor NOR4 (N7136, N7134, N537, N6381, N3326);
and AND4 (N7137, N7109, N1811, N5652, N694);
and AND4 (N7138, N7125, N1456, N2496, N5307);
and AND4 (N7139, N7136, N3256, N5546, N3253);
nor NOR3 (N7140, N7130, N687, N2800);
not NOT1 (N7141, N7129);
nand NAND3 (N7142, N7131, N6166, N1179);
xor XOR2 (N7143, N7140, N6437);
or OR4 (N7144, N7138, N2174, N1094, N1);
nand NAND2 (N7145, N7108, N378);
nor NOR3 (N7146, N7139, N5027, N4427);
nand NAND3 (N7147, N7146, N6850, N1325);
buf BUF1 (N7148, N7141);
xor XOR2 (N7149, N7137, N5498);
nor NOR4 (N7150, N7142, N5896, N650, N4960);
or OR2 (N7151, N7143, N7116);
nor NOR3 (N7152, N7144, N425, N6565);
not NOT1 (N7153, N7152);
or OR4 (N7154, N7145, N1954, N539, N4787);
or OR2 (N7155, N7148, N5816);
not NOT1 (N7156, N7153);
nand NAND2 (N7157, N7132, N5196);
nand NAND3 (N7158, N7135, N4930, N1631);
not NOT1 (N7159, N7158);
and AND4 (N7160, N7155, N1665, N1404, N6924);
nor NOR2 (N7161, N7147, N6989);
and AND4 (N7162, N7133, N2242, N2645, N1713);
or OR3 (N7163, N7162, N1232, N2045);
xor XOR2 (N7164, N7163, N6695);
buf BUF1 (N7165, N7157);
nand NAND3 (N7166, N7149, N6440, N4178);
nand NAND2 (N7167, N7160, N4629);
and AND4 (N7168, N7151, N1615, N600, N3894);
buf BUF1 (N7169, N7164);
not NOT1 (N7170, N7154);
buf BUF1 (N7171, N7170);
or OR4 (N7172, N7156, N6777, N4573, N6025);
not NOT1 (N7173, N7166);
xor XOR2 (N7174, N7165, N6588);
nor NOR2 (N7175, N7150, N3558);
buf BUF1 (N7176, N7161);
nand NAND3 (N7177, N7168, N3611, N6069);
or OR2 (N7178, N7167, N2522);
or OR3 (N7179, N7177, N3776, N1463);
or OR2 (N7180, N7159, N4760);
not NOT1 (N7181, N7174);
not NOT1 (N7182, N7179);
and AND4 (N7183, N7172, N2446, N4579, N2099);
nor NOR4 (N7184, N7176, N2817, N4082, N4419);
nor NOR3 (N7185, N7184, N480, N2475);
buf BUF1 (N7186, N7180);
nand NAND3 (N7187, N7186, N1540, N6892);
xor XOR2 (N7188, N7182, N2149);
not NOT1 (N7189, N7173);
nor NOR4 (N7190, N7181, N2141, N4469, N4236);
or OR4 (N7191, N7178, N1754, N57, N3158);
nand NAND4 (N7192, N7171, N3489, N3651, N3226);
nor NOR4 (N7193, N7191, N1035, N2032, N2439);
nand NAND3 (N7194, N7192, N3976, N4788);
or OR2 (N7195, N7187, N635);
buf BUF1 (N7196, N7175);
buf BUF1 (N7197, N7188);
nand NAND2 (N7198, N7197, N3061);
not NOT1 (N7199, N7194);
nand NAND2 (N7200, N7195, N3874);
not NOT1 (N7201, N7198);
or OR3 (N7202, N7169, N7125, N5907);
buf BUF1 (N7203, N7196);
and AND4 (N7204, N7199, N1362, N297, N2761);
or OR2 (N7205, N7185, N5428);
nor NOR4 (N7206, N7205, N2559, N417, N251);
buf BUF1 (N7207, N7203);
buf BUF1 (N7208, N7201);
or OR2 (N7209, N7206, N4967);
nand NAND3 (N7210, N7202, N4030, N5103);
buf BUF1 (N7211, N7193);
or OR4 (N7212, N7183, N5293, N5267, N2860);
nor NOR3 (N7213, N7212, N454, N1513);
buf BUF1 (N7214, N7213);
and AND2 (N7215, N7210, N6901);
buf BUF1 (N7216, N7214);
xor XOR2 (N7217, N7208, N3440);
nand NAND3 (N7218, N7209, N3681, N373);
buf BUF1 (N7219, N7190);
and AND3 (N7220, N7211, N5808, N1840);
nor NOR2 (N7221, N7220, N3359);
and AND3 (N7222, N7207, N5842, N6711);
xor XOR2 (N7223, N7204, N4956);
buf BUF1 (N7224, N7217);
buf BUF1 (N7225, N7223);
nor NOR3 (N7226, N7222, N2672, N6695);
not NOT1 (N7227, N7219);
nor NOR3 (N7228, N7225, N3954, N5645);
nand NAND2 (N7229, N7215, N4110);
buf BUF1 (N7230, N7227);
not NOT1 (N7231, N7189);
xor XOR2 (N7232, N7228, N1422);
or OR4 (N7233, N7216, N4953, N666, N5209);
buf BUF1 (N7234, N7231);
xor XOR2 (N7235, N7234, N5754);
and AND4 (N7236, N7226, N4246, N6393, N5159);
nor NOR2 (N7237, N7236, N6856);
and AND4 (N7238, N7232, N2153, N3142, N2433);
or OR2 (N7239, N7233, N4770);
nor NOR2 (N7240, N7229, N3422);
nor NOR2 (N7241, N7240, N3665);
nor NOR2 (N7242, N7238, N1304);
or OR3 (N7243, N7241, N4372, N6956);
nor NOR2 (N7244, N7239, N2147);
or OR3 (N7245, N7200, N5119, N2828);
buf BUF1 (N7246, N7242);
xor XOR2 (N7247, N7237, N5353);
nand NAND2 (N7248, N7218, N7200);
not NOT1 (N7249, N7244);
not NOT1 (N7250, N7221);
xor XOR2 (N7251, N7230, N4070);
and AND4 (N7252, N7251, N2475, N3319, N1350);
and AND2 (N7253, N7245, N3229);
xor XOR2 (N7254, N7249, N955);
and AND4 (N7255, N7253, N4280, N2099, N834);
xor XOR2 (N7256, N7255, N7084);
or OR4 (N7257, N7243, N2274, N4628, N6129);
not NOT1 (N7258, N7235);
nand NAND3 (N7259, N7247, N5679, N4870);
nand NAND2 (N7260, N7258, N6786);
nand NAND2 (N7261, N7252, N4121);
nand NAND2 (N7262, N7256, N1258);
or OR3 (N7263, N7261, N4844, N7201);
and AND2 (N7264, N7257, N5524);
buf BUF1 (N7265, N7248);
nand NAND2 (N7266, N7246, N5405);
or OR2 (N7267, N7266, N4855);
nor NOR3 (N7268, N7263, N1237, N2713);
nand NAND2 (N7269, N7254, N2934);
nor NOR4 (N7270, N7262, N1323, N315, N6263);
nor NOR4 (N7271, N7269, N2183, N5246, N4424);
or OR4 (N7272, N7271, N6942, N1519, N2058);
and AND3 (N7273, N7264, N7118, N4759);
xor XOR2 (N7274, N7268, N3304);
nor NOR3 (N7275, N7270, N6078, N862);
buf BUF1 (N7276, N7272);
or OR3 (N7277, N7259, N2830, N2803);
not NOT1 (N7278, N7276);
nor NOR4 (N7279, N7250, N3385, N3992, N3827);
and AND4 (N7280, N7224, N1443, N2814, N6259);
or OR3 (N7281, N7274, N4448, N7199);
or OR2 (N7282, N7277, N2194);
buf BUF1 (N7283, N7273);
nand NAND3 (N7284, N7265, N4745, N6015);
or OR4 (N7285, N7278, N114, N376, N2625);
and AND3 (N7286, N7260, N2394, N2542);
and AND2 (N7287, N7275, N4160);
buf BUF1 (N7288, N7283);
or OR4 (N7289, N7280, N2691, N2488, N574);
buf BUF1 (N7290, N7281);
nor NOR4 (N7291, N7290, N225, N2885, N1974);
nand NAND2 (N7292, N7267, N6170);
and AND4 (N7293, N7288, N940, N6700, N1559);
nand NAND4 (N7294, N7289, N7237, N1830, N2010);
xor XOR2 (N7295, N7279, N716);
buf BUF1 (N7296, N7286);
not NOT1 (N7297, N7291);
nor NOR2 (N7298, N7292, N4685);
buf BUF1 (N7299, N7284);
buf BUF1 (N7300, N7293);
or OR2 (N7301, N7300, N1860);
or OR4 (N7302, N7282, N1555, N1478, N4726);
buf BUF1 (N7303, N7298);
xor XOR2 (N7304, N7301, N3140);
nor NOR4 (N7305, N7297, N5699, N2980, N5558);
not NOT1 (N7306, N7302);
nor NOR4 (N7307, N7295, N5447, N361, N214);
buf BUF1 (N7308, N7304);
or OR2 (N7309, N7285, N3056);
not NOT1 (N7310, N7303);
not NOT1 (N7311, N7307);
and AND2 (N7312, N7294, N7141);
nor NOR2 (N7313, N7287, N1607);
not NOT1 (N7314, N7311);
xor XOR2 (N7315, N7308, N2835);
xor XOR2 (N7316, N7309, N3158);
nand NAND4 (N7317, N7312, N5454, N601, N6276);
or OR4 (N7318, N7317, N2921, N6640, N5256);
and AND2 (N7319, N7313, N3877);
or OR4 (N7320, N7299, N930, N2778, N1546);
and AND3 (N7321, N7320, N2855, N7317);
nand NAND3 (N7322, N7316, N1763, N2494);
xor XOR2 (N7323, N7319, N2658);
nor NOR3 (N7324, N7296, N5272, N1603);
not NOT1 (N7325, N7323);
and AND2 (N7326, N7305, N1191);
and AND4 (N7327, N7318, N4170, N315, N341);
buf BUF1 (N7328, N7310);
not NOT1 (N7329, N7306);
buf BUF1 (N7330, N7326);
or OR2 (N7331, N7321, N5997);
nand NAND3 (N7332, N7327, N4921, N801);
xor XOR2 (N7333, N7331, N3106);
buf BUF1 (N7334, N7328);
and AND2 (N7335, N7329, N2656);
nor NOR2 (N7336, N7332, N873);
nand NAND3 (N7337, N7322, N1497, N230);
not NOT1 (N7338, N7314);
or OR3 (N7339, N7338, N7062, N1710);
nor NOR2 (N7340, N7336, N6744);
buf BUF1 (N7341, N7315);
not NOT1 (N7342, N7341);
not NOT1 (N7343, N7334);
not NOT1 (N7344, N7337);
or OR4 (N7345, N7344, N2944, N2424, N236);
xor XOR2 (N7346, N7345, N7228);
and AND2 (N7347, N7339, N6902);
nor NOR2 (N7348, N7333, N864);
nand NAND4 (N7349, N7347, N6677, N3, N4832);
buf BUF1 (N7350, N7340);
or OR3 (N7351, N7348, N288, N4065);
or OR2 (N7352, N7349, N4007);
buf BUF1 (N7353, N7325);
buf BUF1 (N7354, N7353);
and AND4 (N7355, N7346, N3586, N6098, N503);
nor NOR3 (N7356, N7355, N2683, N112);
xor XOR2 (N7357, N7354, N6104);
nor NOR2 (N7358, N7357, N6685);
xor XOR2 (N7359, N7352, N5846);
xor XOR2 (N7360, N7358, N313);
nand NAND2 (N7361, N7330, N1533);
nor NOR4 (N7362, N7356, N6068, N1006, N7186);
nor NOR2 (N7363, N7350, N160);
nor NOR2 (N7364, N7363, N3371);
not NOT1 (N7365, N7359);
not NOT1 (N7366, N7362);
nor NOR2 (N7367, N7342, N1731);
or OR3 (N7368, N7366, N1540, N5539);
nor NOR4 (N7369, N7324, N59, N1854, N1559);
xor XOR2 (N7370, N7360, N3308);
nor NOR3 (N7371, N7343, N5090, N4201);
xor XOR2 (N7372, N7369, N3928);
xor XOR2 (N7373, N7368, N2144);
or OR2 (N7374, N7371, N4478);
xor XOR2 (N7375, N7374, N4128);
xor XOR2 (N7376, N7372, N3134);
and AND2 (N7377, N7361, N5189);
and AND3 (N7378, N7364, N367, N599);
xor XOR2 (N7379, N7367, N7086);
nand NAND2 (N7380, N7370, N6421);
nor NOR4 (N7381, N7376, N3080, N4817, N6297);
buf BUF1 (N7382, N7379);
xor XOR2 (N7383, N7335, N1748);
and AND4 (N7384, N7373, N3548, N2233, N4525);
nor NOR3 (N7385, N7380, N1886, N3296);
and AND3 (N7386, N7381, N5388, N3591);
xor XOR2 (N7387, N7375, N1521);
nand NAND4 (N7388, N7384, N755, N1080, N7314);
or OR2 (N7389, N7377, N2934);
xor XOR2 (N7390, N7382, N1394);
or OR4 (N7391, N7351, N6299, N7117, N2822);
not NOT1 (N7392, N7385);
or OR2 (N7393, N7389, N1411);
or OR4 (N7394, N7383, N1754, N229, N5576);
not NOT1 (N7395, N7387);
not NOT1 (N7396, N7393);
xor XOR2 (N7397, N7395, N6714);
not NOT1 (N7398, N7388);
not NOT1 (N7399, N7394);
or OR3 (N7400, N7386, N3563, N1812);
xor XOR2 (N7401, N7391, N6510);
or OR2 (N7402, N7397, N2044);
nand NAND3 (N7403, N7365, N3104, N3705);
and AND4 (N7404, N7403, N251, N248, N3034);
buf BUF1 (N7405, N7400);
buf BUF1 (N7406, N7402);
or OR2 (N7407, N7390, N6843);
or OR2 (N7408, N7404, N2503);
xor XOR2 (N7409, N7396, N3533);
and AND4 (N7410, N7408, N2792, N3119, N6529);
and AND2 (N7411, N7407, N988);
xor XOR2 (N7412, N7392, N5309);
or OR3 (N7413, N7411, N2980, N3836);
nand NAND2 (N7414, N7398, N2213);
nor NOR4 (N7415, N7406, N1174, N4260, N1766);
and AND4 (N7416, N7378, N1329, N2055, N1553);
buf BUF1 (N7417, N7399);
and AND4 (N7418, N7405, N4050, N3349, N6821);
nand NAND2 (N7419, N7415, N1749);
nor NOR3 (N7420, N7417, N1430, N129);
or OR2 (N7421, N7401, N7350);
xor XOR2 (N7422, N7418, N4173);
nand NAND4 (N7423, N7420, N4094, N1432, N6547);
nor NOR4 (N7424, N7423, N649, N6740, N3066);
not NOT1 (N7425, N7409);
nor NOR2 (N7426, N7425, N4871);
or OR2 (N7427, N7424, N2951);
not NOT1 (N7428, N7422);
or OR2 (N7429, N7416, N3037);
nand NAND3 (N7430, N7413, N2067, N5180);
xor XOR2 (N7431, N7421, N840);
or OR2 (N7432, N7431, N488);
and AND2 (N7433, N7426, N1110);
nand NAND4 (N7434, N7419, N798, N6794, N719);
nor NOR3 (N7435, N7433, N3983, N2211);
not NOT1 (N7436, N7412);
nor NOR3 (N7437, N7435, N2654, N2648);
and AND4 (N7438, N7427, N4833, N3290, N431);
nor NOR4 (N7439, N7429, N6653, N5820, N5002);
buf BUF1 (N7440, N7439);
buf BUF1 (N7441, N7428);
nand NAND3 (N7442, N7441, N3870, N4912);
buf BUF1 (N7443, N7414);
nor NOR2 (N7444, N7430, N3477);
nand NAND4 (N7445, N7434, N982, N325, N278);
and AND4 (N7446, N7432, N7027, N6010, N5679);
nand NAND4 (N7447, N7443, N2835, N1053, N3671);
and AND2 (N7448, N7444, N303);
buf BUF1 (N7449, N7442);
nor NOR4 (N7450, N7437, N1364, N4399, N5924);
and AND2 (N7451, N7438, N6967);
and AND2 (N7452, N7445, N1638);
nand NAND3 (N7453, N7449, N1931, N6615);
nand NAND3 (N7454, N7453, N6721, N5484);
nand NAND3 (N7455, N7447, N7154, N4257);
nand NAND2 (N7456, N7452, N6618);
or OR2 (N7457, N7450, N1792);
buf BUF1 (N7458, N7446);
xor XOR2 (N7459, N7457, N4496);
or OR2 (N7460, N7456, N1431);
not NOT1 (N7461, N7436);
nand NAND3 (N7462, N7461, N4024, N198);
xor XOR2 (N7463, N7440, N2359);
nor NOR3 (N7464, N7458, N2542, N7383);
not NOT1 (N7465, N7463);
or OR3 (N7466, N7455, N1702, N3530);
not NOT1 (N7467, N7465);
not NOT1 (N7468, N7448);
and AND3 (N7469, N7466, N7431, N4410);
not NOT1 (N7470, N7469);
xor XOR2 (N7471, N7459, N5053);
xor XOR2 (N7472, N7454, N3179);
and AND2 (N7473, N7462, N6947);
or OR4 (N7474, N7470, N5770, N673, N4981);
nor NOR2 (N7475, N7460, N6972);
nor NOR2 (N7476, N7474, N1698);
buf BUF1 (N7477, N7464);
and AND2 (N7478, N7451, N1289);
xor XOR2 (N7479, N7467, N2998);
buf BUF1 (N7480, N7472);
nand NAND3 (N7481, N7410, N7378, N4264);
nor NOR4 (N7482, N7478, N957, N6161, N6562);
nor NOR3 (N7483, N7481, N2924, N6736);
or OR3 (N7484, N7482, N365, N4109);
or OR2 (N7485, N7476, N5540);
nor NOR2 (N7486, N7485, N4700);
nand NAND2 (N7487, N7468, N348);
not NOT1 (N7488, N7479);
nand NAND4 (N7489, N7486, N4294, N5567, N1222);
nand NAND2 (N7490, N7477, N1192);
buf BUF1 (N7491, N7480);
not NOT1 (N7492, N7484);
nand NAND3 (N7493, N7483, N828, N4220);
not NOT1 (N7494, N7473);
xor XOR2 (N7495, N7493, N5488);
nand NAND2 (N7496, N7489, N4399);
xor XOR2 (N7497, N7475, N5675);
or OR2 (N7498, N7491, N98);
and AND2 (N7499, N7471, N3272);
not NOT1 (N7500, N7494);
not NOT1 (N7501, N7495);
or OR2 (N7502, N7492, N4194);
not NOT1 (N7503, N7500);
and AND4 (N7504, N7488, N4828, N6455, N5169);
not NOT1 (N7505, N7498);
or OR3 (N7506, N7490, N1178, N277);
and AND4 (N7507, N7502, N3952, N6998, N7169);
buf BUF1 (N7508, N7506);
xor XOR2 (N7509, N7497, N197);
xor XOR2 (N7510, N7505, N7472);
and AND3 (N7511, N7504, N7410, N6464);
buf BUF1 (N7512, N7508);
nor NOR3 (N7513, N7501, N51, N1875);
and AND2 (N7514, N7509, N5041);
xor XOR2 (N7515, N7511, N6968);
xor XOR2 (N7516, N7512, N1453);
and AND2 (N7517, N7515, N3694);
not NOT1 (N7518, N7503);
not NOT1 (N7519, N7507);
nand NAND2 (N7520, N7499, N2737);
nor NOR2 (N7521, N7510, N5479);
buf BUF1 (N7522, N7514);
buf BUF1 (N7523, N7496);
and AND4 (N7524, N7517, N5345, N5048, N1633);
not NOT1 (N7525, N7522);
nand NAND4 (N7526, N7487, N3488, N3882, N4540);
and AND2 (N7527, N7526, N5089);
xor XOR2 (N7528, N7525, N4117);
xor XOR2 (N7529, N7518, N368);
not NOT1 (N7530, N7527);
and AND2 (N7531, N7520, N1774);
nand NAND3 (N7532, N7531, N5967, N1524);
nor NOR4 (N7533, N7530, N646, N2276, N4441);
nand NAND3 (N7534, N7516, N553, N1748);
or OR4 (N7535, N7523, N3534, N6693, N2932);
or OR3 (N7536, N7533, N7388, N380);
and AND3 (N7537, N7532, N3880, N5646);
buf BUF1 (N7538, N7534);
or OR4 (N7539, N7538, N6087, N475, N1045);
not NOT1 (N7540, N7539);
nand NAND3 (N7541, N7521, N5293, N5363);
and AND4 (N7542, N7535, N5533, N4494, N5965);
not NOT1 (N7543, N7540);
nor NOR3 (N7544, N7537, N4342, N5535);
nand NAND4 (N7545, N7536, N513, N6493, N1680);
nand NAND3 (N7546, N7524, N5355, N5097);
nor NOR3 (N7547, N7542, N3199, N3182);
or OR4 (N7548, N7519, N3738, N5801, N3811);
nor NOR4 (N7549, N7548, N115, N1140, N504);
nand NAND3 (N7550, N7528, N5759, N4569);
nand NAND2 (N7551, N7546, N5632);
buf BUF1 (N7552, N7551);
not NOT1 (N7553, N7545);
or OR4 (N7554, N7541, N4013, N7351, N824);
and AND4 (N7555, N7529, N1218, N5277, N1104);
xor XOR2 (N7556, N7547, N4929);
nand NAND4 (N7557, N7513, N1825, N3276, N5581);
nand NAND2 (N7558, N7554, N2098);
buf BUF1 (N7559, N7549);
not NOT1 (N7560, N7553);
or OR2 (N7561, N7559, N6078);
nand NAND4 (N7562, N7555, N7175, N3150, N3711);
nand NAND3 (N7563, N7550, N1233, N2759);
xor XOR2 (N7564, N7560, N404);
xor XOR2 (N7565, N7544, N4214);
xor XOR2 (N7566, N7552, N3790);
xor XOR2 (N7567, N7562, N1633);
not NOT1 (N7568, N7557);
nand NAND2 (N7569, N7567, N7497);
xor XOR2 (N7570, N7568, N1026);
and AND4 (N7571, N7565, N3934, N4153, N2062);
buf BUF1 (N7572, N7556);
or OR3 (N7573, N7561, N3453, N3103);
xor XOR2 (N7574, N7563, N2332);
or OR4 (N7575, N7571, N5559, N1350, N6449);
buf BUF1 (N7576, N7572);
or OR2 (N7577, N7558, N6597);
xor XOR2 (N7578, N7576, N6992);
not NOT1 (N7579, N7543);
nand NAND2 (N7580, N7577, N4260);
not NOT1 (N7581, N7575);
not NOT1 (N7582, N7581);
nand NAND3 (N7583, N7574, N5933, N4194);
buf BUF1 (N7584, N7566);
buf BUF1 (N7585, N7570);
and AND4 (N7586, N7564, N6371, N5944, N1110);
nor NOR4 (N7587, N7585, N1136, N695, N7454);
and AND2 (N7588, N7569, N1114);
xor XOR2 (N7589, N7583, N4598);
nand NAND3 (N7590, N7573, N1113, N7280);
nand NAND4 (N7591, N7578, N3102, N5945, N1445);
and AND4 (N7592, N7582, N6857, N1782, N3249);
and AND3 (N7593, N7586, N7546, N4956);
and AND2 (N7594, N7590, N6752);
buf BUF1 (N7595, N7587);
and AND4 (N7596, N7588, N7421, N4898, N3785);
and AND2 (N7597, N7579, N4226);
nor NOR3 (N7598, N7596, N2543, N2863);
not NOT1 (N7599, N7592);
not NOT1 (N7600, N7593);
and AND4 (N7601, N7599, N1965, N5594, N4345);
buf BUF1 (N7602, N7601);
xor XOR2 (N7603, N7589, N2388);
buf BUF1 (N7604, N7595);
nor NOR3 (N7605, N7600, N6170, N993);
xor XOR2 (N7606, N7602, N4743);
and AND2 (N7607, N7603, N3836);
nand NAND3 (N7608, N7604, N6796, N3361);
nand NAND4 (N7609, N7584, N6890, N488, N4834);
not NOT1 (N7610, N7598);
and AND3 (N7611, N7606, N4352, N4935);
not NOT1 (N7612, N7597);
not NOT1 (N7613, N7611);
xor XOR2 (N7614, N7613, N2593);
xor XOR2 (N7615, N7610, N1927);
nor NOR3 (N7616, N7608, N6563, N5682);
nor NOR3 (N7617, N7615, N4774, N2352);
nor NOR2 (N7618, N7594, N5284);
buf BUF1 (N7619, N7612);
nor NOR3 (N7620, N7580, N2903, N1792);
buf BUF1 (N7621, N7614);
nand NAND4 (N7622, N7619, N5782, N793, N7011);
buf BUF1 (N7623, N7607);
xor XOR2 (N7624, N7623, N2468);
buf BUF1 (N7625, N7616);
nand NAND3 (N7626, N7621, N3286, N1220);
or OR3 (N7627, N7617, N7219, N7125);
or OR3 (N7628, N7618, N7392, N2441);
nor NOR3 (N7629, N7609, N875, N14);
and AND4 (N7630, N7620, N5561, N3238, N640);
or OR4 (N7631, N7626, N5402, N6164, N7495);
nand NAND2 (N7632, N7631, N5260);
and AND3 (N7633, N7630, N1253, N3112);
not NOT1 (N7634, N7622);
buf BUF1 (N7635, N7591);
nor NOR2 (N7636, N7633, N7320);
not NOT1 (N7637, N7634);
buf BUF1 (N7638, N7629);
nand NAND2 (N7639, N7638, N5224);
nor NOR3 (N7640, N7636, N6857, N4734);
buf BUF1 (N7641, N7624);
nand NAND4 (N7642, N7637, N4558, N927, N4673);
nand NAND4 (N7643, N7625, N7468, N5960, N6761);
not NOT1 (N7644, N7643);
and AND4 (N7645, N7641, N6535, N682, N5611);
not NOT1 (N7646, N7644);
and AND3 (N7647, N7639, N44, N2410);
and AND4 (N7648, N7647, N5264, N2398, N975);
or OR4 (N7649, N7632, N2687, N7117, N2313);
nand NAND3 (N7650, N7605, N5609, N6229);
xor XOR2 (N7651, N7635, N5942);
or OR4 (N7652, N7640, N6082, N921, N826);
buf BUF1 (N7653, N7646);
nor NOR2 (N7654, N7648, N3992);
nor NOR4 (N7655, N7642, N2436, N7488, N3726);
nor NOR4 (N7656, N7649, N1250, N1854, N3233);
buf BUF1 (N7657, N7652);
not NOT1 (N7658, N7653);
xor XOR2 (N7659, N7658, N793);
nor NOR3 (N7660, N7656, N2419, N338);
xor XOR2 (N7661, N7654, N190);
not NOT1 (N7662, N7655);
and AND2 (N7663, N7657, N7507);
and AND3 (N7664, N7627, N3542, N925);
or OR4 (N7665, N7651, N5313, N4602, N5478);
xor XOR2 (N7666, N7665, N1481);
xor XOR2 (N7667, N7664, N3798);
xor XOR2 (N7668, N7659, N7276);
nand NAND3 (N7669, N7661, N4561, N195);
nor NOR2 (N7670, N7669, N5109);
buf BUF1 (N7671, N7668);
not NOT1 (N7672, N7662);
and AND3 (N7673, N7670, N1193, N727);
or OR2 (N7674, N7663, N3912);
not NOT1 (N7675, N7674);
and AND4 (N7676, N7650, N861, N2738, N5459);
nand NAND3 (N7677, N7671, N5787, N5357);
nor NOR4 (N7678, N7666, N7672, N4617, N4255);
not NOT1 (N7679, N671);
buf BUF1 (N7680, N7660);
xor XOR2 (N7681, N7673, N3952);
nand NAND2 (N7682, N7667, N6497);
and AND2 (N7683, N7676, N2790);
xor XOR2 (N7684, N7683, N2393);
nand NAND2 (N7685, N7675, N6423);
buf BUF1 (N7686, N7685);
xor XOR2 (N7687, N7678, N3909);
and AND4 (N7688, N7680, N1083, N3430, N2691);
and AND2 (N7689, N7681, N3224);
not NOT1 (N7690, N7628);
xor XOR2 (N7691, N7689, N6908);
xor XOR2 (N7692, N7645, N1253);
xor XOR2 (N7693, N7692, N2254);
xor XOR2 (N7694, N7690, N7052);
not NOT1 (N7695, N7693);
buf BUF1 (N7696, N7691);
not NOT1 (N7697, N7695);
or OR3 (N7698, N7686, N3900, N3716);
nand NAND2 (N7699, N7688, N1888);
buf BUF1 (N7700, N7679);
and AND4 (N7701, N7697, N6420, N4059, N3308);
or OR4 (N7702, N7684, N5633, N896, N4233);
not NOT1 (N7703, N7682);
and AND3 (N7704, N7702, N3431, N6301);
buf BUF1 (N7705, N7701);
or OR2 (N7706, N7677, N6068);
nand NAND2 (N7707, N7698, N6657);
buf BUF1 (N7708, N7705);
and AND3 (N7709, N7707, N5235, N7558);
or OR2 (N7710, N7699, N2846);
xor XOR2 (N7711, N7709, N5767);
nand NAND4 (N7712, N7694, N7683, N5167, N1150);
and AND3 (N7713, N7706, N6994, N3144);
xor XOR2 (N7714, N7710, N2029);
or OR2 (N7715, N7714, N4935);
not NOT1 (N7716, N7711);
or OR4 (N7717, N7716, N1773, N5195, N1756);
and AND2 (N7718, N7717, N3859);
nand NAND2 (N7719, N7712, N1635);
not NOT1 (N7720, N7708);
not NOT1 (N7721, N7703);
and AND3 (N7722, N7715, N27, N980);
xor XOR2 (N7723, N7721, N4619);
not NOT1 (N7724, N7723);
buf BUF1 (N7725, N7719);
nand NAND4 (N7726, N7696, N902, N5336, N7075);
nand NAND2 (N7727, N7724, N1976);
xor XOR2 (N7728, N7718, N1422);
or OR2 (N7729, N7728, N5721);
nor NOR3 (N7730, N7726, N6840, N236);
nand NAND3 (N7731, N7700, N4171, N243);
buf BUF1 (N7732, N7687);
not NOT1 (N7733, N7727);
nor NOR2 (N7734, N7725, N5079);
or OR2 (N7735, N7730, N651);
buf BUF1 (N7736, N7729);
nand NAND3 (N7737, N7713, N3527, N7065);
nor NOR2 (N7738, N7732, N4717);
nor NOR2 (N7739, N7720, N5898);
nand NAND2 (N7740, N7737, N565);
xor XOR2 (N7741, N7740, N1995);
xor XOR2 (N7742, N7739, N762);
buf BUF1 (N7743, N7735);
not NOT1 (N7744, N7733);
nand NAND2 (N7745, N7741, N5190);
not NOT1 (N7746, N7738);
or OR2 (N7747, N7736, N6627);
buf BUF1 (N7748, N7744);
or OR2 (N7749, N7745, N4512);
or OR4 (N7750, N7731, N1177, N2378, N7301);
and AND3 (N7751, N7722, N5231, N3494);
not NOT1 (N7752, N7749);
and AND4 (N7753, N7704, N1711, N6029, N308);
or OR2 (N7754, N7734, N1651);
buf BUF1 (N7755, N7753);
nor NOR3 (N7756, N7746, N7397, N5782);
buf BUF1 (N7757, N7748);
buf BUF1 (N7758, N7751);
buf BUF1 (N7759, N7747);
nand NAND4 (N7760, N7750, N1883, N2382, N2198);
nor NOR4 (N7761, N7759, N5051, N2408, N6674);
xor XOR2 (N7762, N7760, N4332);
xor XOR2 (N7763, N7755, N435);
or OR2 (N7764, N7752, N6707);
nor NOR3 (N7765, N7758, N5164, N813);
buf BUF1 (N7766, N7763);
not NOT1 (N7767, N7757);
buf BUF1 (N7768, N7754);
not NOT1 (N7769, N7768);
not NOT1 (N7770, N7769);
and AND2 (N7771, N7765, N2713);
and AND3 (N7772, N7766, N6273, N5645);
buf BUF1 (N7773, N7772);
xor XOR2 (N7774, N7771, N2090);
and AND2 (N7775, N7770, N6458);
and AND3 (N7776, N7773, N1287, N3954);
not NOT1 (N7777, N7776);
and AND3 (N7778, N7774, N788, N406);
nand NAND2 (N7779, N7767, N4898);
and AND4 (N7780, N7775, N403, N115, N634);
and AND4 (N7781, N7778, N908, N207, N1436);
or OR2 (N7782, N7780, N6372);
and AND4 (N7783, N7761, N4922, N5664, N3589);
nand NAND2 (N7784, N7782, N6759);
or OR2 (N7785, N7783, N2589);
buf BUF1 (N7786, N7781);
and AND2 (N7787, N7785, N3355);
buf BUF1 (N7788, N7764);
buf BUF1 (N7789, N7787);
not NOT1 (N7790, N7777);
xor XOR2 (N7791, N7789, N3216);
or OR2 (N7792, N7786, N3073);
xor XOR2 (N7793, N7784, N155);
nor NOR2 (N7794, N7791, N2681);
or OR4 (N7795, N7790, N7076, N4237, N4649);
buf BUF1 (N7796, N7779);
not NOT1 (N7797, N7795);
nand NAND3 (N7798, N7762, N4861, N2816);
or OR2 (N7799, N7743, N6899);
xor XOR2 (N7800, N7799, N4213);
buf BUF1 (N7801, N7793);
and AND2 (N7802, N7788, N4914);
or OR3 (N7803, N7756, N4536, N6619);
nor NOR4 (N7804, N7797, N4227, N1612, N5410);
not NOT1 (N7805, N7804);
buf BUF1 (N7806, N7805);
nor NOR2 (N7807, N7803, N976);
nand NAND2 (N7808, N7801, N3937);
buf BUF1 (N7809, N7794);
xor XOR2 (N7810, N7802, N6336);
nor NOR3 (N7811, N7800, N2667, N5698);
xor XOR2 (N7812, N7807, N5031);
nor NOR2 (N7813, N7742, N327);
not NOT1 (N7814, N7796);
xor XOR2 (N7815, N7814, N3650);
and AND3 (N7816, N7792, N2535, N517);
buf BUF1 (N7817, N7811);
nor NOR4 (N7818, N7816, N4385, N4923, N7690);
buf BUF1 (N7819, N7812);
and AND4 (N7820, N7818, N4493, N6582, N4768);
nor NOR2 (N7821, N7808, N3458);
not NOT1 (N7822, N7817);
and AND3 (N7823, N7822, N1535, N6596);
xor XOR2 (N7824, N7798, N5849);
buf BUF1 (N7825, N7815);
nand NAND2 (N7826, N7806, N4652);
nor NOR4 (N7827, N7821, N5879, N1988, N935);
or OR4 (N7828, N7824, N1653, N1491, N1872);
buf BUF1 (N7829, N7810);
xor XOR2 (N7830, N7819, N4338);
not NOT1 (N7831, N7830);
or OR3 (N7832, N7820, N1939, N4809);
xor XOR2 (N7833, N7826, N4934);
buf BUF1 (N7834, N7813);
not NOT1 (N7835, N7832);
not NOT1 (N7836, N7825);
or OR4 (N7837, N7833, N2927, N7473, N2201);
nor NOR2 (N7838, N7835, N5583);
not NOT1 (N7839, N7831);
or OR3 (N7840, N7827, N4754, N2619);
and AND2 (N7841, N7839, N4728);
nand NAND3 (N7842, N7840, N3897, N3146);
nand NAND4 (N7843, N7838, N4913, N6568, N823);
nand NAND3 (N7844, N7842, N5941, N6237);
nor NOR2 (N7845, N7844, N5827);
or OR4 (N7846, N7823, N6574, N237, N3591);
buf BUF1 (N7847, N7828);
nand NAND3 (N7848, N7809, N7019, N1328);
not NOT1 (N7849, N7837);
buf BUF1 (N7850, N7829);
nor NOR4 (N7851, N7834, N5555, N3663, N18);
xor XOR2 (N7852, N7841, N2071);
nor NOR2 (N7853, N7849, N2846);
xor XOR2 (N7854, N7845, N1553);
nand NAND3 (N7855, N7836, N3889, N6716);
not NOT1 (N7856, N7851);
buf BUF1 (N7857, N7846);
xor XOR2 (N7858, N7856, N3551);
not NOT1 (N7859, N7858);
and AND4 (N7860, N7847, N3921, N5898, N6625);
nor NOR2 (N7861, N7854, N3171);
xor XOR2 (N7862, N7843, N7689);
and AND3 (N7863, N7860, N4744, N303);
nor NOR4 (N7864, N7861, N4806, N711, N1069);
xor XOR2 (N7865, N7850, N6898);
and AND3 (N7866, N7863, N3126, N5819);
xor XOR2 (N7867, N7859, N2409);
or OR2 (N7868, N7852, N5812);
nor NOR2 (N7869, N7866, N5449);
not NOT1 (N7870, N7865);
buf BUF1 (N7871, N7867);
xor XOR2 (N7872, N7855, N3428);
or OR3 (N7873, N7862, N6309, N5226);
buf BUF1 (N7874, N7864);
nor NOR3 (N7875, N7869, N5641, N5733);
nand NAND2 (N7876, N7853, N6198);
nor NOR3 (N7877, N7872, N1951, N1553);
nor NOR4 (N7878, N7868, N775, N1192, N1856);
and AND4 (N7879, N7848, N4225, N2094, N1123);
nor NOR4 (N7880, N7871, N3750, N7198, N5245);
xor XOR2 (N7881, N7877, N4614);
nand NAND2 (N7882, N7880, N2312);
or OR2 (N7883, N7874, N4122);
or OR2 (N7884, N7883, N5381);
buf BUF1 (N7885, N7870);
or OR2 (N7886, N7875, N3886);
buf BUF1 (N7887, N7879);
not NOT1 (N7888, N7878);
nor NOR2 (N7889, N7887, N774);
not NOT1 (N7890, N7882);
nor NOR2 (N7891, N7889, N7887);
nor NOR2 (N7892, N7886, N2244);
xor XOR2 (N7893, N7884, N2395);
xor XOR2 (N7894, N7885, N3030);
buf BUF1 (N7895, N7892);
xor XOR2 (N7896, N7890, N6185);
and AND2 (N7897, N7857, N1514);
buf BUF1 (N7898, N7876);
not NOT1 (N7899, N7897);
nor NOR2 (N7900, N7888, N2629);
or OR3 (N7901, N7896, N4421, N5514);
not NOT1 (N7902, N7894);
and AND3 (N7903, N7901, N3582, N2070);
not NOT1 (N7904, N7891);
nand NAND4 (N7905, N7904, N7490, N643, N2127);
and AND2 (N7906, N7873, N6542);
not NOT1 (N7907, N7900);
not NOT1 (N7908, N7907);
nor NOR3 (N7909, N7881, N6978, N2732);
buf BUF1 (N7910, N7909);
nand NAND4 (N7911, N7893, N5396, N5652, N6374);
buf BUF1 (N7912, N7899);
buf BUF1 (N7913, N7905);
xor XOR2 (N7914, N7913, N714);
xor XOR2 (N7915, N7906, N6157);
xor XOR2 (N7916, N7910, N6646);
and AND3 (N7917, N7898, N6616, N239);
not NOT1 (N7918, N7903);
not NOT1 (N7919, N7916);
nand NAND4 (N7920, N7895, N7896, N7830, N5021);
or OR3 (N7921, N7908, N581, N5658);
xor XOR2 (N7922, N7917, N3938);
nand NAND3 (N7923, N7902, N6160, N5369);
not NOT1 (N7924, N7912);
xor XOR2 (N7925, N7914, N4766);
or OR3 (N7926, N7918, N4649, N944);
xor XOR2 (N7927, N7924, N32);
nand NAND4 (N7928, N7919, N1898, N3545, N4517);
and AND3 (N7929, N7926, N974, N3051);
xor XOR2 (N7930, N7925, N3678);
not NOT1 (N7931, N7922);
not NOT1 (N7932, N7927);
nand NAND2 (N7933, N7931, N2071);
nand NAND4 (N7934, N7911, N560, N6518, N7441);
nand NAND2 (N7935, N7932, N2506);
buf BUF1 (N7936, N7920);
or OR2 (N7937, N7915, N6330);
and AND2 (N7938, N7934, N909);
buf BUF1 (N7939, N7930);
or OR3 (N7940, N7939, N1206, N5438);
nor NOR3 (N7941, N7929, N1297, N1350);
and AND4 (N7942, N7935, N3458, N4888, N2213);
nand NAND3 (N7943, N7942, N4958, N5136);
buf BUF1 (N7944, N7928);
nor NOR3 (N7945, N7938, N2541, N6391);
and AND2 (N7946, N7944, N4136);
xor XOR2 (N7947, N7941, N3304);
nand NAND4 (N7948, N7940, N1795, N4305, N5628);
xor XOR2 (N7949, N7946, N7025);
and AND2 (N7950, N7947, N3837);
and AND2 (N7951, N7933, N4738);
buf BUF1 (N7952, N7923);
nand NAND3 (N7953, N7948, N2577, N1388);
buf BUF1 (N7954, N7937);
or OR4 (N7955, N7951, N6414, N6780, N5);
or OR2 (N7956, N7955, N5959);
nor NOR3 (N7957, N7945, N2584, N124);
buf BUF1 (N7958, N7953);
and AND2 (N7959, N7950, N3518);
xor XOR2 (N7960, N7921, N3448);
or OR4 (N7961, N7960, N6974, N6966, N4257);
not NOT1 (N7962, N7959);
not NOT1 (N7963, N7952);
nand NAND3 (N7964, N7949, N4752, N5664);
and AND3 (N7965, N7954, N36, N4634);
xor XOR2 (N7966, N7956, N3719);
or OR4 (N7967, N7964, N1756, N3650, N711);
nor NOR3 (N7968, N7936, N5236, N7501);
nand NAND2 (N7969, N7962, N1863);
nor NOR4 (N7970, N7966, N5451, N4094, N3229);
and AND3 (N7971, N7967, N4703, N6826);
or OR4 (N7972, N7971, N4317, N3038, N3408);
buf BUF1 (N7973, N7958);
nor NOR4 (N7974, N7972, N4193, N7444, N6520);
nand NAND3 (N7975, N7974, N1852, N7223);
nand NAND2 (N7976, N7957, N6560);
xor XOR2 (N7977, N7961, N6528);
xor XOR2 (N7978, N7968, N5513);
or OR2 (N7979, N7973, N4697);
nand NAND2 (N7980, N7965, N6251);
and AND3 (N7981, N7970, N3896, N6546);
xor XOR2 (N7982, N7978, N3996);
and AND3 (N7983, N7943, N1691, N6975);
xor XOR2 (N7984, N7980, N3119);
buf BUF1 (N7985, N7981);
xor XOR2 (N7986, N7985, N7274);
xor XOR2 (N7987, N7979, N7915);
xor XOR2 (N7988, N7983, N3941);
and AND3 (N7989, N7988, N5787, N2604);
not NOT1 (N7990, N7984);
and AND4 (N7991, N7975, N1884, N2714, N2025);
not NOT1 (N7992, N7982);
or OR3 (N7993, N7989, N6055, N4324);
not NOT1 (N7994, N7992);
not NOT1 (N7995, N7986);
buf BUF1 (N7996, N7994);
xor XOR2 (N7997, N7993, N1752);
nor NOR4 (N7998, N7963, N3576, N6785, N5693);
or OR2 (N7999, N7969, N6038);
nand NAND4 (N8000, N7990, N5539, N1917, N4454);
nor NOR2 (N8001, N7996, N4264);
buf BUF1 (N8002, N8000);
nand NAND2 (N8003, N8001, N5567);
xor XOR2 (N8004, N7977, N2260);
buf BUF1 (N8005, N7998);
buf BUF1 (N8006, N8002);
xor XOR2 (N8007, N8005, N509);
nand NAND3 (N8008, N8004, N6189, N5833);
not NOT1 (N8009, N8007);
or OR3 (N8010, N8003, N4970, N2034);
or OR4 (N8011, N7991, N5774, N7783, N3521);
nor NOR2 (N8012, N7987, N7382);
nand NAND4 (N8013, N8006, N4973, N449, N6073);
or OR3 (N8014, N8011, N6848, N5891);
buf BUF1 (N8015, N8013);
and AND4 (N8016, N7976, N2327, N5281, N989);
nor NOR2 (N8017, N7995, N3877);
nor NOR2 (N8018, N8016, N5115);
nor NOR2 (N8019, N8008, N1405);
and AND4 (N8020, N8015, N4625, N6581, N1424);
or OR4 (N8021, N8018, N3067, N3765, N5802);
xor XOR2 (N8022, N8019, N5268);
nand NAND2 (N8023, N8022, N3504);
not NOT1 (N8024, N8017);
nor NOR4 (N8025, N8023, N4095, N7991, N5756);
buf BUF1 (N8026, N8024);
not NOT1 (N8027, N8021);
and AND4 (N8028, N8020, N363, N6997, N6776);
nand NAND3 (N8029, N8009, N2178, N6301);
and AND3 (N8030, N8010, N663, N3409);
nand NAND2 (N8031, N8025, N5951);
xor XOR2 (N8032, N8029, N2869);
or OR4 (N8033, N8026, N2693, N4481, N1266);
nand NAND4 (N8034, N8033, N2623, N5929, N2850);
or OR2 (N8035, N8027, N8025);
not NOT1 (N8036, N8035);
buf BUF1 (N8037, N8014);
not NOT1 (N8038, N8012);
nor NOR2 (N8039, N8032, N3197);
and AND3 (N8040, N8028, N1039, N4579);
buf BUF1 (N8041, N8040);
xor XOR2 (N8042, N8037, N6115);
not NOT1 (N8043, N8041);
not NOT1 (N8044, N8034);
xor XOR2 (N8045, N8036, N7975);
and AND2 (N8046, N8043, N3623);
not NOT1 (N8047, N8039);
not NOT1 (N8048, N8046);
nor NOR3 (N8049, N8044, N1091, N1783);
nand NAND3 (N8050, N8031, N6361, N3899);
not NOT1 (N8051, N8038);
buf BUF1 (N8052, N8047);
buf BUF1 (N8053, N7999);
buf BUF1 (N8054, N8049);
xor XOR2 (N8055, N8042, N150);
and AND2 (N8056, N8055, N681);
not NOT1 (N8057, N8045);
and AND3 (N8058, N8052, N6299, N3624);
nand NAND3 (N8059, N7997, N5689, N190);
buf BUF1 (N8060, N8051);
xor XOR2 (N8061, N8056, N3897);
nor NOR2 (N8062, N8053, N3161);
nand NAND3 (N8063, N8061, N2246, N1957);
and AND2 (N8064, N8058, N2206);
and AND2 (N8065, N8057, N2009);
nand NAND4 (N8066, N8054, N2047, N196, N1598);
buf BUF1 (N8067, N8030);
xor XOR2 (N8068, N8060, N5193);
buf BUF1 (N8069, N8050);
nor NOR3 (N8070, N8066, N7355, N6811);
buf BUF1 (N8071, N8064);
not NOT1 (N8072, N8059);
or OR4 (N8073, N8065, N4765, N2136, N388);
or OR3 (N8074, N8062, N5551, N8018);
nand NAND3 (N8075, N8072, N1188, N5099);
not NOT1 (N8076, N8048);
buf BUF1 (N8077, N8075);
nand NAND3 (N8078, N8076, N2443, N7463);
nand NAND4 (N8079, N8074, N1998, N4170, N245);
not NOT1 (N8080, N8073);
nand NAND2 (N8081, N8071, N6961);
nand NAND3 (N8082, N8079, N6088, N7412);
xor XOR2 (N8083, N8069, N1848);
nor NOR3 (N8084, N8063, N4227, N3006);
buf BUF1 (N8085, N8070);
nand NAND4 (N8086, N8068, N5782, N1679, N2841);
xor XOR2 (N8087, N8085, N2708);
and AND4 (N8088, N8082, N5738, N6271, N5094);
nand NAND2 (N8089, N8067, N6549);
or OR3 (N8090, N8078, N752, N1806);
buf BUF1 (N8091, N8089);
nand NAND4 (N8092, N8084, N5154, N6149, N5623);
not NOT1 (N8093, N8077);
nor NOR3 (N8094, N8088, N1241, N371);
not NOT1 (N8095, N8083);
xor XOR2 (N8096, N8081, N2331);
xor XOR2 (N8097, N8080, N1607);
xor XOR2 (N8098, N8090, N1184);
or OR4 (N8099, N8092, N1911, N2379, N4971);
nand NAND3 (N8100, N8095, N7761, N336);
or OR4 (N8101, N8091, N4403, N2032, N6499);
xor XOR2 (N8102, N8098, N7423);
and AND2 (N8103, N8102, N5218);
xor XOR2 (N8104, N8096, N1503);
nor NOR3 (N8105, N8094, N7130, N5444);
and AND2 (N8106, N8093, N4460);
nand NAND3 (N8107, N8105, N213, N5485);
nand NAND4 (N8108, N8100, N7430, N1512, N7233);
nand NAND4 (N8109, N8087, N5639, N234, N5186);
buf BUF1 (N8110, N8103);
buf BUF1 (N8111, N8109);
nor NOR2 (N8112, N8110, N7956);
buf BUF1 (N8113, N8106);
and AND2 (N8114, N8111, N1661);
not NOT1 (N8115, N8097);
nand NAND3 (N8116, N8104, N4311, N2512);
nor NOR3 (N8117, N8114, N5000, N565);
and AND3 (N8118, N8108, N1787, N2561);
nand NAND4 (N8119, N8086, N7901, N391, N5864);
not NOT1 (N8120, N8119);
nor NOR4 (N8121, N8107, N7014, N4475, N1499);
nor NOR3 (N8122, N8116, N61, N7038);
not NOT1 (N8123, N8122);
nand NAND2 (N8124, N8120, N5409);
and AND3 (N8125, N8101, N3428, N621);
not NOT1 (N8126, N8113);
buf BUF1 (N8127, N8112);
or OR3 (N8128, N8123, N5141, N2034);
nor NOR4 (N8129, N8118, N4026, N7031, N6423);
and AND3 (N8130, N8127, N7600, N3725);
or OR2 (N8131, N8126, N2773);
and AND4 (N8132, N8121, N4319, N2066, N2974);
nand NAND3 (N8133, N8124, N5489, N3368);
nand NAND4 (N8134, N8131, N5947, N6267, N4404);
xor XOR2 (N8135, N8129, N3185);
nand NAND2 (N8136, N8125, N4191);
buf BUF1 (N8137, N8099);
nand NAND4 (N8138, N8130, N6727, N4311, N3183);
nor NOR2 (N8139, N8138, N3717);
or OR3 (N8140, N8135, N1378, N3998);
nand NAND2 (N8141, N8115, N310);
nor NOR2 (N8142, N8134, N1879);
nor NOR2 (N8143, N8141, N4352);
buf BUF1 (N8144, N8136);
not NOT1 (N8145, N8143);
xor XOR2 (N8146, N8144, N2990);
buf BUF1 (N8147, N8145);
xor XOR2 (N8148, N8140, N4256);
and AND3 (N8149, N8148, N6884, N3798);
or OR2 (N8150, N8137, N58);
xor XOR2 (N8151, N8142, N4600);
or OR4 (N8152, N8117, N2062, N1258, N5230);
buf BUF1 (N8153, N8150);
and AND2 (N8154, N8152, N2227);
xor XOR2 (N8155, N8147, N3025);
not NOT1 (N8156, N8153);
not NOT1 (N8157, N8154);
not NOT1 (N8158, N8157);
not NOT1 (N8159, N8128);
nand NAND4 (N8160, N8155, N2926, N7532, N70);
nor NOR3 (N8161, N8151, N6695, N2410);
or OR3 (N8162, N8132, N8108, N2);
or OR2 (N8163, N8162, N1686);
not NOT1 (N8164, N8158);
nor NOR3 (N8165, N8146, N7096, N1385);
nand NAND3 (N8166, N8161, N3109, N6132);
nor NOR3 (N8167, N8163, N193, N2074);
and AND4 (N8168, N8159, N6180, N4936, N5864);
xor XOR2 (N8169, N8139, N5249);
not NOT1 (N8170, N8168);
and AND4 (N8171, N8165, N6172, N8160, N2092);
nand NAND3 (N8172, N8009, N7924, N1321);
buf BUF1 (N8173, N8133);
nor NOR4 (N8174, N8166, N3194, N2349, N886);
not NOT1 (N8175, N8167);
nand NAND3 (N8176, N8172, N24, N3051);
nor NOR4 (N8177, N8164, N4748, N2071, N5652);
nand NAND3 (N8178, N8174, N1665, N6572);
not NOT1 (N8179, N8156);
buf BUF1 (N8180, N8176);
xor XOR2 (N8181, N8173, N4646);
buf BUF1 (N8182, N8149);
buf BUF1 (N8183, N8178);
and AND3 (N8184, N8182, N749, N3681);
not NOT1 (N8185, N8170);
and AND4 (N8186, N8175, N3158, N7559, N6118);
buf BUF1 (N8187, N8184);
xor XOR2 (N8188, N8183, N5224);
and AND4 (N8189, N8185, N2181, N6578, N512);
nand NAND4 (N8190, N8189, N4782, N3165, N1043);
not NOT1 (N8191, N8171);
buf BUF1 (N8192, N8181);
xor XOR2 (N8193, N8169, N6574);
nor NOR2 (N8194, N8179, N6178);
and AND4 (N8195, N8180, N5847, N1556, N1311);
buf BUF1 (N8196, N8188);
xor XOR2 (N8197, N8192, N5216);
and AND2 (N8198, N8195, N2448);
not NOT1 (N8199, N8187);
buf BUF1 (N8200, N8186);
nor NOR2 (N8201, N8190, N953);
and AND4 (N8202, N8177, N580, N3221, N1967);
or OR2 (N8203, N8202, N5455);
xor XOR2 (N8204, N8201, N2164);
and AND2 (N8205, N8199, N4822);
nor NOR4 (N8206, N8193, N3913, N7665, N1401);
and AND4 (N8207, N8194, N7064, N1586, N4146);
nand NAND4 (N8208, N8200, N6938, N8003, N7217);
xor XOR2 (N8209, N8205, N2389);
xor XOR2 (N8210, N8197, N2957);
buf BUF1 (N8211, N8198);
and AND3 (N8212, N8209, N754, N2023);
not NOT1 (N8213, N8203);
and AND4 (N8214, N8213, N1025, N3661, N7425);
nand NAND2 (N8215, N8191, N7789);
or OR4 (N8216, N8210, N5180, N606, N2819);
not NOT1 (N8217, N8211);
nor NOR3 (N8218, N8217, N7538, N6435);
xor XOR2 (N8219, N8218, N834);
nor NOR3 (N8220, N8206, N1713, N7202);
xor XOR2 (N8221, N8219, N1258);
xor XOR2 (N8222, N8204, N4238);
and AND2 (N8223, N8216, N66);
not NOT1 (N8224, N8196);
and AND4 (N8225, N8220, N7291, N1421, N201);
and AND2 (N8226, N8208, N139);
buf BUF1 (N8227, N8225);
xor XOR2 (N8228, N8227, N2547);
nand NAND2 (N8229, N8226, N7701);
not NOT1 (N8230, N8215);
not NOT1 (N8231, N8229);
xor XOR2 (N8232, N8214, N5345);
nand NAND3 (N8233, N8224, N6509, N7290);
or OR3 (N8234, N8221, N158, N6423);
nand NAND3 (N8235, N8231, N1283, N1925);
nand NAND4 (N8236, N8223, N1139, N6846, N8045);
not NOT1 (N8237, N8207);
and AND4 (N8238, N8222, N2180, N2450, N7458);
nand NAND3 (N8239, N8237, N5335, N7682);
not NOT1 (N8240, N8232);
nand NAND3 (N8241, N8239, N6647, N4566);
xor XOR2 (N8242, N8236, N5183);
nor NOR2 (N8243, N8233, N7809);
xor XOR2 (N8244, N8212, N3100);
nand NAND2 (N8245, N8238, N1752);
xor XOR2 (N8246, N8241, N6319);
not NOT1 (N8247, N8240);
or OR3 (N8248, N8242, N5019, N6725);
nor NOR4 (N8249, N8246, N78, N3590, N2364);
nand NAND4 (N8250, N8245, N3700, N3807, N8225);
nor NOR3 (N8251, N8228, N4815, N6103);
nor NOR3 (N8252, N8234, N5555, N4091);
and AND2 (N8253, N8247, N6120);
or OR4 (N8254, N8248, N1034, N6541, N4926);
buf BUF1 (N8255, N8252);
xor XOR2 (N8256, N8250, N3804);
nor NOR4 (N8257, N8230, N5867, N8234, N75);
nand NAND4 (N8258, N8254, N976, N128, N5189);
nor NOR2 (N8259, N8257, N5043);
nand NAND4 (N8260, N8244, N3882, N1532, N7787);
xor XOR2 (N8261, N8258, N7317);
nor NOR3 (N8262, N8235, N2074, N4568);
not NOT1 (N8263, N8260);
nand NAND4 (N8264, N8256, N7536, N4330, N2620);
xor XOR2 (N8265, N8251, N803);
and AND2 (N8266, N8261, N6327);
xor XOR2 (N8267, N8243, N327);
buf BUF1 (N8268, N8262);
or OR4 (N8269, N8266, N8135, N2819, N1966);
xor XOR2 (N8270, N8268, N4787);
not NOT1 (N8271, N8255);
or OR2 (N8272, N8264, N2117);
or OR2 (N8273, N8271, N4273);
or OR3 (N8274, N8249, N249, N1480);
nor NOR2 (N8275, N8263, N3538);
or OR3 (N8276, N8267, N5471, N1095);
and AND3 (N8277, N8273, N4577, N3176);
nand NAND2 (N8278, N8253, N3392);
buf BUF1 (N8279, N8276);
buf BUF1 (N8280, N8275);
not NOT1 (N8281, N8280);
and AND3 (N8282, N8278, N7441, N4906);
not NOT1 (N8283, N8272);
nor NOR2 (N8284, N8265, N82);
xor XOR2 (N8285, N8259, N981);
xor XOR2 (N8286, N8269, N490);
not NOT1 (N8287, N8277);
buf BUF1 (N8288, N8285);
or OR2 (N8289, N8281, N2561);
buf BUF1 (N8290, N8274);
or OR3 (N8291, N8270, N953, N3918);
and AND4 (N8292, N8291, N7782, N334, N258);
and AND2 (N8293, N8279, N1451);
nor NOR4 (N8294, N8290, N4527, N392, N1904);
buf BUF1 (N8295, N8293);
not NOT1 (N8296, N8289);
nor NOR4 (N8297, N8287, N3614, N7687, N7863);
or OR3 (N8298, N8282, N8003, N6971);
and AND3 (N8299, N8283, N3513, N6453);
nand NAND2 (N8300, N8284, N4565);
nand NAND3 (N8301, N8297, N941, N5814);
nand NAND4 (N8302, N8288, N1853, N2265, N422);
not NOT1 (N8303, N8302);
nor NOR3 (N8304, N8301, N8214, N1695);
or OR2 (N8305, N8295, N6430);
nor NOR2 (N8306, N8292, N2064);
or OR4 (N8307, N8294, N953, N7287, N6965);
not NOT1 (N8308, N8296);
and AND2 (N8309, N8308, N8229);
not NOT1 (N8310, N8300);
xor XOR2 (N8311, N8303, N934);
not NOT1 (N8312, N8309);
buf BUF1 (N8313, N8310);
and AND2 (N8314, N8312, N5211);
buf BUF1 (N8315, N8286);
or OR4 (N8316, N8304, N6610, N1708, N7452);
not NOT1 (N8317, N8315);
nor NOR3 (N8318, N8298, N3786, N4480);
not NOT1 (N8319, N8317);
xor XOR2 (N8320, N8307, N4907);
not NOT1 (N8321, N8316);
nor NOR4 (N8322, N8305, N7405, N2181, N684);
and AND4 (N8323, N8306, N2123, N6580, N1230);
xor XOR2 (N8324, N8318, N4004);
xor XOR2 (N8325, N8314, N4348);
and AND3 (N8326, N8323, N2239, N2467);
and AND4 (N8327, N8299, N3772, N561, N6702);
buf BUF1 (N8328, N8325);
not NOT1 (N8329, N8326);
xor XOR2 (N8330, N8321, N5353);
or OR4 (N8331, N8311, N1559, N6620, N3565);
nand NAND2 (N8332, N8313, N3944);
or OR2 (N8333, N8329, N2893);
buf BUF1 (N8334, N8327);
buf BUF1 (N8335, N8319);
not NOT1 (N8336, N8330);
nand NAND4 (N8337, N8328, N6529, N2107, N400);
and AND4 (N8338, N8333, N5012, N7811, N3309);
nor NOR3 (N8339, N8337, N3866, N1147);
xor XOR2 (N8340, N8332, N5897);
buf BUF1 (N8341, N8338);
or OR2 (N8342, N8331, N4821);
nand NAND3 (N8343, N8335, N6570, N2401);
xor XOR2 (N8344, N8320, N8036);
xor XOR2 (N8345, N8344, N7357);
not NOT1 (N8346, N8343);
not NOT1 (N8347, N8334);
buf BUF1 (N8348, N8346);
nand NAND3 (N8349, N8324, N1446, N1387);
not NOT1 (N8350, N8336);
nand NAND2 (N8351, N8348, N820);
not NOT1 (N8352, N8351);
and AND4 (N8353, N8345, N6556, N3178, N653);
nand NAND3 (N8354, N8342, N4706, N3432);
not NOT1 (N8355, N8347);
and AND4 (N8356, N8341, N7335, N2576, N5319);
xor XOR2 (N8357, N8355, N1663);
nand NAND4 (N8358, N8322, N4280, N5948, N2230);
nand NAND4 (N8359, N8353, N1695, N2489, N2165);
and AND3 (N8360, N8357, N4217, N4506);
or OR2 (N8361, N8360, N4383);
xor XOR2 (N8362, N8361, N5534);
nor NOR2 (N8363, N8339, N3295);
xor XOR2 (N8364, N8359, N6227);
xor XOR2 (N8365, N8340, N8319);
buf BUF1 (N8366, N8363);
xor XOR2 (N8367, N8349, N3182);
nor NOR3 (N8368, N8366, N2290, N1916);
or OR4 (N8369, N8354, N6461, N2493, N6544);
not NOT1 (N8370, N8368);
xor XOR2 (N8371, N8352, N3831);
not NOT1 (N8372, N8364);
xor XOR2 (N8373, N8358, N5552);
buf BUF1 (N8374, N8369);
nand NAND4 (N8375, N8374, N6473, N3872, N1583);
nand NAND2 (N8376, N8367, N1067);
nand NAND4 (N8377, N8350, N2674, N6834, N6362);
and AND2 (N8378, N8372, N4418);
and AND2 (N8379, N8376, N1045);
and AND2 (N8380, N8362, N1701);
buf BUF1 (N8381, N8380);
nand NAND2 (N8382, N8379, N1044);
nor NOR2 (N8383, N8371, N8291);
nor NOR4 (N8384, N8375, N6693, N2935, N5734);
buf BUF1 (N8385, N8370);
or OR2 (N8386, N8377, N2468);
buf BUF1 (N8387, N8365);
not NOT1 (N8388, N8384);
nand NAND3 (N8389, N8387, N8233, N5078);
xor XOR2 (N8390, N8382, N7538);
buf BUF1 (N8391, N8386);
not NOT1 (N8392, N8381);
nor NOR4 (N8393, N8378, N3790, N6404, N820);
or OR3 (N8394, N8389, N6486, N3694);
nand NAND4 (N8395, N8393, N1519, N2806, N3187);
nand NAND4 (N8396, N8383, N3180, N2835, N946);
buf BUF1 (N8397, N8356);
buf BUF1 (N8398, N8391);
xor XOR2 (N8399, N8388, N4316);
nand NAND3 (N8400, N8394, N3958, N1704);
xor XOR2 (N8401, N8392, N4686);
not NOT1 (N8402, N8390);
and AND2 (N8403, N8396, N2621);
or OR2 (N8404, N8373, N1658);
nand NAND4 (N8405, N8398, N5795, N2132, N4536);
xor XOR2 (N8406, N8397, N1627);
xor XOR2 (N8407, N8395, N297);
xor XOR2 (N8408, N8402, N391);
buf BUF1 (N8409, N8385);
buf BUF1 (N8410, N8399);
buf BUF1 (N8411, N8405);
or OR2 (N8412, N8400, N2023);
or OR4 (N8413, N8408, N6083, N6696, N5532);
not NOT1 (N8414, N8409);
nand NAND2 (N8415, N8404, N7589);
nor NOR4 (N8416, N8415, N3671, N1076, N1297);
xor XOR2 (N8417, N8416, N7882);
xor XOR2 (N8418, N8411, N660);
xor XOR2 (N8419, N8414, N4619);
nor NOR4 (N8420, N8403, N6774, N4859, N8408);
buf BUF1 (N8421, N8418);
nor NOR3 (N8422, N8417, N1411, N6384);
and AND3 (N8423, N8406, N6333, N1902);
nor NOR2 (N8424, N8420, N7611);
xor XOR2 (N8425, N8419, N1929);
nand NAND2 (N8426, N8424, N6312);
and AND4 (N8427, N8407, N5755, N2422, N6618);
and AND4 (N8428, N8425, N7913, N6410, N5851);
nor NOR4 (N8429, N8413, N5247, N8063, N7419);
or OR2 (N8430, N8422, N2314);
nor NOR2 (N8431, N8429, N4566);
nor NOR2 (N8432, N8412, N2307);
or OR3 (N8433, N8426, N2829, N8044);
xor XOR2 (N8434, N8401, N4102);
not NOT1 (N8435, N8430);
xor XOR2 (N8436, N8427, N4556);
nor NOR3 (N8437, N8421, N4997, N2650);
xor XOR2 (N8438, N8434, N2208);
not NOT1 (N8439, N8428);
not NOT1 (N8440, N8423);
and AND3 (N8441, N8410, N3272, N4353);
nand NAND2 (N8442, N8439, N3677);
nor NOR3 (N8443, N8433, N3029, N3968);
and AND2 (N8444, N8431, N577);
xor XOR2 (N8445, N8440, N882);
nor NOR4 (N8446, N8445, N4495, N568, N1240);
nor NOR4 (N8447, N8432, N827, N1022, N4200);
and AND2 (N8448, N8442, N2340);
buf BUF1 (N8449, N8444);
nand NAND4 (N8450, N8437, N6555, N4961, N3504);
xor XOR2 (N8451, N8446, N5050);
not NOT1 (N8452, N8449);
nand NAND3 (N8453, N8435, N3376, N536);
nor NOR4 (N8454, N8441, N1288, N6069, N5876);
nor NOR3 (N8455, N8454, N5799, N4361);
or OR3 (N8456, N8450, N3258, N6973);
or OR3 (N8457, N8452, N1066, N508);
buf BUF1 (N8458, N8453);
xor XOR2 (N8459, N8447, N7689);
and AND2 (N8460, N8458, N2107);
nor NOR4 (N8461, N8438, N7934, N5838, N4829);
and AND4 (N8462, N8460, N7684, N3491, N5469);
nor NOR4 (N8463, N8459, N8289, N8304, N5309);
not NOT1 (N8464, N8463);
not NOT1 (N8465, N8455);
not NOT1 (N8466, N8464);
and AND3 (N8467, N8461, N3008, N6322);
or OR4 (N8468, N8436, N4552, N5464, N6689);
buf BUF1 (N8469, N8462);
buf BUF1 (N8470, N8468);
nand NAND2 (N8471, N8466, N1141);
buf BUF1 (N8472, N8467);
buf BUF1 (N8473, N8469);
not NOT1 (N8474, N8473);
buf BUF1 (N8475, N8448);
not NOT1 (N8476, N8443);
xor XOR2 (N8477, N8457, N2101);
and AND4 (N8478, N8451, N1642, N3599, N6819);
buf BUF1 (N8479, N8471);
nor NOR3 (N8480, N8477, N2798, N4706);
buf BUF1 (N8481, N8474);
xor XOR2 (N8482, N8470, N113);
nor NOR3 (N8483, N8480, N6377, N1865);
nor NOR4 (N8484, N8479, N7624, N4199, N3722);
nor NOR2 (N8485, N8465, N3470);
xor XOR2 (N8486, N8481, N2726);
nand NAND4 (N8487, N8486, N7217, N5482, N6454);
xor XOR2 (N8488, N8472, N2487);
nor NOR2 (N8489, N8475, N674);
and AND2 (N8490, N8489, N5006);
xor XOR2 (N8491, N8482, N4158);
and AND4 (N8492, N8487, N5198, N1156, N8398);
buf BUF1 (N8493, N8492);
not NOT1 (N8494, N8483);
nand NAND3 (N8495, N8484, N4887, N5889);
or OR3 (N8496, N8488, N7414, N1928);
nand NAND3 (N8497, N8490, N7749, N661);
nand NAND4 (N8498, N8478, N757, N6245, N5300);
nand NAND4 (N8499, N8497, N7648, N7400, N3274);
not NOT1 (N8500, N8496);
nor NOR4 (N8501, N8493, N4683, N7376, N7);
nor NOR3 (N8502, N8500, N4761, N6387);
not NOT1 (N8503, N8485);
nand NAND3 (N8504, N8495, N6130, N1464);
nand NAND2 (N8505, N8504, N1098);
not NOT1 (N8506, N8498);
xor XOR2 (N8507, N8499, N7891);
nor NOR2 (N8508, N8491, N2018);
or OR4 (N8509, N8507, N2163, N4810, N6783);
not NOT1 (N8510, N8506);
nand NAND4 (N8511, N8494, N6848, N3187, N7958);
not NOT1 (N8512, N8510);
and AND2 (N8513, N8501, N2466);
nand NAND4 (N8514, N8511, N6901, N4450, N6974);
xor XOR2 (N8515, N8513, N1390);
buf BUF1 (N8516, N8505);
nand NAND2 (N8517, N8512, N7827);
nand NAND4 (N8518, N8515, N728, N1667, N6769);
and AND4 (N8519, N8509, N4777, N4708, N7733);
and AND2 (N8520, N8476, N6149);
buf BUF1 (N8521, N8503);
nand NAND4 (N8522, N8521, N3900, N6923, N7152);
not NOT1 (N8523, N8514);
not NOT1 (N8524, N8502);
not NOT1 (N8525, N8524);
nor NOR4 (N8526, N8508, N3060, N7073, N2359);
nor NOR2 (N8527, N8518, N4614);
and AND4 (N8528, N8525, N517, N5460, N796);
nand NAND2 (N8529, N8517, N5973);
nand NAND2 (N8530, N8456, N4395);
and AND4 (N8531, N8528, N4327, N6593, N4875);
not NOT1 (N8532, N8530);
nand NAND4 (N8533, N8529, N4036, N456, N5981);
or OR4 (N8534, N8520, N5164, N2872, N7891);
buf BUF1 (N8535, N8534);
xor XOR2 (N8536, N8522, N2790);
nor NOR2 (N8537, N8533, N3440);
nand NAND2 (N8538, N8526, N5664);
or OR2 (N8539, N8537, N328);
or OR4 (N8540, N8536, N3376, N8275, N4743);
nor NOR3 (N8541, N8538, N6758, N3409);
and AND2 (N8542, N8540, N4294);
not NOT1 (N8543, N8539);
not NOT1 (N8544, N8531);
and AND2 (N8545, N8523, N3448);
nand NAND2 (N8546, N8519, N1369);
or OR3 (N8547, N8543, N3285, N201);
or OR2 (N8548, N8527, N5609);
buf BUF1 (N8549, N8548);
nand NAND4 (N8550, N8549, N303, N1719, N7871);
nor NOR4 (N8551, N8545, N4083, N3176, N6812);
nand NAND2 (N8552, N8551, N8378);
buf BUF1 (N8553, N8542);
and AND2 (N8554, N8552, N1848);
xor XOR2 (N8555, N8535, N462);
or OR2 (N8556, N8541, N2977);
or OR2 (N8557, N8547, N2859);
buf BUF1 (N8558, N8550);
xor XOR2 (N8559, N8544, N8473);
and AND4 (N8560, N8555, N1972, N899, N7768);
or OR4 (N8561, N8557, N6928, N8284, N848);
and AND4 (N8562, N8554, N1226, N6457, N2921);
nor NOR3 (N8563, N8559, N2991, N505);
nor NOR2 (N8564, N8516, N4340);
xor XOR2 (N8565, N8532, N8469);
nand NAND3 (N8566, N8553, N559, N282);
nor NOR4 (N8567, N8566, N2676, N3322, N7146);
nor NOR2 (N8568, N8565, N5051);
buf BUF1 (N8569, N8564);
not NOT1 (N8570, N8567);
nor NOR4 (N8571, N8558, N848, N7001, N7690);
nand NAND3 (N8572, N8569, N1028, N6383);
and AND3 (N8573, N8572, N2723, N7612);
xor XOR2 (N8574, N8546, N5487);
and AND2 (N8575, N8570, N8238);
xor XOR2 (N8576, N8575, N6889);
nand NAND2 (N8577, N8560, N4145);
buf BUF1 (N8578, N8574);
nand NAND4 (N8579, N8562, N5668, N5212, N5420);
buf BUF1 (N8580, N8578);
and AND2 (N8581, N8579, N6091);
xor XOR2 (N8582, N8573, N4772);
buf BUF1 (N8583, N8571);
or OR4 (N8584, N8580, N6644, N4688, N5122);
not NOT1 (N8585, N8584);
nor NOR4 (N8586, N8582, N2593, N4991, N4214);
nor NOR4 (N8587, N8583, N655, N5548, N8090);
nand NAND4 (N8588, N8586, N5525, N5360, N5908);
and AND2 (N8589, N8576, N2158);
buf BUF1 (N8590, N8577);
buf BUF1 (N8591, N8588);
and AND2 (N8592, N8581, N5348);
nand NAND3 (N8593, N8561, N2475, N6312);
or OR4 (N8594, N8591, N2707, N3373, N6035);
not NOT1 (N8595, N8592);
buf BUF1 (N8596, N8585);
nor NOR3 (N8597, N8563, N6088, N4202);
not NOT1 (N8598, N8556);
not NOT1 (N8599, N8594);
and AND3 (N8600, N8595, N6409, N5741);
buf BUF1 (N8601, N8590);
and AND4 (N8602, N8597, N1511, N707, N166);
not NOT1 (N8603, N8598);
nand NAND4 (N8604, N8568, N261, N355, N4888);
buf BUF1 (N8605, N8602);
or OR2 (N8606, N8600, N5451);
not NOT1 (N8607, N8589);
nor NOR3 (N8608, N8596, N7150, N5047);
or OR4 (N8609, N8593, N7608, N5785, N3246);
and AND4 (N8610, N8587, N7648, N8261, N4203);
nand NAND3 (N8611, N8610, N5924, N5);
xor XOR2 (N8612, N8599, N1307);
xor XOR2 (N8613, N8601, N3790);
nand NAND4 (N8614, N8609, N2945, N4348, N6414);
or OR4 (N8615, N8608, N5347, N8027, N8046);
nor NOR4 (N8616, N8607, N2328, N6467, N6096);
nor NOR4 (N8617, N8604, N6516, N5992, N5180);
or OR3 (N8618, N8605, N7468, N6966);
nand NAND2 (N8619, N8614, N7420);
nor NOR3 (N8620, N8603, N767, N7664);
and AND4 (N8621, N8619, N4998, N4960, N179);
and AND2 (N8622, N8615, N2765);
xor XOR2 (N8623, N8611, N4229);
xor XOR2 (N8624, N8622, N1109);
nand NAND3 (N8625, N8621, N2205, N5987);
buf BUF1 (N8626, N8624);
buf BUF1 (N8627, N8617);
and AND2 (N8628, N8620, N4742);
nand NAND2 (N8629, N8618, N6884);
nor NOR4 (N8630, N8628, N5005, N2920, N5348);
buf BUF1 (N8631, N8627);
nor NOR4 (N8632, N8606, N3784, N8413, N7996);
or OR4 (N8633, N8632, N665, N2487, N4464);
xor XOR2 (N8634, N8613, N4463);
and AND2 (N8635, N8612, N3415);
xor XOR2 (N8636, N8629, N2167);
and AND2 (N8637, N8634, N8429);
nand NAND4 (N8638, N8616, N3793, N4818, N6387);
and AND2 (N8639, N8637, N3687);
nand NAND2 (N8640, N8630, N2113);
not NOT1 (N8641, N8631);
not NOT1 (N8642, N8633);
not NOT1 (N8643, N8635);
nor NOR4 (N8644, N8643, N2474, N938, N6795);
nand NAND4 (N8645, N8636, N7739, N2207, N8358);
nor NOR4 (N8646, N8645, N1208, N5500, N2778);
xor XOR2 (N8647, N8626, N2445);
nor NOR4 (N8648, N8646, N2794, N8478, N7396);
xor XOR2 (N8649, N8640, N5399);
buf BUF1 (N8650, N8639);
and AND3 (N8651, N8650, N4141, N2083);
xor XOR2 (N8652, N8648, N633);
buf BUF1 (N8653, N8625);
nand NAND4 (N8654, N8644, N4803, N3407, N983);
or OR4 (N8655, N8623, N2690, N6440, N5977);
not NOT1 (N8656, N8649);
or OR4 (N8657, N8655, N7347, N5284, N4339);
and AND3 (N8658, N8654, N3733, N615);
xor XOR2 (N8659, N8653, N3774);
not NOT1 (N8660, N8657);
and AND3 (N8661, N8659, N2393, N3013);
and AND2 (N8662, N8642, N3262);
buf BUF1 (N8663, N8647);
and AND3 (N8664, N8651, N5007, N1031);
and AND4 (N8665, N8658, N6367, N3389, N3356);
nand NAND4 (N8666, N8662, N7645, N5149, N2507);
buf BUF1 (N8667, N8641);
or OR3 (N8668, N8667, N8555, N4243);
buf BUF1 (N8669, N8661);
or OR3 (N8670, N8665, N3059, N4227);
xor XOR2 (N8671, N8660, N829);
and AND2 (N8672, N8671, N331);
not NOT1 (N8673, N8652);
xor XOR2 (N8674, N8664, N6001);
buf BUF1 (N8675, N8674);
xor XOR2 (N8676, N8670, N4932);
xor XOR2 (N8677, N8666, N1971);
buf BUF1 (N8678, N8669);
not NOT1 (N8679, N8656);
buf BUF1 (N8680, N8673);
and AND4 (N8681, N8676, N6354, N1841, N4299);
nand NAND2 (N8682, N8680, N2388);
or OR4 (N8683, N8682, N6794, N7005, N4287);
nand NAND2 (N8684, N8663, N1852);
and AND2 (N8685, N8681, N2251);
nor NOR2 (N8686, N8685, N6533);
buf BUF1 (N8687, N8683);
nor NOR4 (N8688, N8678, N1510, N6546, N2850);
buf BUF1 (N8689, N8638);
and AND2 (N8690, N8689, N650);
not NOT1 (N8691, N8672);
xor XOR2 (N8692, N8691, N7473);
xor XOR2 (N8693, N8679, N2992);
and AND4 (N8694, N8693, N2237, N5186, N4944);
nor NOR2 (N8695, N8688, N1942);
and AND4 (N8696, N8668, N2332, N1740, N2042);
buf BUF1 (N8697, N8690);
or OR3 (N8698, N8687, N7466, N1604);
nor NOR3 (N8699, N8695, N1637, N7317);
nand NAND3 (N8700, N8698, N1151, N7009);
and AND4 (N8701, N8699, N6517, N2533, N2327);
nor NOR3 (N8702, N8696, N4850, N392);
or OR3 (N8703, N8700, N5803, N5680);
xor XOR2 (N8704, N8692, N2112);
buf BUF1 (N8705, N8675);
xor XOR2 (N8706, N8684, N3448);
xor XOR2 (N8707, N8702, N666);
buf BUF1 (N8708, N8686);
and AND3 (N8709, N8703, N7644, N5201);
not NOT1 (N8710, N8709);
or OR3 (N8711, N8707, N528, N5065);
nand NAND4 (N8712, N8694, N5977, N7349, N875);
or OR4 (N8713, N8711, N4423, N1838, N2471);
nor NOR3 (N8714, N8701, N6239, N6257);
xor XOR2 (N8715, N8710, N4795);
nor NOR3 (N8716, N8677, N6052, N5931);
nor NOR3 (N8717, N8715, N5343, N7730);
and AND4 (N8718, N8714, N6701, N4276, N3364);
and AND3 (N8719, N8697, N8312, N5866);
nor NOR4 (N8720, N8719, N2797, N1744, N618);
or OR4 (N8721, N8717, N6083, N8545, N6136);
or OR2 (N8722, N8712, N8545);
or OR2 (N8723, N8721, N997);
buf BUF1 (N8724, N8705);
nand NAND4 (N8725, N8724, N6892, N4804, N6294);
and AND3 (N8726, N8706, N5561, N2735);
and AND2 (N8727, N8725, N5768);
xor XOR2 (N8728, N8708, N6878);
or OR4 (N8729, N8718, N3857, N6804, N8029);
or OR4 (N8730, N8727, N8582, N1026, N1943);
buf BUF1 (N8731, N8729);
buf BUF1 (N8732, N8722);
xor XOR2 (N8733, N8713, N7189);
nand NAND3 (N8734, N8730, N6139, N8499);
nand NAND2 (N8735, N8716, N841);
nor NOR3 (N8736, N8720, N2941, N8538);
nor NOR2 (N8737, N8735, N2010);
and AND4 (N8738, N8704, N7369, N3867, N6981);
or OR3 (N8739, N8728, N5621, N973);
and AND4 (N8740, N8737, N7816, N3688, N29);
xor XOR2 (N8741, N8740, N8712);
nand NAND2 (N8742, N8736, N34);
nor NOR2 (N8743, N8726, N7609);
or OR4 (N8744, N8739, N6610, N8688, N3352);
not NOT1 (N8745, N8732);
xor XOR2 (N8746, N8733, N3984);
not NOT1 (N8747, N8742);
or OR2 (N8748, N8744, N2907);
or OR3 (N8749, N8748, N4195, N8208);
nand NAND4 (N8750, N8731, N3497, N5428, N4022);
or OR4 (N8751, N8750, N4380, N6094, N768);
buf BUF1 (N8752, N8747);
buf BUF1 (N8753, N8738);
buf BUF1 (N8754, N8741);
buf BUF1 (N8755, N8743);
or OR4 (N8756, N8745, N3202, N6592, N2397);
buf BUF1 (N8757, N8752);
nand NAND3 (N8758, N8734, N5478, N2835);
buf BUF1 (N8759, N8751);
buf BUF1 (N8760, N8749);
xor XOR2 (N8761, N8759, N5695);
not NOT1 (N8762, N8760);
nand NAND2 (N8763, N8757, N6800);
not NOT1 (N8764, N8756);
not NOT1 (N8765, N8746);
nor NOR4 (N8766, N8723, N5296, N83, N6615);
xor XOR2 (N8767, N8764, N3823);
xor XOR2 (N8768, N8765, N4935);
xor XOR2 (N8769, N8768, N791);
xor XOR2 (N8770, N8767, N3348);
nor NOR3 (N8771, N8769, N7956, N7944);
or OR3 (N8772, N8753, N7002, N1315);
nand NAND4 (N8773, N8755, N4061, N1588, N1652);
and AND3 (N8774, N8772, N290, N6591);
nand NAND3 (N8775, N8773, N3543, N2175);
buf BUF1 (N8776, N8762);
buf BUF1 (N8777, N8761);
not NOT1 (N8778, N8776);
not NOT1 (N8779, N8771);
xor XOR2 (N8780, N8778, N7443);
xor XOR2 (N8781, N8780, N924);
and AND4 (N8782, N8763, N8320, N3424, N6766);
nand NAND2 (N8783, N8782, N6126);
not NOT1 (N8784, N8783);
buf BUF1 (N8785, N8775);
xor XOR2 (N8786, N8774, N2521);
and AND2 (N8787, N8766, N4289);
or OR4 (N8788, N8787, N2440, N1657, N2723);
xor XOR2 (N8789, N8754, N3574);
or OR3 (N8790, N8770, N3754, N2335);
xor XOR2 (N8791, N8788, N1345);
and AND2 (N8792, N8786, N341);
xor XOR2 (N8793, N8789, N1537);
nand NAND3 (N8794, N8791, N2452, N2121);
not NOT1 (N8795, N8790);
nand NAND3 (N8796, N8779, N1271, N4364);
not NOT1 (N8797, N8781);
and AND4 (N8798, N8784, N4653, N5005, N7114);
nand NAND2 (N8799, N8794, N8353);
not NOT1 (N8800, N8785);
nand NAND3 (N8801, N8758, N8616, N7638);
nor NOR3 (N8802, N8792, N5677, N1291);
nor NOR3 (N8803, N8793, N4812, N2784);
and AND2 (N8804, N8801, N1888);
or OR2 (N8805, N8777, N5394);
and AND2 (N8806, N8805, N3127);
buf BUF1 (N8807, N8800);
buf BUF1 (N8808, N8806);
nand NAND2 (N8809, N8796, N8142);
not NOT1 (N8810, N8809);
nor NOR2 (N8811, N8802, N284);
nand NAND4 (N8812, N8811, N4921, N7846, N2708);
and AND2 (N8813, N8798, N7177);
not NOT1 (N8814, N8799);
nand NAND2 (N8815, N8810, N7763);
nor NOR4 (N8816, N8815, N7339, N1298, N1943);
nor NOR3 (N8817, N8812, N3374, N6313);
nand NAND3 (N8818, N8804, N2464, N2377);
nor NOR3 (N8819, N8817, N7799, N6773);
nor NOR2 (N8820, N8807, N6622);
nand NAND2 (N8821, N8808, N1198);
nor NOR2 (N8822, N8803, N7622);
buf BUF1 (N8823, N8816);
nand NAND3 (N8824, N8821, N4927, N442);
buf BUF1 (N8825, N8797);
nor NOR4 (N8826, N8820, N5477, N4188, N7587);
buf BUF1 (N8827, N8822);
nor NOR4 (N8828, N8826, N3443, N725, N1741);
or OR4 (N8829, N8795, N3290, N513, N1091);
and AND2 (N8830, N8829, N8261);
buf BUF1 (N8831, N8824);
buf BUF1 (N8832, N8827);
xor XOR2 (N8833, N8823, N7741);
nand NAND4 (N8834, N8828, N2297, N879, N2001);
nand NAND2 (N8835, N8825, N6003);
xor XOR2 (N8836, N8832, N507);
nor NOR2 (N8837, N8834, N3322);
buf BUF1 (N8838, N8833);
or OR3 (N8839, N8813, N1139, N5258);
buf BUF1 (N8840, N8831);
not NOT1 (N8841, N8839);
or OR4 (N8842, N8840, N885, N917, N7469);
nand NAND2 (N8843, N8836, N2457);
or OR2 (N8844, N8837, N7874);
nand NAND2 (N8845, N8841, N138);
nor NOR2 (N8846, N8818, N6103);
not NOT1 (N8847, N8814);
and AND2 (N8848, N8845, N3910);
buf BUF1 (N8849, N8838);
or OR2 (N8850, N8849, N5031);
nor NOR2 (N8851, N8843, N8846);
nor NOR3 (N8852, N606, N6290, N5685);
nor NOR3 (N8853, N8844, N102, N8760);
buf BUF1 (N8854, N8851);
or OR4 (N8855, N8848, N191, N217, N4234);
buf BUF1 (N8856, N8855);
nand NAND3 (N8857, N8856, N4724, N5334);
not NOT1 (N8858, N8850);
or OR4 (N8859, N8858, N6669, N3396, N4162);
not NOT1 (N8860, N8857);
buf BUF1 (N8861, N8842);
xor XOR2 (N8862, N8835, N1474);
or OR2 (N8863, N8853, N7811);
nand NAND2 (N8864, N8854, N7215);
nand NAND3 (N8865, N8860, N1505, N6692);
not NOT1 (N8866, N8847);
nor NOR3 (N8867, N8864, N6388, N5963);
or OR3 (N8868, N8852, N6849, N713);
and AND4 (N8869, N8866, N4461, N4882, N7162);
nand NAND2 (N8870, N8861, N7769);
or OR4 (N8871, N8859, N8677, N6420, N260);
nor NOR3 (N8872, N8830, N4881, N1802);
buf BUF1 (N8873, N8871);
buf BUF1 (N8874, N8863);
and AND4 (N8875, N8869, N6322, N2949, N3638);
or OR2 (N8876, N8865, N3805);
nand NAND2 (N8877, N8875, N4348);
buf BUF1 (N8878, N8862);
buf BUF1 (N8879, N8868);
xor XOR2 (N8880, N8878, N2168);
nor NOR2 (N8881, N8870, N4943);
and AND2 (N8882, N8873, N8197);
and AND2 (N8883, N8877, N7505);
not NOT1 (N8884, N8876);
buf BUF1 (N8885, N8880);
not NOT1 (N8886, N8884);
nand NAND4 (N8887, N8872, N2063, N4843, N1465);
or OR4 (N8888, N8885, N7069, N7133, N798);
or OR2 (N8889, N8867, N728);
nand NAND4 (N8890, N8874, N7913, N7382, N1895);
nand NAND3 (N8891, N8881, N1531, N8486);
buf BUF1 (N8892, N8891);
buf BUF1 (N8893, N8890);
and AND4 (N8894, N8886, N1132, N1140, N6883);
not NOT1 (N8895, N8879);
or OR4 (N8896, N8888, N3269, N748, N6991);
buf BUF1 (N8897, N8892);
nand NAND2 (N8898, N8893, N1792);
nor NOR4 (N8899, N8889, N240, N3711, N8437);
xor XOR2 (N8900, N8897, N6502);
buf BUF1 (N8901, N8899);
not NOT1 (N8902, N8883);
nand NAND4 (N8903, N8898, N1493, N7583, N4158);
or OR3 (N8904, N8895, N956, N1533);
and AND2 (N8905, N8900, N4427);
xor XOR2 (N8906, N8882, N2107);
buf BUF1 (N8907, N8905);
xor XOR2 (N8908, N8887, N5399);
not NOT1 (N8909, N8901);
xor XOR2 (N8910, N8902, N1299);
or OR4 (N8911, N8904, N5669, N8231, N801);
nor NOR3 (N8912, N8896, N7250, N6053);
nor NOR2 (N8913, N8911, N3967);
and AND3 (N8914, N8819, N7880, N5024);
buf BUF1 (N8915, N8910);
and AND2 (N8916, N8912, N8631);
nor NOR3 (N8917, N8909, N6367, N214);
xor XOR2 (N8918, N8917, N6934);
nor NOR2 (N8919, N8903, N1671);
not NOT1 (N8920, N8915);
nor NOR4 (N8921, N8919, N4241, N7169, N5150);
and AND2 (N8922, N8913, N3659);
nor NOR3 (N8923, N8922, N4059, N6882);
nor NOR4 (N8924, N8914, N2684, N3668, N6058);
or OR4 (N8925, N8908, N6564, N808, N3064);
and AND3 (N8926, N8921, N112, N3391);
buf BUF1 (N8927, N8924);
and AND2 (N8928, N8926, N5370);
not NOT1 (N8929, N8916);
buf BUF1 (N8930, N8894);
nand NAND4 (N8931, N8907, N1544, N440, N4825);
not NOT1 (N8932, N8918);
buf BUF1 (N8933, N8920);
and AND3 (N8934, N8906, N5070, N1799);
nand NAND3 (N8935, N8932, N1623, N901);
nand NAND4 (N8936, N8923, N8532, N7495, N1502);
nand NAND2 (N8937, N8927, N8158);
not NOT1 (N8938, N8934);
nand NAND3 (N8939, N8930, N4192, N1284);
or OR4 (N8940, N8928, N1353, N5189, N5203);
not NOT1 (N8941, N8936);
or OR4 (N8942, N8931, N6660, N3815, N4431);
xor XOR2 (N8943, N8939, N2963);
nand NAND3 (N8944, N8940, N7399, N2764);
nor NOR2 (N8945, N8935, N8740);
buf BUF1 (N8946, N8933);
nor NOR3 (N8947, N8942, N5932, N2176);
and AND3 (N8948, N8941, N7024, N1856);
nand NAND4 (N8949, N8943, N4692, N8261, N5561);
nor NOR4 (N8950, N8949, N3085, N5123, N6912);
not NOT1 (N8951, N8938);
nor NOR3 (N8952, N8929, N352, N2937);
nor NOR3 (N8953, N8945, N6625, N1461);
xor XOR2 (N8954, N8952, N2576);
nor NOR3 (N8955, N8946, N166, N2339);
not NOT1 (N8956, N8944);
not NOT1 (N8957, N8956);
xor XOR2 (N8958, N8953, N4165);
xor XOR2 (N8959, N8947, N3748);
buf BUF1 (N8960, N8950);
not NOT1 (N8961, N8951);
or OR2 (N8962, N8937, N3509);
and AND2 (N8963, N8955, N3412);
nand NAND4 (N8964, N8963, N122, N7058, N1171);
or OR3 (N8965, N8964, N811, N8227);
nand NAND3 (N8966, N8959, N2591, N46);
xor XOR2 (N8967, N8948, N7742);
nor NOR4 (N8968, N8966, N5543, N6660, N6637);
and AND4 (N8969, N8957, N4809, N190, N8072);
buf BUF1 (N8970, N8958);
or OR4 (N8971, N8961, N5956, N8552, N1019);
nand NAND2 (N8972, N8962, N1592);
and AND4 (N8973, N8970, N7383, N145, N4446);
buf BUF1 (N8974, N8967);
buf BUF1 (N8975, N8925);
not NOT1 (N8976, N8968);
buf BUF1 (N8977, N8973);
nor NOR3 (N8978, N8976, N4640, N8105);
and AND3 (N8979, N8977, N4273, N2842);
nand NAND2 (N8980, N8974, N8778);
and AND2 (N8981, N8972, N7877);
and AND4 (N8982, N8979, N6360, N2072, N6087);
not NOT1 (N8983, N8981);
buf BUF1 (N8984, N8980);
nand NAND2 (N8985, N8960, N4171);
xor XOR2 (N8986, N8983, N4475);
or OR3 (N8987, N8969, N2128, N7962);
and AND3 (N8988, N8982, N1694, N5252);
not NOT1 (N8989, N8975);
xor XOR2 (N8990, N8989, N4580);
or OR3 (N8991, N8985, N3571, N6063);
nor NOR4 (N8992, N8988, N6588, N4571, N3140);
nor NOR2 (N8993, N8978, N426);
nand NAND2 (N8994, N8971, N3756);
nand NAND4 (N8995, N8992, N5348, N6958, N3259);
xor XOR2 (N8996, N8954, N3527);
nor NOR4 (N8997, N8986, N8147, N3918, N2303);
xor XOR2 (N8998, N8994, N7537);
not NOT1 (N8999, N8990);
buf BUF1 (N9000, N8984);
not NOT1 (N9001, N8999);
or OR2 (N9002, N8995, N340);
or OR2 (N9003, N9002, N301);
and AND2 (N9004, N8965, N7224);
or OR3 (N9005, N8987, N6701, N6008);
xor XOR2 (N9006, N9001, N643);
nor NOR4 (N9007, N9000, N8258, N7419, N1186);
nand NAND4 (N9008, N8991, N4160, N867, N4542);
xor XOR2 (N9009, N9003, N470);
buf BUF1 (N9010, N9004);
not NOT1 (N9011, N8997);
not NOT1 (N9012, N9009);
and AND3 (N9013, N9012, N624, N3575);
buf BUF1 (N9014, N9007);
xor XOR2 (N9015, N8998, N335);
nand NAND4 (N9016, N9008, N2045, N1491, N2052);
or OR4 (N9017, N9010, N4219, N863, N4610);
nand NAND4 (N9018, N9006, N4613, N3159, N565);
xor XOR2 (N9019, N9011, N4205);
nand NAND3 (N9020, N9018, N3757, N6277);
xor XOR2 (N9021, N9014, N743);
or OR2 (N9022, N9017, N2909);
buf BUF1 (N9023, N9015);
buf BUF1 (N9024, N9019);
buf BUF1 (N9025, N9021);
and AND2 (N9026, N8993, N6350);
buf BUF1 (N9027, N9023);
xor XOR2 (N9028, N9016, N3288);
or OR2 (N9029, N9028, N8891);
xor XOR2 (N9030, N9020, N5836);
not NOT1 (N9031, N9026);
xor XOR2 (N9032, N9027, N8559);
buf BUF1 (N9033, N8996);
not NOT1 (N9034, N9013);
xor XOR2 (N9035, N9025, N3596);
or OR4 (N9036, N9030, N4809, N1831, N3816);
buf BUF1 (N9037, N9032);
or OR3 (N9038, N9037, N3251, N8518);
nor NOR2 (N9039, N9031, N781);
nor NOR2 (N9040, N9022, N1923);
buf BUF1 (N9041, N9024);
not NOT1 (N9042, N9041);
buf BUF1 (N9043, N9029);
nand NAND3 (N9044, N9043, N7149, N4496);
buf BUF1 (N9045, N9044);
buf BUF1 (N9046, N9005);
nand NAND4 (N9047, N9038, N7083, N801, N2482);
not NOT1 (N9048, N9046);
nand NAND3 (N9049, N9042, N301, N3991);
or OR3 (N9050, N9047, N8448, N875);
xor XOR2 (N9051, N9045, N8900);
nor NOR4 (N9052, N9050, N2861, N744, N1013);
buf BUF1 (N9053, N9051);
and AND3 (N9054, N9035, N5658, N7260);
nand NAND2 (N9055, N9034, N8462);
xor XOR2 (N9056, N9054, N6816);
buf BUF1 (N9057, N9048);
not NOT1 (N9058, N9049);
nand NAND3 (N9059, N9058, N2698, N2086);
and AND3 (N9060, N9033, N986, N2280);
xor XOR2 (N9061, N9052, N6250);
or OR2 (N9062, N9057, N5300);
nand NAND2 (N9063, N9059, N5948);
xor XOR2 (N9064, N9063, N6453);
nand NAND2 (N9065, N9061, N5008);
or OR4 (N9066, N9062, N712, N7260, N816);
or OR2 (N9067, N9040, N3935);
buf BUF1 (N9068, N9056);
xor XOR2 (N9069, N9060, N8043);
not NOT1 (N9070, N9065);
not NOT1 (N9071, N9053);
nand NAND3 (N9072, N9036, N3637, N5141);
or OR2 (N9073, N9066, N652);
xor XOR2 (N9074, N9064, N6496);
nor NOR3 (N9075, N9055, N370, N7601);
buf BUF1 (N9076, N9071);
nand NAND3 (N9077, N9070, N2015, N2719);
not NOT1 (N9078, N9077);
xor XOR2 (N9079, N9039, N1497);
or OR3 (N9080, N9067, N1786, N6388);
nor NOR4 (N9081, N9076, N2271, N3022, N8048);
xor XOR2 (N9082, N9068, N490);
buf BUF1 (N9083, N9075);
nor NOR2 (N9084, N9079, N594);
nand NAND2 (N9085, N9072, N5644);
not NOT1 (N9086, N9073);
or OR2 (N9087, N9080, N7444);
and AND4 (N9088, N9069, N728, N2720, N1134);
nand NAND4 (N9089, N9087, N7862, N890, N7464);
not NOT1 (N9090, N9082);
and AND2 (N9091, N9078, N6220);
or OR3 (N9092, N9088, N7062, N6013);
nand NAND3 (N9093, N9084, N3109, N7591);
buf BUF1 (N9094, N9090);
and AND3 (N9095, N9086, N1533, N5824);
nand NAND2 (N9096, N9074, N3717);
nand NAND3 (N9097, N9095, N8454, N5579);
xor XOR2 (N9098, N9096, N2731);
or OR3 (N9099, N9097, N7100, N207);
xor XOR2 (N9100, N9093, N755);
buf BUF1 (N9101, N9081);
buf BUF1 (N9102, N9089);
or OR2 (N9103, N9085, N6873);
buf BUF1 (N9104, N9083);
xor XOR2 (N9105, N9103, N434);
buf BUF1 (N9106, N9094);
nand NAND3 (N9107, N9100, N3129, N6549);
and AND2 (N9108, N9098, N7214);
and AND4 (N9109, N9108, N7951, N1707, N7554);
nor NOR2 (N9110, N9106, N8545);
buf BUF1 (N9111, N9099);
nand NAND4 (N9112, N9092, N8064, N8246, N1318);
nor NOR3 (N9113, N9105, N175, N7282);
xor XOR2 (N9114, N9104, N1626);
and AND2 (N9115, N9111, N1131);
or OR4 (N9116, N9115, N7901, N7435, N4973);
xor XOR2 (N9117, N9107, N2083);
nor NOR4 (N9118, N9109, N8783, N7009, N608);
nor NOR3 (N9119, N9101, N5339, N2965);
nor NOR4 (N9120, N9118, N5068, N1257, N4736);
xor XOR2 (N9121, N9112, N5720);
nor NOR3 (N9122, N9120, N5813, N2856);
buf BUF1 (N9123, N9102);
buf BUF1 (N9124, N9116);
buf BUF1 (N9125, N9114);
xor XOR2 (N9126, N9122, N7910);
nor NOR2 (N9127, N9110, N4402);
and AND2 (N9128, N9113, N2988);
buf BUF1 (N9129, N9123);
nor NOR4 (N9130, N9128, N7248, N8667, N6690);
and AND2 (N9131, N9117, N8430);
not NOT1 (N9132, N9130);
buf BUF1 (N9133, N9119);
or OR2 (N9134, N9127, N2913);
and AND4 (N9135, N9134, N8186, N6742, N36);
not NOT1 (N9136, N9125);
not NOT1 (N9137, N9124);
xor XOR2 (N9138, N9129, N8568);
not NOT1 (N9139, N9133);
not NOT1 (N9140, N9139);
buf BUF1 (N9141, N9131);
nor NOR3 (N9142, N9141, N6178, N2219);
or OR2 (N9143, N9136, N3845);
buf BUF1 (N9144, N9091);
nor NOR3 (N9145, N9144, N4192, N5981);
xor XOR2 (N9146, N9135, N6433);
buf BUF1 (N9147, N9132);
nor NOR2 (N9148, N9143, N6944);
nand NAND4 (N9149, N9147, N2217, N5602, N7163);
nor NOR3 (N9150, N9142, N3615, N8328);
nand NAND3 (N9151, N9150, N4304, N7391);
nand NAND3 (N9152, N9137, N3561, N691);
buf BUF1 (N9153, N9151);
or OR3 (N9154, N9148, N2296, N6253);
not NOT1 (N9155, N9146);
buf BUF1 (N9156, N9138);
not NOT1 (N9157, N9154);
and AND4 (N9158, N9156, N909, N1494, N1015);
nand NAND4 (N9159, N9121, N7855, N2288, N5437);
nor NOR4 (N9160, N9157, N1818, N2458, N7477);
not NOT1 (N9161, N9145);
buf BUF1 (N9162, N9152);
nor NOR3 (N9163, N9158, N2638, N4265);
buf BUF1 (N9164, N9149);
xor XOR2 (N9165, N9155, N2549);
nand NAND4 (N9166, N9160, N526, N919, N1069);
buf BUF1 (N9167, N9159);
nor NOR4 (N9168, N9163, N709, N820, N4542);
and AND3 (N9169, N9140, N6260, N6549);
not NOT1 (N9170, N9165);
not NOT1 (N9171, N9126);
not NOT1 (N9172, N9161);
nor NOR2 (N9173, N9170, N4673);
nand NAND3 (N9174, N9164, N6741, N4744);
nor NOR4 (N9175, N9173, N7293, N7133, N1968);
or OR2 (N9176, N9175, N5356);
nor NOR3 (N9177, N9166, N3310, N6543);
and AND4 (N9178, N9168, N6677, N5828, N9137);
not NOT1 (N9179, N9153);
buf BUF1 (N9180, N9176);
and AND2 (N9181, N9178, N8063);
xor XOR2 (N9182, N9169, N3550);
nand NAND2 (N9183, N9172, N1096);
or OR3 (N9184, N9167, N6260, N7445);
xor XOR2 (N9185, N9171, N4308);
xor XOR2 (N9186, N9180, N5902);
not NOT1 (N9187, N9185);
xor XOR2 (N9188, N9187, N6074);
and AND3 (N9189, N9182, N4259, N3533);
not NOT1 (N9190, N9186);
xor XOR2 (N9191, N9184, N5489);
xor XOR2 (N9192, N9188, N8270);
not NOT1 (N9193, N9192);
xor XOR2 (N9194, N9189, N4256);
nand NAND4 (N9195, N9183, N4935, N6623, N7037);
nor NOR4 (N9196, N9177, N7426, N5953, N2586);
xor XOR2 (N9197, N9194, N6597);
nand NAND3 (N9198, N9196, N8082, N555);
and AND2 (N9199, N9174, N8961);
or OR3 (N9200, N9179, N7704, N5949);
or OR3 (N9201, N9197, N6916, N8909);
buf BUF1 (N9202, N9200);
nand NAND2 (N9203, N9202, N872);
nand NAND4 (N9204, N9195, N6914, N4582, N3327);
xor XOR2 (N9205, N9199, N4077);
nor NOR2 (N9206, N9191, N5527);
not NOT1 (N9207, N9198);
nand NAND3 (N9208, N9203, N7508, N2856);
nor NOR4 (N9209, N9206, N4590, N2034, N2750);
nand NAND3 (N9210, N9162, N7778, N5243);
nand NAND2 (N9211, N9201, N604);
buf BUF1 (N9212, N9207);
not NOT1 (N9213, N9212);
nor NOR4 (N9214, N9210, N7565, N6072, N519);
nor NOR4 (N9215, N9208, N58, N2701, N7304);
nand NAND2 (N9216, N9213, N1796);
buf BUF1 (N9217, N9190);
or OR2 (N9218, N9204, N6669);
nor NOR3 (N9219, N9217, N9191, N532);
nor NOR2 (N9220, N9219, N6352);
nand NAND4 (N9221, N9218, N1567, N5519, N7747);
or OR4 (N9222, N9221, N5651, N4779, N8379);
nand NAND3 (N9223, N9215, N8900, N5064);
or OR2 (N9224, N9222, N8768);
nor NOR3 (N9225, N9211, N3413, N1403);
xor XOR2 (N9226, N9220, N2277);
nand NAND3 (N9227, N9181, N1856, N1273);
xor XOR2 (N9228, N9226, N7999);
not NOT1 (N9229, N9223);
or OR3 (N9230, N9209, N5740, N2389);
xor XOR2 (N9231, N9216, N4503);
not NOT1 (N9232, N9214);
xor XOR2 (N9233, N9227, N8571);
nand NAND2 (N9234, N9230, N5392);
or OR2 (N9235, N9205, N2177);
buf BUF1 (N9236, N9231);
or OR3 (N9237, N9228, N8991, N8071);
nor NOR4 (N9238, N9233, N1580, N1776, N6258);
buf BUF1 (N9239, N9224);
not NOT1 (N9240, N9229);
not NOT1 (N9241, N9240);
and AND2 (N9242, N9236, N2816);
nand NAND4 (N9243, N9193, N7616, N3713, N4693);
buf BUF1 (N9244, N9238);
nor NOR3 (N9245, N9243, N2123, N1897);
or OR3 (N9246, N9239, N1736, N2769);
nor NOR4 (N9247, N9232, N5517, N3331, N6077);
or OR3 (N9248, N9244, N7624, N1287);
nor NOR4 (N9249, N9246, N3090, N6406, N4738);
nand NAND4 (N9250, N9237, N5629, N2951, N5316);
or OR2 (N9251, N9225, N8672);
not NOT1 (N9252, N9250);
buf BUF1 (N9253, N9245);
and AND4 (N9254, N9253, N3924, N8799, N5066);
and AND2 (N9255, N9254, N4822);
or OR3 (N9256, N9255, N7632, N6657);
not NOT1 (N9257, N9234);
xor XOR2 (N9258, N9252, N2395);
and AND3 (N9259, N9242, N2849, N119);
or OR4 (N9260, N9241, N6889, N5092, N4455);
xor XOR2 (N9261, N9251, N1958);
nor NOR4 (N9262, N9249, N4761, N7304, N7593);
not NOT1 (N9263, N9259);
or OR4 (N9264, N9248, N714, N1935, N2613);
and AND2 (N9265, N9263, N6849);
or OR3 (N9266, N9256, N3289, N2897);
nor NOR3 (N9267, N9264, N3918, N6657);
buf BUF1 (N9268, N9261);
not NOT1 (N9269, N9268);
xor XOR2 (N9270, N9267, N4546);
nor NOR3 (N9271, N9265, N3529, N1743);
xor XOR2 (N9272, N9271, N6292);
and AND3 (N9273, N9272, N381, N678);
buf BUF1 (N9274, N9266);
or OR4 (N9275, N9260, N6156, N7777, N7119);
not NOT1 (N9276, N9262);
nor NOR2 (N9277, N9275, N8070);
buf BUF1 (N9278, N9277);
xor XOR2 (N9279, N9270, N8887);
nand NAND2 (N9280, N9274, N2534);
nor NOR4 (N9281, N9278, N7934, N2063, N1099);
not NOT1 (N9282, N9247);
nand NAND4 (N9283, N9269, N2112, N2636, N6875);
buf BUF1 (N9284, N9273);
or OR2 (N9285, N9284, N1585);
not NOT1 (N9286, N9280);
nor NOR2 (N9287, N9258, N4777);
not NOT1 (N9288, N9281);
or OR2 (N9289, N9286, N1090);
xor XOR2 (N9290, N9285, N4848);
and AND4 (N9291, N9235, N180, N6616, N6404);
nor NOR4 (N9292, N9290, N8759, N6906, N8289);
nor NOR4 (N9293, N9287, N8750, N7824, N1543);
not NOT1 (N9294, N9288);
xor XOR2 (N9295, N9282, N4053);
not NOT1 (N9296, N9294);
or OR4 (N9297, N9276, N942, N210, N1446);
or OR3 (N9298, N9279, N6387, N7275);
nand NAND4 (N9299, N9295, N3275, N823, N7507);
and AND4 (N9300, N9297, N7182, N2086, N4566);
and AND4 (N9301, N9257, N2919, N3332, N3772);
and AND3 (N9302, N9289, N832, N3448);
nor NOR3 (N9303, N9293, N7503, N4167);
nand NAND2 (N9304, N9291, N3609);
or OR4 (N9305, N9298, N8728, N5872, N5191);
nor NOR2 (N9306, N9304, N1351);
and AND2 (N9307, N9296, N3617);
or OR3 (N9308, N9292, N2982, N4664);
not NOT1 (N9309, N9308);
or OR3 (N9310, N9303, N4112, N152);
nand NAND3 (N9311, N9307, N4221, N34);
or OR3 (N9312, N9309, N9110, N2083);
nor NOR4 (N9313, N9302, N3270, N6727, N4623);
and AND2 (N9314, N9306, N8744);
and AND4 (N9315, N9299, N7519, N4347, N421);
and AND4 (N9316, N9301, N5688, N1873, N1691);
nor NOR2 (N9317, N9311, N681);
buf BUF1 (N9318, N9283);
not NOT1 (N9319, N9300);
buf BUF1 (N9320, N9317);
not NOT1 (N9321, N9315);
xor XOR2 (N9322, N9312, N3016);
nor NOR2 (N9323, N9318, N493);
not NOT1 (N9324, N9305);
not NOT1 (N9325, N9322);
nand NAND2 (N9326, N9319, N7525);
not NOT1 (N9327, N9314);
buf BUF1 (N9328, N9310);
or OR3 (N9329, N9324, N5176, N6069);
or OR3 (N9330, N9328, N5826, N8696);
nor NOR2 (N9331, N9330, N3453);
or OR4 (N9332, N9323, N4282, N7772, N4042);
xor XOR2 (N9333, N9320, N7164);
nor NOR3 (N9334, N9333, N3646, N1972);
and AND3 (N9335, N9313, N7307, N6985);
nor NOR2 (N9336, N9334, N6943);
buf BUF1 (N9337, N9327);
xor XOR2 (N9338, N9316, N417);
not NOT1 (N9339, N9336);
and AND3 (N9340, N9325, N4897, N2613);
or OR2 (N9341, N9321, N8498);
not NOT1 (N9342, N9332);
nand NAND4 (N9343, N9331, N7299, N8925, N7423);
nand NAND4 (N9344, N9343, N8312, N6762, N2563);
nand NAND3 (N9345, N9326, N9264, N5941);
xor XOR2 (N9346, N9339, N4509);
and AND3 (N9347, N9329, N781, N43);
buf BUF1 (N9348, N9344);
xor XOR2 (N9349, N9341, N3316);
nand NAND4 (N9350, N9348, N1743, N8926, N2849);
not NOT1 (N9351, N9346);
or OR4 (N9352, N9349, N3832, N5329, N8230);
buf BUF1 (N9353, N9350);
buf BUF1 (N9354, N9338);
nand NAND2 (N9355, N9342, N9118);
or OR3 (N9356, N9352, N3293, N4716);
nand NAND4 (N9357, N9345, N3571, N571, N2408);
buf BUF1 (N9358, N9354);
nor NOR3 (N9359, N9337, N8720, N4661);
nor NOR3 (N9360, N9347, N1679, N8576);
nor NOR2 (N9361, N9357, N3269);
xor XOR2 (N9362, N9358, N8644);
nor NOR4 (N9363, N9351, N58, N3427, N764);
not NOT1 (N9364, N9361);
xor XOR2 (N9365, N9364, N9212);
not NOT1 (N9366, N9335);
and AND4 (N9367, N9355, N7621, N4831, N1327);
xor XOR2 (N9368, N9367, N8784);
nand NAND2 (N9369, N9365, N5479);
buf BUF1 (N9370, N9369);
nand NAND4 (N9371, N9359, N1910, N5307, N1720);
or OR4 (N9372, N9366, N5065, N4737, N8155);
xor XOR2 (N9373, N9353, N2294);
nand NAND3 (N9374, N9371, N2068, N8740);
not NOT1 (N9375, N9374);
not NOT1 (N9376, N9375);
nand NAND2 (N9377, N9360, N4246);
xor XOR2 (N9378, N9377, N3754);
nor NOR3 (N9379, N9370, N6210, N693);
buf BUF1 (N9380, N9378);
nor NOR2 (N9381, N9372, N4666);
not NOT1 (N9382, N9373);
not NOT1 (N9383, N9362);
or OR2 (N9384, N9382, N7240);
buf BUF1 (N9385, N9384);
and AND2 (N9386, N9356, N4542);
and AND2 (N9387, N9381, N1842);
not NOT1 (N9388, N9380);
xor XOR2 (N9389, N9386, N8290);
not NOT1 (N9390, N9387);
not NOT1 (N9391, N9389);
xor XOR2 (N9392, N9340, N6041);
or OR2 (N9393, N9385, N6870);
not NOT1 (N9394, N9391);
xor XOR2 (N9395, N9388, N2101);
and AND4 (N9396, N9390, N9377, N4867, N1015);
nor NOR2 (N9397, N9383, N7909);
not NOT1 (N9398, N9395);
nand NAND3 (N9399, N9379, N195, N3111);
and AND4 (N9400, N9376, N1586, N1654, N5316);
nor NOR4 (N9401, N9368, N2317, N37, N2978);
xor XOR2 (N9402, N9392, N2803);
nand NAND2 (N9403, N9399, N8107);
buf BUF1 (N9404, N9397);
nand NAND3 (N9405, N9403, N6732, N4386);
and AND4 (N9406, N9393, N1011, N4340, N3249);
and AND2 (N9407, N9400, N3923);
xor XOR2 (N9408, N9407, N3922);
nor NOR3 (N9409, N9402, N1195, N1147);
and AND4 (N9410, N9404, N4900, N991, N6725);
buf BUF1 (N9411, N9406);
buf BUF1 (N9412, N9409);
and AND4 (N9413, N9396, N2950, N673, N8529);
nor NOR2 (N9414, N9408, N9383);
nor NOR3 (N9415, N9411, N3925, N6001);
not NOT1 (N9416, N9394);
xor XOR2 (N9417, N9413, N8019);
and AND4 (N9418, N9414, N8725, N733, N2866);
not NOT1 (N9419, N9363);
or OR4 (N9420, N9410, N9224, N2192, N3006);
buf BUF1 (N9421, N9419);
and AND4 (N9422, N9401, N9299, N1334, N319);
nor NOR2 (N9423, N9418, N9277);
and AND3 (N9424, N9405, N2373, N5924);
buf BUF1 (N9425, N9415);
nor NOR3 (N9426, N9416, N3927, N968);
and AND3 (N9427, N9426, N2308, N4);
xor XOR2 (N9428, N9424, N7402);
buf BUF1 (N9429, N9421);
xor XOR2 (N9430, N9429, N2036);
and AND4 (N9431, N9428, N6680, N598, N8964);
and AND2 (N9432, N9431, N866);
nor NOR3 (N9433, N9430, N472, N5163);
buf BUF1 (N9434, N9433);
and AND2 (N9435, N9434, N413);
buf BUF1 (N9436, N9423);
nand NAND2 (N9437, N9398, N8518);
or OR4 (N9438, N9435, N8001, N3979, N3734);
buf BUF1 (N9439, N9432);
nor NOR2 (N9440, N9420, N5476);
nor NOR3 (N9441, N9412, N4, N8221);
not NOT1 (N9442, N9425);
nor NOR3 (N9443, N9438, N5537, N5372);
nor NOR4 (N9444, N9437, N6953, N4231, N1411);
buf BUF1 (N9445, N9443);
xor XOR2 (N9446, N9427, N3362);
and AND4 (N9447, N9439, N2427, N8015, N8213);
buf BUF1 (N9448, N9417);
not NOT1 (N9449, N9442);
xor XOR2 (N9450, N9448, N2792);
buf BUF1 (N9451, N9441);
nor NOR3 (N9452, N9422, N2468, N3696);
or OR2 (N9453, N9447, N3297);
or OR2 (N9454, N9436, N5119);
or OR4 (N9455, N9440, N6746, N1464, N7985);
not NOT1 (N9456, N9454);
and AND2 (N9457, N9444, N6143);
not NOT1 (N9458, N9446);
nor NOR3 (N9459, N9452, N5786, N780);
buf BUF1 (N9460, N9455);
buf BUF1 (N9461, N9445);
or OR3 (N9462, N9457, N1523, N1209);
not NOT1 (N9463, N9459);
or OR2 (N9464, N9451, N8637);
or OR2 (N9465, N9449, N8738);
xor XOR2 (N9466, N9464, N2861);
nor NOR4 (N9467, N9450, N4024, N8781, N4515);
or OR2 (N9468, N9465, N51);
and AND4 (N9469, N9460, N5310, N2669, N8134);
or OR3 (N9470, N9458, N1920, N6936);
xor XOR2 (N9471, N9453, N8178);
and AND4 (N9472, N9467, N9380, N3831, N3452);
and AND3 (N9473, N9470, N2518, N4474);
xor XOR2 (N9474, N9456, N576);
xor XOR2 (N9475, N9473, N4851);
nor NOR4 (N9476, N9472, N5565, N262, N709);
xor XOR2 (N9477, N9471, N3964);
nand NAND4 (N9478, N9468, N2478, N4002, N1721);
nand NAND3 (N9479, N9469, N4681, N6496);
and AND4 (N9480, N9463, N6248, N4218, N549);
not NOT1 (N9481, N9476);
nor NOR3 (N9482, N9477, N627, N1553);
nor NOR3 (N9483, N9461, N3986, N2784);
nand NAND3 (N9484, N9466, N9065, N2754);
not NOT1 (N9485, N9479);
buf BUF1 (N9486, N9462);
nor NOR2 (N9487, N9484, N5545);
buf BUF1 (N9488, N9482);
buf BUF1 (N9489, N9486);
nor NOR4 (N9490, N9488, N8259, N4254, N2030);
nor NOR2 (N9491, N9480, N7552);
not NOT1 (N9492, N9474);
nand NAND2 (N9493, N9478, N3242);
xor XOR2 (N9494, N9492, N1845);
not NOT1 (N9495, N9487);
and AND4 (N9496, N9485, N3418, N8780, N5510);
not NOT1 (N9497, N9491);
buf BUF1 (N9498, N9489);
and AND4 (N9499, N9494, N4089, N1555, N830);
nor NOR4 (N9500, N9495, N4662, N1807, N1505);
xor XOR2 (N9501, N9497, N965);
buf BUF1 (N9502, N9499);
or OR2 (N9503, N9500, N8847);
not NOT1 (N9504, N9501);
not NOT1 (N9505, N9483);
and AND3 (N9506, N9493, N9135, N337);
buf BUF1 (N9507, N9505);
not NOT1 (N9508, N9504);
not NOT1 (N9509, N9507);
nor NOR3 (N9510, N9506, N2155, N4678);
not NOT1 (N9511, N9509);
and AND4 (N9512, N9496, N4911, N3004, N5362);
xor XOR2 (N9513, N9503, N8348);
xor XOR2 (N9514, N9513, N3645);
and AND3 (N9515, N9508, N6525, N3743);
nor NOR4 (N9516, N9502, N6303, N8246, N6534);
not NOT1 (N9517, N9510);
and AND4 (N9518, N9498, N7441, N119, N7849);
xor XOR2 (N9519, N9517, N1357);
and AND2 (N9520, N9490, N6456);
or OR2 (N9521, N9475, N4909);
nand NAND3 (N9522, N9519, N8980, N2838);
nand NAND3 (N9523, N9516, N7424, N1303);
not NOT1 (N9524, N9521);
xor XOR2 (N9525, N9518, N7496);
not NOT1 (N9526, N9511);
nand NAND3 (N9527, N9524, N4387, N7411);
nand NAND2 (N9528, N9526, N1441);
buf BUF1 (N9529, N9523);
not NOT1 (N9530, N9525);
nor NOR4 (N9531, N9527, N636, N5833, N8181);
or OR2 (N9532, N9481, N5247);
nor NOR2 (N9533, N9512, N1792);
and AND2 (N9534, N9530, N7791);
buf BUF1 (N9535, N9514);
nor NOR4 (N9536, N9533, N9266, N6085, N3111);
buf BUF1 (N9537, N9520);
xor XOR2 (N9538, N9528, N477);
buf BUF1 (N9539, N9537);
nand NAND4 (N9540, N9531, N15, N2123, N4944);
nor NOR2 (N9541, N9536, N9519);
buf BUF1 (N9542, N9539);
and AND3 (N9543, N9535, N6597, N7241);
or OR2 (N9544, N9542, N2629);
not NOT1 (N9545, N9515);
buf BUF1 (N9546, N9532);
nand NAND3 (N9547, N9534, N5644, N1592);
or OR4 (N9548, N9538, N1509, N1223, N6840);
nor NOR2 (N9549, N9548, N3727);
or OR3 (N9550, N9549, N6989, N5631);
nor NOR2 (N9551, N9529, N9497);
nand NAND3 (N9552, N9550, N1050, N2010);
and AND4 (N9553, N9540, N5040, N5727, N774);
not NOT1 (N9554, N9545);
not NOT1 (N9555, N9546);
xor XOR2 (N9556, N9544, N5422);
not NOT1 (N9557, N9543);
not NOT1 (N9558, N9541);
or OR2 (N9559, N9555, N1632);
nor NOR2 (N9560, N9558, N69);
nor NOR3 (N9561, N9522, N5524, N7372);
and AND3 (N9562, N9552, N1446, N5782);
buf BUF1 (N9563, N9560);
nand NAND2 (N9564, N9553, N7397);
nor NOR2 (N9565, N9562, N8224);
not NOT1 (N9566, N9557);
nor NOR2 (N9567, N9566, N4323);
or OR4 (N9568, N9547, N5472, N925, N4959);
xor XOR2 (N9569, N9567, N8413);
or OR4 (N9570, N9559, N4212, N3394, N2008);
xor XOR2 (N9571, N9565, N8089);
xor XOR2 (N9572, N9568, N8907);
buf BUF1 (N9573, N9563);
nor NOR4 (N9574, N9554, N9170, N2721, N932);
buf BUF1 (N9575, N9572);
and AND4 (N9576, N9571, N2954, N5721, N3190);
and AND3 (N9577, N9576, N9212, N2402);
and AND2 (N9578, N9551, N5760);
not NOT1 (N9579, N9569);
buf BUF1 (N9580, N9564);
not NOT1 (N9581, N9573);
not NOT1 (N9582, N9561);
nor NOR4 (N9583, N9574, N4957, N7813, N2672);
nor NOR2 (N9584, N9582, N441);
nor NOR4 (N9585, N9578, N2710, N7742, N6670);
xor XOR2 (N9586, N9583, N1364);
or OR3 (N9587, N9570, N2825, N6172);
xor XOR2 (N9588, N9587, N1530);
and AND2 (N9589, N9579, N7058);
and AND4 (N9590, N9577, N3998, N8560, N4200);
or OR4 (N9591, N9575, N4236, N3488, N8850);
and AND2 (N9592, N9556, N9247);
buf BUF1 (N9593, N9590);
not NOT1 (N9594, N9586);
nor NOR2 (N9595, N9584, N6470);
and AND3 (N9596, N9594, N6674, N8855);
or OR2 (N9597, N9580, N3947);
buf BUF1 (N9598, N9596);
or OR2 (N9599, N9593, N6670);
nor NOR3 (N9600, N9592, N5162, N5246);
nor NOR3 (N9601, N9597, N1744, N4035);
xor XOR2 (N9602, N9598, N74);
xor XOR2 (N9603, N9591, N5480);
or OR2 (N9604, N9600, N4359);
not NOT1 (N9605, N9588);
and AND2 (N9606, N9601, N1717);
buf BUF1 (N9607, N9603);
and AND2 (N9608, N9581, N3920);
nand NAND4 (N9609, N9599, N8385, N693, N2156);
or OR2 (N9610, N9595, N6174);
buf BUF1 (N9611, N9609);
not NOT1 (N9612, N9610);
and AND3 (N9613, N9585, N5882, N1922);
and AND3 (N9614, N9607, N1965, N6354);
nor NOR2 (N9615, N9604, N7131);
nor NOR4 (N9616, N9611, N6789, N2141, N5491);
nor NOR3 (N9617, N9589, N4440, N1902);
nor NOR2 (N9618, N9613, N2826);
nand NAND2 (N9619, N9615, N5281);
not NOT1 (N9620, N9619);
nand NAND3 (N9621, N9614, N4085, N4587);
and AND2 (N9622, N9617, N1185);
and AND4 (N9623, N9621, N2518, N571, N573);
nor NOR4 (N9624, N9616, N3840, N4057, N1096);
or OR3 (N9625, N9624, N8367, N8212);
not NOT1 (N9626, N9625);
and AND2 (N9627, N9612, N5060);
or OR3 (N9628, N9606, N2957, N763);
nand NAND2 (N9629, N9608, N1617);
buf BUF1 (N9630, N9620);
nor NOR4 (N9631, N9602, N115, N6369, N5079);
xor XOR2 (N9632, N9629, N7258);
not NOT1 (N9633, N9627);
buf BUF1 (N9634, N9628);
nand NAND2 (N9635, N9632, N2560);
not NOT1 (N9636, N9635);
buf BUF1 (N9637, N9634);
nand NAND3 (N9638, N9631, N1466, N9355);
xor XOR2 (N9639, N9626, N3531);
nor NOR4 (N9640, N9638, N1146, N1472, N7702);
xor XOR2 (N9641, N9639, N7201);
buf BUF1 (N9642, N9623);
or OR4 (N9643, N9630, N5186, N52, N4724);
nor NOR4 (N9644, N9641, N8379, N6746, N5285);
xor XOR2 (N9645, N9633, N2728);
xor XOR2 (N9646, N9645, N643);
not NOT1 (N9647, N9646);
nor NOR4 (N9648, N9622, N9021, N7995, N3050);
xor XOR2 (N9649, N9642, N4884);
nand NAND3 (N9650, N9605, N5700, N2026);
nand NAND2 (N9651, N9650, N2063);
xor XOR2 (N9652, N9651, N5395);
buf BUF1 (N9653, N9637);
nor NOR3 (N9654, N9643, N67, N7797);
nor NOR4 (N9655, N9618, N3136, N1318, N3969);
not NOT1 (N9656, N9654);
xor XOR2 (N9657, N9640, N4667);
not NOT1 (N9658, N9647);
not NOT1 (N9659, N9648);
or OR2 (N9660, N9658, N2746);
nor NOR2 (N9661, N9653, N5313);
not NOT1 (N9662, N9636);
or OR2 (N9663, N9661, N7010);
or OR4 (N9664, N9657, N739, N759, N5776);
or OR4 (N9665, N9656, N8198, N9500, N9344);
not NOT1 (N9666, N9652);
buf BUF1 (N9667, N9663);
and AND4 (N9668, N9660, N3255, N2264, N6592);
nor NOR2 (N9669, N9659, N375);
nand NAND2 (N9670, N9668, N7573);
and AND2 (N9671, N9669, N5716);
and AND3 (N9672, N9655, N1870, N486);
or OR2 (N9673, N9649, N3657);
not NOT1 (N9674, N9662);
xor XOR2 (N9675, N9671, N8880);
xor XOR2 (N9676, N9667, N2277);
xor XOR2 (N9677, N9670, N7328);
xor XOR2 (N9678, N9665, N8941);
nor NOR2 (N9679, N9673, N2935);
buf BUF1 (N9680, N9664);
xor XOR2 (N9681, N9644, N6583);
and AND2 (N9682, N9677, N4593);
and AND3 (N9683, N9674, N264, N8794);
buf BUF1 (N9684, N9679);
nor NOR4 (N9685, N9675, N9354, N8677, N6545);
nand NAND2 (N9686, N9685, N7496);
or OR2 (N9687, N9680, N4923);
nand NAND2 (N9688, N9684, N5694);
nor NOR3 (N9689, N9687, N8339, N4110);
or OR4 (N9690, N9683, N3740, N7075, N8336);
nor NOR2 (N9691, N9682, N2633);
or OR2 (N9692, N9690, N473);
and AND3 (N9693, N9691, N1789, N2896);
xor XOR2 (N9694, N9689, N4781);
not NOT1 (N9695, N9694);
nor NOR2 (N9696, N9666, N8295);
not NOT1 (N9697, N9696);
not NOT1 (N9698, N9678);
nor NOR2 (N9699, N9688, N436);
buf BUF1 (N9700, N9681);
nor NOR4 (N9701, N9699, N4817, N8976, N4227);
nand NAND4 (N9702, N9695, N1467, N5913, N1055);
or OR4 (N9703, N9697, N9440, N8238, N5288);
nor NOR3 (N9704, N9672, N1827, N1353);
or OR4 (N9705, N9701, N4952, N4393, N5622);
nor NOR3 (N9706, N9705, N4903, N6103);
nor NOR2 (N9707, N9676, N8659);
or OR2 (N9708, N9706, N1874);
or OR3 (N9709, N9704, N505, N2493);
nor NOR2 (N9710, N9686, N9543);
not NOT1 (N9711, N9710);
nor NOR4 (N9712, N9702, N6097, N256, N175);
nor NOR4 (N9713, N9708, N8340, N5905, N745);
xor XOR2 (N9714, N9698, N6422);
and AND2 (N9715, N9709, N7624);
and AND3 (N9716, N9713, N7077, N2419);
buf BUF1 (N9717, N9707);
nand NAND4 (N9718, N9711, N4874, N5036, N7287);
nand NAND4 (N9719, N9717, N3390, N4855, N277);
nand NAND3 (N9720, N9715, N7157, N4856);
buf BUF1 (N9721, N9700);
or OR4 (N9722, N9720, N7511, N4385, N3389);
nand NAND3 (N9723, N9693, N6659, N6090);
xor XOR2 (N9724, N9723, N3958);
or OR4 (N9725, N9712, N1998, N1909, N1435);
nand NAND2 (N9726, N9722, N7031);
xor XOR2 (N9727, N9721, N1717);
and AND3 (N9728, N9703, N7338, N7937);
not NOT1 (N9729, N9728);
nand NAND4 (N9730, N9724, N5925, N9547, N8844);
buf BUF1 (N9731, N9718);
buf BUF1 (N9732, N9692);
nor NOR2 (N9733, N9714, N2048);
nand NAND3 (N9734, N9719, N3564, N6828);
buf BUF1 (N9735, N9725);
nand NAND4 (N9736, N9731, N1458, N235, N236);
or OR4 (N9737, N9730, N4979, N5032, N5577);
buf BUF1 (N9738, N9716);
nor NOR4 (N9739, N9736, N1827, N95, N8640);
xor XOR2 (N9740, N9729, N7598);
nor NOR3 (N9741, N9740, N7227, N4867);
not NOT1 (N9742, N9739);
xor XOR2 (N9743, N9735, N3515);
nor NOR3 (N9744, N9726, N9267, N7827);
nor NOR4 (N9745, N9734, N714, N4726, N3572);
nand NAND3 (N9746, N9738, N9189, N6516);
and AND3 (N9747, N9744, N9033, N2028);
buf BUF1 (N9748, N9745);
or OR4 (N9749, N9747, N835, N1901, N9359);
and AND2 (N9750, N9742, N5212);
nand NAND2 (N9751, N9732, N6762);
xor XOR2 (N9752, N9748, N1071);
xor XOR2 (N9753, N9741, N7087);
nor NOR3 (N9754, N9751, N1393, N5247);
xor XOR2 (N9755, N9746, N1087);
and AND4 (N9756, N9749, N8416, N4932, N1744);
and AND3 (N9757, N9756, N5270, N4018);
buf BUF1 (N9758, N9755);
not NOT1 (N9759, N9753);
buf BUF1 (N9760, N9737);
not NOT1 (N9761, N9760);
xor XOR2 (N9762, N9759, N1613);
not NOT1 (N9763, N9752);
nor NOR4 (N9764, N9757, N5439, N708, N9706);
or OR2 (N9765, N9764, N6183);
xor XOR2 (N9766, N9754, N5164);
and AND3 (N9767, N9763, N8476, N8730);
nand NAND3 (N9768, N9761, N3407, N6011);
xor XOR2 (N9769, N9727, N5904);
or OR3 (N9770, N9758, N9230, N67);
not NOT1 (N9771, N9769);
nor NOR4 (N9772, N9770, N5971, N5888, N4472);
not NOT1 (N9773, N9766);
or OR2 (N9774, N9743, N7573);
buf BUF1 (N9775, N9762);
or OR2 (N9776, N9765, N9631);
not NOT1 (N9777, N9771);
nor NOR3 (N9778, N9774, N3586, N4504);
nor NOR3 (N9779, N9767, N9379, N5590);
and AND4 (N9780, N9773, N3014, N561, N274);
not NOT1 (N9781, N9775);
and AND3 (N9782, N9777, N471, N8870);
buf BUF1 (N9783, N9781);
buf BUF1 (N9784, N9776);
and AND3 (N9785, N9784, N9309, N9302);
xor XOR2 (N9786, N9779, N8984);
buf BUF1 (N9787, N9786);
and AND2 (N9788, N9783, N720);
xor XOR2 (N9789, N9782, N1078);
nand NAND3 (N9790, N9785, N990, N9547);
and AND3 (N9791, N9787, N3015, N3985);
xor XOR2 (N9792, N9780, N6550);
not NOT1 (N9793, N9788);
or OR4 (N9794, N9778, N5764, N5872, N5594);
not NOT1 (N9795, N9768);
not NOT1 (N9796, N9750);
and AND2 (N9797, N9733, N323);
buf BUF1 (N9798, N9793);
or OR4 (N9799, N9796, N7216, N7202, N8172);
buf BUF1 (N9800, N9795);
xor XOR2 (N9801, N9790, N6930);
not NOT1 (N9802, N9792);
not NOT1 (N9803, N9802);
nor NOR2 (N9804, N9798, N6150);
buf BUF1 (N9805, N9794);
xor XOR2 (N9806, N9772, N8958);
or OR2 (N9807, N9805, N9014);
not NOT1 (N9808, N9801);
not NOT1 (N9809, N9808);
buf BUF1 (N9810, N9800);
and AND3 (N9811, N9804, N5173, N9469);
nand NAND3 (N9812, N9806, N1318, N8373);
nand NAND3 (N9813, N9797, N4777, N8193);
buf BUF1 (N9814, N9803);
or OR2 (N9815, N9812, N2387);
buf BUF1 (N9816, N9813);
nor NOR2 (N9817, N9810, N7399);
xor XOR2 (N9818, N9817, N3493);
and AND3 (N9819, N9799, N25, N8901);
buf BUF1 (N9820, N9807);
or OR4 (N9821, N9816, N7106, N7678, N4330);
xor XOR2 (N9822, N9809, N2482);
nor NOR3 (N9823, N9815, N6517, N7467);
and AND4 (N9824, N9811, N928, N8076, N1064);
nand NAND3 (N9825, N9818, N3075, N3085);
and AND2 (N9826, N9825, N5610);
not NOT1 (N9827, N9819);
and AND3 (N9828, N9822, N4602, N858);
not NOT1 (N9829, N9814);
not NOT1 (N9830, N9823);
nand NAND3 (N9831, N9827, N5136, N4388);
not NOT1 (N9832, N9821);
nand NAND3 (N9833, N9791, N1334, N303);
or OR4 (N9834, N9832, N9374, N1448, N4819);
or OR2 (N9835, N9831, N2854);
xor XOR2 (N9836, N9828, N4545);
nor NOR3 (N9837, N9829, N8080, N5705);
nor NOR4 (N9838, N9837, N713, N1820, N4632);
nand NAND2 (N9839, N9820, N5582);
not NOT1 (N9840, N9836);
or OR4 (N9841, N9826, N3247, N6180, N986);
and AND4 (N9842, N9833, N2682, N4794, N3345);
nand NAND3 (N9843, N9838, N4763, N5776);
xor XOR2 (N9844, N9834, N7743);
xor XOR2 (N9845, N9843, N2535);
and AND3 (N9846, N9845, N8903, N4192);
and AND4 (N9847, N9789, N1766, N2871, N245);
and AND4 (N9848, N9844, N3927, N4441, N8365);
nor NOR4 (N9849, N9841, N5565, N3152, N4640);
or OR2 (N9850, N9849, N4293);
not NOT1 (N9851, N9846);
and AND2 (N9852, N9847, N2052);
nand NAND3 (N9853, N9848, N680, N2403);
xor XOR2 (N9854, N9850, N4228);
not NOT1 (N9855, N9842);
and AND2 (N9856, N9840, N7566);
nand NAND3 (N9857, N9853, N2442, N1750);
nand NAND2 (N9858, N9852, N8289);
buf BUF1 (N9859, N9856);
xor XOR2 (N9860, N9835, N3028);
buf BUF1 (N9861, N9859);
nand NAND2 (N9862, N9851, N4554);
not NOT1 (N9863, N9861);
not NOT1 (N9864, N9857);
not NOT1 (N9865, N9839);
or OR3 (N9866, N9830, N5432, N1653);
and AND4 (N9867, N9864, N6637, N6668, N8149);
nand NAND2 (N9868, N9855, N7971);
buf BUF1 (N9869, N9866);
or OR4 (N9870, N9858, N2595, N6327, N6269);
not NOT1 (N9871, N9867);
and AND4 (N9872, N9869, N4949, N867, N7892);
or OR2 (N9873, N9824, N309);
or OR2 (N9874, N9862, N1253);
and AND4 (N9875, N9860, N4521, N4929, N7151);
and AND3 (N9876, N9872, N9288, N8286);
buf BUF1 (N9877, N9871);
nor NOR3 (N9878, N9875, N6678, N4003);
nand NAND3 (N9879, N9870, N3746, N2371);
nor NOR4 (N9880, N9854, N2524, N3620, N9612);
xor XOR2 (N9881, N9878, N4040);
or OR4 (N9882, N9868, N7113, N9578, N1022);
and AND3 (N9883, N9876, N9587, N4214);
buf BUF1 (N9884, N9877);
buf BUF1 (N9885, N9879);
xor XOR2 (N9886, N9865, N5409);
buf BUF1 (N9887, N9886);
nand NAND2 (N9888, N9874, N7999);
nand NAND2 (N9889, N9873, N7179);
and AND3 (N9890, N9888, N3124, N7561);
not NOT1 (N9891, N9887);
buf BUF1 (N9892, N9883);
not NOT1 (N9893, N9882);
buf BUF1 (N9894, N9881);
nand NAND3 (N9895, N9893, N2461, N3919);
xor XOR2 (N9896, N9891, N5074);
or OR2 (N9897, N9889, N4378);
buf BUF1 (N9898, N9863);
buf BUF1 (N9899, N9894);
xor XOR2 (N9900, N9880, N8402);
or OR2 (N9901, N9890, N2543);
nand NAND2 (N9902, N9892, N673);
not NOT1 (N9903, N9899);
nor NOR3 (N9904, N9898, N6071, N1788);
xor XOR2 (N9905, N9900, N9695);
xor XOR2 (N9906, N9896, N774);
not NOT1 (N9907, N9903);
or OR2 (N9908, N9906, N444);
and AND3 (N9909, N9905, N4104, N9068);
not NOT1 (N9910, N9908);
not NOT1 (N9911, N9885);
and AND2 (N9912, N9897, N3637);
xor XOR2 (N9913, N9910, N552);
nand NAND2 (N9914, N9904, N2585);
nand NAND3 (N9915, N9914, N4825, N4096);
not NOT1 (N9916, N9913);
or OR4 (N9917, N9884, N167, N9241, N5113);
buf BUF1 (N9918, N9902);
and AND2 (N9919, N9918, N9288);
and AND4 (N9920, N9901, N5685, N926, N8337);
not NOT1 (N9921, N9909);
not NOT1 (N9922, N9895);
or OR3 (N9923, N9907, N7861, N315);
nand NAND4 (N9924, N9916, N3201, N7825, N8658);
or OR4 (N9925, N9923, N9416, N8147, N1198);
nand NAND2 (N9926, N9922, N5157);
xor XOR2 (N9927, N9926, N6691);
buf BUF1 (N9928, N9925);
and AND3 (N9929, N9915, N2797, N6227);
nand NAND3 (N9930, N9929, N2421, N5889);
and AND3 (N9931, N9924, N5663, N4462);
buf BUF1 (N9932, N9912);
xor XOR2 (N9933, N9919, N1271);
nand NAND3 (N9934, N9917, N1059, N1268);
not NOT1 (N9935, N9911);
and AND4 (N9936, N9928, N2240, N96, N8667);
buf BUF1 (N9937, N9933);
not NOT1 (N9938, N9937);
nor NOR2 (N9939, N9927, N3213);
xor XOR2 (N9940, N9931, N3081);
nor NOR4 (N9941, N9930, N3580, N5801, N7);
and AND4 (N9942, N9934, N4243, N9105, N3432);
and AND4 (N9943, N9938, N9483, N6036, N8655);
or OR3 (N9944, N9939, N646, N3661);
or OR3 (N9945, N9944, N8566, N3341);
xor XOR2 (N9946, N9936, N4805);
xor XOR2 (N9947, N9921, N8323);
buf BUF1 (N9948, N9932);
nor NOR2 (N9949, N9945, N9669);
and AND2 (N9950, N9920, N1132);
buf BUF1 (N9951, N9935);
nand NAND4 (N9952, N9947, N3472, N8430, N56);
xor XOR2 (N9953, N9946, N8429);
or OR3 (N9954, N9948, N8804, N2951);
not NOT1 (N9955, N9952);
not NOT1 (N9956, N9951);
or OR2 (N9957, N9941, N9759);
not NOT1 (N9958, N9957);
buf BUF1 (N9959, N9956);
not NOT1 (N9960, N9958);
nor NOR4 (N9961, N9950, N8103, N194, N2199);
buf BUF1 (N9962, N9953);
nand NAND3 (N9963, N9954, N7474, N8332);
xor XOR2 (N9964, N9942, N3493);
nand NAND3 (N9965, N9961, N29, N9002);
and AND3 (N9966, N9959, N8235, N1153);
xor XOR2 (N9967, N9949, N7027);
nor NOR2 (N9968, N9943, N2350);
xor XOR2 (N9969, N9962, N7396);
xor XOR2 (N9970, N9960, N7978);
not NOT1 (N9971, N9940);
buf BUF1 (N9972, N9964);
nor NOR2 (N9973, N9970, N4200);
buf BUF1 (N9974, N9967);
and AND2 (N9975, N9955, N3129);
buf BUF1 (N9976, N9963);
buf BUF1 (N9977, N9972);
not NOT1 (N9978, N9965);
xor XOR2 (N9979, N9974, N5886);
not NOT1 (N9980, N9978);
and AND3 (N9981, N9979, N5149, N8576);
nand NAND2 (N9982, N9980, N2000);
nand NAND3 (N9983, N9977, N3037, N6776);
xor XOR2 (N9984, N9976, N5649);
or OR4 (N9985, N9984, N8352, N476, N1074);
xor XOR2 (N9986, N9981, N6492);
or OR3 (N9987, N9968, N2612, N6564);
and AND2 (N9988, N9985, N3529);
or OR2 (N9989, N9987, N2677);
not NOT1 (N9990, N9983);
not NOT1 (N9991, N9975);
nor NOR3 (N9992, N9971, N6290, N3403);
xor XOR2 (N9993, N9969, N4698);
not NOT1 (N9994, N9973);
or OR4 (N9995, N9994, N6175, N8958, N7751);
or OR3 (N9996, N9991, N1284, N6224);
or OR4 (N9997, N9992, N289, N273, N1253);
and AND4 (N9998, N9988, N8776, N3463, N3561);
or OR3 (N9999, N9966, N4250, N1506);
or OR2 (N10000, N9989, N9135);
and AND3 (N10001, N9990, N1369, N321);
not NOT1 (N10002, N10001);
not NOT1 (N10003, N9982);
or OR2 (N10004, N10003, N283);
nor NOR2 (N10005, N9999, N1081);
not NOT1 (N10006, N10002);
and AND4 (N10007, N9998, N5871, N4937, N7295);
nand NAND4 (N10008, N9997, N11, N9705, N5147);
or OR2 (N10009, N9995, N8102);
nor NOR2 (N10010, N10000, N1898);
nand NAND3 (N10011, N10007, N6310, N5797);
nand NAND4 (N10012, N9996, N8118, N7691, N6489);
or OR2 (N10013, N10004, N1198);
nand NAND3 (N10014, N10009, N6916, N7578);
and AND3 (N10015, N9993, N7178, N3823);
buf BUF1 (N10016, N10005);
buf BUF1 (N10017, N10013);
buf BUF1 (N10018, N10014);
xor XOR2 (N10019, N9986, N6906);
xor XOR2 (N10020, N10008, N8615);
and AND4 (N10021, N10006, N5408, N6453, N6893);
and AND4 (N10022, N10018, N3784, N2454, N5560);
nand NAND2 (N10023, N10019, N71);
and AND4 (N10024, N10023, N8512, N8730, N3363);
buf BUF1 (N10025, N10015);
not NOT1 (N10026, N10010);
nor NOR3 (N10027, N10020, N4169, N6445);
xor XOR2 (N10028, N10027, N2720);
and AND2 (N10029, N10021, N4544);
nor NOR4 (N10030, N10011, N5887, N1677, N9520);
and AND2 (N10031, N10022, N5453);
or OR3 (N10032, N10025, N8901, N9082);
xor XOR2 (N10033, N10032, N2696);
and AND2 (N10034, N10024, N2553);
nor NOR3 (N10035, N10016, N1123, N6785);
buf BUF1 (N10036, N10017);
nor NOR4 (N10037, N10026, N3640, N7247, N2616);
nor NOR4 (N10038, N10035, N9612, N2247, N2861);
nand NAND2 (N10039, N10033, N2821);
nand NAND3 (N10040, N10037, N1497, N8107);
or OR4 (N10041, N10034, N3968, N4798, N9862);
buf BUF1 (N10042, N10028);
nor NOR2 (N10043, N10039, N2456);
not NOT1 (N10044, N10030);
not NOT1 (N10045, N10031);
xor XOR2 (N10046, N10042, N6997);
xor XOR2 (N10047, N10046, N4335);
nor NOR2 (N10048, N10040, N120);
xor XOR2 (N10049, N10029, N5325);
nor NOR4 (N10050, N10012, N7460, N5539, N7805);
xor XOR2 (N10051, N10045, N4397);
nand NAND4 (N10052, N10043, N9771, N9283, N3671);
not NOT1 (N10053, N10047);
nand NAND2 (N10054, N10038, N9714);
not NOT1 (N10055, N10048);
buf BUF1 (N10056, N10036);
not NOT1 (N10057, N10050);
xor XOR2 (N10058, N10049, N4591);
buf BUF1 (N10059, N10053);
or OR2 (N10060, N10059, N7140);
nor NOR4 (N10061, N10055, N8986, N1865, N9477);
and AND2 (N10062, N10041, N7021);
not NOT1 (N10063, N10062);
nand NAND3 (N10064, N10057, N8980, N1978);
buf BUF1 (N10065, N10060);
and AND3 (N10066, N10056, N4456, N4655);
buf BUF1 (N10067, N10066);
buf BUF1 (N10068, N10067);
nor NOR3 (N10069, N10061, N2904, N6558);
and AND3 (N10070, N10065, N7710, N6873);
not NOT1 (N10071, N10058);
nand NAND4 (N10072, N10051, N6115, N943, N9153);
and AND3 (N10073, N10063, N6078, N6648);
and AND3 (N10074, N10071, N9320, N2022);
not NOT1 (N10075, N10069);
not NOT1 (N10076, N10068);
xor XOR2 (N10077, N10072, N3226);
buf BUF1 (N10078, N10054);
and AND2 (N10079, N10078, N5648);
and AND2 (N10080, N10074, N8402);
nor NOR2 (N10081, N10076, N8484);
nand NAND3 (N10082, N10079, N932, N9770);
buf BUF1 (N10083, N10052);
nand NAND3 (N10084, N10080, N8680, N6234);
xor XOR2 (N10085, N10073, N5203);
buf BUF1 (N10086, N10075);
buf BUF1 (N10087, N10086);
or OR4 (N10088, N10077, N7364, N3181, N6775);
nand NAND3 (N10089, N10044, N6055, N6272);
xor XOR2 (N10090, N10083, N1303);
not NOT1 (N10091, N10070);
or OR2 (N10092, N10089, N4747);
buf BUF1 (N10093, N10092);
not NOT1 (N10094, N10085);
or OR4 (N10095, N10093, N3237, N6185, N647);
nor NOR3 (N10096, N10081, N6868, N2467);
nand NAND4 (N10097, N10096, N1076, N1147, N961);
and AND2 (N10098, N10095, N1654);
buf BUF1 (N10099, N10088);
buf BUF1 (N10100, N10098);
nand NAND4 (N10101, N10082, N9215, N6347, N4104);
xor XOR2 (N10102, N10064, N4517);
nor NOR2 (N10103, N10087, N7182);
nand NAND3 (N10104, N10097, N10042, N9479);
or OR4 (N10105, N10104, N8240, N4914, N1842);
nand NAND3 (N10106, N10102, N6515, N8007);
or OR4 (N10107, N10106, N4174, N7910, N1051);
nor NOR2 (N10108, N10101, N5943);
buf BUF1 (N10109, N10100);
xor XOR2 (N10110, N10109, N5384);
not NOT1 (N10111, N10094);
buf BUF1 (N10112, N10108);
and AND2 (N10113, N10107, N4411);
buf BUF1 (N10114, N10111);
nor NOR4 (N10115, N10091, N1596, N2944, N6071);
or OR2 (N10116, N10112, N1499);
and AND3 (N10117, N10113, N3786, N6768);
nand NAND3 (N10118, N10115, N5793, N6307);
not NOT1 (N10119, N10099);
or OR2 (N10120, N10118, N7744);
buf BUF1 (N10121, N10084);
xor XOR2 (N10122, N10110, N326);
and AND2 (N10123, N10121, N2614);
not NOT1 (N10124, N10090);
and AND3 (N10125, N10114, N7940, N3997);
not NOT1 (N10126, N10122);
nand NAND4 (N10127, N10117, N4550, N3934, N3566);
buf BUF1 (N10128, N10124);
and AND3 (N10129, N10120, N6767, N7145);
nor NOR2 (N10130, N10119, N1975);
or OR2 (N10131, N10126, N5955);
xor XOR2 (N10132, N10129, N3217);
not NOT1 (N10133, N10125);
nor NOR2 (N10134, N10127, N2518);
not NOT1 (N10135, N10123);
buf BUF1 (N10136, N10105);
xor XOR2 (N10137, N10133, N5074);
or OR2 (N10138, N10135, N4271);
nand NAND4 (N10139, N10136, N8363, N7529, N8408);
or OR2 (N10140, N10137, N8310);
nor NOR2 (N10141, N10131, N961);
nor NOR3 (N10142, N10103, N6839, N3331);
or OR3 (N10143, N10116, N3301, N9715);
xor XOR2 (N10144, N10141, N6003);
or OR2 (N10145, N10143, N4445);
xor XOR2 (N10146, N10128, N9441);
not NOT1 (N10147, N10140);
nand NAND4 (N10148, N10144, N4817, N1048, N3025);
buf BUF1 (N10149, N10139);
buf BUF1 (N10150, N10148);
not NOT1 (N10151, N10145);
buf BUF1 (N10152, N10147);
or OR2 (N10153, N10149, N40);
buf BUF1 (N10154, N10132);
and AND3 (N10155, N10153, N4793, N6252);
not NOT1 (N10156, N10142);
nor NOR4 (N10157, N10151, N5995, N8921, N7415);
nor NOR4 (N10158, N10157, N8774, N3986, N5227);
nor NOR4 (N10159, N10158, N6160, N6806, N4906);
nor NOR2 (N10160, N10138, N3950);
xor XOR2 (N10161, N10150, N524);
buf BUF1 (N10162, N10160);
and AND3 (N10163, N10154, N3527, N6172);
or OR4 (N10164, N10163, N3966, N5836, N3285);
and AND2 (N10165, N10152, N7857);
nor NOR3 (N10166, N10155, N5651, N2826);
nor NOR2 (N10167, N10161, N6540);
nand NAND4 (N10168, N10167, N6579, N4669, N4892);
not NOT1 (N10169, N10166);
nor NOR2 (N10170, N10162, N9057);
nor NOR4 (N10171, N10169, N1820, N4586, N5746);
nor NOR4 (N10172, N10168, N5693, N4023, N9125);
and AND3 (N10173, N10130, N4372, N2307);
nor NOR2 (N10174, N10164, N5750);
not NOT1 (N10175, N10174);
nand NAND2 (N10176, N10171, N3041);
buf BUF1 (N10177, N10176);
or OR3 (N10178, N10156, N33, N765);
or OR3 (N10179, N10159, N571, N3195);
or OR2 (N10180, N10178, N3084);
and AND3 (N10181, N10175, N8098, N9491);
nor NOR4 (N10182, N10165, N6357, N5207, N8086);
not NOT1 (N10183, N10146);
buf BUF1 (N10184, N10179);
buf BUF1 (N10185, N10134);
not NOT1 (N10186, N10181);
not NOT1 (N10187, N10173);
nand NAND3 (N10188, N10185, N4178, N748);
and AND3 (N10189, N10183, N4468, N7539);
and AND3 (N10190, N10184, N5649, N2415);
nor NOR4 (N10191, N10186, N5170, N6998, N2136);
nand NAND4 (N10192, N10187, N6719, N10162, N5376);
or OR4 (N10193, N10189, N115, N7420, N2157);
buf BUF1 (N10194, N10193);
not NOT1 (N10195, N10172);
xor XOR2 (N10196, N10182, N4690);
nor NOR2 (N10197, N10180, N7189);
buf BUF1 (N10198, N10197);
and AND3 (N10199, N10191, N2103, N9571);
nor NOR2 (N10200, N10198, N7122);
and AND4 (N10201, N10190, N5702, N5360, N9268);
nor NOR2 (N10202, N10196, N9007);
not NOT1 (N10203, N10199);
xor XOR2 (N10204, N10177, N4595);
and AND4 (N10205, N10202, N4759, N6449, N5115);
not NOT1 (N10206, N10195);
nand NAND2 (N10207, N10200, N4209);
not NOT1 (N10208, N10194);
nor NOR3 (N10209, N10206, N5613, N3406);
xor XOR2 (N10210, N10204, N7855);
and AND2 (N10211, N10210, N9690);
nand NAND3 (N10212, N10211, N9607, N6039);
nor NOR2 (N10213, N10208, N7557);
or OR4 (N10214, N10188, N9381, N6694, N4869);
nand NAND4 (N10215, N10203, N6895, N3975, N4825);
or OR2 (N10216, N10205, N3561);
not NOT1 (N10217, N10192);
or OR2 (N10218, N10170, N4944);
not NOT1 (N10219, N10216);
buf BUF1 (N10220, N10207);
not NOT1 (N10221, N10213);
nand NAND3 (N10222, N10219, N1741, N7614);
or OR3 (N10223, N10221, N6618, N7866);
and AND2 (N10224, N10215, N8168);
xor XOR2 (N10225, N10220, N5164);
xor XOR2 (N10226, N10224, N1585);
buf BUF1 (N10227, N10218);
or OR3 (N10228, N10217, N5936, N5684);
nor NOR4 (N10229, N10227, N9120, N1175, N5663);
nor NOR2 (N10230, N10223, N2201);
nor NOR3 (N10231, N10214, N2112, N3310);
and AND4 (N10232, N10231, N10045, N4564, N7734);
and AND2 (N10233, N10226, N9445);
and AND3 (N10234, N10229, N10181, N2057);
buf BUF1 (N10235, N10209);
buf BUF1 (N10236, N10222);
not NOT1 (N10237, N10233);
nor NOR4 (N10238, N10237, N8861, N4628, N906);
nor NOR3 (N10239, N10234, N7439, N6828);
or OR3 (N10240, N10235, N6596, N6456);
and AND4 (N10241, N10228, N8245, N9092, N8404);
buf BUF1 (N10242, N10236);
buf BUF1 (N10243, N10238);
xor XOR2 (N10244, N10239, N10210);
not NOT1 (N10245, N10240);
not NOT1 (N10246, N10244);
not NOT1 (N10247, N10241);
nor NOR3 (N10248, N10247, N6707, N918);
or OR2 (N10249, N10242, N1017);
or OR3 (N10250, N10232, N7915, N2013);
nand NAND3 (N10251, N10250, N6588, N9993);
and AND3 (N10252, N10246, N1986, N7898);
buf BUF1 (N10253, N10230);
and AND2 (N10254, N10252, N4504);
or OR2 (N10255, N10251, N7846);
xor XOR2 (N10256, N10254, N1809);
xor XOR2 (N10257, N10245, N1646);
nor NOR2 (N10258, N10243, N2741);
and AND2 (N10259, N10225, N4895);
xor XOR2 (N10260, N10248, N2554);
and AND4 (N10261, N10260, N1144, N8453, N6985);
nor NOR4 (N10262, N10259, N2396, N4813, N9414);
nand NAND2 (N10263, N10257, N9746);
nor NOR3 (N10264, N10255, N7814, N785);
nor NOR4 (N10265, N10263, N1145, N4166, N2081);
buf BUF1 (N10266, N10262);
nand NAND3 (N10267, N10212, N6081, N2016);
xor XOR2 (N10268, N10253, N10214);
and AND2 (N10269, N10261, N6303);
nor NOR2 (N10270, N10258, N5644);
and AND4 (N10271, N10269, N4631, N6105, N2419);
nor NOR3 (N10272, N10249, N7131, N6906);
buf BUF1 (N10273, N10271);
nand NAND2 (N10274, N10265, N4963);
not NOT1 (N10275, N10256);
nand NAND3 (N10276, N10274, N7476, N4183);
xor XOR2 (N10277, N10276, N5448);
or OR4 (N10278, N10273, N4522, N3114, N600);
or OR3 (N10279, N10266, N9678, N245);
and AND2 (N10280, N10272, N9171);
buf BUF1 (N10281, N10264);
xor XOR2 (N10282, N10277, N8233);
nor NOR2 (N10283, N10268, N2193);
nor NOR3 (N10284, N10201, N2045, N8684);
not NOT1 (N10285, N10267);
buf BUF1 (N10286, N10284);
or OR2 (N10287, N10281, N3059);
nand NAND2 (N10288, N10285, N1215);
nand NAND4 (N10289, N10288, N8828, N6468, N1078);
nor NOR3 (N10290, N10278, N2172, N3739);
nand NAND4 (N10291, N10286, N8302, N4217, N6041);
and AND2 (N10292, N10291, N9195);
xor XOR2 (N10293, N10290, N8356);
and AND2 (N10294, N10279, N5055);
or OR2 (N10295, N10280, N4760);
xor XOR2 (N10296, N10275, N78);
and AND2 (N10297, N10292, N1031);
not NOT1 (N10298, N10282);
nor NOR2 (N10299, N10295, N10173);
buf BUF1 (N10300, N10270);
buf BUF1 (N10301, N10289);
nor NOR4 (N10302, N10297, N3698, N8766, N339);
not NOT1 (N10303, N10294);
and AND3 (N10304, N10293, N5136, N8761);
and AND4 (N10305, N10304, N9139, N1369, N7783);
nor NOR2 (N10306, N10287, N9836);
nor NOR2 (N10307, N10283, N3499);
buf BUF1 (N10308, N10300);
not NOT1 (N10309, N10298);
or OR4 (N10310, N10308, N6722, N3413, N7719);
nand NAND3 (N10311, N10301, N7039, N4028);
nor NOR2 (N10312, N10306, N7253);
or OR2 (N10313, N10305, N2303);
nand NAND4 (N10314, N10313, N2740, N738, N6743);
not NOT1 (N10315, N10311);
or OR3 (N10316, N10315, N2523, N4070);
or OR3 (N10317, N10310, N1538, N6454);
nor NOR2 (N10318, N10314, N7075);
nor NOR3 (N10319, N10317, N6891, N8330);
xor XOR2 (N10320, N10319, N4843);
nor NOR4 (N10321, N10299, N8415, N4686, N4894);
nor NOR3 (N10322, N10309, N10279, N5195);
buf BUF1 (N10323, N10316);
and AND2 (N10324, N10320, N9895);
xor XOR2 (N10325, N10321, N6628);
or OR3 (N10326, N10312, N5895, N5817);
and AND4 (N10327, N10325, N2762, N539, N6126);
not NOT1 (N10328, N10318);
and AND2 (N10329, N10296, N8019);
and AND4 (N10330, N10324, N1224, N3165, N7788);
or OR2 (N10331, N10323, N7898);
or OR4 (N10332, N10328, N3046, N8384, N58);
xor XOR2 (N10333, N10327, N4563);
and AND4 (N10334, N10331, N5442, N7068, N2472);
nor NOR3 (N10335, N10330, N8643, N4145);
nor NOR2 (N10336, N10302, N18);
xor XOR2 (N10337, N10332, N2777);
or OR4 (N10338, N10337, N9987, N1390, N7298);
nand NAND2 (N10339, N10303, N5265);
buf BUF1 (N10340, N10329);
or OR4 (N10341, N10307, N1759, N5730, N10040);
nor NOR3 (N10342, N10335, N5950, N5687);
xor XOR2 (N10343, N10333, N6560);
buf BUF1 (N10344, N10340);
not NOT1 (N10345, N10341);
xor XOR2 (N10346, N10336, N5187);
nor NOR4 (N10347, N10326, N6741, N356, N1566);
xor XOR2 (N10348, N10322, N2788);
nand NAND4 (N10349, N10343, N4814, N2989, N7630);
xor XOR2 (N10350, N10347, N5621);
nor NOR4 (N10351, N10338, N4694, N99, N8859);
xor XOR2 (N10352, N10351, N8869);
xor XOR2 (N10353, N10349, N3144);
nor NOR3 (N10354, N10334, N13, N3825);
and AND3 (N10355, N10350, N8020, N329);
buf BUF1 (N10356, N10339);
or OR4 (N10357, N10354, N6292, N1041, N5280);
buf BUF1 (N10358, N10355);
xor XOR2 (N10359, N10346, N9611);
buf BUF1 (N10360, N10348);
buf BUF1 (N10361, N10356);
not NOT1 (N10362, N10352);
buf BUF1 (N10363, N10360);
not NOT1 (N10364, N10357);
and AND3 (N10365, N10363, N3580, N449);
nand NAND2 (N10366, N10344, N9570);
nor NOR3 (N10367, N10359, N1673, N6922);
or OR2 (N10368, N10358, N8989);
and AND3 (N10369, N10342, N5014, N6380);
nor NOR3 (N10370, N10365, N6747, N9016);
xor XOR2 (N10371, N10367, N3754);
nand NAND3 (N10372, N10362, N10187, N339);
or OR3 (N10373, N10370, N10235, N2010);
nand NAND4 (N10374, N10371, N9474, N7432, N3538);
nand NAND4 (N10375, N10364, N2193, N1255, N9822);
not NOT1 (N10376, N10369);
nor NOR2 (N10377, N10345, N5058);
not NOT1 (N10378, N10377);
or OR3 (N10379, N10353, N10052, N686);
xor XOR2 (N10380, N10375, N7697);
nor NOR2 (N10381, N10373, N6638);
or OR2 (N10382, N10368, N4660);
xor XOR2 (N10383, N10378, N5023);
not NOT1 (N10384, N10361);
nor NOR2 (N10385, N10381, N8509);
buf BUF1 (N10386, N10383);
buf BUF1 (N10387, N10384);
nand NAND2 (N10388, N10372, N8651);
or OR2 (N10389, N10387, N10100);
or OR2 (N10390, N10380, N821);
buf BUF1 (N10391, N10374);
xor XOR2 (N10392, N10366, N7113);
xor XOR2 (N10393, N10390, N5087);
buf BUF1 (N10394, N10379);
nand NAND3 (N10395, N10385, N3061, N7557);
nand NAND3 (N10396, N10392, N9503, N8299);
and AND4 (N10397, N10391, N226, N3569, N9261);
xor XOR2 (N10398, N10393, N942);
or OR3 (N10399, N10395, N9963, N1919);
nand NAND4 (N10400, N10399, N721, N7601, N534);
xor XOR2 (N10401, N10400, N9266);
not NOT1 (N10402, N10376);
not NOT1 (N10403, N10397);
nand NAND4 (N10404, N10386, N732, N9329, N1105);
and AND2 (N10405, N10389, N4471);
and AND2 (N10406, N10404, N3486);
or OR3 (N10407, N10403, N4202, N8433);
xor XOR2 (N10408, N10394, N9090);
nand NAND2 (N10409, N10398, N6466);
or OR2 (N10410, N10405, N4379);
nor NOR2 (N10411, N10410, N3192);
and AND2 (N10412, N10382, N5610);
and AND2 (N10413, N10409, N5951);
and AND4 (N10414, N10412, N9088, N1462, N62);
xor XOR2 (N10415, N10401, N9679);
buf BUF1 (N10416, N10408);
or OR4 (N10417, N10416, N5248, N1962, N6974);
not NOT1 (N10418, N10396);
nor NOR3 (N10419, N10388, N7920, N8857);
and AND3 (N10420, N10402, N5796, N8763);
or OR4 (N10421, N10407, N43, N3527, N8968);
nor NOR2 (N10422, N10414, N5209);
nand NAND2 (N10423, N10419, N6455);
and AND2 (N10424, N10415, N10187);
nand NAND3 (N10425, N10423, N1930, N8724);
and AND3 (N10426, N10421, N4805, N157);
buf BUF1 (N10427, N10426);
nor NOR3 (N10428, N10420, N3108, N1006);
or OR4 (N10429, N10428, N4689, N2255, N6994);
nor NOR3 (N10430, N10417, N369, N8050);
and AND3 (N10431, N10413, N7024, N1343);
buf BUF1 (N10432, N10431);
xor XOR2 (N10433, N10432, N8273);
not NOT1 (N10434, N10424);
nor NOR4 (N10435, N10427, N2053, N7833, N8348);
xor XOR2 (N10436, N10429, N8804);
and AND2 (N10437, N10434, N4382);
and AND4 (N10438, N10435, N7948, N3265, N7154);
not NOT1 (N10439, N10425);
nor NOR3 (N10440, N10430, N398, N216);
xor XOR2 (N10441, N10439, N1924);
and AND3 (N10442, N10436, N4208, N6177);
and AND3 (N10443, N10422, N5250, N6416);
or OR3 (N10444, N10437, N9935, N8716);
nor NOR2 (N10445, N10411, N1971);
xor XOR2 (N10446, N10444, N9244);
not NOT1 (N10447, N10446);
not NOT1 (N10448, N10441);
buf BUF1 (N10449, N10433);
nand NAND2 (N10450, N10442, N8758);
not NOT1 (N10451, N10449);
nand NAND3 (N10452, N10448, N2136, N7903);
or OR3 (N10453, N10450, N2796, N5349);
not NOT1 (N10454, N10445);
buf BUF1 (N10455, N10438);
nand NAND3 (N10456, N10454, N5678, N8679);
and AND4 (N10457, N10453, N2251, N4662, N5496);
not NOT1 (N10458, N10406);
nor NOR3 (N10459, N10440, N4288, N3555);
buf BUF1 (N10460, N10457);
and AND3 (N10461, N10458, N1302, N10132);
nor NOR3 (N10462, N10443, N1842, N2891);
xor XOR2 (N10463, N10447, N6568);
nand NAND3 (N10464, N10452, N10252, N369);
or OR2 (N10465, N10461, N5745);
buf BUF1 (N10466, N10463);
or OR3 (N10467, N10465, N1365, N3476);
nand NAND3 (N10468, N10467, N2213, N7885);
not NOT1 (N10469, N10466);
or OR3 (N10470, N10468, N5756, N1685);
nor NOR4 (N10471, N10451, N9175, N1395, N6120);
xor XOR2 (N10472, N10460, N1395);
nand NAND3 (N10473, N10469, N2757, N8614);
nor NOR3 (N10474, N10472, N3226, N9408);
or OR3 (N10475, N10456, N753, N4550);
or OR2 (N10476, N10464, N7500);
nand NAND2 (N10477, N10476, N10327);
and AND4 (N10478, N10462, N9593, N10239, N8623);
nand NAND3 (N10479, N10471, N5306, N5436);
xor XOR2 (N10480, N10473, N1678);
or OR2 (N10481, N10479, N9773);
and AND2 (N10482, N10475, N3332);
nor NOR2 (N10483, N10418, N1138);
buf BUF1 (N10484, N10455);
xor XOR2 (N10485, N10478, N7184);
and AND2 (N10486, N10485, N8146);
nand NAND4 (N10487, N10481, N1992, N8477, N653);
nor NOR3 (N10488, N10482, N10400, N8214);
and AND2 (N10489, N10470, N9206);
not NOT1 (N10490, N10483);
nand NAND3 (N10491, N10459, N5100, N5771);
or OR2 (N10492, N10480, N2046);
or OR2 (N10493, N10491, N5078);
nor NOR2 (N10494, N10488, N1807);
buf BUF1 (N10495, N10484);
not NOT1 (N10496, N10493);
buf BUF1 (N10497, N10474);
buf BUF1 (N10498, N10496);
not NOT1 (N10499, N10490);
buf BUF1 (N10500, N10497);
xor XOR2 (N10501, N10486, N5339);
nor NOR4 (N10502, N10494, N1315, N9174, N269);
and AND4 (N10503, N10499, N3692, N2791, N3281);
and AND4 (N10504, N10489, N6280, N5100, N2956);
and AND3 (N10505, N10501, N1785, N2906);
xor XOR2 (N10506, N10495, N6188);
nor NOR3 (N10507, N10502, N5262, N6037);
nand NAND4 (N10508, N10477, N3241, N8708, N2162);
nand NAND2 (N10509, N10506, N6904);
or OR4 (N10510, N10507, N6299, N3045, N3023);
nor NOR2 (N10511, N10510, N8041);
and AND2 (N10512, N10503, N3919);
not NOT1 (N10513, N10498);
and AND4 (N10514, N10492, N4587, N1046, N2246);
or OR2 (N10515, N10511, N6746);
nand NAND2 (N10516, N10509, N8356);
not NOT1 (N10517, N10516);
and AND4 (N10518, N10487, N3290, N2000, N7181);
not NOT1 (N10519, N10517);
or OR3 (N10520, N10518, N5845, N7807);
xor XOR2 (N10521, N10514, N8608);
nor NOR4 (N10522, N10521, N5577, N1286, N8546);
or OR2 (N10523, N10500, N2421);
and AND3 (N10524, N10504, N8690, N2356);
buf BUF1 (N10525, N10523);
nor NOR2 (N10526, N10515, N6630);
nand NAND2 (N10527, N10508, N2246);
nand NAND2 (N10528, N10505, N4833);
and AND4 (N10529, N10527, N1257, N1393, N3331);
buf BUF1 (N10530, N10525);
and AND3 (N10531, N10512, N9314, N10085);
nor NOR2 (N10532, N10529, N4250);
buf BUF1 (N10533, N10530);
or OR3 (N10534, N10528, N6287, N9385);
and AND2 (N10535, N10522, N2544);
and AND4 (N10536, N10535, N5499, N9520, N802);
nand NAND4 (N10537, N10526, N7388, N9148, N5406);
not NOT1 (N10538, N10533);
nand NAND3 (N10539, N10536, N8226, N6710);
buf BUF1 (N10540, N10539);
and AND2 (N10541, N10531, N10475);
and AND2 (N10542, N10524, N7925);
xor XOR2 (N10543, N10532, N7578);
nand NAND4 (N10544, N10540, N9820, N3740, N3057);
nor NOR3 (N10545, N10543, N6347, N271);
nor NOR2 (N10546, N10542, N7006);
or OR3 (N10547, N10519, N5838, N7298);
buf BUF1 (N10548, N10537);
nor NOR2 (N10549, N10534, N3723);
or OR3 (N10550, N10544, N288, N8060);
or OR3 (N10551, N10546, N4007, N9831);
and AND4 (N10552, N10541, N7946, N8319, N4603);
nand NAND3 (N10553, N10513, N6007, N5475);
xor XOR2 (N10554, N10553, N1673);
or OR3 (N10555, N10554, N9777, N1467);
and AND3 (N10556, N10545, N10425, N6306);
nor NOR3 (N10557, N10552, N7907, N6855);
nor NOR2 (N10558, N10551, N1644);
nand NAND4 (N10559, N10556, N10305, N7347, N8604);
nor NOR4 (N10560, N10548, N2835, N555, N1490);
nor NOR4 (N10561, N10520, N756, N789, N9675);
nand NAND4 (N10562, N10550, N4292, N6486, N3246);
nor NOR3 (N10563, N10547, N3292, N5673);
xor XOR2 (N10564, N10538, N4131);
nand NAND2 (N10565, N10558, N7355);
xor XOR2 (N10566, N10564, N6042);
buf BUF1 (N10567, N10563);
nand NAND2 (N10568, N10565, N3584);
not NOT1 (N10569, N10560);
nand NAND2 (N10570, N10566, N544);
buf BUF1 (N10571, N10561);
nor NOR2 (N10572, N10562, N6813);
nor NOR3 (N10573, N10555, N1670, N5697);
nand NAND4 (N10574, N10572, N5239, N5891, N7003);
buf BUF1 (N10575, N10574);
not NOT1 (N10576, N10568);
nor NOR2 (N10577, N10559, N166);
or OR3 (N10578, N10557, N4676, N10547);
and AND4 (N10579, N10575, N9303, N8015, N5994);
and AND2 (N10580, N10569, N5451);
not NOT1 (N10581, N10573);
nand NAND2 (N10582, N10567, N259);
nor NOR4 (N10583, N10570, N8927, N583, N50);
nor NOR2 (N10584, N10571, N4427);
not NOT1 (N10585, N10576);
and AND4 (N10586, N10579, N9848, N5005, N1814);
and AND4 (N10587, N10578, N3830, N6410, N7218);
nand NAND4 (N10588, N10583, N8055, N4778, N3062);
or OR3 (N10589, N10581, N1289, N3789);
not NOT1 (N10590, N10586);
and AND3 (N10591, N10587, N6680, N1291);
not NOT1 (N10592, N10580);
not NOT1 (N10593, N10592);
buf BUF1 (N10594, N10591);
or OR2 (N10595, N10584, N5362);
not NOT1 (N10596, N10594);
nor NOR2 (N10597, N10585, N1716);
buf BUF1 (N10598, N10589);
not NOT1 (N10599, N10596);
nor NOR4 (N10600, N10599, N10360, N5587, N1745);
xor XOR2 (N10601, N10593, N3036);
buf BUF1 (N10602, N10577);
buf BUF1 (N10603, N10549);
xor XOR2 (N10604, N10602, N562);
nand NAND4 (N10605, N10582, N9988, N1578, N1483);
and AND3 (N10606, N10600, N9337, N1785);
buf BUF1 (N10607, N10598);
nor NOR4 (N10608, N10601, N2475, N2251, N2651);
nor NOR2 (N10609, N10605, N10382);
buf BUF1 (N10610, N10595);
not NOT1 (N10611, N10606);
nor NOR4 (N10612, N10588, N2594, N7519, N6527);
xor XOR2 (N10613, N10609, N4190);
buf BUF1 (N10614, N10604);
nor NOR2 (N10615, N10608, N4007);
buf BUF1 (N10616, N10614);
not NOT1 (N10617, N10615);
nor NOR4 (N10618, N10607, N4942, N2111, N7015);
buf BUF1 (N10619, N10590);
and AND4 (N10620, N10597, N6246, N10165, N6902);
nand NAND2 (N10621, N10611, N581);
nand NAND2 (N10622, N10603, N260);
nor NOR2 (N10623, N10617, N4485);
or OR3 (N10624, N10622, N9496, N9263);
not NOT1 (N10625, N10619);
not NOT1 (N10626, N10624);
and AND3 (N10627, N10620, N7873, N4889);
nor NOR3 (N10628, N10623, N3375, N8718);
nand NAND4 (N10629, N10628, N8311, N6271, N3308);
and AND4 (N10630, N10618, N1638, N10393, N6309);
buf BUF1 (N10631, N10621);
nor NOR4 (N10632, N10613, N7640, N2768, N4069);
not NOT1 (N10633, N10610);
and AND2 (N10634, N10616, N8078);
nand NAND2 (N10635, N10629, N4044);
nand NAND3 (N10636, N10635, N9732, N7051);
or OR2 (N10637, N10627, N2380);
nand NAND4 (N10638, N10626, N3494, N3945, N59);
or OR4 (N10639, N10625, N4577, N7096, N3826);
not NOT1 (N10640, N10633);
not NOT1 (N10641, N10612);
nor NOR2 (N10642, N10640, N5399);
or OR3 (N10643, N10630, N10564, N2683);
nor NOR2 (N10644, N10638, N2947);
or OR2 (N10645, N10634, N8262);
nor NOR3 (N10646, N10639, N1453, N8647);
xor XOR2 (N10647, N10637, N8021);
and AND4 (N10648, N10631, N4001, N4734, N5396);
or OR4 (N10649, N10644, N2754, N10511, N10086);
nor NOR4 (N10650, N10632, N10508, N7246, N5278);
and AND3 (N10651, N10643, N5413, N10405);
and AND2 (N10652, N10649, N6100);
not NOT1 (N10653, N10652);
buf BUF1 (N10654, N10636);
nor NOR3 (N10655, N10646, N8270, N9613);
xor XOR2 (N10656, N10641, N4062);
xor XOR2 (N10657, N10650, N810);
or OR4 (N10658, N10645, N2170, N3395, N6436);
xor XOR2 (N10659, N10647, N3834);
or OR4 (N10660, N10659, N8517, N10481, N7078);
and AND4 (N10661, N10660, N10108, N7298, N4663);
not NOT1 (N10662, N10642);
buf BUF1 (N10663, N10661);
nand NAND3 (N10664, N10653, N4968, N481);
nor NOR2 (N10665, N10662, N7653);
nand NAND2 (N10666, N10654, N4866);
not NOT1 (N10667, N10656);
or OR2 (N10668, N10648, N8674);
or OR4 (N10669, N10667, N2222, N802, N6589);
nor NOR2 (N10670, N10663, N9481);
nor NOR2 (N10671, N10670, N7298);
buf BUF1 (N10672, N10658);
nor NOR4 (N10673, N10665, N6210, N3717, N1489);
xor XOR2 (N10674, N10669, N307);
buf BUF1 (N10675, N10671);
not NOT1 (N10676, N10672);
buf BUF1 (N10677, N10651);
and AND4 (N10678, N10664, N3621, N7234, N7044);
or OR4 (N10679, N10677, N10229, N6684, N4976);
buf BUF1 (N10680, N10668);
buf BUF1 (N10681, N10666);
and AND2 (N10682, N10674, N1385);
buf BUF1 (N10683, N10676);
and AND3 (N10684, N10675, N9341, N5872);
not NOT1 (N10685, N10655);
nand NAND3 (N10686, N10657, N1537, N1528);
and AND4 (N10687, N10684, N2240, N10516, N3081);
or OR2 (N10688, N10686, N4819);
not NOT1 (N10689, N10687);
buf BUF1 (N10690, N10673);
xor XOR2 (N10691, N10683, N4687);
xor XOR2 (N10692, N10678, N9333);
and AND2 (N10693, N10681, N3940);
or OR4 (N10694, N10682, N2976, N722, N4936);
nor NOR3 (N10695, N10689, N6332, N9119);
buf BUF1 (N10696, N10693);
buf BUF1 (N10697, N10691);
buf BUF1 (N10698, N10679);
not NOT1 (N10699, N10695);
nor NOR2 (N10700, N10688, N1564);
buf BUF1 (N10701, N10698);
buf BUF1 (N10702, N10696);
not NOT1 (N10703, N10699);
nor NOR4 (N10704, N10694, N7122, N1155, N3396);
or OR4 (N10705, N10700, N5949, N4508, N4968);
or OR3 (N10706, N10692, N4166, N6217);
buf BUF1 (N10707, N10703);
and AND2 (N10708, N10707, N8349);
not NOT1 (N10709, N10705);
xor XOR2 (N10710, N10709, N8435);
nand NAND2 (N10711, N10701, N10502);
not NOT1 (N10712, N10690);
or OR2 (N10713, N10697, N4750);
and AND2 (N10714, N10685, N4832);
nand NAND2 (N10715, N10702, N7335);
xor XOR2 (N10716, N10708, N5068);
or OR2 (N10717, N10706, N3397);
xor XOR2 (N10718, N10704, N9557);
or OR3 (N10719, N10711, N9602, N8716);
and AND4 (N10720, N10719, N3942, N4194, N3594);
xor XOR2 (N10721, N10714, N9720);
and AND3 (N10722, N10721, N1471, N5637);
buf BUF1 (N10723, N10722);
or OR2 (N10724, N10715, N10459);
xor XOR2 (N10725, N10720, N1634);
nor NOR3 (N10726, N10725, N5436, N3311);
or OR4 (N10727, N10680, N7058, N9552, N5440);
xor XOR2 (N10728, N10717, N9811);
nor NOR3 (N10729, N10723, N2601, N9975);
nor NOR2 (N10730, N10713, N1146);
nand NAND3 (N10731, N10730, N6913, N545);
xor XOR2 (N10732, N10726, N5602);
and AND3 (N10733, N10728, N1197, N8566);
or OR3 (N10734, N10716, N2282, N6888);
buf BUF1 (N10735, N10733);
xor XOR2 (N10736, N10727, N6348);
xor XOR2 (N10737, N10732, N5951);
nor NOR2 (N10738, N10724, N3653);
and AND3 (N10739, N10718, N3138, N10487);
or OR2 (N10740, N10739, N10691);
and AND2 (N10741, N10737, N4134);
or OR4 (N10742, N10741, N7671, N7462, N9803);
nand NAND2 (N10743, N10738, N2773);
nand NAND2 (N10744, N10743, N9066);
or OR2 (N10745, N10736, N8564);
or OR2 (N10746, N10740, N9309);
nand NAND2 (N10747, N10710, N9155);
nor NOR2 (N10748, N10744, N7141);
xor XOR2 (N10749, N10745, N8711);
and AND2 (N10750, N10729, N9033);
or OR4 (N10751, N10734, N1544, N432, N7045);
nand NAND2 (N10752, N10751, N913);
nor NOR2 (N10753, N10731, N5568);
xor XOR2 (N10754, N10753, N1754);
nand NAND3 (N10755, N10735, N10200, N3710);
and AND2 (N10756, N10746, N6661);
nor NOR3 (N10757, N10752, N9344, N9332);
buf BUF1 (N10758, N10712);
nand NAND3 (N10759, N10742, N6671, N10600);
buf BUF1 (N10760, N10755);
xor XOR2 (N10761, N10750, N4731);
and AND3 (N10762, N10754, N5205, N1097);
buf BUF1 (N10763, N10749);
xor XOR2 (N10764, N10757, N4329);
buf BUF1 (N10765, N10756);
buf BUF1 (N10766, N10761);
and AND2 (N10767, N10762, N7736);
nand NAND2 (N10768, N10764, N8791);
buf BUF1 (N10769, N10748);
nand NAND2 (N10770, N10759, N6377);
buf BUF1 (N10771, N10768);
and AND3 (N10772, N10771, N10531, N8729);
xor XOR2 (N10773, N10767, N1303);
buf BUF1 (N10774, N10769);
nand NAND4 (N10775, N10760, N1848, N3381, N6486);
xor XOR2 (N10776, N10765, N9890);
and AND2 (N10777, N10766, N64);
nand NAND3 (N10778, N10770, N4076, N7598);
xor XOR2 (N10779, N10747, N7417);
nand NAND2 (N10780, N10777, N487);
nor NOR2 (N10781, N10780, N2122);
and AND4 (N10782, N10779, N3470, N2839, N4506);
buf BUF1 (N10783, N10775);
nor NOR2 (N10784, N10778, N3);
buf BUF1 (N10785, N10772);
or OR4 (N10786, N10763, N3315, N402, N12);
and AND2 (N10787, N10781, N604);
and AND3 (N10788, N10783, N10543, N9998);
xor XOR2 (N10789, N10784, N3477);
or OR2 (N10790, N10758, N756);
nand NAND3 (N10791, N10782, N8678, N1542);
not NOT1 (N10792, N10787);
not NOT1 (N10793, N10789);
or OR4 (N10794, N10791, N3080, N3130, N10771);
nor NOR3 (N10795, N10786, N4317, N1520);
nand NAND4 (N10796, N10793, N10516, N2309, N7856);
and AND4 (N10797, N10785, N9630, N6238, N3053);
and AND4 (N10798, N10792, N7256, N10144, N6380);
or OR4 (N10799, N10790, N7707, N8876, N4392);
or OR4 (N10800, N10774, N4129, N10193, N4004);
buf BUF1 (N10801, N10800);
or OR2 (N10802, N10795, N9600);
xor XOR2 (N10803, N10797, N233);
not NOT1 (N10804, N10776);
xor XOR2 (N10805, N10798, N9093);
nand NAND4 (N10806, N10805, N3645, N10469, N1079);
buf BUF1 (N10807, N10799);
xor XOR2 (N10808, N10794, N8187);
buf BUF1 (N10809, N10801);
or OR3 (N10810, N10807, N3632, N4460);
buf BUF1 (N10811, N10808);
and AND2 (N10812, N10810, N10586);
nand NAND3 (N10813, N10788, N8830, N5582);
nand NAND2 (N10814, N10811, N1897);
not NOT1 (N10815, N10802);
nand NAND2 (N10816, N10812, N3561);
not NOT1 (N10817, N10803);
or OR3 (N10818, N10806, N1366, N5453);
not NOT1 (N10819, N10796);
buf BUF1 (N10820, N10813);
and AND4 (N10821, N10818, N7256, N6884, N382);
not NOT1 (N10822, N10821);
or OR2 (N10823, N10817, N284);
and AND2 (N10824, N10815, N7860);
not NOT1 (N10825, N10816);
nor NOR4 (N10826, N10820, N6389, N6085, N9594);
xor XOR2 (N10827, N10814, N8359);
not NOT1 (N10828, N10819);
and AND2 (N10829, N10825, N5809);
buf BUF1 (N10830, N10824);
nand NAND3 (N10831, N10773, N3920, N9421);
xor XOR2 (N10832, N10809, N6424);
xor XOR2 (N10833, N10804, N913);
nand NAND4 (N10834, N10828, N7429, N8615, N6129);
xor XOR2 (N10835, N10832, N6588);
buf BUF1 (N10836, N10831);
nor NOR4 (N10837, N10829, N8343, N2090, N8222);
nor NOR2 (N10838, N10827, N837);
or OR3 (N10839, N10822, N4631, N2318);
or OR2 (N10840, N10837, N8254);
nand NAND3 (N10841, N10839, N3267, N9029);
and AND2 (N10842, N10835, N53);
buf BUF1 (N10843, N10838);
nor NOR4 (N10844, N10834, N10816, N6377, N6315);
buf BUF1 (N10845, N10836);
nand NAND3 (N10846, N10842, N7519, N10136);
or OR4 (N10847, N10830, N8470, N6842, N7640);
buf BUF1 (N10848, N10843);
and AND3 (N10849, N10841, N5727, N10306);
and AND2 (N10850, N10847, N9435);
and AND2 (N10851, N10826, N7473);
or OR4 (N10852, N10849, N5642, N5226, N2026);
not NOT1 (N10853, N10850);
nor NOR3 (N10854, N10844, N4197, N5400);
or OR2 (N10855, N10852, N2934);
xor XOR2 (N10856, N10840, N8239);
or OR3 (N10857, N10845, N5455, N2118);
nor NOR4 (N10858, N10855, N9314, N7161, N1671);
nor NOR3 (N10859, N10857, N3989, N7403);
nor NOR2 (N10860, N10858, N6201);
and AND4 (N10861, N10833, N6571, N3283, N2054);
nand NAND4 (N10862, N10856, N6896, N2610, N9151);
nand NAND2 (N10863, N10848, N1331);
nand NAND4 (N10864, N10823, N3270, N6733, N7827);
or OR3 (N10865, N10860, N5287, N10280);
buf BUF1 (N10866, N10853);
nand NAND4 (N10867, N10862, N8292, N1202, N3872);
buf BUF1 (N10868, N10854);
not NOT1 (N10869, N10846);
not NOT1 (N10870, N10863);
nor NOR4 (N10871, N10851, N8668, N8772, N844);
nor NOR3 (N10872, N10868, N5778, N8438);
nand NAND4 (N10873, N10864, N5575, N2147, N5811);
buf BUF1 (N10874, N10869);
nor NOR3 (N10875, N10866, N3827, N6518);
not NOT1 (N10876, N10870);
and AND3 (N10877, N10865, N1096, N7343);
nand NAND3 (N10878, N10877, N9257, N1079);
buf BUF1 (N10879, N10867);
buf BUF1 (N10880, N10873);
not NOT1 (N10881, N10875);
nor NOR3 (N10882, N10874, N7459, N9972);
and AND2 (N10883, N10859, N2508);
nor NOR3 (N10884, N10876, N6400, N4598);
nand NAND2 (N10885, N10882, N10852);
xor XOR2 (N10886, N10879, N463);
and AND3 (N10887, N10878, N5275, N3064);
nand NAND3 (N10888, N10861, N9145, N5816);
and AND2 (N10889, N10881, N1032);
and AND2 (N10890, N10887, N2484);
nor NOR2 (N10891, N10872, N2996);
not NOT1 (N10892, N10885);
nor NOR4 (N10893, N10888, N2017, N9656, N1777);
xor XOR2 (N10894, N10871, N9349);
and AND2 (N10895, N10893, N10696);
xor XOR2 (N10896, N10880, N7248);
or OR2 (N10897, N10886, N9331);
nor NOR2 (N10898, N10884, N5769);
and AND2 (N10899, N10894, N902);
buf BUF1 (N10900, N10899);
nand NAND2 (N10901, N10889, N8114);
nor NOR4 (N10902, N10900, N404, N6199, N9040);
nor NOR3 (N10903, N10897, N3759, N9182);
nand NAND3 (N10904, N10895, N10052, N2398);
nand NAND2 (N10905, N10892, N1129);
or OR4 (N10906, N10905, N1369, N7415, N5392);
nor NOR3 (N10907, N10898, N584, N1856);
or OR4 (N10908, N10891, N5889, N5645, N9121);
buf BUF1 (N10909, N10883);
xor XOR2 (N10910, N10903, N6273);
not NOT1 (N10911, N10906);
or OR2 (N10912, N10904, N6195);
buf BUF1 (N10913, N10912);
or OR4 (N10914, N10911, N9256, N3886, N10595);
not NOT1 (N10915, N10909);
or OR2 (N10916, N10907, N1980);
not NOT1 (N10917, N10908);
xor XOR2 (N10918, N10916, N6907);
nor NOR4 (N10919, N10917, N1288, N8129, N4500);
not NOT1 (N10920, N10914);
and AND2 (N10921, N10910, N3017);
nor NOR3 (N10922, N10890, N6417, N8942);
or OR4 (N10923, N10921, N10739, N2032, N138);
xor XOR2 (N10924, N10896, N3635);
buf BUF1 (N10925, N10919);
nand NAND2 (N10926, N10924, N4651);
buf BUF1 (N10927, N10918);
or OR2 (N10928, N10925, N5391);
buf BUF1 (N10929, N10926);
nor NOR3 (N10930, N10920, N1681, N8273);
nor NOR3 (N10931, N10901, N8402, N5110);
nor NOR3 (N10932, N10913, N4207, N3972);
or OR3 (N10933, N10902, N4946, N9101);
or OR2 (N10934, N10932, N5689);
not NOT1 (N10935, N10930);
nand NAND4 (N10936, N10923, N1699, N6485, N10630);
xor XOR2 (N10937, N10922, N1725);
nand NAND4 (N10938, N10936, N6411, N8744, N6866);
not NOT1 (N10939, N10929);
nand NAND4 (N10940, N10933, N7129, N6405, N6457);
buf BUF1 (N10941, N10935);
buf BUF1 (N10942, N10927);
nor NOR3 (N10943, N10931, N7617, N5319);
xor XOR2 (N10944, N10942, N7617);
and AND3 (N10945, N10944, N938, N3780);
buf BUF1 (N10946, N10941);
xor XOR2 (N10947, N10939, N9182);
and AND3 (N10948, N10943, N3938, N6557);
buf BUF1 (N10949, N10915);
buf BUF1 (N10950, N10940);
xor XOR2 (N10951, N10947, N2080);
nand NAND4 (N10952, N10928, N1893, N8138, N5188);
xor XOR2 (N10953, N10938, N8282);
nand NAND3 (N10954, N10937, N9588, N164);
and AND4 (N10955, N10945, N7645, N6414, N8445);
xor XOR2 (N10956, N10934, N5128);
not NOT1 (N10957, N10954);
not NOT1 (N10958, N10952);
nor NOR3 (N10959, N10958, N1268, N9443);
or OR4 (N10960, N10949, N5272, N7791, N10383);
buf BUF1 (N10961, N10959);
nor NOR3 (N10962, N10961, N7823, N3353);
xor XOR2 (N10963, N10953, N6821);
nor NOR3 (N10964, N10963, N6609, N2495);
or OR4 (N10965, N10957, N3995, N7836, N8891);
nand NAND2 (N10966, N10955, N4521);
buf BUF1 (N10967, N10950);
xor XOR2 (N10968, N10965, N8048);
not NOT1 (N10969, N10968);
nor NOR4 (N10970, N10948, N2977, N9214, N583);
buf BUF1 (N10971, N10946);
nand NAND2 (N10972, N10971, N2411);
nand NAND3 (N10973, N10962, N8106, N833);
nand NAND2 (N10974, N10966, N4121);
xor XOR2 (N10975, N10972, N162);
xor XOR2 (N10976, N10967, N5872);
or OR2 (N10977, N10960, N7345);
buf BUF1 (N10978, N10951);
not NOT1 (N10979, N10978);
buf BUF1 (N10980, N10973);
and AND3 (N10981, N10980, N10369, N7966);
xor XOR2 (N10982, N10969, N2255);
buf BUF1 (N10983, N10975);
or OR2 (N10984, N10974, N782);
and AND4 (N10985, N10956, N6968, N7621, N2660);
buf BUF1 (N10986, N10977);
or OR4 (N10987, N10985, N4798, N9976, N926);
nor NOR3 (N10988, N10987, N4634, N4378);
not NOT1 (N10989, N10984);
nand NAND3 (N10990, N10982, N5707, N9924);
buf BUF1 (N10991, N10976);
and AND2 (N10992, N10964, N10868);
buf BUF1 (N10993, N10979);
xor XOR2 (N10994, N10990, N8968);
and AND3 (N10995, N10991, N6151, N802);
not NOT1 (N10996, N10993);
or OR4 (N10997, N10994, N5737, N1605, N3604);
or OR3 (N10998, N10995, N3510, N9249);
nor NOR3 (N10999, N10996, N733, N9238);
nor NOR4 (N11000, N10992, N10755, N965, N6476);
buf BUF1 (N11001, N10989);
xor XOR2 (N11002, N10986, N5692);
not NOT1 (N11003, N10988);
and AND4 (N11004, N11000, N7143, N4179, N8621);
or OR4 (N11005, N11004, N9506, N4724, N5365);
nor NOR4 (N11006, N11003, N2398, N8660, N4887);
xor XOR2 (N11007, N10981, N7729);
or OR3 (N11008, N11005, N6179, N9798);
nand NAND4 (N11009, N11002, N4134, N1027, N5545);
or OR3 (N11010, N10998, N6133, N2753);
not NOT1 (N11011, N11010);
and AND3 (N11012, N11011, N10746, N4845);
not NOT1 (N11013, N11008);
or OR4 (N11014, N11013, N6432, N814, N6793);
and AND4 (N11015, N10983, N5530, N8134, N7541);
not NOT1 (N11016, N10999);
not NOT1 (N11017, N11007);
buf BUF1 (N11018, N11015);
xor XOR2 (N11019, N11016, N9008);
not NOT1 (N11020, N11006);
nand NAND4 (N11021, N11009, N8852, N8585, N7630);
buf BUF1 (N11022, N11012);
buf BUF1 (N11023, N11021);
xor XOR2 (N11024, N11017, N8920);
not NOT1 (N11025, N10997);
nand NAND2 (N11026, N11019, N6732);
not NOT1 (N11027, N11018);
buf BUF1 (N11028, N10970);
xor XOR2 (N11029, N11027, N1998);
nand NAND3 (N11030, N11024, N1199, N4213);
xor XOR2 (N11031, N11001, N3085);
xor XOR2 (N11032, N11029, N6600);
nand NAND3 (N11033, N11014, N5978, N8451);
not NOT1 (N11034, N11026);
xor XOR2 (N11035, N11030, N10034);
not NOT1 (N11036, N11033);
buf BUF1 (N11037, N11034);
buf BUF1 (N11038, N11023);
nor NOR3 (N11039, N11032, N8206, N4205);
nor NOR2 (N11040, N11020, N805);
or OR4 (N11041, N11040, N522, N1006, N3598);
xor XOR2 (N11042, N11035, N3313);
nand NAND2 (N11043, N11036, N3655);
or OR3 (N11044, N11031, N9767, N6380);
and AND3 (N11045, N11044, N7526, N5684);
buf BUF1 (N11046, N11045);
nand NAND3 (N11047, N11042, N6663, N6520);
nor NOR2 (N11048, N11028, N7984);
buf BUF1 (N11049, N11037);
nor NOR2 (N11050, N11039, N7519);
buf BUF1 (N11051, N11049);
and AND4 (N11052, N11025, N4827, N9798, N8123);
nand NAND2 (N11053, N11046, N8615);
nand NAND2 (N11054, N11038, N10580);
xor XOR2 (N11055, N11050, N801);
nand NAND2 (N11056, N11054, N4653);
nand NAND4 (N11057, N11051, N1167, N3513, N1088);
or OR2 (N11058, N11048, N10308);
buf BUF1 (N11059, N11047);
xor XOR2 (N11060, N11059, N8027);
nand NAND2 (N11061, N11053, N6534);
or OR2 (N11062, N11041, N944);
nor NOR2 (N11063, N11056, N3279);
or OR2 (N11064, N11060, N8957);
and AND3 (N11065, N11063, N3676, N3479);
nand NAND3 (N11066, N11064, N9068, N6476);
buf BUF1 (N11067, N11061);
nand NAND4 (N11068, N11066, N2691, N5245, N9348);
xor XOR2 (N11069, N11052, N8931);
buf BUF1 (N11070, N11043);
nor NOR3 (N11071, N11062, N1968, N3357);
nand NAND2 (N11072, N11068, N7814);
not NOT1 (N11073, N11065);
xor XOR2 (N11074, N11071, N11000);
or OR2 (N11075, N11067, N3964);
xor XOR2 (N11076, N11057, N1264);
not NOT1 (N11077, N11022);
or OR2 (N11078, N11069, N1831);
nand NAND3 (N11079, N11072, N9966, N2735);
buf BUF1 (N11080, N11074);
buf BUF1 (N11081, N11055);
not NOT1 (N11082, N11078);
buf BUF1 (N11083, N11082);
or OR2 (N11084, N11070, N9432);
not NOT1 (N11085, N11075);
nand NAND3 (N11086, N11073, N8610, N6193);
nor NOR2 (N11087, N11084, N3375);
xor XOR2 (N11088, N11076, N3178);
nand NAND4 (N11089, N11087, N9299, N6742, N2164);
buf BUF1 (N11090, N11089);
buf BUF1 (N11091, N11077);
and AND4 (N11092, N11083, N7124, N7251, N1286);
not NOT1 (N11093, N11085);
and AND2 (N11094, N11092, N5316);
not NOT1 (N11095, N11081);
xor XOR2 (N11096, N11094, N2969);
buf BUF1 (N11097, N11079);
or OR3 (N11098, N11097, N4387, N8330);
and AND2 (N11099, N11090, N9669);
not NOT1 (N11100, N11093);
nand NAND3 (N11101, N11095, N763, N3582);
and AND4 (N11102, N11098, N3970, N5919, N7581);
buf BUF1 (N11103, N11088);
or OR4 (N11104, N11080, N2762, N4559, N7561);
and AND3 (N11105, N11101, N9927, N5864);
buf BUF1 (N11106, N11086);
and AND4 (N11107, N11099, N5897, N6028, N10599);
nand NAND2 (N11108, N11103, N5351);
and AND3 (N11109, N11096, N10914, N6268);
nor NOR3 (N11110, N11102, N10417, N1104);
buf BUF1 (N11111, N11110);
xor XOR2 (N11112, N11108, N7738);
buf BUF1 (N11113, N11100);
nor NOR4 (N11114, N11107, N8888, N1784, N6795);
or OR4 (N11115, N11104, N6045, N685, N9670);
nor NOR2 (N11116, N11058, N9541);
nand NAND4 (N11117, N11105, N4988, N6050, N4486);
xor XOR2 (N11118, N11112, N10760);
nor NOR3 (N11119, N11113, N3726, N5263);
not NOT1 (N11120, N11109);
buf BUF1 (N11121, N11120);
nand NAND2 (N11122, N11116, N8487);
buf BUF1 (N11123, N11121);
nand NAND2 (N11124, N11115, N7262);
xor XOR2 (N11125, N11117, N2999);
nor NOR4 (N11126, N11125, N2665, N10983, N10268);
not NOT1 (N11127, N11118);
and AND3 (N11128, N11111, N6171, N8046);
buf BUF1 (N11129, N11123);
and AND3 (N11130, N11127, N9500, N4957);
xor XOR2 (N11131, N11130, N7029);
and AND2 (N11132, N11122, N4153);
buf BUF1 (N11133, N11132);
or OR2 (N11134, N11091, N842);
not NOT1 (N11135, N11133);
nand NAND4 (N11136, N11135, N3538, N1331, N9031);
or OR2 (N11137, N11136, N7518);
or OR4 (N11138, N11124, N3110, N7617, N5137);
or OR4 (N11139, N11126, N4709, N11006, N2814);
and AND3 (N11140, N11139, N2030, N10536);
nand NAND2 (N11141, N11131, N5244);
or OR2 (N11142, N11106, N3602);
or OR3 (N11143, N11142, N7166, N3927);
or OR4 (N11144, N11128, N7271, N6608, N4262);
xor XOR2 (N11145, N11129, N3987);
or OR3 (N11146, N11137, N2001, N801);
and AND3 (N11147, N11134, N695, N2248);
xor XOR2 (N11148, N11147, N11056);
buf BUF1 (N11149, N11145);
xor XOR2 (N11150, N11148, N3853);
buf BUF1 (N11151, N11144);
buf BUF1 (N11152, N11119);
and AND4 (N11153, N11141, N7934, N8257, N2028);
nand NAND2 (N11154, N11149, N3761);
or OR2 (N11155, N11138, N2948);
nand NAND4 (N11156, N11155, N6505, N116, N10072);
and AND3 (N11157, N11156, N2144, N5210);
nand NAND2 (N11158, N11151, N7097);
buf BUF1 (N11159, N11153);
and AND4 (N11160, N11158, N6960, N10361, N2761);
and AND3 (N11161, N11152, N4737, N7761);
nand NAND3 (N11162, N11161, N4587, N4413);
nand NAND3 (N11163, N11159, N10985, N2565);
xor XOR2 (N11164, N11162, N4706);
not NOT1 (N11165, N11163);
buf BUF1 (N11166, N11157);
nor NOR2 (N11167, N11146, N1207);
xor XOR2 (N11168, N11154, N7109);
nand NAND4 (N11169, N11114, N3740, N1841, N1912);
nor NOR4 (N11170, N11143, N1356, N10150, N2173);
nor NOR3 (N11171, N11167, N10293, N9174);
nand NAND3 (N11172, N11166, N9253, N10598);
nor NOR2 (N11173, N11172, N2072);
not NOT1 (N11174, N11165);
nor NOR3 (N11175, N11164, N1024, N1399);
nor NOR2 (N11176, N11173, N2672);
not NOT1 (N11177, N11169);
or OR4 (N11178, N11160, N9615, N3390, N3850);
nor NOR2 (N11179, N11178, N2425);
not NOT1 (N11180, N11177);
buf BUF1 (N11181, N11170);
nor NOR4 (N11182, N11181, N9327, N1496, N7756);
xor XOR2 (N11183, N11140, N10539);
nor NOR2 (N11184, N11179, N3279);
buf BUF1 (N11185, N11182);
and AND2 (N11186, N11174, N6482);
not NOT1 (N11187, N11186);
or OR2 (N11188, N11185, N5950);
nor NOR4 (N11189, N11187, N9050, N6491, N9936);
nor NOR4 (N11190, N11184, N11153, N10598, N8255);
or OR4 (N11191, N11190, N5061, N9583, N8709);
nor NOR2 (N11192, N11189, N10402);
xor XOR2 (N11193, N11192, N4081);
not NOT1 (N11194, N11193);
xor XOR2 (N11195, N11176, N2849);
buf BUF1 (N11196, N11195);
not NOT1 (N11197, N11168);
nand NAND2 (N11198, N11197, N1430);
xor XOR2 (N11199, N11150, N869);
xor XOR2 (N11200, N11183, N4086);
buf BUF1 (N11201, N11198);
xor XOR2 (N11202, N11175, N7826);
nor NOR3 (N11203, N11201, N4685, N3830);
nand NAND4 (N11204, N11196, N2536, N1064, N5177);
or OR3 (N11205, N11200, N832, N1285);
not NOT1 (N11206, N11171);
and AND4 (N11207, N11204, N3786, N5677, N1484);
nand NAND4 (N11208, N11202, N6503, N7901, N10279);
xor XOR2 (N11209, N11208, N7554);
nand NAND3 (N11210, N11180, N5931, N1139);
nor NOR4 (N11211, N11188, N4304, N192, N919);
or OR3 (N11212, N11211, N9317, N2430);
nor NOR2 (N11213, N11209, N10772);
buf BUF1 (N11214, N11213);
nor NOR4 (N11215, N11206, N9302, N3739, N6605);
and AND4 (N11216, N11214, N7356, N7720, N10897);
not NOT1 (N11217, N11216);
nor NOR2 (N11218, N11203, N9833);
buf BUF1 (N11219, N11191);
nor NOR4 (N11220, N11205, N7623, N3604, N6069);
nor NOR3 (N11221, N11220, N6872, N1994);
or OR3 (N11222, N11217, N600, N5683);
and AND4 (N11223, N11212, N6594, N3147, N8098);
not NOT1 (N11224, N11219);
nor NOR2 (N11225, N11215, N6693);
or OR2 (N11226, N11224, N3003);
buf BUF1 (N11227, N11225);
nor NOR2 (N11228, N11218, N5044);
not NOT1 (N11229, N11227);
not NOT1 (N11230, N11199);
nor NOR4 (N11231, N11221, N5111, N8709, N8569);
xor XOR2 (N11232, N11228, N8270);
or OR2 (N11233, N11232, N8440);
buf BUF1 (N11234, N11230);
xor XOR2 (N11235, N11223, N1989);
not NOT1 (N11236, N11222);
nand NAND4 (N11237, N11194, N8153, N8394, N1156);
buf BUF1 (N11238, N11210);
and AND4 (N11239, N11238, N10292, N4988, N8392);
buf BUF1 (N11240, N11234);
buf BUF1 (N11241, N11231);
xor XOR2 (N11242, N11235, N9057);
nor NOR2 (N11243, N11226, N7703);
and AND3 (N11244, N11240, N1773, N4992);
nand NAND2 (N11245, N11244, N6398);
and AND4 (N11246, N11243, N2936, N8783, N2854);
xor XOR2 (N11247, N11239, N10870);
and AND3 (N11248, N11207, N4797, N5075);
nand NAND4 (N11249, N11241, N1515, N3505, N3805);
or OR4 (N11250, N11247, N9584, N6430, N8412);
or OR3 (N11251, N11236, N7702, N10938);
or OR2 (N11252, N11237, N684);
and AND3 (N11253, N11249, N6138, N6158);
nand NAND4 (N11254, N11252, N5892, N6071, N5833);
and AND2 (N11255, N11251, N3699);
nor NOR2 (N11256, N11233, N6725);
nor NOR2 (N11257, N11246, N3);
nand NAND4 (N11258, N11229, N6329, N6683, N10789);
or OR2 (N11259, N11245, N3952);
xor XOR2 (N11260, N11253, N11119);
and AND3 (N11261, N11259, N10996, N481);
nor NOR4 (N11262, N11257, N6556, N6945, N3006);
nand NAND3 (N11263, N11260, N3493, N1294);
and AND2 (N11264, N11250, N6467);
xor XOR2 (N11265, N11258, N9100);
and AND4 (N11266, N11263, N2314, N485, N5165);
nand NAND2 (N11267, N11242, N7110);
or OR4 (N11268, N11266, N10194, N1335, N937);
not NOT1 (N11269, N11264);
and AND3 (N11270, N11268, N8136, N2826);
nand NAND3 (N11271, N11254, N3044, N3300);
not NOT1 (N11272, N11261);
and AND2 (N11273, N11271, N2548);
xor XOR2 (N11274, N11248, N8846);
nor NOR3 (N11275, N11255, N6542, N4893);
or OR4 (N11276, N11262, N1153, N10722, N4660);
nand NAND2 (N11277, N11276, N5264);
or OR4 (N11278, N11256, N5425, N4348, N7205);
or OR3 (N11279, N11272, N7299, N2356);
nand NAND2 (N11280, N11278, N10194);
or OR3 (N11281, N11279, N854, N1334);
xor XOR2 (N11282, N11277, N2393);
nor NOR2 (N11283, N11282, N1975);
not NOT1 (N11284, N11283);
or OR2 (N11285, N11267, N2040);
nor NOR4 (N11286, N11275, N2947, N9485, N3394);
not NOT1 (N11287, N11274);
or OR2 (N11288, N11265, N1594);
and AND3 (N11289, N11280, N1262, N4590);
xor XOR2 (N11290, N11285, N4797);
xor XOR2 (N11291, N11286, N7525);
nand NAND2 (N11292, N11289, N2180);
xor XOR2 (N11293, N11273, N10320);
buf BUF1 (N11294, N11290);
and AND4 (N11295, N11270, N3010, N9818, N1170);
or OR3 (N11296, N11294, N10913, N1736);
xor XOR2 (N11297, N11269, N8726);
nor NOR4 (N11298, N11287, N7705, N1665, N7233);
not NOT1 (N11299, N11288);
buf BUF1 (N11300, N11299);
and AND4 (N11301, N11296, N2493, N661, N50);
and AND2 (N11302, N11281, N7023);
nand NAND3 (N11303, N11295, N2010, N11091);
nand NAND2 (N11304, N11303, N3145);
nand NAND4 (N11305, N11304, N2683, N2823, N192);
buf BUF1 (N11306, N11301);
not NOT1 (N11307, N11302);
buf BUF1 (N11308, N11306);
and AND2 (N11309, N11308, N11173);
or OR4 (N11310, N11284, N4267, N10265, N1073);
xor XOR2 (N11311, N11293, N1132);
nor NOR2 (N11312, N11309, N7546);
not NOT1 (N11313, N11297);
and AND2 (N11314, N11307, N4833);
xor XOR2 (N11315, N11305, N3448);
buf BUF1 (N11316, N11292);
nor NOR3 (N11317, N11312, N6072, N4777);
buf BUF1 (N11318, N11317);
nand NAND4 (N11319, N11300, N7394, N10113, N6922);
or OR3 (N11320, N11311, N7802, N7230);
xor XOR2 (N11321, N11314, N9979);
nor NOR3 (N11322, N11313, N4607, N9995);
nand NAND2 (N11323, N11298, N9664);
and AND2 (N11324, N11320, N2497);
nand NAND3 (N11325, N11291, N3141, N5429);
nand NAND4 (N11326, N11321, N665, N9533, N4519);
nand NAND2 (N11327, N11323, N4029);
or OR2 (N11328, N11322, N1521);
xor XOR2 (N11329, N11327, N10931);
xor XOR2 (N11330, N11319, N7476);
nor NOR2 (N11331, N11330, N6772);
buf BUF1 (N11332, N11331);
or OR3 (N11333, N11329, N322, N1152);
buf BUF1 (N11334, N11315);
nor NOR4 (N11335, N11324, N4884, N980, N1486);
nand NAND3 (N11336, N11318, N4697, N1643);
and AND2 (N11337, N11334, N1098);
and AND3 (N11338, N11326, N7935, N287);
nand NAND2 (N11339, N11338, N2175);
xor XOR2 (N11340, N11328, N2270);
or OR3 (N11341, N11333, N950, N6208);
and AND2 (N11342, N11310, N7269);
buf BUF1 (N11343, N11340);
and AND4 (N11344, N11336, N8044, N8851, N2389);
or OR2 (N11345, N11316, N9136);
and AND4 (N11346, N11339, N1905, N175, N1769);
nor NOR4 (N11347, N11332, N5179, N3914, N4319);
buf BUF1 (N11348, N11343);
and AND2 (N11349, N11347, N9902);
buf BUF1 (N11350, N11341);
nor NOR3 (N11351, N11346, N9548, N6011);
and AND3 (N11352, N11349, N1249, N10563);
and AND4 (N11353, N11345, N2286, N4967, N10683);
not NOT1 (N11354, N11325);
or OR2 (N11355, N11348, N2154);
nand NAND4 (N11356, N11337, N7768, N6574, N7826);
nand NAND3 (N11357, N11356, N9298, N495);
nor NOR2 (N11358, N11352, N1285);
or OR3 (N11359, N11344, N2377, N825);
and AND4 (N11360, N11351, N4979, N5620, N9187);
xor XOR2 (N11361, N11354, N3697);
nand NAND3 (N11362, N11353, N4476, N5531);
and AND3 (N11363, N11362, N7540, N1679);
nor NOR3 (N11364, N11361, N10030, N6693);
buf BUF1 (N11365, N11355);
nor NOR2 (N11366, N11364, N8920);
nor NOR2 (N11367, N11350, N2375);
xor XOR2 (N11368, N11357, N4978);
nor NOR2 (N11369, N11342, N7708);
or OR3 (N11370, N11359, N2395, N6727);
nor NOR4 (N11371, N11366, N4833, N1864, N4507);
not NOT1 (N11372, N11360);
and AND3 (N11373, N11369, N114, N4885);
and AND2 (N11374, N11358, N11373);
buf BUF1 (N11375, N10999);
nor NOR3 (N11376, N11375, N10837, N8177);
xor XOR2 (N11377, N11372, N8465);
or OR4 (N11378, N11371, N7444, N11201, N9018);
nor NOR2 (N11379, N11368, N1830);
nand NAND3 (N11380, N11374, N8497, N7458);
buf BUF1 (N11381, N11377);
and AND4 (N11382, N11379, N4309, N9311, N6857);
xor XOR2 (N11383, N11370, N8367);
nand NAND2 (N11384, N11381, N5633);
nor NOR2 (N11385, N11382, N7374);
nor NOR2 (N11386, N11383, N1097);
not NOT1 (N11387, N11376);
xor XOR2 (N11388, N11365, N2765);
not NOT1 (N11389, N11378);
or OR3 (N11390, N11386, N1807, N8379);
nor NOR2 (N11391, N11389, N5435);
and AND2 (N11392, N11388, N6802);
buf BUF1 (N11393, N11363);
or OR2 (N11394, N11367, N11191);
nand NAND2 (N11395, N11392, N696);
xor XOR2 (N11396, N11387, N190);
or OR2 (N11397, N11385, N11325);
xor XOR2 (N11398, N11380, N8616);
nand NAND2 (N11399, N11391, N2067);
nor NOR2 (N11400, N11335, N4384);
buf BUF1 (N11401, N11398);
nand NAND3 (N11402, N11399, N10885, N3826);
nor NOR2 (N11403, N11400, N5199);
or OR2 (N11404, N11395, N6088);
nor NOR3 (N11405, N11403, N6202, N4179);
buf BUF1 (N11406, N11396);
and AND4 (N11407, N11402, N8871, N2239, N4413);
or OR2 (N11408, N11406, N1453);
xor XOR2 (N11409, N11384, N8960);
nand NAND2 (N11410, N11405, N2689);
buf BUF1 (N11411, N11408);
nand NAND3 (N11412, N11410, N159, N6432);
nand NAND2 (N11413, N11393, N2769);
nor NOR4 (N11414, N11404, N112, N2493, N8398);
buf BUF1 (N11415, N11397);
or OR2 (N11416, N11414, N9116);
not NOT1 (N11417, N11394);
not NOT1 (N11418, N11407);
nand NAND3 (N11419, N11413, N2940, N10651);
not NOT1 (N11420, N11411);
xor XOR2 (N11421, N11416, N8146);
nor NOR4 (N11422, N11420, N6900, N7565, N7609);
or OR2 (N11423, N11412, N7630);
not NOT1 (N11424, N11422);
or OR2 (N11425, N11418, N7465);
xor XOR2 (N11426, N11415, N9258);
or OR3 (N11427, N11419, N230, N875);
not NOT1 (N11428, N11421);
or OR2 (N11429, N11409, N7128);
buf BUF1 (N11430, N11390);
nor NOR4 (N11431, N11417, N4048, N6064, N7738);
buf BUF1 (N11432, N11430);
not NOT1 (N11433, N11424);
buf BUF1 (N11434, N11426);
and AND2 (N11435, N11401, N555);
buf BUF1 (N11436, N11435);
buf BUF1 (N11437, N11434);
xor XOR2 (N11438, N11431, N3535);
xor XOR2 (N11439, N11437, N1994);
and AND2 (N11440, N11429, N9170);
not NOT1 (N11441, N11428);
not NOT1 (N11442, N11425);
not NOT1 (N11443, N11433);
xor XOR2 (N11444, N11443, N3942);
xor XOR2 (N11445, N11439, N4105);
nor NOR2 (N11446, N11427, N6428);
or OR3 (N11447, N11446, N10100, N6387);
nand NAND2 (N11448, N11444, N5982);
nor NOR2 (N11449, N11438, N210);
or OR2 (N11450, N11436, N6929);
xor XOR2 (N11451, N11432, N1510);
or OR4 (N11452, N11448, N9755, N7193, N1726);
nor NOR3 (N11453, N11451, N1871, N1956);
and AND2 (N11454, N11449, N2757);
xor XOR2 (N11455, N11442, N9401);
or OR2 (N11456, N11450, N1458);
and AND2 (N11457, N11453, N2343);
and AND3 (N11458, N11454, N11164, N7065);
xor XOR2 (N11459, N11456, N5284);
nor NOR3 (N11460, N11459, N10370, N5542);
not NOT1 (N11461, N11458);
nand NAND3 (N11462, N11452, N3171, N7480);
nand NAND4 (N11463, N11461, N4919, N2095, N4546);
and AND4 (N11464, N11423, N11183, N3544, N7453);
nand NAND2 (N11465, N11445, N1836);
and AND2 (N11466, N11440, N8554);
xor XOR2 (N11467, N11455, N3656);
or OR3 (N11468, N11462, N5667, N10238);
xor XOR2 (N11469, N11464, N1315);
nand NAND2 (N11470, N11457, N5305);
xor XOR2 (N11471, N11470, N7472);
or OR2 (N11472, N11467, N7931);
not NOT1 (N11473, N11447);
nor NOR2 (N11474, N11463, N1779);
xor XOR2 (N11475, N11468, N9819);
xor XOR2 (N11476, N11441, N1894);
buf BUF1 (N11477, N11465);
or OR2 (N11478, N11466, N5940);
not NOT1 (N11479, N11476);
xor XOR2 (N11480, N11460, N8686);
xor XOR2 (N11481, N11475, N4959);
buf BUF1 (N11482, N11474);
nor NOR3 (N11483, N11478, N805, N8829);
buf BUF1 (N11484, N11483);
nor NOR2 (N11485, N11477, N4640);
buf BUF1 (N11486, N11471);
and AND4 (N11487, N11481, N6747, N212, N3521);
and AND2 (N11488, N11472, N181);
xor XOR2 (N11489, N11485, N10674);
and AND4 (N11490, N11489, N6851, N6721, N9468);
not NOT1 (N11491, N11490);
buf BUF1 (N11492, N11482);
or OR2 (N11493, N11479, N1975);
buf BUF1 (N11494, N11469);
xor XOR2 (N11495, N11494, N6429);
nand NAND2 (N11496, N11484, N5322);
or OR3 (N11497, N11473, N996, N7068);
or OR4 (N11498, N11486, N1196, N990, N3999);
nor NOR3 (N11499, N11487, N10168, N8355);
nor NOR4 (N11500, N11488, N2785, N1201, N3139);
buf BUF1 (N11501, N11497);
or OR4 (N11502, N11500, N4715, N8745, N7973);
and AND3 (N11503, N11480, N7434, N8543);
not NOT1 (N11504, N11493);
or OR2 (N11505, N11501, N1969);
nand NAND2 (N11506, N11492, N5032);
or OR2 (N11507, N11499, N7940);
not NOT1 (N11508, N11498);
xor XOR2 (N11509, N11502, N7103);
or OR3 (N11510, N11506, N9696, N2074);
nor NOR2 (N11511, N11510, N3619);
xor XOR2 (N11512, N11508, N6935);
nand NAND2 (N11513, N11496, N1511);
not NOT1 (N11514, N11491);
xor XOR2 (N11515, N11507, N4274);
buf BUF1 (N11516, N11515);
and AND4 (N11517, N11505, N7135, N2131, N8914);
and AND3 (N11518, N11503, N8580, N2250);
buf BUF1 (N11519, N11511);
buf BUF1 (N11520, N11514);
nor NOR2 (N11521, N11504, N4386);
nor NOR4 (N11522, N11513, N6341, N8752, N814);
or OR3 (N11523, N11512, N8989, N7460);
xor XOR2 (N11524, N11509, N10392);
and AND3 (N11525, N11524, N7103, N1571);
xor XOR2 (N11526, N11521, N2331);
buf BUF1 (N11527, N11495);
xor XOR2 (N11528, N11520, N2715);
or OR3 (N11529, N11527, N5722, N2574);
not NOT1 (N11530, N11528);
nor NOR2 (N11531, N11525, N4536);
buf BUF1 (N11532, N11529);
and AND4 (N11533, N11518, N548, N10893, N2672);
nor NOR4 (N11534, N11519, N3594, N11139, N10348);
buf BUF1 (N11535, N11522);
buf BUF1 (N11536, N11535);
and AND2 (N11537, N11526, N3934);
or OR2 (N11538, N11532, N4744);
or OR4 (N11539, N11530, N1581, N11288, N7306);
not NOT1 (N11540, N11537);
nand NAND4 (N11541, N11533, N10882, N5870, N8748);
and AND4 (N11542, N11517, N5754, N5362, N7424);
xor XOR2 (N11543, N11536, N8773);
buf BUF1 (N11544, N11541);
not NOT1 (N11545, N11539);
buf BUF1 (N11546, N11531);
buf BUF1 (N11547, N11516);
nor NOR3 (N11548, N11542, N2847, N9417);
not NOT1 (N11549, N11543);
xor XOR2 (N11550, N11540, N4426);
buf BUF1 (N11551, N11523);
xor XOR2 (N11552, N11546, N7989);
nor NOR3 (N11553, N11548, N3648, N4118);
and AND4 (N11554, N11544, N515, N3367, N117);
and AND2 (N11555, N11545, N7216);
and AND2 (N11556, N11552, N5059);
not NOT1 (N11557, N11555);
not NOT1 (N11558, N11538);
or OR2 (N11559, N11549, N5829);
not NOT1 (N11560, N11558);
not NOT1 (N11561, N11547);
xor XOR2 (N11562, N11559, N4541);
not NOT1 (N11563, N11553);
nand NAND2 (N11564, N11560, N476);
and AND4 (N11565, N11562, N1635, N109, N194);
and AND2 (N11566, N11551, N2656);
not NOT1 (N11567, N11561);
buf BUF1 (N11568, N11554);
not NOT1 (N11569, N11566);
buf BUF1 (N11570, N11564);
nor NOR2 (N11571, N11570, N9593);
buf BUF1 (N11572, N11534);
xor XOR2 (N11573, N11563, N10723);
not NOT1 (N11574, N11572);
nor NOR4 (N11575, N11550, N10346, N665, N2172);
buf BUF1 (N11576, N11565);
nor NOR2 (N11577, N11574, N2759);
buf BUF1 (N11578, N11568);
nor NOR4 (N11579, N11569, N8099, N7660, N3234);
xor XOR2 (N11580, N11573, N4786);
or OR4 (N11581, N11567, N5065, N1221, N3720);
xor XOR2 (N11582, N11581, N7744);
or OR3 (N11583, N11580, N4769, N5121);
or OR3 (N11584, N11576, N9634, N5434);
buf BUF1 (N11585, N11577);
and AND4 (N11586, N11583, N4723, N2657, N8062);
nand NAND2 (N11587, N11575, N6867);
and AND3 (N11588, N11556, N9544, N10536);
xor XOR2 (N11589, N11579, N4706);
nand NAND4 (N11590, N11588, N10953, N4787, N5330);
buf BUF1 (N11591, N11557);
not NOT1 (N11592, N11586);
buf BUF1 (N11593, N11578);
nand NAND3 (N11594, N11589, N11494, N5453);
or OR3 (N11595, N11585, N3605, N6579);
or OR2 (N11596, N11571, N2997);
nor NOR2 (N11597, N11596, N11335);
or OR3 (N11598, N11595, N4593, N2035);
nor NOR3 (N11599, N11597, N2565, N2816);
or OR4 (N11600, N11587, N9159, N4111, N651);
buf BUF1 (N11601, N11582);
not NOT1 (N11602, N11594);
or OR3 (N11603, N11584, N8562, N3667);
nand NAND4 (N11604, N11591, N7359, N2169, N3621);
nor NOR2 (N11605, N11604, N10964);
nor NOR3 (N11606, N11592, N8659, N6980);
or OR3 (N11607, N11606, N11228, N1258);
nor NOR2 (N11608, N11603, N9525);
nor NOR2 (N11609, N11602, N5165);
nand NAND4 (N11610, N11598, N10350, N9595, N4516);
and AND3 (N11611, N11599, N6802, N10312);
buf BUF1 (N11612, N11601);
or OR3 (N11613, N11607, N9078, N4322);
nand NAND2 (N11614, N11593, N6496);
not NOT1 (N11615, N11590);
buf BUF1 (N11616, N11600);
not NOT1 (N11617, N11608);
xor XOR2 (N11618, N11611, N6444);
buf BUF1 (N11619, N11617);
not NOT1 (N11620, N11619);
and AND3 (N11621, N11616, N1215, N10579);
nand NAND4 (N11622, N11605, N10352, N1180, N5285);
nor NOR4 (N11623, N11610, N1374, N5292, N1530);
or OR2 (N11624, N11612, N3021);
not NOT1 (N11625, N11615);
nand NAND4 (N11626, N11622, N8454, N8004, N7454);
nand NAND2 (N11627, N11613, N189);
and AND2 (N11628, N11623, N4444);
or OR4 (N11629, N11626, N1501, N5594, N6221);
nor NOR3 (N11630, N11624, N8115, N6361);
buf BUF1 (N11631, N11620);
buf BUF1 (N11632, N11629);
nor NOR2 (N11633, N11628, N10099);
not NOT1 (N11634, N11625);
and AND2 (N11635, N11609, N10318);
not NOT1 (N11636, N11633);
or OR3 (N11637, N11635, N4537, N746);
and AND3 (N11638, N11632, N9968, N2598);
nand NAND3 (N11639, N11637, N4330, N9586);
nand NAND2 (N11640, N11634, N7844);
xor XOR2 (N11641, N11631, N8776);
not NOT1 (N11642, N11640);
xor XOR2 (N11643, N11614, N7497);
not NOT1 (N11644, N11636);
and AND3 (N11645, N11639, N3288, N8278);
and AND3 (N11646, N11618, N270, N8207);
buf BUF1 (N11647, N11630);
and AND3 (N11648, N11642, N3470, N8862);
or OR3 (N11649, N11627, N11220, N8732);
nor NOR3 (N11650, N11646, N7038, N11073);
xor XOR2 (N11651, N11643, N9151);
and AND2 (N11652, N11641, N7729);
buf BUF1 (N11653, N11651);
not NOT1 (N11654, N11644);
and AND2 (N11655, N11621, N585);
xor XOR2 (N11656, N11649, N2159);
or OR4 (N11657, N11647, N395, N7045, N6006);
buf BUF1 (N11658, N11650);
buf BUF1 (N11659, N11653);
not NOT1 (N11660, N11645);
nor NOR4 (N11661, N11648, N10002, N10849, N1292);
nor NOR3 (N11662, N11658, N6296, N7520);
xor XOR2 (N11663, N11661, N6229);
or OR3 (N11664, N11638, N8025, N6180);
xor XOR2 (N11665, N11655, N10657);
and AND2 (N11666, N11657, N4530);
buf BUF1 (N11667, N11664);
or OR2 (N11668, N11662, N11290);
buf BUF1 (N11669, N11659);
not NOT1 (N11670, N11652);
xor XOR2 (N11671, N11665, N2571);
xor XOR2 (N11672, N11670, N913);
not NOT1 (N11673, N11667);
and AND4 (N11674, N11654, N111, N11639, N7684);
or OR3 (N11675, N11656, N1497, N7108);
xor XOR2 (N11676, N11666, N10061);
buf BUF1 (N11677, N11671);
or OR2 (N11678, N11660, N634);
not NOT1 (N11679, N11677);
nor NOR3 (N11680, N11668, N8156, N5540);
not NOT1 (N11681, N11675);
not NOT1 (N11682, N11674);
xor XOR2 (N11683, N11672, N11165);
and AND3 (N11684, N11673, N1685, N5938);
not NOT1 (N11685, N11680);
or OR4 (N11686, N11679, N3918, N6079, N7716);
nand NAND2 (N11687, N11682, N752);
not NOT1 (N11688, N11685);
or OR4 (N11689, N11684, N257, N11082, N6935);
and AND2 (N11690, N11689, N8682);
not NOT1 (N11691, N11681);
nand NAND4 (N11692, N11686, N2468, N9357, N731);
nor NOR2 (N11693, N11678, N3874);
xor XOR2 (N11694, N11688, N4799);
xor XOR2 (N11695, N11676, N7379);
nand NAND3 (N11696, N11669, N1443, N8727);
nand NAND3 (N11697, N11694, N8674, N953);
nand NAND2 (N11698, N11692, N7350);
buf BUF1 (N11699, N11697);
or OR4 (N11700, N11696, N2380, N2021, N4165);
nand NAND3 (N11701, N11683, N4223, N7848);
nand NAND2 (N11702, N11691, N11332);
and AND4 (N11703, N11695, N7149, N9222, N11667);
nand NAND4 (N11704, N11690, N8888, N212, N7398);
buf BUF1 (N11705, N11693);
and AND3 (N11706, N11702, N1008, N7654);
buf BUF1 (N11707, N11705);
nor NOR2 (N11708, N11663, N8995);
not NOT1 (N11709, N11699);
buf BUF1 (N11710, N11708);
nor NOR3 (N11711, N11707, N8534, N9906);
and AND4 (N11712, N11700, N9014, N10613, N3626);
or OR4 (N11713, N11712, N10829, N10143, N7121);
not NOT1 (N11714, N11709);
nor NOR3 (N11715, N11713, N6810, N11098);
buf BUF1 (N11716, N11715);
nand NAND4 (N11717, N11703, N4210, N11510, N6975);
nand NAND4 (N11718, N11687, N7998, N7464, N10201);
xor XOR2 (N11719, N11706, N839);
buf BUF1 (N11720, N11716);
xor XOR2 (N11721, N11701, N7284);
and AND4 (N11722, N11714, N3198, N9391, N1252);
buf BUF1 (N11723, N11717);
xor XOR2 (N11724, N11698, N4293);
nor NOR3 (N11725, N11720, N7436, N3093);
xor XOR2 (N11726, N11711, N11025);
not NOT1 (N11727, N11704);
or OR4 (N11728, N11710, N6046, N3964, N10087);
xor XOR2 (N11729, N11724, N4224);
or OR2 (N11730, N11725, N6659);
not NOT1 (N11731, N11728);
buf BUF1 (N11732, N11719);
xor XOR2 (N11733, N11718, N4152);
buf BUF1 (N11734, N11731);
xor XOR2 (N11735, N11733, N11195);
xor XOR2 (N11736, N11726, N10444);
and AND3 (N11737, N11721, N9477, N6772);
xor XOR2 (N11738, N11722, N539);
nor NOR2 (N11739, N11736, N4798);
or OR2 (N11740, N11732, N7263);
nor NOR3 (N11741, N11735, N2520, N7005);
xor XOR2 (N11742, N11729, N2057);
nor NOR3 (N11743, N11727, N4527, N7910);
and AND2 (N11744, N11740, N392);
not NOT1 (N11745, N11723);
not NOT1 (N11746, N11737);
or OR2 (N11747, N11734, N9917);
not NOT1 (N11748, N11743);
nand NAND3 (N11749, N11746, N2457, N4453);
nor NOR2 (N11750, N11748, N3065);
nor NOR3 (N11751, N11730, N7571, N2910);
xor XOR2 (N11752, N11751, N6505);
xor XOR2 (N11753, N11741, N4087);
or OR2 (N11754, N11747, N11366);
not NOT1 (N11755, N11752);
buf BUF1 (N11756, N11742);
nor NOR2 (N11757, N11739, N5955);
or OR4 (N11758, N11754, N3043, N10165, N1224);
nor NOR2 (N11759, N11738, N4928);
not NOT1 (N11760, N11753);
or OR3 (N11761, N11750, N3264, N4701);
xor XOR2 (N11762, N11755, N1017);
not NOT1 (N11763, N11759);
xor XOR2 (N11764, N11758, N1824);
or OR2 (N11765, N11760, N2854);
nor NOR4 (N11766, N11756, N2617, N4076, N10168);
and AND3 (N11767, N11745, N10229, N10641);
nand NAND2 (N11768, N11766, N8475);
nor NOR3 (N11769, N11749, N4788, N10770);
buf BUF1 (N11770, N11763);
xor XOR2 (N11771, N11762, N11383);
nor NOR3 (N11772, N11769, N6004, N7350);
xor XOR2 (N11773, N11771, N5970);
buf BUF1 (N11774, N11767);
buf BUF1 (N11775, N11744);
nand NAND2 (N11776, N11773, N8940);
nand NAND2 (N11777, N11770, N4578);
and AND4 (N11778, N11777, N6601, N11018, N5094);
nand NAND4 (N11779, N11768, N9870, N1037, N11274);
xor XOR2 (N11780, N11764, N9322);
not NOT1 (N11781, N11765);
not NOT1 (N11782, N11775);
xor XOR2 (N11783, N11778, N466);
buf BUF1 (N11784, N11776);
not NOT1 (N11785, N11782);
and AND3 (N11786, N11785, N11759, N11395);
or OR3 (N11787, N11772, N8356, N11388);
nor NOR3 (N11788, N11774, N10474, N9573);
and AND4 (N11789, N11787, N7397, N1198, N707);
buf BUF1 (N11790, N11779);
nand NAND2 (N11791, N11788, N1196);
nand NAND2 (N11792, N11780, N4835);
and AND4 (N11793, N11757, N1926, N10059, N10327);
and AND4 (N11794, N11792, N4825, N10669, N9957);
or OR3 (N11795, N11794, N9739, N2602);
and AND2 (N11796, N11795, N11050);
or OR3 (N11797, N11786, N1419, N1827);
or OR3 (N11798, N11761, N7276, N6586);
nor NOR3 (N11799, N11798, N5515, N1293);
buf BUF1 (N11800, N11796);
nand NAND3 (N11801, N11790, N8689, N8634);
not NOT1 (N11802, N11800);
or OR3 (N11803, N11802, N6751, N9079);
not NOT1 (N11804, N11783);
or OR2 (N11805, N11781, N3751);
nor NOR4 (N11806, N11793, N8693, N6735, N7531);
not NOT1 (N11807, N11805);
and AND3 (N11808, N11806, N6190, N11628);
nand NAND2 (N11809, N11801, N11330);
nor NOR3 (N11810, N11804, N20, N1500);
buf BUF1 (N11811, N11799);
or OR2 (N11812, N11789, N4162);
nor NOR4 (N11813, N11803, N10688, N4140, N5034);
not NOT1 (N11814, N11812);
nand NAND3 (N11815, N11797, N832, N395);
buf BUF1 (N11816, N11814);
nand NAND3 (N11817, N11815, N9565, N11344);
not NOT1 (N11818, N11813);
buf BUF1 (N11819, N11808);
not NOT1 (N11820, N11784);
nand NAND2 (N11821, N11810, N4471);
buf BUF1 (N11822, N11811);
xor XOR2 (N11823, N11821, N2156);
buf BUF1 (N11824, N11822);
and AND2 (N11825, N11809, N932);
nand NAND4 (N11826, N11817, N3066, N5292, N3326);
nand NAND3 (N11827, N11823, N884, N10237);
nand NAND2 (N11828, N11825, N455);
or OR2 (N11829, N11824, N8240);
nor NOR3 (N11830, N11829, N9058, N4800);
nand NAND2 (N11831, N11816, N7279);
and AND4 (N11832, N11791, N5181, N6294, N7366);
nand NAND4 (N11833, N11831, N8872, N16, N11646);
nor NOR4 (N11834, N11827, N5387, N10639, N3482);
nor NOR2 (N11835, N11807, N11117);
not NOT1 (N11836, N11835);
not NOT1 (N11837, N11818);
or OR2 (N11838, N11837, N9582);
nor NOR3 (N11839, N11826, N7412, N4009);
not NOT1 (N11840, N11838);
and AND2 (N11841, N11834, N3867);
and AND3 (N11842, N11832, N2320, N2280);
xor XOR2 (N11843, N11841, N3515);
or OR3 (N11844, N11820, N6495, N5117);
or OR4 (N11845, N11833, N5377, N10494, N4215);
or OR2 (N11846, N11844, N10066);
nand NAND2 (N11847, N11846, N10899);
xor XOR2 (N11848, N11845, N8393);
not NOT1 (N11849, N11830);
nand NAND4 (N11850, N11848, N6919, N2674, N6133);
nor NOR2 (N11851, N11849, N4187);
buf BUF1 (N11852, N11840);
nor NOR3 (N11853, N11850, N4650, N4187);
nand NAND3 (N11854, N11852, N8353, N11334);
not NOT1 (N11855, N11842);
nand NAND4 (N11856, N11851, N9057, N8382, N2204);
buf BUF1 (N11857, N11839);
or OR3 (N11858, N11819, N5515, N6600);
and AND2 (N11859, N11856, N7022);
buf BUF1 (N11860, N11855);
nand NAND4 (N11861, N11847, N8009, N6418, N2855);
nand NAND2 (N11862, N11854, N3469);
xor XOR2 (N11863, N11861, N6685);
buf BUF1 (N11864, N11858);
buf BUF1 (N11865, N11863);
not NOT1 (N11866, N11828);
buf BUF1 (N11867, N11860);
nand NAND4 (N11868, N11853, N10717, N2122, N3073);
nand NAND3 (N11869, N11859, N59, N10201);
xor XOR2 (N11870, N11836, N606);
nor NOR2 (N11871, N11862, N295);
xor XOR2 (N11872, N11857, N10143);
not NOT1 (N11873, N11866);
nand NAND3 (N11874, N11869, N10363, N11460);
nor NOR3 (N11875, N11843, N10890, N2937);
buf BUF1 (N11876, N11872);
and AND4 (N11877, N11867, N3192, N11642, N295);
and AND3 (N11878, N11870, N4849, N3842);
xor XOR2 (N11879, N11873, N9194);
nand NAND2 (N11880, N11871, N8592);
or OR3 (N11881, N11876, N3600, N8157);
xor XOR2 (N11882, N11864, N967);
and AND2 (N11883, N11879, N4736);
nor NOR4 (N11884, N11880, N303, N8219, N10544);
xor XOR2 (N11885, N11874, N3470);
nand NAND3 (N11886, N11884, N2479, N11863);
or OR4 (N11887, N11881, N344, N3320, N3833);
not NOT1 (N11888, N11877);
not NOT1 (N11889, N11868);
and AND4 (N11890, N11883, N5439, N4540, N277);
not NOT1 (N11891, N11890);
buf BUF1 (N11892, N11878);
and AND2 (N11893, N11885, N4605);
or OR2 (N11894, N11889, N4935);
buf BUF1 (N11895, N11891);
or OR2 (N11896, N11892, N1067);
xor XOR2 (N11897, N11888, N6533);
not NOT1 (N11898, N11882);
not NOT1 (N11899, N11865);
nand NAND4 (N11900, N11894, N84, N400, N7937);
nand NAND4 (N11901, N11875, N3059, N4328, N10921);
not NOT1 (N11902, N11899);
nor NOR2 (N11903, N11886, N7642);
nor NOR4 (N11904, N11900, N6589, N743, N11446);
and AND2 (N11905, N11897, N9385);
xor XOR2 (N11906, N11902, N2266);
nor NOR4 (N11907, N11893, N6113, N9029, N4372);
nor NOR3 (N11908, N11896, N5626, N10713);
nand NAND4 (N11909, N11901, N8783, N5511, N2049);
or OR4 (N11910, N11906, N10515, N6017, N9937);
not NOT1 (N11911, N11887);
nand NAND3 (N11912, N11904, N2133, N7722);
nor NOR3 (N11913, N11912, N5550, N1547);
xor XOR2 (N11914, N11909, N3220);
not NOT1 (N11915, N11895);
or OR2 (N11916, N11898, N8438);
buf BUF1 (N11917, N11907);
and AND4 (N11918, N11913, N7725, N9821, N7607);
not NOT1 (N11919, N11905);
nor NOR2 (N11920, N11916, N53);
and AND2 (N11921, N11920, N3938);
buf BUF1 (N11922, N11914);
nor NOR4 (N11923, N11910, N2652, N3101, N1885);
and AND2 (N11924, N11921, N11615);
buf BUF1 (N11925, N11919);
and AND3 (N11926, N11908, N3225, N1366);
not NOT1 (N11927, N11915);
xor XOR2 (N11928, N11911, N10624);
or OR3 (N11929, N11926, N4556, N3027);
nand NAND2 (N11930, N11903, N1539);
and AND3 (N11931, N11928, N7625, N591);
xor XOR2 (N11932, N11917, N8182);
and AND3 (N11933, N11931, N5332, N9666);
nand NAND3 (N11934, N11930, N2132, N3231);
not NOT1 (N11935, N11925);
not NOT1 (N11936, N11918);
nand NAND4 (N11937, N11933, N8741, N10051, N11737);
xor XOR2 (N11938, N11934, N3634);
not NOT1 (N11939, N11923);
or OR2 (N11940, N11939, N6623);
not NOT1 (N11941, N11927);
not NOT1 (N11942, N11938);
xor XOR2 (N11943, N11932, N8155);
buf BUF1 (N11944, N11943);
xor XOR2 (N11945, N11937, N8186);
nand NAND3 (N11946, N11922, N11231, N10851);
and AND2 (N11947, N11936, N2091);
and AND2 (N11948, N11945, N495);
and AND2 (N11949, N11948, N6619);
nand NAND2 (N11950, N11947, N9045);
xor XOR2 (N11951, N11944, N8882);
xor XOR2 (N11952, N11929, N7276);
not NOT1 (N11953, N11949);
nor NOR2 (N11954, N11941, N7165);
not NOT1 (N11955, N11954);
and AND3 (N11956, N11955, N4243, N9403);
nor NOR4 (N11957, N11956, N9170, N6434, N347);
and AND2 (N11958, N11924, N6480);
not NOT1 (N11959, N11935);
or OR2 (N11960, N11940, N1793);
or OR4 (N11961, N11951, N6697, N4954, N2144);
nand NAND2 (N11962, N11946, N441);
nor NOR2 (N11963, N11957, N4340);
nand NAND4 (N11964, N11961, N321, N3749, N2289);
or OR2 (N11965, N11958, N1881);
xor XOR2 (N11966, N11942, N11806);
nand NAND4 (N11967, N11962, N8197, N187, N6171);
or OR2 (N11968, N11966, N10509);
nand NAND2 (N11969, N11968, N9541);
not NOT1 (N11970, N11965);
and AND4 (N11971, N11969, N10073, N3935, N8388);
or OR2 (N11972, N11963, N11179);
and AND2 (N11973, N11952, N4886);
buf BUF1 (N11974, N11972);
buf BUF1 (N11975, N11953);
buf BUF1 (N11976, N11950);
not NOT1 (N11977, N11967);
xor XOR2 (N11978, N11976, N9032);
xor XOR2 (N11979, N11964, N10822);
nor NOR4 (N11980, N11979, N1862, N5545, N5695);
nand NAND4 (N11981, N11960, N5505, N1186, N198);
buf BUF1 (N11982, N11973);
buf BUF1 (N11983, N11977);
not NOT1 (N11984, N11980);
xor XOR2 (N11985, N11959, N2930);
xor XOR2 (N11986, N11982, N428);
not NOT1 (N11987, N11970);
or OR2 (N11988, N11978, N4275);
nor NOR3 (N11989, N11971, N3468, N9723);
nor NOR2 (N11990, N11983, N5045);
nand NAND4 (N11991, N11975, N4982, N11130, N9832);
not NOT1 (N11992, N11985);
nor NOR2 (N11993, N11984, N6125);
not NOT1 (N11994, N11991);
and AND2 (N11995, N11981, N7134);
not NOT1 (N11996, N11988);
not NOT1 (N11997, N11974);
or OR2 (N11998, N11995, N1295);
or OR3 (N11999, N11989, N6213, N7940);
nand NAND3 (N12000, N11993, N3103, N8059);
nand NAND4 (N12001, N11986, N790, N3540, N9290);
and AND3 (N12002, N11999, N8208, N2475);
buf BUF1 (N12003, N11987);
nand NAND2 (N12004, N11997, N6520);
buf BUF1 (N12005, N12004);
and AND4 (N12006, N11996, N6605, N5901, N7936);
and AND3 (N12007, N12006, N2646, N9983);
nor NOR3 (N12008, N12005, N7459, N6229);
xor XOR2 (N12009, N12008, N3893);
nor NOR3 (N12010, N12001, N4661, N8167);
and AND3 (N12011, N12002, N8513, N8561);
xor XOR2 (N12012, N11998, N6621);
xor XOR2 (N12013, N12003, N2246);
nor NOR4 (N12014, N11990, N9066, N33, N5128);
nand NAND4 (N12015, N11992, N7706, N4807, N6882);
and AND3 (N12016, N12012, N985, N8109);
nand NAND3 (N12017, N12011, N4682, N4274);
nand NAND3 (N12018, N12000, N7340, N2406);
buf BUF1 (N12019, N12014);
not NOT1 (N12020, N12013);
nor NOR2 (N12021, N12018, N6352);
or OR3 (N12022, N12010, N10190, N10530);
or OR4 (N12023, N12021, N6590, N11703, N9472);
not NOT1 (N12024, N12007);
not NOT1 (N12025, N11994);
and AND4 (N12026, N12024, N7200, N973, N170);
nand NAND4 (N12027, N12023, N506, N194, N6730);
buf BUF1 (N12028, N12022);
xor XOR2 (N12029, N12009, N5858);
or OR4 (N12030, N12015, N6123, N3627, N2229);
xor XOR2 (N12031, N12019, N5868);
not NOT1 (N12032, N12025);
not NOT1 (N12033, N12016);
or OR2 (N12034, N12027, N1587);
or OR4 (N12035, N12017, N3239, N3482, N5901);
xor XOR2 (N12036, N12026, N10142);
and AND2 (N12037, N12032, N10458);
and AND3 (N12038, N12035, N878, N5752);
buf BUF1 (N12039, N12031);
buf BUF1 (N12040, N12037);
not NOT1 (N12041, N12029);
and AND3 (N12042, N12034, N11368, N785);
not NOT1 (N12043, N12020);
nand NAND2 (N12044, N12041, N5335);
and AND4 (N12045, N12042, N2363, N9150, N3841);
nand NAND3 (N12046, N12043, N347, N9737);
not NOT1 (N12047, N12028);
nor NOR4 (N12048, N12040, N5491, N6838, N5193);
and AND3 (N12049, N12048, N2063, N5178);
and AND4 (N12050, N12049, N7543, N4561, N3982);
buf BUF1 (N12051, N12050);
or OR3 (N12052, N12030, N2448, N526);
or OR4 (N12053, N12052, N10772, N4961, N4302);
or OR3 (N12054, N12046, N6787, N11921);
xor XOR2 (N12055, N12047, N6198);
or OR2 (N12056, N12055, N5550);
nand NAND3 (N12057, N12053, N9930, N8727);
nand NAND4 (N12058, N12044, N5995, N9597, N1712);
and AND3 (N12059, N12039, N94, N4019);
not NOT1 (N12060, N12038);
not NOT1 (N12061, N12036);
and AND3 (N12062, N12051, N11290, N465);
or OR4 (N12063, N12060, N3631, N2331, N22);
not NOT1 (N12064, N12045);
or OR4 (N12065, N12054, N7139, N2003, N2606);
xor XOR2 (N12066, N12061, N824);
xor XOR2 (N12067, N12065, N7438);
xor XOR2 (N12068, N12062, N4079);
and AND2 (N12069, N12066, N9581);
not NOT1 (N12070, N12064);
xor XOR2 (N12071, N12059, N1046);
xor XOR2 (N12072, N12068, N11248);
and AND3 (N12073, N12071, N6402, N7412);
nand NAND2 (N12074, N12067, N9787);
nand NAND2 (N12075, N12057, N5891);
or OR4 (N12076, N12070, N7457, N7292, N11550);
or OR2 (N12077, N12069, N8439);
xor XOR2 (N12078, N12075, N7988);
nand NAND4 (N12079, N12073, N11462, N6963, N4046);
and AND2 (N12080, N12079, N9591);
xor XOR2 (N12081, N12076, N4210);
or OR4 (N12082, N12063, N10279, N7008, N5033);
nor NOR3 (N12083, N12081, N936, N6343);
buf BUF1 (N12084, N12080);
buf BUF1 (N12085, N12058);
buf BUF1 (N12086, N12083);
xor XOR2 (N12087, N12072, N11753);
or OR4 (N12088, N12074, N2949, N10813, N9231);
nor NOR4 (N12089, N12033, N10211, N346, N9339);
not NOT1 (N12090, N12086);
buf BUF1 (N12091, N12082);
or OR2 (N12092, N12090, N5176);
nand NAND3 (N12093, N12078, N8244, N1275);
xor XOR2 (N12094, N12093, N8363);
and AND3 (N12095, N12077, N5152, N11294);
or OR4 (N12096, N12089, N723, N6084, N2200);
nand NAND2 (N12097, N12096, N10804);
buf BUF1 (N12098, N12085);
nor NOR4 (N12099, N12095, N6415, N3424, N11879);
xor XOR2 (N12100, N12088, N8437);
or OR2 (N12101, N12091, N6668);
nand NAND4 (N12102, N12101, N7025, N6873, N8740);
nor NOR2 (N12103, N12100, N1978);
or OR4 (N12104, N12084, N5525, N7066, N11196);
buf BUF1 (N12105, N12087);
nor NOR3 (N12106, N12056, N10190, N1571);
not NOT1 (N12107, N12103);
xor XOR2 (N12108, N12107, N2090);
nor NOR3 (N12109, N12106, N7265, N3416);
nor NOR3 (N12110, N12102, N3688, N6784);
not NOT1 (N12111, N12097);
and AND4 (N12112, N12092, N7829, N7805, N11855);
nor NOR3 (N12113, N12104, N10889, N4219);
or OR4 (N12114, N12111, N3366, N7410, N10146);
nor NOR2 (N12115, N12094, N7691);
nand NAND3 (N12116, N12113, N5244, N7520);
nor NOR4 (N12117, N12098, N8851, N4106, N8444);
nor NOR4 (N12118, N12105, N11914, N12041, N10996);
buf BUF1 (N12119, N12110);
nand NAND4 (N12120, N12108, N2423, N9713, N10232);
nand NAND2 (N12121, N12099, N3786);
and AND2 (N12122, N12119, N5727);
or OR4 (N12123, N12121, N3360, N3231, N5303);
buf BUF1 (N12124, N12123);
xor XOR2 (N12125, N12112, N3463);
nand NAND4 (N12126, N12124, N6474, N1801, N621);
nor NOR2 (N12127, N12126, N7437);
not NOT1 (N12128, N12122);
and AND2 (N12129, N12114, N4776);
nand NAND2 (N12130, N12109, N994);
nor NOR2 (N12131, N12117, N6332);
nor NOR2 (N12132, N12128, N6287);
or OR2 (N12133, N12120, N8073);
nor NOR3 (N12134, N12133, N4173, N198);
buf BUF1 (N12135, N12129);
not NOT1 (N12136, N12134);
nand NAND3 (N12137, N12132, N2184, N11284);
buf BUF1 (N12138, N12125);
or OR2 (N12139, N12131, N681);
xor XOR2 (N12140, N12118, N8879);
or OR3 (N12141, N12116, N5160, N508);
xor XOR2 (N12142, N12115, N6908);
xor XOR2 (N12143, N12127, N6370);
nor NOR3 (N12144, N12141, N7871, N2496);
buf BUF1 (N12145, N12137);
nor NOR2 (N12146, N12130, N8608);
not NOT1 (N12147, N12139);
buf BUF1 (N12148, N12135);
and AND2 (N12149, N12140, N3155);
buf BUF1 (N12150, N12147);
nor NOR3 (N12151, N12145, N4359, N4974);
and AND3 (N12152, N12143, N9761, N11283);
and AND4 (N12153, N12148, N2447, N6302, N4833);
nand NAND2 (N12154, N12144, N6545);
and AND4 (N12155, N12149, N6297, N11730, N7798);
or OR2 (N12156, N12152, N6602);
not NOT1 (N12157, N12156);
buf BUF1 (N12158, N12153);
nand NAND2 (N12159, N12151, N2093);
or OR3 (N12160, N12158, N11790, N55);
and AND2 (N12161, N12160, N3009);
and AND2 (N12162, N12159, N10943);
buf BUF1 (N12163, N12162);
nor NOR3 (N12164, N12146, N11703, N9734);
and AND4 (N12165, N12136, N1824, N11749, N8356);
not NOT1 (N12166, N12155);
or OR4 (N12167, N12166, N11845, N5052, N5039);
nor NOR2 (N12168, N12163, N10333);
or OR2 (N12169, N12154, N693);
nor NOR2 (N12170, N12168, N11010);
nor NOR4 (N12171, N12170, N899, N11496, N3022);
nand NAND3 (N12172, N12138, N8477, N5850);
nand NAND2 (N12173, N12157, N7622);
or OR3 (N12174, N12161, N5608, N7750);
nand NAND4 (N12175, N12169, N10277, N9598, N5708);
not NOT1 (N12176, N12175);
nand NAND3 (N12177, N12173, N1280, N11083);
buf BUF1 (N12178, N12142);
nor NOR3 (N12179, N12150, N6429, N7911);
nor NOR4 (N12180, N12164, N8717, N1762, N4475);
not NOT1 (N12181, N12171);
nor NOR4 (N12182, N12167, N817, N29, N2606);
and AND2 (N12183, N12182, N9794);
nand NAND4 (N12184, N12183, N11017, N209, N8616);
or OR4 (N12185, N12178, N974, N3338, N5494);
xor XOR2 (N12186, N12180, N2626);
or OR3 (N12187, N12174, N4995, N2667);
or OR4 (N12188, N12185, N1544, N8587, N932);
nor NOR3 (N12189, N12179, N6149, N630);
or OR2 (N12190, N12188, N4450);
and AND3 (N12191, N12165, N8563, N8301);
and AND4 (N12192, N12172, N10923, N8361, N5305);
buf BUF1 (N12193, N12190);
or OR4 (N12194, N12186, N11428, N5281, N6034);
nand NAND4 (N12195, N12187, N9764, N6533, N4838);
not NOT1 (N12196, N12191);
buf BUF1 (N12197, N12196);
xor XOR2 (N12198, N12197, N10658);
or OR2 (N12199, N12181, N3998);
and AND2 (N12200, N12194, N7783);
xor XOR2 (N12201, N12177, N1136);
nor NOR2 (N12202, N12189, N8412);
not NOT1 (N12203, N12202);
buf BUF1 (N12204, N12201);
not NOT1 (N12205, N12184);
not NOT1 (N12206, N12193);
nor NOR2 (N12207, N12195, N10711);
nor NOR2 (N12208, N12203, N4158);
buf BUF1 (N12209, N12200);
xor XOR2 (N12210, N12208, N8507);
xor XOR2 (N12211, N12207, N10380);
nand NAND4 (N12212, N12204, N6075, N7897, N4140);
buf BUF1 (N12213, N12212);
not NOT1 (N12214, N12176);
xor XOR2 (N12215, N12192, N11764);
buf BUF1 (N12216, N12199);
nand NAND4 (N12217, N12211, N10804, N1193, N9894);
and AND2 (N12218, N12205, N4485);
and AND4 (N12219, N12215, N2557, N515, N449);
or OR4 (N12220, N12217, N886, N6614, N2773);
or OR3 (N12221, N12198, N2997, N7076);
nand NAND4 (N12222, N12209, N12004, N5729, N2512);
xor XOR2 (N12223, N12216, N284);
xor XOR2 (N12224, N12221, N2126);
not NOT1 (N12225, N12214);
and AND3 (N12226, N12225, N10962, N11520);
xor XOR2 (N12227, N12206, N2673);
or OR3 (N12228, N12210, N3504, N7196);
nor NOR4 (N12229, N12228, N88, N10932, N11350);
not NOT1 (N12230, N12229);
nor NOR3 (N12231, N12224, N3622, N11639);
buf BUF1 (N12232, N12220);
nand NAND2 (N12233, N12213, N5430);
nor NOR3 (N12234, N12232, N4783, N6021);
or OR3 (N12235, N12222, N11479, N8056);
or OR4 (N12236, N12230, N10912, N4425, N11013);
xor XOR2 (N12237, N12236, N3087);
or OR3 (N12238, N12227, N8376, N10853);
xor XOR2 (N12239, N12238, N2827);
buf BUF1 (N12240, N12234);
nand NAND3 (N12241, N12240, N12023, N2710);
buf BUF1 (N12242, N12235);
buf BUF1 (N12243, N12237);
buf BUF1 (N12244, N12233);
and AND3 (N12245, N12226, N1953, N4580);
xor XOR2 (N12246, N12239, N6396);
nand NAND2 (N12247, N12218, N9986);
and AND3 (N12248, N12246, N3107, N7439);
and AND4 (N12249, N12243, N4512, N11451, N7952);
buf BUF1 (N12250, N12244);
and AND4 (N12251, N12250, N2145, N6781, N2312);
and AND3 (N12252, N12247, N11408, N12146);
nor NOR2 (N12253, N12242, N10031);
xor XOR2 (N12254, N12231, N5883);
buf BUF1 (N12255, N12245);
and AND4 (N12256, N12253, N6843, N9863, N11854);
or OR2 (N12257, N12251, N3044);
nand NAND4 (N12258, N12256, N8634, N628, N6638);
or OR3 (N12259, N12219, N9456, N2098);
nor NOR4 (N12260, N12258, N10743, N1432, N10045);
buf BUF1 (N12261, N12252);
nand NAND4 (N12262, N12254, N3615, N5436, N10524);
nor NOR2 (N12263, N12260, N7687);
xor XOR2 (N12264, N12249, N5213);
and AND2 (N12265, N12262, N468);
nand NAND3 (N12266, N12255, N2304, N6638);
xor XOR2 (N12267, N12264, N7919);
buf BUF1 (N12268, N12267);
or OR4 (N12269, N12248, N12239, N9972, N8846);
or OR2 (N12270, N12268, N74);
nor NOR2 (N12271, N12269, N1447);
not NOT1 (N12272, N12270);
xor XOR2 (N12273, N12259, N3307);
nand NAND3 (N12274, N12261, N8974, N9580);
nand NAND4 (N12275, N12271, N11633, N7861, N6752);
and AND2 (N12276, N12265, N10171);
nand NAND3 (N12277, N12263, N5840, N12006);
nand NAND3 (N12278, N12275, N4916, N8998);
xor XOR2 (N12279, N12257, N11363);
not NOT1 (N12280, N12278);
not NOT1 (N12281, N12279);
xor XOR2 (N12282, N12280, N9697);
nand NAND2 (N12283, N12281, N5935);
buf BUF1 (N12284, N12277);
or OR4 (N12285, N12276, N5061, N2194, N11566);
nor NOR2 (N12286, N12274, N2224);
or OR4 (N12287, N12273, N8033, N6139, N6038);
nand NAND3 (N12288, N12282, N5999, N7901);
buf BUF1 (N12289, N12288);
nor NOR4 (N12290, N12266, N1584, N7336, N12094);
not NOT1 (N12291, N12285);
buf BUF1 (N12292, N12284);
nor NOR3 (N12293, N12286, N9487, N3247);
buf BUF1 (N12294, N12223);
nor NOR3 (N12295, N12293, N3487, N2790);
nor NOR3 (N12296, N12292, N1679, N10907);
or OR2 (N12297, N12296, N11657);
buf BUF1 (N12298, N12295);
nor NOR2 (N12299, N12272, N2129);
nand NAND2 (N12300, N12291, N8787);
buf BUF1 (N12301, N12241);
buf BUF1 (N12302, N12298);
nand NAND4 (N12303, N12283, N7364, N5845, N4259);
nor NOR2 (N12304, N12299, N8640);
nor NOR3 (N12305, N12301, N1828, N10066);
nor NOR2 (N12306, N12305, N7246);
not NOT1 (N12307, N12290);
not NOT1 (N12308, N12302);
not NOT1 (N12309, N12287);
nand NAND4 (N12310, N12289, N2470, N4663, N3890);
xor XOR2 (N12311, N12303, N10846);
xor XOR2 (N12312, N12311, N4590);
and AND3 (N12313, N12306, N9074, N11505);
xor XOR2 (N12314, N12308, N3058);
buf BUF1 (N12315, N12312);
buf BUF1 (N12316, N12315);
or OR3 (N12317, N12316, N9819, N4634);
xor XOR2 (N12318, N12310, N159);
or OR3 (N12319, N12313, N2207, N2573);
xor XOR2 (N12320, N12318, N11300);
or OR2 (N12321, N12304, N2639);
or OR2 (N12322, N12300, N8507);
buf BUF1 (N12323, N12319);
or OR2 (N12324, N12309, N9404);
buf BUF1 (N12325, N12314);
and AND2 (N12326, N12307, N4630);
and AND4 (N12327, N12321, N9859, N7938, N914);
or OR2 (N12328, N12320, N90);
or OR4 (N12329, N12323, N4243, N162, N8344);
or OR3 (N12330, N12317, N1799, N8518);
not NOT1 (N12331, N12322);
buf BUF1 (N12332, N12328);
not NOT1 (N12333, N12329);
nor NOR2 (N12334, N12294, N11786);
xor XOR2 (N12335, N12332, N10752);
nor NOR3 (N12336, N12325, N1591, N7086);
nor NOR3 (N12337, N12330, N7167, N7655);
or OR2 (N12338, N12324, N5394);
buf BUF1 (N12339, N12336);
nor NOR3 (N12340, N12331, N4891, N4839);
not NOT1 (N12341, N12334);
or OR2 (N12342, N12297, N551);
xor XOR2 (N12343, N12342, N1658);
or OR4 (N12344, N12335, N4763, N2964, N9503);
or OR4 (N12345, N12338, N6313, N8786, N2623);
not NOT1 (N12346, N12337);
buf BUF1 (N12347, N12345);
xor XOR2 (N12348, N12333, N8480);
nand NAND3 (N12349, N12346, N10138, N3520);
or OR2 (N12350, N12348, N2245);
buf BUF1 (N12351, N12349);
buf BUF1 (N12352, N12344);
nor NOR4 (N12353, N12351, N6819, N2722, N9277);
not NOT1 (N12354, N12341);
and AND4 (N12355, N12350, N2253, N11084, N5837);
xor XOR2 (N12356, N12353, N5126);
or OR4 (N12357, N12352, N12145, N9410, N4886);
or OR4 (N12358, N12354, N1674, N10733, N9001);
and AND2 (N12359, N12339, N7666);
nor NOR3 (N12360, N12358, N6830, N6890);
not NOT1 (N12361, N12356);
not NOT1 (N12362, N12360);
buf BUF1 (N12363, N12355);
nor NOR3 (N12364, N12359, N3804, N10241);
or OR4 (N12365, N12340, N11296, N8346, N1870);
buf BUF1 (N12366, N12327);
buf BUF1 (N12367, N12363);
xor XOR2 (N12368, N12364, N9968);
and AND3 (N12369, N12357, N9173, N6164);
buf BUF1 (N12370, N12347);
not NOT1 (N12371, N12362);
xor XOR2 (N12372, N12326, N9851);
buf BUF1 (N12373, N12370);
not NOT1 (N12374, N12361);
nor NOR2 (N12375, N12373, N9404);
xor XOR2 (N12376, N12343, N5631);
buf BUF1 (N12377, N12372);
nand NAND2 (N12378, N12368, N5410);
buf BUF1 (N12379, N12378);
buf BUF1 (N12380, N12365);
nor NOR3 (N12381, N12371, N9555, N6645);
or OR4 (N12382, N12380, N2257, N7754, N11006);
buf BUF1 (N12383, N12374);
or OR3 (N12384, N12382, N6045, N11211);
xor XOR2 (N12385, N12375, N12153);
or OR3 (N12386, N12381, N7714, N8701);
or OR3 (N12387, N12385, N985, N6053);
not NOT1 (N12388, N12383);
buf BUF1 (N12389, N12384);
nand NAND2 (N12390, N12366, N6167);
buf BUF1 (N12391, N12389);
or OR2 (N12392, N12386, N473);
nor NOR4 (N12393, N12388, N7064, N4864, N2843);
and AND4 (N12394, N12376, N7482, N7106, N3265);
nand NAND3 (N12395, N12392, N2844, N11087);
and AND3 (N12396, N12387, N5334, N5440);
buf BUF1 (N12397, N12396);
nand NAND4 (N12398, N12390, N3487, N8791, N9236);
and AND4 (N12399, N12379, N11299, N10692, N5966);
nor NOR3 (N12400, N12397, N233, N12134);
not NOT1 (N12401, N12369);
xor XOR2 (N12402, N12391, N864);
or OR4 (N12403, N12402, N11242, N4453, N6875);
and AND3 (N12404, N12377, N3531, N11281);
or OR3 (N12405, N12393, N10748, N1641);
nand NAND3 (N12406, N12405, N3931, N6261);
buf BUF1 (N12407, N12398);
xor XOR2 (N12408, N12367, N1857);
or OR4 (N12409, N12394, N12054, N6415, N6768);
buf BUF1 (N12410, N12401);
nand NAND2 (N12411, N12400, N8388);
nand NAND4 (N12412, N12395, N174, N2778, N9864);
nand NAND4 (N12413, N12407, N807, N6147, N11779);
or OR4 (N12414, N12411, N2594, N111, N11297);
nor NOR4 (N12415, N12399, N9688, N9211, N4742);
nor NOR4 (N12416, N12413, N5037, N843, N3820);
xor XOR2 (N12417, N12409, N1821);
nand NAND3 (N12418, N12408, N8444, N8497);
not NOT1 (N12419, N12404);
not NOT1 (N12420, N12418);
or OR4 (N12421, N12403, N2879, N1189, N546);
and AND4 (N12422, N12414, N9748, N889, N5681);
not NOT1 (N12423, N12412);
nand NAND4 (N12424, N12421, N2219, N11556, N5847);
nor NOR2 (N12425, N12419, N10717);
nand NAND4 (N12426, N12422, N3691, N12127, N9355);
and AND4 (N12427, N12424, N7193, N12340, N6994);
not NOT1 (N12428, N12410);
buf BUF1 (N12429, N12406);
or OR3 (N12430, N12427, N737, N7361);
not NOT1 (N12431, N12415);
not NOT1 (N12432, N12426);
nand NAND4 (N12433, N12423, N4418, N7373, N1321);
not NOT1 (N12434, N12428);
not NOT1 (N12435, N12429);
not NOT1 (N12436, N12417);
or OR4 (N12437, N12434, N9502, N3783, N2825);
buf BUF1 (N12438, N12416);
and AND2 (N12439, N12420, N12316);
not NOT1 (N12440, N12439);
nand NAND3 (N12441, N12438, N1929, N3538);
xor XOR2 (N12442, N12431, N420);
buf BUF1 (N12443, N12432);
nor NOR4 (N12444, N12425, N6799, N2183, N6463);
nand NAND2 (N12445, N12435, N5240);
and AND3 (N12446, N12437, N7438, N8830);
nor NOR3 (N12447, N12440, N757, N9229);
nor NOR4 (N12448, N12446, N7988, N256, N8258);
or OR2 (N12449, N12442, N7963);
nor NOR3 (N12450, N12448, N4049, N5285);
or OR3 (N12451, N12436, N8538, N12136);
xor XOR2 (N12452, N12444, N1871);
nor NOR2 (N12453, N12445, N5716);
buf BUF1 (N12454, N12441);
nor NOR4 (N12455, N12453, N4527, N10431, N3989);
buf BUF1 (N12456, N12447);
nor NOR4 (N12457, N12454, N1794, N7336, N6533);
or OR3 (N12458, N12451, N11214, N5082);
nor NOR3 (N12459, N12458, N1618, N9165);
or OR2 (N12460, N12455, N10695);
not NOT1 (N12461, N12430);
not NOT1 (N12462, N12452);
not NOT1 (N12463, N12456);
and AND4 (N12464, N12457, N1868, N1328, N1202);
xor XOR2 (N12465, N12450, N9661);
and AND4 (N12466, N12460, N5703, N1997, N7244);
nand NAND4 (N12467, N12463, N2921, N3725, N8877);
or OR3 (N12468, N12461, N11949, N6192);
and AND4 (N12469, N12459, N2070, N1756, N3182);
and AND4 (N12470, N12449, N6880, N1782, N10023);
xor XOR2 (N12471, N12443, N8271);
not NOT1 (N12472, N12466);
or OR4 (N12473, N12462, N1846, N10301, N3392);
not NOT1 (N12474, N12465);
and AND4 (N12475, N12469, N4239, N11913, N4022);
or OR4 (N12476, N12433, N2207, N2042, N999);
buf BUF1 (N12477, N12467);
or OR2 (N12478, N12470, N11584);
xor XOR2 (N12479, N12473, N599);
buf BUF1 (N12480, N12472);
not NOT1 (N12481, N12474);
and AND4 (N12482, N12481, N7538, N9343, N4261);
not NOT1 (N12483, N12475);
and AND2 (N12484, N12479, N9883);
not NOT1 (N12485, N12468);
nand NAND4 (N12486, N12482, N8162, N6520, N10020);
nor NOR3 (N12487, N12484, N4204, N6172);
not NOT1 (N12488, N12486);
not NOT1 (N12489, N12477);
not NOT1 (N12490, N12488);
or OR2 (N12491, N12490, N12489);
nor NOR4 (N12492, N2443, N2354, N7537, N3399);
buf BUF1 (N12493, N12491);
nand NAND3 (N12494, N12493, N1148, N11728);
xor XOR2 (N12495, N12480, N10759);
nand NAND3 (N12496, N12492, N4840, N11014);
xor XOR2 (N12497, N12485, N7636);
nand NAND4 (N12498, N12496, N8572, N9110, N3379);
buf BUF1 (N12499, N12476);
xor XOR2 (N12500, N12495, N1116);
nor NOR4 (N12501, N12464, N8419, N6280, N11419);
not NOT1 (N12502, N12501);
xor XOR2 (N12503, N12483, N6842);
not NOT1 (N12504, N12494);
nor NOR2 (N12505, N12497, N3608);
nand NAND3 (N12506, N12503, N1034, N9117);
nor NOR4 (N12507, N12504, N10463, N2781, N6552);
xor XOR2 (N12508, N12471, N11453);
and AND2 (N12509, N12499, N11758);
nand NAND4 (N12510, N12507, N9038, N6066, N1971);
buf BUF1 (N12511, N12487);
nand NAND4 (N12512, N12509, N5871, N5746, N1452);
nand NAND3 (N12513, N12510, N4616, N1929);
xor XOR2 (N12514, N12498, N11034);
and AND3 (N12515, N12512, N8314, N9743);
xor XOR2 (N12516, N12506, N11085);
nor NOR2 (N12517, N12502, N11354);
and AND4 (N12518, N12478, N2938, N8428, N12312);
not NOT1 (N12519, N12505);
not NOT1 (N12520, N12508);
buf BUF1 (N12521, N12513);
or OR4 (N12522, N12515, N4540, N1652, N10683);
buf BUF1 (N12523, N12519);
not NOT1 (N12524, N12500);
and AND4 (N12525, N12518, N2725, N5270, N5480);
not NOT1 (N12526, N12523);
buf BUF1 (N12527, N12522);
nand NAND2 (N12528, N12524, N9354);
buf BUF1 (N12529, N12517);
or OR2 (N12530, N12514, N4781);
nand NAND2 (N12531, N12526, N5333);
nor NOR3 (N12532, N12529, N8073, N7656);
buf BUF1 (N12533, N12528);
or OR4 (N12534, N12521, N7410, N3393, N6085);
nor NOR4 (N12535, N12531, N7487, N9734, N7034);
not NOT1 (N12536, N12511);
and AND4 (N12537, N12535, N2285, N8492, N3514);
or OR2 (N12538, N12537, N2455);
not NOT1 (N12539, N12536);
xor XOR2 (N12540, N12530, N7449);
buf BUF1 (N12541, N12540);
nand NAND3 (N12542, N12516, N8334, N868);
buf BUF1 (N12543, N12539);
and AND4 (N12544, N12534, N4978, N8263, N9144);
not NOT1 (N12545, N12542);
buf BUF1 (N12546, N12532);
xor XOR2 (N12547, N12527, N11824);
xor XOR2 (N12548, N12538, N8276);
not NOT1 (N12549, N12541);
nor NOR4 (N12550, N12548, N3777, N10292, N1882);
or OR2 (N12551, N12525, N9615);
and AND3 (N12552, N12545, N4874, N5745);
and AND3 (N12553, N12550, N1624, N10031);
and AND4 (N12554, N12533, N863, N8635, N9020);
xor XOR2 (N12555, N12544, N7013);
nor NOR3 (N12556, N12546, N1025, N4929);
or OR4 (N12557, N12547, N4456, N1899, N5552);
not NOT1 (N12558, N12549);
not NOT1 (N12559, N12556);
and AND3 (N12560, N12551, N85, N4856);
buf BUF1 (N12561, N12553);
not NOT1 (N12562, N12554);
nor NOR2 (N12563, N12555, N6201);
nand NAND3 (N12564, N12562, N6638, N5931);
nand NAND4 (N12565, N12552, N5899, N6922, N12434);
or OR2 (N12566, N12564, N6479);
nor NOR3 (N12567, N12560, N1249, N11997);
xor XOR2 (N12568, N12557, N236);
not NOT1 (N12569, N12543);
and AND2 (N12570, N12569, N10327);
buf BUF1 (N12571, N12566);
nor NOR4 (N12572, N12565, N11512, N6167, N4689);
xor XOR2 (N12573, N12567, N4220);
nand NAND4 (N12574, N12568, N9224, N6672, N3064);
and AND2 (N12575, N12558, N1199);
buf BUF1 (N12576, N12559);
nor NOR2 (N12577, N12573, N6811);
xor XOR2 (N12578, N12561, N6694);
and AND3 (N12579, N12576, N9531, N5391);
and AND4 (N12580, N12563, N6223, N9665, N8659);
xor XOR2 (N12581, N12572, N12062);
nor NOR4 (N12582, N12579, N11267, N9929, N7709);
and AND2 (N12583, N12581, N8571);
buf BUF1 (N12584, N12583);
nand NAND3 (N12585, N12575, N8344, N7188);
or OR4 (N12586, N12520, N3498, N1945, N10787);
or OR2 (N12587, N12585, N7222);
nand NAND4 (N12588, N12570, N10471, N2078, N2145);
not NOT1 (N12589, N12580);
or OR3 (N12590, N12574, N3813, N10104);
not NOT1 (N12591, N12584);
not NOT1 (N12592, N12590);
nor NOR2 (N12593, N12578, N2835);
and AND3 (N12594, N12593, N1218, N7979);
not NOT1 (N12595, N12591);
buf BUF1 (N12596, N12588);
or OR2 (N12597, N12582, N10328);
nand NAND2 (N12598, N12587, N10580);
and AND2 (N12599, N12589, N10747);
nand NAND3 (N12600, N12599, N10708, N1436);
not NOT1 (N12601, N12598);
buf BUF1 (N12602, N12596);
not NOT1 (N12603, N12577);
nand NAND4 (N12604, N12586, N8704, N5327, N8658);
xor XOR2 (N12605, N12597, N1169);
nor NOR4 (N12606, N12603, N8408, N830, N4894);
buf BUF1 (N12607, N12600);
and AND3 (N12608, N12605, N4724, N451);
and AND4 (N12609, N12595, N974, N985, N4539);
not NOT1 (N12610, N12604);
and AND4 (N12611, N12571, N10642, N517, N362);
buf BUF1 (N12612, N12608);
nor NOR3 (N12613, N12602, N9507, N9616);
or OR3 (N12614, N12610, N6801, N10450);
nand NAND3 (N12615, N12607, N1383, N3131);
buf BUF1 (N12616, N12592);
nor NOR4 (N12617, N12609, N9634, N2331, N9147);
buf BUF1 (N12618, N12594);
not NOT1 (N12619, N12613);
buf BUF1 (N12620, N12614);
buf BUF1 (N12621, N12601);
buf BUF1 (N12622, N12612);
and AND3 (N12623, N12616, N5032, N1393);
buf BUF1 (N12624, N12619);
xor XOR2 (N12625, N12615, N3222);
and AND2 (N12626, N12624, N3594);
not NOT1 (N12627, N12625);
and AND2 (N12628, N12623, N3468);
and AND4 (N12629, N12622, N11227, N9795, N1808);
not NOT1 (N12630, N12611);
not NOT1 (N12631, N12606);
and AND4 (N12632, N12617, N6930, N10890, N1580);
xor XOR2 (N12633, N12629, N10725);
and AND2 (N12634, N12628, N7913);
nand NAND2 (N12635, N12630, N8212);
nand NAND3 (N12636, N12631, N8864, N3348);
nor NOR3 (N12637, N12633, N9002, N5547);
xor XOR2 (N12638, N12618, N7392);
buf BUF1 (N12639, N12636);
not NOT1 (N12640, N12637);
buf BUF1 (N12641, N12620);
not NOT1 (N12642, N12627);
buf BUF1 (N12643, N12641);
or OR4 (N12644, N12639, N4682, N8407, N2855);
xor XOR2 (N12645, N12644, N10801);
nand NAND4 (N12646, N12632, N11704, N2118, N6978);
not NOT1 (N12647, N12646);
or OR2 (N12648, N12634, N10368);
xor XOR2 (N12649, N12648, N6179);
buf BUF1 (N12650, N12638);
nor NOR3 (N12651, N12621, N1217, N10681);
or OR4 (N12652, N12640, N170, N4762, N7560);
nor NOR3 (N12653, N12649, N6233, N70);
xor XOR2 (N12654, N12647, N12443);
nor NOR2 (N12655, N12653, N4961);
buf BUF1 (N12656, N12654);
and AND3 (N12657, N12650, N7925, N8171);
nand NAND3 (N12658, N12642, N10840, N87);
buf BUF1 (N12659, N12635);
xor XOR2 (N12660, N12657, N10673);
nand NAND2 (N12661, N12651, N1673);
or OR3 (N12662, N12643, N5290, N3411);
or OR3 (N12663, N12655, N4072, N4929);
nand NAND3 (N12664, N12662, N10142, N6657);
nand NAND3 (N12665, N12652, N2564, N4889);
buf BUF1 (N12666, N12661);
or OR2 (N12667, N12666, N7178);
nor NOR2 (N12668, N12660, N4177);
xor XOR2 (N12669, N12664, N2400);
or OR3 (N12670, N12659, N12214, N6344);
not NOT1 (N12671, N12665);
and AND4 (N12672, N12670, N9645, N1561, N10238);
or OR2 (N12673, N12671, N6146);
not NOT1 (N12674, N12626);
and AND3 (N12675, N12668, N10532, N11711);
and AND2 (N12676, N12645, N6284);
not NOT1 (N12677, N12676);
xor XOR2 (N12678, N12667, N23);
and AND2 (N12679, N12656, N10081);
xor XOR2 (N12680, N12679, N4683);
nand NAND4 (N12681, N12678, N2226, N12177, N10598);
nand NAND3 (N12682, N12669, N7899, N5513);
or OR4 (N12683, N12663, N4550, N5668, N12164);
nand NAND2 (N12684, N12677, N6092);
nor NOR2 (N12685, N12675, N1516);
not NOT1 (N12686, N12681);
xor XOR2 (N12687, N12672, N5160);
and AND4 (N12688, N12680, N1266, N1232, N5451);
xor XOR2 (N12689, N12673, N5309);
buf BUF1 (N12690, N12658);
xor XOR2 (N12691, N12690, N1056);
nand NAND4 (N12692, N12687, N11617, N5860, N5958);
buf BUF1 (N12693, N12686);
nand NAND3 (N12694, N12688, N9099, N10573);
xor XOR2 (N12695, N12683, N591);
not NOT1 (N12696, N12682);
or OR2 (N12697, N12695, N12577);
and AND2 (N12698, N12674, N9873);
not NOT1 (N12699, N12697);
or OR2 (N12700, N12694, N12384);
or OR2 (N12701, N12698, N7301);
xor XOR2 (N12702, N12689, N8924);
and AND4 (N12703, N12691, N1108, N10743, N7847);
buf BUF1 (N12704, N12684);
nor NOR4 (N12705, N12693, N2713, N11028, N9915);
nand NAND3 (N12706, N12703, N11134, N10657);
nor NOR2 (N12707, N12696, N11444);
nor NOR4 (N12708, N12705, N6492, N7698, N8753);
not NOT1 (N12709, N12706);
and AND4 (N12710, N12699, N7838, N5649, N2508);
xor XOR2 (N12711, N12685, N278);
buf BUF1 (N12712, N12708);
and AND2 (N12713, N12702, N10580);
buf BUF1 (N12714, N12713);
and AND3 (N12715, N12704, N2141, N6983);
buf BUF1 (N12716, N12700);
xor XOR2 (N12717, N12707, N9757);
nand NAND4 (N12718, N12715, N8104, N1472, N10874);
and AND2 (N12719, N12712, N6520);
nor NOR2 (N12720, N12719, N1288);
or OR4 (N12721, N12718, N3779, N8391, N7799);
not NOT1 (N12722, N12714);
not NOT1 (N12723, N12711);
and AND4 (N12724, N12720, N11820, N8527, N9307);
nand NAND3 (N12725, N12710, N3538, N7484);
nand NAND3 (N12726, N12701, N12279, N3012);
not NOT1 (N12727, N12692);
and AND2 (N12728, N12709, N7887);
buf BUF1 (N12729, N12725);
nand NAND4 (N12730, N12727, N3551, N4710, N12179);
nor NOR3 (N12731, N12729, N8630, N8289);
not NOT1 (N12732, N12722);
nand NAND2 (N12733, N12716, N12651);
not NOT1 (N12734, N12730);
buf BUF1 (N12735, N12726);
xor XOR2 (N12736, N12735, N6918);
and AND4 (N12737, N12733, N12030, N6141, N10707);
and AND3 (N12738, N12731, N12286, N4336);
nand NAND4 (N12739, N12734, N6716, N4803, N3620);
nand NAND4 (N12740, N12739, N480, N11150, N3365);
and AND4 (N12741, N12732, N9973, N3154, N8121);
or OR3 (N12742, N12741, N8666, N625);
nand NAND3 (N12743, N12742, N4133, N5456);
nor NOR2 (N12744, N12736, N12548);
xor XOR2 (N12745, N12737, N6700);
xor XOR2 (N12746, N12728, N1078);
and AND2 (N12747, N12721, N6044);
or OR2 (N12748, N12740, N10797);
and AND3 (N12749, N12724, N11056, N9372);
not NOT1 (N12750, N12717);
not NOT1 (N12751, N12748);
buf BUF1 (N12752, N12744);
and AND4 (N12753, N12745, N278, N7429, N606);
xor XOR2 (N12754, N12723, N10384);
xor XOR2 (N12755, N12738, N4832);
buf BUF1 (N12756, N12749);
not NOT1 (N12757, N12754);
or OR2 (N12758, N12756, N3775);
xor XOR2 (N12759, N12755, N9727);
and AND2 (N12760, N12751, N12736);
and AND3 (N12761, N12757, N3707, N4581);
xor XOR2 (N12762, N12753, N8128);
nand NAND2 (N12763, N12762, N7521);
nand NAND2 (N12764, N12761, N465);
xor XOR2 (N12765, N12758, N620);
nand NAND3 (N12766, N12750, N11759, N6284);
buf BUF1 (N12767, N12747);
and AND3 (N12768, N12760, N4347, N11604);
or OR3 (N12769, N12765, N120, N12301);
xor XOR2 (N12770, N12766, N6994);
or OR3 (N12771, N12769, N7644, N2049);
nor NOR3 (N12772, N12759, N5481, N9493);
xor XOR2 (N12773, N12771, N8122);
nor NOR2 (N12774, N12767, N9126);
buf BUF1 (N12775, N12772);
not NOT1 (N12776, N12763);
nand NAND3 (N12777, N12764, N3565, N3549);
or OR3 (N12778, N12752, N7861, N4882);
not NOT1 (N12779, N12768);
or OR2 (N12780, N12774, N7990);
and AND4 (N12781, N12773, N583, N7959, N12729);
nor NOR3 (N12782, N12775, N7805, N9509);
buf BUF1 (N12783, N12743);
xor XOR2 (N12784, N12781, N5775);
buf BUF1 (N12785, N12746);
or OR3 (N12786, N12783, N11735, N6747);
buf BUF1 (N12787, N12782);
not NOT1 (N12788, N12780);
nor NOR3 (N12789, N12776, N9789, N10252);
not NOT1 (N12790, N12787);
not NOT1 (N12791, N12779);
not NOT1 (N12792, N12778);
and AND3 (N12793, N12777, N6449, N8254);
buf BUF1 (N12794, N12791);
buf BUF1 (N12795, N12784);
buf BUF1 (N12796, N12770);
xor XOR2 (N12797, N12796, N10854);
xor XOR2 (N12798, N12797, N1402);
nor NOR2 (N12799, N12788, N6652);
and AND2 (N12800, N12785, N4602);
nor NOR4 (N12801, N12798, N1873, N12759, N9597);
not NOT1 (N12802, N12795);
not NOT1 (N12803, N12801);
buf BUF1 (N12804, N12803);
and AND4 (N12805, N12793, N6914, N5657, N2770);
xor XOR2 (N12806, N12805, N10468);
or OR4 (N12807, N12789, N4719, N8579, N1338);
or OR4 (N12808, N12790, N2280, N8885, N872);
xor XOR2 (N12809, N12804, N11664);
and AND4 (N12810, N12809, N757, N6558, N4708);
not NOT1 (N12811, N12792);
xor XOR2 (N12812, N12811, N7412);
nor NOR3 (N12813, N12808, N2378, N1983);
and AND4 (N12814, N12810, N4690, N10103, N3238);
not NOT1 (N12815, N12794);
nor NOR2 (N12816, N12815, N3503);
or OR3 (N12817, N12816, N6119, N800);
buf BUF1 (N12818, N12806);
not NOT1 (N12819, N12814);
not NOT1 (N12820, N12799);
and AND2 (N12821, N12818, N5569);
xor XOR2 (N12822, N12821, N5227);
buf BUF1 (N12823, N12822);
nor NOR2 (N12824, N12813, N5176);
and AND4 (N12825, N12819, N2251, N5358, N8292);
not NOT1 (N12826, N12800);
nand NAND2 (N12827, N12807, N7648);
nor NOR3 (N12828, N12826, N6814, N8578);
nor NOR3 (N12829, N12802, N10305, N6625);
and AND3 (N12830, N12827, N10416, N10588);
and AND2 (N12831, N12830, N3373);
buf BUF1 (N12832, N12817);
not NOT1 (N12833, N12812);
xor XOR2 (N12834, N12823, N6708);
not NOT1 (N12835, N12786);
nand NAND3 (N12836, N12834, N2728, N2763);
buf BUF1 (N12837, N12836);
and AND4 (N12838, N12820, N7633, N5976, N12322);
nand NAND2 (N12839, N12833, N3182);
or OR4 (N12840, N12838, N4079, N10439, N8119);
xor XOR2 (N12841, N12824, N1542);
xor XOR2 (N12842, N12832, N2255);
nor NOR3 (N12843, N12829, N4843, N5233);
nor NOR3 (N12844, N12837, N9147, N9343);
not NOT1 (N12845, N12825);
nand NAND4 (N12846, N12840, N1190, N10120, N3848);
nand NAND4 (N12847, N12845, N11069, N12182, N8864);
not NOT1 (N12848, N12841);
nand NAND2 (N12849, N12844, N5249);
and AND3 (N12850, N12842, N3119, N10666);
xor XOR2 (N12851, N12849, N6506);
xor XOR2 (N12852, N12843, N5020);
buf BUF1 (N12853, N12839);
nand NAND2 (N12854, N12853, N5271);
nor NOR4 (N12855, N12850, N10636, N6620, N6238);
xor XOR2 (N12856, N12846, N9173);
xor XOR2 (N12857, N12856, N4130);
xor XOR2 (N12858, N12847, N3448);
buf BUF1 (N12859, N12852);
buf BUF1 (N12860, N12831);
not NOT1 (N12861, N12848);
not NOT1 (N12862, N12858);
buf BUF1 (N12863, N12862);
nand NAND2 (N12864, N12857, N6542);
nor NOR2 (N12865, N12835, N1868);
not NOT1 (N12866, N12854);
or OR3 (N12867, N12828, N8916, N7908);
nor NOR3 (N12868, N12866, N6044, N1312);
buf BUF1 (N12869, N12861);
and AND2 (N12870, N12851, N6759);
nor NOR2 (N12871, N12860, N2022);
or OR4 (N12872, N12859, N9434, N5146, N8057);
nand NAND3 (N12873, N12872, N10781, N6569);
and AND3 (N12874, N12869, N4681, N9146);
and AND4 (N12875, N12867, N2165, N11537, N8297);
or OR4 (N12876, N12868, N9535, N12120, N6301);
xor XOR2 (N12877, N12871, N11921);
not NOT1 (N12878, N12865);
buf BUF1 (N12879, N12870);
buf BUF1 (N12880, N12878);
and AND2 (N12881, N12863, N5939);
not NOT1 (N12882, N12877);
buf BUF1 (N12883, N12880);
nor NOR2 (N12884, N12875, N11158);
not NOT1 (N12885, N12879);
not NOT1 (N12886, N12864);
xor XOR2 (N12887, N12883, N8054);
and AND2 (N12888, N12885, N6161);
nor NOR2 (N12889, N12874, N12320);
or OR4 (N12890, N12855, N1227, N2091, N11421);
or OR3 (N12891, N12886, N10972, N11173);
and AND4 (N12892, N12882, N7103, N12120, N10941);
nand NAND4 (N12893, N12892, N8600, N11933, N4465);
nor NOR4 (N12894, N12873, N1358, N11216, N6516);
xor XOR2 (N12895, N12881, N6288);
xor XOR2 (N12896, N12894, N10344);
not NOT1 (N12897, N12895);
nand NAND2 (N12898, N12887, N8438);
and AND4 (N12899, N12898, N10117, N1827, N5293);
and AND3 (N12900, N12884, N10274, N12364);
buf BUF1 (N12901, N12876);
xor XOR2 (N12902, N12890, N12502);
or OR4 (N12903, N12888, N11679, N5292, N5158);
buf BUF1 (N12904, N12889);
xor XOR2 (N12905, N12897, N8760);
xor XOR2 (N12906, N12900, N7964);
and AND4 (N12907, N12905, N12364, N11436, N11440);
not NOT1 (N12908, N12902);
and AND2 (N12909, N12907, N5264);
buf BUF1 (N12910, N12901);
buf BUF1 (N12911, N12893);
not NOT1 (N12912, N12896);
not NOT1 (N12913, N12908);
nor NOR3 (N12914, N12912, N2454, N10190);
nor NOR2 (N12915, N12899, N8025);
buf BUF1 (N12916, N12903);
or OR3 (N12917, N12891, N8442, N7856);
xor XOR2 (N12918, N12909, N5945);
or OR4 (N12919, N12906, N11312, N847, N11671);
nand NAND4 (N12920, N12916, N4730, N9352, N12880);
buf BUF1 (N12921, N12920);
and AND3 (N12922, N12904, N1406, N614);
xor XOR2 (N12923, N12910, N9455);
buf BUF1 (N12924, N12915);
not NOT1 (N12925, N12914);
buf BUF1 (N12926, N12923);
buf BUF1 (N12927, N12926);
nor NOR2 (N12928, N12918, N1892);
xor XOR2 (N12929, N12925, N3263);
and AND4 (N12930, N12917, N7286, N6729, N2263);
buf BUF1 (N12931, N12927);
and AND2 (N12932, N12924, N3106);
not NOT1 (N12933, N12931);
not NOT1 (N12934, N12928);
nor NOR4 (N12935, N12933, N9551, N1094, N1012);
and AND2 (N12936, N12929, N6725);
or OR3 (N12937, N12919, N12927, N2120);
nor NOR4 (N12938, N12930, N2748, N6131, N11973);
buf BUF1 (N12939, N12935);
buf BUF1 (N12940, N12913);
or OR4 (N12941, N12936, N5052, N10942, N4742);
buf BUF1 (N12942, N12932);
not NOT1 (N12943, N12941);
or OR3 (N12944, N12940, N2636, N1227);
nor NOR4 (N12945, N12934, N11192, N6482, N2943);
xor XOR2 (N12946, N12939, N2798);
buf BUF1 (N12947, N12944);
nand NAND4 (N12948, N12911, N3365, N12152, N1385);
and AND4 (N12949, N12937, N380, N2712, N5702);
not NOT1 (N12950, N12921);
buf BUF1 (N12951, N12946);
nor NOR4 (N12952, N12947, N3646, N2081, N2392);
nor NOR3 (N12953, N12922, N7303, N11449);
nor NOR4 (N12954, N12952, N507, N7250, N12410);
xor XOR2 (N12955, N12945, N2709);
or OR3 (N12956, N12942, N9467, N12508);
or OR3 (N12957, N12943, N1048, N1209);
nand NAND4 (N12958, N12957, N9330, N7806, N8015);
not NOT1 (N12959, N12949);
buf BUF1 (N12960, N12953);
not NOT1 (N12961, N12938);
not NOT1 (N12962, N12955);
not NOT1 (N12963, N12950);
or OR3 (N12964, N12961, N9993, N4293);
not NOT1 (N12965, N12959);
nand NAND3 (N12966, N12965, N3961, N1756);
buf BUF1 (N12967, N12963);
and AND4 (N12968, N12967, N7196, N4617, N10357);
or OR4 (N12969, N12948, N6541, N12309, N3234);
buf BUF1 (N12970, N12966);
buf BUF1 (N12971, N12970);
nor NOR2 (N12972, N12971, N6819);
and AND2 (N12973, N12968, N9970);
not NOT1 (N12974, N12951);
nand NAND3 (N12975, N12964, N12602, N6156);
nor NOR2 (N12976, N12962, N1904);
or OR3 (N12977, N12969, N5426, N9402);
nand NAND3 (N12978, N12960, N6485, N6162);
nor NOR4 (N12979, N12958, N12349, N2548, N6541);
and AND4 (N12980, N12956, N5551, N8844, N2962);
nor NOR3 (N12981, N12975, N7316, N9051);
nor NOR4 (N12982, N12973, N3339, N7033, N8006);
not NOT1 (N12983, N12974);
and AND4 (N12984, N12979, N3540, N1647, N5542);
nand NAND2 (N12985, N12981, N12403);
not NOT1 (N12986, N12984);
buf BUF1 (N12987, N12977);
and AND3 (N12988, N12976, N3079, N10550);
xor XOR2 (N12989, N12972, N5031);
and AND3 (N12990, N12954, N8545, N149);
not NOT1 (N12991, N12987);
not NOT1 (N12992, N12990);
not NOT1 (N12993, N12992);
or OR3 (N12994, N12982, N5757, N11514);
xor XOR2 (N12995, N12988, N2818);
buf BUF1 (N12996, N12983);
buf BUF1 (N12997, N12985);
nand NAND4 (N12998, N12989, N9595, N11969, N1758);
nor NOR4 (N12999, N12986, N1831, N2860, N1530);
xor XOR2 (N13000, N12991, N10045);
xor XOR2 (N13001, N12994, N12918);
or OR4 (N13002, N12998, N10688, N354, N5613);
nor NOR2 (N13003, N12993, N12205);
nand NAND4 (N13004, N13003, N5371, N2677, N11265);
buf BUF1 (N13005, N12996);
not NOT1 (N13006, N13004);
nor NOR4 (N13007, N13006, N4544, N11096, N8101);
nor NOR3 (N13008, N13005, N7449, N192);
nor NOR3 (N13009, N13008, N1113, N10492);
nor NOR3 (N13010, N12995, N6367, N2673);
nor NOR2 (N13011, N12980, N10444);
xor XOR2 (N13012, N13011, N5477);
nand NAND4 (N13013, N13001, N11883, N11569, N4165);
not NOT1 (N13014, N13007);
nand NAND4 (N13015, N13013, N304, N1675, N7596);
nor NOR3 (N13016, N13002, N9553, N12626);
or OR3 (N13017, N13009, N7703, N2638);
nor NOR3 (N13018, N13016, N3633, N6974);
or OR3 (N13019, N13010, N4323, N1787);
not NOT1 (N13020, N13014);
nand NAND3 (N13021, N12999, N889, N3779);
buf BUF1 (N13022, N13020);
not NOT1 (N13023, N12978);
buf BUF1 (N13024, N12997);
and AND3 (N13025, N13000, N8753, N4248);
and AND4 (N13026, N13021, N11350, N1382, N2597);
or OR4 (N13027, N13025, N531, N11335, N7253);
or OR4 (N13028, N13012, N8795, N9688, N423);
or OR3 (N13029, N13023, N2390, N4525);
not NOT1 (N13030, N13017);
or OR2 (N13031, N13027, N6816);
not NOT1 (N13032, N13028);
and AND3 (N13033, N13022, N11087, N5479);
not NOT1 (N13034, N13030);
and AND4 (N13035, N13015, N4536, N9923, N2855);
nor NOR3 (N13036, N13024, N3854, N5966);
not NOT1 (N13037, N13032);
xor XOR2 (N13038, N13035, N5998);
and AND2 (N13039, N13038, N8854);
nor NOR3 (N13040, N13034, N11029, N28);
and AND2 (N13041, N13029, N1771);
and AND4 (N13042, N13026, N12463, N9063, N4569);
nor NOR4 (N13043, N13018, N6551, N6107, N10720);
or OR2 (N13044, N13040, N4946);
nor NOR2 (N13045, N13044, N5324);
not NOT1 (N13046, N13042);
or OR4 (N13047, N13039, N6485, N4470, N2100);
not NOT1 (N13048, N13036);
xor XOR2 (N13049, N13048, N2799);
nand NAND3 (N13050, N13031, N1198, N3241);
and AND3 (N13051, N13041, N8927, N10269);
buf BUF1 (N13052, N13050);
not NOT1 (N13053, N13045);
buf BUF1 (N13054, N13033);
buf BUF1 (N13055, N13053);
and AND2 (N13056, N13055, N5862);
not NOT1 (N13057, N13037);
xor XOR2 (N13058, N13052, N1665);
nor NOR3 (N13059, N13058, N8708, N8273);
or OR3 (N13060, N13051, N11312, N11578);
buf BUF1 (N13061, N13046);
and AND4 (N13062, N13054, N12051, N9275, N9515);
nor NOR2 (N13063, N13043, N2248);
nand NAND2 (N13064, N13061, N7758);
xor XOR2 (N13065, N13047, N11363);
or OR3 (N13066, N13019, N2286, N7723);
xor XOR2 (N13067, N13062, N7381);
or OR2 (N13068, N13049, N643);
nor NOR4 (N13069, N13056, N4195, N7141, N10079);
nand NAND4 (N13070, N13066, N10567, N4232, N3973);
or OR4 (N13071, N13069, N7931, N2413, N1109);
or OR4 (N13072, N13060, N12032, N10260, N2133);
nor NOR3 (N13073, N13059, N10545, N583);
xor XOR2 (N13074, N13073, N8538);
not NOT1 (N13075, N13070);
and AND2 (N13076, N13064, N2283);
not NOT1 (N13077, N13075);
xor XOR2 (N13078, N13063, N8944);
nor NOR2 (N13079, N13074, N1298);
xor XOR2 (N13080, N13076, N11825);
nor NOR3 (N13081, N13077, N9222, N4996);
nand NAND3 (N13082, N13065, N7212, N12162);
buf BUF1 (N13083, N13078);
and AND4 (N13084, N13068, N5114, N2402, N1299);
nor NOR3 (N13085, N13067, N2576, N785);
or OR4 (N13086, N13071, N3417, N12906, N9067);
not NOT1 (N13087, N13082);
buf BUF1 (N13088, N13086);
not NOT1 (N13089, N13081);
xor XOR2 (N13090, N13088, N2714);
nor NOR3 (N13091, N13085, N6728, N6707);
not NOT1 (N13092, N13089);
not NOT1 (N13093, N13090);
nor NOR3 (N13094, N13091, N2578, N7117);
not NOT1 (N13095, N13057);
buf BUF1 (N13096, N13083);
nand NAND4 (N13097, N13092, N8849, N12110, N10437);
buf BUF1 (N13098, N13079);
and AND2 (N13099, N13093, N2511);
buf BUF1 (N13100, N13098);
xor XOR2 (N13101, N13072, N9119);
and AND3 (N13102, N13101, N7110, N377);
xor XOR2 (N13103, N13096, N12991);
buf BUF1 (N13104, N13097);
not NOT1 (N13105, N13100);
buf BUF1 (N13106, N13080);
or OR3 (N13107, N13087, N10719, N12713);
not NOT1 (N13108, N13107);
or OR3 (N13109, N13104, N11232, N1162);
nand NAND4 (N13110, N13109, N6675, N1457, N12376);
and AND2 (N13111, N13103, N7571);
nand NAND2 (N13112, N13084, N10813);
nand NAND3 (N13113, N13106, N5245, N4650);
not NOT1 (N13114, N13105);
xor XOR2 (N13115, N13114, N10760);
and AND4 (N13116, N13113, N7713, N3632, N3939);
xor XOR2 (N13117, N13108, N12079);
xor XOR2 (N13118, N13094, N6385);
not NOT1 (N13119, N13112);
nand NAND4 (N13120, N13095, N8196, N10328, N1029);
buf BUF1 (N13121, N13119);
or OR3 (N13122, N13121, N8304, N12461);
nor NOR4 (N13123, N13111, N9031, N2820, N4357);
xor XOR2 (N13124, N13116, N1725);
or OR4 (N13125, N13117, N3377, N11305, N1288);
nor NOR3 (N13126, N13099, N571, N8144);
xor XOR2 (N13127, N13125, N10940);
xor XOR2 (N13128, N13110, N1894);
nand NAND3 (N13129, N13126, N7119, N5273);
xor XOR2 (N13130, N13118, N5007);
buf BUF1 (N13131, N13115);
nor NOR3 (N13132, N13127, N11883, N7491);
nand NAND3 (N13133, N13130, N9600, N5868);
nor NOR3 (N13134, N13124, N8883, N11422);
and AND4 (N13135, N13132, N1042, N10164, N3068);
nor NOR2 (N13136, N13129, N2619);
nand NAND2 (N13137, N13120, N10068);
and AND4 (N13138, N13137, N5308, N4607, N9947);
nor NOR2 (N13139, N13122, N9320);
not NOT1 (N13140, N13138);
nand NAND2 (N13141, N13135, N12359);
buf BUF1 (N13142, N13134);
or OR4 (N13143, N13140, N6072, N1031, N3601);
not NOT1 (N13144, N13141);
buf BUF1 (N13145, N13131);
xor XOR2 (N13146, N13144, N2543);
not NOT1 (N13147, N13143);
and AND2 (N13148, N13142, N5735);
xor XOR2 (N13149, N13133, N2734);
and AND3 (N13150, N13149, N759, N9392);
nor NOR3 (N13151, N13147, N11969, N6036);
or OR3 (N13152, N13148, N11284, N1705);
or OR4 (N13153, N13152, N447, N1706, N9922);
nand NAND3 (N13154, N13139, N11922, N10886);
or OR3 (N13155, N13136, N7264, N8474);
or OR4 (N13156, N13150, N2825, N1060, N1196);
not NOT1 (N13157, N13102);
xor XOR2 (N13158, N13155, N9789);
not NOT1 (N13159, N13151);
buf BUF1 (N13160, N13146);
and AND3 (N13161, N13157, N426, N10012);
buf BUF1 (N13162, N13159);
xor XOR2 (N13163, N13123, N11384);
xor XOR2 (N13164, N13128, N764);
and AND4 (N13165, N13154, N4295, N1074, N6006);
or OR4 (N13166, N13158, N4756, N7478, N647);
nand NAND4 (N13167, N13164, N4420, N2298, N5976);
and AND3 (N13168, N13160, N2489, N7358);
nand NAND4 (N13169, N13166, N8784, N7218, N7815);
or OR3 (N13170, N13165, N9619, N8846);
nand NAND2 (N13171, N13169, N1021);
buf BUF1 (N13172, N13171);
xor XOR2 (N13173, N13163, N9645);
not NOT1 (N13174, N13153);
not NOT1 (N13175, N13170);
or OR3 (N13176, N13172, N12358, N6491);
or OR4 (N13177, N13168, N4634, N8288, N2163);
or OR2 (N13178, N13145, N3971);
nand NAND2 (N13179, N13176, N634);
and AND2 (N13180, N13178, N3283);
nand NAND3 (N13181, N13167, N4687, N2263);
buf BUF1 (N13182, N13174);
xor XOR2 (N13183, N13179, N1581);
or OR4 (N13184, N13162, N13062, N9024, N4838);
buf BUF1 (N13185, N13180);
and AND4 (N13186, N13161, N12412, N3630, N5497);
buf BUF1 (N13187, N13182);
not NOT1 (N13188, N13184);
nor NOR3 (N13189, N13181, N5108, N11421);
xor XOR2 (N13190, N13156, N89);
nor NOR2 (N13191, N13183, N11534);
and AND3 (N13192, N13175, N8309, N12301);
buf BUF1 (N13193, N13190);
and AND3 (N13194, N13186, N7265, N4949);
not NOT1 (N13195, N13177);
xor XOR2 (N13196, N13189, N8206);
xor XOR2 (N13197, N13191, N5640);
buf BUF1 (N13198, N13192);
or OR2 (N13199, N13173, N6614);
xor XOR2 (N13200, N13193, N2697);
buf BUF1 (N13201, N13188);
nand NAND4 (N13202, N13185, N2331, N2582, N7971);
xor XOR2 (N13203, N13201, N7811);
and AND4 (N13204, N13194, N869, N9288, N863);
and AND3 (N13205, N13197, N9169, N8449);
not NOT1 (N13206, N13187);
and AND4 (N13207, N13200, N13114, N9581, N8330);
or OR2 (N13208, N13206, N7660);
and AND4 (N13209, N13205, N6946, N8304, N291);
nand NAND4 (N13210, N13198, N4527, N2400, N6736);
xor XOR2 (N13211, N13196, N4299);
buf BUF1 (N13212, N13210);
nand NAND2 (N13213, N13203, N8517);
or OR3 (N13214, N13202, N8805, N4726);
not NOT1 (N13215, N13204);
buf BUF1 (N13216, N13199);
nand NAND4 (N13217, N13211, N4410, N942, N2190);
or OR2 (N13218, N13213, N12073);
and AND3 (N13219, N13216, N8036, N6297);
buf BUF1 (N13220, N13219);
nor NOR4 (N13221, N13217, N9382, N12867, N9084);
nand NAND3 (N13222, N13208, N2581, N3053);
nor NOR4 (N13223, N13214, N1417, N9245, N6892);
not NOT1 (N13224, N13209);
not NOT1 (N13225, N13221);
buf BUF1 (N13226, N13195);
xor XOR2 (N13227, N13207, N7205);
nand NAND3 (N13228, N13226, N11471, N9708);
buf BUF1 (N13229, N13223);
nor NOR3 (N13230, N13220, N2055, N11132);
buf BUF1 (N13231, N13228);
nand NAND3 (N13232, N13225, N5218, N1856);
nand NAND3 (N13233, N13230, N7868, N7242);
or OR2 (N13234, N13227, N2604);
nor NOR3 (N13235, N13234, N4001, N1314);
nand NAND2 (N13236, N13232, N2136);
nand NAND2 (N13237, N13215, N11263);
nor NOR3 (N13238, N13212, N4263, N11669);
and AND3 (N13239, N13238, N5298, N3963);
buf BUF1 (N13240, N13239);
nor NOR3 (N13241, N13229, N165, N12874);
and AND4 (N13242, N13222, N7483, N1095, N10812);
nor NOR3 (N13243, N13241, N5337, N12727);
not NOT1 (N13244, N13224);
buf BUF1 (N13245, N13237);
nand NAND4 (N13246, N13242, N8981, N6083, N11802);
and AND2 (N13247, N13245, N2990);
buf BUF1 (N13248, N13236);
not NOT1 (N13249, N13231);
or OR4 (N13250, N13235, N5545, N12162, N499);
not NOT1 (N13251, N13248);
and AND3 (N13252, N13244, N6307, N5984);
not NOT1 (N13253, N13240);
and AND2 (N13254, N13252, N9088);
and AND3 (N13255, N13249, N8594, N9332);
and AND2 (N13256, N13246, N4008);
nor NOR2 (N13257, N13247, N2798);
buf BUF1 (N13258, N13257);
not NOT1 (N13259, N13251);
or OR3 (N13260, N13254, N5883, N6889);
nand NAND3 (N13261, N13218, N8172, N4290);
not NOT1 (N13262, N13253);
buf BUF1 (N13263, N13256);
nand NAND4 (N13264, N13260, N2653, N12618, N1194);
not NOT1 (N13265, N13250);
or OR3 (N13266, N13262, N5529, N11411);
nand NAND4 (N13267, N13258, N8783, N5538, N12214);
not NOT1 (N13268, N13261);
or OR2 (N13269, N13259, N4107);
not NOT1 (N13270, N13268);
nand NAND4 (N13271, N13266, N11154, N75, N9736);
buf BUF1 (N13272, N13267);
xor XOR2 (N13273, N13265, N7826);
not NOT1 (N13274, N13263);
and AND3 (N13275, N13271, N103, N3252);
or OR3 (N13276, N13255, N12530, N8471);
nor NOR3 (N13277, N13270, N12927, N11842);
nor NOR3 (N13278, N13276, N6846, N8440);
or OR4 (N13279, N13269, N12885, N2102, N8469);
not NOT1 (N13280, N13264);
not NOT1 (N13281, N13272);
or OR3 (N13282, N13278, N9445, N7854);
nor NOR2 (N13283, N13279, N8821);
not NOT1 (N13284, N13273);
not NOT1 (N13285, N13284);
xor XOR2 (N13286, N13281, N4772);
not NOT1 (N13287, N13243);
nor NOR2 (N13288, N13274, N11391);
xor XOR2 (N13289, N13282, N2822);
nand NAND4 (N13290, N13286, N6731, N8477, N800);
xor XOR2 (N13291, N13277, N3656);
or OR3 (N13292, N13275, N8598, N6167);
not NOT1 (N13293, N13285);
or OR4 (N13294, N13290, N6457, N12894, N4971);
xor XOR2 (N13295, N13294, N12915);
and AND4 (N13296, N13292, N1470, N5620, N66);
or OR4 (N13297, N13283, N9683, N6167, N7200);
nand NAND2 (N13298, N13297, N12753);
nor NOR4 (N13299, N13295, N5620, N7852, N12972);
or OR3 (N13300, N13289, N1220, N10408);
and AND2 (N13301, N13287, N11980);
xor XOR2 (N13302, N13280, N11693);
and AND2 (N13303, N13299, N2488);
xor XOR2 (N13304, N13301, N6454);
buf BUF1 (N13305, N13291);
nand NAND3 (N13306, N13298, N3539, N7895);
buf BUF1 (N13307, N13306);
nand NAND4 (N13308, N13304, N2765, N4133, N9177);
and AND3 (N13309, N13308, N2444, N3867);
nor NOR3 (N13310, N13293, N6765, N13181);
and AND2 (N13311, N13303, N3281);
nor NOR4 (N13312, N13233, N7672, N9415, N8199);
and AND3 (N13313, N13309, N7938, N677);
buf BUF1 (N13314, N13296);
buf BUF1 (N13315, N13312);
xor XOR2 (N13316, N13313, N3723);
or OR2 (N13317, N13311, N8251);
nor NOR3 (N13318, N13315, N6034, N544);
nor NOR4 (N13319, N13318, N7770, N5650, N5261);
xor XOR2 (N13320, N13317, N5503);
xor XOR2 (N13321, N13302, N1725);
nor NOR2 (N13322, N13288, N1374);
and AND2 (N13323, N13300, N2759);
buf BUF1 (N13324, N13322);
or OR4 (N13325, N13305, N1227, N9262, N8294);
not NOT1 (N13326, N13320);
nand NAND4 (N13327, N13307, N6620, N9109, N10544);
nand NAND2 (N13328, N13321, N10687);
not NOT1 (N13329, N13316);
and AND2 (N13330, N13327, N994);
not NOT1 (N13331, N13326);
or OR3 (N13332, N13331, N2947, N8519);
or OR2 (N13333, N13314, N1883);
xor XOR2 (N13334, N13323, N775);
nor NOR3 (N13335, N13330, N9642, N7628);
buf BUF1 (N13336, N13333);
and AND3 (N13337, N13328, N12099, N9538);
nand NAND4 (N13338, N13335, N5520, N11083, N8287);
or OR3 (N13339, N13329, N13078, N4815);
buf BUF1 (N13340, N13324);
nand NAND4 (N13341, N13337, N10116, N8049, N8116);
not NOT1 (N13342, N13334);
nand NAND3 (N13343, N13338, N3061, N10532);
or OR4 (N13344, N13310, N7990, N367, N2357);
or OR2 (N13345, N13319, N4485);
xor XOR2 (N13346, N13339, N4643);
nor NOR2 (N13347, N13332, N12874);
xor XOR2 (N13348, N13343, N4985);
not NOT1 (N13349, N13340);
and AND4 (N13350, N13348, N6775, N11789, N2931);
nand NAND2 (N13351, N13341, N4884);
and AND2 (N13352, N13325, N2994);
buf BUF1 (N13353, N13336);
or OR3 (N13354, N13353, N2285, N10514);
xor XOR2 (N13355, N13346, N7911);
or OR3 (N13356, N13344, N9031, N7410);
not NOT1 (N13357, N13352);
not NOT1 (N13358, N13349);
or OR3 (N13359, N13342, N4121, N6602);
buf BUF1 (N13360, N13347);
or OR4 (N13361, N13350, N51, N6447, N3013);
and AND2 (N13362, N13356, N9621);
and AND3 (N13363, N13351, N6192, N9758);
nand NAND4 (N13364, N13358, N11978, N13127, N7636);
nor NOR2 (N13365, N13359, N9982);
or OR2 (N13366, N13354, N5094);
or OR3 (N13367, N13345, N11363, N7094);
xor XOR2 (N13368, N13361, N9563);
and AND3 (N13369, N13362, N9731, N9562);
nor NOR3 (N13370, N13357, N9792, N2676);
not NOT1 (N13371, N13365);
not NOT1 (N13372, N13368);
or OR4 (N13373, N13364, N9181, N6266, N10412);
xor XOR2 (N13374, N13371, N9079);
and AND2 (N13375, N13374, N8307);
and AND3 (N13376, N13367, N5820, N3184);
or OR2 (N13377, N13373, N6208);
buf BUF1 (N13378, N13369);
nand NAND3 (N13379, N13360, N5239, N5721);
and AND2 (N13380, N13375, N2826);
not NOT1 (N13381, N13366);
xor XOR2 (N13382, N13376, N7767);
buf BUF1 (N13383, N13382);
buf BUF1 (N13384, N13372);
nand NAND4 (N13385, N13370, N624, N4389, N10989);
nor NOR4 (N13386, N13379, N5283, N11510, N502);
buf BUF1 (N13387, N13378);
buf BUF1 (N13388, N13355);
buf BUF1 (N13389, N13385);
or OR4 (N13390, N13386, N13063, N12927, N7101);
and AND3 (N13391, N13389, N8731, N9466);
nor NOR2 (N13392, N13390, N4442);
buf BUF1 (N13393, N13383);
buf BUF1 (N13394, N13381);
and AND2 (N13395, N13391, N3255);
not NOT1 (N13396, N13392);
xor XOR2 (N13397, N13394, N9961);
buf BUF1 (N13398, N13397);
or OR4 (N13399, N13393, N3287, N10183, N6696);
not NOT1 (N13400, N13363);
nand NAND4 (N13401, N13388, N4127, N7165, N4219);
nand NAND3 (N13402, N13399, N6046, N7532);
buf BUF1 (N13403, N13396);
xor XOR2 (N13404, N13380, N7147);
or OR4 (N13405, N13404, N7263, N11088, N4398);
buf BUF1 (N13406, N13405);
and AND3 (N13407, N13401, N11947, N2634);
nor NOR3 (N13408, N13398, N13243, N1330);
not NOT1 (N13409, N13384);
or OR2 (N13410, N13395, N719);
not NOT1 (N13411, N13403);
xor XOR2 (N13412, N13406, N3990);
buf BUF1 (N13413, N13402);
nor NOR2 (N13414, N13413, N5638);
nor NOR3 (N13415, N13387, N7825, N7216);
or OR4 (N13416, N13407, N8428, N11097, N7303);
not NOT1 (N13417, N13414);
xor XOR2 (N13418, N13415, N429);
nor NOR2 (N13419, N13409, N11977);
buf BUF1 (N13420, N13419);
buf BUF1 (N13421, N13411);
or OR3 (N13422, N13412, N341, N10655);
and AND2 (N13423, N13400, N11379);
buf BUF1 (N13424, N13410);
or OR4 (N13425, N13408, N5165, N11399, N491);
xor XOR2 (N13426, N13423, N9163);
or OR4 (N13427, N13416, N11849, N5441, N2836);
nor NOR4 (N13428, N13417, N10930, N10903, N4585);
not NOT1 (N13429, N13377);
nand NAND3 (N13430, N13425, N7902, N6671);
or OR2 (N13431, N13421, N143);
and AND2 (N13432, N13420, N11604);
or OR4 (N13433, N13431, N12368, N8425, N4829);
xor XOR2 (N13434, N13427, N2977);
xor XOR2 (N13435, N13429, N6092);
nor NOR4 (N13436, N13428, N12574, N7120, N6706);
and AND4 (N13437, N13435, N4805, N8111, N9917);
xor XOR2 (N13438, N13434, N10776);
nand NAND3 (N13439, N13426, N7041, N5292);
buf BUF1 (N13440, N13438);
and AND4 (N13441, N13432, N8187, N11745, N1686);
buf BUF1 (N13442, N13440);
or OR2 (N13443, N13436, N5331);
nand NAND2 (N13444, N13439, N3620);
or OR3 (N13445, N13444, N6040, N12473);
not NOT1 (N13446, N13433);
xor XOR2 (N13447, N13445, N11638);
buf BUF1 (N13448, N13437);
nor NOR3 (N13449, N13447, N7099, N2000);
nor NOR2 (N13450, N13446, N7693);
not NOT1 (N13451, N13441);
buf BUF1 (N13452, N13422);
nor NOR2 (N13453, N13449, N10618);
and AND4 (N13454, N13443, N4871, N2472, N8769);
or OR4 (N13455, N13442, N10717, N12746, N5880);
buf BUF1 (N13456, N13448);
or OR4 (N13457, N13452, N5319, N395, N8222);
nand NAND3 (N13458, N13424, N3909, N8976);
xor XOR2 (N13459, N13451, N3695);
buf BUF1 (N13460, N13454);
nor NOR2 (N13461, N13459, N274);
and AND3 (N13462, N13458, N9658, N10532);
not NOT1 (N13463, N13455);
or OR3 (N13464, N13418, N8471, N5696);
xor XOR2 (N13465, N13461, N9060);
and AND4 (N13466, N13463, N6952, N3521, N2826);
not NOT1 (N13467, N13460);
nor NOR2 (N13468, N13462, N6625);
buf BUF1 (N13469, N13468);
buf BUF1 (N13470, N13456);
and AND3 (N13471, N13466, N9647, N11904);
nor NOR2 (N13472, N13465, N1813);
buf BUF1 (N13473, N13469);
xor XOR2 (N13474, N13464, N1163);
not NOT1 (N13475, N13473);
not NOT1 (N13476, N13453);
buf BUF1 (N13477, N13476);
or OR4 (N13478, N13474, N10021, N8523, N11546);
nor NOR3 (N13479, N13472, N5964, N12421);
not NOT1 (N13480, N13477);
buf BUF1 (N13481, N13467);
nand NAND2 (N13482, N13470, N1615);
buf BUF1 (N13483, N13480);
and AND3 (N13484, N13479, N9602, N4121);
not NOT1 (N13485, N13482);
buf BUF1 (N13486, N13471);
nor NOR3 (N13487, N13475, N2708, N7171);
nand NAND4 (N13488, N13485, N11229, N10589, N10590);
or OR2 (N13489, N13486, N7968);
nand NAND3 (N13490, N13489, N356, N6471);
not NOT1 (N13491, N13484);
not NOT1 (N13492, N13478);
and AND4 (N13493, N13487, N3026, N4561, N7763);
nor NOR3 (N13494, N13430, N4800, N4751);
nand NAND4 (N13495, N13494, N5020, N8818, N3871);
xor XOR2 (N13496, N13481, N9967);
not NOT1 (N13497, N13483);
buf BUF1 (N13498, N13496);
not NOT1 (N13499, N13457);
nand NAND2 (N13500, N13495, N1828);
xor XOR2 (N13501, N13490, N12757);
nor NOR2 (N13502, N13488, N12697);
buf BUF1 (N13503, N13500);
and AND4 (N13504, N13497, N7934, N10637, N6748);
buf BUF1 (N13505, N13504);
xor XOR2 (N13506, N13499, N4114);
buf BUF1 (N13507, N13493);
not NOT1 (N13508, N13506);
not NOT1 (N13509, N13507);
and AND3 (N13510, N13503, N9459, N3525);
nand NAND4 (N13511, N13492, N9505, N10476, N8695);
buf BUF1 (N13512, N13450);
buf BUF1 (N13513, N13512);
nor NOR4 (N13514, N13509, N7610, N881, N707);
buf BUF1 (N13515, N13514);
xor XOR2 (N13516, N13513, N10034);
not NOT1 (N13517, N13508);
nand NAND2 (N13518, N13511, N11366);
or OR3 (N13519, N13501, N10671, N7215);
nand NAND4 (N13520, N13517, N6043, N12580, N9961);
nor NOR3 (N13521, N13510, N11226, N5224);
xor XOR2 (N13522, N13502, N7465);
buf BUF1 (N13523, N13515);
xor XOR2 (N13524, N13519, N4635);
and AND3 (N13525, N13523, N6688, N7884);
xor XOR2 (N13526, N13524, N2077);
or OR3 (N13527, N13526, N6697, N8756);
or OR2 (N13528, N13516, N13323);
not NOT1 (N13529, N13521);
nand NAND4 (N13530, N13525, N10551, N9445, N5669);
nor NOR4 (N13531, N13505, N11784, N5224, N9476);
or OR4 (N13532, N13531, N2257, N2976, N3681);
and AND2 (N13533, N13518, N3121);
buf BUF1 (N13534, N13529);
or OR3 (N13535, N13534, N11484, N13149);
not NOT1 (N13536, N13498);
buf BUF1 (N13537, N13527);
nor NOR4 (N13538, N13522, N13490, N11653, N8309);
nor NOR2 (N13539, N13528, N8107);
and AND3 (N13540, N13539, N1919, N5266);
nand NAND3 (N13541, N13520, N7563, N1834);
nand NAND4 (N13542, N13533, N11088, N6401, N3598);
or OR4 (N13543, N13537, N2073, N12166, N8026);
nor NOR4 (N13544, N13543, N10836, N5086, N11160);
not NOT1 (N13545, N13544);
not NOT1 (N13546, N13541);
xor XOR2 (N13547, N13530, N7899);
and AND2 (N13548, N13532, N5149);
not NOT1 (N13549, N13546);
buf BUF1 (N13550, N13548);
nand NAND4 (N13551, N13540, N11224, N5353, N420);
buf BUF1 (N13552, N13547);
or OR4 (N13553, N13550, N1954, N9393, N3423);
and AND4 (N13554, N13536, N8322, N12333, N778);
not NOT1 (N13555, N13552);
or OR4 (N13556, N13554, N6388, N9072, N10772);
nand NAND2 (N13557, N13549, N9623);
nor NOR3 (N13558, N13538, N8720, N9740);
not NOT1 (N13559, N13545);
xor XOR2 (N13560, N13542, N2926);
xor XOR2 (N13561, N13555, N3690);
or OR2 (N13562, N13558, N11409);
or OR3 (N13563, N13535, N7549, N5079);
nand NAND3 (N13564, N13561, N2046, N3711);
buf BUF1 (N13565, N13559);
xor XOR2 (N13566, N13491, N6584);
buf BUF1 (N13567, N13556);
nand NAND4 (N13568, N13553, N2490, N53, N8542);
nand NAND2 (N13569, N13563, N6768);
buf BUF1 (N13570, N13569);
xor XOR2 (N13571, N13562, N8847);
xor XOR2 (N13572, N13571, N13014);
xor XOR2 (N13573, N13570, N9261);
nor NOR2 (N13574, N13573, N6628);
or OR2 (N13575, N13551, N8148);
and AND3 (N13576, N13565, N1837, N11853);
nand NAND3 (N13577, N13575, N4114, N2499);
nor NOR4 (N13578, N13566, N1465, N7161, N3416);
nor NOR2 (N13579, N13567, N3194);
buf BUF1 (N13580, N13579);
not NOT1 (N13581, N13557);
xor XOR2 (N13582, N13564, N1180);
buf BUF1 (N13583, N13580);
and AND2 (N13584, N13572, N2106);
nor NOR4 (N13585, N13582, N768, N4870, N8542);
not NOT1 (N13586, N13584);
and AND4 (N13587, N13574, N5047, N5098, N6288);
buf BUF1 (N13588, N13587);
nand NAND4 (N13589, N13576, N11948, N5026, N5633);
or OR2 (N13590, N13560, N12184);
not NOT1 (N13591, N13588);
and AND3 (N13592, N13589, N7945, N13069);
nand NAND2 (N13593, N13581, N3398);
or OR4 (N13594, N13593, N5844, N12922, N7507);
nor NOR2 (N13595, N13578, N5196);
not NOT1 (N13596, N13577);
nor NOR3 (N13597, N13590, N4488, N9854);
nor NOR3 (N13598, N13595, N13147, N248);
xor XOR2 (N13599, N13592, N4341);
nor NOR3 (N13600, N13583, N7073, N2109);
xor XOR2 (N13601, N13599, N5930);
or OR2 (N13602, N13601, N1749);
xor XOR2 (N13603, N13568, N8805);
nor NOR2 (N13604, N13594, N1744);
nand NAND3 (N13605, N13597, N8539, N11711);
and AND3 (N13606, N13585, N6106, N5460);
and AND3 (N13607, N13606, N10460, N766);
not NOT1 (N13608, N13605);
and AND4 (N13609, N13598, N10579, N657, N13082);
not NOT1 (N13610, N13586);
nor NOR2 (N13611, N13604, N3134);
xor XOR2 (N13612, N13591, N5325);
nand NAND3 (N13613, N13612, N7099, N11931);
nor NOR3 (N13614, N13607, N12037, N11745);
nand NAND4 (N13615, N13608, N8190, N389, N5850);
not NOT1 (N13616, N13613);
buf BUF1 (N13617, N13602);
not NOT1 (N13618, N13611);
nand NAND2 (N13619, N13617, N7833);
nor NOR3 (N13620, N13603, N10491, N5638);
nor NOR2 (N13621, N13615, N6371);
not NOT1 (N13622, N13616);
nand NAND4 (N13623, N13610, N13106, N12053, N11055);
and AND2 (N13624, N13609, N6091);
xor XOR2 (N13625, N13622, N4406);
nor NOR2 (N13626, N13624, N12804);
buf BUF1 (N13627, N13620);
or OR2 (N13628, N13625, N5481);
and AND2 (N13629, N13623, N3035);
and AND3 (N13630, N13618, N12515, N3997);
xor XOR2 (N13631, N13626, N8490);
nand NAND3 (N13632, N13614, N2746, N2226);
nor NOR3 (N13633, N13631, N5180, N7061);
nor NOR3 (N13634, N13627, N12213, N5064);
buf BUF1 (N13635, N13596);
buf BUF1 (N13636, N13628);
not NOT1 (N13637, N13621);
and AND2 (N13638, N13633, N1084);
xor XOR2 (N13639, N13632, N2717);
buf BUF1 (N13640, N13619);
not NOT1 (N13641, N13635);
or OR2 (N13642, N13637, N5744);
or OR4 (N13643, N13629, N10309, N3734, N9407);
xor XOR2 (N13644, N13636, N11105);
nand NAND4 (N13645, N13641, N2206, N11091, N2505);
buf BUF1 (N13646, N13644);
not NOT1 (N13647, N13638);
buf BUF1 (N13648, N13645);
buf BUF1 (N13649, N13642);
nor NOR4 (N13650, N13630, N6002, N991, N3957);
nand NAND3 (N13651, N13600, N9374, N89);
nand NAND3 (N13652, N13639, N8171, N5219);
xor XOR2 (N13653, N13649, N5484);
buf BUF1 (N13654, N13648);
nand NAND2 (N13655, N13647, N10566);
nor NOR4 (N13656, N13643, N4555, N3952, N7531);
buf BUF1 (N13657, N13650);
buf BUF1 (N13658, N13640);
buf BUF1 (N13659, N13651);
nor NOR3 (N13660, N13656, N7894, N4178);
nor NOR3 (N13661, N13660, N6816, N12861);
xor XOR2 (N13662, N13659, N8063);
not NOT1 (N13663, N13653);
nand NAND4 (N13664, N13662, N6403, N8332, N2790);
xor XOR2 (N13665, N13658, N1620);
nor NOR4 (N13666, N13655, N12684, N6423, N13069);
not NOT1 (N13667, N13646);
and AND4 (N13668, N13657, N5389, N8528, N3576);
nand NAND3 (N13669, N13652, N2685, N1746);
xor XOR2 (N13670, N13665, N9619);
xor XOR2 (N13671, N13666, N7110);
not NOT1 (N13672, N13670);
nor NOR3 (N13673, N13634, N9684, N9712);
or OR3 (N13674, N13661, N455, N7048);
or OR2 (N13675, N13672, N2060);
buf BUF1 (N13676, N13669);
not NOT1 (N13677, N13668);
not NOT1 (N13678, N13671);
xor XOR2 (N13679, N13654, N2336);
xor XOR2 (N13680, N13676, N6447);
or OR4 (N13681, N13680, N10079, N8876, N7605);
or OR2 (N13682, N13679, N6707);
not NOT1 (N13683, N13664);
nor NOR3 (N13684, N13675, N9997, N707);
buf BUF1 (N13685, N13678);
nand NAND2 (N13686, N13673, N1639);
or OR2 (N13687, N13674, N10075);
or OR4 (N13688, N13667, N4886, N7683, N1103);
not NOT1 (N13689, N13677);
not NOT1 (N13690, N13684);
nand NAND2 (N13691, N13682, N10203);
and AND2 (N13692, N13681, N2357);
and AND2 (N13693, N13692, N557);
buf BUF1 (N13694, N13687);
nor NOR4 (N13695, N13663, N10071, N8491, N10746);
nor NOR2 (N13696, N13689, N4005);
buf BUF1 (N13697, N13695);
xor XOR2 (N13698, N13688, N13365);
or OR3 (N13699, N13690, N12837, N331);
nand NAND4 (N13700, N13698, N1569, N7258, N7768);
or OR2 (N13701, N13693, N8344);
nand NAND2 (N13702, N13683, N4269);
nand NAND3 (N13703, N13702, N11147, N1646);
xor XOR2 (N13704, N13701, N2877);
xor XOR2 (N13705, N13697, N2830);
nor NOR3 (N13706, N13704, N4855, N13471);
not NOT1 (N13707, N13694);
not NOT1 (N13708, N13706);
not NOT1 (N13709, N13708);
buf BUF1 (N13710, N13686);
or OR3 (N13711, N13691, N4463, N7094);
xor XOR2 (N13712, N13699, N2891);
not NOT1 (N13713, N13700);
nand NAND2 (N13714, N13707, N13440);
not NOT1 (N13715, N13696);
nor NOR4 (N13716, N13711, N13616, N9232, N1588);
buf BUF1 (N13717, N13715);
buf BUF1 (N13718, N13714);
and AND2 (N13719, N13713, N6367);
nand NAND4 (N13720, N13709, N7892, N8594, N5071);
not NOT1 (N13721, N13705);
xor XOR2 (N13722, N13720, N10569);
and AND3 (N13723, N13703, N5882, N9728);
nand NAND3 (N13724, N13717, N7702, N4802);
xor XOR2 (N13725, N13723, N5676);
or OR4 (N13726, N13718, N12132, N12974, N13324);
xor XOR2 (N13727, N13710, N1992);
nor NOR2 (N13728, N13712, N10326);
buf BUF1 (N13729, N13724);
nor NOR4 (N13730, N13721, N1208, N13569, N13188);
not NOT1 (N13731, N13727);
nor NOR4 (N13732, N13685, N2821, N12794, N5617);
buf BUF1 (N13733, N13732);
buf BUF1 (N13734, N13730);
nor NOR2 (N13735, N13729, N291);
or OR4 (N13736, N13722, N7394, N12563, N1699);
buf BUF1 (N13737, N13731);
buf BUF1 (N13738, N13726);
nand NAND2 (N13739, N13728, N12689);
xor XOR2 (N13740, N13737, N7777);
and AND4 (N13741, N13735, N8682, N10117, N3996);
nand NAND2 (N13742, N13739, N6715);
xor XOR2 (N13743, N13725, N7817);
not NOT1 (N13744, N13733);
nand NAND4 (N13745, N13719, N344, N8012, N5556);
buf BUF1 (N13746, N13743);
nand NAND3 (N13747, N13740, N3779, N2589);
not NOT1 (N13748, N13745);
and AND3 (N13749, N13747, N6150, N11553);
not NOT1 (N13750, N13716);
nor NOR4 (N13751, N13734, N10006, N2701, N2105);
nor NOR2 (N13752, N13736, N883);
buf BUF1 (N13753, N13746);
buf BUF1 (N13754, N13752);
nand NAND3 (N13755, N13750, N8892, N6918);
or OR2 (N13756, N13755, N1453);
buf BUF1 (N13757, N13756);
nor NOR3 (N13758, N13744, N12999, N6648);
and AND2 (N13759, N13741, N11918);
or OR3 (N13760, N13757, N8173, N9030);
nor NOR4 (N13761, N13758, N1573, N8569, N9147);
nor NOR4 (N13762, N13749, N4970, N10298, N1585);
or OR4 (N13763, N13753, N6573, N11936, N4052);
nor NOR4 (N13764, N13754, N10842, N8381, N504);
not NOT1 (N13765, N13751);
or OR2 (N13766, N13764, N1338);
buf BUF1 (N13767, N13761);
or OR4 (N13768, N13762, N5862, N2597, N7712);
buf BUF1 (N13769, N13760);
or OR4 (N13770, N13769, N12973, N424, N12413);
not NOT1 (N13771, N13763);
not NOT1 (N13772, N13771);
nand NAND4 (N13773, N13759, N4653, N3387, N2013);
xor XOR2 (N13774, N13766, N3645);
or OR3 (N13775, N13738, N12875, N12119);
not NOT1 (N13776, N13765);
and AND2 (N13777, N13768, N4024);
not NOT1 (N13778, N13748);
or OR3 (N13779, N13775, N8383, N11406);
nand NAND2 (N13780, N13767, N4586);
nor NOR3 (N13781, N13776, N11415, N2484);
nor NOR3 (N13782, N13774, N13081, N7430);
xor XOR2 (N13783, N13778, N12574);
and AND2 (N13784, N13772, N2504);
xor XOR2 (N13785, N13784, N11295);
nor NOR3 (N13786, N13770, N8608, N37);
and AND3 (N13787, N13779, N11609, N10353);
nor NOR4 (N13788, N13742, N9677, N3775, N9829);
nand NAND4 (N13789, N13781, N12032, N9221, N7028);
buf BUF1 (N13790, N13785);
or OR4 (N13791, N13777, N13285, N5132, N9918);
buf BUF1 (N13792, N13783);
nand NAND2 (N13793, N13782, N6102);
xor XOR2 (N13794, N13788, N3532);
nand NAND3 (N13795, N13786, N2171, N12561);
not NOT1 (N13796, N13792);
not NOT1 (N13797, N13795);
buf BUF1 (N13798, N13791);
xor XOR2 (N13799, N13780, N7261);
buf BUF1 (N13800, N13789);
nor NOR2 (N13801, N13796, N13311);
xor XOR2 (N13802, N13801, N1700);
and AND2 (N13803, N13800, N9853);
or OR2 (N13804, N13794, N10019);
not NOT1 (N13805, N13804);
nand NAND3 (N13806, N13799, N234, N2616);
and AND4 (N13807, N13793, N9496, N2884, N4933);
nand NAND2 (N13808, N13803, N9437);
not NOT1 (N13809, N13787);
nor NOR4 (N13810, N13808, N13568, N6101, N4650);
or OR2 (N13811, N13805, N5348);
and AND3 (N13812, N13806, N9318, N7586);
buf BUF1 (N13813, N13802);
and AND2 (N13814, N13813, N4817);
not NOT1 (N13815, N13811);
buf BUF1 (N13816, N13815);
xor XOR2 (N13817, N13809, N9601);
not NOT1 (N13818, N13773);
not NOT1 (N13819, N13818);
and AND4 (N13820, N13807, N918, N12410, N6391);
and AND4 (N13821, N13817, N9506, N4787, N3476);
xor XOR2 (N13822, N13797, N9630);
nand NAND2 (N13823, N13814, N13282);
and AND4 (N13824, N13810, N8413, N2893, N12997);
or OR4 (N13825, N13824, N13038, N2629, N3798);
not NOT1 (N13826, N13825);
or OR4 (N13827, N13790, N8256, N10774, N738);
nor NOR3 (N13828, N13827, N5630, N9743);
xor XOR2 (N13829, N13816, N7914);
xor XOR2 (N13830, N13829, N5979);
buf BUF1 (N13831, N13826);
buf BUF1 (N13832, N13828);
not NOT1 (N13833, N13820);
nor NOR3 (N13834, N13822, N6037, N5499);
not NOT1 (N13835, N13823);
not NOT1 (N13836, N13832);
buf BUF1 (N13837, N13830);
or OR3 (N13838, N13819, N3183, N13346);
or OR2 (N13839, N13831, N6082);
buf BUF1 (N13840, N13812);
or OR2 (N13841, N13798, N9236);
nor NOR2 (N13842, N13840, N352);
buf BUF1 (N13843, N13821);
not NOT1 (N13844, N13837);
not NOT1 (N13845, N13841);
xor XOR2 (N13846, N13844, N1624);
and AND4 (N13847, N13833, N10078, N7459, N5548);
and AND4 (N13848, N13836, N2885, N5333, N12333);
buf BUF1 (N13849, N13845);
or OR4 (N13850, N13848, N9462, N12606, N4823);
not NOT1 (N13851, N13849);
nand NAND3 (N13852, N13847, N10606, N3591);
not NOT1 (N13853, N13843);
buf BUF1 (N13854, N13851);
nor NOR3 (N13855, N13834, N12190, N3714);
nor NOR3 (N13856, N13852, N11119, N284);
or OR3 (N13857, N13856, N5081, N6922);
not NOT1 (N13858, N13838);
not NOT1 (N13859, N13853);
nand NAND3 (N13860, N13835, N7504, N6501);
buf BUF1 (N13861, N13854);
nor NOR3 (N13862, N13839, N8501, N6123);
buf BUF1 (N13863, N13842);
buf BUF1 (N13864, N13859);
or OR3 (N13865, N13846, N9086, N866);
or OR3 (N13866, N13865, N3819, N7665);
nand NAND3 (N13867, N13858, N3163, N9098);
not NOT1 (N13868, N13862);
or OR3 (N13869, N13861, N2103, N6901);
and AND2 (N13870, N13850, N2866);
xor XOR2 (N13871, N13870, N4328);
nor NOR4 (N13872, N13863, N8886, N12367, N9788);
nand NAND3 (N13873, N13872, N6721, N551);
or OR3 (N13874, N13857, N10856, N3278);
or OR3 (N13875, N13855, N2881, N7542);
or OR4 (N13876, N13875, N13638, N4371, N1955);
xor XOR2 (N13877, N13860, N11050);
and AND2 (N13878, N13868, N3233);
not NOT1 (N13879, N13877);
and AND2 (N13880, N13874, N3975);
xor XOR2 (N13881, N13879, N5763);
or OR3 (N13882, N13867, N4433, N1288);
nand NAND4 (N13883, N13878, N3184, N6563, N9275);
nand NAND3 (N13884, N13873, N2698, N2582);
or OR4 (N13885, N13880, N445, N2245, N2216);
nor NOR3 (N13886, N13871, N3823, N12508);
xor XOR2 (N13887, N13882, N13673);
nand NAND3 (N13888, N13885, N6564, N9044);
nor NOR2 (N13889, N13869, N425);
or OR4 (N13890, N13884, N5496, N12706, N13165);
buf BUF1 (N13891, N13866);
nand NAND4 (N13892, N13881, N7504, N1186, N3591);
xor XOR2 (N13893, N13888, N3304);
nor NOR2 (N13894, N13886, N8729);
nor NOR3 (N13895, N13893, N9532, N5782);
or OR3 (N13896, N13876, N10220, N12229);
buf BUF1 (N13897, N13887);
and AND2 (N13898, N13897, N11220);
and AND3 (N13899, N13883, N1759, N3720);
nor NOR2 (N13900, N13890, N11490);
xor XOR2 (N13901, N13898, N12010);
or OR4 (N13902, N13899, N4468, N11590, N6265);
or OR2 (N13903, N13894, N13791);
nand NAND2 (N13904, N13902, N3595);
nor NOR2 (N13905, N13900, N860);
xor XOR2 (N13906, N13904, N3643);
or OR3 (N13907, N13901, N5461, N6607);
nand NAND4 (N13908, N13896, N6936, N5536, N99);
nor NOR3 (N13909, N13907, N10921, N1094);
nor NOR4 (N13910, N13906, N6049, N13527, N795);
buf BUF1 (N13911, N13892);
or OR3 (N13912, N13908, N5928, N5261);
not NOT1 (N13913, N13905);
nor NOR4 (N13914, N13895, N11983, N7423, N9317);
nand NAND3 (N13915, N13911, N4534, N4998);
nand NAND4 (N13916, N13912, N4107, N1645, N5873);
nor NOR4 (N13917, N13889, N12955, N7104, N12915);
and AND3 (N13918, N13917, N3929, N7962);
nor NOR3 (N13919, N13914, N131, N13859);
nor NOR2 (N13920, N13891, N4927);
nand NAND4 (N13921, N13920, N3143, N9263, N3311);
or OR4 (N13922, N13916, N529, N4175, N13185);
nor NOR3 (N13923, N13918, N2003, N13226);
nor NOR2 (N13924, N13919, N10479);
not NOT1 (N13925, N13923);
buf BUF1 (N13926, N13915);
nor NOR3 (N13927, N13913, N9996, N5807);
buf BUF1 (N13928, N13924);
or OR4 (N13929, N13864, N5646, N5539, N371);
or OR2 (N13930, N13921, N11115);
not NOT1 (N13931, N13903);
buf BUF1 (N13932, N13928);
xor XOR2 (N13933, N13926, N3298);
not NOT1 (N13934, N13910);
buf BUF1 (N13935, N13932);
nor NOR4 (N13936, N13925, N6159, N1737, N4652);
xor XOR2 (N13937, N13933, N9914);
or OR3 (N13938, N13936, N7759, N12012);
buf BUF1 (N13939, N13935);
and AND4 (N13940, N13909, N12806, N12368, N5194);
or OR4 (N13941, N13938, N8813, N5379, N2938);
buf BUF1 (N13942, N13931);
and AND4 (N13943, N13934, N1154, N11280, N12877);
and AND3 (N13944, N13941, N8286, N9381);
not NOT1 (N13945, N13929);
and AND2 (N13946, N13939, N2324);
nor NOR2 (N13947, N13940, N5073);
xor XOR2 (N13948, N13942, N7536);
not NOT1 (N13949, N13927);
nand NAND3 (N13950, N13943, N1451, N10684);
or OR2 (N13951, N13950, N11075);
nand NAND3 (N13952, N13949, N3146, N3343);
nand NAND3 (N13953, N13947, N13886, N4044);
not NOT1 (N13954, N13937);
buf BUF1 (N13955, N13922);
xor XOR2 (N13956, N13948, N12408);
or OR4 (N13957, N13944, N3996, N1799, N9940);
nand NAND2 (N13958, N13952, N3390);
not NOT1 (N13959, N13956);
not NOT1 (N13960, N13958);
nand NAND3 (N13961, N13930, N184, N9636);
or OR4 (N13962, N13954, N12312, N7071, N2934);
buf BUF1 (N13963, N13959);
or OR3 (N13964, N13951, N6220, N4308);
or OR4 (N13965, N13962, N3109, N13932, N9162);
nor NOR4 (N13966, N13953, N2100, N13881, N9993);
buf BUF1 (N13967, N13945);
or OR4 (N13968, N13963, N6808, N1618, N13147);
not NOT1 (N13969, N13967);
buf BUF1 (N13970, N13964);
or OR4 (N13971, N13955, N11129, N8483, N8595);
buf BUF1 (N13972, N13971);
or OR4 (N13973, N13966, N10194, N9494, N13552);
xor XOR2 (N13974, N13972, N5925);
not NOT1 (N13975, N13946);
and AND4 (N13976, N13968, N877, N1981, N10551);
and AND2 (N13977, N13969, N3938);
or OR4 (N13978, N13975, N12265, N12048, N5617);
not NOT1 (N13979, N13961);
nand NAND4 (N13980, N13974, N406, N22, N7101);
or OR3 (N13981, N13970, N5991, N1087);
not NOT1 (N13982, N13973);
nand NAND3 (N13983, N13965, N2834, N958);
nor NOR3 (N13984, N13983, N11999, N1597);
nor NOR4 (N13985, N13979, N13768, N13476, N8494);
not NOT1 (N13986, N13985);
buf BUF1 (N13987, N13981);
nand NAND2 (N13988, N13977, N10818);
nor NOR3 (N13989, N13957, N4009, N6343);
and AND3 (N13990, N13989, N8838, N9941);
not NOT1 (N13991, N13987);
nor NOR2 (N13992, N13980, N2006);
xor XOR2 (N13993, N13982, N3771);
not NOT1 (N13994, N13992);
xor XOR2 (N13995, N13960, N10445);
not NOT1 (N13996, N13986);
or OR3 (N13997, N13984, N2651, N7126);
nand NAND3 (N13998, N13988, N6644, N3503);
nor NOR2 (N13999, N13994, N8751);
or OR4 (N14000, N13997, N13724, N1012, N11608);
buf BUF1 (N14001, N13991);
nand NAND4 (N14002, N13998, N1917, N5618, N13702);
nand NAND2 (N14003, N14001, N8141);
or OR4 (N14004, N13976, N3369, N5167, N2911);
nor NOR3 (N14005, N13990, N13706, N4058);
xor XOR2 (N14006, N13993, N11204);
nand NAND3 (N14007, N14004, N9037, N2532);
nand NAND4 (N14008, N13996, N1084, N9137, N13155);
xor XOR2 (N14009, N14000, N8577);
and AND4 (N14010, N13995, N13416, N7075, N12477);
not NOT1 (N14011, N13978);
and AND2 (N14012, N14002, N3703);
nand NAND4 (N14013, N14003, N838, N4296, N9319);
and AND2 (N14014, N13999, N8436);
nor NOR3 (N14015, N14014, N11102, N325);
not NOT1 (N14016, N14008);
buf BUF1 (N14017, N14010);
not NOT1 (N14018, N14012);
and AND4 (N14019, N14013, N6920, N13878, N8161);
and AND2 (N14020, N14011, N3831);
xor XOR2 (N14021, N14007, N2269);
nand NAND3 (N14022, N14018, N13956, N12123);
xor XOR2 (N14023, N14016, N5194);
nand NAND4 (N14024, N14020, N6945, N9449, N4561);
not NOT1 (N14025, N14019);
nand NAND3 (N14026, N14017, N10101, N4101);
buf BUF1 (N14027, N14025);
nor NOR4 (N14028, N14021, N9517, N4598, N11126);
xor XOR2 (N14029, N14027, N13623);
nor NOR4 (N14030, N14006, N3395, N245, N539);
or OR3 (N14031, N14024, N8921, N3658);
nand NAND4 (N14032, N14009, N9699, N9769, N12685);
buf BUF1 (N14033, N14022);
not NOT1 (N14034, N14005);
nor NOR3 (N14035, N14026, N8207, N11382);
buf BUF1 (N14036, N14031);
not NOT1 (N14037, N14029);
xor XOR2 (N14038, N14032, N1770);
buf BUF1 (N14039, N14030);
or OR4 (N14040, N14038, N4044, N3973, N13212);
buf BUF1 (N14041, N14034);
xor XOR2 (N14042, N14035, N4320);
or OR3 (N14043, N14015, N12300, N5950);
or OR3 (N14044, N14039, N9625, N12289);
or OR2 (N14045, N14028, N7559);
buf BUF1 (N14046, N14041);
and AND3 (N14047, N14045, N12282, N3204);
not NOT1 (N14048, N14043);
not NOT1 (N14049, N14040);
nor NOR4 (N14050, N14046, N6484, N55, N13742);
and AND4 (N14051, N14050, N2505, N4130, N2411);
buf BUF1 (N14052, N14044);
buf BUF1 (N14053, N14033);
or OR2 (N14054, N14053, N3927);
not NOT1 (N14055, N14052);
and AND4 (N14056, N14048, N10401, N3198, N9395);
nor NOR4 (N14057, N14042, N8533, N3587, N7063);
nor NOR3 (N14058, N14056, N13312, N4423);
xor XOR2 (N14059, N14058, N5699);
nor NOR3 (N14060, N14036, N11421, N3816);
not NOT1 (N14061, N14049);
buf BUF1 (N14062, N14037);
buf BUF1 (N14063, N14057);
and AND2 (N14064, N14023, N9057);
not NOT1 (N14065, N14060);
not NOT1 (N14066, N14054);
buf BUF1 (N14067, N14059);
nor NOR2 (N14068, N14047, N4835);
nor NOR4 (N14069, N14068, N8906, N9377, N1575);
not NOT1 (N14070, N14065);
nor NOR4 (N14071, N14063, N3016, N9669, N7577);
or OR4 (N14072, N14067, N10352, N5566, N13243);
nand NAND3 (N14073, N14072, N3995, N6303);
not NOT1 (N14074, N14055);
xor XOR2 (N14075, N14066, N3122);
buf BUF1 (N14076, N14075);
and AND2 (N14077, N14051, N6662);
or OR2 (N14078, N14064, N8598);
not NOT1 (N14079, N14070);
nor NOR3 (N14080, N14071, N9991, N1316);
nor NOR2 (N14081, N14062, N4125);
and AND3 (N14082, N14078, N3160, N2376);
not NOT1 (N14083, N14081);
not NOT1 (N14084, N14061);
and AND4 (N14085, N14083, N7391, N2417, N8672);
nand NAND4 (N14086, N14082, N5451, N3577, N3201);
xor XOR2 (N14087, N14079, N10544);
nand NAND4 (N14088, N14074, N1878, N5611, N11198);
or OR4 (N14089, N14088, N5990, N3898, N5377);
nand NAND4 (N14090, N14076, N676, N8932, N1442);
nor NOR2 (N14091, N14089, N12313);
nor NOR3 (N14092, N14086, N2391, N12944);
and AND3 (N14093, N14087, N12094, N10417);
or OR3 (N14094, N14090, N13354, N8159);
xor XOR2 (N14095, N14091, N781);
xor XOR2 (N14096, N14077, N5123);
not NOT1 (N14097, N14096);
xor XOR2 (N14098, N14080, N13929);
nor NOR3 (N14099, N14092, N3115, N9266);
buf BUF1 (N14100, N14073);
and AND2 (N14101, N14069, N3548);
buf BUF1 (N14102, N14095);
nor NOR3 (N14103, N14085, N1772, N7414);
buf BUF1 (N14104, N14097);
or OR2 (N14105, N14100, N5259);
and AND4 (N14106, N14102, N10114, N4122, N6571);
xor XOR2 (N14107, N14101, N1899);
buf BUF1 (N14108, N14094);
xor XOR2 (N14109, N14099, N2335);
xor XOR2 (N14110, N14103, N12143);
buf BUF1 (N14111, N14106);
or OR2 (N14112, N14084, N8849);
nor NOR4 (N14113, N14098, N8092, N623, N8034);
nand NAND4 (N14114, N14105, N13889, N2558, N13102);
and AND4 (N14115, N14112, N4622, N792, N4523);
nor NOR4 (N14116, N14113, N3768, N4493, N2049);
nand NAND4 (N14117, N14116, N10802, N2778, N11500);
not NOT1 (N14118, N14114);
nand NAND2 (N14119, N14118, N11325);
or OR3 (N14120, N14109, N7833, N1767);
and AND2 (N14121, N14110, N3766);
or OR4 (N14122, N14093, N1046, N4471, N1224);
not NOT1 (N14123, N14111);
nand NAND4 (N14124, N14119, N9189, N2333, N2311);
xor XOR2 (N14125, N14115, N5892);
xor XOR2 (N14126, N14124, N11249);
nand NAND3 (N14127, N14107, N790, N10733);
or OR2 (N14128, N14122, N3422);
nor NOR4 (N14129, N14123, N6899, N13900, N1968);
nand NAND2 (N14130, N14125, N13275);
or OR2 (N14131, N14108, N11063);
or OR3 (N14132, N14130, N4126, N2380);
not NOT1 (N14133, N14132);
nand NAND3 (N14134, N14131, N9839, N9142);
xor XOR2 (N14135, N14117, N3459);
buf BUF1 (N14136, N14133);
buf BUF1 (N14137, N14136);
nor NOR3 (N14138, N14120, N12480, N8010);
nand NAND2 (N14139, N14126, N12413);
nor NOR4 (N14140, N14104, N2593, N344, N10608);
buf BUF1 (N14141, N14121);
and AND4 (N14142, N14135, N9715, N8139, N1989);
nor NOR2 (N14143, N14128, N4594);
xor XOR2 (N14144, N14143, N2636);
nor NOR3 (N14145, N14137, N5256, N7255);
nand NAND2 (N14146, N14141, N7848);
xor XOR2 (N14147, N14134, N9679);
buf BUF1 (N14148, N14140);
nand NAND2 (N14149, N14145, N1588);
or OR4 (N14150, N14147, N5387, N8291, N7209);
xor XOR2 (N14151, N14138, N6326);
nor NOR4 (N14152, N14144, N9364, N2609, N5540);
xor XOR2 (N14153, N14152, N8498);
or OR3 (N14154, N14149, N9366, N232);
nor NOR2 (N14155, N14148, N9487);
and AND4 (N14156, N14127, N3965, N26, N6808);
nand NAND3 (N14157, N14146, N4411, N5766);
nor NOR4 (N14158, N14153, N5885, N9460, N6600);
xor XOR2 (N14159, N14154, N14106);
nand NAND4 (N14160, N14142, N12893, N2646, N3999);
and AND2 (N14161, N14156, N10296);
and AND2 (N14162, N14159, N8458);
buf BUF1 (N14163, N14129);
and AND2 (N14164, N14161, N10747);
xor XOR2 (N14165, N14157, N12159);
xor XOR2 (N14166, N14158, N11810);
not NOT1 (N14167, N14160);
nand NAND4 (N14168, N14151, N4892, N3454, N11244);
or OR3 (N14169, N14168, N11481, N4393);
or OR4 (N14170, N14162, N3292, N11329, N6588);
xor XOR2 (N14171, N14150, N7577);
nor NOR2 (N14172, N14169, N1053);
buf BUF1 (N14173, N14165);
and AND2 (N14174, N14155, N384);
xor XOR2 (N14175, N14174, N7083);
not NOT1 (N14176, N14175);
nand NAND2 (N14177, N14173, N5904);
or OR3 (N14178, N14139, N5094, N1567);
nor NOR4 (N14179, N14166, N7449, N13975, N1894);
not NOT1 (N14180, N14178);
nor NOR3 (N14181, N14171, N542, N7976);
or OR4 (N14182, N14163, N9813, N10797, N9820);
or OR4 (N14183, N14167, N1841, N13819, N3282);
or OR2 (N14184, N14183, N13962);
xor XOR2 (N14185, N14181, N9109);
and AND2 (N14186, N14184, N4720);
buf BUF1 (N14187, N14164);
and AND3 (N14188, N14177, N7736, N9945);
or OR3 (N14189, N14187, N3025, N3227);
or OR4 (N14190, N14180, N3704, N13201, N5097);
not NOT1 (N14191, N14176);
and AND4 (N14192, N14182, N11120, N1694, N11976);
and AND3 (N14193, N14172, N7008, N3164);
nand NAND3 (N14194, N14191, N4503, N14192);
or OR2 (N14195, N10174, N181);
and AND2 (N14196, N14189, N9163);
nor NOR3 (N14197, N14190, N12956, N6531);
not NOT1 (N14198, N14196);
and AND3 (N14199, N14179, N8282, N2783);
buf BUF1 (N14200, N14195);
buf BUF1 (N14201, N14199);
not NOT1 (N14202, N14198);
nand NAND2 (N14203, N14186, N9014);
and AND2 (N14204, N14185, N13878);
not NOT1 (N14205, N14200);
buf BUF1 (N14206, N14201);
buf BUF1 (N14207, N14170);
buf BUF1 (N14208, N14206);
nor NOR3 (N14209, N14203, N9777, N8115);
xor XOR2 (N14210, N14188, N11357);
buf BUF1 (N14211, N14209);
nor NOR2 (N14212, N14194, N2479);
buf BUF1 (N14213, N14202);
or OR3 (N14214, N14197, N7976, N6496);
xor XOR2 (N14215, N14205, N8997);
buf BUF1 (N14216, N14212);
xor XOR2 (N14217, N14207, N11357);
or OR2 (N14218, N14208, N13969);
or OR3 (N14219, N14216, N2563, N8309);
and AND3 (N14220, N14210, N3353, N2917);
buf BUF1 (N14221, N14211);
and AND3 (N14222, N14220, N11666, N11725);
nor NOR2 (N14223, N14219, N853);
nand NAND4 (N14224, N14221, N12472, N14201, N6857);
and AND2 (N14225, N14213, N3289);
not NOT1 (N14226, N14225);
nand NAND2 (N14227, N14204, N8186);
xor XOR2 (N14228, N14215, N10282);
nand NAND4 (N14229, N14228, N14141, N10708, N14052);
nand NAND2 (N14230, N14223, N13672);
nor NOR2 (N14231, N14226, N5770);
xor XOR2 (N14232, N14224, N4340);
nand NAND3 (N14233, N14214, N10278, N11294);
nor NOR2 (N14234, N14222, N4690);
xor XOR2 (N14235, N14218, N8126);
nor NOR3 (N14236, N14235, N7282, N3954);
not NOT1 (N14237, N14193);
nor NOR4 (N14238, N14217, N8864, N3613, N4703);
buf BUF1 (N14239, N14227);
xor XOR2 (N14240, N14237, N7841);
nand NAND4 (N14241, N14240, N10756, N13577, N3391);
nor NOR2 (N14242, N14229, N1064);
xor XOR2 (N14243, N14238, N2148);
and AND2 (N14244, N14233, N11493);
buf BUF1 (N14245, N14243);
nor NOR2 (N14246, N14232, N8256);
and AND3 (N14247, N14244, N11830, N3180);
or OR3 (N14248, N14245, N2428, N7268);
or OR2 (N14249, N14236, N2602);
and AND4 (N14250, N14248, N7628, N10763, N10449);
buf BUF1 (N14251, N14234);
buf BUF1 (N14252, N14251);
or OR4 (N14253, N14249, N4404, N7165, N4032);
nor NOR3 (N14254, N14252, N7962, N6741);
nor NOR4 (N14255, N14246, N8361, N2858, N1109);
not NOT1 (N14256, N14247);
not NOT1 (N14257, N14255);
xor XOR2 (N14258, N14254, N13078);
nand NAND2 (N14259, N14250, N6432);
nor NOR4 (N14260, N14242, N2755, N4692, N6928);
and AND4 (N14261, N14230, N3552, N11971, N11251);
or OR2 (N14262, N14259, N11008);
nor NOR3 (N14263, N14256, N3916, N7686);
nor NOR2 (N14264, N14263, N14014);
nor NOR4 (N14265, N14264, N2673, N2929, N5859);
xor XOR2 (N14266, N14261, N682);
buf BUF1 (N14267, N14266);
nor NOR3 (N14268, N14258, N2716, N8824);
buf BUF1 (N14269, N14267);
not NOT1 (N14270, N14265);
xor XOR2 (N14271, N14241, N13190);
or OR2 (N14272, N14239, N4776);
and AND4 (N14273, N14271, N863, N14202, N2145);
and AND2 (N14274, N14231, N1747);
nand NAND2 (N14275, N14269, N7729);
nand NAND4 (N14276, N14270, N8473, N10013, N13261);
or OR3 (N14277, N14276, N14022, N10649);
or OR3 (N14278, N14275, N606, N14155);
nor NOR4 (N14279, N14272, N536, N1772, N9962);
nor NOR2 (N14280, N14260, N10534);
xor XOR2 (N14281, N14262, N11392);
and AND4 (N14282, N14278, N14062, N13789, N3718);
buf BUF1 (N14283, N14273);
or OR3 (N14284, N14281, N13181, N3157);
or OR4 (N14285, N14279, N11063, N5604, N14215);
buf BUF1 (N14286, N14280);
not NOT1 (N14287, N14286);
xor XOR2 (N14288, N14285, N5850);
xor XOR2 (N14289, N14288, N14225);
not NOT1 (N14290, N14287);
xor XOR2 (N14291, N14274, N481);
or OR4 (N14292, N14290, N7115, N10958, N8406);
nand NAND4 (N14293, N14268, N2668, N7892, N4000);
and AND4 (N14294, N14282, N518, N11980, N7350);
not NOT1 (N14295, N14291);
not NOT1 (N14296, N14277);
nand NAND2 (N14297, N14296, N13312);
buf BUF1 (N14298, N14293);
not NOT1 (N14299, N14284);
nand NAND2 (N14300, N14294, N12905);
xor XOR2 (N14301, N14300, N12144);
not NOT1 (N14302, N14292);
or OR3 (N14303, N14289, N7781, N6272);
or OR3 (N14304, N14257, N803, N7589);
and AND3 (N14305, N14298, N4112, N4182);
and AND3 (N14306, N14301, N6669, N11358);
nor NOR2 (N14307, N14306, N8308);
xor XOR2 (N14308, N14295, N12453);
or OR2 (N14309, N14307, N11554);
buf BUF1 (N14310, N14299);
xor XOR2 (N14311, N14309, N9869);
xor XOR2 (N14312, N14308, N13576);
buf BUF1 (N14313, N14312);
nor NOR2 (N14314, N14303, N1346);
and AND3 (N14315, N14297, N10986, N22);
not NOT1 (N14316, N14310);
and AND2 (N14317, N14304, N12260);
nor NOR3 (N14318, N14314, N14148, N5932);
or OR3 (N14319, N14315, N11938, N2064);
buf BUF1 (N14320, N14305);
not NOT1 (N14321, N14320);
xor XOR2 (N14322, N14318, N13684);
buf BUF1 (N14323, N14253);
nand NAND4 (N14324, N14313, N3521, N7470, N3716);
buf BUF1 (N14325, N14316);
nor NOR2 (N14326, N14317, N715);
xor XOR2 (N14327, N14326, N4215);
not NOT1 (N14328, N14302);
or OR3 (N14329, N14328, N9752, N12665);
nand NAND2 (N14330, N14325, N3697);
or OR3 (N14331, N14324, N11131, N3801);
nor NOR2 (N14332, N14322, N7552);
nor NOR2 (N14333, N14330, N2306);
nand NAND4 (N14334, N14331, N6901, N277, N1956);
or OR2 (N14335, N14333, N1917);
not NOT1 (N14336, N14283);
and AND3 (N14337, N14319, N1677, N9374);
buf BUF1 (N14338, N14327);
not NOT1 (N14339, N14338);
xor XOR2 (N14340, N14335, N12855);
not NOT1 (N14341, N14321);
buf BUF1 (N14342, N14336);
buf BUF1 (N14343, N14329);
nand NAND3 (N14344, N14339, N12857, N10676);
and AND3 (N14345, N14332, N4312, N13545);
nor NOR4 (N14346, N14337, N10107, N4979, N6241);
nand NAND2 (N14347, N14334, N6658);
not NOT1 (N14348, N14340);
buf BUF1 (N14349, N14323);
xor XOR2 (N14350, N14343, N10129);
or OR3 (N14351, N14349, N8677, N9482);
nor NOR2 (N14352, N14350, N6042);
buf BUF1 (N14353, N14348);
or OR2 (N14354, N14311, N13844);
nand NAND2 (N14355, N14342, N10250);
buf BUF1 (N14356, N14355);
xor XOR2 (N14357, N14347, N6799);
buf BUF1 (N14358, N14357);
nand NAND4 (N14359, N14345, N10259, N3151, N2746);
or OR4 (N14360, N14341, N1458, N14187, N9533);
nor NOR3 (N14361, N14354, N1861, N2781);
buf BUF1 (N14362, N14360);
xor XOR2 (N14363, N14359, N12739);
nor NOR2 (N14364, N14353, N6856);
nor NOR4 (N14365, N14361, N5880, N2507, N13398);
xor XOR2 (N14366, N14356, N7362);
and AND3 (N14367, N14363, N6665, N10918);
and AND4 (N14368, N14351, N12300, N9936, N12473);
xor XOR2 (N14369, N14352, N3532);
or OR4 (N14370, N14366, N195, N5605, N5873);
xor XOR2 (N14371, N14367, N74);
xor XOR2 (N14372, N14344, N12068);
or OR4 (N14373, N14368, N8288, N11165, N2377);
or OR2 (N14374, N14371, N5545);
or OR4 (N14375, N14374, N12993, N8599, N1506);
buf BUF1 (N14376, N14346);
buf BUF1 (N14377, N14375);
nor NOR2 (N14378, N14376, N13712);
not NOT1 (N14379, N14373);
and AND4 (N14380, N14379, N11915, N1947, N12);
buf BUF1 (N14381, N14378);
nand NAND3 (N14382, N14369, N9395, N9161);
xor XOR2 (N14383, N14365, N13088);
buf BUF1 (N14384, N14383);
or OR2 (N14385, N14381, N5800);
buf BUF1 (N14386, N14362);
nand NAND3 (N14387, N14382, N12446, N6094);
nand NAND3 (N14388, N14370, N10745, N2410);
xor XOR2 (N14389, N14372, N8208);
nand NAND4 (N14390, N14380, N560, N1028, N4850);
not NOT1 (N14391, N14389);
or OR2 (N14392, N14364, N8671);
buf BUF1 (N14393, N14384);
nand NAND2 (N14394, N14388, N13404);
xor XOR2 (N14395, N14391, N10574);
or OR4 (N14396, N14387, N59, N5391, N11697);
or OR2 (N14397, N14358, N10602);
nor NOR2 (N14398, N14377, N3280);
nand NAND4 (N14399, N14394, N8371, N6588, N308);
xor XOR2 (N14400, N14386, N7916);
not NOT1 (N14401, N14395);
nand NAND2 (N14402, N14399, N11539);
nand NAND2 (N14403, N14396, N3666);
buf BUF1 (N14404, N14397);
buf BUF1 (N14405, N14400);
or OR2 (N14406, N14385, N6762);
and AND4 (N14407, N14405, N9633, N456, N3800);
and AND3 (N14408, N14407, N11703, N14363);
or OR2 (N14409, N14401, N9900);
not NOT1 (N14410, N14406);
buf BUF1 (N14411, N14410);
or OR4 (N14412, N14411, N611, N9333, N6727);
or OR4 (N14413, N14409, N1197, N9036, N4644);
nor NOR3 (N14414, N14390, N4625, N5038);
xor XOR2 (N14415, N14403, N8);
nor NOR2 (N14416, N14392, N5401);
xor XOR2 (N14417, N14416, N1026);
or OR4 (N14418, N14412, N8133, N14194, N12352);
or OR4 (N14419, N14417, N8062, N12620, N12285);
buf BUF1 (N14420, N14398);
nand NAND2 (N14421, N14408, N7050);
nor NOR4 (N14422, N14404, N12145, N11288, N3833);
buf BUF1 (N14423, N14420);
not NOT1 (N14424, N14413);
nor NOR3 (N14425, N14415, N5582, N128);
xor XOR2 (N14426, N14418, N10122);
buf BUF1 (N14427, N14393);
buf BUF1 (N14428, N14422);
and AND3 (N14429, N14426, N5626, N4729);
buf BUF1 (N14430, N14428);
and AND3 (N14431, N14419, N5003, N4463);
not NOT1 (N14432, N14427);
and AND2 (N14433, N14431, N7608);
buf BUF1 (N14434, N14414);
nor NOR4 (N14435, N14434, N3266, N9225, N9330);
nand NAND4 (N14436, N14433, N3674, N11224, N10803);
and AND4 (N14437, N14435, N3065, N28, N12681);
not NOT1 (N14438, N14429);
nand NAND2 (N14439, N14436, N5994);
nand NAND3 (N14440, N14432, N6485, N13536);
nand NAND4 (N14441, N14421, N8461, N6848, N10443);
nor NOR2 (N14442, N14440, N2059);
nor NOR4 (N14443, N14438, N3538, N13685, N3974);
xor XOR2 (N14444, N14423, N6137);
not NOT1 (N14445, N14444);
or OR2 (N14446, N14443, N9745);
not NOT1 (N14447, N14442);
buf BUF1 (N14448, N14445);
nor NOR2 (N14449, N14448, N12229);
or OR2 (N14450, N14437, N12261);
and AND2 (N14451, N14439, N1566);
or OR2 (N14452, N14451, N1227);
or OR2 (N14453, N14449, N7570);
buf BUF1 (N14454, N14425);
xor XOR2 (N14455, N14447, N10629);
buf BUF1 (N14456, N14454);
nor NOR2 (N14457, N14456, N10601);
buf BUF1 (N14458, N14450);
xor XOR2 (N14459, N14441, N13057);
xor XOR2 (N14460, N14459, N13953);
or OR3 (N14461, N14455, N710, N8672);
and AND3 (N14462, N14453, N4307, N13833);
or OR3 (N14463, N14446, N8368, N13494);
nor NOR2 (N14464, N14462, N3910);
nand NAND2 (N14465, N14452, N12500);
not NOT1 (N14466, N14424);
nor NOR3 (N14467, N14466, N7897, N12409);
nand NAND4 (N14468, N14467, N13403, N6295, N5532);
and AND3 (N14469, N14402, N2318, N14425);
nand NAND3 (N14470, N14430, N10701, N13699);
or OR2 (N14471, N14461, N14064);
nand NAND3 (N14472, N14458, N11025, N8577);
xor XOR2 (N14473, N14465, N5405);
buf BUF1 (N14474, N14464);
nand NAND3 (N14475, N14463, N13402, N5258);
nor NOR4 (N14476, N14475, N8689, N12289, N25);
xor XOR2 (N14477, N14460, N3583);
xor XOR2 (N14478, N14473, N8263);
not NOT1 (N14479, N14477);
or OR3 (N14480, N14474, N4847, N8052);
nor NOR3 (N14481, N14469, N11049, N11756);
and AND2 (N14482, N14476, N9683);
or OR4 (N14483, N14470, N4923, N9200, N3191);
or OR3 (N14484, N14472, N10074, N893);
not NOT1 (N14485, N14479);
and AND4 (N14486, N14482, N5770, N8061, N4373);
buf BUF1 (N14487, N14468);
buf BUF1 (N14488, N14485);
buf BUF1 (N14489, N14471);
nor NOR3 (N14490, N14481, N4098, N4958);
or OR3 (N14491, N14457, N13381, N2943);
and AND2 (N14492, N14480, N10149);
nor NOR4 (N14493, N14478, N10655, N6401, N8159);
nor NOR4 (N14494, N14483, N4185, N9546, N4537);
buf BUF1 (N14495, N14487);
not NOT1 (N14496, N14494);
nor NOR2 (N14497, N14496, N9018);
or OR4 (N14498, N14489, N12419, N3388, N8923);
nor NOR3 (N14499, N14488, N12422, N9214);
or OR4 (N14500, N14499, N6705, N4651, N13192);
or OR3 (N14501, N14484, N9036, N11719);
xor XOR2 (N14502, N14493, N14248);
or OR2 (N14503, N14486, N8112);
nand NAND2 (N14504, N14503, N266);
xor XOR2 (N14505, N14500, N2744);
and AND3 (N14506, N14504, N7139, N5208);
xor XOR2 (N14507, N14495, N13471);
nand NAND4 (N14508, N14497, N2143, N6036, N9246);
nand NAND4 (N14509, N14490, N10682, N7892, N6301);
buf BUF1 (N14510, N14507);
and AND2 (N14511, N14509, N1589);
and AND3 (N14512, N14501, N3420, N9841);
xor XOR2 (N14513, N14512, N11056);
buf BUF1 (N14514, N14505);
or OR4 (N14515, N14492, N5523, N4746, N13632);
buf BUF1 (N14516, N14508);
xor XOR2 (N14517, N14498, N4385);
xor XOR2 (N14518, N14513, N2130);
xor XOR2 (N14519, N14491, N523);
nand NAND3 (N14520, N14517, N14069, N915);
nand NAND2 (N14521, N14520, N13030);
buf BUF1 (N14522, N14506);
or OR2 (N14523, N14511, N10361);
not NOT1 (N14524, N14519);
xor XOR2 (N14525, N14524, N11617);
and AND3 (N14526, N14515, N340, N5592);
or OR3 (N14527, N14518, N5785, N483);
buf BUF1 (N14528, N14510);
buf BUF1 (N14529, N14516);
xor XOR2 (N14530, N14529, N4985);
xor XOR2 (N14531, N14521, N7697);
nand NAND2 (N14532, N14525, N4914);
and AND3 (N14533, N14526, N13758, N8675);
and AND2 (N14534, N14531, N409);
buf BUF1 (N14535, N14522);
or OR2 (N14536, N14530, N8375);
or OR2 (N14537, N14502, N4746);
xor XOR2 (N14538, N14534, N2941);
or OR3 (N14539, N14535, N4823, N14531);
and AND2 (N14540, N14528, N3872);
and AND4 (N14541, N14533, N2534, N12899, N9445);
nor NOR3 (N14542, N14523, N9556, N6352);
nand NAND3 (N14543, N14537, N2391, N12923);
not NOT1 (N14544, N14532);
xor XOR2 (N14545, N14540, N304);
xor XOR2 (N14546, N14539, N4724);
or OR2 (N14547, N14542, N6676);
nor NOR3 (N14548, N14547, N98, N5025);
not NOT1 (N14549, N14545);
or OR4 (N14550, N14548, N7197, N13280, N386);
or OR2 (N14551, N14544, N13973);
nor NOR4 (N14552, N14541, N13864, N6117, N11956);
nand NAND3 (N14553, N14550, N11853, N1940);
not NOT1 (N14554, N14543);
nand NAND2 (N14555, N14536, N9779);
or OR2 (N14556, N14538, N6785);
nor NOR2 (N14557, N14514, N2426);
nor NOR2 (N14558, N14554, N12595);
or OR2 (N14559, N14558, N10533);
not NOT1 (N14560, N14557);
nor NOR4 (N14561, N14527, N12955, N5625, N6558);
or OR4 (N14562, N14546, N9419, N8193, N8117);
not NOT1 (N14563, N14562);
buf BUF1 (N14564, N14555);
nand NAND4 (N14565, N14564, N13219, N3186, N13438);
or OR2 (N14566, N14553, N711);
xor XOR2 (N14567, N14559, N12308);
and AND2 (N14568, N14549, N675);
not NOT1 (N14569, N14561);
nor NOR2 (N14570, N14563, N195);
not NOT1 (N14571, N14568);
nor NOR2 (N14572, N14560, N9226);
nor NOR4 (N14573, N14570, N223, N9241, N1862);
nand NAND3 (N14574, N14552, N12834, N12944);
buf BUF1 (N14575, N14556);
and AND3 (N14576, N14569, N4136, N6319);
buf BUF1 (N14577, N14572);
not NOT1 (N14578, N14566);
nand NAND2 (N14579, N14577, N5399);
or OR2 (N14580, N14565, N6360);
or OR4 (N14581, N14579, N6275, N7590, N6905);
not NOT1 (N14582, N14567);
buf BUF1 (N14583, N14573);
and AND2 (N14584, N14583, N11953);
not NOT1 (N14585, N14581);
or OR3 (N14586, N14576, N1834, N13736);
buf BUF1 (N14587, N14551);
not NOT1 (N14588, N14582);
buf BUF1 (N14589, N14578);
nand NAND2 (N14590, N14587, N1349);
buf BUF1 (N14591, N14571);
and AND4 (N14592, N14585, N10611, N1805, N5169);
or OR2 (N14593, N14588, N4747);
not NOT1 (N14594, N14574);
xor XOR2 (N14595, N14575, N1381);
or OR3 (N14596, N14592, N8052, N7422);
xor XOR2 (N14597, N14590, N14332);
not NOT1 (N14598, N14596);
nor NOR4 (N14599, N14598, N3215, N9638, N8437);
or OR3 (N14600, N14595, N3280, N11498);
xor XOR2 (N14601, N14599, N4332);
xor XOR2 (N14602, N14586, N8588);
not NOT1 (N14603, N14602);
or OR3 (N14604, N14580, N14112, N1600);
or OR4 (N14605, N14604, N2129, N5160, N10512);
nor NOR4 (N14606, N14605, N9098, N12868, N13658);
and AND4 (N14607, N14603, N3779, N5300, N14489);
not NOT1 (N14608, N14591);
or OR3 (N14609, N14589, N6188, N7534);
nand NAND3 (N14610, N14609, N5105, N7019);
or OR2 (N14611, N14606, N1082);
buf BUF1 (N14612, N14584);
buf BUF1 (N14613, N14611);
nand NAND4 (N14614, N14593, N1617, N5035, N13338);
xor XOR2 (N14615, N14597, N2956);
and AND3 (N14616, N14612, N1576, N12872);
buf BUF1 (N14617, N14616);
or OR2 (N14618, N14614, N2047);
nand NAND2 (N14619, N14613, N11877);
or OR3 (N14620, N14617, N2638, N12827);
or OR2 (N14621, N14594, N1899);
nand NAND3 (N14622, N14600, N11779, N2485);
nor NOR4 (N14623, N14618, N11175, N7006, N9920);
nor NOR4 (N14624, N14615, N1058, N8118, N4421);
nand NAND3 (N14625, N14624, N8957, N8708);
nor NOR2 (N14626, N14621, N14170);
nor NOR4 (N14627, N14623, N10515, N2675, N11098);
or OR3 (N14628, N14610, N3815, N11518);
nor NOR3 (N14629, N14620, N8635, N12321);
not NOT1 (N14630, N14607);
buf BUF1 (N14631, N14626);
nor NOR2 (N14632, N14601, N6102);
nand NAND3 (N14633, N14622, N9435, N9963);
xor XOR2 (N14634, N14631, N1915);
nand NAND4 (N14635, N14630, N9373, N6201, N7375);
xor XOR2 (N14636, N14625, N7688);
xor XOR2 (N14637, N14628, N14636);
and AND4 (N14638, N8102, N8491, N9921, N11166);
xor XOR2 (N14639, N14637, N6872);
and AND4 (N14640, N14608, N6651, N9420, N12370);
buf BUF1 (N14641, N14639);
nand NAND3 (N14642, N14627, N12384, N3905);
or OR3 (N14643, N14619, N13582, N3530);
buf BUF1 (N14644, N14629);
nand NAND2 (N14645, N14632, N11808);
and AND2 (N14646, N14635, N7619);
nor NOR4 (N14647, N14646, N9241, N8458, N421);
and AND2 (N14648, N14638, N4074);
nand NAND4 (N14649, N14642, N11659, N1223, N1053);
or OR4 (N14650, N14647, N9027, N3425, N14486);
buf BUF1 (N14651, N14640);
nand NAND4 (N14652, N14648, N11585, N10235, N6788);
not NOT1 (N14653, N14644);
buf BUF1 (N14654, N14645);
nor NOR4 (N14655, N14643, N10555, N4081, N12255);
nand NAND2 (N14656, N14652, N5772);
xor XOR2 (N14657, N14654, N7821);
nor NOR3 (N14658, N14649, N7256, N8519);
or OR3 (N14659, N14655, N12124, N5648);
not NOT1 (N14660, N14659);
nor NOR3 (N14661, N14657, N11898, N8324);
and AND3 (N14662, N14656, N11431, N956);
or OR3 (N14663, N14658, N11678, N7956);
buf BUF1 (N14664, N14661);
xor XOR2 (N14665, N14633, N13606);
xor XOR2 (N14666, N14663, N9002);
nand NAND3 (N14667, N14650, N178, N13616);
not NOT1 (N14668, N14641);
or OR4 (N14669, N14667, N14533, N13453, N9282);
nor NOR4 (N14670, N14660, N8378, N5197, N5234);
buf BUF1 (N14671, N14665);
nand NAND2 (N14672, N14651, N11842);
nor NOR3 (N14673, N14672, N8181, N14595);
not NOT1 (N14674, N14668);
and AND4 (N14675, N14671, N12049, N6664, N12943);
nor NOR2 (N14676, N14664, N1139);
and AND4 (N14677, N14666, N3967, N13029, N5058);
xor XOR2 (N14678, N14634, N6020);
nor NOR4 (N14679, N14678, N6758, N7787, N5698);
xor XOR2 (N14680, N14677, N11982);
not NOT1 (N14681, N14662);
and AND4 (N14682, N14669, N14413, N2683, N10635);
not NOT1 (N14683, N14676);
xor XOR2 (N14684, N14682, N13437);
nor NOR3 (N14685, N14681, N9775, N6085);
and AND3 (N14686, N14673, N13886, N4729);
and AND3 (N14687, N14653, N8733, N5421);
and AND4 (N14688, N14679, N7145, N6713, N2408);
and AND2 (N14689, N14686, N10042);
or OR3 (N14690, N14689, N3996, N13135);
buf BUF1 (N14691, N14674);
not NOT1 (N14692, N14687);
or OR4 (N14693, N14680, N7372, N4835, N10211);
or OR4 (N14694, N14684, N1279, N729, N6527);
nand NAND4 (N14695, N14675, N7288, N10925, N11231);
or OR3 (N14696, N14683, N13082, N4010);
or OR3 (N14697, N14692, N4836, N13731);
and AND3 (N14698, N14685, N10441, N4392);
not NOT1 (N14699, N14691);
xor XOR2 (N14700, N14695, N2538);
buf BUF1 (N14701, N14697);
not NOT1 (N14702, N14670);
or OR4 (N14703, N14696, N6832, N8161, N9070);
nand NAND2 (N14704, N14702, N5487);
nor NOR4 (N14705, N14704, N11517, N6026, N12941);
buf BUF1 (N14706, N14701);
or OR2 (N14707, N14688, N955);
buf BUF1 (N14708, N14698);
xor XOR2 (N14709, N14699, N3407);
or OR4 (N14710, N14700, N4048, N7273, N4782);
buf BUF1 (N14711, N14703);
xor XOR2 (N14712, N14708, N1727);
and AND2 (N14713, N14690, N3283);
nor NOR3 (N14714, N14694, N165, N10230);
and AND4 (N14715, N14712, N9370, N10957, N9696);
buf BUF1 (N14716, N14705);
or OR3 (N14717, N14714, N9765, N14348);
or OR2 (N14718, N14717, N8356);
or OR3 (N14719, N14718, N5095, N1393);
buf BUF1 (N14720, N14716);
xor XOR2 (N14721, N14706, N9631);
nor NOR3 (N14722, N14711, N11515, N5510);
and AND3 (N14723, N14709, N14481, N5285);
and AND3 (N14724, N14722, N14467, N11429);
or OR3 (N14725, N14707, N13147, N1696);
xor XOR2 (N14726, N14723, N7577);
nor NOR4 (N14727, N14720, N8948, N7642, N11882);
and AND3 (N14728, N14719, N2728, N14707);
or OR3 (N14729, N14726, N773, N12247);
nand NAND4 (N14730, N14724, N9906, N3856, N4404);
nor NOR3 (N14731, N14730, N4383, N3476);
xor XOR2 (N14732, N14728, N1149);
nor NOR3 (N14733, N14715, N3593, N6289);
nor NOR4 (N14734, N14729, N4255, N611, N5047);
nand NAND4 (N14735, N14693, N12938, N1959, N3045);
not NOT1 (N14736, N14721);
xor XOR2 (N14737, N14725, N6903);
and AND4 (N14738, N14733, N11613, N12742, N1523);
or OR2 (N14739, N14736, N7064);
or OR2 (N14740, N14737, N1417);
or OR3 (N14741, N14734, N1764, N707);
and AND2 (N14742, N14740, N6040);
nor NOR2 (N14743, N14741, N3072);
and AND3 (N14744, N14732, N3053, N12154);
buf BUF1 (N14745, N14710);
xor XOR2 (N14746, N14739, N3260);
buf BUF1 (N14747, N14743);
and AND2 (N14748, N14742, N980);
and AND3 (N14749, N14748, N9864, N2559);
not NOT1 (N14750, N14738);
nor NOR2 (N14751, N14746, N5499);
buf BUF1 (N14752, N14744);
nand NAND2 (N14753, N14752, N13190);
not NOT1 (N14754, N14753);
and AND2 (N14755, N14713, N14031);
not NOT1 (N14756, N14750);
xor XOR2 (N14757, N14731, N4024);
xor XOR2 (N14758, N14754, N7727);
xor XOR2 (N14759, N14745, N8246);
nand NAND4 (N14760, N14755, N7458, N13465, N10699);
xor XOR2 (N14761, N14747, N11857);
or OR3 (N14762, N14760, N8628, N9031);
or OR4 (N14763, N14757, N13433, N5568, N1056);
xor XOR2 (N14764, N14727, N7730);
not NOT1 (N14765, N14756);
xor XOR2 (N14766, N14763, N14229);
and AND4 (N14767, N14758, N13400, N5443, N3081);
and AND4 (N14768, N14759, N11397, N11449, N12248);
and AND4 (N14769, N14749, N373, N11923, N608);
nand NAND3 (N14770, N14769, N7072, N6904);
or OR3 (N14771, N14768, N5238, N7458);
and AND3 (N14772, N14735, N386, N7095);
nor NOR3 (N14773, N14766, N6414, N10987);
nor NOR3 (N14774, N14767, N8358, N12039);
buf BUF1 (N14775, N14751);
nand NAND4 (N14776, N14771, N6909, N14127, N1068);
and AND2 (N14777, N14765, N3551);
buf BUF1 (N14778, N14774);
nand NAND2 (N14779, N14777, N3117);
xor XOR2 (N14780, N14764, N12473);
nor NOR4 (N14781, N14772, N7584, N9180, N1513);
and AND4 (N14782, N14770, N9563, N3004, N4598);
nor NOR2 (N14783, N14780, N12445);
xor XOR2 (N14784, N14776, N9936);
buf BUF1 (N14785, N14773);
not NOT1 (N14786, N14762);
xor XOR2 (N14787, N14779, N6649);
and AND4 (N14788, N14786, N14257, N13265, N10457);
xor XOR2 (N14789, N14783, N11436);
xor XOR2 (N14790, N14775, N8742);
buf BUF1 (N14791, N14788);
not NOT1 (N14792, N14790);
and AND2 (N14793, N14761, N9948);
nor NOR4 (N14794, N14781, N6682, N8532, N14568);
nand NAND3 (N14795, N14792, N13859, N10900);
nand NAND3 (N14796, N14787, N1542, N4317);
or OR3 (N14797, N14782, N10597, N4073);
or OR3 (N14798, N14794, N12237, N14714);
not NOT1 (N14799, N14789);
and AND3 (N14800, N14795, N5817, N13069);
not NOT1 (N14801, N14796);
nand NAND4 (N14802, N14791, N1577, N1787, N14139);
not NOT1 (N14803, N14785);
nand NAND3 (N14804, N14801, N4633, N11474);
not NOT1 (N14805, N14784);
buf BUF1 (N14806, N14803);
nor NOR3 (N14807, N14793, N9806, N2440);
xor XOR2 (N14808, N14799, N5774);
and AND2 (N14809, N14805, N3802);
and AND3 (N14810, N14807, N8396, N13621);
nor NOR2 (N14811, N14778, N12363);
not NOT1 (N14812, N14800);
and AND2 (N14813, N14812, N3608);
and AND4 (N14814, N14802, N12319, N1451, N5044);
nor NOR4 (N14815, N14810, N6301, N9008, N4316);
or OR3 (N14816, N14815, N6933, N488);
or OR3 (N14817, N14813, N8861, N5652);
xor XOR2 (N14818, N14798, N5197);
or OR3 (N14819, N14814, N9361, N7335);
buf BUF1 (N14820, N14808);
not NOT1 (N14821, N14817);
nor NOR3 (N14822, N14804, N7541, N6691);
xor XOR2 (N14823, N14806, N3149);
nand NAND3 (N14824, N14816, N1638, N7051);
and AND3 (N14825, N14821, N11113, N11534);
nand NAND3 (N14826, N14820, N264, N9676);
nand NAND2 (N14827, N14825, N2771);
xor XOR2 (N14828, N14826, N9822);
nor NOR2 (N14829, N14818, N993);
and AND2 (N14830, N14823, N8423);
not NOT1 (N14831, N14829);
nor NOR3 (N14832, N14811, N4410, N5123);
or OR3 (N14833, N14832, N13383, N8263);
or OR3 (N14834, N14819, N2270, N5760);
not NOT1 (N14835, N14822);
or OR2 (N14836, N14828, N13626);
and AND4 (N14837, N14836, N12971, N11369, N772);
and AND3 (N14838, N14834, N13179, N11027);
xor XOR2 (N14839, N14797, N14591);
nor NOR4 (N14840, N14838, N8184, N9161, N1370);
not NOT1 (N14841, N14809);
xor XOR2 (N14842, N14837, N11379);
xor XOR2 (N14843, N14833, N4010);
or OR2 (N14844, N14835, N6445);
not NOT1 (N14845, N14827);
or OR4 (N14846, N14839, N14057, N13401, N11086);
xor XOR2 (N14847, N14843, N8038);
buf BUF1 (N14848, N14831);
buf BUF1 (N14849, N14841);
buf BUF1 (N14850, N14847);
buf BUF1 (N14851, N14844);
not NOT1 (N14852, N14846);
not NOT1 (N14853, N14848);
xor XOR2 (N14854, N14849, N8590);
buf BUF1 (N14855, N14830);
buf BUF1 (N14856, N14850);
nand NAND2 (N14857, N14840, N5030);
not NOT1 (N14858, N14851);
and AND2 (N14859, N14856, N3814);
and AND2 (N14860, N14855, N7023);
buf BUF1 (N14861, N14824);
xor XOR2 (N14862, N14845, N5599);
xor XOR2 (N14863, N14859, N4173);
buf BUF1 (N14864, N14842);
xor XOR2 (N14865, N14863, N2820);
not NOT1 (N14866, N14862);
nand NAND2 (N14867, N14857, N2871);
nand NAND4 (N14868, N14854, N8763, N7544, N8448);
xor XOR2 (N14869, N14866, N366);
not NOT1 (N14870, N14860);
or OR3 (N14871, N14861, N2854, N4463);
xor XOR2 (N14872, N14868, N3840);
not NOT1 (N14873, N14871);
and AND3 (N14874, N14853, N13635, N12417);
nand NAND4 (N14875, N14852, N6810, N10093, N9464);
or OR4 (N14876, N14872, N8609, N8482, N2244);
buf BUF1 (N14877, N14864);
or OR4 (N14878, N14874, N8485, N8910, N1770);
nand NAND2 (N14879, N14877, N5848);
nand NAND2 (N14880, N14875, N4463);
nor NOR2 (N14881, N14879, N8589);
or OR2 (N14882, N14881, N9976);
nand NAND4 (N14883, N14873, N10741, N5750, N1272);
buf BUF1 (N14884, N14869);
xor XOR2 (N14885, N14884, N14183);
and AND3 (N14886, N14885, N752, N10759);
xor XOR2 (N14887, N14867, N10436);
and AND2 (N14888, N14882, N11574);
nor NOR3 (N14889, N14858, N11549, N4987);
buf BUF1 (N14890, N14880);
buf BUF1 (N14891, N14878);
or OR2 (N14892, N14889, N8608);
buf BUF1 (N14893, N14870);
nand NAND4 (N14894, N14892, N11975, N5418, N9357);
nor NOR4 (N14895, N14893, N14369, N10810, N5853);
xor XOR2 (N14896, N14895, N14868);
nand NAND4 (N14897, N14894, N7443, N10772, N8609);
not NOT1 (N14898, N14891);
xor XOR2 (N14899, N14886, N5262);
not NOT1 (N14900, N14865);
buf BUF1 (N14901, N14898);
nand NAND4 (N14902, N14890, N2580, N12587, N8619);
nor NOR2 (N14903, N14896, N8761);
and AND2 (N14904, N14897, N6839);
and AND4 (N14905, N14903, N12627, N7037, N3581);
not NOT1 (N14906, N14887);
nor NOR4 (N14907, N14901, N2336, N581, N8586);
or OR4 (N14908, N14899, N416, N9388, N8672);
and AND2 (N14909, N14905, N7605);
buf BUF1 (N14910, N14888);
nor NOR4 (N14911, N14904, N13068, N7940, N286);
nor NOR3 (N14912, N14908, N1851, N596);
nor NOR2 (N14913, N14909, N11363);
nand NAND3 (N14914, N14910, N7159, N14720);
nor NOR4 (N14915, N14914, N1969, N8179, N13929);
nand NAND3 (N14916, N14906, N8228, N12397);
buf BUF1 (N14917, N14907);
xor XOR2 (N14918, N14902, N3746);
nand NAND3 (N14919, N14883, N14805, N3805);
nand NAND4 (N14920, N14918, N50, N4316, N13199);
xor XOR2 (N14921, N14913, N10214);
nor NOR2 (N14922, N14921, N6737);
xor XOR2 (N14923, N14900, N4561);
or OR4 (N14924, N14917, N7063, N6075, N8996);
xor XOR2 (N14925, N14923, N14494);
not NOT1 (N14926, N14915);
and AND4 (N14927, N14920, N2528, N12261, N14381);
not NOT1 (N14928, N14912);
or OR3 (N14929, N14919, N11283, N2535);
buf BUF1 (N14930, N14927);
or OR3 (N14931, N14922, N11427, N5214);
nor NOR4 (N14932, N14924, N11590, N13056, N7853);
nand NAND2 (N14933, N14911, N9271);
buf BUF1 (N14934, N14932);
and AND2 (N14935, N14925, N12452);
nor NOR2 (N14936, N14876, N11435);
nor NOR2 (N14937, N14935, N1783);
nand NAND2 (N14938, N14930, N4090);
and AND2 (N14939, N14936, N5826);
not NOT1 (N14940, N14926);
buf BUF1 (N14941, N14940);
and AND3 (N14942, N14941, N9173, N9323);
not NOT1 (N14943, N14938);
not NOT1 (N14944, N14942);
or OR2 (N14945, N14916, N10509);
xor XOR2 (N14946, N14928, N1525);
buf BUF1 (N14947, N14933);
nor NOR3 (N14948, N14937, N13348, N8842);
or OR4 (N14949, N14948, N13576, N52, N14644);
not NOT1 (N14950, N14947);
nor NOR2 (N14951, N14931, N5916);
not NOT1 (N14952, N14929);
xor XOR2 (N14953, N14944, N7126);
buf BUF1 (N14954, N14946);
nor NOR4 (N14955, N14945, N5793, N10599, N3954);
or OR3 (N14956, N14955, N7005, N9061);
nand NAND4 (N14957, N14939, N5838, N5486, N12541);
or OR4 (N14958, N14953, N4776, N13496, N11918);
nand NAND4 (N14959, N14952, N13556, N14321, N11092);
buf BUF1 (N14960, N14957);
and AND2 (N14961, N14951, N7839);
nor NOR4 (N14962, N14960, N7798, N4374, N6877);
not NOT1 (N14963, N14956);
buf BUF1 (N14964, N14962);
and AND4 (N14965, N14958, N3235, N2800, N14215);
or OR2 (N14966, N14954, N9914);
xor XOR2 (N14967, N14966, N9976);
or OR3 (N14968, N14950, N8156, N14799);
not NOT1 (N14969, N14943);
buf BUF1 (N14970, N14965);
xor XOR2 (N14971, N14961, N4262);
nand NAND4 (N14972, N14963, N7440, N708, N10852);
buf BUF1 (N14973, N14959);
not NOT1 (N14974, N14973);
or OR4 (N14975, N14934, N6814, N6582, N3800);
not NOT1 (N14976, N14969);
and AND4 (N14977, N14974, N1704, N10537, N14658);
or OR3 (N14978, N14972, N6932, N12335);
or OR4 (N14979, N14978, N7724, N3930, N3454);
nor NOR2 (N14980, N14967, N6621);
nand NAND3 (N14981, N14968, N1027, N8386);
or OR3 (N14982, N14964, N6996, N9208);
and AND2 (N14983, N14970, N7863);
nand NAND2 (N14984, N14976, N12255);
buf BUF1 (N14985, N14971);
and AND3 (N14986, N14982, N14315, N14947);
and AND2 (N14987, N14986, N6702);
nor NOR4 (N14988, N14987, N1862, N10034, N4602);
or OR4 (N14989, N14983, N14970, N13767, N9074);
and AND4 (N14990, N14977, N7850, N10648, N14402);
and AND2 (N14991, N14988, N13527);
xor XOR2 (N14992, N14949, N13333);
buf BUF1 (N14993, N14975);
and AND3 (N14994, N14989, N10217, N5535);
nor NOR3 (N14995, N14991, N64, N10079);
not NOT1 (N14996, N14984);
xor XOR2 (N14997, N14995, N2481);
not NOT1 (N14998, N14980);
and AND2 (N14999, N14998, N1126);
xor XOR2 (N15000, N14994, N2236);
nand NAND4 (N15001, N14981, N11098, N13259, N7447);
nand NAND4 (N15002, N14996, N12987, N13091, N11864);
xor XOR2 (N15003, N15001, N6831);
nor NOR3 (N15004, N14997, N7138, N12318);
xor XOR2 (N15005, N14985, N8857);
xor XOR2 (N15006, N14990, N10497);
or OR2 (N15007, N15006, N6678);
not NOT1 (N15008, N15002);
and AND2 (N15009, N15008, N3059);
nor NOR4 (N15010, N14993, N5976, N10606, N295);
and AND3 (N15011, N15003, N6938, N14770);
xor XOR2 (N15012, N15011, N4263);
xor XOR2 (N15013, N14999, N13945);
buf BUF1 (N15014, N15012);
and AND4 (N15015, N15000, N15001, N14815, N11273);
and AND4 (N15016, N15015, N5522, N4996, N14041);
xor XOR2 (N15017, N15013, N10625);
or OR3 (N15018, N15017, N6650, N1893);
and AND3 (N15019, N14992, N2076, N3132);
and AND3 (N15020, N15004, N14972, N14994);
not NOT1 (N15021, N15007);
nor NOR4 (N15022, N15010, N12647, N12669, N5974);
buf BUF1 (N15023, N15014);
or OR4 (N15024, N15016, N6800, N13871, N11688);
not NOT1 (N15025, N15023);
and AND2 (N15026, N15024, N9072);
nand NAND4 (N15027, N15018, N1787, N8843, N14385);
or OR4 (N15028, N15021, N14020, N2621, N2637);
nor NOR4 (N15029, N15019, N1978, N8549, N4655);
and AND2 (N15030, N15029, N2872);
buf BUF1 (N15031, N15028);
nand NAND4 (N15032, N15022, N8607, N5356, N2097);
buf BUF1 (N15033, N15032);
and AND3 (N15034, N15026, N14795, N3150);
or OR2 (N15035, N15020, N7225);
or OR3 (N15036, N15031, N11260, N3607);
not NOT1 (N15037, N15025);
nor NOR4 (N15038, N15037, N9964, N9144, N5252);
and AND4 (N15039, N15027, N8356, N6067, N5546);
nand NAND2 (N15040, N15005, N7393);
and AND2 (N15041, N15039, N7899);
or OR3 (N15042, N15030, N10888, N3602);
nor NOR2 (N15043, N14979, N5566);
xor XOR2 (N15044, N15035, N9812);
buf BUF1 (N15045, N15043);
buf BUF1 (N15046, N15044);
nand NAND4 (N15047, N15042, N2908, N9166, N8235);
nand NAND4 (N15048, N15046, N4770, N930, N3919);
not NOT1 (N15049, N15047);
nand NAND3 (N15050, N15040, N4657, N5221);
nand NAND2 (N15051, N15049, N557);
or OR3 (N15052, N15051, N551, N9390);
buf BUF1 (N15053, N15045);
not NOT1 (N15054, N15041);
nand NAND4 (N15055, N15034, N9598, N10438, N14299);
buf BUF1 (N15056, N15048);
and AND4 (N15057, N15009, N1118, N7789, N3552);
nand NAND4 (N15058, N15050, N11328, N3099, N3678);
nor NOR3 (N15059, N15053, N8502, N2396);
xor XOR2 (N15060, N15054, N5040);
buf BUF1 (N15061, N15055);
and AND2 (N15062, N15036, N3560);
nand NAND3 (N15063, N15062, N12779, N14417);
not NOT1 (N15064, N15063);
buf BUF1 (N15065, N15058);
nor NOR3 (N15066, N15060, N13830, N1646);
and AND2 (N15067, N15064, N715);
not NOT1 (N15068, N15065);
or OR2 (N15069, N15033, N3692);
buf BUF1 (N15070, N15052);
nor NOR4 (N15071, N15056, N6488, N14078, N12992);
or OR3 (N15072, N15070, N6341, N14386);
and AND4 (N15073, N15061, N11752, N10204, N8420);
and AND3 (N15074, N15072, N14615, N6719);
xor XOR2 (N15075, N15057, N12946);
or OR4 (N15076, N15067, N36, N168, N7122);
nor NOR3 (N15077, N15066, N14745, N6541);
nand NAND2 (N15078, N15038, N12195);
and AND3 (N15079, N15075, N1842, N13703);
buf BUF1 (N15080, N15071);
and AND2 (N15081, N15079, N12697);
xor XOR2 (N15082, N15080, N479);
nand NAND4 (N15083, N15082, N5059, N10091, N10591);
not NOT1 (N15084, N15083);
and AND4 (N15085, N15073, N6618, N2950, N14983);
nor NOR3 (N15086, N15077, N13480, N11018);
and AND3 (N15087, N15081, N7777, N11849);
xor XOR2 (N15088, N15076, N5465);
not NOT1 (N15089, N15069);
or OR3 (N15090, N15088, N14185, N4139);
xor XOR2 (N15091, N15090, N11860);
xor XOR2 (N15092, N15087, N12630);
not NOT1 (N15093, N15092);
or OR3 (N15094, N15068, N6166, N7838);
not NOT1 (N15095, N15086);
nor NOR3 (N15096, N15091, N10945, N8962);
or OR2 (N15097, N15078, N7120);
buf BUF1 (N15098, N15059);
and AND3 (N15099, N15074, N14730, N14976);
xor XOR2 (N15100, N15089, N1148);
nor NOR2 (N15101, N15095, N13659);
nand NAND2 (N15102, N15101, N5786);
not NOT1 (N15103, N15102);
or OR2 (N15104, N15085, N14852);
or OR2 (N15105, N15103, N7622);
nor NOR4 (N15106, N15093, N4774, N5085, N14928);
nand NAND2 (N15107, N15097, N10629);
xor XOR2 (N15108, N15105, N11155);
xor XOR2 (N15109, N15104, N10449);
or OR4 (N15110, N15098, N2496, N14748, N426);
nand NAND2 (N15111, N15107, N10822);
buf BUF1 (N15112, N15099);
xor XOR2 (N15113, N15084, N6676);
buf BUF1 (N15114, N15110);
nand NAND2 (N15115, N15114, N3154);
nand NAND2 (N15116, N15096, N9181);
not NOT1 (N15117, N15108);
or OR3 (N15118, N15117, N15100, N11787);
not NOT1 (N15119, N3257);
not NOT1 (N15120, N15116);
not NOT1 (N15121, N15109);
buf BUF1 (N15122, N15113);
nand NAND4 (N15123, N15118, N14316, N4879, N11067);
not NOT1 (N15124, N15121);
and AND2 (N15125, N15094, N10007);
or OR4 (N15126, N15123, N1235, N13641, N10103);
buf BUF1 (N15127, N15119);
nor NOR3 (N15128, N15125, N13268, N14481);
xor XOR2 (N15129, N15112, N1415);
not NOT1 (N15130, N15115);
not NOT1 (N15131, N15127);
and AND3 (N15132, N15106, N12283, N14940);
nand NAND4 (N15133, N15120, N13458, N2692, N6183);
buf BUF1 (N15134, N15133);
not NOT1 (N15135, N15126);
nor NOR4 (N15136, N15124, N8841, N1911, N9694);
nand NAND3 (N15137, N15130, N13368, N264);
or OR2 (N15138, N15122, N14624);
or OR3 (N15139, N15134, N2742, N12849);
nand NAND2 (N15140, N15138, N11090);
and AND4 (N15141, N15129, N14095, N8916, N11523);
and AND4 (N15142, N15137, N5043, N6006, N6785);
nor NOR2 (N15143, N15135, N11784);
xor XOR2 (N15144, N15111, N4295);
and AND3 (N15145, N15142, N10638, N13612);
nor NOR3 (N15146, N15139, N10185, N6979);
buf BUF1 (N15147, N15145);
not NOT1 (N15148, N15143);
nand NAND4 (N15149, N15141, N14938, N1808, N12962);
or OR4 (N15150, N15144, N3685, N7371, N3121);
xor XOR2 (N15151, N15131, N6672);
buf BUF1 (N15152, N15147);
nor NOR4 (N15153, N15136, N2521, N12674, N9071);
nor NOR4 (N15154, N15151, N14836, N6264, N682);
not NOT1 (N15155, N15132);
nand NAND3 (N15156, N15146, N1520, N2412);
nor NOR2 (N15157, N15149, N3142);
nand NAND3 (N15158, N15153, N3710, N6641);
not NOT1 (N15159, N15128);
and AND2 (N15160, N15152, N10273);
nand NAND4 (N15161, N15140, N1329, N11876, N2702);
or OR4 (N15162, N15158, N7650, N280, N3619);
and AND3 (N15163, N15159, N5686, N5215);
or OR3 (N15164, N15160, N6975, N9720);
nor NOR2 (N15165, N15161, N6372);
nor NOR2 (N15166, N15150, N7654);
xor XOR2 (N15167, N15156, N15133);
buf BUF1 (N15168, N15164);
or OR2 (N15169, N15166, N11463);
nand NAND3 (N15170, N15169, N11649, N13304);
nor NOR3 (N15171, N15168, N6472, N12749);
xor XOR2 (N15172, N15170, N11027);
nor NOR2 (N15173, N15163, N1363);
and AND3 (N15174, N15154, N7455, N10204);
nand NAND4 (N15175, N15174, N11903, N11834, N6053);
xor XOR2 (N15176, N15165, N9036);
or OR4 (N15177, N15176, N13079, N2524, N106);
nand NAND3 (N15178, N15171, N1026, N346);
xor XOR2 (N15179, N15178, N5770);
and AND4 (N15180, N15162, N2874, N10679, N14056);
nand NAND2 (N15181, N15167, N12115);
and AND3 (N15182, N15179, N7164, N12802);
not NOT1 (N15183, N15177);
nand NAND2 (N15184, N15172, N4240);
and AND2 (N15185, N15181, N11129);
not NOT1 (N15186, N15157);
or OR3 (N15187, N15180, N2303, N4260);
buf BUF1 (N15188, N15187);
or OR3 (N15189, N15188, N5711, N2171);
buf BUF1 (N15190, N15148);
or OR4 (N15191, N15184, N14532, N10134, N1641);
buf BUF1 (N15192, N15155);
nand NAND2 (N15193, N15189, N9945);
and AND4 (N15194, N15173, N8723, N2131, N3808);
nand NAND3 (N15195, N15175, N10310, N9727);
and AND2 (N15196, N15193, N13959);
and AND2 (N15197, N15183, N8473);
xor XOR2 (N15198, N15194, N569);
not NOT1 (N15199, N15196);
nor NOR4 (N15200, N15186, N13650, N1925, N3568);
nand NAND2 (N15201, N15198, N10542);
xor XOR2 (N15202, N15190, N3070);
or OR4 (N15203, N15185, N791, N4680, N9134);
buf BUF1 (N15204, N15195);
nor NOR3 (N15205, N15182, N468, N8479);
xor XOR2 (N15206, N15202, N9254);
buf BUF1 (N15207, N15206);
buf BUF1 (N15208, N15192);
or OR4 (N15209, N15207, N14614, N6179, N2398);
nand NAND3 (N15210, N15201, N2635, N6075);
xor XOR2 (N15211, N15200, N666);
xor XOR2 (N15212, N15197, N9280);
nor NOR4 (N15213, N15199, N7622, N8532, N3676);
and AND2 (N15214, N15213, N12128);
nor NOR2 (N15215, N15208, N11893);
nor NOR3 (N15216, N15191, N4582, N12264);
nand NAND3 (N15217, N15209, N1712, N5977);
nand NAND3 (N15218, N15204, N9777, N4995);
and AND4 (N15219, N15211, N13697, N6965, N14761);
nor NOR4 (N15220, N15212, N4673, N8204, N6141);
xor XOR2 (N15221, N15214, N7253);
or OR4 (N15222, N15205, N10701, N13530, N10070);
nor NOR3 (N15223, N15219, N6258, N12622);
and AND3 (N15224, N15220, N14585, N1442);
nand NAND3 (N15225, N15215, N3556, N7043);
and AND4 (N15226, N15217, N10889, N14094, N9026);
buf BUF1 (N15227, N15226);
not NOT1 (N15228, N15225);
not NOT1 (N15229, N15203);
and AND3 (N15230, N15228, N13172, N13437);
nor NOR3 (N15231, N15222, N12255, N9428);
or OR2 (N15232, N15216, N8397);
not NOT1 (N15233, N15230);
not NOT1 (N15234, N15227);
not NOT1 (N15235, N15233);
not NOT1 (N15236, N15235);
nand NAND3 (N15237, N15221, N14350, N3510);
not NOT1 (N15238, N15232);
or OR2 (N15239, N15224, N9759);
nand NAND4 (N15240, N15231, N1533, N6878, N9820);
and AND3 (N15241, N15238, N12960, N7002);
buf BUF1 (N15242, N15241);
xor XOR2 (N15243, N15236, N5618);
buf BUF1 (N15244, N15210);
and AND4 (N15245, N15239, N7438, N1130, N4603);
nor NOR3 (N15246, N15218, N8948, N15085);
not NOT1 (N15247, N15234);
and AND2 (N15248, N15247, N7301);
and AND3 (N15249, N15244, N8158, N799);
buf BUF1 (N15250, N15242);
and AND4 (N15251, N15229, N10367, N3365, N9108);
and AND2 (N15252, N15248, N6856);
or OR4 (N15253, N15252, N7575, N14512, N8762);
buf BUF1 (N15254, N15240);
buf BUF1 (N15255, N15243);
buf BUF1 (N15256, N15246);
buf BUF1 (N15257, N15250);
nand NAND3 (N15258, N15251, N4774, N14516);
nand NAND4 (N15259, N15256, N9098, N12822, N8867);
nand NAND3 (N15260, N15245, N12654, N3661);
and AND2 (N15261, N15255, N7955);
nand NAND2 (N15262, N15254, N1684);
or OR3 (N15263, N15259, N7072, N12308);
nor NOR4 (N15264, N15263, N5982, N11865, N14197);
or OR4 (N15265, N15237, N7935, N13429, N7646);
xor XOR2 (N15266, N15265, N5297);
xor XOR2 (N15267, N15253, N13486);
xor XOR2 (N15268, N15223, N6227);
nor NOR4 (N15269, N15266, N2817, N12746, N7801);
xor XOR2 (N15270, N15261, N4249);
or OR4 (N15271, N15257, N5909, N2003, N11107);
buf BUF1 (N15272, N15270);
not NOT1 (N15273, N15268);
xor XOR2 (N15274, N15249, N9022);
not NOT1 (N15275, N15267);
xor XOR2 (N15276, N15271, N13229);
nand NAND4 (N15277, N15273, N10064, N14969, N1679);
xor XOR2 (N15278, N15277, N9447);
not NOT1 (N15279, N15260);
nor NOR2 (N15280, N15264, N9313);
nand NAND4 (N15281, N15279, N7383, N345, N13913);
nand NAND3 (N15282, N15280, N757, N11194);
and AND4 (N15283, N15281, N5262, N5304, N9888);
or OR3 (N15284, N15262, N6526, N9170);
nor NOR3 (N15285, N15274, N8224, N12683);
not NOT1 (N15286, N15258);
not NOT1 (N15287, N15285);
and AND3 (N15288, N15286, N2926, N5728);
buf BUF1 (N15289, N15282);
or OR2 (N15290, N15284, N10069);
xor XOR2 (N15291, N15287, N12825);
nand NAND2 (N15292, N15283, N12519);
or OR2 (N15293, N15276, N3215);
buf BUF1 (N15294, N15288);
xor XOR2 (N15295, N15272, N12424);
xor XOR2 (N15296, N15292, N4651);
and AND2 (N15297, N15269, N12263);
and AND3 (N15298, N15289, N3706, N6383);
nor NOR4 (N15299, N15295, N11993, N3924, N11911);
xor XOR2 (N15300, N15296, N5681);
not NOT1 (N15301, N15300);
nand NAND2 (N15302, N15291, N13582);
nor NOR3 (N15303, N15299, N7123, N6216);
buf BUF1 (N15304, N15301);
and AND2 (N15305, N15294, N9583);
xor XOR2 (N15306, N15304, N14417);
nand NAND2 (N15307, N15290, N3706);
xor XOR2 (N15308, N15293, N8063);
nor NOR2 (N15309, N15298, N12482);
buf BUF1 (N15310, N15306);
nor NOR4 (N15311, N15309, N10622, N9490, N6142);
nor NOR4 (N15312, N15311, N9682, N2567, N7166);
nand NAND4 (N15313, N15310, N10208, N9886, N11268);
nand NAND3 (N15314, N15312, N3143, N7621);
nor NOR3 (N15315, N15275, N3064, N9016);
or OR4 (N15316, N15305, N2375, N5345, N2021);
buf BUF1 (N15317, N15302);
and AND2 (N15318, N15316, N1799);
not NOT1 (N15319, N15314);
xor XOR2 (N15320, N15278, N836);
or OR3 (N15321, N15297, N14780, N3694);
nor NOR2 (N15322, N15318, N1753);
buf BUF1 (N15323, N15315);
buf BUF1 (N15324, N15307);
and AND2 (N15325, N15313, N8569);
or OR4 (N15326, N15325, N10189, N6724, N14597);
and AND3 (N15327, N15321, N13176, N13542);
xor XOR2 (N15328, N15303, N2404);
or OR4 (N15329, N15326, N9867, N2150, N9883);
buf BUF1 (N15330, N15317);
buf BUF1 (N15331, N15330);
or OR4 (N15332, N15328, N6552, N10090, N7783);
or OR4 (N15333, N15308, N628, N15215, N1276);
not NOT1 (N15334, N15320);
or OR3 (N15335, N15334, N14229, N1972);
xor XOR2 (N15336, N15327, N14537);
xor XOR2 (N15337, N15319, N9409);
xor XOR2 (N15338, N15336, N3818);
or OR3 (N15339, N15331, N10945, N2109);
nor NOR4 (N15340, N15329, N440, N6892, N6573);
nand NAND4 (N15341, N15322, N15277, N6351, N2434);
and AND3 (N15342, N15340, N320, N14241);
nor NOR2 (N15343, N15338, N10325);
xor XOR2 (N15344, N15343, N3673);
and AND3 (N15345, N15337, N14028, N77);
xor XOR2 (N15346, N15324, N10712);
nor NOR2 (N15347, N15341, N13775);
xor XOR2 (N15348, N15345, N3889);
xor XOR2 (N15349, N15348, N2406);
xor XOR2 (N15350, N15346, N1602);
not NOT1 (N15351, N15344);
buf BUF1 (N15352, N15333);
not NOT1 (N15353, N15335);
or OR2 (N15354, N15332, N9971);
and AND4 (N15355, N15349, N4067, N3875, N7561);
nor NOR3 (N15356, N15353, N4377, N7662);
not NOT1 (N15357, N15323);
nand NAND3 (N15358, N15350, N1606, N8803);
or OR3 (N15359, N15351, N2139, N12416);
nor NOR4 (N15360, N15356, N2643, N5026, N433);
or OR4 (N15361, N15339, N7940, N8127, N8244);
not NOT1 (N15362, N15347);
not NOT1 (N15363, N15358);
nand NAND3 (N15364, N15357, N14916, N3448);
nand NAND3 (N15365, N15363, N8768, N8142);
buf BUF1 (N15366, N15352);
and AND2 (N15367, N15355, N5319);
nor NOR2 (N15368, N15360, N1053);
buf BUF1 (N15369, N15362);
or OR3 (N15370, N15368, N15321, N6796);
xor XOR2 (N15371, N15369, N10441);
and AND2 (N15372, N15371, N4781);
nor NOR4 (N15373, N15361, N4477, N1351, N5879);
not NOT1 (N15374, N15342);
xor XOR2 (N15375, N15354, N2880);
buf BUF1 (N15376, N15359);
nor NOR3 (N15377, N15375, N10164, N10375);
buf BUF1 (N15378, N15377);
xor XOR2 (N15379, N15367, N4564);
nor NOR2 (N15380, N15378, N941);
nand NAND4 (N15381, N15372, N10994, N8034, N12485);
buf BUF1 (N15382, N15376);
and AND3 (N15383, N15379, N15286, N650);
buf BUF1 (N15384, N15374);
or OR4 (N15385, N15383, N14683, N5243, N11040);
xor XOR2 (N15386, N15384, N7780);
xor XOR2 (N15387, N15366, N4875);
and AND3 (N15388, N15365, N10123, N1167);
nand NAND2 (N15389, N15373, N2307);
not NOT1 (N15390, N15387);
and AND2 (N15391, N15389, N12288);
or OR2 (N15392, N15385, N11936);
xor XOR2 (N15393, N15392, N9584);
nand NAND2 (N15394, N15370, N14248);
and AND2 (N15395, N15391, N15388);
buf BUF1 (N15396, N1639);
and AND2 (N15397, N15364, N9963);
nor NOR3 (N15398, N15380, N1904, N11205);
or OR3 (N15399, N15394, N14019, N4005);
nand NAND2 (N15400, N15393, N2180);
nand NAND3 (N15401, N15386, N10641, N14875);
not NOT1 (N15402, N15382);
or OR4 (N15403, N15400, N3142, N12465, N6355);
not NOT1 (N15404, N15399);
nand NAND3 (N15405, N15397, N2228, N11815);
xor XOR2 (N15406, N15381, N11201);
nand NAND4 (N15407, N15404, N11395, N10393, N12254);
nand NAND4 (N15408, N15395, N12587, N2816, N6711);
nor NOR3 (N15409, N15403, N14418, N11673);
not NOT1 (N15410, N15408);
not NOT1 (N15411, N15396);
xor XOR2 (N15412, N15407, N1010);
not NOT1 (N15413, N15405);
xor XOR2 (N15414, N15406, N6905);
xor XOR2 (N15415, N15402, N10668);
not NOT1 (N15416, N15414);
nor NOR2 (N15417, N15401, N8136);
nand NAND3 (N15418, N15410, N10720, N4521);
and AND3 (N15419, N15415, N10692, N11520);
nor NOR3 (N15420, N15411, N875, N12921);
not NOT1 (N15421, N15416);
nor NOR4 (N15422, N15421, N5817, N7404, N11693);
not NOT1 (N15423, N15417);
xor XOR2 (N15424, N15409, N4201);
xor XOR2 (N15425, N15422, N7575);
nor NOR2 (N15426, N15424, N10006);
nor NOR2 (N15427, N15426, N974);
nand NAND2 (N15428, N15419, N4277);
xor XOR2 (N15429, N15398, N4484);
not NOT1 (N15430, N15418);
nand NAND4 (N15431, N15412, N6508, N8027, N3562);
and AND4 (N15432, N15430, N282, N13835, N4346);
or OR4 (N15433, N15420, N11120, N6808, N7727);
nand NAND3 (N15434, N15429, N9592, N7189);
or OR3 (N15435, N15390, N522, N6491);
not NOT1 (N15436, N15433);
or OR4 (N15437, N15427, N3443, N13846, N9304);
or OR4 (N15438, N15423, N1104, N8186, N14044);
buf BUF1 (N15439, N15413);
or OR2 (N15440, N15439, N1773);
and AND4 (N15441, N15435, N14854, N10337, N893);
buf BUF1 (N15442, N15431);
not NOT1 (N15443, N15425);
or OR2 (N15444, N15441, N4985);
nor NOR3 (N15445, N15436, N4675, N3564);
xor XOR2 (N15446, N15445, N11707);
buf BUF1 (N15447, N15446);
xor XOR2 (N15448, N15442, N13499);
nor NOR4 (N15449, N15428, N9498, N2485, N13144);
nand NAND4 (N15450, N15440, N6134, N1938, N5712);
nand NAND4 (N15451, N15448, N3980, N13749, N10847);
nand NAND2 (N15452, N15437, N1201);
xor XOR2 (N15453, N15449, N294);
nor NOR3 (N15454, N15438, N3269, N5035);
xor XOR2 (N15455, N15452, N1251);
xor XOR2 (N15456, N15434, N3865);
nor NOR3 (N15457, N15443, N12353, N9602);
and AND3 (N15458, N15451, N7776, N1820);
and AND2 (N15459, N15432, N7243);
nand NAND3 (N15460, N15459, N8761, N4644);
or OR4 (N15461, N15460, N863, N8177, N6785);
and AND3 (N15462, N15450, N2969, N2784);
xor XOR2 (N15463, N15458, N13385);
not NOT1 (N15464, N15444);
nor NOR2 (N15465, N15463, N1255);
and AND2 (N15466, N15454, N14634);
nor NOR4 (N15467, N15447, N9430, N14243, N8124);
or OR3 (N15468, N15462, N14457, N2414);
buf BUF1 (N15469, N15456);
nor NOR4 (N15470, N15457, N10681, N7556, N3700);
xor XOR2 (N15471, N15467, N6576);
buf BUF1 (N15472, N15471);
nand NAND3 (N15473, N15461, N6473, N2474);
and AND2 (N15474, N15464, N14205);
xor XOR2 (N15475, N15473, N8472);
buf BUF1 (N15476, N15468);
not NOT1 (N15477, N15474);
and AND2 (N15478, N15472, N8811);
or OR3 (N15479, N15469, N9858, N14926);
or OR3 (N15480, N15478, N10467, N107);
not NOT1 (N15481, N15479);
not NOT1 (N15482, N15480);
and AND4 (N15483, N15475, N7966, N2981, N12825);
and AND3 (N15484, N15477, N12539, N13914);
nor NOR4 (N15485, N15470, N14160, N8406, N10634);
buf BUF1 (N15486, N15481);
and AND2 (N15487, N15466, N8457);
nor NOR2 (N15488, N15455, N7934);
nor NOR4 (N15489, N15453, N11957, N6914, N2600);
or OR3 (N15490, N15489, N14381, N7700);
not NOT1 (N15491, N15486);
nand NAND2 (N15492, N15482, N7452);
xor XOR2 (N15493, N15484, N1097);
xor XOR2 (N15494, N15485, N8080);
xor XOR2 (N15495, N15488, N5306);
not NOT1 (N15496, N15490);
not NOT1 (N15497, N15465);
nor NOR2 (N15498, N15495, N14333);
nand NAND2 (N15499, N15476, N10386);
buf BUF1 (N15500, N15492);
or OR3 (N15501, N15497, N3319, N11248);
nand NAND2 (N15502, N15483, N9561);
not NOT1 (N15503, N15500);
and AND4 (N15504, N15503, N2396, N3979, N5408);
nor NOR4 (N15505, N15493, N7749, N3531, N6047);
nor NOR2 (N15506, N15502, N2306);
or OR3 (N15507, N15496, N4414, N13357);
or OR2 (N15508, N15487, N7959);
buf BUF1 (N15509, N15499);
and AND3 (N15510, N15498, N8126, N12546);
nand NAND2 (N15511, N15508, N1528);
xor XOR2 (N15512, N15491, N1860);
or OR3 (N15513, N15506, N5784, N14894);
nor NOR4 (N15514, N15513, N13020, N2568, N3606);
and AND2 (N15515, N15510, N10282);
and AND3 (N15516, N15512, N11625, N14395);
nand NAND3 (N15517, N15505, N12976, N1933);
nand NAND4 (N15518, N15514, N13135, N3191, N11593);
xor XOR2 (N15519, N15515, N7267);
xor XOR2 (N15520, N15504, N12664);
and AND2 (N15521, N15501, N1401);
and AND3 (N15522, N15519, N4136, N15458);
not NOT1 (N15523, N15516);
buf BUF1 (N15524, N15523);
and AND2 (N15525, N15511, N12168);
not NOT1 (N15526, N15494);
nand NAND4 (N15527, N15520, N2823, N7760, N3158);
or OR3 (N15528, N15522, N2383, N4829);
and AND4 (N15529, N15507, N12946, N15295, N4413);
or OR2 (N15530, N15518, N5217);
or OR2 (N15531, N15509, N8922);
xor XOR2 (N15532, N15525, N319);
nand NAND2 (N15533, N15532, N13049);
buf BUF1 (N15534, N15521);
buf BUF1 (N15535, N15524);
nand NAND4 (N15536, N15527, N5439, N9151, N14540);
buf BUF1 (N15537, N15531);
buf BUF1 (N15538, N15529);
xor XOR2 (N15539, N15535, N14486);
nor NOR2 (N15540, N15528, N7705);
not NOT1 (N15541, N15539);
xor XOR2 (N15542, N15537, N5342);
and AND2 (N15543, N15530, N9875);
and AND3 (N15544, N15543, N256, N5786);
nand NAND2 (N15545, N15534, N4669);
nor NOR3 (N15546, N15526, N9071, N3222);
nor NOR4 (N15547, N15538, N15013, N5350, N2408);
xor XOR2 (N15548, N15517, N6502);
not NOT1 (N15549, N15547);
or OR4 (N15550, N15544, N7879, N12698, N6621);
not NOT1 (N15551, N15546);
not NOT1 (N15552, N15541);
and AND4 (N15553, N15545, N13031, N642, N12464);
nor NOR2 (N15554, N15553, N1882);
buf BUF1 (N15555, N15542);
nor NOR2 (N15556, N15550, N1618);
and AND2 (N15557, N15555, N5336);
xor XOR2 (N15558, N15552, N12835);
buf BUF1 (N15559, N15536);
and AND4 (N15560, N15556, N13569, N1167, N102);
xor XOR2 (N15561, N15558, N4866);
xor XOR2 (N15562, N15560, N2089);
nor NOR4 (N15563, N15551, N8022, N2590, N5588);
and AND2 (N15564, N15554, N5683);
or OR4 (N15565, N15561, N2848, N8633, N13561);
buf BUF1 (N15566, N15559);
and AND4 (N15567, N15548, N1394, N1289, N14763);
and AND4 (N15568, N15563, N12874, N1057, N2257);
nand NAND2 (N15569, N15557, N10625);
buf BUF1 (N15570, N15549);
not NOT1 (N15571, N15568);
nor NOR3 (N15572, N15540, N11721, N5510);
and AND4 (N15573, N15533, N11225, N7014, N7382);
nand NAND2 (N15574, N15572, N2765);
buf BUF1 (N15575, N15574);
or OR4 (N15576, N15566, N1878, N2452, N12846);
and AND3 (N15577, N15571, N1839, N14171);
nor NOR4 (N15578, N15564, N13474, N7978, N1665);
not NOT1 (N15579, N15576);
or OR2 (N15580, N15578, N400);
not NOT1 (N15581, N15577);
or OR4 (N15582, N15581, N1133, N14228, N6577);
xor XOR2 (N15583, N15569, N4752);
buf BUF1 (N15584, N15567);
nor NOR4 (N15585, N15580, N5461, N7478, N5856);
not NOT1 (N15586, N15570);
and AND2 (N15587, N15583, N1751);
nand NAND4 (N15588, N15582, N10061, N5639, N12464);
xor XOR2 (N15589, N15588, N14830);
nor NOR4 (N15590, N15579, N1988, N11525, N1454);
buf BUF1 (N15591, N15587);
buf BUF1 (N15592, N15562);
xor XOR2 (N15593, N15585, N3410);
xor XOR2 (N15594, N15586, N5953);
nor NOR4 (N15595, N15590, N7486, N7455, N9609);
xor XOR2 (N15596, N15591, N5247);
xor XOR2 (N15597, N15596, N4512);
nand NAND3 (N15598, N15589, N1758, N9958);
nor NOR3 (N15599, N15594, N8401, N11153);
buf BUF1 (N15600, N15575);
and AND4 (N15601, N15597, N1966, N1811, N2293);
xor XOR2 (N15602, N15601, N11407);
xor XOR2 (N15603, N15593, N6941);
not NOT1 (N15604, N15599);
nand NAND4 (N15605, N15595, N4365, N12798, N12217);
and AND2 (N15606, N15584, N10061);
or OR3 (N15607, N15604, N9511, N3093);
not NOT1 (N15608, N15573);
buf BUF1 (N15609, N15602);
buf BUF1 (N15610, N15605);
and AND3 (N15611, N15592, N3708, N6);
buf BUF1 (N15612, N15610);
not NOT1 (N15613, N15609);
xor XOR2 (N15614, N15607, N14723);
nand NAND3 (N15615, N15565, N15385, N310);
or OR3 (N15616, N15611, N8726, N10658);
nand NAND3 (N15617, N15600, N3844, N11994);
or OR4 (N15618, N15612, N15265, N13371, N15233);
xor XOR2 (N15619, N15617, N11766);
buf BUF1 (N15620, N15613);
not NOT1 (N15621, N15620);
not NOT1 (N15622, N15608);
buf BUF1 (N15623, N15598);
not NOT1 (N15624, N15606);
nor NOR2 (N15625, N15616, N8658);
and AND2 (N15626, N15603, N7926);
nor NOR3 (N15627, N15621, N12460, N10658);
or OR2 (N15628, N15627, N12266);
buf BUF1 (N15629, N15622);
not NOT1 (N15630, N15624);
or OR2 (N15631, N15623, N912);
xor XOR2 (N15632, N15618, N15434);
nand NAND3 (N15633, N15615, N7772, N271);
and AND2 (N15634, N15628, N6510);
nor NOR4 (N15635, N15630, N15004, N12272, N4081);
not NOT1 (N15636, N15625);
and AND3 (N15637, N15631, N36, N12100);
xor XOR2 (N15638, N15636, N2363);
nand NAND4 (N15639, N15638, N6716, N3555, N2950);
not NOT1 (N15640, N15632);
xor XOR2 (N15641, N15637, N824);
xor XOR2 (N15642, N15634, N6640);
xor XOR2 (N15643, N15640, N2192);
or OR4 (N15644, N15639, N13373, N2570, N13243);
and AND4 (N15645, N15644, N12296, N13605, N2972);
xor XOR2 (N15646, N15633, N8669);
not NOT1 (N15647, N15614);
buf BUF1 (N15648, N15629);
buf BUF1 (N15649, N15626);
nor NOR4 (N15650, N15643, N4113, N14021, N11516);
not NOT1 (N15651, N15646);
nand NAND2 (N15652, N15647, N1058);
not NOT1 (N15653, N15648);
xor XOR2 (N15654, N15649, N7141);
nand NAND2 (N15655, N15653, N8576);
not NOT1 (N15656, N15650);
and AND2 (N15657, N15642, N7104);
xor XOR2 (N15658, N15652, N12843);
and AND2 (N15659, N15619, N3651);
or OR4 (N15660, N15657, N8466, N15457, N1784);
not NOT1 (N15661, N15658);
not NOT1 (N15662, N15645);
or OR2 (N15663, N15641, N6144);
and AND4 (N15664, N15663, N1505, N14201, N13413);
not NOT1 (N15665, N15660);
nor NOR4 (N15666, N15635, N7485, N7467, N932);
buf BUF1 (N15667, N15654);
or OR4 (N15668, N15665, N10014, N15537, N14028);
and AND4 (N15669, N15662, N13895, N7157, N6690);
nand NAND4 (N15670, N15668, N11165, N758, N2135);
buf BUF1 (N15671, N15655);
not NOT1 (N15672, N15669);
not NOT1 (N15673, N15671);
and AND3 (N15674, N15661, N9759, N12160);
nand NAND4 (N15675, N15656, N10391, N13524, N14613);
buf BUF1 (N15676, N15664);
nor NOR2 (N15677, N15675, N10494);
or OR4 (N15678, N15667, N4185, N4620, N3680);
nor NOR2 (N15679, N15673, N14037);
xor XOR2 (N15680, N15678, N13237);
nand NAND4 (N15681, N15670, N1902, N12537, N12703);
nor NOR4 (N15682, N15681, N5176, N11790, N13465);
xor XOR2 (N15683, N15659, N12738);
not NOT1 (N15684, N15651);
nand NAND3 (N15685, N15683, N6070, N3737);
xor XOR2 (N15686, N15666, N12925);
nand NAND4 (N15687, N15685, N14682, N10226, N4931);
xor XOR2 (N15688, N15686, N10438);
xor XOR2 (N15689, N15688, N13311);
xor XOR2 (N15690, N15680, N743);
xor XOR2 (N15691, N15672, N6955);
xor XOR2 (N15692, N15684, N14609);
not NOT1 (N15693, N15682);
nand NAND2 (N15694, N15689, N9733);
not NOT1 (N15695, N15676);
buf BUF1 (N15696, N15674);
nand NAND3 (N15697, N15693, N11755, N2399);
or OR3 (N15698, N15687, N14868, N7654);
buf BUF1 (N15699, N15691);
not NOT1 (N15700, N15695);
xor XOR2 (N15701, N15696, N15618);
and AND4 (N15702, N15677, N10567, N6440, N4828);
and AND3 (N15703, N15700, N11888, N15644);
nand NAND4 (N15704, N15692, N1518, N6366, N12099);
xor XOR2 (N15705, N15697, N15458);
and AND4 (N15706, N15699, N852, N2713, N9674);
xor XOR2 (N15707, N15706, N15416);
xor XOR2 (N15708, N15690, N4950);
or OR3 (N15709, N15705, N2996, N10863);
nor NOR3 (N15710, N15694, N14218, N14989);
nand NAND3 (N15711, N15704, N5676, N4401);
buf BUF1 (N15712, N15710);
nor NOR2 (N15713, N15712, N9810);
buf BUF1 (N15714, N15713);
or OR3 (N15715, N15711, N9711, N11478);
or OR2 (N15716, N15707, N11406);
buf BUF1 (N15717, N15703);
and AND3 (N15718, N15716, N15037, N7528);
nand NAND3 (N15719, N15679, N10098, N1804);
not NOT1 (N15720, N15719);
nand NAND3 (N15721, N15715, N13071, N14376);
or OR4 (N15722, N15708, N5458, N15093, N9839);
not NOT1 (N15723, N15718);
nor NOR3 (N15724, N15722, N6920, N2233);
nand NAND2 (N15725, N15701, N8289);
nand NAND2 (N15726, N15714, N2796);
xor XOR2 (N15727, N15709, N2311);
xor XOR2 (N15728, N15727, N2373);
and AND2 (N15729, N15721, N14165);
nor NOR4 (N15730, N15729, N13414, N7457, N7221);
not NOT1 (N15731, N15723);
xor XOR2 (N15732, N15702, N6263);
or OR2 (N15733, N15726, N790);
nand NAND2 (N15734, N15698, N10617);
xor XOR2 (N15735, N15734, N10408);
not NOT1 (N15736, N15720);
xor XOR2 (N15737, N15736, N491);
nor NOR3 (N15738, N15724, N6889, N6278);
not NOT1 (N15739, N15733);
or OR3 (N15740, N15732, N14865, N28);
xor XOR2 (N15741, N15728, N14458);
nand NAND2 (N15742, N15730, N14648);
and AND2 (N15743, N15739, N7144);
not NOT1 (N15744, N15735);
or OR3 (N15745, N15744, N3458, N14402);
not NOT1 (N15746, N15742);
and AND2 (N15747, N15745, N10891);
xor XOR2 (N15748, N15741, N14882);
not NOT1 (N15749, N15740);
xor XOR2 (N15750, N15738, N3323);
or OR3 (N15751, N15747, N3292, N1082);
buf BUF1 (N15752, N15749);
nand NAND4 (N15753, N15717, N10984, N9128, N1514);
or OR2 (N15754, N15731, N12559);
or OR4 (N15755, N15746, N6961, N11345, N12437);
nor NOR4 (N15756, N15743, N10549, N12567, N2278);
nor NOR3 (N15757, N15725, N1565, N3839);
buf BUF1 (N15758, N15751);
nor NOR2 (N15759, N15753, N13806);
nor NOR4 (N15760, N15748, N7606, N7600, N5155);
and AND3 (N15761, N15754, N1975, N137);
xor XOR2 (N15762, N15761, N3476);
xor XOR2 (N15763, N15758, N7707);
nor NOR3 (N15764, N15737, N12536, N4649);
buf BUF1 (N15765, N15764);
not NOT1 (N15766, N15756);
xor XOR2 (N15767, N15752, N8540);
and AND2 (N15768, N15760, N9234);
xor XOR2 (N15769, N15767, N12062);
xor XOR2 (N15770, N15763, N5386);
and AND3 (N15771, N15768, N8062, N8059);
buf BUF1 (N15772, N15765);
or OR3 (N15773, N15772, N10482, N4285);
nor NOR2 (N15774, N15755, N131);
xor XOR2 (N15775, N15762, N9756);
buf BUF1 (N15776, N15770);
or OR4 (N15777, N15775, N4189, N9725, N12773);
or OR4 (N15778, N15771, N4285, N2561, N162);
not NOT1 (N15779, N15778);
xor XOR2 (N15780, N15773, N908);
nor NOR2 (N15781, N15750, N80);
buf BUF1 (N15782, N15769);
not NOT1 (N15783, N15757);
or OR3 (N15784, N15779, N13252, N3798);
not NOT1 (N15785, N15766);
nor NOR2 (N15786, N15776, N5041);
nand NAND4 (N15787, N15782, N2303, N11423, N3817);
nor NOR2 (N15788, N15787, N8685);
buf BUF1 (N15789, N15783);
buf BUF1 (N15790, N15759);
nand NAND3 (N15791, N15790, N2050, N9478);
buf BUF1 (N15792, N15781);
nor NOR2 (N15793, N15777, N3542);
not NOT1 (N15794, N15774);
xor XOR2 (N15795, N15788, N980);
nor NOR2 (N15796, N15780, N12759);
xor XOR2 (N15797, N15792, N8031);
and AND2 (N15798, N15793, N6335);
not NOT1 (N15799, N15791);
xor XOR2 (N15800, N15796, N14959);
nand NAND3 (N15801, N15800, N9224, N10076);
and AND2 (N15802, N15784, N4049);
not NOT1 (N15803, N15794);
nor NOR3 (N15804, N15803, N15006, N14777);
buf BUF1 (N15805, N15786);
nor NOR2 (N15806, N15785, N4565);
or OR2 (N15807, N15799, N7253);
xor XOR2 (N15808, N15802, N8954);
buf BUF1 (N15809, N15797);
and AND3 (N15810, N15808, N2965, N7307);
buf BUF1 (N15811, N15789);
xor XOR2 (N15812, N15805, N3177);
or OR2 (N15813, N15812, N3552);
or OR2 (N15814, N15806, N12877);
nand NAND2 (N15815, N15813, N13411);
xor XOR2 (N15816, N15804, N969);
xor XOR2 (N15817, N15811, N13564);
nor NOR3 (N15818, N15815, N7872, N13259);
or OR4 (N15819, N15795, N3799, N8573, N9806);
not NOT1 (N15820, N15807);
buf BUF1 (N15821, N15818);
nor NOR3 (N15822, N15816, N6618, N3515);
nor NOR4 (N15823, N15819, N7972, N15077, N9234);
or OR2 (N15824, N15809, N14550);
nor NOR3 (N15825, N15817, N14677, N5337);
or OR3 (N15826, N15822, N4058, N13697);
and AND4 (N15827, N15810, N15347, N13808, N14820);
xor XOR2 (N15828, N15824, N13021);
not NOT1 (N15829, N15828);
and AND3 (N15830, N15821, N6105, N6304);
not NOT1 (N15831, N15826);
nand NAND2 (N15832, N15801, N8942);
nand NAND2 (N15833, N15814, N11385);
nor NOR3 (N15834, N15832, N4989, N14475);
nand NAND2 (N15835, N15830, N1403);
and AND3 (N15836, N15831, N7322, N4950);
and AND2 (N15837, N15820, N3367);
nor NOR2 (N15838, N15834, N8216);
or OR4 (N15839, N15825, N603, N3517, N10794);
nand NAND2 (N15840, N15837, N4932);
buf BUF1 (N15841, N15833);
not NOT1 (N15842, N15827);
or OR4 (N15843, N15823, N4169, N11283, N6329);
not NOT1 (N15844, N15840);
nor NOR4 (N15845, N15836, N1619, N15570, N3408);
buf BUF1 (N15846, N15838);
or OR3 (N15847, N15841, N2372, N11391);
and AND3 (N15848, N15829, N14985, N9911);
not NOT1 (N15849, N15835);
nand NAND3 (N15850, N15848, N3725, N5228);
xor XOR2 (N15851, N15849, N7288);
nand NAND2 (N15852, N15851, N9043);
nor NOR4 (N15853, N15846, N5678, N5278, N15627);
xor XOR2 (N15854, N15845, N4734);
buf BUF1 (N15855, N15853);
nor NOR3 (N15856, N15854, N927, N6174);
buf BUF1 (N15857, N15844);
nand NAND2 (N15858, N15798, N1607);
and AND2 (N15859, N15847, N11731);
or OR4 (N15860, N15856, N7471, N7568, N11713);
and AND3 (N15861, N15843, N6915, N15028);
nand NAND2 (N15862, N15842, N6761);
xor XOR2 (N15863, N15859, N6442);
xor XOR2 (N15864, N15857, N14244);
buf BUF1 (N15865, N15855);
nand NAND4 (N15866, N15863, N8998, N15065, N11658);
xor XOR2 (N15867, N15862, N4485);
nor NOR3 (N15868, N15852, N1400, N15505);
nand NAND2 (N15869, N15866, N6066);
or OR3 (N15870, N15858, N6759, N14042);
buf BUF1 (N15871, N15870);
buf BUF1 (N15872, N15865);
nand NAND4 (N15873, N15869, N5981, N13958, N1192);
or OR4 (N15874, N15850, N6091, N8145, N14282);
nand NAND4 (N15875, N15860, N1570, N15286, N14992);
or OR3 (N15876, N15872, N2132, N13521);
buf BUF1 (N15877, N15875);
or OR2 (N15878, N15877, N1255);
not NOT1 (N15879, N15861);
buf BUF1 (N15880, N15878);
nand NAND4 (N15881, N15879, N10713, N1990, N3545);
not NOT1 (N15882, N15874);
not NOT1 (N15883, N15864);
buf BUF1 (N15884, N15881);
and AND4 (N15885, N15871, N6973, N12119, N14558);
xor XOR2 (N15886, N15839, N10457);
and AND4 (N15887, N15876, N4952, N13608, N10170);
buf BUF1 (N15888, N15883);
and AND4 (N15889, N15868, N12497, N8147, N5345);
buf BUF1 (N15890, N15886);
not NOT1 (N15891, N15884);
nor NOR4 (N15892, N15880, N11857, N10488, N7490);
xor XOR2 (N15893, N15885, N4690);
or OR4 (N15894, N15891, N8812, N792, N2103);
xor XOR2 (N15895, N15890, N6081);
or OR4 (N15896, N15888, N10393, N11234, N5915);
nor NOR2 (N15897, N15887, N12607);
not NOT1 (N15898, N15892);
nor NOR3 (N15899, N15894, N11922, N801);
xor XOR2 (N15900, N15898, N7487);
xor XOR2 (N15901, N15895, N6865);
nand NAND3 (N15902, N15899, N6934, N8998);
or OR3 (N15903, N15867, N9633, N6039);
xor XOR2 (N15904, N15873, N4369);
buf BUF1 (N15905, N15882);
or OR3 (N15906, N15896, N4714, N14022);
and AND2 (N15907, N15902, N7981);
nand NAND2 (N15908, N15901, N12917);
or OR4 (N15909, N15905, N11405, N9041, N11121);
nand NAND4 (N15910, N15903, N3598, N1096, N3049);
or OR2 (N15911, N15893, N2518);
and AND3 (N15912, N15910, N442, N15739);
and AND2 (N15913, N15889, N11597);
buf BUF1 (N15914, N15900);
not NOT1 (N15915, N15913);
nand NAND2 (N15916, N15911, N13495);
not NOT1 (N15917, N15912);
nand NAND4 (N15918, N15915, N11580, N10136, N7330);
nor NOR3 (N15919, N15897, N8568, N13207);
not NOT1 (N15920, N15914);
not NOT1 (N15921, N15904);
xor XOR2 (N15922, N15908, N4218);
xor XOR2 (N15923, N15922, N10687);
and AND4 (N15924, N15909, N1028, N10995, N337);
and AND2 (N15925, N15917, N13374);
nor NOR4 (N15926, N15921, N15330, N3448, N6088);
and AND3 (N15927, N15925, N284, N2447);
nor NOR4 (N15928, N15923, N5845, N1891, N9153);
nand NAND3 (N15929, N15906, N10445, N9361);
or OR2 (N15930, N15927, N5377);
buf BUF1 (N15931, N15928);
and AND3 (N15932, N15919, N2035, N339);
buf BUF1 (N15933, N15918);
buf BUF1 (N15934, N15920);
and AND4 (N15935, N15926, N10126, N2853, N4419);
nand NAND3 (N15936, N15932, N6891, N39);
or OR2 (N15937, N15935, N2647);
nand NAND4 (N15938, N15933, N15809, N7436, N9607);
or OR2 (N15939, N15930, N3632);
nand NAND4 (N15940, N15924, N8189, N11548, N15411);
not NOT1 (N15941, N15937);
nor NOR4 (N15942, N15929, N13580, N15306, N5001);
nor NOR2 (N15943, N15941, N13062);
and AND4 (N15944, N15934, N2806, N14582, N9617);
and AND3 (N15945, N15942, N7434, N10810);
and AND4 (N15946, N15939, N13646, N7447, N334);
or OR4 (N15947, N15938, N10513, N12207, N4067);
xor XOR2 (N15948, N15947, N12975);
not NOT1 (N15949, N15946);
buf BUF1 (N15950, N15949);
and AND3 (N15951, N15931, N4001, N1638);
nand NAND2 (N15952, N15943, N14833);
or OR2 (N15953, N15952, N4581);
nand NAND4 (N15954, N15944, N9472, N14126, N5207);
not NOT1 (N15955, N15948);
nor NOR3 (N15956, N15955, N11491, N1480);
nand NAND4 (N15957, N15950, N782, N12012, N5531);
buf BUF1 (N15958, N15936);
or OR3 (N15959, N15916, N6380, N12452);
and AND3 (N15960, N15907, N15630, N14335);
and AND2 (N15961, N15960, N12108);
and AND3 (N15962, N15958, N12953, N14372);
xor XOR2 (N15963, N15951, N7116);
not NOT1 (N15964, N15954);
xor XOR2 (N15965, N15962, N13685);
not NOT1 (N15966, N15940);
and AND3 (N15967, N15966, N6445, N6401);
xor XOR2 (N15968, N15953, N11452);
xor XOR2 (N15969, N15965, N3110);
nor NOR3 (N15970, N15957, N4217, N1458);
buf BUF1 (N15971, N15961);
not NOT1 (N15972, N15963);
xor XOR2 (N15973, N15968, N15570);
nand NAND4 (N15974, N15956, N11401, N2474, N14084);
nand NAND3 (N15975, N15964, N2246, N13551);
not NOT1 (N15976, N15974);
or OR4 (N15977, N15967, N7533, N15008, N14261);
nand NAND3 (N15978, N15975, N12161, N6276);
nand NAND4 (N15979, N15970, N1230, N4199, N7371);
or OR3 (N15980, N15973, N10090, N4917);
nor NOR2 (N15981, N15979, N15509);
or OR2 (N15982, N15972, N9903);
not NOT1 (N15983, N15971);
not NOT1 (N15984, N15969);
nor NOR4 (N15985, N15945, N8806, N9541, N15234);
nor NOR4 (N15986, N15977, N11609, N3035, N2413);
and AND3 (N15987, N15983, N2437, N12015);
xor XOR2 (N15988, N15982, N6930);
or OR3 (N15989, N15976, N3813, N7191);
nor NOR3 (N15990, N15987, N14521, N8495);
xor XOR2 (N15991, N15978, N3922);
and AND2 (N15992, N15959, N23);
and AND2 (N15993, N15989, N9454);
and AND3 (N15994, N15988, N12527, N12470);
buf BUF1 (N15995, N15984);
or OR3 (N15996, N15993, N6758, N925);
buf BUF1 (N15997, N15994);
xor XOR2 (N15998, N15985, N10406);
xor XOR2 (N15999, N15997, N6201);
nor NOR2 (N16000, N15990, N3596);
xor XOR2 (N16001, N15996, N8112);
nand NAND3 (N16002, N15980, N5254, N1777);
and AND2 (N16003, N15998, N11113);
nor NOR3 (N16004, N16001, N6098, N2909);
not NOT1 (N16005, N16002);
xor XOR2 (N16006, N16000, N11675);
xor XOR2 (N16007, N16003, N9052);
nand NAND2 (N16008, N15995, N4639);
not NOT1 (N16009, N15999);
and AND2 (N16010, N15992, N7543);
nor NOR2 (N16011, N16004, N9265);
nand NAND4 (N16012, N16008, N1831, N2265, N12462);
and AND3 (N16013, N16007, N11457, N6566);
xor XOR2 (N16014, N16010, N2586);
buf BUF1 (N16015, N15991);
buf BUF1 (N16016, N15986);
endmodule