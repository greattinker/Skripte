// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23;

output N12821,N12815,N12818,N12813,N12781,N12814,N12820,N12822,N12819,N12823;

or OR2 (N24, N12, N19);
buf BUF1 (N25, N14);
xor XOR2 (N26, N21, N25);
xor XOR2 (N27, N14, N8);
or OR3 (N28, N22, N14, N1);
buf BUF1 (N29, N5);
nor NOR4 (N30, N4, N8, N2, N6);
xor XOR2 (N31, N22, N8);
not NOT1 (N32, N1);
not NOT1 (N33, N3);
or OR3 (N34, N30, N24, N9);
or OR2 (N35, N16, N3);
xor XOR2 (N36, N30, N11);
xor XOR2 (N37, N28, N25);
or OR3 (N38, N29, N10, N17);
or OR4 (N39, N36, N13, N20, N17);
buf BUF1 (N40, N38);
nor NOR2 (N41, N35, N8);
or OR2 (N42, N40, N20);
xor XOR2 (N43, N32, N15);
or OR3 (N44, N31, N15, N23);
not NOT1 (N45, N33);
not NOT1 (N46, N37);
xor XOR2 (N47, N45, N39);
or OR4 (N48, N44, N5, N16, N28);
nand NAND4 (N49, N35, N31, N29, N1);
not NOT1 (N50, N27);
or OR3 (N51, N34, N16, N21);
not NOT1 (N52, N51);
nor NOR4 (N53, N46, N18, N30, N52);
xor XOR2 (N54, N9, N13);
nor NOR4 (N55, N41, N52, N16, N2);
and AND2 (N56, N54, N53);
nand NAND2 (N57, N49, N16);
or OR4 (N58, N21, N43, N17, N4);
nand NAND2 (N59, N43, N3);
xor XOR2 (N60, N59, N6);
xor XOR2 (N61, N47, N28);
and AND4 (N62, N61, N32, N30, N35);
and AND3 (N63, N62, N43, N34);
nor NOR2 (N64, N60, N34);
nor NOR4 (N65, N56, N32, N11, N18);
nand NAND3 (N66, N57, N57, N45);
not NOT1 (N67, N58);
nand NAND3 (N68, N55, N15, N61);
buf BUF1 (N69, N26);
nor NOR2 (N70, N50, N62);
nor NOR3 (N71, N64, N20, N41);
and AND3 (N72, N42, N64, N2);
nor NOR2 (N73, N67, N1);
or OR4 (N74, N72, N22, N55, N11);
nand NAND4 (N75, N73, N1, N62, N74);
and AND3 (N76, N66, N21, N48);
and AND3 (N77, N3, N30, N17);
xor XOR2 (N78, N31, N1);
not NOT1 (N79, N78);
or OR2 (N80, N69, N10);
buf BUF1 (N81, N63);
nor NOR3 (N82, N65, N41, N71);
nand NAND3 (N83, N64, N18, N22);
and AND3 (N84, N77, N30, N39);
or OR2 (N85, N80, N18);
buf BUF1 (N86, N70);
xor XOR2 (N87, N81, N71);
or OR3 (N88, N75, N51, N18);
not NOT1 (N89, N85);
or OR4 (N90, N83, N85, N31, N72);
and AND3 (N91, N88, N20, N20);
xor XOR2 (N92, N86, N46);
or OR4 (N93, N82, N49, N70, N83);
or OR3 (N94, N68, N71, N3);
nand NAND4 (N95, N94, N65, N94, N29);
not NOT1 (N96, N79);
not NOT1 (N97, N91);
buf BUF1 (N98, N87);
or OR2 (N99, N97, N50);
not NOT1 (N100, N95);
nand NAND4 (N101, N98, N62, N3, N27);
nand NAND3 (N102, N93, N33, N42);
xor XOR2 (N103, N92, N47);
buf BUF1 (N104, N101);
buf BUF1 (N105, N102);
not NOT1 (N106, N100);
and AND3 (N107, N96, N13, N2);
nor NOR2 (N108, N84, N80);
nand NAND3 (N109, N105, N71, N43);
nor NOR3 (N110, N103, N33, N75);
and AND2 (N111, N107, N10);
and AND3 (N112, N76, N111, N5);
not NOT1 (N113, N89);
not NOT1 (N114, N89);
or OR2 (N115, N99, N104);
and AND4 (N116, N27, N82, N95, N41);
xor XOR2 (N117, N114, N53);
and AND4 (N118, N106, N77, N111, N106);
or OR2 (N119, N108, N10);
buf BUF1 (N120, N116);
buf BUF1 (N121, N117);
xor XOR2 (N122, N119, N96);
not NOT1 (N123, N122);
not NOT1 (N124, N110);
nand NAND2 (N125, N115, N60);
nand NAND2 (N126, N124, N83);
xor XOR2 (N127, N123, N36);
nand NAND4 (N128, N127, N119, N124, N75);
xor XOR2 (N129, N128, N4);
nor NOR3 (N130, N118, N73, N13);
not NOT1 (N131, N125);
nor NOR3 (N132, N120, N102, N79);
nor NOR2 (N133, N131, N80);
buf BUF1 (N134, N109);
xor XOR2 (N135, N129, N96);
and AND4 (N136, N126, N102, N101, N115);
not NOT1 (N137, N90);
or OR4 (N138, N121, N80, N16, N4);
not NOT1 (N139, N135);
not NOT1 (N140, N133);
nor NOR4 (N141, N113, N8, N113, N60);
not NOT1 (N142, N130);
buf BUF1 (N143, N132);
xor XOR2 (N144, N136, N134);
xor XOR2 (N145, N130, N130);
not NOT1 (N146, N139);
nand NAND3 (N147, N144, N144, N38);
xor XOR2 (N148, N145, N18);
buf BUF1 (N149, N148);
nor NOR3 (N150, N147, N108, N50);
nor NOR4 (N151, N140, N16, N4, N122);
not NOT1 (N152, N143);
not NOT1 (N153, N149);
or OR4 (N154, N138, N113, N96, N63);
not NOT1 (N155, N112);
xor XOR2 (N156, N142, N121);
nor NOR4 (N157, N156, N97, N40, N72);
xor XOR2 (N158, N153, N52);
buf BUF1 (N159, N158);
xor XOR2 (N160, N154, N146);
xor XOR2 (N161, N119, N133);
not NOT1 (N162, N161);
not NOT1 (N163, N157);
nand NAND3 (N164, N152, N55, N25);
buf BUF1 (N165, N155);
nand NAND2 (N166, N164, N72);
xor XOR2 (N167, N141, N122);
not NOT1 (N168, N167);
xor XOR2 (N169, N159, N105);
nor NOR2 (N170, N163, N135);
nand NAND2 (N171, N168, N50);
nor NOR2 (N172, N151, N41);
nor NOR2 (N173, N172, N95);
or OR2 (N174, N162, N168);
nor NOR3 (N175, N166, N35, N161);
buf BUF1 (N176, N174);
nor NOR3 (N177, N171, N13, N141);
and AND2 (N178, N160, N106);
nor NOR4 (N179, N177, N97, N32, N107);
nand NAND2 (N180, N176, N59);
buf BUF1 (N181, N150);
or OR3 (N182, N170, N149, N19);
buf BUF1 (N183, N175);
nor NOR3 (N184, N179, N84, N144);
and AND2 (N185, N181, N31);
and AND4 (N186, N184, N48, N47, N89);
xor XOR2 (N187, N178, N109);
or OR3 (N188, N185, N88, N62);
buf BUF1 (N189, N180);
nor NOR3 (N190, N188, N35, N144);
nor NOR4 (N191, N183, N123, N134, N11);
or OR4 (N192, N191, N191, N162, N10);
nor NOR2 (N193, N169, N38);
or OR3 (N194, N190, N40, N183);
nand NAND3 (N195, N192, N47, N142);
nand NAND2 (N196, N173, N159);
and AND3 (N197, N165, N52, N89);
nand NAND3 (N198, N189, N17, N171);
xor XOR2 (N199, N193, N63);
nor NOR2 (N200, N199, N93);
nand NAND4 (N201, N187, N59, N150, N200);
xor XOR2 (N202, N3, N113);
nand NAND3 (N203, N186, N133, N110);
nor NOR3 (N204, N194, N48, N125);
not NOT1 (N205, N204);
not NOT1 (N206, N197);
nor NOR4 (N207, N201, N111, N106, N93);
xor XOR2 (N208, N206, N3);
not NOT1 (N209, N203);
xor XOR2 (N210, N196, N114);
xor XOR2 (N211, N198, N201);
and AND3 (N212, N195, N186, N28);
nand NAND2 (N213, N137, N210);
not NOT1 (N214, N191);
or OR2 (N215, N212, N133);
not NOT1 (N216, N215);
buf BUF1 (N217, N202);
xor XOR2 (N218, N213, N43);
not NOT1 (N219, N207);
or OR3 (N220, N209, N149, N187);
nor NOR2 (N221, N205, N53);
nor NOR3 (N222, N211, N143, N160);
or OR2 (N223, N218, N43);
nand NAND4 (N224, N216, N14, N190, N171);
not NOT1 (N225, N223);
xor XOR2 (N226, N214, N199);
nor NOR4 (N227, N222, N223, N179, N24);
nand NAND3 (N228, N221, N59, N109);
or OR3 (N229, N182, N130, N61);
nor NOR4 (N230, N225, N150, N172, N30);
xor XOR2 (N231, N230, N12);
nor NOR4 (N232, N224, N229, N158, N131);
nand NAND3 (N233, N86, N55, N213);
nand NAND4 (N234, N220, N114, N33, N214);
or OR3 (N235, N208, N191, N132);
nor NOR3 (N236, N219, N59, N36);
nand NAND3 (N237, N233, N35, N6);
buf BUF1 (N238, N227);
or OR4 (N239, N232, N69, N55, N137);
and AND2 (N240, N236, N43);
xor XOR2 (N241, N228, N8);
buf BUF1 (N242, N241);
xor XOR2 (N243, N217, N88);
xor XOR2 (N244, N226, N85);
xor XOR2 (N245, N231, N44);
nand NAND2 (N246, N238, N14);
or OR4 (N247, N239, N59, N227, N146);
nand NAND2 (N248, N237, N104);
buf BUF1 (N249, N234);
nor NOR2 (N250, N245, N174);
not NOT1 (N251, N247);
nand NAND3 (N252, N248, N198, N12);
buf BUF1 (N253, N249);
nand NAND2 (N254, N242, N29);
buf BUF1 (N255, N246);
nand NAND3 (N256, N250, N54, N251);
or OR2 (N257, N24, N210);
or OR2 (N258, N257, N38);
not NOT1 (N259, N240);
buf BUF1 (N260, N253);
buf BUF1 (N261, N244);
nand NAND2 (N262, N260, N155);
nor NOR3 (N263, N256, N195, N123);
and AND3 (N264, N261, N44, N162);
nor NOR4 (N265, N243, N153, N135, N166);
and AND2 (N266, N262, N43);
not NOT1 (N267, N235);
nor NOR4 (N268, N252, N136, N45, N34);
and AND4 (N269, N258, N179, N213, N79);
xor XOR2 (N270, N254, N230);
and AND4 (N271, N268, N196, N267, N191);
nand NAND4 (N272, N107, N20, N176, N33);
not NOT1 (N273, N259);
nand NAND2 (N274, N266, N57);
nand NAND3 (N275, N274, N146, N225);
nor NOR4 (N276, N275, N259, N212, N138);
buf BUF1 (N277, N271);
buf BUF1 (N278, N265);
or OR3 (N279, N263, N160, N278);
nand NAND3 (N280, N149, N153, N132);
nand NAND3 (N281, N279, N153, N126);
nand NAND3 (N282, N272, N221, N98);
nand NAND2 (N283, N273, N96);
nand NAND3 (N284, N277, N171, N24);
buf BUF1 (N285, N264);
nand NAND3 (N286, N285, N38, N196);
nand NAND4 (N287, N280, N257, N162, N116);
nor NOR2 (N288, N269, N64);
not NOT1 (N289, N281);
nand NAND2 (N290, N276, N222);
and AND2 (N291, N284, N29);
nor NOR3 (N292, N288, N245, N259);
not NOT1 (N293, N286);
nand NAND2 (N294, N283, N7);
and AND3 (N295, N291, N116, N65);
buf BUF1 (N296, N293);
buf BUF1 (N297, N290);
or OR3 (N298, N270, N70, N9);
buf BUF1 (N299, N298);
nand NAND2 (N300, N289, N181);
nand NAND4 (N301, N255, N60, N279, N285);
and AND2 (N302, N295, N96);
nor NOR2 (N303, N302, N14);
nand NAND2 (N304, N294, N25);
nor NOR2 (N305, N287, N62);
and AND4 (N306, N299, N113, N232, N130);
xor XOR2 (N307, N303, N9);
nor NOR4 (N308, N307, N253, N159, N59);
xor XOR2 (N309, N306, N277);
buf BUF1 (N310, N296);
and AND4 (N311, N300, N304, N42, N107);
buf BUF1 (N312, N132);
buf BUF1 (N313, N310);
nand NAND3 (N314, N311, N53, N104);
nor NOR3 (N315, N313, N156, N216);
xor XOR2 (N316, N282, N305);
or OR4 (N317, N104, N58, N127, N57);
nor NOR4 (N318, N301, N54, N195, N109);
or OR4 (N319, N312, N91, N259, N205);
nor NOR3 (N320, N309, N257, N15);
and AND2 (N321, N314, N164);
not NOT1 (N322, N321);
not NOT1 (N323, N308);
or OR4 (N324, N316, N78, N176, N177);
nor NOR2 (N325, N318, N199);
nor NOR2 (N326, N319, N210);
not NOT1 (N327, N297);
xor XOR2 (N328, N324, N84);
or OR2 (N329, N328, N288);
not NOT1 (N330, N317);
nor NOR4 (N331, N315, N16, N313, N262);
buf BUF1 (N332, N329);
and AND3 (N333, N323, N159, N140);
and AND4 (N334, N326, N66, N298, N34);
and AND2 (N335, N327, N17);
buf BUF1 (N336, N335);
not NOT1 (N337, N334);
and AND2 (N338, N292, N319);
not NOT1 (N339, N338);
buf BUF1 (N340, N322);
nor NOR3 (N341, N332, N176, N150);
xor XOR2 (N342, N330, N56);
xor XOR2 (N343, N341, N143);
buf BUF1 (N344, N342);
xor XOR2 (N345, N339, N260);
nor NOR3 (N346, N333, N165, N275);
or OR4 (N347, N320, N22, N244, N84);
or OR4 (N348, N347, N246, N194, N268);
and AND3 (N349, N325, N235, N114);
and AND3 (N350, N349, N66, N253);
or OR4 (N351, N346, N12, N203, N317);
nand NAND4 (N352, N344, N299, N324, N335);
not NOT1 (N353, N331);
nand NAND2 (N354, N340, N229);
and AND3 (N355, N337, N202, N208);
nor NOR3 (N356, N351, N342, N324);
buf BUF1 (N357, N353);
or OR4 (N358, N352, N47, N209, N2);
xor XOR2 (N359, N348, N6);
buf BUF1 (N360, N343);
not NOT1 (N361, N355);
not NOT1 (N362, N356);
and AND2 (N363, N350, N178);
or OR4 (N364, N358, N226, N237, N217);
buf BUF1 (N365, N354);
nor NOR2 (N366, N357, N117);
buf BUF1 (N367, N366);
buf BUF1 (N368, N345);
not NOT1 (N369, N365);
not NOT1 (N370, N368);
or OR3 (N371, N361, N54, N103);
and AND2 (N372, N370, N298);
nor NOR2 (N373, N359, N139);
not NOT1 (N374, N371);
nand NAND3 (N375, N372, N52, N36);
or OR3 (N376, N369, N176, N320);
and AND3 (N377, N360, N47, N163);
xor XOR2 (N378, N373, N117);
nand NAND2 (N379, N364, N29);
xor XOR2 (N380, N336, N331);
not NOT1 (N381, N380);
nor NOR2 (N382, N377, N18);
xor XOR2 (N383, N367, N159);
buf BUF1 (N384, N375);
nand NAND2 (N385, N363, N17);
nand NAND4 (N386, N384, N43, N364, N97);
and AND3 (N387, N378, N237, N242);
buf BUF1 (N388, N386);
nand NAND2 (N389, N383, N74);
or OR3 (N390, N374, N218, N247);
buf BUF1 (N391, N389);
not NOT1 (N392, N376);
buf BUF1 (N393, N392);
buf BUF1 (N394, N362);
nor NOR2 (N395, N391, N197);
xor XOR2 (N396, N390, N234);
and AND4 (N397, N388, N30, N366, N132);
nand NAND4 (N398, N396, N4, N204, N180);
buf BUF1 (N399, N382);
or OR2 (N400, N379, N110);
nor NOR3 (N401, N394, N370, N87);
xor XOR2 (N402, N399, N88);
xor XOR2 (N403, N387, N318);
xor XOR2 (N404, N398, N137);
nand NAND2 (N405, N400, N79);
or OR4 (N406, N404, N263, N111, N132);
and AND3 (N407, N395, N13, N138);
buf BUF1 (N408, N397);
buf BUF1 (N409, N381);
buf BUF1 (N410, N409);
xor XOR2 (N411, N402, N122);
not NOT1 (N412, N385);
and AND4 (N413, N406, N351, N181, N83);
not NOT1 (N414, N408);
xor XOR2 (N415, N411, N322);
nor NOR2 (N416, N410, N400);
nor NOR2 (N417, N415, N129);
buf BUF1 (N418, N413);
or OR3 (N419, N407, N21, N289);
or OR4 (N420, N419, N73, N240, N238);
or OR4 (N421, N401, N16, N42, N360);
nor NOR2 (N422, N420, N7);
or OR2 (N423, N393, N65);
or OR3 (N424, N416, N366, N278);
or OR2 (N425, N412, N93);
xor XOR2 (N426, N422, N151);
nor NOR2 (N427, N425, N337);
and AND3 (N428, N417, N170, N290);
buf BUF1 (N429, N403);
and AND3 (N430, N424, N429, N321);
nor NOR3 (N431, N75, N58, N415);
or OR3 (N432, N427, N211, N429);
nor NOR3 (N433, N423, N322, N27);
buf BUF1 (N434, N433);
and AND4 (N435, N434, N324, N184, N399);
nor NOR4 (N436, N414, N10, N305, N5);
not NOT1 (N437, N421);
nor NOR3 (N438, N405, N197, N280);
nand NAND3 (N439, N432, N8, N364);
and AND3 (N440, N437, N163, N182);
not NOT1 (N441, N428);
and AND3 (N442, N436, N170, N419);
or OR3 (N443, N435, N72, N106);
buf BUF1 (N444, N439);
buf BUF1 (N445, N438);
nor NOR4 (N446, N418, N139, N293, N397);
xor XOR2 (N447, N443, N174);
not NOT1 (N448, N430);
nor NOR2 (N449, N446, N62);
xor XOR2 (N450, N440, N198);
nand NAND2 (N451, N426, N449);
or OR3 (N452, N104, N126, N255);
xor XOR2 (N453, N448, N327);
nand NAND2 (N454, N431, N289);
or OR2 (N455, N451, N219);
or OR4 (N456, N447, N396, N256, N241);
not NOT1 (N457, N450);
nand NAND4 (N458, N444, N106, N414, N276);
or OR3 (N459, N452, N420, N238);
nor NOR2 (N460, N455, N410);
nor NOR2 (N461, N453, N361);
nor NOR4 (N462, N459, N60, N184, N415);
buf BUF1 (N463, N462);
nor NOR3 (N464, N457, N62, N401);
or OR4 (N465, N460, N184, N29, N181);
or OR4 (N466, N454, N285, N10, N279);
nand NAND4 (N467, N461, N140, N52, N175);
nor NOR4 (N468, N456, N5, N101, N402);
not NOT1 (N469, N441);
nor NOR3 (N470, N468, N33, N91);
nor NOR2 (N471, N445, N201);
nor NOR2 (N472, N467, N218);
nor NOR3 (N473, N472, N112, N468);
nor NOR4 (N474, N464, N115, N277, N259);
xor XOR2 (N475, N473, N144);
and AND3 (N476, N463, N239, N201);
nor NOR4 (N477, N474, N355, N298, N9);
or OR4 (N478, N477, N304, N432, N214);
nand NAND2 (N479, N465, N75);
buf BUF1 (N480, N458);
nand NAND2 (N481, N478, N96);
or OR2 (N482, N476, N384);
or OR2 (N483, N469, N225);
not NOT1 (N484, N481);
nand NAND3 (N485, N475, N438, N271);
or OR3 (N486, N483, N332, N311);
nand NAND2 (N487, N485, N160);
or OR3 (N488, N484, N465, N102);
or OR4 (N489, N482, N346, N440, N461);
and AND2 (N490, N470, N143);
nor NOR4 (N491, N490, N469, N269, N415);
buf BUF1 (N492, N471);
or OR4 (N493, N466, N327, N409, N32);
buf BUF1 (N494, N487);
xor XOR2 (N495, N494, N305);
not NOT1 (N496, N488);
buf BUF1 (N497, N489);
nor NOR3 (N498, N479, N147, N497);
not NOT1 (N499, N59);
or OR4 (N500, N498, N298, N279, N314);
nor NOR2 (N501, N492, N59);
xor XOR2 (N502, N496, N372);
or OR4 (N503, N495, N428, N486, N49);
nand NAND4 (N504, N473, N213, N5, N408);
or OR3 (N505, N442, N317, N448);
nand NAND4 (N506, N502, N340, N354, N138);
nand NAND3 (N507, N493, N6, N443);
buf BUF1 (N508, N500);
buf BUF1 (N509, N501);
and AND3 (N510, N499, N491, N29);
xor XOR2 (N511, N443, N301);
buf BUF1 (N512, N480);
and AND2 (N513, N504, N214);
xor XOR2 (N514, N507, N457);
and AND2 (N515, N510, N431);
nand NAND2 (N516, N512, N404);
not NOT1 (N517, N516);
nand NAND2 (N518, N514, N95);
xor XOR2 (N519, N505, N191);
not NOT1 (N520, N517);
not NOT1 (N521, N520);
nand NAND2 (N522, N508, N504);
and AND4 (N523, N519, N364, N157, N380);
nand NAND3 (N524, N522, N103, N373);
nand NAND3 (N525, N518, N128, N428);
or OR3 (N526, N513, N363, N241);
or OR3 (N527, N511, N515, N302);
and AND3 (N528, N15, N442, N423);
buf BUF1 (N529, N524);
or OR2 (N530, N525, N89);
nand NAND3 (N531, N506, N401, N234);
nand NAND3 (N532, N521, N24, N219);
buf BUF1 (N533, N529);
nand NAND3 (N534, N526, N126, N171);
nor NOR3 (N535, N523, N92, N385);
xor XOR2 (N536, N531, N232);
or OR4 (N537, N530, N254, N81, N237);
nor NOR4 (N538, N527, N365, N428, N266);
or OR3 (N539, N535, N368, N143);
buf BUF1 (N540, N528);
not NOT1 (N541, N540);
or OR4 (N542, N534, N246, N294, N278);
not NOT1 (N543, N542);
nor NOR4 (N544, N543, N34, N146, N540);
nand NAND2 (N545, N538, N436);
nand NAND2 (N546, N537, N432);
and AND2 (N547, N536, N286);
buf BUF1 (N548, N509);
nand NAND3 (N549, N539, N345, N476);
not NOT1 (N550, N549);
and AND4 (N551, N548, N95, N17, N208);
or OR3 (N552, N550, N47, N49);
or OR2 (N553, N503, N283);
and AND2 (N554, N551, N27);
xor XOR2 (N555, N552, N503);
not NOT1 (N556, N541);
nand NAND2 (N557, N544, N488);
or OR4 (N558, N545, N422, N292, N94);
nor NOR4 (N559, N554, N16, N473, N117);
nor NOR3 (N560, N547, N290, N47);
xor XOR2 (N561, N557, N438);
not NOT1 (N562, N561);
or OR4 (N563, N532, N328, N149, N263);
nor NOR4 (N564, N559, N416, N419, N441);
not NOT1 (N565, N564);
and AND3 (N566, N565, N433, N526);
xor XOR2 (N567, N533, N55);
nor NOR3 (N568, N558, N242, N26);
buf BUF1 (N569, N553);
nand NAND3 (N570, N568, N465, N43);
and AND4 (N571, N566, N406, N58, N202);
and AND4 (N572, N556, N32, N521, N272);
xor XOR2 (N573, N567, N109);
and AND4 (N574, N572, N243, N142, N104);
and AND2 (N575, N555, N371);
or OR3 (N576, N570, N448, N370);
or OR2 (N577, N571, N131);
nor NOR2 (N578, N560, N47);
buf BUF1 (N579, N563);
or OR3 (N580, N579, N412, N560);
and AND4 (N581, N562, N557, N117, N426);
and AND2 (N582, N546, N344);
buf BUF1 (N583, N576);
nor NOR3 (N584, N578, N68, N549);
buf BUF1 (N585, N577);
xor XOR2 (N586, N583, N329);
and AND2 (N587, N585, N300);
or OR2 (N588, N573, N509);
not NOT1 (N589, N575);
nor NOR4 (N590, N584, N489, N376, N326);
and AND3 (N591, N569, N197, N93);
not NOT1 (N592, N581);
and AND2 (N593, N582, N391);
xor XOR2 (N594, N574, N247);
nor NOR4 (N595, N594, N442, N22, N281);
not NOT1 (N596, N589);
nand NAND3 (N597, N587, N173, N156);
nand NAND2 (N598, N590, N497);
nor NOR3 (N599, N588, N311, N554);
xor XOR2 (N600, N580, N105);
nand NAND3 (N601, N600, N12, N237);
not NOT1 (N602, N599);
nor NOR2 (N603, N596, N3);
nor NOR3 (N604, N601, N299, N520);
nand NAND3 (N605, N586, N378, N237);
nor NOR3 (N606, N592, N109, N434);
nor NOR2 (N607, N598, N273);
nand NAND4 (N608, N602, N445, N208, N382);
not NOT1 (N609, N605);
nand NAND4 (N610, N609, N309, N135, N390);
nand NAND2 (N611, N597, N507);
buf BUF1 (N612, N607);
not NOT1 (N613, N611);
and AND3 (N614, N591, N439, N482);
and AND4 (N615, N604, N214, N83, N299);
nand NAND2 (N616, N603, N282);
nand NAND3 (N617, N616, N372, N301);
xor XOR2 (N618, N595, N142);
buf BUF1 (N619, N610);
xor XOR2 (N620, N619, N256);
nor NOR4 (N621, N614, N465, N614, N498);
nand NAND3 (N622, N620, N218, N262);
xor XOR2 (N623, N621, N467);
xor XOR2 (N624, N623, N239);
nor NOR3 (N625, N617, N574, N569);
nor NOR2 (N626, N625, N240);
and AND3 (N627, N626, N8, N271);
xor XOR2 (N628, N615, N260);
nor NOR3 (N629, N613, N4, N30);
buf BUF1 (N630, N593);
and AND3 (N631, N627, N511, N498);
or OR4 (N632, N612, N223, N94, N113);
not NOT1 (N633, N624);
and AND4 (N634, N629, N609, N11, N317);
and AND4 (N635, N606, N381, N89, N225);
buf BUF1 (N636, N635);
nand NAND4 (N637, N608, N255, N51, N399);
buf BUF1 (N638, N637);
or OR2 (N639, N638, N40);
xor XOR2 (N640, N636, N220);
xor XOR2 (N641, N630, N3);
buf BUF1 (N642, N618);
nor NOR2 (N643, N633, N31);
nor NOR4 (N644, N639, N403, N402, N95);
not NOT1 (N645, N631);
nand NAND4 (N646, N640, N109, N148, N368);
nand NAND4 (N647, N646, N591, N460, N361);
or OR4 (N648, N632, N234, N466, N441);
nor NOR4 (N649, N648, N22, N162, N473);
nor NOR4 (N650, N643, N403, N645, N339);
nor NOR4 (N651, N190, N316, N202, N26);
or OR3 (N652, N628, N288, N61);
nor NOR3 (N653, N642, N546, N419);
and AND4 (N654, N634, N344, N566, N447);
nor NOR4 (N655, N622, N10, N393, N258);
or OR4 (N656, N655, N382, N140, N216);
or OR2 (N657, N649, N467);
xor XOR2 (N658, N654, N445);
nand NAND3 (N659, N647, N216, N373);
not NOT1 (N660, N657);
nor NOR2 (N661, N656, N243);
nand NAND3 (N662, N659, N133, N234);
or OR2 (N663, N644, N411);
xor XOR2 (N664, N662, N392);
nand NAND3 (N665, N658, N654, N566);
or OR4 (N666, N661, N585, N564, N342);
not NOT1 (N667, N666);
or OR2 (N668, N650, N554);
and AND3 (N669, N667, N516, N83);
and AND3 (N670, N641, N329, N661);
and AND4 (N671, N669, N501, N320, N497);
not NOT1 (N672, N665);
or OR4 (N673, N670, N140, N591, N324);
nand NAND2 (N674, N664, N75);
xor XOR2 (N675, N663, N417);
buf BUF1 (N676, N652);
or OR4 (N677, N672, N361, N449, N492);
nor NOR3 (N678, N674, N354, N184);
nor NOR4 (N679, N675, N614, N7, N1);
and AND3 (N680, N673, N137, N313);
xor XOR2 (N681, N680, N141);
or OR3 (N682, N668, N153, N301);
xor XOR2 (N683, N651, N103);
xor XOR2 (N684, N683, N39);
buf BUF1 (N685, N677);
nand NAND3 (N686, N676, N246, N463);
nor NOR2 (N687, N653, N168);
not NOT1 (N688, N686);
nor NOR3 (N689, N679, N137, N605);
or OR4 (N690, N660, N613, N328, N388);
buf BUF1 (N691, N671);
not NOT1 (N692, N688);
nor NOR3 (N693, N684, N314, N629);
or OR2 (N694, N693, N328);
not NOT1 (N695, N691);
nand NAND4 (N696, N692, N154, N188, N527);
not NOT1 (N697, N687);
xor XOR2 (N698, N681, N262);
nor NOR3 (N699, N678, N407, N277);
or OR3 (N700, N690, N439, N87);
and AND3 (N701, N700, N459, N465);
and AND3 (N702, N699, N100, N173);
not NOT1 (N703, N701);
xor XOR2 (N704, N698, N509);
buf BUF1 (N705, N696);
xor XOR2 (N706, N703, N604);
nand NAND3 (N707, N685, N9, N683);
buf BUF1 (N708, N704);
nand NAND2 (N709, N705, N397);
xor XOR2 (N710, N709, N95);
and AND2 (N711, N694, N330);
nor NOR3 (N712, N682, N335, N167);
or OR3 (N713, N695, N432, N652);
and AND4 (N714, N689, N250, N437, N536);
nand NAND3 (N715, N706, N230, N608);
or OR3 (N716, N713, N499, N186);
xor XOR2 (N717, N707, N358);
nor NOR2 (N718, N702, N716);
nand NAND4 (N719, N199, N327, N184, N696);
or OR4 (N720, N719, N306, N322, N708);
xor XOR2 (N721, N278, N43);
or OR3 (N722, N710, N477, N611);
xor XOR2 (N723, N717, N77);
nand NAND3 (N724, N722, N674, N345);
nand NAND4 (N725, N718, N715, N707, N203);
or OR3 (N726, N302, N406, N567);
and AND2 (N727, N720, N313);
xor XOR2 (N728, N724, N324);
xor XOR2 (N729, N725, N355);
xor XOR2 (N730, N711, N31);
or OR2 (N731, N714, N518);
not NOT1 (N732, N712);
not NOT1 (N733, N729);
or OR4 (N734, N728, N53, N712, N158);
not NOT1 (N735, N721);
xor XOR2 (N736, N733, N418);
nor NOR2 (N737, N723, N481);
and AND3 (N738, N732, N192, N87);
xor XOR2 (N739, N730, N706);
and AND2 (N740, N727, N105);
and AND4 (N741, N737, N524, N30, N306);
not NOT1 (N742, N741);
nand NAND2 (N743, N726, N157);
or OR4 (N744, N740, N166, N712, N104);
nand NAND4 (N745, N739, N714, N548, N451);
nand NAND2 (N746, N734, N29);
buf BUF1 (N747, N738);
and AND4 (N748, N743, N332, N438, N457);
not NOT1 (N749, N744);
or OR3 (N750, N747, N711, N437);
and AND4 (N751, N736, N158, N721, N558);
xor XOR2 (N752, N750, N438);
or OR2 (N753, N749, N72);
xor XOR2 (N754, N735, N123);
nand NAND2 (N755, N746, N533);
xor XOR2 (N756, N752, N621);
and AND4 (N757, N745, N704, N698, N3);
xor XOR2 (N758, N751, N104);
xor XOR2 (N759, N748, N699);
and AND4 (N760, N757, N5, N317, N514);
not NOT1 (N761, N753);
nor NOR3 (N762, N731, N616, N657);
buf BUF1 (N763, N758);
nor NOR3 (N764, N742, N170, N334);
and AND4 (N765, N697, N650, N478, N641);
not NOT1 (N766, N764);
or OR3 (N767, N754, N649, N268);
not NOT1 (N768, N766);
xor XOR2 (N769, N756, N582);
buf BUF1 (N770, N761);
buf BUF1 (N771, N759);
not NOT1 (N772, N771);
buf BUF1 (N773, N768);
nand NAND2 (N774, N765, N67);
buf BUF1 (N775, N767);
and AND2 (N776, N775, N290);
nand NAND2 (N777, N774, N203);
or OR2 (N778, N769, N494);
buf BUF1 (N779, N762);
nand NAND2 (N780, N778, N478);
xor XOR2 (N781, N777, N535);
xor XOR2 (N782, N779, N401);
nand NAND3 (N783, N782, N596, N108);
buf BUF1 (N784, N776);
or OR2 (N785, N780, N622);
nor NOR2 (N786, N783, N259);
xor XOR2 (N787, N786, N3);
buf BUF1 (N788, N785);
buf BUF1 (N789, N760);
not NOT1 (N790, N787);
xor XOR2 (N791, N772, N521);
nand NAND4 (N792, N781, N730, N578, N568);
and AND2 (N793, N763, N676);
and AND2 (N794, N755, N645);
not NOT1 (N795, N793);
or OR4 (N796, N789, N515, N50, N97);
xor XOR2 (N797, N794, N178);
nor NOR4 (N798, N784, N202, N360, N501);
not NOT1 (N799, N796);
buf BUF1 (N800, N795);
or OR3 (N801, N800, N726, N217);
and AND4 (N802, N790, N446, N797, N224);
buf BUF1 (N803, N776);
buf BUF1 (N804, N802);
xor XOR2 (N805, N798, N107);
nor NOR2 (N806, N803, N553);
buf BUF1 (N807, N792);
nand NAND4 (N808, N805, N682, N417, N66);
not NOT1 (N809, N799);
or OR4 (N810, N788, N399, N182, N276);
buf BUF1 (N811, N770);
or OR3 (N812, N810, N237, N489);
and AND4 (N813, N807, N69, N615, N75);
buf BUF1 (N814, N791);
buf BUF1 (N815, N813);
xor XOR2 (N816, N773, N308);
and AND4 (N817, N804, N326, N128, N375);
not NOT1 (N818, N808);
and AND2 (N819, N816, N656);
xor XOR2 (N820, N811, N433);
nand NAND3 (N821, N820, N354, N455);
xor XOR2 (N822, N821, N94);
buf BUF1 (N823, N817);
xor XOR2 (N824, N818, N564);
xor XOR2 (N825, N823, N23);
or OR4 (N826, N824, N226, N608, N435);
buf BUF1 (N827, N812);
and AND2 (N828, N819, N262);
not NOT1 (N829, N828);
and AND3 (N830, N806, N785, N418);
and AND4 (N831, N829, N341, N689, N468);
not NOT1 (N832, N826);
or OR2 (N833, N825, N796);
and AND2 (N834, N822, N419);
or OR4 (N835, N831, N687, N280, N624);
or OR2 (N836, N833, N267);
nor NOR3 (N837, N809, N719, N678);
not NOT1 (N838, N815);
or OR4 (N839, N837, N620, N550, N486);
buf BUF1 (N840, N827);
nor NOR4 (N841, N839, N476, N484, N202);
and AND4 (N842, N830, N184, N568, N637);
or OR2 (N843, N842, N184);
not NOT1 (N844, N843);
xor XOR2 (N845, N814, N796);
nor NOR4 (N846, N801, N593, N701, N53);
nor NOR3 (N847, N844, N402, N619);
not NOT1 (N848, N840);
not NOT1 (N849, N841);
not NOT1 (N850, N838);
or OR4 (N851, N846, N317, N373, N389);
buf BUF1 (N852, N849);
xor XOR2 (N853, N851, N629);
nor NOR3 (N854, N853, N84, N361);
or OR3 (N855, N850, N493, N721);
xor XOR2 (N856, N832, N593);
or OR2 (N857, N848, N285);
nor NOR2 (N858, N856, N7);
xor XOR2 (N859, N858, N520);
and AND3 (N860, N857, N121, N361);
nand NAND2 (N861, N852, N676);
nor NOR4 (N862, N836, N443, N491, N353);
or OR2 (N863, N855, N277);
not NOT1 (N864, N845);
not NOT1 (N865, N862);
xor XOR2 (N866, N861, N789);
nor NOR3 (N867, N864, N697, N265);
not NOT1 (N868, N854);
and AND3 (N869, N834, N453, N718);
nor NOR3 (N870, N835, N244, N769);
or OR3 (N871, N869, N99, N391);
nand NAND2 (N872, N859, N391);
not NOT1 (N873, N868);
buf BUF1 (N874, N865);
nand NAND4 (N875, N866, N311, N347, N716);
not NOT1 (N876, N871);
nand NAND4 (N877, N872, N70, N596, N105);
buf BUF1 (N878, N860);
nand NAND2 (N879, N870, N713);
buf BUF1 (N880, N878);
or OR4 (N881, N863, N549, N196, N312);
nor NOR2 (N882, N881, N669);
nand NAND3 (N883, N882, N112, N112);
nand NAND2 (N884, N867, N479);
not NOT1 (N885, N879);
nor NOR4 (N886, N875, N633, N818, N394);
and AND4 (N887, N883, N595, N1, N105);
nand NAND3 (N888, N877, N206, N34);
nand NAND4 (N889, N885, N228, N630, N500);
or OR2 (N890, N880, N610);
and AND2 (N891, N890, N213);
xor XOR2 (N892, N889, N801);
buf BUF1 (N893, N886);
nand NAND3 (N894, N873, N421, N716);
xor XOR2 (N895, N876, N104);
nor NOR4 (N896, N888, N405, N879, N420);
nand NAND2 (N897, N847, N145);
xor XOR2 (N898, N896, N344);
xor XOR2 (N899, N891, N117);
buf BUF1 (N900, N898);
or OR4 (N901, N897, N832, N110, N552);
or OR3 (N902, N892, N375, N901);
nand NAND2 (N903, N390, N308);
not NOT1 (N904, N902);
buf BUF1 (N905, N884);
buf BUF1 (N906, N887);
nand NAND2 (N907, N899, N768);
or OR3 (N908, N900, N183, N287);
not NOT1 (N909, N908);
buf BUF1 (N910, N874);
not NOT1 (N911, N895);
xor XOR2 (N912, N905, N222);
or OR4 (N913, N912, N524, N813, N625);
buf BUF1 (N914, N911);
nor NOR3 (N915, N914, N119, N90);
xor XOR2 (N916, N915, N247);
nand NAND2 (N917, N903, N534);
or OR3 (N918, N910, N95, N869);
nor NOR4 (N919, N907, N80, N726, N67);
buf BUF1 (N920, N909);
not NOT1 (N921, N906);
nand NAND3 (N922, N918, N116, N12);
or OR4 (N923, N921, N754, N203, N214);
nand NAND4 (N924, N893, N272, N215, N427);
or OR4 (N925, N924, N921, N669, N721);
xor XOR2 (N926, N917, N712);
not NOT1 (N927, N920);
or OR2 (N928, N919, N253);
and AND4 (N929, N926, N633, N831, N928);
buf BUF1 (N930, N376);
nor NOR4 (N931, N923, N654, N125, N813);
nand NAND4 (N932, N904, N46, N101, N664);
and AND3 (N933, N927, N560, N302);
or OR3 (N934, N931, N86, N576);
and AND3 (N935, N933, N579, N740);
nor NOR4 (N936, N929, N935, N746, N702);
xor XOR2 (N937, N178, N578);
not NOT1 (N938, N932);
nor NOR2 (N939, N938, N291);
xor XOR2 (N940, N936, N209);
buf BUF1 (N941, N934);
xor XOR2 (N942, N916, N145);
or OR3 (N943, N941, N511, N246);
not NOT1 (N944, N894);
or OR2 (N945, N942, N169);
not NOT1 (N946, N943);
and AND3 (N947, N925, N916, N646);
and AND2 (N948, N930, N247);
buf BUF1 (N949, N913);
not NOT1 (N950, N922);
nor NOR2 (N951, N945, N616);
not NOT1 (N952, N949);
and AND3 (N953, N950, N148, N933);
xor XOR2 (N954, N946, N916);
xor XOR2 (N955, N940, N456);
not NOT1 (N956, N947);
nand NAND4 (N957, N955, N28, N146, N533);
nor NOR2 (N958, N957, N190);
buf BUF1 (N959, N952);
buf BUF1 (N960, N954);
xor XOR2 (N961, N951, N568);
or OR3 (N962, N956, N909, N679);
xor XOR2 (N963, N937, N922);
xor XOR2 (N964, N962, N111);
nor NOR3 (N965, N939, N165, N309);
or OR3 (N966, N959, N530, N727);
nand NAND3 (N967, N966, N141, N514);
and AND3 (N968, N967, N780, N123);
not NOT1 (N969, N963);
nand NAND2 (N970, N969, N485);
xor XOR2 (N971, N965, N352);
xor XOR2 (N972, N958, N80);
or OR4 (N973, N970, N252, N176, N189);
and AND4 (N974, N968, N309, N439, N486);
nand NAND2 (N975, N944, N700);
xor XOR2 (N976, N973, N461);
nor NOR2 (N977, N974, N954);
xor XOR2 (N978, N960, N25);
buf BUF1 (N979, N978);
and AND3 (N980, N975, N761, N620);
not NOT1 (N981, N972);
and AND2 (N982, N971, N30);
buf BUF1 (N983, N977);
or OR4 (N984, N953, N275, N194, N90);
not NOT1 (N985, N964);
nor NOR2 (N986, N961, N6);
not NOT1 (N987, N980);
and AND3 (N988, N948, N486, N197);
nand NAND4 (N989, N984, N340, N607, N221);
nand NAND2 (N990, N989, N99);
xor XOR2 (N991, N982, N634);
buf BUF1 (N992, N983);
and AND3 (N993, N981, N631, N610);
nand NAND2 (N994, N979, N897);
and AND4 (N995, N987, N466, N615, N311);
nand NAND4 (N996, N992, N87, N201, N601);
buf BUF1 (N997, N986);
not NOT1 (N998, N995);
nor NOR4 (N999, N996, N845, N802, N975);
nor NOR4 (N1000, N997, N157, N568, N117);
and AND2 (N1001, N994, N557);
not NOT1 (N1002, N988);
xor XOR2 (N1003, N999, N272);
and AND2 (N1004, N991, N12);
buf BUF1 (N1005, N990);
nor NOR4 (N1006, N998, N934, N122, N122);
or OR4 (N1007, N993, N483, N47, N103);
and AND3 (N1008, N1002, N609, N190);
buf BUF1 (N1009, N1000);
not NOT1 (N1010, N1001);
nand NAND2 (N1011, N1007, N462);
buf BUF1 (N1012, N1008);
buf BUF1 (N1013, N1005);
not NOT1 (N1014, N1003);
or OR3 (N1015, N1009, N221, N154);
nor NOR4 (N1016, N1012, N191, N786, N485);
and AND4 (N1017, N1006, N378, N700, N791);
nand NAND2 (N1018, N1004, N232);
and AND2 (N1019, N976, N127);
and AND2 (N1020, N1016, N413);
and AND2 (N1021, N985, N716);
not NOT1 (N1022, N1010);
buf BUF1 (N1023, N1014);
nor NOR4 (N1024, N1021, N182, N161, N848);
buf BUF1 (N1025, N1017);
xor XOR2 (N1026, N1020, N236);
nor NOR2 (N1027, N1013, N1021);
or OR3 (N1028, N1026, N594, N970);
buf BUF1 (N1029, N1011);
xor XOR2 (N1030, N1024, N292);
buf BUF1 (N1031, N1029);
and AND2 (N1032, N1027, N736);
nand NAND2 (N1033, N1018, N829);
nand NAND2 (N1034, N1033, N1007);
nand NAND2 (N1035, N1028, N230);
not NOT1 (N1036, N1022);
not NOT1 (N1037, N1015);
nand NAND3 (N1038, N1019, N150, N883);
buf BUF1 (N1039, N1023);
or OR4 (N1040, N1025, N940, N709, N17);
not NOT1 (N1041, N1040);
and AND2 (N1042, N1031, N348);
not NOT1 (N1043, N1032);
buf BUF1 (N1044, N1041);
buf BUF1 (N1045, N1044);
nand NAND4 (N1046, N1034, N277, N126, N57);
and AND2 (N1047, N1038, N491);
nor NOR2 (N1048, N1047, N463);
xor XOR2 (N1049, N1036, N732);
not NOT1 (N1050, N1042);
and AND3 (N1051, N1039, N447, N499);
or OR2 (N1052, N1035, N921);
xor XOR2 (N1053, N1030, N96);
xor XOR2 (N1054, N1051, N639);
buf BUF1 (N1055, N1054);
nor NOR3 (N1056, N1046, N565, N307);
and AND3 (N1057, N1055, N760, N419);
not NOT1 (N1058, N1052);
nand NAND2 (N1059, N1049, N736);
and AND4 (N1060, N1057, N230, N986, N638);
buf BUF1 (N1061, N1058);
nor NOR2 (N1062, N1053, N851);
xor XOR2 (N1063, N1037, N289);
or OR3 (N1064, N1059, N972, N866);
xor XOR2 (N1065, N1061, N258);
or OR2 (N1066, N1056, N256);
nand NAND2 (N1067, N1043, N96);
nand NAND3 (N1068, N1067, N343, N520);
nor NOR4 (N1069, N1066, N842, N745, N236);
nor NOR2 (N1070, N1050, N470);
nand NAND3 (N1071, N1064, N442, N320);
nor NOR4 (N1072, N1069, N102, N714, N896);
buf BUF1 (N1073, N1065);
nor NOR3 (N1074, N1070, N831, N882);
and AND2 (N1075, N1045, N173);
nor NOR3 (N1076, N1073, N252, N484);
and AND4 (N1077, N1072, N754, N983, N256);
or OR2 (N1078, N1062, N213);
xor XOR2 (N1079, N1068, N188);
nand NAND2 (N1080, N1048, N258);
buf BUF1 (N1081, N1071);
xor XOR2 (N1082, N1074, N438);
and AND4 (N1083, N1079, N671, N936, N846);
buf BUF1 (N1084, N1077);
buf BUF1 (N1085, N1060);
xor XOR2 (N1086, N1063, N920);
xor XOR2 (N1087, N1078, N828);
not NOT1 (N1088, N1086);
xor XOR2 (N1089, N1085, N711);
or OR2 (N1090, N1088, N292);
xor XOR2 (N1091, N1076, N804);
and AND2 (N1092, N1083, N992);
nor NOR4 (N1093, N1075, N192, N891, N19);
xor XOR2 (N1094, N1091, N807);
or OR2 (N1095, N1090, N371);
and AND4 (N1096, N1084, N608, N13, N760);
xor XOR2 (N1097, N1096, N580);
not NOT1 (N1098, N1081);
xor XOR2 (N1099, N1094, N1097);
not NOT1 (N1100, N732);
nand NAND3 (N1101, N1087, N632, N693);
xor XOR2 (N1102, N1093, N310);
buf BUF1 (N1103, N1099);
or OR2 (N1104, N1095, N158);
or OR4 (N1105, N1102, N510, N681, N464);
buf BUF1 (N1106, N1105);
buf BUF1 (N1107, N1082);
nor NOR2 (N1108, N1092, N773);
and AND3 (N1109, N1103, N164, N611);
nand NAND3 (N1110, N1106, N526, N94);
buf BUF1 (N1111, N1107);
xor XOR2 (N1112, N1098, N697);
or OR3 (N1113, N1104, N19, N403);
or OR4 (N1114, N1080, N175, N344, N268);
buf BUF1 (N1115, N1112);
or OR4 (N1116, N1110, N1102, N505, N138);
nand NAND4 (N1117, N1115, N283, N934, N1081);
buf BUF1 (N1118, N1101);
buf BUF1 (N1119, N1100);
and AND3 (N1120, N1117, N682, N328);
nor NOR4 (N1121, N1120, N359, N537, N461);
and AND3 (N1122, N1116, N225, N760);
nor NOR4 (N1123, N1114, N1116, N536, N248);
not NOT1 (N1124, N1109);
buf BUF1 (N1125, N1111);
or OR3 (N1126, N1121, N293, N1027);
nor NOR4 (N1127, N1123, N413, N1024, N986);
xor XOR2 (N1128, N1108, N141);
nor NOR2 (N1129, N1125, N1018);
buf BUF1 (N1130, N1129);
or OR4 (N1131, N1122, N827, N360, N499);
not NOT1 (N1132, N1127);
xor XOR2 (N1133, N1089, N196);
not NOT1 (N1134, N1126);
and AND3 (N1135, N1133, N952, N550);
or OR2 (N1136, N1132, N169);
xor XOR2 (N1137, N1119, N185);
nand NAND3 (N1138, N1130, N24, N776);
nor NOR3 (N1139, N1131, N740, N808);
nand NAND4 (N1140, N1137, N989, N227, N729);
buf BUF1 (N1141, N1128);
nand NAND4 (N1142, N1136, N1046, N833, N1086);
not NOT1 (N1143, N1142);
xor XOR2 (N1144, N1124, N356);
nor NOR2 (N1145, N1134, N323);
buf BUF1 (N1146, N1140);
nand NAND3 (N1147, N1141, N327, N18);
and AND4 (N1148, N1147, N248, N1070, N164);
not NOT1 (N1149, N1146);
buf BUF1 (N1150, N1139);
and AND4 (N1151, N1148, N895, N44, N433);
buf BUF1 (N1152, N1144);
nand NAND2 (N1153, N1149, N681);
not NOT1 (N1154, N1145);
nor NOR3 (N1155, N1152, N307, N1120);
and AND4 (N1156, N1155, N207, N482, N726);
or OR2 (N1157, N1118, N81);
buf BUF1 (N1158, N1143);
buf BUF1 (N1159, N1138);
nand NAND4 (N1160, N1151, N281, N476, N542);
nor NOR3 (N1161, N1157, N224, N182);
nor NOR4 (N1162, N1159, N528, N942, N422);
xor XOR2 (N1163, N1156, N461);
or OR4 (N1164, N1158, N1142, N273, N664);
and AND2 (N1165, N1113, N472);
not NOT1 (N1166, N1164);
xor XOR2 (N1167, N1166, N378);
or OR3 (N1168, N1135, N525, N940);
xor XOR2 (N1169, N1153, N841);
not NOT1 (N1170, N1165);
not NOT1 (N1171, N1161);
or OR2 (N1172, N1168, N396);
xor XOR2 (N1173, N1169, N1114);
and AND3 (N1174, N1172, N986, N96);
xor XOR2 (N1175, N1173, N702);
nor NOR3 (N1176, N1150, N49, N362);
or OR4 (N1177, N1175, N549, N195, N363);
nand NAND3 (N1178, N1162, N569, N936);
and AND2 (N1179, N1154, N446);
nand NAND2 (N1180, N1167, N161);
nand NAND4 (N1181, N1177, N672, N552, N507);
nand NAND3 (N1182, N1178, N851, N1026);
not NOT1 (N1183, N1171);
xor XOR2 (N1184, N1183, N120);
not NOT1 (N1185, N1176);
buf BUF1 (N1186, N1179);
buf BUF1 (N1187, N1182);
and AND2 (N1188, N1185, N820);
nand NAND4 (N1189, N1187, N688, N335, N731);
nand NAND2 (N1190, N1188, N1158);
not NOT1 (N1191, N1163);
and AND3 (N1192, N1190, N382, N884);
xor XOR2 (N1193, N1186, N48);
xor XOR2 (N1194, N1160, N579);
not NOT1 (N1195, N1174);
and AND4 (N1196, N1189, N619, N267, N809);
buf BUF1 (N1197, N1180);
nand NAND3 (N1198, N1195, N312, N257);
and AND4 (N1199, N1170, N689, N169, N969);
nor NOR2 (N1200, N1197, N139);
not NOT1 (N1201, N1181);
not NOT1 (N1202, N1192);
nor NOR2 (N1203, N1201, N514);
xor XOR2 (N1204, N1199, N650);
xor XOR2 (N1205, N1203, N877);
not NOT1 (N1206, N1184);
buf BUF1 (N1207, N1194);
not NOT1 (N1208, N1193);
and AND4 (N1209, N1202, N582, N924, N660);
and AND3 (N1210, N1208, N63, N821);
nor NOR2 (N1211, N1200, N228);
buf BUF1 (N1212, N1209);
nor NOR2 (N1213, N1204, N976);
buf BUF1 (N1214, N1207);
buf BUF1 (N1215, N1191);
nor NOR4 (N1216, N1196, N75, N51, N1005);
or OR2 (N1217, N1198, N374);
or OR2 (N1218, N1216, N645);
and AND4 (N1219, N1210, N1076, N344, N143);
not NOT1 (N1220, N1218);
buf BUF1 (N1221, N1217);
and AND3 (N1222, N1219, N642, N60);
not NOT1 (N1223, N1211);
xor XOR2 (N1224, N1220, N165);
nor NOR2 (N1225, N1221, N272);
and AND4 (N1226, N1223, N679, N174, N741);
and AND3 (N1227, N1206, N1029, N571);
not NOT1 (N1228, N1226);
not NOT1 (N1229, N1228);
nand NAND2 (N1230, N1225, N377);
not NOT1 (N1231, N1205);
nor NOR3 (N1232, N1214, N664, N592);
nand NAND2 (N1233, N1231, N1042);
buf BUF1 (N1234, N1224);
nor NOR4 (N1235, N1232, N819, N765, N901);
nor NOR4 (N1236, N1235, N1201, N222, N631);
nand NAND2 (N1237, N1234, N828);
nor NOR3 (N1238, N1213, N965, N280);
buf BUF1 (N1239, N1222);
buf BUF1 (N1240, N1212);
xor XOR2 (N1241, N1230, N1033);
buf BUF1 (N1242, N1239);
nand NAND2 (N1243, N1237, N362);
and AND2 (N1244, N1227, N438);
buf BUF1 (N1245, N1215);
nor NOR4 (N1246, N1244, N1245, N1069, N91);
not NOT1 (N1247, N115);
or OR4 (N1248, N1236, N1079, N259, N1127);
and AND4 (N1249, N1246, N819, N1025, N6);
buf BUF1 (N1250, N1229);
and AND4 (N1251, N1242, N553, N588, N1055);
buf BUF1 (N1252, N1240);
nor NOR3 (N1253, N1251, N193, N1059);
buf BUF1 (N1254, N1233);
nor NOR2 (N1255, N1253, N523);
xor XOR2 (N1256, N1247, N853);
nand NAND3 (N1257, N1256, N338, N578);
buf BUF1 (N1258, N1255);
not NOT1 (N1259, N1258);
not NOT1 (N1260, N1243);
not NOT1 (N1261, N1241);
not NOT1 (N1262, N1257);
and AND4 (N1263, N1260, N572, N748, N365);
xor XOR2 (N1264, N1254, N55);
not NOT1 (N1265, N1248);
not NOT1 (N1266, N1264);
nor NOR2 (N1267, N1249, N1167);
and AND2 (N1268, N1259, N469);
nand NAND3 (N1269, N1268, N569, N8);
or OR2 (N1270, N1265, N441);
nor NOR4 (N1271, N1269, N42, N257, N786);
nor NOR4 (N1272, N1238, N505, N885, N1260);
buf BUF1 (N1273, N1271);
buf BUF1 (N1274, N1273);
nor NOR4 (N1275, N1252, N867, N1121, N738);
nor NOR2 (N1276, N1250, N380);
not NOT1 (N1277, N1274);
xor XOR2 (N1278, N1267, N612);
not NOT1 (N1279, N1277);
not NOT1 (N1280, N1275);
nor NOR4 (N1281, N1279, N638, N438, N1062);
or OR4 (N1282, N1281, N1214, N517, N711);
and AND2 (N1283, N1261, N761);
xor XOR2 (N1284, N1266, N1116);
xor XOR2 (N1285, N1280, N552);
or OR2 (N1286, N1282, N226);
nor NOR4 (N1287, N1285, N166, N381, N1243);
xor XOR2 (N1288, N1283, N718);
buf BUF1 (N1289, N1270);
nor NOR4 (N1290, N1289, N1255, N707, N360);
nor NOR4 (N1291, N1284, N233, N757, N1062);
nor NOR4 (N1292, N1272, N78, N399, N376);
not NOT1 (N1293, N1288);
buf BUF1 (N1294, N1290);
buf BUF1 (N1295, N1276);
buf BUF1 (N1296, N1287);
nand NAND4 (N1297, N1294, N1010, N479, N811);
xor XOR2 (N1298, N1293, N82);
nor NOR3 (N1299, N1291, N1221, N578);
nor NOR3 (N1300, N1298, N465, N318);
xor XOR2 (N1301, N1296, N1145);
xor XOR2 (N1302, N1263, N647);
or OR3 (N1303, N1286, N43, N220);
or OR4 (N1304, N1301, N919, N26, N908);
xor XOR2 (N1305, N1292, N375);
nor NOR3 (N1306, N1304, N401, N824);
nor NOR3 (N1307, N1302, N1222, N135);
and AND2 (N1308, N1305, N107);
buf BUF1 (N1309, N1299);
xor XOR2 (N1310, N1306, N1205);
not NOT1 (N1311, N1303);
buf BUF1 (N1312, N1307);
xor XOR2 (N1313, N1297, N208);
xor XOR2 (N1314, N1278, N1106);
not NOT1 (N1315, N1312);
not NOT1 (N1316, N1295);
buf BUF1 (N1317, N1314);
or OR4 (N1318, N1310, N111, N869, N1100);
and AND4 (N1319, N1300, N829, N379, N982);
nor NOR4 (N1320, N1262, N729, N89, N35);
and AND2 (N1321, N1313, N869);
nand NAND4 (N1322, N1321, N20, N701, N672);
not NOT1 (N1323, N1311);
buf BUF1 (N1324, N1317);
nand NAND3 (N1325, N1319, N759, N674);
and AND3 (N1326, N1320, N384, N920);
buf BUF1 (N1327, N1325);
and AND4 (N1328, N1318, N238, N604, N1165);
buf BUF1 (N1329, N1326);
xor XOR2 (N1330, N1327, N221);
xor XOR2 (N1331, N1308, N1139);
nor NOR4 (N1332, N1323, N471, N163, N337);
xor XOR2 (N1333, N1309, N1277);
nor NOR2 (N1334, N1316, N1238);
or OR4 (N1335, N1324, N193, N1280, N87);
or OR3 (N1336, N1333, N1272, N170);
nand NAND4 (N1337, N1328, N710, N1108, N592);
and AND3 (N1338, N1337, N125, N525);
buf BUF1 (N1339, N1332);
buf BUF1 (N1340, N1338);
buf BUF1 (N1341, N1336);
xor XOR2 (N1342, N1330, N1280);
buf BUF1 (N1343, N1329);
xor XOR2 (N1344, N1335, N1017);
and AND2 (N1345, N1339, N99);
and AND3 (N1346, N1341, N362, N340);
and AND2 (N1347, N1334, N851);
nand NAND2 (N1348, N1343, N1208);
and AND3 (N1349, N1331, N822, N670);
xor XOR2 (N1350, N1347, N539);
or OR2 (N1351, N1344, N33);
buf BUF1 (N1352, N1349);
and AND3 (N1353, N1315, N1162, N1245);
or OR4 (N1354, N1350, N547, N1303, N1105);
or OR2 (N1355, N1340, N431);
xor XOR2 (N1356, N1345, N823);
and AND2 (N1357, N1355, N109);
or OR4 (N1358, N1348, N943, N1103, N150);
not NOT1 (N1359, N1353);
xor XOR2 (N1360, N1322, N1314);
buf BUF1 (N1361, N1352);
and AND3 (N1362, N1356, N537, N1350);
xor XOR2 (N1363, N1359, N1000);
nor NOR2 (N1364, N1351, N707);
nor NOR2 (N1365, N1342, N662);
nor NOR3 (N1366, N1357, N295, N360);
xor XOR2 (N1367, N1361, N192);
or OR2 (N1368, N1366, N429);
and AND4 (N1369, N1365, N446, N1089, N227);
or OR3 (N1370, N1360, N480, N123);
not NOT1 (N1371, N1369);
or OR2 (N1372, N1362, N250);
xor XOR2 (N1373, N1364, N237);
and AND4 (N1374, N1346, N141, N1367, N1023);
buf BUF1 (N1375, N59);
and AND3 (N1376, N1371, N647, N179);
not NOT1 (N1377, N1370);
or OR2 (N1378, N1354, N1349);
and AND3 (N1379, N1374, N818, N268);
not NOT1 (N1380, N1373);
and AND3 (N1381, N1358, N470, N1205);
xor XOR2 (N1382, N1363, N855);
or OR3 (N1383, N1368, N1346, N571);
and AND4 (N1384, N1381, N587, N1190, N70);
not NOT1 (N1385, N1376);
nor NOR4 (N1386, N1382, N515, N1308, N740);
nand NAND4 (N1387, N1383, N1194, N354, N1032);
and AND2 (N1388, N1384, N341);
buf BUF1 (N1389, N1388);
xor XOR2 (N1390, N1372, N1233);
xor XOR2 (N1391, N1380, N1056);
not NOT1 (N1392, N1390);
buf BUF1 (N1393, N1392);
buf BUF1 (N1394, N1391);
nor NOR3 (N1395, N1389, N1334, N1107);
xor XOR2 (N1396, N1386, N32);
xor XOR2 (N1397, N1387, N437);
not NOT1 (N1398, N1397);
nor NOR4 (N1399, N1396, N760, N1086, N359);
not NOT1 (N1400, N1379);
or OR4 (N1401, N1393, N1377, N302, N1110);
and AND4 (N1402, N227, N659, N292, N1130);
or OR3 (N1403, N1400, N995, N1359);
and AND4 (N1404, N1403, N983, N737, N862);
or OR2 (N1405, N1378, N796);
buf BUF1 (N1406, N1375);
nand NAND3 (N1407, N1405, N374, N715);
not NOT1 (N1408, N1404);
nor NOR4 (N1409, N1401, N325, N1162, N397);
nor NOR2 (N1410, N1398, N526);
nor NOR3 (N1411, N1399, N294, N777);
nand NAND2 (N1412, N1402, N989);
buf BUF1 (N1413, N1407);
nand NAND2 (N1414, N1410, N1356);
nor NOR2 (N1415, N1412, N844);
or OR3 (N1416, N1413, N19, N1250);
not NOT1 (N1417, N1409);
not NOT1 (N1418, N1406);
xor XOR2 (N1419, N1417, N986);
or OR4 (N1420, N1416, N207, N379, N840);
nand NAND2 (N1421, N1415, N740);
nand NAND2 (N1422, N1408, N581);
not NOT1 (N1423, N1385);
or OR3 (N1424, N1422, N313, N747);
or OR2 (N1425, N1411, N1310);
nand NAND2 (N1426, N1395, N524);
xor XOR2 (N1427, N1414, N366);
nor NOR2 (N1428, N1418, N1099);
and AND3 (N1429, N1427, N983, N569);
nand NAND4 (N1430, N1420, N1153, N870, N1153);
nand NAND4 (N1431, N1423, N1125, N276, N1426);
nor NOR3 (N1432, N1260, N1189, N343);
or OR4 (N1433, N1424, N781, N560, N1129);
not NOT1 (N1434, N1421);
nor NOR2 (N1435, N1428, N313);
xor XOR2 (N1436, N1434, N1167);
and AND2 (N1437, N1425, N279);
not NOT1 (N1438, N1431);
not NOT1 (N1439, N1438);
not NOT1 (N1440, N1429);
or OR2 (N1441, N1433, N1228);
and AND3 (N1442, N1440, N427, N289);
nor NOR3 (N1443, N1419, N50, N150);
nor NOR4 (N1444, N1439, N1093, N1198, N586);
nand NAND3 (N1445, N1430, N856, N1121);
nor NOR2 (N1446, N1435, N1262);
and AND4 (N1447, N1436, N1128, N109, N437);
xor XOR2 (N1448, N1444, N1424);
nand NAND3 (N1449, N1394, N634, N1176);
buf BUF1 (N1450, N1449);
not NOT1 (N1451, N1446);
nor NOR3 (N1452, N1448, N1356, N411);
nor NOR3 (N1453, N1452, N1255, N942);
nor NOR2 (N1454, N1443, N851);
and AND3 (N1455, N1451, N396, N268);
or OR3 (N1456, N1447, N584, N551);
nand NAND3 (N1457, N1456, N595, N942);
and AND4 (N1458, N1450, N953, N995, N623);
xor XOR2 (N1459, N1454, N972);
and AND3 (N1460, N1457, N962, N1106);
buf BUF1 (N1461, N1453);
or OR2 (N1462, N1461, N1318);
and AND2 (N1463, N1437, N929);
not NOT1 (N1464, N1459);
nor NOR4 (N1465, N1441, N1116, N283, N1048);
xor XOR2 (N1466, N1462, N1103);
buf BUF1 (N1467, N1458);
buf BUF1 (N1468, N1442);
and AND3 (N1469, N1468, N1160, N1201);
buf BUF1 (N1470, N1463);
or OR4 (N1471, N1470, N1029, N374, N1213);
nor NOR3 (N1472, N1467, N661, N382);
buf BUF1 (N1473, N1465);
xor XOR2 (N1474, N1471, N354);
nor NOR4 (N1475, N1445, N514, N314, N429);
not NOT1 (N1476, N1464);
and AND3 (N1477, N1469, N1439, N693);
nor NOR4 (N1478, N1460, N1131, N1253, N580);
not NOT1 (N1479, N1455);
buf BUF1 (N1480, N1475);
not NOT1 (N1481, N1472);
nand NAND4 (N1482, N1479, N710, N1218, N719);
xor XOR2 (N1483, N1466, N757);
buf BUF1 (N1484, N1477);
xor XOR2 (N1485, N1474, N294);
and AND4 (N1486, N1478, N1145, N22, N1475);
nor NOR4 (N1487, N1482, N606, N1127, N1103);
not NOT1 (N1488, N1487);
nand NAND3 (N1489, N1432, N730, N816);
or OR4 (N1490, N1483, N800, N935, N452);
xor XOR2 (N1491, N1480, N253);
or OR2 (N1492, N1484, N965);
and AND4 (N1493, N1476, N777, N487, N661);
and AND3 (N1494, N1481, N1188, N83);
nor NOR3 (N1495, N1490, N1122, N352);
nand NAND2 (N1496, N1494, N297);
xor XOR2 (N1497, N1493, N836);
xor XOR2 (N1498, N1492, N965);
and AND2 (N1499, N1496, N160);
not NOT1 (N1500, N1473);
xor XOR2 (N1501, N1488, N178);
nand NAND4 (N1502, N1485, N1345, N895, N330);
or OR3 (N1503, N1489, N802, N830);
or OR3 (N1504, N1491, N1477, N434);
and AND4 (N1505, N1498, N641, N977, N690);
and AND2 (N1506, N1497, N255);
or OR3 (N1507, N1502, N211, N55);
nand NAND2 (N1508, N1501, N509);
nor NOR3 (N1509, N1503, N531, N835);
buf BUF1 (N1510, N1500);
xor XOR2 (N1511, N1506, N979);
nor NOR4 (N1512, N1507, N530, N382, N102);
not NOT1 (N1513, N1512);
nand NAND3 (N1514, N1510, N905, N1335);
or OR2 (N1515, N1505, N479);
nor NOR3 (N1516, N1504, N166, N1111);
and AND4 (N1517, N1486, N585, N1010, N1349);
nand NAND3 (N1518, N1508, N1012, N1509);
buf BUF1 (N1519, N1375);
xor XOR2 (N1520, N1495, N1396);
or OR2 (N1521, N1519, N1383);
nand NAND4 (N1522, N1514, N994, N501, N218);
not NOT1 (N1523, N1511);
buf BUF1 (N1524, N1520);
xor XOR2 (N1525, N1515, N1491);
or OR4 (N1526, N1521, N1460, N928, N1114);
buf BUF1 (N1527, N1517);
or OR2 (N1528, N1516, N1327);
xor XOR2 (N1529, N1526, N16);
nand NAND3 (N1530, N1499, N188, N1054);
nor NOR2 (N1531, N1513, N471);
and AND2 (N1532, N1527, N1161);
xor XOR2 (N1533, N1522, N388);
not NOT1 (N1534, N1529);
nand NAND3 (N1535, N1534, N1192, N167);
or OR4 (N1536, N1530, N321, N1155, N387);
or OR2 (N1537, N1528, N1227);
buf BUF1 (N1538, N1536);
buf BUF1 (N1539, N1533);
xor XOR2 (N1540, N1535, N963);
or OR2 (N1541, N1523, N757);
buf BUF1 (N1542, N1537);
nor NOR2 (N1543, N1540, N1103);
nor NOR4 (N1544, N1542, N1295, N64, N706);
xor XOR2 (N1545, N1532, N69);
not NOT1 (N1546, N1531);
or OR4 (N1547, N1544, N606, N371, N179);
nand NAND3 (N1548, N1543, N1122, N778);
not NOT1 (N1549, N1548);
and AND4 (N1550, N1546, N3, N1370, N1252);
buf BUF1 (N1551, N1539);
nand NAND2 (N1552, N1551, N497);
and AND3 (N1553, N1524, N474, N1448);
nand NAND2 (N1554, N1538, N431);
and AND4 (N1555, N1553, N1213, N51, N321);
nand NAND2 (N1556, N1541, N1034);
xor XOR2 (N1557, N1556, N226);
buf BUF1 (N1558, N1518);
not NOT1 (N1559, N1557);
not NOT1 (N1560, N1549);
and AND4 (N1561, N1545, N861, N496, N678);
xor XOR2 (N1562, N1547, N577);
nor NOR3 (N1563, N1555, N1245, N421);
not NOT1 (N1564, N1563);
nand NAND2 (N1565, N1558, N619);
not NOT1 (N1566, N1550);
xor XOR2 (N1567, N1525, N614);
nor NOR4 (N1568, N1559, N1075, N821, N1123);
and AND3 (N1569, N1567, N743, N1034);
nor NOR4 (N1570, N1560, N773, N974, N1251);
buf BUF1 (N1571, N1569);
nor NOR2 (N1572, N1570, N1514);
or OR2 (N1573, N1562, N698);
not NOT1 (N1574, N1568);
xor XOR2 (N1575, N1565, N1235);
or OR4 (N1576, N1561, N1098, N709, N1499);
buf BUF1 (N1577, N1573);
buf BUF1 (N1578, N1571);
buf BUF1 (N1579, N1566);
nor NOR3 (N1580, N1576, N244, N69);
buf BUF1 (N1581, N1579);
or OR3 (N1582, N1578, N1127, N382);
and AND4 (N1583, N1564, N1328, N29, N946);
xor XOR2 (N1584, N1572, N349);
buf BUF1 (N1585, N1554);
buf BUF1 (N1586, N1577);
not NOT1 (N1587, N1586);
xor XOR2 (N1588, N1583, N9);
buf BUF1 (N1589, N1584);
xor XOR2 (N1590, N1588, N611);
and AND4 (N1591, N1575, N1589, N1045, N1260);
not NOT1 (N1592, N1360);
and AND3 (N1593, N1574, N679, N853);
nor NOR2 (N1594, N1592, N754);
and AND3 (N1595, N1593, N1426, N381);
or OR4 (N1596, N1585, N34, N1358, N984);
nand NAND4 (N1597, N1581, N85, N1532, N942);
xor XOR2 (N1598, N1590, N659);
xor XOR2 (N1599, N1587, N939);
not NOT1 (N1600, N1595);
xor XOR2 (N1601, N1598, N975);
and AND3 (N1602, N1594, N222, N666);
or OR2 (N1603, N1602, N432);
nor NOR4 (N1604, N1582, N783, N740, N90);
and AND2 (N1605, N1600, N128);
not NOT1 (N1606, N1580);
buf BUF1 (N1607, N1603);
and AND2 (N1608, N1604, N1511);
or OR2 (N1609, N1606, N519);
and AND4 (N1610, N1608, N704, N632, N920);
and AND3 (N1611, N1601, N530, N773);
nand NAND2 (N1612, N1605, N1485);
buf BUF1 (N1613, N1552);
and AND4 (N1614, N1591, N1367, N1393, N246);
nand NAND3 (N1615, N1597, N1303, N224);
and AND4 (N1616, N1615, N1288, N76, N343);
buf BUF1 (N1617, N1596);
and AND2 (N1618, N1614, N995);
buf BUF1 (N1619, N1611);
not NOT1 (N1620, N1617);
not NOT1 (N1621, N1607);
and AND2 (N1622, N1620, N9);
buf BUF1 (N1623, N1621);
and AND4 (N1624, N1612, N511, N1042, N485);
and AND4 (N1625, N1618, N1213, N1282, N236);
buf BUF1 (N1626, N1623);
nor NOR2 (N1627, N1622, N241);
nand NAND2 (N1628, N1625, N399);
buf BUF1 (N1629, N1610);
or OR4 (N1630, N1629, N655, N73, N1602);
and AND4 (N1631, N1619, N1596, N1572, N1360);
and AND4 (N1632, N1613, N1009, N621, N703);
not NOT1 (N1633, N1630);
and AND4 (N1634, N1609, N890, N749, N582);
nand NAND2 (N1635, N1626, N1464);
nor NOR3 (N1636, N1633, N1022, N1121);
buf BUF1 (N1637, N1627);
or OR3 (N1638, N1635, N359, N1115);
nor NOR2 (N1639, N1634, N569);
buf BUF1 (N1640, N1628);
xor XOR2 (N1641, N1631, N878);
and AND2 (N1642, N1640, N966);
xor XOR2 (N1643, N1616, N288);
and AND4 (N1644, N1638, N919, N96, N698);
xor XOR2 (N1645, N1632, N726);
buf BUF1 (N1646, N1642);
xor XOR2 (N1647, N1637, N896);
not NOT1 (N1648, N1644);
and AND3 (N1649, N1646, N781, N1314);
and AND3 (N1650, N1624, N1442, N552);
or OR4 (N1651, N1649, N609, N331, N478);
or OR3 (N1652, N1645, N1651, N1413);
nand NAND3 (N1653, N1272, N1591, N724);
buf BUF1 (N1654, N1643);
or OR2 (N1655, N1599, N324);
and AND3 (N1656, N1636, N507, N1613);
and AND4 (N1657, N1654, N532, N546, N326);
nand NAND2 (N1658, N1647, N1072);
nor NOR4 (N1659, N1658, N1423, N929, N431);
nor NOR3 (N1660, N1652, N272, N1520);
not NOT1 (N1661, N1659);
xor XOR2 (N1662, N1657, N1389);
not NOT1 (N1663, N1641);
or OR2 (N1664, N1648, N125);
or OR3 (N1665, N1655, N108, N369);
buf BUF1 (N1666, N1661);
buf BUF1 (N1667, N1664);
buf BUF1 (N1668, N1639);
and AND4 (N1669, N1650, N494, N494, N677);
not NOT1 (N1670, N1665);
or OR3 (N1671, N1660, N228, N1338);
xor XOR2 (N1672, N1666, N1559);
nor NOR3 (N1673, N1670, N981, N851);
not NOT1 (N1674, N1656);
xor XOR2 (N1675, N1668, N863);
buf BUF1 (N1676, N1672);
or OR4 (N1677, N1673, N1277, N1116, N1350);
xor XOR2 (N1678, N1653, N1055);
and AND2 (N1679, N1678, N1171);
and AND3 (N1680, N1679, N694, N626);
or OR3 (N1681, N1674, N1002, N398);
buf BUF1 (N1682, N1677);
or OR2 (N1683, N1663, N1631);
nand NAND4 (N1684, N1681, N972, N681, N801);
nand NAND2 (N1685, N1675, N759);
xor XOR2 (N1686, N1667, N190);
nor NOR4 (N1687, N1682, N695, N1052, N188);
nand NAND2 (N1688, N1671, N1136);
nor NOR3 (N1689, N1688, N1397, N1206);
and AND2 (N1690, N1684, N1058);
and AND3 (N1691, N1680, N97, N1261);
nand NAND4 (N1692, N1683, N1093, N1640, N1);
not NOT1 (N1693, N1662);
nor NOR2 (N1694, N1689, N1094);
and AND2 (N1695, N1693, N372);
and AND3 (N1696, N1690, N419, N1249);
and AND2 (N1697, N1687, N1004);
xor XOR2 (N1698, N1686, N1082);
and AND4 (N1699, N1694, N322, N1164, N508);
xor XOR2 (N1700, N1697, N535);
nand NAND4 (N1701, N1691, N608, N732, N240);
buf BUF1 (N1702, N1692);
buf BUF1 (N1703, N1701);
nand NAND4 (N1704, N1700, N126, N34, N1600);
nor NOR3 (N1705, N1704, N966, N1632);
xor XOR2 (N1706, N1703, N1184);
and AND3 (N1707, N1706, N385, N234);
buf BUF1 (N1708, N1707);
nor NOR3 (N1709, N1698, N525, N1055);
nand NAND2 (N1710, N1705, N727);
or OR2 (N1711, N1695, N342);
buf BUF1 (N1712, N1709);
and AND2 (N1713, N1696, N1387);
xor XOR2 (N1714, N1713, N1556);
not NOT1 (N1715, N1702);
nor NOR2 (N1716, N1699, N1686);
or OR4 (N1717, N1715, N116, N498, N19);
not NOT1 (N1718, N1676);
nor NOR3 (N1719, N1711, N1473, N119);
not NOT1 (N1720, N1685);
and AND4 (N1721, N1712, N734, N1337, N1558);
buf BUF1 (N1722, N1669);
xor XOR2 (N1723, N1717, N753);
not NOT1 (N1724, N1718);
xor XOR2 (N1725, N1720, N1057);
or OR2 (N1726, N1725, N1299);
buf BUF1 (N1727, N1719);
and AND3 (N1728, N1716, N775, N710);
not NOT1 (N1729, N1727);
nand NAND3 (N1730, N1723, N955, N379);
nor NOR2 (N1731, N1729, N805);
nand NAND4 (N1732, N1708, N1358, N1335, N74);
nor NOR2 (N1733, N1714, N519);
and AND4 (N1734, N1728, N867, N1076, N761);
or OR3 (N1735, N1734, N1665, N679);
or OR2 (N1736, N1722, N328);
and AND4 (N1737, N1733, N1079, N1296, N586);
or OR3 (N1738, N1724, N1522, N984);
or OR2 (N1739, N1730, N1578);
xor XOR2 (N1740, N1735, N1059);
and AND3 (N1741, N1732, N1736, N1361);
nand NAND3 (N1742, N458, N912, N844);
or OR2 (N1743, N1710, N1649);
buf BUF1 (N1744, N1721);
nor NOR4 (N1745, N1738, N1143, N610, N452);
nor NOR3 (N1746, N1744, N1472, N1003);
xor XOR2 (N1747, N1746, N1708);
nor NOR3 (N1748, N1739, N867, N1413);
nor NOR4 (N1749, N1740, N1568, N494, N656);
not NOT1 (N1750, N1743);
and AND3 (N1751, N1747, N1592, N1517);
nand NAND4 (N1752, N1741, N465, N1397, N759);
and AND2 (N1753, N1748, N640);
buf BUF1 (N1754, N1750);
nand NAND3 (N1755, N1726, N1050, N273);
nand NAND2 (N1756, N1754, N820);
or OR3 (N1757, N1753, N6, N1549);
and AND2 (N1758, N1757, N1686);
buf BUF1 (N1759, N1752);
and AND3 (N1760, N1759, N183, N1375);
buf BUF1 (N1761, N1755);
not NOT1 (N1762, N1761);
xor XOR2 (N1763, N1731, N1551);
not NOT1 (N1764, N1763);
nand NAND3 (N1765, N1758, N535, N1109);
nor NOR4 (N1766, N1749, N1571, N1761, N1031);
nand NAND4 (N1767, N1756, N1122, N871, N542);
nand NAND4 (N1768, N1765, N740, N750, N1211);
or OR4 (N1769, N1760, N320, N796, N1233);
nor NOR4 (N1770, N1742, N1678, N615, N1398);
not NOT1 (N1771, N1737);
nand NAND2 (N1772, N1768, N1756);
buf BUF1 (N1773, N1772);
nand NAND2 (N1774, N1751, N510);
nand NAND4 (N1775, N1769, N566, N837, N1140);
nand NAND2 (N1776, N1766, N509);
not NOT1 (N1777, N1776);
and AND3 (N1778, N1767, N1688, N1585);
nor NOR3 (N1779, N1773, N1433, N1755);
not NOT1 (N1780, N1777);
or OR3 (N1781, N1762, N988, N249);
and AND2 (N1782, N1780, N1321);
not NOT1 (N1783, N1779);
not NOT1 (N1784, N1764);
nand NAND3 (N1785, N1745, N948, N265);
and AND4 (N1786, N1784, N773, N401, N133);
or OR3 (N1787, N1781, N1484, N835);
not NOT1 (N1788, N1782);
xor XOR2 (N1789, N1778, N40);
not NOT1 (N1790, N1788);
nand NAND4 (N1791, N1785, N854, N1325, N68);
xor XOR2 (N1792, N1789, N1370);
and AND3 (N1793, N1774, N1373, N1702);
nand NAND4 (N1794, N1770, N1643, N1640, N283);
and AND4 (N1795, N1793, N677, N1424, N436);
and AND4 (N1796, N1792, N1008, N1589, N1684);
and AND4 (N1797, N1783, N368, N981, N1652);
nor NOR4 (N1798, N1786, N1487, N809, N879);
xor XOR2 (N1799, N1771, N1124);
nor NOR3 (N1800, N1795, N1560, N863);
buf BUF1 (N1801, N1787);
buf BUF1 (N1802, N1791);
not NOT1 (N1803, N1796);
xor XOR2 (N1804, N1790, N715);
xor XOR2 (N1805, N1802, N1343);
xor XOR2 (N1806, N1800, N1292);
and AND2 (N1807, N1775, N1052);
buf BUF1 (N1808, N1806);
nor NOR4 (N1809, N1808, N1524, N787, N1123);
or OR4 (N1810, N1799, N1477, N669, N97);
or OR3 (N1811, N1803, N760, N178);
xor XOR2 (N1812, N1797, N1656);
xor XOR2 (N1813, N1812, N1217);
xor XOR2 (N1814, N1809, N605);
nand NAND4 (N1815, N1794, N225, N1420, N960);
or OR3 (N1816, N1815, N520, N647);
or OR4 (N1817, N1798, N1691, N785, N48);
xor XOR2 (N1818, N1811, N920);
not NOT1 (N1819, N1818);
nand NAND3 (N1820, N1810, N461, N1412);
buf BUF1 (N1821, N1813);
or OR3 (N1822, N1816, N921, N513);
nand NAND3 (N1823, N1817, N1451, N105);
not NOT1 (N1824, N1805);
and AND3 (N1825, N1807, N1088, N989);
nor NOR2 (N1826, N1822, N850);
not NOT1 (N1827, N1804);
nand NAND4 (N1828, N1825, N1052, N894, N1701);
nor NOR4 (N1829, N1824, N549, N45, N90);
nand NAND2 (N1830, N1814, N1405);
buf BUF1 (N1831, N1830);
nand NAND3 (N1832, N1826, N925, N768);
nor NOR3 (N1833, N1801, N1623, N1371);
and AND4 (N1834, N1832, N1761, N1493, N475);
not NOT1 (N1835, N1820);
or OR4 (N1836, N1834, N452, N769, N1224);
and AND4 (N1837, N1836, N1513, N1296, N78);
nand NAND2 (N1838, N1835, N359);
buf BUF1 (N1839, N1837);
nand NAND2 (N1840, N1838, N452);
and AND2 (N1841, N1840, N77);
buf BUF1 (N1842, N1821);
nand NAND2 (N1843, N1842, N1160);
nor NOR2 (N1844, N1827, N1693);
or OR3 (N1845, N1829, N497, N690);
nand NAND4 (N1846, N1831, N369, N1732, N1166);
nand NAND2 (N1847, N1839, N69);
or OR3 (N1848, N1846, N1357, N1545);
xor XOR2 (N1849, N1845, N223);
and AND2 (N1850, N1828, N1696);
buf BUF1 (N1851, N1847);
nor NOR4 (N1852, N1848, N660, N1275, N462);
buf BUF1 (N1853, N1833);
and AND3 (N1854, N1851, N1430, N1307);
not NOT1 (N1855, N1852);
nand NAND4 (N1856, N1823, N340, N121, N1344);
and AND3 (N1857, N1819, N939, N1125);
xor XOR2 (N1858, N1841, N1387);
not NOT1 (N1859, N1858);
buf BUF1 (N1860, N1855);
and AND4 (N1861, N1859, N1542, N1171, N457);
buf BUF1 (N1862, N1861);
nor NOR4 (N1863, N1856, N292, N812, N1545);
not NOT1 (N1864, N1849);
nor NOR2 (N1865, N1862, N569);
buf BUF1 (N1866, N1843);
not NOT1 (N1867, N1866);
xor XOR2 (N1868, N1854, N273);
buf BUF1 (N1869, N1867);
xor XOR2 (N1870, N1869, N173);
buf BUF1 (N1871, N1868);
or OR4 (N1872, N1853, N230, N550, N1172);
xor XOR2 (N1873, N1863, N1153);
nand NAND3 (N1874, N1857, N953, N124);
or OR2 (N1875, N1871, N593);
nor NOR4 (N1876, N1870, N1174, N435, N1251);
not NOT1 (N1877, N1874);
and AND4 (N1878, N1864, N1466, N63, N893);
buf BUF1 (N1879, N1878);
buf BUF1 (N1880, N1844);
buf BUF1 (N1881, N1873);
buf BUF1 (N1882, N1880);
or OR2 (N1883, N1872, N1477);
nand NAND2 (N1884, N1875, N1732);
nor NOR2 (N1885, N1884, N125);
and AND4 (N1886, N1850, N1552, N908, N1202);
not NOT1 (N1887, N1886);
not NOT1 (N1888, N1860);
buf BUF1 (N1889, N1881);
not NOT1 (N1890, N1879);
nor NOR2 (N1891, N1877, N1344);
nor NOR2 (N1892, N1885, N1589);
or OR3 (N1893, N1889, N503, N701);
buf BUF1 (N1894, N1882);
buf BUF1 (N1895, N1888);
nor NOR3 (N1896, N1876, N651, N696);
nor NOR3 (N1897, N1892, N197, N1361);
nor NOR2 (N1898, N1897, N1020);
xor XOR2 (N1899, N1865, N702);
buf BUF1 (N1900, N1896);
or OR2 (N1901, N1883, N1463);
xor XOR2 (N1902, N1895, N1471);
nand NAND3 (N1903, N1887, N236, N159);
and AND2 (N1904, N1890, N1826);
nor NOR4 (N1905, N1893, N740, N452, N300);
nand NAND2 (N1906, N1894, N1413);
nor NOR2 (N1907, N1901, N839);
not NOT1 (N1908, N1891);
buf BUF1 (N1909, N1907);
xor XOR2 (N1910, N1908, N906);
not NOT1 (N1911, N1906);
and AND2 (N1912, N1904, N982);
or OR3 (N1913, N1911, N1150, N693);
or OR2 (N1914, N1903, N669);
nor NOR4 (N1915, N1910, N1836, N815, N827);
or OR4 (N1916, N1905, N202, N1010, N141);
not NOT1 (N1917, N1912);
buf BUF1 (N1918, N1909);
buf BUF1 (N1919, N1898);
nand NAND3 (N1920, N1916, N1258, N1172);
nand NAND2 (N1921, N1919, N818);
not NOT1 (N1922, N1920);
or OR4 (N1923, N1899, N1238, N1440, N999);
buf BUF1 (N1924, N1915);
buf BUF1 (N1925, N1917);
xor XOR2 (N1926, N1923, N1116);
buf BUF1 (N1927, N1913);
xor XOR2 (N1928, N1902, N140);
xor XOR2 (N1929, N1927, N1472);
nor NOR4 (N1930, N1918, N1681, N29, N1007);
buf BUF1 (N1931, N1900);
not NOT1 (N1932, N1921);
buf BUF1 (N1933, N1929);
buf BUF1 (N1934, N1914);
nor NOR3 (N1935, N1922, N954, N1415);
nand NAND2 (N1936, N1932, N763);
or OR2 (N1937, N1930, N18);
or OR4 (N1938, N1924, N972, N1466, N314);
buf BUF1 (N1939, N1925);
or OR3 (N1940, N1926, N67, N1143);
buf BUF1 (N1941, N1939);
or OR2 (N1942, N1937, N668);
and AND4 (N1943, N1942, N1337, N996, N1831);
nor NOR4 (N1944, N1931, N548, N227, N1099);
buf BUF1 (N1945, N1940);
nand NAND3 (N1946, N1933, N1548, N264);
nand NAND3 (N1947, N1938, N1497, N805);
xor XOR2 (N1948, N1935, N1584);
xor XOR2 (N1949, N1948, N536);
and AND2 (N1950, N1947, N1326);
buf BUF1 (N1951, N1950);
nand NAND4 (N1952, N1945, N1770, N828, N319);
not NOT1 (N1953, N1928);
nand NAND3 (N1954, N1949, N88, N617);
nor NOR3 (N1955, N1954, N406, N37);
or OR3 (N1956, N1944, N1827, N10);
or OR2 (N1957, N1934, N141);
not NOT1 (N1958, N1955);
xor XOR2 (N1959, N1957, N1794);
and AND2 (N1960, N1956, N90);
buf BUF1 (N1961, N1951);
and AND3 (N1962, N1936, N1651, N1719);
xor XOR2 (N1963, N1960, N1508);
and AND2 (N1964, N1962, N1377);
nor NOR2 (N1965, N1953, N1765);
nor NOR3 (N1966, N1952, N1209, N162);
buf BUF1 (N1967, N1961);
nand NAND2 (N1968, N1959, N1619);
nand NAND4 (N1969, N1965, N1115, N833, N1234);
and AND2 (N1970, N1941, N1363);
or OR3 (N1971, N1943, N1703, N286);
not NOT1 (N1972, N1967);
nor NOR4 (N1973, N1966, N1466, N1422, N714);
nor NOR3 (N1974, N1968, N1763, N118);
nor NOR4 (N1975, N1964, N742, N1675, N1477);
nor NOR3 (N1976, N1969, N751, N1901);
not NOT1 (N1977, N1970);
buf BUF1 (N1978, N1976);
buf BUF1 (N1979, N1977);
or OR3 (N1980, N1972, N1853, N1630);
xor XOR2 (N1981, N1975, N966);
or OR4 (N1982, N1958, N116, N170, N59);
not NOT1 (N1983, N1980);
not NOT1 (N1984, N1982);
buf BUF1 (N1985, N1946);
nor NOR4 (N1986, N1984, N1205, N1319, N143);
buf BUF1 (N1987, N1974);
and AND3 (N1988, N1978, N441, N1065);
not NOT1 (N1989, N1979);
or OR2 (N1990, N1973, N1968);
or OR4 (N1991, N1981, N567, N1501, N919);
and AND4 (N1992, N1986, N526, N95, N929);
or OR2 (N1993, N1990, N252);
nor NOR4 (N1994, N1985, N535, N629, N1827);
nor NOR2 (N1995, N1993, N671);
xor XOR2 (N1996, N1983, N682);
xor XOR2 (N1997, N1992, N565);
not NOT1 (N1998, N1995);
nand NAND4 (N1999, N1991, N233, N660, N1395);
and AND2 (N2000, N1996, N555);
nand NAND4 (N2001, N1989, N916, N330, N1120);
and AND2 (N2002, N1971, N1186);
nand NAND2 (N2003, N1994, N1694);
xor XOR2 (N2004, N1999, N965);
xor XOR2 (N2005, N2001, N894);
and AND4 (N2006, N2002, N284, N1153, N1690);
not NOT1 (N2007, N2004);
xor XOR2 (N2008, N1963, N1328);
not NOT1 (N2009, N2008);
nand NAND4 (N2010, N2000, N17, N1746, N1002);
nand NAND3 (N2011, N2003, N724, N1717);
nor NOR4 (N2012, N2006, N869, N1007, N1307);
buf BUF1 (N2013, N1998);
or OR2 (N2014, N2005, N816);
buf BUF1 (N2015, N2014);
or OR2 (N2016, N2011, N859);
nand NAND3 (N2017, N2010, N425, N1604);
buf BUF1 (N2018, N1987);
not NOT1 (N2019, N2015);
or OR4 (N2020, N1997, N1421, N382, N156);
not NOT1 (N2021, N2017);
buf BUF1 (N2022, N2013);
or OR3 (N2023, N2019, N1183, N476);
buf BUF1 (N2024, N2007);
and AND4 (N2025, N1988, N1980, N1916, N942);
xor XOR2 (N2026, N2020, N675);
or OR4 (N2027, N2024, N778, N1160, N627);
or OR2 (N2028, N2016, N1157);
nand NAND3 (N2029, N2027, N1063, N686);
buf BUF1 (N2030, N2021);
and AND4 (N2031, N2028, N2003, N83, N552);
buf BUF1 (N2032, N2009);
or OR4 (N2033, N2022, N1852, N318, N54);
nand NAND2 (N2034, N2033, N76);
nor NOR4 (N2035, N2023, N1642, N547, N1896);
xor XOR2 (N2036, N2018, N1003);
not NOT1 (N2037, N2026);
buf BUF1 (N2038, N2035);
nor NOR4 (N2039, N2012, N425, N745, N873);
buf BUF1 (N2040, N2034);
nand NAND4 (N2041, N2031, N1355, N1533, N1348);
buf BUF1 (N2042, N2030);
and AND4 (N2043, N2032, N109, N554, N84);
and AND4 (N2044, N2038, N443, N1238, N769);
and AND2 (N2045, N2036, N798);
or OR4 (N2046, N2025, N1398, N1243, N2033);
nor NOR2 (N2047, N2040, N173);
not NOT1 (N2048, N2029);
not NOT1 (N2049, N2039);
buf BUF1 (N2050, N2046);
and AND4 (N2051, N2047, N761, N1610, N940);
nand NAND4 (N2052, N2048, N1781, N780, N1126);
or OR4 (N2053, N2043, N7, N1782, N1625);
not NOT1 (N2054, N2050);
and AND3 (N2055, N2054, N223, N2014);
nand NAND4 (N2056, N2053, N1782, N1376, N824);
nor NOR2 (N2057, N2042, N148);
nor NOR4 (N2058, N2055, N754, N173, N952);
nand NAND4 (N2059, N2049, N759, N278, N318);
nand NAND4 (N2060, N2056, N1045, N1, N14);
nand NAND4 (N2061, N2041, N384, N1178, N1069);
buf BUF1 (N2062, N2037);
or OR4 (N2063, N2044, N1718, N851, N1947);
not NOT1 (N2064, N2057);
nand NAND4 (N2065, N2060, N1799, N1192, N562);
xor XOR2 (N2066, N2051, N703);
nor NOR2 (N2067, N2062, N503);
or OR3 (N2068, N2067, N54, N1426);
nand NAND3 (N2069, N2052, N1924, N32);
not NOT1 (N2070, N2066);
or OR3 (N2071, N2068, N668, N1187);
nand NAND2 (N2072, N2070, N255);
or OR2 (N2073, N2061, N939);
nand NAND3 (N2074, N2045, N1876, N339);
xor XOR2 (N2075, N2059, N938);
nand NAND2 (N2076, N2073, N785);
or OR3 (N2077, N2069, N1050, N97);
nor NOR2 (N2078, N2071, N789);
not NOT1 (N2079, N2076);
nor NOR3 (N2080, N2058, N1427, N1499);
or OR4 (N2081, N2078, N1002, N662, N399);
or OR3 (N2082, N2064, N1676, N981);
nand NAND3 (N2083, N2074, N822, N1517);
xor XOR2 (N2084, N2082, N321);
and AND2 (N2085, N2063, N1200);
nand NAND4 (N2086, N2083, N414, N1324, N74);
nand NAND2 (N2087, N2079, N1995);
nand NAND4 (N2088, N2077, N173, N287, N1039);
or OR3 (N2089, N2085, N288, N1328);
and AND4 (N2090, N2072, N957, N455, N1810);
buf BUF1 (N2091, N2080);
or OR3 (N2092, N2089, N499, N1131);
nand NAND3 (N2093, N2087, N1829, N431);
or OR2 (N2094, N2093, N1271);
and AND2 (N2095, N2091, N200);
nor NOR4 (N2096, N2086, N21, N1658, N219);
not NOT1 (N2097, N2065);
buf BUF1 (N2098, N2084);
xor XOR2 (N2099, N2094, N533);
buf BUF1 (N2100, N2095);
xor XOR2 (N2101, N2090, N1653);
nor NOR3 (N2102, N2100, N88, N1061);
and AND2 (N2103, N2097, N1182);
not NOT1 (N2104, N2103);
not NOT1 (N2105, N2088);
xor XOR2 (N2106, N2081, N533);
and AND3 (N2107, N2096, N1870, N1630);
nor NOR3 (N2108, N2092, N1327, N1503);
buf BUF1 (N2109, N2102);
and AND4 (N2110, N2109, N1381, N1418, N919);
and AND2 (N2111, N2108, N1634);
nand NAND4 (N2112, N2101, N115, N1233, N1542);
nor NOR4 (N2113, N2112, N661, N2035, N28);
nand NAND2 (N2114, N2111, N28);
and AND3 (N2115, N2107, N1322, N1995);
or OR3 (N2116, N2098, N8, N1409);
not NOT1 (N2117, N2105);
xor XOR2 (N2118, N2106, N1208);
not NOT1 (N2119, N2114);
nor NOR4 (N2120, N2116, N1518, N248, N1600);
and AND4 (N2121, N2099, N1361, N1999, N1303);
buf BUF1 (N2122, N2119);
nor NOR4 (N2123, N2075, N1611, N219, N1539);
or OR3 (N2124, N2120, N1298, N146);
or OR2 (N2125, N2122, N379);
xor XOR2 (N2126, N2121, N1026);
not NOT1 (N2127, N2113);
xor XOR2 (N2128, N2126, N1727);
and AND3 (N2129, N2117, N696, N394);
nand NAND2 (N2130, N2124, N1826);
nor NOR2 (N2131, N2127, N1881);
and AND3 (N2132, N2128, N781, N348);
nand NAND2 (N2133, N2132, N14);
nand NAND4 (N2134, N2110, N653, N2013, N377);
nand NAND3 (N2135, N2131, N201, N224);
buf BUF1 (N2136, N2115);
nand NAND2 (N2137, N2118, N241);
or OR4 (N2138, N2136, N268, N1175, N309);
nand NAND2 (N2139, N2125, N532);
buf BUF1 (N2140, N2104);
xor XOR2 (N2141, N2130, N519);
nand NAND3 (N2142, N2129, N116, N2122);
or OR4 (N2143, N2134, N1804, N16, N90);
or OR4 (N2144, N2140, N1564, N1725, N271);
not NOT1 (N2145, N2142);
and AND4 (N2146, N2139, N151, N1260, N360);
xor XOR2 (N2147, N2138, N1355);
and AND3 (N2148, N2143, N1131, N972);
or OR3 (N2149, N2133, N1297, N18);
and AND2 (N2150, N2148, N464);
nor NOR2 (N2151, N2135, N264);
or OR4 (N2152, N2151, N1783, N797, N1119);
buf BUF1 (N2153, N2144);
buf BUF1 (N2154, N2150);
buf BUF1 (N2155, N2153);
xor XOR2 (N2156, N2123, N1319);
not NOT1 (N2157, N2154);
and AND4 (N2158, N2145, N1609, N388, N1655);
not NOT1 (N2159, N2141);
not NOT1 (N2160, N2159);
not NOT1 (N2161, N2157);
not NOT1 (N2162, N2147);
and AND3 (N2163, N2156, N1309, N226);
or OR4 (N2164, N2149, N1150, N1200, N2103);
xor XOR2 (N2165, N2161, N1375);
or OR3 (N2166, N2152, N2040, N2049);
not NOT1 (N2167, N2164);
or OR4 (N2168, N2158, N711, N449, N1592);
nand NAND3 (N2169, N2146, N1886, N1281);
nor NOR4 (N2170, N2169, N1881, N101, N1220);
buf BUF1 (N2171, N2166);
nor NOR4 (N2172, N2170, N1676, N498, N1420);
and AND3 (N2173, N2172, N1689, N1246);
and AND3 (N2174, N2165, N392, N1126);
nand NAND3 (N2175, N2167, N984, N973);
not NOT1 (N2176, N2160);
buf BUF1 (N2177, N2171);
nor NOR4 (N2178, N2173, N668, N1897, N1072);
or OR3 (N2179, N2168, N1274, N430);
nor NOR2 (N2180, N2179, N595);
or OR4 (N2181, N2180, N1879, N2037, N584);
nor NOR3 (N2182, N2137, N1594, N574);
or OR4 (N2183, N2155, N470, N1904, N160);
nand NAND2 (N2184, N2178, N1542);
xor XOR2 (N2185, N2175, N1680);
nand NAND3 (N2186, N2177, N747, N1143);
not NOT1 (N2187, N2163);
or OR4 (N2188, N2174, N871, N1688, N1861);
and AND3 (N2189, N2183, N1517, N1777);
and AND2 (N2190, N2185, N1298);
xor XOR2 (N2191, N2182, N179);
nand NAND4 (N2192, N2189, N927, N2022, N848);
and AND4 (N2193, N2162, N1830, N604, N2173);
buf BUF1 (N2194, N2184);
nand NAND3 (N2195, N2192, N430, N722);
buf BUF1 (N2196, N2176);
xor XOR2 (N2197, N2186, N34);
not NOT1 (N2198, N2193);
not NOT1 (N2199, N2194);
xor XOR2 (N2200, N2187, N1609);
or OR3 (N2201, N2191, N946, N1929);
xor XOR2 (N2202, N2197, N496);
and AND3 (N2203, N2196, N1841, N1688);
and AND3 (N2204, N2202, N1712, N1337);
buf BUF1 (N2205, N2188);
or OR4 (N2206, N2190, N418, N2048, N1511);
nand NAND2 (N2207, N2204, N2014);
or OR4 (N2208, N2181, N837, N399, N995);
nand NAND3 (N2209, N2200, N308, N652);
or OR3 (N2210, N2209, N899, N1568);
not NOT1 (N2211, N2210);
buf BUF1 (N2212, N2208);
and AND2 (N2213, N2201, N1980);
and AND4 (N2214, N2195, N1781, N1590, N1601);
xor XOR2 (N2215, N2213, N1495);
xor XOR2 (N2216, N2215, N665);
nand NAND2 (N2217, N2206, N1721);
xor XOR2 (N2218, N2212, N226);
nand NAND2 (N2219, N2199, N1288);
not NOT1 (N2220, N2203);
buf BUF1 (N2221, N2219);
buf BUF1 (N2222, N2205);
and AND4 (N2223, N2220, N1141, N580, N1226);
and AND3 (N2224, N2216, N1720, N631);
nor NOR2 (N2225, N2211, N1878);
nand NAND2 (N2226, N2222, N1887);
not NOT1 (N2227, N2223);
nor NOR4 (N2228, N2226, N1947, N1214, N747);
not NOT1 (N2229, N2221);
or OR4 (N2230, N2198, N1028, N1863, N599);
and AND3 (N2231, N2229, N1664, N1886);
and AND4 (N2232, N2231, N1568, N44, N1716);
and AND4 (N2233, N2230, N332, N2162, N1871);
or OR2 (N2234, N2227, N2048);
nor NOR3 (N2235, N2228, N1814, N1465);
nor NOR2 (N2236, N2218, N1196);
nor NOR3 (N2237, N2235, N485, N1632);
or OR3 (N2238, N2225, N20, N960);
xor XOR2 (N2239, N2238, N1850);
nor NOR4 (N2240, N2233, N705, N879, N470);
xor XOR2 (N2241, N2232, N757);
nand NAND3 (N2242, N2214, N1292, N2138);
not NOT1 (N2243, N2240);
or OR3 (N2244, N2217, N1596, N1428);
and AND2 (N2245, N2243, N154);
not NOT1 (N2246, N2224);
nand NAND4 (N2247, N2234, N975, N1144, N1872);
nand NAND2 (N2248, N2247, N979);
not NOT1 (N2249, N2239);
or OR3 (N2250, N2249, N962, N1551);
xor XOR2 (N2251, N2237, N1131);
not NOT1 (N2252, N2207);
not NOT1 (N2253, N2236);
buf BUF1 (N2254, N2250);
nand NAND3 (N2255, N2254, N1772, N228);
and AND3 (N2256, N2252, N2108, N450);
nor NOR2 (N2257, N2253, N198);
xor XOR2 (N2258, N2256, N969);
not NOT1 (N2259, N2257);
or OR4 (N2260, N2251, N250, N382, N144);
buf BUF1 (N2261, N2241);
not NOT1 (N2262, N2246);
buf BUF1 (N2263, N2260);
nor NOR4 (N2264, N2259, N1660, N103, N1353);
nand NAND3 (N2265, N2262, N542, N988);
and AND4 (N2266, N2248, N574, N1913, N83);
and AND3 (N2267, N2255, N748, N515);
buf BUF1 (N2268, N2245);
or OR4 (N2269, N2244, N2011, N1803, N227);
not NOT1 (N2270, N2265);
xor XOR2 (N2271, N2263, N1248);
buf BUF1 (N2272, N2242);
or OR3 (N2273, N2271, N1389, N1234);
not NOT1 (N2274, N2269);
or OR2 (N2275, N2264, N1228);
xor XOR2 (N2276, N2270, N770);
not NOT1 (N2277, N2272);
nand NAND2 (N2278, N2261, N106);
buf BUF1 (N2279, N2258);
nand NAND4 (N2280, N2266, N807, N2168, N2138);
not NOT1 (N2281, N2268);
or OR4 (N2282, N2279, N1947, N1488, N278);
not NOT1 (N2283, N2277);
not NOT1 (N2284, N2275);
buf BUF1 (N2285, N2276);
nand NAND4 (N2286, N2284, N1337, N1514, N1424);
nor NOR3 (N2287, N2267, N1941, N119);
xor XOR2 (N2288, N2287, N150);
or OR4 (N2289, N2281, N962, N1123, N989);
or OR2 (N2290, N2280, N1642);
or OR4 (N2291, N2282, N824, N1080, N1091);
or OR3 (N2292, N2288, N199, N347);
not NOT1 (N2293, N2278);
or OR3 (N2294, N2273, N1759, N829);
or OR2 (N2295, N2289, N1806);
and AND2 (N2296, N2286, N1321);
or OR4 (N2297, N2290, N376, N391, N892);
not NOT1 (N2298, N2283);
nand NAND2 (N2299, N2293, N499);
and AND2 (N2300, N2297, N687);
or OR3 (N2301, N2295, N2176, N1750);
xor XOR2 (N2302, N2296, N1584);
and AND3 (N2303, N2301, N2071, N824);
xor XOR2 (N2304, N2294, N1715);
or OR4 (N2305, N2291, N1912, N1817, N1348);
nand NAND3 (N2306, N2304, N1688, N1776);
xor XOR2 (N2307, N2303, N1289);
nand NAND3 (N2308, N2292, N916, N851);
nand NAND3 (N2309, N2274, N1847, N254);
and AND3 (N2310, N2306, N1574, N726);
xor XOR2 (N2311, N2300, N1651);
nor NOR4 (N2312, N2310, N2277, N493, N1401);
not NOT1 (N2313, N2308);
buf BUF1 (N2314, N2312);
buf BUF1 (N2315, N2313);
nand NAND3 (N2316, N2302, N211, N1838);
nand NAND2 (N2317, N2298, N2307);
buf BUF1 (N2318, N1314);
nor NOR3 (N2319, N2311, N313, N2052);
or OR2 (N2320, N2309, N1961);
and AND2 (N2321, N2318, N21);
nand NAND4 (N2322, N2320, N381, N1518, N2309);
nand NAND4 (N2323, N2321, N735, N822, N1378);
or OR4 (N2324, N2314, N212, N1367, N2002);
not NOT1 (N2325, N2315);
nand NAND3 (N2326, N2317, N566, N1017);
or OR4 (N2327, N2326, N595, N1943, N1050);
buf BUF1 (N2328, N2322);
nand NAND3 (N2329, N2305, N2062, N1665);
and AND2 (N2330, N2328, N869);
and AND2 (N2331, N2323, N2304);
buf BUF1 (N2332, N2331);
nand NAND3 (N2333, N2316, N340, N1751);
xor XOR2 (N2334, N2329, N2160);
nor NOR3 (N2335, N2332, N2280, N540);
or OR4 (N2336, N2324, N177, N1235, N25);
or OR4 (N2337, N2299, N1856, N332, N1636);
not NOT1 (N2338, N2335);
buf BUF1 (N2339, N2327);
nor NOR4 (N2340, N2336, N440, N2038, N879);
and AND3 (N2341, N2334, N2311, N1238);
or OR2 (N2342, N2341, N1553);
buf BUF1 (N2343, N2340);
nor NOR2 (N2344, N2330, N596);
xor XOR2 (N2345, N2337, N2172);
nand NAND2 (N2346, N2342, N296);
xor XOR2 (N2347, N2343, N1408);
xor XOR2 (N2348, N2339, N2246);
or OR4 (N2349, N2348, N2337, N195, N110);
nand NAND3 (N2350, N2347, N1182, N863);
xor XOR2 (N2351, N2319, N1301);
xor XOR2 (N2352, N2344, N1763);
buf BUF1 (N2353, N2333);
nor NOR2 (N2354, N2351, N98);
buf BUF1 (N2355, N2350);
nor NOR4 (N2356, N2355, N1398, N2132, N548);
and AND2 (N2357, N2325, N533);
not NOT1 (N2358, N2346);
nor NOR3 (N2359, N2349, N1484, N1950);
not NOT1 (N2360, N2345);
xor XOR2 (N2361, N2358, N1762);
or OR2 (N2362, N2353, N2217);
or OR4 (N2363, N2357, N209, N1099, N241);
xor XOR2 (N2364, N2352, N698);
nor NOR3 (N2365, N2360, N706, N359);
or OR4 (N2366, N2356, N1203, N104, N1869);
nand NAND3 (N2367, N2362, N655, N1886);
or OR3 (N2368, N2364, N1257, N1696);
and AND2 (N2369, N2367, N266);
buf BUF1 (N2370, N2359);
not NOT1 (N2371, N2338);
buf BUF1 (N2372, N2365);
nand NAND2 (N2373, N2369, N1280);
nor NOR2 (N2374, N2370, N1400);
xor XOR2 (N2375, N2374, N864);
and AND2 (N2376, N2354, N261);
buf BUF1 (N2377, N2371);
or OR3 (N2378, N2361, N1117, N1333);
xor XOR2 (N2379, N2363, N1639);
or OR4 (N2380, N2375, N1954, N2330, N778);
nand NAND2 (N2381, N2377, N1860);
and AND3 (N2382, N2372, N1965, N1539);
nor NOR3 (N2383, N2381, N1203, N1639);
nand NAND3 (N2384, N2379, N1939, N775);
nor NOR4 (N2385, N2285, N597, N468, N2308);
nor NOR3 (N2386, N2383, N1769, N860);
not NOT1 (N2387, N2378);
or OR3 (N2388, N2380, N1907, N351);
nor NOR2 (N2389, N2373, N1188);
and AND3 (N2390, N2388, N665, N2171);
not NOT1 (N2391, N2387);
nand NAND3 (N2392, N2368, N1484, N20);
not NOT1 (N2393, N2384);
xor XOR2 (N2394, N2386, N640);
not NOT1 (N2395, N2393);
xor XOR2 (N2396, N2389, N1029);
nand NAND4 (N2397, N2391, N694, N2116, N1882);
nand NAND3 (N2398, N2395, N181, N1774);
xor XOR2 (N2399, N2376, N1550);
nor NOR4 (N2400, N2390, N353, N382, N1666);
not NOT1 (N2401, N2396);
nand NAND4 (N2402, N2398, N2102, N2199, N1108);
xor XOR2 (N2403, N2402, N1197);
and AND4 (N2404, N2385, N1226, N2108, N349);
nor NOR2 (N2405, N2404, N974);
and AND2 (N2406, N2405, N1802);
and AND2 (N2407, N2399, N282);
nand NAND4 (N2408, N2397, N849, N1998, N419);
or OR3 (N2409, N2408, N251, N1035);
not NOT1 (N2410, N2394);
nand NAND3 (N2411, N2401, N295, N809);
nor NOR3 (N2412, N2382, N1255, N268);
nor NOR3 (N2413, N2403, N317, N2248);
not NOT1 (N2414, N2412);
nor NOR3 (N2415, N2411, N1072, N2187);
buf BUF1 (N2416, N2414);
or OR4 (N2417, N2415, N1701, N1896, N1839);
buf BUF1 (N2418, N2417);
and AND3 (N2419, N2392, N343, N645);
nand NAND2 (N2420, N2407, N1336);
nand NAND3 (N2421, N2418, N806, N690);
and AND3 (N2422, N2410, N964, N380);
nor NOR2 (N2423, N2416, N659);
nand NAND2 (N2424, N2406, N912);
xor XOR2 (N2425, N2422, N613);
nor NOR2 (N2426, N2420, N1464);
and AND4 (N2427, N2421, N1764, N172, N2201);
buf BUF1 (N2428, N2366);
xor XOR2 (N2429, N2423, N1797);
not NOT1 (N2430, N2419);
nand NAND3 (N2431, N2426, N1162, N972);
and AND4 (N2432, N2429, N576, N219, N1337);
not NOT1 (N2433, N2400);
and AND3 (N2434, N2425, N2233, N1220);
and AND4 (N2435, N2432, N2238, N480, N1364);
xor XOR2 (N2436, N2434, N2386);
buf BUF1 (N2437, N2428);
buf BUF1 (N2438, N2427);
nor NOR2 (N2439, N2431, N2306);
not NOT1 (N2440, N2409);
xor XOR2 (N2441, N2413, N110);
nor NOR4 (N2442, N2437, N352, N1973, N807);
not NOT1 (N2443, N2442);
buf BUF1 (N2444, N2443);
or OR4 (N2445, N2430, N2265, N1610, N542);
nor NOR2 (N2446, N2436, N109);
or OR2 (N2447, N2439, N320);
xor XOR2 (N2448, N2441, N2179);
nor NOR2 (N2449, N2440, N1712);
buf BUF1 (N2450, N2424);
nor NOR3 (N2451, N2445, N11, N590);
xor XOR2 (N2452, N2449, N1260);
not NOT1 (N2453, N2452);
nand NAND4 (N2454, N2435, N150, N624, N1013);
or OR2 (N2455, N2444, N1010);
xor XOR2 (N2456, N2453, N2310);
and AND3 (N2457, N2446, N2275, N1755);
buf BUF1 (N2458, N2447);
xor XOR2 (N2459, N2455, N1825);
nor NOR2 (N2460, N2459, N1745);
not NOT1 (N2461, N2460);
xor XOR2 (N2462, N2451, N54);
and AND2 (N2463, N2433, N432);
nor NOR4 (N2464, N2454, N2231, N1658, N1056);
or OR3 (N2465, N2461, N1721, N2355);
nor NOR2 (N2466, N2465, N315);
or OR4 (N2467, N2462, N1813, N1502, N1292);
buf BUF1 (N2468, N2438);
buf BUF1 (N2469, N2458);
not NOT1 (N2470, N2464);
and AND4 (N2471, N2470, N2408, N1349, N1908);
not NOT1 (N2472, N2463);
and AND3 (N2473, N2448, N668, N1685);
or OR4 (N2474, N2456, N844, N1564, N1164);
not NOT1 (N2475, N2450);
and AND3 (N2476, N2471, N947, N1262);
not NOT1 (N2477, N2468);
or OR2 (N2478, N2466, N819);
nand NAND3 (N2479, N2478, N1222, N734);
nor NOR4 (N2480, N2474, N1796, N1589, N2351);
nand NAND2 (N2481, N2476, N1157);
nand NAND4 (N2482, N2473, N1018, N1870, N2038);
or OR2 (N2483, N2467, N2408);
and AND2 (N2484, N2481, N1143);
buf BUF1 (N2485, N2472);
xor XOR2 (N2486, N2483, N2055);
buf BUF1 (N2487, N2477);
and AND3 (N2488, N2479, N1664, N1923);
buf BUF1 (N2489, N2482);
buf BUF1 (N2490, N2485);
or OR3 (N2491, N2484, N1795, N36);
nand NAND4 (N2492, N2469, N733, N300, N1963);
not NOT1 (N2493, N2489);
not NOT1 (N2494, N2480);
nand NAND3 (N2495, N2488, N895, N965);
and AND4 (N2496, N2486, N1307, N1605, N189);
or OR4 (N2497, N2496, N919, N482, N2469);
buf BUF1 (N2498, N2494);
nor NOR2 (N2499, N2487, N2293);
nand NAND4 (N2500, N2497, N1221, N2414, N619);
nor NOR2 (N2501, N2490, N1691);
nor NOR3 (N2502, N2493, N768, N227);
nand NAND4 (N2503, N2495, N1427, N807, N2331);
nand NAND2 (N2504, N2475, N956);
nor NOR4 (N2505, N2500, N1368, N1899, N1568);
buf BUF1 (N2506, N2504);
nor NOR4 (N2507, N2457, N2008, N2068, N1772);
not NOT1 (N2508, N2501);
nor NOR3 (N2509, N2502, N1776, N810);
and AND4 (N2510, N2499, N863, N438, N1620);
nand NAND2 (N2511, N2492, N2094);
or OR2 (N2512, N2509, N2509);
buf BUF1 (N2513, N2508);
xor XOR2 (N2514, N2503, N2415);
not NOT1 (N2515, N2507);
nand NAND4 (N2516, N2515, N2507, N1191, N1034);
nor NOR3 (N2517, N2498, N120, N1735);
nor NOR4 (N2518, N2512, N1214, N1577, N1109);
nor NOR3 (N2519, N2511, N2267, N11);
and AND3 (N2520, N2517, N2480, N2320);
not NOT1 (N2521, N2519);
or OR3 (N2522, N2491, N858, N1325);
xor XOR2 (N2523, N2522, N122);
or OR3 (N2524, N2516, N1531, N323);
xor XOR2 (N2525, N2518, N1140);
or OR2 (N2526, N2524, N860);
and AND2 (N2527, N2526, N1128);
xor XOR2 (N2528, N2513, N1918);
xor XOR2 (N2529, N2521, N1804);
not NOT1 (N2530, N2525);
nor NOR2 (N2531, N2506, N2484);
nand NAND3 (N2532, N2514, N1839, N232);
xor XOR2 (N2533, N2505, N2177);
not NOT1 (N2534, N2533);
or OR4 (N2535, N2532, N1338, N2228, N1568);
nand NAND4 (N2536, N2531, N1265, N279, N1166);
xor XOR2 (N2537, N2520, N585);
or OR4 (N2538, N2528, N2458, N2450, N537);
or OR2 (N2539, N2530, N875);
buf BUF1 (N2540, N2539);
or OR4 (N2541, N2529, N1019, N1278, N1649);
not NOT1 (N2542, N2523);
and AND4 (N2543, N2534, N1409, N8, N352);
nor NOR4 (N2544, N2510, N2489, N1407, N2340);
xor XOR2 (N2545, N2538, N897);
nor NOR2 (N2546, N2543, N1728);
not NOT1 (N2547, N2535);
xor XOR2 (N2548, N2546, N1055);
nand NAND4 (N2549, N2537, N2435, N423, N1098);
or OR2 (N2550, N2547, N1774);
xor XOR2 (N2551, N2527, N121);
and AND3 (N2552, N2541, N739, N465);
xor XOR2 (N2553, N2544, N1043);
nand NAND2 (N2554, N2553, N2428);
not NOT1 (N2555, N2536);
and AND2 (N2556, N2551, N1250);
and AND2 (N2557, N2556, N1046);
not NOT1 (N2558, N2549);
or OR4 (N2559, N2554, N2455, N1186, N196);
buf BUF1 (N2560, N2548);
or OR3 (N2561, N2560, N2244, N2375);
or OR2 (N2562, N2558, N2031);
or OR3 (N2563, N2545, N478, N1576);
xor XOR2 (N2564, N2561, N1796);
xor XOR2 (N2565, N2559, N1717);
nand NAND2 (N2566, N2550, N2099);
and AND2 (N2567, N2562, N1797);
buf BUF1 (N2568, N2557);
nand NAND4 (N2569, N2555, N1825, N157, N2366);
xor XOR2 (N2570, N2569, N2324);
nand NAND4 (N2571, N2568, N1516, N1285, N2401);
nor NOR4 (N2572, N2570, N348, N998, N1188);
and AND4 (N2573, N2563, N1431, N810, N1445);
or OR3 (N2574, N2542, N760, N113);
or OR2 (N2575, N2573, N1229);
or OR4 (N2576, N2564, N1438, N847, N348);
nand NAND4 (N2577, N2566, N677, N1860, N365);
buf BUF1 (N2578, N2574);
not NOT1 (N2579, N2567);
not NOT1 (N2580, N2540);
and AND4 (N2581, N2572, N1393, N100, N422);
xor XOR2 (N2582, N2579, N1038);
nor NOR2 (N2583, N2577, N1309);
or OR4 (N2584, N2552, N1639, N1170, N2067);
not NOT1 (N2585, N2580);
or OR2 (N2586, N2575, N704);
not NOT1 (N2587, N2581);
or OR4 (N2588, N2578, N1700, N1418, N1367);
not NOT1 (N2589, N2571);
buf BUF1 (N2590, N2576);
and AND2 (N2591, N2583, N1770);
nand NAND2 (N2592, N2582, N387);
and AND3 (N2593, N2591, N1926, N2460);
nand NAND2 (N2594, N2590, N1392);
xor XOR2 (N2595, N2593, N1520);
xor XOR2 (N2596, N2585, N2272);
xor XOR2 (N2597, N2565, N2312);
buf BUF1 (N2598, N2586);
buf BUF1 (N2599, N2589);
not NOT1 (N2600, N2584);
xor XOR2 (N2601, N2596, N971);
xor XOR2 (N2602, N2587, N832);
nand NAND4 (N2603, N2598, N1458, N1865, N744);
nor NOR4 (N2604, N2597, N833, N1474, N1660);
not NOT1 (N2605, N2599);
and AND2 (N2606, N2601, N1430);
nor NOR2 (N2607, N2605, N1900);
buf BUF1 (N2608, N2588);
xor XOR2 (N2609, N2595, N1829);
or OR4 (N2610, N2592, N1530, N653, N664);
xor XOR2 (N2611, N2608, N2075);
and AND4 (N2612, N2610, N1744, N72, N1202);
xor XOR2 (N2613, N2604, N494);
or OR2 (N2614, N2609, N1210);
and AND3 (N2615, N2602, N1264, N1103);
and AND2 (N2616, N2612, N2495);
or OR4 (N2617, N2594, N2427, N371, N901);
not NOT1 (N2618, N2606);
not NOT1 (N2619, N2611);
not NOT1 (N2620, N2615);
nor NOR2 (N2621, N2614, N1388);
xor XOR2 (N2622, N2619, N2014);
nand NAND3 (N2623, N2600, N190, N1484);
or OR3 (N2624, N2618, N758, N2423);
nor NOR4 (N2625, N2617, N445, N1229, N2196);
xor XOR2 (N2626, N2620, N165);
nand NAND3 (N2627, N2616, N2020, N823);
and AND4 (N2628, N2623, N2255, N155, N396);
and AND3 (N2629, N2627, N2588, N2386);
buf BUF1 (N2630, N2622);
and AND3 (N2631, N2613, N278, N331);
xor XOR2 (N2632, N2626, N236);
or OR4 (N2633, N2628, N1995, N2063, N2007);
not NOT1 (N2634, N2607);
buf BUF1 (N2635, N2625);
nor NOR4 (N2636, N2634, N2453, N2230, N2251);
and AND3 (N2637, N2629, N2253, N1541);
nand NAND3 (N2638, N2636, N1436, N1671);
buf BUF1 (N2639, N2635);
or OR4 (N2640, N2624, N1989, N2546, N609);
nor NOR4 (N2641, N2632, N794, N331, N863);
nor NOR2 (N2642, N2631, N1440);
or OR3 (N2643, N2638, N1540, N1662);
buf BUF1 (N2644, N2637);
buf BUF1 (N2645, N2643);
not NOT1 (N2646, N2645);
and AND4 (N2647, N2644, N1699, N1720, N276);
and AND3 (N2648, N2641, N1714, N1448);
not NOT1 (N2649, N2603);
nor NOR4 (N2650, N2649, N2418, N320, N231);
buf BUF1 (N2651, N2647);
nor NOR3 (N2652, N2633, N468, N2142);
nor NOR4 (N2653, N2650, N1632, N2302, N643);
not NOT1 (N2654, N2630);
nor NOR2 (N2655, N2621, N557);
nor NOR2 (N2656, N2640, N452);
and AND3 (N2657, N2652, N2507, N737);
nand NAND4 (N2658, N2657, N541, N662, N1552);
or OR2 (N2659, N2646, N2267);
not NOT1 (N2660, N2651);
not NOT1 (N2661, N2654);
or OR4 (N2662, N2648, N759, N250, N442);
or OR3 (N2663, N2655, N1790, N890);
xor XOR2 (N2664, N2642, N1038);
xor XOR2 (N2665, N2661, N618);
nand NAND2 (N2666, N2658, N1831);
or OR3 (N2667, N2656, N2423, N487);
and AND4 (N2668, N2667, N1098, N1823, N1170);
or OR3 (N2669, N2660, N7, N1804);
xor XOR2 (N2670, N2665, N217);
xor XOR2 (N2671, N2669, N2378);
xor XOR2 (N2672, N2671, N2323);
and AND3 (N2673, N2639, N153, N1819);
nand NAND3 (N2674, N2664, N1291, N2560);
nor NOR4 (N2675, N2673, N597, N1403, N2305);
and AND3 (N2676, N2666, N2124, N2420);
and AND3 (N2677, N2676, N331, N216);
nand NAND2 (N2678, N2672, N1844);
or OR4 (N2679, N2674, N1120, N1456, N2573);
nand NAND4 (N2680, N2663, N2670, N1158, N124);
nand NAND4 (N2681, N2581, N2527, N351, N417);
nor NOR3 (N2682, N2653, N1120, N924);
buf BUF1 (N2683, N2679);
xor XOR2 (N2684, N2677, N1987);
or OR2 (N2685, N2678, N2020);
buf BUF1 (N2686, N2675);
not NOT1 (N2687, N2686);
or OR4 (N2688, N2681, N1076, N1678, N383);
nor NOR2 (N2689, N2662, N2020);
not NOT1 (N2690, N2685);
buf BUF1 (N2691, N2668);
not NOT1 (N2692, N2691);
nand NAND3 (N2693, N2690, N1192, N607);
nor NOR2 (N2694, N2687, N21);
and AND3 (N2695, N2688, N52, N818);
not NOT1 (N2696, N2680);
nor NOR2 (N2697, N2659, N1082);
not NOT1 (N2698, N2682);
and AND3 (N2699, N2684, N694, N2529);
nor NOR3 (N2700, N2689, N1749, N2680);
xor XOR2 (N2701, N2697, N1867);
nor NOR4 (N2702, N2701, N1730, N1545, N2664);
xor XOR2 (N2703, N2694, N1117);
nand NAND3 (N2704, N2700, N1833, N884);
nand NAND3 (N2705, N2692, N2524, N540);
buf BUF1 (N2706, N2702);
xor XOR2 (N2707, N2706, N2689);
xor XOR2 (N2708, N2705, N2561);
and AND2 (N2709, N2695, N1469);
nand NAND2 (N2710, N2704, N1759);
not NOT1 (N2711, N2707);
or OR2 (N2712, N2683, N1776);
xor XOR2 (N2713, N2699, N365);
buf BUF1 (N2714, N2712);
nand NAND2 (N2715, N2693, N2680);
and AND2 (N2716, N2714, N103);
and AND4 (N2717, N2716, N1806, N37, N2029);
nor NOR4 (N2718, N2708, N989, N64, N2508);
xor XOR2 (N2719, N2713, N1360);
xor XOR2 (N2720, N2717, N2022);
or OR3 (N2721, N2720, N2476, N948);
buf BUF1 (N2722, N2711);
nand NAND4 (N2723, N2698, N574, N1806, N222);
or OR4 (N2724, N2696, N2091, N1575, N1180);
buf BUF1 (N2725, N2722);
nor NOR3 (N2726, N2710, N2586, N2038);
nor NOR3 (N2727, N2721, N1564, N2472);
and AND4 (N2728, N2719, N1662, N240, N1742);
buf BUF1 (N2729, N2728);
and AND4 (N2730, N2703, N2290, N93, N616);
not NOT1 (N2731, N2715);
and AND3 (N2732, N2729, N2467, N710);
or OR3 (N2733, N2724, N418, N1670);
buf BUF1 (N2734, N2709);
buf BUF1 (N2735, N2732);
xor XOR2 (N2736, N2727, N27);
not NOT1 (N2737, N2730);
not NOT1 (N2738, N2718);
buf BUF1 (N2739, N2737);
or OR4 (N2740, N2733, N1896, N1990, N2488);
nor NOR2 (N2741, N2734, N2183);
not NOT1 (N2742, N2735);
or OR4 (N2743, N2726, N233, N2200, N1317);
xor XOR2 (N2744, N2741, N16);
nand NAND3 (N2745, N2740, N1108, N329);
nand NAND3 (N2746, N2743, N2502, N1795);
xor XOR2 (N2747, N2742, N490);
not NOT1 (N2748, N2745);
and AND3 (N2749, N2723, N2208, N37);
xor XOR2 (N2750, N2736, N283);
nor NOR4 (N2751, N2725, N1761, N788, N1332);
buf BUF1 (N2752, N2744);
xor XOR2 (N2753, N2747, N1631);
xor XOR2 (N2754, N2731, N1907);
and AND4 (N2755, N2748, N879, N2152, N1818);
xor XOR2 (N2756, N2754, N1053);
xor XOR2 (N2757, N2755, N2299);
not NOT1 (N2758, N2749);
or OR3 (N2759, N2757, N916, N487);
buf BUF1 (N2760, N2752);
buf BUF1 (N2761, N2751);
or OR3 (N2762, N2758, N1515, N151);
or OR4 (N2763, N2738, N2035, N92, N902);
not NOT1 (N2764, N2750);
buf BUF1 (N2765, N2764);
buf BUF1 (N2766, N2761);
and AND4 (N2767, N2762, N2315, N86, N1828);
not NOT1 (N2768, N2739);
xor XOR2 (N2769, N2753, N2538);
nand NAND4 (N2770, N2766, N1767, N2089, N422);
buf BUF1 (N2771, N2759);
and AND3 (N2772, N2767, N867, N2627);
or OR3 (N2773, N2756, N1708, N1766);
nor NOR3 (N2774, N2769, N2422, N1210);
not NOT1 (N2775, N2746);
nand NAND2 (N2776, N2765, N2708);
or OR3 (N2777, N2760, N2038, N1620);
nand NAND4 (N2778, N2770, N1447, N2758, N303);
or OR3 (N2779, N2778, N1216, N2657);
and AND2 (N2780, N2775, N1300);
nand NAND3 (N2781, N2768, N2610, N138);
and AND3 (N2782, N2772, N643, N597);
and AND4 (N2783, N2774, N209, N420, N1305);
nand NAND3 (N2784, N2776, N30, N786);
xor XOR2 (N2785, N2782, N1053);
nor NOR4 (N2786, N2771, N1248, N1420, N2241);
nor NOR2 (N2787, N2783, N1737);
xor XOR2 (N2788, N2784, N2174);
and AND4 (N2789, N2773, N247, N766, N327);
or OR4 (N2790, N2787, N560, N1122, N910);
or OR4 (N2791, N2781, N56, N1134, N931);
nand NAND2 (N2792, N2790, N667);
nor NOR4 (N2793, N2791, N83, N2471, N778);
not NOT1 (N2794, N2789);
nand NAND3 (N2795, N2779, N433, N302);
xor XOR2 (N2796, N2793, N1849);
not NOT1 (N2797, N2780);
buf BUF1 (N2798, N2795);
or OR4 (N2799, N2794, N2592, N1549, N1463);
nor NOR3 (N2800, N2797, N435, N1266);
nand NAND4 (N2801, N2777, N2101, N2467, N655);
nand NAND4 (N2802, N2798, N2470, N2446, N2416);
xor XOR2 (N2803, N2785, N1538);
xor XOR2 (N2804, N2763, N900);
buf BUF1 (N2805, N2792);
buf BUF1 (N2806, N2786);
or OR4 (N2807, N2803, N39, N2753, N2036);
buf BUF1 (N2808, N2801);
nor NOR4 (N2809, N2800, N866, N1604, N2731);
not NOT1 (N2810, N2796);
nor NOR3 (N2811, N2805, N1971, N499);
buf BUF1 (N2812, N2808);
nand NAND4 (N2813, N2804, N757, N678, N1401);
nand NAND2 (N2814, N2802, N2753);
buf BUF1 (N2815, N2813);
and AND4 (N2816, N2799, N1338, N2623, N1799);
nor NOR4 (N2817, N2807, N2090, N1941, N435);
buf BUF1 (N2818, N2788);
nand NAND4 (N2819, N2818, N1617, N2313, N1441);
nand NAND2 (N2820, N2812, N35);
nor NOR3 (N2821, N2806, N2463, N1440);
and AND2 (N2822, N2809, N1067);
xor XOR2 (N2823, N2819, N2612);
not NOT1 (N2824, N2810);
or OR2 (N2825, N2824, N1065);
not NOT1 (N2826, N2820);
buf BUF1 (N2827, N2823);
nor NOR3 (N2828, N2822, N2731, N1541);
nand NAND4 (N2829, N2816, N243, N2305, N683);
buf BUF1 (N2830, N2829);
nand NAND2 (N2831, N2815, N2078);
or OR2 (N2832, N2825, N69);
buf BUF1 (N2833, N2830);
buf BUF1 (N2834, N2833);
xor XOR2 (N2835, N2814, N2139);
not NOT1 (N2836, N2811);
and AND2 (N2837, N2835, N1746);
or OR4 (N2838, N2826, N1573, N875, N990);
or OR3 (N2839, N2831, N357, N2355);
and AND3 (N2840, N2827, N737, N162);
or OR4 (N2841, N2821, N705, N2291, N607);
or OR4 (N2842, N2838, N136, N1073, N1087);
not NOT1 (N2843, N2836);
nand NAND2 (N2844, N2843, N806);
nand NAND3 (N2845, N2837, N2117, N848);
not NOT1 (N2846, N2828);
buf BUF1 (N2847, N2845);
buf BUF1 (N2848, N2841);
or OR4 (N2849, N2844, N968, N1153, N1045);
not NOT1 (N2850, N2817);
nor NOR3 (N2851, N2849, N1611, N189);
or OR4 (N2852, N2834, N439, N1528, N2325);
xor XOR2 (N2853, N2847, N1928);
nand NAND4 (N2854, N2842, N1245, N1605, N2219);
not NOT1 (N2855, N2854);
and AND3 (N2856, N2840, N1651, N2066);
nand NAND2 (N2857, N2832, N818);
nor NOR3 (N2858, N2855, N2029, N1044);
buf BUF1 (N2859, N2848);
xor XOR2 (N2860, N2856, N1704);
nand NAND4 (N2861, N2846, N1661, N2117, N2813);
nand NAND2 (N2862, N2860, N360);
or OR2 (N2863, N2852, N872);
not NOT1 (N2864, N2861);
nor NOR2 (N2865, N2863, N1665);
not NOT1 (N2866, N2862);
not NOT1 (N2867, N2864);
and AND2 (N2868, N2857, N1191);
nor NOR3 (N2869, N2853, N1738, N389);
nor NOR4 (N2870, N2859, N2739, N120, N2822);
xor XOR2 (N2871, N2867, N1300);
nor NOR4 (N2872, N2839, N428, N1219, N368);
and AND3 (N2873, N2869, N1562, N144);
or OR2 (N2874, N2868, N1148);
not NOT1 (N2875, N2866);
xor XOR2 (N2876, N2872, N245);
nand NAND3 (N2877, N2871, N1587, N2172);
xor XOR2 (N2878, N2875, N2144);
nor NOR3 (N2879, N2874, N841, N1572);
or OR2 (N2880, N2858, N2743);
not NOT1 (N2881, N2870);
xor XOR2 (N2882, N2877, N1575);
not NOT1 (N2883, N2851);
xor XOR2 (N2884, N2881, N197);
not NOT1 (N2885, N2878);
nand NAND4 (N2886, N2882, N1459, N448, N2415);
and AND3 (N2887, N2876, N545, N187);
nor NOR4 (N2888, N2883, N1840, N2469, N247);
nor NOR4 (N2889, N2880, N2074, N2020, N99);
nand NAND3 (N2890, N2885, N2333, N1730);
and AND4 (N2891, N2873, N182, N2718, N2222);
not NOT1 (N2892, N2888);
not NOT1 (N2893, N2891);
nand NAND3 (N2894, N2879, N2135, N982);
nand NAND3 (N2895, N2865, N1862, N1327);
not NOT1 (N2896, N2892);
or OR3 (N2897, N2893, N2616, N2103);
and AND2 (N2898, N2850, N38);
nand NAND4 (N2899, N2889, N1599, N1872, N2513);
and AND2 (N2900, N2897, N1692);
or OR3 (N2901, N2896, N2119, N2839);
buf BUF1 (N2902, N2899);
or OR4 (N2903, N2886, N1673, N2660, N531);
not NOT1 (N2904, N2898);
not NOT1 (N2905, N2903);
xor XOR2 (N2906, N2894, N174);
buf BUF1 (N2907, N2900);
nand NAND2 (N2908, N2895, N663);
xor XOR2 (N2909, N2884, N2233);
nand NAND3 (N2910, N2890, N2211, N1402);
nand NAND4 (N2911, N2908, N345, N2794, N1892);
and AND2 (N2912, N2887, N1724);
buf BUF1 (N2913, N2906);
xor XOR2 (N2914, N2905, N636);
nor NOR4 (N2915, N2909, N1511, N2749, N436);
buf BUF1 (N2916, N2915);
and AND4 (N2917, N2916, N2698, N218, N2130);
or OR4 (N2918, N2901, N1367, N198, N838);
not NOT1 (N2919, N2902);
nand NAND4 (N2920, N2907, N157, N2609, N550);
nor NOR4 (N2921, N2910, N470, N1255, N1847);
xor XOR2 (N2922, N2914, N528);
nor NOR4 (N2923, N2922, N519, N1529, N2079);
nor NOR4 (N2924, N2904, N748, N309, N1150);
xor XOR2 (N2925, N2924, N2046);
buf BUF1 (N2926, N2912);
or OR4 (N2927, N2921, N1880, N1257, N166);
not NOT1 (N2928, N2923);
or OR2 (N2929, N2926, N1838);
xor XOR2 (N2930, N2919, N424);
or OR4 (N2931, N2911, N1354, N1748, N607);
xor XOR2 (N2932, N2927, N2092);
nor NOR4 (N2933, N2930, N101, N1465, N460);
and AND3 (N2934, N2933, N1992, N631);
not NOT1 (N2935, N2917);
not NOT1 (N2936, N2929);
not NOT1 (N2937, N2935);
not NOT1 (N2938, N2928);
nor NOR4 (N2939, N2913, N1401, N1692, N1173);
nor NOR2 (N2940, N2932, N1921);
nor NOR4 (N2941, N2934, N2118, N2633, N2436);
nand NAND4 (N2942, N2925, N1047, N2303, N1622);
not NOT1 (N2943, N2939);
nor NOR4 (N2944, N2941, N1, N153, N2698);
nor NOR3 (N2945, N2938, N1253, N1479);
not NOT1 (N2946, N2937);
xor XOR2 (N2947, N2946, N2179);
xor XOR2 (N2948, N2931, N856);
and AND4 (N2949, N2944, N188, N247, N2063);
or OR4 (N2950, N2940, N2093, N550, N965);
buf BUF1 (N2951, N2918);
xor XOR2 (N2952, N2947, N2012);
not NOT1 (N2953, N2950);
nand NAND2 (N2954, N2948, N2049);
nor NOR4 (N2955, N2953, N2460, N2536, N1490);
nor NOR4 (N2956, N2951, N1279, N102, N174);
nor NOR4 (N2957, N2942, N1501, N260, N2768);
nand NAND2 (N2958, N2954, N128);
xor XOR2 (N2959, N2956, N1484);
buf BUF1 (N2960, N2959);
nor NOR4 (N2961, N2957, N635, N2231, N1647);
nor NOR4 (N2962, N2952, N1523, N371, N2297);
xor XOR2 (N2963, N2949, N63);
xor XOR2 (N2964, N2943, N1169);
not NOT1 (N2965, N2960);
not NOT1 (N2966, N2920);
not NOT1 (N2967, N2958);
or OR2 (N2968, N2963, N219);
xor XOR2 (N2969, N2961, N2473);
nand NAND2 (N2970, N2965, N1815);
and AND4 (N2971, N2936, N1694, N2630, N909);
xor XOR2 (N2972, N2967, N1973);
nor NOR3 (N2973, N2966, N2425, N1061);
buf BUF1 (N2974, N2973);
or OR3 (N2975, N2968, N1096, N2596);
and AND4 (N2976, N2975, N744, N712, N2354);
nand NAND3 (N2977, N2969, N2759, N2403);
nand NAND3 (N2978, N2972, N299, N1135);
and AND4 (N2979, N2974, N2159, N215, N2692);
xor XOR2 (N2980, N2978, N105);
nand NAND2 (N2981, N2955, N121);
nor NOR2 (N2982, N2977, N1984);
or OR4 (N2983, N2979, N1100, N890, N976);
or OR3 (N2984, N2982, N2750, N439);
buf BUF1 (N2985, N2945);
nor NOR3 (N2986, N2976, N1049, N2485);
not NOT1 (N2987, N2962);
and AND4 (N2988, N2971, N2325, N1862, N826);
and AND3 (N2989, N2985, N1471, N852);
xor XOR2 (N2990, N2983, N2553);
nand NAND2 (N2991, N2988, N1175);
not NOT1 (N2992, N2964);
xor XOR2 (N2993, N2984, N706);
buf BUF1 (N2994, N2993);
and AND2 (N2995, N2989, N2306);
and AND2 (N2996, N2991, N2201);
xor XOR2 (N2997, N2990, N2194);
nand NAND3 (N2998, N2987, N2357, N2613);
nand NAND3 (N2999, N2981, N1611, N2599);
nand NAND2 (N3000, N2999, N2268);
and AND3 (N3001, N2998, N548, N2114);
nor NOR4 (N3002, N3001, N1291, N1219, N400);
or OR3 (N3003, N2992, N2814, N1664);
nand NAND3 (N3004, N2980, N767, N948);
not NOT1 (N3005, N3003);
or OR4 (N3006, N3005, N2023, N238, N1109);
not NOT1 (N3007, N2970);
not NOT1 (N3008, N2996);
nand NAND3 (N3009, N3004, N1529, N1769);
nand NAND4 (N3010, N3006, N1305, N45, N1824);
and AND3 (N3011, N2986, N19, N1777);
nand NAND2 (N3012, N3007, N855);
and AND4 (N3013, N2995, N1191, N2404, N2247);
buf BUF1 (N3014, N3013);
nor NOR4 (N3015, N2994, N2853, N1685, N52);
not NOT1 (N3016, N3000);
nand NAND4 (N3017, N3002, N1797, N1847, N907);
or OR4 (N3018, N3016, N1561, N1255, N2856);
or OR3 (N3019, N3015, N2746, N471);
nor NOR2 (N3020, N3011, N2312);
and AND3 (N3021, N2997, N2911, N1206);
buf BUF1 (N3022, N3010);
or OR4 (N3023, N3017, N2557, N2151, N585);
or OR4 (N3024, N3012, N816, N1552, N1038);
xor XOR2 (N3025, N3014, N2835);
buf BUF1 (N3026, N3019);
nor NOR4 (N3027, N3023, N586, N17, N1569);
or OR4 (N3028, N3021, N54, N2035, N2105);
or OR3 (N3029, N3008, N2903, N1944);
nand NAND4 (N3030, N3025, N605, N245, N249);
buf BUF1 (N3031, N3027);
and AND2 (N3032, N3020, N1929);
buf BUF1 (N3033, N3029);
nor NOR3 (N3034, N3022, N641, N1141);
nand NAND3 (N3035, N3034, N561, N2896);
and AND2 (N3036, N3024, N219);
buf BUF1 (N3037, N3032);
not NOT1 (N3038, N3037);
nor NOR3 (N3039, N3028, N1149, N2086);
nor NOR2 (N3040, N3035, N2368);
or OR2 (N3041, N3030, N1925);
and AND2 (N3042, N3038, N1464);
buf BUF1 (N3043, N3036);
buf BUF1 (N3044, N3033);
buf BUF1 (N3045, N3009);
not NOT1 (N3046, N3045);
buf BUF1 (N3047, N3044);
and AND3 (N3048, N3046, N1394, N851);
xor XOR2 (N3049, N3047, N2057);
buf BUF1 (N3050, N3031);
or OR4 (N3051, N3049, N2514, N1901, N3049);
not NOT1 (N3052, N3048);
or OR3 (N3053, N3042, N727, N1911);
xor XOR2 (N3054, N3052, N2780);
and AND3 (N3055, N3018, N796, N594);
and AND4 (N3056, N3026, N2481, N614, N116);
nor NOR2 (N3057, N3051, N2797);
buf BUF1 (N3058, N3057);
xor XOR2 (N3059, N3054, N1492);
not NOT1 (N3060, N3040);
not NOT1 (N3061, N3059);
and AND4 (N3062, N3058, N2520, N695, N413);
xor XOR2 (N3063, N3043, N605);
nand NAND3 (N3064, N3060, N1570, N2419);
not NOT1 (N3065, N3062);
nor NOR2 (N3066, N3055, N2295);
and AND2 (N3067, N3050, N862);
nor NOR3 (N3068, N3066, N2722, N1300);
and AND4 (N3069, N3065, N1398, N2925, N1364);
nand NAND3 (N3070, N3068, N1914, N997);
buf BUF1 (N3071, N3041);
buf BUF1 (N3072, N3056);
nor NOR3 (N3073, N3072, N382, N1427);
xor XOR2 (N3074, N3069, N2348);
nand NAND2 (N3075, N3064, N376);
not NOT1 (N3076, N3075);
and AND2 (N3077, N3063, N2959);
nand NAND3 (N3078, N3073, N2115, N692);
nor NOR2 (N3079, N3039, N486);
and AND4 (N3080, N3074, N972, N267, N991);
or OR3 (N3081, N3078, N1837, N556);
xor XOR2 (N3082, N3081, N3064);
nand NAND2 (N3083, N3077, N1758);
nand NAND4 (N3084, N3080, N2923, N936, N2902);
and AND3 (N3085, N3083, N182, N1048);
buf BUF1 (N3086, N3079);
and AND3 (N3087, N3067, N617, N1213);
buf BUF1 (N3088, N3071);
or OR2 (N3089, N3085, N1442);
and AND2 (N3090, N3053, N575);
or OR2 (N3091, N3087, N827);
nor NOR2 (N3092, N3061, N1259);
buf BUF1 (N3093, N3070);
and AND3 (N3094, N3092, N974, N2450);
or OR2 (N3095, N3094, N1698);
nor NOR2 (N3096, N3091, N1793);
and AND4 (N3097, N3076, N2476, N1693, N2816);
nor NOR4 (N3098, N3093, N1195, N2291, N1057);
not NOT1 (N3099, N3086);
and AND2 (N3100, N3095, N3024);
nand NAND3 (N3101, N3089, N2825, N504);
xor XOR2 (N3102, N3084, N1484);
and AND2 (N3103, N3088, N2019);
nor NOR4 (N3104, N3103, N3090, N1569, N1400);
nand NAND3 (N3105, N1863, N2550, N738);
buf BUF1 (N3106, N3096);
buf BUF1 (N3107, N3100);
or OR3 (N3108, N3097, N1310, N2065);
buf BUF1 (N3109, N3108);
and AND4 (N3110, N3102, N2122, N1549, N1566);
nand NAND2 (N3111, N3106, N464);
not NOT1 (N3112, N3109);
nand NAND2 (N3113, N3111, N473);
not NOT1 (N3114, N3082);
buf BUF1 (N3115, N3098);
not NOT1 (N3116, N3107);
not NOT1 (N3117, N3099);
or OR4 (N3118, N3116, N2665, N2525, N492);
nand NAND2 (N3119, N3112, N2920);
or OR2 (N3120, N3115, N1743);
nand NAND2 (N3121, N3118, N1289);
or OR4 (N3122, N3113, N748, N1043, N1311);
not NOT1 (N3123, N3104);
buf BUF1 (N3124, N3120);
and AND4 (N3125, N3105, N2134, N3028, N2610);
or OR3 (N3126, N3101, N820, N2163);
xor XOR2 (N3127, N3119, N978);
nor NOR3 (N3128, N3126, N1039, N1047);
buf BUF1 (N3129, N3121);
nor NOR4 (N3130, N3123, N1851, N44, N2683);
nor NOR2 (N3131, N3125, N2577);
and AND4 (N3132, N3127, N2938, N422, N287);
nor NOR2 (N3133, N3110, N2423);
not NOT1 (N3134, N3122);
and AND2 (N3135, N3114, N2296);
or OR2 (N3136, N3128, N721);
buf BUF1 (N3137, N3130);
nand NAND4 (N3138, N3129, N1306, N298, N2831);
nand NAND2 (N3139, N3124, N2515);
xor XOR2 (N3140, N3134, N1525);
nand NAND3 (N3141, N3137, N2272, N1087);
or OR4 (N3142, N3139, N1658, N1143, N2697);
not NOT1 (N3143, N3140);
and AND3 (N3144, N3141, N975, N188);
not NOT1 (N3145, N3143);
nand NAND4 (N3146, N3135, N3018, N1133, N3078);
and AND3 (N3147, N3142, N2178, N1630);
xor XOR2 (N3148, N3146, N2244);
xor XOR2 (N3149, N3148, N881);
xor XOR2 (N3150, N3138, N556);
and AND2 (N3151, N3145, N2606);
not NOT1 (N3152, N3144);
or OR3 (N3153, N3152, N807, N2992);
buf BUF1 (N3154, N3153);
or OR3 (N3155, N3132, N1132, N2607);
nand NAND2 (N3156, N3149, N1050);
or OR2 (N3157, N3151, N2521);
nand NAND3 (N3158, N3131, N2616, N467);
not NOT1 (N3159, N3155);
buf BUF1 (N3160, N3159);
xor XOR2 (N3161, N3157, N2959);
xor XOR2 (N3162, N3154, N1408);
nand NAND3 (N3163, N3161, N2359, N773);
nor NOR4 (N3164, N3160, N128, N1180, N3120);
nand NAND4 (N3165, N3156, N2097, N537, N332);
nand NAND4 (N3166, N3133, N389, N1976, N719);
and AND2 (N3167, N3163, N34);
nand NAND2 (N3168, N3166, N1390);
not NOT1 (N3169, N3158);
buf BUF1 (N3170, N3117);
nor NOR4 (N3171, N3164, N2930, N2090, N2563);
nand NAND3 (N3172, N3167, N458, N2475);
not NOT1 (N3173, N3171);
nor NOR4 (N3174, N3147, N2691, N627, N892);
xor XOR2 (N3175, N3170, N2629);
not NOT1 (N3176, N3175);
nor NOR4 (N3177, N3162, N1182, N3105, N166);
and AND4 (N3178, N3173, N1823, N2429, N2294);
buf BUF1 (N3179, N3177);
xor XOR2 (N3180, N3179, N2325);
nand NAND2 (N3181, N3168, N754);
and AND2 (N3182, N3169, N994);
nand NAND4 (N3183, N3181, N3012, N1761, N262);
nand NAND3 (N3184, N3150, N2056, N1600);
buf BUF1 (N3185, N3178);
not NOT1 (N3186, N3176);
or OR4 (N3187, N3172, N3069, N1970, N2758);
and AND2 (N3188, N3180, N2958);
nor NOR3 (N3189, N3136, N3148, N2338);
xor XOR2 (N3190, N3186, N1208);
nand NAND2 (N3191, N3185, N1540);
xor XOR2 (N3192, N3182, N2795);
not NOT1 (N3193, N3192);
not NOT1 (N3194, N3189);
nand NAND4 (N3195, N3187, N937, N1895, N1804);
buf BUF1 (N3196, N3184);
nand NAND4 (N3197, N3196, N58, N2008, N134);
not NOT1 (N3198, N3195);
nand NAND4 (N3199, N3174, N1914, N1327, N1747);
xor XOR2 (N3200, N3188, N1995);
buf BUF1 (N3201, N3194);
not NOT1 (N3202, N3200);
buf BUF1 (N3203, N3197);
nor NOR3 (N3204, N3190, N1811, N1866);
or OR4 (N3205, N3201, N987, N1303, N393);
nand NAND3 (N3206, N3199, N315, N1033);
not NOT1 (N3207, N3203);
not NOT1 (N3208, N3191);
xor XOR2 (N3209, N3193, N1156);
nand NAND2 (N3210, N3205, N748);
nor NOR4 (N3211, N3202, N2135, N1471, N1589);
nor NOR4 (N3212, N3207, N325, N1027, N2132);
not NOT1 (N3213, N3210);
nor NOR4 (N3214, N3211, N1166, N1437, N995);
and AND3 (N3215, N3183, N1283, N1836);
or OR4 (N3216, N3209, N1362, N2962, N3193);
and AND2 (N3217, N3208, N2529);
nor NOR4 (N3218, N3198, N1564, N2338, N27);
nor NOR3 (N3219, N3215, N2504, N218);
nand NAND3 (N3220, N3219, N1869, N2226);
or OR3 (N3221, N3217, N2076, N741);
nand NAND2 (N3222, N3212, N1864);
nand NAND2 (N3223, N3218, N684);
buf BUF1 (N3224, N3221);
and AND2 (N3225, N3223, N2212);
not NOT1 (N3226, N3204);
nor NOR3 (N3227, N3216, N1962, N1903);
and AND2 (N3228, N3225, N112);
xor XOR2 (N3229, N3213, N2891);
xor XOR2 (N3230, N3206, N258);
or OR4 (N3231, N3224, N261, N2940, N162);
not NOT1 (N3232, N3230);
nor NOR3 (N3233, N3220, N1008, N1012);
or OR2 (N3234, N3227, N1935);
not NOT1 (N3235, N3226);
nand NAND4 (N3236, N3234, N1787, N1847, N3016);
buf BUF1 (N3237, N3236);
xor XOR2 (N3238, N3232, N3029);
not NOT1 (N3239, N3237);
nor NOR2 (N3240, N3229, N1789);
or OR2 (N3241, N3235, N3157);
buf BUF1 (N3242, N3222);
nand NAND2 (N3243, N3240, N1429);
nand NAND3 (N3244, N3231, N3067, N606);
nand NAND2 (N3245, N3242, N2362);
or OR3 (N3246, N3165, N1240, N1168);
not NOT1 (N3247, N3214);
nor NOR3 (N3248, N3238, N397, N559);
and AND4 (N3249, N3244, N627, N576, N3245);
nor NOR3 (N3250, N324, N1724, N3187);
buf BUF1 (N3251, N3247);
xor XOR2 (N3252, N3239, N1701);
nand NAND4 (N3253, N3243, N1382, N2142, N1209);
nor NOR4 (N3254, N3233, N2791, N3136, N1451);
buf BUF1 (N3255, N3252);
nor NOR3 (N3256, N3249, N2619, N2434);
not NOT1 (N3257, N3250);
not NOT1 (N3258, N3248);
and AND2 (N3259, N3241, N1072);
buf BUF1 (N3260, N3246);
buf BUF1 (N3261, N3255);
nand NAND4 (N3262, N3260, N2488, N3224, N1080);
nand NAND3 (N3263, N3262, N258, N802);
not NOT1 (N3264, N3254);
and AND2 (N3265, N3253, N1489);
nor NOR2 (N3266, N3259, N1698);
xor XOR2 (N3267, N3261, N3065);
not NOT1 (N3268, N3257);
and AND2 (N3269, N3267, N1948);
and AND3 (N3270, N3256, N1120, N259);
and AND4 (N3271, N3268, N2432, N63, N2488);
nor NOR4 (N3272, N3270, N279, N2088, N1051);
nor NOR4 (N3273, N3272, N869, N661, N2560);
buf BUF1 (N3274, N3266);
xor XOR2 (N3275, N3273, N2623);
nor NOR2 (N3276, N3251, N360);
or OR4 (N3277, N3271, N1638, N2835, N1035);
xor XOR2 (N3278, N3264, N1122);
buf BUF1 (N3279, N3265);
and AND2 (N3280, N3278, N2477);
and AND4 (N3281, N3228, N2870, N1223, N1683);
nor NOR2 (N3282, N3269, N1000);
nand NAND2 (N3283, N3263, N809);
nor NOR3 (N3284, N3283, N1225, N1946);
xor XOR2 (N3285, N3275, N3250);
buf BUF1 (N3286, N3276);
buf BUF1 (N3287, N3277);
and AND2 (N3288, N3258, N2170);
not NOT1 (N3289, N3282);
and AND3 (N3290, N3287, N1986, N1018);
or OR4 (N3291, N3289, N3056, N1258, N1770);
or OR3 (N3292, N3281, N2453, N1132);
xor XOR2 (N3293, N3288, N779);
nor NOR3 (N3294, N3279, N1947, N3011);
buf BUF1 (N3295, N3290);
nand NAND4 (N3296, N3291, N429, N2077, N3099);
or OR3 (N3297, N3292, N2747, N343);
or OR3 (N3298, N3297, N452, N1935);
or OR2 (N3299, N3298, N271);
nor NOR2 (N3300, N3296, N1623);
and AND2 (N3301, N3274, N302);
not NOT1 (N3302, N3285);
or OR2 (N3303, N3286, N388);
and AND3 (N3304, N3303, N3164, N3237);
and AND2 (N3305, N3299, N2958);
xor XOR2 (N3306, N3305, N2134);
not NOT1 (N3307, N3280);
buf BUF1 (N3308, N3294);
or OR4 (N3309, N3300, N2795, N1610, N3144);
xor XOR2 (N3310, N3293, N860);
nand NAND2 (N3311, N3310, N934);
not NOT1 (N3312, N3308);
not NOT1 (N3313, N3301);
xor XOR2 (N3314, N3304, N2444);
not NOT1 (N3315, N3306);
buf BUF1 (N3316, N3295);
or OR3 (N3317, N3314, N504, N155);
or OR4 (N3318, N3316, N1136, N2534, N1328);
xor XOR2 (N3319, N3315, N2166);
buf BUF1 (N3320, N3319);
and AND4 (N3321, N3309, N530, N1014, N1032);
not NOT1 (N3322, N3312);
not NOT1 (N3323, N3320);
and AND4 (N3324, N3321, N2928, N720, N348);
buf BUF1 (N3325, N3307);
nand NAND4 (N3326, N3317, N447, N1640, N682);
nor NOR3 (N3327, N3325, N1069, N2244);
nor NOR2 (N3328, N3318, N2236);
and AND3 (N3329, N3313, N3104, N2808);
not NOT1 (N3330, N3324);
or OR2 (N3331, N3328, N175);
buf BUF1 (N3332, N3331);
xor XOR2 (N3333, N3330, N2482);
xor XOR2 (N3334, N3284, N886);
xor XOR2 (N3335, N3333, N2148);
xor XOR2 (N3336, N3334, N1102);
not NOT1 (N3337, N3323);
or OR2 (N3338, N3332, N2330);
and AND4 (N3339, N3302, N2676, N533, N318);
nor NOR4 (N3340, N3329, N130, N1293, N325);
buf BUF1 (N3341, N3336);
xor XOR2 (N3342, N3341, N2834);
nand NAND2 (N3343, N3337, N3133);
not NOT1 (N3344, N3322);
or OR4 (N3345, N3335, N2465, N2047, N2120);
buf BUF1 (N3346, N3326);
and AND4 (N3347, N3343, N1574, N2255, N455);
or OR3 (N3348, N3327, N731, N1788);
nand NAND3 (N3349, N3345, N2379, N2550);
nand NAND4 (N3350, N3344, N1873, N1347, N1604);
nand NAND2 (N3351, N3348, N2535);
nor NOR4 (N3352, N3349, N1977, N1618, N1591);
nor NOR2 (N3353, N3347, N1839);
nor NOR4 (N3354, N3346, N1211, N1643, N1080);
buf BUF1 (N3355, N3311);
and AND3 (N3356, N3355, N1978, N1011);
nand NAND3 (N3357, N3351, N1020, N489);
xor XOR2 (N3358, N3340, N1023);
buf BUF1 (N3359, N3358);
nand NAND3 (N3360, N3338, N1855, N3081);
buf BUF1 (N3361, N3357);
buf BUF1 (N3362, N3339);
nor NOR3 (N3363, N3361, N1136, N1117);
nand NAND3 (N3364, N3360, N3223, N1255);
or OR2 (N3365, N3356, N2422);
buf BUF1 (N3366, N3354);
nand NAND2 (N3367, N3362, N2215);
nor NOR2 (N3368, N3359, N661);
buf BUF1 (N3369, N3366);
and AND4 (N3370, N3342, N1246, N1896, N3142);
xor XOR2 (N3371, N3363, N1202);
nand NAND2 (N3372, N3370, N2116);
and AND3 (N3373, N3372, N1993, N1022);
xor XOR2 (N3374, N3368, N2363);
and AND2 (N3375, N3369, N968);
nand NAND4 (N3376, N3373, N2193, N1797, N2405);
and AND2 (N3377, N3350, N3213);
not NOT1 (N3378, N3352);
and AND2 (N3379, N3353, N396);
buf BUF1 (N3380, N3364);
or OR2 (N3381, N3376, N1285);
buf BUF1 (N3382, N3375);
buf BUF1 (N3383, N3365);
or OR4 (N3384, N3381, N2548, N2207, N1633);
buf BUF1 (N3385, N3384);
not NOT1 (N3386, N3379);
buf BUF1 (N3387, N3377);
nor NOR2 (N3388, N3382, N2917);
buf BUF1 (N3389, N3385);
or OR3 (N3390, N3371, N225, N2133);
and AND2 (N3391, N3387, N2300);
xor XOR2 (N3392, N3389, N846);
xor XOR2 (N3393, N3383, N1757);
nor NOR3 (N3394, N3388, N2672, N2608);
xor XOR2 (N3395, N3390, N504);
nor NOR4 (N3396, N3394, N15, N330, N2866);
not NOT1 (N3397, N3396);
and AND4 (N3398, N3395, N1519, N2418, N2213);
nand NAND2 (N3399, N3392, N1153);
nand NAND2 (N3400, N3391, N536);
buf BUF1 (N3401, N3374);
nand NAND3 (N3402, N3367, N2327, N967);
buf BUF1 (N3403, N3380);
and AND2 (N3404, N3401, N2252);
and AND3 (N3405, N3402, N974, N402);
nor NOR2 (N3406, N3378, N3326);
xor XOR2 (N3407, N3386, N1774);
nand NAND2 (N3408, N3393, N2460);
or OR3 (N3409, N3403, N1776, N892);
nor NOR2 (N3410, N3406, N2595);
buf BUF1 (N3411, N3400);
and AND2 (N3412, N3411, N880);
and AND2 (N3413, N3410, N2703);
and AND4 (N3414, N3408, N3225, N2807, N905);
or OR4 (N3415, N3413, N1006, N253, N612);
nor NOR2 (N3416, N3407, N2730);
nand NAND4 (N3417, N3405, N2179, N2728, N534);
xor XOR2 (N3418, N3399, N1817);
xor XOR2 (N3419, N3414, N262);
nand NAND3 (N3420, N3417, N2978, N1180);
nand NAND2 (N3421, N3412, N2063);
xor XOR2 (N3422, N3419, N1744);
or OR2 (N3423, N3416, N929);
xor XOR2 (N3424, N3423, N2081);
xor XOR2 (N3425, N3415, N1837);
xor XOR2 (N3426, N3420, N2937);
buf BUF1 (N3427, N3418);
and AND2 (N3428, N3422, N2150);
and AND2 (N3429, N3428, N2942);
not NOT1 (N3430, N3398);
not NOT1 (N3431, N3424);
or OR3 (N3432, N3427, N579, N2435);
and AND2 (N3433, N3404, N1836);
nand NAND2 (N3434, N3431, N2541);
not NOT1 (N3435, N3426);
or OR3 (N3436, N3432, N41, N2287);
not NOT1 (N3437, N3425);
or OR3 (N3438, N3429, N299, N1369);
xor XOR2 (N3439, N3433, N966);
buf BUF1 (N3440, N3437);
and AND4 (N3441, N3440, N1874, N635, N1955);
and AND3 (N3442, N3434, N446, N3196);
buf BUF1 (N3443, N3438);
nand NAND3 (N3444, N3409, N220, N1342);
nand NAND4 (N3445, N3435, N2681, N3078, N2762);
buf BUF1 (N3446, N3397);
nor NOR4 (N3447, N3444, N3290, N1424, N1665);
nor NOR4 (N3448, N3445, N1233, N2361, N1954);
nand NAND3 (N3449, N3446, N1289, N2246);
nor NOR4 (N3450, N3441, N2855, N2930, N603);
not NOT1 (N3451, N3436);
and AND4 (N3452, N3448, N3339, N866, N2039);
or OR3 (N3453, N3442, N1342, N1871);
buf BUF1 (N3454, N3443);
or OR3 (N3455, N3449, N3264, N1661);
and AND3 (N3456, N3447, N2952, N2126);
nand NAND4 (N3457, N3450, N55, N159, N1155);
nor NOR3 (N3458, N3453, N2526, N1588);
nand NAND2 (N3459, N3455, N3291);
or OR4 (N3460, N3454, N2192, N2566, N435);
not NOT1 (N3461, N3451);
and AND3 (N3462, N3430, N2301, N2311);
not NOT1 (N3463, N3461);
nor NOR4 (N3464, N3421, N1414, N1678, N2316);
not NOT1 (N3465, N3457);
nand NAND3 (N3466, N3452, N2410, N1879);
not NOT1 (N3467, N3464);
and AND3 (N3468, N3465, N855, N82);
or OR2 (N3469, N3468, N1214);
not NOT1 (N3470, N3463);
not NOT1 (N3471, N3459);
buf BUF1 (N3472, N3462);
nand NAND4 (N3473, N3469, N97, N2241, N1129);
nand NAND3 (N3474, N3458, N671, N135);
not NOT1 (N3475, N3456);
nand NAND4 (N3476, N3439, N3161, N1150, N1345);
buf BUF1 (N3477, N3474);
not NOT1 (N3478, N3466);
not NOT1 (N3479, N3460);
nor NOR3 (N3480, N3479, N328, N608);
nor NOR4 (N3481, N3467, N934, N1987, N1797);
or OR2 (N3482, N3472, N715);
and AND4 (N3483, N3480, N3054, N1390, N570);
nand NAND3 (N3484, N3475, N1414, N724);
and AND2 (N3485, N3470, N20);
buf BUF1 (N3486, N3471);
or OR4 (N3487, N3484, N3354, N279, N31);
nand NAND4 (N3488, N3487, N272, N1908, N2317);
xor XOR2 (N3489, N3473, N972);
and AND4 (N3490, N3489, N2437, N1477, N835);
not NOT1 (N3491, N3478);
xor XOR2 (N3492, N3483, N3176);
not NOT1 (N3493, N3488);
or OR4 (N3494, N3492, N3012, N3373, N413);
nand NAND3 (N3495, N3493, N1814, N2102);
nor NOR3 (N3496, N3490, N1378, N2113);
and AND2 (N3497, N3485, N2357);
xor XOR2 (N3498, N3497, N2635);
nor NOR3 (N3499, N3481, N1041, N3083);
not NOT1 (N3500, N3494);
nand NAND2 (N3501, N3500, N1995);
xor XOR2 (N3502, N3498, N3160);
nand NAND4 (N3503, N3502, N2438, N2636, N1152);
not NOT1 (N3504, N3482);
nor NOR3 (N3505, N3499, N374, N1513);
nor NOR3 (N3506, N3476, N1441, N3305);
and AND3 (N3507, N3477, N2800, N2253);
xor XOR2 (N3508, N3504, N1955);
and AND4 (N3509, N3495, N2055, N3117, N2867);
and AND4 (N3510, N3503, N867, N2340, N1940);
buf BUF1 (N3511, N3501);
nor NOR4 (N3512, N3496, N1521, N2109, N1276);
buf BUF1 (N3513, N3491);
buf BUF1 (N3514, N3505);
buf BUF1 (N3515, N3512);
xor XOR2 (N3516, N3511, N2765);
or OR2 (N3517, N3509, N2870);
buf BUF1 (N3518, N3514);
nor NOR3 (N3519, N3518, N1188, N722);
not NOT1 (N3520, N3508);
nor NOR3 (N3521, N3519, N3382, N3030);
nor NOR3 (N3522, N3486, N2317, N2770);
and AND3 (N3523, N3522, N758, N2632);
xor XOR2 (N3524, N3506, N1240);
not NOT1 (N3525, N3523);
nand NAND2 (N3526, N3516, N1992);
xor XOR2 (N3527, N3513, N3263);
nor NOR2 (N3528, N3521, N2690);
nand NAND3 (N3529, N3526, N2409, N2340);
xor XOR2 (N3530, N3525, N2105);
not NOT1 (N3531, N3515);
buf BUF1 (N3532, N3530);
buf BUF1 (N3533, N3527);
or OR4 (N3534, N3531, N356, N1478, N1860);
buf BUF1 (N3535, N3533);
nand NAND4 (N3536, N3529, N3088, N1450, N3079);
buf BUF1 (N3537, N3507);
not NOT1 (N3538, N3535);
nand NAND2 (N3539, N3532, N754);
and AND2 (N3540, N3539, N2126);
nor NOR3 (N3541, N3528, N1981, N1707);
not NOT1 (N3542, N3541);
nor NOR3 (N3543, N3537, N2868, N715);
not NOT1 (N3544, N3510);
or OR3 (N3545, N3536, N3335, N2173);
xor XOR2 (N3546, N3520, N1797);
nand NAND4 (N3547, N3540, N2717, N1201, N3263);
or OR4 (N3548, N3524, N55, N8, N1507);
not NOT1 (N3549, N3538);
buf BUF1 (N3550, N3548);
buf BUF1 (N3551, N3549);
and AND4 (N3552, N3544, N3111, N833, N1200);
or OR4 (N3553, N3543, N2578, N1951, N48);
nor NOR3 (N3554, N3551, N1764, N1061);
buf BUF1 (N3555, N3545);
nand NAND3 (N3556, N3553, N3261, N463);
and AND3 (N3557, N3550, N1887, N2976);
xor XOR2 (N3558, N3557, N3138);
not NOT1 (N3559, N3542);
xor XOR2 (N3560, N3555, N1542);
not NOT1 (N3561, N3554);
xor XOR2 (N3562, N3534, N2764);
or OR3 (N3563, N3558, N903, N1573);
buf BUF1 (N3564, N3552);
buf BUF1 (N3565, N3546);
buf BUF1 (N3566, N3559);
not NOT1 (N3567, N3517);
and AND2 (N3568, N3556, N241);
and AND3 (N3569, N3566, N2630, N1586);
nor NOR4 (N3570, N3560, N3508, N1054, N1928);
nor NOR3 (N3571, N3563, N3300, N3506);
xor XOR2 (N3572, N3561, N2128);
nor NOR4 (N3573, N3567, N3018, N1921, N27);
xor XOR2 (N3574, N3564, N1798);
xor XOR2 (N3575, N3547, N2692);
or OR3 (N3576, N3573, N120, N3471);
and AND2 (N3577, N3565, N2157);
nand NAND4 (N3578, N3571, N337, N1421, N136);
buf BUF1 (N3579, N3575);
nor NOR2 (N3580, N3577, N2426);
or OR3 (N3581, N3570, N3161, N1677);
nor NOR4 (N3582, N3576, N1598, N600, N3119);
nand NAND2 (N3583, N3579, N2921);
and AND2 (N3584, N3578, N1351);
not NOT1 (N3585, N3581);
or OR3 (N3586, N3580, N204, N115);
nand NAND2 (N3587, N3574, N2160);
xor XOR2 (N3588, N3572, N1179);
xor XOR2 (N3589, N3582, N370);
xor XOR2 (N3590, N3588, N2087);
not NOT1 (N3591, N3587);
buf BUF1 (N3592, N3585);
not NOT1 (N3593, N3562);
xor XOR2 (N3594, N3584, N1590);
and AND2 (N3595, N3590, N185);
xor XOR2 (N3596, N3593, N2778);
or OR4 (N3597, N3596, N2106, N3233, N1939);
not NOT1 (N3598, N3583);
and AND4 (N3599, N3598, N3537, N1208, N506);
and AND3 (N3600, N3569, N1326, N2372);
not NOT1 (N3601, N3597);
and AND2 (N3602, N3592, N545);
not NOT1 (N3603, N3595);
buf BUF1 (N3604, N3589);
or OR2 (N3605, N3601, N94);
not NOT1 (N3606, N3591);
buf BUF1 (N3607, N3603);
and AND4 (N3608, N3600, N2574, N2050, N1412);
xor XOR2 (N3609, N3586, N1865);
nand NAND4 (N3610, N3602, N2920, N447, N2671);
buf BUF1 (N3611, N3607);
and AND2 (N3612, N3599, N1612);
xor XOR2 (N3613, N3606, N671);
not NOT1 (N3614, N3594);
nor NOR3 (N3615, N3613, N2337, N3346);
nand NAND4 (N3616, N3608, N2118, N958, N1710);
and AND4 (N3617, N3616, N491, N2985, N1248);
not NOT1 (N3618, N3605);
buf BUF1 (N3619, N3568);
buf BUF1 (N3620, N3619);
nor NOR2 (N3621, N3614, N3519);
and AND3 (N3622, N3604, N3585, N1767);
nor NOR3 (N3623, N3620, N2441, N1455);
nand NAND4 (N3624, N3617, N2016, N243, N2064);
nand NAND4 (N3625, N3622, N1321, N701, N3492);
not NOT1 (N3626, N3623);
and AND3 (N3627, N3621, N702, N1847);
and AND4 (N3628, N3615, N1004, N2528, N466);
xor XOR2 (N3629, N3627, N1987);
buf BUF1 (N3630, N3626);
buf BUF1 (N3631, N3611);
xor XOR2 (N3632, N3631, N2066);
not NOT1 (N3633, N3625);
and AND4 (N3634, N3628, N2276, N3193, N2952);
xor XOR2 (N3635, N3630, N2041);
xor XOR2 (N3636, N3609, N3577);
or OR2 (N3637, N3629, N1917);
not NOT1 (N3638, N3635);
nor NOR4 (N3639, N3624, N923, N1610, N2118);
buf BUF1 (N3640, N3633);
buf BUF1 (N3641, N3632);
not NOT1 (N3642, N3637);
nor NOR2 (N3643, N3638, N2312);
buf BUF1 (N3644, N3642);
nor NOR4 (N3645, N3636, N2629, N640, N2732);
nand NAND2 (N3646, N3618, N3316);
nor NOR4 (N3647, N3643, N2712, N938, N1633);
nand NAND4 (N3648, N3645, N1845, N1878, N1185);
xor XOR2 (N3649, N3641, N1358);
and AND2 (N3650, N3612, N712);
nor NOR4 (N3651, N3634, N2915, N843, N2494);
nor NOR3 (N3652, N3647, N1047, N769);
and AND2 (N3653, N3639, N2796);
not NOT1 (N3654, N3652);
buf BUF1 (N3655, N3640);
not NOT1 (N3656, N3644);
xor XOR2 (N3657, N3646, N2350);
nand NAND2 (N3658, N3649, N3612);
and AND4 (N3659, N3657, N1437, N2394, N2959);
and AND4 (N3660, N3654, N3645, N115, N2555);
nor NOR3 (N3661, N3659, N811, N3154);
not NOT1 (N3662, N3610);
not NOT1 (N3663, N3660);
xor XOR2 (N3664, N3648, N1940);
xor XOR2 (N3665, N3663, N3636);
xor XOR2 (N3666, N3662, N1157);
buf BUF1 (N3667, N3664);
and AND3 (N3668, N3665, N2550, N1646);
nand NAND3 (N3669, N3661, N735, N2902);
and AND3 (N3670, N3668, N3429, N3547);
buf BUF1 (N3671, N3666);
xor XOR2 (N3672, N3658, N957);
not NOT1 (N3673, N3671);
xor XOR2 (N3674, N3653, N2845);
nand NAND2 (N3675, N3667, N2874);
xor XOR2 (N3676, N3650, N2703);
or OR4 (N3677, N3673, N3166, N2430, N2096);
nand NAND3 (N3678, N3656, N1632, N3212);
or OR4 (N3679, N3672, N897, N1258, N2692);
buf BUF1 (N3680, N3669);
xor XOR2 (N3681, N3674, N611);
not NOT1 (N3682, N3677);
nor NOR3 (N3683, N3679, N2509, N550);
or OR3 (N3684, N3651, N225, N1999);
nor NOR3 (N3685, N3680, N2675, N654);
buf BUF1 (N3686, N3678);
xor XOR2 (N3687, N3684, N117);
and AND2 (N3688, N3686, N2093);
xor XOR2 (N3689, N3687, N1962);
nor NOR4 (N3690, N3688, N1461, N1154, N1550);
nor NOR2 (N3691, N3683, N3462);
and AND2 (N3692, N3676, N1912);
or OR2 (N3693, N3692, N3507);
nor NOR4 (N3694, N3693, N3332, N3228, N3122);
buf BUF1 (N3695, N3685);
buf BUF1 (N3696, N3681);
or OR2 (N3697, N3696, N825);
not NOT1 (N3698, N3670);
not NOT1 (N3699, N3694);
xor XOR2 (N3700, N3690, N164);
nor NOR3 (N3701, N3675, N1043, N2809);
nand NAND3 (N3702, N3695, N137, N906);
or OR3 (N3703, N3698, N417, N2436);
and AND3 (N3704, N3655, N2567, N774);
and AND2 (N3705, N3691, N1494);
nand NAND2 (N3706, N3704, N2507);
not NOT1 (N3707, N3702);
xor XOR2 (N3708, N3701, N1434);
not NOT1 (N3709, N3700);
buf BUF1 (N3710, N3706);
nand NAND4 (N3711, N3703, N2978, N1177, N2571);
nand NAND4 (N3712, N3689, N3591, N3080, N1850);
nor NOR2 (N3713, N3712, N113);
and AND2 (N3714, N3697, N1406);
and AND3 (N3715, N3711, N2316, N534);
xor XOR2 (N3716, N3710, N900);
or OR4 (N3717, N3714, N2851, N618, N3458);
or OR2 (N3718, N3717, N1177);
buf BUF1 (N3719, N3709);
nor NOR4 (N3720, N3719, N2215, N3574, N707);
nor NOR4 (N3721, N3707, N2447, N1892, N3422);
buf BUF1 (N3722, N3716);
nor NOR4 (N3723, N3721, N2158, N2693, N2676);
nand NAND3 (N3724, N3718, N699, N2902);
nor NOR3 (N3725, N3715, N1860, N3572);
nand NAND2 (N3726, N3708, N51);
and AND2 (N3727, N3726, N3187);
xor XOR2 (N3728, N3682, N3672);
nand NAND3 (N3729, N3724, N3684, N1220);
buf BUF1 (N3730, N3728);
not NOT1 (N3731, N3699);
and AND4 (N3732, N3720, N2618, N1513, N1894);
and AND3 (N3733, N3729, N2294, N2847);
not NOT1 (N3734, N3727);
xor XOR2 (N3735, N3731, N480);
nor NOR4 (N3736, N3723, N3269, N614, N3217);
buf BUF1 (N3737, N3705);
nor NOR2 (N3738, N3735, N175);
nand NAND4 (N3739, N3725, N1581, N3466, N2444);
and AND4 (N3740, N3732, N1670, N1319, N129);
nand NAND4 (N3741, N3734, N1782, N677, N536);
or OR3 (N3742, N3741, N565, N2042);
or OR2 (N3743, N3740, N363);
and AND3 (N3744, N3730, N3511, N3638);
buf BUF1 (N3745, N3742);
nand NAND3 (N3746, N3738, N1057, N35);
nand NAND3 (N3747, N3736, N3450, N1051);
xor XOR2 (N3748, N3733, N1890);
not NOT1 (N3749, N3744);
nand NAND4 (N3750, N3722, N2215, N3305, N1774);
or OR3 (N3751, N3747, N1817, N2476);
or OR2 (N3752, N3746, N1676);
nand NAND3 (N3753, N3737, N2590, N836);
xor XOR2 (N3754, N3750, N486);
or OR3 (N3755, N3754, N161, N2879);
and AND2 (N3756, N3713, N999);
xor XOR2 (N3757, N3739, N456);
nor NOR4 (N3758, N3752, N3345, N2, N3716);
or OR4 (N3759, N3756, N1375, N2202, N1593);
xor XOR2 (N3760, N3758, N3283);
not NOT1 (N3761, N3759);
and AND3 (N3762, N3753, N1892, N3073);
or OR3 (N3763, N3755, N1234, N1488);
not NOT1 (N3764, N3757);
or OR2 (N3765, N3743, N176);
nor NOR3 (N3766, N3764, N624, N1455);
not NOT1 (N3767, N3748);
and AND2 (N3768, N3745, N383);
nand NAND2 (N3769, N3749, N2077);
not NOT1 (N3770, N3760);
not NOT1 (N3771, N3766);
not NOT1 (N3772, N3769);
xor XOR2 (N3773, N3772, N1610);
xor XOR2 (N3774, N3771, N2143);
nand NAND4 (N3775, N3774, N2885, N830, N2175);
nor NOR2 (N3776, N3762, N2765);
and AND3 (N3777, N3773, N2252, N681);
xor XOR2 (N3778, N3761, N507);
nand NAND2 (N3779, N3767, N115);
not NOT1 (N3780, N3768);
or OR3 (N3781, N3770, N1975, N662);
xor XOR2 (N3782, N3765, N2593);
nor NOR2 (N3783, N3779, N2315);
and AND4 (N3784, N3783, N802, N2300, N3203);
nand NAND2 (N3785, N3781, N2577);
buf BUF1 (N3786, N3782);
not NOT1 (N3787, N3784);
xor XOR2 (N3788, N3786, N2543);
or OR4 (N3789, N3787, N2911, N1861, N598);
not NOT1 (N3790, N3775);
or OR4 (N3791, N3776, N1008, N337, N106);
and AND3 (N3792, N3791, N1212, N1712);
nor NOR3 (N3793, N3778, N963, N1851);
nor NOR2 (N3794, N3777, N1630);
not NOT1 (N3795, N3788);
nand NAND3 (N3796, N3793, N2563, N3606);
nand NAND4 (N3797, N3789, N788, N3162, N612);
and AND2 (N3798, N3794, N449);
and AND2 (N3799, N3751, N437);
nor NOR3 (N3800, N3792, N607, N336);
or OR2 (N3801, N3763, N5);
xor XOR2 (N3802, N3797, N3218);
nor NOR4 (N3803, N3780, N2245, N2497, N1931);
nor NOR3 (N3804, N3802, N2672, N75);
or OR4 (N3805, N3804, N1632, N92, N1679);
xor XOR2 (N3806, N3796, N804);
nand NAND4 (N3807, N3806, N1784, N2304, N2681);
buf BUF1 (N3808, N3795);
buf BUF1 (N3809, N3790);
xor XOR2 (N3810, N3798, N1781);
or OR4 (N3811, N3810, N2233, N1957, N100);
nand NAND4 (N3812, N3809, N1202, N777, N1375);
not NOT1 (N3813, N3812);
or OR2 (N3814, N3785, N2128);
and AND2 (N3815, N3801, N1927);
xor XOR2 (N3816, N3815, N275);
nand NAND2 (N3817, N3807, N1145);
not NOT1 (N3818, N3814);
and AND4 (N3819, N3805, N712, N2835, N2433);
nand NAND3 (N3820, N3813, N3110, N2954);
nand NAND2 (N3821, N3819, N1774);
xor XOR2 (N3822, N3799, N195);
nand NAND3 (N3823, N3818, N1817, N2833);
xor XOR2 (N3824, N3822, N471);
and AND3 (N3825, N3803, N785, N3554);
nor NOR3 (N3826, N3811, N1172, N2387);
not NOT1 (N3827, N3817);
nor NOR2 (N3828, N3821, N342);
nor NOR3 (N3829, N3828, N2218, N3461);
nand NAND3 (N3830, N3823, N1602, N526);
xor XOR2 (N3831, N3808, N414);
and AND3 (N3832, N3800, N2531, N1601);
nand NAND3 (N3833, N3816, N2886, N3164);
xor XOR2 (N3834, N3820, N673);
and AND4 (N3835, N3833, N2597, N2842, N1034);
buf BUF1 (N3836, N3829);
or OR4 (N3837, N3824, N1825, N1307, N2686);
buf BUF1 (N3838, N3835);
nand NAND4 (N3839, N3827, N2934, N721, N89);
or OR2 (N3840, N3834, N510);
or OR2 (N3841, N3831, N2668);
xor XOR2 (N3842, N3838, N2311);
nor NOR4 (N3843, N3830, N511, N3116, N3367);
buf BUF1 (N3844, N3840);
nor NOR3 (N3845, N3837, N2604, N2262);
buf BUF1 (N3846, N3825);
or OR2 (N3847, N3844, N3365);
and AND3 (N3848, N3847, N53, N2143);
xor XOR2 (N3849, N3842, N2478);
and AND4 (N3850, N3845, N1066, N2784, N1078);
nand NAND2 (N3851, N3846, N3708);
or OR2 (N3852, N3850, N3243);
nor NOR3 (N3853, N3843, N1997, N3517);
nor NOR2 (N3854, N3832, N2278);
nor NOR3 (N3855, N3851, N2360, N2606);
not NOT1 (N3856, N3855);
not NOT1 (N3857, N3856);
or OR3 (N3858, N3836, N2720, N1484);
or OR2 (N3859, N3852, N3649);
buf BUF1 (N3860, N3857);
or OR4 (N3861, N3853, N3377, N387, N229);
nand NAND4 (N3862, N3849, N3096, N3045, N286);
or OR3 (N3863, N3841, N3628, N1109);
xor XOR2 (N3864, N3862, N803);
buf BUF1 (N3865, N3861);
nand NAND3 (N3866, N3858, N1833, N1314);
nand NAND4 (N3867, N3866, N1199, N2863, N1764);
and AND4 (N3868, N3826, N397, N3795, N3052);
nand NAND4 (N3869, N3860, N1609, N2781, N1978);
and AND3 (N3870, N3854, N1969, N2840);
or OR4 (N3871, N3864, N3082, N2381, N640);
or OR4 (N3872, N3870, N1990, N3849, N2275);
or OR3 (N3873, N3872, N524, N243);
or OR2 (N3874, N3867, N2033);
buf BUF1 (N3875, N3868);
nor NOR2 (N3876, N3848, N1850);
xor XOR2 (N3877, N3865, N2733);
nor NOR3 (N3878, N3874, N1113, N847);
or OR3 (N3879, N3839, N127, N1906);
nand NAND3 (N3880, N3859, N3237, N1168);
nor NOR2 (N3881, N3880, N2056);
buf BUF1 (N3882, N3881);
not NOT1 (N3883, N3882);
or OR2 (N3884, N3873, N1433);
or OR3 (N3885, N3877, N1845, N503);
not NOT1 (N3886, N3885);
not NOT1 (N3887, N3886);
buf BUF1 (N3888, N3878);
nor NOR2 (N3889, N3879, N687);
not NOT1 (N3890, N3875);
and AND3 (N3891, N3869, N1638, N2831);
xor XOR2 (N3892, N3884, N1578);
xor XOR2 (N3893, N3891, N3254);
nor NOR3 (N3894, N3887, N1355, N3012);
nand NAND2 (N3895, N3893, N3021);
xor XOR2 (N3896, N3895, N2988);
or OR3 (N3897, N3883, N731, N367);
nor NOR3 (N3898, N3896, N1189, N3636);
and AND2 (N3899, N3892, N944);
xor XOR2 (N3900, N3888, N1849);
not NOT1 (N3901, N3889);
buf BUF1 (N3902, N3863);
nor NOR3 (N3903, N3900, N205, N836);
nor NOR3 (N3904, N3901, N556, N268);
nand NAND2 (N3905, N3890, N2071);
or OR2 (N3906, N3898, N1739);
and AND4 (N3907, N3876, N3793, N3373, N1412);
or OR4 (N3908, N3871, N545, N1331, N283);
xor XOR2 (N3909, N3907, N2069);
nor NOR2 (N3910, N3905, N3786);
buf BUF1 (N3911, N3903);
nor NOR3 (N3912, N3909, N576, N2397);
nor NOR3 (N3913, N3906, N2021, N3378);
and AND3 (N3914, N3913, N1593, N927);
or OR2 (N3915, N3902, N2224);
xor XOR2 (N3916, N3915, N2728);
xor XOR2 (N3917, N3897, N2686);
or OR3 (N3918, N3910, N2503, N1980);
nand NAND3 (N3919, N3904, N2435, N2995);
and AND2 (N3920, N3912, N1387);
nand NAND4 (N3921, N3894, N3919, N3568, N1653);
nor NOR2 (N3922, N2888, N3245);
nand NAND2 (N3923, N3916, N1856);
or OR4 (N3924, N3918, N2983, N3436, N2606);
buf BUF1 (N3925, N3922);
and AND3 (N3926, N3923, N2444, N2331);
or OR4 (N3927, N3899, N2664, N1040, N3446);
nor NOR4 (N3928, N3920, N3260, N3593, N1531);
nor NOR2 (N3929, N3908, N2251);
not NOT1 (N3930, N3914);
or OR2 (N3931, N3917, N1160);
xor XOR2 (N3932, N3928, N1726);
xor XOR2 (N3933, N3930, N1236);
xor XOR2 (N3934, N3927, N3535);
nor NOR4 (N3935, N3926, N3741, N154, N2916);
xor XOR2 (N3936, N3934, N1868);
and AND3 (N3937, N3931, N2330, N1354);
buf BUF1 (N3938, N3911);
and AND4 (N3939, N3932, N3484, N2195, N3532);
nand NAND4 (N3940, N3936, N2553, N356, N1050);
buf BUF1 (N3941, N3924);
nor NOR4 (N3942, N3921, N3512, N3834, N704);
nor NOR3 (N3943, N3942, N1076, N3312);
and AND4 (N3944, N3925, N2301, N722, N227);
buf BUF1 (N3945, N3933);
buf BUF1 (N3946, N3943);
buf BUF1 (N3947, N3944);
and AND4 (N3948, N3935, N2029, N2982, N3743);
and AND3 (N3949, N3937, N2219, N674);
nand NAND2 (N3950, N3929, N817);
or OR2 (N3951, N3949, N3015);
and AND3 (N3952, N3939, N3231, N1646);
not NOT1 (N3953, N3945);
nor NOR2 (N3954, N3952, N708);
xor XOR2 (N3955, N3947, N661);
and AND3 (N3956, N3938, N1642, N936);
or OR3 (N3957, N3951, N1856, N1908);
nand NAND2 (N3958, N3956, N3442);
and AND2 (N3959, N3948, N656);
xor XOR2 (N3960, N3950, N2854);
not NOT1 (N3961, N3946);
not NOT1 (N3962, N3960);
not NOT1 (N3963, N3955);
buf BUF1 (N3964, N3958);
buf BUF1 (N3965, N3941);
nand NAND2 (N3966, N3965, N684);
nor NOR3 (N3967, N3954, N2787, N1949);
nand NAND4 (N3968, N3964, N1109, N1546, N1720);
and AND2 (N3969, N3959, N1865);
nor NOR2 (N3970, N3968, N3803);
nor NOR4 (N3971, N3969, N2280, N2025, N1574);
and AND4 (N3972, N3940, N1281, N2495, N1520);
not NOT1 (N3973, N3967);
xor XOR2 (N3974, N3961, N1815);
nand NAND2 (N3975, N3972, N1106);
nand NAND2 (N3976, N3973, N1514);
and AND4 (N3977, N3976, N3304, N824, N3630);
and AND3 (N3978, N3953, N3241, N3595);
xor XOR2 (N3979, N3977, N3702);
or OR2 (N3980, N3979, N3358);
or OR2 (N3981, N3978, N948);
buf BUF1 (N3982, N3970);
not NOT1 (N3983, N3962);
buf BUF1 (N3984, N3980);
xor XOR2 (N3985, N3957, N2107);
not NOT1 (N3986, N3963);
or OR3 (N3987, N3985, N2616, N50);
nand NAND3 (N3988, N3975, N3784, N3724);
and AND4 (N3989, N3981, N1940, N2199, N647);
buf BUF1 (N3990, N3983);
or OR4 (N3991, N3966, N3088, N3885, N2254);
nor NOR3 (N3992, N3984, N128, N374);
nand NAND4 (N3993, N3974, N1048, N2939, N3830);
buf BUF1 (N3994, N3993);
not NOT1 (N3995, N3982);
and AND4 (N3996, N3989, N932, N3015, N593);
nand NAND4 (N3997, N3991, N360, N521, N416);
buf BUF1 (N3998, N3988);
nor NOR2 (N3999, N3971, N1165);
and AND4 (N4000, N3998, N2516, N783, N2848);
xor XOR2 (N4001, N3994, N2189);
or OR2 (N4002, N3996, N1488);
not NOT1 (N4003, N4000);
nand NAND4 (N4004, N4003, N1118, N905, N2580);
xor XOR2 (N4005, N4004, N832);
nor NOR4 (N4006, N3992, N636, N1130, N2352);
or OR3 (N4007, N4002, N3293, N213);
xor XOR2 (N4008, N3995, N1712);
nand NAND3 (N4009, N4006, N534, N1245);
nor NOR4 (N4010, N4001, N2306, N236, N1074);
not NOT1 (N4011, N4010);
not NOT1 (N4012, N4008);
not NOT1 (N4013, N4005);
nor NOR3 (N4014, N3987, N1406, N1871);
not NOT1 (N4015, N4013);
nor NOR4 (N4016, N4012, N7, N3443, N3034);
not NOT1 (N4017, N4011);
not NOT1 (N4018, N4009);
and AND4 (N4019, N3997, N1673, N1473, N3479);
xor XOR2 (N4020, N3999, N280);
nand NAND3 (N4021, N3986, N2594, N840);
buf BUF1 (N4022, N4018);
not NOT1 (N4023, N4021);
nand NAND4 (N4024, N4016, N179, N710, N616);
nand NAND3 (N4025, N4024, N1056, N1513);
not NOT1 (N4026, N4007);
and AND4 (N4027, N3990, N254, N2736, N2826);
or OR3 (N4028, N4022, N2921, N85);
and AND4 (N4029, N4020, N657, N1613, N2129);
buf BUF1 (N4030, N4019);
nand NAND2 (N4031, N4027, N2832);
or OR4 (N4032, N4014, N2501, N94, N726);
or OR2 (N4033, N4026, N3339);
nor NOR4 (N4034, N4015, N2810, N1679, N1363);
nand NAND3 (N4035, N4029, N3571, N3202);
buf BUF1 (N4036, N4017);
or OR3 (N4037, N4023, N3915, N1244);
nand NAND2 (N4038, N4025, N3251);
buf BUF1 (N4039, N4033);
or OR3 (N4040, N4031, N2710, N1914);
not NOT1 (N4041, N4038);
buf BUF1 (N4042, N4041);
xor XOR2 (N4043, N4034, N3783);
nand NAND2 (N4044, N4036, N2290);
buf BUF1 (N4045, N4030);
and AND3 (N4046, N4042, N1276, N2216);
not NOT1 (N4047, N4028);
nor NOR4 (N4048, N4040, N2159, N138, N584);
xor XOR2 (N4049, N4043, N2258);
nor NOR2 (N4050, N4047, N2271);
and AND2 (N4051, N4046, N2027);
buf BUF1 (N4052, N4051);
nand NAND4 (N4053, N4045, N1998, N3414, N3031);
nand NAND3 (N4054, N4048, N1427, N2577);
not NOT1 (N4055, N4032);
or OR3 (N4056, N4044, N3507, N1458);
nor NOR3 (N4057, N4053, N3713, N3550);
and AND3 (N4058, N4054, N2284, N2506);
buf BUF1 (N4059, N4058);
not NOT1 (N4060, N4057);
nor NOR4 (N4061, N4050, N1361, N1169, N3712);
nand NAND3 (N4062, N4039, N1736, N2704);
and AND2 (N4063, N4062, N1216);
buf BUF1 (N4064, N4055);
xor XOR2 (N4065, N4052, N672);
xor XOR2 (N4066, N4063, N3985);
buf BUF1 (N4067, N4060);
xor XOR2 (N4068, N4066, N670);
not NOT1 (N4069, N4037);
and AND3 (N4070, N4067, N4038, N802);
and AND3 (N4071, N4069, N3342, N3493);
xor XOR2 (N4072, N4035, N3398);
and AND2 (N4073, N4070, N3329);
nor NOR3 (N4074, N4064, N1385, N2810);
nor NOR4 (N4075, N4072, N1311, N3950, N3029);
or OR3 (N4076, N4061, N3676, N1749);
buf BUF1 (N4077, N4068);
not NOT1 (N4078, N4073);
and AND3 (N4079, N4076, N362, N2195);
and AND3 (N4080, N4077, N3216, N347);
xor XOR2 (N4081, N4074, N3359);
and AND3 (N4082, N4065, N3778, N861);
nor NOR3 (N4083, N4071, N3161, N1887);
nor NOR4 (N4084, N4080, N335, N1373, N3836);
buf BUF1 (N4085, N4078);
buf BUF1 (N4086, N4083);
or OR2 (N4087, N4082, N3398);
xor XOR2 (N4088, N4049, N3931);
or OR3 (N4089, N4056, N2330, N3909);
and AND4 (N4090, N4088, N3056, N3762, N245);
nand NAND2 (N4091, N4079, N3980);
xor XOR2 (N4092, N4091, N471);
nor NOR3 (N4093, N4090, N781, N3680);
xor XOR2 (N4094, N4086, N2669);
not NOT1 (N4095, N4094);
xor XOR2 (N4096, N4087, N3113);
buf BUF1 (N4097, N4096);
and AND4 (N4098, N4075, N1719, N577, N2340);
and AND2 (N4099, N4097, N1180);
xor XOR2 (N4100, N4085, N2002);
nand NAND4 (N4101, N4089, N739, N3181, N2950);
and AND4 (N4102, N4092, N2806, N3904, N985);
and AND4 (N4103, N4093, N4041, N1895, N3718);
not NOT1 (N4104, N4102);
and AND2 (N4105, N4101, N4051);
not NOT1 (N4106, N4105);
xor XOR2 (N4107, N4098, N1505);
not NOT1 (N4108, N4104);
not NOT1 (N4109, N4107);
and AND4 (N4110, N4095, N367, N63, N97);
nor NOR2 (N4111, N4100, N2511);
nor NOR2 (N4112, N4111, N2616);
and AND4 (N4113, N4108, N47, N1312, N3127);
xor XOR2 (N4114, N4103, N1274);
and AND3 (N4115, N4084, N556, N3975);
nand NAND2 (N4116, N4099, N3505);
or OR3 (N4117, N4110, N1210, N971);
xor XOR2 (N4118, N4114, N3116);
nand NAND4 (N4119, N4116, N1323, N1770, N2000);
or OR2 (N4120, N4059, N1093);
buf BUF1 (N4121, N4109);
or OR3 (N4122, N4119, N3560, N1320);
xor XOR2 (N4123, N4106, N1381);
or OR3 (N4124, N4120, N2884, N3445);
nand NAND4 (N4125, N4124, N1085, N734, N3541);
buf BUF1 (N4126, N4123);
not NOT1 (N4127, N4081);
or OR3 (N4128, N4115, N429, N2647);
buf BUF1 (N4129, N4113);
nor NOR2 (N4130, N4112, N2156);
buf BUF1 (N4131, N4129);
xor XOR2 (N4132, N4126, N409);
nand NAND4 (N4133, N4131, N3266, N3473, N2277);
buf BUF1 (N4134, N4122);
or OR3 (N4135, N4130, N3533, N1227);
nand NAND3 (N4136, N4132, N163, N3699);
nand NAND4 (N4137, N4136, N1252, N2637, N3701);
xor XOR2 (N4138, N4118, N3220);
and AND4 (N4139, N4134, N3930, N1166, N28);
nor NOR3 (N4140, N4128, N2757, N982);
nor NOR4 (N4141, N4133, N2095, N2960, N1487);
nor NOR3 (N4142, N4125, N2557, N3620);
nor NOR4 (N4143, N4140, N458, N147, N4077);
or OR4 (N4144, N4138, N2326, N3553, N1868);
not NOT1 (N4145, N4141);
not NOT1 (N4146, N4135);
xor XOR2 (N4147, N4117, N2388);
buf BUF1 (N4148, N4145);
nand NAND4 (N4149, N4147, N52, N1869, N2420);
and AND4 (N4150, N4143, N1721, N801, N875);
and AND4 (N4151, N4142, N2355, N3563, N1800);
nor NOR2 (N4152, N4150, N430);
and AND2 (N4153, N4137, N702);
not NOT1 (N4154, N4144);
nor NOR2 (N4155, N4146, N1274);
nand NAND4 (N4156, N4152, N1236, N1763, N1182);
nor NOR2 (N4157, N4121, N2513);
not NOT1 (N4158, N4148);
or OR4 (N4159, N4157, N3204, N2561, N3416);
or OR2 (N4160, N4158, N3502);
or OR3 (N4161, N4159, N2956, N13);
xor XOR2 (N4162, N4139, N1459);
not NOT1 (N4163, N4149);
or OR4 (N4164, N4156, N1168, N95, N3084);
or OR3 (N4165, N4151, N3427, N3734);
nor NOR4 (N4166, N4161, N3900, N3644, N51);
nand NAND2 (N4167, N4154, N740);
not NOT1 (N4168, N4162);
not NOT1 (N4169, N4165);
buf BUF1 (N4170, N4163);
buf BUF1 (N4171, N4164);
nand NAND2 (N4172, N4160, N921);
xor XOR2 (N4173, N4166, N417);
or OR4 (N4174, N4167, N322, N1752, N1511);
xor XOR2 (N4175, N4127, N1193);
buf BUF1 (N4176, N4169);
nand NAND2 (N4177, N4153, N2627);
nor NOR4 (N4178, N4176, N1576, N1900, N3987);
xor XOR2 (N4179, N4171, N1461);
and AND3 (N4180, N4168, N1863, N812);
and AND4 (N4181, N4177, N3276, N2986, N1341);
nand NAND3 (N4182, N4181, N345, N2830);
and AND4 (N4183, N4172, N3614, N2784, N3366);
xor XOR2 (N4184, N4155, N816);
not NOT1 (N4185, N4174);
and AND3 (N4186, N4175, N1763, N2811);
xor XOR2 (N4187, N4170, N3044);
nand NAND4 (N4188, N4185, N201, N611, N3160);
nor NOR2 (N4189, N4186, N4111);
xor XOR2 (N4190, N4179, N4076);
xor XOR2 (N4191, N4188, N2080);
buf BUF1 (N4192, N4189);
not NOT1 (N4193, N4187);
or OR2 (N4194, N4182, N1565);
or OR2 (N4195, N4194, N3877);
and AND2 (N4196, N4178, N1503);
xor XOR2 (N4197, N4191, N2246);
and AND2 (N4198, N4195, N2283);
nor NOR2 (N4199, N4192, N1698);
nor NOR3 (N4200, N4193, N520, N976);
buf BUF1 (N4201, N4199);
xor XOR2 (N4202, N4184, N3572);
not NOT1 (N4203, N4202);
and AND3 (N4204, N4183, N140, N3351);
not NOT1 (N4205, N4204);
nand NAND3 (N4206, N4198, N778, N506);
xor XOR2 (N4207, N4196, N554);
nand NAND4 (N4208, N4197, N3718, N3931, N2352);
or OR2 (N4209, N4201, N3409);
and AND3 (N4210, N4207, N4027, N699);
xor XOR2 (N4211, N4210, N3058);
buf BUF1 (N4212, N4173);
not NOT1 (N4213, N4205);
not NOT1 (N4214, N4206);
nor NOR3 (N4215, N4180, N3029, N1715);
nor NOR2 (N4216, N4214, N3802);
nor NOR3 (N4217, N4200, N3278, N869);
not NOT1 (N4218, N4212);
buf BUF1 (N4219, N4190);
and AND2 (N4220, N4218, N2999);
nor NOR3 (N4221, N4203, N239, N3430);
or OR3 (N4222, N4215, N478, N2862);
or OR2 (N4223, N4208, N591);
nand NAND4 (N4224, N4217, N1704, N4125, N1434);
nor NOR3 (N4225, N4222, N3046, N610);
buf BUF1 (N4226, N4213);
and AND4 (N4227, N4225, N357, N2216, N677);
not NOT1 (N4228, N4227);
not NOT1 (N4229, N4216);
xor XOR2 (N4230, N4226, N3555);
xor XOR2 (N4231, N4229, N3414);
nand NAND2 (N4232, N4223, N3281);
and AND4 (N4233, N4231, N424, N1031, N13);
and AND4 (N4234, N4220, N4129, N2952, N1192);
or OR4 (N4235, N4209, N2928, N1298, N702);
buf BUF1 (N4236, N4224);
or OR2 (N4237, N4221, N3513);
buf BUF1 (N4238, N4233);
and AND2 (N4239, N4236, N1174);
not NOT1 (N4240, N4228);
not NOT1 (N4241, N4238);
or OR2 (N4242, N4240, N1498);
not NOT1 (N4243, N4235);
nor NOR2 (N4244, N4234, N2148);
or OR4 (N4245, N4211, N3274, N3611, N1986);
not NOT1 (N4246, N4239);
or OR3 (N4247, N4246, N3020, N1081);
xor XOR2 (N4248, N4247, N3524);
buf BUF1 (N4249, N4242);
nor NOR4 (N4250, N4248, N884, N4102, N1391);
and AND2 (N4251, N4241, N3195);
or OR3 (N4252, N4243, N1557, N2790);
and AND2 (N4253, N4244, N2422);
buf BUF1 (N4254, N4251);
nand NAND3 (N4255, N4253, N1693, N2271);
or OR2 (N4256, N4252, N1633);
or OR4 (N4257, N4237, N249, N3858, N1629);
or OR2 (N4258, N4254, N2732);
buf BUF1 (N4259, N4219);
and AND4 (N4260, N4250, N3606, N4042, N4219);
nor NOR3 (N4261, N4232, N116, N527);
and AND2 (N4262, N4256, N3038);
nand NAND2 (N4263, N4230, N282);
not NOT1 (N4264, N4257);
nand NAND4 (N4265, N4263, N3400, N4261, N1767);
nor NOR3 (N4266, N1508, N2512, N2305);
nand NAND4 (N4267, N4260, N1920, N4243, N1190);
xor XOR2 (N4268, N4259, N1550);
buf BUF1 (N4269, N4266);
buf BUF1 (N4270, N4249);
or OR4 (N4271, N4265, N1240, N2763, N1427);
or OR4 (N4272, N4268, N2514, N1523, N1111);
xor XOR2 (N4273, N4255, N1161);
not NOT1 (N4274, N4245);
or OR2 (N4275, N4274, N3596);
xor XOR2 (N4276, N4267, N2480);
and AND3 (N4277, N4275, N3254, N573);
xor XOR2 (N4278, N4271, N1348);
buf BUF1 (N4279, N4277);
or OR3 (N4280, N4262, N2997, N2755);
nor NOR4 (N4281, N4278, N3750, N1033, N1759);
xor XOR2 (N4282, N4281, N1861);
not NOT1 (N4283, N4258);
nand NAND3 (N4284, N4282, N91, N2364);
or OR2 (N4285, N4272, N1888);
nor NOR4 (N4286, N4276, N884, N20, N650);
nand NAND4 (N4287, N4285, N3501, N3806, N3172);
nor NOR3 (N4288, N4264, N677, N495);
nand NAND3 (N4289, N4279, N2682, N2133);
nor NOR3 (N4290, N4288, N3109, N2011);
nor NOR4 (N4291, N4269, N740, N2632, N3633);
and AND2 (N4292, N4273, N3696);
buf BUF1 (N4293, N4270);
or OR4 (N4294, N4291, N3412, N741, N3511);
xor XOR2 (N4295, N4293, N2594);
xor XOR2 (N4296, N4283, N183);
xor XOR2 (N4297, N4280, N792);
xor XOR2 (N4298, N4290, N2970);
nand NAND3 (N4299, N4296, N3247, N2873);
nor NOR4 (N4300, N4284, N1406, N1521, N184);
nor NOR3 (N4301, N4286, N2693, N1839);
nor NOR3 (N4302, N4299, N1213, N1606);
or OR4 (N4303, N4292, N3799, N3576, N1204);
or OR4 (N4304, N4300, N1074, N919, N980);
buf BUF1 (N4305, N4297);
buf BUF1 (N4306, N4287);
or OR2 (N4307, N4303, N915);
or OR4 (N4308, N4289, N3866, N3766, N2721);
buf BUF1 (N4309, N4306);
or OR4 (N4310, N4294, N3621, N2820, N3743);
nand NAND2 (N4311, N4308, N3077);
nand NAND2 (N4312, N4310, N3272);
xor XOR2 (N4313, N4305, N4279);
xor XOR2 (N4314, N4301, N3832);
xor XOR2 (N4315, N4313, N1384);
and AND3 (N4316, N4302, N791, N1020);
xor XOR2 (N4317, N4307, N3782);
xor XOR2 (N4318, N4315, N2262);
xor XOR2 (N4319, N4317, N1319);
and AND3 (N4320, N4304, N3863, N2459);
xor XOR2 (N4321, N4298, N2181);
or OR4 (N4322, N4316, N1553, N2274, N990);
nor NOR4 (N4323, N4321, N1894, N3647, N1764);
xor XOR2 (N4324, N4312, N1818);
buf BUF1 (N4325, N4323);
xor XOR2 (N4326, N4309, N3224);
nand NAND2 (N4327, N4324, N2275);
or OR2 (N4328, N4318, N3410);
and AND4 (N4329, N4314, N2153, N3162, N2678);
nand NAND2 (N4330, N4319, N349);
or OR2 (N4331, N4326, N4209);
nand NAND4 (N4332, N4322, N548, N1955, N2116);
nand NAND2 (N4333, N4330, N2374);
nand NAND2 (N4334, N4329, N3043);
not NOT1 (N4335, N4334);
not NOT1 (N4336, N4320);
buf BUF1 (N4337, N4333);
buf BUF1 (N4338, N4327);
nor NOR3 (N4339, N4311, N1181, N610);
nor NOR4 (N4340, N4335, N2205, N472, N2183);
nor NOR2 (N4341, N4332, N2565);
buf BUF1 (N4342, N4337);
or OR4 (N4343, N4295, N298, N1561, N4081);
not NOT1 (N4344, N4325);
nand NAND4 (N4345, N4343, N245, N4104, N1752);
nand NAND4 (N4346, N4345, N3816, N3290, N3927);
xor XOR2 (N4347, N4344, N1771);
or OR4 (N4348, N4328, N3294, N3387, N2479);
xor XOR2 (N4349, N4342, N3823);
xor XOR2 (N4350, N4339, N3747);
and AND2 (N4351, N4341, N2223);
nand NAND3 (N4352, N4336, N3667, N1272);
not NOT1 (N4353, N4350);
nor NOR4 (N4354, N4340, N1136, N3630, N2865);
or OR3 (N4355, N4346, N3315, N603);
xor XOR2 (N4356, N4338, N1375);
nor NOR4 (N4357, N4356, N54, N2291, N360);
nor NOR3 (N4358, N4353, N2596, N2551);
and AND3 (N4359, N4354, N364, N1181);
and AND4 (N4360, N4352, N3470, N1477, N1404);
nor NOR3 (N4361, N4355, N3863, N345);
xor XOR2 (N4362, N4351, N3118);
not NOT1 (N4363, N4331);
not NOT1 (N4364, N4362);
or OR2 (N4365, N4361, N1342);
nor NOR4 (N4366, N4358, N3934, N1433, N3268);
and AND4 (N4367, N4359, N2826, N1325, N1239);
not NOT1 (N4368, N4366);
buf BUF1 (N4369, N4367);
buf BUF1 (N4370, N4363);
or OR3 (N4371, N4348, N2511, N2339);
xor XOR2 (N4372, N4368, N927);
xor XOR2 (N4373, N4370, N1565);
nand NAND2 (N4374, N4364, N1357);
or OR4 (N4375, N4360, N1467, N3857, N2945);
and AND4 (N4376, N4349, N127, N4179, N1348);
buf BUF1 (N4377, N4357);
nand NAND2 (N4378, N4365, N802);
xor XOR2 (N4379, N4369, N249);
not NOT1 (N4380, N4371);
nand NAND3 (N4381, N4347, N1926, N1280);
nor NOR3 (N4382, N4381, N3259, N1573);
nor NOR4 (N4383, N4377, N742, N198, N1169);
buf BUF1 (N4384, N4382);
nand NAND3 (N4385, N4384, N2243, N56);
nand NAND2 (N4386, N4378, N59);
xor XOR2 (N4387, N4375, N3150);
xor XOR2 (N4388, N4376, N692);
or OR3 (N4389, N4383, N397, N1736);
nor NOR4 (N4390, N4386, N4013, N3006, N3046);
nor NOR3 (N4391, N4372, N978, N2978);
and AND3 (N4392, N4390, N2157, N3040);
or OR3 (N4393, N4392, N3346, N3267);
xor XOR2 (N4394, N4393, N487);
xor XOR2 (N4395, N4373, N249);
and AND2 (N4396, N4395, N1087);
or OR3 (N4397, N4380, N3629, N87);
nand NAND3 (N4398, N4388, N2395, N2893);
xor XOR2 (N4399, N4374, N3117);
not NOT1 (N4400, N4379);
or OR2 (N4401, N4394, N3201);
and AND4 (N4402, N4397, N1509, N2836, N942);
nor NOR3 (N4403, N4389, N1913, N111);
nor NOR2 (N4404, N4385, N632);
nand NAND3 (N4405, N4398, N3224, N3530);
or OR4 (N4406, N4405, N2773, N1670, N3898);
and AND3 (N4407, N4387, N3746, N2375);
nand NAND2 (N4408, N4401, N2488);
not NOT1 (N4409, N4402);
buf BUF1 (N4410, N4396);
and AND3 (N4411, N4410, N3563, N2049);
and AND2 (N4412, N4411, N2061);
xor XOR2 (N4413, N4403, N1647);
xor XOR2 (N4414, N4408, N2590);
and AND2 (N4415, N4406, N1839);
buf BUF1 (N4416, N4414);
nand NAND3 (N4417, N4415, N3449, N2947);
xor XOR2 (N4418, N4412, N2329);
nand NAND3 (N4419, N4404, N2537, N1853);
nand NAND3 (N4420, N4413, N36, N3337);
xor XOR2 (N4421, N4407, N3234);
or OR2 (N4422, N4421, N1085);
xor XOR2 (N4423, N4418, N1337);
buf BUF1 (N4424, N4399);
nand NAND2 (N4425, N4400, N3168);
buf BUF1 (N4426, N4416);
not NOT1 (N4427, N4424);
not NOT1 (N4428, N4420);
or OR2 (N4429, N4425, N3469);
nand NAND2 (N4430, N4429, N1973);
or OR3 (N4431, N4428, N497, N451);
not NOT1 (N4432, N4430);
or OR4 (N4433, N4417, N2731, N4237, N4376);
or OR2 (N4434, N4423, N3592);
not NOT1 (N4435, N4409);
buf BUF1 (N4436, N4391);
buf BUF1 (N4437, N4422);
buf BUF1 (N4438, N4434);
not NOT1 (N4439, N4427);
not NOT1 (N4440, N4426);
buf BUF1 (N4441, N4431);
nor NOR4 (N4442, N4435, N1752, N2667, N1744);
buf BUF1 (N4443, N4439);
buf BUF1 (N4444, N4441);
nand NAND2 (N4445, N4443, N1728);
not NOT1 (N4446, N4436);
not NOT1 (N4447, N4432);
nor NOR4 (N4448, N4444, N1095, N3821, N3293);
and AND2 (N4449, N4438, N2207);
not NOT1 (N4450, N4448);
nand NAND2 (N4451, N4440, N4210);
nand NAND2 (N4452, N4447, N158);
buf BUF1 (N4453, N4449);
or OR3 (N4454, N4450, N3550, N1043);
xor XOR2 (N4455, N4453, N3086);
nand NAND3 (N4456, N4454, N3051, N2101);
nand NAND2 (N4457, N4437, N2488);
xor XOR2 (N4458, N4455, N841);
nand NAND3 (N4459, N4451, N75, N1382);
nor NOR4 (N4460, N4456, N753, N2019, N526);
and AND4 (N4461, N4419, N165, N3769, N1834);
nand NAND4 (N4462, N4445, N165, N4188, N3361);
not NOT1 (N4463, N4461);
or OR3 (N4464, N4459, N3024, N3235);
not NOT1 (N4465, N4460);
nor NOR3 (N4466, N4446, N373, N1421);
nand NAND3 (N4467, N4433, N3104, N2958);
and AND3 (N4468, N4457, N73, N418);
nand NAND4 (N4469, N4467, N585, N3581, N1457);
not NOT1 (N4470, N4464);
or OR2 (N4471, N4470, N471);
nor NOR2 (N4472, N4466, N3872);
nand NAND3 (N4473, N4442, N2466, N2336);
nor NOR2 (N4474, N4462, N1565);
buf BUF1 (N4475, N4472);
nor NOR2 (N4476, N4475, N2539);
buf BUF1 (N4477, N4476);
buf BUF1 (N4478, N4465);
not NOT1 (N4479, N4478);
or OR3 (N4480, N4474, N262, N4316);
not NOT1 (N4481, N4469);
xor XOR2 (N4482, N4473, N1436);
and AND2 (N4483, N4479, N3404);
nor NOR3 (N4484, N4477, N4432, N3492);
nor NOR3 (N4485, N4481, N4436, N4390);
buf BUF1 (N4486, N4458);
nor NOR4 (N4487, N4483, N980, N4258, N2331);
not NOT1 (N4488, N4482);
or OR3 (N4489, N4487, N1669, N4189);
or OR4 (N4490, N4468, N1660, N592, N2567);
not NOT1 (N4491, N4484);
nand NAND2 (N4492, N4463, N4023);
nor NOR3 (N4493, N4491, N1891, N1391);
xor XOR2 (N4494, N4493, N364);
nand NAND2 (N4495, N4471, N3254);
and AND4 (N4496, N4486, N3344, N1652, N3329);
not NOT1 (N4497, N4495);
xor XOR2 (N4498, N4494, N2893);
not NOT1 (N4499, N4496);
nor NOR4 (N4500, N4492, N2047, N2158, N2444);
nand NAND2 (N4501, N4488, N2088);
and AND4 (N4502, N4490, N390, N2251, N3242);
or OR4 (N4503, N4502, N1455, N126, N4460);
xor XOR2 (N4504, N4489, N872);
xor XOR2 (N4505, N4504, N3751);
xor XOR2 (N4506, N4498, N495);
and AND2 (N4507, N4503, N3695);
nor NOR4 (N4508, N4505, N1946, N4347, N3778);
nand NAND3 (N4509, N4508, N2759, N3871);
not NOT1 (N4510, N4507);
xor XOR2 (N4511, N4452, N2941);
or OR4 (N4512, N4511, N1322, N962, N2091);
xor XOR2 (N4513, N4506, N2614);
xor XOR2 (N4514, N4512, N1433);
nand NAND4 (N4515, N4514, N982, N8, N3225);
and AND3 (N4516, N4485, N1698, N623);
or OR2 (N4517, N4497, N838);
and AND4 (N4518, N4515, N1347, N206, N2591);
nand NAND2 (N4519, N4509, N596);
xor XOR2 (N4520, N4510, N2468);
nor NOR4 (N4521, N4499, N1058, N1535, N577);
not NOT1 (N4522, N4516);
or OR3 (N4523, N4522, N3244, N3065);
not NOT1 (N4524, N4519);
and AND4 (N4525, N4524, N1739, N1690, N4026);
buf BUF1 (N4526, N4520);
or OR3 (N4527, N4500, N902, N530);
xor XOR2 (N4528, N4518, N3657);
and AND2 (N4529, N4517, N1443);
nor NOR3 (N4530, N4525, N1627, N1929);
or OR2 (N4531, N4527, N3750);
and AND3 (N4532, N4526, N1556, N138);
nor NOR2 (N4533, N4529, N3126);
or OR4 (N4534, N4523, N1454, N2813, N4437);
buf BUF1 (N4535, N4528);
nand NAND4 (N4536, N4513, N3689, N2352, N1666);
not NOT1 (N4537, N4530);
and AND4 (N4538, N4532, N2159, N9, N3710);
buf BUF1 (N4539, N4531);
or OR4 (N4540, N4537, N2002, N1252, N1254);
or OR4 (N4541, N4521, N3664, N2741, N3411);
nand NAND4 (N4542, N4538, N2176, N294, N3396);
nor NOR2 (N4543, N4535, N747);
buf BUF1 (N4544, N4480);
buf BUF1 (N4545, N4534);
and AND3 (N4546, N4545, N2151, N4149);
xor XOR2 (N4547, N4542, N2149);
or OR4 (N4548, N4539, N1462, N4420, N2906);
or OR3 (N4549, N4540, N450, N605);
nor NOR2 (N4550, N4546, N119);
not NOT1 (N4551, N4550);
buf BUF1 (N4552, N4551);
or OR3 (N4553, N4501, N3118, N3074);
nor NOR4 (N4554, N4533, N785, N4426, N3161);
xor XOR2 (N4555, N4553, N2068);
not NOT1 (N4556, N4547);
and AND3 (N4557, N4554, N2460, N2902);
and AND3 (N4558, N4557, N2999, N2886);
not NOT1 (N4559, N4548);
or OR3 (N4560, N4536, N551, N541);
and AND3 (N4561, N4558, N3624, N686);
or OR3 (N4562, N4541, N232, N704);
or OR4 (N4563, N4555, N530, N3783, N3835);
not NOT1 (N4564, N4559);
and AND4 (N4565, N4543, N2615, N3650, N2621);
nor NOR4 (N4566, N4544, N2196, N2598, N4240);
and AND2 (N4567, N4561, N1854);
xor XOR2 (N4568, N4549, N1029);
nor NOR3 (N4569, N4564, N3599, N2468);
buf BUF1 (N4570, N4552);
nor NOR3 (N4571, N4570, N2928, N1234);
not NOT1 (N4572, N4571);
nor NOR4 (N4573, N4565, N2063, N4219, N607);
xor XOR2 (N4574, N4560, N3765);
or OR3 (N4575, N4562, N1878, N3946);
nand NAND3 (N4576, N4574, N1937, N1402);
and AND4 (N4577, N4568, N3956, N1633, N228);
nand NAND3 (N4578, N4563, N3028, N1674);
not NOT1 (N4579, N4575);
nand NAND3 (N4580, N4566, N3076, N2481);
buf BUF1 (N4581, N4576);
xor XOR2 (N4582, N4572, N2090);
nand NAND4 (N4583, N4556, N805, N1236, N3300);
nand NAND2 (N4584, N4580, N4344);
not NOT1 (N4585, N4581);
nand NAND3 (N4586, N4578, N3142, N3330);
or OR4 (N4587, N4582, N3944, N3656, N4044);
nor NOR4 (N4588, N4569, N131, N3522, N2350);
xor XOR2 (N4589, N4583, N4397);
not NOT1 (N4590, N4584);
xor XOR2 (N4591, N4579, N1287);
nand NAND3 (N4592, N4567, N4001, N3613);
buf BUF1 (N4593, N4585);
or OR4 (N4594, N4587, N4235, N3627, N732);
not NOT1 (N4595, N4586);
not NOT1 (N4596, N4589);
nor NOR3 (N4597, N4594, N885, N4119);
not NOT1 (N4598, N4593);
and AND2 (N4599, N4598, N2001);
and AND2 (N4600, N4599, N713);
or OR3 (N4601, N4591, N1847, N3553);
buf BUF1 (N4602, N4597);
nand NAND2 (N4603, N4592, N3991);
or OR3 (N4604, N4588, N2949, N2491);
buf BUF1 (N4605, N4577);
xor XOR2 (N4606, N4573, N632);
or OR3 (N4607, N4600, N3803, N1269);
and AND4 (N4608, N4590, N991, N1059, N2950);
not NOT1 (N4609, N4602);
not NOT1 (N4610, N4604);
or OR4 (N4611, N4606, N1081, N4294, N3860);
xor XOR2 (N4612, N4603, N3016);
and AND3 (N4613, N4596, N2790, N3195);
buf BUF1 (N4614, N4601);
nand NAND3 (N4615, N4613, N488, N3240);
and AND3 (N4616, N4595, N2941, N1135);
or OR3 (N4617, N4608, N4599, N4086);
or OR4 (N4618, N4612, N2456, N2018, N3102);
nand NAND2 (N4619, N4611, N3378);
nand NAND2 (N4620, N4609, N2877);
and AND2 (N4621, N4618, N1093);
nor NOR3 (N4622, N4621, N2189, N2730);
not NOT1 (N4623, N4610);
nand NAND3 (N4624, N4623, N2236, N2181);
buf BUF1 (N4625, N4616);
or OR4 (N4626, N4605, N1944, N1040, N1074);
nor NOR2 (N4627, N4626, N1748);
not NOT1 (N4628, N4619);
not NOT1 (N4629, N4617);
nand NAND4 (N4630, N4624, N495, N4184, N3591);
and AND2 (N4631, N4622, N2549);
nor NOR2 (N4632, N4607, N3054);
not NOT1 (N4633, N4631);
buf BUF1 (N4634, N4630);
not NOT1 (N4635, N4633);
nand NAND4 (N4636, N4615, N2500, N899, N986);
nor NOR4 (N4637, N4634, N923, N1584, N3186);
not NOT1 (N4638, N4628);
xor XOR2 (N4639, N4625, N56);
nor NOR2 (N4640, N4638, N4449);
buf BUF1 (N4641, N4627);
not NOT1 (N4642, N4632);
or OR4 (N4643, N4641, N1782, N4061, N3297);
nand NAND2 (N4644, N4639, N2898);
nand NAND3 (N4645, N4620, N3584, N4006);
or OR3 (N4646, N4614, N317, N1289);
and AND4 (N4647, N4643, N4032, N2221, N4390);
nor NOR3 (N4648, N4640, N601, N1682);
or OR2 (N4649, N4636, N1952);
xor XOR2 (N4650, N4644, N94);
and AND4 (N4651, N4647, N3883, N3612, N3268);
nand NAND4 (N4652, N4637, N2563, N2901, N4279);
xor XOR2 (N4653, N4635, N4355);
xor XOR2 (N4654, N4645, N299);
and AND2 (N4655, N4648, N2461);
or OR2 (N4656, N4642, N1431);
not NOT1 (N4657, N4654);
or OR4 (N4658, N4651, N4321, N820, N4373);
and AND2 (N4659, N4652, N3223);
buf BUF1 (N4660, N4659);
nand NAND4 (N4661, N4650, N2852, N1793, N781);
buf BUF1 (N4662, N4658);
or OR3 (N4663, N4649, N3770, N3154);
not NOT1 (N4664, N4653);
nor NOR2 (N4665, N4629, N3684);
and AND4 (N4666, N4661, N1071, N4591, N3337);
buf BUF1 (N4667, N4660);
xor XOR2 (N4668, N4657, N947);
and AND3 (N4669, N4662, N2101, N1329);
nand NAND4 (N4670, N4646, N3021, N2710, N1603);
and AND3 (N4671, N4665, N2376, N1733);
nand NAND2 (N4672, N4664, N1577);
xor XOR2 (N4673, N4671, N2699);
nor NOR2 (N4674, N4666, N1908);
nor NOR2 (N4675, N4672, N3338);
and AND2 (N4676, N4668, N469);
nand NAND4 (N4677, N4673, N583, N2106, N3149);
nor NOR4 (N4678, N4655, N4207, N1097, N4025);
or OR3 (N4679, N4667, N3885, N1134);
or OR4 (N4680, N4677, N2412, N968, N2702);
buf BUF1 (N4681, N4678);
or OR3 (N4682, N4656, N528, N355);
not NOT1 (N4683, N4680);
not NOT1 (N4684, N4670);
xor XOR2 (N4685, N4681, N901);
or OR4 (N4686, N4683, N2912, N1173, N1997);
and AND2 (N4687, N4669, N1629);
buf BUF1 (N4688, N4684);
nor NOR3 (N4689, N4676, N4249, N40);
buf BUF1 (N4690, N4679);
not NOT1 (N4691, N4682);
nor NOR4 (N4692, N4674, N842, N263, N2368);
or OR3 (N4693, N4686, N1888, N3938);
or OR2 (N4694, N4687, N2545);
not NOT1 (N4695, N4693);
or OR2 (N4696, N4692, N3869);
not NOT1 (N4697, N4696);
not NOT1 (N4698, N4675);
nor NOR3 (N4699, N4663, N3947, N460);
or OR4 (N4700, N4689, N11, N1877, N2852);
not NOT1 (N4701, N4694);
xor XOR2 (N4702, N4685, N2128);
and AND3 (N4703, N4700, N2773, N2519);
nand NAND3 (N4704, N4701, N2725, N4073);
nor NOR4 (N4705, N4698, N1970, N228, N1259);
not NOT1 (N4706, N4688);
buf BUF1 (N4707, N4703);
xor XOR2 (N4708, N4695, N4194);
nor NOR3 (N4709, N4704, N4314, N2469);
not NOT1 (N4710, N4699);
nor NOR3 (N4711, N4710, N4142, N1701);
nor NOR4 (N4712, N4705, N1175, N3458, N1316);
and AND4 (N4713, N4711, N3386, N1711, N359);
not NOT1 (N4714, N4702);
or OR4 (N4715, N4709, N374, N2684, N3887);
and AND4 (N4716, N4707, N3507, N88, N734);
or OR4 (N4717, N4706, N2550, N155, N2069);
and AND2 (N4718, N4712, N240);
nor NOR4 (N4719, N4713, N836, N3120, N3885);
buf BUF1 (N4720, N4714);
nand NAND3 (N4721, N4720, N799, N1406);
nand NAND3 (N4722, N4717, N1684, N4264);
buf BUF1 (N4723, N4716);
nand NAND3 (N4724, N4708, N72, N4524);
buf BUF1 (N4725, N4690);
xor XOR2 (N4726, N4697, N4442);
xor XOR2 (N4727, N4724, N1601);
and AND2 (N4728, N4722, N1750);
xor XOR2 (N4729, N4718, N1770);
xor XOR2 (N4730, N4729, N3945);
xor XOR2 (N4731, N4730, N2373);
or OR3 (N4732, N4723, N3589, N2030);
xor XOR2 (N4733, N4719, N2802);
nand NAND3 (N4734, N4691, N1607, N3879);
and AND4 (N4735, N4734, N1007, N3560, N416);
not NOT1 (N4736, N4731);
not NOT1 (N4737, N4726);
and AND3 (N4738, N4728, N1296, N890);
not NOT1 (N4739, N4736);
or OR4 (N4740, N4721, N4236, N2443, N647);
and AND4 (N4741, N4725, N4425, N2950, N373);
not NOT1 (N4742, N4740);
nand NAND4 (N4743, N4715, N1484, N686, N3216);
buf BUF1 (N4744, N4735);
xor XOR2 (N4745, N4738, N1777);
buf BUF1 (N4746, N4732);
buf BUF1 (N4747, N4742);
not NOT1 (N4748, N4743);
nand NAND2 (N4749, N4746, N596);
nand NAND3 (N4750, N4739, N3057, N4098);
or OR4 (N4751, N4737, N745, N4663, N2280);
nor NOR3 (N4752, N4727, N66, N1974);
buf BUF1 (N4753, N4745);
and AND4 (N4754, N4749, N227, N3185, N2576);
xor XOR2 (N4755, N4741, N89);
buf BUF1 (N4756, N4751);
nand NAND3 (N4757, N4754, N140, N3476);
nand NAND2 (N4758, N4757, N2241);
xor XOR2 (N4759, N4753, N2553);
and AND2 (N4760, N4752, N2215);
buf BUF1 (N4761, N4750);
not NOT1 (N4762, N4748);
and AND4 (N4763, N4744, N3899, N3944, N1852);
xor XOR2 (N4764, N4762, N1906);
and AND4 (N4765, N4761, N3528, N3471, N3769);
or OR4 (N4766, N4763, N2871, N4359, N2209);
or OR3 (N4767, N4755, N3246, N121);
nor NOR2 (N4768, N4733, N2410);
nor NOR2 (N4769, N4758, N2129);
buf BUF1 (N4770, N4767);
nor NOR2 (N4771, N4765, N577);
nand NAND4 (N4772, N4766, N420, N4717, N875);
xor XOR2 (N4773, N4768, N4171);
xor XOR2 (N4774, N4747, N2228);
and AND3 (N4775, N4772, N3622, N4466);
or OR2 (N4776, N4760, N3413);
or OR2 (N4777, N4771, N3625);
and AND4 (N4778, N4775, N1935, N1077, N4601);
and AND4 (N4779, N4773, N2769, N2188, N1332);
and AND4 (N4780, N4759, N2366, N304, N996);
nand NAND4 (N4781, N4770, N2526, N3945, N1647);
not NOT1 (N4782, N4776);
nand NAND3 (N4783, N4774, N394, N4064);
xor XOR2 (N4784, N4769, N2024);
xor XOR2 (N4785, N4783, N3056);
xor XOR2 (N4786, N4784, N3899);
and AND4 (N4787, N4764, N3998, N2938, N940);
nand NAND4 (N4788, N4787, N4735, N4486, N2485);
nor NOR4 (N4789, N4777, N108, N4669, N2536);
and AND3 (N4790, N4789, N3970, N605);
nand NAND3 (N4791, N4756, N1000, N2685);
nand NAND3 (N4792, N4779, N3350, N4415);
xor XOR2 (N4793, N4778, N1478);
nor NOR4 (N4794, N4785, N1666, N313, N4157);
buf BUF1 (N4795, N4793);
and AND2 (N4796, N4792, N3624);
or OR2 (N4797, N4790, N2844);
or OR4 (N4798, N4780, N3187, N3863, N2045);
and AND4 (N4799, N4782, N1866, N2421, N3643);
not NOT1 (N4800, N4781);
xor XOR2 (N4801, N4788, N2429);
buf BUF1 (N4802, N4791);
not NOT1 (N4803, N4802);
xor XOR2 (N4804, N4803, N1236);
buf BUF1 (N4805, N4797);
not NOT1 (N4806, N4794);
and AND2 (N4807, N4801, N3849);
buf BUF1 (N4808, N4804);
xor XOR2 (N4809, N4786, N1655);
or OR4 (N4810, N4808, N1089, N3999, N3006);
not NOT1 (N4811, N4795);
not NOT1 (N4812, N4796);
buf BUF1 (N4813, N4799);
nand NAND4 (N4814, N4807, N4360, N4713, N484);
xor XOR2 (N4815, N4805, N861);
xor XOR2 (N4816, N4810, N2035);
and AND2 (N4817, N4813, N1867);
not NOT1 (N4818, N4811);
and AND4 (N4819, N4815, N3265, N83, N1140);
or OR4 (N4820, N4816, N1245, N4542, N2454);
or OR4 (N4821, N4818, N222, N1433, N3460);
not NOT1 (N4822, N4800);
xor XOR2 (N4823, N4820, N313);
or OR2 (N4824, N4806, N690);
or OR4 (N4825, N4819, N3337, N2771, N3670);
nor NOR3 (N4826, N4809, N4523, N2339);
nor NOR2 (N4827, N4798, N3639);
or OR2 (N4828, N4827, N799);
nand NAND3 (N4829, N4817, N177, N3129);
not NOT1 (N4830, N4821);
not NOT1 (N4831, N4828);
or OR2 (N4832, N4823, N2171);
buf BUF1 (N4833, N4824);
not NOT1 (N4834, N4822);
or OR2 (N4835, N4812, N1221);
nor NOR4 (N4836, N4832, N1167, N2549, N103);
and AND2 (N4837, N4829, N3549);
buf BUF1 (N4838, N4835);
nand NAND4 (N4839, N4814, N2608, N4587, N1544);
buf BUF1 (N4840, N4837);
nand NAND4 (N4841, N4833, N3054, N4041, N4824);
xor XOR2 (N4842, N4830, N1741);
nor NOR4 (N4843, N4831, N634, N4247, N962);
nand NAND2 (N4844, N4841, N147);
or OR4 (N4845, N4843, N1940, N1030, N595);
buf BUF1 (N4846, N4836);
nand NAND2 (N4847, N4826, N3137);
nor NOR3 (N4848, N4846, N2028, N1915);
and AND3 (N4849, N4842, N4289, N4599);
nor NOR3 (N4850, N4825, N4005, N1760);
and AND2 (N4851, N4844, N317);
buf BUF1 (N4852, N4834);
or OR3 (N4853, N4838, N2105, N839);
or OR4 (N4854, N4850, N3260, N310, N2831);
nand NAND4 (N4855, N4845, N2189, N4645, N794);
nand NAND2 (N4856, N4847, N1684);
buf BUF1 (N4857, N4849);
buf BUF1 (N4858, N4840);
xor XOR2 (N4859, N4852, N306);
nor NOR4 (N4860, N4856, N927, N2430, N1871);
xor XOR2 (N4861, N4860, N2872);
and AND4 (N4862, N4853, N3660, N4699, N1244);
buf BUF1 (N4863, N4862);
or OR4 (N4864, N4851, N865, N530, N2198);
xor XOR2 (N4865, N4855, N4321);
and AND3 (N4866, N4864, N3179, N549);
buf BUF1 (N4867, N4857);
nor NOR4 (N4868, N4865, N1191, N1179, N4390);
or OR2 (N4869, N4854, N210);
not NOT1 (N4870, N4858);
and AND4 (N4871, N4870, N267, N67, N4055);
or OR2 (N4872, N4868, N3925);
and AND3 (N4873, N4869, N2922, N4646);
nor NOR4 (N4874, N4866, N4633, N985, N683);
or OR2 (N4875, N4839, N1957);
not NOT1 (N4876, N4873);
or OR4 (N4877, N4872, N2610, N3182, N1196);
xor XOR2 (N4878, N4859, N4392);
or OR3 (N4879, N4876, N1070, N2360);
nor NOR4 (N4880, N4879, N263, N2271, N1352);
xor XOR2 (N4881, N4878, N3297);
nor NOR2 (N4882, N4880, N728);
and AND2 (N4883, N4848, N1933);
and AND3 (N4884, N4881, N967, N814);
buf BUF1 (N4885, N4884);
nand NAND3 (N4886, N4867, N4627, N2912);
nand NAND2 (N4887, N4882, N1179);
nor NOR2 (N4888, N4883, N3666);
nor NOR4 (N4889, N4887, N1150, N3556, N2977);
or OR4 (N4890, N4886, N1760, N3878, N3982);
nor NOR4 (N4891, N4875, N2167, N1061, N4324);
buf BUF1 (N4892, N4891);
xor XOR2 (N4893, N4861, N1105);
nor NOR4 (N4894, N4893, N524, N1942, N920);
nor NOR3 (N4895, N4871, N2541, N1684);
nand NAND2 (N4896, N4874, N4498);
xor XOR2 (N4897, N4896, N1671);
nand NAND4 (N4898, N4897, N4870, N4675, N254);
nor NOR4 (N4899, N4888, N52, N1744, N184);
or OR3 (N4900, N4877, N1168, N2266);
not NOT1 (N4901, N4895);
not NOT1 (N4902, N4863);
nand NAND2 (N4903, N4892, N2524);
buf BUF1 (N4904, N4903);
buf BUF1 (N4905, N4899);
nor NOR2 (N4906, N4902, N4310);
xor XOR2 (N4907, N4906, N506);
buf BUF1 (N4908, N4901);
nand NAND3 (N4909, N4905, N2962, N44);
or OR2 (N4910, N4898, N2888);
nand NAND4 (N4911, N4900, N3565, N2791, N3781);
xor XOR2 (N4912, N4910, N164);
or OR3 (N4913, N4907, N4447, N2766);
not NOT1 (N4914, N4909);
xor XOR2 (N4915, N4914, N1486);
nand NAND4 (N4916, N4894, N2732, N3739, N4738);
xor XOR2 (N4917, N4889, N3988);
and AND4 (N4918, N4890, N1048, N1712, N2634);
xor XOR2 (N4919, N4916, N4569);
nor NOR3 (N4920, N4917, N1932, N2386);
or OR3 (N4921, N4913, N733, N3637);
and AND4 (N4922, N4918, N442, N2610, N2046);
nor NOR3 (N4923, N4922, N3547, N722);
not NOT1 (N4924, N4911);
buf BUF1 (N4925, N4924);
and AND2 (N4926, N4919, N2602);
xor XOR2 (N4927, N4885, N3992);
and AND3 (N4928, N4921, N616, N2574);
not NOT1 (N4929, N4927);
nor NOR4 (N4930, N4915, N1949, N16, N2908);
nor NOR2 (N4931, N4923, N932);
nor NOR4 (N4932, N4904, N2186, N4131, N1125);
nor NOR4 (N4933, N4931, N1291, N1760, N1534);
nand NAND3 (N4934, N4908, N2665, N3347);
nand NAND4 (N4935, N4929, N486, N3302, N1227);
and AND3 (N4936, N4930, N3233, N361);
nand NAND4 (N4937, N4932, N1942, N1857, N190);
not NOT1 (N4938, N4935);
and AND3 (N4939, N4933, N630, N1805);
and AND4 (N4940, N4925, N1024, N775, N66);
buf BUF1 (N4941, N4940);
xor XOR2 (N4942, N4938, N3184);
xor XOR2 (N4943, N4934, N1118);
nor NOR2 (N4944, N4920, N2187);
and AND3 (N4945, N4912, N557, N217);
or OR2 (N4946, N4939, N3478);
or OR4 (N4947, N4941, N4916, N2999, N1596);
xor XOR2 (N4948, N4928, N4848);
nand NAND4 (N4949, N4942, N954, N2264, N1769);
and AND4 (N4950, N4937, N1960, N4703, N708);
buf BUF1 (N4951, N4949);
xor XOR2 (N4952, N4926, N126);
or OR4 (N4953, N4950, N239, N2102, N1879);
nor NOR2 (N4954, N4948, N105);
or OR4 (N4955, N4953, N76, N1645, N1330);
nor NOR4 (N4956, N4943, N1624, N758, N2988);
xor XOR2 (N4957, N4945, N4873);
xor XOR2 (N4958, N4946, N4490);
nand NAND2 (N4959, N4944, N4589);
nor NOR4 (N4960, N4947, N2183, N1147, N4436);
buf BUF1 (N4961, N4951);
buf BUF1 (N4962, N4936);
and AND4 (N4963, N4958, N2995, N3649, N3535);
buf BUF1 (N4964, N4960);
nor NOR3 (N4965, N4955, N701, N1823);
xor XOR2 (N4966, N4962, N2159);
xor XOR2 (N4967, N4966, N4411);
xor XOR2 (N4968, N4965, N662);
and AND3 (N4969, N4952, N4568, N2642);
xor XOR2 (N4970, N4956, N2497);
nor NOR4 (N4971, N4954, N3861, N4497, N229);
not NOT1 (N4972, N4963);
and AND2 (N4973, N4959, N4296);
or OR2 (N4974, N4972, N4333);
and AND3 (N4975, N4961, N1335, N3768);
nor NOR3 (N4976, N4971, N3168, N758);
not NOT1 (N4977, N4973);
buf BUF1 (N4978, N4957);
nor NOR4 (N4979, N4968, N2357, N242, N71);
xor XOR2 (N4980, N4979, N3888);
xor XOR2 (N4981, N4969, N1851);
xor XOR2 (N4982, N4977, N1456);
buf BUF1 (N4983, N4970);
nand NAND4 (N4984, N4975, N2180, N495, N475);
nor NOR3 (N4985, N4982, N274, N524);
buf BUF1 (N4986, N4981);
or OR3 (N4987, N4974, N2842, N132);
nor NOR4 (N4988, N4980, N3129, N3576, N3608);
nand NAND4 (N4989, N4985, N1010, N4765, N1658);
buf BUF1 (N4990, N4967);
xor XOR2 (N4991, N4988, N3848);
nor NOR2 (N4992, N4990, N1374);
or OR2 (N4993, N4976, N1726);
and AND4 (N4994, N4986, N4380, N4422, N4492);
not NOT1 (N4995, N4987);
xor XOR2 (N4996, N4964, N4516);
or OR4 (N4997, N4993, N2920, N2242, N3595);
nor NOR4 (N4998, N4984, N4191, N2689, N4699);
and AND3 (N4999, N4978, N139, N4226);
not NOT1 (N5000, N4989);
nor NOR2 (N5001, N4994, N2567);
buf BUF1 (N5002, N4995);
and AND3 (N5003, N4983, N1548, N1802);
buf BUF1 (N5004, N5001);
xor XOR2 (N5005, N5003, N4120);
and AND3 (N5006, N5002, N3179, N2821);
nand NAND2 (N5007, N4992, N611);
and AND3 (N5008, N4996, N2825, N1970);
not NOT1 (N5009, N4991);
buf BUF1 (N5010, N5009);
and AND3 (N5011, N5008, N2094, N3742);
not NOT1 (N5012, N4997);
xor XOR2 (N5013, N4999, N1235);
xor XOR2 (N5014, N5007, N2369);
nand NAND2 (N5015, N5014, N357);
nand NAND3 (N5016, N5004, N880, N3585);
nand NAND2 (N5017, N5012, N3167);
and AND2 (N5018, N5000, N4495);
or OR4 (N5019, N5006, N2509, N2102, N3821);
nand NAND4 (N5020, N5016, N2086, N4153, N2102);
buf BUF1 (N5021, N5018);
nand NAND3 (N5022, N5017, N3542, N116);
nand NAND4 (N5023, N5015, N2817, N1791, N579);
buf BUF1 (N5024, N5005);
nand NAND3 (N5025, N5021, N340, N2291);
nand NAND2 (N5026, N5023, N3816);
nor NOR3 (N5027, N5025, N291, N4054);
xor XOR2 (N5028, N5010, N957);
buf BUF1 (N5029, N5027);
not NOT1 (N5030, N5013);
xor XOR2 (N5031, N5029, N3119);
buf BUF1 (N5032, N5019);
nor NOR3 (N5033, N4998, N4952, N2803);
or OR4 (N5034, N5033, N3053, N3471, N4930);
nand NAND2 (N5035, N5034, N4288);
and AND4 (N5036, N5035, N2219, N381, N1414);
and AND2 (N5037, N5020, N3305);
or OR2 (N5038, N5024, N3044);
or OR3 (N5039, N5011, N3291, N2567);
xor XOR2 (N5040, N5028, N2454);
nand NAND2 (N5041, N5036, N3273);
nand NAND3 (N5042, N5026, N145, N157);
or OR4 (N5043, N5041, N3466, N4960, N3900);
buf BUF1 (N5044, N5042);
and AND3 (N5045, N5040, N2567, N36);
and AND4 (N5046, N5032, N2538, N2646, N3819);
not NOT1 (N5047, N5037);
or OR2 (N5048, N5038, N4725);
or OR3 (N5049, N5030, N4522, N3083);
buf BUF1 (N5050, N5047);
or OR4 (N5051, N5022, N473, N3399, N1196);
buf BUF1 (N5052, N5049);
and AND4 (N5053, N5048, N944, N932, N5044);
buf BUF1 (N5054, N1084);
or OR4 (N5055, N5045, N4851, N2581, N921);
and AND4 (N5056, N5055, N2561, N1082, N2534);
nand NAND4 (N5057, N5043, N2202, N1937, N4098);
and AND2 (N5058, N5056, N2916);
buf BUF1 (N5059, N5053);
nor NOR4 (N5060, N5059, N3052, N4546, N3591);
not NOT1 (N5061, N5054);
or OR2 (N5062, N5039, N4834);
nor NOR2 (N5063, N5062, N1500);
and AND3 (N5064, N5060, N515, N953);
xor XOR2 (N5065, N5061, N3346);
and AND4 (N5066, N5064, N2002, N1412, N1960);
or OR3 (N5067, N5051, N4894, N1064);
buf BUF1 (N5068, N5063);
buf BUF1 (N5069, N5046);
and AND3 (N5070, N5031, N1883, N1496);
buf BUF1 (N5071, N5066);
or OR3 (N5072, N5052, N2311, N3642);
buf BUF1 (N5073, N5069);
or OR3 (N5074, N5065, N4970, N3223);
xor XOR2 (N5075, N5058, N2486);
buf BUF1 (N5076, N5073);
nand NAND4 (N5077, N5057, N295, N4041, N2443);
and AND2 (N5078, N5072, N4872);
nand NAND4 (N5079, N5068, N3917, N1308, N4278);
buf BUF1 (N5080, N5071);
and AND2 (N5081, N5079, N1845);
xor XOR2 (N5082, N5076, N507);
and AND3 (N5083, N5077, N3161, N955);
nand NAND3 (N5084, N5050, N2704, N5073);
and AND4 (N5085, N5074, N4626, N4277, N3195);
xor XOR2 (N5086, N5070, N2288);
or OR3 (N5087, N5080, N4835, N1421);
xor XOR2 (N5088, N5087, N2783);
nor NOR4 (N5089, N5088, N3118, N3776, N4303);
buf BUF1 (N5090, N5089);
not NOT1 (N5091, N5083);
or OR3 (N5092, N5082, N1638, N4756);
buf BUF1 (N5093, N5067);
nand NAND4 (N5094, N5084, N2642, N3212, N4778);
and AND3 (N5095, N5093, N3802, N1904);
nor NOR2 (N5096, N5095, N1857);
xor XOR2 (N5097, N5085, N4082);
buf BUF1 (N5098, N5091);
and AND4 (N5099, N5096, N3030, N4091, N4956);
nand NAND4 (N5100, N5081, N1202, N2877, N4237);
or OR4 (N5101, N5092, N4080, N46, N880);
xor XOR2 (N5102, N5099, N1633);
nand NAND4 (N5103, N5102, N2485, N985, N4232);
nand NAND3 (N5104, N5086, N2099, N838);
nor NOR4 (N5105, N5094, N2920, N3270, N1271);
nand NAND4 (N5106, N5100, N3739, N1678, N4120);
or OR4 (N5107, N5101, N2509, N2667, N3910);
or OR2 (N5108, N5090, N3392);
nor NOR2 (N5109, N5078, N1587);
nand NAND2 (N5110, N5103, N3870);
buf BUF1 (N5111, N5106);
not NOT1 (N5112, N5097);
not NOT1 (N5113, N5104);
buf BUF1 (N5114, N5075);
xor XOR2 (N5115, N5111, N2453);
xor XOR2 (N5116, N5109, N2380);
buf BUF1 (N5117, N5116);
nor NOR3 (N5118, N5117, N757, N3067);
or OR4 (N5119, N5118, N1575, N2470, N3134);
buf BUF1 (N5120, N5110);
nand NAND2 (N5121, N5108, N257);
xor XOR2 (N5122, N5115, N4455);
not NOT1 (N5123, N5098);
or OR4 (N5124, N5112, N4060, N673, N986);
or OR3 (N5125, N5121, N2584, N4014);
or OR2 (N5126, N5105, N620);
buf BUF1 (N5127, N5107);
xor XOR2 (N5128, N5127, N1020);
nor NOR4 (N5129, N5125, N3248, N1494, N1124);
or OR2 (N5130, N5128, N3759);
not NOT1 (N5131, N5129);
and AND4 (N5132, N5130, N168, N4261, N48);
or OR4 (N5133, N5124, N1643, N4091, N4749);
nand NAND2 (N5134, N5120, N87);
nor NOR2 (N5135, N5122, N3209);
xor XOR2 (N5136, N5114, N3300);
nand NAND4 (N5137, N5132, N1785, N36, N848);
xor XOR2 (N5138, N5137, N3116);
and AND3 (N5139, N5138, N1740, N918);
nand NAND2 (N5140, N5133, N3955);
xor XOR2 (N5141, N5134, N3667);
buf BUF1 (N5142, N5126);
or OR4 (N5143, N5140, N1991, N4997, N4154);
nand NAND3 (N5144, N5131, N551, N3506);
and AND4 (N5145, N5113, N4732, N1362, N2239);
not NOT1 (N5146, N5119);
buf BUF1 (N5147, N5145);
and AND2 (N5148, N5144, N3024);
xor XOR2 (N5149, N5143, N839);
nand NAND2 (N5150, N5147, N1824);
not NOT1 (N5151, N5136);
nand NAND3 (N5152, N5151, N296, N1627);
and AND2 (N5153, N5148, N3572);
nand NAND2 (N5154, N5139, N5006);
buf BUF1 (N5155, N5141);
buf BUF1 (N5156, N5135);
or OR2 (N5157, N5155, N1026);
nand NAND3 (N5158, N5146, N4433, N1099);
nor NOR2 (N5159, N5153, N3782);
and AND2 (N5160, N5150, N1926);
not NOT1 (N5161, N5152);
not NOT1 (N5162, N5154);
and AND4 (N5163, N5158, N4172, N4990, N5135);
nand NAND3 (N5164, N5149, N3526, N3318);
and AND2 (N5165, N5162, N2438);
not NOT1 (N5166, N5159);
xor XOR2 (N5167, N5163, N3284);
nand NAND3 (N5168, N5156, N4183, N1275);
nor NOR2 (N5169, N5161, N3459);
or OR4 (N5170, N5167, N3835, N4725, N3693);
and AND4 (N5171, N5142, N4418, N925, N4059);
and AND3 (N5172, N5164, N4979, N879);
or OR2 (N5173, N5166, N559);
or OR4 (N5174, N5123, N2052, N2528, N2265);
buf BUF1 (N5175, N5169);
not NOT1 (N5176, N5168);
buf BUF1 (N5177, N5174);
not NOT1 (N5178, N5177);
or OR3 (N5179, N5173, N2329, N5);
not NOT1 (N5180, N5178);
and AND2 (N5181, N5157, N4534);
xor XOR2 (N5182, N5171, N4085);
buf BUF1 (N5183, N5182);
nor NOR3 (N5184, N5180, N3879, N973);
and AND4 (N5185, N5183, N165, N2385, N1201);
xor XOR2 (N5186, N5172, N4730);
nor NOR3 (N5187, N5179, N3590, N3267);
nand NAND4 (N5188, N5160, N1979, N4201, N4006);
nand NAND4 (N5189, N5185, N2467, N862, N2618);
nand NAND4 (N5190, N5187, N5070, N4175, N4371);
xor XOR2 (N5191, N5170, N3568);
nor NOR3 (N5192, N5176, N216, N1346);
xor XOR2 (N5193, N5190, N3436);
not NOT1 (N5194, N5192);
nand NAND4 (N5195, N5165, N1763, N556, N4931);
or OR3 (N5196, N5194, N2025, N388);
or OR3 (N5197, N5188, N2645, N4613);
xor XOR2 (N5198, N5196, N1076);
or OR2 (N5199, N5198, N603);
nand NAND2 (N5200, N5199, N1781);
and AND4 (N5201, N5186, N3130, N2104, N4436);
xor XOR2 (N5202, N5191, N619);
nand NAND2 (N5203, N5201, N3130);
buf BUF1 (N5204, N5193);
nand NAND3 (N5205, N5200, N77, N680);
or OR2 (N5206, N5203, N2828);
xor XOR2 (N5207, N5204, N2594);
not NOT1 (N5208, N5197);
xor XOR2 (N5209, N5205, N413);
nand NAND2 (N5210, N5181, N3612);
or OR4 (N5211, N5210, N4567, N1042, N2223);
nor NOR3 (N5212, N5202, N1690, N148);
or OR4 (N5213, N5175, N2840, N4942, N3353);
not NOT1 (N5214, N5208);
and AND4 (N5215, N5189, N4335, N3742, N2853);
or OR3 (N5216, N5212, N2910, N3804);
nor NOR3 (N5217, N5216, N1940, N4303);
not NOT1 (N5218, N5213);
and AND4 (N5219, N5207, N1144, N445, N832);
or OR4 (N5220, N5209, N3700, N1076, N1786);
not NOT1 (N5221, N5215);
xor XOR2 (N5222, N5219, N2657);
buf BUF1 (N5223, N5221);
buf BUF1 (N5224, N5214);
xor XOR2 (N5225, N5217, N1939);
nor NOR2 (N5226, N5220, N1000);
xor XOR2 (N5227, N5222, N4891);
nand NAND4 (N5228, N5225, N312, N2982, N2952);
xor XOR2 (N5229, N5227, N1852);
not NOT1 (N5230, N5228);
and AND3 (N5231, N5223, N3060, N3338);
buf BUF1 (N5232, N5231);
buf BUF1 (N5233, N5195);
and AND2 (N5234, N5230, N3127);
xor XOR2 (N5235, N5226, N207);
nand NAND3 (N5236, N5234, N749, N1482);
xor XOR2 (N5237, N5235, N4972);
and AND2 (N5238, N5218, N2371);
or OR2 (N5239, N5206, N4058);
or OR2 (N5240, N5224, N705);
not NOT1 (N5241, N5236);
not NOT1 (N5242, N5240);
nand NAND3 (N5243, N5232, N1396, N3712);
nand NAND2 (N5244, N5184, N2068);
not NOT1 (N5245, N5233);
xor XOR2 (N5246, N5244, N2836);
or OR3 (N5247, N5243, N1427, N159);
buf BUF1 (N5248, N5239);
xor XOR2 (N5249, N5211, N166);
nand NAND3 (N5250, N5242, N4764, N4308);
nor NOR4 (N5251, N5237, N3118, N536, N2714);
nand NAND2 (N5252, N5250, N2577);
and AND4 (N5253, N5249, N2797, N2536, N61);
buf BUF1 (N5254, N5253);
or OR2 (N5255, N5247, N4023);
nand NAND4 (N5256, N5245, N1596, N1011, N3356);
nand NAND4 (N5257, N5251, N4526, N4169, N2496);
xor XOR2 (N5258, N5256, N1630);
nand NAND4 (N5259, N5229, N1498, N4842, N5068);
or OR3 (N5260, N5254, N1146, N2911);
nor NOR3 (N5261, N5252, N809, N3051);
not NOT1 (N5262, N5258);
nand NAND2 (N5263, N5257, N2481);
nor NOR4 (N5264, N5263, N4302, N3958, N4909);
buf BUF1 (N5265, N5248);
buf BUF1 (N5266, N5262);
nor NOR4 (N5267, N5246, N4590, N4830, N886);
xor XOR2 (N5268, N5266, N5238);
and AND4 (N5269, N2105, N629, N3524, N3178);
buf BUF1 (N5270, N5267);
or OR2 (N5271, N5260, N642);
nand NAND4 (N5272, N5255, N3711, N2372, N5009);
and AND3 (N5273, N5272, N380, N4988);
buf BUF1 (N5274, N5241);
nand NAND3 (N5275, N5268, N4530, N1100);
or OR3 (N5276, N5265, N4899, N2945);
nand NAND3 (N5277, N5261, N4301, N1500);
nor NOR2 (N5278, N5276, N1186);
xor XOR2 (N5279, N5275, N1171);
not NOT1 (N5280, N5271);
xor XOR2 (N5281, N5259, N2662);
or OR3 (N5282, N5281, N1775, N177);
xor XOR2 (N5283, N5280, N2921);
or OR2 (N5284, N5282, N4725);
or OR4 (N5285, N5278, N2603, N4050, N889);
and AND2 (N5286, N5284, N4065);
nand NAND4 (N5287, N5264, N481, N4820, N459);
buf BUF1 (N5288, N5286);
nor NOR2 (N5289, N5277, N538);
nand NAND4 (N5290, N5288, N2895, N578, N5123);
not NOT1 (N5291, N5270);
xor XOR2 (N5292, N5290, N3223);
and AND2 (N5293, N5279, N2357);
nand NAND2 (N5294, N5269, N4580);
or OR4 (N5295, N5293, N864, N2926, N917);
or OR2 (N5296, N5287, N2706);
or OR3 (N5297, N5291, N5002, N4122);
and AND3 (N5298, N5285, N5211, N1728);
and AND2 (N5299, N5289, N2818);
and AND4 (N5300, N5298, N3707, N3713, N2891);
xor XOR2 (N5301, N5300, N4222);
xor XOR2 (N5302, N5295, N1176);
and AND4 (N5303, N5273, N1461, N2173, N3866);
buf BUF1 (N5304, N5303);
not NOT1 (N5305, N5304);
or OR2 (N5306, N5274, N3371);
and AND2 (N5307, N5296, N1615);
or OR2 (N5308, N5302, N2967);
nand NAND3 (N5309, N5305, N2652, N349);
nor NOR2 (N5310, N5309, N3707);
or OR3 (N5311, N5308, N2662, N4196);
not NOT1 (N5312, N5307);
not NOT1 (N5313, N5311);
buf BUF1 (N5314, N5283);
nand NAND3 (N5315, N5294, N795, N2113);
nor NOR2 (N5316, N5297, N3309);
or OR3 (N5317, N5313, N1538, N5129);
nand NAND2 (N5318, N5315, N1778);
and AND3 (N5319, N5301, N3481, N1358);
nor NOR3 (N5320, N5316, N4430, N1606);
not NOT1 (N5321, N5310);
buf BUF1 (N5322, N5317);
xor XOR2 (N5323, N5312, N2824);
xor XOR2 (N5324, N5318, N3266);
nor NOR4 (N5325, N5321, N4631, N4929, N284);
or OR3 (N5326, N5322, N4697, N339);
or OR3 (N5327, N5326, N3102, N2960);
nand NAND4 (N5328, N5320, N636, N1575, N5003);
xor XOR2 (N5329, N5324, N947);
buf BUF1 (N5330, N5327);
or OR4 (N5331, N5314, N3259, N1408, N2966);
buf BUF1 (N5332, N5319);
and AND4 (N5333, N5292, N2362, N3571, N3075);
xor XOR2 (N5334, N5328, N5089);
and AND2 (N5335, N5325, N657);
nand NAND4 (N5336, N5299, N860, N1176, N341);
or OR4 (N5337, N5323, N760, N5094, N2160);
or OR3 (N5338, N5333, N3103, N3465);
and AND2 (N5339, N5332, N4233);
and AND3 (N5340, N5306, N4158, N129);
xor XOR2 (N5341, N5336, N4266);
and AND4 (N5342, N5337, N2596, N329, N3035);
not NOT1 (N5343, N5338);
not NOT1 (N5344, N5340);
nand NAND3 (N5345, N5329, N1427, N3596);
or OR4 (N5346, N5330, N1970, N1764, N1639);
xor XOR2 (N5347, N5341, N449);
and AND2 (N5348, N5346, N4651);
buf BUF1 (N5349, N5342);
nand NAND4 (N5350, N5334, N3599, N1945, N4659);
nand NAND3 (N5351, N5350, N2875, N3025);
xor XOR2 (N5352, N5351, N3586);
nor NOR2 (N5353, N5345, N4913);
nand NAND2 (N5354, N5343, N4739);
and AND2 (N5355, N5335, N3350);
xor XOR2 (N5356, N5355, N4919);
or OR3 (N5357, N5339, N4209, N2731);
nand NAND4 (N5358, N5356, N1692, N2914, N4582);
buf BUF1 (N5359, N5357);
xor XOR2 (N5360, N5359, N1176);
or OR4 (N5361, N5344, N4377, N526, N3969);
or OR3 (N5362, N5348, N4306, N4478);
nand NAND2 (N5363, N5354, N317);
or OR2 (N5364, N5331, N3056);
or OR2 (N5365, N5362, N349);
not NOT1 (N5366, N5365);
xor XOR2 (N5367, N5364, N3427);
nand NAND4 (N5368, N5367, N4987, N650, N4926);
not NOT1 (N5369, N5366);
not NOT1 (N5370, N5363);
xor XOR2 (N5371, N5370, N1559);
not NOT1 (N5372, N5368);
xor XOR2 (N5373, N5372, N3114);
or OR2 (N5374, N5360, N2479);
nand NAND3 (N5375, N5353, N2564, N3854);
nand NAND2 (N5376, N5373, N1056);
xor XOR2 (N5377, N5358, N3415);
nor NOR3 (N5378, N5374, N1294, N4215);
nor NOR4 (N5379, N5377, N1652, N824, N1602);
nor NOR4 (N5380, N5352, N1062, N4708, N2172);
buf BUF1 (N5381, N5380);
xor XOR2 (N5382, N5381, N1916);
buf BUF1 (N5383, N5378);
not NOT1 (N5384, N5375);
or OR2 (N5385, N5349, N1474);
buf BUF1 (N5386, N5382);
xor XOR2 (N5387, N5376, N4626);
and AND3 (N5388, N5383, N5202, N4683);
not NOT1 (N5389, N5371);
buf BUF1 (N5390, N5361);
and AND2 (N5391, N5379, N5026);
nor NOR4 (N5392, N5386, N835, N1883, N5348);
xor XOR2 (N5393, N5347, N949);
or OR2 (N5394, N5369, N2235);
nand NAND3 (N5395, N5385, N134, N2731);
not NOT1 (N5396, N5387);
not NOT1 (N5397, N5391);
xor XOR2 (N5398, N5384, N657);
and AND2 (N5399, N5392, N4125);
not NOT1 (N5400, N5390);
and AND2 (N5401, N5399, N3405);
xor XOR2 (N5402, N5394, N3209);
buf BUF1 (N5403, N5393);
nor NOR4 (N5404, N5401, N2700, N389, N1960);
buf BUF1 (N5405, N5388);
xor XOR2 (N5406, N5397, N1159);
not NOT1 (N5407, N5403);
buf BUF1 (N5408, N5400);
buf BUF1 (N5409, N5405);
nor NOR4 (N5410, N5408, N5312, N2964, N3488);
and AND2 (N5411, N5404, N4727);
nor NOR3 (N5412, N5395, N976, N3702);
nor NOR4 (N5413, N5411, N3891, N5203, N584);
or OR3 (N5414, N5398, N2027, N2406);
and AND3 (N5415, N5396, N4294, N4683);
and AND3 (N5416, N5412, N2793, N979);
not NOT1 (N5417, N5416);
buf BUF1 (N5418, N5413);
xor XOR2 (N5419, N5415, N2510);
not NOT1 (N5420, N5409);
nand NAND3 (N5421, N5410, N5034, N1457);
and AND2 (N5422, N5420, N5252);
and AND3 (N5423, N5406, N2047, N3304);
and AND3 (N5424, N5414, N4963, N3);
not NOT1 (N5425, N5419);
buf BUF1 (N5426, N5425);
not NOT1 (N5427, N5407);
buf BUF1 (N5428, N5422);
and AND2 (N5429, N5427, N1056);
or OR2 (N5430, N5421, N1579);
nor NOR2 (N5431, N5389, N1479);
xor XOR2 (N5432, N5429, N801);
not NOT1 (N5433, N5418);
buf BUF1 (N5434, N5428);
not NOT1 (N5435, N5426);
nor NOR4 (N5436, N5424, N2497, N603, N3884);
and AND4 (N5437, N5431, N4939, N1202, N4540);
or OR2 (N5438, N5434, N4632);
xor XOR2 (N5439, N5423, N2908);
not NOT1 (N5440, N5436);
nand NAND2 (N5441, N5439, N1947);
or OR4 (N5442, N5432, N235, N1514, N2430);
or OR3 (N5443, N5435, N1295, N2433);
not NOT1 (N5444, N5402);
buf BUF1 (N5445, N5442);
and AND3 (N5446, N5417, N1139, N2421);
and AND4 (N5447, N5437, N2678, N2193, N638);
not NOT1 (N5448, N5438);
or OR4 (N5449, N5445, N4269, N1359, N287);
not NOT1 (N5450, N5449);
not NOT1 (N5451, N5433);
not NOT1 (N5452, N5448);
not NOT1 (N5453, N5452);
xor XOR2 (N5454, N5443, N2200);
nor NOR4 (N5455, N5446, N4647, N3884, N247);
or OR2 (N5456, N5453, N503);
nor NOR4 (N5457, N5451, N2365, N4217, N1367);
not NOT1 (N5458, N5454);
xor XOR2 (N5459, N5450, N645);
not NOT1 (N5460, N5455);
nor NOR2 (N5461, N5457, N3562);
not NOT1 (N5462, N5458);
xor XOR2 (N5463, N5441, N481);
buf BUF1 (N5464, N5447);
not NOT1 (N5465, N5461);
nand NAND3 (N5466, N5460, N2501, N5069);
and AND4 (N5467, N5430, N3566, N4496, N3916);
buf BUF1 (N5468, N5463);
not NOT1 (N5469, N5462);
or OR4 (N5470, N5464, N3469, N1340, N1027);
nor NOR3 (N5471, N5456, N5166, N1269);
buf BUF1 (N5472, N5465);
not NOT1 (N5473, N5444);
nand NAND2 (N5474, N5440, N4005);
not NOT1 (N5475, N5459);
not NOT1 (N5476, N5473);
nor NOR3 (N5477, N5467, N3692, N5421);
buf BUF1 (N5478, N5469);
nand NAND3 (N5479, N5470, N2664, N1634);
or OR2 (N5480, N5477, N4743);
nor NOR4 (N5481, N5479, N1848, N2208, N1616);
not NOT1 (N5482, N5481);
and AND3 (N5483, N5482, N5187, N982);
and AND2 (N5484, N5476, N2137);
nand NAND4 (N5485, N5472, N862, N3616, N3078);
nand NAND2 (N5486, N5480, N2008);
or OR3 (N5487, N5483, N4781, N4223);
and AND4 (N5488, N5485, N501, N3984, N1408);
and AND2 (N5489, N5486, N2367);
buf BUF1 (N5490, N5471);
xor XOR2 (N5491, N5475, N3536);
xor XOR2 (N5492, N5484, N1014);
nor NOR4 (N5493, N5466, N118, N3325, N2628);
buf BUF1 (N5494, N5487);
nand NAND2 (N5495, N5494, N3112);
nor NOR4 (N5496, N5495, N1993, N130, N2816);
xor XOR2 (N5497, N5478, N3422);
nor NOR4 (N5498, N5496, N4461, N245, N373);
and AND3 (N5499, N5492, N1416, N58);
and AND3 (N5500, N5489, N5114, N214);
and AND4 (N5501, N5498, N45, N793, N1202);
and AND3 (N5502, N5497, N2176, N84);
buf BUF1 (N5503, N5493);
and AND2 (N5504, N5501, N3189);
buf BUF1 (N5505, N5504);
xor XOR2 (N5506, N5491, N2545);
or OR2 (N5507, N5488, N622);
or OR3 (N5508, N5490, N3330, N1937);
xor XOR2 (N5509, N5505, N5172);
xor XOR2 (N5510, N5468, N1641);
or OR3 (N5511, N5500, N749, N198);
nor NOR2 (N5512, N5474, N3903);
nand NAND3 (N5513, N5499, N3269, N4409);
nand NAND2 (N5514, N5512, N1532);
buf BUF1 (N5515, N5508);
not NOT1 (N5516, N5506);
nor NOR4 (N5517, N5507, N5459, N148, N902);
not NOT1 (N5518, N5509);
not NOT1 (N5519, N5516);
buf BUF1 (N5520, N5510);
nor NOR3 (N5521, N5514, N1273, N689);
nand NAND3 (N5522, N5521, N2965, N4828);
nor NOR3 (N5523, N5518, N5108, N2961);
not NOT1 (N5524, N5503);
nor NOR3 (N5525, N5520, N3756, N1127);
and AND3 (N5526, N5524, N3495, N2715);
xor XOR2 (N5527, N5525, N4567);
and AND4 (N5528, N5515, N613, N3068, N720);
xor XOR2 (N5529, N5517, N4011);
xor XOR2 (N5530, N5502, N5290);
nand NAND2 (N5531, N5530, N4839);
and AND2 (N5532, N5526, N5010);
and AND4 (N5533, N5519, N3915, N1305, N4323);
nor NOR3 (N5534, N5532, N4843, N4090);
or OR4 (N5535, N5528, N3598, N4138, N5220);
xor XOR2 (N5536, N5513, N3910);
nand NAND4 (N5537, N5523, N971, N2667, N574);
and AND2 (N5538, N5535, N5010);
nor NOR4 (N5539, N5533, N3003, N3351, N3910);
or OR2 (N5540, N5527, N4360);
not NOT1 (N5541, N5537);
not NOT1 (N5542, N5529);
buf BUF1 (N5543, N5538);
nand NAND4 (N5544, N5534, N126, N3877, N1691);
or OR2 (N5545, N5540, N5212);
not NOT1 (N5546, N5544);
not NOT1 (N5547, N5543);
nor NOR3 (N5548, N5511, N3770, N587);
nor NOR2 (N5549, N5531, N5183);
not NOT1 (N5550, N5546);
nor NOR4 (N5551, N5522, N965, N3464, N2216);
xor XOR2 (N5552, N5551, N1359);
xor XOR2 (N5553, N5541, N4076);
xor XOR2 (N5554, N5553, N768);
xor XOR2 (N5555, N5536, N1444);
nor NOR2 (N5556, N5550, N3642);
nand NAND3 (N5557, N5556, N3873, N2980);
nand NAND3 (N5558, N5547, N4410, N8);
xor XOR2 (N5559, N5554, N3433);
not NOT1 (N5560, N5539);
and AND4 (N5561, N5555, N4151, N5224, N3912);
nor NOR2 (N5562, N5549, N1821);
nand NAND3 (N5563, N5552, N2735, N806);
not NOT1 (N5564, N5558);
not NOT1 (N5565, N5561);
and AND4 (N5566, N5542, N3549, N3659, N4171);
and AND3 (N5567, N5565, N929, N2747);
or OR4 (N5568, N5567, N2201, N4415, N5097);
nand NAND2 (N5569, N5548, N4255);
and AND4 (N5570, N5545, N3488, N1038, N2884);
and AND4 (N5571, N5557, N1918, N2133, N865);
nand NAND2 (N5572, N5563, N1308);
and AND3 (N5573, N5570, N5239, N5200);
xor XOR2 (N5574, N5562, N3698);
not NOT1 (N5575, N5566);
buf BUF1 (N5576, N5559);
buf BUF1 (N5577, N5576);
buf BUF1 (N5578, N5571);
xor XOR2 (N5579, N5569, N62);
buf BUF1 (N5580, N5560);
not NOT1 (N5581, N5575);
buf BUF1 (N5582, N5564);
xor XOR2 (N5583, N5573, N3998);
not NOT1 (N5584, N5568);
buf BUF1 (N5585, N5580);
xor XOR2 (N5586, N5578, N3591);
nor NOR2 (N5587, N5584, N5239);
nor NOR3 (N5588, N5583, N1522, N3931);
or OR2 (N5589, N5574, N4396);
or OR3 (N5590, N5585, N202, N3017);
nor NOR3 (N5591, N5590, N2809, N3470);
and AND3 (N5592, N5581, N1537, N4496);
and AND2 (N5593, N5577, N5002);
buf BUF1 (N5594, N5591);
buf BUF1 (N5595, N5579);
and AND4 (N5596, N5588, N4073, N1758, N1678);
not NOT1 (N5597, N5582);
nor NOR3 (N5598, N5589, N2000, N3179);
nand NAND4 (N5599, N5598, N4602, N3799, N3456);
nor NOR4 (N5600, N5599, N639, N1968, N1970);
buf BUF1 (N5601, N5592);
and AND3 (N5602, N5601, N4000, N3246);
buf BUF1 (N5603, N5600);
nand NAND3 (N5604, N5597, N356, N1969);
not NOT1 (N5605, N5603);
not NOT1 (N5606, N5605);
not NOT1 (N5607, N5596);
buf BUF1 (N5608, N5572);
buf BUF1 (N5609, N5594);
not NOT1 (N5610, N5602);
nor NOR4 (N5611, N5606, N2869, N1893, N5545);
and AND4 (N5612, N5593, N4434, N3675, N1259);
nand NAND4 (N5613, N5612, N2159, N710, N2636);
or OR2 (N5614, N5607, N3058);
buf BUF1 (N5615, N5614);
or OR2 (N5616, N5604, N3590);
and AND2 (N5617, N5609, N2847);
nor NOR3 (N5618, N5610, N1283, N334);
buf BUF1 (N5619, N5611);
nor NOR4 (N5620, N5617, N2301, N79, N4818);
or OR3 (N5621, N5613, N450, N805);
buf BUF1 (N5622, N5615);
buf BUF1 (N5623, N5618);
not NOT1 (N5624, N5587);
nor NOR2 (N5625, N5620, N5422);
nor NOR2 (N5626, N5625, N4650);
nor NOR2 (N5627, N5616, N945);
or OR3 (N5628, N5627, N3617, N843);
nand NAND2 (N5629, N5623, N1070);
not NOT1 (N5630, N5628);
nor NOR3 (N5631, N5586, N4597, N3927);
nand NAND4 (N5632, N5608, N4180, N2115, N574);
nand NAND4 (N5633, N5595, N4720, N2023, N4359);
not NOT1 (N5634, N5631);
or OR2 (N5635, N5621, N164);
nand NAND3 (N5636, N5630, N5229, N2522);
not NOT1 (N5637, N5636);
not NOT1 (N5638, N5633);
not NOT1 (N5639, N5632);
and AND2 (N5640, N5624, N1059);
nor NOR3 (N5641, N5640, N260, N929);
nand NAND4 (N5642, N5626, N5038, N2605, N2557);
xor XOR2 (N5643, N5637, N4064);
not NOT1 (N5644, N5622);
not NOT1 (N5645, N5635);
nand NAND3 (N5646, N5645, N2633, N1914);
and AND4 (N5647, N5639, N3430, N2207, N766);
buf BUF1 (N5648, N5619);
nand NAND3 (N5649, N5643, N4815, N1562);
not NOT1 (N5650, N5646);
xor XOR2 (N5651, N5634, N3042);
or OR3 (N5652, N5638, N473, N1028);
and AND4 (N5653, N5648, N4267, N1241, N21);
or OR3 (N5654, N5652, N3457, N1633);
nand NAND4 (N5655, N5651, N3184, N3375, N5564);
nand NAND4 (N5656, N5653, N1059, N4322, N2184);
nand NAND2 (N5657, N5650, N1222);
xor XOR2 (N5658, N5629, N5070);
or OR2 (N5659, N5641, N1425);
buf BUF1 (N5660, N5658);
or OR2 (N5661, N5660, N2626);
not NOT1 (N5662, N5644);
not NOT1 (N5663, N5662);
not NOT1 (N5664, N5663);
buf BUF1 (N5665, N5659);
or OR2 (N5666, N5654, N2663);
xor XOR2 (N5667, N5661, N3379);
nor NOR2 (N5668, N5665, N5647);
not NOT1 (N5669, N530);
and AND4 (N5670, N5655, N382, N5025, N2839);
nand NAND2 (N5671, N5649, N4088);
or OR2 (N5672, N5642, N4317);
xor XOR2 (N5673, N5664, N1633);
xor XOR2 (N5674, N5667, N1660);
xor XOR2 (N5675, N5673, N895);
nor NOR2 (N5676, N5672, N3530);
xor XOR2 (N5677, N5676, N4842);
xor XOR2 (N5678, N5656, N1216);
or OR3 (N5679, N5677, N3669, N2226);
xor XOR2 (N5680, N5679, N3957);
and AND4 (N5681, N5657, N2133, N2446, N4391);
nand NAND4 (N5682, N5681, N154, N2902, N3823);
nor NOR3 (N5683, N5669, N171, N1483);
and AND2 (N5684, N5675, N2692);
xor XOR2 (N5685, N5684, N3276);
xor XOR2 (N5686, N5668, N1449);
buf BUF1 (N5687, N5671);
and AND2 (N5688, N5670, N2811);
xor XOR2 (N5689, N5678, N175);
buf BUF1 (N5690, N5674);
and AND2 (N5691, N5687, N1783);
xor XOR2 (N5692, N5689, N284);
not NOT1 (N5693, N5688);
nor NOR4 (N5694, N5683, N3218, N1698, N1928);
buf BUF1 (N5695, N5666);
not NOT1 (N5696, N5680);
or OR3 (N5697, N5692, N1378, N3761);
xor XOR2 (N5698, N5696, N4340);
nor NOR3 (N5699, N5698, N163, N3530);
buf BUF1 (N5700, N5695);
or OR3 (N5701, N5694, N5149, N1907);
xor XOR2 (N5702, N5701, N1617);
or OR4 (N5703, N5699, N2537, N528, N2649);
not NOT1 (N5704, N5700);
nand NAND2 (N5705, N5693, N2781);
nor NOR2 (N5706, N5704, N5452);
nand NAND3 (N5707, N5686, N5385, N2662);
buf BUF1 (N5708, N5707);
buf BUF1 (N5709, N5706);
not NOT1 (N5710, N5682);
buf BUF1 (N5711, N5708);
nor NOR4 (N5712, N5691, N5306, N1333, N5552);
not NOT1 (N5713, N5685);
xor XOR2 (N5714, N5709, N2966);
xor XOR2 (N5715, N5710, N5285);
nor NOR4 (N5716, N5712, N666, N33, N2116);
nand NAND3 (N5717, N5702, N2468, N5690);
and AND3 (N5718, N2246, N2897, N2701);
not NOT1 (N5719, N5717);
and AND3 (N5720, N5711, N3089, N2388);
nor NOR2 (N5721, N5720, N3714);
nand NAND2 (N5722, N5703, N1144);
or OR3 (N5723, N5716, N1541, N480);
nand NAND2 (N5724, N5723, N2688);
or OR3 (N5725, N5722, N2257, N3282);
and AND4 (N5726, N5715, N2520, N249, N5000);
xor XOR2 (N5727, N5719, N3624);
and AND3 (N5728, N5705, N4189, N4271);
nand NAND4 (N5729, N5713, N4964, N5028, N394);
buf BUF1 (N5730, N5721);
not NOT1 (N5731, N5729);
nand NAND3 (N5732, N5724, N431, N2463);
and AND2 (N5733, N5697, N3416);
not NOT1 (N5734, N5733);
nand NAND2 (N5735, N5734, N4965);
buf BUF1 (N5736, N5714);
or OR2 (N5737, N5726, N4901);
or OR3 (N5738, N5731, N4367, N2344);
nor NOR2 (N5739, N5737, N3282);
not NOT1 (N5740, N5725);
nand NAND2 (N5741, N5727, N1844);
buf BUF1 (N5742, N5718);
xor XOR2 (N5743, N5736, N5527);
and AND3 (N5744, N5741, N2702, N94);
and AND3 (N5745, N5744, N3933, N3050);
not NOT1 (N5746, N5739);
or OR3 (N5747, N5745, N2733, N4152);
and AND4 (N5748, N5730, N1964, N120, N2752);
xor XOR2 (N5749, N5742, N485);
buf BUF1 (N5750, N5732);
or OR3 (N5751, N5746, N590, N298);
and AND3 (N5752, N5748, N5069, N4999);
xor XOR2 (N5753, N5751, N955);
xor XOR2 (N5754, N5743, N2263);
and AND2 (N5755, N5752, N2993);
nand NAND2 (N5756, N5738, N3190);
and AND4 (N5757, N5756, N786, N4317, N4876);
nand NAND3 (N5758, N5757, N4113, N512);
nor NOR2 (N5759, N5740, N5758);
not NOT1 (N5760, N863);
not NOT1 (N5761, N5755);
nor NOR4 (N5762, N5759, N1838, N4286, N3038);
not NOT1 (N5763, N5728);
buf BUF1 (N5764, N5754);
xor XOR2 (N5765, N5764, N5505);
and AND2 (N5766, N5749, N1075);
nor NOR4 (N5767, N5750, N2406, N3995, N1374);
nand NAND3 (N5768, N5767, N949, N1129);
and AND4 (N5769, N5761, N460, N3848, N4149);
nand NAND4 (N5770, N5763, N1930, N3723, N1455);
nor NOR3 (N5771, N5762, N4968, N2067);
nand NAND2 (N5772, N5753, N5547);
nor NOR3 (N5773, N5768, N1903, N5141);
not NOT1 (N5774, N5773);
and AND2 (N5775, N5760, N2659);
and AND4 (N5776, N5772, N4304, N1552, N5151);
or OR3 (N5777, N5770, N2547, N2331);
xor XOR2 (N5778, N5771, N1760);
xor XOR2 (N5779, N5766, N3973);
buf BUF1 (N5780, N5735);
nand NAND4 (N5781, N5780, N5265, N1705, N1284);
not NOT1 (N5782, N5769);
buf BUF1 (N5783, N5775);
nand NAND4 (N5784, N5765, N4072, N750, N2985);
nand NAND4 (N5785, N5747, N1883, N1682, N5282);
xor XOR2 (N5786, N5779, N84);
buf BUF1 (N5787, N5777);
nand NAND4 (N5788, N5782, N3066, N2908, N2235);
nand NAND3 (N5789, N5781, N1218, N3203);
and AND2 (N5790, N5788, N1518);
not NOT1 (N5791, N5774);
xor XOR2 (N5792, N5785, N5029);
or OR2 (N5793, N5790, N4557);
buf BUF1 (N5794, N5784);
and AND2 (N5795, N5793, N993);
buf BUF1 (N5796, N5794);
xor XOR2 (N5797, N5796, N1322);
nand NAND3 (N5798, N5783, N3042, N5649);
not NOT1 (N5799, N5787);
and AND4 (N5800, N5792, N4272, N2958, N1045);
nand NAND3 (N5801, N5800, N3519, N5716);
not NOT1 (N5802, N5786);
nand NAND2 (N5803, N5776, N2495);
nand NAND4 (N5804, N5803, N3363, N4361, N1311);
not NOT1 (N5805, N5789);
or OR4 (N5806, N5802, N1234, N39, N4045);
buf BUF1 (N5807, N5778);
xor XOR2 (N5808, N5806, N3188);
nand NAND2 (N5809, N5799, N2407);
nand NAND2 (N5810, N5809, N4780);
nor NOR2 (N5811, N5804, N3221);
xor XOR2 (N5812, N5808, N5144);
not NOT1 (N5813, N5791);
nand NAND4 (N5814, N5813, N1948, N1968, N1508);
and AND4 (N5815, N5811, N4615, N4456, N2234);
xor XOR2 (N5816, N5801, N613);
or OR4 (N5817, N5805, N3743, N1649, N3366);
nand NAND4 (N5818, N5797, N2576, N4537, N3387);
not NOT1 (N5819, N5810);
not NOT1 (N5820, N5815);
nand NAND2 (N5821, N5819, N168);
xor XOR2 (N5822, N5814, N1043);
xor XOR2 (N5823, N5818, N3858);
or OR3 (N5824, N5823, N1096, N837);
not NOT1 (N5825, N5795);
buf BUF1 (N5826, N5807);
buf BUF1 (N5827, N5821);
buf BUF1 (N5828, N5816);
not NOT1 (N5829, N5822);
nand NAND4 (N5830, N5817, N699, N5811, N1969);
xor XOR2 (N5831, N5824, N555);
or OR3 (N5832, N5831, N4614, N3885);
and AND2 (N5833, N5828, N1897);
nand NAND3 (N5834, N5833, N4422, N3152);
and AND3 (N5835, N5829, N2398, N5050);
nand NAND4 (N5836, N5820, N4152, N4740, N4706);
buf BUF1 (N5837, N5834);
buf BUF1 (N5838, N5812);
nor NOR4 (N5839, N5827, N1761, N791, N635);
not NOT1 (N5840, N5835);
not NOT1 (N5841, N5839);
or OR4 (N5842, N5832, N5011, N957, N5018);
buf BUF1 (N5843, N5840);
not NOT1 (N5844, N5841);
or OR2 (N5845, N5825, N682);
nand NAND2 (N5846, N5845, N1519);
or OR4 (N5847, N5836, N1177, N4799, N4376);
not NOT1 (N5848, N5830);
nor NOR2 (N5849, N5847, N4150);
nor NOR3 (N5850, N5844, N322, N306);
nand NAND3 (N5851, N5849, N809, N2777);
and AND4 (N5852, N5851, N3460, N107, N2293);
nand NAND3 (N5853, N5852, N480, N2726);
or OR2 (N5854, N5798, N412);
or OR3 (N5855, N5848, N1870, N2610);
and AND4 (N5856, N5837, N3701, N233, N4612);
nand NAND4 (N5857, N5846, N3225, N4712, N5362);
nor NOR4 (N5858, N5857, N2271, N3708, N119);
not NOT1 (N5859, N5850);
nand NAND4 (N5860, N5842, N3699, N349, N3864);
not NOT1 (N5861, N5853);
not NOT1 (N5862, N5859);
buf BUF1 (N5863, N5854);
and AND2 (N5864, N5862, N5391);
nand NAND3 (N5865, N5863, N5492, N2788);
and AND3 (N5866, N5864, N307, N114);
or OR4 (N5867, N5856, N1137, N3703, N2881);
and AND4 (N5868, N5838, N5622, N2899, N3783);
buf BUF1 (N5869, N5867);
or OR2 (N5870, N5858, N1786);
buf BUF1 (N5871, N5860);
not NOT1 (N5872, N5869);
and AND2 (N5873, N5868, N4021);
and AND4 (N5874, N5865, N5172, N1074, N3476);
or OR2 (N5875, N5872, N3550);
nand NAND3 (N5876, N5866, N2028, N4454);
nand NAND2 (N5877, N5876, N3933);
buf BUF1 (N5878, N5861);
and AND2 (N5879, N5870, N1126);
nand NAND2 (N5880, N5855, N4476);
nor NOR4 (N5881, N5871, N5550, N829, N1243);
and AND2 (N5882, N5843, N944);
or OR3 (N5883, N5878, N5248, N2841);
not NOT1 (N5884, N5873);
nand NAND2 (N5885, N5884, N5716);
and AND3 (N5886, N5880, N1499, N4412);
nor NOR3 (N5887, N5826, N3903, N2145);
and AND2 (N5888, N5879, N4748);
nand NAND3 (N5889, N5882, N3026, N5500);
not NOT1 (N5890, N5883);
not NOT1 (N5891, N5888);
buf BUF1 (N5892, N5889);
and AND2 (N5893, N5881, N1283);
nand NAND4 (N5894, N5890, N862, N1042, N2100);
or OR2 (N5895, N5885, N205);
nor NOR3 (N5896, N5894, N5872, N1757);
buf BUF1 (N5897, N5887);
not NOT1 (N5898, N5897);
or OR2 (N5899, N5886, N4477);
xor XOR2 (N5900, N5898, N5170);
nand NAND4 (N5901, N5874, N255, N445, N1673);
or OR2 (N5902, N5895, N5515);
or OR3 (N5903, N5901, N1468, N4951);
not NOT1 (N5904, N5900);
nand NAND4 (N5905, N5902, N5067, N826, N611);
nand NAND2 (N5906, N5892, N4984);
or OR2 (N5907, N5905, N505);
not NOT1 (N5908, N5904);
nor NOR4 (N5909, N5908, N4930, N4081, N2099);
nand NAND3 (N5910, N5906, N2455, N4901);
nor NOR4 (N5911, N5909, N1223, N3873, N4752);
and AND4 (N5912, N5877, N5755, N2640, N5693);
nor NOR2 (N5913, N5907, N1815);
xor XOR2 (N5914, N5899, N1925);
buf BUF1 (N5915, N5903);
and AND3 (N5916, N5910, N2609, N3823);
nor NOR4 (N5917, N5915, N1422, N3526, N2998);
nor NOR2 (N5918, N5917, N4611);
buf BUF1 (N5919, N5896);
or OR4 (N5920, N5875, N4732, N3626, N1589);
not NOT1 (N5921, N5911);
and AND4 (N5922, N5921, N1578, N4216, N905);
and AND2 (N5923, N5916, N5601);
or OR4 (N5924, N5912, N447, N2397, N2537);
or OR4 (N5925, N5924, N516, N394, N2728);
nand NAND4 (N5926, N5891, N2932, N1436, N3048);
nor NOR3 (N5927, N5920, N2282, N1133);
not NOT1 (N5928, N5927);
not NOT1 (N5929, N5928);
buf BUF1 (N5930, N5918);
not NOT1 (N5931, N5914);
not NOT1 (N5932, N5930);
xor XOR2 (N5933, N5922, N4864);
or OR3 (N5934, N5923, N496, N4434);
xor XOR2 (N5935, N5931, N3314);
and AND3 (N5936, N5919, N5846, N5401);
buf BUF1 (N5937, N5913);
not NOT1 (N5938, N5933);
not NOT1 (N5939, N5926);
and AND4 (N5940, N5934, N3333, N4326, N959);
nor NOR4 (N5941, N5925, N1745, N4380, N5282);
buf BUF1 (N5942, N5932);
nor NOR4 (N5943, N5937, N1120, N5753, N1991);
xor XOR2 (N5944, N5936, N1603);
nor NOR4 (N5945, N5938, N3411, N3048, N508);
buf BUF1 (N5946, N5944);
not NOT1 (N5947, N5935);
not NOT1 (N5948, N5939);
xor XOR2 (N5949, N5946, N5195);
buf BUF1 (N5950, N5929);
and AND2 (N5951, N5943, N1965);
not NOT1 (N5952, N5942);
or OR2 (N5953, N5948, N1242);
and AND2 (N5954, N5953, N286);
buf BUF1 (N5955, N5950);
nor NOR2 (N5956, N5955, N1806);
or OR3 (N5957, N5956, N1221, N2470);
nand NAND3 (N5958, N5949, N5722, N2883);
xor XOR2 (N5959, N5957, N474);
not NOT1 (N5960, N5947);
nand NAND4 (N5961, N5951, N603, N4071, N4600);
and AND3 (N5962, N5941, N2657, N5661);
nor NOR2 (N5963, N5893, N2565);
or OR3 (N5964, N5960, N5963, N5256);
nor NOR2 (N5965, N2410, N2083);
and AND2 (N5966, N5965, N501);
nor NOR4 (N5967, N5945, N3846, N25, N88);
buf BUF1 (N5968, N5952);
and AND2 (N5969, N5961, N5786);
xor XOR2 (N5970, N5969, N783);
xor XOR2 (N5971, N5959, N4653);
or OR4 (N5972, N5970, N4541, N1731, N4330);
xor XOR2 (N5973, N5958, N1440);
xor XOR2 (N5974, N5972, N2242);
not NOT1 (N5975, N5967);
buf BUF1 (N5976, N5954);
not NOT1 (N5977, N5976);
nor NOR4 (N5978, N5974, N5819, N5595, N2772);
and AND2 (N5979, N5940, N2680);
not NOT1 (N5980, N5978);
not NOT1 (N5981, N5964);
not NOT1 (N5982, N5962);
nor NOR2 (N5983, N5973, N3461);
nor NOR2 (N5984, N5980, N1396);
or OR3 (N5985, N5984, N3164, N279);
nand NAND3 (N5986, N5985, N5518, N358);
nand NAND3 (N5987, N5982, N109, N5075);
not NOT1 (N5988, N5966);
not NOT1 (N5989, N5988);
not NOT1 (N5990, N5979);
buf BUF1 (N5991, N5987);
buf BUF1 (N5992, N5989);
buf BUF1 (N5993, N5983);
nor NOR3 (N5994, N5993, N4952, N4320);
xor XOR2 (N5995, N5981, N1093);
and AND2 (N5996, N5994, N2023);
xor XOR2 (N5997, N5977, N1777);
nor NOR4 (N5998, N5986, N3212, N1209, N925);
nor NOR3 (N5999, N5995, N946, N2556);
or OR3 (N6000, N5975, N2841, N5021);
buf BUF1 (N6001, N5971);
xor XOR2 (N6002, N5997, N2961);
nor NOR3 (N6003, N6002, N1501, N5722);
nand NAND4 (N6004, N6000, N3321, N2563, N5032);
nor NOR4 (N6005, N6001, N5080, N3491, N1729);
xor XOR2 (N6006, N6005, N1673);
and AND2 (N6007, N6003, N3858);
and AND3 (N6008, N5996, N3737, N2163);
nor NOR4 (N6009, N6004, N2911, N3191, N2092);
nor NOR3 (N6010, N5999, N2068, N3604);
nand NAND4 (N6011, N5990, N440, N4033, N3779);
not NOT1 (N6012, N5998);
nand NAND2 (N6013, N6012, N5260);
nor NOR2 (N6014, N6006, N3114);
buf BUF1 (N6015, N5968);
buf BUF1 (N6016, N6015);
xor XOR2 (N6017, N5991, N5955);
xor XOR2 (N6018, N6009, N1886);
nor NOR2 (N6019, N6016, N3220);
not NOT1 (N6020, N6019);
nor NOR4 (N6021, N6007, N2428, N5197, N3196);
xor XOR2 (N6022, N6013, N1355);
or OR4 (N6023, N6018, N6008, N4496, N5689);
and AND3 (N6024, N2258, N3042, N4672);
buf BUF1 (N6025, N5992);
not NOT1 (N6026, N6025);
nand NAND4 (N6027, N6026, N5261, N1757, N1930);
or OR3 (N6028, N6020, N1792, N2652);
buf BUF1 (N6029, N6024);
buf BUF1 (N6030, N6014);
nor NOR2 (N6031, N6010, N2861);
nor NOR3 (N6032, N6022, N5092, N5730);
not NOT1 (N6033, N6028);
nand NAND2 (N6034, N6033, N5025);
nor NOR4 (N6035, N6017, N3858, N3027, N1760);
buf BUF1 (N6036, N6027);
not NOT1 (N6037, N6021);
not NOT1 (N6038, N6030);
not NOT1 (N6039, N6029);
not NOT1 (N6040, N6036);
nor NOR4 (N6041, N6023, N3621, N3727, N1960);
and AND2 (N6042, N6041, N562);
buf BUF1 (N6043, N6037);
and AND4 (N6044, N6011, N4197, N5300, N1931);
not NOT1 (N6045, N6040);
or OR3 (N6046, N6035, N4516, N38);
nor NOR3 (N6047, N6045, N646, N4674);
nand NAND4 (N6048, N6047, N2823, N4702, N4485);
not NOT1 (N6049, N6034);
xor XOR2 (N6050, N6049, N1372);
nand NAND2 (N6051, N6048, N130);
not NOT1 (N6052, N6043);
buf BUF1 (N6053, N6042);
nor NOR4 (N6054, N6038, N162, N4705, N3986);
xor XOR2 (N6055, N6044, N2649);
buf BUF1 (N6056, N6031);
or OR3 (N6057, N6056, N2755, N3314);
xor XOR2 (N6058, N6054, N1891);
or OR3 (N6059, N6057, N4314, N3878);
nand NAND4 (N6060, N6032, N2394, N4486, N670);
or OR3 (N6061, N6051, N1508, N3161);
or OR4 (N6062, N6061, N1613, N4085, N4853);
buf BUF1 (N6063, N6052);
xor XOR2 (N6064, N6063, N4795);
nor NOR2 (N6065, N6039, N2085);
buf BUF1 (N6066, N6062);
nor NOR3 (N6067, N6059, N4455, N4979);
buf BUF1 (N6068, N6055);
or OR3 (N6069, N6068, N1744, N1923);
or OR2 (N6070, N6066, N4981);
and AND3 (N6071, N6069, N633, N501);
xor XOR2 (N6072, N6064, N3555);
nand NAND2 (N6073, N6058, N2277);
and AND2 (N6074, N6046, N3042);
not NOT1 (N6075, N6072);
and AND3 (N6076, N6073, N5252, N5077);
nor NOR2 (N6077, N6074, N5080);
xor XOR2 (N6078, N6065, N1733);
nand NAND2 (N6079, N6071, N3901);
or OR4 (N6080, N6079, N801, N958, N5339);
and AND4 (N6081, N6050, N3769, N1683, N5039);
nand NAND3 (N6082, N6076, N3546, N4686);
nand NAND4 (N6083, N6067, N34, N2214, N4186);
not NOT1 (N6084, N6070);
nor NOR3 (N6085, N6053, N552, N3045);
buf BUF1 (N6086, N6078);
nor NOR4 (N6087, N6080, N5162, N28, N1940);
nand NAND3 (N6088, N6060, N1711, N4803);
not NOT1 (N6089, N6082);
buf BUF1 (N6090, N6081);
not NOT1 (N6091, N6090);
or OR3 (N6092, N6084, N4130, N3773);
buf BUF1 (N6093, N6083);
not NOT1 (N6094, N6088);
nand NAND3 (N6095, N6087, N5905, N4548);
nand NAND3 (N6096, N6093, N4757, N3417);
not NOT1 (N6097, N6089);
buf BUF1 (N6098, N6086);
or OR4 (N6099, N6094, N4279, N2101, N3537);
buf BUF1 (N6100, N6092);
nor NOR3 (N6101, N6099, N1543, N3345);
not NOT1 (N6102, N6098);
xor XOR2 (N6103, N6095, N2677);
xor XOR2 (N6104, N6085, N3946);
xor XOR2 (N6105, N6102, N5694);
buf BUF1 (N6106, N6101);
not NOT1 (N6107, N6106);
or OR2 (N6108, N6103, N144);
not NOT1 (N6109, N6104);
and AND4 (N6110, N6109, N3805, N5031, N699);
xor XOR2 (N6111, N6110, N4705);
nand NAND3 (N6112, N6091, N5844, N5730);
nand NAND4 (N6113, N6096, N297, N290, N3535);
xor XOR2 (N6114, N6077, N3228);
xor XOR2 (N6115, N6108, N280);
or OR4 (N6116, N6113, N4091, N2130, N3023);
nor NOR3 (N6117, N6105, N5138, N5550);
nor NOR3 (N6118, N6115, N2868, N6082);
nand NAND4 (N6119, N6107, N5327, N963, N3250);
nand NAND4 (N6120, N6075, N2653, N3032, N428);
xor XOR2 (N6121, N6097, N5096);
xor XOR2 (N6122, N6121, N1197);
nand NAND2 (N6123, N6118, N5300);
not NOT1 (N6124, N6100);
nand NAND2 (N6125, N6112, N2170);
or OR3 (N6126, N6122, N372, N5812);
and AND3 (N6127, N6125, N6072, N4510);
nand NAND3 (N6128, N6120, N5595, N4946);
or OR4 (N6129, N6116, N1298, N3285, N3611);
or OR2 (N6130, N6128, N1559);
not NOT1 (N6131, N6129);
and AND2 (N6132, N6123, N3634);
buf BUF1 (N6133, N6126);
buf BUF1 (N6134, N6131);
xor XOR2 (N6135, N6127, N1341);
and AND4 (N6136, N6111, N3643, N4830, N2737);
xor XOR2 (N6137, N6119, N2390);
nor NOR3 (N6138, N6135, N2282, N6096);
or OR4 (N6139, N6130, N765, N1766, N2223);
nor NOR4 (N6140, N6117, N3207, N6132, N1736);
not NOT1 (N6141, N4357);
not NOT1 (N6142, N6114);
not NOT1 (N6143, N6142);
nor NOR4 (N6144, N6133, N83, N3682, N1252);
nand NAND3 (N6145, N6134, N4353, N5026);
buf BUF1 (N6146, N6144);
buf BUF1 (N6147, N6124);
and AND4 (N6148, N6143, N4605, N3233, N2246);
not NOT1 (N6149, N6146);
nor NOR4 (N6150, N6138, N4958, N243, N2363);
buf BUF1 (N6151, N6147);
not NOT1 (N6152, N6151);
or OR2 (N6153, N6149, N2507);
xor XOR2 (N6154, N6140, N5790);
not NOT1 (N6155, N6150);
buf BUF1 (N6156, N6148);
and AND2 (N6157, N6141, N3491);
not NOT1 (N6158, N6139);
buf BUF1 (N6159, N6153);
xor XOR2 (N6160, N6155, N4130);
and AND4 (N6161, N6159, N4940, N3837, N3545);
buf BUF1 (N6162, N6156);
buf BUF1 (N6163, N6137);
or OR3 (N6164, N6158, N5897, N3266);
buf BUF1 (N6165, N6161);
nand NAND3 (N6166, N6152, N306, N1865);
not NOT1 (N6167, N6136);
not NOT1 (N6168, N6160);
nor NOR2 (N6169, N6166, N2424);
not NOT1 (N6170, N6157);
or OR4 (N6171, N6168, N1686, N4039, N5219);
nor NOR2 (N6172, N6165, N3029);
or OR3 (N6173, N6170, N3665, N4277);
nor NOR4 (N6174, N6173, N274, N4884, N3656);
nand NAND2 (N6175, N6167, N4328);
nor NOR4 (N6176, N6154, N591, N5183, N2011);
xor XOR2 (N6177, N6163, N1678);
nand NAND2 (N6178, N6172, N4945);
nor NOR3 (N6179, N6174, N2454, N5285);
buf BUF1 (N6180, N6177);
and AND2 (N6181, N6179, N5154);
nand NAND4 (N6182, N6175, N1298, N1403, N332);
buf BUF1 (N6183, N6145);
not NOT1 (N6184, N6183);
buf BUF1 (N6185, N6184);
not NOT1 (N6186, N6164);
and AND4 (N6187, N6182, N3686, N4248, N3553);
nand NAND4 (N6188, N6185, N4881, N2519, N5220);
and AND3 (N6189, N6188, N3217, N5184);
not NOT1 (N6190, N6189);
or OR4 (N6191, N6171, N2478, N5619, N5690);
xor XOR2 (N6192, N6191, N2566);
not NOT1 (N6193, N6180);
buf BUF1 (N6194, N6178);
buf BUF1 (N6195, N6181);
xor XOR2 (N6196, N6192, N2188);
nor NOR4 (N6197, N6194, N1190, N2999, N2120);
or OR4 (N6198, N6195, N5981, N1462, N5999);
and AND4 (N6199, N6193, N1377, N1153, N4204);
buf BUF1 (N6200, N6187);
or OR4 (N6201, N6197, N365, N6128, N1026);
and AND2 (N6202, N6201, N4886);
not NOT1 (N6203, N6202);
or OR4 (N6204, N6198, N1688, N3435, N3950);
buf BUF1 (N6205, N6204);
or OR3 (N6206, N6186, N212, N1883);
nor NOR3 (N6207, N6199, N2369, N3186);
not NOT1 (N6208, N6200);
or OR2 (N6209, N6162, N4678);
xor XOR2 (N6210, N6169, N4659);
not NOT1 (N6211, N6206);
and AND3 (N6212, N6209, N1040, N2119);
buf BUF1 (N6213, N6210);
xor XOR2 (N6214, N6196, N3893);
not NOT1 (N6215, N6190);
and AND4 (N6216, N6212, N1804, N1573, N3766);
not NOT1 (N6217, N6215);
and AND4 (N6218, N6217, N2072, N9, N3123);
nor NOR2 (N6219, N6207, N16);
nor NOR2 (N6220, N6213, N4622);
nand NAND4 (N6221, N6205, N4551, N2461, N3744);
nor NOR2 (N6222, N6216, N1123);
nand NAND3 (N6223, N6176, N4457, N5668);
or OR2 (N6224, N6208, N557);
not NOT1 (N6225, N6214);
nand NAND2 (N6226, N6224, N4175);
nand NAND4 (N6227, N6203, N2595, N4934, N726);
nor NOR2 (N6228, N6219, N1722);
buf BUF1 (N6229, N6218);
buf BUF1 (N6230, N6222);
not NOT1 (N6231, N6230);
buf BUF1 (N6232, N6211);
nor NOR2 (N6233, N6220, N4573);
xor XOR2 (N6234, N6228, N1719);
not NOT1 (N6235, N6232);
and AND4 (N6236, N6231, N1099, N5009, N4676);
or OR4 (N6237, N6227, N1937, N4898, N4203);
not NOT1 (N6238, N6226);
nand NAND3 (N6239, N6233, N1869, N1606);
xor XOR2 (N6240, N6235, N751);
buf BUF1 (N6241, N6234);
and AND4 (N6242, N6229, N4521, N4059, N404);
xor XOR2 (N6243, N6236, N552);
and AND4 (N6244, N6242, N388, N572, N4895);
xor XOR2 (N6245, N6237, N1352);
and AND2 (N6246, N6243, N2879);
and AND3 (N6247, N6244, N4141, N4759);
or OR3 (N6248, N6241, N5448, N3502);
and AND3 (N6249, N6238, N5181, N2775);
nand NAND2 (N6250, N6247, N3070);
xor XOR2 (N6251, N6250, N4224);
not NOT1 (N6252, N6223);
buf BUF1 (N6253, N6240);
xor XOR2 (N6254, N6245, N3357);
and AND4 (N6255, N6253, N4962, N1940, N1648);
buf BUF1 (N6256, N6221);
xor XOR2 (N6257, N6256, N1022);
or OR4 (N6258, N6255, N5441, N1524, N6123);
or OR2 (N6259, N6252, N4417);
nand NAND2 (N6260, N6248, N905);
buf BUF1 (N6261, N6254);
not NOT1 (N6262, N6258);
nor NOR2 (N6263, N6249, N5126);
and AND3 (N6264, N6263, N173, N4662);
buf BUF1 (N6265, N6239);
and AND4 (N6266, N6251, N6184, N3774, N681);
and AND4 (N6267, N6257, N4278, N4858, N3044);
not NOT1 (N6268, N6259);
nor NOR3 (N6269, N6261, N5541, N4399);
nor NOR4 (N6270, N6265, N5249, N1625, N125);
buf BUF1 (N6271, N6246);
buf BUF1 (N6272, N6225);
nand NAND4 (N6273, N6272, N4709, N1737, N4242);
nor NOR2 (N6274, N6267, N4671);
not NOT1 (N6275, N6262);
xor XOR2 (N6276, N6270, N2767);
nand NAND4 (N6277, N6260, N2529, N4539, N675);
buf BUF1 (N6278, N6266);
nand NAND3 (N6279, N6269, N5872, N3997);
or OR2 (N6280, N6275, N1441);
xor XOR2 (N6281, N6279, N3475);
nor NOR3 (N6282, N6271, N1706, N255);
nand NAND3 (N6283, N6276, N1688, N4083);
nor NOR3 (N6284, N6273, N1384, N4630);
nor NOR3 (N6285, N6264, N5915, N4779);
not NOT1 (N6286, N6274);
nor NOR4 (N6287, N6286, N1244, N843, N3);
nor NOR4 (N6288, N6287, N1850, N751, N2366);
or OR2 (N6289, N6278, N1800);
nand NAND2 (N6290, N6289, N3740);
xor XOR2 (N6291, N6282, N1765);
xor XOR2 (N6292, N6281, N3772);
nand NAND3 (N6293, N6291, N5032, N6051);
buf BUF1 (N6294, N6285);
not NOT1 (N6295, N6284);
nand NAND4 (N6296, N6294, N5660, N2399, N4350);
nand NAND3 (N6297, N6283, N2850, N2158);
or OR3 (N6298, N6290, N4483, N554);
nand NAND4 (N6299, N6292, N3697, N4385, N5940);
not NOT1 (N6300, N6295);
buf BUF1 (N6301, N6288);
and AND4 (N6302, N6280, N3525, N4834, N4922);
nand NAND2 (N6303, N6300, N3734);
buf BUF1 (N6304, N6302);
not NOT1 (N6305, N6277);
xor XOR2 (N6306, N6299, N2790);
nand NAND4 (N6307, N6298, N5138, N5590, N2900);
nand NAND3 (N6308, N6306, N2250, N5459);
xor XOR2 (N6309, N6268, N6054);
and AND4 (N6310, N6296, N2435, N5492, N1624);
not NOT1 (N6311, N6293);
nand NAND3 (N6312, N6305, N5488, N4214);
xor XOR2 (N6313, N6297, N3917);
and AND3 (N6314, N6311, N5994, N2274);
or OR4 (N6315, N6314, N4312, N5943, N2281);
or OR2 (N6316, N6303, N1569);
xor XOR2 (N6317, N6304, N2751);
xor XOR2 (N6318, N6310, N1002);
not NOT1 (N6319, N6308);
xor XOR2 (N6320, N6316, N2688);
nand NAND4 (N6321, N6313, N5617, N4181, N3075);
nor NOR3 (N6322, N6312, N3148, N2777);
or OR3 (N6323, N6315, N2049, N5003);
or OR3 (N6324, N6301, N6192, N692);
buf BUF1 (N6325, N6309);
nor NOR4 (N6326, N6307, N3577, N1457, N3317);
not NOT1 (N6327, N6319);
or OR2 (N6328, N6318, N5573);
nor NOR2 (N6329, N6323, N4365);
and AND3 (N6330, N6324, N376, N4366);
nand NAND2 (N6331, N6320, N145);
and AND4 (N6332, N6322, N1988, N3529, N2006);
not NOT1 (N6333, N6332);
xor XOR2 (N6334, N6327, N4881);
not NOT1 (N6335, N6325);
not NOT1 (N6336, N6328);
nor NOR4 (N6337, N6334, N4071, N6308, N5486);
xor XOR2 (N6338, N6321, N1253);
buf BUF1 (N6339, N6330);
or OR2 (N6340, N6326, N2544);
buf BUF1 (N6341, N6317);
buf BUF1 (N6342, N6331);
xor XOR2 (N6343, N6339, N3969);
not NOT1 (N6344, N6340);
nor NOR2 (N6345, N6343, N1774);
buf BUF1 (N6346, N6345);
not NOT1 (N6347, N6341);
nand NAND3 (N6348, N6347, N3479, N2394);
nand NAND2 (N6349, N6344, N3878);
xor XOR2 (N6350, N6342, N3045);
nand NAND2 (N6351, N6337, N694);
and AND4 (N6352, N6335, N4672, N2920, N1731);
nand NAND3 (N6353, N6348, N4072, N2053);
or OR2 (N6354, N6329, N3222);
buf BUF1 (N6355, N6351);
nor NOR2 (N6356, N6333, N2686);
and AND2 (N6357, N6338, N1118);
nor NOR3 (N6358, N6353, N3533, N3421);
not NOT1 (N6359, N6355);
and AND3 (N6360, N6346, N813, N1578);
and AND4 (N6361, N6336, N504, N4055, N3261);
nand NAND2 (N6362, N6358, N3398);
buf BUF1 (N6363, N6360);
not NOT1 (N6364, N6356);
nand NAND3 (N6365, N6361, N3233, N1583);
and AND4 (N6366, N6354, N2014, N4303, N4698);
not NOT1 (N6367, N6363);
buf BUF1 (N6368, N6359);
xor XOR2 (N6369, N6364, N4040);
and AND4 (N6370, N6369, N4261, N3274, N136);
and AND3 (N6371, N6350, N2134, N3764);
nand NAND3 (N6372, N6365, N1399, N1370);
nand NAND3 (N6373, N6372, N4148, N1506);
nor NOR4 (N6374, N6373, N533, N902, N4167);
not NOT1 (N6375, N6368);
not NOT1 (N6376, N6374);
buf BUF1 (N6377, N6362);
xor XOR2 (N6378, N6370, N5272);
buf BUF1 (N6379, N6376);
xor XOR2 (N6380, N6349, N5017);
or OR2 (N6381, N6367, N3812);
xor XOR2 (N6382, N6366, N2602);
buf BUF1 (N6383, N6357);
not NOT1 (N6384, N6352);
and AND3 (N6385, N6384, N3178, N3599);
buf BUF1 (N6386, N6380);
buf BUF1 (N6387, N6379);
and AND4 (N6388, N6385, N789, N5112, N4623);
buf BUF1 (N6389, N6377);
nor NOR2 (N6390, N6389, N1154);
buf BUF1 (N6391, N6375);
nand NAND2 (N6392, N6381, N5838);
xor XOR2 (N6393, N6392, N1898);
or OR3 (N6394, N6391, N1918, N1447);
nand NAND2 (N6395, N6371, N5582);
not NOT1 (N6396, N6394);
not NOT1 (N6397, N6386);
nor NOR3 (N6398, N6396, N6133, N5351);
and AND2 (N6399, N6387, N411);
and AND3 (N6400, N6397, N2060, N340);
or OR3 (N6401, N6400, N1797, N3506);
buf BUF1 (N6402, N6401);
or OR2 (N6403, N6388, N3073);
not NOT1 (N6404, N6399);
and AND2 (N6405, N6390, N1413);
not NOT1 (N6406, N6404);
nand NAND3 (N6407, N6383, N1468, N3175);
buf BUF1 (N6408, N6378);
buf BUF1 (N6409, N6398);
nor NOR2 (N6410, N6407, N1922);
xor XOR2 (N6411, N6405, N4800);
and AND2 (N6412, N6410, N4329);
nor NOR4 (N6413, N6403, N5904, N5764, N2554);
xor XOR2 (N6414, N6382, N794);
xor XOR2 (N6415, N6411, N6314);
not NOT1 (N6416, N6406);
buf BUF1 (N6417, N6412);
xor XOR2 (N6418, N6402, N72);
nand NAND4 (N6419, N6413, N2065, N2591, N6229);
xor XOR2 (N6420, N6418, N1173);
nor NOR2 (N6421, N6408, N3695);
not NOT1 (N6422, N6414);
not NOT1 (N6423, N6395);
and AND4 (N6424, N6409, N661, N5324, N6315);
nand NAND2 (N6425, N6417, N2808);
nand NAND3 (N6426, N6416, N1354, N5632);
nand NAND3 (N6427, N6424, N159, N3363);
nand NAND2 (N6428, N6422, N2471);
nand NAND3 (N6429, N6426, N3825, N2732);
and AND2 (N6430, N6427, N2799);
or OR2 (N6431, N6429, N6199);
or OR4 (N6432, N6393, N5762, N5825, N5347);
xor XOR2 (N6433, N6428, N1924);
buf BUF1 (N6434, N6420);
nor NOR3 (N6435, N6415, N4826, N5656);
nand NAND2 (N6436, N6423, N4404);
xor XOR2 (N6437, N6421, N1076);
nand NAND3 (N6438, N6432, N2916, N2240);
xor XOR2 (N6439, N6430, N1524);
xor XOR2 (N6440, N6438, N5259);
and AND4 (N6441, N6433, N6399, N5410, N3039);
or OR3 (N6442, N6439, N5291, N17);
or OR2 (N6443, N6436, N4949);
nor NOR4 (N6444, N6437, N5614, N4879, N4628);
nor NOR2 (N6445, N6434, N3435);
nor NOR4 (N6446, N6431, N6189, N4676, N1228);
nand NAND4 (N6447, N6425, N568, N2465, N4400);
or OR4 (N6448, N6443, N5437, N6214, N1497);
nand NAND4 (N6449, N6435, N5371, N5835, N440);
and AND3 (N6450, N6440, N1762, N4510);
nand NAND2 (N6451, N6442, N542);
nor NOR2 (N6452, N6445, N6172);
not NOT1 (N6453, N6451);
or OR3 (N6454, N6449, N520, N5941);
buf BUF1 (N6455, N6441);
or OR4 (N6456, N6452, N1985, N1160, N6264);
not NOT1 (N6457, N6444);
not NOT1 (N6458, N6454);
not NOT1 (N6459, N6419);
or OR4 (N6460, N6453, N2385, N5191, N3482);
nand NAND4 (N6461, N6446, N3292, N514, N3160);
not NOT1 (N6462, N6458);
nand NAND4 (N6463, N6459, N5124, N4650, N5542);
nand NAND4 (N6464, N6447, N2249, N3300, N2124);
buf BUF1 (N6465, N6461);
xor XOR2 (N6466, N6463, N4741);
xor XOR2 (N6467, N6455, N3386);
not NOT1 (N6468, N6450);
nor NOR2 (N6469, N6468, N1789);
and AND4 (N6470, N6464, N6044, N3038, N1742);
nand NAND3 (N6471, N6448, N5501, N1123);
and AND2 (N6472, N6470, N1612);
not NOT1 (N6473, N6472);
not NOT1 (N6474, N6465);
or OR3 (N6475, N6467, N4818, N81);
and AND4 (N6476, N6469, N4351, N6145, N1125);
not NOT1 (N6477, N6462);
xor XOR2 (N6478, N6460, N2758);
nand NAND3 (N6479, N6457, N4442, N5800);
not NOT1 (N6480, N6477);
buf BUF1 (N6481, N6478);
and AND2 (N6482, N6471, N5756);
xor XOR2 (N6483, N6466, N4670);
and AND3 (N6484, N6456, N5754, N2589);
nand NAND2 (N6485, N6484, N1476);
buf BUF1 (N6486, N6485);
nand NAND4 (N6487, N6476, N4578, N5742, N2739);
nor NOR2 (N6488, N6474, N2985);
not NOT1 (N6489, N6486);
and AND2 (N6490, N6480, N533);
and AND2 (N6491, N6487, N5772);
nand NAND3 (N6492, N6475, N683, N610);
and AND3 (N6493, N6489, N5301, N5382);
buf BUF1 (N6494, N6482);
nor NOR4 (N6495, N6493, N31, N4818, N1676);
or OR3 (N6496, N6492, N708, N6386);
and AND2 (N6497, N6473, N733);
xor XOR2 (N6498, N6488, N4958);
buf BUF1 (N6499, N6496);
nand NAND2 (N6500, N6499, N4651);
nand NAND4 (N6501, N6500, N6082, N3555, N4925);
nor NOR4 (N6502, N6491, N768, N5567, N1790);
not NOT1 (N6503, N6483);
and AND3 (N6504, N6490, N4840, N5726);
nand NAND3 (N6505, N6479, N5297, N6061);
nor NOR2 (N6506, N6501, N782);
and AND3 (N6507, N6494, N4067, N3252);
not NOT1 (N6508, N6498);
or OR2 (N6509, N6503, N6489);
or OR2 (N6510, N6495, N1492);
or OR3 (N6511, N6506, N2137, N5929);
xor XOR2 (N6512, N6511, N410);
and AND2 (N6513, N6508, N4216);
and AND3 (N6514, N6509, N3273, N2637);
buf BUF1 (N6515, N6497);
not NOT1 (N6516, N6515);
not NOT1 (N6517, N6513);
not NOT1 (N6518, N6516);
or OR4 (N6519, N6502, N4476, N934, N5747);
xor XOR2 (N6520, N6510, N2061);
buf BUF1 (N6521, N6517);
or OR4 (N6522, N6504, N4846, N3210, N1904);
and AND4 (N6523, N6518, N2232, N418, N6461);
and AND2 (N6524, N6514, N4739);
nor NOR4 (N6525, N6505, N2999, N4366, N2069);
nand NAND2 (N6526, N6525, N4731);
and AND4 (N6527, N6507, N2513, N5796, N1837);
nor NOR2 (N6528, N6527, N4004);
or OR4 (N6529, N6521, N23, N117, N2476);
nand NAND2 (N6530, N6529, N4940);
or OR4 (N6531, N6523, N4414, N4148, N3393);
and AND3 (N6532, N6526, N3538, N4053);
or OR3 (N6533, N6522, N1453, N2547);
and AND4 (N6534, N6528, N4060, N257, N701);
and AND4 (N6535, N6534, N1363, N688, N4967);
nand NAND2 (N6536, N6524, N74);
or OR3 (N6537, N6512, N578, N2817);
nor NOR4 (N6538, N6537, N801, N5254, N4228);
nand NAND4 (N6539, N6520, N2880, N872, N3026);
and AND2 (N6540, N6532, N2853);
buf BUF1 (N6541, N6539);
not NOT1 (N6542, N6536);
nand NAND3 (N6543, N6541, N3017, N1458);
and AND2 (N6544, N6543, N228);
and AND2 (N6545, N6531, N4204);
xor XOR2 (N6546, N6542, N2714);
xor XOR2 (N6547, N6481, N6184);
buf BUF1 (N6548, N6545);
or OR2 (N6549, N6546, N3962);
xor XOR2 (N6550, N6548, N5609);
nor NOR3 (N6551, N6533, N1859, N4396);
nor NOR2 (N6552, N6535, N4771);
xor XOR2 (N6553, N6551, N286);
xor XOR2 (N6554, N6530, N5813);
buf BUF1 (N6555, N6547);
or OR4 (N6556, N6554, N4142, N4255, N1913);
or OR2 (N6557, N6556, N670);
nand NAND2 (N6558, N6540, N3708);
nor NOR2 (N6559, N6558, N418);
and AND3 (N6560, N6544, N4309, N3133);
or OR2 (N6561, N6552, N2716);
nand NAND2 (N6562, N6560, N748);
and AND4 (N6563, N6519, N559, N2815, N2576);
buf BUF1 (N6564, N6553);
or OR3 (N6565, N6557, N4441, N3475);
nor NOR3 (N6566, N6563, N710, N4785);
nand NAND3 (N6567, N6562, N2729, N644);
nand NAND4 (N6568, N6567, N6044, N2875, N4649);
and AND4 (N6569, N6555, N1885, N2291, N3379);
xor XOR2 (N6570, N6564, N3427);
or OR4 (N6571, N6550, N4953, N1361, N5651);
and AND3 (N6572, N6538, N5431, N2008);
nand NAND4 (N6573, N6561, N6384, N4596, N3690);
not NOT1 (N6574, N6571);
xor XOR2 (N6575, N6559, N777);
and AND4 (N6576, N6574, N6255, N1909, N2630);
not NOT1 (N6577, N6569);
buf BUF1 (N6578, N6576);
and AND2 (N6579, N6573, N730);
and AND4 (N6580, N6566, N4920, N2089, N2072);
buf BUF1 (N6581, N6570);
or OR2 (N6582, N6578, N498);
not NOT1 (N6583, N6575);
buf BUF1 (N6584, N6582);
xor XOR2 (N6585, N6577, N4590);
not NOT1 (N6586, N6580);
nand NAND4 (N6587, N6572, N305, N2431, N6033);
not NOT1 (N6588, N6585);
not NOT1 (N6589, N6568);
or OR3 (N6590, N6586, N4831, N4356);
xor XOR2 (N6591, N6587, N5644);
xor XOR2 (N6592, N6565, N3523);
or OR2 (N6593, N6581, N3213);
or OR2 (N6594, N6590, N4457);
buf BUF1 (N6595, N6589);
or OR3 (N6596, N6549, N3852, N1225);
not NOT1 (N6597, N6595);
nor NOR2 (N6598, N6593, N1551);
or OR2 (N6599, N6596, N2681);
not NOT1 (N6600, N6579);
nand NAND4 (N6601, N6591, N4521, N1432, N3107);
buf BUF1 (N6602, N6597);
or OR4 (N6603, N6592, N5969, N608, N2169);
or OR3 (N6604, N6599, N5692, N6373);
nand NAND3 (N6605, N6588, N2032, N4848);
buf BUF1 (N6606, N6605);
and AND3 (N6607, N6598, N1515, N534);
not NOT1 (N6608, N6584);
nor NOR3 (N6609, N6602, N5837, N1400);
buf BUF1 (N6610, N6594);
buf BUF1 (N6611, N6583);
or OR4 (N6612, N6601, N3276, N37, N5649);
nor NOR2 (N6613, N6608, N4987);
and AND2 (N6614, N6604, N552);
and AND4 (N6615, N6610, N1495, N3836, N2511);
and AND2 (N6616, N6607, N6360);
nand NAND3 (N6617, N6613, N4146, N67);
nand NAND2 (N6618, N6614, N2665);
and AND3 (N6619, N6615, N2786, N2390);
buf BUF1 (N6620, N6617);
not NOT1 (N6621, N6612);
nor NOR2 (N6622, N6606, N5293);
and AND2 (N6623, N6621, N451);
and AND3 (N6624, N6603, N1419, N1908);
xor XOR2 (N6625, N6623, N5881);
nand NAND3 (N6626, N6622, N5589, N4315);
buf BUF1 (N6627, N6624);
xor XOR2 (N6628, N6616, N4385);
not NOT1 (N6629, N6600);
nor NOR3 (N6630, N6629, N5491, N6131);
buf BUF1 (N6631, N6628);
buf BUF1 (N6632, N6630);
xor XOR2 (N6633, N6632, N6445);
buf BUF1 (N6634, N6626);
nand NAND4 (N6635, N6619, N2837, N1530, N3131);
and AND3 (N6636, N6611, N5150, N4175);
not NOT1 (N6637, N6635);
and AND3 (N6638, N6627, N2143, N5988);
nand NAND2 (N6639, N6638, N2607);
xor XOR2 (N6640, N6633, N5800);
nor NOR4 (N6641, N6631, N2921, N3940, N70);
buf BUF1 (N6642, N6640);
and AND2 (N6643, N6634, N3805);
nand NAND2 (N6644, N6636, N495);
xor XOR2 (N6645, N6609, N4291);
or OR2 (N6646, N6644, N6170);
nand NAND4 (N6647, N6639, N4396, N3610, N3292);
and AND2 (N6648, N6642, N1649);
nand NAND2 (N6649, N6641, N2381);
and AND4 (N6650, N6646, N3908, N1141, N2968);
not NOT1 (N6651, N6648);
not NOT1 (N6652, N6651);
buf BUF1 (N6653, N6649);
nor NOR3 (N6654, N6618, N1377, N688);
not NOT1 (N6655, N6643);
buf BUF1 (N6656, N6620);
not NOT1 (N6657, N6654);
or OR3 (N6658, N6653, N1967, N2819);
not NOT1 (N6659, N6637);
buf BUF1 (N6660, N6658);
nand NAND4 (N6661, N6660, N457, N2810, N771);
and AND3 (N6662, N6657, N5648, N5654);
nor NOR2 (N6663, N6652, N975);
not NOT1 (N6664, N6655);
buf BUF1 (N6665, N6663);
and AND3 (N6666, N6661, N6058, N4331);
or OR3 (N6667, N6625, N768, N777);
and AND2 (N6668, N6665, N4273);
xor XOR2 (N6669, N6666, N5769);
and AND2 (N6670, N6669, N3898);
or OR3 (N6671, N6659, N2034, N6123);
not NOT1 (N6672, N6647);
or OR3 (N6673, N6671, N3531, N4401);
not NOT1 (N6674, N6668);
nand NAND4 (N6675, N6670, N2105, N1378, N2371);
nand NAND2 (N6676, N6673, N3376);
or OR3 (N6677, N6650, N670, N6457);
or OR4 (N6678, N6645, N3690, N2899, N774);
xor XOR2 (N6679, N6656, N3930);
and AND2 (N6680, N6677, N6231);
not NOT1 (N6681, N6678);
and AND2 (N6682, N6662, N4831);
nand NAND4 (N6683, N6664, N2566, N3440, N6258);
nand NAND2 (N6684, N6681, N3702);
nand NAND2 (N6685, N6679, N2832);
and AND3 (N6686, N6684, N1725, N6177);
nor NOR4 (N6687, N6680, N199, N1461, N5014);
xor XOR2 (N6688, N6672, N5354);
nor NOR3 (N6689, N6683, N3724, N724);
nand NAND2 (N6690, N6675, N4682);
not NOT1 (N6691, N6686);
xor XOR2 (N6692, N6687, N5213);
xor XOR2 (N6693, N6676, N309);
xor XOR2 (N6694, N6689, N1303);
or OR2 (N6695, N6674, N3925);
xor XOR2 (N6696, N6695, N6349);
or OR3 (N6697, N6685, N440, N1598);
and AND2 (N6698, N6692, N2484);
and AND4 (N6699, N6667, N2935, N6292, N1540);
xor XOR2 (N6700, N6691, N5319);
and AND4 (N6701, N6693, N3172, N6178, N3490);
nor NOR3 (N6702, N6700, N2698, N600);
nand NAND2 (N6703, N6682, N5330);
or OR2 (N6704, N6697, N2094);
not NOT1 (N6705, N6690);
nor NOR3 (N6706, N6703, N3870, N1762);
not NOT1 (N6707, N6706);
xor XOR2 (N6708, N6702, N3061);
buf BUF1 (N6709, N6694);
nand NAND4 (N6710, N6708, N6182, N3312, N1886);
nand NAND3 (N6711, N6696, N6137, N6458);
not NOT1 (N6712, N6709);
nand NAND4 (N6713, N6701, N3245, N1770, N4526);
or OR4 (N6714, N6704, N2263, N5004, N1186);
buf BUF1 (N6715, N6712);
nor NOR3 (N6716, N6707, N330, N1873);
buf BUF1 (N6717, N6716);
not NOT1 (N6718, N6688);
or OR2 (N6719, N6714, N3988);
not NOT1 (N6720, N6711);
nor NOR4 (N6721, N6710, N2908, N3043, N1955);
or OR2 (N6722, N6720, N1298);
nor NOR3 (N6723, N6719, N6427, N2444);
xor XOR2 (N6724, N6705, N2884);
nor NOR2 (N6725, N6722, N6365);
not NOT1 (N6726, N6723);
buf BUF1 (N6727, N6724);
and AND4 (N6728, N6715, N6668, N4848, N835);
and AND3 (N6729, N6727, N712, N1101);
or OR4 (N6730, N6718, N4203, N5774, N4174);
or OR4 (N6731, N6728, N971, N894, N3403);
and AND2 (N6732, N6729, N5629);
nor NOR2 (N6733, N6713, N6073);
buf BUF1 (N6734, N6732);
or OR4 (N6735, N6731, N2720, N907, N5594);
buf BUF1 (N6736, N6726);
xor XOR2 (N6737, N6698, N1724);
not NOT1 (N6738, N6717);
or OR2 (N6739, N6737, N3416);
nand NAND2 (N6740, N6699, N4509);
nand NAND4 (N6741, N6725, N373, N554, N31);
or OR3 (N6742, N6740, N39, N6331);
nor NOR2 (N6743, N6735, N3266);
not NOT1 (N6744, N6738);
and AND3 (N6745, N6734, N4572, N1812);
nand NAND4 (N6746, N6730, N1563, N1283, N2862);
xor XOR2 (N6747, N6721, N5460);
xor XOR2 (N6748, N6744, N6603);
xor XOR2 (N6749, N6733, N2679);
and AND2 (N6750, N6749, N2624);
not NOT1 (N6751, N6745);
xor XOR2 (N6752, N6750, N3347);
nand NAND4 (N6753, N6747, N1607, N1295, N3189);
xor XOR2 (N6754, N6739, N6388);
or OR4 (N6755, N6754, N4475, N931, N5615);
buf BUF1 (N6756, N6746);
buf BUF1 (N6757, N6756);
and AND4 (N6758, N6741, N1730, N4709, N5500);
buf BUF1 (N6759, N6758);
buf BUF1 (N6760, N6757);
buf BUF1 (N6761, N6742);
nor NOR3 (N6762, N6751, N5462, N384);
xor XOR2 (N6763, N6760, N3472);
or OR2 (N6764, N6743, N4608);
and AND4 (N6765, N6762, N6721, N1003, N676);
and AND3 (N6766, N6752, N3006, N3979);
and AND3 (N6767, N6748, N6428, N828);
xor XOR2 (N6768, N6755, N1201);
buf BUF1 (N6769, N6763);
and AND2 (N6770, N6769, N2505);
buf BUF1 (N6771, N6767);
or OR2 (N6772, N6766, N3384);
or OR2 (N6773, N6736, N5862);
nand NAND4 (N6774, N6773, N4345, N4690, N68);
xor XOR2 (N6775, N6765, N5657);
xor XOR2 (N6776, N6753, N1762);
nand NAND3 (N6777, N6759, N2645, N1950);
xor XOR2 (N6778, N6776, N273);
not NOT1 (N6779, N6775);
or OR3 (N6780, N6761, N1538, N2307);
and AND4 (N6781, N6764, N5760, N3270, N5317);
not NOT1 (N6782, N6781);
xor XOR2 (N6783, N6778, N4691);
buf BUF1 (N6784, N6772);
nand NAND2 (N6785, N6779, N3419);
buf BUF1 (N6786, N6771);
nand NAND4 (N6787, N6780, N5252, N5238, N6689);
nand NAND3 (N6788, N6785, N2632, N853);
not NOT1 (N6789, N6784);
nor NOR3 (N6790, N6777, N1829, N6593);
nand NAND4 (N6791, N6770, N5183, N4923, N1579);
nand NAND3 (N6792, N6790, N2954, N483);
xor XOR2 (N6793, N6782, N2153);
or OR4 (N6794, N6787, N382, N1252, N2777);
and AND4 (N6795, N6792, N214, N1222, N3652);
not NOT1 (N6796, N6791);
and AND3 (N6797, N6788, N2764, N2626);
not NOT1 (N6798, N6783);
buf BUF1 (N6799, N6794);
nand NAND4 (N6800, N6768, N3726, N3851, N2593);
nand NAND4 (N6801, N6796, N2390, N6095, N3056);
buf BUF1 (N6802, N6801);
not NOT1 (N6803, N6798);
nand NAND4 (N6804, N6799, N6683, N2728, N2308);
xor XOR2 (N6805, N6786, N2653);
nor NOR2 (N6806, N6804, N6456);
xor XOR2 (N6807, N6805, N1850);
not NOT1 (N6808, N6774);
nand NAND3 (N6809, N6806, N162, N4235);
or OR3 (N6810, N6802, N5837, N4739);
and AND2 (N6811, N6789, N2634);
buf BUF1 (N6812, N6809);
nand NAND4 (N6813, N6797, N3204, N291, N343);
buf BUF1 (N6814, N6810);
buf BUF1 (N6815, N6808);
nor NOR3 (N6816, N6814, N3098, N4097);
nand NAND4 (N6817, N6800, N5753, N263, N22);
nand NAND2 (N6818, N6795, N2185);
nand NAND3 (N6819, N6812, N5155, N2521);
buf BUF1 (N6820, N6811);
nor NOR3 (N6821, N6820, N6542, N1357);
nor NOR3 (N6822, N6817, N2863, N2764);
and AND2 (N6823, N6813, N5508);
nor NOR3 (N6824, N6807, N4783, N3312);
buf BUF1 (N6825, N6803);
nor NOR3 (N6826, N6821, N1432, N4461);
xor XOR2 (N6827, N6815, N1188);
buf BUF1 (N6828, N6793);
nand NAND2 (N6829, N6816, N6019);
and AND2 (N6830, N6823, N5642);
nor NOR2 (N6831, N6830, N5075);
xor XOR2 (N6832, N6818, N1908);
or OR3 (N6833, N6832, N3411, N4013);
nand NAND2 (N6834, N6829, N5484);
and AND4 (N6835, N6819, N290, N2527, N2796);
buf BUF1 (N6836, N6822);
nand NAND3 (N6837, N6833, N4649, N2770);
xor XOR2 (N6838, N6837, N2361);
not NOT1 (N6839, N6838);
xor XOR2 (N6840, N6836, N5245);
nor NOR4 (N6841, N6825, N1477, N6678, N4366);
and AND4 (N6842, N6839, N5159, N4683, N5193);
nand NAND3 (N6843, N6828, N2573, N1205);
nor NOR4 (N6844, N6831, N2100, N1139, N4952);
nand NAND3 (N6845, N6840, N1129, N1914);
or OR2 (N6846, N6827, N5334);
xor XOR2 (N6847, N6844, N5289);
xor XOR2 (N6848, N6847, N5253);
or OR4 (N6849, N6846, N5028, N5083, N6186);
nand NAND3 (N6850, N6826, N1600, N495);
and AND3 (N6851, N6824, N977, N3714);
nand NAND3 (N6852, N6851, N4257, N659);
or OR4 (N6853, N6849, N2756, N1907, N3350);
buf BUF1 (N6854, N6842);
and AND4 (N6855, N6834, N2948, N4014, N2024);
xor XOR2 (N6856, N6852, N6262);
or OR4 (N6857, N6843, N6117, N4099, N6057);
nor NOR2 (N6858, N6853, N6382);
or OR4 (N6859, N6845, N6655, N5716, N238);
not NOT1 (N6860, N6855);
nand NAND2 (N6861, N6848, N629);
nor NOR3 (N6862, N6856, N581, N3259);
or OR2 (N6863, N6841, N6143);
buf BUF1 (N6864, N6863);
and AND2 (N6865, N6857, N5288);
or OR4 (N6866, N6860, N4499, N3143, N6701);
and AND4 (N6867, N6858, N3017, N3471, N5897);
nor NOR4 (N6868, N6859, N829, N55, N1495);
not NOT1 (N6869, N6866);
xor XOR2 (N6870, N6850, N6007);
or OR3 (N6871, N6870, N744, N3644);
nor NOR3 (N6872, N6835, N4695, N5406);
or OR4 (N6873, N6872, N6031, N6710, N3180);
nor NOR2 (N6874, N6869, N4635);
or OR2 (N6875, N6867, N6318);
not NOT1 (N6876, N6873);
nand NAND4 (N6877, N6875, N4388, N2173, N2336);
xor XOR2 (N6878, N6861, N4471);
buf BUF1 (N6879, N6874);
or OR3 (N6880, N6864, N139, N2186);
nor NOR3 (N6881, N6878, N3650, N3117);
buf BUF1 (N6882, N6877);
and AND3 (N6883, N6879, N65, N1342);
not NOT1 (N6884, N6865);
and AND3 (N6885, N6880, N5744, N5764);
nor NOR2 (N6886, N6883, N1268);
or OR4 (N6887, N6884, N1125, N3950, N5433);
buf BUF1 (N6888, N6881);
and AND3 (N6889, N6887, N3397, N5203);
nand NAND4 (N6890, N6868, N5411, N1812, N229);
or OR3 (N6891, N6876, N4544, N3655);
nor NOR4 (N6892, N6885, N5086, N3393, N6074);
and AND4 (N6893, N6854, N292, N3037, N960);
and AND4 (N6894, N6893, N5401, N3699, N317);
xor XOR2 (N6895, N6882, N306);
or OR2 (N6896, N6891, N5928);
not NOT1 (N6897, N6889);
and AND2 (N6898, N6862, N4722);
and AND3 (N6899, N6898, N1750, N3030);
or OR4 (N6900, N6890, N5576, N2541, N554);
buf BUF1 (N6901, N6892);
not NOT1 (N6902, N6901);
xor XOR2 (N6903, N6896, N3988);
xor XOR2 (N6904, N6888, N3923);
or OR3 (N6905, N6894, N215, N5919);
nand NAND4 (N6906, N6902, N5737, N4974, N4964);
nand NAND3 (N6907, N6903, N2786, N6466);
nand NAND2 (N6908, N6899, N3743);
or OR4 (N6909, N6871, N6861, N4057, N2401);
not NOT1 (N6910, N6909);
nor NOR2 (N6911, N6906, N3070);
buf BUF1 (N6912, N6908);
buf BUF1 (N6913, N6910);
xor XOR2 (N6914, N6895, N4294);
nand NAND3 (N6915, N6912, N2990, N1448);
not NOT1 (N6916, N6897);
xor XOR2 (N6917, N6900, N4269);
not NOT1 (N6918, N6914);
nand NAND2 (N6919, N6916, N4540);
xor XOR2 (N6920, N6915, N4280);
xor XOR2 (N6921, N6905, N3255);
not NOT1 (N6922, N6917);
xor XOR2 (N6923, N6907, N2420);
nor NOR3 (N6924, N6921, N6073, N6433);
and AND2 (N6925, N6918, N4695);
nor NOR3 (N6926, N6925, N1348, N6452);
or OR2 (N6927, N6920, N6266);
xor XOR2 (N6928, N6924, N4027);
nand NAND2 (N6929, N6919, N5075);
or OR2 (N6930, N6904, N2782);
not NOT1 (N6931, N6886);
and AND2 (N6932, N6930, N5829);
and AND3 (N6933, N6923, N5103, N878);
or OR4 (N6934, N6926, N1811, N5912, N3831);
and AND4 (N6935, N6913, N5651, N239, N935);
xor XOR2 (N6936, N6931, N6329);
and AND2 (N6937, N6929, N954);
buf BUF1 (N6938, N6927);
or OR2 (N6939, N6936, N6833);
nand NAND4 (N6940, N6911, N1714, N2849, N6772);
and AND2 (N6941, N6922, N2584);
and AND3 (N6942, N6940, N5908, N5270);
and AND4 (N6943, N6938, N3800, N385, N3697);
xor XOR2 (N6944, N6928, N6682);
and AND2 (N6945, N6941, N705);
or OR4 (N6946, N6944, N3867, N4223, N6462);
nor NOR3 (N6947, N6937, N3191, N3829);
not NOT1 (N6948, N6942);
not NOT1 (N6949, N6933);
or OR3 (N6950, N6934, N5870, N4442);
nand NAND2 (N6951, N6949, N1718);
or OR2 (N6952, N6935, N5900);
nand NAND4 (N6953, N6948, N4923, N3935, N6158);
nand NAND2 (N6954, N6950, N2523);
buf BUF1 (N6955, N6946);
nand NAND4 (N6956, N6951, N2767, N2922, N554);
buf BUF1 (N6957, N6939);
or OR3 (N6958, N6943, N2964, N689);
nand NAND4 (N6959, N6958, N5730, N2696, N5002);
buf BUF1 (N6960, N6959);
or OR2 (N6961, N6945, N4856);
and AND3 (N6962, N6955, N6917, N6027);
nand NAND3 (N6963, N6956, N2609, N1036);
xor XOR2 (N6964, N6954, N2002);
or OR3 (N6965, N6962, N2565, N5428);
and AND2 (N6966, N6932, N2737);
nand NAND4 (N6967, N6963, N1793, N2583, N4008);
and AND2 (N6968, N6961, N6467);
not NOT1 (N6969, N6960);
nand NAND4 (N6970, N6969, N6002, N1145, N591);
and AND2 (N6971, N6957, N690);
or OR4 (N6972, N6966, N6872, N6618, N2510);
not NOT1 (N6973, N6965);
nor NOR2 (N6974, N6971, N2627);
and AND2 (N6975, N6973, N6758);
nor NOR4 (N6976, N6967, N1801, N705, N4292);
or OR3 (N6977, N6964, N1078, N4868);
nand NAND2 (N6978, N6970, N3234);
nand NAND3 (N6979, N6975, N5688, N5517);
buf BUF1 (N6980, N6976);
nand NAND4 (N6981, N6952, N3914, N5069, N6007);
nand NAND4 (N6982, N6974, N6097, N2640, N4710);
nor NOR2 (N6983, N6968, N946);
nor NOR2 (N6984, N6980, N1014);
or OR4 (N6985, N6984, N105, N781, N3880);
nand NAND3 (N6986, N6982, N6557, N362);
buf BUF1 (N6987, N6979);
nor NOR3 (N6988, N6985, N5034, N6219);
xor XOR2 (N6989, N6988, N4999);
nand NAND2 (N6990, N6989, N5662);
nor NOR4 (N6991, N6986, N2044, N1238, N2878);
nand NAND2 (N6992, N6987, N4363);
nand NAND4 (N6993, N6990, N1933, N6844, N2303);
xor XOR2 (N6994, N6993, N420);
not NOT1 (N6995, N6977);
nor NOR2 (N6996, N6992, N3936);
not NOT1 (N6997, N6953);
xor XOR2 (N6998, N6972, N2076);
xor XOR2 (N6999, N6995, N5294);
xor XOR2 (N7000, N6981, N6982);
nand NAND2 (N7001, N7000, N3100);
buf BUF1 (N7002, N7001);
and AND3 (N7003, N6991, N6694, N6221);
and AND2 (N7004, N6983, N5161);
or OR4 (N7005, N6947, N4586, N1060, N5384);
or OR4 (N7006, N6999, N2811, N3291, N4468);
buf BUF1 (N7007, N7003);
xor XOR2 (N7008, N6997, N2611);
nor NOR3 (N7009, N7005, N2017, N4106);
nor NOR3 (N7010, N6998, N6799, N6008);
buf BUF1 (N7011, N7008);
nor NOR4 (N7012, N6996, N217, N3380, N5748);
buf BUF1 (N7013, N7010);
nand NAND2 (N7014, N6994, N5512);
not NOT1 (N7015, N7007);
not NOT1 (N7016, N7013);
and AND2 (N7017, N7006, N3136);
not NOT1 (N7018, N7012);
and AND2 (N7019, N7014, N5806);
nor NOR2 (N7020, N7016, N2388);
nand NAND3 (N7021, N7002, N3961, N473);
or OR2 (N7022, N7020, N2331);
buf BUF1 (N7023, N7011);
nor NOR2 (N7024, N7022, N2731);
nand NAND2 (N7025, N7019, N1026);
or OR4 (N7026, N7018, N4079, N1913, N738);
nand NAND3 (N7027, N7024, N4950, N4646);
nor NOR2 (N7028, N7021, N6500);
nand NAND3 (N7029, N7017, N5962, N5199);
buf BUF1 (N7030, N7015);
not NOT1 (N7031, N6978);
or OR2 (N7032, N7023, N6797);
not NOT1 (N7033, N7031);
not NOT1 (N7034, N7029);
xor XOR2 (N7035, N7004, N1236);
or OR3 (N7036, N7032, N6942, N6185);
not NOT1 (N7037, N7026);
xor XOR2 (N7038, N7030, N2435);
nor NOR4 (N7039, N7035, N1526, N745, N2549);
nand NAND4 (N7040, N7034, N6562, N3417, N715);
or OR2 (N7041, N7036, N6536);
and AND2 (N7042, N7038, N606);
xor XOR2 (N7043, N7037, N1555);
nor NOR4 (N7044, N7043, N2182, N2278, N86);
and AND2 (N7045, N7041, N1240);
not NOT1 (N7046, N7009);
and AND3 (N7047, N7039, N1064, N335);
or OR4 (N7048, N7044, N4911, N1400, N382);
buf BUF1 (N7049, N7042);
buf BUF1 (N7050, N7045);
nor NOR2 (N7051, N7050, N4458);
or OR3 (N7052, N7047, N3113, N1696);
nand NAND4 (N7053, N7040, N4794, N5302, N2243);
buf BUF1 (N7054, N7049);
buf BUF1 (N7055, N7028);
and AND2 (N7056, N7051, N2557);
and AND4 (N7057, N7027, N4884, N5824, N4627);
and AND4 (N7058, N7053, N4336, N2878, N2280);
xor XOR2 (N7059, N7046, N6633);
buf BUF1 (N7060, N7052);
or OR2 (N7061, N7048, N5028);
or OR2 (N7062, N7055, N1133);
buf BUF1 (N7063, N7061);
and AND2 (N7064, N7063, N4890);
and AND3 (N7065, N7025, N1110, N691);
xor XOR2 (N7066, N7056, N6703);
buf BUF1 (N7067, N7065);
buf BUF1 (N7068, N7060);
xor XOR2 (N7069, N7058, N5757);
xor XOR2 (N7070, N7067, N6482);
and AND4 (N7071, N7069, N4333, N4723, N6181);
not NOT1 (N7072, N7057);
xor XOR2 (N7073, N7033, N2455);
buf BUF1 (N7074, N7054);
xor XOR2 (N7075, N7071, N4538);
and AND2 (N7076, N7068, N5238);
xor XOR2 (N7077, N7064, N2084);
not NOT1 (N7078, N7062);
not NOT1 (N7079, N7059);
not NOT1 (N7080, N7075);
and AND3 (N7081, N7072, N4842, N5239);
and AND2 (N7082, N7077, N4700);
and AND4 (N7083, N7074, N6830, N5041, N4896);
nand NAND4 (N7084, N7070, N3552, N51, N3962);
nor NOR3 (N7085, N7082, N744, N3676);
xor XOR2 (N7086, N7079, N5739);
not NOT1 (N7087, N7081);
and AND3 (N7088, N7083, N2940, N4378);
not NOT1 (N7089, N7084);
nor NOR3 (N7090, N7066, N6840, N615);
or OR3 (N7091, N7086, N3928, N6970);
nor NOR2 (N7092, N7080, N1857);
nand NAND4 (N7093, N7085, N5190, N953, N2995);
or OR2 (N7094, N7091, N4254);
and AND3 (N7095, N7092, N2948, N458);
nand NAND2 (N7096, N7094, N3108);
nand NAND4 (N7097, N7073, N6101, N5762, N3812);
and AND3 (N7098, N7090, N5298, N1435);
nor NOR2 (N7099, N7096, N5766);
nor NOR4 (N7100, N7078, N370, N1827, N544);
nand NAND2 (N7101, N7093, N7077);
nor NOR2 (N7102, N7076, N710);
buf BUF1 (N7103, N7087);
or OR2 (N7104, N7095, N1466);
or OR3 (N7105, N7098, N5715, N3112);
nand NAND2 (N7106, N7088, N6177);
nand NAND2 (N7107, N7089, N2151);
or OR3 (N7108, N7106, N3721, N3840);
or OR3 (N7109, N7104, N5914, N1026);
xor XOR2 (N7110, N7101, N207);
nor NOR2 (N7111, N7099, N1029);
nor NOR3 (N7112, N7107, N575, N5118);
or OR4 (N7113, N7105, N1818, N6573, N7018);
not NOT1 (N7114, N7100);
xor XOR2 (N7115, N7111, N5634);
nor NOR2 (N7116, N7115, N1175);
nor NOR4 (N7117, N7116, N3497, N2253, N6019);
nand NAND3 (N7118, N7110, N7016, N353);
xor XOR2 (N7119, N7112, N1845);
nand NAND2 (N7120, N7117, N6506);
buf BUF1 (N7121, N7097);
nor NOR4 (N7122, N7113, N4046, N5815, N91);
or OR3 (N7123, N7114, N5411, N1944);
nand NAND3 (N7124, N7118, N4708, N4739);
and AND3 (N7125, N7108, N2838, N751);
buf BUF1 (N7126, N7119);
or OR3 (N7127, N7103, N5867, N6496);
nor NOR3 (N7128, N7127, N1855, N4419);
not NOT1 (N7129, N7125);
nor NOR4 (N7130, N7121, N4596, N247, N5751);
or OR3 (N7131, N7109, N5840, N6103);
and AND2 (N7132, N7124, N3965);
or OR2 (N7133, N7123, N1807);
nor NOR2 (N7134, N7120, N1938);
xor XOR2 (N7135, N7132, N3149);
not NOT1 (N7136, N7133);
xor XOR2 (N7137, N7131, N6083);
buf BUF1 (N7138, N7129);
or OR2 (N7139, N7138, N5756);
nor NOR4 (N7140, N7137, N5186, N6609, N950);
nor NOR3 (N7141, N7135, N5276, N2590);
and AND2 (N7142, N7102, N3977);
and AND4 (N7143, N7139, N6959, N4965, N1941);
nor NOR3 (N7144, N7126, N5071, N824);
nand NAND2 (N7145, N7134, N6676);
buf BUF1 (N7146, N7128);
or OR2 (N7147, N7145, N5737);
buf BUF1 (N7148, N7142);
xor XOR2 (N7149, N7143, N2799);
buf BUF1 (N7150, N7149);
xor XOR2 (N7151, N7146, N5303);
nand NAND2 (N7152, N7140, N4500);
nand NAND4 (N7153, N7130, N6754, N6596, N1879);
buf BUF1 (N7154, N7151);
xor XOR2 (N7155, N7150, N4984);
and AND3 (N7156, N7155, N1283, N2595);
nor NOR3 (N7157, N7147, N620, N1532);
nand NAND3 (N7158, N7122, N4572, N5220);
not NOT1 (N7159, N7141);
nand NAND4 (N7160, N7153, N6493, N309, N4569);
nand NAND2 (N7161, N7160, N630);
not NOT1 (N7162, N7159);
buf BUF1 (N7163, N7157);
nand NAND2 (N7164, N7152, N4321);
and AND4 (N7165, N7148, N5233, N6810, N3036);
not NOT1 (N7166, N7163);
xor XOR2 (N7167, N7162, N5272);
buf BUF1 (N7168, N7144);
or OR2 (N7169, N7165, N4647);
xor XOR2 (N7170, N7156, N5820);
not NOT1 (N7171, N7167);
xor XOR2 (N7172, N7136, N5750);
not NOT1 (N7173, N7164);
buf BUF1 (N7174, N7154);
nand NAND4 (N7175, N7169, N7145, N5619, N987);
nor NOR3 (N7176, N7170, N2775, N4487);
nand NAND3 (N7177, N7158, N5137, N3318);
and AND4 (N7178, N7175, N1991, N4457, N4321);
and AND3 (N7179, N7174, N1465, N2330);
buf BUF1 (N7180, N7177);
or OR4 (N7181, N7166, N2916, N2248, N112);
buf BUF1 (N7182, N7171);
xor XOR2 (N7183, N7178, N92);
nor NOR4 (N7184, N7161, N2804, N5575, N5758);
buf BUF1 (N7185, N7179);
nand NAND4 (N7186, N7168, N864, N3266, N3673);
and AND2 (N7187, N7181, N2966);
buf BUF1 (N7188, N7176);
xor XOR2 (N7189, N7184, N6311);
or OR4 (N7190, N7180, N1733, N3682, N1208);
nand NAND2 (N7191, N7187, N1365);
not NOT1 (N7192, N7191);
or OR3 (N7193, N7186, N915, N4295);
not NOT1 (N7194, N7189);
buf BUF1 (N7195, N7194);
not NOT1 (N7196, N7173);
buf BUF1 (N7197, N7188);
or OR3 (N7198, N7196, N5966, N5218);
buf BUF1 (N7199, N7197);
nand NAND4 (N7200, N7190, N6260, N2918, N359);
nand NAND2 (N7201, N7185, N1660);
buf BUF1 (N7202, N7199);
or OR4 (N7203, N7193, N6770, N2501, N4804);
xor XOR2 (N7204, N7202, N77);
buf BUF1 (N7205, N7198);
or OR4 (N7206, N7192, N4548, N6768, N4639);
not NOT1 (N7207, N7204);
not NOT1 (N7208, N7172);
and AND4 (N7209, N7195, N3607, N2522, N1541);
buf BUF1 (N7210, N7203);
nor NOR3 (N7211, N7207, N4616, N2506);
or OR2 (N7212, N7211, N3331);
nand NAND3 (N7213, N7205, N2029, N5130);
not NOT1 (N7214, N7213);
or OR4 (N7215, N7209, N5501, N3931, N5546);
nor NOR4 (N7216, N7212, N6412, N4358, N6467);
nand NAND2 (N7217, N7206, N2224);
and AND4 (N7218, N7210, N4512, N1928, N1533);
or OR4 (N7219, N7183, N1855, N4391, N6051);
nand NAND3 (N7220, N7208, N2942, N6690);
not NOT1 (N7221, N7218);
nand NAND3 (N7222, N7215, N4232, N3753);
or OR4 (N7223, N7222, N1951, N5858, N4299);
and AND3 (N7224, N7216, N6080, N1480);
buf BUF1 (N7225, N7217);
xor XOR2 (N7226, N7219, N5828);
xor XOR2 (N7227, N7225, N5481);
nand NAND4 (N7228, N7201, N794, N1924, N1635);
nor NOR2 (N7229, N7228, N5013);
buf BUF1 (N7230, N7220);
not NOT1 (N7231, N7229);
xor XOR2 (N7232, N7223, N871);
not NOT1 (N7233, N7231);
xor XOR2 (N7234, N7224, N6876);
and AND2 (N7235, N7230, N6658);
nor NOR4 (N7236, N7214, N6482, N4694, N4620);
and AND4 (N7237, N7232, N3584, N6036, N2307);
buf BUF1 (N7238, N7227);
nand NAND4 (N7239, N7182, N3178, N1247, N2389);
nand NAND2 (N7240, N7233, N5538);
or OR4 (N7241, N7239, N2323, N4345, N499);
xor XOR2 (N7242, N7234, N2858);
nand NAND3 (N7243, N7236, N854, N2002);
and AND2 (N7244, N7240, N2312);
or OR4 (N7245, N7200, N3425, N4141, N1715);
nor NOR2 (N7246, N7245, N4361);
nor NOR3 (N7247, N7242, N2780, N748);
and AND4 (N7248, N7246, N597, N108, N2550);
or OR2 (N7249, N7244, N3267);
buf BUF1 (N7250, N7235);
nor NOR4 (N7251, N7243, N4688, N2920, N6803);
or OR3 (N7252, N7250, N3032, N1107);
nand NAND2 (N7253, N7241, N5682);
and AND2 (N7254, N7247, N3650);
nor NOR3 (N7255, N7249, N3353, N2489);
buf BUF1 (N7256, N7221);
not NOT1 (N7257, N7238);
buf BUF1 (N7258, N7255);
buf BUF1 (N7259, N7237);
nor NOR3 (N7260, N7257, N1529, N5814);
nor NOR3 (N7261, N7259, N5332, N6468);
or OR3 (N7262, N7254, N2558, N1996);
not NOT1 (N7263, N7258);
buf BUF1 (N7264, N7263);
buf BUF1 (N7265, N7248);
and AND2 (N7266, N7226, N4220);
or OR3 (N7267, N7261, N3287, N1998);
nor NOR4 (N7268, N7256, N6582, N1911, N2770);
not NOT1 (N7269, N7264);
xor XOR2 (N7270, N7265, N1569);
or OR3 (N7271, N7251, N6612, N5083);
nor NOR4 (N7272, N7268, N2375, N6049, N2675);
nor NOR2 (N7273, N7262, N47);
and AND2 (N7274, N7269, N1131);
or OR2 (N7275, N7272, N5244);
or OR4 (N7276, N7266, N3487, N3527, N4156);
buf BUF1 (N7277, N7275);
buf BUF1 (N7278, N7271);
or OR3 (N7279, N7277, N6049, N4066);
and AND3 (N7280, N7276, N5855, N3875);
nand NAND2 (N7281, N7267, N2112);
and AND4 (N7282, N7281, N5040, N4712, N6816);
or OR4 (N7283, N7279, N6018, N6210, N3774);
buf BUF1 (N7284, N7253);
buf BUF1 (N7285, N7273);
nor NOR2 (N7286, N7282, N4176);
or OR2 (N7287, N7274, N4837);
nor NOR4 (N7288, N7286, N1754, N566, N6328);
not NOT1 (N7289, N7283);
not NOT1 (N7290, N7284);
nor NOR4 (N7291, N7280, N5719, N3084, N6244);
nand NAND4 (N7292, N7285, N4949, N772, N5418);
or OR4 (N7293, N7291, N879, N5551, N1892);
nand NAND2 (N7294, N7278, N3706);
nand NAND3 (N7295, N7292, N2991, N3383);
buf BUF1 (N7296, N7288);
nor NOR3 (N7297, N7289, N1815, N4222);
not NOT1 (N7298, N7295);
not NOT1 (N7299, N7294);
xor XOR2 (N7300, N7293, N1181);
and AND3 (N7301, N7296, N6234, N1804);
xor XOR2 (N7302, N7301, N966);
and AND4 (N7303, N7287, N1429, N145, N6663);
buf BUF1 (N7304, N7297);
xor XOR2 (N7305, N7298, N5448);
or OR3 (N7306, N7302, N5297, N201);
or OR2 (N7307, N7252, N3560);
buf BUF1 (N7308, N7304);
or OR2 (N7309, N7303, N5324);
or OR4 (N7310, N7299, N2539, N1961, N986);
xor XOR2 (N7311, N7305, N5492);
and AND3 (N7312, N7270, N6593, N5609);
and AND3 (N7313, N7300, N2908, N570);
buf BUF1 (N7314, N7306);
and AND3 (N7315, N7314, N3250, N542);
nand NAND2 (N7316, N7310, N5503);
or OR4 (N7317, N7307, N6682, N6685, N493);
buf BUF1 (N7318, N7260);
not NOT1 (N7319, N7308);
and AND2 (N7320, N7313, N5048);
xor XOR2 (N7321, N7316, N2027);
and AND3 (N7322, N7319, N1258, N5026);
xor XOR2 (N7323, N7322, N399);
or OR2 (N7324, N7321, N2220);
and AND3 (N7325, N7312, N2767, N2323);
and AND2 (N7326, N7320, N2338);
nand NAND4 (N7327, N7325, N5326, N1370, N3434);
not NOT1 (N7328, N7315);
or OR2 (N7329, N7326, N2846);
or OR4 (N7330, N7317, N6035, N4862, N1306);
or OR4 (N7331, N7323, N6860, N1284, N4478);
not NOT1 (N7332, N7309);
nand NAND4 (N7333, N7329, N4982, N6659, N3784);
nand NAND4 (N7334, N7311, N5870, N4870, N510);
nor NOR4 (N7335, N7330, N4913, N2627, N4970);
nand NAND3 (N7336, N7328, N6121, N1853);
xor XOR2 (N7337, N7290, N3515);
or OR3 (N7338, N7333, N6827, N5972);
xor XOR2 (N7339, N7332, N6001);
buf BUF1 (N7340, N7327);
buf BUF1 (N7341, N7336);
xor XOR2 (N7342, N7318, N7183);
or OR4 (N7343, N7340, N2276, N6720, N354);
nor NOR4 (N7344, N7341, N5623, N3722, N7263);
nor NOR4 (N7345, N7324, N983, N4766, N4285);
nor NOR4 (N7346, N7331, N4010, N2172, N3183);
nand NAND3 (N7347, N7343, N5847, N2717);
nand NAND3 (N7348, N7334, N5086, N1871);
and AND3 (N7349, N7344, N4812, N2072);
and AND2 (N7350, N7337, N6955);
nand NAND3 (N7351, N7339, N7135, N1745);
nor NOR3 (N7352, N7350, N4909, N5115);
or OR2 (N7353, N7351, N2224);
nor NOR3 (N7354, N7342, N5134, N2351);
xor XOR2 (N7355, N7345, N3242);
and AND3 (N7356, N7338, N1233, N6899);
nand NAND4 (N7357, N7348, N5077, N1090, N670);
xor XOR2 (N7358, N7357, N3089);
nand NAND4 (N7359, N7335, N1018, N6957, N4458);
xor XOR2 (N7360, N7354, N6962);
xor XOR2 (N7361, N7353, N6415);
and AND3 (N7362, N7360, N4842, N6420);
nor NOR3 (N7363, N7361, N3129, N4887);
not NOT1 (N7364, N7346);
nor NOR3 (N7365, N7352, N1395, N904);
not NOT1 (N7366, N7347);
xor XOR2 (N7367, N7358, N7220);
not NOT1 (N7368, N7364);
and AND2 (N7369, N7359, N4325);
nand NAND4 (N7370, N7355, N6184, N4217, N4808);
buf BUF1 (N7371, N7367);
buf BUF1 (N7372, N7368);
nand NAND2 (N7373, N7371, N522);
nor NOR3 (N7374, N7362, N5549, N5013);
and AND3 (N7375, N7366, N4568, N4746);
or OR2 (N7376, N7356, N4155);
not NOT1 (N7377, N7374);
and AND2 (N7378, N7369, N3733);
not NOT1 (N7379, N7365);
not NOT1 (N7380, N7373);
buf BUF1 (N7381, N7370);
or OR4 (N7382, N7379, N4360, N5640, N2457);
nand NAND2 (N7383, N7349, N4729);
and AND3 (N7384, N7377, N4353, N5967);
not NOT1 (N7385, N7381);
buf BUF1 (N7386, N7378);
buf BUF1 (N7387, N7375);
nor NOR3 (N7388, N7372, N7175, N1101);
or OR3 (N7389, N7382, N1433, N6797);
and AND3 (N7390, N7380, N4580, N6646);
nand NAND4 (N7391, N7384, N6980, N5870, N4213);
xor XOR2 (N7392, N7391, N773);
nor NOR3 (N7393, N7392, N2674, N3852);
not NOT1 (N7394, N7376);
xor XOR2 (N7395, N7394, N5972);
nand NAND2 (N7396, N7393, N5722);
buf BUF1 (N7397, N7387);
or OR3 (N7398, N7383, N7166, N6215);
xor XOR2 (N7399, N7397, N5744);
or OR2 (N7400, N7385, N6004);
nor NOR4 (N7401, N7389, N1581, N2253, N2132);
buf BUF1 (N7402, N7401);
not NOT1 (N7403, N7390);
not NOT1 (N7404, N7386);
or OR4 (N7405, N7396, N5825, N3615, N5195);
xor XOR2 (N7406, N7388, N2561);
and AND2 (N7407, N7406, N6353);
not NOT1 (N7408, N7404);
or OR2 (N7409, N7398, N1942);
not NOT1 (N7410, N7405);
xor XOR2 (N7411, N7402, N5529);
xor XOR2 (N7412, N7410, N6432);
nor NOR3 (N7413, N7395, N4694, N6461);
and AND2 (N7414, N7411, N6869);
xor XOR2 (N7415, N7407, N1434);
buf BUF1 (N7416, N7412);
xor XOR2 (N7417, N7399, N1172);
nand NAND3 (N7418, N7414, N1500, N2150);
xor XOR2 (N7419, N7363, N5625);
and AND2 (N7420, N7408, N814);
and AND3 (N7421, N7418, N7395, N6887);
nor NOR4 (N7422, N7419, N5048, N1917, N2015);
or OR3 (N7423, N7413, N5984, N4303);
xor XOR2 (N7424, N7423, N119);
buf BUF1 (N7425, N7415);
nor NOR2 (N7426, N7417, N5795);
buf BUF1 (N7427, N7403);
xor XOR2 (N7428, N7426, N2219);
not NOT1 (N7429, N7409);
xor XOR2 (N7430, N7400, N3010);
not NOT1 (N7431, N7428);
nor NOR3 (N7432, N7422, N7080, N6439);
not NOT1 (N7433, N7429);
nand NAND2 (N7434, N7424, N1689);
and AND3 (N7435, N7416, N2283, N1368);
nor NOR3 (N7436, N7427, N1452, N6112);
or OR2 (N7437, N7434, N2393);
and AND2 (N7438, N7435, N531);
buf BUF1 (N7439, N7420);
not NOT1 (N7440, N7421);
nor NOR2 (N7441, N7439, N1733);
nand NAND2 (N7442, N7436, N2685);
nand NAND4 (N7443, N7432, N4859, N2080, N3438);
nand NAND3 (N7444, N7430, N346, N3997);
or OR2 (N7445, N7425, N5818);
not NOT1 (N7446, N7431);
and AND2 (N7447, N7446, N1578);
xor XOR2 (N7448, N7433, N4436);
xor XOR2 (N7449, N7443, N1842);
buf BUF1 (N7450, N7448);
not NOT1 (N7451, N7440);
xor XOR2 (N7452, N7447, N704);
nand NAND4 (N7453, N7442, N7436, N4005, N514);
nor NOR2 (N7454, N7452, N6621);
nor NOR4 (N7455, N7451, N6618, N346, N5754);
xor XOR2 (N7456, N7445, N3312);
nor NOR2 (N7457, N7449, N4907);
not NOT1 (N7458, N7456);
buf BUF1 (N7459, N7450);
nor NOR3 (N7460, N7438, N472, N502);
buf BUF1 (N7461, N7460);
nor NOR2 (N7462, N7441, N4778);
or OR2 (N7463, N7455, N4355);
buf BUF1 (N7464, N7437);
or OR3 (N7465, N7458, N2672, N27);
nor NOR3 (N7466, N7459, N4086, N1821);
and AND3 (N7467, N7453, N5836, N449);
nor NOR4 (N7468, N7467, N6714, N1662, N2376);
xor XOR2 (N7469, N7462, N2667);
or OR4 (N7470, N7465, N944, N7134, N5135);
not NOT1 (N7471, N7468);
buf BUF1 (N7472, N7464);
buf BUF1 (N7473, N7470);
not NOT1 (N7474, N7472);
nand NAND3 (N7475, N7471, N5605, N1702);
and AND2 (N7476, N7473, N4577);
or OR2 (N7477, N7454, N722);
not NOT1 (N7478, N7469);
buf BUF1 (N7479, N7474);
xor XOR2 (N7480, N7479, N77);
xor XOR2 (N7481, N7457, N444);
not NOT1 (N7482, N7466);
not NOT1 (N7483, N7477);
not NOT1 (N7484, N7475);
nand NAND3 (N7485, N7484, N3107, N1246);
nand NAND3 (N7486, N7444, N2357, N7395);
buf BUF1 (N7487, N7476);
and AND3 (N7488, N7486, N5399, N2618);
or OR4 (N7489, N7482, N5458, N4989, N3251);
or OR3 (N7490, N7483, N7423, N6185);
nor NOR2 (N7491, N7487, N2122);
or OR2 (N7492, N7491, N1229);
not NOT1 (N7493, N7461);
xor XOR2 (N7494, N7485, N5548);
xor XOR2 (N7495, N7494, N6599);
not NOT1 (N7496, N7492);
not NOT1 (N7497, N7489);
and AND4 (N7498, N7463, N1189, N25, N2275);
xor XOR2 (N7499, N7488, N3114);
nor NOR2 (N7500, N7498, N7244);
nand NAND2 (N7501, N7495, N3560);
and AND4 (N7502, N7490, N4631, N5954, N79);
not NOT1 (N7503, N7499);
nand NAND4 (N7504, N7493, N7457, N4648, N416);
or OR4 (N7505, N7501, N7422, N329, N2561);
nand NAND4 (N7506, N7502, N62, N7486, N1064);
buf BUF1 (N7507, N7481);
and AND4 (N7508, N7478, N2118, N1128, N6353);
not NOT1 (N7509, N7507);
or OR4 (N7510, N7504, N5301, N550, N1863);
or OR3 (N7511, N7497, N7323, N3743);
nor NOR3 (N7512, N7480, N4674, N4644);
or OR3 (N7513, N7509, N397, N5909);
nand NAND4 (N7514, N7496, N4231, N6453, N6448);
or OR3 (N7515, N7508, N2876, N4813);
xor XOR2 (N7516, N7503, N4853);
not NOT1 (N7517, N7500);
or OR4 (N7518, N7514, N75, N3421, N6071);
nor NOR2 (N7519, N7515, N1528);
nand NAND4 (N7520, N7510, N5953, N3863, N426);
buf BUF1 (N7521, N7511);
xor XOR2 (N7522, N7517, N3867);
xor XOR2 (N7523, N7518, N3334);
buf BUF1 (N7524, N7513);
nand NAND4 (N7525, N7519, N5475, N2795, N7335);
buf BUF1 (N7526, N7525);
nor NOR2 (N7527, N7506, N3380);
xor XOR2 (N7528, N7520, N2860);
and AND2 (N7529, N7516, N2714);
nor NOR3 (N7530, N7523, N6331, N2477);
buf BUF1 (N7531, N7529);
and AND4 (N7532, N7521, N931, N4163, N7272);
nand NAND3 (N7533, N7512, N7048, N188);
nor NOR4 (N7534, N7531, N3594, N5079, N6104);
buf BUF1 (N7535, N7505);
not NOT1 (N7536, N7527);
not NOT1 (N7537, N7534);
buf BUF1 (N7538, N7526);
nand NAND4 (N7539, N7533, N4764, N3931, N6637);
nor NOR4 (N7540, N7528, N5794, N6159, N246);
and AND2 (N7541, N7540, N3316);
not NOT1 (N7542, N7524);
not NOT1 (N7543, N7537);
xor XOR2 (N7544, N7522, N817);
not NOT1 (N7545, N7541);
nor NOR3 (N7546, N7535, N4577, N6895);
not NOT1 (N7547, N7544);
xor XOR2 (N7548, N7542, N6281);
and AND2 (N7549, N7536, N5246);
buf BUF1 (N7550, N7530);
not NOT1 (N7551, N7549);
nor NOR4 (N7552, N7551, N937, N1522, N1752);
not NOT1 (N7553, N7547);
xor XOR2 (N7554, N7532, N5789);
xor XOR2 (N7555, N7550, N2644);
buf BUF1 (N7556, N7538);
xor XOR2 (N7557, N7556, N4619);
not NOT1 (N7558, N7552);
nand NAND3 (N7559, N7539, N1676, N4802);
nor NOR2 (N7560, N7558, N5169);
buf BUF1 (N7561, N7548);
not NOT1 (N7562, N7557);
xor XOR2 (N7563, N7559, N3847);
buf BUF1 (N7564, N7545);
or OR3 (N7565, N7543, N1169, N6382);
nand NAND2 (N7566, N7565, N6725);
buf BUF1 (N7567, N7555);
not NOT1 (N7568, N7564);
xor XOR2 (N7569, N7562, N7184);
not NOT1 (N7570, N7554);
buf BUF1 (N7571, N7553);
xor XOR2 (N7572, N7570, N4174);
not NOT1 (N7573, N7567);
buf BUF1 (N7574, N7560);
buf BUF1 (N7575, N7569);
nand NAND4 (N7576, N7561, N3350, N3106, N2517);
xor XOR2 (N7577, N7568, N2713);
nor NOR3 (N7578, N7573, N3428, N4450);
not NOT1 (N7579, N7571);
xor XOR2 (N7580, N7577, N3072);
nand NAND2 (N7581, N7580, N3272);
and AND3 (N7582, N7579, N3478, N6775);
and AND2 (N7583, N7575, N2470);
xor XOR2 (N7584, N7583, N2310);
and AND3 (N7585, N7582, N1789, N6789);
nor NOR4 (N7586, N7566, N135, N7041, N686);
xor XOR2 (N7587, N7546, N1553);
nand NAND2 (N7588, N7581, N1343);
and AND3 (N7589, N7585, N6088, N633);
buf BUF1 (N7590, N7587);
and AND2 (N7591, N7578, N3614);
nand NAND3 (N7592, N7574, N66, N1373);
or OR3 (N7593, N7563, N6774, N336);
nand NAND4 (N7594, N7591, N4288, N1875, N5845);
and AND4 (N7595, N7592, N5731, N1517, N4230);
nand NAND2 (N7596, N7584, N3863);
nand NAND2 (N7597, N7586, N2995);
nor NOR4 (N7598, N7596, N5193, N2924, N5049);
nand NAND2 (N7599, N7589, N2632);
nor NOR4 (N7600, N7588, N3823, N7158, N2871);
not NOT1 (N7601, N7595);
or OR3 (N7602, N7593, N2557, N2795);
not NOT1 (N7603, N7601);
and AND2 (N7604, N7590, N1719);
not NOT1 (N7605, N7594);
xor XOR2 (N7606, N7604, N5423);
nand NAND4 (N7607, N7576, N3858, N5953, N2700);
xor XOR2 (N7608, N7572, N1842);
and AND2 (N7609, N7602, N4846);
xor XOR2 (N7610, N7607, N5664);
and AND2 (N7611, N7605, N5202);
nand NAND4 (N7612, N7600, N3616, N3570, N4135);
nand NAND4 (N7613, N7598, N3102, N6077, N6401);
xor XOR2 (N7614, N7613, N4384);
not NOT1 (N7615, N7608);
buf BUF1 (N7616, N7610);
buf BUF1 (N7617, N7609);
buf BUF1 (N7618, N7614);
or OR2 (N7619, N7616, N5065);
nor NOR3 (N7620, N7606, N1600, N6806);
buf BUF1 (N7621, N7615);
or OR4 (N7622, N7599, N1874, N1750, N7044);
xor XOR2 (N7623, N7622, N502);
not NOT1 (N7624, N7619);
xor XOR2 (N7625, N7621, N3032);
nor NOR4 (N7626, N7624, N6064, N4694, N6157);
and AND3 (N7627, N7611, N6542, N754);
nor NOR4 (N7628, N7597, N4289, N292, N2160);
not NOT1 (N7629, N7617);
and AND2 (N7630, N7627, N4948);
xor XOR2 (N7631, N7618, N6771);
nand NAND4 (N7632, N7620, N2291, N2755, N6918);
or OR4 (N7633, N7612, N2207, N6258, N5685);
not NOT1 (N7634, N7632);
and AND2 (N7635, N7630, N2070);
or OR4 (N7636, N7629, N6081, N4071, N6619);
buf BUF1 (N7637, N7626);
xor XOR2 (N7638, N7634, N1367);
and AND2 (N7639, N7635, N3461);
buf BUF1 (N7640, N7637);
and AND3 (N7641, N7631, N734, N6050);
nor NOR2 (N7642, N7638, N5831);
buf BUF1 (N7643, N7639);
buf BUF1 (N7644, N7636);
and AND3 (N7645, N7643, N2467, N4069);
nand NAND4 (N7646, N7633, N884, N2403, N6620);
not NOT1 (N7647, N7641);
not NOT1 (N7648, N7645);
not NOT1 (N7649, N7628);
or OR2 (N7650, N7644, N6467);
or OR4 (N7651, N7640, N4482, N6751, N6207);
nor NOR2 (N7652, N7648, N6289);
buf BUF1 (N7653, N7649);
nand NAND2 (N7654, N7642, N2559);
or OR2 (N7655, N7651, N2551);
buf BUF1 (N7656, N7646);
nand NAND3 (N7657, N7603, N2324, N12);
nor NOR2 (N7658, N7655, N3198);
nand NAND2 (N7659, N7623, N2874);
buf BUF1 (N7660, N7656);
buf BUF1 (N7661, N7650);
or OR4 (N7662, N7647, N2954, N6331, N4448);
buf BUF1 (N7663, N7625);
and AND3 (N7664, N7658, N235, N5425);
or OR2 (N7665, N7661, N6355);
and AND3 (N7666, N7653, N1572, N7368);
nand NAND3 (N7667, N7654, N6111, N5319);
or OR2 (N7668, N7659, N3650);
or OR3 (N7669, N7660, N2927, N1670);
nand NAND4 (N7670, N7652, N2665, N6939, N2458);
buf BUF1 (N7671, N7663);
nand NAND4 (N7672, N7669, N7174, N4073, N1233);
or OR3 (N7673, N7672, N3209, N1380);
nor NOR2 (N7674, N7670, N1516);
not NOT1 (N7675, N7665);
or OR4 (N7676, N7666, N1957, N4454, N7047);
and AND4 (N7677, N7664, N4405, N7659, N55);
and AND3 (N7678, N7657, N4663, N1243);
nand NAND3 (N7679, N7662, N4396, N4204);
nor NOR2 (N7680, N7673, N3729);
xor XOR2 (N7681, N7667, N3810);
or OR4 (N7682, N7675, N2508, N944, N3993);
or OR4 (N7683, N7679, N7521, N6454, N6595);
xor XOR2 (N7684, N7677, N309);
or OR4 (N7685, N7684, N4632, N2863, N5364);
nor NOR3 (N7686, N7671, N5599, N1382);
xor XOR2 (N7687, N7681, N4598);
nand NAND4 (N7688, N7683, N5519, N3595, N252);
nor NOR2 (N7689, N7676, N665);
or OR2 (N7690, N7678, N5895);
or OR2 (N7691, N7685, N3155);
nor NOR2 (N7692, N7687, N4891);
xor XOR2 (N7693, N7674, N6649);
and AND4 (N7694, N7668, N3804, N3048, N1936);
or OR4 (N7695, N7689, N584, N2030, N4916);
not NOT1 (N7696, N7686);
nand NAND4 (N7697, N7692, N1389, N2417, N4049);
buf BUF1 (N7698, N7697);
not NOT1 (N7699, N7690);
not NOT1 (N7700, N7695);
and AND4 (N7701, N7691, N6102, N6208, N3851);
or OR4 (N7702, N7688, N7383, N1316, N2706);
nor NOR2 (N7703, N7702, N1482);
nor NOR3 (N7704, N7703, N2727, N2727);
xor XOR2 (N7705, N7682, N299);
and AND3 (N7706, N7700, N6890, N6513);
buf BUF1 (N7707, N7699);
nand NAND4 (N7708, N7693, N3743, N6490, N4999);
and AND3 (N7709, N7704, N2865, N1112);
or OR4 (N7710, N7696, N4230, N2387, N7466);
buf BUF1 (N7711, N7694);
and AND4 (N7712, N7707, N5086, N582, N7670);
nor NOR2 (N7713, N7710, N2284);
nor NOR4 (N7714, N7711, N3260, N940, N3703);
or OR4 (N7715, N7706, N4336, N2919, N6453);
nand NAND4 (N7716, N7713, N3524, N6923, N5780);
and AND2 (N7717, N7709, N170);
or OR3 (N7718, N7715, N2641, N5622);
xor XOR2 (N7719, N7698, N482);
buf BUF1 (N7720, N7717);
buf BUF1 (N7721, N7719);
and AND4 (N7722, N7712, N6749, N4397, N4363);
xor XOR2 (N7723, N7721, N3979);
and AND3 (N7724, N7723, N7539, N6537);
or OR4 (N7725, N7680, N2954, N7498, N394);
nor NOR3 (N7726, N7705, N6524, N3008);
buf BUF1 (N7727, N7708);
and AND4 (N7728, N7701, N3801, N6092, N4977);
and AND4 (N7729, N7725, N4257, N2454, N4739);
buf BUF1 (N7730, N7727);
not NOT1 (N7731, N7714);
and AND2 (N7732, N7718, N3137);
and AND2 (N7733, N7731, N2985);
not NOT1 (N7734, N7732);
and AND4 (N7735, N7729, N7650, N4339, N3853);
xor XOR2 (N7736, N7734, N3860);
not NOT1 (N7737, N7736);
buf BUF1 (N7738, N7726);
xor XOR2 (N7739, N7724, N1743);
buf BUF1 (N7740, N7730);
and AND2 (N7741, N7720, N537);
or OR2 (N7742, N7738, N6347);
not NOT1 (N7743, N7722);
or OR4 (N7744, N7728, N7373, N411, N2836);
nor NOR3 (N7745, N7741, N758, N833);
or OR4 (N7746, N7716, N5306, N2592, N7234);
not NOT1 (N7747, N7739);
buf BUF1 (N7748, N7735);
nor NOR3 (N7749, N7740, N3608, N5239);
and AND3 (N7750, N7737, N6850, N2196);
buf BUF1 (N7751, N7749);
xor XOR2 (N7752, N7750, N1678);
not NOT1 (N7753, N7751);
nand NAND2 (N7754, N7752, N5655);
nand NAND2 (N7755, N7753, N1217);
xor XOR2 (N7756, N7742, N3991);
xor XOR2 (N7757, N7744, N5618);
nand NAND2 (N7758, N7757, N2984);
not NOT1 (N7759, N7748);
or OR4 (N7760, N7747, N5143, N3996, N2864);
xor XOR2 (N7761, N7746, N7603);
and AND3 (N7762, N7756, N3365, N796);
or OR4 (N7763, N7743, N4035, N7508, N826);
buf BUF1 (N7764, N7745);
nand NAND3 (N7765, N7759, N4698, N5006);
and AND4 (N7766, N7764, N6700, N7685, N2525);
not NOT1 (N7767, N7755);
and AND2 (N7768, N7758, N2368);
and AND2 (N7769, N7754, N3697);
xor XOR2 (N7770, N7767, N806);
and AND4 (N7771, N7733, N4514, N2045, N2993);
buf BUF1 (N7772, N7769);
nand NAND4 (N7773, N7762, N6887, N615, N6288);
and AND3 (N7774, N7768, N7492, N2222);
nor NOR3 (N7775, N7763, N1705, N7559);
buf BUF1 (N7776, N7766);
nand NAND2 (N7777, N7772, N3222);
buf BUF1 (N7778, N7773);
buf BUF1 (N7779, N7776);
not NOT1 (N7780, N7761);
nand NAND4 (N7781, N7771, N5937, N3529, N5648);
and AND2 (N7782, N7780, N7653);
or OR2 (N7783, N7774, N3293);
buf BUF1 (N7784, N7778);
nand NAND2 (N7785, N7784, N6206);
nand NAND3 (N7786, N7760, N6211, N7653);
buf BUF1 (N7787, N7786);
not NOT1 (N7788, N7779);
and AND4 (N7789, N7775, N3030, N3821, N5731);
xor XOR2 (N7790, N7788, N1506);
buf BUF1 (N7791, N7781);
and AND3 (N7792, N7789, N1004, N5319);
not NOT1 (N7793, N7791);
buf BUF1 (N7794, N7765);
xor XOR2 (N7795, N7777, N5146);
nand NAND2 (N7796, N7785, N7535);
or OR3 (N7797, N7770, N5025, N1991);
xor XOR2 (N7798, N7783, N4580);
not NOT1 (N7799, N7795);
or OR4 (N7800, N7787, N7234, N7131, N5913);
not NOT1 (N7801, N7782);
buf BUF1 (N7802, N7796);
buf BUF1 (N7803, N7799);
xor XOR2 (N7804, N7797, N2906);
or OR4 (N7805, N7798, N6118, N2455, N6880);
or OR3 (N7806, N7793, N6177, N1380);
buf BUF1 (N7807, N7792);
buf BUF1 (N7808, N7804);
nand NAND4 (N7809, N7808, N6926, N329, N5797);
nor NOR3 (N7810, N7805, N7614, N4999);
or OR3 (N7811, N7807, N959, N1558);
buf BUF1 (N7812, N7803);
buf BUF1 (N7813, N7809);
and AND3 (N7814, N7813, N262, N856);
xor XOR2 (N7815, N7800, N6687);
xor XOR2 (N7816, N7794, N7070);
not NOT1 (N7817, N7790);
or OR3 (N7818, N7806, N243, N5091);
xor XOR2 (N7819, N7814, N5404);
or OR4 (N7820, N7818, N7726, N1618, N7704);
and AND3 (N7821, N7801, N683, N5659);
or OR3 (N7822, N7819, N2806, N388);
or OR4 (N7823, N7816, N7511, N3801, N2808);
nand NAND2 (N7824, N7812, N3927);
xor XOR2 (N7825, N7817, N7601);
buf BUF1 (N7826, N7802);
buf BUF1 (N7827, N7824);
nor NOR2 (N7828, N7825, N1241);
nand NAND3 (N7829, N7815, N7231, N1219);
and AND3 (N7830, N7821, N4420, N1732);
and AND2 (N7831, N7823, N3116);
or OR4 (N7832, N7828, N2121, N500, N7613);
or OR2 (N7833, N7822, N4081);
nor NOR3 (N7834, N7830, N6294, N3147);
nor NOR4 (N7835, N7827, N4535, N795, N6253);
buf BUF1 (N7836, N7810);
nand NAND4 (N7837, N7832, N6516, N3215, N905);
and AND2 (N7838, N7835, N5415);
buf BUF1 (N7839, N7829);
nor NOR2 (N7840, N7837, N1807);
xor XOR2 (N7841, N7840, N6891);
xor XOR2 (N7842, N7834, N7544);
not NOT1 (N7843, N7820);
nor NOR4 (N7844, N7842, N226, N2925, N5519);
buf BUF1 (N7845, N7839);
and AND3 (N7846, N7838, N674, N6155);
xor XOR2 (N7847, N7836, N3358);
xor XOR2 (N7848, N7845, N396);
or OR3 (N7849, N7848, N3332, N5528);
xor XOR2 (N7850, N7831, N1488);
xor XOR2 (N7851, N7850, N4029);
and AND2 (N7852, N7846, N7436);
or OR3 (N7853, N7851, N4753, N2745);
nand NAND3 (N7854, N7853, N2254, N7042);
not NOT1 (N7855, N7826);
nor NOR4 (N7856, N7854, N4956, N4124, N3682);
or OR2 (N7857, N7856, N1518);
and AND2 (N7858, N7855, N1547);
or OR2 (N7859, N7857, N4993);
and AND3 (N7860, N7859, N7463, N2191);
or OR4 (N7861, N7811, N4362, N6438, N3971);
not NOT1 (N7862, N7841);
xor XOR2 (N7863, N7852, N4681);
nand NAND4 (N7864, N7858, N3238, N4224, N6762);
or OR3 (N7865, N7863, N6384, N4312);
nor NOR3 (N7866, N7864, N5924, N4399);
buf BUF1 (N7867, N7843);
xor XOR2 (N7868, N7862, N1090);
xor XOR2 (N7869, N7849, N2846);
nor NOR2 (N7870, N7860, N7840);
buf BUF1 (N7871, N7870);
xor XOR2 (N7872, N7861, N4986);
and AND4 (N7873, N7865, N7327, N6669, N5786);
and AND3 (N7874, N7844, N390, N1553);
nand NAND4 (N7875, N7868, N737, N806, N1683);
nor NOR2 (N7876, N7833, N6057);
or OR2 (N7877, N7873, N5742);
and AND4 (N7878, N7869, N1037, N112, N958);
buf BUF1 (N7879, N7866);
or OR2 (N7880, N7867, N7642);
xor XOR2 (N7881, N7878, N2102);
and AND3 (N7882, N7847, N7807, N5391);
or OR3 (N7883, N7881, N5755, N831);
nand NAND4 (N7884, N7875, N4745, N6927, N5362);
buf BUF1 (N7885, N7880);
nand NAND4 (N7886, N7874, N7795, N7295, N3892);
or OR4 (N7887, N7879, N6554, N4255, N1983);
and AND3 (N7888, N7882, N3496, N6547);
buf BUF1 (N7889, N7887);
or OR3 (N7890, N7885, N2670, N7295);
buf BUF1 (N7891, N7890);
nor NOR2 (N7892, N7886, N1121);
and AND2 (N7893, N7876, N4979);
or OR3 (N7894, N7883, N6569, N4744);
nand NAND4 (N7895, N7872, N5497, N2506, N2129);
xor XOR2 (N7896, N7877, N5662);
xor XOR2 (N7897, N7893, N4432);
nand NAND4 (N7898, N7889, N7788, N2339, N5981);
xor XOR2 (N7899, N7898, N2204);
or OR4 (N7900, N7891, N790, N7171, N5602);
and AND4 (N7901, N7884, N1919, N4265, N614);
xor XOR2 (N7902, N7899, N2396);
or OR2 (N7903, N7871, N3678);
or OR4 (N7904, N7897, N7040, N5296, N1225);
or OR3 (N7905, N7888, N6693, N4414);
not NOT1 (N7906, N7894);
and AND3 (N7907, N7903, N2545, N4896);
or OR2 (N7908, N7900, N4470);
nor NOR3 (N7909, N7906, N3704, N2274);
xor XOR2 (N7910, N7908, N5126);
not NOT1 (N7911, N7909);
not NOT1 (N7912, N7902);
buf BUF1 (N7913, N7910);
or OR4 (N7914, N7892, N1658, N675, N5761);
or OR4 (N7915, N7905, N6962, N4276, N6283);
buf BUF1 (N7916, N7896);
buf BUF1 (N7917, N7916);
xor XOR2 (N7918, N7914, N7374);
not NOT1 (N7919, N7912);
and AND2 (N7920, N7918, N6983);
or OR4 (N7921, N7920, N122, N1048, N1429);
and AND4 (N7922, N7921, N1156, N7640, N4564);
nor NOR4 (N7923, N7901, N1530, N4721, N3087);
and AND3 (N7924, N7923, N3920, N3823);
nor NOR2 (N7925, N7917, N4034);
nor NOR2 (N7926, N7915, N670);
xor XOR2 (N7927, N7919, N130);
not NOT1 (N7928, N7907);
xor XOR2 (N7929, N7895, N2020);
or OR2 (N7930, N7904, N3980);
not NOT1 (N7931, N7927);
buf BUF1 (N7932, N7930);
nand NAND3 (N7933, N7913, N4280, N2114);
and AND4 (N7934, N7925, N166, N3129, N7313);
or OR2 (N7935, N7926, N5893);
not NOT1 (N7936, N7911);
nor NOR3 (N7937, N7922, N5321, N5925);
or OR4 (N7938, N7932, N5560, N1398, N2296);
and AND4 (N7939, N7924, N1177, N497, N96);
and AND3 (N7940, N7929, N6467, N3326);
nor NOR2 (N7941, N7928, N6053);
buf BUF1 (N7942, N7938);
or OR4 (N7943, N7939, N6916, N148, N4069);
nor NOR2 (N7944, N7943, N5792);
buf BUF1 (N7945, N7940);
xor XOR2 (N7946, N7934, N834);
nor NOR3 (N7947, N7936, N7933, N7309);
xor XOR2 (N7948, N3532, N329);
or OR2 (N7949, N7944, N3802);
xor XOR2 (N7950, N7941, N6851);
nand NAND4 (N7951, N7946, N3730, N3106, N4237);
or OR3 (N7952, N7937, N463, N6249);
not NOT1 (N7953, N7931);
and AND2 (N7954, N7952, N3512);
and AND4 (N7955, N7954, N938, N7583, N4353);
xor XOR2 (N7956, N7947, N4770);
or OR4 (N7957, N7956, N6088, N6050, N11);
xor XOR2 (N7958, N7953, N3927);
xor XOR2 (N7959, N7942, N3518);
nand NAND4 (N7960, N7958, N3611, N2140, N1954);
or OR3 (N7961, N7948, N954, N7313);
not NOT1 (N7962, N7955);
nand NAND2 (N7963, N7959, N6003);
and AND3 (N7964, N7950, N5633, N7528);
xor XOR2 (N7965, N7961, N5105);
or OR2 (N7966, N7965, N4922);
xor XOR2 (N7967, N7963, N5751);
xor XOR2 (N7968, N7945, N7492);
and AND2 (N7969, N7949, N3315);
buf BUF1 (N7970, N7969);
not NOT1 (N7971, N7935);
or OR3 (N7972, N7968, N1984, N1786);
nand NAND2 (N7973, N7971, N6904);
and AND3 (N7974, N7951, N7059, N2516);
nor NOR3 (N7975, N7964, N5858, N3212);
and AND3 (N7976, N7972, N6393, N3467);
nor NOR2 (N7977, N7962, N6998);
nand NAND2 (N7978, N7957, N2657);
buf BUF1 (N7979, N7970);
xor XOR2 (N7980, N7966, N97);
buf BUF1 (N7981, N7978);
buf BUF1 (N7982, N7975);
xor XOR2 (N7983, N7976, N5216);
not NOT1 (N7984, N7980);
nand NAND2 (N7985, N7974, N5613);
and AND2 (N7986, N7967, N5449);
nand NAND4 (N7987, N7960, N2993, N7147, N2939);
nand NAND3 (N7988, N7981, N6476, N6021);
or OR2 (N7989, N7986, N7260);
nor NOR4 (N7990, N7988, N7066, N6271, N4462);
nor NOR4 (N7991, N7987, N886, N4585, N354);
xor XOR2 (N7992, N7973, N5207);
and AND3 (N7993, N7989, N697, N3071);
not NOT1 (N7994, N7985);
and AND4 (N7995, N7992, N1091, N4441, N384);
nand NAND3 (N7996, N7994, N3852, N4011);
xor XOR2 (N7997, N7984, N7032);
nand NAND2 (N7998, N7995, N7608);
and AND2 (N7999, N7977, N3124);
and AND2 (N8000, N7999, N557);
or OR2 (N8001, N7991, N6485);
not NOT1 (N8002, N7990);
nand NAND2 (N8003, N7983, N2193);
xor XOR2 (N8004, N7996, N7930);
nor NOR3 (N8005, N7979, N7203, N7411);
nor NOR2 (N8006, N7993, N1916);
buf BUF1 (N8007, N8002);
xor XOR2 (N8008, N7997, N1453);
xor XOR2 (N8009, N8005, N2747);
or OR2 (N8010, N8001, N3899);
xor XOR2 (N8011, N8010, N1096);
not NOT1 (N8012, N8009);
buf BUF1 (N8013, N8000);
and AND3 (N8014, N7982, N2158, N6698);
nand NAND4 (N8015, N8013, N7151, N6454, N1525);
nand NAND2 (N8016, N7998, N6246);
buf BUF1 (N8017, N8012);
and AND2 (N8018, N8006, N2701);
nand NAND3 (N8019, N8017, N4055, N1272);
or OR2 (N8020, N8015, N5663);
not NOT1 (N8021, N8020);
nand NAND2 (N8022, N8021, N1093);
or OR2 (N8023, N8003, N3514);
or OR2 (N8024, N8014, N1907);
not NOT1 (N8025, N8004);
nor NOR4 (N8026, N8019, N7924, N1952, N686);
nor NOR3 (N8027, N8008, N1157, N6295);
nand NAND4 (N8028, N8016, N4127, N852, N7446);
buf BUF1 (N8029, N8011);
xor XOR2 (N8030, N8027, N5711);
xor XOR2 (N8031, N8007, N2761);
nand NAND2 (N8032, N8024, N6265);
xor XOR2 (N8033, N8031, N5653);
or OR4 (N8034, N8022, N5554, N47, N318);
xor XOR2 (N8035, N8034, N4059);
and AND3 (N8036, N8030, N629, N1624);
buf BUF1 (N8037, N8026);
buf BUF1 (N8038, N8023);
nand NAND4 (N8039, N8035, N4349, N2915, N5972);
nand NAND3 (N8040, N8033, N7835, N6298);
buf BUF1 (N8041, N8036);
nor NOR2 (N8042, N8040, N4923);
not NOT1 (N8043, N8025);
not NOT1 (N8044, N8018);
xor XOR2 (N8045, N8039, N1765);
and AND2 (N8046, N8037, N5161);
and AND3 (N8047, N8038, N7073, N767);
nor NOR4 (N8048, N8028, N7795, N3883, N4808);
xor XOR2 (N8049, N8041, N2123);
or OR2 (N8050, N8044, N527);
buf BUF1 (N8051, N8029);
nand NAND3 (N8052, N8050, N712, N4246);
nor NOR2 (N8053, N8048, N6635);
nand NAND3 (N8054, N8049, N5037, N6539);
not NOT1 (N8055, N8047);
nand NAND4 (N8056, N8042, N583, N656, N67);
or OR2 (N8057, N8053, N4317);
nand NAND4 (N8058, N8043, N1815, N5331, N1265);
nor NOR2 (N8059, N8052, N4413);
buf BUF1 (N8060, N8032);
nor NOR2 (N8061, N8057, N820);
nor NOR2 (N8062, N8054, N4372);
or OR3 (N8063, N8061, N4823, N6984);
and AND4 (N8064, N8051, N7892, N5942, N1211);
xor XOR2 (N8065, N8063, N3126);
buf BUF1 (N8066, N8056);
nor NOR2 (N8067, N8060, N3104);
or OR2 (N8068, N8046, N6859);
xor XOR2 (N8069, N8068, N6896);
xor XOR2 (N8070, N8062, N3574);
and AND4 (N8071, N8065, N7967, N3644, N6320);
nand NAND2 (N8072, N8066, N3695);
xor XOR2 (N8073, N8071, N7657);
and AND4 (N8074, N8059, N5240, N4166, N1205);
and AND3 (N8075, N8073, N6729, N7460);
not NOT1 (N8076, N8072);
and AND2 (N8077, N8045, N1560);
not NOT1 (N8078, N8070);
or OR3 (N8079, N8055, N6298, N4519);
or OR3 (N8080, N8077, N3338, N5208);
or OR2 (N8081, N8075, N7655);
xor XOR2 (N8082, N8067, N723);
buf BUF1 (N8083, N8078);
buf BUF1 (N8084, N8079);
and AND2 (N8085, N8064, N264);
buf BUF1 (N8086, N8069);
and AND4 (N8087, N8086, N1769, N4022, N7104);
and AND3 (N8088, N8083, N3941, N2600);
and AND4 (N8089, N8081, N6935, N7071, N3319);
nand NAND4 (N8090, N8089, N4420, N156, N7419);
buf BUF1 (N8091, N8074);
xor XOR2 (N8092, N8076, N7141);
xor XOR2 (N8093, N8084, N3137);
not NOT1 (N8094, N8088);
xor XOR2 (N8095, N8092, N2905);
not NOT1 (N8096, N8085);
or OR2 (N8097, N8096, N4441);
buf BUF1 (N8098, N8087);
or OR2 (N8099, N8058, N3496);
nand NAND3 (N8100, N8080, N1654, N6500);
xor XOR2 (N8101, N8093, N3326);
nand NAND2 (N8102, N8091, N3922);
not NOT1 (N8103, N8102);
and AND3 (N8104, N8103, N7985, N6602);
or OR4 (N8105, N8082, N1465, N3626, N2632);
nor NOR4 (N8106, N8095, N794, N2336, N4364);
and AND2 (N8107, N8104, N1877);
nand NAND2 (N8108, N8090, N4076);
and AND2 (N8109, N8106, N3848);
not NOT1 (N8110, N8105);
or OR4 (N8111, N8100, N7906, N6497, N3375);
or OR4 (N8112, N8094, N499, N7436, N7744);
xor XOR2 (N8113, N8112, N376);
nand NAND4 (N8114, N8098, N3311, N6017, N6984);
and AND4 (N8115, N8097, N7695, N5137, N7929);
and AND2 (N8116, N8113, N6076);
not NOT1 (N8117, N8116);
xor XOR2 (N8118, N8107, N3881);
nor NOR3 (N8119, N8109, N2583, N6444);
nor NOR4 (N8120, N8114, N3893, N3842, N2232);
or OR3 (N8121, N8101, N557, N7574);
not NOT1 (N8122, N8119);
nand NAND2 (N8123, N8115, N1329);
nor NOR2 (N8124, N8118, N4970);
xor XOR2 (N8125, N8108, N739);
and AND2 (N8126, N8125, N8103);
nand NAND4 (N8127, N8117, N3896, N7959, N3470);
or OR4 (N8128, N8111, N2994, N5210, N6103);
and AND3 (N8129, N8099, N3432, N4583);
and AND4 (N8130, N8129, N6839, N7581, N154);
or OR2 (N8131, N8123, N6907);
buf BUF1 (N8132, N8128);
xor XOR2 (N8133, N8122, N1830);
buf BUF1 (N8134, N8130);
buf BUF1 (N8135, N8131);
xor XOR2 (N8136, N8120, N2126);
and AND3 (N8137, N8134, N2019, N818);
not NOT1 (N8138, N8126);
xor XOR2 (N8139, N8127, N5270);
nor NOR2 (N8140, N8110, N5359);
and AND4 (N8141, N8138, N7991, N6711, N1636);
or OR2 (N8142, N8124, N5143);
buf BUF1 (N8143, N8133);
and AND3 (N8144, N8135, N7207, N4688);
nand NAND2 (N8145, N8121, N8090);
xor XOR2 (N8146, N8137, N2406);
buf BUF1 (N8147, N8144);
xor XOR2 (N8148, N8140, N8020);
xor XOR2 (N8149, N8136, N5965);
or OR3 (N8150, N8149, N1502, N8001);
or OR2 (N8151, N8146, N2359);
not NOT1 (N8152, N8142);
nor NOR2 (N8153, N8148, N8056);
buf BUF1 (N8154, N8153);
buf BUF1 (N8155, N8141);
nor NOR2 (N8156, N8139, N1608);
nor NOR2 (N8157, N8156, N279);
nand NAND2 (N8158, N8150, N6924);
or OR3 (N8159, N8147, N7692, N2913);
xor XOR2 (N8160, N8152, N6938);
not NOT1 (N8161, N8160);
nand NAND2 (N8162, N8143, N2973);
buf BUF1 (N8163, N8132);
and AND2 (N8164, N8145, N1693);
not NOT1 (N8165, N8157);
xor XOR2 (N8166, N8155, N4199);
not NOT1 (N8167, N8166);
buf BUF1 (N8168, N8162);
or OR4 (N8169, N8161, N7493, N6014, N2686);
not NOT1 (N8170, N8158);
xor XOR2 (N8171, N8167, N7611);
or OR2 (N8172, N8169, N3349);
and AND4 (N8173, N8163, N2098, N4237, N2069);
nor NOR3 (N8174, N8159, N4927, N5679);
not NOT1 (N8175, N8154);
nor NOR3 (N8176, N8173, N7784, N5822);
nand NAND3 (N8177, N8175, N5202, N7317);
nor NOR2 (N8178, N8171, N4532);
nand NAND2 (N8179, N8168, N4072);
not NOT1 (N8180, N8164);
and AND4 (N8181, N8179, N2188, N3234, N4702);
nor NOR3 (N8182, N8181, N1110, N6366);
or OR2 (N8183, N8170, N921);
xor XOR2 (N8184, N8165, N4902);
not NOT1 (N8185, N8184);
not NOT1 (N8186, N8185);
nor NOR3 (N8187, N8178, N2917, N5877);
buf BUF1 (N8188, N8187);
xor XOR2 (N8189, N8174, N3264);
nor NOR2 (N8190, N8183, N3682);
buf BUF1 (N8191, N8188);
or OR3 (N8192, N8151, N6497, N2121);
buf BUF1 (N8193, N8180);
nand NAND2 (N8194, N8193, N102);
nor NOR2 (N8195, N8176, N4812);
buf BUF1 (N8196, N8194);
or OR2 (N8197, N8177, N4503);
buf BUF1 (N8198, N8186);
or OR3 (N8199, N8192, N861, N1095);
xor XOR2 (N8200, N8199, N2355);
not NOT1 (N8201, N8198);
xor XOR2 (N8202, N8195, N1535);
nand NAND4 (N8203, N8172, N2744, N7236, N6008);
nand NAND4 (N8204, N8197, N2433, N7649, N2838);
or OR2 (N8205, N8196, N5750);
and AND4 (N8206, N8189, N3574, N79, N6663);
and AND3 (N8207, N8190, N837, N5984);
or OR3 (N8208, N8200, N2550, N5578);
nor NOR3 (N8209, N8203, N4884, N1859);
nor NOR4 (N8210, N8202, N1454, N8085, N171);
nor NOR3 (N8211, N8205, N1394, N2932);
or OR4 (N8212, N8211, N7976, N1297, N5301);
nand NAND3 (N8213, N8201, N7537, N3099);
nand NAND3 (N8214, N8204, N4486, N5253);
and AND4 (N8215, N8210, N7842, N4592, N7631);
and AND3 (N8216, N8206, N4698, N4618);
or OR3 (N8217, N8182, N2157, N3469);
or OR3 (N8218, N8208, N954, N5047);
nand NAND4 (N8219, N8213, N6000, N6356, N172);
buf BUF1 (N8220, N8218);
nor NOR4 (N8221, N8209, N7184, N5920, N5905);
nand NAND3 (N8222, N8220, N6368, N6176);
or OR2 (N8223, N8215, N3676);
nor NOR4 (N8224, N8212, N6210, N5231, N491);
buf BUF1 (N8225, N8219);
buf BUF1 (N8226, N8207);
not NOT1 (N8227, N8224);
nor NOR2 (N8228, N8222, N7528);
or OR4 (N8229, N8223, N659, N4848, N4530);
and AND4 (N8230, N8226, N1426, N3361, N7517);
and AND3 (N8231, N8227, N6583, N92);
nor NOR3 (N8232, N8214, N4310, N4388);
and AND3 (N8233, N8217, N2303, N2679);
buf BUF1 (N8234, N8225);
buf BUF1 (N8235, N8230);
and AND2 (N8236, N8232, N3880);
and AND2 (N8237, N8216, N3457);
not NOT1 (N8238, N8233);
and AND4 (N8239, N8236, N6834, N2893, N3045);
xor XOR2 (N8240, N8191, N3968);
and AND4 (N8241, N8238, N7332, N7672, N2515);
nand NAND4 (N8242, N8221, N7919, N2672, N8010);
not NOT1 (N8243, N8239);
or OR4 (N8244, N8235, N8168, N2068, N3382);
or OR4 (N8245, N8241, N8145, N1365, N1549);
nand NAND2 (N8246, N8228, N4407);
or OR3 (N8247, N8243, N5647, N4960);
xor XOR2 (N8248, N8237, N1726);
nand NAND2 (N8249, N8240, N6903);
and AND3 (N8250, N8246, N2742, N1464);
buf BUF1 (N8251, N8234);
or OR3 (N8252, N8242, N7978, N1479);
buf BUF1 (N8253, N8229);
nand NAND2 (N8254, N8253, N7416);
nand NAND3 (N8255, N8254, N3275, N6054);
buf BUF1 (N8256, N8248);
and AND3 (N8257, N8256, N6875, N2647);
xor XOR2 (N8258, N8252, N6685);
xor XOR2 (N8259, N8250, N3215);
not NOT1 (N8260, N8257);
nand NAND2 (N8261, N8251, N4646);
nor NOR2 (N8262, N8245, N3750);
and AND4 (N8263, N8259, N5975, N5429, N2331);
xor XOR2 (N8264, N8260, N3134);
not NOT1 (N8265, N8247);
not NOT1 (N8266, N8265);
buf BUF1 (N8267, N8249);
nor NOR4 (N8268, N8244, N4442, N6006, N3250);
xor XOR2 (N8269, N8263, N1884);
buf BUF1 (N8270, N8255);
buf BUF1 (N8271, N8269);
buf BUF1 (N8272, N8262);
and AND2 (N8273, N8231, N3732);
buf BUF1 (N8274, N8268);
xor XOR2 (N8275, N8258, N1465);
not NOT1 (N8276, N8264);
nand NAND3 (N8277, N8271, N720, N5084);
xor XOR2 (N8278, N8275, N6499);
buf BUF1 (N8279, N8273);
not NOT1 (N8280, N8274);
nor NOR2 (N8281, N8280, N6689);
not NOT1 (N8282, N8272);
xor XOR2 (N8283, N8267, N5369);
nand NAND3 (N8284, N8277, N1367, N5115);
buf BUF1 (N8285, N8278);
nand NAND2 (N8286, N8281, N7238);
or OR4 (N8287, N8261, N483, N6645, N2461);
nand NAND3 (N8288, N8286, N7262, N5425);
nor NOR2 (N8289, N8287, N1872);
nor NOR2 (N8290, N8266, N1953);
xor XOR2 (N8291, N8276, N4344);
not NOT1 (N8292, N8290);
nand NAND4 (N8293, N8285, N2870, N1450, N4976);
or OR3 (N8294, N8279, N7980, N1778);
xor XOR2 (N8295, N8292, N5075);
and AND4 (N8296, N8282, N8093, N3764, N955);
and AND3 (N8297, N8288, N3697, N7279);
nor NOR4 (N8298, N8294, N327, N2852, N3550);
buf BUF1 (N8299, N8270);
not NOT1 (N8300, N8284);
nor NOR4 (N8301, N8291, N5059, N3752, N2586);
buf BUF1 (N8302, N8300);
and AND4 (N8303, N8299, N1656, N5101, N579);
xor XOR2 (N8304, N8297, N5512);
or OR2 (N8305, N8304, N1360);
nand NAND2 (N8306, N8283, N5262);
or OR3 (N8307, N8289, N2751, N7363);
not NOT1 (N8308, N8305);
nor NOR4 (N8309, N8293, N1300, N5548, N638);
not NOT1 (N8310, N8301);
nand NAND2 (N8311, N8309, N4569);
buf BUF1 (N8312, N8311);
buf BUF1 (N8313, N8298);
nor NOR3 (N8314, N8312, N3917, N370);
nor NOR4 (N8315, N8303, N8281, N5028, N1400);
xor XOR2 (N8316, N8313, N1113);
or OR4 (N8317, N8316, N3920, N1843, N7483);
nor NOR2 (N8318, N8307, N161);
and AND4 (N8319, N8302, N7064, N6635, N2656);
nor NOR2 (N8320, N8308, N194);
not NOT1 (N8321, N8318);
not NOT1 (N8322, N8317);
nor NOR2 (N8323, N8315, N2880);
nor NOR3 (N8324, N8314, N5178, N6520);
xor XOR2 (N8325, N8320, N1154);
buf BUF1 (N8326, N8321);
nor NOR3 (N8327, N8326, N7855, N2651);
buf BUF1 (N8328, N8323);
or OR4 (N8329, N8306, N23, N5976, N8048);
and AND3 (N8330, N8329, N5579, N7439);
xor XOR2 (N8331, N8296, N3379);
and AND4 (N8332, N8330, N2388, N6374, N2886);
buf BUF1 (N8333, N8325);
nor NOR4 (N8334, N8322, N2044, N2246, N6760);
nor NOR2 (N8335, N8310, N6261);
not NOT1 (N8336, N8327);
nor NOR2 (N8337, N8332, N4531);
nand NAND3 (N8338, N8319, N7414, N7939);
and AND4 (N8339, N8336, N5080, N6264, N5887);
not NOT1 (N8340, N8337);
nor NOR3 (N8341, N8339, N700, N4172);
or OR3 (N8342, N8324, N560, N637);
buf BUF1 (N8343, N8295);
not NOT1 (N8344, N8335);
nand NAND3 (N8345, N8333, N7239, N4128);
nand NAND2 (N8346, N8342, N540);
nand NAND2 (N8347, N8346, N4509);
xor XOR2 (N8348, N8347, N7472);
buf BUF1 (N8349, N8338);
not NOT1 (N8350, N8343);
and AND3 (N8351, N8349, N3327, N2613);
nor NOR3 (N8352, N8334, N7791, N1412);
or OR4 (N8353, N8331, N5645, N7006, N1098);
xor XOR2 (N8354, N8341, N6339);
and AND2 (N8355, N8340, N6703);
nor NOR3 (N8356, N8355, N178, N1765);
nand NAND2 (N8357, N8356, N6985);
nor NOR3 (N8358, N8353, N6740, N2);
buf BUF1 (N8359, N8351);
nor NOR2 (N8360, N8358, N474);
and AND4 (N8361, N8357, N5184, N5248, N3979);
nor NOR3 (N8362, N8328, N5780, N3790);
not NOT1 (N8363, N8344);
nor NOR3 (N8364, N8348, N4580, N3091);
nand NAND4 (N8365, N8350, N6951, N8120, N3321);
and AND3 (N8366, N8364, N3180, N5737);
nor NOR4 (N8367, N8360, N6799, N6269, N7473);
and AND2 (N8368, N8363, N5440);
and AND2 (N8369, N8361, N6671);
nand NAND4 (N8370, N8368, N235, N1025, N5721);
buf BUF1 (N8371, N8354);
or OR4 (N8372, N8371, N5466, N7396, N5841);
buf BUF1 (N8373, N8370);
nor NOR3 (N8374, N8366, N2367, N8145);
and AND4 (N8375, N8359, N1653, N1560, N2734);
nor NOR3 (N8376, N8372, N1826, N7745);
buf BUF1 (N8377, N8352);
buf BUF1 (N8378, N8345);
nor NOR3 (N8379, N8362, N5465, N806);
not NOT1 (N8380, N8376);
xor XOR2 (N8381, N8374, N1634);
nand NAND4 (N8382, N8365, N3475, N3430, N1482);
nand NAND4 (N8383, N8379, N1997, N5145, N7272);
and AND4 (N8384, N8375, N475, N7104, N3117);
or OR4 (N8385, N8373, N7538, N751, N5566);
nor NOR3 (N8386, N8382, N7821, N1373);
xor XOR2 (N8387, N8367, N3848);
and AND4 (N8388, N8369, N5885, N2843, N6854);
nand NAND3 (N8389, N8381, N6482, N84);
or OR3 (N8390, N8388, N6164, N1596);
not NOT1 (N8391, N8383);
not NOT1 (N8392, N8390);
and AND4 (N8393, N8378, N2396, N7054, N2742);
nand NAND2 (N8394, N8386, N283);
xor XOR2 (N8395, N8393, N3823);
or OR3 (N8396, N8395, N2041, N5676);
nor NOR2 (N8397, N8384, N4796);
nand NAND3 (N8398, N8385, N2904, N3414);
buf BUF1 (N8399, N8392);
not NOT1 (N8400, N8398);
or OR4 (N8401, N8397, N8052, N942, N272);
nor NOR2 (N8402, N8401, N1833);
buf BUF1 (N8403, N8389);
xor XOR2 (N8404, N8377, N2528);
nand NAND4 (N8405, N8400, N7160, N4753, N851);
or OR3 (N8406, N8396, N2658, N7332);
or OR3 (N8407, N8391, N115, N8);
buf BUF1 (N8408, N8380);
and AND4 (N8409, N8408, N6577, N7080, N5410);
xor XOR2 (N8410, N8402, N5096);
or OR2 (N8411, N8410, N6360);
or OR2 (N8412, N8405, N2851);
not NOT1 (N8413, N8404);
and AND3 (N8414, N8406, N2907, N2833);
nand NAND2 (N8415, N8413, N4663);
not NOT1 (N8416, N8399);
nand NAND4 (N8417, N8412, N1663, N3509, N3085);
or OR4 (N8418, N8417, N7892, N4989, N5526);
or OR4 (N8419, N8387, N484, N2575, N6100);
and AND2 (N8420, N8407, N1205);
nor NOR2 (N8421, N8409, N5923);
nand NAND3 (N8422, N8403, N4033, N3908);
and AND3 (N8423, N8420, N679, N6066);
or OR3 (N8424, N8421, N5556, N8365);
buf BUF1 (N8425, N8416);
or OR4 (N8426, N8414, N2167, N6722, N1339);
and AND2 (N8427, N8415, N4659);
xor XOR2 (N8428, N8423, N225);
nor NOR3 (N8429, N8428, N5742, N5273);
and AND3 (N8430, N8422, N2123, N6161);
not NOT1 (N8431, N8394);
buf BUF1 (N8432, N8430);
or OR4 (N8433, N8419, N1585, N3491, N2652);
xor XOR2 (N8434, N8424, N692);
nand NAND4 (N8435, N8418, N6599, N8025, N1444);
not NOT1 (N8436, N8435);
nand NAND2 (N8437, N8434, N3264);
and AND4 (N8438, N8436, N2742, N1929, N3709);
buf BUF1 (N8439, N8433);
buf BUF1 (N8440, N8425);
not NOT1 (N8441, N8437);
or OR2 (N8442, N8426, N644);
or OR4 (N8443, N8441, N6580, N6642, N7626);
buf BUF1 (N8444, N8440);
and AND3 (N8445, N8431, N186, N30);
nand NAND4 (N8446, N8427, N694, N7637, N2537);
nand NAND2 (N8447, N8444, N140);
buf BUF1 (N8448, N8439);
nor NOR2 (N8449, N8429, N3025);
not NOT1 (N8450, N8443);
xor XOR2 (N8451, N8446, N7648);
nor NOR2 (N8452, N8449, N1709);
xor XOR2 (N8453, N8411, N5863);
and AND2 (N8454, N8442, N282);
nor NOR3 (N8455, N8445, N7628, N6763);
xor XOR2 (N8456, N8453, N4675);
and AND3 (N8457, N8455, N4647, N3339);
xor XOR2 (N8458, N8438, N478);
nand NAND3 (N8459, N8457, N7764, N2600);
buf BUF1 (N8460, N8447);
nor NOR3 (N8461, N8450, N6122, N3654);
xor XOR2 (N8462, N8448, N7761);
not NOT1 (N8463, N8456);
and AND3 (N8464, N8452, N3392, N7204);
or OR2 (N8465, N8451, N4662);
nor NOR3 (N8466, N8458, N1535, N4893);
xor XOR2 (N8467, N8459, N4426);
nand NAND3 (N8468, N8467, N4022, N6079);
not NOT1 (N8469, N8454);
and AND3 (N8470, N8465, N1861, N2879);
nor NOR3 (N8471, N8464, N3419, N1496);
nor NOR2 (N8472, N8463, N1162);
and AND2 (N8473, N8462, N4953);
or OR2 (N8474, N8466, N2014);
buf BUF1 (N8475, N8472);
nor NOR3 (N8476, N8474, N3373, N4129);
or OR3 (N8477, N8432, N6715, N2686);
or OR4 (N8478, N8473, N5478, N4372, N3465);
nor NOR4 (N8479, N8476, N7938, N7310, N2124);
nand NAND4 (N8480, N8468, N2308, N7995, N7701);
or OR4 (N8481, N8475, N1790, N6897, N3301);
buf BUF1 (N8482, N8481);
xor XOR2 (N8483, N8482, N516);
nand NAND4 (N8484, N8477, N7279, N7593, N612);
nor NOR2 (N8485, N8484, N376);
or OR3 (N8486, N8478, N6884, N8346);
and AND3 (N8487, N8485, N7591, N5823);
and AND4 (N8488, N8480, N4077, N3759, N2680);
xor XOR2 (N8489, N8470, N1605);
nor NOR4 (N8490, N8479, N6306, N2077, N2844);
nor NOR2 (N8491, N8469, N1142);
xor XOR2 (N8492, N8471, N4816);
nor NOR2 (N8493, N8489, N1142);
buf BUF1 (N8494, N8461);
nand NAND2 (N8495, N8492, N1713);
nor NOR3 (N8496, N8491, N929, N4993);
nor NOR3 (N8497, N8488, N6623, N3392);
nand NAND4 (N8498, N8483, N286, N3689, N2448);
nor NOR2 (N8499, N8460, N5000);
buf BUF1 (N8500, N8487);
or OR3 (N8501, N8493, N4065, N889);
xor XOR2 (N8502, N8486, N7435);
not NOT1 (N8503, N8498);
xor XOR2 (N8504, N8495, N4625);
or OR4 (N8505, N8502, N972, N6481, N1765);
or OR3 (N8506, N8499, N2787, N3593);
and AND2 (N8507, N8500, N1752);
xor XOR2 (N8508, N8505, N3794);
or OR4 (N8509, N8507, N248, N2825, N1805);
and AND2 (N8510, N8509, N3879);
nand NAND3 (N8511, N8506, N4351, N7620);
or OR3 (N8512, N8510, N7486, N1991);
xor XOR2 (N8513, N8504, N8301);
and AND2 (N8514, N8512, N4533);
not NOT1 (N8515, N8513);
and AND4 (N8516, N8511, N2768, N1, N3066);
xor XOR2 (N8517, N8514, N8373);
nor NOR4 (N8518, N8516, N878, N5383, N1954);
buf BUF1 (N8519, N8515);
not NOT1 (N8520, N8490);
nor NOR3 (N8521, N8518, N6499, N8486);
or OR2 (N8522, N8501, N8439);
nor NOR3 (N8523, N8520, N5354, N186);
not NOT1 (N8524, N8494);
and AND3 (N8525, N8517, N893, N7901);
not NOT1 (N8526, N8519);
nand NAND3 (N8527, N8525, N2979, N8091);
nor NOR2 (N8528, N8497, N2591);
nand NAND4 (N8529, N8522, N6398, N4627, N2585);
nand NAND4 (N8530, N8521, N4945, N3418, N550);
nor NOR3 (N8531, N8524, N6249, N1883);
nor NOR2 (N8532, N8530, N384);
xor XOR2 (N8533, N8532, N7929);
not NOT1 (N8534, N8503);
not NOT1 (N8535, N8531);
not NOT1 (N8536, N8523);
buf BUF1 (N8537, N8535);
or OR2 (N8538, N8526, N3744);
buf BUF1 (N8539, N8527);
nor NOR2 (N8540, N8536, N2037);
or OR4 (N8541, N8539, N1277, N6818, N1262);
nor NOR3 (N8542, N8508, N2446, N6440);
not NOT1 (N8543, N8542);
and AND4 (N8544, N8538, N5421, N7329, N6893);
and AND2 (N8545, N8543, N1076);
and AND3 (N8546, N8544, N2809, N3207);
nand NAND4 (N8547, N8533, N6906, N2119, N4879);
or OR3 (N8548, N8537, N2482, N6432);
nand NAND4 (N8549, N8496, N3926, N34, N2015);
not NOT1 (N8550, N8541);
buf BUF1 (N8551, N8546);
not NOT1 (N8552, N8534);
nand NAND3 (N8553, N8548, N7767, N4682);
buf BUF1 (N8554, N8550);
buf BUF1 (N8555, N8529);
xor XOR2 (N8556, N8528, N2045);
buf BUF1 (N8557, N8540);
nand NAND3 (N8558, N8549, N3681, N8012);
not NOT1 (N8559, N8552);
or OR3 (N8560, N8556, N4444, N6525);
or OR2 (N8561, N8545, N2186);
or OR2 (N8562, N8553, N5277);
nor NOR2 (N8563, N8561, N6379);
or OR2 (N8564, N8555, N8067);
or OR4 (N8565, N8563, N3965, N3916, N8457);
nor NOR3 (N8566, N8551, N113, N4162);
nand NAND3 (N8567, N8557, N7499, N1934);
and AND4 (N8568, N8559, N1694, N903, N7337);
or OR2 (N8569, N8558, N2224);
nor NOR3 (N8570, N8566, N4717, N6937);
and AND4 (N8571, N8568, N2793, N3037, N4658);
and AND2 (N8572, N8565, N5433);
nor NOR4 (N8573, N8554, N2925, N4771, N453);
and AND2 (N8574, N8569, N509);
nor NOR2 (N8575, N8570, N3995);
xor XOR2 (N8576, N8574, N5926);
or OR3 (N8577, N8576, N7444, N6826);
xor XOR2 (N8578, N8572, N3586);
not NOT1 (N8579, N8577);
and AND4 (N8580, N8578, N2451, N7517, N7387);
or OR4 (N8581, N8571, N5131, N5673, N692);
or OR4 (N8582, N8581, N8067, N4985, N3086);
buf BUF1 (N8583, N8580);
buf BUF1 (N8584, N8579);
xor XOR2 (N8585, N8562, N2295);
nand NAND3 (N8586, N8547, N7761, N6635);
buf BUF1 (N8587, N8586);
xor XOR2 (N8588, N8585, N5179);
not NOT1 (N8589, N8564);
xor XOR2 (N8590, N8588, N7476);
nand NAND2 (N8591, N8575, N2880);
and AND3 (N8592, N8560, N1687, N8168);
nor NOR3 (N8593, N8591, N4272, N923);
buf BUF1 (N8594, N8573);
or OR2 (N8595, N8584, N8327);
not NOT1 (N8596, N8590);
nor NOR4 (N8597, N8594, N8057, N3124, N7935);
nor NOR2 (N8598, N8582, N7054);
buf BUF1 (N8599, N8567);
nand NAND2 (N8600, N8593, N2514);
and AND3 (N8601, N8598, N2660, N6181);
nand NAND3 (N8602, N8595, N3233, N521);
nor NOR4 (N8603, N8600, N2296, N2646, N772);
not NOT1 (N8604, N8592);
xor XOR2 (N8605, N8589, N328);
nor NOR4 (N8606, N8596, N4182, N5854, N790);
nand NAND4 (N8607, N8606, N7677, N906, N7285);
nor NOR2 (N8608, N8583, N1343);
not NOT1 (N8609, N8602);
or OR4 (N8610, N8608, N4376, N8397, N6263);
xor XOR2 (N8611, N8601, N55);
not NOT1 (N8612, N8599);
nand NAND3 (N8613, N8604, N7826, N4556);
not NOT1 (N8614, N8612);
nand NAND2 (N8615, N8603, N4011);
or OR2 (N8616, N8609, N5287);
buf BUF1 (N8617, N8605);
xor XOR2 (N8618, N8610, N1568);
nand NAND4 (N8619, N8613, N8541, N3935, N2075);
not NOT1 (N8620, N8617);
not NOT1 (N8621, N8618);
nor NOR3 (N8622, N8611, N2692, N4969);
buf BUF1 (N8623, N8616);
or OR2 (N8624, N8597, N6451);
nand NAND2 (N8625, N8587, N1811);
and AND2 (N8626, N8623, N2293);
or OR3 (N8627, N8607, N4913, N7458);
and AND4 (N8628, N8622, N4417, N2823, N5927);
nor NOR3 (N8629, N8625, N6346, N1507);
xor XOR2 (N8630, N8615, N4940);
nand NAND3 (N8631, N8624, N6337, N4341);
or OR3 (N8632, N8630, N450, N1145);
buf BUF1 (N8633, N8632);
and AND3 (N8634, N8633, N5646, N5482);
xor XOR2 (N8635, N8634, N7609);
not NOT1 (N8636, N8614);
buf BUF1 (N8637, N8629);
not NOT1 (N8638, N8626);
xor XOR2 (N8639, N8619, N6451);
not NOT1 (N8640, N8628);
xor XOR2 (N8641, N8631, N3847);
nand NAND4 (N8642, N8641, N2907, N6020, N6634);
buf BUF1 (N8643, N8621);
buf BUF1 (N8644, N8639);
nor NOR2 (N8645, N8642, N4160);
nor NOR4 (N8646, N8635, N7197, N6038, N808);
nor NOR2 (N8647, N8646, N3388);
buf BUF1 (N8648, N8620);
or OR2 (N8649, N8643, N7162);
or OR4 (N8650, N8627, N4957, N6548, N5920);
nand NAND2 (N8651, N8644, N6642);
nor NOR4 (N8652, N8650, N4003, N7619, N7836);
and AND2 (N8653, N8640, N7299);
nand NAND2 (N8654, N8637, N5734);
not NOT1 (N8655, N8653);
buf BUF1 (N8656, N8645);
xor XOR2 (N8657, N8652, N75);
or OR3 (N8658, N8647, N2001, N3941);
nand NAND2 (N8659, N8655, N2664);
or OR3 (N8660, N8658, N3336, N5151);
and AND3 (N8661, N8654, N2725, N5149);
and AND3 (N8662, N8649, N4387, N5003);
and AND4 (N8663, N8638, N1117, N2714, N889);
xor XOR2 (N8664, N8656, N5402);
or OR4 (N8665, N8663, N990, N7736, N203);
buf BUF1 (N8666, N8661);
and AND3 (N8667, N8659, N970, N438);
not NOT1 (N8668, N8666);
buf BUF1 (N8669, N8667);
nand NAND3 (N8670, N8669, N3405, N2740);
xor XOR2 (N8671, N8657, N7764);
nor NOR4 (N8672, N8662, N3500, N7133, N6602);
nand NAND3 (N8673, N8648, N6635, N8014);
not NOT1 (N8674, N8636);
and AND4 (N8675, N8671, N6477, N3556, N6291);
buf BUF1 (N8676, N8670);
nand NAND4 (N8677, N8668, N4935, N1377, N3730);
xor XOR2 (N8678, N8672, N2256);
nand NAND3 (N8679, N8678, N5586, N7343);
nand NAND2 (N8680, N8676, N4812);
or OR4 (N8681, N8677, N796, N1904, N6695);
nor NOR2 (N8682, N8673, N6504);
buf BUF1 (N8683, N8675);
and AND3 (N8684, N8682, N1249, N5841);
or OR3 (N8685, N8651, N6252, N5734);
nand NAND3 (N8686, N8683, N6205, N6836);
buf BUF1 (N8687, N8679);
or OR4 (N8688, N8686, N7397, N8183, N2695);
buf BUF1 (N8689, N8681);
and AND4 (N8690, N8664, N7652, N853, N4507);
not NOT1 (N8691, N8687);
buf BUF1 (N8692, N8685);
nand NAND2 (N8693, N8665, N3906);
nand NAND3 (N8694, N8690, N4112, N7872);
nor NOR3 (N8695, N8691, N4982, N5330);
xor XOR2 (N8696, N8680, N2041);
not NOT1 (N8697, N8674);
not NOT1 (N8698, N8684);
not NOT1 (N8699, N8697);
xor XOR2 (N8700, N8699, N4071);
buf BUF1 (N8701, N8688);
xor XOR2 (N8702, N8689, N3244);
xor XOR2 (N8703, N8700, N4305);
nand NAND2 (N8704, N8693, N1158);
nand NAND3 (N8705, N8695, N2867, N6647);
not NOT1 (N8706, N8701);
buf BUF1 (N8707, N8704);
nand NAND3 (N8708, N8692, N6093, N3832);
buf BUF1 (N8709, N8707);
and AND2 (N8710, N8696, N6293);
xor XOR2 (N8711, N8660, N2923);
not NOT1 (N8712, N8702);
xor XOR2 (N8713, N8698, N5761);
and AND3 (N8714, N8713, N3567, N3867);
not NOT1 (N8715, N8711);
or OR3 (N8716, N8714, N2606, N5501);
nor NOR2 (N8717, N8716, N5980);
nand NAND4 (N8718, N8710, N3358, N6801, N4281);
not NOT1 (N8719, N8703);
buf BUF1 (N8720, N8718);
or OR4 (N8721, N8719, N6278, N478, N506);
xor XOR2 (N8722, N8706, N570);
nand NAND3 (N8723, N8694, N8712, N762);
xor XOR2 (N8724, N1942, N275);
nand NAND4 (N8725, N8708, N6218, N4752, N5829);
or OR2 (N8726, N8717, N4196);
nand NAND3 (N8727, N8725, N6671, N6069);
not NOT1 (N8728, N8720);
xor XOR2 (N8729, N8709, N4479);
not NOT1 (N8730, N8722);
buf BUF1 (N8731, N8721);
and AND2 (N8732, N8705, N1512);
nand NAND4 (N8733, N8729, N883, N3804, N416);
xor XOR2 (N8734, N8715, N4438);
not NOT1 (N8735, N8732);
xor XOR2 (N8736, N8724, N6667);
nand NAND2 (N8737, N8735, N8543);
or OR4 (N8738, N8726, N8188, N1164, N7570);
buf BUF1 (N8739, N8723);
xor XOR2 (N8740, N8728, N3425);
buf BUF1 (N8741, N8740);
buf BUF1 (N8742, N8737);
nand NAND4 (N8743, N8736, N5967, N6352, N2086);
nor NOR3 (N8744, N8742, N1637, N7372);
nand NAND4 (N8745, N8730, N2605, N1125, N7492);
not NOT1 (N8746, N8745);
xor XOR2 (N8747, N8741, N3116);
buf BUF1 (N8748, N8743);
nand NAND3 (N8749, N8748, N3004, N8263);
buf BUF1 (N8750, N8733);
or OR4 (N8751, N8749, N7859, N3065, N3281);
nand NAND2 (N8752, N8746, N2795);
and AND4 (N8753, N8727, N5828, N5039, N8568);
nand NAND2 (N8754, N8751, N878);
not NOT1 (N8755, N8747);
nand NAND4 (N8756, N8731, N6731, N7929, N3262);
and AND2 (N8757, N8756, N2575);
or OR4 (N8758, N8750, N2163, N2096, N5921);
nor NOR4 (N8759, N8744, N3861, N1475, N5582);
buf BUF1 (N8760, N8757);
buf BUF1 (N8761, N8753);
nor NOR4 (N8762, N8759, N7028, N7636, N2134);
and AND4 (N8763, N8758, N7284, N5308, N7218);
or OR2 (N8764, N8739, N309);
and AND2 (N8765, N8752, N8154);
nand NAND2 (N8766, N8761, N2883);
nor NOR3 (N8767, N8755, N81, N7338);
nor NOR2 (N8768, N8760, N7749);
or OR2 (N8769, N8767, N5342);
buf BUF1 (N8770, N8763);
and AND3 (N8771, N8765, N7227, N7209);
or OR2 (N8772, N8766, N6641);
and AND2 (N8773, N8769, N7371);
nor NOR4 (N8774, N8770, N3153, N211, N7009);
xor XOR2 (N8775, N8738, N8500);
and AND2 (N8776, N8775, N2109);
xor XOR2 (N8777, N8764, N7877);
nor NOR4 (N8778, N8762, N4347, N1987, N1491);
nand NAND4 (N8779, N8734, N8662, N4931, N3603);
or OR2 (N8780, N8768, N1900);
nor NOR2 (N8781, N8772, N19);
or OR2 (N8782, N8754, N757);
not NOT1 (N8783, N8774);
nor NOR2 (N8784, N8781, N177);
nor NOR3 (N8785, N8779, N5414, N924);
nand NAND2 (N8786, N8780, N3050);
xor XOR2 (N8787, N8782, N849);
not NOT1 (N8788, N8787);
not NOT1 (N8789, N8784);
xor XOR2 (N8790, N8785, N7238);
xor XOR2 (N8791, N8788, N1411);
or OR2 (N8792, N8776, N7136);
nor NOR3 (N8793, N8771, N6255, N5761);
buf BUF1 (N8794, N8778);
not NOT1 (N8795, N8789);
or OR2 (N8796, N8792, N506);
or OR4 (N8797, N8794, N6581, N7556, N1972);
xor XOR2 (N8798, N8786, N3080);
nand NAND4 (N8799, N8783, N8377, N5912, N270);
and AND3 (N8800, N8798, N4790, N8059);
or OR3 (N8801, N8795, N6161, N1195);
and AND3 (N8802, N8777, N6621, N822);
or OR2 (N8803, N8796, N6789);
xor XOR2 (N8804, N8799, N5939);
not NOT1 (N8805, N8773);
nor NOR3 (N8806, N8791, N5035, N7616);
nand NAND4 (N8807, N8801, N8007, N94, N8449);
and AND4 (N8808, N8793, N6774, N7509, N5861);
or OR2 (N8809, N8808, N4496);
nand NAND4 (N8810, N8797, N6239, N7295, N4989);
or OR4 (N8811, N8804, N2913, N8280, N4062);
xor XOR2 (N8812, N8811, N1708);
xor XOR2 (N8813, N8800, N3840);
buf BUF1 (N8814, N8813);
xor XOR2 (N8815, N8802, N3595);
and AND3 (N8816, N8790, N8145, N5606);
nand NAND3 (N8817, N8814, N1820, N4459);
or OR3 (N8818, N8805, N7631, N1670);
nor NOR2 (N8819, N8815, N6932);
xor XOR2 (N8820, N8803, N2903);
buf BUF1 (N8821, N8818);
or OR2 (N8822, N8812, N4150);
nor NOR4 (N8823, N8819, N7063, N3471, N7884);
xor XOR2 (N8824, N8806, N2088);
nand NAND2 (N8825, N8821, N4809);
nor NOR2 (N8826, N8823, N8028);
and AND3 (N8827, N8826, N217, N8694);
and AND4 (N8828, N8817, N8718, N6145, N1879);
xor XOR2 (N8829, N8809, N4159);
xor XOR2 (N8830, N8807, N267);
or OR2 (N8831, N8828, N1737);
nand NAND2 (N8832, N8825, N710);
xor XOR2 (N8833, N8820, N4642);
and AND3 (N8834, N8832, N6256, N7536);
nor NOR2 (N8835, N8829, N3092);
not NOT1 (N8836, N8831);
and AND2 (N8837, N8816, N188);
xor XOR2 (N8838, N8824, N2609);
or OR4 (N8839, N8830, N3180, N6094, N7033);
not NOT1 (N8840, N8839);
nand NAND4 (N8841, N8840, N2189, N7147, N4797);
buf BUF1 (N8842, N8838);
not NOT1 (N8843, N8834);
or OR3 (N8844, N8835, N1901, N6505);
nor NOR2 (N8845, N8842, N5108);
xor XOR2 (N8846, N8836, N5712);
nor NOR4 (N8847, N8837, N222, N3905, N2068);
or OR2 (N8848, N8841, N3697);
buf BUF1 (N8849, N8822);
and AND4 (N8850, N8849, N3939, N6999, N3029);
xor XOR2 (N8851, N8848, N1298);
not NOT1 (N8852, N8850);
buf BUF1 (N8853, N8833);
and AND3 (N8854, N8827, N2424, N110);
nor NOR3 (N8855, N8847, N7665, N5483);
xor XOR2 (N8856, N8846, N7875);
nand NAND4 (N8857, N8856, N304, N1546, N1018);
nor NOR4 (N8858, N8845, N8407, N4393, N8500);
nand NAND2 (N8859, N8810, N6750);
and AND4 (N8860, N8859, N5679, N3681, N7731);
buf BUF1 (N8861, N8860);
not NOT1 (N8862, N8861);
nor NOR2 (N8863, N8851, N8118);
nand NAND4 (N8864, N8844, N1350, N375, N4129);
and AND3 (N8865, N8862, N5843, N254);
nand NAND3 (N8866, N8855, N3734, N3826);
nor NOR3 (N8867, N8863, N4436, N3653);
not NOT1 (N8868, N8866);
and AND3 (N8869, N8843, N608, N2915);
xor XOR2 (N8870, N8865, N8365);
or OR4 (N8871, N8869, N7267, N6717, N1716);
buf BUF1 (N8872, N8871);
and AND4 (N8873, N8857, N1804, N749, N7535);
and AND2 (N8874, N8867, N853);
nand NAND4 (N8875, N8858, N6052, N8841, N4502);
nand NAND2 (N8876, N8854, N3072);
nor NOR4 (N8877, N8852, N7913, N6584, N8875);
nand NAND4 (N8878, N1631, N734, N1365, N325);
buf BUF1 (N8879, N8877);
and AND2 (N8880, N8853, N5116);
and AND4 (N8881, N8878, N6619, N935, N7359);
or OR2 (N8882, N8864, N8524);
xor XOR2 (N8883, N8879, N1179);
or OR2 (N8884, N8868, N3712);
buf BUF1 (N8885, N8876);
buf BUF1 (N8886, N8870);
nor NOR2 (N8887, N8884, N1410);
nor NOR3 (N8888, N8872, N3820, N631);
nand NAND2 (N8889, N8883, N7039);
nor NOR4 (N8890, N8889, N6780, N7237, N1481);
nand NAND3 (N8891, N8885, N5308, N4808);
nor NOR4 (N8892, N8881, N2977, N557, N3413);
nor NOR3 (N8893, N8890, N5430, N562);
xor XOR2 (N8894, N8887, N6653);
xor XOR2 (N8895, N8892, N8737);
not NOT1 (N8896, N8882);
xor XOR2 (N8897, N8896, N4123);
nand NAND2 (N8898, N8874, N3920);
and AND2 (N8899, N8886, N4416);
nor NOR2 (N8900, N8873, N1596);
buf BUF1 (N8901, N8894);
not NOT1 (N8902, N8897);
buf BUF1 (N8903, N8895);
nor NOR3 (N8904, N8900, N3777, N2937);
xor XOR2 (N8905, N8891, N2689);
and AND2 (N8906, N8905, N7768);
buf BUF1 (N8907, N8888);
or OR2 (N8908, N8880, N5646);
not NOT1 (N8909, N8893);
and AND4 (N8910, N8909, N2692, N4971, N1553);
nand NAND2 (N8911, N8904, N3826);
nand NAND2 (N8912, N8906, N8652);
nor NOR3 (N8913, N8899, N6687, N3301);
buf BUF1 (N8914, N8913);
not NOT1 (N8915, N8914);
nand NAND3 (N8916, N8911, N3664, N2602);
not NOT1 (N8917, N8910);
xor XOR2 (N8918, N8898, N4429);
xor XOR2 (N8919, N8903, N5300);
buf BUF1 (N8920, N8916);
not NOT1 (N8921, N8918);
and AND3 (N8922, N8901, N4929, N3665);
and AND3 (N8923, N8917, N6929, N522);
nor NOR2 (N8924, N8919, N6652);
nor NOR3 (N8925, N8902, N3501, N8366);
xor XOR2 (N8926, N8923, N2058);
nand NAND4 (N8927, N8926, N173, N3183, N4641);
or OR3 (N8928, N8920, N3985, N931);
xor XOR2 (N8929, N8907, N1607);
xor XOR2 (N8930, N8915, N8670);
or OR3 (N8931, N8912, N1025, N7054);
or OR4 (N8932, N8931, N6632, N8215, N2992);
or OR3 (N8933, N8925, N2915, N1893);
nand NAND2 (N8934, N8908, N6640);
not NOT1 (N8935, N8921);
not NOT1 (N8936, N8922);
nor NOR4 (N8937, N8930, N8075, N5382, N2217);
nor NOR4 (N8938, N8934, N1058, N553, N2445);
nand NAND4 (N8939, N8935, N6079, N7907, N597);
nand NAND3 (N8940, N8927, N8042, N3880);
or OR2 (N8941, N8932, N6114);
xor XOR2 (N8942, N8940, N794);
nand NAND4 (N8943, N8937, N6205, N775, N3976);
or OR4 (N8944, N8943, N3249, N1043, N5167);
xor XOR2 (N8945, N8941, N8909);
buf BUF1 (N8946, N8928);
nor NOR2 (N8947, N8945, N4391);
or OR2 (N8948, N8933, N2233);
nor NOR4 (N8949, N8924, N98, N6142, N3986);
buf BUF1 (N8950, N8949);
nand NAND3 (N8951, N8950, N6347, N5868);
not NOT1 (N8952, N8946);
nor NOR4 (N8953, N8944, N1567, N7169, N4936);
buf BUF1 (N8954, N8953);
nand NAND4 (N8955, N8942, N3167, N7499, N8554);
or OR4 (N8956, N8948, N7144, N4443, N8891);
xor XOR2 (N8957, N8947, N5803);
or OR2 (N8958, N8957, N5001);
buf BUF1 (N8959, N8952);
buf BUF1 (N8960, N8956);
nor NOR3 (N8961, N8938, N7765, N2211);
xor XOR2 (N8962, N8960, N1101);
nand NAND4 (N8963, N8939, N202, N4221, N7013);
xor XOR2 (N8964, N8961, N7424);
not NOT1 (N8965, N8955);
buf BUF1 (N8966, N8954);
xor XOR2 (N8967, N8959, N7738);
not NOT1 (N8968, N8958);
nand NAND2 (N8969, N8966, N3929);
nand NAND2 (N8970, N8967, N2345);
not NOT1 (N8971, N8963);
not NOT1 (N8972, N8971);
not NOT1 (N8973, N8970);
xor XOR2 (N8974, N8962, N7901);
not NOT1 (N8975, N8974);
or OR2 (N8976, N8964, N799);
xor XOR2 (N8977, N8965, N636);
buf BUF1 (N8978, N8936);
nor NOR4 (N8979, N8951, N7705, N4898, N8824);
or OR3 (N8980, N8929, N1995, N2612);
not NOT1 (N8981, N8977);
and AND3 (N8982, N8976, N6547, N8181);
xor XOR2 (N8983, N8979, N4709);
xor XOR2 (N8984, N8980, N7598);
and AND3 (N8985, N8968, N7173, N2408);
nand NAND4 (N8986, N8973, N3869, N4660, N5909);
and AND2 (N8987, N8972, N8253);
not NOT1 (N8988, N8983);
xor XOR2 (N8989, N8975, N6210);
nor NOR3 (N8990, N8988, N5458, N6164);
nand NAND2 (N8991, N8990, N6073);
nand NAND2 (N8992, N8981, N6595);
nand NAND3 (N8993, N8991, N1912, N7145);
nand NAND4 (N8994, N8992, N4935, N331, N2621);
nor NOR2 (N8995, N8986, N203);
xor XOR2 (N8996, N8978, N4928);
and AND2 (N8997, N8994, N6108);
nor NOR4 (N8998, N8969, N8228, N999, N7038);
and AND4 (N8999, N8996, N6917, N8859, N2846);
buf BUF1 (N9000, N8993);
buf BUF1 (N9001, N8997);
and AND3 (N9002, N9000, N2805, N8691);
xor XOR2 (N9003, N8999, N1760);
nand NAND4 (N9004, N8989, N5249, N3894, N6499);
or OR4 (N9005, N9004, N3839, N6925, N8728);
nand NAND2 (N9006, N8998, N206);
nand NAND2 (N9007, N8982, N6773);
not NOT1 (N9008, N9003);
buf BUF1 (N9009, N8987);
xor XOR2 (N9010, N8995, N7592);
buf BUF1 (N9011, N9002);
xor XOR2 (N9012, N9010, N8270);
xor XOR2 (N9013, N8985, N2828);
nand NAND3 (N9014, N8984, N2664, N5294);
not NOT1 (N9015, N9001);
nand NAND4 (N9016, N9011, N8057, N878, N6474);
and AND2 (N9017, N9005, N1153);
or OR4 (N9018, N9012, N6247, N732, N4069);
not NOT1 (N9019, N9018);
and AND2 (N9020, N9019, N930);
and AND2 (N9021, N9016, N5643);
nor NOR3 (N9022, N9009, N2648, N2671);
nor NOR4 (N9023, N9021, N2156, N6905, N7322);
and AND3 (N9024, N9023, N1585, N3835);
not NOT1 (N9025, N9022);
or OR3 (N9026, N9024, N2389, N8134);
nor NOR4 (N9027, N9017, N8047, N7339, N989);
buf BUF1 (N9028, N9008);
buf BUF1 (N9029, N9014);
and AND3 (N9030, N9025, N3971, N6140);
and AND4 (N9031, N9026, N1082, N4440, N2957);
not NOT1 (N9032, N9015);
and AND4 (N9033, N9028, N4509, N4046, N3898);
and AND2 (N9034, N9030, N8946);
nor NOR2 (N9035, N9020, N664);
nor NOR3 (N9036, N9027, N6466, N1713);
nor NOR3 (N9037, N9033, N4928, N496);
xor XOR2 (N9038, N9029, N3411);
xor XOR2 (N9039, N9031, N2419);
xor XOR2 (N9040, N9006, N8055);
or OR2 (N9041, N9037, N1266);
not NOT1 (N9042, N9035);
or OR3 (N9043, N9038, N2371, N1716);
and AND3 (N9044, N9007, N3985, N7637);
and AND3 (N9045, N9044, N8219, N4823);
xor XOR2 (N9046, N9045, N4771);
xor XOR2 (N9047, N9032, N8897);
or OR4 (N9048, N9043, N2195, N1312, N4455);
nand NAND4 (N9049, N9042, N8613, N198, N3922);
or OR4 (N9050, N9039, N5023, N8832, N4357);
nor NOR3 (N9051, N9036, N4097, N943);
or OR2 (N9052, N9046, N4153);
not NOT1 (N9053, N9050);
not NOT1 (N9054, N9041);
xor XOR2 (N9055, N9049, N6064);
xor XOR2 (N9056, N9013, N7157);
nand NAND3 (N9057, N9040, N6690, N61);
and AND2 (N9058, N9048, N5443);
nor NOR4 (N9059, N9051, N9017, N1731, N5438);
not NOT1 (N9060, N9047);
nand NAND2 (N9061, N9034, N1057);
and AND4 (N9062, N9056, N8950, N7012, N56);
nor NOR4 (N9063, N9061, N4336, N853, N5727);
or OR3 (N9064, N9053, N6353, N2195);
nand NAND3 (N9065, N9058, N6985, N872);
and AND4 (N9066, N9064, N4327, N3145, N7201);
not NOT1 (N9067, N9062);
and AND4 (N9068, N9063, N6057, N1980, N1049);
not NOT1 (N9069, N9060);
xor XOR2 (N9070, N9069, N645);
or OR2 (N9071, N9059, N344);
or OR2 (N9072, N9052, N8939);
and AND3 (N9073, N9070, N2725, N6563);
nand NAND3 (N9074, N9067, N2664, N3022);
buf BUF1 (N9075, N9066);
not NOT1 (N9076, N9075);
xor XOR2 (N9077, N9073, N2003);
or OR2 (N9078, N9054, N2003);
nor NOR2 (N9079, N9068, N5846);
nand NAND3 (N9080, N9076, N3754, N5081);
or OR4 (N9081, N9080, N2511, N7810, N7927);
xor XOR2 (N9082, N9077, N209);
buf BUF1 (N9083, N9057);
xor XOR2 (N9084, N9079, N7082);
and AND2 (N9085, N9082, N7105);
or OR2 (N9086, N9078, N6681);
buf BUF1 (N9087, N9071);
and AND4 (N9088, N9087, N2859, N1869, N2586);
nand NAND4 (N9089, N9065, N1761, N6163, N1093);
xor XOR2 (N9090, N9088, N7704);
buf BUF1 (N9091, N9086);
nand NAND4 (N9092, N9089, N8012, N5440, N3967);
buf BUF1 (N9093, N9091);
nand NAND2 (N9094, N9072, N5524);
buf BUF1 (N9095, N9084);
nand NAND4 (N9096, N9090, N6396, N7786, N1762);
buf BUF1 (N9097, N9074);
xor XOR2 (N9098, N9093, N8909);
or OR4 (N9099, N9098, N4974, N8088, N8697);
and AND3 (N9100, N9085, N6649, N5750);
nand NAND2 (N9101, N9081, N5973);
or OR4 (N9102, N9095, N2947, N2897, N4907);
nand NAND3 (N9103, N9096, N2810, N1973);
and AND4 (N9104, N9103, N4291, N1086, N2581);
nor NOR4 (N9105, N9083, N7990, N7178, N4863);
or OR4 (N9106, N9100, N119, N6302, N2911);
or OR2 (N9107, N9105, N342);
nand NAND4 (N9108, N9102, N5530, N5460, N8191);
buf BUF1 (N9109, N9107);
nand NAND4 (N9110, N9094, N6721, N7025, N3901);
nor NOR4 (N9111, N9109, N1662, N8654, N11);
nor NOR3 (N9112, N9055, N2473, N685);
or OR2 (N9113, N9092, N5802);
nor NOR4 (N9114, N9112, N2815, N8673, N7163);
and AND4 (N9115, N9101, N5037, N4169, N2293);
buf BUF1 (N9116, N9114);
nor NOR4 (N9117, N9113, N7104, N2533, N1315);
xor XOR2 (N9118, N9097, N4157);
or OR4 (N9119, N9115, N2250, N8379, N5782);
nand NAND2 (N9120, N9118, N238);
nand NAND4 (N9121, N9120, N418, N8308, N5159);
nand NAND4 (N9122, N9116, N69, N8054, N3415);
not NOT1 (N9123, N9121);
xor XOR2 (N9124, N9110, N6331);
not NOT1 (N9125, N9124);
or OR2 (N9126, N9119, N6943);
not NOT1 (N9127, N9108);
or OR4 (N9128, N9104, N59, N1131, N4982);
not NOT1 (N9129, N9123);
not NOT1 (N9130, N9129);
nand NAND2 (N9131, N9130, N7405);
xor XOR2 (N9132, N9131, N3732);
nor NOR2 (N9133, N9132, N1516);
and AND4 (N9134, N9099, N8352, N5912, N8345);
buf BUF1 (N9135, N9126);
not NOT1 (N9136, N9117);
and AND3 (N9137, N9125, N2913, N3431);
xor XOR2 (N9138, N9134, N3755);
or OR3 (N9139, N9136, N6406, N4800);
nand NAND2 (N9140, N9111, N5861);
and AND4 (N9141, N9133, N1599, N1272, N6025);
nor NOR4 (N9142, N9139, N794, N644, N8245);
nor NOR4 (N9143, N9128, N4558, N631, N177);
buf BUF1 (N9144, N9142);
or OR3 (N9145, N9141, N7631, N7624);
and AND4 (N9146, N9140, N8001, N6358, N634);
and AND3 (N9147, N9143, N6130, N871);
xor XOR2 (N9148, N9135, N2735);
or OR4 (N9149, N9146, N155, N8286, N1294);
or OR2 (N9150, N9144, N525);
xor XOR2 (N9151, N9127, N1114);
or OR4 (N9152, N9106, N9053, N8348, N3454);
xor XOR2 (N9153, N9147, N4354);
and AND2 (N9154, N9149, N8368);
nor NOR3 (N9155, N9153, N5736, N2619);
nand NAND2 (N9156, N9151, N3936);
buf BUF1 (N9157, N9152);
xor XOR2 (N9158, N9122, N6755);
or OR2 (N9159, N9158, N3310);
and AND3 (N9160, N9150, N4966, N6759);
or OR3 (N9161, N9160, N2513, N4169);
nand NAND4 (N9162, N9145, N2647, N985, N23);
nand NAND4 (N9163, N9157, N6727, N2325, N8712);
nand NAND4 (N9164, N9156, N4356, N8631, N5331);
not NOT1 (N9165, N9161);
not NOT1 (N9166, N9159);
buf BUF1 (N9167, N9166);
or OR3 (N9168, N9167, N458, N6671);
nor NOR4 (N9169, N9148, N787, N4362, N6127);
or OR3 (N9170, N9168, N6275, N3932);
not NOT1 (N9171, N9154);
nand NAND2 (N9172, N9163, N3979);
nand NAND2 (N9173, N9172, N384);
buf BUF1 (N9174, N9169);
and AND2 (N9175, N9138, N6984);
or OR3 (N9176, N9137, N695, N369);
buf BUF1 (N9177, N9165);
nand NAND3 (N9178, N9162, N932, N2245);
or OR4 (N9179, N9171, N8691, N1638, N7247);
nand NAND4 (N9180, N9164, N2777, N845, N4549);
nor NOR3 (N9181, N9173, N7008, N9034);
not NOT1 (N9182, N9180);
buf BUF1 (N9183, N9177);
xor XOR2 (N9184, N9155, N6728);
nand NAND4 (N9185, N9175, N4623, N2274, N2260);
buf BUF1 (N9186, N9185);
not NOT1 (N9187, N9181);
nor NOR4 (N9188, N9174, N274, N7603, N5812);
and AND2 (N9189, N9186, N1898);
xor XOR2 (N9190, N9176, N3916);
nor NOR4 (N9191, N9187, N7678, N8908, N7340);
and AND4 (N9192, N9170, N7742, N2345, N6564);
and AND2 (N9193, N9179, N7289);
xor XOR2 (N9194, N9183, N2968);
and AND4 (N9195, N9184, N726, N4304, N111);
nand NAND3 (N9196, N9193, N897, N2474);
nor NOR4 (N9197, N9194, N4779, N3483, N8002);
nor NOR2 (N9198, N9191, N7084);
xor XOR2 (N9199, N9197, N8519);
xor XOR2 (N9200, N9182, N6855);
buf BUF1 (N9201, N9190);
xor XOR2 (N9202, N9196, N3863);
buf BUF1 (N9203, N9192);
or OR4 (N9204, N9202, N7691, N4395, N750);
not NOT1 (N9205, N9198);
and AND2 (N9206, N9188, N4540);
buf BUF1 (N9207, N9201);
xor XOR2 (N9208, N9207, N1296);
nand NAND3 (N9209, N9203, N3100, N6131);
nand NAND4 (N9210, N9200, N7072, N2759, N8530);
or OR2 (N9211, N9189, N6409);
xor XOR2 (N9212, N9195, N2666);
nand NAND3 (N9213, N9206, N8113, N6722);
xor XOR2 (N9214, N9209, N8355);
nor NOR2 (N9215, N9208, N7364);
buf BUF1 (N9216, N9213);
or OR3 (N9217, N9178, N6619, N8190);
nand NAND4 (N9218, N9204, N5664, N8649, N2194);
nand NAND3 (N9219, N9214, N4245, N8567);
and AND2 (N9220, N9212, N2887);
buf BUF1 (N9221, N9215);
xor XOR2 (N9222, N9205, N9121);
not NOT1 (N9223, N9211);
nor NOR2 (N9224, N9222, N5730);
or OR2 (N9225, N9217, N6341);
and AND3 (N9226, N9199, N4406, N4091);
xor XOR2 (N9227, N9221, N1313);
not NOT1 (N9228, N9210);
not NOT1 (N9229, N9226);
nand NAND4 (N9230, N9223, N6829, N8055, N4424);
nand NAND2 (N9231, N9228, N8764);
xor XOR2 (N9232, N9216, N1853);
nand NAND3 (N9233, N9220, N5507, N9193);
not NOT1 (N9234, N9233);
and AND3 (N9235, N9224, N5330, N7324);
and AND3 (N9236, N9225, N8754, N7341);
and AND2 (N9237, N9231, N8317);
or OR4 (N9238, N9236, N3114, N3343, N1930);
xor XOR2 (N9239, N9235, N3987);
and AND3 (N9240, N9234, N8479, N6649);
or OR3 (N9241, N9219, N7151, N1629);
nor NOR3 (N9242, N9239, N1536, N8405);
buf BUF1 (N9243, N9229);
buf BUF1 (N9244, N9227);
nor NOR2 (N9245, N9232, N6870);
buf BUF1 (N9246, N9218);
and AND4 (N9247, N9230, N2298, N3189, N3890);
not NOT1 (N9248, N9238);
not NOT1 (N9249, N9243);
not NOT1 (N9250, N9244);
xor XOR2 (N9251, N9248, N7623);
buf BUF1 (N9252, N9245);
nand NAND2 (N9253, N9241, N1012);
nor NOR2 (N9254, N9237, N4904);
or OR2 (N9255, N9242, N1880);
nor NOR3 (N9256, N9254, N7976, N2635);
nor NOR2 (N9257, N9252, N3632);
xor XOR2 (N9258, N9249, N8670);
nand NAND4 (N9259, N9256, N2848, N4179, N7309);
buf BUF1 (N9260, N9251);
not NOT1 (N9261, N9257);
xor XOR2 (N9262, N9247, N7674);
and AND3 (N9263, N9246, N6552, N4483);
nor NOR3 (N9264, N9259, N9141, N6240);
or OR2 (N9265, N9240, N8318);
xor XOR2 (N9266, N9260, N7139);
buf BUF1 (N9267, N9250);
xor XOR2 (N9268, N9253, N8056);
or OR4 (N9269, N9266, N3020, N1642, N1291);
or OR2 (N9270, N9258, N7345);
xor XOR2 (N9271, N9262, N9060);
buf BUF1 (N9272, N9267);
or OR3 (N9273, N9261, N5771, N4694);
and AND2 (N9274, N9255, N7337);
buf BUF1 (N9275, N9270);
nand NAND3 (N9276, N9275, N2762, N8181);
not NOT1 (N9277, N9264);
buf BUF1 (N9278, N9263);
not NOT1 (N9279, N9277);
buf BUF1 (N9280, N9279);
nand NAND4 (N9281, N9272, N1545, N2944, N2137);
and AND4 (N9282, N9274, N3487, N6937, N5657);
not NOT1 (N9283, N9265);
xor XOR2 (N9284, N9269, N1069);
buf BUF1 (N9285, N9268);
nor NOR2 (N9286, N9271, N549);
nor NOR4 (N9287, N9276, N3404, N1798, N4214);
not NOT1 (N9288, N9284);
buf BUF1 (N9289, N9286);
nand NAND3 (N9290, N9289, N6119, N8989);
buf BUF1 (N9291, N9288);
nor NOR4 (N9292, N9285, N6670, N2918, N7895);
or OR3 (N9293, N9290, N4678, N4447);
nand NAND3 (N9294, N9287, N8768, N5690);
nand NAND4 (N9295, N9283, N2285, N559, N4);
or OR4 (N9296, N9273, N1520, N4918, N7004);
not NOT1 (N9297, N9281);
or OR2 (N9298, N9296, N813);
nand NAND3 (N9299, N9293, N2515, N655);
nand NAND4 (N9300, N9278, N6075, N6058, N952);
not NOT1 (N9301, N9297);
or OR4 (N9302, N9292, N823, N5245, N5457);
nand NAND4 (N9303, N9295, N1486, N6677, N1906);
not NOT1 (N9304, N9294);
nand NAND3 (N9305, N9300, N577, N2732);
and AND3 (N9306, N9302, N1043, N5866);
and AND3 (N9307, N9282, N9172, N7859);
nor NOR2 (N9308, N9301, N9162);
and AND2 (N9309, N9291, N7495);
not NOT1 (N9310, N9303);
and AND4 (N9311, N9310, N6678, N6739, N8612);
and AND2 (N9312, N9280, N6026);
not NOT1 (N9313, N9309);
buf BUF1 (N9314, N9312);
and AND3 (N9315, N9314, N2305, N5574);
not NOT1 (N9316, N9307);
buf BUF1 (N9317, N9304);
and AND3 (N9318, N9317, N2170, N4079);
nand NAND4 (N9319, N9316, N631, N4489, N2944);
and AND3 (N9320, N9298, N5619, N2382);
nor NOR3 (N9321, N9308, N2941, N2393);
or OR3 (N9322, N9299, N5262, N6153);
nor NOR4 (N9323, N9306, N1594, N6252, N6971);
xor XOR2 (N9324, N9323, N8514);
or OR3 (N9325, N9320, N2595, N6990);
nand NAND2 (N9326, N9318, N5900);
xor XOR2 (N9327, N9322, N4534);
nor NOR4 (N9328, N9315, N5425, N9247, N6211);
or OR4 (N9329, N9328, N635, N8547, N6266);
buf BUF1 (N9330, N9326);
or OR2 (N9331, N9325, N5094);
not NOT1 (N9332, N9329);
xor XOR2 (N9333, N9305, N8847);
and AND3 (N9334, N9327, N5763, N4046);
not NOT1 (N9335, N9324);
or OR4 (N9336, N9333, N6200, N8824, N662);
xor XOR2 (N9337, N9331, N7381);
buf BUF1 (N9338, N9337);
xor XOR2 (N9339, N9319, N722);
and AND2 (N9340, N9338, N6287);
xor XOR2 (N9341, N9334, N1074);
nor NOR2 (N9342, N9321, N9122);
nand NAND2 (N9343, N9336, N8053);
not NOT1 (N9344, N9343);
xor XOR2 (N9345, N9335, N1665);
and AND2 (N9346, N9341, N3654);
nor NOR3 (N9347, N9313, N1656, N106);
nor NOR4 (N9348, N9342, N4435, N6736, N657);
nor NOR3 (N9349, N9347, N7467, N7341);
not NOT1 (N9350, N9330);
xor XOR2 (N9351, N9340, N6101);
or OR4 (N9352, N9344, N28, N8476, N6597);
or OR3 (N9353, N9311, N8604, N9314);
or OR4 (N9354, N9349, N2233, N5221, N6971);
or OR4 (N9355, N9345, N1369, N7724, N2849);
and AND3 (N9356, N9352, N8678, N2331);
nand NAND2 (N9357, N9332, N8823);
and AND3 (N9358, N9351, N297, N970);
buf BUF1 (N9359, N9354);
xor XOR2 (N9360, N9346, N3322);
and AND2 (N9361, N9358, N7966);
or OR4 (N9362, N9361, N8301, N3916, N4760);
nor NOR3 (N9363, N9339, N6250, N7009);
not NOT1 (N9364, N9363);
nor NOR3 (N9365, N9360, N4745, N345);
xor XOR2 (N9366, N9350, N6363);
not NOT1 (N9367, N9353);
and AND3 (N9368, N9365, N1310, N648);
xor XOR2 (N9369, N9366, N7093);
and AND2 (N9370, N9357, N6834);
xor XOR2 (N9371, N9355, N7440);
or OR3 (N9372, N9364, N7671, N3986);
nand NAND2 (N9373, N9367, N7068);
not NOT1 (N9374, N9362);
xor XOR2 (N9375, N9373, N779);
not NOT1 (N9376, N9368);
not NOT1 (N9377, N9370);
buf BUF1 (N9378, N9369);
and AND2 (N9379, N9378, N1463);
nor NOR3 (N9380, N9379, N8560, N1136);
and AND4 (N9381, N9377, N5216, N2630, N4756);
xor XOR2 (N9382, N9372, N1476);
nand NAND2 (N9383, N9380, N2969);
nor NOR4 (N9384, N9376, N1607, N4764, N6322);
xor XOR2 (N9385, N9359, N7859);
xor XOR2 (N9386, N9381, N5426);
and AND3 (N9387, N9348, N7334, N7900);
buf BUF1 (N9388, N9385);
nor NOR2 (N9389, N9382, N3324);
nand NAND2 (N9390, N9383, N3612);
xor XOR2 (N9391, N9384, N5770);
xor XOR2 (N9392, N9387, N1046);
nor NOR3 (N9393, N9374, N6785, N4101);
nor NOR4 (N9394, N9392, N2085, N6147, N3877);
or OR2 (N9395, N9394, N6137);
nand NAND3 (N9396, N9356, N6751, N8311);
and AND4 (N9397, N9389, N792, N8816, N7801);
not NOT1 (N9398, N9391);
not NOT1 (N9399, N9371);
and AND3 (N9400, N9396, N520, N4120);
or OR3 (N9401, N9398, N5251, N584);
or OR2 (N9402, N9397, N8667);
buf BUF1 (N9403, N9390);
not NOT1 (N9404, N9393);
xor XOR2 (N9405, N9395, N4413);
nor NOR2 (N9406, N9404, N4160);
xor XOR2 (N9407, N9399, N1325);
or OR2 (N9408, N9386, N2160);
not NOT1 (N9409, N9407);
or OR4 (N9410, N9402, N275, N2094, N2931);
or OR2 (N9411, N9388, N795);
and AND3 (N9412, N9401, N2437, N2590);
buf BUF1 (N9413, N9409);
nand NAND2 (N9414, N9375, N9024);
and AND2 (N9415, N9408, N1978);
and AND3 (N9416, N9414, N5489, N4124);
nor NOR3 (N9417, N9403, N8860, N5826);
nand NAND4 (N9418, N9400, N9346, N5968, N3746);
nand NAND3 (N9419, N9415, N3515, N89);
nand NAND2 (N9420, N9417, N1446);
buf BUF1 (N9421, N9413);
xor XOR2 (N9422, N9412, N9309);
and AND4 (N9423, N9421, N6178, N3484, N5759);
or OR2 (N9424, N9416, N5875);
buf BUF1 (N9425, N9410);
or OR2 (N9426, N9423, N6511);
or OR4 (N9427, N9405, N7264, N7651, N402);
or OR3 (N9428, N9424, N8629, N2409);
xor XOR2 (N9429, N9425, N5109);
nand NAND4 (N9430, N9428, N1224, N4186, N4103);
not NOT1 (N9431, N9430);
or OR4 (N9432, N9406, N6491, N8031, N6491);
buf BUF1 (N9433, N9419);
nor NOR2 (N9434, N9426, N7173);
and AND4 (N9435, N9429, N4620, N319, N1301);
nand NAND4 (N9436, N9433, N6829, N9233, N3987);
nand NAND2 (N9437, N9420, N1713);
or OR3 (N9438, N9422, N3438, N5397);
or OR4 (N9439, N9435, N475, N2150, N3760);
nand NAND4 (N9440, N9427, N1363, N5088, N1366);
buf BUF1 (N9441, N9439);
nor NOR2 (N9442, N9431, N3620);
nor NOR2 (N9443, N9441, N3378);
and AND3 (N9444, N9440, N3689, N4936);
not NOT1 (N9445, N9432);
or OR2 (N9446, N9444, N5662);
and AND4 (N9447, N9434, N3816, N4125, N9224);
or OR3 (N9448, N9446, N1473, N5116);
not NOT1 (N9449, N9418);
not NOT1 (N9450, N9445);
and AND3 (N9451, N9438, N2521, N2789);
not NOT1 (N9452, N9449);
nor NOR2 (N9453, N9450, N7733);
nand NAND4 (N9454, N9451, N150, N4598, N2722);
buf BUF1 (N9455, N9452);
nor NOR2 (N9456, N9454, N6431);
not NOT1 (N9457, N9411);
buf BUF1 (N9458, N9436);
not NOT1 (N9459, N9443);
nand NAND3 (N9460, N9458, N6668, N6875);
and AND3 (N9461, N9447, N7839, N8743);
xor XOR2 (N9462, N9457, N1882);
nor NOR3 (N9463, N9462, N156, N7468);
buf BUF1 (N9464, N9437);
and AND3 (N9465, N9460, N6186, N7809);
and AND3 (N9466, N9463, N1413, N7246);
or OR2 (N9467, N9448, N1184);
nor NOR3 (N9468, N9461, N1675, N1236);
nor NOR3 (N9469, N9466, N9099, N6641);
not NOT1 (N9470, N9465);
and AND4 (N9471, N9442, N5019, N6146, N7405);
nand NAND2 (N9472, N9467, N8069);
xor XOR2 (N9473, N9470, N5233);
nand NAND3 (N9474, N9473, N3446, N6654);
buf BUF1 (N9475, N9456);
not NOT1 (N9476, N9474);
nand NAND4 (N9477, N9476, N8296, N2966, N4899);
buf BUF1 (N9478, N9471);
xor XOR2 (N9479, N9464, N6318);
buf BUF1 (N9480, N9468);
not NOT1 (N9481, N9479);
buf BUF1 (N9482, N9478);
and AND3 (N9483, N9455, N5096, N7625);
and AND4 (N9484, N9475, N4635, N163, N2138);
and AND3 (N9485, N9482, N2829, N8630);
or OR4 (N9486, N9453, N1879, N1363, N6796);
nand NAND3 (N9487, N9483, N4253, N7024);
nand NAND2 (N9488, N9487, N5023);
buf BUF1 (N9489, N9486);
or OR3 (N9490, N9484, N4451, N2548);
nand NAND4 (N9491, N9481, N5676, N2056, N4336);
nor NOR4 (N9492, N9477, N6540, N5902, N3984);
xor XOR2 (N9493, N9489, N6706);
nand NAND2 (N9494, N9493, N7208);
not NOT1 (N9495, N9488);
not NOT1 (N9496, N9494);
nor NOR3 (N9497, N9459, N7216, N5791);
nand NAND4 (N9498, N9485, N5153, N4831, N5049);
not NOT1 (N9499, N9497);
nor NOR3 (N9500, N9472, N6319, N1108);
nand NAND4 (N9501, N9496, N1043, N6101, N1138);
and AND3 (N9502, N9492, N5261, N1279);
nor NOR2 (N9503, N9490, N8115);
nor NOR2 (N9504, N9491, N1314);
and AND4 (N9505, N9499, N5068, N3849, N2355);
nor NOR3 (N9506, N9501, N4490, N4009);
nand NAND4 (N9507, N9498, N3395, N8712, N4780);
nand NAND3 (N9508, N9503, N8061, N1517);
and AND3 (N9509, N9480, N3695, N7378);
nor NOR3 (N9510, N9495, N2349, N7521);
xor XOR2 (N9511, N9506, N4748);
or OR3 (N9512, N9504, N3069, N2826);
or OR3 (N9513, N9500, N3319, N5580);
xor XOR2 (N9514, N9512, N5523);
xor XOR2 (N9515, N9505, N1124);
nand NAND2 (N9516, N9513, N1718);
xor XOR2 (N9517, N9502, N1383);
not NOT1 (N9518, N9507);
and AND4 (N9519, N9508, N2733, N4499, N6165);
not NOT1 (N9520, N9517);
xor XOR2 (N9521, N9516, N7548);
nand NAND2 (N9522, N9519, N6601);
nor NOR4 (N9523, N9510, N3633, N2751, N3388);
nand NAND2 (N9524, N9511, N3436);
or OR4 (N9525, N9524, N9101, N5265, N8688);
nand NAND3 (N9526, N9515, N7144, N1301);
nor NOR3 (N9527, N9469, N1211, N76);
nor NOR2 (N9528, N9525, N9006);
not NOT1 (N9529, N9514);
and AND2 (N9530, N9521, N5763);
xor XOR2 (N9531, N9522, N8856);
nand NAND3 (N9532, N9518, N1626, N4083);
and AND3 (N9533, N9528, N2886, N1990);
and AND4 (N9534, N9520, N1969, N626, N6494);
or OR4 (N9535, N9527, N7909, N1019, N9501);
and AND2 (N9536, N9534, N1865);
or OR3 (N9537, N9509, N5253, N4559);
nand NAND2 (N9538, N9533, N3936);
xor XOR2 (N9539, N9531, N2101);
nor NOR4 (N9540, N9529, N2429, N8394, N7409);
or OR3 (N9541, N9526, N5111, N2190);
not NOT1 (N9542, N9536);
nor NOR2 (N9543, N9540, N5017);
or OR2 (N9544, N9542, N8420);
nor NOR4 (N9545, N9544, N2167, N9212, N1848);
or OR3 (N9546, N9539, N936, N7473);
not NOT1 (N9547, N9546);
or OR3 (N9548, N9541, N983, N6651);
not NOT1 (N9549, N9545);
xor XOR2 (N9550, N9547, N2118);
and AND4 (N9551, N9538, N6437, N5598, N6641);
nand NAND3 (N9552, N9532, N5009, N2730);
not NOT1 (N9553, N9549);
or OR4 (N9554, N9537, N2532, N7158, N2385);
or OR2 (N9555, N9552, N4038);
buf BUF1 (N9556, N9553);
nand NAND4 (N9557, N9543, N2792, N397, N5390);
not NOT1 (N9558, N9556);
nor NOR4 (N9559, N9535, N8995, N2821, N2632);
and AND2 (N9560, N9548, N8603);
nor NOR4 (N9561, N9555, N7243, N853, N5748);
xor XOR2 (N9562, N9560, N3774);
buf BUF1 (N9563, N9523);
buf BUF1 (N9564, N9561);
buf BUF1 (N9565, N9563);
and AND3 (N9566, N9551, N2592, N4613);
or OR4 (N9567, N9530, N2269, N3524, N1188);
xor XOR2 (N9568, N9566, N2321);
or OR4 (N9569, N9550, N697, N2557, N4895);
and AND3 (N9570, N9558, N2228, N3855);
not NOT1 (N9571, N9557);
nor NOR4 (N9572, N9564, N626, N3944, N2367);
or OR3 (N9573, N9569, N532, N7957);
nor NOR4 (N9574, N9568, N4949, N2338, N1573);
or OR4 (N9575, N9565, N7221, N2781, N1337);
nand NAND3 (N9576, N9567, N4385, N9358);
xor XOR2 (N9577, N9559, N5761);
buf BUF1 (N9578, N9575);
not NOT1 (N9579, N9574);
xor XOR2 (N9580, N9572, N6523);
and AND2 (N9581, N9573, N6383);
and AND2 (N9582, N9571, N2151);
nand NAND3 (N9583, N9554, N5124, N5026);
nand NAND4 (N9584, N9580, N2805, N8274, N2905);
xor XOR2 (N9585, N9578, N2784);
not NOT1 (N9586, N9579);
not NOT1 (N9587, N9583);
xor XOR2 (N9588, N9585, N4173);
and AND3 (N9589, N9582, N3977, N1313);
and AND3 (N9590, N9577, N5655, N2472);
nand NAND3 (N9591, N9588, N130, N534);
not NOT1 (N9592, N9590);
and AND4 (N9593, N9570, N8484, N146, N177);
and AND2 (N9594, N9586, N3474);
buf BUF1 (N9595, N9581);
xor XOR2 (N9596, N9593, N6959);
nor NOR2 (N9597, N9595, N9089);
buf BUF1 (N9598, N9592);
not NOT1 (N9599, N9594);
xor XOR2 (N9600, N9562, N9111);
nand NAND2 (N9601, N9599, N3797);
nand NAND3 (N9602, N9584, N4303, N873);
nand NAND3 (N9603, N9587, N6009, N2416);
buf BUF1 (N9604, N9576);
nor NOR3 (N9605, N9597, N6432, N6840);
buf BUF1 (N9606, N9605);
not NOT1 (N9607, N9600);
and AND2 (N9608, N9603, N4203);
or OR2 (N9609, N9601, N7559);
or OR3 (N9610, N9609, N1437, N5148);
and AND4 (N9611, N9610, N6160, N1753, N7241);
xor XOR2 (N9612, N9598, N559);
or OR4 (N9613, N9607, N4318, N2297, N5322);
nand NAND2 (N9614, N9604, N9430);
xor XOR2 (N9615, N9611, N1357);
and AND4 (N9616, N9613, N8262, N8454, N5528);
or OR3 (N9617, N9596, N943, N1132);
and AND2 (N9618, N9589, N8109);
buf BUF1 (N9619, N9591);
or OR4 (N9620, N9612, N281, N4563, N2347);
or OR4 (N9621, N9620, N6089, N7200, N2647);
not NOT1 (N9622, N9602);
buf BUF1 (N9623, N9615);
buf BUF1 (N9624, N9614);
not NOT1 (N9625, N9621);
buf BUF1 (N9626, N9617);
buf BUF1 (N9627, N9608);
not NOT1 (N9628, N9606);
nand NAND3 (N9629, N9623, N637, N7106);
buf BUF1 (N9630, N9619);
buf BUF1 (N9631, N9616);
nor NOR2 (N9632, N9618, N7071);
and AND2 (N9633, N9625, N9199);
buf BUF1 (N9634, N9626);
or OR4 (N9635, N9622, N7749, N4463, N5557);
nand NAND4 (N9636, N9633, N2604, N8620, N9110);
or OR4 (N9637, N9632, N8903, N3114, N425);
and AND3 (N9638, N9627, N8097, N7646);
xor XOR2 (N9639, N9635, N8863);
buf BUF1 (N9640, N9631);
nand NAND3 (N9641, N9640, N2298, N8121);
and AND2 (N9642, N9630, N5853);
or OR4 (N9643, N9634, N3242, N481, N5167);
xor XOR2 (N9644, N9628, N5060);
nand NAND4 (N9645, N9639, N6808, N868, N4597);
xor XOR2 (N9646, N9629, N1162);
not NOT1 (N9647, N9643);
or OR3 (N9648, N9647, N4266, N8946);
buf BUF1 (N9649, N9646);
nor NOR4 (N9650, N9641, N950, N533, N3845);
not NOT1 (N9651, N9648);
or OR2 (N9652, N9637, N8460);
and AND3 (N9653, N9624, N8312, N5327);
nor NOR4 (N9654, N9652, N2728, N5771, N2021);
nor NOR4 (N9655, N9638, N8257, N1204, N5804);
not NOT1 (N9656, N9654);
nor NOR2 (N9657, N9649, N2203);
xor XOR2 (N9658, N9651, N3341);
and AND3 (N9659, N9653, N7691, N9293);
or OR3 (N9660, N9650, N5492, N6384);
or OR4 (N9661, N9656, N1555, N3604, N2490);
and AND3 (N9662, N9659, N3520, N833);
buf BUF1 (N9663, N9657);
not NOT1 (N9664, N9636);
buf BUF1 (N9665, N9642);
xor XOR2 (N9666, N9645, N7035);
nand NAND4 (N9667, N9662, N5794, N6793, N2357);
not NOT1 (N9668, N9664);
nor NOR4 (N9669, N9655, N185, N4477, N811);
nand NAND4 (N9670, N9644, N5241, N6023, N8993);
xor XOR2 (N9671, N9661, N8399);
and AND4 (N9672, N9670, N8676, N7456, N6383);
and AND2 (N9673, N9666, N1132);
nor NOR3 (N9674, N9660, N8035, N4422);
not NOT1 (N9675, N9669);
and AND3 (N9676, N9668, N591, N8996);
or OR2 (N9677, N9667, N1373);
xor XOR2 (N9678, N9676, N4717);
nand NAND3 (N9679, N9672, N1774, N4206);
or OR4 (N9680, N9658, N4833, N778, N1666);
nand NAND3 (N9681, N9675, N2914, N7101);
not NOT1 (N9682, N9665);
nand NAND4 (N9683, N9680, N7090, N1227, N3652);
or OR2 (N9684, N9677, N5161);
and AND3 (N9685, N9682, N871, N4286);
nor NOR4 (N9686, N9681, N5285, N7995, N6096);
xor XOR2 (N9687, N9685, N3466);
or OR2 (N9688, N9679, N3702);
and AND3 (N9689, N9684, N8590, N987);
nor NOR4 (N9690, N9683, N393, N2056, N3482);
nor NOR3 (N9691, N9687, N9296, N8803);
and AND2 (N9692, N9689, N5225);
and AND4 (N9693, N9688, N4377, N7752, N2128);
buf BUF1 (N9694, N9678);
buf BUF1 (N9695, N9663);
xor XOR2 (N9696, N9692, N7174);
xor XOR2 (N9697, N9674, N8866);
xor XOR2 (N9698, N9671, N2322);
buf BUF1 (N9699, N9673);
buf BUF1 (N9700, N9698);
not NOT1 (N9701, N9694);
nor NOR2 (N9702, N9701, N3285);
not NOT1 (N9703, N9691);
xor XOR2 (N9704, N9699, N8098);
and AND3 (N9705, N9704, N2401, N2366);
xor XOR2 (N9706, N9693, N1024);
xor XOR2 (N9707, N9705, N8996);
or OR2 (N9708, N9702, N4553);
nor NOR4 (N9709, N9697, N4728, N5354, N5031);
xor XOR2 (N9710, N9709, N6444);
and AND2 (N9711, N9706, N4283);
xor XOR2 (N9712, N9686, N8515);
buf BUF1 (N9713, N9707);
not NOT1 (N9714, N9708);
buf BUF1 (N9715, N9711);
nor NOR3 (N9716, N9700, N5982, N1023);
not NOT1 (N9717, N9695);
buf BUF1 (N9718, N9712);
and AND4 (N9719, N9703, N6327, N7608, N7707);
xor XOR2 (N9720, N9713, N7707);
nor NOR3 (N9721, N9716, N2344, N5393);
or OR4 (N9722, N9721, N5617, N855, N3137);
not NOT1 (N9723, N9714);
buf BUF1 (N9724, N9722);
nor NOR3 (N9725, N9723, N3258, N1695);
and AND3 (N9726, N9696, N3993, N3203);
or OR2 (N9727, N9710, N8793);
xor XOR2 (N9728, N9715, N7281);
nor NOR2 (N9729, N9719, N788);
buf BUF1 (N9730, N9718);
xor XOR2 (N9731, N9727, N8421);
nor NOR3 (N9732, N9725, N7565, N7681);
and AND4 (N9733, N9731, N2684, N3185, N7162);
buf BUF1 (N9734, N9717);
not NOT1 (N9735, N9734);
nor NOR2 (N9736, N9728, N4901);
or OR4 (N9737, N9735, N6285, N2721, N3228);
xor XOR2 (N9738, N9726, N8238);
not NOT1 (N9739, N9733);
buf BUF1 (N9740, N9738);
or OR4 (N9741, N9690, N9461, N8693, N8952);
xor XOR2 (N9742, N9736, N112);
xor XOR2 (N9743, N9741, N479);
nand NAND4 (N9744, N9720, N3099, N6562, N7262);
or OR2 (N9745, N9744, N2351);
xor XOR2 (N9746, N9729, N7160);
not NOT1 (N9747, N9743);
buf BUF1 (N9748, N9737);
nand NAND4 (N9749, N9745, N4624, N74, N7254);
and AND2 (N9750, N9740, N1049);
nand NAND3 (N9751, N9749, N7550, N7332);
and AND4 (N9752, N9739, N2679, N2379, N7643);
not NOT1 (N9753, N9730);
and AND4 (N9754, N9753, N5969, N349, N2307);
not NOT1 (N9755, N9732);
and AND4 (N9756, N9724, N7303, N3647, N9572);
and AND3 (N9757, N9746, N373, N2514);
or OR2 (N9758, N9755, N523);
xor XOR2 (N9759, N9751, N3957);
xor XOR2 (N9760, N9754, N1696);
buf BUF1 (N9761, N9758);
nand NAND3 (N9762, N9760, N2880, N7047);
buf BUF1 (N9763, N9756);
buf BUF1 (N9764, N9748);
nand NAND2 (N9765, N9757, N783);
or OR2 (N9766, N9764, N1913);
nor NOR2 (N9767, N9765, N9296);
or OR2 (N9768, N9752, N612);
nand NAND2 (N9769, N9768, N1002);
xor XOR2 (N9770, N9759, N2185);
nor NOR3 (N9771, N9766, N2403, N5453);
nand NAND2 (N9772, N9763, N3424);
nand NAND4 (N9773, N9770, N3687, N3469, N6713);
not NOT1 (N9774, N9750);
nor NOR4 (N9775, N9773, N8552, N3095, N6611);
and AND4 (N9776, N9775, N8413, N2602, N3377);
nand NAND4 (N9777, N9761, N4030, N7485, N1072);
or OR4 (N9778, N9747, N4498, N4936, N147);
buf BUF1 (N9779, N9777);
or OR2 (N9780, N9778, N8865);
nand NAND3 (N9781, N9772, N3393, N9079);
and AND3 (N9782, N9780, N4174, N3464);
and AND3 (N9783, N9779, N6592, N8126);
nor NOR4 (N9784, N9742, N4914, N8698, N1084);
nand NAND2 (N9785, N9769, N207);
nand NAND2 (N9786, N9776, N9397);
xor XOR2 (N9787, N9785, N724);
not NOT1 (N9788, N9781);
nand NAND3 (N9789, N9783, N6977, N6);
and AND2 (N9790, N9767, N2650);
nor NOR3 (N9791, N9787, N8575, N854);
or OR4 (N9792, N9791, N9670, N3613, N8909);
xor XOR2 (N9793, N9792, N1792);
buf BUF1 (N9794, N9771);
buf BUF1 (N9795, N9794);
buf BUF1 (N9796, N9782);
nand NAND4 (N9797, N9795, N7709, N5177, N9445);
or OR2 (N9798, N9786, N4928);
nor NOR2 (N9799, N9762, N9022);
buf BUF1 (N9800, N9798);
xor XOR2 (N9801, N9800, N2913);
and AND3 (N9802, N9797, N8242, N5247);
xor XOR2 (N9803, N9789, N5855);
not NOT1 (N9804, N9803);
or OR2 (N9805, N9801, N951);
not NOT1 (N9806, N9804);
not NOT1 (N9807, N9784);
or OR3 (N9808, N9805, N3210, N1085);
and AND3 (N9809, N9793, N7133, N7933);
buf BUF1 (N9810, N9799);
xor XOR2 (N9811, N9808, N1814);
not NOT1 (N9812, N9806);
buf BUF1 (N9813, N9788);
xor XOR2 (N9814, N9807, N8753);
not NOT1 (N9815, N9790);
not NOT1 (N9816, N9814);
and AND2 (N9817, N9796, N6676);
buf BUF1 (N9818, N9811);
and AND4 (N9819, N9817, N5233, N6622, N5382);
or OR4 (N9820, N9816, N7796, N459, N7711);
xor XOR2 (N9821, N9819, N578);
or OR3 (N9822, N9810, N9545, N5920);
nor NOR2 (N9823, N9809, N5754);
nor NOR2 (N9824, N9774, N6380);
buf BUF1 (N9825, N9813);
or OR4 (N9826, N9812, N8832, N5268, N8144);
buf BUF1 (N9827, N9824);
or OR2 (N9828, N9820, N6909);
buf BUF1 (N9829, N9823);
and AND3 (N9830, N9815, N4938, N3679);
nor NOR3 (N9831, N9802, N440, N2975);
xor XOR2 (N9832, N9822, N6139);
nor NOR4 (N9833, N9826, N6547, N5871, N1028);
buf BUF1 (N9834, N9833);
xor XOR2 (N9835, N9830, N6046);
buf BUF1 (N9836, N9827);
nor NOR2 (N9837, N9831, N9624);
not NOT1 (N9838, N9828);
and AND4 (N9839, N9834, N4710, N4538, N2830);
nor NOR4 (N9840, N9837, N2896, N8956, N7871);
nor NOR4 (N9841, N9825, N9666, N3569, N6996);
nand NAND4 (N9842, N9836, N8576, N7582, N3827);
xor XOR2 (N9843, N9829, N1603);
nor NOR3 (N9844, N9818, N1770, N9094);
nor NOR2 (N9845, N9843, N1622);
and AND4 (N9846, N9839, N3583, N9075, N6944);
buf BUF1 (N9847, N9841);
not NOT1 (N9848, N9845);
or OR4 (N9849, N9846, N4892, N8348, N5300);
not NOT1 (N9850, N9821);
nand NAND4 (N9851, N9844, N5849, N93, N6575);
or OR2 (N9852, N9832, N9454);
buf BUF1 (N9853, N9842);
nor NOR4 (N9854, N9848, N3987, N3857, N8740);
and AND4 (N9855, N9853, N5982, N4058, N3406);
xor XOR2 (N9856, N9847, N5105);
and AND3 (N9857, N9840, N1930, N9706);
or OR4 (N9858, N9838, N7641, N2259, N9056);
nor NOR3 (N9859, N9857, N9074, N5850);
nor NOR3 (N9860, N9849, N4507, N3146);
buf BUF1 (N9861, N9835);
nand NAND4 (N9862, N9861, N9618, N2209, N1465);
buf BUF1 (N9863, N9854);
buf BUF1 (N9864, N9850);
or OR4 (N9865, N9855, N2420, N7964, N1146);
xor XOR2 (N9866, N9864, N7816);
not NOT1 (N9867, N9863);
or OR2 (N9868, N9859, N8401);
buf BUF1 (N9869, N9868);
nand NAND4 (N9870, N9851, N1473, N9096, N1899);
or OR4 (N9871, N9862, N3389, N8332, N1015);
and AND4 (N9872, N9858, N9662, N8405, N5854);
not NOT1 (N9873, N9870);
buf BUF1 (N9874, N9873);
xor XOR2 (N9875, N9860, N9056);
and AND2 (N9876, N9875, N2283);
nand NAND4 (N9877, N9869, N3516, N6860, N6995);
and AND2 (N9878, N9865, N5605);
and AND2 (N9879, N9874, N1198);
not NOT1 (N9880, N9867);
buf BUF1 (N9881, N9877);
nand NAND4 (N9882, N9878, N8894, N5339, N7018);
xor XOR2 (N9883, N9856, N1395);
xor XOR2 (N9884, N9871, N9765);
xor XOR2 (N9885, N9883, N5161);
or OR4 (N9886, N9852, N8190, N8537, N8657);
nand NAND4 (N9887, N9882, N7999, N8952, N7594);
and AND2 (N9888, N9885, N6035);
xor XOR2 (N9889, N9876, N6303);
not NOT1 (N9890, N9872);
not NOT1 (N9891, N9884);
not NOT1 (N9892, N9886);
xor XOR2 (N9893, N9881, N2926);
xor XOR2 (N9894, N9880, N1038);
and AND2 (N9895, N9894, N9583);
nor NOR4 (N9896, N9889, N2624, N3325, N768);
or OR3 (N9897, N9866, N6416, N4235);
or OR3 (N9898, N9890, N9725, N209);
nand NAND4 (N9899, N9896, N8140, N1752, N744);
and AND4 (N9900, N9897, N1576, N3788, N7323);
buf BUF1 (N9901, N9879);
or OR3 (N9902, N9891, N3572, N8818);
buf BUF1 (N9903, N9892);
and AND2 (N9904, N9895, N7454);
nor NOR2 (N9905, N9887, N1495);
xor XOR2 (N9906, N9899, N1899);
nor NOR4 (N9907, N9906, N4182, N5768, N2838);
and AND2 (N9908, N9900, N1869);
xor XOR2 (N9909, N9903, N8621);
nand NAND2 (N9910, N9905, N2730);
xor XOR2 (N9911, N9909, N8352);
not NOT1 (N9912, N9907);
nor NOR2 (N9913, N9893, N3704);
nor NOR4 (N9914, N9901, N2436, N3497, N2020);
nor NOR4 (N9915, N9913, N231, N6731, N6383);
xor XOR2 (N9916, N9888, N9314);
xor XOR2 (N9917, N9910, N8599);
nor NOR3 (N9918, N9914, N1787, N7373);
xor XOR2 (N9919, N9902, N7994);
or OR2 (N9920, N9908, N9886);
xor XOR2 (N9921, N9915, N5489);
not NOT1 (N9922, N9898);
nand NAND2 (N9923, N9920, N4675);
nor NOR2 (N9924, N9918, N8008);
nand NAND4 (N9925, N9924, N3093, N771, N473);
buf BUF1 (N9926, N9922);
not NOT1 (N9927, N9923);
nor NOR4 (N9928, N9925, N5399, N4931, N9646);
xor XOR2 (N9929, N9904, N7420);
and AND2 (N9930, N9928, N2738);
nor NOR4 (N9931, N9916, N485, N8364, N4377);
nor NOR2 (N9932, N9929, N4824);
nor NOR2 (N9933, N9932, N5091);
nor NOR4 (N9934, N9921, N8780, N3384, N9595);
and AND3 (N9935, N9912, N2315, N3974);
and AND4 (N9936, N9934, N3522, N313, N5696);
buf BUF1 (N9937, N9926);
nor NOR4 (N9938, N9927, N8446, N9273, N8476);
nor NOR4 (N9939, N9937, N5507, N9565, N5199);
not NOT1 (N9940, N9911);
and AND4 (N9941, N9935, N8132, N8974, N1080);
not NOT1 (N9942, N9919);
or OR3 (N9943, N9933, N4939, N9060);
nor NOR4 (N9944, N9942, N50, N5214, N5423);
buf BUF1 (N9945, N9941);
not NOT1 (N9946, N9943);
xor XOR2 (N9947, N9944, N8679);
or OR4 (N9948, N9939, N5629, N1203, N3520);
xor XOR2 (N9949, N9940, N9553);
and AND2 (N9950, N9949, N7497);
nor NOR4 (N9951, N9948, N7650, N7564, N6822);
not NOT1 (N9952, N9930);
not NOT1 (N9953, N9938);
nor NOR2 (N9954, N9936, N872);
xor XOR2 (N9955, N9945, N277);
or OR3 (N9956, N9954, N6884, N800);
or OR4 (N9957, N9950, N7822, N3278, N5487);
buf BUF1 (N9958, N9951);
or OR3 (N9959, N9947, N4559, N8451);
and AND4 (N9960, N9931, N1745, N6689, N5221);
and AND3 (N9961, N9958, N1047, N8159);
or OR3 (N9962, N9959, N1970, N461);
buf BUF1 (N9963, N9960);
or OR4 (N9964, N9953, N4949, N3543, N4861);
and AND2 (N9965, N9963, N7809);
not NOT1 (N9966, N9965);
or OR2 (N9967, N9917, N8670);
or OR2 (N9968, N9966, N9473);
buf BUF1 (N9969, N9961);
and AND3 (N9970, N9969, N5777, N7657);
or OR3 (N9971, N9956, N4218, N2719);
buf BUF1 (N9972, N9962);
buf BUF1 (N9973, N9955);
xor XOR2 (N9974, N9970, N8842);
or OR4 (N9975, N9964, N6945, N274, N884);
nor NOR3 (N9976, N9974, N1384, N8088);
or OR4 (N9977, N9971, N4979, N5614, N1163);
nor NOR2 (N9978, N9973, N7702);
and AND2 (N9979, N9946, N276);
buf BUF1 (N9980, N9979);
nand NAND3 (N9981, N9968, N1717, N8918);
not NOT1 (N9982, N9978);
xor XOR2 (N9983, N9952, N8643);
and AND2 (N9984, N9976, N8927);
not NOT1 (N9985, N9975);
or OR4 (N9986, N9977, N6266, N3073, N5615);
not NOT1 (N9987, N9983);
and AND4 (N9988, N9982, N946, N2142, N571);
buf BUF1 (N9989, N9987);
and AND3 (N9990, N9967, N2074, N1846);
buf BUF1 (N9991, N9990);
nand NAND4 (N9992, N9981, N8959, N1760, N1544);
xor XOR2 (N9993, N9989, N8284);
xor XOR2 (N9994, N9985, N8885);
not NOT1 (N9995, N9984);
nand NAND4 (N9996, N9995, N1519, N9188, N4605);
or OR4 (N9997, N9986, N3041, N7570, N9265);
and AND3 (N9998, N9991, N2920, N2398);
and AND4 (N9999, N9972, N5752, N357, N9166);
and AND2 (N10000, N9957, N5230);
and AND3 (N10001, N9996, N2407, N161);
xor XOR2 (N10002, N9980, N662);
xor XOR2 (N10003, N9999, N5351);
nand NAND2 (N10004, N9988, N9355);
not NOT1 (N10005, N10004);
not NOT1 (N10006, N10002);
buf BUF1 (N10007, N9993);
and AND2 (N10008, N10001, N4031);
nand NAND4 (N10009, N9998, N69, N771, N5273);
nand NAND3 (N10010, N10005, N6009, N3358);
and AND4 (N10011, N10006, N6556, N3377, N7220);
nand NAND2 (N10012, N10010, N5832);
not NOT1 (N10013, N10003);
and AND2 (N10014, N10013, N8521);
xor XOR2 (N10015, N10014, N8590);
nor NOR2 (N10016, N10015, N3738);
nand NAND3 (N10017, N9997, N4258, N2747);
buf BUF1 (N10018, N10016);
not NOT1 (N10019, N10017);
nand NAND4 (N10020, N10009, N622, N9372, N2300);
nand NAND4 (N10021, N10007, N6382, N2787, N5739);
xor XOR2 (N10022, N10012, N8248);
or OR2 (N10023, N9994, N7540);
and AND3 (N10024, N10008, N5089, N4160);
nor NOR4 (N10025, N10022, N5832, N7158, N6365);
buf BUF1 (N10026, N10018);
and AND3 (N10027, N10019, N5563, N3659);
nor NOR3 (N10028, N10011, N3771, N6529);
not NOT1 (N10029, N10023);
nand NAND4 (N10030, N10020, N839, N4385, N2489);
nand NAND2 (N10031, N10029, N9919);
and AND4 (N10032, N10025, N3988, N458, N7862);
buf BUF1 (N10033, N9992);
or OR4 (N10034, N10030, N6754, N4768, N5879);
nand NAND4 (N10035, N10031, N207, N4565, N2098);
nand NAND3 (N10036, N10000, N4855, N3395);
xor XOR2 (N10037, N10035, N9297);
xor XOR2 (N10038, N10034, N5188);
xor XOR2 (N10039, N10026, N6983);
nor NOR4 (N10040, N10037, N7715, N8194, N444);
and AND2 (N10041, N10032, N961);
xor XOR2 (N10042, N10038, N58);
nand NAND2 (N10043, N10041, N7631);
buf BUF1 (N10044, N10028);
and AND3 (N10045, N10044, N1860, N8087);
not NOT1 (N10046, N10027);
xor XOR2 (N10047, N10021, N3456);
buf BUF1 (N10048, N10047);
and AND2 (N10049, N10042, N6032);
buf BUF1 (N10050, N10048);
buf BUF1 (N10051, N10039);
nand NAND2 (N10052, N10043, N4071);
xor XOR2 (N10053, N10040, N4424);
nand NAND3 (N10054, N10024, N7845, N6275);
and AND2 (N10055, N10054, N4090);
buf BUF1 (N10056, N10051);
xor XOR2 (N10057, N10050, N7381);
xor XOR2 (N10058, N10045, N7117);
nor NOR3 (N10059, N10055, N772, N2461);
not NOT1 (N10060, N10059);
and AND2 (N10061, N10060, N7597);
buf BUF1 (N10062, N10053);
and AND3 (N10063, N10056, N375, N8670);
nand NAND4 (N10064, N10057, N260, N984, N2028);
buf BUF1 (N10065, N10036);
or OR3 (N10066, N10049, N9064, N9933);
not NOT1 (N10067, N10062);
nand NAND2 (N10068, N10063, N1944);
nand NAND2 (N10069, N10058, N3688);
or OR4 (N10070, N10067, N2316, N5523, N7596);
xor XOR2 (N10071, N10068, N597);
xor XOR2 (N10072, N10046, N1548);
xor XOR2 (N10073, N10033, N8831);
nand NAND2 (N10074, N10070, N1896);
not NOT1 (N10075, N10073);
not NOT1 (N10076, N10061);
and AND3 (N10077, N10071, N4320, N3376);
and AND3 (N10078, N10074, N7948, N3699);
buf BUF1 (N10079, N10069);
not NOT1 (N10080, N10066);
buf BUF1 (N10081, N10072);
xor XOR2 (N10082, N10077, N130);
and AND2 (N10083, N10080, N5938);
nor NOR2 (N10084, N10082, N6281);
buf BUF1 (N10085, N10075);
or OR2 (N10086, N10052, N2364);
nor NOR2 (N10087, N10084, N491);
nor NOR3 (N10088, N10065, N5901, N961);
xor XOR2 (N10089, N10079, N7322);
not NOT1 (N10090, N10078);
xor XOR2 (N10091, N10076, N4971);
or OR2 (N10092, N10083, N6112);
and AND3 (N10093, N10088, N9912, N3719);
nand NAND2 (N10094, N10093, N5939);
xor XOR2 (N10095, N10064, N3030);
not NOT1 (N10096, N10092);
nand NAND3 (N10097, N10085, N1684, N2276);
nor NOR2 (N10098, N10086, N7341);
nor NOR4 (N10099, N10095, N4671, N414, N5491);
or OR3 (N10100, N10098, N4033, N6582);
nand NAND3 (N10101, N10100, N8829, N6151);
nand NAND3 (N10102, N10081, N6848, N8808);
nor NOR3 (N10103, N10099, N3462, N4859);
not NOT1 (N10104, N10090);
nor NOR4 (N10105, N10094, N4363, N8016, N796);
or OR3 (N10106, N10101, N4117, N8758);
nor NOR2 (N10107, N10091, N4624);
and AND4 (N10108, N10105, N5762, N5666, N791);
or OR3 (N10109, N10102, N1744, N2976);
nor NOR2 (N10110, N10087, N6218);
xor XOR2 (N10111, N10108, N5246);
nand NAND2 (N10112, N10111, N3417);
nor NOR4 (N10113, N10089, N8718, N9556, N7176);
and AND3 (N10114, N10097, N8, N6628);
or OR2 (N10115, N10110, N242);
nand NAND3 (N10116, N10114, N3093, N3013);
and AND3 (N10117, N10113, N662, N3581);
xor XOR2 (N10118, N10107, N5519);
nand NAND3 (N10119, N10104, N2815, N4805);
buf BUF1 (N10120, N10116);
not NOT1 (N10121, N10112);
and AND4 (N10122, N10115, N8114, N6747, N852);
or OR3 (N10123, N10118, N10041, N4922);
nand NAND4 (N10124, N10109, N3560, N3728, N7656);
nor NOR4 (N10125, N10119, N5850, N7647, N4904);
not NOT1 (N10126, N10106);
or OR3 (N10127, N10126, N7285, N5890);
and AND3 (N10128, N10117, N5157, N1447);
and AND4 (N10129, N10124, N1224, N2580, N9686);
nand NAND3 (N10130, N10103, N9934, N5628);
nor NOR4 (N10131, N10130, N9622, N2807, N1734);
nand NAND2 (N10132, N10128, N3520);
nor NOR3 (N10133, N10132, N5621, N8415);
xor XOR2 (N10134, N10121, N9820);
and AND3 (N10135, N10131, N9710, N3553);
nor NOR2 (N10136, N10120, N81);
nor NOR3 (N10137, N10125, N2296, N7759);
nor NOR2 (N10138, N10129, N6925);
or OR4 (N10139, N10137, N7488, N4603, N3747);
and AND4 (N10140, N10136, N1996, N6275, N5697);
or OR4 (N10141, N10134, N194, N4797, N4273);
or OR2 (N10142, N10138, N6068);
xor XOR2 (N10143, N10142, N6111);
nand NAND2 (N10144, N10140, N4705);
buf BUF1 (N10145, N10144);
nor NOR2 (N10146, N10143, N6207);
and AND2 (N10147, N10123, N1382);
xor XOR2 (N10148, N10139, N7516);
not NOT1 (N10149, N10096);
buf BUF1 (N10150, N10127);
or OR2 (N10151, N10141, N4724);
and AND4 (N10152, N10150, N6786, N3725, N2327);
buf BUF1 (N10153, N10152);
and AND3 (N10154, N10146, N4158, N3477);
or OR2 (N10155, N10154, N4875);
buf BUF1 (N10156, N10147);
nor NOR2 (N10157, N10122, N8908);
not NOT1 (N10158, N10148);
or OR4 (N10159, N10145, N8545, N3588, N864);
nor NOR3 (N10160, N10153, N1367, N7955);
and AND2 (N10161, N10135, N9610);
nor NOR3 (N10162, N10160, N1661, N3462);
or OR3 (N10163, N10151, N2645, N8526);
or OR2 (N10164, N10163, N5972);
or OR4 (N10165, N10155, N398, N868, N7247);
xor XOR2 (N10166, N10157, N1040);
nand NAND4 (N10167, N10149, N9560, N369, N709);
nand NAND4 (N10168, N10162, N1577, N9309, N7509);
nand NAND3 (N10169, N10156, N5386, N6706);
and AND3 (N10170, N10166, N4701, N1387);
or OR2 (N10171, N10165, N3936);
nor NOR2 (N10172, N10159, N1702);
or OR3 (N10173, N10169, N53, N2076);
nor NOR3 (N10174, N10170, N7174, N6099);
buf BUF1 (N10175, N10174);
not NOT1 (N10176, N10158);
and AND4 (N10177, N10171, N3607, N3857, N10131);
nand NAND4 (N10178, N10173, N4896, N6907, N8851);
and AND4 (N10179, N10168, N362, N8256, N7805);
nor NOR4 (N10180, N10179, N4406, N2480, N2580);
not NOT1 (N10181, N10178);
or OR4 (N10182, N10164, N9369, N3548, N733);
buf BUF1 (N10183, N10175);
or OR2 (N10184, N10180, N6525);
xor XOR2 (N10185, N10177, N7665);
nor NOR4 (N10186, N10167, N1517, N9757, N9243);
nand NAND2 (N10187, N10186, N1946);
or OR4 (N10188, N10161, N283, N4450, N489);
nand NAND2 (N10189, N10133, N5882);
nor NOR4 (N10190, N10185, N6508, N7553, N5093);
not NOT1 (N10191, N10190);
xor XOR2 (N10192, N10191, N6602);
nor NOR3 (N10193, N10182, N9340, N1696);
not NOT1 (N10194, N10187);
not NOT1 (N10195, N10183);
nand NAND4 (N10196, N10192, N9394, N7599, N2314);
nor NOR2 (N10197, N10194, N4374);
nand NAND4 (N10198, N10172, N631, N1457, N5553);
buf BUF1 (N10199, N10193);
xor XOR2 (N10200, N10176, N7613);
nand NAND4 (N10201, N10198, N2279, N7427, N4486);
or OR3 (N10202, N10199, N6544, N7303);
and AND4 (N10203, N10196, N3829, N7777, N86);
buf BUF1 (N10204, N10203);
nor NOR2 (N10205, N10197, N37);
nand NAND3 (N10206, N10205, N1330, N8648);
and AND2 (N10207, N10184, N8062);
or OR3 (N10208, N10189, N3716, N4720);
and AND2 (N10209, N10195, N847);
not NOT1 (N10210, N10188);
buf BUF1 (N10211, N10210);
nand NAND2 (N10212, N10207, N8349);
nor NOR4 (N10213, N10204, N4044, N1579, N6823);
nand NAND4 (N10214, N10213, N718, N1826, N3247);
nand NAND4 (N10215, N10202, N79, N6133, N4306);
nand NAND2 (N10216, N10200, N5436);
buf BUF1 (N10217, N10216);
buf BUF1 (N10218, N10215);
buf BUF1 (N10219, N10212);
nor NOR2 (N10220, N10211, N7898);
not NOT1 (N10221, N10208);
not NOT1 (N10222, N10209);
buf BUF1 (N10223, N10220);
nand NAND2 (N10224, N10201, N5233);
nor NOR2 (N10225, N10217, N9652);
xor XOR2 (N10226, N10223, N3015);
not NOT1 (N10227, N10206);
xor XOR2 (N10228, N10222, N5121);
and AND4 (N10229, N10224, N8215, N1109, N7642);
nor NOR3 (N10230, N10214, N1905, N8282);
or OR4 (N10231, N10227, N152, N6971, N2383);
nor NOR4 (N10232, N10229, N9385, N5417, N1702);
or OR3 (N10233, N10232, N6462, N8092);
nand NAND4 (N10234, N10218, N3802, N9709, N10006);
buf BUF1 (N10235, N10226);
nor NOR4 (N10236, N10230, N9933, N203, N6988);
or OR2 (N10237, N10231, N3218);
or OR4 (N10238, N10221, N3060, N4955, N6699);
and AND4 (N10239, N10237, N1608, N4697, N3090);
and AND3 (N10240, N10233, N1237, N1848);
nand NAND3 (N10241, N10234, N404, N6594);
and AND3 (N10242, N10219, N661, N7249);
or OR2 (N10243, N10236, N9818);
not NOT1 (N10244, N10243);
not NOT1 (N10245, N10235);
and AND3 (N10246, N10244, N9953, N7351);
not NOT1 (N10247, N10242);
xor XOR2 (N10248, N10240, N957);
buf BUF1 (N10249, N10228);
buf BUF1 (N10250, N10241);
nand NAND3 (N10251, N10181, N9309, N10165);
nor NOR3 (N10252, N10246, N4561, N6187);
and AND4 (N10253, N10238, N6644, N10218, N1801);
buf BUF1 (N10254, N10250);
not NOT1 (N10255, N10225);
nand NAND4 (N10256, N10251, N5965, N1546, N9224);
nor NOR3 (N10257, N10256, N9185, N840);
xor XOR2 (N10258, N10245, N749);
not NOT1 (N10259, N10249);
buf BUF1 (N10260, N10254);
not NOT1 (N10261, N10257);
nand NAND4 (N10262, N10260, N2033, N7944, N8142);
or OR2 (N10263, N10253, N4784);
not NOT1 (N10264, N10247);
nor NOR4 (N10265, N10248, N4805, N5928, N1845);
buf BUF1 (N10266, N10239);
xor XOR2 (N10267, N10258, N5270);
nand NAND4 (N10268, N10255, N7490, N7722, N413);
or OR4 (N10269, N10266, N9120, N8508, N1053);
nand NAND4 (N10270, N10263, N4692, N5994, N9983);
xor XOR2 (N10271, N10262, N9676);
nor NOR4 (N10272, N10261, N5075, N10011, N142);
xor XOR2 (N10273, N10265, N5114);
and AND2 (N10274, N10269, N484);
not NOT1 (N10275, N10273);
not NOT1 (N10276, N10267);
or OR3 (N10277, N10259, N5582, N6216);
xor XOR2 (N10278, N10271, N1773);
or OR2 (N10279, N10272, N4911);
and AND2 (N10280, N10276, N2035);
and AND4 (N10281, N10268, N9993, N4551, N6729);
and AND3 (N10282, N10279, N2691, N5528);
xor XOR2 (N10283, N10280, N6523);
nor NOR2 (N10284, N10264, N1533);
buf BUF1 (N10285, N10277);
buf BUF1 (N10286, N10285);
buf BUF1 (N10287, N10274);
nand NAND4 (N10288, N10281, N7993, N8256, N3754);
xor XOR2 (N10289, N10270, N3476);
nand NAND3 (N10290, N10288, N6320, N3448);
nor NOR4 (N10291, N10283, N874, N7581, N8751);
and AND2 (N10292, N10289, N10233);
buf BUF1 (N10293, N10275);
and AND2 (N10294, N10278, N4353);
not NOT1 (N10295, N10286);
buf BUF1 (N10296, N10287);
and AND4 (N10297, N10294, N4456, N1630, N1000);
or OR2 (N10298, N10292, N6477);
buf BUF1 (N10299, N10282);
xor XOR2 (N10300, N10252, N1048);
or OR4 (N10301, N10299, N6701, N2477, N5781);
xor XOR2 (N10302, N10297, N1771);
and AND3 (N10303, N10291, N9027, N3014);
nand NAND3 (N10304, N10301, N9703, N1771);
and AND2 (N10305, N10295, N4362);
xor XOR2 (N10306, N10298, N3583);
and AND4 (N10307, N10300, N1111, N5611, N8801);
or OR3 (N10308, N10284, N1783, N8104);
nand NAND2 (N10309, N10304, N5103);
buf BUF1 (N10310, N10309);
nor NOR3 (N10311, N10303, N7829, N7063);
nor NOR4 (N10312, N10293, N7894, N6891, N8308);
not NOT1 (N10313, N10302);
or OR2 (N10314, N10307, N8527);
and AND2 (N10315, N10314, N10230);
nor NOR3 (N10316, N10296, N1273, N9493);
nor NOR3 (N10317, N10316, N270, N10234);
and AND3 (N10318, N10310, N796, N10077);
and AND3 (N10319, N10290, N3888, N2555);
nand NAND4 (N10320, N10313, N5877, N975, N1974);
nor NOR2 (N10321, N10311, N1101);
nand NAND2 (N10322, N10312, N6724);
nor NOR3 (N10323, N10322, N7595, N10114);
buf BUF1 (N10324, N10319);
buf BUF1 (N10325, N10320);
nor NOR4 (N10326, N10315, N6352, N1055, N573);
nor NOR3 (N10327, N10317, N1932, N6947);
buf BUF1 (N10328, N10323);
buf BUF1 (N10329, N10325);
nor NOR2 (N10330, N10328, N4220);
buf BUF1 (N10331, N10305);
nand NAND2 (N10332, N10321, N1365);
xor XOR2 (N10333, N10308, N8043);
nor NOR2 (N10334, N10333, N1104);
or OR2 (N10335, N10330, N7939);
and AND3 (N10336, N10318, N1914, N1457);
buf BUF1 (N10337, N10336);
and AND3 (N10338, N10324, N8946, N1759);
nor NOR2 (N10339, N10332, N5998);
not NOT1 (N10340, N10327);
or OR3 (N10341, N10337, N8132, N8915);
nor NOR3 (N10342, N10338, N5241, N2188);
not NOT1 (N10343, N10341);
and AND2 (N10344, N10335, N2000);
and AND3 (N10345, N10306, N8145, N75);
xor XOR2 (N10346, N10340, N3592);
buf BUF1 (N10347, N10346);
and AND4 (N10348, N10339, N10216, N9109, N2498);
not NOT1 (N10349, N10345);
and AND2 (N10350, N10329, N3710);
nor NOR2 (N10351, N10342, N8669);
xor XOR2 (N10352, N10349, N1167);
nand NAND2 (N10353, N10352, N10241);
nand NAND4 (N10354, N10343, N6500, N1585, N9342);
nand NAND4 (N10355, N10354, N4691, N5092, N3147);
or OR2 (N10356, N10355, N9739);
and AND4 (N10357, N10331, N5522, N6853, N5718);
not NOT1 (N10358, N10334);
and AND3 (N10359, N10358, N7758, N2835);
or OR3 (N10360, N10326, N6761, N10284);
or OR3 (N10361, N10357, N6599, N10283);
or OR2 (N10362, N10347, N8388);
and AND4 (N10363, N10348, N9065, N3794, N6376);
not NOT1 (N10364, N10362);
nand NAND3 (N10365, N10359, N9936, N7192);
or OR4 (N10366, N10344, N1221, N3062, N3011);
and AND2 (N10367, N10356, N427);
buf BUF1 (N10368, N10350);
xor XOR2 (N10369, N10351, N7324);
nor NOR4 (N10370, N10369, N300, N6284, N3825);
nand NAND2 (N10371, N10370, N1471);
xor XOR2 (N10372, N10365, N8456);
and AND4 (N10373, N10367, N7655, N55, N4277);
xor XOR2 (N10374, N10353, N5644);
buf BUF1 (N10375, N10368);
and AND4 (N10376, N10373, N10373, N9274, N1637);
and AND2 (N10377, N10363, N65);
or OR4 (N10378, N10366, N8502, N5621, N5577);
xor XOR2 (N10379, N10377, N2826);
nand NAND2 (N10380, N10364, N9861);
not NOT1 (N10381, N10361);
buf BUF1 (N10382, N10374);
buf BUF1 (N10383, N10382);
or OR2 (N10384, N10381, N8493);
or OR2 (N10385, N10383, N2713);
or OR3 (N10386, N10372, N6502, N7562);
and AND3 (N10387, N10376, N4422, N4743);
or OR4 (N10388, N10371, N3098, N6750, N8797);
buf BUF1 (N10389, N10387);
buf BUF1 (N10390, N10379);
or OR4 (N10391, N10380, N9605, N4868, N9385);
xor XOR2 (N10392, N10384, N2420);
nor NOR4 (N10393, N10389, N7617, N9195, N2505);
nor NOR2 (N10394, N10378, N7796);
and AND4 (N10395, N10360, N937, N3579, N4355);
buf BUF1 (N10396, N10392);
or OR2 (N10397, N10395, N5845);
not NOT1 (N10398, N10397);
buf BUF1 (N10399, N10388);
nor NOR3 (N10400, N10386, N5044, N5793);
nor NOR4 (N10401, N10394, N5021, N3649, N8341);
buf BUF1 (N10402, N10391);
not NOT1 (N10403, N10402);
and AND2 (N10404, N10400, N5366);
xor XOR2 (N10405, N10390, N8942);
nor NOR4 (N10406, N10393, N9364, N8084, N5346);
or OR3 (N10407, N10401, N8197, N5060);
buf BUF1 (N10408, N10396);
nor NOR4 (N10409, N10398, N7496, N515, N1505);
or OR4 (N10410, N10408, N9765, N9007, N6226);
not NOT1 (N10411, N10405);
or OR3 (N10412, N10409, N9648, N5205);
nor NOR2 (N10413, N10406, N2436);
nor NOR4 (N10414, N10412, N1923, N10284, N2337);
and AND4 (N10415, N10385, N404, N838, N7480);
not NOT1 (N10416, N10414);
nand NAND4 (N10417, N10416, N2238, N725, N9631);
not NOT1 (N10418, N10404);
xor XOR2 (N10419, N10413, N2343);
nor NOR2 (N10420, N10417, N10171);
or OR2 (N10421, N10407, N4263);
xor XOR2 (N10422, N10403, N62);
not NOT1 (N10423, N10421);
buf BUF1 (N10424, N10420);
and AND2 (N10425, N10423, N1255);
not NOT1 (N10426, N10419);
buf BUF1 (N10427, N10411);
not NOT1 (N10428, N10427);
nand NAND3 (N10429, N10418, N9435, N6765);
nor NOR4 (N10430, N10429, N7570, N9979, N37);
nor NOR3 (N10431, N10415, N5334, N10349);
nor NOR2 (N10432, N10426, N4336);
buf BUF1 (N10433, N10399);
nor NOR4 (N10434, N10410, N2598, N1320, N7737);
or OR2 (N10435, N10431, N10019);
not NOT1 (N10436, N10432);
and AND4 (N10437, N10434, N2371, N6665, N7805);
xor XOR2 (N10438, N10436, N82);
nor NOR3 (N10439, N10438, N2545, N4432);
or OR3 (N10440, N10422, N9411, N5163);
buf BUF1 (N10441, N10430);
nor NOR3 (N10442, N10440, N9284, N8944);
or OR4 (N10443, N10442, N7120, N1199, N4836);
or OR2 (N10444, N10425, N6698);
nand NAND2 (N10445, N10424, N5398);
xor XOR2 (N10446, N10441, N2771);
nand NAND3 (N10447, N10443, N5442, N5016);
and AND4 (N10448, N10446, N1965, N9905, N5956);
and AND2 (N10449, N10437, N3068);
not NOT1 (N10450, N10435);
not NOT1 (N10451, N10445);
nor NOR4 (N10452, N10375, N7812, N3181, N221);
buf BUF1 (N10453, N10451);
buf BUF1 (N10454, N10428);
not NOT1 (N10455, N10449);
not NOT1 (N10456, N10452);
nor NOR2 (N10457, N10444, N3730);
xor XOR2 (N10458, N10448, N10187);
or OR2 (N10459, N10450, N9782);
nand NAND4 (N10460, N10457, N10042, N6889, N916);
not NOT1 (N10461, N10453);
nand NAND4 (N10462, N10433, N1418, N633, N8781);
nand NAND3 (N10463, N10439, N7343, N10200);
not NOT1 (N10464, N10459);
nand NAND2 (N10465, N10447, N8083);
nand NAND4 (N10466, N10465, N8368, N1979, N5486);
nand NAND2 (N10467, N10455, N1964);
nor NOR4 (N10468, N10460, N77, N5843, N5962);
nor NOR2 (N10469, N10454, N7872);
or OR4 (N10470, N10466, N8564, N5922, N7990);
not NOT1 (N10471, N10470);
buf BUF1 (N10472, N10461);
nor NOR2 (N10473, N10472, N4080);
not NOT1 (N10474, N10467);
nor NOR4 (N10475, N10469, N1352, N7942, N476);
xor XOR2 (N10476, N10471, N6712);
nor NOR4 (N10477, N10464, N7676, N7937, N10188);
not NOT1 (N10478, N10463);
nand NAND4 (N10479, N10456, N5923, N6576, N1612);
and AND4 (N10480, N10477, N9969, N4442, N4790);
nand NAND2 (N10481, N10475, N1286);
nor NOR4 (N10482, N10474, N1733, N349, N6295);
buf BUF1 (N10483, N10480);
not NOT1 (N10484, N10481);
nand NAND2 (N10485, N10458, N8415);
xor XOR2 (N10486, N10476, N7299);
buf BUF1 (N10487, N10473);
and AND4 (N10488, N10483, N6978, N2734, N2605);
or OR2 (N10489, N10468, N5002);
nor NOR2 (N10490, N10485, N1798);
xor XOR2 (N10491, N10487, N5083);
nor NOR3 (N10492, N10489, N5321, N7656);
nor NOR4 (N10493, N10492, N962, N356, N7680);
not NOT1 (N10494, N10490);
or OR2 (N10495, N10462, N3698);
and AND2 (N10496, N10484, N3020);
buf BUF1 (N10497, N10482);
buf BUF1 (N10498, N10488);
not NOT1 (N10499, N10498);
not NOT1 (N10500, N10495);
nor NOR3 (N10501, N10479, N6767, N10315);
not NOT1 (N10502, N10486);
not NOT1 (N10503, N10501);
or OR4 (N10504, N10478, N5853, N5184, N3651);
buf BUF1 (N10505, N10496);
or OR4 (N10506, N10502, N581, N3841, N3056);
buf BUF1 (N10507, N10503);
or OR3 (N10508, N10506, N2470, N806);
not NOT1 (N10509, N10497);
nor NOR4 (N10510, N10505, N923, N5151, N10337);
and AND3 (N10511, N10510, N7036, N9400);
and AND3 (N10512, N10504, N271, N9049);
nor NOR4 (N10513, N10507, N2566, N9990, N3565);
buf BUF1 (N10514, N10491);
nor NOR2 (N10515, N10512, N5465);
nand NAND2 (N10516, N10494, N2863);
and AND2 (N10517, N10499, N7231);
or OR4 (N10518, N10514, N4346, N10072, N6875);
buf BUF1 (N10519, N10517);
or OR4 (N10520, N10509, N8235, N371, N2984);
or OR2 (N10521, N10493, N8925);
nor NOR2 (N10522, N10518, N1623);
xor XOR2 (N10523, N10508, N273);
not NOT1 (N10524, N10521);
not NOT1 (N10525, N10500);
buf BUF1 (N10526, N10522);
buf BUF1 (N10527, N10524);
buf BUF1 (N10528, N10513);
xor XOR2 (N10529, N10526, N1111);
not NOT1 (N10530, N10516);
not NOT1 (N10531, N10515);
or OR3 (N10532, N10529, N8976, N3950);
or OR2 (N10533, N10519, N7358);
nor NOR3 (N10534, N10533, N10251, N3415);
not NOT1 (N10535, N10520);
nand NAND4 (N10536, N10531, N9949, N5183, N8456);
and AND3 (N10537, N10535, N664, N3985);
or OR2 (N10538, N10534, N3893);
and AND4 (N10539, N10530, N789, N7752, N6250);
nand NAND3 (N10540, N10532, N21, N4071);
buf BUF1 (N10541, N10511);
not NOT1 (N10542, N10538);
xor XOR2 (N10543, N10539, N3421);
or OR4 (N10544, N10541, N7014, N8790, N1852);
xor XOR2 (N10545, N10525, N7642);
buf BUF1 (N10546, N10540);
xor XOR2 (N10547, N10542, N9322);
or OR2 (N10548, N10537, N2579);
or OR2 (N10549, N10527, N7505);
xor XOR2 (N10550, N10547, N10360);
nor NOR3 (N10551, N10549, N3692, N1126);
and AND2 (N10552, N10528, N1627);
nand NAND4 (N10553, N10546, N3887, N322, N9169);
or OR2 (N10554, N10545, N6334);
buf BUF1 (N10555, N10550);
nand NAND4 (N10556, N10544, N8335, N3301, N1503);
and AND2 (N10557, N10551, N7505);
buf BUF1 (N10558, N10556);
or OR2 (N10559, N10558, N4466);
xor XOR2 (N10560, N10555, N2323);
nor NOR2 (N10561, N10548, N2687);
nand NAND3 (N10562, N10561, N8625, N800);
buf BUF1 (N10563, N10557);
nor NOR2 (N10564, N10560, N1459);
xor XOR2 (N10565, N10552, N2787);
or OR2 (N10566, N10536, N9345);
buf BUF1 (N10567, N10565);
or OR2 (N10568, N10554, N1294);
nand NAND2 (N10569, N10568, N7014);
buf BUF1 (N10570, N10569);
buf BUF1 (N10571, N10523);
xor XOR2 (N10572, N10553, N3430);
nor NOR2 (N10573, N10572, N2487);
nand NAND2 (N10574, N10567, N3129);
buf BUF1 (N10575, N10563);
nor NOR2 (N10576, N10570, N4472);
nor NOR3 (N10577, N10566, N1086, N7736);
nor NOR3 (N10578, N10574, N7199, N5582);
or OR2 (N10579, N10562, N9880);
buf BUF1 (N10580, N10577);
nand NAND4 (N10581, N10580, N2449, N9306, N3706);
or OR4 (N10582, N10576, N6673, N7469, N3698);
xor XOR2 (N10583, N10579, N3234);
not NOT1 (N10584, N10571);
or OR4 (N10585, N10582, N4783, N5701, N5989);
nor NOR2 (N10586, N10573, N10520);
xor XOR2 (N10587, N10585, N7919);
xor XOR2 (N10588, N10587, N10223);
nor NOR4 (N10589, N10578, N9181, N7276, N72);
buf BUF1 (N10590, N10583);
nand NAND4 (N10591, N10575, N8007, N7235, N2978);
not NOT1 (N10592, N10590);
or OR3 (N10593, N10589, N7275, N2233);
or OR4 (N10594, N10592, N2425, N7588, N7086);
buf BUF1 (N10595, N10564);
nand NAND4 (N10596, N10586, N495, N7953, N4978);
buf BUF1 (N10597, N10581);
or OR2 (N10598, N10591, N9269);
or OR3 (N10599, N10596, N2265, N3933);
nand NAND3 (N10600, N10599, N771, N9426);
not NOT1 (N10601, N10593);
nand NAND4 (N10602, N10594, N1523, N1281, N5405);
and AND4 (N10603, N10601, N4861, N6051, N1258);
and AND2 (N10604, N10588, N7832);
buf BUF1 (N10605, N10559);
and AND2 (N10606, N10605, N4711);
not NOT1 (N10607, N10604);
buf BUF1 (N10608, N10584);
nor NOR3 (N10609, N10600, N7582, N3);
nor NOR2 (N10610, N10608, N4499);
not NOT1 (N10611, N10610);
and AND4 (N10612, N10607, N2849, N18, N2889);
or OR3 (N10613, N10597, N3020, N590);
nand NAND2 (N10614, N10606, N5413);
xor XOR2 (N10615, N10609, N9847);
nand NAND3 (N10616, N10613, N296, N5711);
nand NAND2 (N10617, N10615, N5801);
or OR4 (N10618, N10602, N4027, N772, N3405);
and AND2 (N10619, N10595, N6546);
xor XOR2 (N10620, N10543, N2005);
or OR2 (N10621, N10614, N1555);
xor XOR2 (N10622, N10618, N7812);
and AND4 (N10623, N10598, N6662, N7769, N337);
or OR2 (N10624, N10623, N6790);
or OR3 (N10625, N10620, N1999, N433);
nor NOR3 (N10626, N10625, N8632, N1936);
buf BUF1 (N10627, N10611);
or OR4 (N10628, N10617, N1607, N5871, N1347);
and AND4 (N10629, N10616, N2188, N5300, N2742);
or OR3 (N10630, N10624, N4981, N1178);
buf BUF1 (N10631, N10621);
nand NAND3 (N10632, N10626, N4561, N7044);
and AND4 (N10633, N10628, N9979, N8775, N6404);
not NOT1 (N10634, N10612);
xor XOR2 (N10635, N10631, N4472);
xor XOR2 (N10636, N10635, N2053);
xor XOR2 (N10637, N10622, N5512);
and AND3 (N10638, N10627, N7269, N10390);
not NOT1 (N10639, N10603);
and AND3 (N10640, N10639, N1525, N4925);
nand NAND4 (N10641, N10632, N1383, N2815, N6281);
or OR4 (N10642, N10629, N10146, N6374, N1952);
xor XOR2 (N10643, N10640, N7367);
xor XOR2 (N10644, N10642, N9454);
and AND3 (N10645, N10633, N8502, N10573);
buf BUF1 (N10646, N10630);
buf BUF1 (N10647, N10644);
nor NOR2 (N10648, N10637, N7687);
not NOT1 (N10649, N10646);
or OR2 (N10650, N10648, N4236);
buf BUF1 (N10651, N10641);
buf BUF1 (N10652, N10634);
and AND3 (N10653, N10647, N9993, N782);
not NOT1 (N10654, N10619);
and AND3 (N10655, N10650, N8791, N268);
or OR2 (N10656, N10655, N4191);
nand NAND2 (N10657, N10656, N1146);
nand NAND3 (N10658, N10649, N9911, N4645);
buf BUF1 (N10659, N10658);
nand NAND3 (N10660, N10636, N4334, N10636);
nor NOR4 (N10661, N10654, N10257, N806, N1473);
nor NOR2 (N10662, N10645, N10256);
nand NAND2 (N10663, N10659, N4565);
not NOT1 (N10664, N10643);
and AND4 (N10665, N10652, N10613, N4439, N10146);
not NOT1 (N10666, N10665);
nand NAND3 (N10667, N10662, N9041, N4990);
xor XOR2 (N10668, N10661, N9669);
or OR4 (N10669, N10666, N5171, N6337, N5423);
nor NOR4 (N10670, N10651, N1030, N3374, N6212);
not NOT1 (N10671, N10667);
buf BUF1 (N10672, N10660);
and AND4 (N10673, N10657, N5201, N7520, N72);
and AND2 (N10674, N10638, N3003);
and AND4 (N10675, N10668, N8276, N9132, N1059);
buf BUF1 (N10676, N10674);
and AND3 (N10677, N10672, N1719, N1543);
or OR4 (N10678, N10664, N9758, N9313, N8305);
not NOT1 (N10679, N10673);
xor XOR2 (N10680, N10653, N4763);
and AND4 (N10681, N10663, N5033, N10187, N6581);
not NOT1 (N10682, N10669);
and AND4 (N10683, N10680, N1248, N1487, N7593);
nor NOR2 (N10684, N10678, N7438);
nand NAND4 (N10685, N10684, N102, N2556, N1526);
and AND3 (N10686, N10670, N4924, N6478);
xor XOR2 (N10687, N10676, N5347);
buf BUF1 (N10688, N10677);
not NOT1 (N10689, N10679);
not NOT1 (N10690, N10686);
not NOT1 (N10691, N10690);
xor XOR2 (N10692, N10691, N8316);
nor NOR3 (N10693, N10692, N3491, N5423);
xor XOR2 (N10694, N10681, N2037);
and AND3 (N10695, N10683, N1695, N5914);
or OR2 (N10696, N10693, N4685);
buf BUF1 (N10697, N10671);
or OR2 (N10698, N10687, N7813);
not NOT1 (N10699, N10675);
not NOT1 (N10700, N10696);
nor NOR3 (N10701, N10694, N316, N2455);
or OR2 (N10702, N10695, N5573);
not NOT1 (N10703, N10702);
and AND2 (N10704, N10699, N5922);
not NOT1 (N10705, N10682);
or OR3 (N10706, N10697, N9635, N9678);
not NOT1 (N10707, N10706);
not NOT1 (N10708, N10703);
nand NAND2 (N10709, N10704, N9550);
xor XOR2 (N10710, N10689, N1784);
xor XOR2 (N10711, N10698, N4553);
not NOT1 (N10712, N10685);
or OR4 (N10713, N10711, N4849, N7848, N8092);
or OR3 (N10714, N10707, N5595, N9873);
nand NAND3 (N10715, N10700, N7024, N3719);
buf BUF1 (N10716, N10713);
or OR4 (N10717, N10701, N731, N5615, N1013);
buf BUF1 (N10718, N10705);
or OR4 (N10719, N10718, N4220, N1114, N8659);
xor XOR2 (N10720, N10708, N3106);
or OR2 (N10721, N10710, N5024);
xor XOR2 (N10722, N10714, N8686);
and AND3 (N10723, N10688, N5834, N6577);
nor NOR2 (N10724, N10721, N2914);
xor XOR2 (N10725, N10719, N10365);
nor NOR3 (N10726, N10715, N2862, N8754);
or OR2 (N10727, N10709, N2533);
not NOT1 (N10728, N10723);
nand NAND4 (N10729, N10726, N3322, N3937, N5022);
not NOT1 (N10730, N10712);
nand NAND2 (N10731, N10725, N3272);
and AND2 (N10732, N10727, N7903);
or OR3 (N10733, N10732, N3593, N5465);
buf BUF1 (N10734, N10728);
nor NOR3 (N10735, N10717, N4272, N7937);
not NOT1 (N10736, N10731);
xor XOR2 (N10737, N10720, N5098);
nor NOR3 (N10738, N10735, N955, N8669);
nor NOR2 (N10739, N10729, N840);
and AND4 (N10740, N10730, N411, N677, N3355);
and AND3 (N10741, N10739, N6895, N5787);
or OR3 (N10742, N10716, N1989, N9230);
and AND4 (N10743, N10742, N396, N6940, N2315);
buf BUF1 (N10744, N10724);
not NOT1 (N10745, N10741);
not NOT1 (N10746, N10734);
or OR2 (N10747, N10745, N9538);
nor NOR4 (N10748, N10722, N2675, N968, N4696);
and AND4 (N10749, N10743, N2933, N6153, N438);
nor NOR3 (N10750, N10736, N9011, N8502);
and AND3 (N10751, N10744, N5658, N1086);
or OR3 (N10752, N10750, N1755, N9410);
nand NAND3 (N10753, N10738, N2627, N4894);
nor NOR4 (N10754, N10752, N286, N5058, N8519);
buf BUF1 (N10755, N10754);
nor NOR3 (N10756, N10746, N5391, N5254);
or OR3 (N10757, N10733, N1673, N1165);
nor NOR3 (N10758, N10755, N5126, N6699);
buf BUF1 (N10759, N10751);
nor NOR3 (N10760, N10740, N6356, N5483);
not NOT1 (N10761, N10756);
nor NOR3 (N10762, N10757, N3219, N4392);
nor NOR3 (N10763, N10761, N2386, N7013);
buf BUF1 (N10764, N10763);
buf BUF1 (N10765, N10748);
or OR4 (N10766, N10765, N9203, N4780, N6600);
buf BUF1 (N10767, N10747);
not NOT1 (N10768, N10764);
buf BUF1 (N10769, N10768);
and AND4 (N10770, N10749, N8685, N2363, N515);
xor XOR2 (N10771, N10769, N10672);
nor NOR3 (N10772, N10753, N2229, N7814);
not NOT1 (N10773, N10771);
nand NAND4 (N10774, N10737, N9480, N9402, N5633);
buf BUF1 (N10775, N10773);
nand NAND4 (N10776, N10770, N7145, N5137, N8293);
and AND2 (N10777, N10772, N30);
nor NOR2 (N10778, N10775, N2160);
nand NAND4 (N10779, N10776, N2427, N7442, N6805);
and AND3 (N10780, N10774, N1686, N89);
nor NOR2 (N10781, N10777, N319);
xor XOR2 (N10782, N10778, N9832);
nand NAND3 (N10783, N10759, N4671, N10313);
or OR4 (N10784, N10783, N6074, N6206, N4875);
nand NAND2 (N10785, N10766, N4251);
buf BUF1 (N10786, N10781);
or OR4 (N10787, N10784, N2951, N6935, N5888);
or OR2 (N10788, N10786, N2532);
nand NAND2 (N10789, N10762, N4122);
nor NOR4 (N10790, N10779, N7851, N7873, N4160);
or OR3 (N10791, N10760, N5163, N4432);
nor NOR3 (N10792, N10785, N7154, N8971);
nor NOR4 (N10793, N10758, N1186, N6474, N1090);
and AND3 (N10794, N10767, N2773, N966);
not NOT1 (N10795, N10787);
buf BUF1 (N10796, N10782);
buf BUF1 (N10797, N10795);
or OR4 (N10798, N10797, N2283, N5156, N985);
nor NOR3 (N10799, N10796, N4317, N7575);
nand NAND2 (N10800, N10799, N3843);
nor NOR4 (N10801, N10792, N552, N10353, N2801);
buf BUF1 (N10802, N10788);
buf BUF1 (N10803, N10789);
nand NAND4 (N10804, N10794, N5034, N1030, N2304);
not NOT1 (N10805, N10793);
xor XOR2 (N10806, N10803, N9523);
not NOT1 (N10807, N10806);
nand NAND2 (N10808, N10798, N4079);
not NOT1 (N10809, N10780);
buf BUF1 (N10810, N10791);
and AND2 (N10811, N10808, N2046);
buf BUF1 (N10812, N10801);
buf BUF1 (N10813, N10790);
nand NAND3 (N10814, N10807, N8288, N5566);
nand NAND3 (N10815, N10805, N7263, N6176);
nand NAND2 (N10816, N10804, N3345);
and AND2 (N10817, N10800, N1346);
not NOT1 (N10818, N10809);
buf BUF1 (N10819, N10812);
xor XOR2 (N10820, N10818, N2121);
buf BUF1 (N10821, N10817);
buf BUF1 (N10822, N10816);
nor NOR2 (N10823, N10822, N5325);
not NOT1 (N10824, N10821);
xor XOR2 (N10825, N10811, N5321);
or OR2 (N10826, N10814, N9391);
not NOT1 (N10827, N10820);
xor XOR2 (N10828, N10825, N2963);
buf BUF1 (N10829, N10826);
buf BUF1 (N10830, N10823);
not NOT1 (N10831, N10813);
xor XOR2 (N10832, N10810, N5642);
xor XOR2 (N10833, N10831, N2940);
or OR2 (N10834, N10833, N9746);
buf BUF1 (N10835, N10828);
nand NAND2 (N10836, N10834, N950);
xor XOR2 (N10837, N10835, N3208);
or OR2 (N10838, N10815, N2627);
xor XOR2 (N10839, N10836, N7005);
nor NOR3 (N10840, N10839, N9118, N2852);
or OR3 (N10841, N10832, N8380, N2807);
xor XOR2 (N10842, N10824, N1291);
nand NAND2 (N10843, N10840, N6681);
or OR4 (N10844, N10829, N3854, N307, N2873);
xor XOR2 (N10845, N10844, N4439);
nor NOR4 (N10846, N10830, N7337, N8568, N1833);
not NOT1 (N10847, N10843);
nor NOR2 (N10848, N10827, N1954);
nand NAND4 (N10849, N10842, N2328, N3705, N2597);
nor NOR2 (N10850, N10849, N3463);
not NOT1 (N10851, N10841);
nor NOR4 (N10852, N10851, N6943, N10503, N1149);
buf BUF1 (N10853, N10845);
or OR2 (N10854, N10853, N10068);
nor NOR4 (N10855, N10837, N792, N9511, N2214);
nand NAND2 (N10856, N10838, N5533);
or OR3 (N10857, N10850, N4714, N4446);
xor XOR2 (N10858, N10856, N3461);
nor NOR3 (N10859, N10847, N8096, N10437);
or OR2 (N10860, N10852, N5473);
nor NOR2 (N10861, N10854, N6098);
xor XOR2 (N10862, N10855, N3323);
buf BUF1 (N10863, N10857);
xor XOR2 (N10864, N10819, N10015);
or OR3 (N10865, N10846, N4895, N8471);
nor NOR4 (N10866, N10861, N6282, N8632, N265);
xor XOR2 (N10867, N10863, N2118);
and AND3 (N10868, N10865, N1406, N10481);
not NOT1 (N10869, N10859);
xor XOR2 (N10870, N10868, N2990);
nor NOR2 (N10871, N10870, N3547);
nor NOR2 (N10872, N10869, N2573);
not NOT1 (N10873, N10872);
buf BUF1 (N10874, N10802);
nand NAND3 (N10875, N10873, N8237, N1714);
or OR3 (N10876, N10871, N4875, N9660);
nor NOR2 (N10877, N10864, N2943);
and AND2 (N10878, N10848, N7071);
buf BUF1 (N10879, N10860);
or OR3 (N10880, N10866, N7879, N6474);
not NOT1 (N10881, N10877);
nor NOR2 (N10882, N10858, N10268);
buf BUF1 (N10883, N10876);
nor NOR3 (N10884, N10874, N7440, N10247);
nor NOR2 (N10885, N10883, N10803);
xor XOR2 (N10886, N10867, N5022);
or OR3 (N10887, N10881, N295, N5919);
not NOT1 (N10888, N10879);
or OR4 (N10889, N10862, N7688, N6720, N5672);
xor XOR2 (N10890, N10882, N4455);
xor XOR2 (N10891, N10875, N5805);
nor NOR2 (N10892, N10888, N8916);
nor NOR2 (N10893, N10880, N1584);
or OR3 (N10894, N10884, N8014, N1665);
not NOT1 (N10895, N10885);
nor NOR4 (N10896, N10891, N5165, N273, N5019);
or OR2 (N10897, N10893, N2807);
or OR2 (N10898, N10878, N1575);
xor XOR2 (N10899, N10897, N900);
not NOT1 (N10900, N10887);
xor XOR2 (N10901, N10889, N4018);
and AND3 (N10902, N10886, N363, N10760);
or OR3 (N10903, N10902, N58, N10893);
and AND4 (N10904, N10899, N5819, N10754, N1359);
nor NOR2 (N10905, N10898, N6634);
nor NOR3 (N10906, N10900, N1673, N7646);
xor XOR2 (N10907, N10903, N1372);
nor NOR4 (N10908, N10906, N992, N1151, N7499);
nor NOR2 (N10909, N10907, N10826);
not NOT1 (N10910, N10896);
and AND4 (N10911, N10910, N8043, N862, N6556);
buf BUF1 (N10912, N10909);
xor XOR2 (N10913, N10912, N1326);
xor XOR2 (N10914, N10894, N3593);
nand NAND4 (N10915, N10895, N4803, N8391, N4078);
or OR3 (N10916, N10913, N5410, N4803);
or OR2 (N10917, N10901, N3233);
not NOT1 (N10918, N10917);
buf BUF1 (N10919, N10892);
buf BUF1 (N10920, N10918);
or OR4 (N10921, N10919, N6688, N10023, N3852);
and AND4 (N10922, N10911, N2136, N10111, N9407);
buf BUF1 (N10923, N10914);
not NOT1 (N10924, N10904);
xor XOR2 (N10925, N10921, N3842);
xor XOR2 (N10926, N10905, N10360);
not NOT1 (N10927, N10924);
not NOT1 (N10928, N10925);
and AND3 (N10929, N10890, N7686, N6693);
buf BUF1 (N10930, N10915);
and AND3 (N10931, N10923, N5380, N9970);
not NOT1 (N10932, N10929);
nand NAND4 (N10933, N10927, N7085, N7276, N10146);
not NOT1 (N10934, N10922);
or OR2 (N10935, N10928, N3949);
nor NOR2 (N10936, N10934, N3072);
or OR2 (N10937, N10930, N1219);
xor XOR2 (N10938, N10936, N2349);
nor NOR4 (N10939, N10932, N3302, N10759, N789);
not NOT1 (N10940, N10935);
not NOT1 (N10941, N10933);
buf BUF1 (N10942, N10920);
buf BUF1 (N10943, N10939);
not NOT1 (N10944, N10940);
and AND3 (N10945, N10943, N683, N90);
buf BUF1 (N10946, N10945);
xor XOR2 (N10947, N10931, N5918);
nand NAND3 (N10948, N10938, N2134, N5730);
not NOT1 (N10949, N10946);
and AND4 (N10950, N10916, N6506, N8453, N8910);
nand NAND2 (N10951, N10908, N8491);
buf BUF1 (N10952, N10926);
buf BUF1 (N10953, N10951);
not NOT1 (N10954, N10944);
buf BUF1 (N10955, N10950);
nand NAND3 (N10956, N10947, N10893, N1505);
and AND4 (N10957, N10948, N7328, N5570, N655);
and AND2 (N10958, N10949, N620);
nor NOR2 (N10959, N10953, N8297);
not NOT1 (N10960, N10941);
and AND2 (N10961, N10959, N7164);
and AND4 (N10962, N10942, N847, N6276, N5720);
or OR4 (N10963, N10961, N581, N7608, N662);
nor NOR3 (N10964, N10937, N1328, N9882);
nand NAND3 (N10965, N10956, N3418, N1778);
nand NAND4 (N10966, N10952, N1503, N1785, N2205);
nor NOR2 (N10967, N10962, N5286);
or OR4 (N10968, N10955, N7418, N3436, N5118);
nor NOR4 (N10969, N10957, N5504, N4125, N3337);
nand NAND3 (N10970, N10960, N4538, N8366);
not NOT1 (N10971, N10967);
not NOT1 (N10972, N10958);
nand NAND3 (N10973, N10968, N2483, N2081);
buf BUF1 (N10974, N10954);
not NOT1 (N10975, N10969);
nor NOR4 (N10976, N10964, N1203, N10722, N3332);
nor NOR4 (N10977, N10966, N1247, N4903, N8205);
buf BUF1 (N10978, N10970);
nor NOR3 (N10979, N10976, N2090, N7131);
and AND2 (N10980, N10971, N1596);
nor NOR3 (N10981, N10973, N4670, N6298);
not NOT1 (N10982, N10977);
or OR3 (N10983, N10981, N10532, N7952);
not NOT1 (N10984, N10980);
nand NAND2 (N10985, N10982, N2330);
xor XOR2 (N10986, N10975, N967);
buf BUF1 (N10987, N10963);
not NOT1 (N10988, N10986);
or OR3 (N10989, N10972, N1862, N9297);
buf BUF1 (N10990, N10978);
nand NAND3 (N10991, N10979, N1030, N1233);
nor NOR3 (N10992, N10985, N5859, N8329);
buf BUF1 (N10993, N10992);
and AND3 (N10994, N10990, N5883, N9831);
buf BUF1 (N10995, N10991);
nand NAND4 (N10996, N10974, N10531, N6551, N1759);
nor NOR3 (N10997, N10965, N2899, N1898);
or OR3 (N10998, N10988, N6072, N2705);
nand NAND4 (N10999, N10989, N3695, N602, N9235);
or OR4 (N11000, N10998, N434, N7798, N28);
not NOT1 (N11001, N10997);
nor NOR2 (N11002, N11001, N6671);
and AND2 (N11003, N10994, N5500);
buf BUF1 (N11004, N10996);
not NOT1 (N11005, N10995);
nor NOR3 (N11006, N11000, N2353, N686);
buf BUF1 (N11007, N10987);
and AND4 (N11008, N11002, N10338, N8658, N7309);
nand NAND3 (N11009, N11003, N8832, N6792);
nand NAND2 (N11010, N11005, N5977);
buf BUF1 (N11011, N11009);
xor XOR2 (N11012, N11004, N7621);
or OR2 (N11013, N11011, N9205);
or OR3 (N11014, N10983, N1474, N7494);
nand NAND4 (N11015, N11008, N3403, N9253, N3062);
nand NAND2 (N11016, N10984, N7913);
nor NOR3 (N11017, N11007, N9220, N5267);
nand NAND4 (N11018, N11017, N4954, N7592, N3736);
xor XOR2 (N11019, N11014, N759);
nand NAND2 (N11020, N10993, N372);
nand NAND3 (N11021, N11016, N253, N3228);
not NOT1 (N11022, N11010);
xor XOR2 (N11023, N11021, N4388);
buf BUF1 (N11024, N11022);
xor XOR2 (N11025, N11015, N5294);
nor NOR3 (N11026, N11024, N2708, N1002);
buf BUF1 (N11027, N11020);
and AND4 (N11028, N10999, N7155, N7043, N10933);
xor XOR2 (N11029, N11023, N6321);
nand NAND4 (N11030, N11027, N3532, N4572, N6544);
xor XOR2 (N11031, N11025, N10174);
or OR4 (N11032, N11026, N8310, N2065, N1125);
and AND3 (N11033, N11018, N6719, N562);
not NOT1 (N11034, N11029);
buf BUF1 (N11035, N11034);
or OR4 (N11036, N11012, N8426, N3818, N10483);
nand NAND4 (N11037, N11019, N3765, N9413, N7696);
nand NAND3 (N11038, N11013, N6388, N9771);
nor NOR4 (N11039, N11033, N5647, N6595, N3636);
xor XOR2 (N11040, N11031, N2999);
nor NOR2 (N11041, N11006, N7623);
nor NOR4 (N11042, N11028, N5920, N5246, N4514);
nor NOR2 (N11043, N11030, N7345);
and AND3 (N11044, N11035, N2156, N1720);
not NOT1 (N11045, N11037);
nand NAND3 (N11046, N11044, N10474, N7083);
nand NAND3 (N11047, N11040, N420, N6792);
buf BUF1 (N11048, N11045);
not NOT1 (N11049, N11032);
and AND2 (N11050, N11042, N8463);
not NOT1 (N11051, N11038);
not NOT1 (N11052, N11049);
or OR2 (N11053, N11039, N126);
nor NOR3 (N11054, N11043, N219, N4301);
buf BUF1 (N11055, N11053);
nor NOR3 (N11056, N11048, N3785, N9778);
or OR3 (N11057, N11055, N6907, N2181);
buf BUF1 (N11058, N11052);
nor NOR4 (N11059, N11046, N769, N5229, N334);
buf BUF1 (N11060, N11050);
nor NOR3 (N11061, N11036, N8803, N270);
not NOT1 (N11062, N11057);
not NOT1 (N11063, N11051);
and AND3 (N11064, N11058, N6991, N4026);
not NOT1 (N11065, N11062);
and AND2 (N11066, N11041, N4603);
and AND4 (N11067, N11056, N5465, N5529, N9800);
nand NAND2 (N11068, N11059, N337);
or OR4 (N11069, N11047, N8303, N1780, N8442);
or OR4 (N11070, N11064, N6364, N811, N3699);
nand NAND3 (N11071, N11060, N6340, N10518);
buf BUF1 (N11072, N11068);
and AND3 (N11073, N11065, N9050, N9651);
xor XOR2 (N11074, N11073, N2199);
and AND3 (N11075, N11074, N9857, N7857);
buf BUF1 (N11076, N11067);
not NOT1 (N11077, N11066);
nand NAND3 (N11078, N11063, N22, N5112);
nand NAND2 (N11079, N11078, N4830);
and AND4 (N11080, N11070, N8082, N9066, N9768);
not NOT1 (N11081, N11069);
xor XOR2 (N11082, N11072, N1497);
not NOT1 (N11083, N11061);
buf BUF1 (N11084, N11082);
nor NOR3 (N11085, N11080, N9809, N7305);
buf BUF1 (N11086, N11085);
nand NAND2 (N11087, N11081, N9676);
and AND2 (N11088, N11054, N2091);
xor XOR2 (N11089, N11083, N9226);
and AND4 (N11090, N11088, N6127, N810, N10374);
and AND4 (N11091, N11087, N6777, N10767, N6064);
and AND3 (N11092, N11075, N1617, N639);
xor XOR2 (N11093, N11071, N3575);
and AND2 (N11094, N11092, N5906);
and AND3 (N11095, N11089, N8398, N8333);
nor NOR4 (N11096, N11079, N5128, N1852, N6873);
or OR3 (N11097, N11091, N2132, N7834);
and AND3 (N11098, N11076, N2756, N446);
nor NOR2 (N11099, N11090, N5722);
xor XOR2 (N11100, N11098, N8883);
nand NAND4 (N11101, N11096, N9021, N9621, N7961);
nor NOR3 (N11102, N11077, N3943, N2018);
xor XOR2 (N11103, N11084, N1284);
not NOT1 (N11104, N11100);
nor NOR4 (N11105, N11103, N2480, N5978, N5427);
or OR4 (N11106, N11101, N1988, N2734, N6218);
xor XOR2 (N11107, N11095, N10100);
nor NOR4 (N11108, N11097, N9633, N953, N4601);
not NOT1 (N11109, N11108);
xor XOR2 (N11110, N11093, N8037);
not NOT1 (N11111, N11106);
nand NAND3 (N11112, N11104, N547, N5709);
and AND2 (N11113, N11107, N2532);
nand NAND3 (N11114, N11094, N9091, N7832);
buf BUF1 (N11115, N11114);
and AND4 (N11116, N11086, N4498, N1421, N4855);
xor XOR2 (N11117, N11110, N1156);
nor NOR4 (N11118, N11102, N1020, N1456, N6116);
or OR2 (N11119, N11112, N10300);
buf BUF1 (N11120, N11115);
not NOT1 (N11121, N11116);
nor NOR2 (N11122, N11117, N9432);
nand NAND3 (N11123, N11109, N9695, N7478);
buf BUF1 (N11124, N11111);
or OR2 (N11125, N11099, N6759);
and AND2 (N11126, N11123, N4182);
nand NAND2 (N11127, N11121, N4617);
nor NOR4 (N11128, N11105, N1810, N10679, N419);
nor NOR4 (N11129, N11125, N9619, N132, N8292);
not NOT1 (N11130, N11124);
nor NOR3 (N11131, N11113, N4304, N9557);
nor NOR3 (N11132, N11120, N212, N6911);
buf BUF1 (N11133, N11129);
and AND2 (N11134, N11118, N1115);
nand NAND4 (N11135, N11127, N501, N1788, N7439);
nor NOR3 (N11136, N11130, N4399, N5692);
or OR3 (N11137, N11128, N7911, N2137);
or OR4 (N11138, N11137, N8356, N8277, N3671);
or OR4 (N11139, N11138, N1283, N10074, N10734);
nand NAND2 (N11140, N11131, N8867);
not NOT1 (N11141, N11122);
nand NAND4 (N11142, N11136, N5538, N5525, N2319);
nor NOR3 (N11143, N11126, N7107, N1233);
and AND4 (N11144, N11132, N10647, N3038, N5426);
buf BUF1 (N11145, N11142);
and AND3 (N11146, N11140, N7348, N254);
and AND2 (N11147, N11134, N7592);
and AND4 (N11148, N11144, N2342, N9196, N6499);
or OR4 (N11149, N11141, N2050, N3259, N5563);
nand NAND4 (N11150, N11135, N9230, N10479, N6260);
not NOT1 (N11151, N11143);
xor XOR2 (N11152, N11119, N2883);
not NOT1 (N11153, N11133);
buf BUF1 (N11154, N11146);
not NOT1 (N11155, N11154);
or OR4 (N11156, N11150, N7545, N135, N468);
xor XOR2 (N11157, N11152, N2673);
xor XOR2 (N11158, N11157, N9872);
or OR4 (N11159, N11153, N566, N5219, N9147);
nand NAND4 (N11160, N11156, N4947, N352, N2870);
xor XOR2 (N11161, N11149, N6727);
or OR3 (N11162, N11161, N2814, N2104);
or OR2 (N11163, N11162, N7080);
or OR3 (N11164, N11158, N8045, N3698);
or OR4 (N11165, N11139, N7861, N3122, N5363);
xor XOR2 (N11166, N11163, N10570);
and AND3 (N11167, N11151, N7903, N11074);
or OR3 (N11168, N11155, N2865, N4257);
xor XOR2 (N11169, N11148, N2626);
and AND3 (N11170, N11145, N4713, N7396);
nand NAND3 (N11171, N11165, N8485, N4118);
and AND4 (N11172, N11167, N6082, N2645, N3720);
nor NOR2 (N11173, N11169, N9979);
or OR4 (N11174, N11164, N6363, N1950, N5633);
or OR4 (N11175, N11173, N8704, N2305, N6734);
and AND2 (N11176, N11175, N3018);
not NOT1 (N11177, N11147);
not NOT1 (N11178, N11177);
nand NAND4 (N11179, N11172, N6960, N4670, N3395);
not NOT1 (N11180, N11160);
or OR3 (N11181, N11179, N2070, N5261);
nand NAND4 (N11182, N11171, N10196, N1602, N8998);
nand NAND2 (N11183, N11170, N10569);
xor XOR2 (N11184, N11174, N7161);
and AND2 (N11185, N11181, N9748);
nand NAND2 (N11186, N11180, N912);
and AND3 (N11187, N11159, N271, N4459);
nand NAND2 (N11188, N11185, N5273);
not NOT1 (N11189, N11188);
nand NAND2 (N11190, N11168, N8969);
not NOT1 (N11191, N11166);
not NOT1 (N11192, N11191);
not NOT1 (N11193, N11182);
nor NOR3 (N11194, N11184, N1387, N4907);
xor XOR2 (N11195, N11192, N7183);
and AND4 (N11196, N11186, N5436, N3832, N758);
and AND4 (N11197, N11194, N10925, N7500, N7451);
and AND2 (N11198, N11196, N6451);
xor XOR2 (N11199, N11187, N7435);
nand NAND4 (N11200, N11189, N4843, N3454, N9733);
xor XOR2 (N11201, N11183, N9133);
not NOT1 (N11202, N11198);
nor NOR3 (N11203, N11195, N9677, N7099);
buf BUF1 (N11204, N11178);
nand NAND4 (N11205, N11199, N6897, N11085, N2032);
xor XOR2 (N11206, N11176, N4419);
nor NOR3 (N11207, N11193, N4298, N7715);
nand NAND2 (N11208, N11207, N2312);
buf BUF1 (N11209, N11206);
xor XOR2 (N11210, N11205, N10807);
and AND2 (N11211, N11204, N3966);
nor NOR3 (N11212, N11202, N3959, N4257);
xor XOR2 (N11213, N11208, N4034);
xor XOR2 (N11214, N11212, N7314);
and AND3 (N11215, N11190, N1655, N6738);
buf BUF1 (N11216, N11215);
not NOT1 (N11217, N11210);
nor NOR3 (N11218, N11213, N8869, N8052);
not NOT1 (N11219, N11201);
nand NAND4 (N11220, N11209, N5164, N6796, N9472);
and AND2 (N11221, N11203, N1370);
and AND3 (N11222, N11217, N2759, N618);
and AND2 (N11223, N11214, N2793);
or OR4 (N11224, N11222, N2211, N1067, N2543);
nor NOR4 (N11225, N11223, N5444, N6295, N8433);
not NOT1 (N11226, N11216);
xor XOR2 (N11227, N11200, N6006);
xor XOR2 (N11228, N11224, N2954);
buf BUF1 (N11229, N11218);
and AND4 (N11230, N11225, N336, N8965, N8146);
nand NAND3 (N11231, N11219, N9153, N9048);
and AND4 (N11232, N11197, N1187, N4178, N4889);
buf BUF1 (N11233, N11228);
not NOT1 (N11234, N11221);
nand NAND3 (N11235, N11226, N3817, N1350);
xor XOR2 (N11236, N11211, N4117);
and AND4 (N11237, N11227, N4672, N5646, N7431);
or OR2 (N11238, N11231, N4639);
buf BUF1 (N11239, N11220);
nand NAND3 (N11240, N11229, N4814, N7804);
and AND2 (N11241, N11239, N1570);
and AND2 (N11242, N11240, N5623);
and AND2 (N11243, N11241, N8766);
and AND3 (N11244, N11234, N7490, N7479);
not NOT1 (N11245, N11230);
nand NAND3 (N11246, N11242, N9836, N6747);
nor NOR4 (N11247, N11243, N3949, N11137, N8711);
not NOT1 (N11248, N11238);
nor NOR2 (N11249, N11244, N8823);
xor XOR2 (N11250, N11235, N8113);
nand NAND4 (N11251, N11232, N8047, N2007, N185);
buf BUF1 (N11252, N11248);
xor XOR2 (N11253, N11237, N1110);
or OR3 (N11254, N11249, N10174, N672);
or OR2 (N11255, N11246, N3020);
not NOT1 (N11256, N11255);
nand NAND4 (N11257, N11252, N6629, N2922, N3863);
nand NAND2 (N11258, N11257, N11044);
nand NAND4 (N11259, N11251, N5238, N431, N2534);
not NOT1 (N11260, N11236);
not NOT1 (N11261, N11256);
nand NAND3 (N11262, N11258, N3356, N7532);
buf BUF1 (N11263, N11260);
and AND4 (N11264, N11245, N2166, N10245, N6381);
and AND3 (N11265, N11264, N9427, N785);
not NOT1 (N11266, N11261);
nor NOR3 (N11267, N11253, N11123, N2767);
and AND4 (N11268, N11254, N2353, N6463, N5180);
xor XOR2 (N11269, N11247, N9086);
nand NAND3 (N11270, N11259, N3698, N2167);
nand NAND2 (N11271, N11233, N4123);
buf BUF1 (N11272, N11265);
not NOT1 (N11273, N11266);
xor XOR2 (N11274, N11270, N1861);
or OR2 (N11275, N11268, N6331);
nand NAND4 (N11276, N11274, N5026, N9232, N1273);
nor NOR2 (N11277, N11263, N8121);
xor XOR2 (N11278, N11271, N8248);
nor NOR4 (N11279, N11262, N6496, N11084, N2811);
or OR3 (N11280, N11250, N6056, N9935);
not NOT1 (N11281, N11277);
xor XOR2 (N11282, N11280, N2319);
and AND4 (N11283, N11276, N1856, N1926, N8906);
not NOT1 (N11284, N11267);
not NOT1 (N11285, N11282);
and AND2 (N11286, N11285, N4762);
buf BUF1 (N11287, N11275);
or OR4 (N11288, N11279, N2582, N11076, N351);
nand NAND4 (N11289, N11284, N8830, N562, N9228);
not NOT1 (N11290, N11272);
buf BUF1 (N11291, N11287);
or OR3 (N11292, N11289, N9275, N7466);
buf BUF1 (N11293, N11269);
buf BUF1 (N11294, N11278);
xor XOR2 (N11295, N11293, N1566);
or OR4 (N11296, N11281, N5964, N5743, N4865);
nand NAND4 (N11297, N11290, N3948, N10950, N8808);
nor NOR3 (N11298, N11286, N9902, N3918);
buf BUF1 (N11299, N11291);
and AND2 (N11300, N11294, N6282);
nor NOR2 (N11301, N11292, N6540);
nand NAND3 (N11302, N11297, N2185, N4289);
buf BUF1 (N11303, N11273);
or OR2 (N11304, N11301, N2624);
nand NAND3 (N11305, N11303, N7202, N469);
not NOT1 (N11306, N11295);
nand NAND3 (N11307, N11299, N9743, N10596);
nor NOR4 (N11308, N11300, N8703, N9677, N5364);
buf BUF1 (N11309, N11283);
xor XOR2 (N11310, N11306, N5726);
xor XOR2 (N11311, N11308, N11126);
buf BUF1 (N11312, N11288);
and AND2 (N11313, N11305, N100);
nand NAND4 (N11314, N11310, N7426, N7941, N9911);
nand NAND2 (N11315, N11313, N1580);
nor NOR4 (N11316, N11298, N5145, N493, N221);
nor NOR2 (N11317, N11311, N4390);
or OR4 (N11318, N11315, N1905, N7916, N10913);
nor NOR4 (N11319, N11317, N9046, N2944, N1759);
not NOT1 (N11320, N11312);
buf BUF1 (N11321, N11316);
xor XOR2 (N11322, N11321, N7141);
or OR4 (N11323, N11302, N4672, N2525, N8564);
buf BUF1 (N11324, N11314);
not NOT1 (N11325, N11319);
xor XOR2 (N11326, N11318, N887);
buf BUF1 (N11327, N11325);
not NOT1 (N11328, N11323);
xor XOR2 (N11329, N11307, N5370);
or OR2 (N11330, N11320, N324);
xor XOR2 (N11331, N11304, N838);
nor NOR3 (N11332, N11309, N6424, N1877);
not NOT1 (N11333, N11327);
nand NAND4 (N11334, N11332, N5952, N1619, N9726);
nand NAND2 (N11335, N11322, N9093);
buf BUF1 (N11336, N11335);
xor XOR2 (N11337, N11336, N1104);
xor XOR2 (N11338, N11326, N6027);
xor XOR2 (N11339, N11296, N2165);
nor NOR2 (N11340, N11337, N9786);
nand NAND2 (N11341, N11328, N1843);
and AND3 (N11342, N11340, N3459, N5561);
or OR3 (N11343, N11330, N3061, N10883);
xor XOR2 (N11344, N11329, N3056);
or OR2 (N11345, N11342, N6219);
nor NOR4 (N11346, N11338, N6439, N4916, N11175);
and AND4 (N11347, N11341, N3634, N7742, N8432);
xor XOR2 (N11348, N11334, N6001);
buf BUF1 (N11349, N11346);
and AND4 (N11350, N11348, N5110, N5665, N3115);
or OR4 (N11351, N11345, N11221, N3587, N10950);
nand NAND3 (N11352, N11347, N9762, N1020);
buf BUF1 (N11353, N11333);
and AND2 (N11354, N11353, N9412);
or OR2 (N11355, N11349, N10227);
or OR4 (N11356, N11339, N2916, N3070, N8505);
buf BUF1 (N11357, N11350);
nor NOR3 (N11358, N11356, N4902, N37);
buf BUF1 (N11359, N11358);
buf BUF1 (N11360, N11324);
or OR3 (N11361, N11352, N7945, N3866);
or OR2 (N11362, N11331, N5300);
not NOT1 (N11363, N11351);
xor XOR2 (N11364, N11359, N2800);
nor NOR2 (N11365, N11360, N7209);
xor XOR2 (N11366, N11344, N8251);
and AND2 (N11367, N11361, N3691);
xor XOR2 (N11368, N11366, N10919);
nand NAND3 (N11369, N11364, N7827, N3576);
nand NAND3 (N11370, N11369, N5153, N4220);
and AND4 (N11371, N11355, N45, N5964, N9052);
or OR4 (N11372, N11362, N100, N9519, N5036);
and AND3 (N11373, N11372, N4761, N10668);
buf BUF1 (N11374, N11357);
buf BUF1 (N11375, N11371);
nor NOR2 (N11376, N11370, N5171);
nor NOR3 (N11377, N11367, N5176, N6762);
buf BUF1 (N11378, N11368);
not NOT1 (N11379, N11374);
or OR2 (N11380, N11379, N9722);
or OR3 (N11381, N11363, N6069, N2023);
buf BUF1 (N11382, N11373);
not NOT1 (N11383, N11343);
not NOT1 (N11384, N11376);
and AND2 (N11385, N11377, N4043);
not NOT1 (N11386, N11381);
buf BUF1 (N11387, N11386);
not NOT1 (N11388, N11375);
nor NOR4 (N11389, N11365, N2745, N9222, N6361);
or OR4 (N11390, N11378, N4733, N4037, N5064);
nand NAND2 (N11391, N11389, N6966);
nand NAND4 (N11392, N11391, N5261, N1475, N574);
not NOT1 (N11393, N11385);
or OR4 (N11394, N11392, N7834, N3162, N8596);
not NOT1 (N11395, N11388);
buf BUF1 (N11396, N11383);
and AND4 (N11397, N11387, N2789, N3555, N2266);
nand NAND2 (N11398, N11397, N693);
xor XOR2 (N11399, N11394, N3331);
or OR2 (N11400, N11399, N6214);
nand NAND3 (N11401, N11380, N9685, N10670);
not NOT1 (N11402, N11384);
or OR2 (N11403, N11382, N1482);
or OR2 (N11404, N11400, N5794);
nor NOR3 (N11405, N11398, N1827, N572);
xor XOR2 (N11406, N11404, N146);
nor NOR3 (N11407, N11396, N6707, N724);
nor NOR2 (N11408, N11407, N6977);
nor NOR3 (N11409, N11406, N8542, N994);
not NOT1 (N11410, N11401);
nor NOR3 (N11411, N11393, N7883, N11276);
and AND2 (N11412, N11408, N10974);
and AND3 (N11413, N11390, N4734, N7530);
buf BUF1 (N11414, N11403);
xor XOR2 (N11415, N11412, N6446);
xor XOR2 (N11416, N11409, N7454);
and AND2 (N11417, N11354, N3700);
not NOT1 (N11418, N11410);
buf BUF1 (N11419, N11411);
not NOT1 (N11420, N11417);
and AND2 (N11421, N11419, N6004);
buf BUF1 (N11422, N11402);
xor XOR2 (N11423, N11415, N8764);
and AND3 (N11424, N11413, N1939, N59);
buf BUF1 (N11425, N11422);
or OR2 (N11426, N11423, N6402);
or OR2 (N11427, N11421, N1457);
nor NOR3 (N11428, N11424, N9888, N7780);
not NOT1 (N11429, N11426);
nor NOR4 (N11430, N11416, N3032, N6735, N1299);
xor XOR2 (N11431, N11414, N2597);
nand NAND2 (N11432, N11395, N8097);
buf BUF1 (N11433, N11428);
buf BUF1 (N11434, N11432);
xor XOR2 (N11435, N11431, N5478);
or OR2 (N11436, N11434, N8537);
and AND4 (N11437, N11420, N1297, N3446, N1684);
nand NAND4 (N11438, N11427, N2053, N9633, N664);
and AND2 (N11439, N11418, N4114);
not NOT1 (N11440, N11435);
buf BUF1 (N11441, N11430);
and AND4 (N11442, N11433, N7518, N369, N295);
xor XOR2 (N11443, N11439, N6985);
and AND3 (N11444, N11438, N2551, N7656);
and AND4 (N11445, N11405, N6335, N7392, N2525);
nor NOR3 (N11446, N11442, N10141, N8868);
or OR4 (N11447, N11425, N376, N4755, N3922);
not NOT1 (N11448, N11447);
and AND2 (N11449, N11437, N5483);
not NOT1 (N11450, N11445);
or OR4 (N11451, N11450, N7396, N10143, N5014);
xor XOR2 (N11452, N11451, N6438);
xor XOR2 (N11453, N11452, N5986);
xor XOR2 (N11454, N11441, N7655);
xor XOR2 (N11455, N11453, N5392);
xor XOR2 (N11456, N11448, N10191);
nor NOR3 (N11457, N11456, N2074, N10976);
nor NOR2 (N11458, N11429, N6981);
not NOT1 (N11459, N11449);
nor NOR3 (N11460, N11443, N9083, N4855);
xor XOR2 (N11461, N11454, N9242);
nand NAND2 (N11462, N11457, N2068);
nand NAND4 (N11463, N11458, N4013, N1327, N8196);
not NOT1 (N11464, N11436);
xor XOR2 (N11465, N11459, N11248);
not NOT1 (N11466, N11465);
and AND4 (N11467, N11444, N3910, N802, N6866);
buf BUF1 (N11468, N11464);
not NOT1 (N11469, N11468);
or OR2 (N11470, N11455, N5529);
or OR4 (N11471, N11462, N5316, N3575, N10969);
or OR4 (N11472, N11460, N643, N7920, N6784);
nand NAND3 (N11473, N11463, N3757, N2486);
or OR4 (N11474, N11471, N4891, N3725, N9945);
nor NOR2 (N11475, N11461, N6042);
nor NOR2 (N11476, N11469, N1465);
not NOT1 (N11477, N11474);
or OR3 (N11478, N11440, N6747, N1189);
nor NOR4 (N11479, N11473, N8169, N8414, N1586);
not NOT1 (N11480, N11477);
not NOT1 (N11481, N11476);
or OR2 (N11482, N11472, N6214);
xor XOR2 (N11483, N11482, N4589);
and AND2 (N11484, N11467, N11149);
nand NAND4 (N11485, N11470, N8486, N1057, N663);
nor NOR4 (N11486, N11485, N1718, N1772, N3535);
buf BUF1 (N11487, N11483);
xor XOR2 (N11488, N11475, N8225);
xor XOR2 (N11489, N11481, N5290);
xor XOR2 (N11490, N11488, N8325);
or OR2 (N11491, N11478, N617);
buf BUF1 (N11492, N11480);
or OR4 (N11493, N11446, N7619, N8459, N8395);
or OR3 (N11494, N11479, N6239, N580);
not NOT1 (N11495, N11492);
buf BUF1 (N11496, N11495);
xor XOR2 (N11497, N11489, N728);
not NOT1 (N11498, N11487);
xor XOR2 (N11499, N11498, N3405);
and AND3 (N11500, N11499, N10732, N6679);
nor NOR2 (N11501, N11484, N3716);
xor XOR2 (N11502, N11500, N9804);
or OR2 (N11503, N11501, N2697);
nor NOR3 (N11504, N11466, N5341, N7780);
nor NOR3 (N11505, N11504, N3111, N8050);
xor XOR2 (N11506, N11493, N1956);
nor NOR4 (N11507, N11502, N3494, N6974, N8517);
xor XOR2 (N11508, N11507, N5174);
nand NAND4 (N11509, N11490, N9097, N2879, N6982);
nand NAND3 (N11510, N11505, N8309, N4836);
xor XOR2 (N11511, N11506, N9423);
nand NAND4 (N11512, N11503, N5294, N6126, N1736);
buf BUF1 (N11513, N11491);
xor XOR2 (N11514, N11486, N7952);
nor NOR2 (N11515, N11510, N9871);
nor NOR4 (N11516, N11509, N4503, N3206, N3242);
nand NAND4 (N11517, N11513, N10986, N7774, N4663);
xor XOR2 (N11518, N11512, N2026);
nor NOR4 (N11519, N11516, N4861, N11489, N4322);
nand NAND4 (N11520, N11511, N9712, N5162, N10063);
buf BUF1 (N11521, N11515);
nand NAND2 (N11522, N11494, N558);
or OR4 (N11523, N11497, N10991, N10752, N3543);
buf BUF1 (N11524, N11496);
and AND3 (N11525, N11522, N10267, N7008);
and AND2 (N11526, N11517, N802);
nor NOR4 (N11527, N11524, N1071, N1736, N8472);
xor XOR2 (N11528, N11521, N9717);
buf BUF1 (N11529, N11523);
nand NAND2 (N11530, N11518, N6903);
xor XOR2 (N11531, N11530, N4874);
nor NOR4 (N11532, N11519, N8539, N2719, N1114);
and AND2 (N11533, N11520, N7947);
or OR2 (N11534, N11525, N2259);
buf BUF1 (N11535, N11526);
nor NOR3 (N11536, N11514, N7063, N708);
not NOT1 (N11537, N11533);
nor NOR3 (N11538, N11531, N9943, N3382);
or OR4 (N11539, N11536, N4863, N7159, N7484);
xor XOR2 (N11540, N11539, N8172);
xor XOR2 (N11541, N11537, N8437);
buf BUF1 (N11542, N11538);
xor XOR2 (N11543, N11528, N5262);
xor XOR2 (N11544, N11540, N4023);
xor XOR2 (N11545, N11532, N6229);
not NOT1 (N11546, N11545);
nor NOR2 (N11547, N11542, N5354);
nand NAND4 (N11548, N11547, N11078, N7880, N9468);
not NOT1 (N11549, N11548);
or OR2 (N11550, N11508, N6534);
buf BUF1 (N11551, N11550);
buf BUF1 (N11552, N11529);
not NOT1 (N11553, N11535);
xor XOR2 (N11554, N11527, N9469);
or OR2 (N11555, N11554, N5569);
not NOT1 (N11556, N11546);
nor NOR3 (N11557, N11551, N7600, N4997);
xor XOR2 (N11558, N11549, N7085);
xor XOR2 (N11559, N11553, N9558);
buf BUF1 (N11560, N11555);
nor NOR4 (N11561, N11559, N8444, N8461, N5340);
buf BUF1 (N11562, N11552);
and AND3 (N11563, N11557, N9698, N11370);
nand NAND4 (N11564, N11562, N7506, N93, N10068);
xor XOR2 (N11565, N11564, N2346);
and AND3 (N11566, N11543, N7361, N8901);
buf BUF1 (N11567, N11534);
or OR4 (N11568, N11565, N5292, N180, N3396);
and AND4 (N11569, N11541, N6481, N6049, N621);
not NOT1 (N11570, N11544);
nor NOR2 (N11571, N11560, N9471);
or OR3 (N11572, N11563, N5018, N8459);
nand NAND2 (N11573, N11572, N3396);
or OR2 (N11574, N11558, N11216);
nor NOR3 (N11575, N11574, N10779, N1679);
buf BUF1 (N11576, N11571);
buf BUF1 (N11577, N11566);
xor XOR2 (N11578, N11570, N8801);
nand NAND3 (N11579, N11569, N10811, N11351);
buf BUF1 (N11580, N11578);
buf BUF1 (N11581, N11576);
and AND2 (N11582, N11579, N8739);
and AND4 (N11583, N11577, N3597, N4677, N1555);
xor XOR2 (N11584, N11561, N4307);
not NOT1 (N11585, N11556);
nor NOR4 (N11586, N11585, N8057, N6866, N8988);
nor NOR2 (N11587, N11584, N9188);
and AND3 (N11588, N11583, N3477, N548);
nand NAND2 (N11589, N11588, N4610);
xor XOR2 (N11590, N11589, N370);
nand NAND4 (N11591, N11582, N10062, N10544, N9768);
buf BUF1 (N11592, N11581);
buf BUF1 (N11593, N11573);
or OR3 (N11594, N11590, N758, N240);
not NOT1 (N11595, N11568);
or OR4 (N11596, N11587, N3377, N6392, N2888);
or OR3 (N11597, N11567, N1821, N5416);
nor NOR4 (N11598, N11597, N7851, N1310, N2046);
and AND4 (N11599, N11580, N1728, N7037, N7463);
xor XOR2 (N11600, N11593, N2359);
nor NOR2 (N11601, N11595, N7171);
not NOT1 (N11602, N11586);
xor XOR2 (N11603, N11602, N2790);
or OR3 (N11604, N11594, N2314, N9786);
or OR2 (N11605, N11601, N1169);
or OR3 (N11606, N11596, N10073, N4832);
not NOT1 (N11607, N11575);
nor NOR4 (N11608, N11605, N10698, N10993, N9415);
nor NOR3 (N11609, N11604, N5301, N5652);
nand NAND4 (N11610, N11608, N4949, N2331, N7590);
not NOT1 (N11611, N11591);
not NOT1 (N11612, N11592);
buf BUF1 (N11613, N11600);
and AND4 (N11614, N11611, N5551, N6685, N7158);
not NOT1 (N11615, N11613);
xor XOR2 (N11616, N11615, N4798);
xor XOR2 (N11617, N11599, N8710);
nor NOR3 (N11618, N11617, N5453, N1576);
or OR3 (N11619, N11606, N9186, N2647);
xor XOR2 (N11620, N11598, N7099);
not NOT1 (N11621, N11616);
nor NOR4 (N11622, N11619, N27, N4272, N155);
buf BUF1 (N11623, N11622);
nand NAND4 (N11624, N11623, N4793, N2613, N8944);
nand NAND4 (N11625, N11607, N2476, N8892, N10802);
and AND4 (N11626, N11624, N6299, N11421, N9997);
and AND3 (N11627, N11612, N5521, N9365);
xor XOR2 (N11628, N11618, N3938);
buf BUF1 (N11629, N11621);
nand NAND4 (N11630, N11610, N9433, N5508, N2113);
and AND2 (N11631, N11629, N9937);
or OR3 (N11632, N11627, N4684, N10283);
xor XOR2 (N11633, N11614, N8247);
not NOT1 (N11634, N11632);
and AND2 (N11635, N11628, N5794);
nand NAND3 (N11636, N11609, N193, N7949);
nor NOR2 (N11637, N11633, N308);
or OR4 (N11638, N11620, N9911, N6087, N2349);
not NOT1 (N11639, N11626);
and AND4 (N11640, N11638, N3184, N11633, N6817);
nand NAND4 (N11641, N11634, N45, N6484, N1709);
nor NOR3 (N11642, N11625, N5522, N8845);
nor NOR4 (N11643, N11603, N1584, N2284, N157);
xor XOR2 (N11644, N11640, N6126);
not NOT1 (N11645, N11631);
not NOT1 (N11646, N11645);
nor NOR4 (N11647, N11639, N11344, N8070, N9541);
xor XOR2 (N11648, N11644, N6779);
buf BUF1 (N11649, N11647);
xor XOR2 (N11650, N11642, N5303);
xor XOR2 (N11651, N11637, N1395);
or OR3 (N11652, N11630, N9444, N9814);
nor NOR2 (N11653, N11648, N3670);
nand NAND3 (N11654, N11651, N5336, N10685);
nor NOR2 (N11655, N11652, N9971);
or OR4 (N11656, N11636, N2071, N5214, N10234);
nor NOR2 (N11657, N11654, N7719);
or OR3 (N11658, N11649, N11257, N6784);
xor XOR2 (N11659, N11656, N3724);
nor NOR2 (N11660, N11653, N10612);
xor XOR2 (N11661, N11646, N9146);
nor NOR2 (N11662, N11658, N6721);
and AND4 (N11663, N11655, N11030, N9894, N98);
buf BUF1 (N11664, N11643);
or OR3 (N11665, N11661, N4025, N8676);
nand NAND2 (N11666, N11660, N6914);
nor NOR2 (N11667, N11665, N11316);
nand NAND2 (N11668, N11662, N1685);
or OR3 (N11669, N11668, N354, N4817);
not NOT1 (N11670, N11659);
not NOT1 (N11671, N11650);
buf BUF1 (N11672, N11667);
nor NOR4 (N11673, N11663, N8123, N8165, N10241);
and AND4 (N11674, N11664, N10333, N53, N7388);
not NOT1 (N11675, N11670);
nand NAND4 (N11676, N11657, N6175, N689, N8839);
or OR2 (N11677, N11666, N8258);
not NOT1 (N11678, N11635);
or OR3 (N11679, N11674, N4095, N446);
nand NAND4 (N11680, N11672, N3032, N9665, N10639);
xor XOR2 (N11681, N11641, N5601);
buf BUF1 (N11682, N11680);
not NOT1 (N11683, N11678);
buf BUF1 (N11684, N11681);
and AND2 (N11685, N11673, N8243);
xor XOR2 (N11686, N11669, N4371);
not NOT1 (N11687, N11683);
nor NOR3 (N11688, N11684, N716, N5338);
nand NAND2 (N11689, N11671, N44);
and AND2 (N11690, N11685, N8019);
buf BUF1 (N11691, N11682);
and AND2 (N11692, N11677, N5305);
buf BUF1 (N11693, N11690);
or OR3 (N11694, N11691, N10819, N11546);
buf BUF1 (N11695, N11693);
xor XOR2 (N11696, N11675, N264);
and AND4 (N11697, N11679, N10066, N3895, N11545);
not NOT1 (N11698, N11687);
nor NOR4 (N11699, N11698, N4719, N8823, N6133);
nor NOR4 (N11700, N11699, N3404, N358, N3026);
or OR2 (N11701, N11686, N4643);
or OR2 (N11702, N11676, N3326);
not NOT1 (N11703, N11694);
xor XOR2 (N11704, N11697, N5703);
buf BUF1 (N11705, N11700);
nor NOR2 (N11706, N11701, N2597);
nand NAND2 (N11707, N11704, N9529);
or OR4 (N11708, N11688, N7980, N6545, N10745);
or OR3 (N11709, N11695, N3870, N8087);
not NOT1 (N11710, N11708);
buf BUF1 (N11711, N11702);
nor NOR3 (N11712, N11692, N7112, N678);
xor XOR2 (N11713, N11710, N8909);
nor NOR2 (N11714, N11706, N4373);
nor NOR3 (N11715, N11709, N7420, N3720);
buf BUF1 (N11716, N11703);
nor NOR4 (N11717, N11696, N8652, N1672, N9428);
not NOT1 (N11718, N11712);
xor XOR2 (N11719, N11716, N8345);
not NOT1 (N11720, N11711);
not NOT1 (N11721, N11689);
not NOT1 (N11722, N11719);
and AND3 (N11723, N11718, N9290, N7652);
nand NAND2 (N11724, N11714, N9850);
not NOT1 (N11725, N11717);
nand NAND4 (N11726, N11721, N8915, N10950, N2943);
nand NAND2 (N11727, N11723, N2642);
not NOT1 (N11728, N11707);
and AND3 (N11729, N11727, N781, N10078);
nor NOR4 (N11730, N11728, N4053, N10328, N7749);
xor XOR2 (N11731, N11726, N8730);
not NOT1 (N11732, N11724);
and AND3 (N11733, N11732, N3815, N9031);
not NOT1 (N11734, N11731);
not NOT1 (N11735, N11730);
buf BUF1 (N11736, N11722);
or OR3 (N11737, N11725, N11011, N8089);
xor XOR2 (N11738, N11735, N10508);
or OR2 (N11739, N11713, N3386);
nor NOR4 (N11740, N11733, N10758, N5995, N6715);
or OR4 (N11741, N11705, N9358, N8052, N1467);
xor XOR2 (N11742, N11739, N2325);
or OR3 (N11743, N11738, N4315, N7535);
buf BUF1 (N11744, N11720);
or OR4 (N11745, N11744, N5736, N7845, N1618);
buf BUF1 (N11746, N11729);
not NOT1 (N11747, N11741);
buf BUF1 (N11748, N11743);
buf BUF1 (N11749, N11748);
not NOT1 (N11750, N11715);
nor NOR2 (N11751, N11749, N9104);
not NOT1 (N11752, N11742);
nand NAND3 (N11753, N11740, N10046, N7100);
nor NOR4 (N11754, N11737, N2955, N3044, N8140);
or OR2 (N11755, N11754, N3667);
nor NOR4 (N11756, N11746, N6393, N4528, N10332);
not NOT1 (N11757, N11752);
nand NAND3 (N11758, N11755, N3527, N7261);
nand NAND4 (N11759, N11734, N10202, N5901, N8635);
nand NAND2 (N11760, N11750, N8687);
or OR4 (N11761, N11756, N10995, N6247, N7545);
nand NAND3 (N11762, N11759, N8427, N11313);
not NOT1 (N11763, N11753);
nor NOR4 (N11764, N11758, N8434, N9075, N7725);
buf BUF1 (N11765, N11747);
or OR3 (N11766, N11745, N11640, N4075);
xor XOR2 (N11767, N11757, N6234);
and AND4 (N11768, N11762, N290, N83, N1167);
and AND3 (N11769, N11765, N4239, N7429);
nor NOR4 (N11770, N11751, N10441, N682, N11306);
and AND4 (N11771, N11770, N4877, N11615, N7148);
buf BUF1 (N11772, N11767);
nand NAND4 (N11773, N11760, N5027, N10413, N10710);
xor XOR2 (N11774, N11766, N4894);
xor XOR2 (N11775, N11774, N5271);
buf BUF1 (N11776, N11763);
buf BUF1 (N11777, N11772);
nand NAND2 (N11778, N11761, N2833);
nor NOR4 (N11779, N11769, N5268, N3155, N10752);
xor XOR2 (N11780, N11736, N6785);
nor NOR3 (N11781, N11764, N9031, N5464);
and AND4 (N11782, N11776, N8878, N10775, N6800);
buf BUF1 (N11783, N11778);
nand NAND2 (N11784, N11773, N10020);
not NOT1 (N11785, N11777);
xor XOR2 (N11786, N11782, N4273);
or OR4 (N11787, N11785, N10757, N2319, N10298);
not NOT1 (N11788, N11771);
buf BUF1 (N11789, N11768);
not NOT1 (N11790, N11786);
buf BUF1 (N11791, N11780);
nand NAND3 (N11792, N11789, N5444, N7906);
or OR3 (N11793, N11781, N7455, N10454);
or OR2 (N11794, N11779, N8019);
nand NAND4 (N11795, N11784, N11672, N10670, N11699);
xor XOR2 (N11796, N11790, N1955);
not NOT1 (N11797, N11787);
or OR3 (N11798, N11775, N1792, N5481);
or OR3 (N11799, N11796, N7802, N1948);
and AND2 (N11800, N11793, N8826);
not NOT1 (N11801, N11800);
not NOT1 (N11802, N11788);
and AND4 (N11803, N11798, N4079, N11647, N11580);
and AND2 (N11804, N11797, N4722);
xor XOR2 (N11805, N11795, N8463);
buf BUF1 (N11806, N11803);
not NOT1 (N11807, N11792);
not NOT1 (N11808, N11804);
nand NAND2 (N11809, N11799, N9448);
and AND4 (N11810, N11809, N8197, N3102, N11744);
not NOT1 (N11811, N11810);
and AND4 (N11812, N11805, N10907, N8593, N8378);
not NOT1 (N11813, N11808);
or OR3 (N11814, N11811, N4311, N5844);
nand NAND4 (N11815, N11802, N7088, N11698, N3653);
nor NOR2 (N11816, N11812, N3812);
and AND2 (N11817, N11813, N11618);
and AND3 (N11818, N11801, N2240, N9473);
buf BUF1 (N11819, N11791);
and AND2 (N11820, N11783, N10493);
nor NOR4 (N11821, N11817, N6862, N10529, N2744);
buf BUF1 (N11822, N11818);
or OR2 (N11823, N11819, N4084);
or OR2 (N11824, N11820, N10109);
nand NAND3 (N11825, N11794, N1888, N1363);
nor NOR4 (N11826, N11807, N4419, N1828, N1482);
and AND3 (N11827, N11823, N7724, N9805);
xor XOR2 (N11828, N11822, N1882);
not NOT1 (N11829, N11821);
nand NAND4 (N11830, N11806, N1703, N5229, N111);
not NOT1 (N11831, N11815);
xor XOR2 (N11832, N11830, N1643);
buf BUF1 (N11833, N11826);
nor NOR3 (N11834, N11831, N7055, N3462);
or OR3 (N11835, N11814, N4371, N3688);
or OR4 (N11836, N11833, N6724, N1180, N1856);
buf BUF1 (N11837, N11825);
and AND4 (N11838, N11828, N694, N6350, N10351);
and AND4 (N11839, N11829, N10769, N5891, N7357);
nor NOR2 (N11840, N11832, N9829);
and AND4 (N11841, N11838, N375, N9217, N3479);
not NOT1 (N11842, N11841);
or OR2 (N11843, N11836, N2955);
or OR3 (N11844, N11834, N4516, N6627);
buf BUF1 (N11845, N11840);
and AND3 (N11846, N11844, N10686, N939);
xor XOR2 (N11847, N11839, N6433);
buf BUF1 (N11848, N11837);
buf BUF1 (N11849, N11835);
xor XOR2 (N11850, N11827, N1960);
nor NOR3 (N11851, N11843, N4195, N11517);
and AND4 (N11852, N11850, N9310, N371, N3028);
buf BUF1 (N11853, N11849);
nand NAND2 (N11854, N11846, N10808);
not NOT1 (N11855, N11824);
buf BUF1 (N11856, N11854);
not NOT1 (N11857, N11842);
xor XOR2 (N11858, N11851, N1552);
not NOT1 (N11859, N11856);
xor XOR2 (N11860, N11816, N4382);
buf BUF1 (N11861, N11848);
xor XOR2 (N11862, N11861, N4007);
or OR3 (N11863, N11852, N8630, N980);
or OR2 (N11864, N11863, N6955);
buf BUF1 (N11865, N11859);
or OR2 (N11866, N11853, N555);
and AND4 (N11867, N11865, N8061, N6366, N2969);
xor XOR2 (N11868, N11855, N9724);
not NOT1 (N11869, N11860);
nand NAND4 (N11870, N11866, N3826, N5833, N9526);
not NOT1 (N11871, N11867);
xor XOR2 (N11872, N11869, N11215);
buf BUF1 (N11873, N11864);
nand NAND4 (N11874, N11845, N1007, N2567, N2791);
buf BUF1 (N11875, N11857);
and AND3 (N11876, N11873, N10573, N11342);
buf BUF1 (N11877, N11847);
nor NOR3 (N11878, N11872, N8641, N7411);
nor NOR2 (N11879, N11871, N157);
xor XOR2 (N11880, N11875, N8318);
not NOT1 (N11881, N11878);
not NOT1 (N11882, N11879);
or OR4 (N11883, N11870, N7939, N7299, N8400);
and AND2 (N11884, N11880, N3213);
nand NAND2 (N11885, N11862, N7738);
and AND4 (N11886, N11882, N7432, N8136, N5479);
nor NOR3 (N11887, N11883, N6082, N7377);
or OR4 (N11888, N11884, N2175, N10623, N5911);
nor NOR4 (N11889, N11876, N11460, N6812, N5677);
or OR3 (N11890, N11874, N9865, N8829);
nor NOR3 (N11891, N11868, N2284, N266);
nand NAND2 (N11892, N11888, N4415);
nand NAND3 (N11893, N11890, N10429, N576);
not NOT1 (N11894, N11881);
and AND3 (N11895, N11893, N1429, N3071);
nand NAND2 (N11896, N11886, N9808);
buf BUF1 (N11897, N11877);
not NOT1 (N11898, N11897);
buf BUF1 (N11899, N11889);
buf BUF1 (N11900, N11899);
nand NAND4 (N11901, N11858, N9184, N2023, N4915);
nand NAND2 (N11902, N11895, N11679);
or OR2 (N11903, N11894, N10628);
xor XOR2 (N11904, N11902, N7128);
buf BUF1 (N11905, N11901);
and AND4 (N11906, N11885, N7692, N6666, N9420);
nor NOR3 (N11907, N11891, N6734, N3395);
nor NOR2 (N11908, N11900, N5207);
not NOT1 (N11909, N11906);
or OR3 (N11910, N11903, N1017, N2124);
or OR3 (N11911, N11905, N10288, N1565);
or OR2 (N11912, N11887, N4002);
or OR3 (N11913, N11898, N2779, N5634);
and AND4 (N11914, N11912, N4247, N6317, N8195);
and AND2 (N11915, N11907, N4551);
nor NOR4 (N11916, N11896, N8351, N3730, N5864);
nand NAND2 (N11917, N11915, N2487);
nand NAND4 (N11918, N11911, N7615, N2799, N5110);
buf BUF1 (N11919, N11914);
nand NAND3 (N11920, N11917, N5053, N10199);
or OR2 (N11921, N11916, N8802);
not NOT1 (N11922, N11904);
nand NAND3 (N11923, N11919, N161, N11542);
and AND3 (N11924, N11908, N2664, N1525);
or OR3 (N11925, N11924, N4677, N9153);
nor NOR3 (N11926, N11913, N622, N6909);
buf BUF1 (N11927, N11926);
and AND3 (N11928, N11918, N7266, N3931);
not NOT1 (N11929, N11920);
nand NAND4 (N11930, N11910, N7343, N6246, N9121);
nand NAND4 (N11931, N11921, N10876, N5715, N7877);
not NOT1 (N11932, N11922);
xor XOR2 (N11933, N11925, N4710);
nand NAND3 (N11934, N11909, N6286, N1451);
or OR2 (N11935, N11923, N463);
nor NOR4 (N11936, N11931, N6975, N1996, N2589);
nand NAND2 (N11937, N11934, N10617);
buf BUF1 (N11938, N11937);
xor XOR2 (N11939, N11935, N9763);
or OR2 (N11940, N11936, N6733);
nor NOR4 (N11941, N11927, N9560, N10113, N6665);
xor XOR2 (N11942, N11930, N10451);
not NOT1 (N11943, N11941);
nor NOR3 (N11944, N11943, N2317, N11280);
and AND4 (N11945, N11932, N543, N810, N4864);
nand NAND3 (N11946, N11928, N6819, N3153);
not NOT1 (N11947, N11940);
xor XOR2 (N11948, N11946, N3300);
not NOT1 (N11949, N11939);
nor NOR3 (N11950, N11944, N4723, N5305);
not NOT1 (N11951, N11948);
or OR3 (N11952, N11929, N4013, N7270);
not NOT1 (N11953, N11942);
or OR4 (N11954, N11950, N5463, N8051, N8194);
not NOT1 (N11955, N11952);
xor XOR2 (N11956, N11947, N3497);
xor XOR2 (N11957, N11949, N9093);
buf BUF1 (N11958, N11945);
and AND2 (N11959, N11892, N5059);
xor XOR2 (N11960, N11959, N11777);
buf BUF1 (N11961, N11938);
not NOT1 (N11962, N11960);
buf BUF1 (N11963, N11962);
and AND2 (N11964, N11954, N9789);
nand NAND4 (N11965, N11961, N3495, N2412, N3930);
xor XOR2 (N11966, N11965, N6509);
nand NAND2 (N11967, N11956, N3313);
xor XOR2 (N11968, N11955, N3756);
xor XOR2 (N11969, N11966, N10945);
nor NOR3 (N11970, N11958, N9117, N8904);
not NOT1 (N11971, N11951);
not NOT1 (N11972, N11967);
not NOT1 (N11973, N11972);
or OR2 (N11974, N11953, N6607);
buf BUF1 (N11975, N11974);
nand NAND4 (N11976, N11964, N4665, N10483, N5687);
buf BUF1 (N11977, N11957);
nand NAND4 (N11978, N11971, N7670, N11228, N5693);
nor NOR4 (N11979, N11933, N7657, N9907, N3175);
or OR4 (N11980, N11979, N980, N5615, N4021);
nor NOR3 (N11981, N11977, N344, N2380);
nor NOR2 (N11982, N11978, N4152);
and AND2 (N11983, N11969, N11734);
and AND2 (N11984, N11973, N1365);
not NOT1 (N11985, N11982);
and AND3 (N11986, N11975, N516, N1108);
xor XOR2 (N11987, N11968, N8568);
not NOT1 (N11988, N11981);
nor NOR2 (N11989, N11984, N6200);
or OR3 (N11990, N11987, N5033, N7529);
or OR4 (N11991, N11990, N366, N1838, N8916);
not NOT1 (N11992, N11976);
not NOT1 (N11993, N11989);
xor XOR2 (N11994, N11991, N4530);
buf BUF1 (N11995, N11993);
nand NAND2 (N11996, N11988, N5277);
and AND3 (N11997, N11963, N11201, N3390);
or OR2 (N11998, N11995, N5895);
xor XOR2 (N11999, N11998, N11319);
xor XOR2 (N12000, N11994, N6813);
buf BUF1 (N12001, N11986);
or OR3 (N12002, N11999, N1371, N10460);
nor NOR4 (N12003, N11992, N9574, N4313, N9034);
nor NOR3 (N12004, N12001, N9042, N6744);
not NOT1 (N12005, N12002);
nor NOR2 (N12006, N11980, N3271);
and AND3 (N12007, N12004, N2801, N2837);
nand NAND4 (N12008, N11983, N4507, N3567, N4998);
or OR3 (N12009, N12006, N10002, N2947);
or OR2 (N12010, N11970, N3144);
nor NOR3 (N12011, N11985, N6112, N1074);
and AND3 (N12012, N12010, N9816, N6137);
or OR4 (N12013, N12000, N2008, N10841, N967);
buf BUF1 (N12014, N12012);
xor XOR2 (N12015, N12005, N11894);
and AND2 (N12016, N12015, N10866);
not NOT1 (N12017, N12007);
xor XOR2 (N12018, N12017, N7681);
and AND2 (N12019, N12011, N8819);
not NOT1 (N12020, N12019);
xor XOR2 (N12021, N12016, N5021);
xor XOR2 (N12022, N12018, N11358);
buf BUF1 (N12023, N12008);
nand NAND4 (N12024, N12021, N330, N10679, N10170);
and AND3 (N12025, N12014, N4682, N8397);
buf BUF1 (N12026, N12009);
xor XOR2 (N12027, N12013, N4253);
nand NAND4 (N12028, N12023, N4423, N10359, N6933);
xor XOR2 (N12029, N12025, N10296);
or OR4 (N12030, N12024, N9145, N11755, N6236);
not NOT1 (N12031, N11996);
xor XOR2 (N12032, N12022, N1985);
buf BUF1 (N12033, N12003);
not NOT1 (N12034, N12027);
not NOT1 (N12035, N12032);
xor XOR2 (N12036, N12031, N5923);
nand NAND3 (N12037, N12035, N2289, N8126);
not NOT1 (N12038, N12030);
nand NAND2 (N12039, N12020, N3551);
buf BUF1 (N12040, N12038);
not NOT1 (N12041, N12037);
not NOT1 (N12042, N12039);
nand NAND3 (N12043, N12042, N6990, N4924);
not NOT1 (N12044, N12026);
and AND3 (N12045, N11997, N1195, N225);
nand NAND3 (N12046, N12043, N8169, N3182);
or OR3 (N12047, N12045, N10028, N6523);
and AND4 (N12048, N12028, N6841, N7492, N11401);
nand NAND3 (N12049, N12047, N11515, N2298);
xor XOR2 (N12050, N12046, N11223);
buf BUF1 (N12051, N12044);
xor XOR2 (N12052, N12029, N11571);
or OR2 (N12053, N12033, N4033);
or OR3 (N12054, N12041, N10578, N431);
not NOT1 (N12055, N12050);
nand NAND2 (N12056, N12051, N10676);
or OR4 (N12057, N12056, N9470, N5149, N4372);
buf BUF1 (N12058, N12053);
nor NOR3 (N12059, N12054, N346, N10681);
or OR4 (N12060, N12058, N9798, N2837, N4475);
nand NAND3 (N12061, N12040, N4803, N7636);
nor NOR2 (N12062, N12049, N7602);
xor XOR2 (N12063, N12055, N4918);
xor XOR2 (N12064, N12057, N11439);
and AND3 (N12065, N12064, N3555, N5093);
xor XOR2 (N12066, N12060, N9031);
not NOT1 (N12067, N12036);
or OR2 (N12068, N12062, N891);
and AND3 (N12069, N12061, N2527, N6212);
not NOT1 (N12070, N12066);
xor XOR2 (N12071, N12067, N10239);
and AND3 (N12072, N12063, N7163, N8312);
nand NAND2 (N12073, N12071, N4983);
nor NOR4 (N12074, N12073, N857, N2531, N11159);
nand NAND2 (N12075, N12065, N9805);
not NOT1 (N12076, N12059);
not NOT1 (N12077, N12072);
or OR2 (N12078, N12048, N11670);
nor NOR4 (N12079, N12075, N4037, N8910, N10198);
and AND4 (N12080, N12034, N1544, N5004, N10435);
nand NAND4 (N12081, N12069, N11862, N6865, N1516);
xor XOR2 (N12082, N12080, N1374);
and AND2 (N12083, N12082, N6585);
xor XOR2 (N12084, N12070, N5849);
not NOT1 (N12085, N12084);
or OR2 (N12086, N12078, N2548);
nor NOR3 (N12087, N12083, N3089, N8733);
or OR3 (N12088, N12077, N5247, N11366);
xor XOR2 (N12089, N12052, N6810);
not NOT1 (N12090, N12085);
nor NOR2 (N12091, N12088, N7747);
not NOT1 (N12092, N12087);
nand NAND2 (N12093, N12081, N1016);
not NOT1 (N12094, N12076);
xor XOR2 (N12095, N12091, N9270);
or OR2 (N12096, N12079, N8669);
not NOT1 (N12097, N12094);
xor XOR2 (N12098, N12074, N11535);
and AND3 (N12099, N12098, N10688, N11086);
buf BUF1 (N12100, N12086);
not NOT1 (N12101, N12090);
not NOT1 (N12102, N12093);
nand NAND4 (N12103, N12102, N6428, N10918, N4011);
xor XOR2 (N12104, N12101, N9806);
nand NAND4 (N12105, N12068, N7354, N7358, N6094);
buf BUF1 (N12106, N12097);
or OR3 (N12107, N12089, N10463, N410);
buf BUF1 (N12108, N12100);
and AND4 (N12109, N12103, N4741, N6199, N7282);
xor XOR2 (N12110, N12092, N1272);
not NOT1 (N12111, N12108);
not NOT1 (N12112, N12099);
or OR3 (N12113, N12095, N6490, N365);
or OR4 (N12114, N12096, N5682, N4207, N10118);
and AND3 (N12115, N12113, N6173, N6520);
nor NOR3 (N12116, N12109, N5738, N10815);
nor NOR2 (N12117, N12111, N4479);
not NOT1 (N12118, N12112);
not NOT1 (N12119, N12117);
and AND4 (N12120, N12119, N2016, N8306, N8509);
nand NAND2 (N12121, N12110, N879);
xor XOR2 (N12122, N12121, N5335);
and AND4 (N12123, N12122, N7068, N9318, N1945);
buf BUF1 (N12124, N12105);
and AND3 (N12125, N12114, N4437, N3353);
nand NAND2 (N12126, N12106, N6354);
buf BUF1 (N12127, N12123);
or OR4 (N12128, N12126, N4419, N8258, N187);
nor NOR4 (N12129, N12127, N7439, N5882, N4353);
nor NOR4 (N12130, N12120, N6987, N878, N2709);
not NOT1 (N12131, N12130);
not NOT1 (N12132, N12115);
or OR4 (N12133, N12107, N11627, N8460, N7981);
nand NAND4 (N12134, N12125, N10571, N651, N2073);
xor XOR2 (N12135, N12134, N9758);
xor XOR2 (N12136, N12131, N2644);
not NOT1 (N12137, N12129);
buf BUF1 (N12138, N12104);
and AND4 (N12139, N12124, N4233, N4205, N10189);
not NOT1 (N12140, N12135);
xor XOR2 (N12141, N12139, N493);
not NOT1 (N12142, N12118);
nand NAND2 (N12143, N12142, N7795);
xor XOR2 (N12144, N12138, N3611);
or OR4 (N12145, N12133, N5302, N3747, N3190);
buf BUF1 (N12146, N12143);
buf BUF1 (N12147, N12145);
or OR4 (N12148, N12147, N2986, N10932, N10927);
not NOT1 (N12149, N12136);
xor XOR2 (N12150, N12141, N6136);
not NOT1 (N12151, N12132);
nor NOR2 (N12152, N12144, N5449);
or OR3 (N12153, N12151, N10319, N8073);
nand NAND2 (N12154, N12148, N4256);
nand NAND4 (N12155, N12140, N10886, N4059, N5187);
and AND3 (N12156, N12155, N3771, N179);
xor XOR2 (N12157, N12137, N3449);
or OR4 (N12158, N12128, N9267, N8675, N11756);
buf BUF1 (N12159, N12146);
and AND3 (N12160, N12149, N5912, N8145);
or OR4 (N12161, N12157, N2068, N6832, N62);
nor NOR4 (N12162, N12153, N2071, N5989, N703);
buf BUF1 (N12163, N12156);
nor NOR2 (N12164, N12154, N11477);
buf BUF1 (N12165, N12159);
not NOT1 (N12166, N12163);
nand NAND2 (N12167, N12165, N7022);
buf BUF1 (N12168, N12150);
nor NOR4 (N12169, N12166, N11933, N5369, N4551);
nor NOR3 (N12170, N12158, N5723, N9085);
not NOT1 (N12171, N12164);
nor NOR3 (N12172, N12167, N3913, N9756);
nor NOR4 (N12173, N12168, N11832, N1584, N2964);
and AND2 (N12174, N12160, N4615);
nor NOR4 (N12175, N12152, N8119, N11987, N4504);
xor XOR2 (N12176, N12171, N7508);
nand NAND4 (N12177, N12174, N11837, N7963, N7720);
xor XOR2 (N12178, N12173, N11742);
and AND4 (N12179, N12176, N10133, N6148, N2354);
nor NOR3 (N12180, N12161, N2327, N3710);
xor XOR2 (N12181, N12179, N8030);
buf BUF1 (N12182, N12175);
and AND3 (N12183, N12169, N4467, N8989);
buf BUF1 (N12184, N12177);
xor XOR2 (N12185, N12183, N1784);
not NOT1 (N12186, N12116);
not NOT1 (N12187, N12185);
or OR3 (N12188, N12178, N11830, N8072);
not NOT1 (N12189, N12187);
not NOT1 (N12190, N12188);
or OR3 (N12191, N12186, N3322, N2398);
nor NOR2 (N12192, N12184, N11283);
nand NAND3 (N12193, N12191, N1156, N1938);
nor NOR3 (N12194, N12192, N10490, N4316);
xor XOR2 (N12195, N12189, N3299);
nand NAND4 (N12196, N12193, N3071, N1948, N7917);
xor XOR2 (N12197, N12170, N10703);
not NOT1 (N12198, N12195);
not NOT1 (N12199, N12197);
buf BUF1 (N12200, N12194);
and AND4 (N12201, N12198, N985, N5212, N321);
or OR2 (N12202, N12196, N982);
nand NAND2 (N12203, N12190, N11655);
and AND3 (N12204, N12202, N6126, N8575);
or OR2 (N12205, N12180, N5959);
and AND3 (N12206, N12181, N11804, N346);
not NOT1 (N12207, N12206);
buf BUF1 (N12208, N12201);
or OR3 (N12209, N12182, N2094, N4428);
and AND2 (N12210, N12199, N3764);
nand NAND3 (N12211, N12204, N11746, N3036);
not NOT1 (N12212, N12207);
xor XOR2 (N12213, N12205, N2389);
buf BUF1 (N12214, N12211);
xor XOR2 (N12215, N12200, N6620);
nor NOR4 (N12216, N12162, N10905, N10899, N11655);
nor NOR2 (N12217, N12208, N9737);
nand NAND3 (N12218, N12212, N10897, N8298);
or OR4 (N12219, N12210, N2154, N7304, N7146);
or OR4 (N12220, N12216, N2379, N2292, N2363);
and AND3 (N12221, N12218, N6809, N2905);
or OR4 (N12222, N12172, N4251, N4449, N1240);
not NOT1 (N12223, N12213);
nor NOR3 (N12224, N12214, N8317, N507);
nand NAND2 (N12225, N12215, N8577);
nand NAND2 (N12226, N12220, N6740);
buf BUF1 (N12227, N12221);
and AND4 (N12228, N12226, N10212, N3959, N1074);
and AND2 (N12229, N12228, N1238);
not NOT1 (N12230, N12222);
not NOT1 (N12231, N12217);
nor NOR3 (N12232, N12209, N10508, N1896);
or OR2 (N12233, N12232, N4135);
xor XOR2 (N12234, N12233, N6270);
and AND3 (N12235, N12229, N9575, N1840);
and AND3 (N12236, N12223, N1925, N185);
xor XOR2 (N12237, N12203, N5697);
nor NOR2 (N12238, N12219, N4912);
buf BUF1 (N12239, N12236);
and AND3 (N12240, N12238, N5286, N11714);
buf BUF1 (N12241, N12239);
buf BUF1 (N12242, N12235);
or OR4 (N12243, N12237, N2507, N11056, N11546);
or OR2 (N12244, N12230, N976);
xor XOR2 (N12245, N12243, N8132);
and AND3 (N12246, N12244, N5754, N4349);
not NOT1 (N12247, N12246);
xor XOR2 (N12248, N12241, N11657);
not NOT1 (N12249, N12248);
buf BUF1 (N12250, N12242);
nand NAND4 (N12251, N12231, N8703, N1365, N11571);
and AND3 (N12252, N12249, N1233, N2552);
nand NAND3 (N12253, N12252, N11387, N9129);
nor NOR4 (N12254, N12227, N3094, N1328, N2942);
nand NAND4 (N12255, N12251, N873, N8042, N9326);
nor NOR2 (N12256, N12255, N4956);
nor NOR2 (N12257, N12234, N5442);
buf BUF1 (N12258, N12240);
and AND2 (N12259, N12256, N1678);
xor XOR2 (N12260, N12259, N6857);
or OR2 (N12261, N12225, N9753);
xor XOR2 (N12262, N12261, N10124);
buf BUF1 (N12263, N12260);
nor NOR2 (N12264, N12254, N3431);
and AND2 (N12265, N12247, N4577);
and AND3 (N12266, N12263, N1383, N9781);
not NOT1 (N12267, N12264);
nand NAND3 (N12268, N12265, N1034, N4469);
and AND4 (N12269, N12250, N2080, N9917, N8880);
or OR3 (N12270, N12267, N2011, N8857);
nor NOR4 (N12271, N12262, N3662, N8027, N2009);
and AND4 (N12272, N12270, N7402, N6300, N1711);
and AND4 (N12273, N12266, N2798, N7930, N4314);
buf BUF1 (N12274, N12272);
nor NOR3 (N12275, N12257, N10056, N3418);
and AND3 (N12276, N12275, N3099, N6699);
and AND2 (N12277, N12271, N9321);
xor XOR2 (N12278, N12276, N10136);
and AND3 (N12279, N12258, N8158, N2581);
not NOT1 (N12280, N12278);
not NOT1 (N12281, N12279);
buf BUF1 (N12282, N12280);
or OR3 (N12283, N12245, N580, N11668);
xor XOR2 (N12284, N12268, N6676);
nor NOR3 (N12285, N12283, N8371, N1975);
xor XOR2 (N12286, N12277, N2931);
not NOT1 (N12287, N12285);
buf BUF1 (N12288, N12253);
or OR3 (N12289, N12269, N11586, N2511);
nand NAND3 (N12290, N12284, N4576, N9389);
nand NAND3 (N12291, N12273, N5296, N5952);
nand NAND4 (N12292, N12288, N9316, N10514, N3865);
not NOT1 (N12293, N12282);
nand NAND3 (N12294, N12286, N1230, N9529);
or OR4 (N12295, N12292, N6769, N8590, N8519);
not NOT1 (N12296, N12290);
nor NOR4 (N12297, N12287, N11376, N2442, N2277);
and AND4 (N12298, N12295, N3350, N11356, N1776);
nor NOR2 (N12299, N12298, N2907);
or OR3 (N12300, N12293, N6400, N8498);
nand NAND2 (N12301, N12296, N11820);
and AND3 (N12302, N12224, N5638, N259);
buf BUF1 (N12303, N12297);
not NOT1 (N12304, N12281);
nand NAND2 (N12305, N12291, N8591);
and AND3 (N12306, N12303, N3162, N1584);
and AND2 (N12307, N12306, N5567);
buf BUF1 (N12308, N12302);
or OR3 (N12309, N12294, N3603, N5985);
not NOT1 (N12310, N12289);
and AND4 (N12311, N12304, N7394, N9817, N4749);
not NOT1 (N12312, N12299);
and AND3 (N12313, N12308, N2655, N7711);
not NOT1 (N12314, N12300);
and AND3 (N12315, N12312, N7244, N2125);
xor XOR2 (N12316, N12307, N2007);
not NOT1 (N12317, N12301);
and AND2 (N12318, N12317, N104);
not NOT1 (N12319, N12310);
buf BUF1 (N12320, N12315);
xor XOR2 (N12321, N12320, N757);
or OR4 (N12322, N12314, N4542, N7599, N2008);
xor XOR2 (N12323, N12309, N5506);
or OR4 (N12324, N12305, N10323, N962, N4141);
and AND2 (N12325, N12322, N5237);
nand NAND2 (N12326, N12324, N9353);
buf BUF1 (N12327, N12274);
nand NAND4 (N12328, N12318, N9570, N4919, N2837);
xor XOR2 (N12329, N12328, N7834);
buf BUF1 (N12330, N12321);
buf BUF1 (N12331, N12319);
nand NAND2 (N12332, N12325, N8454);
nand NAND2 (N12333, N12327, N5830);
xor XOR2 (N12334, N12331, N11570);
nor NOR2 (N12335, N12316, N8328);
xor XOR2 (N12336, N12313, N8940);
nand NAND2 (N12337, N12326, N7781);
and AND3 (N12338, N12330, N797, N53);
nor NOR2 (N12339, N12311, N10490);
nand NAND2 (N12340, N12337, N10957);
or OR3 (N12341, N12329, N2726, N5938);
xor XOR2 (N12342, N12336, N8249);
not NOT1 (N12343, N12334);
xor XOR2 (N12344, N12333, N2170);
not NOT1 (N12345, N12342);
nand NAND4 (N12346, N12335, N6918, N10859, N4571);
nor NOR3 (N12347, N12338, N1034, N7910);
buf BUF1 (N12348, N12345);
not NOT1 (N12349, N12347);
and AND3 (N12350, N12349, N1946, N11394);
buf BUF1 (N12351, N12348);
buf BUF1 (N12352, N12340);
nor NOR2 (N12353, N12352, N8110);
xor XOR2 (N12354, N12341, N1608);
or OR4 (N12355, N12351, N8875, N2697, N9127);
not NOT1 (N12356, N12332);
buf BUF1 (N12357, N12346);
buf BUF1 (N12358, N12355);
xor XOR2 (N12359, N12344, N3551);
not NOT1 (N12360, N12353);
nand NAND3 (N12361, N12354, N7663, N3112);
buf BUF1 (N12362, N12323);
xor XOR2 (N12363, N12360, N9855);
or OR3 (N12364, N12343, N7012, N764);
or OR2 (N12365, N12359, N5348);
xor XOR2 (N12366, N12356, N2652);
or OR3 (N12367, N12339, N10999, N2781);
nand NAND2 (N12368, N12365, N2972);
nand NAND3 (N12369, N12366, N8990, N9906);
buf BUF1 (N12370, N12364);
or OR4 (N12371, N12350, N10997, N7277, N10064);
and AND4 (N12372, N12370, N10320, N3533, N1712);
nand NAND4 (N12373, N12357, N8795, N7869, N2852);
buf BUF1 (N12374, N12362);
buf BUF1 (N12375, N12373);
and AND4 (N12376, N12358, N2288, N1721, N3453);
buf BUF1 (N12377, N12361);
nor NOR4 (N12378, N12363, N3029, N6188, N2089);
and AND2 (N12379, N12377, N7122);
and AND2 (N12380, N12374, N8064);
nor NOR4 (N12381, N12378, N8849, N968, N745);
nor NOR4 (N12382, N12368, N9149, N7754, N9569);
not NOT1 (N12383, N12372);
nand NAND3 (N12384, N12381, N5778, N9982);
xor XOR2 (N12385, N12382, N7973);
nor NOR3 (N12386, N12380, N1723, N4479);
or OR4 (N12387, N12367, N804, N7037, N6727);
xor XOR2 (N12388, N12379, N2531);
xor XOR2 (N12389, N12371, N3363);
not NOT1 (N12390, N12385);
buf BUF1 (N12391, N12388);
xor XOR2 (N12392, N12375, N2202);
or OR3 (N12393, N12383, N10573, N11393);
buf BUF1 (N12394, N12387);
and AND2 (N12395, N12394, N6793);
or OR3 (N12396, N12376, N7018, N224);
or OR3 (N12397, N12390, N5669, N7321);
or OR2 (N12398, N12384, N3427);
or OR2 (N12399, N12395, N814);
or OR4 (N12400, N12392, N8948, N12066, N1852);
nor NOR4 (N12401, N12391, N619, N11082, N4177);
buf BUF1 (N12402, N12400);
nand NAND3 (N12403, N12397, N7272, N11139);
xor XOR2 (N12404, N12399, N2062);
and AND3 (N12405, N12401, N9554, N2536);
and AND3 (N12406, N12402, N1524, N4566);
xor XOR2 (N12407, N12369, N11825);
xor XOR2 (N12408, N12406, N11016);
buf BUF1 (N12409, N12389);
or OR4 (N12410, N12403, N10070, N5688, N2181);
nor NOR3 (N12411, N12408, N3390, N2467);
nand NAND4 (N12412, N12405, N528, N6752, N10871);
or OR3 (N12413, N12396, N7922, N576);
nor NOR2 (N12414, N12413, N10907);
nor NOR2 (N12415, N12393, N12135);
nor NOR2 (N12416, N12407, N6797);
and AND3 (N12417, N12414, N7036, N8181);
xor XOR2 (N12418, N12417, N1685);
nand NAND4 (N12419, N12416, N10798, N9746, N8889);
not NOT1 (N12420, N12409);
nor NOR4 (N12421, N12412, N5039, N12206, N4078);
or OR3 (N12422, N12411, N7482, N4597);
nor NOR2 (N12423, N12398, N7082);
xor XOR2 (N12424, N12386, N44);
xor XOR2 (N12425, N12418, N10324);
not NOT1 (N12426, N12415);
xor XOR2 (N12427, N12419, N10652);
and AND4 (N12428, N12426, N7658, N10352, N7094);
nor NOR2 (N12429, N12425, N8252);
or OR2 (N12430, N12421, N4554);
or OR4 (N12431, N12428, N9952, N4102, N316);
xor XOR2 (N12432, N12431, N10045);
buf BUF1 (N12433, N12420);
xor XOR2 (N12434, N12423, N5571);
buf BUF1 (N12435, N12424);
not NOT1 (N12436, N12427);
and AND3 (N12437, N12436, N8331, N3134);
xor XOR2 (N12438, N12422, N4889);
and AND4 (N12439, N12432, N5824, N8483, N5270);
and AND3 (N12440, N12437, N11609, N11033);
nand NAND4 (N12441, N12438, N10441, N10316, N8964);
nand NAND2 (N12442, N12433, N746);
xor XOR2 (N12443, N12430, N9189);
and AND3 (N12444, N12441, N12132, N3599);
not NOT1 (N12445, N12410);
xor XOR2 (N12446, N12442, N12347);
buf BUF1 (N12447, N12434);
buf BUF1 (N12448, N12404);
xor XOR2 (N12449, N12440, N3318);
or OR2 (N12450, N12445, N7205);
and AND4 (N12451, N12447, N192, N9317, N9098);
xor XOR2 (N12452, N12429, N3059);
buf BUF1 (N12453, N12435);
nor NOR4 (N12454, N12449, N8096, N3246, N79);
xor XOR2 (N12455, N12446, N2067);
or OR3 (N12456, N12450, N2906, N6203);
xor XOR2 (N12457, N12454, N10780);
nor NOR3 (N12458, N12439, N4771, N1737);
or OR4 (N12459, N12451, N9, N5631, N3251);
and AND3 (N12460, N12459, N11510, N10186);
xor XOR2 (N12461, N12457, N2887);
or OR2 (N12462, N12452, N7096);
xor XOR2 (N12463, N12460, N9989);
nand NAND2 (N12464, N12461, N5052);
nand NAND4 (N12465, N12462, N7247, N2953, N2196);
buf BUF1 (N12466, N12443);
xor XOR2 (N12467, N12456, N6282);
xor XOR2 (N12468, N12466, N5478);
or OR2 (N12469, N12458, N802);
nor NOR2 (N12470, N12444, N8319);
buf BUF1 (N12471, N12455);
xor XOR2 (N12472, N12470, N7388);
xor XOR2 (N12473, N12469, N1349);
buf BUF1 (N12474, N12448);
nand NAND3 (N12475, N12453, N5428, N10005);
nor NOR3 (N12476, N12475, N2170, N5282);
or OR3 (N12477, N12464, N1859, N11054);
xor XOR2 (N12478, N12467, N8519);
not NOT1 (N12479, N12473);
or OR3 (N12480, N12477, N3767, N6321);
nand NAND2 (N12481, N12474, N4277);
and AND2 (N12482, N12468, N12189);
buf BUF1 (N12483, N12465);
xor XOR2 (N12484, N12471, N1894);
nor NOR3 (N12485, N12480, N5976, N1697);
not NOT1 (N12486, N12484);
buf BUF1 (N12487, N12478);
not NOT1 (N12488, N12463);
xor XOR2 (N12489, N12483, N11275);
and AND3 (N12490, N12486, N3974, N12261);
nand NAND2 (N12491, N12487, N3379);
nor NOR4 (N12492, N12479, N11152, N10385, N10268);
not NOT1 (N12493, N12491);
xor XOR2 (N12494, N12482, N1274);
nand NAND4 (N12495, N12472, N2495, N2417, N7850);
nand NAND4 (N12496, N12489, N7335, N10034, N12222);
or OR4 (N12497, N12488, N10385, N5614, N592);
not NOT1 (N12498, N12496);
or OR4 (N12499, N12476, N9254, N6102, N1261);
buf BUF1 (N12500, N12494);
nand NAND4 (N12501, N12493, N2187, N6463, N551);
not NOT1 (N12502, N12500);
and AND2 (N12503, N12501, N4676);
or OR2 (N12504, N12499, N3935);
or OR2 (N12505, N12503, N4960);
xor XOR2 (N12506, N12497, N2033);
or OR2 (N12507, N12485, N7851);
and AND3 (N12508, N12504, N11759, N3689);
and AND4 (N12509, N12498, N9174, N5693, N11538);
not NOT1 (N12510, N12490);
xor XOR2 (N12511, N12510, N4128);
buf BUF1 (N12512, N12492);
or OR4 (N12513, N12509, N6329, N10869, N8077);
or OR2 (N12514, N12508, N2237);
and AND4 (N12515, N12502, N1640, N9641, N5951);
nand NAND3 (N12516, N12495, N4784, N8877);
nor NOR2 (N12517, N12507, N1396);
and AND2 (N12518, N12515, N2916);
nand NAND2 (N12519, N12481, N1371);
nand NAND2 (N12520, N12512, N1938);
nor NOR2 (N12521, N12505, N4921);
nand NAND2 (N12522, N12519, N10723);
not NOT1 (N12523, N12516);
nor NOR2 (N12524, N12514, N10571);
and AND4 (N12525, N12523, N11316, N10677, N11436);
buf BUF1 (N12526, N12517);
xor XOR2 (N12527, N12521, N8482);
nand NAND4 (N12528, N12513, N715, N9220, N1822);
or OR3 (N12529, N12525, N4529, N520);
nand NAND3 (N12530, N12520, N1059, N1271);
or OR4 (N12531, N12506, N1994, N4067, N12364);
buf BUF1 (N12532, N12526);
xor XOR2 (N12533, N12518, N313);
and AND3 (N12534, N12528, N4752, N4967);
nor NOR2 (N12535, N12511, N1467);
xor XOR2 (N12536, N12532, N7880);
or OR4 (N12537, N12536, N9749, N4375, N3633);
nor NOR4 (N12538, N12531, N1695, N4419, N5285);
buf BUF1 (N12539, N12538);
xor XOR2 (N12540, N12534, N1509);
and AND2 (N12541, N12524, N2020);
and AND4 (N12542, N12540, N9074, N2469, N2879);
or OR3 (N12543, N12535, N10036, N3160);
xor XOR2 (N12544, N12530, N8728);
nor NOR2 (N12545, N12543, N185);
not NOT1 (N12546, N12537);
or OR4 (N12547, N12542, N2042, N1496, N7305);
nor NOR3 (N12548, N12545, N10053, N5427);
nor NOR2 (N12549, N12548, N1600);
or OR2 (N12550, N12544, N6121);
and AND4 (N12551, N12546, N12504, N2950, N5201);
or OR4 (N12552, N12522, N2909, N4705, N10739);
and AND3 (N12553, N12533, N11329, N8951);
or OR2 (N12554, N12539, N115);
not NOT1 (N12555, N12554);
xor XOR2 (N12556, N12552, N8992);
buf BUF1 (N12557, N12529);
buf BUF1 (N12558, N12553);
not NOT1 (N12559, N12541);
or OR3 (N12560, N12549, N10639, N1465);
nor NOR3 (N12561, N12527, N2499, N1390);
nor NOR2 (N12562, N12561, N3860);
and AND3 (N12563, N12547, N5410, N9728);
nor NOR2 (N12564, N12555, N7735);
and AND3 (N12565, N12559, N97, N8229);
not NOT1 (N12566, N12562);
nand NAND3 (N12567, N12558, N10823, N10477);
or OR4 (N12568, N12560, N7539, N11156, N9908);
or OR2 (N12569, N12563, N3963);
xor XOR2 (N12570, N12556, N12244);
nand NAND3 (N12571, N12550, N3444, N11656);
and AND4 (N12572, N12569, N1449, N11532, N6505);
not NOT1 (N12573, N12571);
nand NAND2 (N12574, N12565, N8084);
xor XOR2 (N12575, N12568, N8474);
not NOT1 (N12576, N12574);
and AND3 (N12577, N12551, N12136, N4888);
nand NAND3 (N12578, N12576, N10742, N3380);
buf BUF1 (N12579, N12567);
xor XOR2 (N12580, N12564, N2319);
not NOT1 (N12581, N12577);
or OR2 (N12582, N12570, N2176);
or OR4 (N12583, N12582, N7349, N6914, N3310);
nand NAND3 (N12584, N12572, N6344, N567);
buf BUF1 (N12585, N12573);
buf BUF1 (N12586, N12584);
buf BUF1 (N12587, N12557);
not NOT1 (N12588, N12575);
nand NAND3 (N12589, N12578, N8456, N9891);
xor XOR2 (N12590, N12588, N9585);
not NOT1 (N12591, N12589);
not NOT1 (N12592, N12566);
and AND4 (N12593, N12585, N3724, N343, N2324);
or OR2 (N12594, N12590, N4656);
not NOT1 (N12595, N12587);
buf BUF1 (N12596, N12593);
not NOT1 (N12597, N12581);
nand NAND3 (N12598, N12583, N4060, N7168);
nor NOR3 (N12599, N12594, N9537, N6680);
xor XOR2 (N12600, N12595, N227);
xor XOR2 (N12601, N12599, N3007);
or OR2 (N12602, N12592, N12519);
buf BUF1 (N12603, N12596);
and AND2 (N12604, N12601, N9966);
or OR2 (N12605, N12586, N11105);
not NOT1 (N12606, N12604);
or OR4 (N12607, N12580, N4267, N11141, N3902);
and AND3 (N12608, N12579, N4863, N7354);
nand NAND4 (N12609, N12605, N1126, N7672, N7921);
not NOT1 (N12610, N12591);
or OR2 (N12611, N12608, N11357);
nand NAND3 (N12612, N12597, N2041, N12490);
nor NOR4 (N12613, N12606, N5032, N9462, N9030);
nor NOR4 (N12614, N12603, N834, N11441, N387);
buf BUF1 (N12615, N12614);
and AND2 (N12616, N12598, N2029);
xor XOR2 (N12617, N12610, N6064);
buf BUF1 (N12618, N12616);
or OR2 (N12619, N12612, N2480);
xor XOR2 (N12620, N12600, N5017);
and AND2 (N12621, N12613, N6064);
buf BUF1 (N12622, N12618);
not NOT1 (N12623, N12607);
not NOT1 (N12624, N12619);
xor XOR2 (N12625, N12611, N11631);
and AND3 (N12626, N12622, N6476, N10919);
nand NAND3 (N12627, N12625, N12405, N1875);
xor XOR2 (N12628, N12624, N7987);
or OR4 (N12629, N12617, N9352, N6044, N7236);
nand NAND2 (N12630, N12629, N9353);
or OR3 (N12631, N12628, N1336, N8319);
not NOT1 (N12632, N12620);
xor XOR2 (N12633, N12626, N11391);
xor XOR2 (N12634, N12630, N658);
not NOT1 (N12635, N12609);
or OR3 (N12636, N12602, N12443, N3229);
not NOT1 (N12637, N12635);
not NOT1 (N12638, N12634);
buf BUF1 (N12639, N12627);
nor NOR3 (N12640, N12633, N2532, N9010);
and AND3 (N12641, N12636, N8727, N201);
and AND2 (N12642, N12623, N315);
buf BUF1 (N12643, N12632);
xor XOR2 (N12644, N12621, N5309);
nor NOR3 (N12645, N12615, N8649, N6156);
xor XOR2 (N12646, N12645, N8172);
nor NOR3 (N12647, N12641, N10854, N2036);
xor XOR2 (N12648, N12639, N4953);
nand NAND3 (N12649, N12644, N8318, N6517);
nor NOR2 (N12650, N12640, N1331);
or OR2 (N12651, N12650, N2441);
and AND3 (N12652, N12637, N4763, N5681);
or OR3 (N12653, N12652, N248, N5966);
not NOT1 (N12654, N12631);
buf BUF1 (N12655, N12653);
buf BUF1 (N12656, N12638);
nor NOR2 (N12657, N12643, N597);
nor NOR2 (N12658, N12646, N4338);
xor XOR2 (N12659, N12656, N8177);
nor NOR2 (N12660, N12655, N438);
not NOT1 (N12661, N12660);
not NOT1 (N12662, N12648);
nand NAND3 (N12663, N12658, N10005, N7915);
nor NOR3 (N12664, N12662, N10125, N11161);
xor XOR2 (N12665, N12661, N1100);
nand NAND3 (N12666, N12663, N4305, N12512);
nor NOR4 (N12667, N12657, N12413, N8927, N12540);
buf BUF1 (N12668, N12659);
nor NOR2 (N12669, N12665, N7464);
nor NOR2 (N12670, N12647, N3128);
buf BUF1 (N12671, N12667);
nor NOR4 (N12672, N12649, N12500, N6325, N11905);
nor NOR4 (N12673, N12672, N5154, N1327, N12142);
not NOT1 (N12674, N12654);
buf BUF1 (N12675, N12671);
nand NAND2 (N12676, N12673, N9421);
not NOT1 (N12677, N12666);
or OR4 (N12678, N12651, N11878, N10172, N1761);
xor XOR2 (N12679, N12678, N3286);
nor NOR4 (N12680, N12676, N10459, N7864, N5534);
not NOT1 (N12681, N12642);
and AND3 (N12682, N12677, N884, N2530);
not NOT1 (N12683, N12674);
buf BUF1 (N12684, N12675);
not NOT1 (N12685, N12669);
not NOT1 (N12686, N12684);
not NOT1 (N12687, N12686);
nand NAND4 (N12688, N12664, N7959, N9589, N2190);
nor NOR2 (N12689, N12681, N6049);
nand NAND3 (N12690, N12687, N177, N6594);
xor XOR2 (N12691, N12685, N3039);
buf BUF1 (N12692, N12683);
not NOT1 (N12693, N12668);
or OR2 (N12694, N12691, N5312);
and AND3 (N12695, N12693, N3121, N1868);
not NOT1 (N12696, N12688);
and AND4 (N12697, N12692, N10474, N3859, N2323);
nor NOR3 (N12698, N12694, N1869, N4872);
xor XOR2 (N12699, N12695, N1028);
buf BUF1 (N12700, N12682);
nor NOR2 (N12701, N12698, N8294);
xor XOR2 (N12702, N12690, N7842);
nor NOR3 (N12703, N12670, N3921, N5268);
xor XOR2 (N12704, N12679, N5160);
nor NOR2 (N12705, N12701, N11079);
not NOT1 (N12706, N12703);
nor NOR3 (N12707, N12704, N4441, N7632);
xor XOR2 (N12708, N12707, N184);
xor XOR2 (N12709, N12680, N902);
and AND2 (N12710, N12709, N12377);
or OR4 (N12711, N12697, N12703, N806, N5849);
or OR4 (N12712, N12705, N6528, N4374, N5921);
buf BUF1 (N12713, N12708);
nand NAND2 (N12714, N12699, N9401);
or OR4 (N12715, N12700, N6034, N2681, N832);
not NOT1 (N12716, N12713);
or OR3 (N12717, N12702, N6996, N506);
xor XOR2 (N12718, N12717, N7410);
not NOT1 (N12719, N12696);
xor XOR2 (N12720, N12706, N9793);
not NOT1 (N12721, N12718);
nor NOR4 (N12722, N12689, N6804, N12019, N8965);
or OR2 (N12723, N12714, N10389);
not NOT1 (N12724, N12723);
xor XOR2 (N12725, N12722, N1205);
or OR2 (N12726, N12711, N7290);
nor NOR2 (N12727, N12715, N5480);
not NOT1 (N12728, N12712);
nand NAND4 (N12729, N12716, N9347, N7008, N12510);
nor NOR3 (N12730, N12728, N6731, N3223);
or OR2 (N12731, N12729, N8967);
buf BUF1 (N12732, N12720);
nor NOR3 (N12733, N12730, N7684, N245);
xor XOR2 (N12734, N12727, N9084);
and AND4 (N12735, N12724, N9602, N11210, N1023);
nor NOR4 (N12736, N12733, N751, N11668, N5808);
and AND4 (N12737, N12732, N2274, N131, N7602);
or OR4 (N12738, N12719, N5146, N5889, N11844);
not NOT1 (N12739, N12710);
xor XOR2 (N12740, N12736, N7094);
or OR4 (N12741, N12740, N3737, N11057, N1310);
nor NOR4 (N12742, N12739, N2234, N505, N4082);
nand NAND2 (N12743, N12725, N10697);
xor XOR2 (N12744, N12721, N5862);
or OR4 (N12745, N12726, N7176, N4502, N3142);
nand NAND2 (N12746, N12731, N4555);
or OR4 (N12747, N12734, N8108, N7889, N10484);
xor XOR2 (N12748, N12735, N574);
nor NOR3 (N12749, N12745, N2050, N4674);
and AND2 (N12750, N12748, N8681);
buf BUF1 (N12751, N12746);
nand NAND4 (N12752, N12741, N3183, N4892, N1445);
and AND2 (N12753, N12750, N12163);
nand NAND4 (N12754, N12749, N9789, N6420, N2788);
not NOT1 (N12755, N12747);
or OR3 (N12756, N12744, N6979, N5492);
buf BUF1 (N12757, N12752);
nor NOR4 (N12758, N12754, N3257, N11247, N3853);
buf BUF1 (N12759, N12757);
and AND4 (N12760, N12755, N7015, N1786, N10580);
or OR2 (N12761, N12738, N9613);
or OR4 (N12762, N12753, N2793, N8039, N9075);
nor NOR2 (N12763, N12751, N10593);
and AND2 (N12764, N12756, N10990);
and AND3 (N12765, N12761, N10508, N301);
nor NOR4 (N12766, N12742, N7932, N2925, N7814);
xor XOR2 (N12767, N12763, N2245);
buf BUF1 (N12768, N12759);
buf BUF1 (N12769, N12766);
xor XOR2 (N12770, N12769, N4741);
nand NAND2 (N12771, N12764, N6154);
and AND4 (N12772, N12765, N7198, N2350, N8487);
and AND2 (N12773, N12737, N11301);
not NOT1 (N12774, N12760);
nor NOR3 (N12775, N12762, N5894, N7312);
buf BUF1 (N12776, N12767);
buf BUF1 (N12777, N12768);
not NOT1 (N12778, N12743);
and AND3 (N12779, N12758, N2983, N10340);
xor XOR2 (N12780, N12776, N520);
nand NAND4 (N12781, N12774, N11437, N9306, N1766);
and AND2 (N12782, N12775, N5671);
xor XOR2 (N12783, N12782, N2720);
xor XOR2 (N12784, N12778, N1177);
not NOT1 (N12785, N12772);
nand NAND4 (N12786, N12785, N4876, N11688, N10757);
xor XOR2 (N12787, N12780, N1581);
nand NAND2 (N12788, N12783, N3357);
not NOT1 (N12789, N12771);
nand NAND2 (N12790, N12784, N6217);
nor NOR3 (N12791, N12786, N5872, N2737);
xor XOR2 (N12792, N12789, N7130);
and AND3 (N12793, N12790, N3483, N5925);
nor NOR2 (N12794, N12787, N2116);
not NOT1 (N12795, N12779);
nand NAND4 (N12796, N12770, N229, N10905, N2341);
buf BUF1 (N12797, N12796);
or OR2 (N12798, N12792, N7199);
or OR4 (N12799, N12794, N9034, N12671, N6238);
xor XOR2 (N12800, N12773, N10960);
nand NAND4 (N12801, N12798, N8665, N7002, N8555);
buf BUF1 (N12802, N12797);
xor XOR2 (N12803, N12777, N1145);
not NOT1 (N12804, N12793);
xor XOR2 (N12805, N12804, N1579);
and AND2 (N12806, N12802, N6754);
nand NAND2 (N12807, N12799, N4419);
buf BUF1 (N12808, N12806);
nand NAND2 (N12809, N12805, N5136);
xor XOR2 (N12810, N12809, N10093);
not NOT1 (N12811, N12803);
buf BUF1 (N12812, N12807);
xor XOR2 (N12813, N12810, N6220);
or OR4 (N12814, N12791, N1796, N4703, N7696);
not NOT1 (N12815, N12801);
buf BUF1 (N12816, N12808);
xor XOR2 (N12817, N12816, N8624);
not NOT1 (N12818, N12812);
nand NAND3 (N12819, N12817, N5228, N7856);
buf BUF1 (N12820, N12788);
xor XOR2 (N12821, N12795, N5525);
buf BUF1 (N12822, N12811);
nor NOR3 (N12823, N12800, N4184, N11191);
endmodule