// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22;

output N1017,N1021,N1010,N1001,N954,N1020,N1016,N1014,N1011,N1022;

not NOT1 (N23, N3);
nor NOR4 (N24, N18, N3, N20, N8);
or OR4 (N25, N22, N4, N1, N24);
buf BUF1 (N26, N2);
and AND3 (N27, N26, N1, N16);
xor XOR2 (N28, N19, N24);
or OR2 (N29, N2, N15);
xor XOR2 (N30, N1, N23);
buf BUF1 (N31, N5);
nand NAND4 (N32, N11, N12, N8, N17);
buf BUF1 (N33, N24);
nand NAND4 (N34, N22, N20, N25, N33);
and AND2 (N35, N16, N12);
nand NAND4 (N36, N14, N32, N7, N29);
nand NAND4 (N37, N22, N17, N6, N31);
buf BUF1 (N38, N6);
and AND4 (N39, N16, N3, N17, N22);
xor XOR2 (N40, N18, N35);
or OR4 (N41, N11, N6, N6, N38);
or OR3 (N42, N13, N13, N28);
and AND4 (N43, N35, N37, N12, N5);
and AND2 (N44, N18, N27);
or OR3 (N45, N24, N30, N27);
nor NOR3 (N46, N32, N32, N37);
nor NOR2 (N47, N45, N6);
nor NOR2 (N48, N47, N47);
nor NOR3 (N49, N41, N31, N29);
not NOT1 (N50, N49);
and AND4 (N51, N42, N27, N47, N23);
nand NAND4 (N52, N36, N31, N28, N4);
and AND3 (N53, N34, N13, N9);
nand NAND3 (N54, N51, N34, N51);
buf BUF1 (N55, N52);
nand NAND3 (N56, N39, N16, N51);
xor XOR2 (N57, N46, N15);
buf BUF1 (N58, N43);
nand NAND3 (N59, N40, N53, N22);
nor NOR2 (N60, N4, N38);
xor XOR2 (N61, N58, N20);
xor XOR2 (N62, N50, N40);
or OR4 (N63, N54, N31, N52, N61);
not NOT1 (N64, N55);
not NOT1 (N65, N17);
buf BUF1 (N66, N57);
buf BUF1 (N67, N60);
nor NOR4 (N68, N67, N7, N11, N46);
and AND2 (N69, N64, N4);
and AND4 (N70, N66, N42, N62, N13);
nor NOR3 (N71, N70, N58, N44);
not NOT1 (N72, N38);
xor XOR2 (N73, N11, N66);
not NOT1 (N74, N72);
nor NOR4 (N75, N71, N29, N24, N69);
nor NOR3 (N76, N33, N69, N13);
or OR3 (N77, N56, N56, N73);
not NOT1 (N78, N5);
nor NOR2 (N79, N76, N4);
nand NAND3 (N80, N68, N30, N43);
xor XOR2 (N81, N75, N54);
buf BUF1 (N82, N63);
not NOT1 (N83, N59);
buf BUF1 (N84, N82);
not NOT1 (N85, N65);
or OR4 (N86, N85, N42, N59, N78);
buf BUF1 (N87, N23);
nor NOR4 (N88, N74, N79, N49, N44);
buf BUF1 (N89, N70);
nor NOR2 (N90, N88, N18);
and AND4 (N91, N87, N3, N69, N63);
or OR2 (N92, N81, N73);
and AND4 (N93, N83, N64, N16, N5);
and AND2 (N94, N89, N22);
nand NAND2 (N95, N80, N56);
or OR4 (N96, N93, N72, N79, N92);
not NOT1 (N97, N48);
xor XOR2 (N98, N81, N47);
nand NAND4 (N99, N98, N77, N83, N84);
buf BUF1 (N100, N15);
not NOT1 (N101, N26);
buf BUF1 (N102, N97);
nand NAND4 (N103, N86, N70, N92, N75);
or OR2 (N104, N101, N22);
not NOT1 (N105, N90);
and AND2 (N106, N95, N46);
buf BUF1 (N107, N91);
buf BUF1 (N108, N104);
xor XOR2 (N109, N99, N55);
not NOT1 (N110, N105);
not NOT1 (N111, N100);
nand NAND2 (N112, N107, N33);
nand NAND3 (N113, N106, N14, N43);
or OR4 (N114, N102, N11, N31, N20);
buf BUF1 (N115, N112);
and AND4 (N116, N108, N6, N89, N71);
xor XOR2 (N117, N109, N54);
xor XOR2 (N118, N103, N59);
buf BUF1 (N119, N111);
or OR4 (N120, N119, N72, N34, N113);
or OR3 (N121, N17, N63, N77);
or OR4 (N122, N94, N31, N99, N5);
not NOT1 (N123, N116);
nand NAND2 (N124, N120, N64);
nor NOR2 (N125, N114, N21);
nand NAND2 (N126, N121, N125);
nand NAND2 (N127, N58, N94);
or OR4 (N128, N115, N66, N103, N47);
buf BUF1 (N129, N117);
buf BUF1 (N130, N129);
nand NAND2 (N131, N110, N84);
and AND3 (N132, N128, N71, N119);
or OR3 (N133, N126, N99, N104);
xor XOR2 (N134, N133, N18);
or OR4 (N135, N134, N105, N17, N88);
or OR3 (N136, N96, N40, N13);
xor XOR2 (N137, N118, N127);
nand NAND3 (N138, N71, N60, N125);
xor XOR2 (N139, N138, N90);
or OR3 (N140, N122, N82, N115);
nor NOR2 (N141, N132, N15);
buf BUF1 (N142, N135);
not NOT1 (N143, N131);
and AND4 (N144, N136, N51, N131, N1);
and AND2 (N145, N139, N32);
xor XOR2 (N146, N140, N114);
nand NAND3 (N147, N141, N119, N115);
nor NOR4 (N148, N124, N72, N6, N140);
or OR3 (N149, N147, N111, N24);
nand NAND4 (N150, N142, N117, N139, N8);
nor NOR2 (N151, N145, N49);
or OR4 (N152, N144, N1, N37, N78);
nor NOR4 (N153, N123, N102, N16, N26);
xor XOR2 (N154, N146, N94);
xor XOR2 (N155, N154, N55);
nand NAND3 (N156, N153, N30, N4);
xor XOR2 (N157, N152, N24);
and AND3 (N158, N130, N31, N42);
buf BUF1 (N159, N151);
not NOT1 (N160, N158);
and AND4 (N161, N150, N37, N74, N148);
or OR2 (N162, N65, N130);
buf BUF1 (N163, N137);
nor NOR3 (N164, N162, N2, N131);
not NOT1 (N165, N149);
nand NAND4 (N166, N160, N62, N70, N159);
or OR3 (N167, N21, N72, N87);
nand NAND4 (N168, N156, N69, N47, N118);
nand NAND2 (N169, N143, N72);
not NOT1 (N170, N163);
nor NOR3 (N171, N155, N46, N48);
not NOT1 (N172, N171);
not NOT1 (N173, N168);
and AND4 (N174, N157, N99, N127, N7);
nand NAND3 (N175, N165, N166, N48);
nand NAND4 (N176, N11, N116, N25, N142);
xor XOR2 (N177, N170, N46);
or OR4 (N178, N169, N85, N166, N152);
and AND2 (N179, N174, N1);
and AND3 (N180, N177, N53, N34);
and AND2 (N181, N178, N4);
xor XOR2 (N182, N167, N172);
nand NAND2 (N183, N142, N146);
nor NOR3 (N184, N161, N119, N66);
nor NOR3 (N185, N173, N107, N41);
buf BUF1 (N186, N185);
or OR3 (N187, N180, N12, N133);
or OR3 (N188, N176, N76, N159);
xor XOR2 (N189, N182, N181);
xor XOR2 (N190, N64, N35);
nor NOR3 (N191, N183, N82, N121);
nor NOR2 (N192, N186, N189);
buf BUF1 (N193, N25);
or OR3 (N194, N187, N43, N189);
or OR2 (N195, N190, N23);
buf BUF1 (N196, N164);
nand NAND4 (N197, N193, N189, N166, N53);
or OR4 (N198, N195, N21, N120, N95);
xor XOR2 (N199, N198, N193);
nor NOR4 (N200, N197, N17, N51, N41);
nor NOR4 (N201, N199, N73, N11, N38);
xor XOR2 (N202, N175, N1);
nor NOR4 (N203, N179, N109, N138, N200);
buf BUF1 (N204, N161);
or OR3 (N205, N196, N70, N176);
buf BUF1 (N206, N205);
nor NOR2 (N207, N194, N30);
nand NAND2 (N208, N188, N118);
and AND2 (N209, N208, N114);
nor NOR4 (N210, N191, N39, N138, N9);
nor NOR4 (N211, N204, N138, N110, N168);
xor XOR2 (N212, N192, N100);
nand NAND4 (N213, N184, N131, N182, N135);
not NOT1 (N214, N201);
nor NOR2 (N215, N203, N5);
and AND2 (N216, N207, N169);
nand NAND4 (N217, N206, N95, N109, N24);
xor XOR2 (N218, N212, N41);
nor NOR3 (N219, N210, N85, N80);
xor XOR2 (N220, N209, N133);
xor XOR2 (N221, N215, N72);
and AND4 (N222, N213, N28, N191, N184);
nor NOR4 (N223, N218, N39, N134, N25);
not NOT1 (N224, N202);
xor XOR2 (N225, N222, N149);
nor NOR4 (N226, N224, N153, N42, N103);
and AND2 (N227, N220, N222);
nor NOR3 (N228, N227, N127, N62);
nand NAND4 (N229, N211, N189, N171, N196);
not NOT1 (N230, N228);
or OR4 (N231, N217, N22, N163, N225);
nand NAND2 (N232, N13, N210);
buf BUF1 (N233, N216);
nor NOR4 (N234, N230, N120, N135, N81);
nor NOR4 (N235, N214, N95, N60, N60);
not NOT1 (N236, N233);
nor NOR4 (N237, N219, N23, N99, N67);
nand NAND2 (N238, N236, N225);
xor XOR2 (N239, N237, N95);
and AND4 (N240, N223, N134, N42, N171);
or OR3 (N241, N234, N137, N172);
not NOT1 (N242, N238);
not NOT1 (N243, N241);
or OR2 (N244, N232, N161);
xor XOR2 (N245, N244, N99);
not NOT1 (N246, N239);
nor NOR3 (N247, N229, N38, N217);
not NOT1 (N248, N243);
buf BUF1 (N249, N242);
nor NOR2 (N250, N248, N201);
xor XOR2 (N251, N245, N55);
and AND3 (N252, N249, N11, N41);
not NOT1 (N253, N251);
buf BUF1 (N254, N226);
and AND2 (N255, N253, N31);
nor NOR3 (N256, N221, N42, N242);
and AND2 (N257, N235, N46);
not NOT1 (N258, N250);
not NOT1 (N259, N240);
and AND3 (N260, N256, N67, N224);
and AND2 (N261, N260, N170);
or OR2 (N262, N254, N134);
nand NAND4 (N263, N255, N140, N65, N37);
or OR3 (N264, N258, N1, N23);
nor NOR3 (N265, N259, N247, N38);
xor XOR2 (N266, N183, N54);
nand NAND3 (N267, N264, N64, N155);
or OR2 (N268, N257, N34);
xor XOR2 (N269, N231, N168);
nand NAND4 (N270, N263, N30, N224, N36);
or OR2 (N271, N268, N144);
buf BUF1 (N272, N271);
or OR4 (N273, N270, N236, N184, N48);
and AND2 (N274, N262, N196);
xor XOR2 (N275, N273, N106);
nor NOR4 (N276, N252, N265, N265, N162);
or OR3 (N277, N122, N214, N32);
nor NOR3 (N278, N246, N101, N47);
xor XOR2 (N279, N277, N164);
nand NAND3 (N280, N275, N225, N242);
nor NOR3 (N281, N267, N274, N260);
nand NAND2 (N282, N236, N45);
or OR4 (N283, N280, N31, N183, N158);
xor XOR2 (N284, N269, N241);
or OR3 (N285, N261, N38, N73);
xor XOR2 (N286, N276, N204);
nor NOR3 (N287, N282, N259, N50);
nor NOR4 (N288, N287, N15, N185, N120);
and AND3 (N289, N288, N74, N13);
not NOT1 (N290, N285);
not NOT1 (N291, N279);
buf BUF1 (N292, N291);
not NOT1 (N293, N281);
buf BUF1 (N294, N266);
not NOT1 (N295, N289);
and AND3 (N296, N272, N28, N203);
nand NAND4 (N297, N295, N73, N171, N244);
and AND2 (N298, N296, N29);
not NOT1 (N299, N278);
nand NAND4 (N300, N290, N61, N99, N81);
nand NAND2 (N301, N300, N30);
and AND3 (N302, N298, N190, N99);
not NOT1 (N303, N283);
xor XOR2 (N304, N303, N146);
buf BUF1 (N305, N284);
and AND4 (N306, N297, N97, N204, N216);
buf BUF1 (N307, N302);
nor NOR3 (N308, N294, N177, N194);
nand NAND4 (N309, N307, N159, N241, N112);
nand NAND2 (N310, N292, N188);
nor NOR2 (N311, N301, N102);
or OR4 (N312, N293, N5, N215, N268);
and AND3 (N313, N304, N14, N256);
nand NAND3 (N314, N306, N84, N162);
or OR4 (N315, N310, N30, N261, N115);
nand NAND4 (N316, N299, N127, N290, N264);
buf BUF1 (N317, N312);
and AND4 (N318, N311, N148, N110, N41);
xor XOR2 (N319, N286, N219);
and AND2 (N320, N317, N55);
not NOT1 (N321, N308);
or OR2 (N322, N320, N179);
nor NOR4 (N323, N322, N211, N69, N94);
xor XOR2 (N324, N314, N249);
buf BUF1 (N325, N316);
and AND4 (N326, N323, N86, N300, N17);
xor XOR2 (N327, N326, N214);
or OR3 (N328, N309, N192, N322);
nor NOR3 (N329, N321, N11, N133);
xor XOR2 (N330, N305, N247);
or OR4 (N331, N313, N284, N150, N16);
nor NOR4 (N332, N325, N54, N159, N195);
and AND2 (N333, N319, N163);
or OR3 (N334, N333, N257, N212);
or OR3 (N335, N331, N213, N328);
not NOT1 (N336, N40);
and AND4 (N337, N318, N9, N111, N231);
xor XOR2 (N338, N324, N132);
not NOT1 (N339, N329);
not NOT1 (N340, N327);
xor XOR2 (N341, N340, N96);
and AND3 (N342, N330, N151, N107);
buf BUF1 (N343, N339);
xor XOR2 (N344, N341, N244);
nand NAND4 (N345, N343, N74, N340, N224);
buf BUF1 (N346, N334);
not NOT1 (N347, N344);
nand NAND3 (N348, N332, N14, N145);
not NOT1 (N349, N342);
nor NOR3 (N350, N338, N227, N115);
nand NAND4 (N351, N335, N60, N89, N23);
not NOT1 (N352, N345);
and AND4 (N353, N337, N166, N289, N328);
nand NAND2 (N354, N347, N250);
nand NAND2 (N355, N349, N20);
and AND4 (N356, N352, N336, N204, N211);
and AND2 (N357, N298, N341);
buf BUF1 (N358, N356);
nand NAND4 (N359, N358, N79, N35, N37);
not NOT1 (N360, N351);
nand NAND2 (N361, N354, N299);
buf BUF1 (N362, N315);
and AND2 (N363, N357, N265);
or OR2 (N364, N361, N134);
xor XOR2 (N365, N364, N160);
xor XOR2 (N366, N350, N51);
or OR2 (N367, N353, N184);
or OR4 (N368, N365, N106, N292, N163);
not NOT1 (N369, N359);
nor NOR3 (N370, N362, N32, N291);
and AND2 (N371, N370, N172);
nor NOR3 (N372, N371, N333, N88);
and AND4 (N373, N372, N365, N301, N36);
buf BUF1 (N374, N368);
not NOT1 (N375, N374);
nor NOR4 (N376, N348, N19, N274, N210);
nor NOR3 (N377, N360, N265, N152);
and AND3 (N378, N373, N286, N145);
buf BUF1 (N379, N346);
not NOT1 (N380, N378);
and AND2 (N381, N355, N99);
xor XOR2 (N382, N363, N48);
not NOT1 (N383, N377);
nor NOR2 (N384, N380, N383);
xor XOR2 (N385, N190, N52);
nor NOR4 (N386, N381, N66, N258, N224);
buf BUF1 (N387, N367);
nor NOR3 (N388, N385, N115, N212);
buf BUF1 (N389, N382);
or OR2 (N390, N386, N200);
not NOT1 (N391, N375);
not NOT1 (N392, N391);
nand NAND3 (N393, N387, N384, N61);
nor NOR3 (N394, N98, N234, N273);
and AND4 (N395, N379, N1, N353, N65);
nand NAND4 (N396, N369, N194, N99, N360);
and AND2 (N397, N376, N393);
and AND3 (N398, N346, N15, N187);
buf BUF1 (N399, N366);
xor XOR2 (N400, N392, N157);
and AND3 (N401, N398, N145, N92);
buf BUF1 (N402, N401);
nand NAND2 (N403, N389, N171);
buf BUF1 (N404, N402);
nand NAND2 (N405, N396, N221);
and AND4 (N406, N405, N35, N284, N237);
nand NAND2 (N407, N388, N149);
nand NAND4 (N408, N394, N232, N156, N407);
nand NAND4 (N409, N356, N360, N329, N235);
and AND3 (N410, N404, N251, N34);
not NOT1 (N411, N403);
or OR4 (N412, N390, N48, N360, N378);
xor XOR2 (N413, N411, N218);
xor XOR2 (N414, N408, N42);
or OR2 (N415, N400, N318);
nand NAND2 (N416, N414, N286);
nor NOR2 (N417, N415, N143);
buf BUF1 (N418, N417);
not NOT1 (N419, N410);
buf BUF1 (N420, N406);
and AND3 (N421, N397, N175, N247);
and AND4 (N422, N413, N276, N193, N125);
nand NAND3 (N423, N395, N263, N51);
and AND2 (N424, N418, N244);
not NOT1 (N425, N421);
nor NOR2 (N426, N425, N226);
xor XOR2 (N427, N423, N130);
or OR3 (N428, N416, N162, N404);
not NOT1 (N429, N427);
and AND3 (N430, N429, N380, N404);
buf BUF1 (N431, N430);
nand NAND3 (N432, N409, N34, N161);
and AND2 (N433, N422, N30);
nand NAND4 (N434, N420, N189, N116, N35);
buf BUF1 (N435, N428);
nand NAND3 (N436, N434, N332, N378);
buf BUF1 (N437, N412);
not NOT1 (N438, N399);
nand NAND2 (N439, N435, N338);
xor XOR2 (N440, N419, N419);
xor XOR2 (N441, N437, N337);
buf BUF1 (N442, N438);
and AND4 (N443, N432, N143, N360, N357);
nor NOR4 (N444, N433, N150, N308, N328);
nor NOR3 (N445, N443, N200, N414);
nor NOR3 (N446, N424, N196, N18);
or OR2 (N447, N442, N193);
and AND2 (N448, N447, N59);
not NOT1 (N449, N444);
buf BUF1 (N450, N426);
not NOT1 (N451, N431);
nor NOR4 (N452, N440, N309, N194, N264);
or OR4 (N453, N451, N353, N389, N281);
xor XOR2 (N454, N452, N343);
xor XOR2 (N455, N454, N170);
buf BUF1 (N456, N449);
or OR2 (N457, N441, N156);
and AND3 (N458, N450, N28, N179);
not NOT1 (N459, N456);
nand NAND2 (N460, N458, N446);
buf BUF1 (N461, N160);
or OR4 (N462, N448, N131, N431, N455);
and AND2 (N463, N110, N282);
not NOT1 (N464, N459);
buf BUF1 (N465, N460);
not NOT1 (N466, N436);
and AND4 (N467, N445, N46, N265, N355);
nor NOR3 (N468, N439, N420, N253);
not NOT1 (N469, N464);
nor NOR3 (N470, N469, N368, N61);
nor NOR2 (N471, N457, N347);
or OR2 (N472, N463, N374);
and AND3 (N473, N471, N177, N220);
or OR3 (N474, N461, N152, N14);
not NOT1 (N475, N472);
or OR2 (N476, N474, N455);
nor NOR3 (N477, N465, N6, N12);
and AND3 (N478, N477, N53, N413);
buf BUF1 (N479, N468);
xor XOR2 (N480, N466, N49);
or OR3 (N481, N462, N240, N73);
buf BUF1 (N482, N453);
not NOT1 (N483, N480);
and AND2 (N484, N476, N71);
buf BUF1 (N485, N475);
and AND2 (N486, N485, N277);
or OR3 (N487, N478, N195, N143);
and AND4 (N488, N473, N260, N335, N69);
nor NOR3 (N489, N484, N132, N380);
nor NOR3 (N490, N488, N62, N395);
or OR4 (N491, N483, N356, N336, N92);
or OR3 (N492, N487, N183, N385);
nor NOR3 (N493, N467, N75, N441);
and AND2 (N494, N489, N273);
or OR4 (N495, N491, N486, N383, N136);
buf BUF1 (N496, N223);
xor XOR2 (N497, N494, N457);
buf BUF1 (N498, N490);
not NOT1 (N499, N479);
xor XOR2 (N500, N498, N241);
and AND2 (N501, N481, N335);
nor NOR4 (N502, N470, N498, N166, N174);
nor NOR3 (N503, N492, N168, N459);
xor XOR2 (N504, N495, N153);
and AND2 (N505, N500, N487);
nand NAND4 (N506, N493, N114, N382, N50);
nand NAND4 (N507, N501, N124, N80, N356);
nor NOR2 (N508, N496, N466);
and AND3 (N509, N499, N282, N475);
not NOT1 (N510, N506);
or OR3 (N511, N504, N306, N318);
nand NAND4 (N512, N503, N181, N19, N10);
nand NAND2 (N513, N509, N10);
and AND2 (N514, N507, N459);
not NOT1 (N515, N510);
and AND3 (N516, N515, N391, N74);
not NOT1 (N517, N482);
buf BUF1 (N518, N502);
xor XOR2 (N519, N514, N365);
and AND2 (N520, N512, N108);
buf BUF1 (N521, N519);
nand NAND4 (N522, N517, N376, N502, N283);
or OR2 (N523, N505, N318);
or OR3 (N524, N522, N19, N78);
nand NAND2 (N525, N521, N90);
xor XOR2 (N526, N520, N429);
and AND2 (N527, N523, N363);
or OR4 (N528, N527, N329, N55, N266);
not NOT1 (N529, N511);
not NOT1 (N530, N526);
buf BUF1 (N531, N516);
xor XOR2 (N532, N513, N515);
nand NAND2 (N533, N532, N73);
not NOT1 (N534, N518);
xor XOR2 (N535, N533, N47);
and AND2 (N536, N525, N410);
or OR3 (N537, N536, N348, N165);
not NOT1 (N538, N528);
xor XOR2 (N539, N531, N478);
and AND2 (N540, N530, N521);
or OR3 (N541, N529, N523, N209);
nand NAND3 (N542, N497, N16, N326);
buf BUF1 (N543, N508);
or OR4 (N544, N541, N99, N392, N456);
nand NAND3 (N545, N538, N275, N224);
nand NAND4 (N546, N534, N289, N508, N92);
not NOT1 (N547, N543);
not NOT1 (N548, N524);
or OR3 (N549, N539, N119, N323);
nand NAND4 (N550, N545, N225, N519, N549);
xor XOR2 (N551, N154, N128);
xor XOR2 (N552, N551, N40);
buf BUF1 (N553, N540);
not NOT1 (N554, N544);
buf BUF1 (N555, N546);
and AND2 (N556, N553, N208);
xor XOR2 (N557, N547, N438);
or OR2 (N558, N548, N547);
or OR2 (N559, N542, N495);
not NOT1 (N560, N555);
not NOT1 (N561, N559);
xor XOR2 (N562, N556, N518);
not NOT1 (N563, N561);
buf BUF1 (N564, N562);
buf BUF1 (N565, N554);
not NOT1 (N566, N565);
nor NOR2 (N567, N557, N405);
nor NOR2 (N568, N563, N193);
or OR2 (N569, N567, N145);
and AND4 (N570, N550, N460, N90, N250);
or OR4 (N571, N564, N377, N298, N132);
or OR4 (N572, N566, N383, N474, N271);
nor NOR4 (N573, N558, N194, N488, N126);
nor NOR2 (N574, N552, N341);
and AND3 (N575, N574, N259, N13);
buf BUF1 (N576, N568);
nor NOR3 (N577, N535, N104, N170);
not NOT1 (N578, N560);
not NOT1 (N579, N576);
and AND4 (N580, N577, N411, N177, N286);
nor NOR3 (N581, N580, N503, N289);
nor NOR4 (N582, N578, N551, N412, N322);
buf BUF1 (N583, N571);
or OR2 (N584, N573, N123);
not NOT1 (N585, N570);
and AND4 (N586, N581, N240, N253, N384);
nor NOR3 (N587, N579, N481, N111);
not NOT1 (N588, N585);
not NOT1 (N589, N583);
and AND3 (N590, N537, N437, N476);
nor NOR4 (N591, N569, N502, N590, N436);
not NOT1 (N592, N15);
not NOT1 (N593, N582);
buf BUF1 (N594, N588);
not NOT1 (N595, N587);
xor XOR2 (N596, N572, N312);
not NOT1 (N597, N589);
not NOT1 (N598, N594);
nor NOR3 (N599, N596, N286, N198);
xor XOR2 (N600, N598, N260);
nor NOR2 (N601, N597, N141);
or OR4 (N602, N593, N316, N372, N264);
buf BUF1 (N603, N600);
and AND4 (N604, N591, N143, N548, N409);
or OR2 (N605, N601, N443);
xor XOR2 (N606, N575, N107);
nor NOR3 (N607, N602, N90, N605);
xor XOR2 (N608, N327, N403);
nor NOR4 (N609, N604, N282, N254, N335);
nand NAND2 (N610, N607, N250);
xor XOR2 (N611, N610, N425);
xor XOR2 (N612, N609, N134);
or OR3 (N613, N586, N272, N242);
xor XOR2 (N614, N603, N532);
or OR2 (N615, N611, N463);
and AND2 (N616, N615, N353);
and AND4 (N617, N592, N48, N121, N519);
and AND3 (N618, N616, N452, N147);
xor XOR2 (N619, N606, N146);
nor NOR2 (N620, N619, N570);
xor XOR2 (N621, N612, N287);
or OR2 (N622, N614, N266);
and AND4 (N623, N595, N507, N250, N494);
nor NOR4 (N624, N608, N566, N467, N130);
not NOT1 (N625, N599);
or OR2 (N626, N623, N320);
nand NAND4 (N627, N621, N247, N25, N155);
or OR3 (N628, N625, N303, N243);
nor NOR3 (N629, N628, N268, N571);
nand NAND2 (N630, N624, N472);
not NOT1 (N631, N622);
buf BUF1 (N632, N627);
nand NAND3 (N633, N620, N87, N17);
not NOT1 (N634, N613);
or OR4 (N635, N634, N39, N216, N286);
buf BUF1 (N636, N629);
buf BUF1 (N637, N584);
buf BUF1 (N638, N636);
nand NAND4 (N639, N617, N633, N425, N108);
buf BUF1 (N640, N431);
nand NAND4 (N641, N640, N296, N492, N389);
or OR4 (N642, N641, N506, N4, N23);
xor XOR2 (N643, N639, N272);
buf BUF1 (N644, N631);
not NOT1 (N645, N626);
or OR4 (N646, N638, N101, N363, N230);
nor NOR3 (N647, N635, N206, N50);
not NOT1 (N648, N646);
and AND4 (N649, N637, N541, N248, N429);
nand NAND2 (N650, N630, N210);
xor XOR2 (N651, N649, N134);
or OR3 (N652, N642, N27, N231);
nor NOR2 (N653, N618, N13);
xor XOR2 (N654, N644, N205);
not NOT1 (N655, N643);
xor XOR2 (N656, N650, N605);
or OR3 (N657, N656, N226, N542);
and AND3 (N658, N648, N234, N147);
xor XOR2 (N659, N645, N506);
or OR3 (N660, N652, N220, N557);
xor XOR2 (N661, N632, N294);
buf BUF1 (N662, N654);
and AND2 (N663, N651, N489);
nand NAND3 (N664, N661, N475, N326);
or OR2 (N665, N659, N460);
buf BUF1 (N666, N664);
and AND4 (N667, N660, N406, N571, N524);
not NOT1 (N668, N647);
nand NAND4 (N669, N655, N432, N32, N38);
or OR2 (N670, N658, N62);
buf BUF1 (N671, N665);
nor NOR4 (N672, N669, N621, N155, N589);
or OR3 (N673, N653, N76, N65);
nand NAND4 (N674, N668, N142, N200, N591);
not NOT1 (N675, N670);
xor XOR2 (N676, N671, N652);
not NOT1 (N677, N667);
nand NAND4 (N678, N672, N557, N505, N207);
nor NOR3 (N679, N677, N113, N528);
or OR3 (N680, N676, N341, N206);
not NOT1 (N681, N657);
xor XOR2 (N682, N678, N474);
nor NOR4 (N683, N680, N401, N23, N187);
or OR4 (N684, N683, N81, N458, N492);
nor NOR4 (N685, N666, N626, N504, N355);
not NOT1 (N686, N679);
and AND4 (N687, N681, N519, N123, N229);
xor XOR2 (N688, N682, N213);
and AND2 (N689, N662, N166);
not NOT1 (N690, N673);
nor NOR3 (N691, N675, N13, N686);
and AND2 (N692, N293, N194);
nand NAND4 (N693, N690, N621, N257, N460);
nor NOR3 (N694, N693, N65, N37);
nor NOR4 (N695, N692, N246, N458, N404);
nor NOR3 (N696, N689, N158, N305);
nand NAND3 (N697, N684, N139, N639);
nor NOR3 (N698, N695, N230, N136);
buf BUF1 (N699, N694);
nor NOR2 (N700, N699, N406);
not NOT1 (N701, N698);
nor NOR3 (N702, N685, N11, N444);
xor XOR2 (N703, N700, N361);
nor NOR2 (N704, N674, N545);
or OR3 (N705, N687, N375, N465);
nand NAND3 (N706, N691, N280, N109);
and AND3 (N707, N696, N286, N622);
or OR2 (N708, N707, N374);
and AND2 (N709, N708, N610);
nand NAND2 (N710, N703, N589);
nand NAND3 (N711, N705, N341, N523);
buf BUF1 (N712, N701);
xor XOR2 (N713, N697, N649);
and AND4 (N714, N713, N183, N639, N128);
and AND3 (N715, N663, N132, N677);
and AND3 (N716, N715, N283, N326);
or OR4 (N717, N711, N41, N625, N549);
not NOT1 (N718, N688);
nand NAND3 (N719, N716, N318, N361);
nand NAND2 (N720, N719, N128);
and AND2 (N721, N709, N412);
buf BUF1 (N722, N702);
nand NAND3 (N723, N704, N588, N659);
nand NAND4 (N724, N710, N267, N602, N72);
nor NOR3 (N725, N714, N103, N590);
buf BUF1 (N726, N712);
nor NOR4 (N727, N717, N268, N574, N665);
nand NAND3 (N728, N726, N555, N377);
not NOT1 (N729, N706);
not NOT1 (N730, N728);
xor XOR2 (N731, N724, N707);
buf BUF1 (N732, N723);
nand NAND2 (N733, N720, N501);
nor NOR4 (N734, N732, N173, N23, N630);
nor NOR4 (N735, N729, N397, N299, N637);
not NOT1 (N736, N731);
nor NOR4 (N737, N727, N569, N249, N679);
and AND4 (N738, N734, N320, N11, N708);
or OR4 (N739, N718, N470, N156, N421);
nand NAND2 (N740, N725, N229);
or OR4 (N741, N733, N73, N219, N217);
nand NAND4 (N742, N740, N328, N300, N110);
nand NAND3 (N743, N737, N222, N174);
and AND4 (N744, N730, N8, N525, N107);
or OR3 (N745, N742, N508, N397);
buf BUF1 (N746, N722);
xor XOR2 (N747, N736, N436);
and AND4 (N748, N743, N565, N482, N18);
or OR2 (N749, N721, N453);
not NOT1 (N750, N739);
and AND2 (N751, N747, N279);
xor XOR2 (N752, N738, N47);
not NOT1 (N753, N735);
or OR3 (N754, N744, N461, N452);
buf BUF1 (N755, N745);
not NOT1 (N756, N753);
nand NAND3 (N757, N751, N637, N207);
or OR4 (N758, N746, N132, N551, N669);
buf BUF1 (N759, N752);
or OR2 (N760, N750, N253);
and AND4 (N761, N759, N124, N513, N260);
nor NOR2 (N762, N760, N293);
not NOT1 (N763, N749);
not NOT1 (N764, N757);
or OR4 (N765, N741, N520, N133, N546);
nor NOR3 (N766, N762, N443, N57);
and AND2 (N767, N755, N247);
or OR2 (N768, N767, N572);
buf BUF1 (N769, N748);
xor XOR2 (N770, N768, N562);
or OR4 (N771, N756, N356, N241, N761);
xor XOR2 (N772, N98, N266);
not NOT1 (N773, N769);
nand NAND3 (N774, N758, N751, N756);
xor XOR2 (N775, N773, N499);
and AND3 (N776, N774, N675, N498);
nand NAND2 (N777, N763, N169);
and AND2 (N778, N766, N554);
and AND4 (N779, N754, N636, N197, N749);
buf BUF1 (N780, N772);
not NOT1 (N781, N776);
xor XOR2 (N782, N780, N692);
not NOT1 (N783, N781);
not NOT1 (N784, N775);
xor XOR2 (N785, N771, N441);
or OR4 (N786, N785, N634, N5, N633);
nand NAND4 (N787, N782, N28, N574, N786);
and AND3 (N788, N681, N486, N480);
not NOT1 (N789, N770);
or OR2 (N790, N779, N667);
not NOT1 (N791, N790);
nand NAND3 (N792, N787, N296, N45);
buf BUF1 (N793, N778);
buf BUF1 (N794, N765);
xor XOR2 (N795, N777, N170);
not NOT1 (N796, N794);
nand NAND2 (N797, N789, N290);
or OR3 (N798, N796, N691, N680);
not NOT1 (N799, N793);
not NOT1 (N800, N797);
buf BUF1 (N801, N783);
nor NOR4 (N802, N792, N8, N39, N618);
buf BUF1 (N803, N784);
buf BUF1 (N804, N791);
nor NOR4 (N805, N798, N59, N184, N426);
nand NAND4 (N806, N801, N607, N217, N731);
nand NAND2 (N807, N803, N609);
or OR2 (N808, N800, N125);
and AND3 (N809, N799, N611, N27);
xor XOR2 (N810, N808, N287);
xor XOR2 (N811, N804, N72);
buf BUF1 (N812, N811);
and AND2 (N813, N806, N405);
not NOT1 (N814, N788);
and AND2 (N815, N802, N148);
not NOT1 (N816, N814);
xor XOR2 (N817, N809, N234);
nor NOR3 (N818, N816, N706, N613);
xor XOR2 (N819, N764, N141);
or OR2 (N820, N818, N790);
and AND4 (N821, N820, N799, N84, N419);
and AND4 (N822, N795, N712, N40, N695);
or OR3 (N823, N815, N662, N555);
not NOT1 (N824, N812);
not NOT1 (N825, N824);
not NOT1 (N826, N822);
xor XOR2 (N827, N825, N358);
not NOT1 (N828, N807);
and AND2 (N829, N819, N721);
and AND4 (N830, N821, N588, N155, N636);
or OR4 (N831, N817, N335, N784, N87);
nand NAND3 (N832, N826, N391, N773);
and AND3 (N833, N829, N410, N340);
nor NOR4 (N834, N827, N481, N464, N367);
buf BUF1 (N835, N810);
xor XOR2 (N836, N828, N635);
xor XOR2 (N837, N835, N649);
xor XOR2 (N838, N834, N716);
and AND4 (N839, N813, N561, N606, N417);
xor XOR2 (N840, N839, N82);
or OR3 (N841, N823, N397, N352);
or OR3 (N842, N831, N326, N264);
and AND3 (N843, N805, N510, N264);
nand NAND4 (N844, N841, N244, N555, N107);
xor XOR2 (N845, N830, N159);
nand NAND3 (N846, N832, N124, N277);
or OR2 (N847, N836, N101);
nor NOR2 (N848, N846, N547);
and AND3 (N849, N833, N361, N827);
not NOT1 (N850, N848);
nand NAND4 (N851, N842, N261, N634, N576);
nand NAND3 (N852, N844, N222, N708);
not NOT1 (N853, N850);
nand NAND3 (N854, N845, N842, N174);
nor NOR2 (N855, N838, N636);
nand NAND2 (N856, N840, N768);
or OR3 (N857, N856, N561, N317);
or OR4 (N858, N847, N247, N684, N307);
xor XOR2 (N859, N855, N812);
nand NAND2 (N860, N843, N439);
buf BUF1 (N861, N860);
and AND3 (N862, N854, N242, N512);
or OR4 (N863, N849, N651, N461, N571);
or OR4 (N864, N852, N28, N463, N627);
xor XOR2 (N865, N864, N95);
xor XOR2 (N866, N837, N433);
or OR2 (N867, N862, N853);
not NOT1 (N868, N79);
nor NOR3 (N869, N867, N86, N570);
not NOT1 (N870, N861);
nor NOR3 (N871, N868, N552, N38);
nor NOR3 (N872, N859, N12, N543);
buf BUF1 (N873, N857);
or OR2 (N874, N869, N689);
buf BUF1 (N875, N863);
xor XOR2 (N876, N865, N43);
and AND4 (N877, N874, N798, N28, N673);
or OR3 (N878, N873, N538, N553);
not NOT1 (N879, N866);
and AND2 (N880, N879, N848);
buf BUF1 (N881, N876);
not NOT1 (N882, N881);
buf BUF1 (N883, N882);
not NOT1 (N884, N858);
nor NOR4 (N885, N871, N491, N789, N816);
or OR2 (N886, N851, N866);
xor XOR2 (N887, N878, N314);
buf BUF1 (N888, N877);
buf BUF1 (N889, N870);
or OR2 (N890, N872, N22);
and AND3 (N891, N887, N850, N525);
xor XOR2 (N892, N880, N176);
xor XOR2 (N893, N875, N183);
xor XOR2 (N894, N891, N72);
and AND4 (N895, N893, N190, N735, N795);
not NOT1 (N896, N889);
nor NOR2 (N897, N888, N428);
or OR4 (N898, N886, N555, N817, N503);
not NOT1 (N899, N895);
buf BUF1 (N900, N884);
or OR4 (N901, N883, N608, N683, N270);
nand NAND2 (N902, N885, N744);
nor NOR2 (N903, N897, N578);
nand NAND3 (N904, N892, N217, N43);
buf BUF1 (N905, N902);
buf BUF1 (N906, N901);
not NOT1 (N907, N904);
not NOT1 (N908, N905);
not NOT1 (N909, N899);
not NOT1 (N910, N907);
or OR4 (N911, N906, N99, N858, N281);
buf BUF1 (N912, N896);
xor XOR2 (N913, N898, N181);
or OR3 (N914, N900, N159, N853);
and AND3 (N915, N894, N893, N106);
not NOT1 (N916, N909);
buf BUF1 (N917, N913);
or OR2 (N918, N911, N12);
nand NAND2 (N919, N917, N813);
nand NAND4 (N920, N908, N605, N311, N735);
nand NAND4 (N921, N903, N704, N568, N516);
buf BUF1 (N922, N910);
not NOT1 (N923, N912);
buf BUF1 (N924, N919);
not NOT1 (N925, N922);
xor XOR2 (N926, N920, N17);
and AND2 (N927, N914, N290);
or OR2 (N928, N924, N723);
not NOT1 (N929, N918);
not NOT1 (N930, N927);
not NOT1 (N931, N925);
not NOT1 (N932, N890);
and AND3 (N933, N929, N217, N51);
and AND3 (N934, N928, N382, N670);
and AND3 (N935, N930, N261, N224);
and AND2 (N936, N921, N840);
not NOT1 (N937, N926);
xor XOR2 (N938, N915, N184);
or OR4 (N939, N932, N75, N870, N732);
and AND4 (N940, N923, N144, N161, N568);
nand NAND2 (N941, N939, N405);
xor XOR2 (N942, N936, N561);
and AND4 (N943, N937, N402, N905, N785);
xor XOR2 (N944, N931, N188);
or OR2 (N945, N941, N188);
xor XOR2 (N946, N938, N509);
nor NOR3 (N947, N935, N322, N322);
and AND2 (N948, N947, N263);
nor NOR2 (N949, N945, N710);
or OR2 (N950, N934, N527);
and AND4 (N951, N933, N583, N820, N120);
and AND3 (N952, N948, N809, N906);
nand NAND4 (N953, N940, N952, N524, N150);
nor NOR3 (N954, N204, N375, N782);
xor XOR2 (N955, N953, N204);
and AND2 (N956, N950, N350);
not NOT1 (N957, N916);
nand NAND2 (N958, N955, N312);
and AND2 (N959, N957, N349);
or OR3 (N960, N946, N587, N535);
buf BUF1 (N961, N943);
xor XOR2 (N962, N956, N892);
xor XOR2 (N963, N949, N527);
not NOT1 (N964, N942);
xor XOR2 (N965, N960, N304);
buf BUF1 (N966, N944);
xor XOR2 (N967, N963, N472);
nand NAND2 (N968, N966, N30);
nand NAND2 (N969, N962, N443);
not NOT1 (N970, N961);
nand NAND3 (N971, N970, N706, N228);
nor NOR3 (N972, N959, N704, N756);
nand NAND4 (N973, N951, N757, N607, N317);
and AND3 (N974, N964, N294, N14);
or OR3 (N975, N969, N888, N39);
buf BUF1 (N976, N974);
nor NOR4 (N977, N965, N576, N633, N354);
nand NAND3 (N978, N968, N396, N752);
nand NAND2 (N979, N973, N850);
nor NOR2 (N980, N971, N388);
nand NAND4 (N981, N977, N523, N95, N875);
xor XOR2 (N982, N981, N220);
nor NOR4 (N983, N978, N285, N105, N953);
and AND3 (N984, N979, N623, N878);
not NOT1 (N985, N984);
nand NAND2 (N986, N975, N886);
xor XOR2 (N987, N976, N273);
not NOT1 (N988, N967);
not NOT1 (N989, N983);
nand NAND4 (N990, N986, N923, N198, N871);
nor NOR2 (N991, N989, N365);
not NOT1 (N992, N972);
nand NAND4 (N993, N992, N330, N58, N70);
nand NAND3 (N994, N993, N663, N479);
and AND2 (N995, N990, N896);
buf BUF1 (N996, N991);
nand NAND4 (N997, N988, N502, N835, N390);
not NOT1 (N998, N958);
nand NAND3 (N999, N987, N608, N165);
and AND3 (N1000, N982, N354, N543);
nor NOR2 (N1001, N995, N898);
or OR2 (N1002, N999, N201);
buf BUF1 (N1003, N980);
not NOT1 (N1004, N1003);
xor XOR2 (N1005, N1000, N15);
not NOT1 (N1006, N1004);
buf BUF1 (N1007, N985);
not NOT1 (N1008, N994);
not NOT1 (N1009, N1006);
buf BUF1 (N1010, N996);
nand NAND3 (N1011, N998, N831, N466);
or OR4 (N1012, N1009, N252, N797, N729);
buf BUF1 (N1013, N1012);
buf BUF1 (N1014, N1007);
xor XOR2 (N1015, N1002, N102);
buf BUF1 (N1016, N997);
nand NAND2 (N1017, N1005, N1005);
and AND4 (N1018, N1008, N840, N893, N340);
and AND3 (N1019, N1015, N291, N588);
nor NOR2 (N1020, N1013, N907);
nor NOR2 (N1021, N1018, N381);
nor NOR2 (N1022, N1019, N355);
endmodule