// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23;

output N25622,N25615,N25612,N25620,N25617,N25590,N25593,N25616,N25621,N25623;

buf BUF1 (N24, N18);
or OR4 (N25, N20, N18, N20, N3);
or OR3 (N26, N12, N2, N23);
nor NOR4 (N27, N15, N4, N22, N6);
buf BUF1 (N28, N26);
xor XOR2 (N29, N3, N6);
nor NOR4 (N30, N1, N20, N5, N8);
not NOT1 (N31, N21);
and AND2 (N32, N31, N23);
or OR2 (N33, N19, N21);
or OR2 (N34, N30, N17);
or OR3 (N35, N1, N27, N8);
not NOT1 (N36, N9);
nand NAND4 (N37, N8, N7, N27, N1);
nor NOR4 (N38, N24, N9, N16, N25);
or OR4 (N39, N20, N26, N1, N37);
not NOT1 (N40, N26);
or OR3 (N41, N36, N10, N15);
not NOT1 (N42, N39);
and AND3 (N43, N34, N32, N36);
nand NAND3 (N44, N30, N18, N6);
not NOT1 (N45, N38);
not NOT1 (N46, N42);
not NOT1 (N47, N46);
and AND2 (N48, N35, N43);
and AND2 (N49, N39, N4);
not NOT1 (N50, N41);
and AND3 (N51, N50, N26, N4);
nand NAND3 (N52, N40, N25, N41);
nor NOR2 (N53, N51, N43);
not NOT1 (N54, N28);
nand NAND3 (N55, N33, N6, N41);
and AND4 (N56, N47, N33, N51, N23);
not NOT1 (N57, N48);
or OR2 (N58, N49, N23);
and AND2 (N59, N55, N45);
xor XOR2 (N60, N59, N52);
and AND4 (N61, N51, N20, N36, N36);
nand NAND4 (N62, N3, N47, N17, N16);
and AND4 (N63, N29, N60, N41, N48);
or OR4 (N64, N30, N42, N52, N28);
or OR4 (N65, N53, N11, N47, N51);
xor XOR2 (N66, N44, N41);
and AND2 (N67, N63, N11);
nand NAND3 (N68, N58, N5, N8);
buf BUF1 (N69, N54);
not NOT1 (N70, N69);
not NOT1 (N71, N61);
nand NAND4 (N72, N70, N18, N30, N15);
nor NOR3 (N73, N67, N56, N51);
buf BUF1 (N74, N64);
or OR4 (N75, N46, N62, N24, N8);
not NOT1 (N76, N14);
buf BUF1 (N77, N66);
buf BUF1 (N78, N77);
or OR4 (N79, N75, N55, N68, N46);
not NOT1 (N80, N44);
nor NOR2 (N81, N57, N2);
not NOT1 (N82, N80);
buf BUF1 (N83, N65);
nand NAND2 (N84, N73, N10);
buf BUF1 (N85, N71);
and AND2 (N86, N81, N55);
not NOT1 (N87, N79);
nor NOR3 (N88, N72, N52, N34);
or OR4 (N89, N86, N64, N80, N53);
or OR3 (N90, N88, N44, N10);
buf BUF1 (N91, N85);
or OR2 (N92, N90, N36);
not NOT1 (N93, N84);
nand NAND4 (N94, N82, N4, N28, N20);
or OR4 (N95, N93, N49, N13, N55);
buf BUF1 (N96, N94);
and AND4 (N97, N95, N36, N66, N54);
nor NOR3 (N98, N83, N40, N64);
nor NOR3 (N99, N87, N60, N35);
nor NOR3 (N100, N78, N5, N2);
nor NOR4 (N101, N99, N88, N29, N13);
and AND2 (N102, N74, N26);
and AND3 (N103, N97, N30, N97);
nand NAND2 (N104, N103, N23);
nand NAND3 (N105, N92, N97, N1);
or OR4 (N106, N96, N74, N80, N72);
nand NAND4 (N107, N105, N98, N22, N49);
not NOT1 (N108, N15);
nand NAND3 (N109, N101, N47, N51);
or OR2 (N110, N107, N104);
and AND3 (N111, N64, N1, N54);
nor NOR2 (N112, N76, N54);
buf BUF1 (N113, N112);
and AND3 (N114, N91, N34, N65);
buf BUF1 (N115, N108);
xor XOR2 (N116, N114, N74);
xor XOR2 (N117, N110, N115);
nor NOR2 (N118, N56, N74);
and AND2 (N119, N89, N98);
not NOT1 (N120, N111);
or OR3 (N121, N117, N28, N81);
xor XOR2 (N122, N120, N25);
nand NAND3 (N123, N122, N87, N121);
buf BUF1 (N124, N85);
nor NOR2 (N125, N106, N55);
xor XOR2 (N126, N113, N6);
and AND3 (N127, N124, N100, N102);
nand NAND4 (N128, N6, N74, N98, N75);
nor NOR3 (N129, N115, N45, N101);
or OR2 (N130, N127, N112);
or OR4 (N131, N119, N9, N22, N36);
and AND2 (N132, N129, N35);
nand NAND2 (N133, N132, N127);
and AND2 (N134, N118, N82);
xor XOR2 (N135, N126, N100);
not NOT1 (N136, N116);
nor NOR3 (N137, N109, N99, N129);
nor NOR3 (N138, N131, N132, N130);
not NOT1 (N139, N59);
nor NOR2 (N140, N136, N58);
nand NAND2 (N141, N128, N114);
and AND2 (N142, N134, N51);
nand NAND3 (N143, N135, N76, N2);
nor NOR3 (N144, N139, N112, N60);
not NOT1 (N145, N141);
nand NAND3 (N146, N123, N13, N109);
buf BUF1 (N147, N133);
and AND4 (N148, N144, N12, N5, N48);
and AND4 (N149, N145, N128, N101, N10);
nand NAND2 (N150, N137, N69);
or OR2 (N151, N147, N150);
not NOT1 (N152, N121);
xor XOR2 (N153, N148, N133);
nor NOR3 (N154, N149, N91, N50);
nand NAND2 (N155, N142, N7);
buf BUF1 (N156, N152);
xor XOR2 (N157, N125, N143);
nor NOR4 (N158, N110, N23, N43, N33);
nor NOR3 (N159, N154, N15, N30);
and AND2 (N160, N140, N70);
nand NAND2 (N161, N156, N25);
buf BUF1 (N162, N153);
and AND3 (N163, N146, N84, N111);
or OR4 (N164, N151, N3, N114, N64);
nand NAND4 (N165, N162, N19, N128, N120);
nand NAND4 (N166, N163, N43, N164, N58);
nor NOR4 (N167, N76, N9, N7, N85);
buf BUF1 (N168, N155);
nand NAND3 (N169, N158, N100, N140);
not NOT1 (N170, N157);
nand NAND2 (N171, N161, N88);
xor XOR2 (N172, N167, N157);
nor NOR4 (N173, N171, N70, N149, N112);
nor NOR4 (N174, N159, N3, N97, N110);
buf BUF1 (N175, N172);
nor NOR3 (N176, N165, N41, N151);
nor NOR3 (N177, N173, N152, N110);
buf BUF1 (N178, N138);
not NOT1 (N179, N166);
xor XOR2 (N180, N175, N35);
nand NAND3 (N181, N176, N145, N126);
or OR4 (N182, N177, N161, N8, N90);
nand NAND4 (N183, N170, N16, N151, N7);
not NOT1 (N184, N183);
nor NOR3 (N185, N182, N108, N139);
and AND2 (N186, N174, N129);
not NOT1 (N187, N185);
not NOT1 (N188, N181);
buf BUF1 (N189, N169);
and AND4 (N190, N189, N160, N10, N79);
xor XOR2 (N191, N21, N32);
nand NAND3 (N192, N179, N88, N38);
nand NAND4 (N193, N188, N191, N27, N96);
buf BUF1 (N194, N39);
and AND3 (N195, N192, N163, N4);
or OR2 (N196, N187, N132);
nor NOR4 (N197, N193, N117, N85, N160);
buf BUF1 (N198, N194);
nor NOR2 (N199, N178, N173);
xor XOR2 (N200, N199, N57);
or OR2 (N201, N198, N200);
and AND3 (N202, N64, N131, N118);
or OR4 (N203, N201, N15, N135, N70);
nor NOR3 (N204, N203, N199, N173);
not NOT1 (N205, N168);
not NOT1 (N206, N196);
not NOT1 (N207, N204);
nor NOR3 (N208, N190, N56, N88);
or OR4 (N209, N207, N26, N89, N153);
not NOT1 (N210, N197);
xor XOR2 (N211, N195, N141);
nand NAND4 (N212, N186, N82, N99, N28);
or OR2 (N213, N184, N80);
xor XOR2 (N214, N212, N31);
or OR3 (N215, N202, N93, N115);
nor NOR3 (N216, N208, N92, N70);
buf BUF1 (N217, N216);
nand NAND3 (N218, N209, N3, N8);
xor XOR2 (N219, N218, N98);
buf BUF1 (N220, N180);
xor XOR2 (N221, N213, N193);
nor NOR3 (N222, N219, N49, N34);
buf BUF1 (N223, N210);
xor XOR2 (N224, N217, N64);
xor XOR2 (N225, N211, N14);
nand NAND4 (N226, N223, N50, N106, N111);
or OR4 (N227, N225, N41, N196, N138);
nor NOR4 (N228, N220, N172, N161, N28);
nor NOR4 (N229, N221, N120, N133, N40);
and AND3 (N230, N222, N159, N132);
nor NOR2 (N231, N229, N225);
xor XOR2 (N232, N227, N65);
and AND3 (N233, N231, N75, N159);
buf BUF1 (N234, N205);
xor XOR2 (N235, N214, N158);
or OR4 (N236, N226, N112, N92, N121);
not NOT1 (N237, N228);
nor NOR4 (N238, N232, N133, N226, N16);
nand NAND2 (N239, N237, N219);
not NOT1 (N240, N230);
or OR2 (N241, N240, N162);
buf BUF1 (N242, N215);
and AND4 (N243, N224, N35, N60, N53);
nand NAND4 (N244, N235, N168, N38, N166);
not NOT1 (N245, N239);
buf BUF1 (N246, N234);
not NOT1 (N247, N246);
or OR3 (N248, N245, N143, N132);
nor NOR3 (N249, N242, N26, N110);
or OR4 (N250, N206, N72, N157, N190);
nand NAND2 (N251, N248, N101);
nor NOR2 (N252, N236, N31);
and AND2 (N253, N251, N114);
not NOT1 (N254, N233);
buf BUF1 (N255, N253);
xor XOR2 (N256, N249, N156);
buf BUF1 (N257, N256);
and AND2 (N258, N255, N121);
and AND2 (N259, N257, N8);
not NOT1 (N260, N238);
buf BUF1 (N261, N258);
not NOT1 (N262, N259);
nor NOR4 (N263, N244, N243, N164, N12);
nand NAND2 (N264, N96, N46);
not NOT1 (N265, N241);
xor XOR2 (N266, N252, N222);
or OR2 (N267, N266, N126);
xor XOR2 (N268, N267, N92);
nand NAND3 (N269, N254, N120, N10);
nor NOR2 (N270, N261, N203);
or OR2 (N271, N269, N244);
nand NAND4 (N272, N270, N21, N54, N200);
not NOT1 (N273, N272);
nand NAND2 (N274, N247, N75);
and AND4 (N275, N250, N161, N73, N14);
or OR2 (N276, N264, N271);
xor XOR2 (N277, N230, N4);
nor NOR2 (N278, N262, N254);
xor XOR2 (N279, N268, N122);
xor XOR2 (N280, N278, N31);
xor XOR2 (N281, N273, N265);
or OR3 (N282, N212, N220, N147);
nor NOR2 (N283, N277, N15);
nor NOR3 (N284, N274, N73, N178);
or OR4 (N285, N284, N184, N219, N114);
nor NOR3 (N286, N279, N176, N230);
not NOT1 (N287, N276);
buf BUF1 (N288, N280);
xor XOR2 (N289, N275, N83);
buf BUF1 (N290, N263);
or OR3 (N291, N282, N147, N276);
nand NAND4 (N292, N260, N31, N230, N270);
or OR3 (N293, N291, N36, N114);
nand NAND4 (N294, N287, N285, N171, N83);
buf BUF1 (N295, N288);
not NOT1 (N296, N204);
nor NOR3 (N297, N295, N90, N164);
not NOT1 (N298, N290);
xor XOR2 (N299, N297, N293);
and AND3 (N300, N154, N162, N211);
and AND2 (N301, N296, N267);
nor NOR2 (N302, N283, N31);
nand NAND3 (N303, N298, N249, N41);
not NOT1 (N304, N286);
xor XOR2 (N305, N292, N102);
nand NAND3 (N306, N304, N56, N17);
nand NAND2 (N307, N306, N85);
buf BUF1 (N308, N305);
buf BUF1 (N309, N307);
nor NOR4 (N310, N309, N204, N95, N122);
nor NOR4 (N311, N299, N241, N295, N43);
nor NOR4 (N312, N281, N127, N229, N167);
not NOT1 (N313, N301);
nor NOR3 (N314, N289, N306, N301);
nor NOR3 (N315, N311, N90, N91);
and AND2 (N316, N312, N138);
nor NOR4 (N317, N303, N243, N116, N243);
not NOT1 (N318, N315);
not NOT1 (N319, N300);
not NOT1 (N320, N302);
or OR4 (N321, N319, N109, N245, N229);
not NOT1 (N322, N294);
nand NAND3 (N323, N318, N164, N101);
buf BUF1 (N324, N320);
or OR2 (N325, N321, N97);
buf BUF1 (N326, N325);
nand NAND4 (N327, N316, N230, N117, N151);
nand NAND2 (N328, N317, N293);
nand NAND3 (N329, N322, N213, N309);
or OR2 (N330, N323, N291);
xor XOR2 (N331, N310, N138);
not NOT1 (N332, N331);
buf BUF1 (N333, N328);
xor XOR2 (N334, N327, N320);
nand NAND4 (N335, N326, N1, N295, N233);
xor XOR2 (N336, N335, N141);
nor NOR4 (N337, N313, N112, N80, N181);
nor NOR2 (N338, N314, N166);
nor NOR3 (N339, N324, N197, N67);
nand NAND2 (N340, N336, N144);
nand NAND2 (N341, N338, N44);
and AND4 (N342, N308, N183, N57, N319);
buf BUF1 (N343, N340);
xor XOR2 (N344, N332, N183);
nand NAND3 (N345, N339, N69, N261);
not NOT1 (N346, N334);
or OR4 (N347, N345, N99, N195, N174);
or OR4 (N348, N342, N252, N338, N99);
and AND4 (N349, N329, N140, N66, N215);
and AND3 (N350, N344, N88, N99);
xor XOR2 (N351, N348, N150);
or OR2 (N352, N346, N149);
not NOT1 (N353, N341);
nand NAND2 (N354, N343, N175);
nand NAND2 (N355, N330, N250);
not NOT1 (N356, N347);
nand NAND3 (N357, N333, N135, N55);
xor XOR2 (N358, N349, N291);
xor XOR2 (N359, N350, N51);
or OR2 (N360, N354, N135);
buf BUF1 (N361, N337);
xor XOR2 (N362, N356, N2);
or OR4 (N363, N352, N180, N159, N338);
nor NOR4 (N364, N351, N119, N191, N138);
nand NAND3 (N365, N357, N106, N80);
or OR3 (N366, N360, N245, N308);
not NOT1 (N367, N363);
xor XOR2 (N368, N362, N158);
xor XOR2 (N369, N367, N25);
nor NOR4 (N370, N366, N311, N38, N252);
nand NAND3 (N371, N353, N242, N209);
nand NAND2 (N372, N355, N86);
and AND2 (N373, N368, N252);
or OR4 (N374, N370, N163, N236, N160);
buf BUF1 (N375, N358);
or OR3 (N376, N373, N323, N268);
buf BUF1 (N377, N364);
buf BUF1 (N378, N371);
nor NOR2 (N379, N378, N252);
not NOT1 (N380, N359);
nand NAND2 (N381, N374, N79);
or OR4 (N382, N369, N301, N103, N342);
nor NOR3 (N383, N365, N235, N367);
not NOT1 (N384, N379);
nand NAND2 (N385, N377, N292);
not NOT1 (N386, N383);
nand NAND2 (N387, N375, N319);
nand NAND3 (N388, N386, N263, N190);
nand NAND4 (N389, N372, N64, N8, N156);
xor XOR2 (N390, N382, N209);
buf BUF1 (N391, N390);
buf BUF1 (N392, N387);
xor XOR2 (N393, N392, N257);
nor NOR2 (N394, N388, N230);
nand NAND2 (N395, N394, N283);
nand NAND4 (N396, N384, N97, N139, N123);
buf BUF1 (N397, N380);
buf BUF1 (N398, N385);
or OR4 (N399, N393, N85, N357, N251);
xor XOR2 (N400, N399, N325);
buf BUF1 (N401, N376);
or OR4 (N402, N397, N99, N136, N135);
and AND3 (N403, N402, N294, N375);
not NOT1 (N404, N391);
or OR4 (N405, N403, N294, N260, N177);
xor XOR2 (N406, N401, N192);
buf BUF1 (N407, N400);
xor XOR2 (N408, N396, N170);
xor XOR2 (N409, N404, N21);
buf BUF1 (N410, N409);
xor XOR2 (N411, N398, N365);
and AND3 (N412, N389, N312, N64);
not NOT1 (N413, N410);
nor NOR4 (N414, N381, N252, N158, N174);
or OR4 (N415, N413, N297, N190, N295);
buf BUF1 (N416, N405);
buf BUF1 (N417, N411);
xor XOR2 (N418, N412, N216);
nor NOR2 (N419, N361, N51);
xor XOR2 (N420, N416, N147);
buf BUF1 (N421, N415);
or OR4 (N422, N419, N407, N208, N52);
buf BUF1 (N423, N15);
not NOT1 (N424, N422);
and AND2 (N425, N408, N337);
and AND4 (N426, N406, N167, N33, N366);
nor NOR2 (N427, N395, N231);
xor XOR2 (N428, N420, N47);
buf BUF1 (N429, N417);
or OR3 (N430, N423, N327, N32);
buf BUF1 (N431, N414);
buf BUF1 (N432, N418);
xor XOR2 (N433, N431, N151);
and AND4 (N434, N430, N377, N250, N137);
nor NOR4 (N435, N433, N280, N228, N320);
nor NOR2 (N436, N427, N364);
buf BUF1 (N437, N436);
buf BUF1 (N438, N428);
not NOT1 (N439, N429);
not NOT1 (N440, N425);
and AND4 (N441, N426, N406, N206, N322);
or OR3 (N442, N424, N303, N224);
or OR2 (N443, N440, N157);
xor XOR2 (N444, N438, N2);
not NOT1 (N445, N435);
nor NOR4 (N446, N439, N257, N201, N394);
nor NOR3 (N447, N443, N235, N207);
nand NAND2 (N448, N444, N368);
xor XOR2 (N449, N447, N370);
buf BUF1 (N450, N421);
nand NAND2 (N451, N434, N355);
and AND3 (N452, N442, N54, N199);
xor XOR2 (N453, N449, N352);
not NOT1 (N454, N448);
and AND2 (N455, N445, N392);
and AND3 (N456, N446, N158, N390);
not NOT1 (N457, N456);
not NOT1 (N458, N450);
nor NOR3 (N459, N441, N94, N90);
buf BUF1 (N460, N457);
nor NOR3 (N461, N437, N334, N251);
not NOT1 (N462, N461);
buf BUF1 (N463, N454);
and AND2 (N464, N462, N169);
buf BUF1 (N465, N460);
buf BUF1 (N466, N455);
and AND2 (N467, N465, N98);
not NOT1 (N468, N451);
buf BUF1 (N469, N453);
or OR4 (N470, N452, N28, N158, N74);
buf BUF1 (N471, N469);
or OR2 (N472, N470, N101);
nor NOR2 (N473, N463, N369);
xor XOR2 (N474, N472, N459);
or OR4 (N475, N186, N436, N119, N372);
nor NOR4 (N476, N464, N299, N379, N230);
not NOT1 (N477, N468);
and AND3 (N478, N458, N264, N140);
nor NOR2 (N479, N473, N290);
xor XOR2 (N480, N477, N163);
or OR4 (N481, N432, N31, N77, N125);
or OR2 (N482, N467, N232);
nand NAND2 (N483, N474, N324);
nand NAND2 (N484, N482, N122);
xor XOR2 (N485, N476, N339);
nand NAND2 (N486, N483, N258);
xor XOR2 (N487, N466, N473);
or OR4 (N488, N486, N479, N270, N73);
xor XOR2 (N489, N55, N22);
xor XOR2 (N490, N475, N48);
xor XOR2 (N491, N471, N10);
xor XOR2 (N492, N487, N392);
buf BUF1 (N493, N492);
not NOT1 (N494, N488);
or OR3 (N495, N481, N102, N253);
or OR2 (N496, N490, N430);
nand NAND3 (N497, N484, N97, N233);
and AND2 (N498, N496, N189);
nor NOR3 (N499, N480, N461, N279);
xor XOR2 (N500, N497, N143);
and AND4 (N501, N491, N425, N302, N235);
or OR4 (N502, N494, N469, N378, N270);
not NOT1 (N503, N493);
nand NAND3 (N504, N499, N325, N444);
nor NOR3 (N505, N502, N462, N154);
and AND2 (N506, N505, N431);
xor XOR2 (N507, N498, N399);
or OR4 (N508, N495, N494, N496, N445);
nor NOR3 (N509, N485, N395, N44);
nor NOR4 (N510, N501, N327, N129, N140);
xor XOR2 (N511, N509, N347);
xor XOR2 (N512, N511, N74);
or OR3 (N513, N478, N169, N39);
or OR3 (N514, N506, N96, N16);
or OR3 (N515, N512, N315, N181);
nor NOR2 (N516, N510, N229);
nor NOR2 (N517, N515, N450);
not NOT1 (N518, N489);
nor NOR3 (N519, N507, N387, N455);
nor NOR4 (N520, N516, N44, N386, N330);
nand NAND2 (N521, N500, N2);
nor NOR4 (N522, N518, N477, N192, N96);
or OR4 (N523, N520, N16, N395, N414);
nand NAND3 (N524, N521, N204, N230);
nand NAND3 (N525, N519, N499, N28);
or OR4 (N526, N523, N90, N370, N12);
nand NAND3 (N527, N522, N118, N482);
nand NAND2 (N528, N517, N208);
nand NAND2 (N529, N508, N122);
and AND4 (N530, N525, N161, N380, N252);
nor NOR4 (N531, N530, N177, N417, N431);
buf BUF1 (N532, N527);
and AND3 (N533, N524, N193, N284);
nand NAND3 (N534, N526, N75, N307);
nand NAND3 (N535, N532, N237, N47);
or OR3 (N536, N533, N360, N519);
nor NOR2 (N537, N535, N32);
or OR3 (N538, N504, N295, N232);
nand NAND2 (N539, N528, N89);
or OR3 (N540, N538, N225, N22);
and AND2 (N541, N503, N278);
nand NAND2 (N542, N540, N453);
or OR4 (N543, N513, N158, N201, N4);
nand NAND2 (N544, N543, N324);
not NOT1 (N545, N536);
nor NOR3 (N546, N514, N405, N527);
and AND4 (N547, N546, N115, N60, N7);
or OR2 (N548, N537, N135);
and AND2 (N549, N542, N149);
and AND4 (N550, N529, N62, N144, N237);
or OR3 (N551, N541, N50, N144);
and AND4 (N552, N547, N265, N531, N46);
or OR2 (N553, N106, N255);
nor NOR2 (N554, N534, N143);
not NOT1 (N555, N552);
and AND2 (N556, N555, N169);
xor XOR2 (N557, N548, N21);
and AND3 (N558, N557, N523, N309);
nand NAND3 (N559, N551, N256, N335);
or OR2 (N560, N549, N72);
nand NAND3 (N561, N554, N90, N149);
xor XOR2 (N562, N559, N421);
not NOT1 (N563, N562);
nor NOR4 (N564, N544, N356, N409, N195);
nand NAND2 (N565, N560, N300);
and AND3 (N566, N553, N294, N185);
nor NOR4 (N567, N566, N365, N43, N108);
or OR4 (N568, N545, N367, N89, N246);
nor NOR2 (N569, N556, N173);
nor NOR3 (N570, N569, N87, N534);
xor XOR2 (N571, N570, N352);
or OR2 (N572, N564, N172);
not NOT1 (N573, N563);
and AND3 (N574, N572, N17, N182);
xor XOR2 (N575, N550, N24);
nand NAND2 (N576, N539, N360);
and AND4 (N577, N558, N399, N420, N185);
nor NOR2 (N578, N565, N403);
buf BUF1 (N579, N574);
nor NOR2 (N580, N575, N317);
and AND3 (N581, N573, N134, N339);
xor XOR2 (N582, N571, N138);
and AND4 (N583, N577, N484, N324, N543);
not NOT1 (N584, N580);
nand NAND4 (N585, N568, N574, N382, N219);
nor NOR4 (N586, N582, N416, N95, N195);
nor NOR4 (N587, N585, N358, N13, N60);
not NOT1 (N588, N586);
not NOT1 (N589, N576);
or OR2 (N590, N587, N457);
not NOT1 (N591, N583);
and AND2 (N592, N579, N446);
buf BUF1 (N593, N561);
nand NAND2 (N594, N581, N573);
nor NOR3 (N595, N594, N289, N258);
and AND4 (N596, N588, N203, N218, N449);
buf BUF1 (N597, N589);
not NOT1 (N598, N593);
xor XOR2 (N599, N597, N388);
nand NAND2 (N600, N596, N14);
buf BUF1 (N601, N590);
buf BUF1 (N602, N600);
xor XOR2 (N603, N602, N453);
xor XOR2 (N604, N601, N97);
nand NAND2 (N605, N591, N47);
xor XOR2 (N606, N584, N565);
xor XOR2 (N607, N578, N283);
not NOT1 (N608, N598);
not NOT1 (N609, N595);
or OR3 (N610, N607, N578, N91);
buf BUF1 (N611, N603);
xor XOR2 (N612, N606, N446);
and AND2 (N613, N567, N71);
nand NAND3 (N614, N611, N607, N293);
xor XOR2 (N615, N613, N478);
nand NAND3 (N616, N609, N187, N302);
not NOT1 (N617, N592);
or OR4 (N618, N605, N100, N48, N212);
not NOT1 (N619, N612);
nand NAND4 (N620, N614, N412, N413, N290);
xor XOR2 (N621, N617, N245);
xor XOR2 (N622, N604, N100);
not NOT1 (N623, N620);
nor NOR4 (N624, N623, N430, N314, N556);
nand NAND2 (N625, N610, N225);
buf BUF1 (N626, N624);
not NOT1 (N627, N615);
or OR2 (N628, N618, N195);
not NOT1 (N629, N626);
and AND4 (N630, N599, N220, N520, N395);
not NOT1 (N631, N629);
nor NOR3 (N632, N627, N174, N300);
or OR3 (N633, N632, N135, N223);
nand NAND3 (N634, N608, N323, N620);
and AND3 (N635, N634, N148, N147);
not NOT1 (N636, N631);
xor XOR2 (N637, N621, N95);
or OR4 (N638, N635, N75, N473, N368);
nand NAND4 (N639, N637, N335, N63, N465);
and AND4 (N640, N638, N294, N190, N550);
or OR4 (N641, N630, N472, N483, N283);
buf BUF1 (N642, N636);
nor NOR4 (N643, N622, N13, N611, N210);
nor NOR4 (N644, N633, N503, N83, N351);
nor NOR3 (N645, N628, N246, N33);
buf BUF1 (N646, N642);
not NOT1 (N647, N645);
not NOT1 (N648, N646);
not NOT1 (N649, N644);
nand NAND4 (N650, N639, N325, N297, N494);
nor NOR4 (N651, N619, N88, N271, N469);
nor NOR2 (N652, N643, N288);
or OR3 (N653, N640, N220, N473);
nor NOR3 (N654, N651, N183, N320);
buf BUF1 (N655, N653);
and AND3 (N656, N650, N558, N39);
not NOT1 (N657, N616);
xor XOR2 (N658, N648, N174);
nand NAND3 (N659, N656, N540, N296);
xor XOR2 (N660, N647, N144);
nor NOR4 (N661, N649, N374, N493, N312);
nor NOR3 (N662, N655, N632, N218);
not NOT1 (N663, N654);
xor XOR2 (N664, N663, N613);
xor XOR2 (N665, N657, N109);
or OR4 (N666, N661, N647, N250, N28);
and AND2 (N667, N641, N518);
nor NOR4 (N668, N664, N658, N171, N527);
or OR4 (N669, N9, N523, N572, N646);
or OR2 (N670, N662, N507);
nor NOR3 (N671, N666, N376, N217);
nor NOR4 (N672, N668, N512, N422, N169);
buf BUF1 (N673, N671);
or OR2 (N674, N665, N521);
xor XOR2 (N675, N673, N564);
nand NAND3 (N676, N660, N598, N39);
not NOT1 (N677, N659);
xor XOR2 (N678, N670, N560);
nand NAND4 (N679, N652, N507, N623, N415);
or OR4 (N680, N675, N267, N531, N63);
buf BUF1 (N681, N677);
buf BUF1 (N682, N672);
nor NOR2 (N683, N678, N212);
buf BUF1 (N684, N683);
xor XOR2 (N685, N681, N75);
not NOT1 (N686, N680);
not NOT1 (N687, N676);
nor NOR3 (N688, N625, N385, N543);
and AND4 (N689, N674, N268, N470, N284);
not NOT1 (N690, N688);
buf BUF1 (N691, N682);
and AND4 (N692, N684, N451, N96, N50);
not NOT1 (N693, N667);
not NOT1 (N694, N686);
buf BUF1 (N695, N692);
buf BUF1 (N696, N687);
nor NOR2 (N697, N694, N628);
nand NAND3 (N698, N697, N673, N246);
buf BUF1 (N699, N696);
not NOT1 (N700, N685);
buf BUF1 (N701, N695);
not NOT1 (N702, N679);
nor NOR2 (N703, N702, N111);
nand NAND4 (N704, N701, N239, N432, N410);
nor NOR2 (N705, N700, N1);
nor NOR4 (N706, N691, N274, N337, N68);
and AND2 (N707, N705, N22);
and AND3 (N708, N706, N656, N21);
xor XOR2 (N709, N704, N696);
nor NOR2 (N710, N708, N525);
and AND2 (N711, N707, N638);
xor XOR2 (N712, N693, N635);
buf BUF1 (N713, N711);
nor NOR3 (N714, N703, N605, N638);
nand NAND3 (N715, N710, N150, N443);
nor NOR4 (N716, N714, N306, N67, N70);
or OR3 (N717, N699, N712, N318);
or OR2 (N718, N120, N563);
or OR2 (N719, N690, N193);
nor NOR4 (N720, N669, N704, N296, N292);
not NOT1 (N721, N720);
nand NAND3 (N722, N698, N567, N463);
nand NAND2 (N723, N713, N629);
nor NOR4 (N724, N715, N384, N253, N576);
nand NAND4 (N725, N689, N548, N329, N458);
not NOT1 (N726, N719);
and AND2 (N727, N723, N183);
nor NOR3 (N728, N722, N418, N595);
xor XOR2 (N729, N728, N266);
and AND2 (N730, N717, N95);
nor NOR2 (N731, N709, N249);
or OR4 (N732, N727, N611, N501, N2);
nor NOR2 (N733, N718, N620);
nor NOR2 (N734, N731, N44);
or OR3 (N735, N733, N251, N172);
nor NOR2 (N736, N716, N319);
xor XOR2 (N737, N721, N485);
or OR4 (N738, N724, N614, N205, N705);
nor NOR3 (N739, N725, N555, N145);
or OR4 (N740, N736, N323, N716, N264);
buf BUF1 (N741, N737);
nand NAND2 (N742, N735, N37);
or OR4 (N743, N738, N472, N605, N532);
not NOT1 (N744, N726);
not NOT1 (N745, N740);
nor NOR2 (N746, N729, N81);
buf BUF1 (N747, N734);
buf BUF1 (N748, N744);
nand NAND2 (N749, N741, N586);
xor XOR2 (N750, N748, N473);
and AND4 (N751, N747, N609, N164, N204);
nand NAND3 (N752, N739, N459, N587);
xor XOR2 (N753, N730, N578);
nor NOR3 (N754, N743, N127, N563);
xor XOR2 (N755, N742, N295);
nor NOR3 (N756, N745, N299, N40);
and AND3 (N757, N746, N380, N574);
nor NOR4 (N758, N751, N101, N43, N370);
not NOT1 (N759, N749);
or OR2 (N760, N756, N500);
not NOT1 (N761, N732);
nand NAND3 (N762, N754, N92, N59);
nand NAND3 (N763, N761, N636, N82);
and AND2 (N764, N759, N9);
nor NOR2 (N765, N762, N258);
nand NAND3 (N766, N758, N461, N425);
or OR3 (N767, N760, N191, N243);
nor NOR3 (N768, N750, N14, N342);
and AND3 (N769, N766, N681, N42);
or OR2 (N770, N755, N636);
not NOT1 (N771, N752);
not NOT1 (N772, N770);
xor XOR2 (N773, N768, N377);
buf BUF1 (N774, N763);
and AND4 (N775, N757, N373, N548, N769);
nand NAND2 (N776, N589, N59);
nor NOR3 (N777, N775, N328, N241);
nand NAND2 (N778, N771, N292);
nand NAND2 (N779, N772, N328);
nand NAND3 (N780, N778, N12, N430);
not NOT1 (N781, N774);
nand NAND3 (N782, N773, N660, N294);
nand NAND2 (N783, N764, N188);
and AND3 (N784, N753, N62, N377);
nand NAND2 (N785, N765, N707);
nand NAND3 (N786, N780, N243, N460);
nor NOR2 (N787, N776, N51);
xor XOR2 (N788, N781, N715);
buf BUF1 (N789, N785);
xor XOR2 (N790, N783, N689);
and AND3 (N791, N787, N708, N113);
buf BUF1 (N792, N784);
xor XOR2 (N793, N789, N29);
nand NAND3 (N794, N793, N385, N658);
or OR2 (N795, N777, N196);
nor NOR3 (N796, N788, N730, N615);
not NOT1 (N797, N782);
and AND4 (N798, N794, N107, N724, N174);
xor XOR2 (N799, N795, N733);
xor XOR2 (N800, N796, N246);
or OR2 (N801, N791, N592);
not NOT1 (N802, N767);
buf BUF1 (N803, N792);
buf BUF1 (N804, N786);
nand NAND3 (N805, N799, N803, N457);
not NOT1 (N806, N297);
and AND4 (N807, N797, N788, N276, N365);
and AND2 (N808, N800, N14);
xor XOR2 (N809, N798, N264);
not NOT1 (N810, N779);
not NOT1 (N811, N804);
nor NOR4 (N812, N808, N303, N485, N375);
buf BUF1 (N813, N790);
xor XOR2 (N814, N813, N671);
buf BUF1 (N815, N812);
nand NAND3 (N816, N811, N99, N797);
nor NOR3 (N817, N807, N687, N110);
nand NAND4 (N818, N814, N147, N172, N399);
nand NAND4 (N819, N809, N392, N79, N302);
nor NOR3 (N820, N816, N658, N244);
buf BUF1 (N821, N818);
or OR4 (N822, N805, N675, N29, N398);
or OR2 (N823, N802, N300);
nand NAND3 (N824, N823, N100, N107);
nand NAND2 (N825, N822, N350);
nor NOR2 (N826, N810, N777);
and AND4 (N827, N806, N790, N339, N440);
and AND2 (N828, N817, N647);
and AND2 (N829, N827, N89);
buf BUF1 (N830, N819);
buf BUF1 (N831, N815);
nor NOR4 (N832, N829, N343, N138, N712);
not NOT1 (N833, N824);
or OR4 (N834, N833, N26, N278, N699);
not NOT1 (N835, N801);
not NOT1 (N836, N820);
not NOT1 (N837, N835);
not NOT1 (N838, N826);
xor XOR2 (N839, N828, N548);
or OR3 (N840, N839, N356, N300);
or OR3 (N841, N821, N312, N531);
nor NOR2 (N842, N836, N367);
nand NAND3 (N843, N837, N44, N128);
xor XOR2 (N844, N838, N761);
nand NAND3 (N845, N844, N94, N75);
xor XOR2 (N846, N843, N161);
or OR3 (N847, N845, N475, N845);
buf BUF1 (N848, N846);
buf BUF1 (N849, N841);
xor XOR2 (N850, N834, N402);
nand NAND2 (N851, N825, N252);
or OR4 (N852, N832, N38, N248, N544);
nand NAND2 (N853, N850, N723);
not NOT1 (N854, N851);
nand NAND3 (N855, N849, N157, N159);
xor XOR2 (N856, N852, N711);
or OR3 (N857, N854, N133, N578);
not NOT1 (N858, N848);
not NOT1 (N859, N858);
nor NOR4 (N860, N856, N52, N728, N796);
nand NAND3 (N861, N860, N294, N92);
buf BUF1 (N862, N840);
buf BUF1 (N863, N830);
nand NAND3 (N864, N859, N58, N604);
nor NOR3 (N865, N831, N455, N637);
and AND3 (N866, N864, N53, N666);
xor XOR2 (N867, N842, N45);
not NOT1 (N868, N866);
and AND3 (N869, N861, N227, N828);
and AND2 (N870, N847, N629);
and AND4 (N871, N867, N289, N720, N188);
and AND4 (N872, N862, N73, N817, N136);
nor NOR2 (N873, N869, N781);
nand NAND2 (N874, N868, N529);
or OR4 (N875, N863, N564, N506, N2);
nand NAND3 (N876, N872, N117, N276);
and AND3 (N877, N857, N839, N235);
and AND3 (N878, N853, N247, N492);
buf BUF1 (N879, N878);
not NOT1 (N880, N875);
nand NAND4 (N881, N874, N451, N313, N852);
buf BUF1 (N882, N879);
not NOT1 (N883, N881);
not NOT1 (N884, N880);
nor NOR3 (N885, N883, N515, N447);
nand NAND4 (N886, N865, N865, N694, N616);
and AND3 (N887, N870, N621, N730);
xor XOR2 (N888, N887, N456);
buf BUF1 (N889, N886);
or OR3 (N890, N877, N627, N838);
and AND2 (N891, N889, N782);
or OR2 (N892, N885, N405);
buf BUF1 (N893, N884);
xor XOR2 (N894, N888, N337);
buf BUF1 (N895, N882);
nand NAND4 (N896, N876, N354, N416, N223);
and AND2 (N897, N893, N786);
nor NOR3 (N898, N891, N508, N602);
xor XOR2 (N899, N895, N487);
and AND4 (N900, N896, N344, N265, N384);
nand NAND4 (N901, N892, N438, N611, N552);
not NOT1 (N902, N855);
not NOT1 (N903, N899);
nand NAND4 (N904, N900, N880, N380, N315);
nand NAND4 (N905, N901, N98, N12, N555);
or OR2 (N906, N904, N856);
xor XOR2 (N907, N894, N375);
or OR3 (N908, N890, N641, N830);
or OR2 (N909, N903, N49);
or OR4 (N910, N902, N139, N515, N860);
buf BUF1 (N911, N897);
not NOT1 (N912, N910);
buf BUF1 (N913, N907);
buf BUF1 (N914, N873);
nand NAND3 (N915, N908, N606, N146);
buf BUF1 (N916, N898);
not NOT1 (N917, N913);
buf BUF1 (N918, N912);
buf BUF1 (N919, N871);
not NOT1 (N920, N906);
nor NOR2 (N921, N918, N279);
nand NAND4 (N922, N915, N398, N401, N395);
or OR4 (N923, N909, N262, N902, N854);
nor NOR2 (N924, N911, N55);
buf BUF1 (N925, N922);
nor NOR4 (N926, N916, N512, N50, N260);
xor XOR2 (N927, N925, N334);
not NOT1 (N928, N926);
buf BUF1 (N929, N920);
and AND3 (N930, N921, N351, N852);
not NOT1 (N931, N929);
and AND3 (N932, N923, N48, N567);
nand NAND3 (N933, N917, N91, N187);
buf BUF1 (N934, N928);
nor NOR4 (N935, N914, N43, N350, N665);
nand NAND4 (N936, N905, N662, N501, N323);
buf BUF1 (N937, N931);
nor NOR4 (N938, N927, N642, N789, N675);
or OR2 (N939, N932, N770);
buf BUF1 (N940, N936);
not NOT1 (N941, N939);
or OR2 (N942, N937, N808);
nand NAND3 (N943, N941, N862, N215);
xor XOR2 (N944, N919, N274);
nor NOR4 (N945, N924, N892, N317, N626);
nand NAND4 (N946, N944, N1, N753, N437);
nand NAND3 (N947, N935, N769, N605);
nand NAND2 (N948, N940, N284);
buf BUF1 (N949, N947);
not NOT1 (N950, N943);
nand NAND4 (N951, N930, N752, N742, N825);
nor NOR4 (N952, N934, N60, N304, N461);
nor NOR2 (N953, N938, N110);
and AND4 (N954, N946, N798, N845, N257);
buf BUF1 (N955, N933);
xor XOR2 (N956, N945, N117);
and AND2 (N957, N951, N156);
and AND4 (N958, N952, N868, N887, N311);
nor NOR4 (N959, N942, N551, N611, N308);
nor NOR2 (N960, N956, N871);
buf BUF1 (N961, N958);
buf BUF1 (N962, N953);
or OR4 (N963, N961, N5, N938, N408);
and AND2 (N964, N948, N507);
or OR2 (N965, N963, N293);
not NOT1 (N966, N950);
or OR2 (N967, N955, N527);
nor NOR2 (N968, N957, N965);
not NOT1 (N969, N822);
nand NAND4 (N970, N960, N275, N858, N531);
nand NAND2 (N971, N964, N383);
not NOT1 (N972, N970);
not NOT1 (N973, N962);
buf BUF1 (N974, N959);
not NOT1 (N975, N971);
or OR3 (N976, N968, N44, N898);
or OR3 (N977, N954, N545, N550);
buf BUF1 (N978, N972);
nand NAND3 (N979, N949, N361, N719);
and AND3 (N980, N969, N769, N198);
or OR4 (N981, N979, N34, N336, N790);
and AND4 (N982, N967, N138, N965, N867);
not NOT1 (N983, N976);
and AND4 (N984, N982, N654, N8, N264);
nand NAND2 (N985, N981, N512);
xor XOR2 (N986, N977, N148);
xor XOR2 (N987, N966, N299);
xor XOR2 (N988, N980, N714);
and AND3 (N989, N985, N796, N499);
or OR2 (N990, N987, N789);
buf BUF1 (N991, N984);
nor NOR4 (N992, N978, N563, N976, N290);
nor NOR2 (N993, N989, N385);
buf BUF1 (N994, N988);
nand NAND4 (N995, N986, N595, N901, N858);
nand NAND2 (N996, N993, N73);
and AND3 (N997, N994, N230, N541);
or OR3 (N998, N992, N92, N157);
nor NOR4 (N999, N983, N206, N554, N394);
not NOT1 (N1000, N975);
buf BUF1 (N1001, N973);
nand NAND3 (N1002, N991, N866, N705);
nand NAND2 (N1003, N998, N829);
nor NOR2 (N1004, N996, N216);
and AND3 (N1005, N1003, N590, N36);
or OR2 (N1006, N990, N835);
nor NOR4 (N1007, N974, N995, N221, N580);
not NOT1 (N1008, N350);
nor NOR4 (N1009, N999, N286, N593, N318);
buf BUF1 (N1010, N1009);
buf BUF1 (N1011, N1004);
buf BUF1 (N1012, N1007);
buf BUF1 (N1013, N1001);
nor NOR3 (N1014, N1002, N801, N848);
nand NAND2 (N1015, N1008, N1009);
xor XOR2 (N1016, N1006, N466);
xor XOR2 (N1017, N1005, N669);
nor NOR4 (N1018, N1000, N737, N620, N356);
or OR2 (N1019, N1018, N870);
nand NAND3 (N1020, N1014, N628, N339);
not NOT1 (N1021, N1013);
and AND4 (N1022, N1015, N271, N345, N528);
and AND4 (N1023, N1012, N865, N209, N165);
not NOT1 (N1024, N1010);
nor NOR4 (N1025, N1020, N419, N650, N947);
and AND2 (N1026, N1017, N745);
nor NOR2 (N1027, N1024, N440);
nor NOR4 (N1028, N1011, N623, N898, N540);
buf BUF1 (N1029, N1028);
and AND3 (N1030, N1021, N155, N450);
nor NOR4 (N1031, N1016, N258, N248, N807);
nand NAND3 (N1032, N1027, N855, N462);
not NOT1 (N1033, N1019);
not NOT1 (N1034, N997);
or OR3 (N1035, N1029, N22, N413);
buf BUF1 (N1036, N1023);
not NOT1 (N1037, N1033);
nand NAND4 (N1038, N1037, N714, N584, N868);
xor XOR2 (N1039, N1031, N627);
nor NOR2 (N1040, N1026, N839);
nand NAND3 (N1041, N1034, N484, N604);
buf BUF1 (N1042, N1030);
and AND4 (N1043, N1041, N959, N1001, N1017);
nand NAND3 (N1044, N1036, N162, N327);
nor NOR2 (N1045, N1025, N439);
or OR4 (N1046, N1042, N221, N104, N250);
and AND4 (N1047, N1022, N988, N965, N409);
xor XOR2 (N1048, N1035, N662);
or OR3 (N1049, N1039, N879, N307);
xor XOR2 (N1050, N1040, N735);
nor NOR3 (N1051, N1047, N133, N805);
nand NAND3 (N1052, N1051, N963, N649);
nand NAND2 (N1053, N1049, N127);
nand NAND4 (N1054, N1043, N132, N840, N89);
not NOT1 (N1055, N1032);
and AND4 (N1056, N1045, N929, N212, N125);
xor XOR2 (N1057, N1055, N617);
nor NOR2 (N1058, N1050, N917);
nand NAND2 (N1059, N1046, N636);
nand NAND3 (N1060, N1056, N819, N854);
xor XOR2 (N1061, N1052, N946);
xor XOR2 (N1062, N1060, N862);
buf BUF1 (N1063, N1058);
nand NAND2 (N1064, N1059, N109);
xor XOR2 (N1065, N1064, N561);
buf BUF1 (N1066, N1062);
nand NAND4 (N1067, N1057, N418, N40, N899);
xor XOR2 (N1068, N1067, N773);
nand NAND4 (N1069, N1061, N607, N811, N493);
and AND4 (N1070, N1053, N398, N748, N503);
buf BUF1 (N1071, N1048);
buf BUF1 (N1072, N1070);
nor NOR3 (N1073, N1063, N905, N315);
or OR3 (N1074, N1068, N420, N75);
nor NOR3 (N1075, N1065, N302, N221);
and AND4 (N1076, N1066, N1049, N469, N472);
xor XOR2 (N1077, N1054, N377);
nand NAND3 (N1078, N1044, N91, N1002);
or OR4 (N1079, N1072, N830, N32, N901);
or OR4 (N1080, N1076, N1078, N196, N511);
xor XOR2 (N1081, N251, N1035);
nor NOR3 (N1082, N1081, N401, N199);
nor NOR4 (N1083, N1071, N88, N501, N807);
xor XOR2 (N1084, N1079, N3);
or OR3 (N1085, N1069, N567, N830);
buf BUF1 (N1086, N1082);
xor XOR2 (N1087, N1038, N760);
buf BUF1 (N1088, N1086);
nand NAND4 (N1089, N1074, N374, N936, N733);
not NOT1 (N1090, N1083);
and AND4 (N1091, N1087, N747, N309, N618);
and AND3 (N1092, N1090, N106, N245);
xor XOR2 (N1093, N1084, N508);
xor XOR2 (N1094, N1077, N729);
xor XOR2 (N1095, N1075, N734);
buf BUF1 (N1096, N1091);
xor XOR2 (N1097, N1096, N1060);
or OR2 (N1098, N1085, N501);
not NOT1 (N1099, N1094);
nor NOR3 (N1100, N1099, N587, N730);
xor XOR2 (N1101, N1089, N546);
nand NAND2 (N1102, N1095, N122);
buf BUF1 (N1103, N1100);
or OR3 (N1104, N1103, N1009, N933);
or OR3 (N1105, N1097, N465, N869);
buf BUF1 (N1106, N1088);
or OR2 (N1107, N1105, N1013);
or OR3 (N1108, N1093, N179, N598);
xor XOR2 (N1109, N1106, N504);
and AND2 (N1110, N1098, N562);
xor XOR2 (N1111, N1092, N591);
buf BUF1 (N1112, N1107);
not NOT1 (N1113, N1080);
buf BUF1 (N1114, N1110);
not NOT1 (N1115, N1109);
xor XOR2 (N1116, N1111, N746);
or OR3 (N1117, N1115, N617, N902);
buf BUF1 (N1118, N1114);
or OR3 (N1119, N1073, N286, N519);
buf BUF1 (N1120, N1119);
nor NOR2 (N1121, N1108, N187);
nand NAND4 (N1122, N1117, N436, N35, N825);
buf BUF1 (N1123, N1102);
and AND4 (N1124, N1101, N496, N979, N617);
nor NOR4 (N1125, N1124, N972, N300, N435);
xor XOR2 (N1126, N1125, N565);
not NOT1 (N1127, N1121);
and AND3 (N1128, N1104, N773, N16);
or OR4 (N1129, N1128, N606, N1017, N634);
or OR3 (N1130, N1129, N526, N848);
and AND4 (N1131, N1130, N850, N388, N123);
and AND2 (N1132, N1120, N109);
nor NOR2 (N1133, N1122, N9);
nor NOR4 (N1134, N1113, N227, N310, N452);
nor NOR4 (N1135, N1126, N258, N667, N956);
or OR4 (N1136, N1131, N863, N1022, N992);
not NOT1 (N1137, N1132);
buf BUF1 (N1138, N1123);
nor NOR2 (N1139, N1135, N1099);
nor NOR4 (N1140, N1112, N1020, N546, N1127);
xor XOR2 (N1141, N30, N287);
nor NOR2 (N1142, N1139, N521);
nor NOR4 (N1143, N1137, N557, N565, N678);
not NOT1 (N1144, N1116);
nor NOR4 (N1145, N1142, N187, N773, N356);
not NOT1 (N1146, N1143);
and AND2 (N1147, N1138, N1130);
and AND2 (N1148, N1134, N793);
xor XOR2 (N1149, N1148, N717);
or OR2 (N1150, N1144, N39);
or OR3 (N1151, N1136, N361, N716);
not NOT1 (N1152, N1150);
xor XOR2 (N1153, N1149, N411);
buf BUF1 (N1154, N1153);
xor XOR2 (N1155, N1133, N294);
or OR2 (N1156, N1145, N573);
or OR3 (N1157, N1154, N361, N708);
or OR4 (N1158, N1118, N773, N245, N985);
xor XOR2 (N1159, N1155, N322);
xor XOR2 (N1160, N1151, N759);
xor XOR2 (N1161, N1147, N6);
nor NOR2 (N1162, N1140, N72);
buf BUF1 (N1163, N1157);
xor XOR2 (N1164, N1163, N203);
buf BUF1 (N1165, N1141);
or OR2 (N1166, N1156, N872);
not NOT1 (N1167, N1166);
nor NOR3 (N1168, N1158, N464, N309);
or OR4 (N1169, N1167, N253, N1019, N3);
buf BUF1 (N1170, N1168);
xor XOR2 (N1171, N1152, N817);
or OR4 (N1172, N1164, N505, N1025, N906);
xor XOR2 (N1173, N1162, N625);
nor NOR2 (N1174, N1165, N522);
nand NAND4 (N1175, N1174, N590, N1148, N522);
or OR2 (N1176, N1159, N699);
not NOT1 (N1177, N1170);
or OR3 (N1178, N1171, N823, N257);
nor NOR3 (N1179, N1161, N189, N725);
or OR2 (N1180, N1169, N999);
or OR2 (N1181, N1172, N1064);
nand NAND3 (N1182, N1178, N115, N1059);
nand NAND3 (N1183, N1182, N718, N1172);
not NOT1 (N1184, N1173);
not NOT1 (N1185, N1183);
nand NAND2 (N1186, N1177, N479);
xor XOR2 (N1187, N1186, N137);
xor XOR2 (N1188, N1184, N203);
buf BUF1 (N1189, N1179);
xor XOR2 (N1190, N1175, N52);
and AND3 (N1191, N1146, N1008, N334);
xor XOR2 (N1192, N1180, N1045);
not NOT1 (N1193, N1160);
buf BUF1 (N1194, N1191);
or OR3 (N1195, N1193, N649, N551);
nand NAND2 (N1196, N1176, N1090);
and AND3 (N1197, N1196, N661, N591);
nand NAND4 (N1198, N1195, N448, N694, N963);
or OR2 (N1199, N1181, N83);
nor NOR2 (N1200, N1194, N1140);
not NOT1 (N1201, N1200);
buf BUF1 (N1202, N1192);
nor NOR4 (N1203, N1197, N874, N41, N972);
nor NOR3 (N1204, N1190, N338, N1051);
nor NOR2 (N1205, N1187, N582);
or OR3 (N1206, N1185, N303, N1122);
xor XOR2 (N1207, N1206, N912);
nand NAND2 (N1208, N1205, N509);
not NOT1 (N1209, N1208);
and AND2 (N1210, N1198, N118);
or OR2 (N1211, N1201, N192);
xor XOR2 (N1212, N1199, N967);
or OR4 (N1213, N1189, N80, N40, N442);
nor NOR4 (N1214, N1209, N454, N1149, N809);
nor NOR4 (N1215, N1214, N292, N567, N1208);
xor XOR2 (N1216, N1215, N140);
or OR2 (N1217, N1204, N255);
nor NOR3 (N1218, N1212, N1198, N557);
nor NOR3 (N1219, N1203, N168, N886);
and AND4 (N1220, N1213, N10, N350, N565);
not NOT1 (N1221, N1219);
nand NAND4 (N1222, N1188, N1078, N916, N447);
nand NAND3 (N1223, N1211, N1138, N280);
nand NAND2 (N1224, N1220, N1100);
nor NOR4 (N1225, N1210, N948, N253, N569);
nor NOR4 (N1226, N1207, N621, N830, N1101);
xor XOR2 (N1227, N1216, N41);
nand NAND3 (N1228, N1226, N1078, N238);
xor XOR2 (N1229, N1225, N182);
buf BUF1 (N1230, N1228);
nand NAND2 (N1231, N1224, N319);
and AND4 (N1232, N1202, N777, N289, N123);
nor NOR2 (N1233, N1231, N1033);
not NOT1 (N1234, N1232);
and AND4 (N1235, N1217, N862, N906, N1058);
not NOT1 (N1236, N1229);
nor NOR3 (N1237, N1218, N279, N1054);
buf BUF1 (N1238, N1227);
nor NOR4 (N1239, N1230, N1192, N145, N160);
nand NAND4 (N1240, N1238, N652, N166, N646);
nand NAND3 (N1241, N1222, N544, N386);
xor XOR2 (N1242, N1241, N1078);
not NOT1 (N1243, N1233);
nor NOR2 (N1244, N1239, N264);
nor NOR4 (N1245, N1221, N335, N984, N1047);
xor XOR2 (N1246, N1243, N121);
nor NOR4 (N1247, N1242, N274, N962, N37);
and AND4 (N1248, N1235, N612, N210, N318);
nand NAND2 (N1249, N1248, N1213);
nand NAND3 (N1250, N1247, N885, N1061);
nor NOR3 (N1251, N1244, N723, N303);
nand NAND4 (N1252, N1251, N32, N301, N570);
xor XOR2 (N1253, N1246, N197);
nor NOR4 (N1254, N1240, N856, N383, N1237);
not NOT1 (N1255, N201);
xor XOR2 (N1256, N1253, N708);
nand NAND4 (N1257, N1256, N635, N1107, N735);
nor NOR3 (N1258, N1245, N819, N321);
buf BUF1 (N1259, N1257);
nor NOR2 (N1260, N1236, N546);
or OR4 (N1261, N1223, N76, N329, N909);
not NOT1 (N1262, N1258);
and AND3 (N1263, N1259, N844, N754);
or OR3 (N1264, N1254, N978, N359);
buf BUF1 (N1265, N1260);
buf BUF1 (N1266, N1265);
or OR4 (N1267, N1255, N601, N558, N1218);
xor XOR2 (N1268, N1252, N849);
and AND4 (N1269, N1264, N223, N1240, N341);
not NOT1 (N1270, N1261);
and AND4 (N1271, N1270, N492, N458, N941);
and AND3 (N1272, N1263, N1149, N1262);
nor NOR3 (N1273, N1178, N762, N1266);
and AND2 (N1274, N756, N476);
and AND3 (N1275, N1234, N1068, N339);
or OR3 (N1276, N1267, N881, N105);
nor NOR3 (N1277, N1249, N572, N528);
nand NAND4 (N1278, N1250, N309, N1092, N932);
nor NOR3 (N1279, N1274, N122, N938);
buf BUF1 (N1280, N1277);
buf BUF1 (N1281, N1272);
or OR3 (N1282, N1269, N818, N96);
and AND4 (N1283, N1278, N988, N736, N641);
not NOT1 (N1284, N1279);
xor XOR2 (N1285, N1280, N808);
buf BUF1 (N1286, N1282);
nand NAND4 (N1287, N1275, N676, N1209, N824);
and AND3 (N1288, N1271, N576, N319);
or OR3 (N1289, N1286, N809, N721);
nor NOR4 (N1290, N1289, N672, N446, N505);
nand NAND2 (N1291, N1287, N1201);
buf BUF1 (N1292, N1290);
nor NOR4 (N1293, N1292, N75, N905, N368);
not NOT1 (N1294, N1283);
or OR2 (N1295, N1294, N913);
nand NAND3 (N1296, N1276, N353, N776);
buf BUF1 (N1297, N1268);
buf BUF1 (N1298, N1295);
buf BUF1 (N1299, N1293);
nand NAND3 (N1300, N1284, N1020, N1113);
nand NAND2 (N1301, N1273, N171);
nor NOR4 (N1302, N1298, N1227, N954, N984);
or OR2 (N1303, N1302, N69);
and AND3 (N1304, N1297, N27, N160);
nor NOR4 (N1305, N1304, N740, N97, N1253);
not NOT1 (N1306, N1301);
buf BUF1 (N1307, N1306);
and AND4 (N1308, N1296, N701, N590, N188);
or OR4 (N1309, N1288, N158, N753, N1120);
not NOT1 (N1310, N1300);
nand NAND4 (N1311, N1281, N1155, N213, N539);
or OR4 (N1312, N1303, N312, N457, N1282);
xor XOR2 (N1313, N1311, N18);
buf BUF1 (N1314, N1291);
nand NAND2 (N1315, N1314, N378);
not NOT1 (N1316, N1312);
not NOT1 (N1317, N1307);
nor NOR4 (N1318, N1285, N913, N1053, N164);
nand NAND4 (N1319, N1317, N1117, N952, N681);
buf BUF1 (N1320, N1316);
xor XOR2 (N1321, N1309, N692);
buf BUF1 (N1322, N1308);
not NOT1 (N1323, N1322);
nand NAND3 (N1324, N1315, N5, N1147);
or OR4 (N1325, N1299, N263, N533, N708);
and AND3 (N1326, N1320, N1009, N92);
nor NOR2 (N1327, N1319, N562);
or OR2 (N1328, N1326, N669);
not NOT1 (N1329, N1324);
nor NOR4 (N1330, N1328, N127, N1101, N1280);
nand NAND3 (N1331, N1325, N1175, N136);
and AND4 (N1332, N1330, N362, N639, N484);
nand NAND2 (N1333, N1332, N431);
xor XOR2 (N1334, N1333, N1057);
or OR4 (N1335, N1323, N576, N1210, N550);
buf BUF1 (N1336, N1321);
and AND3 (N1337, N1305, N1000, N1086);
nand NAND2 (N1338, N1335, N1124);
nor NOR4 (N1339, N1310, N858, N1312, N266);
or OR4 (N1340, N1336, N490, N1085, N412);
and AND3 (N1341, N1318, N34, N1175);
and AND2 (N1342, N1338, N933);
buf BUF1 (N1343, N1334);
buf BUF1 (N1344, N1339);
nor NOR4 (N1345, N1341, N37, N580, N987);
xor XOR2 (N1346, N1343, N35);
nand NAND3 (N1347, N1331, N1080, N262);
nor NOR3 (N1348, N1329, N723, N637);
xor XOR2 (N1349, N1327, N265);
nor NOR4 (N1350, N1349, N1224, N891, N897);
nor NOR3 (N1351, N1347, N694, N972);
nand NAND4 (N1352, N1342, N675, N996, N507);
xor XOR2 (N1353, N1340, N1291);
nand NAND3 (N1354, N1353, N953, N557);
xor XOR2 (N1355, N1351, N1161);
or OR2 (N1356, N1346, N400);
not NOT1 (N1357, N1345);
xor XOR2 (N1358, N1350, N1135);
buf BUF1 (N1359, N1357);
buf BUF1 (N1360, N1352);
xor XOR2 (N1361, N1358, N1253);
not NOT1 (N1362, N1356);
xor XOR2 (N1363, N1348, N429);
or OR4 (N1364, N1344, N947, N220, N1282);
or OR4 (N1365, N1359, N980, N491, N656);
nor NOR2 (N1366, N1364, N853);
buf BUF1 (N1367, N1365);
nor NOR3 (N1368, N1363, N483, N196);
or OR3 (N1369, N1361, N203, N252);
nand NAND3 (N1370, N1362, N1267, N619);
buf BUF1 (N1371, N1367);
or OR3 (N1372, N1313, N403, N251);
buf BUF1 (N1373, N1354);
nor NOR4 (N1374, N1337, N131, N230, N876);
nand NAND4 (N1375, N1360, N379, N190, N1058);
or OR4 (N1376, N1374, N577, N1151, N1229);
xor XOR2 (N1377, N1369, N308);
or OR2 (N1378, N1376, N792);
buf BUF1 (N1379, N1371);
not NOT1 (N1380, N1378);
and AND3 (N1381, N1373, N1357, N224);
nor NOR2 (N1382, N1372, N478);
xor XOR2 (N1383, N1370, N67);
buf BUF1 (N1384, N1382);
xor XOR2 (N1385, N1379, N478);
not NOT1 (N1386, N1385);
buf BUF1 (N1387, N1386);
xor XOR2 (N1388, N1355, N470);
nand NAND4 (N1389, N1375, N685, N539, N173);
xor XOR2 (N1390, N1389, N699);
and AND3 (N1391, N1381, N553, N1227);
nor NOR2 (N1392, N1390, N1092);
nand NAND2 (N1393, N1391, N1107);
not NOT1 (N1394, N1384);
nor NOR2 (N1395, N1388, N129);
nor NOR2 (N1396, N1368, N648);
nand NAND3 (N1397, N1380, N13, N1169);
not NOT1 (N1398, N1396);
nor NOR4 (N1399, N1394, N1386, N1106, N575);
xor XOR2 (N1400, N1377, N1332);
nand NAND4 (N1401, N1398, N268, N755, N108);
and AND3 (N1402, N1392, N109, N1386);
not NOT1 (N1403, N1402);
and AND3 (N1404, N1383, N493, N988);
or OR3 (N1405, N1403, N537, N204);
xor XOR2 (N1406, N1397, N244);
or OR3 (N1407, N1405, N887, N636);
nor NOR4 (N1408, N1366, N426, N940, N702);
not NOT1 (N1409, N1408);
xor XOR2 (N1410, N1400, N1102);
and AND4 (N1411, N1401, N289, N1325, N871);
nand NAND4 (N1412, N1393, N611, N958, N51);
or OR3 (N1413, N1399, N535, N60);
nor NOR4 (N1414, N1410, N939, N1069, N907);
and AND3 (N1415, N1406, N1283, N492);
xor XOR2 (N1416, N1413, N431);
and AND2 (N1417, N1387, N887);
not NOT1 (N1418, N1417);
nand NAND2 (N1419, N1407, N198);
nand NAND3 (N1420, N1404, N1218, N791);
xor XOR2 (N1421, N1414, N1382);
nor NOR2 (N1422, N1395, N236);
xor XOR2 (N1423, N1411, N291);
nor NOR4 (N1424, N1418, N10, N979, N910);
nor NOR2 (N1425, N1420, N537);
nor NOR3 (N1426, N1421, N1387, N561);
and AND2 (N1427, N1424, N345);
or OR4 (N1428, N1427, N3, N1273, N619);
nor NOR4 (N1429, N1422, N682, N1320, N501);
nand NAND2 (N1430, N1423, N1024);
xor XOR2 (N1431, N1416, N841);
nor NOR3 (N1432, N1412, N1072, N762);
not NOT1 (N1433, N1409);
xor XOR2 (N1434, N1426, N809);
or OR4 (N1435, N1432, N982, N214, N429);
or OR3 (N1436, N1425, N284, N607);
nand NAND2 (N1437, N1431, N881);
and AND3 (N1438, N1429, N98, N503);
or OR4 (N1439, N1437, N120, N257, N1372);
buf BUF1 (N1440, N1419);
buf BUF1 (N1441, N1439);
not NOT1 (N1442, N1430);
and AND2 (N1443, N1442, N621);
buf BUF1 (N1444, N1415);
and AND2 (N1445, N1443, N1110);
buf BUF1 (N1446, N1434);
or OR4 (N1447, N1440, N1260, N696, N872);
xor XOR2 (N1448, N1438, N321);
xor XOR2 (N1449, N1436, N656);
nor NOR4 (N1450, N1449, N1076, N1238, N1094);
xor XOR2 (N1451, N1446, N911);
buf BUF1 (N1452, N1444);
xor XOR2 (N1453, N1435, N85);
xor XOR2 (N1454, N1433, N808);
buf BUF1 (N1455, N1448);
nor NOR3 (N1456, N1453, N816, N897);
or OR3 (N1457, N1447, N6, N36);
or OR4 (N1458, N1441, N136, N776, N481);
and AND3 (N1459, N1451, N640, N838);
buf BUF1 (N1460, N1450);
and AND3 (N1461, N1445, N840, N1132);
nand NAND3 (N1462, N1428, N297, N794);
nor NOR4 (N1463, N1460, N345, N679, N739);
or OR4 (N1464, N1461, N582, N894, N74);
or OR4 (N1465, N1463, N1365, N22, N37);
nand NAND4 (N1466, N1456, N1356, N583, N549);
buf BUF1 (N1467, N1455);
xor XOR2 (N1468, N1462, N963);
nand NAND2 (N1469, N1467, N1050);
and AND3 (N1470, N1464, N925, N328);
nor NOR2 (N1471, N1459, N581);
and AND3 (N1472, N1468, N96, N1148);
buf BUF1 (N1473, N1472);
or OR3 (N1474, N1465, N90, N1054);
buf BUF1 (N1475, N1474);
buf BUF1 (N1476, N1454);
xor XOR2 (N1477, N1473, N1442);
xor XOR2 (N1478, N1469, N784);
or OR4 (N1479, N1477, N823, N758, N1272);
buf BUF1 (N1480, N1476);
or OR3 (N1481, N1452, N191, N866);
and AND2 (N1482, N1481, N906);
and AND2 (N1483, N1480, N306);
not NOT1 (N1484, N1475);
not NOT1 (N1485, N1471);
and AND2 (N1486, N1483, N1229);
nand NAND3 (N1487, N1479, N210, N892);
or OR2 (N1488, N1487, N1103);
nor NOR3 (N1489, N1482, N548, N1436);
and AND3 (N1490, N1484, N933, N1366);
buf BUF1 (N1491, N1488);
nand NAND2 (N1492, N1470, N61);
xor XOR2 (N1493, N1458, N1424);
not NOT1 (N1494, N1492);
not NOT1 (N1495, N1494);
and AND4 (N1496, N1466, N1138, N1236, N503);
xor XOR2 (N1497, N1489, N716);
nor NOR2 (N1498, N1496, N46);
xor XOR2 (N1499, N1485, N733);
or OR4 (N1500, N1499, N1027, N1003, N266);
not NOT1 (N1501, N1500);
nor NOR4 (N1502, N1478, N1082, N513, N557);
nand NAND2 (N1503, N1491, N1111);
and AND3 (N1504, N1490, N475, N161);
xor XOR2 (N1505, N1504, N810);
xor XOR2 (N1506, N1457, N819);
buf BUF1 (N1507, N1498);
buf BUF1 (N1508, N1503);
or OR4 (N1509, N1495, N1217, N1473, N1265);
and AND2 (N1510, N1486, N984);
xor XOR2 (N1511, N1502, N1249);
buf BUF1 (N1512, N1507);
nor NOR4 (N1513, N1511, N1141, N3, N21);
or OR4 (N1514, N1501, N10, N915, N1428);
or OR4 (N1515, N1497, N1050, N1301, N1128);
not NOT1 (N1516, N1505);
nor NOR3 (N1517, N1493, N686, N681);
nand NAND3 (N1518, N1514, N91, N1040);
not NOT1 (N1519, N1518);
xor XOR2 (N1520, N1513, N1119);
and AND4 (N1521, N1506, N87, N1178, N1321);
nor NOR4 (N1522, N1517, N273, N474, N1282);
buf BUF1 (N1523, N1520);
nand NAND2 (N1524, N1523, N1435);
and AND3 (N1525, N1522, N1089, N460);
nand NAND2 (N1526, N1524, N512);
buf BUF1 (N1527, N1519);
xor XOR2 (N1528, N1510, N1410);
and AND3 (N1529, N1528, N1267, N6);
nand NAND4 (N1530, N1516, N532, N63, N1269);
nor NOR2 (N1531, N1515, N22);
and AND3 (N1532, N1521, N539, N1122);
xor XOR2 (N1533, N1532, N585);
buf BUF1 (N1534, N1529);
not NOT1 (N1535, N1508);
not NOT1 (N1536, N1512);
xor XOR2 (N1537, N1531, N896);
or OR4 (N1538, N1537, N1104, N1287, N1155);
nand NAND3 (N1539, N1538, N1208, N1044);
buf BUF1 (N1540, N1530);
or OR3 (N1541, N1535, N827, N1342);
buf BUF1 (N1542, N1534);
nand NAND3 (N1543, N1539, N401, N1517);
xor XOR2 (N1544, N1536, N155);
and AND4 (N1545, N1544, N339, N1538, N1170);
buf BUF1 (N1546, N1533);
and AND2 (N1547, N1542, N625);
xor XOR2 (N1548, N1545, N1169);
or OR3 (N1549, N1541, N52, N1401);
nand NAND4 (N1550, N1509, N1179, N79, N254);
nand NAND2 (N1551, N1543, N1467);
and AND4 (N1552, N1526, N168, N784, N1264);
nor NOR2 (N1553, N1525, N752);
and AND4 (N1554, N1553, N670, N1453, N52);
or OR3 (N1555, N1527, N631, N954);
xor XOR2 (N1556, N1549, N466);
and AND4 (N1557, N1540, N627, N1005, N1177);
xor XOR2 (N1558, N1552, N27);
nor NOR3 (N1559, N1547, N238, N340);
nand NAND4 (N1560, N1548, N404, N1411, N339);
buf BUF1 (N1561, N1558);
buf BUF1 (N1562, N1557);
or OR2 (N1563, N1550, N809);
and AND4 (N1564, N1556, N1554, N291, N1020);
nor NOR2 (N1565, N731, N405);
buf BUF1 (N1566, N1559);
nand NAND4 (N1567, N1565, N1032, N184, N1095);
not NOT1 (N1568, N1546);
not NOT1 (N1569, N1568);
nor NOR4 (N1570, N1563, N1041, N407, N193);
nand NAND4 (N1571, N1570, N27, N653, N1318);
nand NAND2 (N1572, N1564, N9);
nand NAND2 (N1573, N1567, N1475);
xor XOR2 (N1574, N1571, N429);
not NOT1 (N1575, N1555);
and AND2 (N1576, N1575, N620);
and AND3 (N1577, N1569, N162, N11);
buf BUF1 (N1578, N1577);
nor NOR3 (N1579, N1574, N447, N522);
buf BUF1 (N1580, N1566);
and AND2 (N1581, N1573, N295);
nor NOR3 (N1582, N1562, N1336, N1143);
nor NOR2 (N1583, N1579, N567);
buf BUF1 (N1584, N1582);
not NOT1 (N1585, N1576);
buf BUF1 (N1586, N1561);
xor XOR2 (N1587, N1586, N1418);
not NOT1 (N1588, N1580);
not NOT1 (N1589, N1560);
or OR2 (N1590, N1587, N1249);
nor NOR2 (N1591, N1581, N487);
or OR3 (N1592, N1551, N1560, N1262);
or OR4 (N1593, N1591, N755, N270, N369);
nand NAND4 (N1594, N1588, N1217, N1127, N1320);
and AND3 (N1595, N1572, N1203, N1417);
or OR2 (N1596, N1584, N1235);
xor XOR2 (N1597, N1593, N1050);
buf BUF1 (N1598, N1583);
not NOT1 (N1599, N1595);
not NOT1 (N1600, N1598);
xor XOR2 (N1601, N1589, N1169);
nor NOR3 (N1602, N1601, N948, N1549);
buf BUF1 (N1603, N1594);
xor XOR2 (N1604, N1578, N656);
and AND4 (N1605, N1603, N1338, N338, N1060);
buf BUF1 (N1606, N1597);
buf BUF1 (N1607, N1596);
nand NAND2 (N1608, N1604, N1543);
not NOT1 (N1609, N1606);
nand NAND3 (N1610, N1602, N591, N954);
nor NOR4 (N1611, N1610, N802, N685, N858);
or OR3 (N1612, N1611, N1281, N1012);
buf BUF1 (N1613, N1592);
and AND2 (N1614, N1600, N202);
buf BUF1 (N1615, N1609);
or OR2 (N1616, N1612, N232);
and AND3 (N1617, N1613, N226, N1448);
nand NAND2 (N1618, N1615, N840);
nor NOR3 (N1619, N1585, N883, N698);
xor XOR2 (N1620, N1616, N981);
xor XOR2 (N1621, N1617, N322);
not NOT1 (N1622, N1621);
not NOT1 (N1623, N1590);
xor XOR2 (N1624, N1620, N741);
buf BUF1 (N1625, N1608);
nand NAND4 (N1626, N1605, N15, N1190, N808);
or OR2 (N1627, N1599, N52);
not NOT1 (N1628, N1626);
not NOT1 (N1629, N1614);
not NOT1 (N1630, N1628);
or OR3 (N1631, N1619, N928, N469);
nor NOR4 (N1632, N1624, N1521, N1100, N301);
and AND4 (N1633, N1618, N981, N530, N900);
nand NAND4 (N1634, N1625, N1606, N754, N1626);
xor XOR2 (N1635, N1631, N565);
and AND2 (N1636, N1632, N1383);
not NOT1 (N1637, N1635);
nor NOR3 (N1638, N1607, N478, N1141);
nor NOR2 (N1639, N1629, N976);
and AND3 (N1640, N1636, N613, N331);
buf BUF1 (N1641, N1638);
or OR4 (N1642, N1627, N1464, N607, N303);
and AND2 (N1643, N1637, N342);
and AND4 (N1644, N1634, N869, N567, N1509);
not NOT1 (N1645, N1623);
nor NOR3 (N1646, N1630, N621, N1175);
not NOT1 (N1647, N1641);
buf BUF1 (N1648, N1644);
nand NAND2 (N1649, N1639, N1446);
buf BUF1 (N1650, N1648);
nor NOR2 (N1651, N1647, N575);
or OR2 (N1652, N1650, N611);
buf BUF1 (N1653, N1645);
or OR3 (N1654, N1642, N840, N1338);
nand NAND2 (N1655, N1654, N541);
nor NOR3 (N1656, N1633, N334, N912);
not NOT1 (N1657, N1622);
xor XOR2 (N1658, N1643, N182);
not NOT1 (N1659, N1651);
xor XOR2 (N1660, N1658, N1651);
or OR4 (N1661, N1653, N1535, N250, N1083);
and AND2 (N1662, N1646, N1126);
nor NOR2 (N1663, N1662, N1468);
or OR3 (N1664, N1657, N469, N622);
and AND2 (N1665, N1663, N1128);
and AND4 (N1666, N1660, N1284, N39, N407);
xor XOR2 (N1667, N1665, N860);
and AND3 (N1668, N1656, N54, N194);
nand NAND3 (N1669, N1668, N1204, N303);
buf BUF1 (N1670, N1664);
buf BUF1 (N1671, N1659);
not NOT1 (N1672, N1667);
nor NOR4 (N1673, N1661, N1372, N700, N1354);
nand NAND2 (N1674, N1655, N672);
not NOT1 (N1675, N1674);
not NOT1 (N1676, N1652);
nand NAND3 (N1677, N1649, N770, N490);
nand NAND4 (N1678, N1673, N1119, N151, N513);
nand NAND4 (N1679, N1669, N711, N1087, N61);
not NOT1 (N1680, N1675);
xor XOR2 (N1681, N1676, N1664);
nand NAND3 (N1682, N1680, N540, N877);
nor NOR3 (N1683, N1640, N1045, N1345);
not NOT1 (N1684, N1683);
xor XOR2 (N1685, N1677, N979);
and AND4 (N1686, N1681, N955, N1580, N470);
and AND3 (N1687, N1670, N1463, N743);
xor XOR2 (N1688, N1679, N638);
nor NOR3 (N1689, N1685, N1608, N1240);
xor XOR2 (N1690, N1672, N465);
nand NAND4 (N1691, N1682, N583, N566, N1666);
buf BUF1 (N1692, N1501);
nand NAND4 (N1693, N1690, N118, N173, N913);
not NOT1 (N1694, N1671);
nor NOR3 (N1695, N1678, N950, N1285);
not NOT1 (N1696, N1687);
nor NOR2 (N1697, N1693, N325);
or OR3 (N1698, N1696, N383, N1204);
nand NAND3 (N1699, N1695, N1601, N1315);
or OR4 (N1700, N1689, N1621, N921, N88);
not NOT1 (N1701, N1688);
and AND3 (N1702, N1701, N1616, N167);
and AND4 (N1703, N1692, N747, N1598, N233);
not NOT1 (N1704, N1686);
and AND4 (N1705, N1703, N111, N951, N879);
and AND2 (N1706, N1700, N694);
buf BUF1 (N1707, N1699);
or OR3 (N1708, N1694, N258, N845);
nor NOR2 (N1709, N1697, N630);
or OR4 (N1710, N1704, N1674, N111, N494);
not NOT1 (N1711, N1708);
buf BUF1 (N1712, N1706);
xor XOR2 (N1713, N1710, N552);
nor NOR2 (N1714, N1684, N165);
not NOT1 (N1715, N1713);
nor NOR2 (N1716, N1709, N116);
nor NOR3 (N1717, N1712, N643, N1508);
nand NAND4 (N1718, N1711, N661, N1499, N1058);
buf BUF1 (N1719, N1718);
not NOT1 (N1720, N1719);
xor XOR2 (N1721, N1714, N192);
xor XOR2 (N1722, N1691, N1412);
xor XOR2 (N1723, N1705, N171);
not NOT1 (N1724, N1720);
nand NAND2 (N1725, N1722, N449);
buf BUF1 (N1726, N1724);
or OR3 (N1727, N1707, N39, N892);
buf BUF1 (N1728, N1723);
buf BUF1 (N1729, N1726);
and AND4 (N1730, N1728, N212, N383, N386);
or OR4 (N1731, N1702, N1700, N544, N1353);
not NOT1 (N1732, N1730);
and AND2 (N1733, N1721, N1592);
buf BUF1 (N1734, N1733);
and AND3 (N1735, N1725, N1133, N734);
xor XOR2 (N1736, N1727, N22);
xor XOR2 (N1737, N1736, N828);
nand NAND2 (N1738, N1729, N315);
nand NAND3 (N1739, N1738, N1578, N673);
and AND3 (N1740, N1737, N228, N1306);
buf BUF1 (N1741, N1734);
xor XOR2 (N1742, N1717, N1699);
nor NOR4 (N1743, N1731, N959, N545, N496);
not NOT1 (N1744, N1698);
nor NOR3 (N1745, N1743, N1547, N443);
nand NAND2 (N1746, N1716, N884);
and AND2 (N1747, N1735, N742);
xor XOR2 (N1748, N1739, N1635);
nor NOR2 (N1749, N1748, N796);
or OR2 (N1750, N1715, N1577);
not NOT1 (N1751, N1742);
or OR4 (N1752, N1749, N307, N1193, N175);
and AND4 (N1753, N1752, N1139, N1420, N1159);
xor XOR2 (N1754, N1741, N1506);
nand NAND2 (N1755, N1754, N855);
not NOT1 (N1756, N1750);
nand NAND4 (N1757, N1747, N1202, N170, N266);
xor XOR2 (N1758, N1755, N881);
and AND3 (N1759, N1732, N172, N1708);
and AND3 (N1760, N1759, N1693, N1378);
not NOT1 (N1761, N1740);
buf BUF1 (N1762, N1758);
xor XOR2 (N1763, N1760, N967);
not NOT1 (N1764, N1763);
xor XOR2 (N1765, N1753, N379);
or OR4 (N1766, N1745, N368, N1264, N254);
buf BUF1 (N1767, N1761);
xor XOR2 (N1768, N1744, N214);
xor XOR2 (N1769, N1751, N733);
and AND2 (N1770, N1757, N449);
nand NAND3 (N1771, N1768, N74, N1215);
and AND2 (N1772, N1769, N87);
buf BUF1 (N1773, N1772);
not NOT1 (N1774, N1767);
nand NAND3 (N1775, N1773, N115, N869);
or OR4 (N1776, N1765, N1515, N1397, N1237);
nand NAND3 (N1777, N1766, N293, N972);
xor XOR2 (N1778, N1775, N352);
and AND2 (N1779, N1764, N1114);
or OR2 (N1780, N1777, N600);
buf BUF1 (N1781, N1776);
not NOT1 (N1782, N1780);
and AND4 (N1783, N1756, N441, N1278, N1687);
and AND3 (N1784, N1782, N1478, N1321);
nand NAND2 (N1785, N1762, N958);
or OR3 (N1786, N1771, N1598, N40);
xor XOR2 (N1787, N1781, N327);
nor NOR3 (N1788, N1778, N309, N1360);
not NOT1 (N1789, N1787);
xor XOR2 (N1790, N1786, N656);
nor NOR2 (N1791, N1785, N839);
buf BUF1 (N1792, N1774);
buf BUF1 (N1793, N1788);
xor XOR2 (N1794, N1779, N526);
xor XOR2 (N1795, N1794, N888);
nand NAND3 (N1796, N1795, N663, N1669);
xor XOR2 (N1797, N1783, N989);
xor XOR2 (N1798, N1784, N576);
buf BUF1 (N1799, N1789);
nand NAND4 (N1800, N1796, N1038, N1765, N359);
or OR3 (N1801, N1791, N1662, N1712);
not NOT1 (N1802, N1801);
or OR4 (N1803, N1802, N341, N1354, N1355);
or OR4 (N1804, N1790, N1642, N1573, N617);
nand NAND3 (N1805, N1746, N1111, N624);
or OR3 (N1806, N1793, N582, N837);
or OR2 (N1807, N1798, N1503);
nor NOR4 (N1808, N1806, N1161, N1185, N1354);
not NOT1 (N1809, N1797);
not NOT1 (N1810, N1808);
not NOT1 (N1811, N1803);
nand NAND2 (N1812, N1805, N1412);
not NOT1 (N1813, N1811);
buf BUF1 (N1814, N1792);
buf BUF1 (N1815, N1810);
and AND4 (N1816, N1815, N139, N116, N309);
and AND2 (N1817, N1814, N1301);
nand NAND2 (N1818, N1770, N1689);
buf BUF1 (N1819, N1804);
or OR3 (N1820, N1818, N797, N1489);
not NOT1 (N1821, N1819);
nor NOR3 (N1822, N1799, N1431, N626);
nand NAND3 (N1823, N1816, N1133, N134);
not NOT1 (N1824, N1822);
not NOT1 (N1825, N1812);
nor NOR4 (N1826, N1825, N1552, N1040, N1683);
and AND3 (N1827, N1809, N1256, N1119);
or OR2 (N1828, N1820, N147);
nor NOR2 (N1829, N1817, N836);
xor XOR2 (N1830, N1813, N921);
buf BUF1 (N1831, N1807);
nor NOR2 (N1832, N1828, N1620);
nor NOR4 (N1833, N1830, N557, N1423, N621);
and AND2 (N1834, N1831, N66);
nand NAND2 (N1835, N1826, N700);
and AND3 (N1836, N1835, N714, N1141);
not NOT1 (N1837, N1800);
buf BUF1 (N1838, N1832);
and AND3 (N1839, N1838, N1610, N364);
nor NOR2 (N1840, N1839, N917);
or OR2 (N1841, N1829, N557);
nor NOR4 (N1842, N1827, N1198, N154, N787);
not NOT1 (N1843, N1836);
xor XOR2 (N1844, N1824, N303);
buf BUF1 (N1845, N1821);
nand NAND2 (N1846, N1844, N1126);
nand NAND4 (N1847, N1837, N1058, N50, N1564);
xor XOR2 (N1848, N1845, N500);
buf BUF1 (N1849, N1843);
and AND4 (N1850, N1841, N892, N1282, N1204);
and AND3 (N1851, N1849, N712, N41);
or OR4 (N1852, N1848, N1803, N1767, N1543);
not NOT1 (N1853, N1833);
and AND2 (N1854, N1852, N887);
buf BUF1 (N1855, N1854);
buf BUF1 (N1856, N1842);
nand NAND3 (N1857, N1846, N1242, N765);
nand NAND4 (N1858, N1856, N1705, N3, N1461);
and AND4 (N1859, N1834, N309, N338, N1103);
xor XOR2 (N1860, N1823, N1842);
and AND4 (N1861, N1859, N1831, N68, N1354);
nand NAND2 (N1862, N1853, N795);
nand NAND3 (N1863, N1847, N1011, N283);
or OR4 (N1864, N1862, N1751, N1742, N1107);
or OR2 (N1865, N1851, N1385);
not NOT1 (N1866, N1858);
nand NAND4 (N1867, N1863, N452, N1248, N1073);
nand NAND4 (N1868, N1867, N471, N1002, N1058);
buf BUF1 (N1869, N1840);
xor XOR2 (N1870, N1866, N595);
or OR3 (N1871, N1870, N947, N155);
buf BUF1 (N1872, N1861);
or OR4 (N1873, N1850, N860, N409, N1626);
or OR4 (N1874, N1869, N1475, N604, N1429);
xor XOR2 (N1875, N1864, N854);
and AND4 (N1876, N1875, N745, N1835, N433);
not NOT1 (N1877, N1876);
nor NOR3 (N1878, N1868, N212, N1255);
xor XOR2 (N1879, N1873, N916);
nor NOR4 (N1880, N1877, N16, N852, N514);
buf BUF1 (N1881, N1857);
or OR4 (N1882, N1860, N265, N835, N573);
nand NAND3 (N1883, N1871, N960, N193);
not NOT1 (N1884, N1879);
buf BUF1 (N1885, N1865);
and AND4 (N1886, N1883, N404, N1243, N914);
or OR2 (N1887, N1878, N766);
nand NAND2 (N1888, N1886, N1440);
not NOT1 (N1889, N1872);
xor XOR2 (N1890, N1881, N590);
or OR4 (N1891, N1890, N895, N1202, N83);
not NOT1 (N1892, N1874);
and AND2 (N1893, N1892, N420);
nand NAND3 (N1894, N1880, N1250, N784);
and AND4 (N1895, N1888, N668, N1882, N1209);
xor XOR2 (N1896, N650, N911);
not NOT1 (N1897, N1887);
xor XOR2 (N1898, N1893, N1017);
not NOT1 (N1899, N1894);
xor XOR2 (N1900, N1897, N1169);
buf BUF1 (N1901, N1895);
or OR2 (N1902, N1891, N1551);
buf BUF1 (N1903, N1884);
not NOT1 (N1904, N1896);
buf BUF1 (N1905, N1904);
and AND2 (N1906, N1900, N330);
or OR2 (N1907, N1905, N163);
and AND3 (N1908, N1903, N1671, N465);
buf BUF1 (N1909, N1906);
nor NOR2 (N1910, N1889, N927);
nor NOR3 (N1911, N1898, N823, N1356);
nand NAND2 (N1912, N1855, N588);
and AND2 (N1913, N1910, N240);
xor XOR2 (N1914, N1907, N697);
xor XOR2 (N1915, N1911, N1426);
xor XOR2 (N1916, N1885, N1777);
not NOT1 (N1917, N1916);
or OR4 (N1918, N1899, N1742, N625, N683);
buf BUF1 (N1919, N1918);
and AND4 (N1920, N1919, N558, N935, N823);
or OR4 (N1921, N1909, N606, N780, N1741);
xor XOR2 (N1922, N1917, N680);
xor XOR2 (N1923, N1920, N241);
xor XOR2 (N1924, N1913, N1638);
buf BUF1 (N1925, N1922);
or OR4 (N1926, N1908, N1205, N1267, N1627);
not NOT1 (N1927, N1914);
nor NOR3 (N1928, N1912, N1059, N1721);
nand NAND3 (N1929, N1901, N57, N104);
or OR2 (N1930, N1924, N1334);
not NOT1 (N1931, N1928);
not NOT1 (N1932, N1923);
not NOT1 (N1933, N1902);
nand NAND2 (N1934, N1925, N1888);
nor NOR4 (N1935, N1929, N1176, N1537, N931);
buf BUF1 (N1936, N1933);
nor NOR3 (N1937, N1926, N1528, N580);
nand NAND2 (N1938, N1935, N1819);
nor NOR3 (N1939, N1921, N344, N1640);
not NOT1 (N1940, N1938);
buf BUF1 (N1941, N1930);
and AND2 (N1942, N1915, N534);
or OR2 (N1943, N1927, N795);
and AND3 (N1944, N1939, N1560, N1236);
and AND4 (N1945, N1932, N742, N1492, N646);
or OR3 (N1946, N1931, N390, N712);
and AND3 (N1947, N1940, N103, N1622);
nand NAND3 (N1948, N1946, N941, N166);
nor NOR2 (N1949, N1943, N220);
buf BUF1 (N1950, N1945);
nand NAND4 (N1951, N1941, N701, N1620, N1418);
not NOT1 (N1952, N1936);
and AND4 (N1953, N1950, N1469, N402, N1437);
xor XOR2 (N1954, N1934, N1783);
and AND2 (N1955, N1937, N1759);
and AND2 (N1956, N1944, N1149);
xor XOR2 (N1957, N1953, N1586);
not NOT1 (N1958, N1949);
nor NOR2 (N1959, N1955, N1526);
and AND2 (N1960, N1947, N1278);
xor XOR2 (N1961, N1952, N1540);
buf BUF1 (N1962, N1961);
nor NOR3 (N1963, N1957, N1006, N674);
not NOT1 (N1964, N1960);
not NOT1 (N1965, N1956);
xor XOR2 (N1966, N1963, N237);
buf BUF1 (N1967, N1958);
nor NOR2 (N1968, N1948, N572);
nand NAND2 (N1969, N1942, N1753);
or OR3 (N1970, N1967, N417, N1642);
nor NOR3 (N1971, N1951, N780, N580);
buf BUF1 (N1972, N1962);
buf BUF1 (N1973, N1959);
xor XOR2 (N1974, N1965, N1483);
xor XOR2 (N1975, N1973, N1264);
nand NAND2 (N1976, N1972, N1795);
or OR3 (N1977, N1969, N889, N32);
or OR3 (N1978, N1968, N26, N1427);
nand NAND4 (N1979, N1971, N1850, N1437, N1802);
and AND4 (N1980, N1976, N1348, N1531, N1920);
and AND2 (N1981, N1964, N959);
nand NAND4 (N1982, N1980, N599, N1734, N225);
nand NAND3 (N1983, N1979, N337, N1100);
or OR4 (N1984, N1983, N125, N549, N101);
buf BUF1 (N1985, N1981);
xor XOR2 (N1986, N1966, N1846);
nor NOR3 (N1987, N1954, N277, N849);
buf BUF1 (N1988, N1978);
nor NOR3 (N1989, N1984, N751, N157);
nor NOR4 (N1990, N1985, N1189, N1484, N479);
xor XOR2 (N1991, N1977, N1457);
or OR2 (N1992, N1982, N817);
and AND3 (N1993, N1991, N93, N85);
buf BUF1 (N1994, N1970);
or OR2 (N1995, N1986, N969);
or OR3 (N1996, N1988, N713, N1126);
nand NAND2 (N1997, N1993, N1967);
buf BUF1 (N1998, N1996);
xor XOR2 (N1999, N1974, N842);
not NOT1 (N2000, N1995);
or OR2 (N2001, N1998, N1597);
and AND2 (N2002, N2001, N1970);
not NOT1 (N2003, N1994);
buf BUF1 (N2004, N1989);
or OR3 (N2005, N1990, N388, N259);
nor NOR2 (N2006, N1997, N1815);
buf BUF1 (N2007, N1975);
not NOT1 (N2008, N2005);
not NOT1 (N2009, N2002);
or OR3 (N2010, N2007, N785, N923);
not NOT1 (N2011, N2000);
xor XOR2 (N2012, N2003, N1818);
or OR2 (N2013, N2004, N1442);
nand NAND4 (N2014, N2013, N830, N220, N450);
not NOT1 (N2015, N2008);
buf BUF1 (N2016, N2006);
nand NAND3 (N2017, N2016, N73, N1700);
buf BUF1 (N2018, N2011);
nand NAND4 (N2019, N2014, N1317, N300, N168);
buf BUF1 (N2020, N2018);
or OR2 (N2021, N1999, N254);
nand NAND3 (N2022, N2009, N1407, N933);
or OR3 (N2023, N2019, N991, N1183);
buf BUF1 (N2024, N2022);
buf BUF1 (N2025, N2017);
and AND3 (N2026, N2021, N907, N1247);
buf BUF1 (N2027, N2025);
nand NAND3 (N2028, N2020, N1467, N507);
nand NAND2 (N2029, N2010, N1119);
or OR2 (N2030, N2026, N651);
and AND3 (N2031, N2027, N752, N851);
nor NOR2 (N2032, N2029, N1192);
and AND4 (N2033, N1992, N1702, N238, N1958);
not NOT1 (N2034, N2015);
nand NAND2 (N2035, N2030, N1181);
or OR4 (N2036, N2032, N373, N677, N599);
xor XOR2 (N2037, N2024, N771);
or OR2 (N2038, N2036, N299);
not NOT1 (N2039, N2012);
or OR4 (N2040, N2034, N685, N1141, N1840);
or OR2 (N2041, N2039, N1564);
nor NOR3 (N2042, N2035, N1890, N1586);
nor NOR2 (N2043, N2038, N1819);
nor NOR3 (N2044, N2043, N1158, N1513);
nor NOR2 (N2045, N2040, N1003);
buf BUF1 (N2046, N2041);
buf BUF1 (N2047, N1987);
xor XOR2 (N2048, N2046, N573);
not NOT1 (N2049, N2044);
xor XOR2 (N2050, N2037, N1067);
buf BUF1 (N2051, N2023);
nand NAND4 (N2052, N2045, N800, N362, N1691);
xor XOR2 (N2053, N2052, N466);
and AND4 (N2054, N2048, N1342, N1957, N28);
nand NAND2 (N2055, N2031, N97);
or OR2 (N2056, N2051, N760);
not NOT1 (N2057, N2042);
or OR4 (N2058, N2050, N990, N272, N1156);
and AND3 (N2059, N2055, N67, N882);
and AND3 (N2060, N2054, N1360, N1565);
or OR3 (N2061, N2060, N1512, N120);
nand NAND4 (N2062, N2033, N593, N1271, N1629);
xor XOR2 (N2063, N2061, N1022);
xor XOR2 (N2064, N2047, N602);
and AND3 (N2065, N2057, N483, N712);
or OR4 (N2066, N2056, N780, N2021, N1672);
xor XOR2 (N2067, N2049, N625);
xor XOR2 (N2068, N2028, N2027);
and AND4 (N2069, N2063, N514, N1864, N554);
and AND2 (N2070, N2062, N601);
xor XOR2 (N2071, N2068, N1885);
buf BUF1 (N2072, N2070);
or OR2 (N2073, N2059, N1417);
not NOT1 (N2074, N2058);
buf BUF1 (N2075, N2072);
or OR2 (N2076, N2067, N631);
or OR3 (N2077, N2069, N963, N253);
nor NOR4 (N2078, N2064, N1772, N1368, N325);
xor XOR2 (N2079, N2077, N70);
or OR3 (N2080, N2079, N1558, N52);
buf BUF1 (N2081, N2078);
buf BUF1 (N2082, N2074);
nor NOR4 (N2083, N2065, N802, N1885, N1141);
or OR2 (N2084, N2083, N130);
nand NAND3 (N2085, N2073, N1420, N1118);
not NOT1 (N2086, N2076);
xor XOR2 (N2087, N2053, N17);
nor NOR4 (N2088, N2081, N364, N880, N260);
nor NOR2 (N2089, N2080, N167);
buf BUF1 (N2090, N2084);
nand NAND2 (N2091, N2066, N1789);
xor XOR2 (N2092, N2085, N898);
or OR2 (N2093, N2086, N1587);
nor NOR4 (N2094, N2075, N852, N1751, N657);
nor NOR2 (N2095, N2088, N614);
xor XOR2 (N2096, N2091, N1910);
and AND2 (N2097, N2090, N1318);
buf BUF1 (N2098, N2093);
and AND3 (N2099, N2097, N1809, N610);
buf BUF1 (N2100, N2096);
buf BUF1 (N2101, N2100);
nand NAND4 (N2102, N2092, N1252, N139, N545);
xor XOR2 (N2103, N2089, N930);
not NOT1 (N2104, N2099);
not NOT1 (N2105, N2102);
nor NOR4 (N2106, N2105, N2087, N572, N1771);
nor NOR2 (N2107, N1945, N737);
and AND2 (N2108, N2082, N1933);
not NOT1 (N2109, N2098);
or OR4 (N2110, N2107, N1002, N251, N1152);
buf BUF1 (N2111, N2103);
not NOT1 (N2112, N2110);
nand NAND2 (N2113, N2071, N1587);
buf BUF1 (N2114, N2104);
nor NOR3 (N2115, N2114, N1392, N2057);
nor NOR3 (N2116, N2095, N515, N2002);
buf BUF1 (N2117, N2106);
or OR3 (N2118, N2094, N929, N139);
nor NOR2 (N2119, N2101, N942);
and AND4 (N2120, N2112, N1755, N1371, N2086);
nand NAND3 (N2121, N2117, N20, N1065);
xor XOR2 (N2122, N2109, N1010);
not NOT1 (N2123, N2121);
nor NOR3 (N2124, N2111, N743, N1293);
nor NOR4 (N2125, N2113, N1714, N283, N914);
and AND4 (N2126, N2119, N1702, N108, N1708);
and AND3 (N2127, N2123, N18, N848);
or OR2 (N2128, N2127, N1122);
or OR2 (N2129, N2125, N1295);
nand NAND4 (N2130, N2128, N1356, N116, N623);
nor NOR4 (N2131, N2129, N598, N1398, N1365);
buf BUF1 (N2132, N2124);
nand NAND2 (N2133, N2116, N109);
nand NAND2 (N2134, N2131, N1240);
buf BUF1 (N2135, N2133);
not NOT1 (N2136, N2108);
not NOT1 (N2137, N2122);
not NOT1 (N2138, N2130);
buf BUF1 (N2139, N2120);
or OR4 (N2140, N2137, N1848, N617, N361);
or OR2 (N2141, N2135, N1648);
and AND3 (N2142, N2139, N1103, N1052);
not NOT1 (N2143, N2142);
xor XOR2 (N2144, N2136, N1481);
nor NOR2 (N2145, N2143, N1161);
buf BUF1 (N2146, N2115);
xor XOR2 (N2147, N2132, N170);
and AND2 (N2148, N2147, N1837);
nor NOR4 (N2149, N2148, N448, N1598, N1226);
buf BUF1 (N2150, N2144);
not NOT1 (N2151, N2141);
not NOT1 (N2152, N2140);
nor NOR3 (N2153, N2152, N1720, N192);
or OR3 (N2154, N2138, N1501, N1304);
nand NAND4 (N2155, N2153, N530, N731, N1637);
or OR2 (N2156, N2154, N1990);
xor XOR2 (N2157, N2149, N2083);
xor XOR2 (N2158, N2156, N705);
or OR2 (N2159, N2158, N1116);
or OR3 (N2160, N2157, N1562, N1343);
xor XOR2 (N2161, N2145, N449);
nand NAND3 (N2162, N2118, N314, N161);
buf BUF1 (N2163, N2159);
not NOT1 (N2164, N2151);
not NOT1 (N2165, N2126);
buf BUF1 (N2166, N2161);
nand NAND4 (N2167, N2166, N2064, N174, N574);
and AND4 (N2168, N2164, N1736, N866, N260);
buf BUF1 (N2169, N2165);
and AND4 (N2170, N2160, N1257, N270, N807);
nand NAND2 (N2171, N2150, N398);
nor NOR4 (N2172, N2171, N840, N1772, N1424);
xor XOR2 (N2173, N2162, N286);
nand NAND2 (N2174, N2146, N206);
nand NAND4 (N2175, N2170, N751, N2128, N1001);
not NOT1 (N2176, N2168);
or OR2 (N2177, N2174, N1598);
not NOT1 (N2178, N2169);
nor NOR2 (N2179, N2167, N1986);
nor NOR3 (N2180, N2176, N535, N314);
or OR4 (N2181, N2180, N706, N865, N593);
or OR4 (N2182, N2177, N2051, N1130, N823);
xor XOR2 (N2183, N2178, N474);
or OR2 (N2184, N2155, N1400);
nand NAND2 (N2185, N2184, N1732);
nor NOR2 (N2186, N2134, N743);
and AND3 (N2187, N2173, N340, N906);
nor NOR2 (N2188, N2175, N128);
and AND2 (N2189, N2179, N879);
nand NAND4 (N2190, N2172, N1884, N1119, N1480);
not NOT1 (N2191, N2188);
xor XOR2 (N2192, N2186, N572);
xor XOR2 (N2193, N2192, N605);
or OR4 (N2194, N2183, N1717, N548, N636);
nor NOR4 (N2195, N2194, N209, N1459, N1509);
nor NOR3 (N2196, N2195, N839, N2067);
xor XOR2 (N2197, N2182, N413);
nor NOR2 (N2198, N2190, N328);
or OR3 (N2199, N2163, N951, N1056);
xor XOR2 (N2200, N2197, N1281);
or OR2 (N2201, N2189, N2090);
xor XOR2 (N2202, N2181, N634);
and AND4 (N2203, N2196, N2027, N1697, N413);
nor NOR3 (N2204, N2199, N1830, N1669);
nand NAND3 (N2205, N2185, N1694, N1596);
nor NOR4 (N2206, N2193, N1828, N981, N1199);
not NOT1 (N2207, N2206);
not NOT1 (N2208, N2205);
or OR2 (N2209, N2198, N403);
nor NOR4 (N2210, N2187, N1731, N476, N827);
xor XOR2 (N2211, N2204, N1366);
nor NOR3 (N2212, N2203, N602, N1020);
buf BUF1 (N2213, N2201);
buf BUF1 (N2214, N2207);
buf BUF1 (N2215, N2202);
or OR2 (N2216, N2211, N986);
nand NAND2 (N2217, N2191, N1854);
nor NOR2 (N2218, N2208, N40);
buf BUF1 (N2219, N2209);
nor NOR4 (N2220, N2216, N967, N44, N1682);
buf BUF1 (N2221, N2213);
and AND3 (N2222, N2214, N1482, N1084);
nand NAND3 (N2223, N2218, N712, N17);
xor XOR2 (N2224, N2217, N1359);
or OR4 (N2225, N2219, N398, N2079, N729);
and AND2 (N2226, N2215, N1844);
nand NAND2 (N2227, N2223, N1987);
not NOT1 (N2228, N2222);
buf BUF1 (N2229, N2220);
not NOT1 (N2230, N2226);
buf BUF1 (N2231, N2227);
or OR3 (N2232, N2225, N787, N383);
or OR4 (N2233, N2221, N2063, N1042, N717);
nor NOR3 (N2234, N2224, N1302, N1055);
not NOT1 (N2235, N2228);
or OR4 (N2236, N2235, N255, N1346, N112);
xor XOR2 (N2237, N2200, N1305);
xor XOR2 (N2238, N2234, N1033);
buf BUF1 (N2239, N2212);
buf BUF1 (N2240, N2231);
or OR3 (N2241, N2240, N850, N1622);
not NOT1 (N2242, N2237);
nand NAND2 (N2243, N2229, N92);
not NOT1 (N2244, N2232);
xor XOR2 (N2245, N2233, N1146);
nor NOR3 (N2246, N2210, N207, N1813);
nor NOR4 (N2247, N2246, N2165, N1894, N1146);
not NOT1 (N2248, N2238);
or OR4 (N2249, N2241, N755, N628, N1091);
or OR2 (N2250, N2245, N948);
and AND4 (N2251, N2243, N1041, N1863, N100);
nand NAND4 (N2252, N2239, N1827, N92, N946);
or OR3 (N2253, N2244, N1135, N1070);
nor NOR3 (N2254, N2253, N905, N1681);
buf BUF1 (N2255, N2250);
or OR3 (N2256, N2249, N1260, N1801);
nand NAND2 (N2257, N2247, N1375);
not NOT1 (N2258, N2251);
not NOT1 (N2259, N2252);
buf BUF1 (N2260, N2254);
buf BUF1 (N2261, N2257);
xor XOR2 (N2262, N2259, N1383);
and AND2 (N2263, N2260, N1826);
nand NAND2 (N2264, N2261, N519);
nor NOR3 (N2265, N2263, N1795, N456);
buf BUF1 (N2266, N2230);
or OR2 (N2267, N2266, N530);
not NOT1 (N2268, N2262);
buf BUF1 (N2269, N2268);
and AND4 (N2270, N2269, N2108, N2268, N387);
nand NAND4 (N2271, N2242, N1087, N459, N1792);
nor NOR4 (N2272, N2264, N288, N1613, N40);
xor XOR2 (N2273, N2272, N985);
nor NOR4 (N2274, N2248, N677, N1088, N787);
nand NAND3 (N2275, N2255, N27, N1286);
nor NOR2 (N2276, N2271, N491);
xor XOR2 (N2277, N2236, N222);
nand NAND2 (N2278, N2275, N1323);
or OR3 (N2279, N2274, N932, N756);
nand NAND3 (N2280, N2258, N1802, N906);
or OR4 (N2281, N2277, N1546, N385, N1330);
xor XOR2 (N2282, N2276, N305);
nand NAND4 (N2283, N2265, N1899, N1909, N1225);
nand NAND2 (N2284, N2273, N831);
and AND3 (N2285, N2280, N1764, N953);
xor XOR2 (N2286, N2279, N2102);
or OR3 (N2287, N2278, N613, N1641);
nor NOR3 (N2288, N2287, N1256, N2154);
xor XOR2 (N2289, N2284, N1260);
nor NOR3 (N2290, N2281, N2107, N474);
not NOT1 (N2291, N2282);
xor XOR2 (N2292, N2270, N185);
and AND3 (N2293, N2267, N90, N1039);
buf BUF1 (N2294, N2293);
nand NAND2 (N2295, N2283, N700);
xor XOR2 (N2296, N2285, N1048);
nor NOR3 (N2297, N2290, N1260, N1188);
and AND2 (N2298, N2289, N785);
nor NOR4 (N2299, N2291, N468, N2113, N796);
not NOT1 (N2300, N2294);
nand NAND3 (N2301, N2288, N817, N1873);
nand NAND3 (N2302, N2256, N1619, N652);
buf BUF1 (N2303, N2300);
not NOT1 (N2304, N2298);
not NOT1 (N2305, N2292);
xor XOR2 (N2306, N2299, N810);
not NOT1 (N2307, N2305);
nand NAND4 (N2308, N2306, N113, N427, N556);
or OR2 (N2309, N2295, N127);
or OR4 (N2310, N2296, N1139, N569, N1999);
nand NAND4 (N2311, N2297, N1032, N148, N1502);
and AND3 (N2312, N2310, N188, N1290);
buf BUF1 (N2313, N2301);
nor NOR4 (N2314, N2311, N1350, N1493, N1454);
and AND4 (N2315, N2309, N1434, N153, N1803);
nand NAND4 (N2316, N2308, N1887, N974, N1232);
xor XOR2 (N2317, N2307, N697);
buf BUF1 (N2318, N2312);
nor NOR2 (N2319, N2315, N894);
or OR3 (N2320, N2314, N1585, N220);
nor NOR3 (N2321, N2313, N625, N814);
or OR4 (N2322, N2316, N1984, N1726, N1164);
buf BUF1 (N2323, N2302);
nand NAND3 (N2324, N2318, N2223, N2004);
xor XOR2 (N2325, N2324, N1951);
nand NAND3 (N2326, N2303, N861, N919);
nor NOR4 (N2327, N2286, N879, N1411, N1401);
nand NAND3 (N2328, N2320, N2159, N720);
xor XOR2 (N2329, N2322, N202);
buf BUF1 (N2330, N2327);
not NOT1 (N2331, N2319);
buf BUF1 (N2332, N2317);
and AND2 (N2333, N2331, N735);
not NOT1 (N2334, N2326);
nor NOR2 (N2335, N2334, N297);
xor XOR2 (N2336, N2329, N1750);
or OR4 (N2337, N2325, N2098, N1470, N1750);
not NOT1 (N2338, N2335);
buf BUF1 (N2339, N2337);
buf BUF1 (N2340, N2328);
nand NAND4 (N2341, N2323, N483, N1015, N1795);
nor NOR3 (N2342, N2338, N767, N1824);
nand NAND4 (N2343, N2330, N197, N1659, N820);
buf BUF1 (N2344, N2336);
buf BUF1 (N2345, N2332);
nor NOR4 (N2346, N2304, N1483, N1422, N942);
not NOT1 (N2347, N2342);
xor XOR2 (N2348, N2343, N2032);
or OR4 (N2349, N2345, N936, N480, N640);
buf BUF1 (N2350, N2346);
or OR2 (N2351, N2333, N874);
or OR4 (N2352, N2341, N1423, N536, N469);
buf BUF1 (N2353, N2350);
and AND4 (N2354, N2347, N2213, N241, N1700);
and AND3 (N2355, N2351, N1694, N759);
and AND2 (N2356, N2321, N765);
and AND3 (N2357, N2356, N523, N577);
or OR2 (N2358, N2352, N1871);
or OR3 (N2359, N2348, N2010, N1585);
and AND2 (N2360, N2358, N312);
or OR2 (N2361, N2340, N1519);
not NOT1 (N2362, N2353);
not NOT1 (N2363, N2349);
xor XOR2 (N2364, N2361, N506);
and AND2 (N2365, N2363, N229);
nand NAND3 (N2366, N2364, N1210, N708);
nand NAND2 (N2367, N2362, N2082);
not NOT1 (N2368, N2365);
nand NAND3 (N2369, N2357, N1061, N2155);
nor NOR2 (N2370, N2367, N1062);
nand NAND4 (N2371, N2359, N2014, N291, N254);
or OR4 (N2372, N2344, N1577, N598, N184);
nand NAND2 (N2373, N2371, N1213);
xor XOR2 (N2374, N2372, N246);
nor NOR4 (N2375, N2368, N55, N1287, N2022);
buf BUF1 (N2376, N2373);
or OR3 (N2377, N2375, N1697, N1907);
nand NAND2 (N2378, N2374, N1073);
nand NAND3 (N2379, N2360, N858, N571);
nor NOR4 (N2380, N2376, N1329, N1779, N197);
xor XOR2 (N2381, N2370, N350);
xor XOR2 (N2382, N2380, N249);
and AND3 (N2383, N2381, N1442, N213);
not NOT1 (N2384, N2369);
and AND2 (N2385, N2355, N2244);
buf BUF1 (N2386, N2378);
nand NAND3 (N2387, N2383, N507, N705);
nand NAND3 (N2388, N2354, N1295, N1120);
nor NOR4 (N2389, N2386, N515, N1128, N1200);
nand NAND3 (N2390, N2388, N1813, N1391);
buf BUF1 (N2391, N2379);
nor NOR4 (N2392, N2366, N1748, N1794, N1853);
nor NOR3 (N2393, N2384, N1547, N236);
or OR3 (N2394, N2392, N2345, N223);
nor NOR2 (N2395, N2377, N1760);
or OR4 (N2396, N2395, N2268, N428, N1251);
buf BUF1 (N2397, N2394);
not NOT1 (N2398, N2382);
buf BUF1 (N2399, N2385);
buf BUF1 (N2400, N2399);
buf BUF1 (N2401, N2397);
not NOT1 (N2402, N2393);
or OR4 (N2403, N2390, N2349, N50, N2331);
not NOT1 (N2404, N2389);
not NOT1 (N2405, N2387);
nand NAND4 (N2406, N2404, N2209, N1952, N949);
or OR3 (N2407, N2396, N370, N1481);
nand NAND3 (N2408, N2405, N1440, N2029);
or OR2 (N2409, N2391, N204);
and AND4 (N2410, N2403, N1676, N1769, N1601);
xor XOR2 (N2411, N2408, N1769);
xor XOR2 (N2412, N2410, N1515);
nor NOR4 (N2413, N2400, N457, N671, N1766);
buf BUF1 (N2414, N2406);
and AND3 (N2415, N2412, N412, N1060);
or OR4 (N2416, N2415, N1389, N712, N1567);
not NOT1 (N2417, N2416);
xor XOR2 (N2418, N2417, N1749);
buf BUF1 (N2419, N2398);
buf BUF1 (N2420, N2401);
and AND4 (N2421, N2420, N1051, N2348, N2124);
or OR2 (N2422, N2413, N859);
or OR3 (N2423, N2411, N365, N2311);
and AND4 (N2424, N2339, N1378, N1769, N683);
nand NAND2 (N2425, N2423, N215);
or OR2 (N2426, N2409, N894);
and AND3 (N2427, N2422, N2016, N666);
not NOT1 (N2428, N2426);
or OR3 (N2429, N2419, N695, N1594);
nand NAND4 (N2430, N2425, N608, N577, N650);
buf BUF1 (N2431, N2429);
nor NOR2 (N2432, N2427, N1966);
xor XOR2 (N2433, N2428, N931);
and AND4 (N2434, N2407, N469, N380, N2072);
or OR4 (N2435, N2431, N1795, N1760, N1103);
nor NOR4 (N2436, N2402, N1198, N1243, N1858);
nor NOR2 (N2437, N2434, N1212);
or OR4 (N2438, N2432, N1460, N1926, N584);
buf BUF1 (N2439, N2435);
not NOT1 (N2440, N2414);
or OR4 (N2441, N2430, N1388, N1916, N2017);
not NOT1 (N2442, N2437);
not NOT1 (N2443, N2442);
nand NAND4 (N2444, N2441, N2061, N867, N732);
and AND2 (N2445, N2436, N511);
nor NOR3 (N2446, N2440, N135, N2432);
nand NAND2 (N2447, N2439, N1936);
xor XOR2 (N2448, N2447, N207);
or OR4 (N2449, N2443, N1495, N1037, N592);
and AND2 (N2450, N2446, N1959);
not NOT1 (N2451, N2444);
not NOT1 (N2452, N2433);
and AND4 (N2453, N2418, N961, N882, N419);
and AND2 (N2454, N2450, N751);
not NOT1 (N2455, N2448);
or OR3 (N2456, N2445, N594, N1204);
xor XOR2 (N2457, N2455, N1288);
xor XOR2 (N2458, N2449, N2308);
xor XOR2 (N2459, N2457, N1543);
buf BUF1 (N2460, N2458);
or OR4 (N2461, N2424, N25, N1291, N1098);
or OR3 (N2462, N2453, N1093, N570);
not NOT1 (N2463, N2456);
or OR3 (N2464, N2461, N1280, N1712);
xor XOR2 (N2465, N2460, N1754);
xor XOR2 (N2466, N2421, N1191);
not NOT1 (N2467, N2438);
buf BUF1 (N2468, N2467);
buf BUF1 (N2469, N2465);
nor NOR4 (N2470, N2451, N448, N1588, N195);
nor NOR3 (N2471, N2468, N1422, N1495);
xor XOR2 (N2472, N2459, N1623);
or OR2 (N2473, N2462, N294);
or OR3 (N2474, N2471, N763, N1565);
and AND3 (N2475, N2454, N1140, N1901);
buf BUF1 (N2476, N2473);
nor NOR3 (N2477, N2474, N385, N1992);
xor XOR2 (N2478, N2470, N2323);
or OR4 (N2479, N2469, N316, N731, N580);
nor NOR4 (N2480, N2463, N538, N999, N483);
nor NOR3 (N2481, N2480, N261, N1953);
and AND2 (N2482, N2476, N197);
not NOT1 (N2483, N2452);
buf BUF1 (N2484, N2478);
or OR3 (N2485, N2483, N575, N1578);
not NOT1 (N2486, N2484);
nand NAND2 (N2487, N2479, N730);
and AND2 (N2488, N2477, N1968);
nor NOR2 (N2489, N2475, N1181);
nand NAND3 (N2490, N2464, N382, N1814);
xor XOR2 (N2491, N2485, N2399);
buf BUF1 (N2492, N2472);
not NOT1 (N2493, N2487);
buf BUF1 (N2494, N2486);
and AND3 (N2495, N2482, N658, N1143);
nor NOR3 (N2496, N2491, N921, N1553);
or OR3 (N2497, N2466, N2165, N2487);
and AND2 (N2498, N2481, N76);
xor XOR2 (N2499, N2494, N2347);
buf BUF1 (N2500, N2496);
not NOT1 (N2501, N2490);
or OR2 (N2502, N2497, N1034);
buf BUF1 (N2503, N2488);
not NOT1 (N2504, N2492);
not NOT1 (N2505, N2493);
or OR2 (N2506, N2501, N447);
and AND4 (N2507, N2505, N33, N2415, N962);
and AND2 (N2508, N2502, N1317);
nand NAND3 (N2509, N2498, N508, N713);
and AND3 (N2510, N2489, N1896, N2457);
or OR4 (N2511, N2506, N514, N682, N919);
xor XOR2 (N2512, N2504, N2309);
buf BUF1 (N2513, N2508);
xor XOR2 (N2514, N2512, N2263);
buf BUF1 (N2515, N2510);
not NOT1 (N2516, N2511);
nor NOR3 (N2517, N2509, N706, N875);
not NOT1 (N2518, N2500);
nor NOR4 (N2519, N2507, N2079, N2256, N1946);
and AND3 (N2520, N2503, N2346, N1972);
nand NAND3 (N2521, N2516, N545, N1632);
not NOT1 (N2522, N2515);
and AND4 (N2523, N2518, N653, N1753, N550);
nand NAND3 (N2524, N2495, N2295, N783);
buf BUF1 (N2525, N2522);
nand NAND2 (N2526, N2519, N1783);
not NOT1 (N2527, N2521);
and AND2 (N2528, N2520, N718);
and AND4 (N2529, N2525, N861, N933, N1610);
not NOT1 (N2530, N2528);
nor NOR2 (N2531, N2527, N1958);
not NOT1 (N2532, N2514);
or OR4 (N2533, N2529, N355, N1820, N1197);
xor XOR2 (N2534, N2524, N953);
buf BUF1 (N2535, N2526);
nor NOR4 (N2536, N2530, N2231, N2531, N2099);
buf BUF1 (N2537, N2209);
xor XOR2 (N2538, N2513, N1129);
nand NAND4 (N2539, N2533, N1456, N1514, N1354);
nand NAND3 (N2540, N2537, N251, N499);
nand NAND4 (N2541, N2499, N2086, N1098, N2256);
xor XOR2 (N2542, N2523, N788);
or OR4 (N2543, N2540, N2159, N1232, N55);
xor XOR2 (N2544, N2532, N2523);
nand NAND2 (N2545, N2534, N1098);
or OR2 (N2546, N2543, N1520);
and AND4 (N2547, N2538, N2159, N1493, N1984);
nand NAND2 (N2548, N2541, N1655);
and AND3 (N2549, N2545, N1785, N2001);
nand NAND2 (N2550, N2544, N59);
nor NOR4 (N2551, N2535, N2347, N1397, N1363);
nor NOR2 (N2552, N2550, N1261);
nand NAND3 (N2553, N2546, N42, N1614);
buf BUF1 (N2554, N2539);
or OR4 (N2555, N2542, N2101, N67, N714);
nor NOR4 (N2556, N2554, N2180, N2273, N1378);
or OR4 (N2557, N2556, N308, N628, N1552);
not NOT1 (N2558, N2553);
buf BUF1 (N2559, N2558);
not NOT1 (N2560, N2551);
or OR2 (N2561, N2548, N1110);
not NOT1 (N2562, N2555);
xor XOR2 (N2563, N2560, N1495);
buf BUF1 (N2564, N2557);
nor NOR4 (N2565, N2559, N2514, N492, N598);
and AND2 (N2566, N2549, N2564);
nand NAND3 (N2567, N1303, N1433, N111);
nor NOR2 (N2568, N2566, N2453);
and AND3 (N2569, N2562, N10, N299);
or OR3 (N2570, N2547, N1698, N2278);
or OR3 (N2571, N2561, N469, N144);
xor XOR2 (N2572, N2517, N2246);
nand NAND3 (N2573, N2568, N1499, N1258);
nor NOR3 (N2574, N2565, N2400, N211);
buf BUF1 (N2575, N2573);
not NOT1 (N2576, N2574);
xor XOR2 (N2577, N2570, N1806);
nor NOR3 (N2578, N2575, N1755, N1555);
xor XOR2 (N2579, N2572, N2068);
or OR2 (N2580, N2563, N420);
and AND2 (N2581, N2552, N2326);
nand NAND3 (N2582, N2579, N2230, N2411);
xor XOR2 (N2583, N2567, N786);
nand NAND4 (N2584, N2569, N2471, N1066, N1620);
xor XOR2 (N2585, N2576, N1604);
or OR3 (N2586, N2536, N1759, N483);
nor NOR4 (N2587, N2584, N2016, N741, N1168);
not NOT1 (N2588, N2585);
not NOT1 (N2589, N2582);
nor NOR3 (N2590, N2587, N1582, N2427);
or OR3 (N2591, N2580, N2517, N1070);
nor NOR2 (N2592, N2590, N670);
nor NOR2 (N2593, N2577, N2285);
nor NOR2 (N2594, N2592, N1241);
nand NAND2 (N2595, N2593, N268);
xor XOR2 (N2596, N2586, N384);
nand NAND3 (N2597, N2591, N2570, N365);
nand NAND3 (N2598, N2596, N1160, N1136);
or OR4 (N2599, N2588, N803, N572, N669);
nor NOR3 (N2600, N2599, N2140, N2198);
nor NOR3 (N2601, N2578, N806, N1634);
not NOT1 (N2602, N2597);
xor XOR2 (N2603, N2598, N2281);
buf BUF1 (N2604, N2602);
nand NAND3 (N2605, N2595, N2082, N2258);
xor XOR2 (N2606, N2600, N1900);
and AND4 (N2607, N2605, N177, N2082, N2231);
not NOT1 (N2608, N2594);
or OR3 (N2609, N2601, N2273, N984);
or OR3 (N2610, N2608, N523, N1668);
nor NOR3 (N2611, N2571, N2240, N513);
or OR4 (N2612, N2583, N977, N2098, N1838);
nand NAND3 (N2613, N2609, N1243, N2111);
xor XOR2 (N2614, N2612, N1399);
nor NOR3 (N2615, N2611, N2089, N580);
nor NOR4 (N2616, N2613, N2291, N1256, N80);
not NOT1 (N2617, N2615);
xor XOR2 (N2618, N2604, N2414);
xor XOR2 (N2619, N2607, N53);
xor XOR2 (N2620, N2603, N2607);
and AND2 (N2621, N2610, N2543);
buf BUF1 (N2622, N2606);
buf BUF1 (N2623, N2619);
or OR2 (N2624, N2617, N1281);
xor XOR2 (N2625, N2581, N877);
not NOT1 (N2626, N2620);
nand NAND2 (N2627, N2623, N82);
nor NOR3 (N2628, N2627, N327, N943);
and AND2 (N2629, N2621, N325);
buf BUF1 (N2630, N2614);
or OR3 (N2631, N2626, N2508, N2556);
buf BUF1 (N2632, N2618);
xor XOR2 (N2633, N2624, N1229);
not NOT1 (N2634, N2631);
or OR3 (N2635, N2628, N2618, N1787);
or OR4 (N2636, N2622, N2224, N1399, N1048);
buf BUF1 (N2637, N2634);
not NOT1 (N2638, N2589);
buf BUF1 (N2639, N2625);
nand NAND2 (N2640, N2636, N2504);
nand NAND2 (N2641, N2630, N1868);
nor NOR4 (N2642, N2641, N1491, N1545, N2536);
and AND2 (N2643, N2637, N2269);
xor XOR2 (N2644, N2642, N872);
buf BUF1 (N2645, N2629);
and AND2 (N2646, N2639, N1040);
and AND3 (N2647, N2633, N2563, N1332);
and AND4 (N2648, N2645, N1358, N2471, N2246);
not NOT1 (N2649, N2638);
xor XOR2 (N2650, N2635, N1755);
nand NAND4 (N2651, N2644, N1215, N827, N1025);
buf BUF1 (N2652, N2646);
or OR2 (N2653, N2650, N1401);
xor XOR2 (N2654, N2647, N1487);
xor XOR2 (N2655, N2616, N1561);
and AND3 (N2656, N2652, N249, N1180);
not NOT1 (N2657, N2654);
xor XOR2 (N2658, N2649, N1165);
not NOT1 (N2659, N2658);
not NOT1 (N2660, N2657);
xor XOR2 (N2661, N2655, N1152);
or OR3 (N2662, N2643, N572, N2249);
nand NAND4 (N2663, N2660, N1543, N1640, N1071);
xor XOR2 (N2664, N2662, N842);
not NOT1 (N2665, N2661);
buf BUF1 (N2666, N2659);
xor XOR2 (N2667, N2656, N1693);
nor NOR2 (N2668, N2667, N104);
not NOT1 (N2669, N2640);
nor NOR2 (N2670, N2651, N2657);
buf BUF1 (N2671, N2648);
nand NAND2 (N2672, N2665, N2596);
not NOT1 (N2673, N2668);
and AND3 (N2674, N2632, N79, N2254);
not NOT1 (N2675, N2670);
not NOT1 (N2676, N2663);
xor XOR2 (N2677, N2675, N1195);
xor XOR2 (N2678, N2653, N2562);
not NOT1 (N2679, N2671);
nor NOR3 (N2680, N2677, N2401, N927);
not NOT1 (N2681, N2664);
and AND4 (N2682, N2681, N1044, N592, N1448);
and AND2 (N2683, N2674, N1997);
not NOT1 (N2684, N2682);
xor XOR2 (N2685, N2666, N84);
and AND3 (N2686, N2672, N2486, N88);
not NOT1 (N2687, N2673);
xor XOR2 (N2688, N2669, N1838);
not NOT1 (N2689, N2679);
or OR3 (N2690, N2688, N2642, N2118);
buf BUF1 (N2691, N2690);
buf BUF1 (N2692, N2687);
and AND3 (N2693, N2684, N2652, N1369);
buf BUF1 (N2694, N2686);
or OR3 (N2695, N2694, N2282, N2618);
or OR4 (N2696, N2693, N999, N1029, N1548);
nand NAND2 (N2697, N2696, N837);
not NOT1 (N2698, N2697);
or OR3 (N2699, N2685, N455, N447);
not NOT1 (N2700, N2683);
and AND2 (N2701, N2698, N1216);
and AND3 (N2702, N2699, N1071, N2187);
nand NAND4 (N2703, N2676, N957, N2560, N692);
and AND2 (N2704, N2689, N1692);
not NOT1 (N2705, N2691);
and AND2 (N2706, N2678, N1874);
xor XOR2 (N2707, N2703, N2408);
nor NOR3 (N2708, N2702, N2495, N1514);
not NOT1 (N2709, N2707);
nor NOR3 (N2710, N2705, N1231, N2701);
not NOT1 (N2711, N539);
nand NAND2 (N2712, N2709, N1420);
xor XOR2 (N2713, N2704, N1570);
or OR2 (N2714, N2692, N1649);
or OR2 (N2715, N2680, N758);
buf BUF1 (N2716, N2715);
and AND4 (N2717, N2714, N651, N2621, N188);
buf BUF1 (N2718, N2716);
nand NAND2 (N2719, N2718, N1992);
nor NOR2 (N2720, N2711, N2476);
nor NOR4 (N2721, N2706, N448, N1005, N275);
xor XOR2 (N2722, N2713, N1267);
nor NOR2 (N2723, N2700, N1626);
nor NOR2 (N2724, N2695, N929);
xor XOR2 (N2725, N2710, N413);
or OR4 (N2726, N2721, N1407, N2012, N1249);
xor XOR2 (N2727, N2725, N355);
buf BUF1 (N2728, N2726);
or OR4 (N2729, N2717, N472, N2512, N1673);
xor XOR2 (N2730, N2708, N1754);
or OR3 (N2731, N2722, N538, N1601);
nand NAND3 (N2732, N2712, N1024, N71);
xor XOR2 (N2733, N2729, N2036);
not NOT1 (N2734, N2730);
xor XOR2 (N2735, N2734, N2478);
or OR2 (N2736, N2727, N2080);
not NOT1 (N2737, N2724);
and AND2 (N2738, N2732, N2699);
buf BUF1 (N2739, N2728);
nor NOR4 (N2740, N2738, N2157, N152, N1219);
or OR2 (N2741, N2733, N966);
or OR2 (N2742, N2720, N1870);
or OR4 (N2743, N2739, N629, N1386, N2190);
nor NOR2 (N2744, N2719, N1455);
xor XOR2 (N2745, N2731, N196);
buf BUF1 (N2746, N2744);
nand NAND3 (N2747, N2743, N934, N2209);
buf BUF1 (N2748, N2737);
buf BUF1 (N2749, N2748);
buf BUF1 (N2750, N2736);
buf BUF1 (N2751, N2746);
nor NOR4 (N2752, N2740, N1121, N1011, N2694);
nand NAND4 (N2753, N2742, N194, N2433, N1797);
nand NAND4 (N2754, N2745, N121, N799, N2215);
buf BUF1 (N2755, N2753);
xor XOR2 (N2756, N2755, N1327);
not NOT1 (N2757, N2751);
nor NOR3 (N2758, N2747, N1322, N598);
nor NOR2 (N2759, N2749, N2601);
not NOT1 (N2760, N2752);
not NOT1 (N2761, N2754);
nor NOR3 (N2762, N2760, N249, N812);
or OR2 (N2763, N2723, N1187);
and AND4 (N2764, N2759, N1317, N534, N1338);
or OR4 (N2765, N2757, N802, N703, N1440);
and AND2 (N2766, N2763, N2467);
nand NAND3 (N2767, N2764, N702, N564);
or OR2 (N2768, N2766, N937);
buf BUF1 (N2769, N2735);
and AND2 (N2770, N2756, N1070);
not NOT1 (N2771, N2741);
nand NAND4 (N2772, N2770, N1047, N1801, N316);
not NOT1 (N2773, N2761);
buf BUF1 (N2774, N2767);
not NOT1 (N2775, N2771);
nand NAND3 (N2776, N2775, N2620, N189);
nand NAND3 (N2777, N2750, N1441, N1997);
nor NOR4 (N2778, N2772, N2692, N1602, N2635);
buf BUF1 (N2779, N2769);
not NOT1 (N2780, N2758);
nand NAND4 (N2781, N2780, N1560, N2097, N401);
not NOT1 (N2782, N2781);
nand NAND2 (N2783, N2762, N1614);
or OR4 (N2784, N2776, N1287, N1444, N2117);
not NOT1 (N2785, N2778);
and AND4 (N2786, N2785, N1860, N348, N1387);
nor NOR3 (N2787, N2777, N2217, N1857);
and AND4 (N2788, N2787, N2703, N2432, N2410);
nand NAND4 (N2789, N2788, N1190, N93, N2095);
and AND2 (N2790, N2768, N103);
and AND2 (N2791, N2782, N2292);
not NOT1 (N2792, N2779);
buf BUF1 (N2793, N2784);
nor NOR4 (N2794, N2773, N2788, N1404, N2643);
xor XOR2 (N2795, N2783, N2434);
buf BUF1 (N2796, N2792);
and AND2 (N2797, N2774, N1786);
nand NAND4 (N2798, N2796, N294, N385, N1946);
nor NOR3 (N2799, N2793, N200, N2569);
and AND3 (N2800, N2794, N2594, N2441);
not NOT1 (N2801, N2799);
nand NAND2 (N2802, N2789, N301);
buf BUF1 (N2803, N2801);
not NOT1 (N2804, N2800);
or OR3 (N2805, N2802, N1377, N433);
nor NOR2 (N2806, N2804, N2368);
not NOT1 (N2807, N2803);
nand NAND2 (N2808, N2786, N2369);
nor NOR4 (N2809, N2795, N2736, N2172, N139);
nand NAND2 (N2810, N2806, N2203);
and AND4 (N2811, N2791, N1632, N1544, N2175);
xor XOR2 (N2812, N2807, N1168);
nand NAND3 (N2813, N2812, N2670, N703);
buf BUF1 (N2814, N2813);
buf BUF1 (N2815, N2810);
xor XOR2 (N2816, N2815, N2463);
buf BUF1 (N2817, N2808);
and AND2 (N2818, N2765, N1613);
or OR2 (N2819, N2811, N1765);
nor NOR4 (N2820, N2805, N198, N1621, N842);
or OR4 (N2821, N2814, N2094, N19, N752);
nor NOR4 (N2822, N2821, N125, N2627, N547);
nand NAND2 (N2823, N2817, N1588);
nand NAND2 (N2824, N2819, N2032);
buf BUF1 (N2825, N2820);
not NOT1 (N2826, N2824);
or OR4 (N2827, N2822, N1295, N1111, N1723);
and AND2 (N2828, N2809, N2381);
not NOT1 (N2829, N2798);
nor NOR4 (N2830, N2823, N2276, N54, N2594);
not NOT1 (N2831, N2797);
or OR4 (N2832, N2816, N2734, N1836, N2825);
nand NAND4 (N2833, N811, N1093, N874, N2720);
xor XOR2 (N2834, N2790, N2563);
nor NOR4 (N2835, N2818, N304, N1828, N194);
not NOT1 (N2836, N2827);
not NOT1 (N2837, N2836);
nor NOR4 (N2838, N2835, N2333, N618, N1024);
nand NAND3 (N2839, N2832, N2471, N2838);
and AND3 (N2840, N853, N1836, N1960);
not NOT1 (N2841, N2828);
buf BUF1 (N2842, N2834);
xor XOR2 (N2843, N2829, N895);
nand NAND4 (N2844, N2830, N875, N1961, N898);
nor NOR2 (N2845, N2833, N2245);
buf BUF1 (N2846, N2839);
nand NAND2 (N2847, N2843, N2357);
xor XOR2 (N2848, N2831, N2339);
buf BUF1 (N2849, N2844);
buf BUF1 (N2850, N2847);
nor NOR3 (N2851, N2846, N1129, N735);
or OR2 (N2852, N2826, N1486);
xor XOR2 (N2853, N2840, N48);
xor XOR2 (N2854, N2842, N240);
and AND3 (N2855, N2841, N511, N1390);
not NOT1 (N2856, N2849);
not NOT1 (N2857, N2845);
buf BUF1 (N2858, N2848);
xor XOR2 (N2859, N2857, N1802);
xor XOR2 (N2860, N2854, N439);
not NOT1 (N2861, N2858);
not NOT1 (N2862, N2853);
or OR3 (N2863, N2852, N2705, N2670);
nand NAND4 (N2864, N2850, N404, N403, N1668);
xor XOR2 (N2865, N2851, N19);
or OR4 (N2866, N2855, N1818, N1969, N2134);
xor XOR2 (N2867, N2837, N426);
buf BUF1 (N2868, N2867);
not NOT1 (N2869, N2856);
or OR4 (N2870, N2869, N2011, N86, N1705);
or OR2 (N2871, N2865, N1508);
not NOT1 (N2872, N2868);
xor XOR2 (N2873, N2863, N346);
not NOT1 (N2874, N2871);
or OR3 (N2875, N2859, N1235, N2366);
nand NAND2 (N2876, N2866, N2350);
nand NAND3 (N2877, N2864, N750, N423);
and AND3 (N2878, N2874, N2157, N978);
and AND4 (N2879, N2877, N1088, N1614, N1689);
nand NAND4 (N2880, N2879, N2847, N283, N1344);
nand NAND4 (N2881, N2880, N2498, N1416, N1930);
buf BUF1 (N2882, N2881);
not NOT1 (N2883, N2873);
nand NAND4 (N2884, N2882, N788, N488, N563);
or OR3 (N2885, N2884, N2484, N82);
and AND2 (N2886, N2862, N1416);
xor XOR2 (N2887, N2886, N487);
buf BUF1 (N2888, N2875);
xor XOR2 (N2889, N2888, N2020);
and AND2 (N2890, N2860, N667);
nand NAND4 (N2891, N2885, N2120, N464, N1818);
or OR4 (N2892, N2876, N2502, N2652, N2169);
nor NOR4 (N2893, N2887, N1398, N721, N2205);
buf BUF1 (N2894, N2889);
nand NAND2 (N2895, N2870, N285);
buf BUF1 (N2896, N2878);
buf BUF1 (N2897, N2861);
buf BUF1 (N2898, N2897);
nand NAND2 (N2899, N2894, N240);
xor XOR2 (N2900, N2898, N1301);
or OR4 (N2901, N2892, N878, N1149, N2032);
nand NAND2 (N2902, N2896, N966);
nor NOR2 (N2903, N2900, N282);
nor NOR4 (N2904, N2872, N938, N937, N881);
not NOT1 (N2905, N2903);
nor NOR3 (N2906, N2902, N2531, N185);
nor NOR3 (N2907, N2901, N1920, N624);
or OR4 (N2908, N2893, N507, N1965, N1665);
or OR2 (N2909, N2905, N1677);
not NOT1 (N2910, N2908);
nand NAND3 (N2911, N2899, N335, N13);
or OR3 (N2912, N2906, N634, N2823);
buf BUF1 (N2913, N2904);
or OR3 (N2914, N2913, N2258, N818);
or OR2 (N2915, N2909, N362);
nand NAND2 (N2916, N2907, N537);
buf BUF1 (N2917, N2910);
and AND4 (N2918, N2883, N1005, N1379, N2733);
and AND3 (N2919, N2911, N800, N1278);
and AND3 (N2920, N2912, N1966, N2258);
and AND4 (N2921, N2914, N1028, N2642, N1567);
buf BUF1 (N2922, N2919);
nand NAND2 (N2923, N2917, N741);
nor NOR3 (N2924, N2895, N1587, N91);
nand NAND4 (N2925, N2923, N1128, N2556, N2457);
not NOT1 (N2926, N2890);
xor XOR2 (N2927, N2916, N161);
buf BUF1 (N2928, N2915);
xor XOR2 (N2929, N2927, N2340);
nand NAND4 (N2930, N2925, N2100, N1961, N1118);
buf BUF1 (N2931, N2926);
nor NOR4 (N2932, N2920, N467, N1813, N2689);
buf BUF1 (N2933, N2930);
xor XOR2 (N2934, N2932, N2645);
xor XOR2 (N2935, N2891, N800);
or OR3 (N2936, N2918, N1153, N755);
buf BUF1 (N2937, N2933);
nand NAND4 (N2938, N2931, N1822, N1049, N2806);
not NOT1 (N2939, N2935);
nor NOR2 (N2940, N2938, N2429);
and AND2 (N2941, N2921, N347);
buf BUF1 (N2942, N2937);
not NOT1 (N2943, N2924);
or OR2 (N2944, N2936, N1160);
and AND4 (N2945, N2943, N2927, N2144, N526);
xor XOR2 (N2946, N2922, N2388);
or OR3 (N2947, N2944, N462, N129);
nor NOR3 (N2948, N2928, N696, N189);
nand NAND4 (N2949, N2946, N1667, N342, N2295);
and AND4 (N2950, N2942, N2264, N1048, N2795);
buf BUF1 (N2951, N2939);
and AND2 (N2952, N2929, N1822);
and AND3 (N2953, N2952, N1390, N2425);
buf BUF1 (N2954, N2949);
not NOT1 (N2955, N2947);
not NOT1 (N2956, N2945);
or OR2 (N2957, N2951, N545);
buf BUF1 (N2958, N2955);
and AND3 (N2959, N2934, N1664, N1501);
xor XOR2 (N2960, N2957, N1042);
nand NAND2 (N2961, N2954, N1168);
nand NAND2 (N2962, N2941, N233);
buf BUF1 (N2963, N2948);
not NOT1 (N2964, N2958);
buf BUF1 (N2965, N2964);
nand NAND4 (N2966, N2959, N2609, N1010, N2264);
buf BUF1 (N2967, N2956);
or OR3 (N2968, N2940, N884, N2597);
xor XOR2 (N2969, N2960, N739);
or OR4 (N2970, N2950, N2164, N2375, N1970);
nor NOR4 (N2971, N2953, N272, N888, N467);
or OR2 (N2972, N2967, N737);
nor NOR4 (N2973, N2965, N2225, N2912, N50);
buf BUF1 (N2974, N2963);
or OR2 (N2975, N2971, N2703);
nor NOR2 (N2976, N2966, N2346);
not NOT1 (N2977, N2976);
buf BUF1 (N2978, N2962);
buf BUF1 (N2979, N2961);
xor XOR2 (N2980, N2977, N1454);
xor XOR2 (N2981, N2970, N826);
xor XOR2 (N2982, N2973, N2024);
xor XOR2 (N2983, N2969, N1046);
not NOT1 (N2984, N2980);
and AND2 (N2985, N2981, N2586);
or OR4 (N2986, N2984, N2310, N1012, N1999);
xor XOR2 (N2987, N2978, N1107);
buf BUF1 (N2988, N2979);
nor NOR4 (N2989, N2982, N2896, N1116, N2640);
and AND4 (N2990, N2972, N258, N839, N2333);
xor XOR2 (N2991, N2975, N2506);
nor NOR2 (N2992, N2989, N2366);
xor XOR2 (N2993, N2991, N1603);
nor NOR2 (N2994, N2990, N1433);
nor NOR4 (N2995, N2992, N942, N1395, N2709);
buf BUF1 (N2996, N2985);
nor NOR4 (N2997, N2993, N211, N1613, N857);
nor NOR2 (N2998, N2974, N2200);
nand NAND4 (N2999, N2996, N133, N2017, N171);
nor NOR3 (N3000, N2968, N1918, N436);
nor NOR3 (N3001, N2995, N288, N2950);
and AND3 (N3002, N2987, N2093, N291);
buf BUF1 (N3003, N2998);
xor XOR2 (N3004, N3000, N1589);
or OR3 (N3005, N2986, N958, N1736);
or OR2 (N3006, N3005, N723);
nand NAND3 (N3007, N2997, N251, N1389);
nor NOR4 (N3008, N2988, N733, N2647, N505);
not NOT1 (N3009, N3003);
buf BUF1 (N3010, N3006);
and AND2 (N3011, N3002, N2093);
xor XOR2 (N3012, N3009, N2402);
buf BUF1 (N3013, N2999);
not NOT1 (N3014, N3013);
not NOT1 (N3015, N3004);
xor XOR2 (N3016, N2983, N766);
xor XOR2 (N3017, N3001, N2699);
nand NAND3 (N3018, N3016, N576, N1174);
or OR3 (N3019, N2994, N2560, N217);
and AND3 (N3020, N3011, N1494, N1435);
nor NOR4 (N3021, N3007, N2701, N508, N1504);
buf BUF1 (N3022, N3015);
nand NAND4 (N3023, N3018, N2564, N1355, N1303);
nand NAND4 (N3024, N3017, N2406, N120, N1045);
nor NOR4 (N3025, N3008, N1479, N1715, N2436);
not NOT1 (N3026, N3024);
buf BUF1 (N3027, N3014);
not NOT1 (N3028, N3010);
or OR2 (N3029, N3022, N2359);
and AND3 (N3030, N3028, N581, N478);
nor NOR3 (N3031, N3019, N325, N2562);
or OR2 (N3032, N3020, N842);
buf BUF1 (N3033, N3023);
buf BUF1 (N3034, N3032);
nor NOR3 (N3035, N3030, N1236, N1060);
nand NAND3 (N3036, N3035, N82, N2138);
buf BUF1 (N3037, N3025);
not NOT1 (N3038, N3036);
not NOT1 (N3039, N3038);
or OR4 (N3040, N3027, N95, N2854, N1662);
not NOT1 (N3041, N3029);
or OR4 (N3042, N3041, N2025, N1588, N2412);
buf BUF1 (N3043, N3039);
buf BUF1 (N3044, N3031);
nand NAND4 (N3045, N3042, N846, N1886, N270);
and AND2 (N3046, N3040, N52);
or OR3 (N3047, N3034, N1158, N2799);
not NOT1 (N3048, N3046);
or OR4 (N3049, N3045, N1081, N2243, N2907);
and AND2 (N3050, N3026, N2827);
not NOT1 (N3051, N3033);
nand NAND4 (N3052, N3050, N1142, N497, N1223);
not NOT1 (N3053, N3043);
not NOT1 (N3054, N3049);
xor XOR2 (N3055, N3044, N1872);
nand NAND2 (N3056, N3052, N1719);
or OR2 (N3057, N3012, N456);
nor NOR4 (N3058, N3053, N2086, N2225, N1916);
not NOT1 (N3059, N3051);
nor NOR2 (N3060, N3056, N1486);
xor XOR2 (N3061, N3055, N583);
not NOT1 (N3062, N3048);
nor NOR4 (N3063, N3061, N1711, N2157, N692);
nand NAND4 (N3064, N3059, N287, N2486, N1747);
xor XOR2 (N3065, N3047, N2838);
xor XOR2 (N3066, N3060, N1997);
xor XOR2 (N3067, N3064, N212);
buf BUF1 (N3068, N3067);
or OR3 (N3069, N3066, N2863, N960);
and AND2 (N3070, N3021, N1772);
nor NOR4 (N3071, N3063, N2393, N2261, N469);
nor NOR4 (N3072, N3068, N2022, N2978, N1426);
buf BUF1 (N3073, N3037);
and AND4 (N3074, N3062, N685, N888, N1183);
nand NAND3 (N3075, N3054, N3039, N1517);
or OR3 (N3076, N3070, N3069, N2551);
xor XOR2 (N3077, N1539, N1968);
buf BUF1 (N3078, N3076);
buf BUF1 (N3079, N3075);
not NOT1 (N3080, N3074);
or OR2 (N3081, N3073, N2406);
buf BUF1 (N3082, N3065);
not NOT1 (N3083, N3079);
xor XOR2 (N3084, N3081, N1473);
not NOT1 (N3085, N3071);
nand NAND2 (N3086, N3085, N2475);
and AND4 (N3087, N3083, N27, N2072, N2471);
and AND2 (N3088, N3080, N44);
xor XOR2 (N3089, N3082, N2379);
nand NAND2 (N3090, N3088, N1301);
not NOT1 (N3091, N3058);
not NOT1 (N3092, N3078);
buf BUF1 (N3093, N3057);
xor XOR2 (N3094, N3092, N2090);
not NOT1 (N3095, N3077);
or OR4 (N3096, N3094, N2140, N2150, N1805);
and AND3 (N3097, N3086, N210, N324);
or OR3 (N3098, N3089, N2780, N1031);
buf BUF1 (N3099, N3093);
nor NOR2 (N3100, N3099, N137);
not NOT1 (N3101, N3096);
xor XOR2 (N3102, N3101, N2239);
not NOT1 (N3103, N3090);
buf BUF1 (N3104, N3095);
xor XOR2 (N3105, N3091, N2612);
or OR2 (N3106, N3097, N470);
xor XOR2 (N3107, N3105, N1302);
xor XOR2 (N3108, N3106, N99);
nor NOR2 (N3109, N3100, N2234);
xor XOR2 (N3110, N3072, N1754);
buf BUF1 (N3111, N3110);
nand NAND2 (N3112, N3087, N304);
not NOT1 (N3113, N3102);
and AND4 (N3114, N3109, N447, N3075, N2975);
or OR2 (N3115, N3098, N2197);
xor XOR2 (N3116, N3108, N2581);
xor XOR2 (N3117, N3104, N180);
not NOT1 (N3118, N3116);
xor XOR2 (N3119, N3115, N2543);
buf BUF1 (N3120, N3117);
or OR3 (N3121, N3119, N523, N1482);
not NOT1 (N3122, N3107);
xor XOR2 (N3123, N3121, N2662);
nand NAND4 (N3124, N3122, N2687, N2203, N218);
buf BUF1 (N3125, N3114);
nor NOR3 (N3126, N3103, N1265, N2124);
buf BUF1 (N3127, N3118);
nor NOR2 (N3128, N3113, N1743);
or OR3 (N3129, N3123, N2382, N3066);
not NOT1 (N3130, N3129);
nor NOR2 (N3131, N3111, N2647);
nand NAND3 (N3132, N3125, N1742, N1842);
nand NAND3 (N3133, N3128, N1644, N592);
nand NAND3 (N3134, N3112, N1283, N1863);
and AND2 (N3135, N3132, N2902);
not NOT1 (N3136, N3133);
buf BUF1 (N3137, N3131);
or OR4 (N3138, N3137, N1952, N2919, N538);
nor NOR2 (N3139, N3134, N2353);
not NOT1 (N3140, N3084);
buf BUF1 (N3141, N3124);
nor NOR2 (N3142, N3120, N1812);
buf BUF1 (N3143, N3140);
and AND3 (N3144, N3126, N1596, N1001);
not NOT1 (N3145, N3138);
and AND3 (N3146, N3142, N1891, N2569);
buf BUF1 (N3147, N3139);
or OR4 (N3148, N3127, N1766, N2020, N1431);
or OR2 (N3149, N3135, N2959);
nor NOR2 (N3150, N3143, N2987);
buf BUF1 (N3151, N3141);
buf BUF1 (N3152, N3149);
xor XOR2 (N3153, N3152, N865);
not NOT1 (N3154, N3147);
nand NAND2 (N3155, N3153, N698);
not NOT1 (N3156, N3145);
buf BUF1 (N3157, N3136);
xor XOR2 (N3158, N3155, N1534);
and AND2 (N3159, N3146, N570);
nor NOR2 (N3160, N3144, N2079);
buf BUF1 (N3161, N3150);
nand NAND2 (N3162, N3156, N1905);
and AND2 (N3163, N3151, N2178);
not NOT1 (N3164, N3160);
or OR3 (N3165, N3164, N449, N965);
buf BUF1 (N3166, N3163);
xor XOR2 (N3167, N3166, N713);
buf BUF1 (N3168, N3161);
or OR3 (N3169, N3159, N1309, N1365);
not NOT1 (N3170, N3162);
and AND2 (N3171, N3169, N2544);
nor NOR4 (N3172, N3158, N749, N1092, N3069);
xor XOR2 (N3173, N3130, N2217);
or OR3 (N3174, N3172, N2597, N2874);
nor NOR4 (N3175, N3167, N882, N1764, N1316);
nand NAND3 (N3176, N3171, N295, N1142);
buf BUF1 (N3177, N3174);
not NOT1 (N3178, N3168);
and AND3 (N3179, N3157, N1688, N355);
buf BUF1 (N3180, N3175);
not NOT1 (N3181, N3179);
or OR2 (N3182, N3177, N283);
and AND2 (N3183, N3173, N362);
not NOT1 (N3184, N3180);
nand NAND3 (N3185, N3170, N1488, N756);
and AND4 (N3186, N3184, N1436, N136, N2001);
nand NAND4 (N3187, N3148, N2840, N2608, N855);
nand NAND4 (N3188, N3186, N1433, N795, N435);
xor XOR2 (N3189, N3188, N771);
nand NAND4 (N3190, N3176, N442, N855, N2384);
or OR3 (N3191, N3165, N594, N721);
and AND2 (N3192, N3183, N2445);
nand NAND3 (N3193, N3182, N2217, N2446);
buf BUF1 (N3194, N3154);
not NOT1 (N3195, N3190);
nand NAND4 (N3196, N3189, N101, N44, N316);
or OR2 (N3197, N3187, N3043);
xor XOR2 (N3198, N3197, N1202);
or OR2 (N3199, N3196, N181);
nand NAND2 (N3200, N3181, N2152);
or OR3 (N3201, N3178, N1794, N2422);
buf BUF1 (N3202, N3194);
and AND2 (N3203, N3200, N2090);
xor XOR2 (N3204, N3191, N1150);
nand NAND3 (N3205, N3192, N1270, N589);
or OR2 (N3206, N3185, N2314);
nand NAND2 (N3207, N3193, N798);
nor NOR2 (N3208, N3199, N1044);
buf BUF1 (N3209, N3208);
not NOT1 (N3210, N3201);
nand NAND2 (N3211, N3195, N1043);
xor XOR2 (N3212, N3204, N1642);
buf BUF1 (N3213, N3206);
or OR4 (N3214, N3211, N1850, N743, N2398);
not NOT1 (N3215, N3202);
and AND2 (N3216, N3213, N2728);
and AND4 (N3217, N3205, N1683, N2075, N2978);
xor XOR2 (N3218, N3216, N1986);
nor NOR4 (N3219, N3207, N2232, N1077, N1276);
nand NAND4 (N3220, N3198, N2488, N1907, N993);
buf BUF1 (N3221, N3209);
nor NOR3 (N3222, N3215, N1205, N2688);
or OR3 (N3223, N3217, N909, N547);
or OR4 (N3224, N3223, N526, N300, N1889);
buf BUF1 (N3225, N3212);
nand NAND4 (N3226, N3221, N2728, N1887, N1787);
not NOT1 (N3227, N3222);
or OR2 (N3228, N3226, N230);
buf BUF1 (N3229, N3210);
nor NOR4 (N3230, N3203, N2588, N2161, N85);
xor XOR2 (N3231, N3220, N2867);
nor NOR4 (N3232, N3214, N1621, N82, N2895);
buf BUF1 (N3233, N3218);
xor XOR2 (N3234, N3225, N2750);
buf BUF1 (N3235, N3232);
and AND3 (N3236, N3230, N3068, N1912);
and AND4 (N3237, N3233, N2252, N2173, N917);
nor NOR2 (N3238, N3224, N321);
buf BUF1 (N3239, N3219);
or OR4 (N3240, N3235, N2287, N1608, N1182);
and AND2 (N3241, N3231, N1435);
xor XOR2 (N3242, N3236, N1001);
buf BUF1 (N3243, N3238);
or OR4 (N3244, N3229, N1985, N2217, N1223);
and AND4 (N3245, N3239, N1181, N295, N571);
and AND4 (N3246, N3240, N125, N146, N2826);
not NOT1 (N3247, N3246);
and AND2 (N3248, N3245, N1791);
nand NAND4 (N3249, N3248, N1274, N2999, N2534);
xor XOR2 (N3250, N3242, N3173);
xor XOR2 (N3251, N3250, N372);
nor NOR4 (N3252, N3241, N1065, N1724, N1446);
xor XOR2 (N3253, N3237, N1129);
or OR2 (N3254, N3253, N1160);
buf BUF1 (N3255, N3234);
nor NOR2 (N3256, N3251, N2483);
not NOT1 (N3257, N3249);
or OR2 (N3258, N3252, N1004);
and AND3 (N3259, N3255, N2697, N2230);
buf BUF1 (N3260, N3228);
not NOT1 (N3261, N3256);
buf BUF1 (N3262, N3259);
nor NOR3 (N3263, N3244, N2822, N1981);
xor XOR2 (N3264, N3262, N2402);
buf BUF1 (N3265, N3260);
nand NAND4 (N3266, N3263, N1203, N580, N210);
not NOT1 (N3267, N3227);
or OR4 (N3268, N3261, N2722, N68, N1084);
or OR4 (N3269, N3265, N2448, N1882, N2689);
xor XOR2 (N3270, N3257, N1561);
xor XOR2 (N3271, N3254, N429);
not NOT1 (N3272, N3243);
xor XOR2 (N3273, N3268, N1883);
nand NAND2 (N3274, N3267, N1095);
and AND2 (N3275, N3273, N2377);
nand NAND4 (N3276, N3247, N2982, N1151, N293);
xor XOR2 (N3277, N3275, N546);
nand NAND4 (N3278, N3266, N69, N544, N1298);
nor NOR2 (N3279, N3258, N2841);
buf BUF1 (N3280, N3278);
and AND2 (N3281, N3274, N1718);
nor NOR3 (N3282, N3269, N1696, N1240);
buf BUF1 (N3283, N3271);
or OR3 (N3284, N3276, N1350, N874);
buf BUF1 (N3285, N3284);
and AND3 (N3286, N3264, N1744, N868);
nand NAND3 (N3287, N3283, N537, N294);
xor XOR2 (N3288, N3282, N266);
nand NAND3 (N3289, N3270, N2908, N1364);
buf BUF1 (N3290, N3286);
or OR3 (N3291, N3277, N1100, N1293);
or OR3 (N3292, N3291, N2094, N531);
nand NAND2 (N3293, N3292, N505);
nand NAND2 (N3294, N3281, N2925);
nand NAND4 (N3295, N3280, N909, N2626, N30);
nand NAND3 (N3296, N3288, N2593, N3105);
or OR4 (N3297, N3272, N878, N1800, N829);
nor NOR2 (N3298, N3287, N2058);
not NOT1 (N3299, N3294);
nand NAND2 (N3300, N3285, N1169);
or OR3 (N3301, N3299, N706, N381);
and AND4 (N3302, N3293, N1835, N630, N1859);
xor XOR2 (N3303, N3290, N422);
xor XOR2 (N3304, N3298, N789);
nand NAND4 (N3305, N3304, N1779, N788, N340);
not NOT1 (N3306, N3303);
and AND3 (N3307, N3295, N3177, N563);
buf BUF1 (N3308, N3300);
and AND4 (N3309, N3308, N2585, N2715, N180);
not NOT1 (N3310, N3306);
and AND4 (N3311, N3279, N1841, N1141, N3129);
xor XOR2 (N3312, N3310, N42);
not NOT1 (N3313, N3296);
nor NOR2 (N3314, N3301, N2164);
xor XOR2 (N3315, N3297, N1855);
not NOT1 (N3316, N3307);
xor XOR2 (N3317, N3312, N2452);
nor NOR3 (N3318, N3315, N2685, N2505);
buf BUF1 (N3319, N3316);
nand NAND2 (N3320, N3314, N2557);
nand NAND4 (N3321, N3311, N298, N2297, N2491);
or OR4 (N3322, N3320, N1591, N424, N3258);
nor NOR4 (N3323, N3318, N3238, N849, N2917);
and AND4 (N3324, N3289, N2733, N2283, N2478);
or OR2 (N3325, N3309, N1995);
nand NAND2 (N3326, N3324, N263);
xor XOR2 (N3327, N3323, N1912);
and AND3 (N3328, N3327, N1598, N1158);
nand NAND4 (N3329, N3322, N1259, N1090, N148);
buf BUF1 (N3330, N3302);
nor NOR2 (N3331, N3317, N2279);
xor XOR2 (N3332, N3325, N3095);
and AND4 (N3333, N3326, N2235, N2185, N1014);
buf BUF1 (N3334, N3321);
or OR4 (N3335, N3319, N2515, N2749, N1414);
nor NOR2 (N3336, N3331, N592);
buf BUF1 (N3337, N3305);
and AND3 (N3338, N3313, N1860, N2220);
nor NOR3 (N3339, N3329, N2877, N2306);
xor XOR2 (N3340, N3328, N2814);
xor XOR2 (N3341, N3340, N2099);
xor XOR2 (N3342, N3341, N2503);
and AND3 (N3343, N3330, N2536, N2306);
nor NOR3 (N3344, N3338, N1214, N1928);
or OR4 (N3345, N3342, N942, N750, N2289);
and AND4 (N3346, N3336, N1579, N2459, N653);
nor NOR4 (N3347, N3334, N2273, N3300, N234);
buf BUF1 (N3348, N3337);
buf BUF1 (N3349, N3333);
or OR4 (N3350, N3346, N443, N760, N2889);
or OR4 (N3351, N3347, N238, N2131, N1419);
and AND4 (N3352, N3348, N287, N1142, N2554);
buf BUF1 (N3353, N3351);
nor NOR4 (N3354, N3335, N2267, N467, N1079);
and AND2 (N3355, N3353, N3081);
nand NAND2 (N3356, N3345, N748);
nor NOR4 (N3357, N3343, N3248, N2709, N2543);
xor XOR2 (N3358, N3350, N1358);
and AND3 (N3359, N3355, N2637, N1446);
nor NOR4 (N3360, N3339, N1350, N3105, N461);
nor NOR3 (N3361, N3359, N1268, N902);
not NOT1 (N3362, N3349);
or OR2 (N3363, N3357, N1572);
not NOT1 (N3364, N3356);
not NOT1 (N3365, N3358);
buf BUF1 (N3366, N3364);
nand NAND4 (N3367, N3352, N1843, N2301, N2326);
or OR3 (N3368, N3366, N2497, N2648);
nor NOR3 (N3369, N3363, N1217, N106);
nand NAND3 (N3370, N3354, N770, N201);
nand NAND4 (N3371, N3369, N225, N1465, N973);
nand NAND4 (N3372, N3344, N794, N2785, N2002);
not NOT1 (N3373, N3365);
not NOT1 (N3374, N3361);
xor XOR2 (N3375, N3368, N3134);
or OR4 (N3376, N3373, N2483, N1549, N1556);
and AND3 (N3377, N3370, N2658, N3094);
xor XOR2 (N3378, N3374, N1494);
not NOT1 (N3379, N3371);
nand NAND2 (N3380, N3372, N2497);
and AND4 (N3381, N3360, N1207, N2458, N2967);
or OR4 (N3382, N3377, N1337, N1921, N625);
nand NAND4 (N3383, N3378, N1976, N1509, N1061);
buf BUF1 (N3384, N3379);
not NOT1 (N3385, N3362);
not NOT1 (N3386, N3383);
buf BUF1 (N3387, N3386);
and AND2 (N3388, N3385, N195);
xor XOR2 (N3389, N3367, N1206);
or OR2 (N3390, N3381, N1435);
nor NOR2 (N3391, N3375, N2650);
nand NAND3 (N3392, N3387, N2377, N1608);
nor NOR3 (N3393, N3390, N2373, N2621);
and AND3 (N3394, N3384, N2899, N986);
nor NOR3 (N3395, N3389, N3131, N3267);
nand NAND2 (N3396, N3376, N2961);
xor XOR2 (N3397, N3395, N1594);
xor XOR2 (N3398, N3392, N827);
or OR2 (N3399, N3396, N2640);
nand NAND4 (N3400, N3332, N2504, N2917, N355);
or OR4 (N3401, N3397, N3031, N1815, N1551);
buf BUF1 (N3402, N3400);
or OR2 (N3403, N3382, N2803);
not NOT1 (N3404, N3401);
nor NOR3 (N3405, N3399, N2614, N2004);
nand NAND3 (N3406, N3403, N1191, N1021);
not NOT1 (N3407, N3406);
xor XOR2 (N3408, N3394, N948);
nor NOR3 (N3409, N3404, N50, N3327);
nor NOR3 (N3410, N3402, N2283, N2945);
or OR4 (N3411, N3391, N881, N1724, N539);
not NOT1 (N3412, N3393);
or OR4 (N3413, N3410, N2185, N2650, N1022);
nand NAND3 (N3414, N3405, N2450, N2338);
buf BUF1 (N3415, N3414);
buf BUF1 (N3416, N3407);
buf BUF1 (N3417, N3380);
nand NAND4 (N3418, N3398, N933, N1753, N1707);
and AND4 (N3419, N3418, N1787, N3395, N1425);
nand NAND4 (N3420, N3413, N1194, N385, N673);
not NOT1 (N3421, N3409);
buf BUF1 (N3422, N3417);
nor NOR4 (N3423, N3419, N1046, N1073, N2547);
buf BUF1 (N3424, N3408);
not NOT1 (N3425, N3424);
or OR2 (N3426, N3423, N3291);
buf BUF1 (N3427, N3425);
not NOT1 (N3428, N3422);
xor XOR2 (N3429, N3421, N1168);
nor NOR4 (N3430, N3388, N2022, N2508, N154);
nand NAND4 (N3431, N3427, N2620, N1123, N2076);
or OR4 (N3432, N3426, N3260, N483, N669);
xor XOR2 (N3433, N3428, N959);
buf BUF1 (N3434, N3430);
xor XOR2 (N3435, N3411, N2637);
buf BUF1 (N3436, N3431);
nor NOR4 (N3437, N3436, N346, N2454, N2832);
not NOT1 (N3438, N3435);
and AND2 (N3439, N3420, N2903);
nand NAND4 (N3440, N3433, N899, N523, N2006);
nor NOR3 (N3441, N3432, N2671, N3114);
and AND4 (N3442, N3441, N1218, N2406, N3152);
nand NAND3 (N3443, N3439, N1738, N501);
xor XOR2 (N3444, N3440, N3232);
not NOT1 (N3445, N3444);
xor XOR2 (N3446, N3434, N1123);
not NOT1 (N3447, N3438);
buf BUF1 (N3448, N3446);
nor NOR3 (N3449, N3415, N2474, N259);
and AND2 (N3450, N3442, N1755);
buf BUF1 (N3451, N3429);
and AND2 (N3452, N3437, N934);
buf BUF1 (N3453, N3450);
nand NAND2 (N3454, N3447, N83);
or OR4 (N3455, N3412, N2357, N2736, N1539);
buf BUF1 (N3456, N3416);
nor NOR2 (N3457, N3443, N651);
buf BUF1 (N3458, N3453);
not NOT1 (N3459, N3455);
not NOT1 (N3460, N3448);
xor XOR2 (N3461, N3452, N2577);
xor XOR2 (N3462, N3445, N2588);
and AND4 (N3463, N3462, N1709, N551, N943);
nand NAND4 (N3464, N3449, N3100, N3371, N1922);
or OR3 (N3465, N3461, N562, N311);
not NOT1 (N3466, N3457);
and AND4 (N3467, N3460, N951, N3174, N3026);
or OR2 (N3468, N3463, N1503);
xor XOR2 (N3469, N3451, N1390);
nor NOR3 (N3470, N3466, N794, N562);
and AND4 (N3471, N3468, N2198, N2418, N1886);
nor NOR2 (N3472, N3464, N2686);
and AND2 (N3473, N3458, N3040);
and AND4 (N3474, N3470, N2863, N1719, N846);
nand NAND2 (N3475, N3469, N210);
buf BUF1 (N3476, N3473);
buf BUF1 (N3477, N3476);
and AND4 (N3478, N3474, N1124, N3385, N693);
and AND2 (N3479, N3477, N742);
buf BUF1 (N3480, N3478);
nand NAND4 (N3481, N3465, N2269, N2654, N411);
xor XOR2 (N3482, N3475, N1504);
nand NAND3 (N3483, N3471, N437, N1808);
nor NOR4 (N3484, N3472, N2650, N1613, N556);
xor XOR2 (N3485, N3482, N2114);
nor NOR4 (N3486, N3456, N1371, N2619, N1971);
nand NAND2 (N3487, N3467, N3049);
not NOT1 (N3488, N3486);
not NOT1 (N3489, N3479);
xor XOR2 (N3490, N3488, N3213);
or OR3 (N3491, N3454, N66, N3138);
nor NOR2 (N3492, N3459, N1446);
and AND3 (N3493, N3491, N3488, N3150);
nand NAND2 (N3494, N3483, N2930);
nor NOR2 (N3495, N3487, N2076);
nor NOR3 (N3496, N3494, N3434, N2723);
xor XOR2 (N3497, N3492, N186);
buf BUF1 (N3498, N3490);
xor XOR2 (N3499, N3480, N1730);
xor XOR2 (N3500, N3485, N2444);
not NOT1 (N3501, N3489);
nor NOR4 (N3502, N3495, N2183, N501, N2373);
xor XOR2 (N3503, N3502, N1802);
xor XOR2 (N3504, N3484, N1169);
nand NAND4 (N3505, N3501, N3049, N1186, N380);
or OR2 (N3506, N3504, N765);
buf BUF1 (N3507, N3500);
buf BUF1 (N3508, N3497);
nor NOR2 (N3509, N3493, N918);
nand NAND3 (N3510, N3505, N625, N1305);
and AND3 (N3511, N3496, N3086, N179);
xor XOR2 (N3512, N3507, N415);
buf BUF1 (N3513, N3508);
xor XOR2 (N3514, N3513, N2022);
or OR2 (N3515, N3481, N3411);
xor XOR2 (N3516, N3512, N2075);
xor XOR2 (N3517, N3516, N360);
and AND3 (N3518, N3510, N3152, N2992);
xor XOR2 (N3519, N3515, N2020);
nor NOR2 (N3520, N3517, N1908);
xor XOR2 (N3521, N3509, N2291);
nand NAND3 (N3522, N3520, N2088, N163);
nand NAND3 (N3523, N3506, N881, N11);
xor XOR2 (N3524, N3518, N2532);
or OR3 (N3525, N3511, N3349, N1091);
xor XOR2 (N3526, N3523, N2366);
nand NAND4 (N3527, N3498, N3193, N3054, N470);
nand NAND3 (N3528, N3525, N30, N3095);
and AND4 (N3529, N3503, N816, N2303, N1348);
or OR4 (N3530, N3522, N2110, N34, N3265);
nor NOR4 (N3531, N3514, N2716, N2885, N1317);
buf BUF1 (N3532, N3529);
nor NOR4 (N3533, N3521, N842, N2530, N3475);
and AND4 (N3534, N3524, N1069, N1689, N1644);
nor NOR4 (N3535, N3534, N58, N906, N560);
nand NAND4 (N3536, N3533, N3169, N3258, N3010);
and AND2 (N3537, N3519, N1030);
nand NAND2 (N3538, N3536, N1355);
xor XOR2 (N3539, N3499, N3197);
xor XOR2 (N3540, N3538, N2956);
nand NAND4 (N3541, N3527, N2922, N1387, N1547);
nor NOR3 (N3542, N3539, N10, N2026);
not NOT1 (N3543, N3528);
xor XOR2 (N3544, N3542, N564);
nand NAND3 (N3545, N3537, N732, N2605);
buf BUF1 (N3546, N3530);
nand NAND2 (N3547, N3526, N673);
xor XOR2 (N3548, N3545, N122);
buf BUF1 (N3549, N3547);
nor NOR4 (N3550, N3549, N1375, N3035, N1558);
nor NOR3 (N3551, N3548, N1961, N2504);
not NOT1 (N3552, N3550);
or OR4 (N3553, N3532, N1864, N554, N2290);
nor NOR3 (N3554, N3552, N858, N1735);
buf BUF1 (N3555, N3544);
buf BUF1 (N3556, N3540);
and AND2 (N3557, N3556, N860);
nand NAND3 (N3558, N3557, N1459, N1269);
nand NAND2 (N3559, N3554, N964);
or OR3 (N3560, N3555, N1909, N2423);
and AND2 (N3561, N3546, N2515);
not NOT1 (N3562, N3531);
xor XOR2 (N3563, N3541, N2159);
xor XOR2 (N3564, N3535, N1607);
not NOT1 (N3565, N3562);
xor XOR2 (N3566, N3559, N3298);
buf BUF1 (N3567, N3551);
nor NOR3 (N3568, N3565, N2920, N1977);
nor NOR3 (N3569, N3568, N787, N1107);
nand NAND2 (N3570, N3564, N1255);
xor XOR2 (N3571, N3569, N628);
nand NAND2 (N3572, N3560, N2116);
xor XOR2 (N3573, N3566, N2329);
and AND3 (N3574, N3543, N677, N274);
xor XOR2 (N3575, N3571, N3042);
buf BUF1 (N3576, N3567);
nor NOR3 (N3577, N3573, N2020, N2203);
or OR3 (N3578, N3563, N3020, N3056);
not NOT1 (N3579, N3576);
nand NAND2 (N3580, N3561, N286);
not NOT1 (N3581, N3577);
nor NOR2 (N3582, N3575, N1573);
nand NAND3 (N3583, N3570, N424, N1606);
nand NAND2 (N3584, N3579, N1376);
or OR2 (N3585, N3580, N2170);
nor NOR2 (N3586, N3574, N266);
or OR3 (N3587, N3585, N339, N2408);
or OR2 (N3588, N3558, N1435);
nand NAND4 (N3589, N3586, N2524, N1517, N3443);
xor XOR2 (N3590, N3581, N1527);
buf BUF1 (N3591, N3572);
not NOT1 (N3592, N3589);
nand NAND4 (N3593, N3578, N908, N3355, N270);
buf BUF1 (N3594, N3584);
or OR2 (N3595, N3594, N2224);
or OR4 (N3596, N3582, N2910, N2045, N2742);
or OR2 (N3597, N3588, N593);
buf BUF1 (N3598, N3590);
nor NOR3 (N3599, N3587, N585, N648);
and AND3 (N3600, N3599, N3370, N1865);
nand NAND3 (N3601, N3598, N1017, N1187);
nand NAND2 (N3602, N3596, N1289);
or OR2 (N3603, N3601, N2883);
xor XOR2 (N3604, N3583, N244);
or OR2 (N3605, N3595, N3051);
buf BUF1 (N3606, N3597);
nor NOR2 (N3607, N3606, N692);
buf BUF1 (N3608, N3604);
xor XOR2 (N3609, N3605, N1793);
or OR2 (N3610, N3607, N1855);
not NOT1 (N3611, N3608);
buf BUF1 (N3612, N3603);
buf BUF1 (N3613, N3553);
buf BUF1 (N3614, N3602);
nor NOR3 (N3615, N3609, N447, N474);
nor NOR3 (N3616, N3592, N443, N2673);
or OR4 (N3617, N3591, N2452, N1155, N856);
nand NAND2 (N3618, N3600, N1437);
not NOT1 (N3619, N3613);
and AND4 (N3620, N3615, N2403, N2904, N1349);
and AND4 (N3621, N3617, N1165, N3394, N2995);
not NOT1 (N3622, N3616);
or OR2 (N3623, N3610, N3317);
nor NOR4 (N3624, N3612, N2883, N3142, N175);
xor XOR2 (N3625, N3619, N769);
xor XOR2 (N3626, N3623, N1851);
nand NAND2 (N3627, N3618, N354);
buf BUF1 (N3628, N3620);
or OR2 (N3629, N3627, N1826);
or OR3 (N3630, N3611, N2984, N2582);
nor NOR2 (N3631, N3625, N2660);
nor NOR4 (N3632, N3630, N680, N187, N255);
nor NOR3 (N3633, N3631, N576, N1165);
nand NAND3 (N3634, N3628, N1017, N480);
buf BUF1 (N3635, N3634);
not NOT1 (N3636, N3621);
nor NOR4 (N3637, N3614, N2523, N1280, N789);
nor NOR3 (N3638, N3622, N1, N937);
nor NOR3 (N3639, N3638, N3231, N66);
nand NAND3 (N3640, N3636, N608, N2157);
buf BUF1 (N3641, N3640);
or OR4 (N3642, N3624, N323, N2974, N1923);
xor XOR2 (N3643, N3642, N3550);
or OR2 (N3644, N3643, N2978);
and AND4 (N3645, N3593, N2348, N1275, N2485);
not NOT1 (N3646, N3635);
nand NAND3 (N3647, N3646, N1790, N121);
xor XOR2 (N3648, N3637, N1633);
nor NOR2 (N3649, N3626, N841);
not NOT1 (N3650, N3632);
buf BUF1 (N3651, N3647);
and AND2 (N3652, N3641, N1211);
and AND3 (N3653, N3648, N3117, N1568);
nand NAND4 (N3654, N3629, N3617, N581, N1600);
nand NAND2 (N3655, N3645, N1475);
buf BUF1 (N3656, N3644);
nor NOR4 (N3657, N3654, N1047, N722, N2181);
or OR2 (N3658, N3655, N2889);
not NOT1 (N3659, N3656);
nor NOR3 (N3660, N3651, N2727, N1027);
xor XOR2 (N3661, N3657, N2482);
or OR2 (N3662, N3649, N300);
xor XOR2 (N3663, N3658, N1871);
not NOT1 (N3664, N3652);
nor NOR3 (N3665, N3650, N392, N2176);
nor NOR3 (N3666, N3653, N2493, N1832);
nand NAND3 (N3667, N3661, N1374, N3547);
nor NOR2 (N3668, N3666, N1390);
not NOT1 (N3669, N3659);
and AND4 (N3670, N3664, N3312, N1401, N2085);
and AND4 (N3671, N3660, N3231, N1841, N1716);
nor NOR4 (N3672, N3668, N78, N1289, N1735);
xor XOR2 (N3673, N3665, N1650);
or OR4 (N3674, N3670, N1813, N1757, N3291);
nor NOR2 (N3675, N3639, N2266);
or OR2 (N3676, N3672, N1226);
xor XOR2 (N3677, N3662, N560);
nand NAND4 (N3678, N3674, N1555, N2419, N520);
or OR3 (N3679, N3673, N528, N402);
nor NOR4 (N3680, N3678, N331, N3093, N3157);
nor NOR3 (N3681, N3667, N1197, N1559);
not NOT1 (N3682, N3679);
or OR3 (N3683, N3671, N1638, N2144);
buf BUF1 (N3684, N3676);
not NOT1 (N3685, N3669);
nor NOR3 (N3686, N3633, N1127, N2635);
xor XOR2 (N3687, N3677, N1748);
xor XOR2 (N3688, N3686, N127);
nor NOR4 (N3689, N3682, N1459, N2765, N1326);
or OR3 (N3690, N3675, N2702, N3170);
or OR3 (N3691, N3687, N3044, N424);
or OR2 (N3692, N3685, N1117);
nand NAND4 (N3693, N3688, N2181, N1409, N3481);
and AND3 (N3694, N3681, N3094, N140);
buf BUF1 (N3695, N3680);
buf BUF1 (N3696, N3694);
nor NOR3 (N3697, N3683, N1658, N1386);
or OR3 (N3698, N3663, N2015, N2911);
or OR3 (N3699, N3692, N3268, N2490);
nand NAND3 (N3700, N3699, N1443, N1290);
and AND2 (N3701, N3700, N528);
or OR2 (N3702, N3698, N1306);
buf BUF1 (N3703, N3695);
nor NOR3 (N3704, N3691, N484, N3086);
nor NOR4 (N3705, N3693, N292, N152, N126);
xor XOR2 (N3706, N3702, N1995);
or OR4 (N3707, N3697, N2235, N156, N1843);
or OR4 (N3708, N3707, N310, N1062, N429);
and AND3 (N3709, N3705, N1361, N3142);
nand NAND2 (N3710, N3696, N3549);
or OR4 (N3711, N3703, N1850, N360, N1869);
nor NOR2 (N3712, N3704, N2572);
buf BUF1 (N3713, N3709);
or OR4 (N3714, N3689, N1708, N3405, N3411);
not NOT1 (N3715, N3714);
buf BUF1 (N3716, N3715);
not NOT1 (N3717, N3716);
nor NOR4 (N3718, N3690, N1296, N568, N3667);
buf BUF1 (N3719, N3711);
nand NAND2 (N3720, N3717, N1149);
or OR2 (N3721, N3684, N2055);
or OR4 (N3722, N3712, N2976, N1899, N633);
xor XOR2 (N3723, N3701, N2542);
buf BUF1 (N3724, N3713);
or OR4 (N3725, N3706, N161, N802, N3184);
nor NOR4 (N3726, N3710, N1342, N3151, N2410);
nand NAND3 (N3727, N3726, N2518, N3594);
nand NAND4 (N3728, N3720, N963, N556, N2616);
buf BUF1 (N3729, N3719);
not NOT1 (N3730, N3725);
nor NOR4 (N3731, N3730, N685, N2447, N3532);
or OR2 (N3732, N3718, N462);
not NOT1 (N3733, N3728);
xor XOR2 (N3734, N3724, N1117);
and AND3 (N3735, N3723, N500, N2538);
and AND2 (N3736, N3729, N1845);
xor XOR2 (N3737, N3721, N970);
nand NAND3 (N3738, N3736, N477, N1302);
buf BUF1 (N3739, N3727);
nor NOR3 (N3740, N3708, N1438, N2831);
buf BUF1 (N3741, N3722);
buf BUF1 (N3742, N3734);
or OR4 (N3743, N3742, N1682, N526, N29);
buf BUF1 (N3744, N3733);
not NOT1 (N3745, N3738);
not NOT1 (N3746, N3743);
nor NOR3 (N3747, N3739, N3385, N2047);
not NOT1 (N3748, N3741);
nor NOR2 (N3749, N3744, N2482);
not NOT1 (N3750, N3746);
nand NAND4 (N3751, N3750, N52, N3589, N3488);
buf BUF1 (N3752, N3747);
nor NOR4 (N3753, N3732, N1160, N525, N592);
or OR2 (N3754, N3745, N1097);
or OR3 (N3755, N3754, N1152, N3689);
not NOT1 (N3756, N3751);
not NOT1 (N3757, N3737);
nor NOR4 (N3758, N3753, N480, N2468, N1229);
xor XOR2 (N3759, N3756, N1935);
buf BUF1 (N3760, N3731);
nand NAND3 (N3761, N3749, N254, N1788);
nand NAND3 (N3762, N3735, N3115, N10);
and AND4 (N3763, N3752, N465, N2036, N2482);
buf BUF1 (N3764, N3755);
xor XOR2 (N3765, N3763, N3432);
or OR4 (N3766, N3761, N1515, N3389, N2177);
buf BUF1 (N3767, N3748);
xor XOR2 (N3768, N3767, N1766);
or OR4 (N3769, N3757, N3271, N843, N3679);
and AND2 (N3770, N3760, N612);
and AND4 (N3771, N3764, N2570, N187, N2286);
xor XOR2 (N3772, N3768, N454);
and AND3 (N3773, N3740, N74, N2466);
nor NOR2 (N3774, N3766, N1672);
xor XOR2 (N3775, N3773, N2450);
buf BUF1 (N3776, N3775);
not NOT1 (N3777, N3762);
and AND3 (N3778, N3765, N561, N30);
xor XOR2 (N3779, N3776, N778);
not NOT1 (N3780, N3759);
nor NOR2 (N3781, N3772, N1544);
buf BUF1 (N3782, N3779);
buf BUF1 (N3783, N3780);
buf BUF1 (N3784, N3774);
nor NOR4 (N3785, N3770, N3503, N1558, N2839);
not NOT1 (N3786, N3769);
nor NOR3 (N3787, N3785, N1854, N3657);
or OR4 (N3788, N3783, N2364, N3253, N3559);
and AND3 (N3789, N3786, N1132, N3378);
buf BUF1 (N3790, N3778);
or OR2 (N3791, N3790, N68);
nor NOR2 (N3792, N3789, N3044);
and AND3 (N3793, N3784, N1164, N1067);
nand NAND3 (N3794, N3793, N1842, N312);
xor XOR2 (N3795, N3758, N629);
xor XOR2 (N3796, N3771, N2742);
not NOT1 (N3797, N3791);
and AND3 (N3798, N3795, N2620, N1471);
nor NOR2 (N3799, N3796, N2209);
or OR2 (N3800, N3799, N3417);
or OR3 (N3801, N3777, N822, N93);
or OR4 (N3802, N3794, N2415, N1944, N58);
nand NAND3 (N3803, N3798, N3465, N45);
nand NAND4 (N3804, N3787, N409, N2528, N942);
or OR2 (N3805, N3802, N2675);
buf BUF1 (N3806, N3792);
or OR2 (N3807, N3806, N45);
or OR4 (N3808, N3800, N1102, N501, N3593);
nand NAND4 (N3809, N3788, N1151, N1673, N2649);
nor NOR4 (N3810, N3801, N3198, N662, N1582);
nand NAND4 (N3811, N3782, N3645, N2888, N2055);
and AND3 (N3812, N3810, N2571, N2147);
not NOT1 (N3813, N3804);
not NOT1 (N3814, N3807);
xor XOR2 (N3815, N3809, N160);
nor NOR4 (N3816, N3781, N1958, N751, N3395);
nor NOR3 (N3817, N3814, N3428, N1841);
buf BUF1 (N3818, N3816);
or OR4 (N3819, N3811, N1437, N3673, N1546);
and AND3 (N3820, N3818, N1653, N2655);
or OR3 (N3821, N3808, N234, N3392);
and AND3 (N3822, N3817, N1941, N1333);
nor NOR2 (N3823, N3805, N825);
or OR4 (N3824, N3819, N1830, N1654, N1668);
xor XOR2 (N3825, N3815, N1152);
not NOT1 (N3826, N3821);
nor NOR3 (N3827, N3825, N563, N147);
not NOT1 (N3828, N3813);
nand NAND4 (N3829, N3803, N2232, N3466, N194);
and AND3 (N3830, N3823, N1280, N2376);
and AND2 (N3831, N3812, N395);
or OR2 (N3832, N3829, N930);
nor NOR2 (N3833, N3797, N2526);
xor XOR2 (N3834, N3820, N2889);
and AND3 (N3835, N3827, N1212, N2407);
or OR2 (N3836, N3833, N91);
nand NAND2 (N3837, N3826, N691);
xor XOR2 (N3838, N3828, N710);
xor XOR2 (N3839, N3838, N2840);
not NOT1 (N3840, N3822);
or OR2 (N3841, N3831, N1757);
xor XOR2 (N3842, N3839, N2573);
not NOT1 (N3843, N3824);
and AND4 (N3844, N3843, N999, N562, N537);
buf BUF1 (N3845, N3844);
buf BUF1 (N3846, N3842);
nor NOR2 (N3847, N3837, N2157);
xor XOR2 (N3848, N3830, N1370);
nand NAND2 (N3849, N3835, N2066);
nand NAND4 (N3850, N3832, N2406, N3569, N640);
nor NOR2 (N3851, N3836, N3106);
and AND4 (N3852, N3850, N1868, N2212, N824);
or OR2 (N3853, N3834, N3392);
or OR2 (N3854, N3853, N3832);
xor XOR2 (N3855, N3840, N1883);
and AND2 (N3856, N3851, N2121);
buf BUF1 (N3857, N3854);
nand NAND4 (N3858, N3849, N2946, N3659, N3189);
nor NOR3 (N3859, N3847, N972, N1092);
nand NAND2 (N3860, N3858, N2803);
buf BUF1 (N3861, N3852);
buf BUF1 (N3862, N3859);
not NOT1 (N3863, N3861);
and AND2 (N3864, N3863, N1512);
and AND3 (N3865, N3845, N3376, N2819);
or OR4 (N3866, N3841, N3330, N2637, N2796);
xor XOR2 (N3867, N3860, N885);
not NOT1 (N3868, N3848);
nor NOR2 (N3869, N3855, N2090);
nand NAND3 (N3870, N3869, N2203, N2879);
xor XOR2 (N3871, N3862, N2282);
xor XOR2 (N3872, N3866, N430);
or OR4 (N3873, N3872, N1693, N880, N1208);
and AND2 (N3874, N3865, N2772);
xor XOR2 (N3875, N3867, N3380);
xor XOR2 (N3876, N3871, N1238);
xor XOR2 (N3877, N3868, N2611);
and AND2 (N3878, N3856, N3763);
and AND4 (N3879, N3877, N1406, N3838, N269);
nor NOR4 (N3880, N3875, N928, N308, N2463);
xor XOR2 (N3881, N3878, N3452);
and AND2 (N3882, N3876, N1419);
and AND4 (N3883, N3870, N220, N1040, N2240);
xor XOR2 (N3884, N3864, N1612);
nand NAND4 (N3885, N3880, N3028, N3220, N481);
and AND2 (N3886, N3874, N1910);
not NOT1 (N3887, N3881);
xor XOR2 (N3888, N3846, N1759);
xor XOR2 (N3889, N3885, N2520);
nand NAND2 (N3890, N3857, N952);
buf BUF1 (N3891, N3890);
not NOT1 (N3892, N3884);
not NOT1 (N3893, N3879);
xor XOR2 (N3894, N3893, N302);
and AND2 (N3895, N3887, N2519);
nand NAND3 (N3896, N3882, N2759, N934);
nand NAND4 (N3897, N3883, N208, N694, N2523);
buf BUF1 (N3898, N3886);
buf BUF1 (N3899, N3888);
xor XOR2 (N3900, N3899, N122);
nand NAND3 (N3901, N3889, N1420, N935);
nand NAND4 (N3902, N3900, N3292, N3470, N2913);
nor NOR3 (N3903, N3892, N1692, N526);
or OR4 (N3904, N3897, N1381, N789, N3739);
nand NAND2 (N3905, N3896, N1042);
or OR4 (N3906, N3901, N1226, N3612, N244);
nand NAND2 (N3907, N3904, N2357);
xor XOR2 (N3908, N3907, N3103);
buf BUF1 (N3909, N3908);
xor XOR2 (N3910, N3898, N2765);
nor NOR4 (N3911, N3910, N2531, N122, N1320);
nand NAND3 (N3912, N3906, N173, N260);
xor XOR2 (N3913, N3902, N2732);
or OR4 (N3914, N3873, N1303, N2045, N1122);
or OR3 (N3915, N3894, N3461, N704);
xor XOR2 (N3916, N3915, N3325);
and AND2 (N3917, N3903, N3243);
not NOT1 (N3918, N3917);
buf BUF1 (N3919, N3918);
or OR3 (N3920, N3891, N294, N726);
nand NAND4 (N3921, N3895, N2898, N1172, N3705);
xor XOR2 (N3922, N3919, N2648);
xor XOR2 (N3923, N3922, N2988);
not NOT1 (N3924, N3913);
and AND4 (N3925, N3914, N3042, N3025, N509);
or OR2 (N3926, N3912, N3834);
nand NAND3 (N3927, N3916, N3012, N183);
not NOT1 (N3928, N3926);
not NOT1 (N3929, N3920);
nor NOR4 (N3930, N3927, N3639, N1610, N114);
nor NOR2 (N3931, N3911, N485);
xor XOR2 (N3932, N3930, N3046);
nand NAND2 (N3933, N3932, N302);
nand NAND4 (N3934, N3909, N2259, N542, N1611);
nor NOR2 (N3935, N3905, N874);
and AND2 (N3936, N3928, N1813);
buf BUF1 (N3937, N3936);
xor XOR2 (N3938, N3934, N2912);
xor XOR2 (N3939, N3924, N3226);
not NOT1 (N3940, N3935);
xor XOR2 (N3941, N3933, N646);
or OR4 (N3942, N3925, N621, N489, N3801);
xor XOR2 (N3943, N3937, N1481);
or OR3 (N3944, N3938, N3648, N486);
buf BUF1 (N3945, N3940);
or OR4 (N3946, N3921, N200, N515, N1241);
or OR3 (N3947, N3931, N1654, N3143);
not NOT1 (N3948, N3945);
and AND2 (N3949, N3946, N3880);
or OR4 (N3950, N3943, N524, N411, N440);
xor XOR2 (N3951, N3947, N3104);
or OR4 (N3952, N3941, N1312, N492, N2558);
nand NAND2 (N3953, N3952, N2838);
nand NAND4 (N3954, N3953, N873, N1160, N1934);
xor XOR2 (N3955, N3923, N696);
nand NAND4 (N3956, N3942, N2858, N209, N897);
xor XOR2 (N3957, N3956, N3360);
nand NAND3 (N3958, N3948, N3252, N3035);
and AND4 (N3959, N3929, N3059, N2367, N2921);
buf BUF1 (N3960, N3957);
nor NOR4 (N3961, N3939, N2830, N1798, N1102);
or OR2 (N3962, N3961, N2288);
nand NAND4 (N3963, N3951, N925, N1816, N792);
xor XOR2 (N3964, N3944, N2240);
nand NAND3 (N3965, N3950, N1904, N2163);
and AND4 (N3966, N3959, N3918, N3070, N570);
not NOT1 (N3967, N3966);
xor XOR2 (N3968, N3949, N1457);
nand NAND3 (N3969, N3955, N2771, N66);
nand NAND2 (N3970, N3964, N2720);
or OR3 (N3971, N3960, N2516, N1424);
nor NOR3 (N3972, N3963, N2789, N1486);
nor NOR4 (N3973, N3954, N1612, N2262, N3770);
nor NOR2 (N3974, N3969, N808);
xor XOR2 (N3975, N3970, N2811);
buf BUF1 (N3976, N3967);
nand NAND2 (N3977, N3968, N30);
nand NAND3 (N3978, N3958, N2821, N1089);
nor NOR4 (N3979, N3965, N1006, N950, N627);
not NOT1 (N3980, N3974);
not NOT1 (N3981, N3972);
buf BUF1 (N3982, N3975);
nand NAND3 (N3983, N3979, N2939, N242);
and AND4 (N3984, N3971, N1474, N2964, N3234);
nor NOR3 (N3985, N3980, N3871, N1020);
buf BUF1 (N3986, N3962);
nor NOR4 (N3987, N3981, N3631, N1132, N3129);
buf BUF1 (N3988, N3977);
not NOT1 (N3989, N3984);
buf BUF1 (N3990, N3987);
buf BUF1 (N3991, N3982);
and AND3 (N3992, N3988, N2904, N1661);
not NOT1 (N3993, N3973);
nand NAND3 (N3994, N3993, N3371, N634);
and AND3 (N3995, N3990, N1759, N2994);
not NOT1 (N3996, N3976);
and AND2 (N3997, N3985, N3653);
and AND3 (N3998, N3994, N2006, N3698);
or OR4 (N3999, N3996, N3482, N3225, N13);
buf BUF1 (N4000, N3989);
and AND2 (N4001, N4000, N529);
or OR4 (N4002, N3991, N873, N3363, N1214);
and AND2 (N4003, N3978, N1389);
nand NAND4 (N4004, N3997, N3384, N3306, N2623);
not NOT1 (N4005, N3998);
not NOT1 (N4006, N3999);
or OR2 (N4007, N3992, N2175);
nand NAND4 (N4008, N4005, N3946, N1125, N1);
not NOT1 (N4009, N4008);
nor NOR2 (N4010, N3983, N751);
nand NAND4 (N4011, N4003, N3628, N193, N1202);
nand NAND3 (N4012, N4011, N320, N1608);
or OR4 (N4013, N3995, N2682, N1512, N3183);
nor NOR2 (N4014, N4010, N820);
nand NAND3 (N4015, N4001, N3226, N814);
buf BUF1 (N4016, N4007);
and AND2 (N4017, N4015, N1825);
or OR2 (N4018, N4009, N3581);
or OR3 (N4019, N4018, N2129, N3772);
not NOT1 (N4020, N4014);
and AND4 (N4021, N4012, N1291, N2578, N1790);
buf BUF1 (N4022, N4019);
not NOT1 (N4023, N4006);
buf BUF1 (N4024, N4023);
xor XOR2 (N4025, N4017, N2492);
nand NAND2 (N4026, N4002, N1095);
nand NAND3 (N4027, N4022, N3347, N2523);
nand NAND4 (N4028, N4024, N1245, N3708, N1995);
nand NAND2 (N4029, N4020, N3563);
buf BUF1 (N4030, N4027);
buf BUF1 (N4031, N4025);
or OR2 (N4032, N4030, N188);
and AND4 (N4033, N4026, N2851, N265, N2657);
or OR4 (N4034, N4013, N938, N1224, N1636);
and AND4 (N4035, N4033, N2528, N1993, N2711);
and AND2 (N4036, N4016, N2816);
and AND3 (N4037, N3986, N2735, N1960);
not NOT1 (N4038, N4004);
and AND2 (N4039, N4031, N1536);
or OR2 (N4040, N4039, N530);
or OR2 (N4041, N4040, N1553);
not NOT1 (N4042, N4028);
or OR4 (N4043, N4034, N2083, N126, N2452);
and AND3 (N4044, N4036, N1671, N6);
or OR4 (N4045, N4021, N3586, N1790, N233);
or OR4 (N4046, N4037, N2751, N3715, N1299);
and AND4 (N4047, N4041, N3703, N2550, N1234);
buf BUF1 (N4048, N4045);
and AND4 (N4049, N4042, N3181, N679, N2108);
nand NAND3 (N4050, N4047, N1417, N2327);
not NOT1 (N4051, N4035);
buf BUF1 (N4052, N4049);
or OR4 (N4053, N4038, N2367, N1409, N1451);
not NOT1 (N4054, N4050);
or OR4 (N4055, N4043, N2932, N883, N2219);
and AND4 (N4056, N4029, N3387, N3131, N2801);
not NOT1 (N4057, N4048);
or OR3 (N4058, N4054, N68, N1495);
nand NAND3 (N4059, N4052, N1316, N2583);
or OR3 (N4060, N4058, N1074, N3574);
or OR4 (N4061, N4044, N727, N3222, N3109);
nand NAND4 (N4062, N4060, N2878, N217, N145);
nand NAND4 (N4063, N4057, N1598, N1076, N399);
or OR4 (N4064, N4051, N3237, N155, N3575);
and AND4 (N4065, N4032, N117, N3464, N190);
or OR2 (N4066, N4056, N3745);
and AND3 (N4067, N4064, N1321, N1573);
xor XOR2 (N4068, N4062, N2477);
and AND3 (N4069, N4059, N2042, N1225);
nand NAND4 (N4070, N4065, N2345, N2486, N43);
xor XOR2 (N4071, N4069, N441);
buf BUF1 (N4072, N4067);
nor NOR3 (N4073, N4071, N1417, N2813);
nand NAND3 (N4074, N4063, N2029, N2375);
and AND3 (N4075, N4066, N172, N557);
not NOT1 (N4076, N4075);
not NOT1 (N4077, N4046);
nor NOR4 (N4078, N4068, N2764, N1511, N1743);
not NOT1 (N4079, N4077);
nand NAND2 (N4080, N4070, N3312);
xor XOR2 (N4081, N4055, N227);
nand NAND3 (N4082, N4074, N541, N3986);
nand NAND4 (N4083, N4072, N2842, N306, N1558);
nor NOR3 (N4084, N4080, N1149, N412);
nand NAND4 (N4085, N4082, N216, N3519, N2548);
or OR3 (N4086, N4085, N584, N823);
nand NAND3 (N4087, N4084, N980, N3025);
buf BUF1 (N4088, N4087);
xor XOR2 (N4089, N4076, N3270);
and AND2 (N4090, N4061, N3745);
buf BUF1 (N4091, N4088);
not NOT1 (N4092, N4090);
buf BUF1 (N4093, N4053);
or OR2 (N4094, N4089, N922);
nand NAND2 (N4095, N4083, N3948);
nand NAND2 (N4096, N4094, N3967);
nor NOR2 (N4097, N4073, N4054);
buf BUF1 (N4098, N4081);
or OR3 (N4099, N4093, N3848, N2246);
or OR3 (N4100, N4086, N2040, N467);
nor NOR4 (N4101, N4097, N1400, N2434, N3644);
buf BUF1 (N4102, N4095);
nand NAND4 (N4103, N4079, N3412, N1866, N3449);
xor XOR2 (N4104, N4099, N1462);
and AND3 (N4105, N4092, N70, N2527);
and AND3 (N4106, N4100, N1939, N2351);
nand NAND2 (N4107, N4102, N2694);
xor XOR2 (N4108, N4103, N165);
or OR2 (N4109, N4096, N51);
nor NOR3 (N4110, N4091, N3300, N612);
and AND2 (N4111, N4106, N2827);
nand NAND4 (N4112, N4105, N3450, N3507, N1856);
nand NAND4 (N4113, N4104, N1821, N3361, N937);
nand NAND3 (N4114, N4078, N2697, N293);
nand NAND3 (N4115, N4107, N1674, N885);
xor XOR2 (N4116, N4098, N1096);
not NOT1 (N4117, N4111);
not NOT1 (N4118, N4110);
buf BUF1 (N4119, N4118);
nand NAND3 (N4120, N4109, N2835, N3641);
and AND3 (N4121, N4101, N1799, N1671);
buf BUF1 (N4122, N4108);
nand NAND4 (N4123, N4116, N1513, N1696, N2580);
or OR4 (N4124, N4117, N4112, N3144, N3724);
nor NOR2 (N4125, N3511, N4032);
xor XOR2 (N4126, N4115, N1667);
xor XOR2 (N4127, N4124, N3792);
nor NOR3 (N4128, N4126, N2825, N668);
nor NOR2 (N4129, N4113, N3321);
or OR4 (N4130, N4128, N2291, N167, N3943);
not NOT1 (N4131, N4121);
xor XOR2 (N4132, N4123, N594);
and AND4 (N4133, N4129, N2902, N2330, N799);
nand NAND2 (N4134, N4127, N2484);
nand NAND2 (N4135, N4125, N2827);
buf BUF1 (N4136, N4114);
not NOT1 (N4137, N4134);
buf BUF1 (N4138, N4132);
not NOT1 (N4139, N4130);
nor NOR4 (N4140, N4133, N1414, N2360, N958);
or OR2 (N4141, N4135, N3453);
and AND2 (N4142, N4137, N1098);
nand NAND4 (N4143, N4142, N1141, N3566, N3841);
nand NAND3 (N4144, N4131, N1944, N1338);
and AND2 (N4145, N4138, N2136);
xor XOR2 (N4146, N4119, N4064);
nand NAND4 (N4147, N4139, N3770, N3832, N241);
and AND3 (N4148, N4143, N3344, N4129);
nor NOR3 (N4149, N4122, N1686, N139);
not NOT1 (N4150, N4147);
nor NOR2 (N4151, N4149, N272);
or OR4 (N4152, N4150, N1331, N819, N3094);
nor NOR2 (N4153, N4144, N1355);
nor NOR3 (N4154, N4151, N3812, N4056);
buf BUF1 (N4155, N4152);
nand NAND2 (N4156, N4154, N760);
and AND4 (N4157, N4148, N3798, N3287, N1972);
and AND3 (N4158, N4141, N1122, N2385);
nor NOR2 (N4159, N4145, N180);
not NOT1 (N4160, N4140);
or OR3 (N4161, N4159, N1433, N280);
buf BUF1 (N4162, N4158);
nor NOR3 (N4163, N4162, N3931, N1884);
nand NAND2 (N4164, N4155, N245);
nor NOR2 (N4165, N4161, N561);
nor NOR2 (N4166, N4165, N3031);
nor NOR2 (N4167, N4166, N2569);
nand NAND2 (N4168, N4164, N2181);
nand NAND3 (N4169, N4157, N2056, N2126);
xor XOR2 (N4170, N4153, N3587);
nand NAND2 (N4171, N4146, N1907);
nand NAND4 (N4172, N4168, N3425, N369, N609);
xor XOR2 (N4173, N4172, N2935);
nor NOR3 (N4174, N4171, N104, N3386);
and AND4 (N4175, N4169, N4083, N1311, N2547);
nor NOR4 (N4176, N4136, N3873, N536, N3305);
nand NAND4 (N4177, N4160, N977, N1795, N511);
nor NOR4 (N4178, N4174, N1123, N1347, N1054);
nand NAND4 (N4179, N4170, N3999, N2, N3201);
and AND3 (N4180, N4167, N3867, N3605);
not NOT1 (N4181, N4173);
nor NOR4 (N4182, N4179, N1264, N3719, N3763);
nand NAND2 (N4183, N4178, N1070);
nand NAND2 (N4184, N4175, N648);
not NOT1 (N4185, N4180);
nor NOR3 (N4186, N4163, N1721, N2659);
xor XOR2 (N4187, N4156, N1321);
and AND2 (N4188, N4177, N1310);
or OR2 (N4189, N4185, N1186);
nand NAND2 (N4190, N4181, N3945);
or OR4 (N4191, N4183, N3310, N3280, N1308);
nor NOR4 (N4192, N4187, N2638, N349, N937);
nor NOR4 (N4193, N4191, N163, N3336, N3503);
and AND3 (N4194, N4189, N2655, N852);
buf BUF1 (N4195, N4194);
nor NOR3 (N4196, N4188, N2980, N1238);
xor XOR2 (N4197, N4176, N1251);
and AND4 (N4198, N4184, N3359, N2335, N2370);
nor NOR2 (N4199, N4195, N259);
nand NAND3 (N4200, N4190, N1677, N3513);
buf BUF1 (N4201, N4200);
xor XOR2 (N4202, N4120, N2259);
and AND3 (N4203, N4198, N3997, N2150);
or OR2 (N4204, N4203, N3321);
nor NOR2 (N4205, N4182, N2700);
not NOT1 (N4206, N4199);
buf BUF1 (N4207, N4197);
xor XOR2 (N4208, N4207, N1443);
buf BUF1 (N4209, N4202);
nor NOR3 (N4210, N4201, N3932, N892);
not NOT1 (N4211, N4206);
or OR4 (N4212, N4210, N2586, N3384, N801);
and AND2 (N4213, N4196, N3927);
buf BUF1 (N4214, N4186);
nand NAND4 (N4215, N4214, N2634, N1714, N2202);
or OR3 (N4216, N4193, N4077, N3146);
and AND4 (N4217, N4205, N3486, N3383, N1800);
not NOT1 (N4218, N4208);
not NOT1 (N4219, N4209);
nand NAND2 (N4220, N4215, N1218);
xor XOR2 (N4221, N4217, N3285);
nand NAND4 (N4222, N4213, N2911, N1064, N3729);
or OR2 (N4223, N4219, N2626);
xor XOR2 (N4224, N4216, N3697);
nor NOR4 (N4225, N4221, N3749, N1612, N4126);
nand NAND4 (N4226, N4212, N2321, N3371, N977);
xor XOR2 (N4227, N4204, N2880);
xor XOR2 (N4228, N4218, N4105);
or OR2 (N4229, N4223, N3476);
and AND3 (N4230, N4224, N1019, N3170);
nand NAND3 (N4231, N4222, N810, N891);
buf BUF1 (N4232, N4211);
not NOT1 (N4233, N4231);
buf BUF1 (N4234, N4228);
buf BUF1 (N4235, N4232);
xor XOR2 (N4236, N4226, N592);
xor XOR2 (N4237, N4192, N2287);
or OR4 (N4238, N4229, N2824, N1647, N971);
or OR2 (N4239, N4233, N2171);
xor XOR2 (N4240, N4225, N2869);
nor NOR3 (N4241, N4230, N2875, N3625);
buf BUF1 (N4242, N4238);
not NOT1 (N4243, N4234);
and AND2 (N4244, N4227, N964);
nand NAND3 (N4245, N4240, N1298, N359);
nand NAND4 (N4246, N4220, N3630, N3450, N1379);
xor XOR2 (N4247, N4244, N3425);
not NOT1 (N4248, N4243);
nor NOR2 (N4249, N4245, N3818);
nand NAND4 (N4250, N4237, N3349, N964, N20);
not NOT1 (N4251, N4247);
xor XOR2 (N4252, N4239, N469);
and AND3 (N4253, N4246, N644, N159);
nor NOR2 (N4254, N4250, N1963);
and AND3 (N4255, N4236, N2450, N3361);
not NOT1 (N4256, N4253);
not NOT1 (N4257, N4251);
or OR2 (N4258, N4252, N826);
and AND2 (N4259, N4255, N1950);
nand NAND3 (N4260, N4259, N1730, N3974);
xor XOR2 (N4261, N4242, N4239);
nand NAND4 (N4262, N4261, N3780, N1985, N3011);
buf BUF1 (N4263, N4235);
buf BUF1 (N4264, N4258);
not NOT1 (N4265, N4254);
nor NOR2 (N4266, N4241, N438);
not NOT1 (N4267, N4262);
not NOT1 (N4268, N4267);
nor NOR4 (N4269, N4256, N3947, N2496, N3043);
and AND2 (N4270, N4248, N367);
and AND3 (N4271, N4266, N3404, N1124);
or OR4 (N4272, N4249, N3318, N3795, N1741);
xor XOR2 (N4273, N4263, N46);
nand NAND2 (N4274, N4273, N1154);
nand NAND2 (N4275, N4271, N3990);
and AND4 (N4276, N4265, N2679, N3070, N1608);
nand NAND2 (N4277, N4268, N2708);
nor NOR2 (N4278, N4277, N1098);
and AND4 (N4279, N4275, N2853, N2445, N1858);
nand NAND3 (N4280, N4279, N857, N1445);
or OR2 (N4281, N4274, N3224);
or OR2 (N4282, N4278, N1223);
xor XOR2 (N4283, N4282, N3153);
and AND4 (N4284, N4276, N2071, N4265, N3836);
nand NAND2 (N4285, N4257, N954);
and AND2 (N4286, N4285, N778);
and AND2 (N4287, N4280, N2337);
xor XOR2 (N4288, N4287, N2385);
and AND4 (N4289, N4286, N408, N832, N1536);
nand NAND3 (N4290, N4270, N3377, N2029);
not NOT1 (N4291, N4290);
and AND2 (N4292, N4264, N3527);
not NOT1 (N4293, N4284);
nor NOR2 (N4294, N4283, N3056);
xor XOR2 (N4295, N4272, N2961);
nor NOR3 (N4296, N4260, N85, N1090);
xor XOR2 (N4297, N4281, N2822);
nand NAND3 (N4298, N4292, N3573, N504);
and AND4 (N4299, N4269, N4265, N2601, N1325);
xor XOR2 (N4300, N4288, N1394);
and AND2 (N4301, N4300, N4140);
xor XOR2 (N4302, N4293, N3652);
or OR3 (N4303, N4299, N1445, N1584);
not NOT1 (N4304, N4289);
and AND4 (N4305, N4302, N851, N1485, N1721);
or OR2 (N4306, N4297, N1215);
not NOT1 (N4307, N4298);
and AND2 (N4308, N4301, N1907);
nand NAND4 (N4309, N4307, N3051, N576, N2349);
buf BUF1 (N4310, N4295);
and AND4 (N4311, N4306, N1621, N1927, N652);
xor XOR2 (N4312, N4303, N3607);
nor NOR3 (N4313, N4294, N946, N3691);
or OR4 (N4314, N4308, N3463, N3172, N1588);
not NOT1 (N4315, N4311);
buf BUF1 (N4316, N4310);
or OR2 (N4317, N4314, N2936);
or OR2 (N4318, N4309, N4108);
nor NOR2 (N4319, N4296, N2256);
xor XOR2 (N4320, N4319, N1455);
or OR4 (N4321, N4318, N744, N531, N4275);
not NOT1 (N4322, N4317);
xor XOR2 (N4323, N4312, N3531);
nand NAND2 (N4324, N4323, N2671);
nor NOR4 (N4325, N4304, N731, N1271, N2887);
or OR2 (N4326, N4321, N426);
nand NAND2 (N4327, N4322, N3295);
not NOT1 (N4328, N4315);
not NOT1 (N4329, N4320);
nand NAND4 (N4330, N4316, N1137, N708, N1960);
nor NOR2 (N4331, N4327, N2408);
buf BUF1 (N4332, N4329);
xor XOR2 (N4333, N4328, N2612);
not NOT1 (N4334, N4326);
nor NOR4 (N4335, N4291, N3298, N3172, N681);
xor XOR2 (N4336, N4330, N2312);
nand NAND3 (N4337, N4324, N4264, N75);
or OR2 (N4338, N4313, N567);
xor XOR2 (N4339, N4336, N1290);
buf BUF1 (N4340, N4332);
or OR4 (N4341, N4337, N4087, N1917, N3014);
xor XOR2 (N4342, N4340, N4334);
xor XOR2 (N4343, N2143, N198);
or OR2 (N4344, N4342, N3839);
or OR2 (N4345, N4341, N4244);
and AND3 (N4346, N4344, N2196, N3300);
and AND2 (N4347, N4339, N1678);
or OR4 (N4348, N4347, N939, N409, N1380);
and AND4 (N4349, N4335, N4322, N2547, N4125);
and AND2 (N4350, N4333, N1947);
or OR4 (N4351, N4331, N3312, N52, N2973);
or OR2 (N4352, N4338, N97);
or OR4 (N4353, N4349, N2698, N927, N660);
and AND4 (N4354, N4305, N1208, N1873, N891);
not NOT1 (N4355, N4352);
nand NAND2 (N4356, N4353, N540);
buf BUF1 (N4357, N4351);
not NOT1 (N4358, N4348);
not NOT1 (N4359, N4350);
xor XOR2 (N4360, N4343, N1463);
not NOT1 (N4361, N4325);
nor NOR3 (N4362, N4355, N4333, N1271);
and AND4 (N4363, N4362, N2198, N1021, N1656);
not NOT1 (N4364, N4357);
and AND2 (N4365, N4345, N1465);
xor XOR2 (N4366, N4364, N2909);
nor NOR3 (N4367, N4361, N3735, N3331);
and AND4 (N4368, N4360, N2190, N2302, N506);
or OR2 (N4369, N4367, N3988);
nor NOR2 (N4370, N4369, N197);
nand NAND4 (N4371, N4346, N539, N2136, N92);
or OR2 (N4372, N4365, N3380);
buf BUF1 (N4373, N4358);
nand NAND4 (N4374, N4370, N3420, N2587, N3485);
nor NOR4 (N4375, N4368, N3914, N3377, N1535);
or OR2 (N4376, N4372, N1940);
nand NAND2 (N4377, N4371, N1769);
and AND4 (N4378, N4363, N78, N3936, N1349);
not NOT1 (N4379, N4378);
not NOT1 (N4380, N4359);
xor XOR2 (N4381, N4380, N315);
nor NOR3 (N4382, N4374, N4255, N4325);
nor NOR3 (N4383, N4373, N2240, N213);
xor XOR2 (N4384, N4366, N653);
or OR2 (N4385, N4375, N1718);
or OR2 (N4386, N4382, N921);
not NOT1 (N4387, N4376);
xor XOR2 (N4388, N4385, N506);
nand NAND2 (N4389, N4384, N2740);
and AND3 (N4390, N4388, N824, N1226);
nand NAND2 (N4391, N4390, N555);
xor XOR2 (N4392, N4356, N1714);
nand NAND2 (N4393, N4377, N667);
not NOT1 (N4394, N4381);
nor NOR2 (N4395, N4394, N4274);
or OR3 (N4396, N4393, N226, N832);
or OR3 (N4397, N4389, N341, N2244);
xor XOR2 (N4398, N4386, N1643);
xor XOR2 (N4399, N4383, N3500);
not NOT1 (N4400, N4387);
xor XOR2 (N4401, N4398, N726);
or OR3 (N4402, N4400, N3393, N2691);
or OR2 (N4403, N4379, N429);
and AND3 (N4404, N4401, N3684, N2429);
or OR2 (N4405, N4392, N977);
nor NOR2 (N4406, N4395, N779);
nor NOR3 (N4407, N4399, N496, N2951);
nor NOR4 (N4408, N4402, N3004, N168, N1115);
or OR2 (N4409, N4354, N1882);
not NOT1 (N4410, N4404);
not NOT1 (N4411, N4410);
and AND3 (N4412, N4408, N3937, N68);
or OR3 (N4413, N4396, N2715, N2373);
nand NAND2 (N4414, N4413, N393);
buf BUF1 (N4415, N4405);
xor XOR2 (N4416, N4415, N1313);
or OR4 (N4417, N4411, N810, N2110, N2144);
buf BUF1 (N4418, N4397);
and AND4 (N4419, N4407, N1444, N2347, N512);
not NOT1 (N4420, N4417);
nor NOR3 (N4421, N4414, N944, N2049);
nand NAND4 (N4422, N4416, N3293, N42, N2063);
nor NOR4 (N4423, N4412, N31, N1119, N1815);
and AND3 (N4424, N4419, N3918, N904);
not NOT1 (N4425, N4424);
or OR4 (N4426, N4406, N4075, N196, N2901);
xor XOR2 (N4427, N4420, N3667);
xor XOR2 (N4428, N4426, N3665);
and AND2 (N4429, N4422, N948);
buf BUF1 (N4430, N4403);
nor NOR4 (N4431, N4425, N1962, N2122, N4027);
not NOT1 (N4432, N4421);
and AND4 (N4433, N4431, N2121, N763, N3327);
nand NAND2 (N4434, N4429, N370);
or OR3 (N4435, N4432, N237, N125);
nor NOR3 (N4436, N4423, N2153, N4171);
nor NOR4 (N4437, N4428, N658, N4199, N3973);
and AND4 (N4438, N4435, N1579, N4128, N2651);
xor XOR2 (N4439, N4438, N2836);
nor NOR4 (N4440, N4391, N2744, N514, N2825);
not NOT1 (N4441, N4430);
buf BUF1 (N4442, N4441);
xor XOR2 (N4443, N4409, N2998);
and AND4 (N4444, N4443, N1370, N1703, N3437);
xor XOR2 (N4445, N4442, N942);
or OR3 (N4446, N4418, N3516, N1309);
and AND2 (N4447, N4445, N513);
or OR4 (N4448, N4427, N4306, N3692, N280);
not NOT1 (N4449, N4448);
nor NOR3 (N4450, N4447, N435, N1964);
not NOT1 (N4451, N4437);
nand NAND4 (N4452, N4451, N2247, N3481, N3606);
buf BUF1 (N4453, N4434);
nor NOR3 (N4454, N4436, N3372, N1830);
and AND2 (N4455, N4449, N822);
not NOT1 (N4456, N4446);
nor NOR2 (N4457, N4454, N1510);
or OR2 (N4458, N4452, N817);
nand NAND3 (N4459, N4457, N3085, N1572);
not NOT1 (N4460, N4458);
xor XOR2 (N4461, N4460, N4146);
nor NOR2 (N4462, N4461, N2542);
or OR3 (N4463, N4453, N3291, N1028);
nand NAND2 (N4464, N4433, N2779);
xor XOR2 (N4465, N4462, N1924);
not NOT1 (N4466, N4459);
nor NOR2 (N4467, N4450, N2457);
or OR4 (N4468, N4455, N1267, N1587, N3645);
nand NAND4 (N4469, N4465, N3968, N142, N3638);
nand NAND3 (N4470, N4467, N4430, N1114);
buf BUF1 (N4471, N4456);
buf BUF1 (N4472, N4471);
not NOT1 (N4473, N4468);
or OR4 (N4474, N4444, N2321, N2723, N3751);
xor XOR2 (N4475, N4464, N707);
nand NAND4 (N4476, N4473, N3481, N1147, N3567);
or OR2 (N4477, N4463, N2386);
xor XOR2 (N4478, N4474, N778);
xor XOR2 (N4479, N4470, N3086);
not NOT1 (N4480, N4478);
or OR3 (N4481, N4476, N3676, N2788);
and AND2 (N4482, N4440, N1743);
not NOT1 (N4483, N4439);
and AND4 (N4484, N4475, N1386, N4377, N4282);
and AND2 (N4485, N4479, N2122);
not NOT1 (N4486, N4483);
or OR3 (N4487, N4466, N4041, N956);
not NOT1 (N4488, N4480);
not NOT1 (N4489, N4472);
or OR2 (N4490, N4484, N2842);
nor NOR3 (N4491, N4486, N994, N3531);
xor XOR2 (N4492, N4487, N539);
buf BUF1 (N4493, N4489);
nand NAND3 (N4494, N4490, N2037, N700);
or OR4 (N4495, N4494, N1067, N1687, N2907);
buf BUF1 (N4496, N4482);
and AND2 (N4497, N4491, N570);
xor XOR2 (N4498, N4492, N2241);
nand NAND4 (N4499, N4497, N2810, N1025, N375);
nor NOR2 (N4500, N4469, N3275);
or OR4 (N4501, N4481, N2245, N4117, N3052);
xor XOR2 (N4502, N4495, N3397);
nor NOR2 (N4503, N4488, N961);
not NOT1 (N4504, N4493);
or OR2 (N4505, N4496, N1554);
not NOT1 (N4506, N4503);
xor XOR2 (N4507, N4498, N4120);
buf BUF1 (N4508, N4500);
nor NOR2 (N4509, N4508, N2376);
and AND4 (N4510, N4485, N1909, N956, N2854);
not NOT1 (N4511, N4507);
or OR3 (N4512, N4509, N3234, N2535);
and AND4 (N4513, N4511, N4125, N564, N957);
buf BUF1 (N4514, N4501);
nand NAND2 (N4515, N4502, N2293);
nor NOR3 (N4516, N4506, N174, N506);
xor XOR2 (N4517, N4477, N4098);
nand NAND4 (N4518, N4504, N139, N1259, N1592);
nor NOR3 (N4519, N4512, N240, N3826);
nand NAND3 (N4520, N4518, N1884, N433);
or OR3 (N4521, N4516, N4256, N3204);
and AND2 (N4522, N4505, N284);
nand NAND2 (N4523, N4513, N2051);
nor NOR2 (N4524, N4521, N3189);
buf BUF1 (N4525, N4499);
not NOT1 (N4526, N4519);
and AND2 (N4527, N4520, N2920);
and AND3 (N4528, N4526, N1753, N3906);
not NOT1 (N4529, N4523);
nand NAND4 (N4530, N4525, N1903, N4182, N4025);
not NOT1 (N4531, N4514);
nor NOR3 (N4532, N4530, N1327, N161);
or OR3 (N4533, N4522, N1848, N2363);
not NOT1 (N4534, N4517);
buf BUF1 (N4535, N4527);
buf BUF1 (N4536, N4515);
or OR4 (N4537, N4533, N1348, N4066, N2462);
not NOT1 (N4538, N4528);
nor NOR4 (N4539, N4529, N2989, N191, N3549);
or OR2 (N4540, N4524, N803);
nand NAND3 (N4541, N4536, N3142, N256);
not NOT1 (N4542, N4538);
not NOT1 (N4543, N4540);
not NOT1 (N4544, N4542);
and AND2 (N4545, N4544, N2996);
and AND2 (N4546, N4539, N3064);
or OR4 (N4547, N4534, N1564, N2060, N261);
or OR2 (N4548, N4531, N129);
not NOT1 (N4549, N4546);
xor XOR2 (N4550, N4545, N3836);
and AND4 (N4551, N4547, N1604, N2770, N2006);
xor XOR2 (N4552, N4510, N4067);
xor XOR2 (N4553, N4551, N908);
nor NOR3 (N4554, N4537, N1334, N3452);
and AND4 (N4555, N4535, N2655, N3852, N790);
and AND4 (N4556, N4554, N3064, N3049, N3423);
nor NOR2 (N4557, N4553, N2108);
buf BUF1 (N4558, N4543);
xor XOR2 (N4559, N4552, N1059);
xor XOR2 (N4560, N4556, N2252);
nor NOR4 (N4561, N4550, N2261, N3375, N2276);
and AND2 (N4562, N4558, N2486);
not NOT1 (N4563, N4549);
or OR2 (N4564, N4560, N1151);
nand NAND2 (N4565, N4563, N47);
or OR4 (N4566, N4559, N4171, N2976, N1743);
and AND2 (N4567, N4564, N630);
and AND3 (N4568, N4566, N128, N4276);
not NOT1 (N4569, N4548);
and AND4 (N4570, N4557, N525, N4459, N4380);
xor XOR2 (N4571, N4567, N4043);
nor NOR3 (N4572, N4561, N819, N644);
nor NOR2 (N4573, N4555, N747);
and AND4 (N4574, N4573, N3016, N3497, N2187);
not NOT1 (N4575, N4570);
nand NAND3 (N4576, N4541, N4329, N1922);
nor NOR3 (N4577, N4569, N1662, N3133);
xor XOR2 (N4578, N4577, N11);
or OR4 (N4579, N4572, N2667, N3773, N3267);
not NOT1 (N4580, N4578);
nand NAND3 (N4581, N4576, N2119, N632);
nand NAND2 (N4582, N4562, N1435);
xor XOR2 (N4583, N4532, N424);
and AND2 (N4584, N4579, N435);
xor XOR2 (N4585, N4575, N3716);
xor XOR2 (N4586, N4574, N2211);
xor XOR2 (N4587, N4568, N3189);
xor XOR2 (N4588, N4583, N4094);
nand NAND3 (N4589, N4571, N2290, N1945);
not NOT1 (N4590, N4565);
buf BUF1 (N4591, N4587);
or OR4 (N4592, N4589, N232, N4303, N428);
nand NAND2 (N4593, N4584, N111);
and AND4 (N4594, N4593, N1739, N813, N93);
and AND4 (N4595, N4591, N1975, N675, N2064);
and AND3 (N4596, N4585, N4298, N916);
xor XOR2 (N4597, N4590, N1536);
xor XOR2 (N4598, N4596, N1637);
or OR2 (N4599, N4597, N736);
buf BUF1 (N4600, N4592);
or OR4 (N4601, N4600, N290, N2013, N1199);
nor NOR3 (N4602, N4599, N689, N4055);
and AND3 (N4603, N4588, N2229, N4315);
nor NOR4 (N4604, N4586, N3418, N2992, N3221);
and AND2 (N4605, N4601, N3817);
and AND4 (N4606, N4581, N1853, N1897, N1611);
xor XOR2 (N4607, N4602, N3549);
and AND3 (N4608, N4604, N1923, N4118);
nor NOR3 (N4609, N4594, N1850, N3840);
nand NAND4 (N4610, N4603, N1237, N176, N2461);
and AND4 (N4611, N4607, N1204, N3862, N2192);
and AND2 (N4612, N4605, N819);
nand NAND3 (N4613, N4598, N2597, N3231);
xor XOR2 (N4614, N4609, N3201);
not NOT1 (N4615, N4582);
nor NOR2 (N4616, N4611, N1577);
and AND2 (N4617, N4614, N632);
and AND4 (N4618, N4616, N2579, N3136, N3726);
buf BUF1 (N4619, N4608);
and AND3 (N4620, N4606, N2413, N1688);
nor NOR2 (N4621, N4618, N3045);
and AND2 (N4622, N4617, N289);
not NOT1 (N4623, N4612);
nor NOR4 (N4624, N4580, N2324, N4183, N1075);
buf BUF1 (N4625, N4620);
nor NOR3 (N4626, N4622, N2091, N983);
buf BUF1 (N4627, N4621);
nor NOR2 (N4628, N4626, N1422);
xor XOR2 (N4629, N4595, N2921);
not NOT1 (N4630, N4610);
nand NAND4 (N4631, N4630, N1632, N4326, N4247);
nor NOR4 (N4632, N4624, N1104, N1901, N3630);
buf BUF1 (N4633, N4631);
buf BUF1 (N4634, N4619);
nor NOR2 (N4635, N4628, N2054);
not NOT1 (N4636, N4627);
or OR3 (N4637, N4633, N3844, N505);
and AND2 (N4638, N4635, N3201);
nor NOR4 (N4639, N4638, N692, N535, N2665);
or OR4 (N4640, N4623, N91, N687, N453);
not NOT1 (N4641, N4632);
or OR2 (N4642, N4641, N2931);
and AND3 (N4643, N4637, N793, N1505);
nor NOR2 (N4644, N4639, N3802);
or OR3 (N4645, N4625, N1419, N3565);
nor NOR4 (N4646, N4643, N163, N1542, N2017);
nor NOR4 (N4647, N4636, N1140, N1412, N65);
and AND2 (N4648, N4644, N666);
not NOT1 (N4649, N4642);
not NOT1 (N4650, N4634);
xor XOR2 (N4651, N4615, N1126);
nand NAND2 (N4652, N4649, N2282);
buf BUF1 (N4653, N4613);
buf BUF1 (N4654, N4629);
buf BUF1 (N4655, N4650);
xor XOR2 (N4656, N4647, N2474);
xor XOR2 (N4657, N4648, N3231);
xor XOR2 (N4658, N4652, N1268);
not NOT1 (N4659, N4657);
xor XOR2 (N4660, N4653, N1175);
nor NOR2 (N4661, N4659, N1089);
not NOT1 (N4662, N4658);
buf BUF1 (N4663, N4660);
and AND4 (N4664, N4656, N4622, N4540, N739);
xor XOR2 (N4665, N4646, N3443);
not NOT1 (N4666, N4662);
and AND2 (N4667, N4666, N3972);
nand NAND2 (N4668, N4667, N2176);
or OR4 (N4669, N4654, N2568, N878, N4653);
xor XOR2 (N4670, N4663, N2278);
and AND2 (N4671, N4668, N1343);
and AND4 (N4672, N4664, N1035, N267, N2278);
or OR2 (N4673, N4655, N3559);
buf BUF1 (N4674, N4671);
not NOT1 (N4675, N4640);
nor NOR3 (N4676, N4675, N1741, N823);
nand NAND4 (N4677, N4669, N1034, N3912, N4652);
or OR3 (N4678, N4645, N2581, N849);
or OR3 (N4679, N4651, N1503, N3633);
not NOT1 (N4680, N4677);
xor XOR2 (N4681, N4665, N2653);
not NOT1 (N4682, N4679);
not NOT1 (N4683, N4661);
and AND3 (N4684, N4676, N2714, N1002);
not NOT1 (N4685, N4684);
buf BUF1 (N4686, N4678);
and AND4 (N4687, N4670, N1049, N2483, N2278);
buf BUF1 (N4688, N4687);
nor NOR3 (N4689, N4680, N2581, N4438);
or OR4 (N4690, N4674, N3434, N3422, N3327);
and AND4 (N4691, N4673, N1044, N3367, N3815);
xor XOR2 (N4692, N4672, N820);
nor NOR3 (N4693, N4683, N1324, N2908);
or OR4 (N4694, N4681, N898, N3040, N4160);
and AND3 (N4695, N4694, N2354, N2597);
nand NAND2 (N4696, N4685, N2268);
nand NAND2 (N4697, N4686, N4285);
xor XOR2 (N4698, N4697, N4418);
or OR3 (N4699, N4695, N3452, N679);
not NOT1 (N4700, N4682);
nor NOR2 (N4701, N4693, N1369);
or OR4 (N4702, N4699, N1457, N1549, N1039);
buf BUF1 (N4703, N4690);
nor NOR2 (N4704, N4702, N3297);
not NOT1 (N4705, N4701);
not NOT1 (N4706, N4704);
nor NOR2 (N4707, N4705, N3485);
and AND3 (N4708, N4707, N3705, N4247);
or OR4 (N4709, N4703, N4300, N3798, N3493);
xor XOR2 (N4710, N4692, N149);
nand NAND3 (N4711, N4688, N334, N12);
xor XOR2 (N4712, N4696, N1243);
nand NAND2 (N4713, N4698, N3236);
nor NOR2 (N4714, N4706, N4696);
xor XOR2 (N4715, N4708, N4546);
nor NOR4 (N4716, N4709, N1158, N2201, N2134);
or OR3 (N4717, N4714, N3658, N171);
nand NAND2 (N4718, N4700, N1935);
or OR3 (N4719, N4718, N4360, N2022);
xor XOR2 (N4720, N4719, N1614);
nor NOR3 (N4721, N4720, N1488, N3666);
nand NAND2 (N4722, N4716, N2290);
not NOT1 (N4723, N4691);
xor XOR2 (N4724, N4721, N1023);
not NOT1 (N4725, N4724);
buf BUF1 (N4726, N4723);
and AND2 (N4727, N4689, N844);
and AND3 (N4728, N4717, N4317, N4399);
buf BUF1 (N4729, N4726);
buf BUF1 (N4730, N4725);
nand NAND3 (N4731, N4713, N4284, N3421);
nand NAND4 (N4732, N4712, N3406, N312, N4513);
xor XOR2 (N4733, N4711, N3923);
nor NOR4 (N4734, N4728, N3125, N3154, N2485);
xor XOR2 (N4735, N4734, N1455);
xor XOR2 (N4736, N4715, N3899);
not NOT1 (N4737, N4732);
and AND2 (N4738, N4733, N2147);
xor XOR2 (N4739, N4731, N3896);
nor NOR2 (N4740, N4727, N3079);
buf BUF1 (N4741, N4729);
nand NAND2 (N4742, N4710, N454);
nor NOR4 (N4743, N4735, N4112, N1026, N2006);
not NOT1 (N4744, N4722);
and AND3 (N4745, N4742, N3289, N3958);
nand NAND4 (N4746, N4744, N3335, N4646, N2954);
or OR2 (N4747, N4736, N394);
or OR2 (N4748, N4737, N2746);
or OR4 (N4749, N4743, N49, N3215, N1726);
buf BUF1 (N4750, N4747);
nor NOR3 (N4751, N4730, N247, N211);
xor XOR2 (N4752, N4746, N910);
or OR2 (N4753, N4751, N842);
nand NAND4 (N4754, N4738, N4024, N3305, N1086);
or OR3 (N4755, N4752, N1396, N3476);
buf BUF1 (N4756, N4739);
and AND3 (N4757, N4740, N173, N484);
nand NAND2 (N4758, N4741, N4421);
nand NAND2 (N4759, N4754, N239);
xor XOR2 (N4760, N4756, N3809);
nor NOR2 (N4761, N4748, N3771);
not NOT1 (N4762, N4761);
nand NAND4 (N4763, N4749, N473, N3267, N1136);
xor XOR2 (N4764, N4760, N689);
xor XOR2 (N4765, N4764, N2895);
nor NOR3 (N4766, N4753, N3092, N4423);
or OR3 (N4767, N4762, N2011, N3211);
and AND4 (N4768, N4766, N4556, N1118, N1922);
or OR4 (N4769, N4757, N3699, N3760, N2415);
not NOT1 (N4770, N4759);
nor NOR3 (N4771, N4765, N1581, N280);
buf BUF1 (N4772, N4770);
xor XOR2 (N4773, N4745, N133);
and AND2 (N4774, N4771, N4089);
and AND2 (N4775, N4773, N2302);
nand NAND2 (N4776, N4775, N1938);
nand NAND4 (N4777, N4768, N928, N2402, N3284);
buf BUF1 (N4778, N4755);
not NOT1 (N4779, N4769);
buf BUF1 (N4780, N4779);
nor NOR3 (N4781, N4772, N3044, N170);
or OR3 (N4782, N4758, N495, N4255);
nor NOR3 (N4783, N4750, N23, N2268);
or OR4 (N4784, N4774, N3600, N1903, N2553);
or OR3 (N4785, N4767, N4126, N1731);
xor XOR2 (N4786, N4763, N4524);
nand NAND4 (N4787, N4777, N346, N1811, N521);
and AND2 (N4788, N4785, N1414);
not NOT1 (N4789, N4783);
and AND2 (N4790, N4786, N1743);
xor XOR2 (N4791, N4782, N1277);
buf BUF1 (N4792, N4787);
and AND3 (N4793, N4791, N898, N3338);
xor XOR2 (N4794, N4776, N2334);
nor NOR2 (N4795, N4793, N2925);
not NOT1 (N4796, N4778);
and AND2 (N4797, N4792, N30);
or OR2 (N4798, N4796, N4026);
not NOT1 (N4799, N4790);
nand NAND3 (N4800, N4798, N4033, N1541);
nand NAND4 (N4801, N4800, N3844, N1011, N1748);
or OR2 (N4802, N4795, N617);
buf BUF1 (N4803, N4802);
xor XOR2 (N4804, N4781, N1837);
nand NAND4 (N4805, N4803, N3390, N1202, N594);
nand NAND2 (N4806, N4797, N2988);
or OR3 (N4807, N4801, N4357, N1852);
nand NAND2 (N4808, N4799, N1343);
nand NAND2 (N4809, N4807, N3020);
buf BUF1 (N4810, N4808);
and AND3 (N4811, N4810, N411, N2814);
xor XOR2 (N4812, N4805, N2202);
and AND3 (N4813, N4809, N3305, N1296);
not NOT1 (N4814, N4788);
buf BUF1 (N4815, N4789);
and AND3 (N4816, N4812, N4574, N867);
xor XOR2 (N4817, N4794, N341);
xor XOR2 (N4818, N4815, N4042);
nand NAND2 (N4819, N4804, N819);
nand NAND2 (N4820, N4813, N4253);
nand NAND2 (N4821, N4819, N4703);
nand NAND4 (N4822, N4818, N3714, N1510, N1283);
xor XOR2 (N4823, N4806, N3693);
or OR3 (N4824, N4811, N2735, N2933);
and AND2 (N4825, N4823, N63);
nand NAND2 (N4826, N4816, N787);
and AND2 (N4827, N4821, N3371);
and AND2 (N4828, N4827, N1743);
buf BUF1 (N4829, N4828);
and AND2 (N4830, N4826, N747);
nand NAND3 (N4831, N4824, N4233, N73);
not NOT1 (N4832, N4780);
or OR2 (N4833, N4831, N348);
nand NAND2 (N4834, N4830, N2330);
nand NAND3 (N4835, N4825, N2663, N2983);
xor XOR2 (N4836, N4820, N1046);
not NOT1 (N4837, N4832);
nand NAND3 (N4838, N4834, N2010, N2401);
not NOT1 (N4839, N4835);
nand NAND2 (N4840, N4837, N4295);
nand NAND4 (N4841, N4822, N2183, N1383, N3386);
xor XOR2 (N4842, N4839, N2949);
nand NAND3 (N4843, N4814, N3127, N91);
buf BUF1 (N4844, N4784);
buf BUF1 (N4845, N4833);
not NOT1 (N4846, N4844);
xor XOR2 (N4847, N4829, N3698);
nand NAND2 (N4848, N4843, N4160);
nand NAND4 (N4849, N4836, N3141, N1373, N3009);
xor XOR2 (N4850, N4840, N832);
buf BUF1 (N4851, N4849);
buf BUF1 (N4852, N4817);
nand NAND3 (N4853, N4842, N87, N2428);
and AND4 (N4854, N4847, N1803, N715, N871);
or OR2 (N4855, N4853, N1480);
not NOT1 (N4856, N4838);
xor XOR2 (N4857, N4841, N1807);
xor XOR2 (N4858, N4854, N1922);
nor NOR3 (N4859, N4852, N4691, N3270);
buf BUF1 (N4860, N4855);
or OR2 (N4861, N4848, N2835);
xor XOR2 (N4862, N4856, N2453);
and AND4 (N4863, N4859, N931, N4526, N3349);
buf BUF1 (N4864, N4846);
nor NOR2 (N4865, N4851, N1799);
or OR2 (N4866, N4845, N232);
and AND2 (N4867, N4863, N4061);
nor NOR3 (N4868, N4860, N3822, N1574);
nand NAND4 (N4869, N4864, N491, N1211, N1036);
not NOT1 (N4870, N4868);
nand NAND3 (N4871, N4857, N2164, N1993);
nor NOR4 (N4872, N4861, N1635, N207, N3124);
not NOT1 (N4873, N4871);
or OR4 (N4874, N4873, N1703, N2977, N2466);
nor NOR3 (N4875, N4872, N2140, N2328);
not NOT1 (N4876, N4870);
not NOT1 (N4877, N4876);
not NOT1 (N4878, N4866);
xor XOR2 (N4879, N4874, N672);
nand NAND2 (N4880, N4862, N4659);
nand NAND2 (N4881, N4869, N4767);
nand NAND4 (N4882, N4881, N74, N4706, N790);
or OR2 (N4883, N4877, N953);
or OR2 (N4884, N4865, N3501);
not NOT1 (N4885, N4858);
xor XOR2 (N4886, N4878, N4404);
xor XOR2 (N4887, N4875, N2179);
xor XOR2 (N4888, N4850, N2200);
buf BUF1 (N4889, N4885);
nand NAND3 (N4890, N4887, N2174, N2064);
buf BUF1 (N4891, N4883);
xor XOR2 (N4892, N4879, N3650);
nor NOR3 (N4893, N4882, N307, N3536);
not NOT1 (N4894, N4867);
not NOT1 (N4895, N4890);
nand NAND2 (N4896, N4894, N4178);
and AND4 (N4897, N4886, N1314, N3668, N1522);
nor NOR4 (N4898, N4880, N1353, N132, N4132);
xor XOR2 (N4899, N4898, N4701);
and AND4 (N4900, N4892, N1963, N663, N1140);
nand NAND4 (N4901, N4896, N2995, N1350, N4794);
xor XOR2 (N4902, N4900, N867);
xor XOR2 (N4903, N4888, N3468);
buf BUF1 (N4904, N4901);
buf BUF1 (N4905, N4891);
nor NOR4 (N4906, N4893, N2101, N2435, N655);
and AND3 (N4907, N4904, N3363, N3969);
and AND4 (N4908, N4907, N1513, N985, N536);
and AND4 (N4909, N4889, N3859, N1946, N4403);
not NOT1 (N4910, N4905);
nor NOR2 (N4911, N4906, N4752);
nand NAND4 (N4912, N4908, N3384, N2908, N1393);
nor NOR4 (N4913, N4897, N3855, N2273, N2983);
nand NAND2 (N4914, N4902, N1063);
buf BUF1 (N4915, N4909);
nor NOR3 (N4916, N4915, N3291, N2673);
nor NOR3 (N4917, N4916, N2074, N2594);
xor XOR2 (N4918, N4884, N3533);
or OR2 (N4919, N4917, N2782);
buf BUF1 (N4920, N4918);
buf BUF1 (N4921, N4911);
nand NAND4 (N4922, N4895, N3579, N656, N4585);
xor XOR2 (N4923, N4921, N2223);
buf BUF1 (N4924, N4913);
or OR4 (N4925, N4903, N3621, N1503, N4677);
nand NAND4 (N4926, N4910, N3054, N1009, N2012);
buf BUF1 (N4927, N4899);
or OR3 (N4928, N4912, N2303, N3206);
nor NOR3 (N4929, N4919, N4623, N4075);
nor NOR2 (N4930, N4924, N935);
and AND4 (N4931, N4929, N4585, N2319, N2799);
not NOT1 (N4932, N4923);
buf BUF1 (N4933, N4927);
or OR3 (N4934, N4926, N314, N4298);
nor NOR3 (N4935, N4930, N4790, N3027);
xor XOR2 (N4936, N4925, N3697);
and AND4 (N4937, N4932, N4075, N4239, N1556);
xor XOR2 (N4938, N4914, N4795);
xor XOR2 (N4939, N4920, N725);
xor XOR2 (N4940, N4939, N1697);
and AND4 (N4941, N4938, N1026, N534, N4900);
or OR4 (N4942, N4934, N120, N868, N3733);
not NOT1 (N4943, N4936);
xor XOR2 (N4944, N4943, N2792);
nand NAND4 (N4945, N4942, N2637, N1578, N325);
nand NAND3 (N4946, N4928, N196, N4065);
or OR3 (N4947, N4935, N539, N2672);
and AND3 (N4948, N4922, N3423, N4888);
and AND2 (N4949, N4947, N4602);
not NOT1 (N4950, N4945);
not NOT1 (N4951, N4948);
not NOT1 (N4952, N4940);
not NOT1 (N4953, N4946);
and AND3 (N4954, N4953, N2639, N1939);
nand NAND4 (N4955, N4933, N786, N4114, N771);
nor NOR3 (N4956, N4954, N989, N2278);
or OR4 (N4957, N4931, N1025, N96, N1166);
nand NAND4 (N4958, N4950, N2167, N2865, N895);
buf BUF1 (N4959, N4958);
or OR3 (N4960, N4957, N3378, N2705);
and AND4 (N4961, N4949, N1186, N2592, N3172);
nand NAND2 (N4962, N4959, N3405);
not NOT1 (N4963, N4956);
nand NAND4 (N4964, N4952, N4211, N3158, N4321);
and AND4 (N4965, N4962, N743, N4236, N1752);
not NOT1 (N4966, N4941);
or OR3 (N4967, N4966, N3742, N1494);
and AND4 (N4968, N4960, N4845, N1723, N3078);
xor XOR2 (N4969, N4965, N4545);
and AND4 (N4970, N4963, N3923, N358, N306);
not NOT1 (N4971, N4968);
nor NOR3 (N4972, N4964, N4362, N3658);
buf BUF1 (N4973, N4944);
xor XOR2 (N4974, N4967, N827);
nand NAND2 (N4975, N4937, N1498);
nand NAND4 (N4976, N4972, N178, N1699, N1311);
and AND3 (N4977, N4969, N553, N375);
not NOT1 (N4978, N4955);
xor XOR2 (N4979, N4961, N710);
nor NOR3 (N4980, N4971, N1738, N4638);
not NOT1 (N4981, N4978);
nand NAND2 (N4982, N4976, N4353);
or OR3 (N4983, N4974, N1844, N2086);
and AND3 (N4984, N4983, N3942, N4491);
nand NAND2 (N4985, N4982, N3507);
xor XOR2 (N4986, N4975, N636);
xor XOR2 (N4987, N4973, N4521);
or OR3 (N4988, N4984, N2093, N412);
buf BUF1 (N4989, N4970);
or OR3 (N4990, N4986, N4069, N777);
buf BUF1 (N4991, N4990);
and AND4 (N4992, N4981, N2344, N1296, N1943);
or OR4 (N4993, N4985, N3299, N1783, N1534);
xor XOR2 (N4994, N4989, N4634);
and AND3 (N4995, N4979, N3993, N4979);
nor NOR2 (N4996, N4977, N4805);
xor XOR2 (N4997, N4993, N185);
not NOT1 (N4998, N4992);
buf BUF1 (N4999, N4988);
and AND4 (N5000, N4998, N3533, N3809, N1748);
buf BUF1 (N5001, N4980);
not NOT1 (N5002, N4995);
xor XOR2 (N5003, N4996, N4562);
nand NAND4 (N5004, N4991, N1565, N4993, N1107);
nand NAND4 (N5005, N4987, N2069, N4170, N774);
nor NOR4 (N5006, N4994, N1237, N814, N872);
nand NAND4 (N5007, N4997, N1662, N1646, N2038);
xor XOR2 (N5008, N5005, N4138);
or OR4 (N5009, N4999, N3539, N2716, N500);
or OR3 (N5010, N5006, N1956, N931);
nor NOR2 (N5011, N5004, N4302);
buf BUF1 (N5012, N5009);
not NOT1 (N5013, N5002);
xor XOR2 (N5014, N5000, N3302);
and AND2 (N5015, N5012, N939);
xor XOR2 (N5016, N5015, N2379);
buf BUF1 (N5017, N5011);
xor XOR2 (N5018, N5014, N1798);
buf BUF1 (N5019, N5016);
nor NOR4 (N5020, N5013, N2607, N4144, N1631);
nand NAND2 (N5021, N5019, N4486);
nor NOR3 (N5022, N5003, N3249, N3111);
nor NOR3 (N5023, N5020, N2882, N4742);
or OR2 (N5024, N5007, N768);
and AND4 (N5025, N5017, N1569, N4070, N4774);
not NOT1 (N5026, N5023);
buf BUF1 (N5027, N5025);
or OR3 (N5028, N5027, N1808, N2126);
xor XOR2 (N5029, N5028, N79);
buf BUF1 (N5030, N5021);
nor NOR2 (N5031, N5022, N1105);
not NOT1 (N5032, N5031);
xor XOR2 (N5033, N5001, N3872);
or OR2 (N5034, N5026, N2726);
nand NAND4 (N5035, N5024, N1391, N3484, N2522);
nand NAND3 (N5036, N5010, N4847, N2060);
not NOT1 (N5037, N5036);
nand NAND2 (N5038, N5018, N3501);
nand NAND3 (N5039, N4951, N4950, N3602);
nand NAND2 (N5040, N5008, N2046);
and AND3 (N5041, N5032, N1480, N4389);
or OR3 (N5042, N5034, N3060, N1965);
buf BUF1 (N5043, N5038);
buf BUF1 (N5044, N5037);
nand NAND2 (N5045, N5030, N4719);
or OR2 (N5046, N5029, N64);
or OR4 (N5047, N5045, N4034, N3172, N764);
or OR3 (N5048, N5043, N3635, N2190);
nor NOR3 (N5049, N5039, N1581, N4583);
nor NOR4 (N5050, N5042, N2971, N3712, N3548);
xor XOR2 (N5051, N5047, N4789);
nor NOR2 (N5052, N5048, N1339);
and AND2 (N5053, N5052, N40);
xor XOR2 (N5054, N5035, N3544);
or OR2 (N5055, N5053, N645);
nor NOR4 (N5056, N5040, N3479, N4816, N1892);
and AND3 (N5057, N5049, N3063, N2421);
buf BUF1 (N5058, N5041);
and AND3 (N5059, N5055, N2878, N4679);
nand NAND4 (N5060, N5058, N2271, N3262, N1822);
nor NOR4 (N5061, N5044, N4272, N4127, N2360);
buf BUF1 (N5062, N5060);
or OR3 (N5063, N5054, N2468, N3983);
nand NAND2 (N5064, N5061, N3098);
nand NAND4 (N5065, N5051, N1231, N1052, N1207);
not NOT1 (N5066, N5059);
buf BUF1 (N5067, N5065);
not NOT1 (N5068, N5046);
buf BUF1 (N5069, N5062);
xor XOR2 (N5070, N5067, N4);
and AND4 (N5071, N5064, N1515, N1968, N4750);
buf BUF1 (N5072, N5057);
nor NOR4 (N5073, N5063, N4569, N4903, N2991);
nor NOR3 (N5074, N5073, N2022, N2737);
nor NOR2 (N5075, N5068, N4991);
nor NOR2 (N5076, N5069, N905);
buf BUF1 (N5077, N5056);
nor NOR3 (N5078, N5072, N1472, N4595);
not NOT1 (N5079, N5075);
xor XOR2 (N5080, N5078, N1550);
and AND3 (N5081, N5070, N3213, N4673);
not NOT1 (N5082, N5071);
and AND4 (N5083, N5074, N319, N2880, N4951);
and AND3 (N5084, N5066, N4208, N1719);
nor NOR4 (N5085, N5083, N1074, N4534, N1139);
buf BUF1 (N5086, N5084);
not NOT1 (N5087, N5077);
nand NAND4 (N5088, N5079, N2425, N1530, N2144);
or OR3 (N5089, N5076, N2816, N4028);
nand NAND4 (N5090, N5086, N3706, N4007, N4014);
nand NAND3 (N5091, N5033, N2518, N1504);
nand NAND2 (N5092, N5087, N922);
buf BUF1 (N5093, N5085);
and AND2 (N5094, N5088, N4064);
xor XOR2 (N5095, N5082, N4108);
buf BUF1 (N5096, N5081);
buf BUF1 (N5097, N5090);
buf BUF1 (N5098, N5089);
or OR3 (N5099, N5095, N362, N1974);
nor NOR4 (N5100, N5092, N4393, N4997, N2086);
buf BUF1 (N5101, N5096);
or OR3 (N5102, N5100, N2035, N2872);
and AND4 (N5103, N5097, N1945, N1306, N1079);
nor NOR4 (N5104, N5080, N4307, N69, N952);
xor XOR2 (N5105, N5098, N4346);
or OR2 (N5106, N5101, N511);
and AND3 (N5107, N5050, N292, N3815);
and AND2 (N5108, N5103, N1712);
xor XOR2 (N5109, N5107, N447);
and AND4 (N5110, N5104, N3667, N2804, N1405);
xor XOR2 (N5111, N5099, N4336);
nor NOR2 (N5112, N5093, N1386);
nor NOR3 (N5113, N5102, N582, N3548);
xor XOR2 (N5114, N5105, N3345);
and AND4 (N5115, N5110, N1692, N75, N82);
nand NAND3 (N5116, N5091, N3492, N3376);
and AND3 (N5117, N5112, N3751, N4822);
not NOT1 (N5118, N5106);
buf BUF1 (N5119, N5113);
not NOT1 (N5120, N5111);
or OR4 (N5121, N5117, N2741, N2465, N1450);
or OR4 (N5122, N5121, N2564, N3829, N2524);
nor NOR4 (N5123, N5114, N1235, N4981, N3301);
and AND2 (N5124, N5094, N3411);
and AND3 (N5125, N5119, N2865, N865);
xor XOR2 (N5126, N5123, N1285);
buf BUF1 (N5127, N5124);
nor NOR4 (N5128, N5116, N4832, N3928, N4443);
not NOT1 (N5129, N5125);
nor NOR3 (N5130, N5127, N1743, N2093);
not NOT1 (N5131, N5118);
and AND3 (N5132, N5126, N1350, N4796);
or OR4 (N5133, N5128, N2011, N305, N3427);
buf BUF1 (N5134, N5108);
nor NOR2 (N5135, N5115, N1900);
and AND4 (N5136, N5129, N2519, N3771, N56);
nand NAND3 (N5137, N5136, N2170, N791);
not NOT1 (N5138, N5131);
buf BUF1 (N5139, N5130);
not NOT1 (N5140, N5137);
and AND4 (N5141, N5139, N3005, N1083, N2035);
and AND2 (N5142, N5120, N421);
xor XOR2 (N5143, N5138, N1105);
and AND3 (N5144, N5133, N4449, N1819);
not NOT1 (N5145, N5134);
buf BUF1 (N5146, N5132);
and AND2 (N5147, N5122, N4601);
nor NOR2 (N5148, N5146, N2817);
not NOT1 (N5149, N5143);
xor XOR2 (N5150, N5142, N2812);
xor XOR2 (N5151, N5150, N116);
nor NOR3 (N5152, N5147, N240, N3127);
not NOT1 (N5153, N5141);
buf BUF1 (N5154, N5135);
buf BUF1 (N5155, N5152);
nand NAND2 (N5156, N5145, N998);
or OR4 (N5157, N5156, N1947, N460, N2855);
nor NOR3 (N5158, N5157, N131, N1096);
xor XOR2 (N5159, N5154, N4209);
nand NAND3 (N5160, N5153, N588, N4558);
or OR2 (N5161, N5109, N549);
buf BUF1 (N5162, N5148);
or OR3 (N5163, N5144, N4262, N1628);
xor XOR2 (N5164, N5158, N1623);
xor XOR2 (N5165, N5140, N1268);
xor XOR2 (N5166, N5161, N61);
nand NAND2 (N5167, N5155, N4110);
or OR2 (N5168, N5162, N1524);
nand NAND4 (N5169, N5167, N357, N509, N4230);
xor XOR2 (N5170, N5166, N230);
buf BUF1 (N5171, N5168);
buf BUF1 (N5172, N5160);
or OR2 (N5173, N5170, N3309);
and AND2 (N5174, N5172, N3710);
and AND2 (N5175, N5171, N5061);
buf BUF1 (N5176, N5149);
nor NOR3 (N5177, N5173, N2203, N3557);
xor XOR2 (N5178, N5175, N3496);
buf BUF1 (N5179, N5174);
xor XOR2 (N5180, N5178, N1138);
or OR2 (N5181, N5151, N3087);
xor XOR2 (N5182, N5159, N4870);
xor XOR2 (N5183, N5165, N1662);
buf BUF1 (N5184, N5163);
nor NOR3 (N5185, N5164, N882, N1257);
nand NAND3 (N5186, N5184, N333, N4484);
xor XOR2 (N5187, N5176, N4190);
nor NOR4 (N5188, N5182, N2906, N3787, N622);
nand NAND3 (N5189, N5183, N513, N1029);
nand NAND3 (N5190, N5187, N5124, N3043);
buf BUF1 (N5191, N5185);
nor NOR4 (N5192, N5169, N3659, N1426, N3677);
and AND2 (N5193, N5177, N4216);
xor XOR2 (N5194, N5186, N4313);
nor NOR3 (N5195, N5181, N973, N759);
nor NOR3 (N5196, N5192, N2473, N736);
buf BUF1 (N5197, N5180);
and AND2 (N5198, N5197, N4747);
nand NAND4 (N5199, N5191, N2899, N390, N172);
and AND4 (N5200, N5188, N2712, N2814, N4659);
and AND3 (N5201, N5195, N1330, N3274);
buf BUF1 (N5202, N5196);
xor XOR2 (N5203, N5200, N4714);
nand NAND3 (N5204, N5193, N4095, N3811);
not NOT1 (N5205, N5202);
and AND4 (N5206, N5190, N3798, N326, N3916);
or OR3 (N5207, N5204, N2273, N4745);
and AND4 (N5208, N5205, N409, N1777, N4499);
or OR3 (N5209, N5179, N1579, N3823);
not NOT1 (N5210, N5198);
and AND2 (N5211, N5210, N4255);
and AND2 (N5212, N5203, N303);
nand NAND2 (N5213, N5199, N3563);
nand NAND4 (N5214, N5201, N3091, N2363, N3150);
not NOT1 (N5215, N5212);
xor XOR2 (N5216, N5206, N4295);
xor XOR2 (N5217, N5211, N494);
nand NAND2 (N5218, N5213, N2030);
and AND2 (N5219, N5189, N4370);
nand NAND4 (N5220, N5215, N2985, N209, N2897);
xor XOR2 (N5221, N5219, N1208);
nand NAND2 (N5222, N5216, N1911);
nand NAND2 (N5223, N5222, N249);
not NOT1 (N5224, N5214);
xor XOR2 (N5225, N5223, N20);
or OR2 (N5226, N5218, N3609);
not NOT1 (N5227, N5217);
nand NAND3 (N5228, N5207, N305, N3627);
nand NAND4 (N5229, N5228, N4513, N1463, N960);
or OR4 (N5230, N5221, N5146, N111, N1247);
xor XOR2 (N5231, N5226, N276);
not NOT1 (N5232, N5209);
not NOT1 (N5233, N5194);
nor NOR3 (N5234, N5224, N2976, N209);
nand NAND2 (N5235, N5220, N2015);
xor XOR2 (N5236, N5225, N4936);
or OR4 (N5237, N5234, N4255, N365, N5141);
and AND3 (N5238, N5231, N4291, N591);
buf BUF1 (N5239, N5227);
and AND2 (N5240, N5233, N1187);
nand NAND2 (N5241, N5238, N4654);
not NOT1 (N5242, N5241);
not NOT1 (N5243, N5230);
or OR4 (N5244, N5229, N4877, N1517, N4573);
nor NOR3 (N5245, N5243, N1743, N3448);
and AND4 (N5246, N5244, N3379, N1180, N4106);
xor XOR2 (N5247, N5239, N2262);
xor XOR2 (N5248, N5242, N4301);
xor XOR2 (N5249, N5246, N2512);
not NOT1 (N5250, N5208);
or OR4 (N5251, N5235, N1315, N3001, N76);
not NOT1 (N5252, N5236);
buf BUF1 (N5253, N5250);
and AND3 (N5254, N5237, N3582, N4298);
and AND4 (N5255, N5251, N1905, N4979, N1954);
or OR3 (N5256, N5253, N424, N2768);
nor NOR3 (N5257, N5240, N4370, N2774);
or OR3 (N5258, N5249, N950, N4081);
xor XOR2 (N5259, N5255, N4922);
nand NAND4 (N5260, N5257, N5068, N4756, N352);
and AND2 (N5261, N5252, N2565);
nand NAND4 (N5262, N5259, N1760, N562, N1481);
nand NAND3 (N5263, N5258, N4907, N768);
nor NOR2 (N5264, N5262, N1326);
nand NAND3 (N5265, N5256, N1488, N1450);
buf BUF1 (N5266, N5263);
or OR4 (N5267, N5264, N4664, N2243, N3314);
not NOT1 (N5268, N5232);
not NOT1 (N5269, N5254);
xor XOR2 (N5270, N5260, N1968);
nor NOR4 (N5271, N5247, N2751, N2070, N2644);
nor NOR4 (N5272, N5265, N2720, N5057, N717);
not NOT1 (N5273, N5266);
buf BUF1 (N5274, N5273);
not NOT1 (N5275, N5248);
and AND2 (N5276, N5261, N941);
buf BUF1 (N5277, N5276);
nand NAND4 (N5278, N5275, N179, N2743, N1381);
buf BUF1 (N5279, N5272);
and AND2 (N5280, N5277, N1906);
or OR2 (N5281, N5279, N1110);
not NOT1 (N5282, N5271);
xor XOR2 (N5283, N5268, N3425);
xor XOR2 (N5284, N5281, N253);
not NOT1 (N5285, N5278);
nand NAND3 (N5286, N5282, N1978, N2896);
not NOT1 (N5287, N5245);
nor NOR3 (N5288, N5280, N1147, N1869);
or OR4 (N5289, N5284, N1313, N293, N460);
not NOT1 (N5290, N5289);
or OR4 (N5291, N5287, N2941, N143, N3985);
not NOT1 (N5292, N5270);
nand NAND2 (N5293, N5285, N764);
or OR4 (N5294, N5291, N4561, N4145, N3178);
or OR4 (N5295, N5292, N2330, N3349, N2831);
buf BUF1 (N5296, N5267);
or OR2 (N5297, N5290, N463);
buf BUF1 (N5298, N5297);
not NOT1 (N5299, N5296);
not NOT1 (N5300, N5298);
or OR2 (N5301, N5295, N2014);
xor XOR2 (N5302, N5274, N4711);
xor XOR2 (N5303, N5299, N4337);
not NOT1 (N5304, N5294);
or OR4 (N5305, N5303, N4340, N4649, N1139);
and AND2 (N5306, N5283, N318);
nor NOR2 (N5307, N5302, N3205);
nor NOR4 (N5308, N5304, N2424, N944, N4955);
nand NAND2 (N5309, N5269, N1079);
xor XOR2 (N5310, N5309, N567);
buf BUF1 (N5311, N5308);
and AND2 (N5312, N5305, N4400);
nand NAND3 (N5313, N5311, N2387, N2330);
nor NOR2 (N5314, N5286, N4940);
buf BUF1 (N5315, N5307);
not NOT1 (N5316, N5310);
not NOT1 (N5317, N5306);
not NOT1 (N5318, N5314);
buf BUF1 (N5319, N5301);
and AND2 (N5320, N5319, N2589);
nor NOR2 (N5321, N5313, N2662);
nand NAND2 (N5322, N5317, N221);
nor NOR4 (N5323, N5300, N3213, N2817, N2927);
not NOT1 (N5324, N5321);
nand NAND4 (N5325, N5320, N4627, N3793, N4330);
buf BUF1 (N5326, N5293);
nand NAND3 (N5327, N5288, N4221, N2005);
not NOT1 (N5328, N5312);
nor NOR2 (N5329, N5325, N1679);
or OR3 (N5330, N5323, N2285, N1215);
buf BUF1 (N5331, N5322);
or OR4 (N5332, N5316, N4331, N610, N5123);
xor XOR2 (N5333, N5318, N379);
or OR3 (N5334, N5326, N5270, N3262);
and AND4 (N5335, N5327, N4702, N4153, N3058);
buf BUF1 (N5336, N5330);
not NOT1 (N5337, N5332);
not NOT1 (N5338, N5329);
buf BUF1 (N5339, N5333);
or OR2 (N5340, N5338, N1066);
and AND3 (N5341, N5328, N1311, N5033);
nor NOR3 (N5342, N5331, N470, N2457);
and AND2 (N5343, N5340, N1957);
xor XOR2 (N5344, N5341, N3793);
nor NOR2 (N5345, N5337, N4784);
or OR2 (N5346, N5342, N2842);
xor XOR2 (N5347, N5334, N4697);
or OR2 (N5348, N5324, N3401);
xor XOR2 (N5349, N5347, N2351);
xor XOR2 (N5350, N5345, N3899);
xor XOR2 (N5351, N5343, N3416);
not NOT1 (N5352, N5348);
not NOT1 (N5353, N5335);
and AND4 (N5354, N5346, N4352, N2033, N182);
or OR2 (N5355, N5336, N2271);
and AND4 (N5356, N5351, N1406, N5104, N1449);
not NOT1 (N5357, N5349);
or OR3 (N5358, N5352, N226, N3675);
buf BUF1 (N5359, N5355);
buf BUF1 (N5360, N5354);
buf BUF1 (N5361, N5353);
and AND4 (N5362, N5350, N4622, N3396, N5294);
nand NAND3 (N5363, N5361, N2243, N3206);
nor NOR3 (N5364, N5339, N303, N4401);
buf BUF1 (N5365, N5359);
and AND4 (N5366, N5360, N4931, N4384, N403);
not NOT1 (N5367, N5362);
buf BUF1 (N5368, N5366);
not NOT1 (N5369, N5315);
nor NOR3 (N5370, N5344, N1970, N4165);
or OR2 (N5371, N5368, N1431);
or OR2 (N5372, N5371, N1808);
and AND3 (N5373, N5364, N1916, N274);
xor XOR2 (N5374, N5370, N1);
and AND2 (N5375, N5367, N2152);
and AND4 (N5376, N5358, N4198, N5205, N2664);
buf BUF1 (N5377, N5376);
not NOT1 (N5378, N5373);
nand NAND4 (N5379, N5357, N4350, N3423, N2213);
buf BUF1 (N5380, N5365);
not NOT1 (N5381, N5372);
nor NOR2 (N5382, N5377, N1565);
nand NAND2 (N5383, N5381, N2641);
nand NAND2 (N5384, N5369, N54);
xor XOR2 (N5385, N5379, N4129);
or OR2 (N5386, N5356, N4783);
nand NAND4 (N5387, N5375, N357, N1097, N2234);
buf BUF1 (N5388, N5380);
or OR3 (N5389, N5386, N4915, N2393);
and AND4 (N5390, N5378, N1129, N2557, N2919);
not NOT1 (N5391, N5363);
buf BUF1 (N5392, N5384);
and AND3 (N5393, N5392, N4643, N1248);
xor XOR2 (N5394, N5391, N1889);
or OR4 (N5395, N5385, N138, N3025, N1004);
or OR2 (N5396, N5393, N3931);
or OR2 (N5397, N5389, N3107);
and AND3 (N5398, N5395, N3297, N1527);
nor NOR2 (N5399, N5398, N2442);
xor XOR2 (N5400, N5383, N2032);
not NOT1 (N5401, N5400);
and AND2 (N5402, N5397, N4891);
and AND2 (N5403, N5382, N1830);
or OR4 (N5404, N5399, N3959, N1751, N4427);
xor XOR2 (N5405, N5403, N2067);
nand NAND4 (N5406, N5374, N1884, N5266, N900);
nor NOR3 (N5407, N5390, N5356, N2160);
not NOT1 (N5408, N5406);
or OR2 (N5409, N5396, N2453);
nand NAND4 (N5410, N5408, N648, N661, N2457);
buf BUF1 (N5411, N5405);
not NOT1 (N5412, N5407);
buf BUF1 (N5413, N5402);
nor NOR4 (N5414, N5394, N3232, N2063, N2923);
nand NAND2 (N5415, N5413, N5386);
xor XOR2 (N5416, N5414, N2603);
not NOT1 (N5417, N5412);
buf BUF1 (N5418, N5417);
nor NOR2 (N5419, N5415, N3233);
or OR3 (N5420, N5416, N1399, N4104);
and AND2 (N5421, N5409, N4916);
or OR3 (N5422, N5411, N1841, N452);
nand NAND4 (N5423, N5421, N3942, N3599, N937);
nor NOR4 (N5424, N5418, N1389, N3920, N18);
not NOT1 (N5425, N5387);
nand NAND3 (N5426, N5422, N5204, N2556);
xor XOR2 (N5427, N5425, N2053);
nand NAND3 (N5428, N5404, N4851, N682);
or OR4 (N5429, N5410, N1632, N2089, N5019);
buf BUF1 (N5430, N5420);
not NOT1 (N5431, N5401);
buf BUF1 (N5432, N5419);
and AND2 (N5433, N5431, N4187);
nand NAND2 (N5434, N5423, N2142);
and AND3 (N5435, N5432, N4858, N503);
nand NAND3 (N5436, N5427, N1454, N3728);
and AND4 (N5437, N5433, N3469, N4910, N2110);
not NOT1 (N5438, N5434);
buf BUF1 (N5439, N5428);
xor XOR2 (N5440, N5438, N1464);
or OR4 (N5441, N5430, N1167, N874, N1081);
and AND2 (N5442, N5436, N5304);
nor NOR2 (N5443, N5437, N1078);
nor NOR4 (N5444, N5429, N4229, N3969, N1119);
xor XOR2 (N5445, N5444, N3496);
and AND2 (N5446, N5443, N3648);
nand NAND2 (N5447, N5426, N100);
and AND3 (N5448, N5441, N5059, N532);
nand NAND2 (N5449, N5442, N2060);
not NOT1 (N5450, N5446);
not NOT1 (N5451, N5447);
nor NOR2 (N5452, N5450, N2755);
and AND3 (N5453, N5448, N3974, N3403);
nor NOR4 (N5454, N5451, N3088, N389, N865);
buf BUF1 (N5455, N5449);
and AND4 (N5456, N5445, N5382, N5297, N2787);
not NOT1 (N5457, N5439);
and AND3 (N5458, N5440, N2876, N1529);
or OR4 (N5459, N5457, N5345, N1824, N1382);
nor NOR2 (N5460, N5458, N5459);
nand NAND3 (N5461, N5327, N2957, N3055);
or OR3 (N5462, N5435, N371, N5380);
buf BUF1 (N5463, N5453);
not NOT1 (N5464, N5456);
buf BUF1 (N5465, N5464);
and AND2 (N5466, N5462, N2250);
nor NOR3 (N5467, N5455, N3949, N4069);
xor XOR2 (N5468, N5452, N835);
buf BUF1 (N5469, N5388);
xor XOR2 (N5470, N5469, N2098);
or OR2 (N5471, N5470, N762);
nor NOR2 (N5472, N5461, N2013);
buf BUF1 (N5473, N5467);
not NOT1 (N5474, N5466);
nand NAND4 (N5475, N5473, N703, N3066, N4297);
buf BUF1 (N5476, N5460);
and AND2 (N5477, N5475, N209);
and AND2 (N5478, N5472, N2560);
nor NOR4 (N5479, N5465, N3958, N2512, N4767);
nor NOR3 (N5480, N5424, N4482, N1496);
xor XOR2 (N5481, N5468, N576);
xor XOR2 (N5482, N5480, N4491);
nor NOR2 (N5483, N5463, N4896);
xor XOR2 (N5484, N5481, N2657);
and AND3 (N5485, N5479, N2379, N638);
nor NOR3 (N5486, N5484, N4466, N1899);
not NOT1 (N5487, N5482);
xor XOR2 (N5488, N5485, N3700);
buf BUF1 (N5489, N5476);
nand NAND4 (N5490, N5478, N1268, N1670, N3232);
nand NAND3 (N5491, N5474, N4900, N746);
xor XOR2 (N5492, N5483, N443);
buf BUF1 (N5493, N5471);
nand NAND3 (N5494, N5477, N2103, N3520);
nand NAND4 (N5495, N5492, N5070, N3022, N5474);
not NOT1 (N5496, N5490);
nand NAND3 (N5497, N5495, N1370, N3178);
nor NOR2 (N5498, N5488, N239);
or OR2 (N5499, N5493, N4487);
nand NAND3 (N5500, N5499, N627, N1333);
not NOT1 (N5501, N5500);
xor XOR2 (N5502, N5497, N5270);
or OR2 (N5503, N5498, N1263);
nand NAND2 (N5504, N5489, N5104);
or OR4 (N5505, N5503, N1131, N4366, N2336);
buf BUF1 (N5506, N5494);
nand NAND4 (N5507, N5454, N3009, N155, N2605);
nand NAND2 (N5508, N5486, N337);
nand NAND2 (N5509, N5502, N4683);
buf BUF1 (N5510, N5508);
buf BUF1 (N5511, N5509);
or OR4 (N5512, N5510, N5319, N5030, N121);
not NOT1 (N5513, N5487);
buf BUF1 (N5514, N5505);
not NOT1 (N5515, N5513);
nor NOR2 (N5516, N5515, N1042);
not NOT1 (N5517, N5506);
or OR3 (N5518, N5511, N3718, N109);
and AND4 (N5519, N5517, N3464, N3470, N583);
and AND4 (N5520, N5518, N1003, N80, N5412);
or OR4 (N5521, N5514, N4703, N503, N517);
not NOT1 (N5522, N5501);
nand NAND2 (N5523, N5521, N1160);
xor XOR2 (N5524, N5523, N3403);
nor NOR2 (N5525, N5496, N3029);
buf BUF1 (N5526, N5519);
xor XOR2 (N5527, N5504, N1932);
buf BUF1 (N5528, N5525);
xor XOR2 (N5529, N5528, N1462);
or OR3 (N5530, N5491, N4612, N332);
and AND2 (N5531, N5522, N1634);
and AND2 (N5532, N5524, N3609);
nor NOR3 (N5533, N5516, N201, N673);
buf BUF1 (N5534, N5507);
buf BUF1 (N5535, N5529);
xor XOR2 (N5536, N5532, N4474);
not NOT1 (N5537, N5534);
buf BUF1 (N5538, N5520);
xor XOR2 (N5539, N5527, N2070);
xor XOR2 (N5540, N5512, N3413);
nand NAND2 (N5541, N5533, N3522);
xor XOR2 (N5542, N5526, N1184);
xor XOR2 (N5543, N5536, N1927);
nor NOR2 (N5544, N5531, N2547);
xor XOR2 (N5545, N5539, N1645);
not NOT1 (N5546, N5538);
nor NOR3 (N5547, N5546, N3798, N4193);
xor XOR2 (N5548, N5537, N1315);
xor XOR2 (N5549, N5548, N3351);
xor XOR2 (N5550, N5530, N76);
nor NOR3 (N5551, N5549, N3905, N1649);
and AND3 (N5552, N5542, N5434, N3678);
xor XOR2 (N5553, N5550, N5020);
xor XOR2 (N5554, N5545, N4923);
not NOT1 (N5555, N5541);
buf BUF1 (N5556, N5555);
nor NOR2 (N5557, N5552, N3896);
not NOT1 (N5558, N5551);
nand NAND2 (N5559, N5556, N2641);
xor XOR2 (N5560, N5554, N1338);
nor NOR2 (N5561, N5535, N5428);
or OR4 (N5562, N5558, N2208, N1360, N3677);
xor XOR2 (N5563, N5547, N5488);
nor NOR4 (N5564, N5561, N276, N5312, N4517);
buf BUF1 (N5565, N5559);
and AND2 (N5566, N5544, N3375);
nor NOR2 (N5567, N5543, N4006);
nor NOR3 (N5568, N5566, N709, N447);
and AND2 (N5569, N5565, N1345);
nand NAND4 (N5570, N5560, N2235, N5354, N2115);
not NOT1 (N5571, N5569);
nor NOR4 (N5572, N5557, N4527, N5331, N4141);
buf BUF1 (N5573, N5568);
nand NAND3 (N5574, N5563, N3991, N1800);
not NOT1 (N5575, N5572);
and AND4 (N5576, N5570, N4107, N1910, N3941);
and AND2 (N5577, N5540, N3060);
xor XOR2 (N5578, N5573, N2626);
nand NAND3 (N5579, N5576, N1712, N3125);
buf BUF1 (N5580, N5575);
xor XOR2 (N5581, N5577, N2807);
nand NAND4 (N5582, N5580, N1509, N2754, N2399);
nor NOR2 (N5583, N5567, N3950);
nor NOR4 (N5584, N5579, N4630, N3490, N3155);
xor XOR2 (N5585, N5584, N2292);
nor NOR3 (N5586, N5581, N2543, N3883);
xor XOR2 (N5587, N5562, N644);
or OR2 (N5588, N5586, N1724);
not NOT1 (N5589, N5587);
nand NAND2 (N5590, N5564, N3413);
nand NAND2 (N5591, N5553, N2946);
and AND3 (N5592, N5578, N4977, N3946);
nor NOR2 (N5593, N5571, N5183);
buf BUF1 (N5594, N5589);
nand NAND3 (N5595, N5583, N2565, N3426);
buf BUF1 (N5596, N5582);
xor XOR2 (N5597, N5595, N4401);
not NOT1 (N5598, N5590);
nand NAND2 (N5599, N5591, N990);
nand NAND3 (N5600, N5599, N1183, N687);
or OR3 (N5601, N5588, N1979, N404);
not NOT1 (N5602, N5598);
or OR2 (N5603, N5593, N3993);
buf BUF1 (N5604, N5594);
nor NOR2 (N5605, N5604, N3234);
buf BUF1 (N5606, N5605);
nand NAND4 (N5607, N5606, N1588, N345, N2032);
nand NAND4 (N5608, N5596, N4261, N635, N246);
or OR3 (N5609, N5603, N2229, N535);
xor XOR2 (N5610, N5585, N3334);
buf BUF1 (N5611, N5608);
nor NOR2 (N5612, N5600, N739);
xor XOR2 (N5613, N5601, N4037);
nand NAND3 (N5614, N5607, N234, N256);
xor XOR2 (N5615, N5611, N1462);
xor XOR2 (N5616, N5609, N4860);
or OR4 (N5617, N5613, N1116, N3507, N3736);
buf BUF1 (N5618, N5597);
nor NOR3 (N5619, N5618, N1436, N3448);
or OR3 (N5620, N5612, N3958, N5225);
or OR3 (N5621, N5574, N116, N4037);
and AND3 (N5622, N5620, N406, N2529);
not NOT1 (N5623, N5602);
or OR2 (N5624, N5621, N776);
nand NAND2 (N5625, N5610, N4782);
or OR2 (N5626, N5592, N1183);
not NOT1 (N5627, N5622);
and AND4 (N5628, N5614, N5133, N2105, N5433);
nor NOR2 (N5629, N5627, N5281);
xor XOR2 (N5630, N5616, N5175);
and AND2 (N5631, N5617, N5159);
buf BUF1 (N5632, N5631);
nand NAND4 (N5633, N5632, N4759, N5614, N5237);
nor NOR3 (N5634, N5615, N5456, N4994);
not NOT1 (N5635, N5623);
nand NAND2 (N5636, N5634, N1206);
nand NAND2 (N5637, N5629, N1966);
nor NOR3 (N5638, N5626, N4112, N1821);
or OR4 (N5639, N5637, N473, N2832, N1372);
or OR3 (N5640, N5636, N3504, N1077);
nor NOR2 (N5641, N5628, N3570);
or OR2 (N5642, N5639, N2102);
buf BUF1 (N5643, N5633);
not NOT1 (N5644, N5643);
not NOT1 (N5645, N5625);
buf BUF1 (N5646, N5624);
buf BUF1 (N5647, N5646);
nand NAND2 (N5648, N5647, N1409);
not NOT1 (N5649, N5619);
or OR2 (N5650, N5644, N2279);
and AND4 (N5651, N5641, N772, N3803, N680);
and AND2 (N5652, N5635, N1665);
nand NAND2 (N5653, N5638, N4447);
or OR4 (N5654, N5648, N5141, N1735, N3999);
xor XOR2 (N5655, N5640, N4700);
nor NOR4 (N5656, N5650, N1581, N405, N2708);
not NOT1 (N5657, N5645);
xor XOR2 (N5658, N5642, N4955);
xor XOR2 (N5659, N5653, N3670);
or OR4 (N5660, N5657, N5475, N5301, N1863);
nand NAND4 (N5661, N5655, N4407, N3349, N2329);
nor NOR3 (N5662, N5649, N2939, N4240);
or OR3 (N5663, N5658, N497, N2479);
or OR4 (N5664, N5652, N729, N3726, N5652);
buf BUF1 (N5665, N5664);
nand NAND3 (N5666, N5665, N4964, N2577);
and AND2 (N5667, N5661, N351);
and AND3 (N5668, N5651, N3862, N5541);
nor NOR4 (N5669, N5666, N2601, N1247, N1405);
not NOT1 (N5670, N5630);
buf BUF1 (N5671, N5656);
or OR4 (N5672, N5667, N1469, N4436, N194);
nor NOR3 (N5673, N5659, N2475, N4313);
or OR3 (N5674, N5662, N4663, N5435);
nor NOR4 (N5675, N5670, N1958, N751, N2185);
not NOT1 (N5676, N5669);
or OR3 (N5677, N5676, N767, N4462);
xor XOR2 (N5678, N5675, N5454);
not NOT1 (N5679, N5677);
nor NOR2 (N5680, N5654, N4301);
nand NAND4 (N5681, N5673, N326, N2973, N72);
nand NAND2 (N5682, N5668, N2360);
or OR2 (N5683, N5678, N5291);
nand NAND4 (N5684, N5672, N5448, N2179, N3210);
not NOT1 (N5685, N5680);
not NOT1 (N5686, N5683);
not NOT1 (N5687, N5660);
not NOT1 (N5688, N5682);
buf BUF1 (N5689, N5685);
and AND4 (N5690, N5686, N1463, N4563, N153);
nor NOR4 (N5691, N5687, N4089, N3400, N3534);
xor XOR2 (N5692, N5688, N2970);
and AND3 (N5693, N5663, N2832, N2085);
and AND3 (N5694, N5690, N4176, N2267);
or OR3 (N5695, N5689, N3025, N3049);
nor NOR4 (N5696, N5671, N2529, N929, N647);
and AND2 (N5697, N5674, N81);
nand NAND3 (N5698, N5697, N217, N5205);
and AND2 (N5699, N5681, N2572);
and AND2 (N5700, N5693, N4043);
and AND2 (N5701, N5698, N2229);
nor NOR3 (N5702, N5701, N3978, N2950);
and AND2 (N5703, N5699, N2022);
nand NAND4 (N5704, N5684, N1393, N5069, N2476);
nor NOR2 (N5705, N5700, N575);
buf BUF1 (N5706, N5694);
or OR4 (N5707, N5706, N2826, N2427, N1077);
and AND4 (N5708, N5707, N638, N3007, N2987);
nand NAND3 (N5709, N5703, N4146, N2278);
nor NOR3 (N5710, N5702, N4468, N3546);
xor XOR2 (N5711, N5708, N1419);
or OR2 (N5712, N5679, N2668);
and AND3 (N5713, N5692, N3671, N1772);
not NOT1 (N5714, N5695);
or OR3 (N5715, N5713, N3307, N4064);
nand NAND2 (N5716, N5712, N4424);
and AND3 (N5717, N5715, N15, N5466);
xor XOR2 (N5718, N5710, N3976);
nor NOR2 (N5719, N5718, N2609);
buf BUF1 (N5720, N5717);
xor XOR2 (N5721, N5704, N608);
not NOT1 (N5722, N5705);
or OR4 (N5723, N5719, N1536, N2515, N365);
and AND3 (N5724, N5721, N2308, N4910);
not NOT1 (N5725, N5724);
and AND4 (N5726, N5725, N3048, N1313, N4747);
nor NOR4 (N5727, N5726, N3502, N5255, N307);
or OR4 (N5728, N5723, N3751, N3226, N2222);
nor NOR2 (N5729, N5696, N4515);
xor XOR2 (N5730, N5711, N355);
nor NOR3 (N5731, N5714, N5604, N1110);
nand NAND4 (N5732, N5727, N4537, N4184, N371);
and AND2 (N5733, N5716, N4591);
nand NAND3 (N5734, N5733, N3823, N4886);
or OR4 (N5735, N5730, N188, N2836, N2131);
xor XOR2 (N5736, N5729, N2758);
nor NOR2 (N5737, N5728, N3322);
or OR2 (N5738, N5734, N4320);
nand NAND4 (N5739, N5722, N4151, N4838, N5193);
and AND2 (N5740, N5731, N1405);
nand NAND2 (N5741, N5720, N1189);
xor XOR2 (N5742, N5709, N4067);
not NOT1 (N5743, N5737);
or OR4 (N5744, N5735, N987, N4873, N4636);
buf BUF1 (N5745, N5732);
nand NAND4 (N5746, N5745, N1502, N1034, N1126);
buf BUF1 (N5747, N5738);
xor XOR2 (N5748, N5739, N1307);
nand NAND3 (N5749, N5736, N2683, N3733);
or OR4 (N5750, N5747, N1732, N4758, N3951);
xor XOR2 (N5751, N5749, N5059);
not NOT1 (N5752, N5751);
and AND3 (N5753, N5748, N5606, N2537);
xor XOR2 (N5754, N5752, N3239);
or OR3 (N5755, N5744, N2095, N3921);
buf BUF1 (N5756, N5754);
xor XOR2 (N5757, N5753, N3975);
and AND3 (N5758, N5742, N2569, N523);
and AND2 (N5759, N5757, N688);
buf BUF1 (N5760, N5750);
xor XOR2 (N5761, N5741, N4032);
and AND2 (N5762, N5746, N5704);
buf BUF1 (N5763, N5756);
xor XOR2 (N5764, N5758, N3682);
and AND4 (N5765, N5691, N3668, N2425, N81);
not NOT1 (N5766, N5740);
nor NOR2 (N5767, N5766, N131);
xor XOR2 (N5768, N5762, N2919);
or OR3 (N5769, N5767, N5598, N4757);
not NOT1 (N5770, N5764);
and AND4 (N5771, N5770, N624, N4414, N2182);
xor XOR2 (N5772, N5760, N2221);
xor XOR2 (N5773, N5759, N1460);
nor NOR4 (N5774, N5743, N3034, N3587, N2706);
and AND3 (N5775, N5765, N1660, N4345);
nand NAND4 (N5776, N5761, N1974, N945, N1791);
nor NOR4 (N5777, N5776, N438, N3449, N2956);
and AND4 (N5778, N5773, N2398, N1495, N5088);
nand NAND3 (N5779, N5763, N2078, N3118);
buf BUF1 (N5780, N5779);
nor NOR3 (N5781, N5774, N5056, N1927);
buf BUF1 (N5782, N5775);
nor NOR3 (N5783, N5777, N1254, N3426);
buf BUF1 (N5784, N5778);
or OR4 (N5785, N5755, N2204, N1442, N2530);
nor NOR3 (N5786, N5771, N5544, N733);
or OR3 (N5787, N5768, N1784, N2282);
nand NAND2 (N5788, N5782, N3540);
and AND2 (N5789, N5780, N3486);
xor XOR2 (N5790, N5787, N2097);
nor NOR2 (N5791, N5772, N3637);
and AND4 (N5792, N5783, N4618, N4496, N2272);
or OR2 (N5793, N5769, N1642);
and AND3 (N5794, N5792, N4696, N5417);
nor NOR3 (N5795, N5785, N1014, N4607);
buf BUF1 (N5796, N5788);
xor XOR2 (N5797, N5794, N106);
and AND4 (N5798, N5781, N3428, N1590, N3567);
buf BUF1 (N5799, N5790);
xor XOR2 (N5800, N5791, N4937);
nor NOR4 (N5801, N5798, N1727, N4647, N5143);
nor NOR3 (N5802, N5795, N1488, N372);
and AND2 (N5803, N5793, N1730);
nand NAND3 (N5804, N5802, N4850, N4985);
nand NAND2 (N5805, N5801, N1658);
buf BUF1 (N5806, N5784);
nor NOR3 (N5807, N5800, N298, N5744);
nand NAND2 (N5808, N5797, N1825);
buf BUF1 (N5809, N5786);
nor NOR3 (N5810, N5807, N936, N711);
not NOT1 (N5811, N5809);
xor XOR2 (N5812, N5806, N3024);
nand NAND2 (N5813, N5796, N1193);
nor NOR2 (N5814, N5804, N2372);
not NOT1 (N5815, N5811);
nand NAND2 (N5816, N5813, N710);
not NOT1 (N5817, N5816);
nor NOR4 (N5818, N5789, N4558, N5777, N3471);
not NOT1 (N5819, N5810);
not NOT1 (N5820, N5808);
buf BUF1 (N5821, N5805);
not NOT1 (N5822, N5818);
or OR2 (N5823, N5817, N4184);
not NOT1 (N5824, N5820);
and AND3 (N5825, N5815, N5781, N682);
or OR4 (N5826, N5824, N3074, N236, N5110);
nand NAND3 (N5827, N5821, N2889, N1743);
not NOT1 (N5828, N5814);
xor XOR2 (N5829, N5812, N4601);
xor XOR2 (N5830, N5827, N2748);
xor XOR2 (N5831, N5825, N2320);
or OR3 (N5832, N5831, N2404, N5362);
nand NAND3 (N5833, N5823, N4663, N704);
or OR4 (N5834, N5799, N1363, N431, N1094);
xor XOR2 (N5835, N5832, N1630);
not NOT1 (N5836, N5826);
buf BUF1 (N5837, N5828);
not NOT1 (N5838, N5819);
and AND3 (N5839, N5803, N77, N1587);
and AND3 (N5840, N5836, N585, N1504);
nand NAND3 (N5841, N5835, N3196, N699);
and AND2 (N5842, N5841, N3399);
not NOT1 (N5843, N5839);
or OR2 (N5844, N5842, N5489);
or OR3 (N5845, N5829, N5840, N520);
not NOT1 (N5846, N106);
buf BUF1 (N5847, N5843);
not NOT1 (N5848, N5846);
nor NOR3 (N5849, N5830, N43, N2716);
and AND2 (N5850, N5844, N3105);
nor NOR4 (N5851, N5845, N4852, N630, N2145);
xor XOR2 (N5852, N5837, N3477);
nor NOR4 (N5853, N5833, N5135, N4940, N5512);
not NOT1 (N5854, N5851);
or OR2 (N5855, N5854, N1182);
and AND4 (N5856, N5848, N5515, N1338, N1950);
buf BUF1 (N5857, N5849);
nor NOR4 (N5858, N5856, N5847, N2580, N930);
nand NAND2 (N5859, N678, N154);
and AND3 (N5860, N5853, N1745, N1314);
buf BUF1 (N5861, N5855);
buf BUF1 (N5862, N5850);
nand NAND2 (N5863, N5838, N1130);
xor XOR2 (N5864, N5822, N3313);
nand NAND4 (N5865, N5857, N3680, N746, N2443);
nand NAND2 (N5866, N5861, N3157);
not NOT1 (N5867, N5864);
xor XOR2 (N5868, N5852, N3405);
not NOT1 (N5869, N5860);
or OR4 (N5870, N5869, N2481, N3284, N2251);
and AND4 (N5871, N5868, N3945, N5511, N2445);
xor XOR2 (N5872, N5863, N1767);
nor NOR3 (N5873, N5865, N6, N370);
buf BUF1 (N5874, N5834);
nand NAND4 (N5875, N5874, N4257, N2880, N4774);
or OR3 (N5876, N5873, N5002, N4150);
or OR2 (N5877, N5870, N2851);
xor XOR2 (N5878, N5866, N2273);
not NOT1 (N5879, N5871);
not NOT1 (N5880, N5867);
and AND2 (N5881, N5880, N2889);
buf BUF1 (N5882, N5877);
buf BUF1 (N5883, N5876);
nand NAND4 (N5884, N5858, N656, N3214, N820);
nor NOR2 (N5885, N5884, N5090);
not NOT1 (N5886, N5862);
nand NAND2 (N5887, N5875, N4024);
not NOT1 (N5888, N5883);
buf BUF1 (N5889, N5879);
nor NOR4 (N5890, N5887, N2303, N800, N3475);
xor XOR2 (N5891, N5890, N5088);
xor XOR2 (N5892, N5882, N370);
or OR3 (N5893, N5859, N1196, N3011);
nand NAND3 (N5894, N5893, N569, N3407);
nor NOR4 (N5895, N5872, N1456, N2059, N3335);
or OR2 (N5896, N5895, N3151);
and AND2 (N5897, N5891, N5151);
nand NAND2 (N5898, N5888, N4654);
buf BUF1 (N5899, N5897);
not NOT1 (N5900, N5885);
and AND2 (N5901, N5898, N1466);
not NOT1 (N5902, N5881);
nand NAND3 (N5903, N5892, N4867, N1037);
buf BUF1 (N5904, N5878);
not NOT1 (N5905, N5889);
and AND4 (N5906, N5900, N5488, N3539, N2685);
xor XOR2 (N5907, N5886, N4449);
not NOT1 (N5908, N5905);
buf BUF1 (N5909, N5899);
not NOT1 (N5910, N5903);
or OR3 (N5911, N5908, N718, N2309);
or OR2 (N5912, N5902, N5565);
nor NOR2 (N5913, N5912, N243);
buf BUF1 (N5914, N5901);
xor XOR2 (N5915, N5907, N5572);
nand NAND2 (N5916, N5910, N5811);
or OR2 (N5917, N5909, N3310);
nor NOR2 (N5918, N5906, N2511);
nor NOR3 (N5919, N5894, N5245, N2091);
nand NAND4 (N5920, N5911, N4488, N1400, N3672);
nor NOR3 (N5921, N5915, N3919, N1157);
not NOT1 (N5922, N5920);
nand NAND4 (N5923, N5918, N4345, N2860, N1068);
or OR3 (N5924, N5919, N4586, N3388);
and AND3 (N5925, N5913, N5496, N59);
xor XOR2 (N5926, N5922, N4010);
or OR3 (N5927, N5921, N1646, N2898);
not NOT1 (N5928, N5896);
xor XOR2 (N5929, N5923, N5210);
or OR3 (N5930, N5926, N90, N5580);
nand NAND2 (N5931, N5904, N1703);
xor XOR2 (N5932, N5931, N1239);
not NOT1 (N5933, N5917);
xor XOR2 (N5934, N5925, N398);
buf BUF1 (N5935, N5934);
nand NAND2 (N5936, N5932, N3202);
nand NAND3 (N5937, N5930, N5613, N3982);
not NOT1 (N5938, N5916);
nor NOR3 (N5939, N5936, N1184, N298);
or OR4 (N5940, N5924, N4100, N5879, N235);
xor XOR2 (N5941, N5927, N1985);
buf BUF1 (N5942, N5933);
not NOT1 (N5943, N5937);
buf BUF1 (N5944, N5929);
xor XOR2 (N5945, N5940, N5739);
not NOT1 (N5946, N5914);
and AND4 (N5947, N5935, N4018, N3814, N3800);
not NOT1 (N5948, N5943);
and AND2 (N5949, N5947, N2671);
xor XOR2 (N5950, N5939, N4977);
and AND3 (N5951, N5948, N3391, N2971);
or OR3 (N5952, N5951, N3046, N3558);
nor NOR4 (N5953, N5952, N1771, N893, N433);
xor XOR2 (N5954, N5938, N559);
or OR4 (N5955, N5944, N1178, N3188, N5757);
buf BUF1 (N5956, N5950);
buf BUF1 (N5957, N5953);
and AND2 (N5958, N5957, N2700);
xor XOR2 (N5959, N5954, N1616);
xor XOR2 (N5960, N5945, N839);
not NOT1 (N5961, N5959);
and AND4 (N5962, N5928, N1931, N3861, N2497);
buf BUF1 (N5963, N5946);
xor XOR2 (N5964, N5956, N4769);
xor XOR2 (N5965, N5960, N2130);
nor NOR4 (N5966, N5962, N1219, N5711, N2741);
not NOT1 (N5967, N5949);
or OR4 (N5968, N5963, N5559, N4675, N2066);
or OR2 (N5969, N5955, N8);
and AND4 (N5970, N5967, N1895, N4631, N1400);
nor NOR3 (N5971, N5961, N4553, N1574);
and AND3 (N5972, N5942, N961, N5039);
and AND2 (N5973, N5969, N1630);
or OR4 (N5974, N5973, N818, N1145, N3258);
not NOT1 (N5975, N5965);
and AND2 (N5976, N5975, N2656);
and AND3 (N5977, N5971, N5908, N1958);
and AND3 (N5978, N5958, N3968, N2401);
buf BUF1 (N5979, N5970);
nor NOR3 (N5980, N5978, N1404, N5970);
or OR3 (N5981, N5941, N2133, N5765);
nand NAND3 (N5982, N5980, N73, N2272);
not NOT1 (N5983, N5968);
not NOT1 (N5984, N5981);
nand NAND4 (N5985, N5972, N5198, N4660, N5700);
not NOT1 (N5986, N5977);
nand NAND4 (N5987, N5985, N5112, N2427, N3981);
and AND4 (N5988, N5982, N3107, N5485, N2379);
and AND4 (N5989, N5979, N4221, N40, N3733);
not NOT1 (N5990, N5987);
nand NAND3 (N5991, N5964, N5148, N2129);
buf BUF1 (N5992, N5983);
buf BUF1 (N5993, N5966);
and AND3 (N5994, N5986, N3686, N1983);
nor NOR2 (N5995, N5989, N3718);
nor NOR4 (N5996, N5990, N1818, N1741, N5351);
buf BUF1 (N5997, N5993);
buf BUF1 (N5998, N5994);
or OR3 (N5999, N5998, N2084, N4700);
and AND4 (N6000, N5996, N1879, N3203, N882);
or OR4 (N6001, N5991, N3627, N2676, N868);
xor XOR2 (N6002, N5988, N4671);
buf BUF1 (N6003, N5992);
nand NAND3 (N6004, N6000, N4766, N5496);
or OR2 (N6005, N6002, N3149);
nor NOR4 (N6006, N5974, N4869, N2131, N1580);
buf BUF1 (N6007, N6005);
xor XOR2 (N6008, N5995, N5347);
nand NAND4 (N6009, N5997, N3868, N1421, N5691);
nor NOR2 (N6010, N5976, N1661);
or OR3 (N6011, N5999, N2431, N2846);
nand NAND3 (N6012, N6009, N449, N5128);
and AND3 (N6013, N6012, N5207, N3491);
buf BUF1 (N6014, N6004);
nor NOR4 (N6015, N6001, N2459, N1878, N4311);
xor XOR2 (N6016, N6007, N347);
or OR3 (N6017, N5984, N783, N5110);
nand NAND4 (N6018, N6011, N119, N817, N1253);
or OR4 (N6019, N6013, N1409, N5032, N4813);
nor NOR4 (N6020, N6010, N5001, N5020, N1196);
not NOT1 (N6021, N6006);
not NOT1 (N6022, N6016);
not NOT1 (N6023, N6021);
or OR3 (N6024, N6018, N4538, N2738);
not NOT1 (N6025, N6017);
not NOT1 (N6026, N6025);
nand NAND4 (N6027, N6003, N5678, N462, N674);
nand NAND3 (N6028, N6019, N654, N3595);
or OR4 (N6029, N6028, N636, N2739, N3097);
xor XOR2 (N6030, N6020, N5286);
and AND2 (N6031, N6014, N3460);
buf BUF1 (N6032, N6029);
nand NAND4 (N6033, N6008, N2084, N3756, N444);
xor XOR2 (N6034, N6022, N2453);
buf BUF1 (N6035, N6033);
or OR3 (N6036, N6015, N3792, N1310);
nand NAND4 (N6037, N6027, N488, N2912, N3959);
xor XOR2 (N6038, N6031, N4404);
xor XOR2 (N6039, N6037, N995);
not NOT1 (N6040, N6039);
and AND4 (N6041, N6034, N4484, N2048, N3439);
buf BUF1 (N6042, N6026);
buf BUF1 (N6043, N6032);
not NOT1 (N6044, N6038);
xor XOR2 (N6045, N6030, N3577);
nand NAND4 (N6046, N6045, N5820, N492, N566);
or OR2 (N6047, N6023, N1890);
and AND4 (N6048, N6035, N1719, N5678, N3733);
buf BUF1 (N6049, N6024);
nand NAND4 (N6050, N6040, N5875, N3160, N4598);
buf BUF1 (N6051, N6042);
or OR4 (N6052, N6046, N3785, N5690, N3576);
nor NOR3 (N6053, N6048, N5583, N4928);
not NOT1 (N6054, N6052);
nor NOR3 (N6055, N6054, N5381, N4471);
buf BUF1 (N6056, N6055);
nand NAND3 (N6057, N6044, N2563, N2087);
nor NOR2 (N6058, N6057, N544);
buf BUF1 (N6059, N6051);
and AND2 (N6060, N6053, N4677);
and AND4 (N6061, N6056, N5326, N5112, N5254);
and AND2 (N6062, N6041, N1469);
not NOT1 (N6063, N6058);
nand NAND2 (N6064, N6060, N3695);
and AND3 (N6065, N6062, N3318, N4659);
not NOT1 (N6066, N6059);
xor XOR2 (N6067, N6049, N2490);
or OR3 (N6068, N6067, N5496, N1723);
not NOT1 (N6069, N6061);
not NOT1 (N6070, N6050);
not NOT1 (N6071, N6068);
and AND4 (N6072, N6036, N2118, N5257, N3610);
nor NOR2 (N6073, N6063, N4243);
nand NAND3 (N6074, N6047, N5617, N26);
buf BUF1 (N6075, N6073);
nand NAND4 (N6076, N6071, N3837, N1, N5844);
or OR2 (N6077, N6043, N1146);
buf BUF1 (N6078, N6069);
or OR4 (N6079, N6070, N541, N3091, N3703);
not NOT1 (N6080, N6074);
or OR4 (N6081, N6072, N1578, N5300, N714);
not NOT1 (N6082, N6079);
buf BUF1 (N6083, N6082);
and AND3 (N6084, N6081, N3870, N2640);
buf BUF1 (N6085, N6077);
xor XOR2 (N6086, N6085, N752);
xor XOR2 (N6087, N6064, N2376);
nand NAND3 (N6088, N6075, N367, N4130);
buf BUF1 (N6089, N6087);
nand NAND2 (N6090, N6088, N5216);
and AND2 (N6091, N6076, N3456);
and AND4 (N6092, N6091, N1870, N2151, N2695);
not NOT1 (N6093, N6090);
not NOT1 (N6094, N6083);
not NOT1 (N6095, N6065);
buf BUF1 (N6096, N6084);
buf BUF1 (N6097, N6094);
nor NOR4 (N6098, N6089, N2336, N966, N406);
not NOT1 (N6099, N6095);
or OR4 (N6100, N6066, N2102, N1018, N1858);
nand NAND3 (N6101, N6093, N224, N623);
or OR4 (N6102, N6100, N3040, N5368, N1679);
nor NOR4 (N6103, N6099, N1800, N1099, N2141);
xor XOR2 (N6104, N6092, N5258);
or OR3 (N6105, N6096, N79, N5621);
not NOT1 (N6106, N6097);
nand NAND2 (N6107, N6105, N3771);
xor XOR2 (N6108, N6080, N5892);
nor NOR3 (N6109, N6078, N2391, N3047);
nand NAND3 (N6110, N6106, N2857, N5614);
nor NOR4 (N6111, N6102, N3276, N5778, N2002);
and AND3 (N6112, N6086, N4428, N3702);
buf BUF1 (N6113, N6107);
not NOT1 (N6114, N6111);
xor XOR2 (N6115, N6108, N2188);
or OR2 (N6116, N6098, N3884);
not NOT1 (N6117, N6113);
buf BUF1 (N6118, N6117);
not NOT1 (N6119, N6118);
not NOT1 (N6120, N6104);
nand NAND3 (N6121, N6110, N4371, N2062);
xor XOR2 (N6122, N6119, N4972);
or OR2 (N6123, N6112, N2143);
nand NAND2 (N6124, N6123, N4481);
nor NOR2 (N6125, N6122, N2620);
nor NOR3 (N6126, N6120, N1091, N5333);
or OR4 (N6127, N6124, N420, N2059, N1725);
xor XOR2 (N6128, N6126, N1637);
or OR2 (N6129, N6101, N3177);
and AND3 (N6130, N6127, N2515, N3807);
or OR4 (N6131, N6115, N5713, N3221, N3073);
nand NAND2 (N6132, N6130, N5244);
and AND4 (N6133, N6131, N225, N485, N5829);
and AND4 (N6134, N6114, N2168, N5523, N2847);
nand NAND4 (N6135, N6121, N2626, N5016, N4340);
xor XOR2 (N6136, N6103, N779);
nand NAND4 (N6137, N6128, N1809, N4876, N4304);
nand NAND3 (N6138, N6129, N6024, N3609);
or OR3 (N6139, N6125, N5505, N4520);
nor NOR2 (N6140, N6132, N3892);
nand NAND2 (N6141, N6134, N3571);
and AND2 (N6142, N6109, N5942);
nor NOR2 (N6143, N6135, N4480);
nand NAND3 (N6144, N6133, N5375, N461);
nand NAND2 (N6145, N6141, N3072);
xor XOR2 (N6146, N6144, N4995);
buf BUF1 (N6147, N6140);
xor XOR2 (N6148, N6145, N3987);
not NOT1 (N6149, N6147);
not NOT1 (N6150, N6142);
and AND4 (N6151, N6138, N2809, N296, N3884);
buf BUF1 (N6152, N6151);
xor XOR2 (N6153, N6143, N1262);
buf BUF1 (N6154, N6148);
buf BUF1 (N6155, N6146);
and AND2 (N6156, N6150, N3612);
not NOT1 (N6157, N6149);
and AND2 (N6158, N6157, N987);
or OR3 (N6159, N6139, N1664, N3869);
xor XOR2 (N6160, N6116, N4119);
and AND3 (N6161, N6136, N2141, N4372);
not NOT1 (N6162, N6159);
nor NOR3 (N6163, N6160, N1913, N5929);
nand NAND2 (N6164, N6158, N1561);
xor XOR2 (N6165, N6161, N1613);
buf BUF1 (N6166, N6165);
xor XOR2 (N6167, N6164, N5691);
xor XOR2 (N6168, N6156, N107);
or OR2 (N6169, N6166, N5921);
nor NOR2 (N6170, N6167, N5477);
xor XOR2 (N6171, N6170, N2029);
buf BUF1 (N6172, N6153);
and AND2 (N6173, N6163, N4689);
nand NAND4 (N6174, N6173, N1015, N5453, N1039);
or OR4 (N6175, N6154, N38, N3524, N4844);
nor NOR4 (N6176, N6162, N247, N2736, N2356);
or OR4 (N6177, N6172, N6094, N2391, N2894);
or OR3 (N6178, N6175, N5945, N1604);
nand NAND2 (N6179, N6178, N4816);
xor XOR2 (N6180, N6171, N2302);
or OR2 (N6181, N6176, N2729);
buf BUF1 (N6182, N6179);
nand NAND4 (N6183, N6152, N2015, N2169, N1751);
and AND3 (N6184, N6137, N1428, N2826);
not NOT1 (N6185, N6177);
not NOT1 (N6186, N6182);
buf BUF1 (N6187, N6169);
nand NAND2 (N6188, N6155, N1260);
or OR4 (N6189, N6184, N2689, N1086, N330);
xor XOR2 (N6190, N6188, N395);
not NOT1 (N6191, N6186);
not NOT1 (N6192, N6190);
buf BUF1 (N6193, N6180);
nand NAND3 (N6194, N6189, N3415, N5659);
xor XOR2 (N6195, N6193, N3966);
or OR2 (N6196, N6183, N1972);
not NOT1 (N6197, N6185);
nor NOR2 (N6198, N6187, N2035);
or OR2 (N6199, N6174, N3812);
xor XOR2 (N6200, N6198, N144);
nand NAND3 (N6201, N6192, N5650, N4028);
or OR4 (N6202, N6181, N856, N4281, N2844);
nor NOR2 (N6203, N6202, N3204);
nor NOR4 (N6204, N6195, N3479, N5163, N224);
nor NOR3 (N6205, N6201, N2491, N5286);
or OR2 (N6206, N6199, N4135);
xor XOR2 (N6207, N6203, N4658);
or OR4 (N6208, N6191, N4372, N3911, N3314);
nor NOR3 (N6209, N6168, N2812, N1328);
or OR2 (N6210, N6197, N151);
xor XOR2 (N6211, N6207, N1430);
nor NOR4 (N6212, N6206, N5823, N4181, N3231);
or OR3 (N6213, N6212, N1054, N2529);
nand NAND3 (N6214, N6205, N4291, N2699);
nor NOR4 (N6215, N6204, N3194, N3093, N5058);
nor NOR2 (N6216, N6208, N5392);
xor XOR2 (N6217, N6214, N282);
nand NAND4 (N6218, N6216, N3952, N3958, N5253);
nor NOR2 (N6219, N6211, N4383);
buf BUF1 (N6220, N6219);
and AND4 (N6221, N6200, N1133, N3379, N3019);
buf BUF1 (N6222, N6213);
nor NOR2 (N6223, N6209, N716);
not NOT1 (N6224, N6217);
not NOT1 (N6225, N6196);
xor XOR2 (N6226, N6218, N2242);
not NOT1 (N6227, N6223);
nor NOR3 (N6228, N6225, N5102, N3569);
or OR3 (N6229, N6222, N2471, N4529);
nor NOR4 (N6230, N6221, N3045, N4717, N4248);
xor XOR2 (N6231, N6226, N2613);
xor XOR2 (N6232, N6224, N203);
buf BUF1 (N6233, N6227);
buf BUF1 (N6234, N6228);
buf BUF1 (N6235, N6232);
or OR4 (N6236, N6235, N891, N1708, N3970);
nor NOR3 (N6237, N6233, N2813, N419);
not NOT1 (N6238, N6215);
and AND3 (N6239, N6236, N2719, N724);
buf BUF1 (N6240, N6229);
nand NAND4 (N6241, N6210, N2168, N623, N2029);
nor NOR3 (N6242, N6239, N3484, N4457);
buf BUF1 (N6243, N6238);
buf BUF1 (N6244, N6220);
nor NOR2 (N6245, N6234, N5691);
buf BUF1 (N6246, N6242);
or OR3 (N6247, N6230, N2853, N1539);
nand NAND3 (N6248, N6243, N5044, N1250);
nand NAND3 (N6249, N6245, N5353, N500);
or OR4 (N6250, N6231, N1391, N1361, N1255);
buf BUF1 (N6251, N6237);
nand NAND2 (N6252, N6250, N2231);
and AND3 (N6253, N6244, N1167, N2555);
or OR3 (N6254, N6240, N4710, N4535);
not NOT1 (N6255, N6254);
nor NOR2 (N6256, N6249, N492);
nor NOR2 (N6257, N6194, N2556);
nor NOR2 (N6258, N6255, N2760);
or OR4 (N6259, N6251, N6226, N4884, N3969);
and AND3 (N6260, N6241, N3130, N4183);
buf BUF1 (N6261, N6260);
not NOT1 (N6262, N6259);
or OR2 (N6263, N6261, N4799);
and AND2 (N6264, N6246, N289);
nor NOR2 (N6265, N6263, N2168);
nor NOR4 (N6266, N6265, N6103, N5268, N3535);
xor XOR2 (N6267, N6248, N807);
not NOT1 (N6268, N6267);
and AND4 (N6269, N6264, N4947, N3124, N5900);
buf BUF1 (N6270, N6269);
xor XOR2 (N6271, N6257, N35);
not NOT1 (N6272, N6266);
buf BUF1 (N6273, N6272);
xor XOR2 (N6274, N6247, N5691);
buf BUF1 (N6275, N6271);
nand NAND4 (N6276, N6275, N6124, N4738, N3660);
or OR4 (N6277, N6268, N2824, N45, N1527);
xor XOR2 (N6278, N6276, N5799);
or OR4 (N6279, N6273, N2921, N2499, N3179);
buf BUF1 (N6280, N6278);
nand NAND2 (N6281, N6270, N4029);
buf BUF1 (N6282, N6279);
and AND4 (N6283, N6253, N6006, N5135, N3068);
xor XOR2 (N6284, N6280, N2774);
or OR4 (N6285, N6274, N1370, N1967, N4347);
nor NOR4 (N6286, N6281, N4970, N5767, N2174);
and AND3 (N6287, N6285, N1499, N2630);
or OR4 (N6288, N6252, N2445, N3874, N352);
nand NAND4 (N6289, N6287, N4223, N2171, N1000);
or OR4 (N6290, N6282, N5793, N3798, N1368);
nand NAND3 (N6291, N6258, N3187, N1466);
nor NOR4 (N6292, N6277, N4291, N4119, N6157);
buf BUF1 (N6293, N6283);
nor NOR3 (N6294, N6292, N2036, N1650);
not NOT1 (N6295, N6291);
or OR2 (N6296, N6256, N2593);
xor XOR2 (N6297, N6296, N5956);
not NOT1 (N6298, N6290);
xor XOR2 (N6299, N6295, N3152);
not NOT1 (N6300, N6289);
buf BUF1 (N6301, N6286);
not NOT1 (N6302, N6284);
or OR4 (N6303, N6302, N5202, N1068, N11);
xor XOR2 (N6304, N6298, N4681);
xor XOR2 (N6305, N6301, N2743);
nor NOR4 (N6306, N6262, N3632, N2627, N2296);
not NOT1 (N6307, N6304);
and AND2 (N6308, N6306, N246);
not NOT1 (N6309, N6297);
nand NAND4 (N6310, N6300, N2439, N4363, N3898);
and AND4 (N6311, N6308, N2126, N279, N2153);
nor NOR3 (N6312, N6288, N5714, N3547);
or OR4 (N6313, N6312, N4820, N1481, N1741);
nor NOR3 (N6314, N6299, N1001, N5344);
or OR4 (N6315, N6307, N5030, N2507, N2089);
and AND3 (N6316, N6311, N537, N4929);
nor NOR4 (N6317, N6293, N1818, N1599, N3752);
nand NAND3 (N6318, N6315, N4082, N265);
xor XOR2 (N6319, N6314, N4614);
buf BUF1 (N6320, N6303);
or OR2 (N6321, N6309, N2041);
nand NAND4 (N6322, N6320, N3325, N5873, N4050);
xor XOR2 (N6323, N6316, N1713);
xor XOR2 (N6324, N6294, N2979);
not NOT1 (N6325, N6313);
or OR3 (N6326, N6322, N6123, N2280);
xor XOR2 (N6327, N6319, N983);
and AND2 (N6328, N6305, N3937);
xor XOR2 (N6329, N6326, N296);
nand NAND3 (N6330, N6318, N4200, N4795);
xor XOR2 (N6331, N6321, N4248);
not NOT1 (N6332, N6331);
not NOT1 (N6333, N6325);
xor XOR2 (N6334, N6323, N30);
or OR4 (N6335, N6334, N834, N1179, N4002);
not NOT1 (N6336, N6324);
buf BUF1 (N6337, N6329);
buf BUF1 (N6338, N6327);
nand NAND3 (N6339, N6337, N1001, N98);
buf BUF1 (N6340, N6339);
or OR4 (N6341, N6335, N922, N1998, N3086);
nand NAND4 (N6342, N6317, N460, N1220, N5489);
not NOT1 (N6343, N6336);
nor NOR4 (N6344, N6328, N3619, N3159, N4029);
and AND2 (N6345, N6340, N1667);
not NOT1 (N6346, N6341);
nand NAND3 (N6347, N6346, N714, N2361);
or OR2 (N6348, N6338, N2827);
buf BUF1 (N6349, N6310);
nand NAND4 (N6350, N6348, N4087, N1647, N2823);
not NOT1 (N6351, N6349);
xor XOR2 (N6352, N6345, N1053);
xor XOR2 (N6353, N6330, N5502);
nor NOR2 (N6354, N6347, N4504);
and AND4 (N6355, N6352, N2767, N5970, N3337);
and AND4 (N6356, N6332, N4198, N2850, N5870);
not NOT1 (N6357, N6351);
nor NOR3 (N6358, N6355, N5794, N3495);
or OR4 (N6359, N6358, N3171, N2079, N4438);
not NOT1 (N6360, N6342);
nand NAND3 (N6361, N6344, N3596, N5318);
buf BUF1 (N6362, N6343);
nand NAND2 (N6363, N6359, N5184);
xor XOR2 (N6364, N6356, N3466);
xor XOR2 (N6365, N6354, N1542);
not NOT1 (N6366, N6360);
or OR4 (N6367, N6353, N5379, N154, N697);
buf BUF1 (N6368, N6366);
not NOT1 (N6369, N6368);
nand NAND2 (N6370, N6361, N5078);
nand NAND2 (N6371, N6350, N1945);
buf BUF1 (N6372, N6357);
buf BUF1 (N6373, N6371);
xor XOR2 (N6374, N6363, N6156);
nor NOR4 (N6375, N6364, N5512, N3011, N5327);
nor NOR4 (N6376, N6367, N4202, N1738, N2766);
nand NAND2 (N6377, N6362, N2887);
xor XOR2 (N6378, N6372, N2861);
nor NOR2 (N6379, N6370, N1569);
nand NAND2 (N6380, N6373, N2353);
and AND2 (N6381, N6376, N5866);
and AND2 (N6382, N6365, N5250);
not NOT1 (N6383, N6375);
xor XOR2 (N6384, N6379, N2076);
xor XOR2 (N6385, N6374, N5976);
xor XOR2 (N6386, N6383, N486);
nor NOR4 (N6387, N6377, N1933, N4828, N2911);
not NOT1 (N6388, N6386);
nand NAND2 (N6389, N6333, N4148);
xor XOR2 (N6390, N6387, N2647);
nand NAND4 (N6391, N6390, N3390, N4624, N464);
buf BUF1 (N6392, N6384);
not NOT1 (N6393, N6385);
nor NOR2 (N6394, N6393, N2126);
buf BUF1 (N6395, N6394);
or OR4 (N6396, N6395, N5522, N4835, N6365);
and AND3 (N6397, N6380, N6041, N545);
nor NOR2 (N6398, N6369, N2443);
or OR3 (N6399, N6381, N6280, N969);
xor XOR2 (N6400, N6388, N1960);
xor XOR2 (N6401, N6399, N2082);
xor XOR2 (N6402, N6400, N6385);
not NOT1 (N6403, N6392);
nor NOR4 (N6404, N6401, N3995, N4574, N1920);
nand NAND2 (N6405, N6378, N1574);
or OR2 (N6406, N6397, N712);
buf BUF1 (N6407, N6404);
or OR2 (N6408, N6402, N4572);
not NOT1 (N6409, N6407);
not NOT1 (N6410, N6409);
not NOT1 (N6411, N6391);
not NOT1 (N6412, N6408);
nand NAND3 (N6413, N6382, N772, N4657);
buf BUF1 (N6414, N6403);
and AND2 (N6415, N6413, N529);
buf BUF1 (N6416, N6396);
and AND4 (N6417, N6405, N2949, N5994, N4037);
buf BUF1 (N6418, N6389);
nor NOR4 (N6419, N6411, N574, N1994, N1690);
nor NOR4 (N6420, N6412, N5786, N5634, N4520);
or OR4 (N6421, N6415, N3914, N3306, N1018);
buf BUF1 (N6422, N6410);
nand NAND3 (N6423, N6419, N5659, N667);
or OR2 (N6424, N6420, N1735);
nand NAND4 (N6425, N6423, N83, N3753, N4044);
and AND2 (N6426, N6414, N3416);
and AND4 (N6427, N6398, N2455, N5485, N1702);
xor XOR2 (N6428, N6421, N1030);
and AND4 (N6429, N6426, N5035, N1455, N3947);
nor NOR2 (N6430, N6424, N6321);
nor NOR4 (N6431, N6427, N2060, N852, N4558);
xor XOR2 (N6432, N6430, N2577);
xor XOR2 (N6433, N6417, N499);
or OR3 (N6434, N6431, N6109, N1894);
or OR2 (N6435, N6425, N5138);
or OR4 (N6436, N6435, N354, N2720, N6354);
not NOT1 (N6437, N6422);
not NOT1 (N6438, N6434);
and AND2 (N6439, N6428, N6164);
or OR3 (N6440, N6439, N6079, N5997);
and AND2 (N6441, N6433, N3497);
xor XOR2 (N6442, N6416, N6342);
xor XOR2 (N6443, N6436, N2887);
xor XOR2 (N6444, N6406, N4908);
and AND3 (N6445, N6429, N1566, N3526);
and AND2 (N6446, N6445, N2312);
buf BUF1 (N6447, N6432);
not NOT1 (N6448, N6446);
xor XOR2 (N6449, N6438, N1687);
nor NOR4 (N6450, N6449, N404, N1990, N1784);
nand NAND3 (N6451, N6437, N5350, N3651);
nor NOR2 (N6452, N6443, N249);
nor NOR4 (N6453, N6418, N5564, N1537, N623);
not NOT1 (N6454, N6447);
nand NAND4 (N6455, N6454, N2595, N5574, N3457);
nor NOR2 (N6456, N6450, N3368);
and AND4 (N6457, N6455, N4761, N6449, N4770);
nor NOR4 (N6458, N6452, N584, N2173, N5685);
nor NOR4 (N6459, N6440, N1169, N1904, N4472);
and AND4 (N6460, N6456, N3712, N1611, N852);
buf BUF1 (N6461, N6451);
xor XOR2 (N6462, N6457, N1074);
not NOT1 (N6463, N6458);
nand NAND3 (N6464, N6462, N1268, N4892);
buf BUF1 (N6465, N6463);
nand NAND4 (N6466, N6461, N262, N3518, N3623);
xor XOR2 (N6467, N6442, N3522);
buf BUF1 (N6468, N6467);
xor XOR2 (N6469, N6464, N2113);
not NOT1 (N6470, N6469);
nand NAND3 (N6471, N6441, N3306, N2168);
xor XOR2 (N6472, N6471, N1390);
or OR2 (N6473, N6448, N2814);
nor NOR4 (N6474, N6468, N747, N3972, N4313);
and AND3 (N6475, N6470, N1239, N5862);
and AND2 (N6476, N6460, N3968);
nor NOR4 (N6477, N6475, N2551, N1946, N1651);
buf BUF1 (N6478, N6472);
and AND4 (N6479, N6477, N4574, N3945, N5930);
nor NOR4 (N6480, N6465, N3453, N2016, N3676);
or OR3 (N6481, N6459, N2199, N4942);
nand NAND4 (N6482, N6453, N1456, N420, N636);
nor NOR4 (N6483, N6482, N106, N665, N1122);
not NOT1 (N6484, N6476);
buf BUF1 (N6485, N6474);
or OR2 (N6486, N6479, N2987);
nor NOR4 (N6487, N6444, N2231, N2087, N5080);
xor XOR2 (N6488, N6473, N2552);
buf BUF1 (N6489, N6480);
buf BUF1 (N6490, N6478);
xor XOR2 (N6491, N6484, N2115);
not NOT1 (N6492, N6491);
or OR3 (N6493, N6492, N3631, N6475);
buf BUF1 (N6494, N6490);
buf BUF1 (N6495, N6488);
and AND4 (N6496, N6487, N3750, N2132, N62);
nor NOR4 (N6497, N6494, N2121, N5234, N34);
xor XOR2 (N6498, N6495, N3532);
buf BUF1 (N6499, N6466);
and AND4 (N6500, N6483, N5128, N5052, N2294);
or OR4 (N6501, N6493, N3169, N3566, N501);
nor NOR2 (N6502, N6489, N156);
and AND4 (N6503, N6496, N212, N3569, N6441);
nand NAND2 (N6504, N6485, N5928);
nor NOR2 (N6505, N6500, N146);
not NOT1 (N6506, N6503);
nor NOR4 (N6507, N6486, N1999, N5098, N4467);
nor NOR3 (N6508, N6481, N928, N2086);
buf BUF1 (N6509, N6498);
or OR4 (N6510, N6504, N6138, N3293, N594);
buf BUF1 (N6511, N6501);
buf BUF1 (N6512, N6510);
and AND2 (N6513, N6508, N941);
not NOT1 (N6514, N6497);
buf BUF1 (N6515, N6506);
xor XOR2 (N6516, N6514, N434);
nand NAND3 (N6517, N6511, N1088, N1272);
xor XOR2 (N6518, N6507, N6411);
or OR4 (N6519, N6502, N55, N1464, N5727);
xor XOR2 (N6520, N6513, N1533);
buf BUF1 (N6521, N6517);
and AND2 (N6522, N6521, N5512);
buf BUF1 (N6523, N6516);
not NOT1 (N6524, N6499);
and AND4 (N6525, N6512, N3837, N6326, N1223);
not NOT1 (N6526, N6515);
nand NAND4 (N6527, N6522, N4364, N6128, N5718);
not NOT1 (N6528, N6505);
nor NOR4 (N6529, N6519, N4091, N5037, N5264);
buf BUF1 (N6530, N6523);
not NOT1 (N6531, N6528);
nor NOR4 (N6532, N6530, N3114, N5694, N169);
xor XOR2 (N6533, N6524, N4708);
not NOT1 (N6534, N6526);
nand NAND4 (N6535, N6527, N5004, N4200, N6503);
not NOT1 (N6536, N6529);
or OR3 (N6537, N6520, N1366, N6274);
xor XOR2 (N6538, N6532, N3141);
nor NOR3 (N6539, N6538, N5858, N6018);
or OR4 (N6540, N6536, N2406, N4420, N5029);
nor NOR4 (N6541, N6531, N3394, N2629, N4146);
or OR3 (N6542, N6509, N6198, N960);
nand NAND4 (N6543, N6518, N5500, N3655, N5933);
xor XOR2 (N6544, N6537, N2309);
or OR3 (N6545, N6541, N3953, N5814);
not NOT1 (N6546, N6542);
buf BUF1 (N6547, N6545);
nor NOR2 (N6548, N6544, N6043);
buf BUF1 (N6549, N6525);
xor XOR2 (N6550, N6548, N2029);
nor NOR2 (N6551, N6535, N6128);
nand NAND2 (N6552, N6540, N4495);
nor NOR4 (N6553, N6552, N4869, N4503, N2175);
not NOT1 (N6554, N6547);
buf BUF1 (N6555, N6550);
and AND4 (N6556, N6555, N5051, N100, N1732);
nor NOR4 (N6557, N6539, N721, N259, N3426);
not NOT1 (N6558, N6554);
nand NAND3 (N6559, N6534, N5761, N3451);
xor XOR2 (N6560, N6556, N5975);
buf BUF1 (N6561, N6559);
nor NOR4 (N6562, N6553, N2679, N6161, N1875);
or OR3 (N6563, N6546, N4164, N680);
nand NAND4 (N6564, N6563, N392, N2634, N5591);
xor XOR2 (N6565, N6549, N3932);
or OR2 (N6566, N6533, N2640);
not NOT1 (N6567, N6566);
and AND2 (N6568, N6543, N472);
buf BUF1 (N6569, N6562);
and AND3 (N6570, N6557, N2354, N5012);
nor NOR4 (N6571, N6570, N685, N3972, N812);
xor XOR2 (N6572, N6569, N1538);
not NOT1 (N6573, N6567);
or OR2 (N6574, N6571, N5549);
nand NAND3 (N6575, N6560, N3633, N2385);
not NOT1 (N6576, N6564);
nand NAND4 (N6577, N6558, N2967, N1280, N1921);
nand NAND4 (N6578, N6561, N3659, N1984, N950);
not NOT1 (N6579, N6577);
buf BUF1 (N6580, N6572);
buf BUF1 (N6581, N6568);
nand NAND3 (N6582, N6580, N1346, N1540);
nand NAND2 (N6583, N6574, N1735);
nor NOR4 (N6584, N6575, N3759, N1789, N1535);
buf BUF1 (N6585, N6579);
xor XOR2 (N6586, N6565, N1998);
nor NOR3 (N6587, N6584, N2952, N6491);
buf BUF1 (N6588, N6573);
and AND4 (N6589, N6582, N4791, N5781, N1331);
not NOT1 (N6590, N6551);
buf BUF1 (N6591, N6587);
nand NAND2 (N6592, N6591, N6121);
xor XOR2 (N6593, N6586, N3897);
xor XOR2 (N6594, N6576, N5615);
xor XOR2 (N6595, N6578, N6362);
nor NOR3 (N6596, N6595, N4034, N5885);
buf BUF1 (N6597, N6593);
xor XOR2 (N6598, N6583, N5016);
nand NAND2 (N6599, N6596, N6070);
xor XOR2 (N6600, N6592, N1346);
buf BUF1 (N6601, N6588);
and AND2 (N6602, N6597, N6392);
and AND2 (N6603, N6598, N5251);
nor NOR3 (N6604, N6585, N235, N2667);
nor NOR3 (N6605, N6590, N2898, N4497);
not NOT1 (N6606, N6594);
buf BUF1 (N6607, N6602);
nand NAND4 (N6608, N6599, N4874, N5483, N5915);
nand NAND2 (N6609, N6600, N330);
and AND2 (N6610, N6606, N4004);
buf BUF1 (N6611, N6609);
not NOT1 (N6612, N6581);
or OR2 (N6613, N6608, N6413);
or OR4 (N6614, N6601, N6010, N5235, N6002);
buf BUF1 (N6615, N6613);
or OR4 (N6616, N6614, N5656, N3458, N455);
not NOT1 (N6617, N6604);
nor NOR4 (N6618, N6610, N2287, N2354, N3112);
or OR3 (N6619, N6612, N4896, N6160);
buf BUF1 (N6620, N6611);
nor NOR4 (N6621, N6618, N4467, N62, N6161);
nor NOR3 (N6622, N6621, N4487, N1876);
buf BUF1 (N6623, N6622);
nand NAND2 (N6624, N6615, N1233);
and AND2 (N6625, N6619, N3791);
not NOT1 (N6626, N6605);
and AND2 (N6627, N6589, N4761);
and AND2 (N6628, N6607, N672);
buf BUF1 (N6629, N6620);
buf BUF1 (N6630, N6626);
and AND2 (N6631, N6627, N809);
nand NAND4 (N6632, N6630, N1146, N4346, N4555);
or OR2 (N6633, N6603, N2994);
buf BUF1 (N6634, N6624);
or OR2 (N6635, N6628, N15);
and AND3 (N6636, N6634, N724, N540);
or OR4 (N6637, N6635, N2986, N5759, N5314);
nand NAND4 (N6638, N6631, N1093, N3500, N3569);
nor NOR4 (N6639, N6616, N2661, N6196, N1717);
not NOT1 (N6640, N6636);
and AND3 (N6641, N6638, N5798, N4467);
not NOT1 (N6642, N6623);
and AND3 (N6643, N6625, N1415, N4070);
and AND3 (N6644, N6629, N4815, N4735);
nor NOR2 (N6645, N6633, N6429);
xor XOR2 (N6646, N6645, N742);
not NOT1 (N6647, N6646);
nor NOR2 (N6648, N6643, N2581);
or OR3 (N6649, N6632, N3561, N887);
buf BUF1 (N6650, N6617);
or OR4 (N6651, N6649, N5540, N6084, N4975);
xor XOR2 (N6652, N6647, N545);
not NOT1 (N6653, N6652);
nand NAND4 (N6654, N6648, N3530, N3558, N1237);
nor NOR3 (N6655, N6640, N4921, N5714);
nand NAND2 (N6656, N6637, N841);
nor NOR2 (N6657, N6654, N5455);
and AND4 (N6658, N6650, N5617, N5406, N5154);
or OR4 (N6659, N6641, N6642, N71, N5366);
buf BUF1 (N6660, N3907);
xor XOR2 (N6661, N6655, N3899);
or OR3 (N6662, N6660, N5629, N5829);
buf BUF1 (N6663, N6656);
buf BUF1 (N6664, N6658);
nor NOR4 (N6665, N6663, N2331, N4435, N3429);
and AND4 (N6666, N6662, N967, N1052, N2065);
or OR4 (N6667, N6639, N4207, N60, N4013);
nand NAND4 (N6668, N6661, N2297, N4755, N1589);
nor NOR4 (N6669, N6664, N4166, N107, N4580);
nor NOR3 (N6670, N6653, N1373, N1001);
not NOT1 (N6671, N6657);
or OR3 (N6672, N6670, N4772, N4822);
and AND2 (N6673, N6672, N78);
buf BUF1 (N6674, N6644);
and AND3 (N6675, N6673, N3783, N5565);
nand NAND4 (N6676, N6667, N4095, N149, N4231);
xor XOR2 (N6677, N6674, N2562);
xor XOR2 (N6678, N6671, N5414);
buf BUF1 (N6679, N6675);
nand NAND3 (N6680, N6666, N2586, N5796);
nand NAND4 (N6681, N6678, N128, N3241, N3080);
nand NAND4 (N6682, N6681, N2045, N5490, N2584);
nand NAND2 (N6683, N6669, N2178);
or OR2 (N6684, N6679, N3638);
xor XOR2 (N6685, N6659, N1557);
or OR4 (N6686, N6682, N2121, N6433, N1010);
nor NOR3 (N6687, N6668, N3005, N261);
and AND4 (N6688, N6683, N3398, N3409, N6248);
nor NOR4 (N6689, N6688, N5969, N6310, N6575);
xor XOR2 (N6690, N6689, N6319);
buf BUF1 (N6691, N6676);
nand NAND4 (N6692, N6684, N2485, N3615, N1394);
and AND3 (N6693, N6680, N1171, N1960);
and AND3 (N6694, N6692, N3682, N5695);
nand NAND3 (N6695, N6691, N3041, N3571);
buf BUF1 (N6696, N6687);
xor XOR2 (N6697, N6686, N1826);
buf BUF1 (N6698, N6695);
buf BUF1 (N6699, N6685);
or OR3 (N6700, N6690, N4817, N5219);
buf BUF1 (N6701, N6698);
or OR3 (N6702, N6696, N616, N4265);
xor XOR2 (N6703, N6694, N1096);
nor NOR3 (N6704, N6651, N1552, N5857);
or OR2 (N6705, N6702, N5543);
nand NAND2 (N6706, N6699, N1734);
buf BUF1 (N6707, N6665);
not NOT1 (N6708, N6693);
xor XOR2 (N6709, N6708, N348);
or OR4 (N6710, N6697, N3677, N2057, N1213);
nand NAND4 (N6711, N6700, N1622, N2812, N5182);
buf BUF1 (N6712, N6701);
not NOT1 (N6713, N6707);
nor NOR3 (N6714, N6704, N3797, N404);
nor NOR3 (N6715, N6709, N1134, N6305);
not NOT1 (N6716, N6712);
or OR3 (N6717, N6706, N5508, N3074);
nor NOR3 (N6718, N6705, N6277, N882);
nand NAND3 (N6719, N6718, N4061, N4204);
buf BUF1 (N6720, N6710);
not NOT1 (N6721, N6677);
or OR3 (N6722, N6716, N3388, N522);
nand NAND4 (N6723, N6720, N1703, N1757, N5875);
xor XOR2 (N6724, N6703, N5134);
nand NAND2 (N6725, N6714, N3918);
buf BUF1 (N6726, N6725);
or OR2 (N6727, N6722, N694);
xor XOR2 (N6728, N6723, N2413);
nand NAND2 (N6729, N6726, N1724);
not NOT1 (N6730, N6717);
or OR3 (N6731, N6711, N3147, N1110);
nand NAND4 (N6732, N6731, N3648, N3844, N2730);
and AND3 (N6733, N6728, N4352, N5737);
buf BUF1 (N6734, N6715);
buf BUF1 (N6735, N6727);
or OR3 (N6736, N6724, N2429, N5539);
xor XOR2 (N6737, N6736, N6566);
not NOT1 (N6738, N6735);
xor XOR2 (N6739, N6719, N3577);
buf BUF1 (N6740, N6734);
not NOT1 (N6741, N6737);
buf BUF1 (N6742, N6733);
nand NAND4 (N6743, N6738, N2059, N4970, N1129);
and AND4 (N6744, N6742, N5138, N3142, N5097);
nor NOR2 (N6745, N6721, N6729);
buf BUF1 (N6746, N5607);
nand NAND4 (N6747, N6732, N771, N3384, N1214);
or OR2 (N6748, N6740, N3520);
and AND2 (N6749, N6748, N1239);
not NOT1 (N6750, N6741);
xor XOR2 (N6751, N6746, N1032);
and AND4 (N6752, N6743, N6254, N240, N644);
not NOT1 (N6753, N6730);
and AND4 (N6754, N6739, N4271, N5581, N6520);
not NOT1 (N6755, N6745);
buf BUF1 (N6756, N6752);
and AND2 (N6757, N6756, N2580);
nand NAND2 (N6758, N6713, N952);
nor NOR3 (N6759, N6749, N1250, N2787);
nand NAND3 (N6760, N6755, N4857, N3441);
xor XOR2 (N6761, N6747, N5590);
not NOT1 (N6762, N6759);
and AND3 (N6763, N6753, N195, N1767);
not NOT1 (N6764, N6750);
nand NAND4 (N6765, N6744, N430, N951, N2704);
or OR3 (N6766, N6751, N6244, N1375);
buf BUF1 (N6767, N6757);
or OR4 (N6768, N6763, N2231, N5676, N1263);
xor XOR2 (N6769, N6765, N1582);
not NOT1 (N6770, N6762);
buf BUF1 (N6771, N6769);
and AND3 (N6772, N6767, N6231, N1770);
nand NAND3 (N6773, N6772, N3423, N3186);
and AND4 (N6774, N6768, N1281, N5091, N561);
not NOT1 (N6775, N6758);
nand NAND4 (N6776, N6754, N201, N2254, N5629);
or OR2 (N6777, N6773, N66);
not NOT1 (N6778, N6761);
xor XOR2 (N6779, N6775, N1940);
nor NOR4 (N6780, N6778, N6190, N3009, N6215);
nor NOR3 (N6781, N6760, N4040, N5367);
nor NOR3 (N6782, N6766, N950, N4717);
xor XOR2 (N6783, N6774, N1546);
nor NOR2 (N6784, N6770, N2831);
nor NOR3 (N6785, N6779, N579, N1051);
not NOT1 (N6786, N6782);
nor NOR3 (N6787, N6785, N2713, N4213);
nor NOR2 (N6788, N6777, N4058);
nand NAND4 (N6789, N6786, N5293, N1152, N5093);
or OR3 (N6790, N6781, N273, N5726);
nor NOR4 (N6791, N6788, N662, N6691, N633);
xor XOR2 (N6792, N6784, N2872);
buf BUF1 (N6793, N6787);
or OR4 (N6794, N6783, N4656, N3360, N3733);
and AND4 (N6795, N6789, N3645, N3415, N642);
not NOT1 (N6796, N6771);
or OR4 (N6797, N6791, N4850, N5524, N5930);
and AND2 (N6798, N6797, N2378);
nand NAND3 (N6799, N6764, N6767, N3133);
xor XOR2 (N6800, N6794, N1538);
xor XOR2 (N6801, N6795, N180);
or OR4 (N6802, N6790, N5029, N1612, N3144);
or OR4 (N6803, N6780, N3170, N6112, N6382);
or OR4 (N6804, N6800, N1746, N6368, N4617);
not NOT1 (N6805, N6799);
buf BUF1 (N6806, N6776);
buf BUF1 (N6807, N6803);
nor NOR2 (N6808, N6801, N4320);
nand NAND3 (N6809, N6808, N2706, N3073);
buf BUF1 (N6810, N6807);
not NOT1 (N6811, N6792);
not NOT1 (N6812, N6793);
nand NAND3 (N6813, N6806, N4640, N2584);
xor XOR2 (N6814, N6812, N6691);
or OR2 (N6815, N6798, N3546);
nor NOR4 (N6816, N6796, N1243, N391, N3442);
nor NOR2 (N6817, N6810, N4032);
buf BUF1 (N6818, N6809);
nand NAND4 (N6819, N6804, N478, N5062, N1353);
nand NAND2 (N6820, N6811, N5948);
and AND3 (N6821, N6805, N5337, N6562);
nand NAND2 (N6822, N6802, N161);
or OR3 (N6823, N6815, N882, N1433);
not NOT1 (N6824, N6819);
not NOT1 (N6825, N6824);
nor NOR4 (N6826, N6821, N6227, N3019, N4908);
or OR3 (N6827, N6825, N2284, N6059);
or OR2 (N6828, N6817, N4127);
xor XOR2 (N6829, N6820, N3421);
or OR2 (N6830, N6827, N1454);
and AND4 (N6831, N6828, N6288, N3703, N3430);
xor XOR2 (N6832, N6829, N2448);
nor NOR2 (N6833, N6832, N4477);
nand NAND2 (N6834, N6813, N3308);
xor XOR2 (N6835, N6823, N1664);
or OR2 (N6836, N6834, N71);
buf BUF1 (N6837, N6818);
xor XOR2 (N6838, N6830, N5269);
buf BUF1 (N6839, N6837);
or OR2 (N6840, N6836, N3832);
nand NAND3 (N6841, N6822, N5524, N2264);
not NOT1 (N6842, N6831);
or OR3 (N6843, N6826, N6032, N6208);
nor NOR3 (N6844, N6835, N1897, N6425);
buf BUF1 (N6845, N6844);
xor XOR2 (N6846, N6839, N1348);
nor NOR4 (N6847, N6841, N3531, N4509, N1554);
and AND4 (N6848, N6814, N1825, N615, N4084);
or OR4 (N6849, N6816, N6442, N5964, N6521);
not NOT1 (N6850, N6843);
and AND2 (N6851, N6842, N4441);
nor NOR3 (N6852, N6845, N4444, N2984);
nand NAND3 (N6853, N6849, N967, N1841);
not NOT1 (N6854, N6846);
not NOT1 (N6855, N6854);
buf BUF1 (N6856, N6840);
nand NAND4 (N6857, N6850, N5870, N3039, N593);
buf BUF1 (N6858, N6838);
not NOT1 (N6859, N6856);
nor NOR3 (N6860, N6853, N1201, N1699);
nand NAND4 (N6861, N6848, N1072, N5534, N2375);
or OR2 (N6862, N6861, N2839);
nor NOR4 (N6863, N6851, N6812, N1909, N2653);
buf BUF1 (N6864, N6863);
xor XOR2 (N6865, N6833, N1640);
nor NOR2 (N6866, N6864, N1180);
nor NOR2 (N6867, N6862, N3175);
not NOT1 (N6868, N6852);
and AND4 (N6869, N6857, N614, N5491, N4361);
buf BUF1 (N6870, N6855);
not NOT1 (N6871, N6858);
or OR3 (N6872, N6860, N658, N6645);
xor XOR2 (N6873, N6870, N2600);
not NOT1 (N6874, N6866);
not NOT1 (N6875, N6859);
nor NOR3 (N6876, N6865, N276, N1597);
buf BUF1 (N6877, N6871);
buf BUF1 (N6878, N6873);
buf BUF1 (N6879, N6847);
buf BUF1 (N6880, N6877);
and AND2 (N6881, N6868, N1907);
or OR4 (N6882, N6880, N5412, N756, N768);
or OR4 (N6883, N6881, N2367, N3659, N4319);
and AND3 (N6884, N6872, N4280, N4069);
and AND4 (N6885, N6875, N3705, N2892, N859);
buf BUF1 (N6886, N6874);
buf BUF1 (N6887, N6886);
not NOT1 (N6888, N6883);
not NOT1 (N6889, N6885);
nor NOR4 (N6890, N6878, N4010, N4072, N4402);
not NOT1 (N6891, N6887);
or OR4 (N6892, N6890, N5072, N5617, N5711);
and AND2 (N6893, N6869, N2886);
or OR4 (N6894, N6891, N2436, N2841, N5807);
nand NAND2 (N6895, N6876, N4932);
nand NAND4 (N6896, N6882, N4964, N2146, N1728);
or OR4 (N6897, N6894, N1376, N470, N2179);
xor XOR2 (N6898, N6895, N5392);
or OR3 (N6899, N6897, N2661, N5320);
or OR2 (N6900, N6892, N4020);
nand NAND4 (N6901, N6896, N588, N3517, N4174);
and AND2 (N6902, N6893, N6700);
nand NAND2 (N6903, N6899, N3084);
nand NAND2 (N6904, N6879, N5708);
buf BUF1 (N6905, N6884);
or OR3 (N6906, N6889, N5940, N698);
not NOT1 (N6907, N6867);
and AND2 (N6908, N6905, N396);
not NOT1 (N6909, N6888);
not NOT1 (N6910, N6909);
and AND2 (N6911, N6904, N1451);
and AND2 (N6912, N6902, N367);
not NOT1 (N6913, N6910);
nand NAND2 (N6914, N6898, N3880);
not NOT1 (N6915, N6906);
buf BUF1 (N6916, N6912);
nand NAND2 (N6917, N6913, N3611);
xor XOR2 (N6918, N6901, N3232);
nor NOR3 (N6919, N6907, N4674, N3744);
xor XOR2 (N6920, N6914, N1118);
nand NAND2 (N6921, N6903, N6683);
not NOT1 (N6922, N6908);
not NOT1 (N6923, N6921);
buf BUF1 (N6924, N6915);
or OR4 (N6925, N6911, N5065, N3451, N1461);
buf BUF1 (N6926, N6900);
not NOT1 (N6927, N6916);
nand NAND3 (N6928, N6920, N5395, N3336);
buf BUF1 (N6929, N6923);
and AND3 (N6930, N6927, N6504, N3062);
xor XOR2 (N6931, N6925, N4363);
nand NAND2 (N6932, N6918, N3181);
and AND4 (N6933, N6919, N6049, N6008, N5499);
buf BUF1 (N6934, N6926);
buf BUF1 (N6935, N6930);
nand NAND3 (N6936, N6932, N2784, N562);
not NOT1 (N6937, N6931);
and AND2 (N6938, N6937, N733);
nor NOR2 (N6939, N6933, N1740);
nor NOR3 (N6940, N6935, N2789, N4990);
and AND4 (N6941, N6924, N3097, N4086, N422);
xor XOR2 (N6942, N6940, N5687);
nand NAND2 (N6943, N6938, N1868);
not NOT1 (N6944, N6942);
not NOT1 (N6945, N6929);
nor NOR3 (N6946, N6934, N151, N3045);
nand NAND3 (N6947, N6917, N445, N1536);
nor NOR4 (N6948, N6947, N3433, N6844, N2612);
nor NOR4 (N6949, N6941, N207, N6377, N541);
not NOT1 (N6950, N6939);
nor NOR3 (N6951, N6945, N2349, N2731);
not NOT1 (N6952, N6949);
nand NAND3 (N6953, N6950, N2107, N3456);
nand NAND3 (N6954, N6922, N3907, N4375);
or OR4 (N6955, N6936, N6250, N6399, N5418);
nor NOR3 (N6956, N6955, N1261, N5814);
buf BUF1 (N6957, N6944);
and AND3 (N6958, N6954, N5474, N5023);
buf BUF1 (N6959, N6957);
not NOT1 (N6960, N6958);
nand NAND4 (N6961, N6928, N2139, N955, N547);
and AND2 (N6962, N6953, N1938);
and AND2 (N6963, N6948, N653);
and AND3 (N6964, N6963, N1667, N6314);
nor NOR3 (N6965, N6943, N4080, N5506);
buf BUF1 (N6966, N6952);
not NOT1 (N6967, N6946);
buf BUF1 (N6968, N6964);
buf BUF1 (N6969, N6965);
buf BUF1 (N6970, N6968);
buf BUF1 (N6971, N6951);
and AND3 (N6972, N6959, N4628, N5346);
not NOT1 (N6973, N6967);
xor XOR2 (N6974, N6970, N6272);
buf BUF1 (N6975, N6962);
nor NOR2 (N6976, N6971, N6187);
xor XOR2 (N6977, N6961, N3683);
buf BUF1 (N6978, N6969);
and AND2 (N6979, N6974, N3073);
or OR2 (N6980, N6973, N5623);
nand NAND3 (N6981, N6976, N671, N5035);
or OR4 (N6982, N6960, N5748, N2263, N2342);
xor XOR2 (N6983, N6956, N3519);
buf BUF1 (N6984, N6977);
nand NAND4 (N6985, N6981, N1122, N3689, N6892);
and AND4 (N6986, N6984, N2570, N5142, N1209);
or OR3 (N6987, N6972, N2926, N3727);
xor XOR2 (N6988, N6986, N815);
not NOT1 (N6989, N6979);
nor NOR2 (N6990, N6985, N5266);
or OR3 (N6991, N6988, N5946, N5674);
nand NAND4 (N6992, N6991, N359, N6414, N6319);
nor NOR4 (N6993, N6982, N3821, N5334, N4029);
and AND4 (N6994, N6983, N2507, N1325, N3295);
and AND2 (N6995, N6994, N5797);
xor XOR2 (N6996, N6975, N5472);
and AND2 (N6997, N6966, N456);
not NOT1 (N6998, N6980);
or OR2 (N6999, N6978, N3882);
buf BUF1 (N7000, N6990);
buf BUF1 (N7001, N6997);
nand NAND3 (N7002, N6995, N3664, N2015);
xor XOR2 (N7003, N6998, N4667);
nand NAND3 (N7004, N7002, N174, N6968);
or OR4 (N7005, N6996, N159, N1236, N3683);
buf BUF1 (N7006, N6999);
not NOT1 (N7007, N7004);
not NOT1 (N7008, N7007);
buf BUF1 (N7009, N7006);
nor NOR2 (N7010, N6992, N163);
and AND2 (N7011, N6989, N2964);
nor NOR3 (N7012, N6993, N6258, N6542);
and AND3 (N7013, N7003, N1105, N5164);
buf BUF1 (N7014, N7005);
nand NAND2 (N7015, N7012, N996);
and AND4 (N7016, N7000, N355, N1814, N6030);
buf BUF1 (N7017, N7001);
or OR4 (N7018, N7017, N5063, N6358, N3533);
nor NOR4 (N7019, N7015, N503, N3503, N757);
or OR3 (N7020, N7013, N4441, N1254);
nand NAND2 (N7021, N7008, N2834);
nor NOR4 (N7022, N7019, N6528, N3634, N2330);
xor XOR2 (N7023, N7014, N6295);
xor XOR2 (N7024, N7011, N3470);
nor NOR2 (N7025, N7021, N2762);
and AND3 (N7026, N7010, N269, N3148);
not NOT1 (N7027, N7026);
buf BUF1 (N7028, N7022);
buf BUF1 (N7029, N7028);
xor XOR2 (N7030, N7018, N4212);
nand NAND3 (N7031, N7027, N4854, N1488);
or OR3 (N7032, N7009, N6591, N6806);
xor XOR2 (N7033, N7020, N5448);
and AND4 (N7034, N6987, N86, N1902, N6644);
or OR2 (N7035, N7023, N5827);
or OR3 (N7036, N7029, N6455, N736);
nand NAND4 (N7037, N7035, N4265, N5866, N5181);
xor XOR2 (N7038, N7034, N3658);
xor XOR2 (N7039, N7032, N5813);
buf BUF1 (N7040, N7031);
nand NAND3 (N7041, N7033, N5292, N262);
nand NAND2 (N7042, N7030, N5116);
nor NOR2 (N7043, N7037, N758);
nor NOR3 (N7044, N7025, N331, N4119);
or OR2 (N7045, N7039, N1698);
nand NAND3 (N7046, N7045, N2781, N3673);
or OR2 (N7047, N7036, N1251);
nor NOR2 (N7048, N7040, N4439);
xor XOR2 (N7049, N7038, N2927);
buf BUF1 (N7050, N7047);
or OR4 (N7051, N7049, N2664, N2716, N6429);
nor NOR3 (N7052, N7024, N6584, N3256);
or OR3 (N7053, N7051, N3262, N3490);
buf BUF1 (N7054, N7050);
nand NAND3 (N7055, N7042, N4505, N95);
nand NAND4 (N7056, N7046, N3451, N4206, N3288);
buf BUF1 (N7057, N7053);
or OR4 (N7058, N7041, N5611, N3237, N226);
and AND3 (N7059, N7052, N6892, N366);
xor XOR2 (N7060, N7057, N3394);
nand NAND4 (N7061, N7060, N1130, N4829, N5233);
and AND2 (N7062, N7055, N3977);
and AND3 (N7063, N7048, N2010, N1952);
nor NOR2 (N7064, N7044, N4821);
xor XOR2 (N7065, N7064, N6099);
and AND2 (N7066, N7063, N3699);
and AND4 (N7067, N7016, N5260, N2086, N2325);
nor NOR4 (N7068, N7066, N545, N4525, N2827);
nand NAND4 (N7069, N7059, N3139, N6358, N5869);
nand NAND4 (N7070, N7062, N1678, N6895, N6153);
xor XOR2 (N7071, N7070, N1594);
xor XOR2 (N7072, N7056, N6010);
buf BUF1 (N7073, N7058);
buf BUF1 (N7074, N7069);
and AND2 (N7075, N7061, N6709);
nand NAND2 (N7076, N7043, N2884);
or OR2 (N7077, N7072, N5738);
not NOT1 (N7078, N7077);
and AND3 (N7079, N7074, N615, N1235);
not NOT1 (N7080, N7078);
nor NOR2 (N7081, N7071, N3604);
or OR3 (N7082, N7076, N3834, N5917);
and AND3 (N7083, N7068, N6365, N5925);
not NOT1 (N7084, N7080);
nor NOR2 (N7085, N7054, N3279);
not NOT1 (N7086, N7081);
not NOT1 (N7087, N7085);
or OR2 (N7088, N7073, N4004);
buf BUF1 (N7089, N7086);
xor XOR2 (N7090, N7089, N2213);
nand NAND3 (N7091, N7087, N5720, N2673);
and AND2 (N7092, N7065, N3019);
nor NOR2 (N7093, N7084, N86);
xor XOR2 (N7094, N7090, N4151);
or OR4 (N7095, N7067, N3062, N6050, N126);
nor NOR4 (N7096, N7075, N1792, N3778, N47);
xor XOR2 (N7097, N7095, N914);
xor XOR2 (N7098, N7088, N2552);
nand NAND3 (N7099, N7091, N3894, N2179);
buf BUF1 (N7100, N7094);
and AND3 (N7101, N7096, N672, N6546);
nor NOR2 (N7102, N7099, N3412);
nor NOR3 (N7103, N7079, N4347, N849);
and AND2 (N7104, N7083, N3276);
or OR3 (N7105, N7102, N5384, N4499);
nor NOR4 (N7106, N7097, N2128, N6718, N5525);
and AND2 (N7107, N7093, N3588);
not NOT1 (N7108, N7105);
nor NOR3 (N7109, N7100, N3854, N3672);
and AND3 (N7110, N7104, N6472, N3691);
buf BUF1 (N7111, N7106);
xor XOR2 (N7112, N7108, N2430);
or OR3 (N7113, N7092, N4662, N3623);
xor XOR2 (N7114, N7098, N3189);
xor XOR2 (N7115, N7111, N771);
and AND4 (N7116, N7082, N801, N3969, N1303);
buf BUF1 (N7117, N7110);
buf BUF1 (N7118, N7103);
and AND4 (N7119, N7112, N3212, N6530, N729);
and AND2 (N7120, N7101, N1164);
xor XOR2 (N7121, N7114, N3183);
or OR3 (N7122, N7119, N3514, N971);
xor XOR2 (N7123, N7115, N2750);
buf BUF1 (N7124, N7122);
nand NAND4 (N7125, N7107, N356, N1162, N1121);
buf BUF1 (N7126, N7121);
xor XOR2 (N7127, N7113, N3310);
xor XOR2 (N7128, N7116, N5261);
or OR3 (N7129, N7109, N6590, N6048);
buf BUF1 (N7130, N7126);
xor XOR2 (N7131, N7127, N5322);
buf BUF1 (N7132, N7123);
or OR3 (N7133, N7131, N4720, N4550);
xor XOR2 (N7134, N7128, N5472);
nand NAND3 (N7135, N7125, N664, N4575);
or OR3 (N7136, N7133, N984, N5820);
or OR2 (N7137, N7120, N3972);
or OR2 (N7138, N7134, N1363);
and AND3 (N7139, N7129, N5089, N1693);
and AND2 (N7140, N7138, N6381);
xor XOR2 (N7141, N7132, N2369);
not NOT1 (N7142, N7117);
and AND4 (N7143, N7124, N4859, N1399, N4913);
xor XOR2 (N7144, N7140, N5507);
xor XOR2 (N7145, N7137, N604);
or OR3 (N7146, N7141, N5370, N1402);
or OR2 (N7147, N7118, N617);
or OR4 (N7148, N7142, N2926, N2820, N211);
buf BUF1 (N7149, N7144);
or OR3 (N7150, N7147, N5603, N5803);
xor XOR2 (N7151, N7150, N1526);
or OR3 (N7152, N7149, N4918, N34);
xor XOR2 (N7153, N7151, N964);
nor NOR2 (N7154, N7135, N2636);
and AND4 (N7155, N7143, N3998, N1375, N327);
not NOT1 (N7156, N7155);
buf BUF1 (N7157, N7139);
and AND2 (N7158, N7154, N949);
and AND2 (N7159, N7153, N4708);
nand NAND3 (N7160, N7158, N783, N4406);
buf BUF1 (N7161, N7160);
nor NOR4 (N7162, N7157, N1707, N6964, N4548);
nor NOR3 (N7163, N7152, N5451, N6790);
nor NOR3 (N7164, N7146, N3176, N6247);
xor XOR2 (N7165, N7159, N5921);
nand NAND4 (N7166, N7156, N2922, N2549, N5715);
or OR4 (N7167, N7162, N3156, N863, N5315);
and AND4 (N7168, N7164, N183, N2989, N4499);
not NOT1 (N7169, N7168);
buf BUF1 (N7170, N7130);
xor XOR2 (N7171, N7167, N3446);
nand NAND4 (N7172, N7145, N2341, N6317, N3395);
xor XOR2 (N7173, N7136, N5176);
not NOT1 (N7174, N7165);
not NOT1 (N7175, N7172);
buf BUF1 (N7176, N7175);
nor NOR2 (N7177, N7174, N3063);
buf BUF1 (N7178, N7161);
or OR2 (N7179, N7166, N2492);
buf BUF1 (N7180, N7177);
nand NAND4 (N7181, N7180, N5880, N1037, N2323);
xor XOR2 (N7182, N7181, N6052);
buf BUF1 (N7183, N7171);
and AND3 (N7184, N7163, N3303, N4348);
and AND3 (N7185, N7183, N1816, N7090);
or OR4 (N7186, N7178, N4354, N1637, N215);
nor NOR4 (N7187, N7186, N3817, N1176, N6878);
or OR3 (N7188, N7169, N6093, N4715);
and AND4 (N7189, N7176, N325, N3135, N3239);
or OR4 (N7190, N7189, N1870, N5881, N6889);
buf BUF1 (N7191, N7184);
buf BUF1 (N7192, N7188);
or OR2 (N7193, N7182, N4946);
nand NAND4 (N7194, N7173, N7089, N643, N7112);
nand NAND4 (N7195, N7148, N5372, N3063, N3547);
buf BUF1 (N7196, N7170);
nand NAND4 (N7197, N7187, N2589, N294, N324);
not NOT1 (N7198, N7193);
nor NOR3 (N7199, N7190, N4840, N5011);
buf BUF1 (N7200, N7195);
nor NOR3 (N7201, N7200, N6699, N4816);
or OR3 (N7202, N7191, N7147, N6892);
or OR4 (N7203, N7201, N4798, N2557, N525);
nand NAND2 (N7204, N7194, N5889);
not NOT1 (N7205, N7199);
not NOT1 (N7206, N7196);
not NOT1 (N7207, N7192);
xor XOR2 (N7208, N7204, N3304);
nand NAND3 (N7209, N7205, N475, N6435);
or OR3 (N7210, N7202, N5640, N6696);
nand NAND3 (N7211, N7203, N819, N1459);
buf BUF1 (N7212, N7207);
and AND3 (N7213, N7206, N6958, N5262);
xor XOR2 (N7214, N7179, N2859);
or OR3 (N7215, N7212, N4586, N662);
or OR2 (N7216, N7198, N6593);
xor XOR2 (N7217, N7215, N2685);
not NOT1 (N7218, N7185);
xor XOR2 (N7219, N7208, N1450);
xor XOR2 (N7220, N7211, N1339);
not NOT1 (N7221, N7209);
and AND3 (N7222, N7217, N109, N226);
not NOT1 (N7223, N7214);
nand NAND3 (N7224, N7221, N5589, N1384);
not NOT1 (N7225, N7216);
not NOT1 (N7226, N7218);
nand NAND2 (N7227, N7210, N4417);
xor XOR2 (N7228, N7219, N4788);
nand NAND2 (N7229, N7224, N5924);
nor NOR2 (N7230, N7227, N1044);
not NOT1 (N7231, N7197);
buf BUF1 (N7232, N7225);
and AND3 (N7233, N7222, N6188, N4240);
nor NOR2 (N7234, N7228, N782);
or OR2 (N7235, N7231, N3968);
buf BUF1 (N7236, N7213);
buf BUF1 (N7237, N7230);
nor NOR4 (N7238, N7233, N7064, N4092, N1894);
xor XOR2 (N7239, N7234, N805);
not NOT1 (N7240, N7223);
or OR2 (N7241, N7238, N3044);
buf BUF1 (N7242, N7226);
and AND4 (N7243, N7235, N6217, N4939, N5152);
and AND3 (N7244, N7241, N258, N28);
xor XOR2 (N7245, N7239, N3970);
nand NAND3 (N7246, N7244, N6687, N3434);
xor XOR2 (N7247, N7237, N4764);
nand NAND3 (N7248, N7236, N148, N5598);
or OR2 (N7249, N7242, N3650);
nor NOR2 (N7250, N7232, N3193);
nor NOR4 (N7251, N7249, N4395, N6055, N3615);
buf BUF1 (N7252, N7229);
nor NOR2 (N7253, N7248, N1695);
buf BUF1 (N7254, N7245);
nor NOR4 (N7255, N7254, N5595, N4005, N1980);
and AND2 (N7256, N7220, N3487);
buf BUF1 (N7257, N7252);
nor NOR4 (N7258, N7253, N3321, N4014, N2851);
nor NOR2 (N7259, N7258, N2039);
or OR3 (N7260, N7255, N1046, N2292);
nor NOR2 (N7261, N7243, N6364);
buf BUF1 (N7262, N7260);
and AND3 (N7263, N7251, N2838, N4253);
nor NOR4 (N7264, N7257, N6997, N1771, N5356);
xor XOR2 (N7265, N7247, N2519);
nor NOR4 (N7266, N7246, N4616, N3176, N1682);
buf BUF1 (N7267, N7259);
and AND4 (N7268, N7261, N3370, N5592, N2584);
or OR3 (N7269, N7250, N2526, N163);
and AND3 (N7270, N7268, N5015, N6162);
or OR4 (N7271, N7256, N255, N5454, N2203);
nand NAND3 (N7272, N7271, N2836, N2028);
nor NOR4 (N7273, N7262, N5449, N4169, N469);
nor NOR3 (N7274, N7266, N6796, N30);
and AND2 (N7275, N7265, N591);
nand NAND4 (N7276, N7275, N291, N4577, N7186);
and AND3 (N7277, N7264, N4724, N1975);
nand NAND2 (N7278, N7240, N6605);
buf BUF1 (N7279, N7277);
and AND3 (N7280, N7272, N1738, N1016);
and AND4 (N7281, N7279, N3751, N3911, N2073);
xor XOR2 (N7282, N7273, N6825);
buf BUF1 (N7283, N7282);
not NOT1 (N7284, N7267);
xor XOR2 (N7285, N7283, N3104);
buf BUF1 (N7286, N7269);
or OR2 (N7287, N7286, N823);
and AND4 (N7288, N7287, N3878, N4729, N4677);
not NOT1 (N7289, N7285);
nand NAND2 (N7290, N7284, N5200);
not NOT1 (N7291, N7276);
xor XOR2 (N7292, N7274, N6552);
buf BUF1 (N7293, N7291);
and AND4 (N7294, N7289, N6079, N6799, N954);
and AND3 (N7295, N7278, N3803, N5435);
and AND3 (N7296, N7290, N3054, N5813);
buf BUF1 (N7297, N7295);
xor XOR2 (N7298, N7296, N644);
not NOT1 (N7299, N7280);
nand NAND3 (N7300, N7270, N4662, N6540);
nand NAND3 (N7301, N7281, N3674, N1858);
xor XOR2 (N7302, N7294, N2075);
nand NAND3 (N7303, N7299, N5437, N134);
not NOT1 (N7304, N7263);
or OR2 (N7305, N7302, N1169);
xor XOR2 (N7306, N7300, N6887);
and AND4 (N7307, N7303, N5975, N2594, N6051);
nand NAND3 (N7308, N7298, N593, N5730);
and AND4 (N7309, N7307, N5639, N6076, N4504);
and AND3 (N7310, N7306, N4460, N6766);
not NOT1 (N7311, N7288);
or OR4 (N7312, N7304, N6247, N823, N3299);
nor NOR2 (N7313, N7301, N4783);
buf BUF1 (N7314, N7310);
buf BUF1 (N7315, N7293);
buf BUF1 (N7316, N7312);
and AND4 (N7317, N7315, N380, N4178, N2386);
nor NOR2 (N7318, N7313, N6622);
and AND3 (N7319, N7314, N6876, N169);
and AND3 (N7320, N7319, N12, N3332);
buf BUF1 (N7321, N7309);
xor XOR2 (N7322, N7297, N4076);
and AND4 (N7323, N7308, N5098, N6612, N3063);
not NOT1 (N7324, N7322);
nor NOR2 (N7325, N7323, N1788);
and AND3 (N7326, N7317, N4219, N336);
buf BUF1 (N7327, N7292);
nor NOR4 (N7328, N7311, N3099, N3429, N3106);
xor XOR2 (N7329, N7318, N3191);
and AND4 (N7330, N7329, N5180, N2037, N6827);
or OR4 (N7331, N7324, N2908, N2299, N999);
nand NAND3 (N7332, N7328, N1890, N5518);
nand NAND3 (N7333, N7327, N1108, N6277);
buf BUF1 (N7334, N7333);
nor NOR2 (N7335, N7330, N5686);
buf BUF1 (N7336, N7334);
nand NAND3 (N7337, N7321, N4728, N2807);
buf BUF1 (N7338, N7332);
xor XOR2 (N7339, N7325, N6692);
nor NOR3 (N7340, N7326, N2021, N5387);
or OR2 (N7341, N7339, N5012);
buf BUF1 (N7342, N7316);
nor NOR4 (N7343, N7341, N2625, N6282, N499);
or OR4 (N7344, N7340, N4395, N303, N2949);
xor XOR2 (N7345, N7343, N4839);
or OR4 (N7346, N7342, N4948, N6289, N6925);
not NOT1 (N7347, N7331);
nor NOR3 (N7348, N7336, N7031, N2853);
buf BUF1 (N7349, N7305);
nor NOR2 (N7350, N7347, N5131);
or OR4 (N7351, N7350, N4929, N5173, N3807);
xor XOR2 (N7352, N7345, N406);
or OR4 (N7353, N7337, N6050, N233, N6867);
and AND4 (N7354, N7335, N361, N512, N7176);
buf BUF1 (N7355, N7352);
nor NOR2 (N7356, N7338, N2603);
nor NOR3 (N7357, N7355, N885, N6258);
nor NOR3 (N7358, N7344, N6498, N4471);
and AND3 (N7359, N7349, N2356, N6030);
nor NOR2 (N7360, N7356, N4829);
not NOT1 (N7361, N7353);
nor NOR3 (N7362, N7348, N5958, N565);
not NOT1 (N7363, N7357);
nand NAND4 (N7364, N7346, N4883, N1933, N5217);
xor XOR2 (N7365, N7362, N6359);
and AND2 (N7366, N7361, N5866);
nor NOR2 (N7367, N7351, N5462);
xor XOR2 (N7368, N7360, N5658);
or OR3 (N7369, N7363, N4974, N7274);
or OR4 (N7370, N7366, N5442, N1232, N1753);
nand NAND2 (N7371, N7354, N3907);
nor NOR4 (N7372, N7367, N2718, N1536, N2970);
nor NOR2 (N7373, N7370, N3740);
nor NOR2 (N7374, N7358, N4890);
nand NAND2 (N7375, N7373, N1027);
xor XOR2 (N7376, N7368, N518);
nor NOR3 (N7377, N7320, N3165, N3683);
nor NOR4 (N7378, N7365, N5516, N6432, N2711);
not NOT1 (N7379, N7364);
or OR3 (N7380, N7377, N1425, N5178);
nand NAND4 (N7381, N7359, N6552, N5712, N2070);
or OR4 (N7382, N7375, N36, N1679, N645);
and AND3 (N7383, N7382, N6260, N525);
or OR4 (N7384, N7376, N4733, N1215, N4610);
or OR2 (N7385, N7369, N1512);
buf BUF1 (N7386, N7380);
nor NOR3 (N7387, N7386, N6360, N5437);
or OR4 (N7388, N7383, N3289, N5268, N761);
or OR4 (N7389, N7387, N5406, N3499, N3419);
nor NOR4 (N7390, N7388, N403, N2004, N5755);
nand NAND2 (N7391, N7378, N621);
not NOT1 (N7392, N7390);
nor NOR2 (N7393, N7381, N1499);
and AND3 (N7394, N7371, N5323, N3767);
nor NOR2 (N7395, N7384, N2953);
nand NAND4 (N7396, N7374, N1177, N5907, N2980);
or OR2 (N7397, N7372, N289);
or OR4 (N7398, N7394, N447, N804, N1637);
and AND4 (N7399, N7397, N6830, N5295, N4876);
buf BUF1 (N7400, N7389);
nand NAND3 (N7401, N7399, N1158, N191);
nor NOR4 (N7402, N7392, N2535, N1899, N5876);
xor XOR2 (N7403, N7396, N4448);
nand NAND2 (N7404, N7391, N6903);
nand NAND2 (N7405, N7393, N3829);
or OR4 (N7406, N7402, N2688, N6709, N1323);
not NOT1 (N7407, N7385);
not NOT1 (N7408, N7379);
nand NAND2 (N7409, N7400, N20);
nor NOR4 (N7410, N7401, N2083, N1165, N3167);
or OR3 (N7411, N7409, N363, N6453);
nand NAND3 (N7412, N7407, N7206, N89);
or OR4 (N7413, N7395, N3236, N6087, N3309);
xor XOR2 (N7414, N7410, N3791);
buf BUF1 (N7415, N7411);
or OR4 (N7416, N7413, N1881, N6799, N2038);
not NOT1 (N7417, N7404);
nand NAND3 (N7418, N7405, N1811, N2238);
nor NOR3 (N7419, N7406, N4863, N4901);
or OR3 (N7420, N7414, N5779, N478);
nor NOR3 (N7421, N7412, N6966, N2671);
nand NAND4 (N7422, N7420, N6950, N7416, N6928);
nor NOR3 (N7423, N4293, N3913, N6656);
nor NOR3 (N7424, N7418, N4599, N5171);
xor XOR2 (N7425, N7408, N5490);
or OR3 (N7426, N7419, N4225, N4783);
not NOT1 (N7427, N7426);
nand NAND4 (N7428, N7423, N4337, N4211, N5899);
xor XOR2 (N7429, N7424, N4530);
and AND2 (N7430, N7422, N2207);
buf BUF1 (N7431, N7403);
or OR3 (N7432, N7417, N6453, N704);
nand NAND4 (N7433, N7425, N396, N4571, N7128);
nand NAND2 (N7434, N7431, N4856);
nand NAND2 (N7435, N7427, N7383);
nand NAND3 (N7436, N7421, N7108, N6273);
not NOT1 (N7437, N7434);
nand NAND4 (N7438, N7428, N4632, N5869, N2959);
not NOT1 (N7439, N7430);
buf BUF1 (N7440, N7398);
not NOT1 (N7441, N7440);
nand NAND2 (N7442, N7433, N5252);
nand NAND4 (N7443, N7442, N2099, N5841, N4832);
not NOT1 (N7444, N7443);
buf BUF1 (N7445, N7439);
and AND3 (N7446, N7432, N5617, N4234);
nand NAND3 (N7447, N7445, N1953, N2820);
and AND2 (N7448, N7444, N5556);
xor XOR2 (N7449, N7446, N2873);
or OR3 (N7450, N7438, N5871, N6736);
not NOT1 (N7451, N7447);
xor XOR2 (N7452, N7448, N3547);
and AND2 (N7453, N7449, N473);
buf BUF1 (N7454, N7429);
or OR3 (N7455, N7441, N551, N3243);
buf BUF1 (N7456, N7452);
or OR2 (N7457, N7456, N6731);
or OR2 (N7458, N7435, N4510);
not NOT1 (N7459, N7454);
xor XOR2 (N7460, N7455, N629);
xor XOR2 (N7461, N7437, N1415);
or OR2 (N7462, N7453, N4295);
nor NOR3 (N7463, N7461, N6937, N177);
nand NAND2 (N7464, N7415, N4840);
and AND2 (N7465, N7459, N4255);
and AND3 (N7466, N7457, N6188, N5809);
not NOT1 (N7467, N7466);
buf BUF1 (N7468, N7436);
and AND2 (N7469, N7464, N3739);
nor NOR2 (N7470, N7465, N2794);
and AND3 (N7471, N7469, N6615, N1467);
xor XOR2 (N7472, N7451, N3553);
buf BUF1 (N7473, N7470);
and AND3 (N7474, N7463, N290, N1508);
not NOT1 (N7475, N7458);
buf BUF1 (N7476, N7473);
or OR4 (N7477, N7468, N5127, N5021, N2798);
or OR2 (N7478, N7450, N1423);
nor NOR4 (N7479, N7475, N5853, N5463, N2336);
or OR2 (N7480, N7467, N7110);
xor XOR2 (N7481, N7478, N6295);
nor NOR4 (N7482, N7460, N5673, N2252, N2241);
and AND3 (N7483, N7472, N3158, N518);
or OR4 (N7484, N7462, N1746, N631, N3720);
or OR2 (N7485, N7477, N2902);
nand NAND2 (N7486, N7485, N3984);
or OR3 (N7487, N7476, N1440, N2909);
and AND4 (N7488, N7482, N4870, N3505, N7348);
nand NAND3 (N7489, N7486, N3009, N1434);
or OR4 (N7490, N7488, N6546, N1272, N4962);
not NOT1 (N7491, N7484);
not NOT1 (N7492, N7480);
not NOT1 (N7493, N7490);
buf BUF1 (N7494, N7491);
nor NOR3 (N7495, N7494, N6505, N7252);
not NOT1 (N7496, N7495);
or OR2 (N7497, N7493, N2122);
and AND2 (N7498, N7487, N7031);
not NOT1 (N7499, N7483);
xor XOR2 (N7500, N7474, N2848);
and AND2 (N7501, N7498, N7166);
or OR2 (N7502, N7489, N1279);
or OR3 (N7503, N7501, N2241, N886);
or OR3 (N7504, N7481, N1830, N309);
not NOT1 (N7505, N7502);
or OR3 (N7506, N7496, N5990, N4662);
buf BUF1 (N7507, N7503);
nor NOR2 (N7508, N7471, N4125);
and AND2 (N7509, N7504, N3930);
or OR4 (N7510, N7508, N6656, N4398, N6121);
xor XOR2 (N7511, N7500, N3138);
buf BUF1 (N7512, N7497);
buf BUF1 (N7513, N7492);
not NOT1 (N7514, N7507);
nor NOR2 (N7515, N7514, N2230);
and AND4 (N7516, N7509, N4155, N3089, N2509);
or OR2 (N7517, N7515, N3914);
and AND3 (N7518, N7506, N2159, N650);
not NOT1 (N7519, N7513);
xor XOR2 (N7520, N7519, N6521);
nor NOR2 (N7521, N7510, N5982);
xor XOR2 (N7522, N7517, N1033);
nor NOR2 (N7523, N7479, N4810);
xor XOR2 (N7524, N7518, N6684);
nand NAND3 (N7525, N7522, N7505, N4204);
xor XOR2 (N7526, N2918, N6665);
nor NOR2 (N7527, N7520, N769);
nand NAND3 (N7528, N7516, N862, N4895);
or OR4 (N7529, N7528, N4857, N2058, N4671);
nand NAND4 (N7530, N7524, N5868, N5042, N6278);
nand NAND2 (N7531, N7526, N2269);
xor XOR2 (N7532, N7499, N7183);
nor NOR3 (N7533, N7521, N7279, N1469);
xor XOR2 (N7534, N7533, N300);
and AND2 (N7535, N7532, N488);
nor NOR2 (N7536, N7534, N3423);
not NOT1 (N7537, N7527);
buf BUF1 (N7538, N7536);
nor NOR2 (N7539, N7535, N4264);
buf BUF1 (N7540, N7531);
xor XOR2 (N7541, N7523, N713);
or OR3 (N7542, N7530, N4900, N3569);
nand NAND4 (N7543, N7541, N2135, N4456, N3744);
buf BUF1 (N7544, N7537);
or OR4 (N7545, N7543, N975, N1109, N7476);
buf BUF1 (N7546, N7540);
nor NOR3 (N7547, N7511, N4911, N5097);
nor NOR4 (N7548, N7542, N491, N434, N7178);
buf BUF1 (N7549, N7529);
and AND4 (N7550, N7546, N2129, N7478, N6909);
or OR4 (N7551, N7548, N6175, N6231, N762);
and AND3 (N7552, N7512, N1112, N4560);
nor NOR2 (N7553, N7551, N2964);
buf BUF1 (N7554, N7538);
not NOT1 (N7555, N7553);
or OR2 (N7556, N7544, N7537);
buf BUF1 (N7557, N7545);
buf BUF1 (N7558, N7539);
and AND3 (N7559, N7556, N1280, N440);
nor NOR4 (N7560, N7550, N1827, N6190, N1776);
not NOT1 (N7561, N7549);
nor NOR2 (N7562, N7561, N1060);
and AND4 (N7563, N7558, N5995, N2423, N1655);
xor XOR2 (N7564, N7554, N1146);
or OR3 (N7565, N7562, N1414, N5218);
nor NOR2 (N7566, N7547, N1191);
not NOT1 (N7567, N7565);
nand NAND2 (N7568, N7560, N3804);
buf BUF1 (N7569, N7564);
xor XOR2 (N7570, N7563, N369);
and AND4 (N7571, N7552, N2445, N5953, N2057);
xor XOR2 (N7572, N7557, N2481);
xor XOR2 (N7573, N7566, N3584);
nand NAND2 (N7574, N7573, N1717);
not NOT1 (N7575, N7525);
and AND4 (N7576, N7575, N4460, N2865, N538);
and AND3 (N7577, N7574, N1548, N39);
nand NAND3 (N7578, N7571, N2301, N1971);
nand NAND4 (N7579, N7569, N2150, N468, N3532);
nand NAND4 (N7580, N7576, N729, N3685, N2623);
nor NOR3 (N7581, N7570, N6651, N7579);
and AND4 (N7582, N5728, N3941, N1594, N6964);
or OR4 (N7583, N7582, N3784, N529, N4809);
not NOT1 (N7584, N7581);
xor XOR2 (N7585, N7559, N432);
or OR2 (N7586, N7577, N4812);
nor NOR3 (N7587, N7583, N6926, N3538);
nor NOR4 (N7588, N7587, N6209, N1645, N3468);
nor NOR2 (N7589, N7567, N4360);
and AND2 (N7590, N7588, N4698);
nor NOR4 (N7591, N7568, N4864, N3792, N3591);
buf BUF1 (N7592, N7586);
or OR3 (N7593, N7592, N71, N6775);
xor XOR2 (N7594, N7572, N7401);
not NOT1 (N7595, N7589);
and AND3 (N7596, N7594, N362, N6320);
buf BUF1 (N7597, N7593);
or OR4 (N7598, N7591, N719, N5708, N4961);
buf BUF1 (N7599, N7598);
buf BUF1 (N7600, N7584);
not NOT1 (N7601, N7600);
and AND2 (N7602, N7580, N1497);
xor XOR2 (N7603, N7596, N4005);
not NOT1 (N7604, N7595);
xor XOR2 (N7605, N7555, N7050);
buf BUF1 (N7606, N7603);
nand NAND4 (N7607, N7585, N2624, N4673, N339);
buf BUF1 (N7608, N7590);
buf BUF1 (N7609, N7607);
nor NOR3 (N7610, N7608, N5026, N1547);
and AND2 (N7611, N7609, N6432);
not NOT1 (N7612, N7578);
xor XOR2 (N7613, N7605, N2218);
not NOT1 (N7614, N7602);
nor NOR3 (N7615, N7613, N808, N4657);
or OR2 (N7616, N7615, N4302);
nor NOR4 (N7617, N7610, N4348, N4477, N7312);
nor NOR2 (N7618, N7614, N6222);
not NOT1 (N7619, N7597);
nand NAND4 (N7620, N7617, N7156, N2456, N637);
and AND4 (N7621, N7606, N6167, N6497, N6991);
and AND2 (N7622, N7616, N1565);
and AND3 (N7623, N7612, N3342, N7381);
or OR2 (N7624, N7623, N3970);
nand NAND4 (N7625, N7599, N3751, N1403, N958);
or OR2 (N7626, N7622, N3467);
xor XOR2 (N7627, N7618, N1477);
or OR3 (N7628, N7620, N2559, N7185);
buf BUF1 (N7629, N7611);
not NOT1 (N7630, N7626);
nand NAND4 (N7631, N7625, N7354, N7055, N1970);
buf BUF1 (N7632, N7629);
and AND4 (N7633, N7628, N3883, N2112, N5064);
nand NAND2 (N7634, N7619, N1774);
buf BUF1 (N7635, N7634);
xor XOR2 (N7636, N7632, N2004);
xor XOR2 (N7637, N7631, N241);
nor NOR3 (N7638, N7624, N1592, N6263);
nand NAND2 (N7639, N7636, N408);
and AND4 (N7640, N7601, N1595, N7384, N1388);
nor NOR3 (N7641, N7627, N2930, N4534);
buf BUF1 (N7642, N7640);
and AND4 (N7643, N7630, N3102, N4930, N6358);
not NOT1 (N7644, N7635);
nor NOR2 (N7645, N7644, N485);
and AND4 (N7646, N7639, N7213, N72, N1299);
xor XOR2 (N7647, N7641, N1575);
nor NOR4 (N7648, N7621, N307, N7019, N2386);
nor NOR4 (N7649, N7638, N1338, N319, N2059);
xor XOR2 (N7650, N7643, N488);
buf BUF1 (N7651, N7650);
not NOT1 (N7652, N7604);
or OR4 (N7653, N7648, N5008, N1502, N3302);
nor NOR2 (N7654, N7633, N543);
xor XOR2 (N7655, N7642, N2387);
or OR3 (N7656, N7645, N2632, N4006);
nor NOR3 (N7657, N7653, N2431, N1047);
not NOT1 (N7658, N7646);
or OR2 (N7659, N7637, N3885);
or OR3 (N7660, N7647, N4339, N4798);
nand NAND3 (N7661, N7658, N5024, N5758);
and AND2 (N7662, N7660, N7270);
xor XOR2 (N7663, N7656, N6156);
not NOT1 (N7664, N7657);
and AND2 (N7665, N7659, N437);
buf BUF1 (N7666, N7661);
nand NAND3 (N7667, N7651, N4661, N2925);
buf BUF1 (N7668, N7649);
nand NAND3 (N7669, N7655, N6036, N6178);
not NOT1 (N7670, N7664);
xor XOR2 (N7671, N7652, N3104);
nand NAND2 (N7672, N7669, N3990);
xor XOR2 (N7673, N7670, N929);
and AND4 (N7674, N7663, N893, N4213, N356);
not NOT1 (N7675, N7672);
nor NOR2 (N7676, N7668, N4743);
nor NOR2 (N7677, N7676, N7466);
xor XOR2 (N7678, N7662, N1961);
not NOT1 (N7679, N7667);
and AND3 (N7680, N7674, N2146, N3535);
not NOT1 (N7681, N7666);
not NOT1 (N7682, N7665);
nand NAND2 (N7683, N7671, N6359);
nand NAND3 (N7684, N7683, N2013, N5729);
nand NAND4 (N7685, N7684, N5, N5051, N1731);
not NOT1 (N7686, N7685);
and AND4 (N7687, N7654, N57, N6128, N5818);
buf BUF1 (N7688, N7682);
xor XOR2 (N7689, N7677, N5444);
or OR4 (N7690, N7679, N2680, N908, N3095);
xor XOR2 (N7691, N7675, N3417);
xor XOR2 (N7692, N7673, N1692);
or OR4 (N7693, N7688, N162, N1420, N4146);
not NOT1 (N7694, N7687);
nor NOR4 (N7695, N7678, N4018, N3876, N1204);
not NOT1 (N7696, N7695);
or OR2 (N7697, N7686, N4424);
xor XOR2 (N7698, N7689, N5812);
nand NAND2 (N7699, N7681, N359);
and AND4 (N7700, N7694, N3109, N1932, N1849);
and AND3 (N7701, N7699, N1194, N7063);
and AND4 (N7702, N7691, N371, N2593, N1633);
buf BUF1 (N7703, N7696);
and AND4 (N7704, N7703, N2582, N7212, N7174);
xor XOR2 (N7705, N7698, N6842);
buf BUF1 (N7706, N7702);
nor NOR4 (N7707, N7697, N4727, N115, N1179);
nand NAND3 (N7708, N7693, N5354, N3691);
nor NOR2 (N7709, N7706, N3200);
nor NOR3 (N7710, N7690, N3460, N857);
not NOT1 (N7711, N7709);
and AND4 (N7712, N7705, N2210, N5106, N1298);
and AND3 (N7713, N7700, N4639, N2328);
nand NAND4 (N7714, N7701, N6672, N3223, N3262);
nor NOR2 (N7715, N7707, N7526);
buf BUF1 (N7716, N7714);
nor NOR4 (N7717, N7704, N2973, N2747, N140);
and AND4 (N7718, N7680, N6433, N6915, N2020);
and AND3 (N7719, N7692, N1846, N155);
or OR2 (N7720, N7718, N314);
xor XOR2 (N7721, N7719, N4048);
nand NAND4 (N7722, N7708, N6030, N7447, N4576);
not NOT1 (N7723, N7712);
nor NOR4 (N7724, N7722, N698, N2305, N1238);
xor XOR2 (N7725, N7723, N7030);
nand NAND3 (N7726, N7715, N1001, N249);
xor XOR2 (N7727, N7724, N2660);
nand NAND2 (N7728, N7721, N4173);
and AND2 (N7729, N7717, N5748);
or OR4 (N7730, N7720, N7228, N2328, N5866);
nor NOR2 (N7731, N7729, N3518);
nand NAND3 (N7732, N7716, N6188, N5784);
xor XOR2 (N7733, N7726, N7425);
nand NAND2 (N7734, N7733, N4692);
and AND2 (N7735, N7710, N1390);
not NOT1 (N7736, N7711);
nand NAND3 (N7737, N7730, N1532, N205);
buf BUF1 (N7738, N7736);
or OR3 (N7739, N7725, N2717, N5964);
nor NOR4 (N7740, N7738, N2387, N5041, N7135);
not NOT1 (N7741, N7739);
nand NAND3 (N7742, N7734, N7394, N540);
nor NOR3 (N7743, N7732, N5502, N5574);
or OR3 (N7744, N7742, N6127, N1291);
buf BUF1 (N7745, N7713);
or OR4 (N7746, N7727, N5184, N3662, N6408);
nor NOR4 (N7747, N7746, N685, N4530, N3981);
xor XOR2 (N7748, N7731, N7129);
buf BUF1 (N7749, N7745);
buf BUF1 (N7750, N7737);
not NOT1 (N7751, N7735);
and AND4 (N7752, N7744, N184, N1274, N5275);
or OR3 (N7753, N7741, N3027, N2170);
buf BUF1 (N7754, N7750);
nor NOR2 (N7755, N7743, N1673);
nand NAND3 (N7756, N7752, N7415, N663);
buf BUF1 (N7757, N7756);
xor XOR2 (N7758, N7755, N4638);
not NOT1 (N7759, N7757);
xor XOR2 (N7760, N7753, N4996);
xor XOR2 (N7761, N7760, N370);
buf BUF1 (N7762, N7759);
xor XOR2 (N7763, N7728, N2144);
xor XOR2 (N7764, N7751, N7244);
xor XOR2 (N7765, N7754, N5009);
buf BUF1 (N7766, N7749);
buf BUF1 (N7767, N7747);
nor NOR4 (N7768, N7763, N294, N1903, N2237);
or OR4 (N7769, N7758, N3383, N452, N6570);
not NOT1 (N7770, N7740);
and AND3 (N7771, N7768, N6015, N761);
and AND3 (N7772, N7771, N1538, N4159);
xor XOR2 (N7773, N7766, N3376);
and AND2 (N7774, N7765, N5644);
nor NOR2 (N7775, N7770, N1939);
and AND2 (N7776, N7748, N4528);
and AND2 (N7777, N7761, N1164);
buf BUF1 (N7778, N7764);
or OR2 (N7779, N7776, N5909);
nand NAND2 (N7780, N7773, N1031);
buf BUF1 (N7781, N7777);
nor NOR2 (N7782, N7772, N3353);
nor NOR2 (N7783, N7779, N2449);
buf BUF1 (N7784, N7782);
xor XOR2 (N7785, N7762, N3599);
and AND3 (N7786, N7780, N3308, N1029);
nor NOR3 (N7787, N7769, N6621, N7714);
nor NOR4 (N7788, N7783, N4841, N1415, N1651);
or OR2 (N7789, N7774, N5503);
not NOT1 (N7790, N7784);
buf BUF1 (N7791, N7781);
or OR4 (N7792, N7787, N7166, N2238, N4619);
not NOT1 (N7793, N7788);
and AND4 (N7794, N7792, N3819, N334, N3180);
or OR2 (N7795, N7767, N4451);
nor NOR4 (N7796, N7794, N5422, N5738, N4892);
nand NAND3 (N7797, N7790, N6458, N7483);
or OR4 (N7798, N7793, N3757, N2292, N5341);
buf BUF1 (N7799, N7797);
nor NOR4 (N7800, N7778, N5260, N7078, N3926);
buf BUF1 (N7801, N7789);
or OR2 (N7802, N7798, N7782);
or OR4 (N7803, N7785, N7169, N5850, N2736);
and AND2 (N7804, N7800, N7758);
xor XOR2 (N7805, N7795, N4695);
nor NOR4 (N7806, N7803, N5146, N4295, N1473);
buf BUF1 (N7807, N7804);
xor XOR2 (N7808, N7791, N2652);
and AND2 (N7809, N7805, N4368);
or OR2 (N7810, N7801, N5267);
and AND4 (N7811, N7799, N757, N1374, N7677);
nand NAND4 (N7812, N7810, N5148, N163, N270);
buf BUF1 (N7813, N7809);
or OR3 (N7814, N7811, N6900, N2073);
xor XOR2 (N7815, N7812, N847);
nor NOR2 (N7816, N7808, N2326);
buf BUF1 (N7817, N7802);
buf BUF1 (N7818, N7807);
nand NAND3 (N7819, N7815, N5217, N6727);
not NOT1 (N7820, N7814);
or OR2 (N7821, N7796, N2374);
buf BUF1 (N7822, N7818);
buf BUF1 (N7823, N7775);
not NOT1 (N7824, N7813);
or OR3 (N7825, N7816, N264, N5928);
and AND4 (N7826, N7786, N5699, N2256, N2942);
or OR4 (N7827, N7826, N6070, N6696, N7242);
not NOT1 (N7828, N7819);
buf BUF1 (N7829, N7822);
xor XOR2 (N7830, N7821, N56);
and AND4 (N7831, N7820, N6908, N1335, N2026);
or OR4 (N7832, N7817, N4186, N366, N972);
buf BUF1 (N7833, N7830);
or OR4 (N7834, N7828, N715, N1439, N652);
xor XOR2 (N7835, N7829, N2370);
nand NAND4 (N7836, N7831, N2465, N6388, N6332);
nand NAND4 (N7837, N7835, N6240, N3216, N5958);
or OR2 (N7838, N7824, N5386);
or OR4 (N7839, N7806, N4334, N3018, N397);
xor XOR2 (N7840, N7836, N6821);
nor NOR4 (N7841, N7834, N641, N5858, N1660);
nand NAND3 (N7842, N7841, N4111, N855);
nand NAND3 (N7843, N7838, N600, N4370);
xor XOR2 (N7844, N7823, N3382);
and AND4 (N7845, N7825, N1150, N2209, N1020);
buf BUF1 (N7846, N7845);
or OR2 (N7847, N7839, N676);
nor NOR4 (N7848, N7837, N511, N4844, N956);
nor NOR3 (N7849, N7833, N5092, N1253);
not NOT1 (N7850, N7847);
xor XOR2 (N7851, N7827, N5206);
xor XOR2 (N7852, N7843, N7252);
and AND4 (N7853, N7849, N3246, N1672, N6934);
xor XOR2 (N7854, N7852, N2899);
not NOT1 (N7855, N7850);
buf BUF1 (N7856, N7853);
and AND3 (N7857, N7846, N5607, N4067);
not NOT1 (N7858, N7840);
not NOT1 (N7859, N7844);
or OR4 (N7860, N7859, N4324, N2110, N91);
buf BUF1 (N7861, N7856);
nor NOR3 (N7862, N7848, N4948, N1843);
or OR4 (N7863, N7851, N4145, N5683, N6172);
buf BUF1 (N7864, N7863);
or OR4 (N7865, N7864, N6095, N955, N5189);
buf BUF1 (N7866, N7855);
not NOT1 (N7867, N7861);
nor NOR2 (N7868, N7860, N3425);
not NOT1 (N7869, N7857);
nand NAND4 (N7870, N7868, N6178, N2075, N4127);
buf BUF1 (N7871, N7865);
not NOT1 (N7872, N7871);
buf BUF1 (N7873, N7872);
xor XOR2 (N7874, N7870, N4162);
buf BUF1 (N7875, N7862);
and AND3 (N7876, N7874, N3463, N3514);
nor NOR2 (N7877, N7875, N5913);
nand NAND4 (N7878, N7854, N5859, N6257, N3838);
xor XOR2 (N7879, N7873, N5554);
or OR3 (N7880, N7867, N6228, N856);
nor NOR2 (N7881, N7877, N45);
or OR3 (N7882, N7866, N1654, N4046);
not NOT1 (N7883, N7876);
nand NAND3 (N7884, N7882, N1556, N1402);
not NOT1 (N7885, N7858);
nor NOR2 (N7886, N7880, N3090);
nand NAND3 (N7887, N7884, N315, N6920);
and AND4 (N7888, N7885, N3786, N720, N7515);
xor XOR2 (N7889, N7842, N2754);
buf BUF1 (N7890, N7881);
or OR3 (N7891, N7878, N5591, N7375);
xor XOR2 (N7892, N7888, N7315);
nor NOR3 (N7893, N7832, N3184, N3172);
xor XOR2 (N7894, N7891, N2938);
not NOT1 (N7895, N7869);
nor NOR3 (N7896, N7892, N4502, N1499);
or OR4 (N7897, N7889, N1174, N4114, N3005);
nor NOR3 (N7898, N7895, N37, N7247);
and AND4 (N7899, N7890, N4947, N533, N2550);
or OR2 (N7900, N7898, N3174);
nand NAND2 (N7901, N7896, N4776);
not NOT1 (N7902, N7893);
buf BUF1 (N7903, N7900);
buf BUF1 (N7904, N7883);
buf BUF1 (N7905, N7903);
nand NAND4 (N7906, N7887, N2336, N893, N3970);
and AND3 (N7907, N7879, N6392, N7368);
xor XOR2 (N7908, N7905, N6106);
buf BUF1 (N7909, N7897);
not NOT1 (N7910, N7907);
nand NAND3 (N7911, N7908, N3179, N63);
and AND2 (N7912, N7886, N3209);
nand NAND4 (N7913, N7910, N3707, N4083, N4816);
buf BUF1 (N7914, N7906);
not NOT1 (N7915, N7901);
or OR4 (N7916, N7902, N2791, N5824, N6555);
and AND2 (N7917, N7912, N7275);
nand NAND3 (N7918, N7914, N4358, N6076);
not NOT1 (N7919, N7894);
not NOT1 (N7920, N7918);
xor XOR2 (N7921, N7904, N2452);
nor NOR3 (N7922, N7916, N3011, N713);
xor XOR2 (N7923, N7913, N970);
and AND3 (N7924, N7920, N2733, N3762);
xor XOR2 (N7925, N7909, N6868);
nor NOR3 (N7926, N7915, N7561, N4490);
nor NOR3 (N7927, N7926, N1372, N7228);
xor XOR2 (N7928, N7921, N7041);
buf BUF1 (N7929, N7919);
buf BUF1 (N7930, N7924);
nand NAND2 (N7931, N7922, N1099);
xor XOR2 (N7932, N7928, N6346);
nor NOR3 (N7933, N7931, N5374, N5885);
or OR4 (N7934, N7923, N3962, N3486, N665);
or OR3 (N7935, N7925, N6897, N7355);
and AND4 (N7936, N7927, N800, N3167, N1702);
not NOT1 (N7937, N7929);
nor NOR2 (N7938, N7917, N5037);
xor XOR2 (N7939, N7930, N4263);
and AND2 (N7940, N7911, N5725);
and AND3 (N7941, N7936, N1027, N2728);
and AND4 (N7942, N7941, N7919, N410, N6725);
or OR2 (N7943, N7942, N7770);
and AND4 (N7944, N7934, N6295, N5570, N4492);
nor NOR3 (N7945, N7943, N6799, N3704);
and AND2 (N7946, N7944, N1297);
or OR3 (N7947, N7935, N5165, N190);
nor NOR4 (N7948, N7946, N3514, N7037, N7400);
xor XOR2 (N7949, N7947, N6623);
xor XOR2 (N7950, N7938, N4996);
or OR4 (N7951, N7937, N7561, N5744, N3132);
and AND2 (N7952, N7948, N6947);
nor NOR3 (N7953, N7940, N511, N5660);
not NOT1 (N7954, N7939);
nand NAND3 (N7955, N7954, N4427, N7072);
nor NOR3 (N7956, N7953, N188, N4371);
xor XOR2 (N7957, N7955, N3900);
or OR3 (N7958, N7957, N1846, N3849);
buf BUF1 (N7959, N7949);
and AND4 (N7960, N7952, N1330, N476, N5010);
nand NAND2 (N7961, N7959, N1967);
nand NAND4 (N7962, N7956, N5183, N3925, N4059);
or OR4 (N7963, N7950, N3019, N782, N4304);
and AND2 (N7964, N7962, N3112);
xor XOR2 (N7965, N7960, N7869);
nor NOR2 (N7966, N7932, N3337);
nor NOR2 (N7967, N7961, N1257);
nand NAND3 (N7968, N7966, N1362, N4808);
and AND2 (N7969, N7899, N6553);
nand NAND3 (N7970, N7951, N6684, N1908);
or OR3 (N7971, N7945, N2954, N7175);
xor XOR2 (N7972, N7964, N6968);
and AND3 (N7973, N7968, N6869, N2611);
or OR4 (N7974, N7972, N3133, N1101, N5431);
and AND2 (N7975, N7971, N4260);
xor XOR2 (N7976, N7933, N424);
xor XOR2 (N7977, N7974, N4321);
not NOT1 (N7978, N7976);
or OR3 (N7979, N7967, N3646, N5171);
nor NOR2 (N7980, N7979, N5428);
and AND4 (N7981, N7980, N1430, N2625, N226);
xor XOR2 (N7982, N7963, N2769);
and AND3 (N7983, N7977, N5803, N7402);
or OR2 (N7984, N7983, N4448);
not NOT1 (N7985, N7965);
buf BUF1 (N7986, N7982);
not NOT1 (N7987, N7958);
nand NAND3 (N7988, N7970, N5115, N3657);
buf BUF1 (N7989, N7975);
nand NAND4 (N7990, N7978, N2583, N3611, N1822);
buf BUF1 (N7991, N7989);
buf BUF1 (N7992, N7987);
and AND4 (N7993, N7991, N5108, N2716, N4678);
nand NAND4 (N7994, N7986, N2533, N4314, N6388);
and AND3 (N7995, N7973, N3933, N7865);
not NOT1 (N7996, N7990);
xor XOR2 (N7997, N7985, N5767);
nor NOR4 (N7998, N7988, N4412, N7409, N1720);
buf BUF1 (N7999, N7994);
buf BUF1 (N8000, N7996);
xor XOR2 (N8001, N7999, N634);
and AND2 (N8002, N7969, N6784);
nor NOR4 (N8003, N7997, N1833, N6112, N1785);
buf BUF1 (N8004, N8000);
nand NAND2 (N8005, N7993, N5945);
nand NAND4 (N8006, N7984, N1471, N6523, N7290);
and AND2 (N8007, N8006, N3944);
or OR4 (N8008, N7981, N958, N5274, N5366);
or OR4 (N8009, N8003, N259, N493, N1183);
not NOT1 (N8010, N8005);
buf BUF1 (N8011, N7995);
nand NAND3 (N8012, N8008, N4358, N1796);
nand NAND2 (N8013, N7992, N7445);
not NOT1 (N8014, N8001);
xor XOR2 (N8015, N8014, N7431);
buf BUF1 (N8016, N8015);
nor NOR4 (N8017, N8007, N5941, N5126, N2350);
nand NAND4 (N8018, N8009, N7116, N7861, N7198);
and AND2 (N8019, N8004, N5798);
and AND4 (N8020, N8017, N740, N661, N2055);
nor NOR4 (N8021, N8010, N7016, N7666, N6028);
not NOT1 (N8022, N8011);
xor XOR2 (N8023, N8019, N7602);
and AND4 (N8024, N8020, N2589, N4833, N2681);
not NOT1 (N8025, N8016);
nand NAND4 (N8026, N8021, N3650, N1851, N2425);
nor NOR4 (N8027, N8026, N4931, N3171, N6162);
buf BUF1 (N8028, N7998);
buf BUF1 (N8029, N8027);
nor NOR2 (N8030, N8012, N4403);
nand NAND3 (N8031, N8022, N4612, N1634);
and AND2 (N8032, N8028, N3622);
nand NAND2 (N8033, N8032, N3599);
and AND3 (N8034, N8002, N318, N7167);
buf BUF1 (N8035, N8024);
nand NAND2 (N8036, N8018, N4609);
and AND2 (N8037, N8029, N5424);
or OR2 (N8038, N8037, N5455);
not NOT1 (N8039, N8025);
buf BUF1 (N8040, N8013);
not NOT1 (N8041, N8030);
or OR3 (N8042, N8040, N7984, N300);
not NOT1 (N8043, N8034);
and AND3 (N8044, N8041, N7741, N6270);
or OR2 (N8045, N8042, N7613);
not NOT1 (N8046, N8035);
buf BUF1 (N8047, N8044);
nor NOR3 (N8048, N8045, N2426, N3437);
and AND4 (N8049, N8048, N1297, N364, N3872);
nor NOR2 (N8050, N8039, N6999);
xor XOR2 (N8051, N8038, N3281);
nand NAND2 (N8052, N8050, N5727);
nor NOR4 (N8053, N8046, N2299, N448, N4498);
xor XOR2 (N8054, N8053, N5828);
or OR4 (N8055, N8054, N2894, N5744, N7159);
or OR3 (N8056, N8043, N3763, N5976);
not NOT1 (N8057, N8023);
not NOT1 (N8058, N8057);
and AND2 (N8059, N8033, N4388);
or OR3 (N8060, N8056, N3773, N7006);
and AND3 (N8061, N8060, N5314, N474);
and AND2 (N8062, N8055, N4277);
buf BUF1 (N8063, N8031);
or OR3 (N8064, N8059, N7821, N4360);
or OR3 (N8065, N8061, N5597, N1301);
xor XOR2 (N8066, N8052, N3381);
nand NAND4 (N8067, N8066, N7593, N2958, N6682);
not NOT1 (N8068, N8051);
buf BUF1 (N8069, N8036);
not NOT1 (N8070, N8067);
or OR3 (N8071, N8064, N4101, N4235);
buf BUF1 (N8072, N8047);
nor NOR4 (N8073, N8069, N5577, N1218, N3034);
not NOT1 (N8074, N8072);
nand NAND2 (N8075, N8071, N76);
xor XOR2 (N8076, N8070, N930);
or OR3 (N8077, N8075, N7946, N1098);
buf BUF1 (N8078, N8062);
nor NOR4 (N8079, N8076, N571, N8056, N6259);
xor XOR2 (N8080, N8049, N7946);
xor XOR2 (N8081, N8079, N3615);
not NOT1 (N8082, N8063);
xor XOR2 (N8083, N8073, N3960);
buf BUF1 (N8084, N8080);
not NOT1 (N8085, N8083);
buf BUF1 (N8086, N8084);
buf BUF1 (N8087, N8081);
xor XOR2 (N8088, N8078, N3478);
or OR2 (N8089, N8087, N5851);
nor NOR2 (N8090, N8068, N4269);
nand NAND3 (N8091, N8088, N4908, N778);
or OR4 (N8092, N8089, N3020, N7706, N7441);
nand NAND4 (N8093, N8085, N6439, N2179, N1606);
xor XOR2 (N8094, N8074, N5932);
nand NAND4 (N8095, N8092, N460, N953, N2423);
nand NAND2 (N8096, N8094, N6686);
nand NAND3 (N8097, N8082, N3523, N6597);
xor XOR2 (N8098, N8065, N2386);
buf BUF1 (N8099, N8058);
nor NOR4 (N8100, N8090, N1674, N2607, N3231);
xor XOR2 (N8101, N8091, N522);
or OR3 (N8102, N8097, N5606, N6184);
nor NOR4 (N8103, N8101, N6797, N881, N506);
not NOT1 (N8104, N8093);
nand NAND2 (N8105, N8102, N5493);
xor XOR2 (N8106, N8105, N1236);
buf BUF1 (N8107, N8077);
xor XOR2 (N8108, N8098, N1100);
xor XOR2 (N8109, N8086, N4823);
not NOT1 (N8110, N8108);
not NOT1 (N8111, N8099);
xor XOR2 (N8112, N8107, N1733);
nor NOR2 (N8113, N8095, N6739);
buf BUF1 (N8114, N8100);
xor XOR2 (N8115, N8109, N172);
and AND2 (N8116, N8104, N6607);
not NOT1 (N8117, N8114);
buf BUF1 (N8118, N8110);
nand NAND3 (N8119, N8116, N2155, N7086);
nor NOR4 (N8120, N8096, N2325, N5434, N8098);
nand NAND4 (N8121, N8120, N5887, N8049, N1943);
and AND4 (N8122, N8103, N1863, N1795, N7308);
nor NOR3 (N8123, N8117, N6509, N3400);
nand NAND4 (N8124, N8118, N16, N375, N6084);
and AND4 (N8125, N8111, N4120, N3005, N4445);
or OR2 (N8126, N8124, N4602);
nor NOR3 (N8127, N8106, N4284, N3606);
or OR3 (N8128, N8126, N3122, N2689);
or OR2 (N8129, N8128, N198);
nor NOR2 (N8130, N8112, N6819);
nor NOR4 (N8131, N8115, N1475, N5949, N6865);
buf BUF1 (N8132, N8121);
or OR4 (N8133, N8123, N7553, N4039, N6027);
nor NOR3 (N8134, N8125, N6618, N2608);
buf BUF1 (N8135, N8131);
xor XOR2 (N8136, N8132, N4213);
buf BUF1 (N8137, N8119);
buf BUF1 (N8138, N8113);
nor NOR4 (N8139, N8129, N5344, N1905, N2609);
xor XOR2 (N8140, N8135, N2460);
buf BUF1 (N8141, N8136);
nor NOR3 (N8142, N8140, N1243, N6894);
nor NOR3 (N8143, N8127, N5267, N51);
not NOT1 (N8144, N8130);
nand NAND3 (N8145, N8141, N5499, N1672);
or OR3 (N8146, N8133, N7709, N3163);
not NOT1 (N8147, N8146);
buf BUF1 (N8148, N8137);
not NOT1 (N8149, N8138);
buf BUF1 (N8150, N8122);
xor XOR2 (N8151, N8134, N6869);
and AND2 (N8152, N8150, N3175);
nor NOR3 (N8153, N8145, N6044, N4277);
buf BUF1 (N8154, N8139);
nor NOR4 (N8155, N8142, N6819, N2746, N4535);
buf BUF1 (N8156, N8148);
not NOT1 (N8157, N8147);
nor NOR2 (N8158, N8143, N7780);
or OR2 (N8159, N8154, N5);
or OR2 (N8160, N8144, N7721);
nor NOR4 (N8161, N8151, N3692, N2607, N3990);
buf BUF1 (N8162, N8159);
buf BUF1 (N8163, N8155);
nand NAND3 (N8164, N8153, N5393, N769);
or OR2 (N8165, N8163, N4729);
xor XOR2 (N8166, N8160, N7860);
and AND2 (N8167, N8152, N4900);
not NOT1 (N8168, N8149);
nor NOR2 (N8169, N8167, N3332);
nand NAND3 (N8170, N8161, N163, N4723);
nor NOR2 (N8171, N8156, N527);
buf BUF1 (N8172, N8169);
nor NOR4 (N8173, N8170, N2878, N4253, N1152);
not NOT1 (N8174, N8172);
xor XOR2 (N8175, N8171, N5041);
xor XOR2 (N8176, N8175, N2104);
xor XOR2 (N8177, N8174, N5685);
nor NOR4 (N8178, N8177, N8176, N7914, N6786);
nand NAND4 (N8179, N79, N2091, N5459, N1486);
nor NOR2 (N8180, N8165, N6522);
nor NOR3 (N8181, N8173, N7502, N80);
nor NOR3 (N8182, N8157, N1526, N7626);
xor XOR2 (N8183, N8166, N1585);
nor NOR3 (N8184, N8183, N5961, N7695);
or OR3 (N8185, N8178, N2005, N6347);
or OR2 (N8186, N8168, N5827);
xor XOR2 (N8187, N8179, N721);
nor NOR4 (N8188, N8182, N7659, N7093, N6518);
buf BUF1 (N8189, N8181);
buf BUF1 (N8190, N8162);
buf BUF1 (N8191, N8186);
and AND4 (N8192, N8189, N3665, N5791, N4137);
not NOT1 (N8193, N8192);
or OR4 (N8194, N8184, N2745, N4343, N7159);
nand NAND2 (N8195, N8193, N4562);
or OR2 (N8196, N8187, N6684);
or OR2 (N8197, N8195, N2513);
buf BUF1 (N8198, N8191);
nor NOR3 (N8199, N8158, N1642, N2815);
nor NOR2 (N8200, N8197, N3269);
nand NAND4 (N8201, N8199, N4987, N1044, N6787);
not NOT1 (N8202, N8194);
xor XOR2 (N8203, N8188, N3003);
xor XOR2 (N8204, N8180, N5914);
not NOT1 (N8205, N8203);
nor NOR4 (N8206, N8204, N2026, N6233, N4928);
xor XOR2 (N8207, N8200, N1311);
or OR4 (N8208, N8201, N6324, N3845, N5731);
nor NOR2 (N8209, N8190, N1098);
nor NOR2 (N8210, N8164, N1542);
or OR2 (N8211, N8185, N1998);
not NOT1 (N8212, N8205);
not NOT1 (N8213, N8212);
buf BUF1 (N8214, N8213);
not NOT1 (N8215, N8202);
not NOT1 (N8216, N8206);
not NOT1 (N8217, N8209);
xor XOR2 (N8218, N8210, N5981);
buf BUF1 (N8219, N8208);
or OR2 (N8220, N8196, N5798);
not NOT1 (N8221, N8215);
and AND2 (N8222, N8207, N7537);
xor XOR2 (N8223, N8198, N4393);
nor NOR3 (N8224, N8211, N7105, N8104);
and AND2 (N8225, N8224, N2662);
not NOT1 (N8226, N8220);
nand NAND3 (N8227, N8221, N3367, N4092);
buf BUF1 (N8228, N8219);
and AND2 (N8229, N8216, N4835);
nor NOR4 (N8230, N8217, N1791, N1558, N2121);
nand NAND4 (N8231, N8222, N2031, N4628, N6917);
nand NAND2 (N8232, N8214, N4297);
nand NAND4 (N8233, N8231, N1468, N3028, N3415);
buf BUF1 (N8234, N8227);
not NOT1 (N8235, N8225);
not NOT1 (N8236, N8230);
buf BUF1 (N8237, N8226);
buf BUF1 (N8238, N8229);
nor NOR2 (N8239, N8234, N4069);
buf BUF1 (N8240, N8237);
nand NAND2 (N8241, N8233, N7412);
not NOT1 (N8242, N8241);
nand NAND2 (N8243, N8235, N6593);
buf BUF1 (N8244, N8236);
not NOT1 (N8245, N8239);
nor NOR4 (N8246, N8218, N4175, N7243, N4328);
not NOT1 (N8247, N8228);
xor XOR2 (N8248, N8232, N695);
or OR3 (N8249, N8223, N6819, N7468);
buf BUF1 (N8250, N8244);
buf BUF1 (N8251, N8249);
and AND4 (N8252, N8238, N2392, N6976, N6341);
nor NOR2 (N8253, N8242, N398);
or OR3 (N8254, N8248, N3270, N7040);
nor NOR4 (N8255, N8243, N4367, N7899, N4721);
and AND4 (N8256, N8253, N4566, N7873, N4009);
or OR4 (N8257, N8250, N2421, N2363, N2937);
not NOT1 (N8258, N8256);
and AND2 (N8259, N8258, N1548);
buf BUF1 (N8260, N8246);
not NOT1 (N8261, N8245);
and AND4 (N8262, N8257, N7060, N2324, N3458);
nor NOR4 (N8263, N8252, N6056, N5130, N3604);
and AND4 (N8264, N8255, N2166, N7407, N4034);
nor NOR3 (N8265, N8247, N806, N3765);
nor NOR4 (N8266, N8260, N1079, N1965, N2809);
buf BUF1 (N8267, N8263);
or OR2 (N8268, N8254, N5009);
or OR4 (N8269, N8261, N1138, N4867, N7171);
or OR4 (N8270, N8267, N4149, N3324, N357);
nand NAND2 (N8271, N8269, N1097);
nor NOR4 (N8272, N8259, N6413, N341, N2195);
not NOT1 (N8273, N8268);
or OR4 (N8274, N8273, N1205, N6641, N6135);
or OR3 (N8275, N8270, N564, N2301);
not NOT1 (N8276, N8275);
buf BUF1 (N8277, N8262);
and AND2 (N8278, N8251, N5808);
xor XOR2 (N8279, N8266, N804);
buf BUF1 (N8280, N8276);
not NOT1 (N8281, N8278);
or OR4 (N8282, N8281, N49, N5317, N6446);
xor XOR2 (N8283, N8277, N5939);
not NOT1 (N8284, N8283);
not NOT1 (N8285, N8240);
nand NAND4 (N8286, N8274, N5937, N5964, N5384);
and AND2 (N8287, N8286, N5254);
xor XOR2 (N8288, N8279, N6771);
or OR2 (N8289, N8272, N2071);
buf BUF1 (N8290, N8264);
not NOT1 (N8291, N8287);
xor XOR2 (N8292, N8290, N2674);
buf BUF1 (N8293, N8291);
not NOT1 (N8294, N8280);
buf BUF1 (N8295, N8284);
buf BUF1 (N8296, N8265);
xor XOR2 (N8297, N8288, N1596);
nand NAND3 (N8298, N8285, N6366, N3078);
nand NAND2 (N8299, N8271, N4516);
or OR4 (N8300, N8296, N3430, N4436, N7820);
not NOT1 (N8301, N8293);
nand NAND4 (N8302, N8299, N6635, N5946, N1366);
xor XOR2 (N8303, N8289, N6055);
not NOT1 (N8304, N8294);
xor XOR2 (N8305, N8292, N6276);
and AND3 (N8306, N8304, N1440, N5014);
xor XOR2 (N8307, N8298, N4996);
not NOT1 (N8308, N8300);
buf BUF1 (N8309, N8302);
buf BUF1 (N8310, N8307);
buf BUF1 (N8311, N8306);
nor NOR4 (N8312, N8295, N6706, N7262, N6005);
buf BUF1 (N8313, N8312);
or OR3 (N8314, N8297, N5762, N3198);
or OR4 (N8315, N8309, N347, N3586, N5212);
xor XOR2 (N8316, N8311, N8221);
nor NOR2 (N8317, N8316, N4795);
not NOT1 (N8318, N8315);
not NOT1 (N8319, N8303);
not NOT1 (N8320, N8314);
xor XOR2 (N8321, N8313, N2984);
nand NAND3 (N8322, N8318, N1575, N8293);
and AND2 (N8323, N8305, N7318);
not NOT1 (N8324, N8282);
and AND4 (N8325, N8324, N3650, N2084, N7522);
xor XOR2 (N8326, N8323, N1045);
xor XOR2 (N8327, N8326, N2251);
xor XOR2 (N8328, N8320, N2568);
buf BUF1 (N8329, N8317);
and AND4 (N8330, N8329, N1726, N1683, N7196);
not NOT1 (N8331, N8308);
and AND3 (N8332, N8319, N7668, N5025);
and AND2 (N8333, N8330, N5783);
buf BUF1 (N8334, N8322);
not NOT1 (N8335, N8333);
nand NAND2 (N8336, N8327, N3359);
xor XOR2 (N8337, N8332, N1699);
nor NOR2 (N8338, N8310, N7649);
buf BUF1 (N8339, N8321);
or OR4 (N8340, N8328, N6575, N6634, N1764);
nor NOR3 (N8341, N8340, N2981, N1556);
or OR2 (N8342, N8336, N186);
and AND4 (N8343, N8331, N7392, N2175, N7996);
nor NOR2 (N8344, N8339, N1296);
buf BUF1 (N8345, N8344);
not NOT1 (N8346, N8341);
and AND3 (N8347, N8346, N4059, N7418);
nand NAND2 (N8348, N8335, N2894);
xor XOR2 (N8349, N8337, N2873);
xor XOR2 (N8350, N8342, N2348);
nor NOR2 (N8351, N8343, N6506);
buf BUF1 (N8352, N8325);
not NOT1 (N8353, N8334);
xor XOR2 (N8354, N8353, N769);
nor NOR4 (N8355, N8347, N3662, N3500, N8044);
xor XOR2 (N8356, N8351, N1107);
nor NOR4 (N8357, N8301, N2973, N5930, N5238);
and AND3 (N8358, N8348, N2584, N949);
nor NOR2 (N8359, N8357, N1940);
or OR4 (N8360, N8338, N845, N2074, N6460);
not NOT1 (N8361, N8354);
nor NOR4 (N8362, N8361, N4434, N7466, N8181);
not NOT1 (N8363, N8358);
nor NOR3 (N8364, N8355, N6596, N7822);
or OR4 (N8365, N8363, N5936, N4345, N3943);
nand NAND4 (N8366, N8360, N1456, N2103, N3747);
nor NOR2 (N8367, N8364, N1716);
nand NAND4 (N8368, N8350, N6908, N1336, N2149);
not NOT1 (N8369, N8362);
nand NAND4 (N8370, N8345, N7673, N4800, N822);
or OR2 (N8371, N8367, N1172);
xor XOR2 (N8372, N8356, N6857);
buf BUF1 (N8373, N8370);
nor NOR3 (N8374, N8373, N8210, N6288);
xor XOR2 (N8375, N8359, N8320);
nor NOR3 (N8376, N8352, N2632, N5960);
buf BUF1 (N8377, N8365);
nor NOR2 (N8378, N8366, N2698);
buf BUF1 (N8379, N8376);
buf BUF1 (N8380, N8372);
buf BUF1 (N8381, N8380);
nand NAND4 (N8382, N8371, N749, N3589, N868);
buf BUF1 (N8383, N8368);
xor XOR2 (N8384, N8382, N5614);
xor XOR2 (N8385, N8377, N3593);
and AND2 (N8386, N8378, N2723);
buf BUF1 (N8387, N8369);
buf BUF1 (N8388, N8374);
or OR4 (N8389, N8385, N4138, N379, N1203);
or OR2 (N8390, N8375, N7832);
nor NOR3 (N8391, N8390, N8086, N906);
and AND2 (N8392, N8384, N950);
or OR4 (N8393, N8387, N4329, N2723, N4031);
xor XOR2 (N8394, N8389, N8391);
or OR3 (N8395, N7689, N2927, N7381);
nand NAND3 (N8396, N8394, N7625, N8114);
nor NOR2 (N8397, N8393, N3034);
nor NOR4 (N8398, N8396, N6791, N7186, N2763);
nand NAND2 (N8399, N8379, N3481);
and AND3 (N8400, N8398, N7898, N7113);
xor XOR2 (N8401, N8392, N7759);
xor XOR2 (N8402, N8400, N1129);
not NOT1 (N8403, N8381);
nor NOR2 (N8404, N8383, N2730);
not NOT1 (N8405, N8386);
nand NAND4 (N8406, N8404, N7936, N4944, N6073);
buf BUF1 (N8407, N8349);
not NOT1 (N8408, N8397);
nand NAND2 (N8409, N8403, N2807);
nor NOR3 (N8410, N8388, N2465, N6814);
and AND3 (N8411, N8408, N5820, N8325);
and AND3 (N8412, N8395, N6060, N4326);
and AND2 (N8413, N8401, N3655);
and AND4 (N8414, N8412, N7858, N7805, N6716);
or OR3 (N8415, N8409, N699, N1733);
nand NAND2 (N8416, N8402, N2810);
nor NOR3 (N8417, N8413, N7171, N4041);
xor XOR2 (N8418, N8407, N720);
and AND4 (N8419, N8414, N1633, N2485, N5919);
not NOT1 (N8420, N8399);
xor XOR2 (N8421, N8411, N2325);
nor NOR4 (N8422, N8415, N5793, N7341, N4631);
xor XOR2 (N8423, N8421, N3845);
or OR3 (N8424, N8419, N8233, N5632);
nand NAND2 (N8425, N8417, N4671);
nor NOR2 (N8426, N8422, N8360);
buf BUF1 (N8427, N8423);
not NOT1 (N8428, N8427);
nor NOR3 (N8429, N8420, N1882, N8370);
not NOT1 (N8430, N8418);
not NOT1 (N8431, N8406);
and AND4 (N8432, N8424, N585, N1945, N2052);
or OR4 (N8433, N8410, N36, N1109, N620);
or OR4 (N8434, N8429, N5382, N1978, N3630);
xor XOR2 (N8435, N8428, N8332);
buf BUF1 (N8436, N8435);
nor NOR2 (N8437, N8434, N2631);
not NOT1 (N8438, N8425);
nand NAND4 (N8439, N8431, N496, N4283, N68);
not NOT1 (N8440, N8430);
nand NAND4 (N8441, N8433, N6794, N5073, N1243);
not NOT1 (N8442, N8440);
or OR4 (N8443, N8439, N7199, N4521, N6596);
nand NAND3 (N8444, N8426, N113, N3633);
nand NAND4 (N8445, N8438, N8070, N7194, N5033);
xor XOR2 (N8446, N8445, N3988);
xor XOR2 (N8447, N8442, N6007);
not NOT1 (N8448, N8405);
and AND2 (N8449, N8447, N2469);
buf BUF1 (N8450, N8443);
or OR4 (N8451, N8450, N6147, N7096, N7233);
nand NAND2 (N8452, N8432, N1482);
xor XOR2 (N8453, N8448, N2605);
nor NOR2 (N8454, N8437, N4977);
or OR3 (N8455, N8452, N4798, N6481);
buf BUF1 (N8456, N8416);
buf BUF1 (N8457, N8456);
or OR4 (N8458, N8454, N1732, N3543, N2344);
and AND2 (N8459, N8453, N4747);
nor NOR3 (N8460, N8449, N7263, N617);
buf BUF1 (N8461, N8451);
xor XOR2 (N8462, N8444, N7767);
or OR3 (N8463, N8460, N7870, N7845);
xor XOR2 (N8464, N8457, N6602);
and AND3 (N8465, N8463, N8366, N1184);
or OR4 (N8466, N8462, N8364, N5459, N1924);
nand NAND3 (N8467, N8465, N2359, N5400);
nand NAND4 (N8468, N8458, N1201, N2569, N4334);
not NOT1 (N8469, N8468);
and AND2 (N8470, N8466, N4625);
buf BUF1 (N8471, N8455);
not NOT1 (N8472, N8470);
xor XOR2 (N8473, N8459, N3242);
xor XOR2 (N8474, N8471, N7467);
or OR4 (N8475, N8464, N2929, N6942, N8066);
xor XOR2 (N8476, N8473, N5876);
and AND4 (N8477, N8474, N1735, N103, N3665);
and AND2 (N8478, N8441, N2867);
nand NAND4 (N8479, N8469, N7971, N4873, N1345);
nand NAND2 (N8480, N8477, N1098);
not NOT1 (N8481, N8475);
xor XOR2 (N8482, N8461, N5168);
not NOT1 (N8483, N8482);
or OR4 (N8484, N8472, N4394, N781, N1160);
nand NAND4 (N8485, N8476, N1634, N6814, N5576);
or OR4 (N8486, N8484, N8121, N4694, N3628);
or OR3 (N8487, N8446, N5650, N3627);
nor NOR4 (N8488, N8467, N3081, N5974, N5056);
and AND4 (N8489, N8480, N5087, N1076, N3160);
or OR3 (N8490, N8489, N44, N558);
and AND4 (N8491, N8478, N5378, N258, N2858);
xor XOR2 (N8492, N8490, N6557);
or OR3 (N8493, N8486, N3410, N6684);
nand NAND2 (N8494, N8492, N8147);
not NOT1 (N8495, N8491);
and AND4 (N8496, N8487, N2491, N7134, N6665);
nand NAND4 (N8497, N8436, N5157, N524, N798);
or OR4 (N8498, N8494, N4680, N6838, N1838);
buf BUF1 (N8499, N8481);
and AND3 (N8500, N8496, N7332, N7719);
or OR3 (N8501, N8479, N6515, N4476);
not NOT1 (N8502, N8483);
nand NAND2 (N8503, N8493, N1515);
xor XOR2 (N8504, N8501, N3118);
or OR4 (N8505, N8498, N4120, N909, N3146);
and AND2 (N8506, N8497, N6500);
or OR4 (N8507, N8499, N7866, N522, N2397);
xor XOR2 (N8508, N8495, N2221);
or OR4 (N8509, N8500, N7239, N2706, N1466);
or OR4 (N8510, N8504, N6345, N1029, N5591);
not NOT1 (N8511, N8506);
buf BUF1 (N8512, N8509);
or OR2 (N8513, N8505, N2784);
or OR3 (N8514, N8485, N3239, N8459);
or OR3 (N8515, N8511, N3188, N1004);
or OR2 (N8516, N8512, N945);
and AND4 (N8517, N8514, N5359, N3528, N2007);
nand NAND2 (N8518, N8508, N6197);
or OR2 (N8519, N8510, N7445);
and AND3 (N8520, N8516, N2229, N2850);
or OR4 (N8521, N8519, N6992, N4768, N8463);
xor XOR2 (N8522, N8507, N7507);
not NOT1 (N8523, N8522);
buf BUF1 (N8524, N8517);
xor XOR2 (N8525, N8488, N956);
buf BUF1 (N8526, N8513);
and AND2 (N8527, N8521, N2382);
nor NOR2 (N8528, N8518, N198);
xor XOR2 (N8529, N8502, N1927);
and AND3 (N8530, N8528, N139, N7180);
nand NAND3 (N8531, N8503, N469, N2697);
nand NAND4 (N8532, N8529, N6284, N7256, N4965);
buf BUF1 (N8533, N8520);
xor XOR2 (N8534, N8532, N8203);
nor NOR4 (N8535, N8531, N50, N2852, N1245);
or OR4 (N8536, N8535, N5498, N2618, N7890);
xor XOR2 (N8537, N8526, N6237);
buf BUF1 (N8538, N8534);
nand NAND2 (N8539, N8515, N7051);
buf BUF1 (N8540, N8537);
buf BUF1 (N8541, N8524);
and AND2 (N8542, N8540, N7589);
nand NAND2 (N8543, N8538, N3992);
buf BUF1 (N8544, N8523);
and AND4 (N8545, N8536, N6508, N3368, N2817);
and AND2 (N8546, N8543, N4599);
and AND3 (N8547, N8530, N3801, N6056);
or OR3 (N8548, N8544, N6618, N7218);
not NOT1 (N8549, N8527);
nor NOR4 (N8550, N8533, N6913, N5635, N7883);
not NOT1 (N8551, N8547);
nand NAND4 (N8552, N8525, N3103, N7373, N2226);
xor XOR2 (N8553, N8551, N6652);
not NOT1 (N8554, N8553);
and AND4 (N8555, N8548, N2486, N8150, N374);
xor XOR2 (N8556, N8549, N6580);
xor XOR2 (N8557, N8545, N5438);
buf BUF1 (N8558, N8552);
or OR3 (N8559, N8554, N7609, N4095);
xor XOR2 (N8560, N8558, N3714);
not NOT1 (N8561, N8542);
xor XOR2 (N8562, N8561, N7178);
nand NAND3 (N8563, N8546, N7077, N6138);
and AND2 (N8564, N8539, N2302);
xor XOR2 (N8565, N8555, N7282);
buf BUF1 (N8566, N8557);
nand NAND2 (N8567, N8541, N5157);
not NOT1 (N8568, N8565);
xor XOR2 (N8569, N8556, N2885);
xor XOR2 (N8570, N8569, N6208);
buf BUF1 (N8571, N8563);
xor XOR2 (N8572, N8570, N4621);
nor NOR2 (N8573, N8566, N8503);
not NOT1 (N8574, N8564);
or OR4 (N8575, N8562, N3927, N4241, N1227);
nor NOR3 (N8576, N8568, N4141, N5167);
and AND2 (N8577, N8559, N4534);
and AND2 (N8578, N8574, N3745);
not NOT1 (N8579, N8550);
nand NAND3 (N8580, N8571, N2616, N3171);
xor XOR2 (N8581, N8572, N2078);
buf BUF1 (N8582, N8578);
nand NAND4 (N8583, N8573, N7598, N5883, N5457);
and AND3 (N8584, N8567, N7191, N4542);
not NOT1 (N8585, N8577);
buf BUF1 (N8586, N8560);
buf BUF1 (N8587, N8586);
nand NAND2 (N8588, N8583, N2199);
or OR3 (N8589, N8582, N2387, N8186);
xor XOR2 (N8590, N8585, N1836);
not NOT1 (N8591, N8581);
and AND3 (N8592, N8589, N1446, N5165);
buf BUF1 (N8593, N8576);
and AND2 (N8594, N8584, N1161);
nor NOR4 (N8595, N8592, N2564, N5069, N3444);
and AND3 (N8596, N8590, N6055, N6405);
not NOT1 (N8597, N8575);
and AND4 (N8598, N8597, N1667, N5352, N2321);
not NOT1 (N8599, N8598);
xor XOR2 (N8600, N8595, N1243);
and AND2 (N8601, N8596, N5820);
nor NOR3 (N8602, N8601, N3385, N80);
and AND4 (N8603, N8593, N1885, N2309, N7666);
xor XOR2 (N8604, N8599, N7313);
and AND4 (N8605, N8591, N7426, N1469, N7374);
or OR3 (N8606, N8604, N7414, N7060);
and AND2 (N8607, N8603, N3224);
or OR3 (N8608, N8605, N1686, N5925);
not NOT1 (N8609, N8608);
not NOT1 (N8610, N8580);
or OR4 (N8611, N8588, N5058, N6030, N2826);
nand NAND3 (N8612, N8610, N4302, N3731);
nand NAND2 (N8613, N8609, N4212);
not NOT1 (N8614, N8612);
buf BUF1 (N8615, N8606);
nor NOR2 (N8616, N8607, N7878);
nand NAND3 (N8617, N8602, N4449, N4212);
nor NOR2 (N8618, N8613, N3530);
or OR3 (N8619, N8617, N938, N1248);
nand NAND3 (N8620, N8587, N1319, N5147);
nor NOR4 (N8621, N8611, N1719, N7697, N1365);
buf BUF1 (N8622, N8594);
nor NOR4 (N8623, N8621, N7247, N6818, N6918);
nor NOR4 (N8624, N8616, N4953, N937, N2234);
nand NAND2 (N8625, N8619, N4767);
not NOT1 (N8626, N8615);
buf BUF1 (N8627, N8623);
and AND4 (N8628, N8614, N110, N1619, N7135);
and AND3 (N8629, N8620, N1660, N7383);
nor NOR2 (N8630, N8628, N8214);
nand NAND2 (N8631, N8626, N4587);
not NOT1 (N8632, N8625);
not NOT1 (N8633, N8627);
or OR2 (N8634, N8630, N2032);
not NOT1 (N8635, N8632);
nand NAND3 (N8636, N8634, N7534, N6176);
xor XOR2 (N8637, N8618, N6979);
not NOT1 (N8638, N8579);
not NOT1 (N8639, N8637);
and AND2 (N8640, N8635, N1935);
and AND3 (N8641, N8639, N8414, N4265);
xor XOR2 (N8642, N8622, N2915);
buf BUF1 (N8643, N8640);
and AND3 (N8644, N8643, N5156, N7502);
nand NAND3 (N8645, N8644, N8233, N8280);
or OR4 (N8646, N8641, N2747, N4298, N8113);
not NOT1 (N8647, N8646);
buf BUF1 (N8648, N8624);
buf BUF1 (N8649, N8633);
not NOT1 (N8650, N8629);
xor XOR2 (N8651, N8636, N5894);
buf BUF1 (N8652, N8650);
and AND4 (N8653, N8652, N8154, N2347, N5089);
buf BUF1 (N8654, N8631);
nand NAND2 (N8655, N8638, N2943);
buf BUF1 (N8656, N8600);
xor XOR2 (N8657, N8653, N8022);
not NOT1 (N8658, N8654);
xor XOR2 (N8659, N8655, N4367);
and AND3 (N8660, N8656, N427, N4349);
and AND4 (N8661, N8658, N8262, N7297, N213);
xor XOR2 (N8662, N8659, N4528);
nor NOR4 (N8663, N8660, N7627, N5447, N1314);
and AND2 (N8664, N8647, N397);
xor XOR2 (N8665, N8657, N331);
not NOT1 (N8666, N8665);
nor NOR2 (N8667, N8661, N6466);
nor NOR3 (N8668, N8648, N8053, N5275);
or OR4 (N8669, N8642, N6603, N3022, N4246);
nor NOR3 (N8670, N8651, N3559, N8400);
nand NAND4 (N8671, N8663, N5638, N5656, N7494);
or OR2 (N8672, N8671, N225);
buf BUF1 (N8673, N8664);
and AND3 (N8674, N8667, N5456, N6269);
nor NOR2 (N8675, N8666, N1093);
nor NOR3 (N8676, N8673, N3797, N3306);
nand NAND2 (N8677, N8674, N443);
and AND3 (N8678, N8675, N4387, N7945);
nand NAND2 (N8679, N8645, N1188);
xor XOR2 (N8680, N8649, N7553);
nand NAND4 (N8681, N8668, N3556, N8108, N738);
xor XOR2 (N8682, N8669, N3347);
nor NOR3 (N8683, N8676, N2597, N3256);
nor NOR3 (N8684, N8683, N6483, N4929);
or OR3 (N8685, N8682, N7197, N6524);
and AND3 (N8686, N8677, N8592, N8251);
nor NOR4 (N8687, N8680, N3401, N1385, N7833);
buf BUF1 (N8688, N8686);
buf BUF1 (N8689, N8685);
xor XOR2 (N8690, N8670, N1792);
buf BUF1 (N8691, N8681);
xor XOR2 (N8692, N8688, N3719);
xor XOR2 (N8693, N8662, N3961);
and AND4 (N8694, N8679, N2572, N179, N1779);
buf BUF1 (N8695, N8672);
nand NAND4 (N8696, N8691, N3879, N3399, N7665);
nand NAND2 (N8697, N8687, N908);
nor NOR3 (N8698, N8690, N4600, N3579);
or OR3 (N8699, N8689, N274, N3142);
and AND3 (N8700, N8697, N1725, N5485);
buf BUF1 (N8701, N8693);
or OR3 (N8702, N8692, N7157, N5198);
xor XOR2 (N8703, N8700, N5052);
and AND4 (N8704, N8699, N1379, N22, N8185);
or OR2 (N8705, N8704, N7367);
xor XOR2 (N8706, N8684, N6880);
or OR2 (N8707, N8695, N3320);
xor XOR2 (N8708, N8678, N5537);
xor XOR2 (N8709, N8702, N5263);
xor XOR2 (N8710, N8708, N2204);
and AND3 (N8711, N8709, N8646, N3239);
nor NOR2 (N8712, N8698, N5018);
xor XOR2 (N8713, N8694, N2545);
xor XOR2 (N8714, N8703, N3204);
or OR3 (N8715, N8714, N5194, N5386);
or OR2 (N8716, N8701, N5253);
nand NAND3 (N8717, N8716, N703, N8200);
or OR2 (N8718, N8696, N4277);
not NOT1 (N8719, N8711);
and AND3 (N8720, N8707, N2577, N1585);
not NOT1 (N8721, N8710);
buf BUF1 (N8722, N8712);
nor NOR2 (N8723, N8706, N6484);
nor NOR2 (N8724, N8723, N8295);
and AND3 (N8725, N8715, N4156, N3669);
or OR2 (N8726, N8705, N1221);
not NOT1 (N8727, N8724);
not NOT1 (N8728, N8722);
not NOT1 (N8729, N8718);
not NOT1 (N8730, N8717);
and AND2 (N8731, N8727, N2859);
or OR2 (N8732, N8729, N5414);
xor XOR2 (N8733, N8728, N7505);
or OR2 (N8734, N8731, N6948);
xor XOR2 (N8735, N8713, N4628);
nor NOR4 (N8736, N8721, N7504, N2681, N6458);
xor XOR2 (N8737, N8726, N1964);
buf BUF1 (N8738, N8733);
buf BUF1 (N8739, N8738);
or OR4 (N8740, N8725, N1519, N3000, N8229);
not NOT1 (N8741, N8735);
nand NAND4 (N8742, N8739, N6936, N3807, N7700);
not NOT1 (N8743, N8719);
and AND4 (N8744, N8743, N8743, N3699, N4775);
nor NOR4 (N8745, N8734, N1081, N1814, N7667);
not NOT1 (N8746, N8730);
and AND4 (N8747, N8732, N1977, N1536, N1980);
and AND2 (N8748, N8746, N2016);
and AND2 (N8749, N8737, N6386);
not NOT1 (N8750, N8736);
buf BUF1 (N8751, N8742);
nand NAND2 (N8752, N8751, N1606);
nand NAND4 (N8753, N8745, N7305, N8560, N7379);
nand NAND4 (N8754, N8748, N1752, N2647, N7298);
nor NOR4 (N8755, N8720, N2798, N5384, N3781);
nand NAND2 (N8756, N8749, N4147);
or OR3 (N8757, N8755, N4049, N376);
nand NAND4 (N8758, N8744, N2187, N7489, N1070);
nand NAND3 (N8759, N8757, N7542, N3138);
not NOT1 (N8760, N8758);
not NOT1 (N8761, N8756);
and AND4 (N8762, N8761, N1409, N5929, N4162);
xor XOR2 (N8763, N8759, N4626);
nor NOR3 (N8764, N8750, N3602, N6112);
xor XOR2 (N8765, N8763, N8592);
not NOT1 (N8766, N8764);
nor NOR3 (N8767, N8760, N1526, N1877);
buf BUF1 (N8768, N8767);
not NOT1 (N8769, N8747);
or OR2 (N8770, N8766, N6170);
buf BUF1 (N8771, N8752);
nor NOR3 (N8772, N8768, N8704, N6260);
xor XOR2 (N8773, N8772, N7843);
or OR3 (N8774, N8773, N5802, N5044);
and AND3 (N8775, N8765, N7165, N6018);
not NOT1 (N8776, N8753);
and AND3 (N8777, N8771, N3537, N7345);
buf BUF1 (N8778, N8762);
and AND2 (N8779, N8770, N8483);
xor XOR2 (N8780, N8776, N5721);
nor NOR3 (N8781, N8780, N7938, N7121);
and AND3 (N8782, N8779, N5794, N5271);
and AND2 (N8783, N8775, N7910);
nand NAND3 (N8784, N8782, N5918, N3868);
not NOT1 (N8785, N8777);
nor NOR2 (N8786, N8784, N460);
xor XOR2 (N8787, N8778, N7534);
not NOT1 (N8788, N8741);
buf BUF1 (N8789, N8788);
nand NAND2 (N8790, N8769, N3244);
buf BUF1 (N8791, N8740);
buf BUF1 (N8792, N8783);
xor XOR2 (N8793, N8786, N7788);
buf BUF1 (N8794, N8789);
buf BUF1 (N8795, N8793);
nand NAND4 (N8796, N8785, N3716, N3183, N8488);
nand NAND2 (N8797, N8796, N4752);
buf BUF1 (N8798, N8791);
and AND4 (N8799, N8774, N8187, N2714, N6578);
not NOT1 (N8800, N8790);
or OR4 (N8801, N8792, N3049, N2670, N5057);
xor XOR2 (N8802, N8794, N7467);
not NOT1 (N8803, N8797);
not NOT1 (N8804, N8802);
nor NOR2 (N8805, N8798, N6806);
not NOT1 (N8806, N8805);
or OR2 (N8807, N8754, N5978);
xor XOR2 (N8808, N8806, N2533);
or OR2 (N8809, N8804, N2091);
buf BUF1 (N8810, N8800);
buf BUF1 (N8811, N8801);
and AND4 (N8812, N8795, N4503, N6791, N8675);
nor NOR3 (N8813, N8787, N7592, N5040);
or OR4 (N8814, N8812, N4170, N2454, N190);
nor NOR2 (N8815, N8809, N4495);
or OR3 (N8816, N8808, N6963, N2289);
and AND3 (N8817, N8815, N5472, N4202);
buf BUF1 (N8818, N8810);
nor NOR3 (N8819, N8813, N157, N5366);
nand NAND3 (N8820, N8816, N2833, N1295);
buf BUF1 (N8821, N8818);
nor NOR2 (N8822, N8819, N2163);
nor NOR3 (N8823, N8820, N8689, N8537);
xor XOR2 (N8824, N8799, N3182);
xor XOR2 (N8825, N8803, N4388);
nor NOR3 (N8826, N8821, N5553, N4478);
xor XOR2 (N8827, N8824, N4123);
buf BUF1 (N8828, N8825);
nor NOR4 (N8829, N8827, N6416, N3263, N7643);
buf BUF1 (N8830, N8829);
nand NAND4 (N8831, N8811, N8258, N5288, N4208);
or OR2 (N8832, N8781, N4491);
buf BUF1 (N8833, N8822);
or OR2 (N8834, N8830, N3826);
xor XOR2 (N8835, N8831, N8697);
nand NAND3 (N8836, N8833, N7977, N6710);
not NOT1 (N8837, N8807);
not NOT1 (N8838, N8837);
nor NOR2 (N8839, N8832, N6215);
not NOT1 (N8840, N8814);
buf BUF1 (N8841, N8817);
nand NAND3 (N8842, N8841, N1176, N4650);
nand NAND3 (N8843, N8828, N5614, N1630);
nor NOR4 (N8844, N8843, N476, N5474, N1515);
nor NOR3 (N8845, N8826, N2434, N6895);
buf BUF1 (N8846, N8844);
buf BUF1 (N8847, N8839);
nand NAND4 (N8848, N8835, N1593, N4881, N7423);
nor NOR2 (N8849, N8840, N7324);
not NOT1 (N8850, N8847);
or OR2 (N8851, N8823, N6068);
nand NAND4 (N8852, N8850, N5773, N1941, N8293);
not NOT1 (N8853, N8838);
or OR3 (N8854, N8834, N3851, N7800);
xor XOR2 (N8855, N8836, N6643);
or OR2 (N8856, N8848, N360);
nand NAND3 (N8857, N8852, N536, N8244);
nor NOR2 (N8858, N8851, N5437);
buf BUF1 (N8859, N8857);
not NOT1 (N8860, N8856);
and AND4 (N8861, N8845, N695, N285, N5110);
or OR4 (N8862, N8849, N5185, N783, N1273);
nand NAND2 (N8863, N8859, N3972);
or OR2 (N8864, N8860, N8401);
and AND2 (N8865, N8863, N2605);
and AND2 (N8866, N8862, N3470);
and AND2 (N8867, N8864, N5656);
nor NOR3 (N8868, N8842, N8332, N1673);
nand NAND3 (N8869, N8865, N5663, N1944);
nand NAND4 (N8870, N8861, N3726, N3689, N4682);
or OR4 (N8871, N8854, N5862, N7186, N2016);
not NOT1 (N8872, N8869);
buf BUF1 (N8873, N8858);
not NOT1 (N8874, N8868);
nand NAND4 (N8875, N8872, N735, N7014, N6256);
and AND2 (N8876, N8866, N8485);
and AND4 (N8877, N8871, N3062, N3654, N3);
or OR3 (N8878, N8875, N5102, N7282);
nor NOR3 (N8879, N8853, N2442, N3884);
and AND4 (N8880, N8873, N1567, N4449, N7612);
nand NAND2 (N8881, N8874, N2535);
not NOT1 (N8882, N8846);
buf BUF1 (N8883, N8881);
xor XOR2 (N8884, N8876, N4419);
or OR2 (N8885, N8878, N2928);
xor XOR2 (N8886, N8855, N4927);
not NOT1 (N8887, N8879);
nor NOR3 (N8888, N8867, N1870, N3239);
not NOT1 (N8889, N8883);
buf BUF1 (N8890, N8888);
or OR3 (N8891, N8877, N7594, N7117);
and AND3 (N8892, N8880, N121, N5431);
nand NAND3 (N8893, N8886, N8049, N4973);
xor XOR2 (N8894, N8887, N5501);
or OR4 (N8895, N8892, N1426, N1603, N1264);
not NOT1 (N8896, N8884);
and AND2 (N8897, N8893, N3694);
xor XOR2 (N8898, N8897, N6006);
and AND3 (N8899, N8882, N6020, N2468);
not NOT1 (N8900, N8894);
or OR3 (N8901, N8898, N5616, N1649);
or OR3 (N8902, N8895, N3901, N4192);
buf BUF1 (N8903, N8891);
or OR2 (N8904, N8885, N7914);
nand NAND2 (N8905, N8889, N6620);
or OR3 (N8906, N8900, N4781, N8451);
xor XOR2 (N8907, N8896, N6119);
xor XOR2 (N8908, N8905, N8207);
or OR4 (N8909, N8908, N3814, N3896, N5764);
buf BUF1 (N8910, N8909);
nor NOR3 (N8911, N8904, N4960, N7196);
and AND4 (N8912, N8903, N3481, N3068, N7281);
and AND4 (N8913, N8890, N8653, N4078, N7539);
xor XOR2 (N8914, N8906, N8265);
nor NOR3 (N8915, N8913, N461, N1303);
nand NAND3 (N8916, N8902, N8534, N4195);
and AND3 (N8917, N8911, N5427, N494);
not NOT1 (N8918, N8915);
or OR2 (N8919, N8870, N6170);
and AND4 (N8920, N8914, N3402, N5536, N962);
nor NOR3 (N8921, N8912, N4581, N7545);
and AND4 (N8922, N8921, N4209, N1110, N3184);
not NOT1 (N8923, N8916);
nand NAND4 (N8924, N8910, N695, N1273, N81);
and AND2 (N8925, N8923, N7581);
nand NAND2 (N8926, N8907, N2554);
not NOT1 (N8927, N8918);
nor NOR2 (N8928, N8920, N7455);
or OR4 (N8929, N8917, N4894, N508, N2910);
and AND3 (N8930, N8929, N2354, N4487);
xor XOR2 (N8931, N8924, N5850);
buf BUF1 (N8932, N8926);
not NOT1 (N8933, N8901);
nand NAND4 (N8934, N8931, N6855, N3010, N6410);
not NOT1 (N8935, N8919);
and AND2 (N8936, N8935, N1593);
nor NOR3 (N8937, N8933, N985, N2613);
not NOT1 (N8938, N8930);
buf BUF1 (N8939, N8937);
or OR2 (N8940, N8922, N1863);
buf BUF1 (N8941, N8925);
or OR4 (N8942, N8928, N8176, N2301, N8742);
not NOT1 (N8943, N8927);
nand NAND2 (N8944, N8943, N5086);
or OR3 (N8945, N8939, N8803, N2043);
or OR3 (N8946, N8944, N4248, N7276);
or OR3 (N8947, N8942, N5908, N4050);
nor NOR4 (N8948, N8940, N664, N8897, N2655);
xor XOR2 (N8949, N8948, N2528);
nor NOR4 (N8950, N8938, N2456, N2079, N8238);
not NOT1 (N8951, N8941);
nor NOR2 (N8952, N8947, N3384);
not NOT1 (N8953, N8951);
nand NAND3 (N8954, N8950, N1204, N8517);
nand NAND2 (N8955, N8953, N8695);
nor NOR2 (N8956, N8949, N3851);
xor XOR2 (N8957, N8955, N1100);
or OR2 (N8958, N8954, N8025);
or OR3 (N8959, N8946, N3891, N956);
xor XOR2 (N8960, N8934, N8078);
xor XOR2 (N8961, N8958, N469);
nand NAND4 (N8962, N8957, N1918, N3651, N590);
nand NAND2 (N8963, N8962, N2347);
nor NOR2 (N8964, N8899, N1177);
or OR2 (N8965, N8952, N6327);
and AND4 (N8966, N8936, N2203, N7597, N1249);
xor XOR2 (N8967, N8961, N1466);
or OR3 (N8968, N8956, N87, N6924);
or OR3 (N8969, N8945, N5492, N6859);
buf BUF1 (N8970, N8968);
and AND2 (N8971, N8960, N3050);
or OR3 (N8972, N8971, N3331, N7951);
or OR4 (N8973, N8972, N7693, N1814, N6267);
buf BUF1 (N8974, N8970);
buf BUF1 (N8975, N8969);
xor XOR2 (N8976, N8963, N4076);
nand NAND3 (N8977, N8973, N3135, N1495);
xor XOR2 (N8978, N8976, N8256);
xor XOR2 (N8979, N8959, N8893);
not NOT1 (N8980, N8932);
buf BUF1 (N8981, N8979);
nor NOR2 (N8982, N8967, N7559);
and AND4 (N8983, N8978, N4050, N2262, N4213);
or OR2 (N8984, N8981, N2904);
nand NAND3 (N8985, N8974, N4986, N4170);
nor NOR3 (N8986, N8983, N3108, N5649);
and AND3 (N8987, N8984, N4807, N1344);
nor NOR2 (N8988, N8977, N5153);
not NOT1 (N8989, N8980);
nand NAND2 (N8990, N8975, N2678);
nor NOR2 (N8991, N8966, N8411);
xor XOR2 (N8992, N8964, N6063);
xor XOR2 (N8993, N8991, N1422);
and AND3 (N8994, N8989, N7836, N4492);
and AND3 (N8995, N8986, N2898, N290);
nand NAND3 (N8996, N8965, N8704, N534);
not NOT1 (N8997, N8995);
or OR2 (N8998, N8982, N4647);
or OR4 (N8999, N8985, N8104, N2484, N777);
nor NOR4 (N9000, N8987, N7266, N634, N8155);
nand NAND2 (N9001, N8988, N1091);
xor XOR2 (N9002, N8999, N5728);
buf BUF1 (N9003, N8998);
nor NOR2 (N9004, N8994, N3016);
and AND3 (N9005, N9000, N4878, N2357);
not NOT1 (N9006, N8996);
buf BUF1 (N9007, N8993);
or OR4 (N9008, N9003, N3091, N5095, N2313);
or OR4 (N9009, N8992, N43, N4192, N4736);
nor NOR3 (N9010, N9007, N6052, N2204);
or OR2 (N9011, N9004, N2270);
or OR2 (N9012, N9008, N2763);
nor NOR4 (N9013, N9011, N7771, N692, N7914);
nand NAND2 (N9014, N9005, N832);
nor NOR4 (N9015, N9012, N6084, N5036, N7057);
not NOT1 (N9016, N9014);
xor XOR2 (N9017, N9015, N5016);
nand NAND4 (N9018, N9002, N6111, N1978, N1377);
not NOT1 (N9019, N9016);
not NOT1 (N9020, N9013);
buf BUF1 (N9021, N9020);
nand NAND3 (N9022, N9018, N260, N2732);
nor NOR4 (N9023, N9006, N3879, N7248, N4004);
and AND4 (N9024, N8997, N3390, N6601, N3884);
not NOT1 (N9025, N9024);
not NOT1 (N9026, N8990);
and AND4 (N9027, N9017, N3544, N5286, N7604);
nor NOR3 (N9028, N9027, N1194, N2252);
and AND2 (N9029, N9023, N1883);
nand NAND3 (N9030, N9022, N3523, N4096);
nand NAND2 (N9031, N9026, N7599);
nand NAND3 (N9032, N9021, N4272, N5429);
xor XOR2 (N9033, N9019, N4546);
xor XOR2 (N9034, N9009, N5544);
xor XOR2 (N9035, N9030, N3813);
nor NOR3 (N9036, N9035, N874, N4537);
or OR3 (N9037, N9029, N4484, N2486);
or OR2 (N9038, N9034, N1020);
buf BUF1 (N9039, N9033);
xor XOR2 (N9040, N9025, N2349);
or OR3 (N9041, N9037, N3776, N7739);
nor NOR3 (N9042, N9010, N8801, N7201);
and AND4 (N9043, N9031, N179, N8726, N6256);
nand NAND3 (N9044, N9043, N4784, N90);
nand NAND3 (N9045, N9038, N8785, N2324);
nor NOR3 (N9046, N9040, N2286, N8103);
nor NOR4 (N9047, N9036, N2266, N7126, N2457);
not NOT1 (N9048, N9001);
buf BUF1 (N9049, N9042);
nor NOR2 (N9050, N9047, N1376);
nor NOR3 (N9051, N9032, N4378, N8482);
xor XOR2 (N9052, N9046, N7243);
xor XOR2 (N9053, N9045, N5425);
not NOT1 (N9054, N9050);
and AND2 (N9055, N9049, N6154);
buf BUF1 (N9056, N9053);
and AND3 (N9057, N9048, N8473, N8690);
or OR4 (N9058, N9055, N6009, N8050, N3823);
nand NAND3 (N9059, N9054, N458, N5329);
and AND2 (N9060, N9051, N3879);
and AND2 (N9061, N9041, N6349);
nand NAND3 (N9062, N9059, N1339, N5797);
or OR2 (N9063, N9060, N967);
or OR3 (N9064, N9057, N2718, N3493);
nor NOR2 (N9065, N9052, N4786);
or OR2 (N9066, N9058, N572);
or OR3 (N9067, N9039, N629, N2574);
nand NAND4 (N9068, N9063, N7879, N5509, N7886);
buf BUF1 (N9069, N9067);
nor NOR2 (N9070, N9056, N2210);
nor NOR2 (N9071, N9066, N5512);
xor XOR2 (N9072, N9061, N1047);
buf BUF1 (N9073, N9072);
or OR4 (N9074, N9070, N6690, N4844, N2604);
nand NAND3 (N9075, N9062, N5132, N4513);
nand NAND3 (N9076, N9069, N3406, N709);
xor XOR2 (N9077, N9074, N4845);
nor NOR4 (N9078, N9028, N5501, N2429, N5688);
nor NOR3 (N9079, N9064, N4260, N6212);
xor XOR2 (N9080, N9044, N3138);
not NOT1 (N9081, N9080);
not NOT1 (N9082, N9076);
and AND2 (N9083, N9081, N8903);
or OR4 (N9084, N9068, N3514, N3498, N6050);
nand NAND2 (N9085, N9079, N2890);
or OR2 (N9086, N9075, N1663);
buf BUF1 (N9087, N9071);
buf BUF1 (N9088, N9087);
buf BUF1 (N9089, N9086);
not NOT1 (N9090, N9089);
or OR2 (N9091, N9077, N6090);
buf BUF1 (N9092, N9088);
buf BUF1 (N9093, N9083);
not NOT1 (N9094, N9065);
buf BUF1 (N9095, N9094);
nor NOR2 (N9096, N9085, N5539);
or OR3 (N9097, N9073, N3801, N8923);
nand NAND2 (N9098, N9090, N3974);
or OR2 (N9099, N9082, N7918);
nor NOR3 (N9100, N9078, N6915, N1411);
and AND3 (N9101, N9097, N1228, N4353);
and AND4 (N9102, N9084, N5501, N6950, N1994);
xor XOR2 (N9103, N9095, N697);
xor XOR2 (N9104, N9091, N4899);
nand NAND3 (N9105, N9092, N7659, N2759);
xor XOR2 (N9106, N9099, N7063);
xor XOR2 (N9107, N9100, N4490);
not NOT1 (N9108, N9105);
nand NAND3 (N9109, N9107, N390, N810);
buf BUF1 (N9110, N9104);
or OR4 (N9111, N9108, N2040, N4739, N4016);
nor NOR2 (N9112, N9109, N8891);
xor XOR2 (N9113, N9112, N7656);
nand NAND2 (N9114, N9103, N4520);
nand NAND3 (N9115, N9098, N6333, N2014);
or OR2 (N9116, N9113, N4297);
nand NAND2 (N9117, N9093, N1220);
xor XOR2 (N9118, N9115, N2811);
nand NAND4 (N9119, N9106, N3980, N82, N3794);
nand NAND2 (N9120, N9101, N5198);
and AND2 (N9121, N9111, N8298);
or OR2 (N9122, N9120, N2072);
buf BUF1 (N9123, N9102);
nand NAND2 (N9124, N9121, N5266);
or OR2 (N9125, N9124, N3172);
buf BUF1 (N9126, N9117);
nor NOR2 (N9127, N9096, N3455);
or OR2 (N9128, N9127, N7853);
and AND2 (N9129, N9114, N7004);
xor XOR2 (N9130, N9118, N7823);
xor XOR2 (N9131, N9125, N2136);
xor XOR2 (N9132, N9119, N5443);
and AND3 (N9133, N9122, N4127, N6077);
xor XOR2 (N9134, N9126, N8116);
or OR2 (N9135, N9129, N6385);
nor NOR2 (N9136, N9133, N2979);
not NOT1 (N9137, N9128);
nor NOR4 (N9138, N9116, N3881, N1300, N7011);
nor NOR3 (N9139, N9110, N6075, N823);
not NOT1 (N9140, N9135);
or OR3 (N9141, N9123, N2161, N3413);
and AND2 (N9142, N9139, N136);
buf BUF1 (N9143, N9137);
and AND4 (N9144, N9138, N7690, N5983, N5021);
xor XOR2 (N9145, N9136, N78);
nand NAND4 (N9146, N9143, N5548, N2235, N2556);
and AND2 (N9147, N9145, N6082);
and AND2 (N9148, N9147, N3598);
buf BUF1 (N9149, N9130);
and AND3 (N9150, N9142, N1734, N553);
or OR4 (N9151, N9148, N2309, N6520, N7372);
not NOT1 (N9152, N9134);
and AND3 (N9153, N9146, N8030, N120);
nor NOR4 (N9154, N9131, N5969, N2478, N2028);
or OR2 (N9155, N9144, N8824);
not NOT1 (N9156, N9149);
buf BUF1 (N9157, N9141);
not NOT1 (N9158, N9150);
nand NAND4 (N9159, N9153, N3213, N2323, N6364);
or OR2 (N9160, N9132, N835);
nor NOR3 (N9161, N9140, N6558, N8608);
nand NAND2 (N9162, N9157, N2389);
buf BUF1 (N9163, N9152);
and AND4 (N9164, N9161, N8205, N8273, N3587);
xor XOR2 (N9165, N9164, N5895);
nor NOR4 (N9166, N9158, N5423, N1145, N1416);
not NOT1 (N9167, N9151);
nor NOR4 (N9168, N9155, N1141, N6769, N3402);
not NOT1 (N9169, N9166);
not NOT1 (N9170, N9167);
and AND4 (N9171, N9154, N3431, N5702, N6410);
xor XOR2 (N9172, N9159, N6994);
nor NOR3 (N9173, N9172, N2923, N4749);
nand NAND4 (N9174, N9162, N1031, N5260, N6636);
not NOT1 (N9175, N9170);
and AND2 (N9176, N9160, N7315);
buf BUF1 (N9177, N9171);
nand NAND4 (N9178, N9173, N6132, N4290, N4422);
nor NOR3 (N9179, N9176, N8493, N2293);
not NOT1 (N9180, N9165);
buf BUF1 (N9181, N9175);
not NOT1 (N9182, N9169);
nand NAND2 (N9183, N9174, N1394);
buf BUF1 (N9184, N9179);
not NOT1 (N9185, N9183);
nand NAND4 (N9186, N9180, N6627, N3856, N8726);
nand NAND3 (N9187, N9186, N6632, N8204);
buf BUF1 (N9188, N9168);
buf BUF1 (N9189, N9182);
buf BUF1 (N9190, N9156);
xor XOR2 (N9191, N9189, N4333);
nand NAND3 (N9192, N9177, N1200, N8727);
nand NAND2 (N9193, N9185, N908);
buf BUF1 (N9194, N9181);
and AND3 (N9195, N9193, N6664, N551);
xor XOR2 (N9196, N9191, N3058);
nand NAND3 (N9197, N9178, N1190, N2045);
and AND4 (N9198, N9197, N3821, N1672, N9131);
nand NAND3 (N9199, N9198, N3251, N3526);
or OR2 (N9200, N9190, N4481);
not NOT1 (N9201, N9200);
nand NAND3 (N9202, N9201, N8996, N5494);
buf BUF1 (N9203, N9192);
nor NOR4 (N9204, N9194, N4902, N4201, N6080);
nand NAND4 (N9205, N9187, N5616, N5517, N1897);
and AND3 (N9206, N9204, N3493, N7788);
buf BUF1 (N9207, N9163);
xor XOR2 (N9208, N9199, N5693);
buf BUF1 (N9209, N9207);
xor XOR2 (N9210, N9209, N938);
nand NAND2 (N9211, N9208, N6249);
nor NOR2 (N9212, N9195, N7610);
nor NOR2 (N9213, N9188, N561);
or OR4 (N9214, N9196, N7939, N3007, N109);
or OR3 (N9215, N9214, N4951, N8353);
or OR4 (N9216, N9213, N2544, N353, N5977);
buf BUF1 (N9217, N9202);
xor XOR2 (N9218, N9217, N276);
nand NAND3 (N9219, N9211, N5326, N4257);
buf BUF1 (N9220, N9203);
nor NOR2 (N9221, N9205, N9002);
or OR4 (N9222, N9210, N5078, N4278, N3651);
xor XOR2 (N9223, N9222, N1511);
buf BUF1 (N9224, N9221);
and AND3 (N9225, N9215, N1524, N1392);
or OR3 (N9226, N9206, N7000, N3489);
nand NAND2 (N9227, N9220, N3721);
xor XOR2 (N9228, N9219, N7548);
and AND2 (N9229, N9228, N5069);
nor NOR3 (N9230, N9184, N4627, N7419);
and AND2 (N9231, N9224, N6291);
nand NAND4 (N9232, N9223, N2656, N7831, N5648);
xor XOR2 (N9233, N9216, N3657);
or OR3 (N9234, N9212, N7235, N6373);
nor NOR2 (N9235, N9218, N4175);
buf BUF1 (N9236, N9227);
and AND4 (N9237, N9229, N2991, N6012, N1137);
buf BUF1 (N9238, N9234);
and AND2 (N9239, N9237, N1913);
nand NAND2 (N9240, N9226, N6835);
not NOT1 (N9241, N9225);
xor XOR2 (N9242, N9240, N652);
nand NAND4 (N9243, N9232, N2239, N3717, N8394);
nand NAND4 (N9244, N9233, N5089, N7817, N713);
nand NAND3 (N9245, N9235, N5937, N5581);
or OR4 (N9246, N9230, N8541, N5520, N1942);
xor XOR2 (N9247, N9231, N1132);
not NOT1 (N9248, N9246);
nand NAND4 (N9249, N9236, N2865, N7404, N1278);
nand NAND2 (N9250, N9249, N6852);
buf BUF1 (N9251, N9238);
xor XOR2 (N9252, N9239, N1196);
not NOT1 (N9253, N9245);
nand NAND4 (N9254, N9252, N5991, N2163, N2660);
nor NOR2 (N9255, N9254, N6212);
and AND4 (N9256, N9244, N7533, N7175, N7671);
nand NAND4 (N9257, N9248, N4853, N5393, N4181);
nand NAND3 (N9258, N9251, N5744, N1346);
and AND4 (N9259, N9255, N8276, N5830, N2863);
nand NAND2 (N9260, N9258, N6193);
buf BUF1 (N9261, N9256);
nand NAND2 (N9262, N9257, N5830);
not NOT1 (N9263, N9259);
xor XOR2 (N9264, N9242, N12);
nor NOR2 (N9265, N9262, N2582);
or OR3 (N9266, N9264, N206, N3274);
buf BUF1 (N9267, N9263);
and AND3 (N9268, N9265, N3830, N5862);
nand NAND4 (N9269, N9267, N6165, N7422, N2645);
buf BUF1 (N9270, N9266);
xor XOR2 (N9271, N9253, N8241);
nor NOR3 (N9272, N9241, N7102, N2107);
nand NAND3 (N9273, N9268, N4619, N8206);
not NOT1 (N9274, N9261);
and AND4 (N9275, N9247, N2541, N6867, N2278);
buf BUF1 (N9276, N9260);
buf BUF1 (N9277, N9276);
not NOT1 (N9278, N9273);
and AND3 (N9279, N9278, N5492, N6577);
nor NOR2 (N9280, N9269, N7100);
buf BUF1 (N9281, N9279);
or OR4 (N9282, N9275, N7224, N2256, N8297);
buf BUF1 (N9283, N9280);
nor NOR3 (N9284, N9282, N6703, N5654);
buf BUF1 (N9285, N9277);
buf BUF1 (N9286, N9281);
or OR3 (N9287, N9274, N8147, N3896);
xor XOR2 (N9288, N9243, N3944);
buf BUF1 (N9289, N9288);
nor NOR3 (N9290, N9271, N4977, N6622);
or OR3 (N9291, N9286, N1193, N367);
nand NAND2 (N9292, N9285, N3971);
buf BUF1 (N9293, N9284);
buf BUF1 (N9294, N9293);
and AND2 (N9295, N9290, N5657);
and AND3 (N9296, N9283, N4142, N2316);
nor NOR3 (N9297, N9250, N8730, N9146);
and AND2 (N9298, N9289, N7365);
nor NOR2 (N9299, N9291, N1595);
not NOT1 (N9300, N9299);
not NOT1 (N9301, N9287);
or OR3 (N9302, N9296, N5294, N4618);
or OR4 (N9303, N9270, N6573, N1432, N834);
and AND2 (N9304, N9298, N969);
nand NAND2 (N9305, N9272, N4068);
buf BUF1 (N9306, N9300);
or OR3 (N9307, N9301, N1246, N4318);
xor XOR2 (N9308, N9295, N7576);
nor NOR2 (N9309, N9307, N7646);
xor XOR2 (N9310, N9297, N7128);
not NOT1 (N9311, N9309);
and AND2 (N9312, N9308, N1647);
xor XOR2 (N9313, N9311, N862);
nand NAND4 (N9314, N9292, N6191, N4267, N975);
or OR2 (N9315, N9305, N3931);
not NOT1 (N9316, N9314);
not NOT1 (N9317, N9294);
nand NAND2 (N9318, N9316, N9150);
buf BUF1 (N9319, N9310);
buf BUF1 (N9320, N9315);
or OR2 (N9321, N9313, N2089);
xor XOR2 (N9322, N9303, N2180);
nor NOR3 (N9323, N9319, N166, N5366);
xor XOR2 (N9324, N9312, N1324);
nor NOR2 (N9325, N9317, N8195);
or OR4 (N9326, N9325, N2919, N3427, N9175);
or OR2 (N9327, N9304, N6986);
nor NOR4 (N9328, N9322, N6255, N1304, N5706);
and AND3 (N9329, N9326, N813, N6003);
or OR4 (N9330, N9324, N33, N8697, N6471);
nand NAND4 (N9331, N9329, N1970, N6275, N7414);
nor NOR3 (N9332, N9302, N9022, N9187);
nor NOR3 (N9333, N9321, N2840, N2620);
nand NAND3 (N9334, N9320, N2006, N1672);
not NOT1 (N9335, N9328);
nor NOR2 (N9336, N9333, N736);
not NOT1 (N9337, N9335);
nor NOR3 (N9338, N9318, N2259, N998);
nor NOR2 (N9339, N9331, N7033);
buf BUF1 (N9340, N9330);
buf BUF1 (N9341, N9332);
or OR2 (N9342, N9327, N6241);
and AND4 (N9343, N9342, N3804, N1436, N7635);
and AND2 (N9344, N9340, N7056);
and AND2 (N9345, N9343, N6158);
buf BUF1 (N9346, N9323);
and AND3 (N9347, N9337, N7794, N2834);
not NOT1 (N9348, N9334);
and AND2 (N9349, N9341, N468);
nand NAND4 (N9350, N9348, N3252, N3593, N829);
nand NAND3 (N9351, N9306, N2276, N8885);
nor NOR4 (N9352, N9349, N2529, N6337, N3459);
not NOT1 (N9353, N9346);
buf BUF1 (N9354, N9353);
nor NOR4 (N9355, N9351, N3949, N7545, N8006);
buf BUF1 (N9356, N9345);
and AND2 (N9357, N9336, N8868);
nor NOR2 (N9358, N9347, N96);
nand NAND3 (N9359, N9354, N3172, N1660);
buf BUF1 (N9360, N9350);
not NOT1 (N9361, N9344);
buf BUF1 (N9362, N9358);
not NOT1 (N9363, N9339);
and AND3 (N9364, N9352, N6720, N5952);
or OR4 (N9365, N9356, N2517, N6397, N7253);
not NOT1 (N9366, N9357);
xor XOR2 (N9367, N9366, N111);
or OR3 (N9368, N9338, N6860, N1408);
nand NAND3 (N9369, N9359, N6919, N5941);
or OR4 (N9370, N9367, N4207, N9323, N8051);
not NOT1 (N9371, N9361);
xor XOR2 (N9372, N9364, N2070);
nand NAND4 (N9373, N9369, N4333, N1485, N9053);
or OR3 (N9374, N9365, N6793, N6439);
not NOT1 (N9375, N9371);
nand NAND3 (N9376, N9355, N5690, N7871);
nor NOR4 (N9377, N9375, N645, N5057, N2217);
nor NOR2 (N9378, N9374, N3931);
xor XOR2 (N9379, N9372, N904);
xor XOR2 (N9380, N9373, N2446);
buf BUF1 (N9381, N9363);
or OR2 (N9382, N9381, N1282);
nor NOR3 (N9383, N9377, N9259, N4015);
nor NOR2 (N9384, N9379, N3919);
not NOT1 (N9385, N9383);
or OR2 (N9386, N9376, N1137);
or OR2 (N9387, N9378, N7809);
xor XOR2 (N9388, N9384, N1664);
and AND3 (N9389, N9368, N3653, N511);
xor XOR2 (N9390, N9385, N2957);
or OR4 (N9391, N9389, N8768, N1138, N516);
not NOT1 (N9392, N9391);
not NOT1 (N9393, N9392);
xor XOR2 (N9394, N9362, N2343);
not NOT1 (N9395, N9382);
nand NAND2 (N9396, N9380, N7302);
nand NAND3 (N9397, N9390, N6540, N328);
nand NAND2 (N9398, N9360, N315);
or OR4 (N9399, N9386, N4688, N5366, N7162);
not NOT1 (N9400, N9388);
and AND4 (N9401, N9370, N2750, N3918, N2074);
and AND4 (N9402, N9396, N8563, N3721, N8677);
not NOT1 (N9403, N9387);
xor XOR2 (N9404, N9399, N7083);
buf BUF1 (N9405, N9404);
xor XOR2 (N9406, N9398, N2106);
and AND4 (N9407, N9397, N2068, N2943, N7406);
buf BUF1 (N9408, N9394);
and AND4 (N9409, N9405, N4914, N2724, N6545);
not NOT1 (N9410, N9393);
not NOT1 (N9411, N9410);
nand NAND3 (N9412, N9403, N2351, N6931);
nor NOR3 (N9413, N9395, N4718, N2546);
buf BUF1 (N9414, N9413);
xor XOR2 (N9415, N9412, N1965);
buf BUF1 (N9416, N9414);
not NOT1 (N9417, N9400);
or OR2 (N9418, N9406, N8130);
or OR3 (N9419, N9411, N6402, N3845);
nand NAND3 (N9420, N9407, N6434, N5451);
nor NOR3 (N9421, N9415, N1476, N2884);
and AND4 (N9422, N9421, N9097, N8320, N945);
nand NAND3 (N9423, N9401, N2365, N417);
not NOT1 (N9424, N9408);
and AND2 (N9425, N9417, N3575);
or OR4 (N9426, N9422, N1538, N8618, N4767);
xor XOR2 (N9427, N9425, N5908);
nor NOR2 (N9428, N9423, N2359);
and AND3 (N9429, N9416, N8907, N3175);
and AND2 (N9430, N9402, N4373);
buf BUF1 (N9431, N9419);
xor XOR2 (N9432, N9429, N405);
nand NAND4 (N9433, N9427, N8228, N6509, N6872);
nor NOR2 (N9434, N9432, N4026);
or OR4 (N9435, N9424, N6119, N8770, N1275);
and AND2 (N9436, N9426, N535);
nor NOR3 (N9437, N9428, N811, N3916);
buf BUF1 (N9438, N9433);
xor XOR2 (N9439, N9420, N7960);
and AND4 (N9440, N9409, N6448, N6696, N8743);
not NOT1 (N9441, N9438);
and AND4 (N9442, N9439, N2630, N2916, N2330);
or OR3 (N9443, N9437, N1888, N1213);
and AND2 (N9444, N9418, N1348);
not NOT1 (N9445, N9444);
xor XOR2 (N9446, N9435, N2975);
and AND3 (N9447, N9445, N8895, N6635);
and AND2 (N9448, N9436, N7503);
xor XOR2 (N9449, N9431, N8563);
or OR4 (N9450, N9449, N2190, N9183, N2253);
or OR3 (N9451, N9448, N3916, N3158);
and AND3 (N9452, N9451, N1073, N4500);
and AND2 (N9453, N9434, N3683);
xor XOR2 (N9454, N9452, N8743);
nor NOR2 (N9455, N9453, N8849);
xor XOR2 (N9456, N9441, N3270);
or OR2 (N9457, N9454, N4332);
or OR2 (N9458, N9456, N3856);
and AND3 (N9459, N9446, N6725, N252);
not NOT1 (N9460, N9459);
not NOT1 (N9461, N9450);
nand NAND4 (N9462, N9457, N7332, N2736, N6679);
buf BUF1 (N9463, N9461);
nand NAND3 (N9464, N9443, N5358, N2055);
not NOT1 (N9465, N9440);
nor NOR4 (N9466, N9442, N3947, N7281, N112);
nand NAND3 (N9467, N9463, N7127, N9340);
not NOT1 (N9468, N9462);
nand NAND3 (N9469, N9467, N2701, N4611);
not NOT1 (N9470, N9466);
nor NOR2 (N9471, N9430, N6128);
not NOT1 (N9472, N9455);
nand NAND4 (N9473, N9458, N2314, N8753, N3580);
nand NAND3 (N9474, N9447, N2121, N8550);
not NOT1 (N9475, N9465);
nand NAND2 (N9476, N9464, N5355);
xor XOR2 (N9477, N9472, N7924);
not NOT1 (N9478, N9471);
nand NAND4 (N9479, N9469, N1323, N609, N7399);
and AND3 (N9480, N9477, N4515, N2903);
buf BUF1 (N9481, N9476);
and AND3 (N9482, N9473, N9445, N8315);
not NOT1 (N9483, N9482);
buf BUF1 (N9484, N9479);
xor XOR2 (N9485, N9480, N3685);
and AND2 (N9486, N9481, N8141);
buf BUF1 (N9487, N9460);
not NOT1 (N9488, N9483);
and AND2 (N9489, N9484, N6514);
and AND4 (N9490, N9488, N6439, N1320, N7356);
not NOT1 (N9491, N9474);
buf BUF1 (N9492, N9468);
nor NOR2 (N9493, N9478, N531);
nand NAND4 (N9494, N9486, N6469, N4933, N3840);
or OR2 (N9495, N9485, N6548);
not NOT1 (N9496, N9495);
nor NOR3 (N9497, N9490, N8703, N1245);
buf BUF1 (N9498, N9475);
nand NAND4 (N9499, N9494, N704, N3067, N2524);
and AND2 (N9500, N9492, N3242);
not NOT1 (N9501, N9489);
or OR2 (N9502, N9501, N2485);
not NOT1 (N9503, N9502);
xor XOR2 (N9504, N9493, N8364);
buf BUF1 (N9505, N9497);
nor NOR4 (N9506, N9503, N1445, N396, N3833);
nor NOR2 (N9507, N9491, N6893);
xor XOR2 (N9508, N9496, N5739);
buf BUF1 (N9509, N9470);
xor XOR2 (N9510, N9487, N963);
or OR2 (N9511, N9504, N4488);
nor NOR4 (N9512, N9500, N3409, N8708, N7297);
xor XOR2 (N9513, N9506, N4806);
nor NOR3 (N9514, N9513, N2886, N759);
xor XOR2 (N9515, N9507, N1104);
and AND4 (N9516, N9510, N8513, N1318, N8451);
nand NAND4 (N9517, N9516, N2259, N7901, N1174);
nand NAND3 (N9518, N9508, N312, N4866);
nand NAND2 (N9519, N9505, N7614);
xor XOR2 (N9520, N9515, N5042);
nor NOR2 (N9521, N9519, N6147);
nor NOR2 (N9522, N9498, N7193);
buf BUF1 (N9523, N9509);
or OR3 (N9524, N9499, N6753, N3550);
nor NOR4 (N9525, N9511, N4825, N995, N4674);
not NOT1 (N9526, N9524);
not NOT1 (N9527, N9522);
nor NOR4 (N9528, N9514, N423, N9327, N818);
buf BUF1 (N9529, N9518);
xor XOR2 (N9530, N9529, N7079);
xor XOR2 (N9531, N9525, N2432);
nor NOR4 (N9532, N9527, N8182, N4548, N7956);
not NOT1 (N9533, N9523);
buf BUF1 (N9534, N9533);
or OR3 (N9535, N9532, N7272, N3124);
xor XOR2 (N9536, N9530, N2529);
nand NAND3 (N9537, N9534, N7971, N6949);
buf BUF1 (N9538, N9535);
buf BUF1 (N9539, N9538);
nor NOR2 (N9540, N9537, N8816);
and AND3 (N9541, N9531, N3493, N4653);
xor XOR2 (N9542, N9512, N4873);
buf BUF1 (N9543, N9521);
nor NOR4 (N9544, N9528, N7342, N6199, N2717);
or OR2 (N9545, N9540, N249);
nand NAND3 (N9546, N9520, N1935, N6034);
and AND4 (N9547, N9545, N5753, N9499, N2284);
buf BUF1 (N9548, N9542);
nor NOR2 (N9549, N9541, N4870);
nor NOR4 (N9550, N9517, N7413, N2192, N8191);
nand NAND4 (N9551, N9526, N1500, N8952, N7520);
nor NOR2 (N9552, N9544, N1182);
nand NAND4 (N9553, N9536, N9118, N9067, N7494);
nand NAND4 (N9554, N9543, N8923, N7029, N2003);
nor NOR3 (N9555, N9539, N9338, N4151);
not NOT1 (N9556, N9550);
or OR4 (N9557, N9552, N4467, N5091, N3688);
nand NAND3 (N9558, N9549, N8971, N2768);
xor XOR2 (N9559, N9555, N6605);
nand NAND4 (N9560, N9557, N1026, N1965, N3350);
and AND4 (N9561, N9553, N3053, N7733, N3078);
nand NAND2 (N9562, N9551, N2730);
and AND3 (N9563, N9554, N9006, N7094);
xor XOR2 (N9564, N9561, N5654);
or OR4 (N9565, N9560, N4737, N2542, N8871);
or OR4 (N9566, N9564, N6546, N2760, N9464);
xor XOR2 (N9567, N9565, N703);
or OR3 (N9568, N9558, N5278, N6463);
buf BUF1 (N9569, N9548);
or OR4 (N9570, N9568, N7397, N97, N8733);
buf BUF1 (N9571, N9563);
buf BUF1 (N9572, N9562);
nor NOR4 (N9573, N9566, N8397, N1833, N5613);
nand NAND4 (N9574, N9556, N8852, N8860, N3515);
xor XOR2 (N9575, N9547, N3127);
buf BUF1 (N9576, N9570);
or OR3 (N9577, N9572, N1201, N9282);
xor XOR2 (N9578, N9574, N9199);
nand NAND2 (N9579, N9578, N2504);
not NOT1 (N9580, N9571);
or OR4 (N9581, N9559, N2803, N2882, N2630);
and AND3 (N9582, N9567, N345, N6064);
nand NAND3 (N9583, N9577, N6009, N268);
not NOT1 (N9584, N9581);
xor XOR2 (N9585, N9569, N6083);
buf BUF1 (N9586, N9575);
and AND3 (N9587, N9586, N7280, N2375);
or OR3 (N9588, N9573, N6289, N8127);
not NOT1 (N9589, N9546);
or OR3 (N9590, N9587, N2716, N4159);
and AND2 (N9591, N9589, N5302);
and AND2 (N9592, N9576, N3050);
or OR4 (N9593, N9584, N9581, N8377, N6591);
not NOT1 (N9594, N9582);
buf BUF1 (N9595, N9592);
nor NOR3 (N9596, N9588, N5985, N2440);
nand NAND4 (N9597, N9596, N8617, N1783, N2127);
or OR2 (N9598, N9593, N3559);
nor NOR3 (N9599, N9590, N2820, N9471);
nand NAND4 (N9600, N9597, N8880, N352, N7733);
buf BUF1 (N9601, N9583);
nand NAND4 (N9602, N9594, N8002, N5589, N1254);
nor NOR2 (N9603, N9591, N1057);
or OR4 (N9604, N9595, N7972, N7356, N1078);
or OR3 (N9605, N9604, N991, N8899);
nand NAND4 (N9606, N9598, N5950, N1721, N6356);
not NOT1 (N9607, N9606);
nor NOR4 (N9608, N9585, N8637, N7936, N895);
buf BUF1 (N9609, N9605);
and AND4 (N9610, N9603, N2855, N7570, N9251);
and AND4 (N9611, N9610, N2156, N4916, N2467);
buf BUF1 (N9612, N9580);
not NOT1 (N9613, N9579);
nand NAND3 (N9614, N9607, N9340, N8209);
xor XOR2 (N9615, N9613, N1882);
buf BUF1 (N9616, N9601);
nor NOR4 (N9617, N9615, N8228, N4372, N7476);
and AND3 (N9618, N9600, N8162, N9323);
nor NOR2 (N9619, N9611, N9204);
and AND3 (N9620, N9616, N3436, N8967);
nand NAND3 (N9621, N9617, N9035, N6046);
and AND4 (N9622, N9612, N6808, N4549, N2665);
not NOT1 (N9623, N9622);
and AND4 (N9624, N9621, N7568, N6242, N9423);
nor NOR4 (N9625, N9599, N4308, N9263, N2519);
not NOT1 (N9626, N9618);
nand NAND2 (N9627, N9623, N2338);
not NOT1 (N9628, N9625);
xor XOR2 (N9629, N9608, N9225);
or OR2 (N9630, N9609, N6530);
xor XOR2 (N9631, N9614, N8506);
nand NAND3 (N9632, N9630, N4060, N6479);
xor XOR2 (N9633, N9626, N5634);
nor NOR4 (N9634, N9627, N4462, N6982, N4456);
xor XOR2 (N9635, N9624, N1204);
nor NOR4 (N9636, N9634, N2947, N2954, N3051);
not NOT1 (N9637, N9602);
nor NOR4 (N9638, N9633, N3794, N644, N767);
nor NOR3 (N9639, N9619, N2440, N4733);
nand NAND4 (N9640, N9638, N1270, N5982, N8520);
nand NAND4 (N9641, N9640, N5441, N3552, N3672);
not NOT1 (N9642, N9639);
nor NOR3 (N9643, N9636, N5951, N4904);
or OR2 (N9644, N9628, N5041);
and AND4 (N9645, N9642, N5250, N8068, N5764);
or OR4 (N9646, N9631, N4779, N6688, N1114);
or OR4 (N9647, N9645, N1287, N805, N2575);
or OR4 (N9648, N9643, N6029, N5730, N5367);
or OR4 (N9649, N9641, N3294, N3907, N2164);
and AND3 (N9650, N9637, N4743, N3434);
nor NOR2 (N9651, N9629, N1540);
nor NOR4 (N9652, N9651, N5504, N814, N29);
and AND3 (N9653, N9632, N4253, N530);
buf BUF1 (N9654, N9653);
xor XOR2 (N9655, N9647, N7595);
and AND4 (N9656, N9650, N1141, N4228, N5170);
nand NAND3 (N9657, N9656, N4208, N8229);
or OR4 (N9658, N9620, N5198, N5691, N9590);
nor NOR2 (N9659, N9648, N6495);
or OR4 (N9660, N9644, N411, N6971, N7775);
not NOT1 (N9661, N9652);
nand NAND2 (N9662, N9657, N2382);
and AND4 (N9663, N9660, N9479, N1592, N2816);
not NOT1 (N9664, N9649);
nand NAND3 (N9665, N9662, N459, N8083);
nand NAND2 (N9666, N9663, N1024);
nor NOR3 (N9667, N9658, N1621, N1057);
buf BUF1 (N9668, N9661);
nor NOR4 (N9669, N9666, N2491, N1005, N3951);
not NOT1 (N9670, N9646);
nand NAND3 (N9671, N9670, N4161, N2888);
or OR3 (N9672, N9654, N7537, N8630);
buf BUF1 (N9673, N9668);
buf BUF1 (N9674, N9655);
nand NAND2 (N9675, N9673, N1602);
nand NAND2 (N9676, N9664, N7230);
nor NOR2 (N9677, N9674, N6917);
buf BUF1 (N9678, N9675);
or OR4 (N9679, N9672, N5410, N136, N3878);
buf BUF1 (N9680, N9671);
nor NOR3 (N9681, N9669, N690, N1716);
not NOT1 (N9682, N9680);
and AND2 (N9683, N9679, N1544);
or OR3 (N9684, N9681, N414, N1120);
xor XOR2 (N9685, N9684, N2765);
buf BUF1 (N9686, N9635);
nor NOR3 (N9687, N9659, N3993, N5809);
or OR3 (N9688, N9686, N8287, N1464);
nor NOR3 (N9689, N9678, N2751, N171);
not NOT1 (N9690, N9667);
or OR3 (N9691, N9690, N4738, N2025);
buf BUF1 (N9692, N9691);
nor NOR2 (N9693, N9688, N6584);
nand NAND4 (N9694, N9693, N1551, N4298, N6588);
or OR2 (N9695, N9682, N8577);
xor XOR2 (N9696, N9695, N6410);
xor XOR2 (N9697, N9696, N7272);
and AND3 (N9698, N9677, N6316, N4763);
or OR2 (N9699, N9697, N331);
nand NAND4 (N9700, N9676, N1069, N874, N2192);
nor NOR4 (N9701, N9699, N9140, N293, N1539);
nor NOR2 (N9702, N9701, N7807);
nor NOR2 (N9703, N9687, N3107);
nor NOR3 (N9704, N9692, N3360, N4721);
nand NAND2 (N9705, N9703, N4187);
not NOT1 (N9706, N9705);
nor NOR2 (N9707, N9698, N9032);
nand NAND4 (N9708, N9694, N6339, N6907, N5081);
nor NOR2 (N9709, N9702, N3981);
and AND4 (N9710, N9709, N5864, N3833, N5079);
or OR2 (N9711, N9708, N9488);
buf BUF1 (N9712, N9710);
buf BUF1 (N9713, N9712);
or OR2 (N9714, N9711, N7008);
or OR4 (N9715, N9665, N7816, N4396, N8576);
nand NAND3 (N9716, N9685, N972, N8273);
not NOT1 (N9717, N9704);
not NOT1 (N9718, N9714);
or OR2 (N9719, N9716, N9340);
nor NOR3 (N9720, N9718, N9475, N6485);
not NOT1 (N9721, N9713);
not NOT1 (N9722, N9689);
xor XOR2 (N9723, N9683, N821);
not NOT1 (N9724, N9719);
nand NAND2 (N9725, N9706, N6015);
and AND3 (N9726, N9720, N5163, N2965);
xor XOR2 (N9727, N9726, N2712);
nor NOR4 (N9728, N9725, N295, N6292, N1203);
buf BUF1 (N9729, N9721);
nor NOR3 (N9730, N9723, N9026, N6834);
xor XOR2 (N9731, N9717, N3863);
nor NOR3 (N9732, N9700, N4555, N1941);
or OR3 (N9733, N9727, N8577, N1146);
not NOT1 (N9734, N9728);
buf BUF1 (N9735, N9732);
not NOT1 (N9736, N9730);
nor NOR3 (N9737, N9715, N2195, N9699);
nand NAND3 (N9738, N9731, N4170, N1436);
or OR2 (N9739, N9734, N7786);
buf BUF1 (N9740, N9739);
or OR4 (N9741, N9722, N8340, N1978, N5547);
or OR3 (N9742, N9741, N2435, N8409);
xor XOR2 (N9743, N9735, N303);
xor XOR2 (N9744, N9724, N2138);
or OR4 (N9745, N9740, N773, N6666, N6651);
nor NOR4 (N9746, N9742, N1509, N3139, N4963);
or OR4 (N9747, N9733, N7614, N3759, N7220);
not NOT1 (N9748, N9743);
buf BUF1 (N9749, N9745);
buf BUF1 (N9750, N9736);
nor NOR2 (N9751, N9748, N4280);
nand NAND4 (N9752, N9737, N5800, N4144, N3230);
nor NOR3 (N9753, N9738, N6636, N5163);
and AND2 (N9754, N9729, N8025);
not NOT1 (N9755, N9754);
nor NOR4 (N9756, N9744, N1483, N3749, N8713);
nand NAND2 (N9757, N9755, N338);
and AND3 (N9758, N9753, N9288, N6228);
and AND3 (N9759, N9707, N8844, N5359);
buf BUF1 (N9760, N9749);
or OR2 (N9761, N9752, N4535);
nor NOR4 (N9762, N9756, N5568, N144, N1502);
xor XOR2 (N9763, N9759, N127);
or OR2 (N9764, N9750, N6299);
and AND4 (N9765, N9764, N8446, N9044, N4539);
not NOT1 (N9766, N9762);
nand NAND2 (N9767, N9758, N2418);
buf BUF1 (N9768, N9757);
not NOT1 (N9769, N9751);
xor XOR2 (N9770, N9766, N2993);
and AND4 (N9771, N9765, N7232, N634, N8931);
xor XOR2 (N9772, N9761, N5349);
xor XOR2 (N9773, N9770, N4863);
or OR3 (N9774, N9768, N7410, N9283);
not NOT1 (N9775, N9763);
nor NOR2 (N9776, N9774, N5140);
or OR4 (N9777, N9775, N9014, N1472, N546);
and AND4 (N9778, N9746, N3716, N459, N5406);
buf BUF1 (N9779, N9777);
buf BUF1 (N9780, N9771);
and AND2 (N9781, N9760, N1456);
and AND2 (N9782, N9781, N360);
nand NAND2 (N9783, N9747, N688);
and AND3 (N9784, N9776, N8713, N3299);
buf BUF1 (N9785, N9783);
or OR2 (N9786, N9784, N8370);
not NOT1 (N9787, N9780);
or OR4 (N9788, N9779, N3197, N8041, N2547);
not NOT1 (N9789, N9778);
buf BUF1 (N9790, N9772);
and AND2 (N9791, N9773, N4121);
nor NOR3 (N9792, N9787, N1889, N9435);
xor XOR2 (N9793, N9767, N9628);
and AND2 (N9794, N9789, N7499);
buf BUF1 (N9795, N9786);
or OR3 (N9796, N9769, N3726, N2152);
nor NOR2 (N9797, N9792, N2506);
buf BUF1 (N9798, N9793);
not NOT1 (N9799, N9790);
nor NOR3 (N9800, N9785, N8068, N8659);
nand NAND2 (N9801, N9799, N1242);
and AND3 (N9802, N9791, N2687, N5629);
or OR2 (N9803, N9797, N3281);
not NOT1 (N9804, N9802);
nor NOR4 (N9805, N9798, N8540, N1498, N6329);
nor NOR3 (N9806, N9794, N5284, N779);
or OR3 (N9807, N9788, N9168, N9744);
nand NAND2 (N9808, N9805, N8290);
or OR4 (N9809, N9782, N9366, N2667, N7366);
nand NAND4 (N9810, N9801, N1732, N7074, N633);
not NOT1 (N9811, N9800);
not NOT1 (N9812, N9795);
not NOT1 (N9813, N9807);
or OR2 (N9814, N9808, N3711);
buf BUF1 (N9815, N9804);
buf BUF1 (N9816, N9812);
nand NAND3 (N9817, N9814, N3985, N7327);
or OR4 (N9818, N9796, N857, N511, N1017);
not NOT1 (N9819, N9806);
buf BUF1 (N9820, N9816);
nor NOR4 (N9821, N9817, N8629, N8031, N4625);
xor XOR2 (N9822, N9819, N5143);
not NOT1 (N9823, N9821);
and AND4 (N9824, N9815, N8716, N8643, N505);
xor XOR2 (N9825, N9809, N8728);
and AND3 (N9826, N9811, N6767, N7742);
and AND2 (N9827, N9810, N5585);
nand NAND4 (N9828, N9825, N5257, N8649, N586);
and AND4 (N9829, N9820, N3115, N4381, N7726);
nor NOR2 (N9830, N9813, N4199);
buf BUF1 (N9831, N9824);
not NOT1 (N9832, N9827);
and AND3 (N9833, N9828, N7701, N8535);
not NOT1 (N9834, N9803);
nand NAND2 (N9835, N9833, N2091);
xor XOR2 (N9836, N9822, N8392);
or OR2 (N9837, N9834, N8044);
nor NOR2 (N9838, N9837, N7023);
nand NAND3 (N9839, N9835, N4075, N5217);
or OR3 (N9840, N9838, N7094, N820);
nor NOR3 (N9841, N9818, N5703, N1419);
nor NOR3 (N9842, N9832, N7204, N7291);
buf BUF1 (N9843, N9842);
nor NOR4 (N9844, N9836, N1719, N7973, N3086);
buf BUF1 (N9845, N9831);
buf BUF1 (N9846, N9844);
or OR3 (N9847, N9843, N4937, N9306);
or OR2 (N9848, N9840, N1984);
and AND4 (N9849, N9841, N6869, N8990, N7930);
nor NOR4 (N9850, N9839, N3677, N6987, N229);
xor XOR2 (N9851, N9846, N4399);
nor NOR3 (N9852, N9851, N7139, N5334);
xor XOR2 (N9853, N9852, N1832);
xor XOR2 (N9854, N9848, N1512);
or OR4 (N9855, N9853, N2775, N7730, N608);
not NOT1 (N9856, N9849);
nand NAND2 (N9857, N9830, N8145);
nand NAND4 (N9858, N9845, N6643, N9820, N2112);
not NOT1 (N9859, N9823);
and AND3 (N9860, N9855, N6132, N6356);
or OR4 (N9861, N9847, N6210, N1233, N740);
nand NAND3 (N9862, N9850, N934, N4351);
xor XOR2 (N9863, N9861, N6733);
or OR4 (N9864, N9859, N1664, N236, N6173);
xor XOR2 (N9865, N9858, N7530);
xor XOR2 (N9866, N9854, N4149);
nand NAND4 (N9867, N9865, N5523, N6624, N9534);
nor NOR4 (N9868, N9867, N7693, N1916, N8447);
or OR4 (N9869, N9856, N6484, N413, N3927);
nand NAND4 (N9870, N9864, N3832, N5085, N1311);
or OR4 (N9871, N9826, N3218, N1547, N129);
nand NAND4 (N9872, N9866, N2394, N3205, N6754);
buf BUF1 (N9873, N9870);
nand NAND2 (N9874, N9829, N3792);
not NOT1 (N9875, N9869);
xor XOR2 (N9876, N9860, N230);
nand NAND3 (N9877, N9863, N6500, N7499);
not NOT1 (N9878, N9877);
or OR3 (N9879, N9876, N280, N1516);
buf BUF1 (N9880, N9874);
and AND4 (N9881, N9875, N4836, N8082, N9284);
nand NAND4 (N9882, N9868, N7343, N5248, N7995);
or OR4 (N9883, N9862, N7382, N6592, N3885);
nand NAND4 (N9884, N9879, N6245, N1023, N6660);
or OR4 (N9885, N9882, N3221, N2080, N5035);
or OR2 (N9886, N9873, N8697);
buf BUF1 (N9887, N9878);
not NOT1 (N9888, N9871);
or OR4 (N9889, N9885, N208, N4530, N1995);
nand NAND3 (N9890, N9881, N5002, N6117);
and AND2 (N9891, N9872, N1989);
and AND3 (N9892, N9883, N440, N6051);
buf BUF1 (N9893, N9889);
nor NOR4 (N9894, N9857, N1347, N6506, N8058);
nand NAND2 (N9895, N9890, N1468);
not NOT1 (N9896, N9894);
nor NOR2 (N9897, N9892, N8916);
not NOT1 (N9898, N9896);
not NOT1 (N9899, N9891);
xor XOR2 (N9900, N9886, N5410);
and AND2 (N9901, N9880, N5260);
not NOT1 (N9902, N9897);
nor NOR2 (N9903, N9887, N4228);
xor XOR2 (N9904, N9903, N5831);
xor XOR2 (N9905, N9902, N8282);
or OR2 (N9906, N9900, N5274);
buf BUF1 (N9907, N9893);
nor NOR2 (N9908, N9907, N8696);
xor XOR2 (N9909, N9888, N1229);
nand NAND4 (N9910, N9895, N7763, N9566, N4389);
not NOT1 (N9911, N9899);
nand NAND3 (N9912, N9910, N3547, N2173);
buf BUF1 (N9913, N9908);
xor XOR2 (N9914, N9898, N4740);
or OR3 (N9915, N9904, N1778, N1293);
nand NAND3 (N9916, N9914, N1343, N3158);
or OR2 (N9917, N9911, N609);
or OR2 (N9918, N9906, N6653);
not NOT1 (N9919, N9917);
nand NAND3 (N9920, N9912, N9490, N8039);
nand NAND3 (N9921, N9916, N4956, N7915);
xor XOR2 (N9922, N9913, N1090);
buf BUF1 (N9923, N9922);
not NOT1 (N9924, N9919);
and AND3 (N9925, N9918, N5712, N4297);
buf BUF1 (N9926, N9901);
not NOT1 (N9927, N9915);
and AND3 (N9928, N9920, N7127, N2119);
and AND2 (N9929, N9927, N2428);
nand NAND2 (N9930, N9905, N4022);
nor NOR2 (N9931, N9930, N4690);
nand NAND4 (N9932, N9926, N8254, N5264, N5401);
not NOT1 (N9933, N9924);
buf BUF1 (N9934, N9929);
xor XOR2 (N9935, N9933, N5789);
nor NOR4 (N9936, N9928, N1591, N8658, N8272);
and AND2 (N9937, N9936, N9089);
or OR4 (N9938, N9931, N6433, N8589, N7062);
buf BUF1 (N9939, N9923);
nand NAND3 (N9940, N9937, N6423, N3398);
xor XOR2 (N9941, N9938, N7972);
not NOT1 (N9942, N9935);
nand NAND3 (N9943, N9932, N8482, N3798);
and AND3 (N9944, N9942, N2843, N7053);
nor NOR3 (N9945, N9921, N3670, N9802);
nor NOR4 (N9946, N9944, N6910, N4381, N9628);
buf BUF1 (N9947, N9909);
or OR3 (N9948, N9947, N2920, N12);
and AND3 (N9949, N9943, N4421, N584);
or OR4 (N9950, N9946, N5134, N4027, N6556);
buf BUF1 (N9951, N9941);
nor NOR3 (N9952, N9950, N5316, N7349);
buf BUF1 (N9953, N9939);
xor XOR2 (N9954, N9951, N4820);
xor XOR2 (N9955, N9940, N9921);
xor XOR2 (N9956, N9925, N137);
buf BUF1 (N9957, N9953);
not NOT1 (N9958, N9954);
and AND4 (N9959, N9945, N3855, N7418, N1113);
nor NOR3 (N9960, N9959, N7116, N4193);
xor XOR2 (N9961, N9958, N4562);
nand NAND3 (N9962, N9884, N1254, N7500);
buf BUF1 (N9963, N9957);
xor XOR2 (N9964, N9955, N9850);
nor NOR3 (N9965, N9964, N5790, N5620);
and AND4 (N9966, N9948, N6451, N7039, N195);
or OR3 (N9967, N9962, N9029, N8638);
nor NOR2 (N9968, N9965, N1615);
and AND3 (N9969, N9949, N5507, N6609);
buf BUF1 (N9970, N9968);
and AND3 (N9971, N9952, N8547, N6309);
or OR2 (N9972, N9966, N1880);
and AND4 (N9973, N9969, N9927, N5023, N8145);
xor XOR2 (N9974, N9956, N5200);
nor NOR2 (N9975, N9934, N4198);
or OR2 (N9976, N9960, N3272);
nor NOR2 (N9977, N9973, N7824);
xor XOR2 (N9978, N9977, N7217);
or OR4 (N9979, N9963, N5594, N8625, N5945);
xor XOR2 (N9980, N9971, N852);
nor NOR3 (N9981, N9976, N4208, N9057);
xor XOR2 (N9982, N9974, N3143);
nand NAND3 (N9983, N9980, N1375, N7936);
xor XOR2 (N9984, N9979, N358);
xor XOR2 (N9985, N9978, N2875);
buf BUF1 (N9986, N9983);
or OR4 (N9987, N9975, N893, N7662, N1131);
buf BUF1 (N9988, N9986);
buf BUF1 (N9989, N9985);
not NOT1 (N9990, N9981);
and AND4 (N9991, N9967, N3918, N8676, N9344);
nor NOR2 (N9992, N9982, N5664);
nor NOR4 (N9993, N9991, N1606, N2011, N6600);
buf BUF1 (N9994, N9987);
xor XOR2 (N9995, N9984, N7017);
buf BUF1 (N9996, N9972);
buf BUF1 (N9997, N9961);
nand NAND2 (N9998, N9996, N7839);
buf BUF1 (N9999, N9997);
nor NOR4 (N10000, N9999, N195, N6896, N8689);
xor XOR2 (N10001, N9988, N8807);
xor XOR2 (N10002, N9992, N5880);
or OR3 (N10003, N10000, N1624, N7968);
nor NOR4 (N10004, N9970, N7595, N8025, N1407);
nand NAND2 (N10005, N10002, N9855);
xor XOR2 (N10006, N10004, N6091);
nand NAND4 (N10007, N10006, N2194, N3567, N6555);
nor NOR4 (N10008, N9990, N7801, N3857, N834);
nor NOR2 (N10009, N10003, N1829);
and AND3 (N10010, N9989, N6593, N3764);
buf BUF1 (N10011, N10005);
xor XOR2 (N10012, N9994, N926);
nand NAND3 (N10013, N10010, N3035, N9193);
xor XOR2 (N10014, N9998, N1794);
buf BUF1 (N10015, N10009);
or OR4 (N10016, N9993, N8409, N3527, N7060);
not NOT1 (N10017, N10016);
nand NAND2 (N10018, N10008, N4383);
not NOT1 (N10019, N10011);
buf BUF1 (N10020, N9995);
not NOT1 (N10021, N10019);
not NOT1 (N10022, N10001);
buf BUF1 (N10023, N10014);
xor XOR2 (N10024, N10012, N341);
or OR4 (N10025, N10023, N8916, N7993, N6967);
nand NAND2 (N10026, N10024, N505);
xor XOR2 (N10027, N10017, N7393);
and AND2 (N10028, N10018, N444);
nor NOR4 (N10029, N10021, N2592, N1856, N8107);
not NOT1 (N10030, N10027);
nor NOR4 (N10031, N10015, N7780, N2904, N3765);
or OR4 (N10032, N10029, N4165, N7341, N5127);
not NOT1 (N10033, N10026);
xor XOR2 (N10034, N10013, N9319);
xor XOR2 (N10035, N10022, N8735);
nor NOR3 (N10036, N10034, N9976, N9874);
or OR3 (N10037, N10025, N1522, N3366);
nor NOR2 (N10038, N10007, N8821);
nand NAND4 (N10039, N10037, N9517, N2574, N9194);
nor NOR3 (N10040, N10036, N7330, N1398);
buf BUF1 (N10041, N10033);
buf BUF1 (N10042, N10039);
nand NAND2 (N10043, N10030, N9852);
nand NAND2 (N10044, N10038, N6902);
not NOT1 (N10045, N10040);
or OR2 (N10046, N10032, N7064);
buf BUF1 (N10047, N10035);
nand NAND2 (N10048, N10047, N9413);
xor XOR2 (N10049, N10045, N3695);
nand NAND2 (N10050, N10044, N3888);
or OR4 (N10051, N10046, N4247, N5002, N8795);
nand NAND4 (N10052, N10049, N9249, N6659, N3050);
buf BUF1 (N10053, N10050);
buf BUF1 (N10054, N10051);
and AND3 (N10055, N10042, N1165, N6862);
buf BUF1 (N10056, N10028);
and AND3 (N10057, N10048, N470, N1220);
xor XOR2 (N10058, N10031, N3665);
nor NOR4 (N10059, N10053, N3505, N6354, N1370);
and AND4 (N10060, N10020, N2872, N5974, N9737);
nand NAND2 (N10061, N10054, N2917);
xor XOR2 (N10062, N10057, N6193);
nor NOR3 (N10063, N10043, N6776, N5545);
and AND4 (N10064, N10056, N8942, N5347, N7981);
xor XOR2 (N10065, N10063, N6090);
nand NAND2 (N10066, N10062, N4786);
and AND3 (N10067, N10061, N7660, N7475);
not NOT1 (N10068, N10058);
nor NOR3 (N10069, N10068, N458, N620);
nand NAND2 (N10070, N10064, N7040);
not NOT1 (N10071, N10055);
or OR3 (N10072, N10052, N2147, N449);
nor NOR2 (N10073, N10041, N4312);
nor NOR2 (N10074, N10071, N2665);
buf BUF1 (N10075, N10074);
buf BUF1 (N10076, N10072);
nor NOR2 (N10077, N10067, N528);
nand NAND3 (N10078, N10066, N6794, N3154);
nor NOR4 (N10079, N10059, N1119, N4632, N9008);
xor XOR2 (N10080, N10060, N9748);
nor NOR2 (N10081, N10079, N6630);
buf BUF1 (N10082, N10075);
and AND2 (N10083, N10069, N3013);
or OR2 (N10084, N10083, N468);
or OR4 (N10085, N10073, N6965, N5861, N6326);
nand NAND4 (N10086, N10085, N9667, N3088, N7047);
buf BUF1 (N10087, N10070);
nand NAND4 (N10088, N10080, N1539, N6529, N6343);
or OR2 (N10089, N10065, N824);
buf BUF1 (N10090, N10089);
nand NAND4 (N10091, N10090, N3768, N8149, N7503);
not NOT1 (N10092, N10082);
or OR2 (N10093, N10077, N8902);
buf BUF1 (N10094, N10081);
xor XOR2 (N10095, N10086, N4739);
nand NAND4 (N10096, N10094, N3455, N4968, N4567);
and AND2 (N10097, N10087, N1565);
nor NOR3 (N10098, N10078, N4434, N9602);
xor XOR2 (N10099, N10092, N6754);
or OR3 (N10100, N10091, N7640, N7251);
and AND3 (N10101, N10096, N4407, N6603);
nand NAND4 (N10102, N10093, N3105, N2680, N6487);
not NOT1 (N10103, N10100);
or OR4 (N10104, N10097, N2104, N7362, N4430);
or OR2 (N10105, N10104, N6827);
xor XOR2 (N10106, N10076, N6201);
nor NOR3 (N10107, N10106, N5709, N3889);
buf BUF1 (N10108, N10088);
or OR4 (N10109, N10099, N2299, N5590, N4733);
not NOT1 (N10110, N10103);
xor XOR2 (N10111, N10102, N9441);
nand NAND2 (N10112, N10095, N9729);
buf BUF1 (N10113, N10107);
nand NAND2 (N10114, N10112, N4953);
or OR3 (N10115, N10108, N5266, N114);
or OR2 (N10116, N10115, N4020);
not NOT1 (N10117, N10111);
xor XOR2 (N10118, N10110, N7527);
not NOT1 (N10119, N10118);
xor XOR2 (N10120, N10113, N6938);
and AND3 (N10121, N10117, N4200, N5571);
nand NAND4 (N10122, N10098, N9174, N5653, N7529);
xor XOR2 (N10123, N10084, N2457);
xor XOR2 (N10124, N10122, N2400);
nand NAND4 (N10125, N10101, N41, N9768, N8707);
not NOT1 (N10126, N10120);
buf BUF1 (N10127, N10116);
nand NAND2 (N10128, N10114, N6628);
nand NAND4 (N10129, N10127, N4510, N7073, N6641);
not NOT1 (N10130, N10126);
buf BUF1 (N10131, N10105);
xor XOR2 (N10132, N10119, N9102);
xor XOR2 (N10133, N10130, N4042);
or OR4 (N10134, N10129, N6226, N7651, N1765);
nand NAND2 (N10135, N10124, N4453);
buf BUF1 (N10136, N10121);
nand NAND4 (N10137, N10133, N7039, N9848, N239);
not NOT1 (N10138, N10132);
xor XOR2 (N10139, N10125, N6941);
xor XOR2 (N10140, N10134, N9693);
and AND3 (N10141, N10123, N5714, N7340);
or OR2 (N10142, N10109, N7670);
nand NAND4 (N10143, N10139, N5700, N5744, N8755);
nand NAND4 (N10144, N10143, N3979, N2133, N9152);
xor XOR2 (N10145, N10128, N7746);
or OR2 (N10146, N10137, N9318);
not NOT1 (N10147, N10146);
and AND4 (N10148, N10131, N2068, N5443, N35);
or OR2 (N10149, N10136, N3963);
or OR4 (N10150, N10140, N1856, N508, N9757);
buf BUF1 (N10151, N10138);
or OR3 (N10152, N10135, N5983, N1658);
nor NOR2 (N10153, N10148, N1369);
buf BUF1 (N10154, N10144);
or OR2 (N10155, N10152, N769);
or OR2 (N10156, N10142, N2898);
nand NAND2 (N10157, N10145, N541);
buf BUF1 (N10158, N10151);
xor XOR2 (N10159, N10147, N8834);
xor XOR2 (N10160, N10153, N7682);
buf BUF1 (N10161, N10156);
and AND4 (N10162, N10159, N3052, N6503, N5435);
and AND3 (N10163, N10158, N6782, N9708);
nor NOR4 (N10164, N10149, N6164, N2576, N1130);
or OR4 (N10165, N10164, N2311, N3538, N8742);
buf BUF1 (N10166, N10162);
nor NOR2 (N10167, N10150, N2284);
nor NOR4 (N10168, N10161, N6752, N8822, N1124);
buf BUF1 (N10169, N10157);
or OR3 (N10170, N10169, N7541, N8959);
nor NOR2 (N10171, N10165, N2998);
not NOT1 (N10172, N10166);
nand NAND2 (N10173, N10160, N1758);
xor XOR2 (N10174, N10163, N7437);
buf BUF1 (N10175, N10155);
and AND3 (N10176, N10154, N2419, N5362);
or OR2 (N10177, N10170, N6084);
and AND3 (N10178, N10172, N5379, N9967);
xor XOR2 (N10179, N10167, N758);
nand NAND2 (N10180, N10174, N9335);
buf BUF1 (N10181, N10171);
buf BUF1 (N10182, N10141);
nand NAND3 (N10183, N10175, N3100, N8129);
nand NAND4 (N10184, N10168, N4318, N3730, N5000);
nor NOR4 (N10185, N10176, N8250, N3936, N924);
or OR3 (N10186, N10181, N2727, N4040);
nand NAND2 (N10187, N10185, N9688);
buf BUF1 (N10188, N10187);
buf BUF1 (N10189, N10173);
and AND2 (N10190, N10189, N1342);
and AND3 (N10191, N10183, N9337, N102);
nor NOR3 (N10192, N10190, N32, N1439);
and AND3 (N10193, N10182, N5449, N7166);
xor XOR2 (N10194, N10192, N6703);
buf BUF1 (N10195, N10178);
buf BUF1 (N10196, N10193);
and AND4 (N10197, N10195, N9929, N1858, N8233);
nand NAND2 (N10198, N10184, N3935);
or OR3 (N10199, N10196, N2119, N8392);
nand NAND2 (N10200, N10198, N9671);
not NOT1 (N10201, N10191);
buf BUF1 (N10202, N10201);
nor NOR3 (N10203, N10202, N9846, N4222);
not NOT1 (N10204, N10186);
and AND2 (N10205, N10180, N1800);
xor XOR2 (N10206, N10200, N4992);
buf BUF1 (N10207, N10203);
nor NOR4 (N10208, N10204, N3576, N8901, N9730);
nor NOR3 (N10209, N10208, N9929, N9936);
nand NAND4 (N10210, N10197, N8344, N6664, N9815);
buf BUF1 (N10211, N10179);
or OR3 (N10212, N10206, N4114, N9053);
xor XOR2 (N10213, N10210, N3326);
or OR2 (N10214, N10177, N4704);
and AND3 (N10215, N10213, N4626, N8474);
nor NOR4 (N10216, N10211, N8812, N1615, N6513);
nand NAND3 (N10217, N10199, N7942, N9284);
or OR2 (N10218, N10214, N1847);
and AND4 (N10219, N10212, N9239, N8989, N8494);
and AND4 (N10220, N10217, N8734, N2952, N3014);
nand NAND2 (N10221, N10188, N7082);
and AND4 (N10222, N10205, N8875, N3988, N2642);
buf BUF1 (N10223, N10216);
not NOT1 (N10224, N10220);
not NOT1 (N10225, N10224);
xor XOR2 (N10226, N10223, N4563);
xor XOR2 (N10227, N10207, N6688);
or OR3 (N10228, N10218, N6730, N8684);
nand NAND4 (N10229, N10228, N1597, N8811, N319);
buf BUF1 (N10230, N10219);
nand NAND4 (N10231, N10225, N1177, N3431, N4195);
not NOT1 (N10232, N10230);
buf BUF1 (N10233, N10194);
xor XOR2 (N10234, N10209, N2064);
or OR4 (N10235, N10233, N2256, N8392, N4431);
buf BUF1 (N10236, N10221);
or OR4 (N10237, N10227, N4687, N4236, N1836);
not NOT1 (N10238, N10232);
xor XOR2 (N10239, N10231, N593);
nor NOR2 (N10240, N10235, N2988);
buf BUF1 (N10241, N10236);
or OR4 (N10242, N10215, N6468, N607, N3273);
nand NAND2 (N10243, N10229, N9067);
or OR3 (N10244, N10238, N9434, N3261);
or OR2 (N10245, N10241, N10232);
xor XOR2 (N10246, N10226, N3165);
or OR2 (N10247, N10222, N9109);
not NOT1 (N10248, N10245);
buf BUF1 (N10249, N10237);
not NOT1 (N10250, N10240);
nor NOR4 (N10251, N10234, N5557, N5435, N1410);
buf BUF1 (N10252, N10250);
and AND4 (N10253, N10239, N6216, N949, N2666);
and AND2 (N10254, N10252, N587);
and AND3 (N10255, N10243, N7124, N7013);
nand NAND4 (N10256, N10247, N4619, N4695, N6735);
buf BUF1 (N10257, N10242);
and AND3 (N10258, N10251, N2998, N5756);
xor XOR2 (N10259, N10256, N4228);
buf BUF1 (N10260, N10249);
nor NOR2 (N10261, N10253, N3866);
buf BUF1 (N10262, N10248);
and AND3 (N10263, N10261, N8425, N7258);
xor XOR2 (N10264, N10263, N9631);
not NOT1 (N10265, N10258);
and AND2 (N10266, N10255, N5585);
not NOT1 (N10267, N10254);
nor NOR3 (N10268, N10244, N6580, N182);
not NOT1 (N10269, N10267);
buf BUF1 (N10270, N10266);
not NOT1 (N10271, N10264);
not NOT1 (N10272, N10257);
not NOT1 (N10273, N10271);
nand NAND4 (N10274, N10260, N2630, N1202, N4553);
buf BUF1 (N10275, N10262);
not NOT1 (N10276, N10274);
nor NOR2 (N10277, N10273, N3381);
nand NAND4 (N10278, N10246, N4529, N1831, N7401);
or OR2 (N10279, N10269, N5452);
xor XOR2 (N10280, N10265, N4330);
not NOT1 (N10281, N10275);
buf BUF1 (N10282, N10259);
and AND4 (N10283, N10280, N4991, N1067, N2050);
not NOT1 (N10284, N10276);
nand NAND2 (N10285, N10281, N433);
and AND2 (N10286, N10284, N1192);
nand NAND2 (N10287, N10268, N594);
not NOT1 (N10288, N10270);
and AND4 (N10289, N10277, N1489, N1563, N2813);
or OR4 (N10290, N10289, N9456, N9528, N1129);
or OR4 (N10291, N10285, N2816, N1582, N7701);
xor XOR2 (N10292, N10288, N118);
not NOT1 (N10293, N10286);
or OR2 (N10294, N10279, N8596);
and AND3 (N10295, N10291, N8498, N2466);
nor NOR2 (N10296, N10290, N1162);
not NOT1 (N10297, N10287);
and AND2 (N10298, N10282, N3162);
nand NAND3 (N10299, N10293, N7620, N1826);
xor XOR2 (N10300, N10292, N987);
nand NAND3 (N10301, N10278, N3000, N10125);
not NOT1 (N10302, N10294);
buf BUF1 (N10303, N10296);
nand NAND4 (N10304, N10299, N1129, N1961, N2836);
or OR4 (N10305, N10297, N4375, N6020, N3683);
xor XOR2 (N10306, N10272, N8698);
and AND3 (N10307, N10283, N1169, N9347);
nand NAND2 (N10308, N10303, N2741);
xor XOR2 (N10309, N10300, N2507);
or OR2 (N10310, N10306, N527);
and AND4 (N10311, N10305, N5200, N9875, N957);
or OR3 (N10312, N10302, N4300, N2909);
xor XOR2 (N10313, N10304, N3212);
not NOT1 (N10314, N10301);
nand NAND2 (N10315, N10308, N9054);
not NOT1 (N10316, N10315);
buf BUF1 (N10317, N10310);
xor XOR2 (N10318, N10314, N1438);
buf BUF1 (N10319, N10313);
or OR4 (N10320, N10309, N3634, N7785, N7268);
nand NAND2 (N10321, N10311, N4752);
nor NOR3 (N10322, N10321, N9135, N3195);
and AND2 (N10323, N10307, N5084);
xor XOR2 (N10324, N10322, N8885);
buf BUF1 (N10325, N10295);
not NOT1 (N10326, N10319);
or OR3 (N10327, N10317, N4682, N4302);
or OR3 (N10328, N10325, N2504, N3700);
xor XOR2 (N10329, N10324, N759);
not NOT1 (N10330, N10328);
not NOT1 (N10331, N10329);
or OR4 (N10332, N10330, N466, N8451, N3172);
nand NAND3 (N10333, N10332, N145, N7425);
and AND4 (N10334, N10333, N2775, N6958, N10319);
or OR2 (N10335, N10318, N4987);
nand NAND4 (N10336, N10320, N7735, N750, N3558);
nand NAND3 (N10337, N10326, N9922, N9062);
or OR4 (N10338, N10334, N8482, N4611, N4425);
not NOT1 (N10339, N10336);
nor NOR3 (N10340, N10338, N6153, N7636);
not NOT1 (N10341, N10316);
not NOT1 (N10342, N10339);
not NOT1 (N10343, N10335);
and AND4 (N10344, N10341, N9794, N6869, N6824);
buf BUF1 (N10345, N10337);
nand NAND2 (N10346, N10331, N6514);
nand NAND2 (N10347, N10346, N1440);
and AND3 (N10348, N10323, N5351, N595);
not NOT1 (N10349, N10347);
xor XOR2 (N10350, N10348, N10025);
xor XOR2 (N10351, N10343, N2301);
xor XOR2 (N10352, N10340, N1271);
buf BUF1 (N10353, N10342);
nor NOR2 (N10354, N10312, N2501);
nor NOR2 (N10355, N10298, N7301);
or OR2 (N10356, N10327, N2257);
or OR2 (N10357, N10344, N3324);
buf BUF1 (N10358, N10349);
and AND4 (N10359, N10353, N1148, N2838, N5347);
buf BUF1 (N10360, N10355);
nor NOR4 (N10361, N10357, N2380, N4127, N8413);
xor XOR2 (N10362, N10351, N6517);
buf BUF1 (N10363, N10362);
or OR4 (N10364, N10354, N1763, N4403, N8059);
nor NOR2 (N10365, N10359, N10066);
nand NAND4 (N10366, N10364, N6656, N5582, N6192);
nand NAND2 (N10367, N10363, N10194);
or OR3 (N10368, N10360, N387, N9134);
nor NOR2 (N10369, N10367, N75);
buf BUF1 (N10370, N10345);
buf BUF1 (N10371, N10352);
or OR4 (N10372, N10365, N5287, N5601, N10039);
nor NOR3 (N10373, N10350, N9504, N8271);
or OR3 (N10374, N10358, N3221, N8974);
or OR3 (N10375, N10373, N8402, N4793);
or OR4 (N10376, N10369, N7927, N4129, N1979);
xor XOR2 (N10377, N10376, N1356);
not NOT1 (N10378, N10370);
not NOT1 (N10379, N10375);
xor XOR2 (N10380, N10356, N2875);
and AND4 (N10381, N10368, N7983, N3990, N318);
and AND3 (N10382, N10381, N5193, N970);
nand NAND3 (N10383, N10378, N9271, N8143);
and AND2 (N10384, N10372, N3210);
not NOT1 (N10385, N10374);
buf BUF1 (N10386, N10385);
not NOT1 (N10387, N10382);
and AND4 (N10388, N10379, N4134, N8474, N9293);
xor XOR2 (N10389, N10380, N7901);
buf BUF1 (N10390, N10371);
nor NOR2 (N10391, N10361, N9416);
nor NOR2 (N10392, N10388, N931);
nand NAND4 (N10393, N10386, N2395, N1777, N3725);
buf BUF1 (N10394, N10387);
or OR4 (N10395, N10391, N2978, N9446, N9519);
xor XOR2 (N10396, N10390, N2974);
buf BUF1 (N10397, N10377);
nand NAND3 (N10398, N10395, N5127, N7845);
xor XOR2 (N10399, N10394, N10360);
or OR3 (N10400, N10397, N1317, N1243);
nand NAND3 (N10401, N10366, N5047, N8697);
not NOT1 (N10402, N10401);
not NOT1 (N10403, N10392);
not NOT1 (N10404, N10403);
not NOT1 (N10405, N10389);
or OR2 (N10406, N10384, N8657);
not NOT1 (N10407, N10399);
and AND4 (N10408, N10406, N8868, N3980, N8894);
and AND4 (N10409, N10404, N9641, N8412, N6624);
not NOT1 (N10410, N10407);
nor NOR2 (N10411, N10410, N324);
nand NAND4 (N10412, N10383, N7544, N1049, N4881);
not NOT1 (N10413, N10411);
buf BUF1 (N10414, N10396);
nand NAND3 (N10415, N10402, N430, N6773);
buf BUF1 (N10416, N10414);
not NOT1 (N10417, N10393);
and AND2 (N10418, N10416, N3632);
xor XOR2 (N10419, N10412, N10345);
xor XOR2 (N10420, N10419, N3128);
and AND2 (N10421, N10400, N9305);
buf BUF1 (N10422, N10421);
and AND2 (N10423, N10420, N4612);
and AND3 (N10424, N10398, N1428, N7110);
buf BUF1 (N10425, N10405);
or OR4 (N10426, N10415, N6865, N5971, N6882);
buf BUF1 (N10427, N10424);
and AND3 (N10428, N10413, N5810, N638);
nor NOR2 (N10429, N10408, N3559);
nor NOR3 (N10430, N10427, N4338, N1006);
buf BUF1 (N10431, N10429);
and AND2 (N10432, N10422, N6630);
nor NOR2 (N10433, N10426, N8179);
or OR2 (N10434, N10431, N4348);
not NOT1 (N10435, N10418);
nand NAND3 (N10436, N10425, N6448, N7601);
and AND2 (N10437, N10436, N1346);
xor XOR2 (N10438, N10432, N5329);
and AND2 (N10439, N10434, N6267);
not NOT1 (N10440, N10437);
and AND4 (N10441, N10440, N10242, N1087, N4528);
and AND2 (N10442, N10409, N4297);
nand NAND4 (N10443, N10441, N376, N3384, N8597);
or OR4 (N10444, N10442, N7738, N5629, N7757);
not NOT1 (N10445, N10438);
nor NOR2 (N10446, N10435, N9166);
xor XOR2 (N10447, N10417, N9336);
xor XOR2 (N10448, N10443, N7720);
buf BUF1 (N10449, N10445);
nor NOR3 (N10450, N10448, N8420, N2952);
and AND3 (N10451, N10439, N8326, N4954);
nor NOR4 (N10452, N10450, N7645, N9996, N9942);
xor XOR2 (N10453, N10451, N2872);
not NOT1 (N10454, N10433);
xor XOR2 (N10455, N10453, N3071);
buf BUF1 (N10456, N10447);
nor NOR4 (N10457, N10455, N9843, N1292, N855);
xor XOR2 (N10458, N10430, N10081);
nand NAND4 (N10459, N10444, N3848, N7117, N10140);
xor XOR2 (N10460, N10458, N5055);
buf BUF1 (N10461, N10457);
or OR3 (N10462, N10456, N9613, N1631);
nand NAND3 (N10463, N10461, N7558, N7180);
xor XOR2 (N10464, N10460, N1877);
nor NOR4 (N10465, N10459, N2576, N844, N3515);
buf BUF1 (N10466, N10452);
not NOT1 (N10467, N10462);
buf BUF1 (N10468, N10466);
nand NAND2 (N10469, N10465, N5913);
nor NOR3 (N10470, N10467, N3959, N9116);
or OR3 (N10471, N10469, N10100, N9283);
buf BUF1 (N10472, N10428);
buf BUF1 (N10473, N10471);
buf BUF1 (N10474, N10472);
nand NAND3 (N10475, N10473, N1491, N5892);
nand NAND2 (N10476, N10463, N273);
or OR3 (N10477, N10454, N1521, N9247);
nor NOR2 (N10478, N10423, N3404);
buf BUF1 (N10479, N10474);
xor XOR2 (N10480, N10449, N7363);
nor NOR4 (N10481, N10470, N4726, N1871, N2145);
buf BUF1 (N10482, N10475);
xor XOR2 (N10483, N10480, N3564);
and AND3 (N10484, N10468, N8234, N8362);
nor NOR4 (N10485, N10484, N1685, N918, N8506);
and AND2 (N10486, N10478, N8245);
buf BUF1 (N10487, N10482);
buf BUF1 (N10488, N10479);
and AND3 (N10489, N10483, N9152, N83);
or OR3 (N10490, N10477, N9702, N6760);
or OR2 (N10491, N10488, N64);
buf BUF1 (N10492, N10481);
and AND2 (N10493, N10492, N10371);
nor NOR4 (N10494, N10491, N5425, N4350, N8331);
nand NAND2 (N10495, N10446, N1405);
or OR2 (N10496, N10493, N9587);
not NOT1 (N10497, N10464);
or OR4 (N10498, N10495, N2742, N3817, N569);
nand NAND2 (N10499, N10494, N1812);
nand NAND4 (N10500, N10476, N9814, N6018, N764);
and AND4 (N10501, N10485, N5670, N7301, N3240);
nand NAND3 (N10502, N10489, N7918, N3739);
nor NOR4 (N10503, N10487, N9193, N8735, N9020);
nor NOR3 (N10504, N10498, N5115, N5862);
or OR2 (N10505, N10499, N9634);
not NOT1 (N10506, N10496);
xor XOR2 (N10507, N10506, N4704);
xor XOR2 (N10508, N10486, N8498);
xor XOR2 (N10509, N10504, N664);
and AND2 (N10510, N10508, N9273);
nor NOR4 (N10511, N10502, N6834, N62, N9562);
nand NAND2 (N10512, N10507, N5481);
xor XOR2 (N10513, N10511, N7504);
xor XOR2 (N10514, N10509, N5193);
xor XOR2 (N10515, N10503, N812);
nand NAND3 (N10516, N10497, N3162, N8858);
buf BUF1 (N10517, N10516);
buf BUF1 (N10518, N10514);
not NOT1 (N10519, N10513);
nand NAND3 (N10520, N10519, N7013, N4503);
nand NAND3 (N10521, N10518, N697, N5087);
buf BUF1 (N10522, N10501);
not NOT1 (N10523, N10505);
buf BUF1 (N10524, N10510);
nor NOR3 (N10525, N10523, N9696, N4968);
and AND2 (N10526, N10521, N5869);
nor NOR3 (N10527, N10520, N188, N9416);
nor NOR3 (N10528, N10490, N8504, N5058);
not NOT1 (N10529, N10525);
not NOT1 (N10530, N10517);
not NOT1 (N10531, N10528);
or OR2 (N10532, N10531, N9747);
or OR4 (N10533, N10530, N5548, N2706, N9047);
not NOT1 (N10534, N10526);
buf BUF1 (N10535, N10500);
or OR4 (N10536, N10524, N8321, N3476, N6533);
not NOT1 (N10537, N10536);
not NOT1 (N10538, N10535);
nor NOR3 (N10539, N10522, N1315, N9420);
buf BUF1 (N10540, N10515);
or OR2 (N10541, N10533, N9021);
xor XOR2 (N10542, N10538, N6860);
and AND2 (N10543, N10527, N9523);
not NOT1 (N10544, N10529);
xor XOR2 (N10545, N10541, N10206);
xor XOR2 (N10546, N10540, N9071);
nand NAND4 (N10547, N10542, N4722, N6412, N925);
or OR2 (N10548, N10532, N260);
not NOT1 (N10549, N10512);
nand NAND2 (N10550, N10545, N3834);
xor XOR2 (N10551, N10549, N5637);
nand NAND4 (N10552, N10550, N3959, N3175, N7623);
xor XOR2 (N10553, N10552, N6941);
and AND3 (N10554, N10548, N1906, N6179);
nand NAND4 (N10555, N10551, N2187, N4516, N10220);
and AND2 (N10556, N10554, N1075);
buf BUF1 (N10557, N10546);
buf BUF1 (N10558, N10553);
nor NOR3 (N10559, N10547, N8527, N2711);
buf BUF1 (N10560, N10534);
nand NAND3 (N10561, N10560, N5478, N8606);
or OR2 (N10562, N10556, N1423);
buf BUF1 (N10563, N10544);
nor NOR4 (N10564, N10537, N9095, N4365, N3046);
not NOT1 (N10565, N10563);
or OR2 (N10566, N10559, N1318);
not NOT1 (N10567, N10562);
or OR3 (N10568, N10566, N3920, N4598);
or OR4 (N10569, N10555, N2691, N3120, N1867);
nor NOR3 (N10570, N10558, N2917, N3393);
buf BUF1 (N10571, N10570);
nor NOR3 (N10572, N10565, N1878, N2390);
or OR4 (N10573, N10561, N3712, N8913, N1820);
buf BUF1 (N10574, N10564);
nor NOR4 (N10575, N10573, N6355, N7372, N4702);
or OR2 (N10576, N10572, N7131);
not NOT1 (N10577, N10557);
xor XOR2 (N10578, N10539, N7301);
nor NOR2 (N10579, N10543, N8626);
and AND3 (N10580, N10571, N5152, N9747);
xor XOR2 (N10581, N10578, N7482);
and AND4 (N10582, N10580, N4558, N5390, N4861);
not NOT1 (N10583, N10579);
xor XOR2 (N10584, N10582, N5499);
or OR3 (N10585, N10584, N10018, N8724);
not NOT1 (N10586, N10567);
and AND2 (N10587, N10569, N7272);
and AND2 (N10588, N10568, N6759);
or OR2 (N10589, N10575, N2721);
and AND2 (N10590, N10585, N655);
or OR2 (N10591, N10589, N5379);
xor XOR2 (N10592, N10590, N3889);
or OR4 (N10593, N10583, N9056, N3589, N3506);
not NOT1 (N10594, N10592);
not NOT1 (N10595, N10581);
buf BUF1 (N10596, N10586);
or OR4 (N10597, N10595, N8566, N5278, N1526);
xor XOR2 (N10598, N10591, N6590);
xor XOR2 (N10599, N10576, N2958);
and AND4 (N10600, N10594, N1623, N2463, N7790);
and AND4 (N10601, N10593, N2658, N4283, N6846);
nor NOR3 (N10602, N10601, N422, N5399);
nor NOR2 (N10603, N10600, N2432);
not NOT1 (N10604, N10587);
and AND4 (N10605, N10574, N5382, N444, N7236);
nor NOR2 (N10606, N10598, N3872);
xor XOR2 (N10607, N10605, N4400);
nand NAND4 (N10608, N10602, N6420, N2522, N10067);
and AND2 (N10609, N10604, N1445);
nand NAND4 (N10610, N10577, N8840, N54, N1441);
not NOT1 (N10611, N10610);
nor NOR3 (N10612, N10603, N598, N2527);
buf BUF1 (N10613, N10608);
not NOT1 (N10614, N10597);
nor NOR2 (N10615, N10611, N2578);
xor XOR2 (N10616, N10612, N6150);
nand NAND2 (N10617, N10616, N1531);
nand NAND3 (N10618, N10614, N1667, N8429);
buf BUF1 (N10619, N10609);
xor XOR2 (N10620, N10607, N7380);
nand NAND4 (N10621, N10618, N5517, N3301, N4811);
and AND3 (N10622, N10599, N8409, N1400);
xor XOR2 (N10623, N10613, N4903);
nand NAND2 (N10624, N10588, N1114);
buf BUF1 (N10625, N10624);
xor XOR2 (N10626, N10619, N9070);
or OR4 (N10627, N10625, N1266, N733, N6595);
nor NOR2 (N10628, N10623, N7780);
nand NAND2 (N10629, N10596, N2987);
xor XOR2 (N10630, N10606, N8655);
nand NAND3 (N10631, N10626, N4002, N6056);
or OR2 (N10632, N10630, N9964);
buf BUF1 (N10633, N10621);
xor XOR2 (N10634, N10633, N6411);
xor XOR2 (N10635, N10629, N4073);
or OR3 (N10636, N10615, N8870, N2469);
not NOT1 (N10637, N10620);
and AND4 (N10638, N10617, N7614, N10050, N4904);
nand NAND4 (N10639, N10632, N126, N6024, N1859);
nor NOR3 (N10640, N10639, N2188, N2687);
nand NAND3 (N10641, N10622, N2429, N5368);
buf BUF1 (N10642, N10627);
or OR2 (N10643, N10642, N1740);
and AND2 (N10644, N10640, N6078);
and AND3 (N10645, N10641, N10635, N839);
buf BUF1 (N10646, N6593);
buf BUF1 (N10647, N10628);
not NOT1 (N10648, N10643);
xor XOR2 (N10649, N10631, N2228);
xor XOR2 (N10650, N10644, N4730);
nor NOR3 (N10651, N10650, N7385, N8525);
xor XOR2 (N10652, N10651, N3337);
nor NOR4 (N10653, N10638, N2450, N10240, N3125);
nor NOR3 (N10654, N10648, N5817, N206);
or OR3 (N10655, N10653, N2297, N8592);
nor NOR2 (N10656, N10652, N3926);
nand NAND2 (N10657, N10645, N8783);
not NOT1 (N10658, N10657);
not NOT1 (N10659, N10634);
nand NAND4 (N10660, N10647, N9805, N5306, N8078);
and AND4 (N10661, N10658, N5820, N2642, N7760);
nand NAND4 (N10662, N10636, N4836, N5084, N7193);
nor NOR2 (N10663, N10637, N7667);
or OR4 (N10664, N10656, N3850, N10116, N7771);
and AND4 (N10665, N10663, N1374, N322, N849);
and AND4 (N10666, N10649, N7879, N6694, N10164);
xor XOR2 (N10667, N10655, N2244);
or OR2 (N10668, N10664, N2494);
and AND2 (N10669, N10662, N3529);
not NOT1 (N10670, N10646);
or OR2 (N10671, N10668, N8784);
not NOT1 (N10672, N10669);
or OR2 (N10673, N10660, N7728);
buf BUF1 (N10674, N10667);
and AND2 (N10675, N10673, N8467);
buf BUF1 (N10676, N10666);
buf BUF1 (N10677, N10675);
buf BUF1 (N10678, N10671);
and AND3 (N10679, N10672, N2248, N9565);
nor NOR2 (N10680, N10654, N10412);
or OR4 (N10681, N10676, N5387, N8033, N2687);
nor NOR2 (N10682, N10661, N2031);
nor NOR2 (N10683, N10678, N2614);
not NOT1 (N10684, N10683);
nand NAND3 (N10685, N10680, N7531, N7538);
or OR2 (N10686, N10682, N9789);
buf BUF1 (N10687, N10659);
and AND3 (N10688, N10685, N3957, N5040);
nor NOR2 (N10689, N10677, N1682);
xor XOR2 (N10690, N10687, N1707);
buf BUF1 (N10691, N10679);
xor XOR2 (N10692, N10670, N2363);
nor NOR4 (N10693, N10692, N3454, N2117, N5329);
buf BUF1 (N10694, N10674);
or OR4 (N10695, N10686, N1560, N2628, N10564);
xor XOR2 (N10696, N10690, N9043);
nand NAND3 (N10697, N10693, N5824, N2284);
nand NAND3 (N10698, N10681, N8934, N5000);
nand NAND2 (N10699, N10688, N6519);
buf BUF1 (N10700, N10691);
and AND3 (N10701, N10695, N6577, N1000);
nor NOR3 (N10702, N10698, N7583, N842);
buf BUF1 (N10703, N10697);
not NOT1 (N10704, N10696);
not NOT1 (N10705, N10694);
buf BUF1 (N10706, N10702);
and AND3 (N10707, N10706, N3306, N7878);
or OR3 (N10708, N10684, N2718, N6949);
and AND2 (N10709, N10705, N2227);
nand NAND4 (N10710, N10707, N123, N7004, N5072);
or OR2 (N10711, N10710, N6365);
or OR3 (N10712, N10700, N6694, N9778);
nand NAND4 (N10713, N10699, N1995, N6992, N5041);
and AND4 (N10714, N10712, N1660, N3096, N9479);
nor NOR3 (N10715, N10701, N10683, N6251);
xor XOR2 (N10716, N10709, N3020);
not NOT1 (N10717, N10714);
nand NAND2 (N10718, N10704, N5690);
and AND3 (N10719, N10718, N9365, N9238);
buf BUF1 (N10720, N10715);
and AND2 (N10721, N10719, N3124);
not NOT1 (N10722, N10711);
nor NOR2 (N10723, N10713, N6741);
nand NAND4 (N10724, N10721, N5676, N929, N5266);
nand NAND3 (N10725, N10723, N3258, N9691);
and AND4 (N10726, N10722, N6698, N6503, N6031);
not NOT1 (N10727, N10724);
and AND2 (N10728, N10727, N6646);
not NOT1 (N10729, N10720);
or OR3 (N10730, N10729, N6471, N9656);
or OR3 (N10731, N10730, N10717, N2817);
buf BUF1 (N10732, N2732);
and AND3 (N10733, N10703, N2183, N9223);
xor XOR2 (N10734, N10731, N7277);
nand NAND3 (N10735, N10728, N1241, N234);
nand NAND4 (N10736, N10733, N5708, N3682, N8616);
nand NAND2 (N10737, N10716, N655);
nand NAND4 (N10738, N10725, N7188, N4918, N9613);
and AND2 (N10739, N10665, N95);
or OR2 (N10740, N10732, N162);
and AND2 (N10741, N10737, N2395);
nor NOR3 (N10742, N10736, N8124, N6620);
xor XOR2 (N10743, N10738, N6718);
nand NAND2 (N10744, N10739, N7216);
or OR3 (N10745, N10689, N9982, N10006);
not NOT1 (N10746, N10745);
nor NOR2 (N10747, N10740, N3263);
xor XOR2 (N10748, N10747, N1631);
and AND4 (N10749, N10744, N2676, N9023, N4685);
or OR2 (N10750, N10749, N6211);
nor NOR2 (N10751, N10735, N10618);
and AND3 (N10752, N10734, N4312, N6186);
not NOT1 (N10753, N10743);
not NOT1 (N10754, N10742);
and AND4 (N10755, N10753, N4513, N7583, N4286);
nand NAND3 (N10756, N10750, N8437, N1784);
buf BUF1 (N10757, N10752);
nor NOR4 (N10758, N10755, N607, N6984, N3153);
xor XOR2 (N10759, N10751, N7628);
nor NOR4 (N10760, N10759, N8810, N10034, N5072);
not NOT1 (N10761, N10754);
buf BUF1 (N10762, N10726);
buf BUF1 (N10763, N10741);
or OR4 (N10764, N10762, N6001, N55, N6089);
buf BUF1 (N10765, N10746);
buf BUF1 (N10766, N10758);
xor XOR2 (N10767, N10764, N7967);
buf BUF1 (N10768, N10760);
xor XOR2 (N10769, N10763, N3081);
not NOT1 (N10770, N10765);
buf BUF1 (N10771, N10748);
and AND4 (N10772, N10766, N10331, N18, N1534);
buf BUF1 (N10773, N10769);
not NOT1 (N10774, N10757);
xor XOR2 (N10775, N10772, N5208);
buf BUF1 (N10776, N10771);
and AND4 (N10777, N10768, N10397, N6836, N7661);
nor NOR2 (N10778, N10776, N9709);
nand NAND3 (N10779, N10756, N9026, N3124);
and AND4 (N10780, N10774, N1184, N3456, N2920);
not NOT1 (N10781, N10761);
and AND4 (N10782, N10770, N3760, N10332, N52);
xor XOR2 (N10783, N10777, N3498);
xor XOR2 (N10784, N10775, N8153);
and AND4 (N10785, N10782, N7319, N3184, N4498);
buf BUF1 (N10786, N10779);
nand NAND4 (N10787, N10783, N3889, N5601, N8773);
xor XOR2 (N10788, N10780, N8911);
and AND4 (N10789, N10788, N9104, N3326, N6475);
and AND2 (N10790, N10767, N7794);
or OR4 (N10791, N10789, N7025, N1068, N1715);
and AND4 (N10792, N10784, N10713, N2394, N2937);
xor XOR2 (N10793, N10781, N7788);
xor XOR2 (N10794, N10792, N6385);
and AND3 (N10795, N10785, N6220, N4336);
buf BUF1 (N10796, N10791);
or OR2 (N10797, N10793, N427);
and AND4 (N10798, N10794, N3639, N10700, N2820);
or OR4 (N10799, N10797, N8, N5350, N2604);
or OR4 (N10800, N10799, N3387, N3917, N8457);
nand NAND3 (N10801, N10708, N1218, N2330);
not NOT1 (N10802, N10796);
xor XOR2 (N10803, N10795, N1714);
nand NAND3 (N10804, N10787, N3777, N9017);
buf BUF1 (N10805, N10798);
nor NOR4 (N10806, N10790, N8587, N7160, N8304);
xor XOR2 (N10807, N10804, N8304);
xor XOR2 (N10808, N10786, N5041);
not NOT1 (N10809, N10802);
nor NOR4 (N10810, N10806, N3147, N1577, N4804);
xor XOR2 (N10811, N10803, N1757);
not NOT1 (N10812, N10810);
nor NOR4 (N10813, N10808, N3070, N3230, N8093);
nand NAND3 (N10814, N10807, N9937, N8170);
xor XOR2 (N10815, N10809, N1334);
nor NOR2 (N10816, N10811, N7324);
not NOT1 (N10817, N10773);
not NOT1 (N10818, N10815);
not NOT1 (N10819, N10818);
buf BUF1 (N10820, N10816);
not NOT1 (N10821, N10817);
and AND4 (N10822, N10821, N10053, N2968, N4633);
nand NAND3 (N10823, N10819, N8300, N8917);
nand NAND2 (N10824, N10800, N3026);
buf BUF1 (N10825, N10812);
nor NOR2 (N10826, N10825, N168);
not NOT1 (N10827, N10826);
and AND3 (N10828, N10822, N979, N3460);
buf BUF1 (N10829, N10814);
buf BUF1 (N10830, N10778);
and AND2 (N10831, N10824, N6975);
nand NAND4 (N10832, N10827, N3658, N980, N6880);
nand NAND2 (N10833, N10832, N6235);
buf BUF1 (N10834, N10823);
buf BUF1 (N10835, N10831);
not NOT1 (N10836, N10829);
not NOT1 (N10837, N10801);
and AND2 (N10838, N10835, N8128);
or OR2 (N10839, N10838, N706);
or OR4 (N10840, N10805, N4879, N2207, N4405);
and AND2 (N10841, N10840, N254);
buf BUF1 (N10842, N10839);
nor NOR2 (N10843, N10833, N2607);
nand NAND2 (N10844, N10830, N6814);
buf BUF1 (N10845, N10841);
and AND3 (N10846, N10842, N8095, N5339);
and AND4 (N10847, N10837, N3074, N10660, N7631);
or OR3 (N10848, N10828, N2802, N4365);
and AND3 (N10849, N10846, N9474, N728);
nand NAND3 (N10850, N10820, N4110, N4984);
nand NAND2 (N10851, N10850, N1642);
nand NAND4 (N10852, N10834, N5150, N4339, N10172);
buf BUF1 (N10853, N10847);
and AND2 (N10854, N10853, N6026);
and AND3 (N10855, N10854, N3940, N9649);
or OR3 (N10856, N10851, N3311, N5059);
xor XOR2 (N10857, N10855, N339);
nor NOR2 (N10858, N10857, N7559);
or OR4 (N10859, N10856, N9365, N8503, N4768);
xor XOR2 (N10860, N10844, N8486);
and AND3 (N10861, N10858, N6824, N15);
buf BUF1 (N10862, N10849);
and AND4 (N10863, N10859, N8723, N6606, N7211);
or OR3 (N10864, N10860, N8090, N4108);
nand NAND3 (N10865, N10863, N855, N1307);
xor XOR2 (N10866, N10864, N1522);
and AND4 (N10867, N10866, N9370, N3397, N2502);
xor XOR2 (N10868, N10848, N8501);
buf BUF1 (N10869, N10868);
and AND4 (N10870, N10813, N4862, N9887, N10771);
buf BUF1 (N10871, N10869);
nand NAND4 (N10872, N10852, N7741, N3621, N5849);
or OR4 (N10873, N10867, N8290, N8657, N1953);
or OR3 (N10874, N10836, N8938, N9822);
nand NAND2 (N10875, N10862, N6632);
not NOT1 (N10876, N10873);
xor XOR2 (N10877, N10845, N9145);
xor XOR2 (N10878, N10843, N6778);
nor NOR2 (N10879, N10874, N4881);
buf BUF1 (N10880, N10861);
nand NAND4 (N10881, N10878, N4215, N6561, N9633);
buf BUF1 (N10882, N10865);
and AND2 (N10883, N10872, N2115);
nand NAND4 (N10884, N10871, N3399, N2101, N4191);
xor XOR2 (N10885, N10877, N2931);
nor NOR4 (N10886, N10876, N7115, N4538, N3735);
nor NOR4 (N10887, N10882, N10298, N97, N9003);
buf BUF1 (N10888, N10875);
xor XOR2 (N10889, N10885, N2998);
nor NOR4 (N10890, N10888, N10012, N2315, N4590);
or OR2 (N10891, N10886, N3470);
buf BUF1 (N10892, N10880);
or OR4 (N10893, N10881, N9738, N9966, N5546);
buf BUF1 (N10894, N10883);
or OR2 (N10895, N10870, N10524);
buf BUF1 (N10896, N10884);
buf BUF1 (N10897, N10887);
xor XOR2 (N10898, N10879, N7125);
nor NOR3 (N10899, N10891, N10743, N7650);
xor XOR2 (N10900, N10896, N9719);
and AND3 (N10901, N10894, N2118, N4583);
nand NAND3 (N10902, N10897, N467, N6133);
nand NAND4 (N10903, N10892, N5301, N6599, N2814);
and AND2 (N10904, N10893, N7707);
nand NAND2 (N10905, N10890, N5841);
buf BUF1 (N10906, N10903);
nand NAND2 (N10907, N10904, N9085);
or OR4 (N10908, N10901, N9658, N4266, N7636);
not NOT1 (N10909, N10906);
not NOT1 (N10910, N10905);
or OR3 (N10911, N10889, N3137, N3686);
nand NAND2 (N10912, N10898, N3107);
and AND2 (N10913, N10899, N8489);
nor NOR4 (N10914, N10909, N10221, N9156, N7572);
xor XOR2 (N10915, N10895, N10193);
buf BUF1 (N10916, N10913);
xor XOR2 (N10917, N10915, N4636);
not NOT1 (N10918, N10916);
and AND4 (N10919, N10908, N1246, N2235, N4237);
xor XOR2 (N10920, N10919, N9656);
or OR3 (N10921, N10914, N2360, N1534);
xor XOR2 (N10922, N10900, N7108);
and AND2 (N10923, N10917, N5745);
and AND3 (N10924, N10922, N10090, N10260);
nor NOR3 (N10925, N10918, N5126, N1833);
and AND4 (N10926, N10911, N8130, N1288, N7571);
and AND3 (N10927, N10907, N10440, N6486);
not NOT1 (N10928, N10920);
buf BUF1 (N10929, N10925);
buf BUF1 (N10930, N10929);
and AND2 (N10931, N10927, N5811);
nand NAND4 (N10932, N10924, N7951, N9628, N5957);
not NOT1 (N10933, N10932);
xor XOR2 (N10934, N10902, N7862);
nor NOR2 (N10935, N10923, N5130);
nor NOR2 (N10936, N10930, N7236);
or OR2 (N10937, N10928, N9144);
and AND3 (N10938, N10910, N243, N9698);
buf BUF1 (N10939, N10912);
and AND4 (N10940, N10931, N3346, N2986, N6063);
buf BUF1 (N10941, N10940);
nor NOR2 (N10942, N10939, N3876);
nand NAND3 (N10943, N10921, N477, N928);
nand NAND3 (N10944, N10935, N2303, N5222);
xor XOR2 (N10945, N10944, N1316);
nor NOR3 (N10946, N10938, N9294, N5283);
and AND3 (N10947, N10943, N4821, N10451);
xor XOR2 (N10948, N10933, N8787);
and AND3 (N10949, N10926, N10916, N8070);
buf BUF1 (N10950, N10936);
nand NAND3 (N10951, N10941, N6847, N7237);
nor NOR3 (N10952, N10942, N686, N8986);
buf BUF1 (N10953, N10947);
and AND2 (N10954, N10934, N6549);
not NOT1 (N10955, N10954);
nor NOR3 (N10956, N10950, N2447, N5364);
nor NOR3 (N10957, N10948, N9715, N10269);
not NOT1 (N10958, N10953);
and AND3 (N10959, N10956, N3861, N9486);
buf BUF1 (N10960, N10949);
nor NOR3 (N10961, N10952, N5016, N8604);
or OR3 (N10962, N10951, N8600, N1516);
nor NOR2 (N10963, N10962, N294);
buf BUF1 (N10964, N10946);
not NOT1 (N10965, N10963);
or OR2 (N10966, N10960, N10931);
nor NOR4 (N10967, N10945, N4528, N10428, N6177);
nor NOR4 (N10968, N10959, N7768, N2629, N1894);
nand NAND4 (N10969, N10957, N4309, N5545, N319);
xor XOR2 (N10970, N10955, N8308);
buf BUF1 (N10971, N10968);
and AND2 (N10972, N10966, N5156);
nor NOR3 (N10973, N10969, N6456, N8512);
and AND2 (N10974, N10961, N7658);
not NOT1 (N10975, N10972);
and AND4 (N10976, N10967, N1321, N5715, N8149);
nor NOR2 (N10977, N10958, N3333);
nor NOR3 (N10978, N10973, N3305, N3572);
and AND3 (N10979, N10970, N5534, N7580);
buf BUF1 (N10980, N10965);
and AND4 (N10981, N10977, N4014, N9078, N5473);
nor NOR3 (N10982, N10937, N7721, N9133);
and AND2 (N10983, N10981, N10845);
nor NOR4 (N10984, N10975, N9390, N7836, N9875);
nand NAND2 (N10985, N10984, N4560);
buf BUF1 (N10986, N10985);
and AND3 (N10987, N10964, N5109, N1737);
buf BUF1 (N10988, N10971);
buf BUF1 (N10989, N10979);
nand NAND4 (N10990, N10988, N8506, N4881, N4835);
buf BUF1 (N10991, N10976);
buf BUF1 (N10992, N10982);
buf BUF1 (N10993, N10987);
nand NAND2 (N10994, N10978, N2035);
or OR4 (N10995, N10992, N10226, N3195, N4606);
xor XOR2 (N10996, N10991, N8857);
not NOT1 (N10997, N10996);
xor XOR2 (N10998, N10990, N3918);
nand NAND4 (N10999, N10989, N4517, N583, N4939);
nand NAND3 (N11000, N10994, N6253, N1506);
buf BUF1 (N11001, N10997);
not NOT1 (N11002, N10983);
xor XOR2 (N11003, N11002, N2143);
nor NOR2 (N11004, N10980, N1739);
or OR4 (N11005, N10998, N2400, N9334, N1466);
nor NOR4 (N11006, N10999, N5821, N9699, N7588);
nor NOR3 (N11007, N11005, N1770, N2395);
xor XOR2 (N11008, N11001, N4649);
xor XOR2 (N11009, N11007, N10324);
not NOT1 (N11010, N11006);
or OR3 (N11011, N11000, N4908, N5631);
nor NOR3 (N11012, N10995, N10443, N6167);
nand NAND2 (N11013, N11010, N9291);
and AND4 (N11014, N11004, N5776, N2069, N10558);
and AND2 (N11015, N11011, N7617);
nand NAND4 (N11016, N11015, N7251, N4836, N2588);
or OR4 (N11017, N10986, N2522, N7070, N10843);
buf BUF1 (N11018, N10993);
buf BUF1 (N11019, N11003);
or OR3 (N11020, N11012, N4612, N2207);
and AND3 (N11021, N11019, N265, N8836);
or OR4 (N11022, N11017, N1839, N5478, N9543);
and AND3 (N11023, N11008, N685, N5884);
not NOT1 (N11024, N11018);
not NOT1 (N11025, N11024);
buf BUF1 (N11026, N11014);
and AND3 (N11027, N11023, N5633, N3155);
buf BUF1 (N11028, N10974);
buf BUF1 (N11029, N11025);
not NOT1 (N11030, N11021);
xor XOR2 (N11031, N11022, N8954);
xor XOR2 (N11032, N11027, N8762);
buf BUF1 (N11033, N11009);
buf BUF1 (N11034, N11028);
or OR4 (N11035, N11030, N1328, N9156, N9031);
xor XOR2 (N11036, N11029, N8807);
nor NOR2 (N11037, N11036, N2612);
not NOT1 (N11038, N11033);
buf BUF1 (N11039, N11035);
nor NOR3 (N11040, N11039, N3187, N5882);
not NOT1 (N11041, N11020);
xor XOR2 (N11042, N11041, N4782);
and AND2 (N11043, N11032, N6773);
nor NOR3 (N11044, N11038, N4044, N8662);
not NOT1 (N11045, N11026);
nor NOR2 (N11046, N11043, N10542);
nor NOR4 (N11047, N11042, N4393, N10562, N8709);
or OR3 (N11048, N11047, N7645, N7216);
or OR3 (N11049, N11045, N5828, N1123);
or OR4 (N11050, N11013, N1499, N4563, N9759);
buf BUF1 (N11051, N11046);
nor NOR4 (N11052, N11040, N2269, N2607, N10608);
nor NOR4 (N11053, N11044, N4120, N10220, N4885);
or OR2 (N11054, N11050, N3031);
buf BUF1 (N11055, N11053);
and AND3 (N11056, N11055, N9712, N3026);
not NOT1 (N11057, N11034);
buf BUF1 (N11058, N11037);
or OR2 (N11059, N11056, N4366);
nor NOR2 (N11060, N11052, N2700);
and AND2 (N11061, N11048, N3403);
and AND2 (N11062, N11060, N3323);
nor NOR2 (N11063, N11058, N7240);
and AND2 (N11064, N11049, N2121);
nand NAND4 (N11065, N11064, N6368, N701, N6142);
xor XOR2 (N11066, N11065, N6361);
xor XOR2 (N11067, N11061, N2886);
nand NAND2 (N11068, N11062, N2976);
and AND4 (N11069, N11051, N5451, N6741, N703);
nor NOR4 (N11070, N11069, N6431, N163, N181);
or OR3 (N11071, N11016, N8954, N9634);
buf BUF1 (N11072, N11067);
nand NAND2 (N11073, N11054, N2503);
buf BUF1 (N11074, N11073);
buf BUF1 (N11075, N11074);
buf BUF1 (N11076, N11071);
buf BUF1 (N11077, N11059);
nand NAND2 (N11078, N11068, N8752);
not NOT1 (N11079, N11063);
nand NAND4 (N11080, N11072, N8307, N228, N9018);
nand NAND4 (N11081, N11075, N2877, N400, N3849);
nand NAND2 (N11082, N11070, N10882);
not NOT1 (N11083, N11078);
buf BUF1 (N11084, N11077);
buf BUF1 (N11085, N11031);
nor NOR2 (N11086, N11084, N9505);
or OR2 (N11087, N11082, N6299);
buf BUF1 (N11088, N11085);
or OR2 (N11089, N11083, N5891);
not NOT1 (N11090, N11081);
not NOT1 (N11091, N11089);
not NOT1 (N11092, N11086);
buf BUF1 (N11093, N11080);
xor XOR2 (N11094, N11066, N3806);
not NOT1 (N11095, N11092);
nor NOR3 (N11096, N11091, N7620, N10847);
nand NAND2 (N11097, N11093, N1617);
xor XOR2 (N11098, N11090, N834);
not NOT1 (N11099, N11079);
not NOT1 (N11100, N11098);
nand NAND2 (N11101, N11096, N4142);
not NOT1 (N11102, N11095);
nor NOR3 (N11103, N11100, N10887, N1502);
and AND4 (N11104, N11087, N7768, N10585, N5268);
and AND2 (N11105, N11094, N4710);
xor XOR2 (N11106, N11057, N7746);
and AND3 (N11107, N11105, N8172, N5833);
nand NAND4 (N11108, N11107, N2075, N671, N4632);
xor XOR2 (N11109, N11099, N8505);
buf BUF1 (N11110, N11088);
buf BUF1 (N11111, N11102);
not NOT1 (N11112, N11097);
nand NAND3 (N11113, N11104, N5832, N6352);
nor NOR2 (N11114, N11106, N8917);
nand NAND4 (N11115, N11103, N6528, N1131, N6041);
and AND4 (N11116, N11101, N5922, N4802, N7557);
or OR3 (N11117, N11110, N9863, N11106);
nor NOR2 (N11118, N11116, N4962);
nor NOR2 (N11119, N11076, N2518);
xor XOR2 (N11120, N11117, N6400);
xor XOR2 (N11121, N11120, N4437);
or OR2 (N11122, N11109, N1748);
not NOT1 (N11123, N11115);
buf BUF1 (N11124, N11121);
nor NOR2 (N11125, N11114, N5124);
nand NAND4 (N11126, N11118, N7229, N2142, N6978);
nand NAND2 (N11127, N11111, N5248);
and AND3 (N11128, N11125, N3322, N8144);
nand NAND4 (N11129, N11119, N2577, N3250, N6774);
nand NAND4 (N11130, N11108, N3884, N9002, N6084);
not NOT1 (N11131, N11113);
or OR3 (N11132, N11127, N4260, N9495);
xor XOR2 (N11133, N11122, N4185);
nand NAND4 (N11134, N11126, N7407, N6979, N1461);
xor XOR2 (N11135, N11112, N4330);
xor XOR2 (N11136, N11128, N10575);
nand NAND4 (N11137, N11130, N3121, N7045, N7650);
and AND3 (N11138, N11137, N2225, N9062);
nor NOR3 (N11139, N11129, N3062, N2307);
xor XOR2 (N11140, N11138, N11094);
xor XOR2 (N11141, N11140, N9315);
nand NAND4 (N11142, N11124, N1869, N8025, N2274);
not NOT1 (N11143, N11135);
and AND4 (N11144, N11142, N5785, N2305, N9220);
buf BUF1 (N11145, N11136);
nor NOR2 (N11146, N11143, N5563);
nor NOR3 (N11147, N11145, N5632, N3236);
and AND2 (N11148, N11131, N9688);
nand NAND4 (N11149, N11147, N1473, N2663, N2636);
not NOT1 (N11150, N11132);
and AND3 (N11151, N11148, N1314, N1426);
not NOT1 (N11152, N11150);
or OR3 (N11153, N11139, N9749, N4743);
nor NOR3 (N11154, N11134, N2508, N1198);
not NOT1 (N11155, N11151);
and AND4 (N11156, N11141, N7009, N3348, N1327);
not NOT1 (N11157, N11152);
nor NOR3 (N11158, N11153, N3575, N9742);
or OR2 (N11159, N11154, N8027);
nor NOR3 (N11160, N11144, N151, N4556);
nand NAND3 (N11161, N11156, N3728, N8632);
nand NAND2 (N11162, N11133, N2292);
and AND3 (N11163, N11158, N6538, N9569);
and AND4 (N11164, N11146, N9337, N4028, N6665);
or OR2 (N11165, N11164, N5174);
xor XOR2 (N11166, N11149, N7664);
nand NAND3 (N11167, N11165, N438, N9569);
xor XOR2 (N11168, N11155, N10140);
nor NOR4 (N11169, N11157, N3973, N3071, N8844);
buf BUF1 (N11170, N11163);
not NOT1 (N11171, N11170);
nor NOR3 (N11172, N11167, N3019, N10059);
xor XOR2 (N11173, N11169, N10240);
not NOT1 (N11174, N11123);
buf BUF1 (N11175, N11171);
and AND2 (N11176, N11168, N10322);
or OR4 (N11177, N11174, N6875, N10845, N9700);
xor XOR2 (N11178, N11166, N7910);
xor XOR2 (N11179, N11178, N10452);
xor XOR2 (N11180, N11172, N2465);
nor NOR2 (N11181, N11175, N2794);
nand NAND2 (N11182, N11159, N7818);
xor XOR2 (N11183, N11173, N484);
and AND4 (N11184, N11162, N10134, N1431, N1395);
nor NOR2 (N11185, N11182, N4590);
or OR4 (N11186, N11179, N10581, N10288, N540);
nor NOR4 (N11187, N11160, N9326, N5912, N4936);
buf BUF1 (N11188, N11176);
buf BUF1 (N11189, N11186);
or OR4 (N11190, N11184, N4206, N194, N1321);
and AND2 (N11191, N11187, N2686);
and AND4 (N11192, N11181, N2278, N8239, N10177);
xor XOR2 (N11193, N11183, N10044);
xor XOR2 (N11194, N11161, N4986);
xor XOR2 (N11195, N11193, N10201);
xor XOR2 (N11196, N11177, N10471);
not NOT1 (N11197, N11180);
xor XOR2 (N11198, N11185, N5475);
buf BUF1 (N11199, N11198);
not NOT1 (N11200, N11190);
and AND2 (N11201, N11197, N2749);
and AND2 (N11202, N11189, N5068);
or OR2 (N11203, N11195, N1487);
or OR3 (N11204, N11203, N2410, N4867);
nor NOR3 (N11205, N11188, N2685, N11072);
xor XOR2 (N11206, N11204, N10075);
and AND4 (N11207, N11191, N9782, N8477, N9251);
nor NOR3 (N11208, N11207, N5574, N6769);
nor NOR4 (N11209, N11192, N2416, N10130, N9208);
nor NOR3 (N11210, N11199, N8560, N1929);
or OR2 (N11211, N11202, N8686);
not NOT1 (N11212, N11200);
and AND2 (N11213, N11205, N7309);
buf BUF1 (N11214, N11209);
or OR2 (N11215, N11214, N3987);
nor NOR2 (N11216, N11213, N2215);
nand NAND3 (N11217, N11212, N4119, N123);
nand NAND3 (N11218, N11210, N6276, N9583);
or OR3 (N11219, N11217, N2840, N6453);
nand NAND3 (N11220, N11218, N5222, N1772);
not NOT1 (N11221, N11220);
nand NAND2 (N11222, N11208, N754);
and AND3 (N11223, N11222, N6816, N1029);
buf BUF1 (N11224, N11211);
and AND2 (N11225, N11196, N5977);
nand NAND3 (N11226, N11216, N6749, N6149);
not NOT1 (N11227, N11206);
nor NOR3 (N11228, N11226, N10565, N4842);
or OR4 (N11229, N11221, N7875, N9444, N2386);
nand NAND4 (N11230, N11194, N5541, N6207, N10988);
nand NAND3 (N11231, N11215, N1855, N10353);
nand NAND2 (N11232, N11219, N5147);
buf BUF1 (N11233, N11228);
xor XOR2 (N11234, N11229, N1145);
nand NAND2 (N11235, N11225, N10543);
xor XOR2 (N11236, N11232, N8972);
nand NAND3 (N11237, N11231, N10492, N770);
xor XOR2 (N11238, N11236, N10389);
buf BUF1 (N11239, N11227);
buf BUF1 (N11240, N11234);
nand NAND3 (N11241, N11239, N7767, N4903);
or OR4 (N11242, N11240, N3801, N177, N8351);
nor NOR4 (N11243, N11233, N4888, N6953, N6692);
and AND4 (N11244, N11201, N6742, N4058, N7240);
nor NOR2 (N11245, N11224, N9035);
buf BUF1 (N11246, N11230);
nor NOR2 (N11247, N11238, N2501);
xor XOR2 (N11248, N11242, N10020);
nor NOR4 (N11249, N11244, N5239, N165, N5156);
xor XOR2 (N11250, N11223, N3171);
xor XOR2 (N11251, N11247, N4406);
buf BUF1 (N11252, N11251);
or OR4 (N11253, N11246, N7614, N9308, N5717);
or OR2 (N11254, N11245, N3270);
nor NOR2 (N11255, N11235, N9976);
not NOT1 (N11256, N11243);
buf BUF1 (N11257, N11254);
nor NOR3 (N11258, N11256, N1020, N10112);
or OR4 (N11259, N11237, N1578, N7251, N3996);
xor XOR2 (N11260, N11257, N5845);
nand NAND3 (N11261, N11248, N4081, N9068);
xor XOR2 (N11262, N11260, N1375);
or OR2 (N11263, N11261, N10262);
nor NOR4 (N11264, N11241, N5050, N7659, N2332);
nand NAND4 (N11265, N11253, N9141, N4522, N7684);
nor NOR3 (N11266, N11252, N7955, N8247);
and AND2 (N11267, N11249, N6181);
nor NOR2 (N11268, N11264, N127);
buf BUF1 (N11269, N11267);
xor XOR2 (N11270, N11255, N7041);
buf BUF1 (N11271, N11265);
and AND4 (N11272, N11266, N8751, N2074, N130);
not NOT1 (N11273, N11250);
or OR3 (N11274, N11270, N1035, N8338);
buf BUF1 (N11275, N11272);
not NOT1 (N11276, N11275);
buf BUF1 (N11277, N11259);
xor XOR2 (N11278, N11263, N8903);
nand NAND3 (N11279, N11271, N9186, N7338);
and AND4 (N11280, N11273, N9779, N8108, N4395);
or OR2 (N11281, N11268, N9820);
nor NOR3 (N11282, N11280, N185, N6252);
xor XOR2 (N11283, N11277, N9922);
nor NOR4 (N11284, N11274, N651, N1133, N5833);
or OR3 (N11285, N11283, N9202, N6401);
and AND2 (N11286, N11284, N5255);
xor XOR2 (N11287, N11262, N10226);
nor NOR4 (N11288, N11282, N9677, N10717, N7629);
or OR2 (N11289, N11286, N6709);
nand NAND2 (N11290, N11285, N5623);
nor NOR3 (N11291, N11269, N3297, N1516);
buf BUF1 (N11292, N11291);
nand NAND2 (N11293, N11290, N11030);
and AND2 (N11294, N11258, N9437);
or OR4 (N11295, N11294, N2529, N9279, N7640);
and AND3 (N11296, N11276, N1385, N1418);
not NOT1 (N11297, N11288);
xor XOR2 (N11298, N11292, N1696);
and AND2 (N11299, N11278, N3668);
nand NAND3 (N11300, N11297, N9191, N8840);
nand NAND2 (N11301, N11289, N5723);
xor XOR2 (N11302, N11298, N10253);
not NOT1 (N11303, N11287);
and AND2 (N11304, N11281, N322);
or OR4 (N11305, N11295, N6773, N637, N2108);
buf BUF1 (N11306, N11304);
not NOT1 (N11307, N11299);
nor NOR4 (N11308, N11300, N10878, N198, N3378);
xor XOR2 (N11309, N11308, N9576);
nand NAND4 (N11310, N11303, N4720, N6675, N959);
nor NOR4 (N11311, N11309, N5223, N6087, N9821);
xor XOR2 (N11312, N11311, N1363);
or OR2 (N11313, N11302, N3670);
nor NOR4 (N11314, N11296, N5831, N9375, N5686);
or OR4 (N11315, N11306, N3591, N4960, N4472);
nor NOR2 (N11316, N11279, N10209);
buf BUF1 (N11317, N11313);
nor NOR2 (N11318, N11307, N6235);
not NOT1 (N11319, N11305);
or OR4 (N11320, N11319, N4486, N3640, N1313);
buf BUF1 (N11321, N11314);
nand NAND2 (N11322, N11312, N9414);
nor NOR2 (N11323, N11317, N9395);
xor XOR2 (N11324, N11323, N7595);
not NOT1 (N11325, N11321);
not NOT1 (N11326, N11324);
nor NOR4 (N11327, N11320, N1564, N10461, N4511);
buf BUF1 (N11328, N11326);
and AND3 (N11329, N11322, N8222, N7229);
nor NOR2 (N11330, N11329, N6781);
buf BUF1 (N11331, N11310);
or OR3 (N11332, N11316, N7299, N9249);
nor NOR4 (N11333, N11293, N1752, N899, N386);
not NOT1 (N11334, N11330);
nand NAND4 (N11335, N11333, N7472, N3430, N3376);
and AND3 (N11336, N11328, N5430, N2835);
nor NOR4 (N11337, N11332, N8041, N2652, N11281);
buf BUF1 (N11338, N11337);
nand NAND2 (N11339, N11336, N5724);
nand NAND2 (N11340, N11339, N8185);
nor NOR3 (N11341, N11327, N7853, N4710);
and AND3 (N11342, N11301, N5322, N1754);
nor NOR4 (N11343, N11318, N6442, N1988, N362);
nand NAND2 (N11344, N11340, N147);
xor XOR2 (N11345, N11331, N1433);
or OR2 (N11346, N11341, N4714);
buf BUF1 (N11347, N11342);
nand NAND3 (N11348, N11315, N7156, N7038);
nor NOR3 (N11349, N11346, N9204, N5103);
not NOT1 (N11350, N11345);
or OR4 (N11351, N11338, N6419, N9249, N3307);
or OR3 (N11352, N11348, N3052, N5555);
buf BUF1 (N11353, N11344);
xor XOR2 (N11354, N11349, N3248);
and AND4 (N11355, N11350, N11233, N6423, N7616);
buf BUF1 (N11356, N11351);
and AND2 (N11357, N11352, N3223);
or OR3 (N11358, N11325, N469, N5471);
buf BUF1 (N11359, N11347);
buf BUF1 (N11360, N11358);
buf BUF1 (N11361, N11353);
or OR4 (N11362, N11354, N8559, N3054, N4491);
or OR4 (N11363, N11361, N9601, N9186, N4077);
nand NAND2 (N11364, N11334, N9614);
nor NOR2 (N11365, N11335, N10771);
and AND4 (N11366, N11359, N6035, N10212, N1438);
xor XOR2 (N11367, N11363, N4552);
and AND2 (N11368, N11362, N885);
nand NAND2 (N11369, N11356, N11176);
and AND4 (N11370, N11369, N7863, N3824, N3664);
not NOT1 (N11371, N11355);
nand NAND4 (N11372, N11370, N476, N182, N10767);
nand NAND3 (N11373, N11367, N1722, N9157);
not NOT1 (N11374, N11357);
nand NAND4 (N11375, N11373, N6228, N886, N7453);
buf BUF1 (N11376, N11364);
buf BUF1 (N11377, N11376);
and AND2 (N11378, N11372, N6196);
or OR2 (N11379, N11375, N7054);
nor NOR4 (N11380, N11378, N10775, N5412, N7859);
or OR2 (N11381, N11374, N4304);
nor NOR4 (N11382, N11377, N5301, N10982, N5724);
and AND3 (N11383, N11382, N6925, N3164);
buf BUF1 (N11384, N11383);
buf BUF1 (N11385, N11384);
nand NAND2 (N11386, N11381, N7519);
or OR2 (N11387, N11386, N9848);
xor XOR2 (N11388, N11365, N8608);
nor NOR4 (N11389, N11366, N7180, N1460, N599);
nand NAND2 (N11390, N11343, N811);
xor XOR2 (N11391, N11371, N3950);
xor XOR2 (N11392, N11389, N4312);
nor NOR4 (N11393, N11380, N4518, N9956, N5846);
xor XOR2 (N11394, N11385, N3934);
nand NAND3 (N11395, N11390, N6871, N224);
xor XOR2 (N11396, N11360, N9273);
not NOT1 (N11397, N11395);
nor NOR4 (N11398, N11393, N4357, N9123, N5321);
not NOT1 (N11399, N11368);
nand NAND4 (N11400, N11387, N597, N11210, N4444);
nand NAND3 (N11401, N11396, N301, N8546);
nor NOR4 (N11402, N11394, N3590, N10450, N3118);
and AND2 (N11403, N11399, N8667);
or OR2 (N11404, N11379, N4453);
xor XOR2 (N11405, N11401, N9822);
and AND2 (N11406, N11402, N2721);
or OR2 (N11407, N11388, N10743);
not NOT1 (N11408, N11404);
buf BUF1 (N11409, N11400);
xor XOR2 (N11410, N11406, N2102);
not NOT1 (N11411, N11408);
not NOT1 (N11412, N11407);
nand NAND2 (N11413, N11397, N5878);
nand NAND2 (N11414, N11392, N943);
nand NAND2 (N11415, N11403, N10046);
and AND2 (N11416, N11391, N5287);
not NOT1 (N11417, N11409);
and AND2 (N11418, N11414, N1921);
not NOT1 (N11419, N11418);
buf BUF1 (N11420, N11413);
and AND2 (N11421, N11420, N6031);
nand NAND3 (N11422, N11405, N8808, N1133);
or OR4 (N11423, N11421, N6135, N38, N8625);
nor NOR2 (N11424, N11416, N8711);
and AND3 (N11425, N11417, N8005, N4415);
xor XOR2 (N11426, N11412, N6709);
xor XOR2 (N11427, N11419, N10190);
xor XOR2 (N11428, N11424, N3538);
and AND2 (N11429, N11426, N4559);
nor NOR2 (N11430, N11425, N2252);
or OR2 (N11431, N11428, N3523);
nor NOR4 (N11432, N11411, N8801, N8829, N4747);
nor NOR3 (N11433, N11410, N8187, N3539);
buf BUF1 (N11434, N11415);
and AND3 (N11435, N11430, N443, N4665);
buf BUF1 (N11436, N11422);
nor NOR2 (N11437, N11434, N1323);
buf BUF1 (N11438, N11398);
nor NOR3 (N11439, N11431, N5437, N6413);
nand NAND2 (N11440, N11429, N8322);
xor XOR2 (N11441, N11440, N6022);
not NOT1 (N11442, N11437);
nor NOR4 (N11443, N11436, N5490, N10893, N6790);
buf BUF1 (N11444, N11438);
nand NAND3 (N11445, N11442, N3682, N7565);
buf BUF1 (N11446, N11443);
nand NAND4 (N11447, N11432, N673, N4880, N7290);
nor NOR4 (N11448, N11444, N7144, N10453, N5170);
or OR4 (N11449, N11433, N2726, N10292, N6679);
buf BUF1 (N11450, N11439);
xor XOR2 (N11451, N11441, N9784);
or OR2 (N11452, N11451, N7119);
or OR3 (N11453, N11448, N1514, N8083);
nor NOR3 (N11454, N11427, N2723, N2395);
or OR4 (N11455, N11423, N1350, N1831, N11040);
not NOT1 (N11456, N11445);
or OR2 (N11457, N11454, N8160);
or OR4 (N11458, N11449, N7357, N3268, N3899);
nor NOR3 (N11459, N11453, N7939, N94);
not NOT1 (N11460, N11456);
not NOT1 (N11461, N11452);
nand NAND4 (N11462, N11458, N4183, N5118, N4757);
not NOT1 (N11463, N11457);
nor NOR3 (N11464, N11450, N8796, N6746);
nand NAND2 (N11465, N11460, N1485);
nand NAND4 (N11466, N11465, N10054, N10385, N2403);
not NOT1 (N11467, N11466);
or OR2 (N11468, N11459, N4018);
buf BUF1 (N11469, N11461);
nor NOR3 (N11470, N11468, N6044, N1905);
not NOT1 (N11471, N11455);
or OR4 (N11472, N11467, N3723, N2879, N7509);
buf BUF1 (N11473, N11471);
and AND2 (N11474, N11462, N5952);
buf BUF1 (N11475, N11474);
not NOT1 (N11476, N11446);
nor NOR2 (N11477, N11472, N1320);
not NOT1 (N11478, N11470);
and AND4 (N11479, N11469, N8322, N5251, N2981);
nand NAND4 (N11480, N11463, N9088, N5418, N8332);
nor NOR2 (N11481, N11475, N9745);
nand NAND3 (N11482, N11477, N11196, N4888);
buf BUF1 (N11483, N11447);
xor XOR2 (N11484, N11476, N5316);
nand NAND3 (N11485, N11478, N2305, N467);
nand NAND4 (N11486, N11473, N8067, N10300, N6144);
xor XOR2 (N11487, N11480, N2852);
nor NOR4 (N11488, N11484, N199, N3081, N55);
nand NAND4 (N11489, N11479, N7674, N1060, N559);
or OR3 (N11490, N11435, N277, N3676);
not NOT1 (N11491, N11483);
or OR4 (N11492, N11488, N9261, N3344, N6747);
nand NAND2 (N11493, N11492, N837);
xor XOR2 (N11494, N11491, N4975);
nor NOR3 (N11495, N11489, N5694, N4991);
nor NOR4 (N11496, N11495, N5974, N1939, N9756);
not NOT1 (N11497, N11481);
buf BUF1 (N11498, N11496);
not NOT1 (N11499, N11464);
buf BUF1 (N11500, N11485);
and AND3 (N11501, N11490, N1937, N3448);
buf BUF1 (N11502, N11487);
buf BUF1 (N11503, N11500);
or OR3 (N11504, N11493, N10659, N7209);
nor NOR2 (N11505, N11497, N5095);
nand NAND3 (N11506, N11503, N9050, N1088);
and AND4 (N11507, N11486, N3162, N3840, N9331);
nor NOR2 (N11508, N11502, N6851);
or OR4 (N11509, N11482, N7418, N4221, N7128);
or OR2 (N11510, N11505, N9639);
nand NAND3 (N11511, N11506, N4008, N690);
nor NOR3 (N11512, N11501, N10791, N8417);
not NOT1 (N11513, N11508);
nor NOR3 (N11514, N11498, N8192, N6748);
nand NAND2 (N11515, N11512, N7923);
xor XOR2 (N11516, N11499, N3980);
not NOT1 (N11517, N11507);
xor XOR2 (N11518, N11514, N7244);
buf BUF1 (N11519, N11504);
and AND4 (N11520, N11510, N7396, N7484, N5421);
nand NAND2 (N11521, N11520, N1519);
xor XOR2 (N11522, N11516, N438);
nand NAND4 (N11523, N11521, N2182, N5645, N2466);
and AND3 (N11524, N11517, N8230, N9953);
or OR2 (N11525, N11511, N8623);
nor NOR3 (N11526, N11494, N6387, N9499);
nor NOR3 (N11527, N11519, N4278, N2921);
nand NAND4 (N11528, N11526, N5986, N5175, N7072);
buf BUF1 (N11529, N11522);
not NOT1 (N11530, N11509);
buf BUF1 (N11531, N11513);
buf BUF1 (N11532, N11518);
or OR4 (N11533, N11531, N7991, N4554, N10516);
buf BUF1 (N11534, N11515);
xor XOR2 (N11535, N11524, N4582);
xor XOR2 (N11536, N11530, N8310);
or OR3 (N11537, N11533, N2087, N10425);
or OR2 (N11538, N11528, N3900);
xor XOR2 (N11539, N11527, N4153);
nand NAND3 (N11540, N11538, N10845, N10034);
and AND4 (N11541, N11537, N5286, N10524, N3397);
and AND2 (N11542, N11541, N2412);
xor XOR2 (N11543, N11534, N6993);
nand NAND2 (N11544, N11532, N4054);
nand NAND4 (N11545, N11525, N7315, N816, N442);
nand NAND3 (N11546, N11543, N2859, N4728);
nand NAND2 (N11547, N11546, N3622);
nor NOR3 (N11548, N11544, N7007, N850);
nor NOR4 (N11549, N11529, N9237, N4847, N659);
buf BUF1 (N11550, N11545);
not NOT1 (N11551, N11549);
and AND4 (N11552, N11542, N4380, N7353, N4405);
xor XOR2 (N11553, N11535, N5637);
nor NOR2 (N11554, N11550, N6380);
or OR3 (N11555, N11553, N3215, N7322);
xor XOR2 (N11556, N11548, N5904);
not NOT1 (N11557, N11552);
buf BUF1 (N11558, N11539);
not NOT1 (N11559, N11555);
nor NOR3 (N11560, N11557, N569, N1474);
or OR4 (N11561, N11558, N4796, N6093, N3792);
nor NOR4 (N11562, N11523, N3138, N1607, N4929);
xor XOR2 (N11563, N11560, N11158);
not NOT1 (N11564, N11554);
and AND2 (N11565, N11547, N7440);
nor NOR2 (N11566, N11540, N4562);
not NOT1 (N11567, N11556);
nand NAND4 (N11568, N11562, N11264, N8513, N6224);
nand NAND4 (N11569, N11564, N2157, N10605, N8739);
or OR4 (N11570, N11565, N2476, N3495, N3390);
buf BUF1 (N11571, N11559);
or OR4 (N11572, N11568, N4628, N5215, N1984);
and AND2 (N11573, N11566, N2102);
buf BUF1 (N11574, N11573);
xor XOR2 (N11575, N11569, N9398);
or OR3 (N11576, N11536, N9188, N10596);
or OR3 (N11577, N11576, N9423, N3987);
xor XOR2 (N11578, N11561, N193);
buf BUF1 (N11579, N11551);
or OR4 (N11580, N11577, N4672, N512, N6617);
not NOT1 (N11581, N11580);
buf BUF1 (N11582, N11578);
nand NAND2 (N11583, N11567, N9601);
not NOT1 (N11584, N11581);
nand NAND3 (N11585, N11583, N7673, N1911);
and AND3 (N11586, N11582, N3256, N7016);
buf BUF1 (N11587, N11579);
not NOT1 (N11588, N11570);
or OR4 (N11589, N11585, N6709, N9344, N9199);
not NOT1 (N11590, N11589);
buf BUF1 (N11591, N11574);
or OR3 (N11592, N11586, N4760, N7780);
nand NAND4 (N11593, N11563, N565, N7858, N5492);
xor XOR2 (N11594, N11592, N2584);
nand NAND2 (N11595, N11591, N4270);
nor NOR3 (N11596, N11584, N8338, N10216);
nand NAND3 (N11597, N11572, N4331, N4820);
xor XOR2 (N11598, N11596, N7967);
xor XOR2 (N11599, N11598, N6685);
buf BUF1 (N11600, N11587);
and AND4 (N11601, N11594, N8120, N10267, N66);
xor XOR2 (N11602, N11601, N11429);
nand NAND3 (N11603, N11599, N2028, N4171);
not NOT1 (N11604, N11597);
xor XOR2 (N11605, N11603, N11342);
nor NOR4 (N11606, N11604, N7297, N3275, N9390);
xor XOR2 (N11607, N11571, N10695);
or OR4 (N11608, N11595, N5086, N1885, N3562);
nor NOR3 (N11609, N11602, N2304, N4500);
buf BUF1 (N11610, N11607);
nor NOR2 (N11611, N11605, N9133);
and AND2 (N11612, N11575, N9646);
nand NAND4 (N11613, N11600, N1442, N10054, N4052);
and AND4 (N11614, N11606, N3630, N282, N1917);
nor NOR3 (N11615, N11614, N4934, N9522);
and AND2 (N11616, N11611, N306);
nor NOR3 (N11617, N11612, N5195, N5000);
xor XOR2 (N11618, N11616, N523);
nand NAND2 (N11619, N11615, N6349);
xor XOR2 (N11620, N11618, N3782);
not NOT1 (N11621, N11613);
xor XOR2 (N11622, N11608, N313);
and AND3 (N11623, N11620, N2536, N2669);
not NOT1 (N11624, N11617);
nand NAND3 (N11625, N11623, N4051, N9960);
xor XOR2 (N11626, N11621, N6312);
nor NOR4 (N11627, N11590, N7053, N9493, N9594);
xor XOR2 (N11628, N11624, N4637);
nor NOR3 (N11629, N11627, N1585, N8614);
nor NOR4 (N11630, N11622, N6395, N5278, N6390);
xor XOR2 (N11631, N11588, N291);
nor NOR2 (N11632, N11631, N10361);
buf BUF1 (N11633, N11609);
and AND2 (N11634, N11619, N2629);
nand NAND4 (N11635, N11628, N1996, N11615, N2046);
nor NOR2 (N11636, N11593, N4599);
or OR3 (N11637, N11635, N10188, N9918);
xor XOR2 (N11638, N11625, N9124);
nor NOR4 (N11639, N11637, N7936, N4827, N5666);
and AND4 (N11640, N11610, N7904, N2124, N643);
xor XOR2 (N11641, N11629, N8533);
xor XOR2 (N11642, N11640, N2104);
or OR3 (N11643, N11632, N9943, N6064);
xor XOR2 (N11644, N11643, N349);
nor NOR4 (N11645, N11636, N4171, N9970, N2568);
nor NOR4 (N11646, N11641, N10890, N1573, N5403);
or OR4 (N11647, N11630, N1140, N4409, N4225);
xor XOR2 (N11648, N11639, N10385);
nand NAND2 (N11649, N11644, N6175);
or OR3 (N11650, N11646, N4648, N299);
buf BUF1 (N11651, N11626);
nand NAND2 (N11652, N11648, N8054);
and AND4 (N11653, N11633, N220, N8283, N10136);
buf BUF1 (N11654, N11634);
nor NOR3 (N11655, N11645, N5383, N3666);
nor NOR2 (N11656, N11647, N8551);
not NOT1 (N11657, N11650);
nand NAND3 (N11658, N11655, N4642, N1454);
or OR2 (N11659, N11654, N427);
or OR4 (N11660, N11659, N4386, N1435, N10627);
not NOT1 (N11661, N11652);
nand NAND4 (N11662, N11658, N6887, N5393, N9715);
nor NOR2 (N11663, N11649, N10532);
not NOT1 (N11664, N11638);
and AND3 (N11665, N11660, N11137, N2969);
nor NOR4 (N11666, N11656, N4439, N8514, N7382);
or OR2 (N11667, N11651, N6012);
nand NAND2 (N11668, N11667, N11470);
buf BUF1 (N11669, N11657);
or OR2 (N11670, N11665, N10451);
nand NAND3 (N11671, N11642, N824, N5439);
and AND4 (N11672, N11661, N5066, N9808, N7054);
buf BUF1 (N11673, N11668);
and AND4 (N11674, N11663, N3361, N10695, N10520);
buf BUF1 (N11675, N11670);
nand NAND3 (N11676, N11674, N8452, N3610);
not NOT1 (N11677, N11666);
and AND3 (N11678, N11675, N3032, N3889);
nand NAND2 (N11679, N11677, N11303);
or OR4 (N11680, N11662, N3769, N6159, N29);
nand NAND4 (N11681, N11678, N7734, N4896, N6788);
and AND2 (N11682, N11653, N9707);
not NOT1 (N11683, N11671);
or OR2 (N11684, N11682, N11413);
nor NOR3 (N11685, N11681, N7758, N9806);
not NOT1 (N11686, N11683);
nor NOR4 (N11687, N11686, N2230, N10727, N11383);
buf BUF1 (N11688, N11672);
or OR4 (N11689, N11687, N3109, N2271, N9169);
buf BUF1 (N11690, N11673);
nand NAND4 (N11691, N11688, N10250, N894, N11058);
or OR3 (N11692, N11669, N4230, N4766);
nor NOR2 (N11693, N11685, N6570);
nor NOR4 (N11694, N11676, N6871, N7922, N10673);
xor XOR2 (N11695, N11680, N354);
not NOT1 (N11696, N11691);
xor XOR2 (N11697, N11696, N9195);
or OR2 (N11698, N11684, N8874);
and AND2 (N11699, N11679, N3756);
nand NAND4 (N11700, N11695, N310, N2334, N1579);
not NOT1 (N11701, N11664);
or OR4 (N11702, N11689, N10558, N4421, N11299);
buf BUF1 (N11703, N11690);
not NOT1 (N11704, N11699);
nor NOR4 (N11705, N11698, N8490, N9015, N6590);
nand NAND4 (N11706, N11701, N1199, N3457, N5497);
not NOT1 (N11707, N11704);
not NOT1 (N11708, N11702);
nand NAND3 (N11709, N11707, N3846, N3875);
buf BUF1 (N11710, N11697);
xor XOR2 (N11711, N11705, N7121);
nor NOR2 (N11712, N11693, N4294);
nor NOR3 (N11713, N11692, N1236, N6827);
not NOT1 (N11714, N11708);
not NOT1 (N11715, N11703);
nand NAND4 (N11716, N11694, N255, N10378, N1465);
and AND4 (N11717, N11700, N5722, N7012, N8392);
buf BUF1 (N11718, N11706);
buf BUF1 (N11719, N11714);
and AND2 (N11720, N11718, N4868);
xor XOR2 (N11721, N11716, N7964);
xor XOR2 (N11722, N11719, N4135);
or OR3 (N11723, N11717, N1018, N3768);
or OR4 (N11724, N11723, N8360, N6270, N1358);
or OR2 (N11725, N11713, N10764);
not NOT1 (N11726, N11712);
or OR3 (N11727, N11722, N9762, N2223);
nand NAND2 (N11728, N11720, N10222);
or OR3 (N11729, N11727, N6239, N9310);
nand NAND4 (N11730, N11710, N1179, N5819, N5670);
and AND2 (N11731, N11729, N7184);
nand NAND2 (N11732, N11726, N11281);
buf BUF1 (N11733, N11731);
xor XOR2 (N11734, N11711, N550);
nand NAND3 (N11735, N11728, N9818, N7624);
nor NOR2 (N11736, N11709, N6476);
not NOT1 (N11737, N11732);
and AND2 (N11738, N11724, N10408);
and AND4 (N11739, N11736, N105, N3502, N3216);
and AND4 (N11740, N11721, N2845, N10824, N1802);
not NOT1 (N11741, N11715);
buf BUF1 (N11742, N11725);
and AND2 (N11743, N11735, N10052);
nand NAND2 (N11744, N11738, N11711);
xor XOR2 (N11745, N11744, N6363);
and AND4 (N11746, N11734, N10871, N10241, N4084);
buf BUF1 (N11747, N11739);
nor NOR3 (N11748, N11747, N6914, N8681);
nand NAND4 (N11749, N11742, N2375, N1010, N6355);
not NOT1 (N11750, N11740);
buf BUF1 (N11751, N11748);
buf BUF1 (N11752, N11745);
nand NAND3 (N11753, N11743, N2218, N2001);
nor NOR2 (N11754, N11753, N9818);
or OR3 (N11755, N11752, N6989, N9704);
nand NAND3 (N11756, N11741, N11353, N1255);
not NOT1 (N11757, N11750);
nor NOR4 (N11758, N11751, N7220, N1908, N10122);
xor XOR2 (N11759, N11737, N285);
or OR3 (N11760, N11756, N3966, N7275);
not NOT1 (N11761, N11730);
xor XOR2 (N11762, N11733, N10770);
xor XOR2 (N11763, N11758, N3527);
xor XOR2 (N11764, N11762, N6604);
nor NOR4 (N11765, N11755, N8951, N7824, N11195);
nor NOR3 (N11766, N11746, N2966, N3087);
nand NAND4 (N11767, N11766, N11058, N9712, N234);
nor NOR2 (N11768, N11765, N5247);
or OR4 (N11769, N11767, N5082, N7951, N6333);
not NOT1 (N11770, N11757);
not NOT1 (N11771, N11754);
nand NAND2 (N11772, N11764, N6735);
not NOT1 (N11773, N11771);
nor NOR3 (N11774, N11749, N388, N7916);
nand NAND3 (N11775, N11760, N5307, N1909);
nand NAND2 (N11776, N11759, N9356);
xor XOR2 (N11777, N11761, N3966);
xor XOR2 (N11778, N11769, N7719);
buf BUF1 (N11779, N11773);
buf BUF1 (N11780, N11763);
nand NAND4 (N11781, N11774, N3111, N996, N3764);
and AND2 (N11782, N11772, N11736);
and AND2 (N11783, N11768, N7741);
and AND4 (N11784, N11779, N3624, N10665, N1470);
not NOT1 (N11785, N11783);
nand NAND4 (N11786, N11784, N9113, N52, N3453);
xor XOR2 (N11787, N11778, N2829);
nor NOR4 (N11788, N11780, N9447, N6440, N4422);
xor XOR2 (N11789, N11781, N4976);
not NOT1 (N11790, N11775);
xor XOR2 (N11791, N11788, N6956);
nand NAND4 (N11792, N11790, N219, N6773, N5128);
xor XOR2 (N11793, N11785, N1953);
and AND2 (N11794, N11776, N3928);
buf BUF1 (N11795, N11789);
buf BUF1 (N11796, N11793);
nand NAND4 (N11797, N11794, N10976, N1704, N2956);
not NOT1 (N11798, N11787);
nor NOR3 (N11799, N11786, N2945, N2338);
nand NAND3 (N11800, N11770, N5528, N5159);
buf BUF1 (N11801, N11798);
or OR2 (N11802, N11792, N7836);
and AND2 (N11803, N11791, N7051);
nand NAND2 (N11804, N11777, N2224);
nor NOR4 (N11805, N11800, N3689, N4354, N1579);
not NOT1 (N11806, N11802);
buf BUF1 (N11807, N11796);
and AND3 (N11808, N11807, N11598, N4889);
xor XOR2 (N11809, N11797, N11213);
or OR3 (N11810, N11809, N9306, N5756);
buf BUF1 (N11811, N11799);
buf BUF1 (N11812, N11782);
nand NAND2 (N11813, N11805, N4165);
xor XOR2 (N11814, N11810, N11023);
nor NOR4 (N11815, N11804, N6100, N8287, N11329);
xor XOR2 (N11816, N11814, N418);
buf BUF1 (N11817, N11795);
or OR4 (N11818, N11806, N11023, N5939, N3639);
and AND2 (N11819, N11812, N4765);
xor XOR2 (N11820, N11808, N6713);
xor XOR2 (N11821, N11811, N6537);
or OR4 (N11822, N11818, N10789, N7417, N1018);
or OR4 (N11823, N11816, N6969, N9454, N5479);
not NOT1 (N11824, N11819);
or OR3 (N11825, N11824, N3082, N8185);
buf BUF1 (N11826, N11823);
xor XOR2 (N11827, N11825, N7820);
buf BUF1 (N11828, N11827);
nand NAND4 (N11829, N11801, N8251, N10078, N7714);
not NOT1 (N11830, N11821);
nor NOR3 (N11831, N11817, N5287, N1067);
nand NAND3 (N11832, N11829, N7487, N3096);
buf BUF1 (N11833, N11832);
nand NAND2 (N11834, N11833, N8458);
not NOT1 (N11835, N11831);
buf BUF1 (N11836, N11828);
nand NAND3 (N11837, N11820, N491, N8387);
xor XOR2 (N11838, N11803, N4776);
and AND4 (N11839, N11830, N2898, N9604, N11753);
buf BUF1 (N11840, N11835);
buf BUF1 (N11841, N11836);
not NOT1 (N11842, N11838);
xor XOR2 (N11843, N11834, N9142);
xor XOR2 (N11844, N11843, N5610);
xor XOR2 (N11845, N11840, N4352);
or OR2 (N11846, N11815, N10286);
xor XOR2 (N11847, N11839, N6009);
nand NAND3 (N11848, N11841, N1749, N713);
and AND2 (N11849, N11813, N9695);
and AND2 (N11850, N11845, N5756);
nand NAND2 (N11851, N11846, N11265);
nor NOR4 (N11852, N11848, N2916, N4465, N547);
buf BUF1 (N11853, N11852);
nor NOR2 (N11854, N11850, N3302);
xor XOR2 (N11855, N11849, N3734);
and AND4 (N11856, N11847, N9359, N4903, N8583);
not NOT1 (N11857, N11822);
nor NOR4 (N11858, N11844, N7385, N10016, N7974);
xor XOR2 (N11859, N11842, N2307);
xor XOR2 (N11860, N11857, N9589);
and AND2 (N11861, N11837, N8936);
nor NOR4 (N11862, N11853, N9619, N261, N8473);
and AND4 (N11863, N11858, N4016, N5655, N9329);
xor XOR2 (N11864, N11862, N8829);
xor XOR2 (N11865, N11826, N1178);
or OR4 (N11866, N11864, N5771, N1448, N11599);
buf BUF1 (N11867, N11859);
not NOT1 (N11868, N11865);
or OR4 (N11869, N11863, N10177, N9518, N4733);
buf BUF1 (N11870, N11854);
or OR3 (N11871, N11855, N10038, N11685);
buf BUF1 (N11872, N11851);
xor XOR2 (N11873, N11871, N11017);
nor NOR4 (N11874, N11867, N2254, N9488, N4003);
and AND3 (N11875, N11868, N9951, N2720);
not NOT1 (N11876, N11856);
not NOT1 (N11877, N11872);
nor NOR2 (N11878, N11870, N6010);
nor NOR2 (N11879, N11877, N1835);
not NOT1 (N11880, N11869);
nor NOR4 (N11881, N11879, N1088, N9279, N2466);
not NOT1 (N11882, N11878);
xor XOR2 (N11883, N11861, N4019);
or OR3 (N11884, N11873, N7098, N3170);
nand NAND3 (N11885, N11883, N7038, N615);
nand NAND2 (N11886, N11884, N8433);
nand NAND4 (N11887, N11885, N11029, N10677, N2528);
or OR2 (N11888, N11874, N7313);
nor NOR4 (N11889, N11860, N9881, N4719, N2248);
nor NOR2 (N11890, N11881, N2149);
nor NOR2 (N11891, N11882, N8262);
xor XOR2 (N11892, N11887, N1921);
xor XOR2 (N11893, N11888, N770);
and AND2 (N11894, N11880, N10095);
or OR3 (N11895, N11891, N6369, N2697);
or OR4 (N11896, N11876, N11369, N4206, N10780);
not NOT1 (N11897, N11896);
and AND4 (N11898, N11897, N5243, N10013, N8431);
nand NAND3 (N11899, N11866, N5404, N7739);
or OR3 (N11900, N11890, N7868, N1722);
nand NAND2 (N11901, N11892, N11148);
nand NAND3 (N11902, N11900, N4958, N4155);
buf BUF1 (N11903, N11902);
nor NOR4 (N11904, N11875, N8285, N9653, N8152);
nand NAND4 (N11905, N11899, N11096, N1691, N1838);
or OR3 (N11906, N11895, N10225, N10472);
and AND3 (N11907, N11898, N2060, N10123);
buf BUF1 (N11908, N11901);
nand NAND4 (N11909, N11904, N9395, N1427, N3139);
or OR4 (N11910, N11907, N2312, N1996, N10144);
xor XOR2 (N11911, N11894, N2528);
xor XOR2 (N11912, N11893, N5047);
xor XOR2 (N11913, N11909, N3271);
or OR2 (N11914, N11912, N8406);
or OR4 (N11915, N11910, N3282, N11879, N8568);
buf BUF1 (N11916, N11915);
and AND2 (N11917, N11886, N9881);
nand NAND4 (N11918, N11916, N4942, N10228, N9045);
not NOT1 (N11919, N11906);
buf BUF1 (N11920, N11913);
nor NOR3 (N11921, N11911, N6026, N11809);
or OR3 (N11922, N11919, N6453, N3799);
buf BUF1 (N11923, N11917);
and AND4 (N11924, N11918, N6849, N2635, N8434);
nor NOR3 (N11925, N11920, N6491, N6792);
or OR2 (N11926, N11903, N10618);
xor XOR2 (N11927, N11922, N7498);
nor NOR2 (N11928, N11905, N8691);
nand NAND2 (N11929, N11908, N826);
and AND4 (N11930, N11929, N10304, N8102, N8913);
not NOT1 (N11931, N11921);
buf BUF1 (N11932, N11924);
buf BUF1 (N11933, N11926);
xor XOR2 (N11934, N11923, N7741);
nand NAND4 (N11935, N11914, N11018, N9147, N6046);
nand NAND3 (N11936, N11935, N11758, N10338);
nor NOR4 (N11937, N11889, N6315, N5774, N4378);
buf BUF1 (N11938, N11930);
nor NOR4 (N11939, N11927, N7663, N3277, N9908);
nor NOR4 (N11940, N11937, N2989, N4492, N7662);
nand NAND4 (N11941, N11940, N6156, N11066, N5581);
or OR4 (N11942, N11932, N7622, N9030, N11270);
nand NAND3 (N11943, N11938, N743, N11623);
nor NOR2 (N11944, N11928, N4680);
nand NAND2 (N11945, N11934, N2622);
or OR4 (N11946, N11943, N11229, N6802, N6829);
and AND2 (N11947, N11942, N1169);
and AND2 (N11948, N11945, N3102);
nor NOR3 (N11949, N11941, N9519, N1544);
buf BUF1 (N11950, N11939);
nor NOR4 (N11951, N11925, N4536, N3248, N9887);
not NOT1 (N11952, N11949);
nor NOR4 (N11953, N11946, N1881, N10807, N7215);
and AND2 (N11954, N11944, N28);
buf BUF1 (N11955, N11951);
and AND3 (N11956, N11948, N3244, N9115);
xor XOR2 (N11957, N11947, N8919);
and AND2 (N11958, N11954, N7023);
buf BUF1 (N11959, N11936);
buf BUF1 (N11960, N11955);
or OR2 (N11961, N11953, N2445);
and AND2 (N11962, N11933, N5752);
and AND3 (N11963, N11956, N10634, N4427);
nor NOR2 (N11964, N11957, N10748);
nand NAND2 (N11965, N11961, N175);
nand NAND3 (N11966, N11950, N2102, N1887);
not NOT1 (N11967, N11966);
and AND3 (N11968, N11958, N5311, N3541);
not NOT1 (N11969, N11964);
or OR2 (N11970, N11963, N2219);
nor NOR2 (N11971, N11960, N139);
and AND3 (N11972, N11952, N9529, N9521);
xor XOR2 (N11973, N11971, N7835);
buf BUF1 (N11974, N11931);
not NOT1 (N11975, N11970);
not NOT1 (N11976, N11975);
buf BUF1 (N11977, N11976);
not NOT1 (N11978, N11974);
and AND2 (N11979, N11969, N1971);
nand NAND2 (N11980, N11979, N11463);
or OR2 (N11981, N11965, N3884);
or OR4 (N11982, N11959, N10551, N5736, N426);
xor XOR2 (N11983, N11981, N3036);
xor XOR2 (N11984, N11973, N4965);
buf BUF1 (N11985, N11977);
or OR3 (N11986, N11983, N8086, N4540);
or OR3 (N11987, N11980, N8901, N2554);
not NOT1 (N11988, N11982);
nor NOR2 (N11989, N11986, N872);
nand NAND4 (N11990, N11962, N552, N10784, N5550);
and AND4 (N11991, N11984, N2780, N9724, N7725);
not NOT1 (N11992, N11988);
and AND2 (N11993, N11978, N1865);
or OR4 (N11994, N11991, N3344, N8321, N8821);
nand NAND3 (N11995, N11993, N11496, N1598);
nor NOR2 (N11996, N11968, N4412);
not NOT1 (N11997, N11987);
and AND2 (N11998, N11995, N2746);
not NOT1 (N11999, N11997);
nand NAND2 (N12000, N11989, N7994);
xor XOR2 (N12001, N11996, N1462);
buf BUF1 (N12002, N11985);
not NOT1 (N12003, N11990);
or OR2 (N12004, N11998, N8677);
nand NAND3 (N12005, N12004, N7459, N2632);
buf BUF1 (N12006, N12001);
xor XOR2 (N12007, N11967, N6703);
and AND3 (N12008, N12007, N4860, N1348);
or OR2 (N12009, N11972, N9336);
buf BUF1 (N12010, N12003);
nand NAND4 (N12011, N12005, N1933, N492, N6668);
or OR4 (N12012, N12002, N11849, N5209, N615);
not NOT1 (N12013, N11994);
and AND2 (N12014, N12000, N11669);
and AND4 (N12015, N12006, N11407, N8590, N4668);
or OR3 (N12016, N12014, N7750, N6620);
and AND3 (N12017, N12012, N8330, N3104);
and AND4 (N12018, N12011, N11441, N2135, N856);
buf BUF1 (N12019, N12010);
or OR2 (N12020, N12013, N9413);
not NOT1 (N12021, N12017);
nand NAND3 (N12022, N11992, N8443, N6209);
or OR4 (N12023, N12018, N7400, N2602, N7107);
nand NAND2 (N12024, N12020, N6384);
buf BUF1 (N12025, N12024);
buf BUF1 (N12026, N12025);
nor NOR3 (N12027, N12015, N10629, N4032);
buf BUF1 (N12028, N12021);
and AND2 (N12029, N12026, N3664);
buf BUF1 (N12030, N12008);
xor XOR2 (N12031, N12016, N4534);
or OR3 (N12032, N12030, N9653, N4103);
or OR2 (N12033, N12032, N10298);
nor NOR4 (N12034, N12029, N10583, N4908, N6644);
nand NAND4 (N12035, N12034, N9429, N9778, N2579);
buf BUF1 (N12036, N12019);
xor XOR2 (N12037, N11999, N8277);
and AND2 (N12038, N12035, N816);
nand NAND4 (N12039, N12023, N3765, N2614, N4540);
or OR3 (N12040, N12036, N9842, N6508);
xor XOR2 (N12041, N12027, N8523);
xor XOR2 (N12042, N12039, N8107);
and AND2 (N12043, N12037, N6183);
nor NOR2 (N12044, N12028, N6040);
buf BUF1 (N12045, N12031);
or OR2 (N12046, N12044, N9449);
not NOT1 (N12047, N12022);
or OR4 (N12048, N12042, N1011, N3132, N3591);
or OR4 (N12049, N12040, N2056, N5802, N10810);
nand NAND2 (N12050, N12041, N4907);
buf BUF1 (N12051, N12049);
buf BUF1 (N12052, N12009);
or OR4 (N12053, N12043, N7167, N6751, N5055);
and AND2 (N12054, N12045, N3937);
nand NAND3 (N12055, N12052, N5743, N8893);
nor NOR2 (N12056, N12053, N9215);
and AND2 (N12057, N12038, N1363);
and AND2 (N12058, N12048, N5057);
nor NOR4 (N12059, N12033, N6469, N6606, N3360);
or OR2 (N12060, N12051, N11045);
not NOT1 (N12061, N12057);
nand NAND3 (N12062, N12055, N4473, N3305);
nand NAND4 (N12063, N12046, N8021, N7977, N6455);
and AND3 (N12064, N12061, N2167, N915);
buf BUF1 (N12065, N12058);
buf BUF1 (N12066, N12047);
nand NAND3 (N12067, N12050, N3722, N4960);
and AND4 (N12068, N12066, N1487, N1275, N8210);
not NOT1 (N12069, N12056);
nand NAND4 (N12070, N12069, N3647, N6146, N7385);
and AND4 (N12071, N12060, N7610, N11200, N474);
and AND4 (N12072, N12054, N3203, N6159, N1332);
buf BUF1 (N12073, N12071);
buf BUF1 (N12074, N12070);
xor XOR2 (N12075, N12073, N7879);
and AND2 (N12076, N12075, N3266);
nand NAND2 (N12077, N12062, N4705);
xor XOR2 (N12078, N12076, N7344);
buf BUF1 (N12079, N12068);
nor NOR2 (N12080, N12077, N395);
buf BUF1 (N12081, N12064);
not NOT1 (N12082, N12080);
not NOT1 (N12083, N12074);
xor XOR2 (N12084, N12079, N684);
not NOT1 (N12085, N12081);
buf BUF1 (N12086, N12063);
buf BUF1 (N12087, N12078);
buf BUF1 (N12088, N12059);
buf BUF1 (N12089, N12065);
nand NAND2 (N12090, N12086, N9078);
or OR4 (N12091, N12083, N10654, N5628, N6714);
nor NOR2 (N12092, N12084, N1367);
xor XOR2 (N12093, N12089, N7279);
or OR3 (N12094, N12092, N5420, N2259);
nand NAND3 (N12095, N12087, N5749, N8223);
buf BUF1 (N12096, N12082);
nor NOR2 (N12097, N12091, N11707);
xor XOR2 (N12098, N12090, N2220);
nor NOR2 (N12099, N12072, N80);
nand NAND2 (N12100, N12096, N10074);
xor XOR2 (N12101, N12094, N11681);
or OR2 (N12102, N12085, N10070);
and AND4 (N12103, N12067, N5443, N6292, N1210);
nor NOR3 (N12104, N12100, N11225, N9993);
buf BUF1 (N12105, N12099);
nor NOR4 (N12106, N12097, N4529, N3075, N8453);
nand NAND2 (N12107, N12095, N5465);
nor NOR3 (N12108, N12103, N8727, N568);
nand NAND3 (N12109, N12106, N375, N2099);
nor NOR2 (N12110, N12093, N7686);
not NOT1 (N12111, N12101);
nor NOR3 (N12112, N12098, N8715, N1117);
or OR4 (N12113, N12104, N10289, N2403, N2749);
nand NAND2 (N12114, N12111, N7389);
not NOT1 (N12115, N12108);
buf BUF1 (N12116, N12112);
nand NAND4 (N12117, N12115, N553, N10244, N7036);
buf BUF1 (N12118, N12107);
xor XOR2 (N12119, N12110, N10362);
nor NOR2 (N12120, N12102, N1704);
and AND2 (N12121, N12114, N1027);
not NOT1 (N12122, N12116);
nor NOR4 (N12123, N12105, N10461, N11540, N2952);
nand NAND3 (N12124, N12122, N8417, N2419);
or OR4 (N12125, N12123, N2436, N9559, N7934);
buf BUF1 (N12126, N12113);
not NOT1 (N12127, N12118);
nor NOR2 (N12128, N12088, N4309);
and AND3 (N12129, N12124, N6942, N8026);
nand NAND2 (N12130, N12120, N11018);
xor XOR2 (N12131, N12119, N6923);
nor NOR4 (N12132, N12129, N5416, N11196, N1262);
xor XOR2 (N12133, N12130, N10555);
xor XOR2 (N12134, N12131, N10170);
nand NAND2 (N12135, N12128, N3840);
nor NOR3 (N12136, N12126, N6955, N2398);
buf BUF1 (N12137, N12125);
nor NOR3 (N12138, N12135, N7599, N11443);
and AND2 (N12139, N12137, N3201);
and AND4 (N12140, N12127, N7763, N251, N9796);
buf BUF1 (N12141, N12139);
nor NOR4 (N12142, N12134, N793, N4774, N2317);
not NOT1 (N12143, N12141);
not NOT1 (N12144, N12143);
xor XOR2 (N12145, N12138, N794);
or OR3 (N12146, N12144, N9345, N8879);
not NOT1 (N12147, N12142);
xor XOR2 (N12148, N12145, N6705);
or OR2 (N12149, N12133, N7156);
buf BUF1 (N12150, N12146);
not NOT1 (N12151, N12136);
nor NOR2 (N12152, N12147, N2130);
nand NAND3 (N12153, N12152, N5304, N1908);
nand NAND3 (N12154, N12153, N3183, N10604);
not NOT1 (N12155, N12109);
or OR2 (N12156, N12155, N6143);
or OR4 (N12157, N12140, N6628, N511, N7160);
or OR4 (N12158, N12157, N4387, N9254, N1192);
and AND2 (N12159, N12117, N8608);
nor NOR4 (N12160, N12121, N3663, N11664, N2278);
xor XOR2 (N12161, N12159, N10378);
and AND2 (N12162, N12150, N7611);
buf BUF1 (N12163, N12158);
not NOT1 (N12164, N12154);
xor XOR2 (N12165, N12151, N2695);
nor NOR3 (N12166, N12132, N7705, N8136);
or OR2 (N12167, N12163, N611);
or OR3 (N12168, N12161, N1745, N9166);
and AND3 (N12169, N12149, N1748, N10987);
not NOT1 (N12170, N12165);
or OR2 (N12171, N12167, N2023);
and AND4 (N12172, N12169, N6183, N2643, N1261);
not NOT1 (N12173, N12171);
buf BUF1 (N12174, N12168);
buf BUF1 (N12175, N12162);
and AND2 (N12176, N12172, N10898);
buf BUF1 (N12177, N12164);
nand NAND4 (N12178, N12175, N6398, N7303, N9035);
and AND4 (N12179, N12173, N6168, N8042, N1803);
buf BUF1 (N12180, N12166);
not NOT1 (N12181, N12174);
nand NAND4 (N12182, N12148, N5152, N9862, N6099);
not NOT1 (N12183, N12176);
buf BUF1 (N12184, N12183);
and AND3 (N12185, N12184, N1510, N8146);
not NOT1 (N12186, N12170);
or OR2 (N12187, N12185, N10744);
buf BUF1 (N12188, N12178);
or OR4 (N12189, N12188, N3534, N9334, N4734);
nor NOR4 (N12190, N12182, N9628, N6962, N4495);
nor NOR3 (N12191, N12186, N2761, N7105);
nor NOR2 (N12192, N12160, N3908);
and AND3 (N12193, N12192, N6735, N7890);
nor NOR3 (N12194, N12191, N1543, N1762);
xor XOR2 (N12195, N12190, N8518);
nand NAND4 (N12196, N12189, N6587, N2560, N3328);
xor XOR2 (N12197, N12193, N10390);
nand NAND4 (N12198, N12187, N9774, N11621, N4401);
nand NAND4 (N12199, N12197, N3822, N1001, N9501);
or OR2 (N12200, N12195, N8503);
buf BUF1 (N12201, N12196);
or OR2 (N12202, N12200, N9321);
xor XOR2 (N12203, N12202, N1181);
nand NAND2 (N12204, N12203, N2909);
or OR4 (N12205, N12198, N1185, N3800, N11920);
not NOT1 (N12206, N12156);
not NOT1 (N12207, N12194);
nand NAND3 (N12208, N12180, N7332, N346);
nand NAND4 (N12209, N12177, N4624, N4506, N424);
not NOT1 (N12210, N12209);
and AND3 (N12211, N12199, N6583, N5588);
nor NOR4 (N12212, N12206, N11685, N1598, N2444);
buf BUF1 (N12213, N12210);
xor XOR2 (N12214, N12205, N11363);
buf BUF1 (N12215, N12213);
buf BUF1 (N12216, N12181);
xor XOR2 (N12217, N12214, N330);
nand NAND3 (N12218, N12179, N1979, N6613);
nand NAND3 (N12219, N12212, N9047, N5972);
not NOT1 (N12220, N12201);
nor NOR3 (N12221, N12220, N1899, N8898);
buf BUF1 (N12222, N12217);
xor XOR2 (N12223, N12211, N1015);
or OR4 (N12224, N12218, N11405, N5578, N6420);
or OR3 (N12225, N12221, N5709, N5174);
nor NOR3 (N12226, N12222, N939, N9864);
nor NOR2 (N12227, N12207, N6930);
nand NAND3 (N12228, N12215, N505, N709);
xor XOR2 (N12229, N12219, N2012);
not NOT1 (N12230, N12204);
xor XOR2 (N12231, N12223, N9523);
or OR2 (N12232, N12227, N9822);
not NOT1 (N12233, N12226);
xor XOR2 (N12234, N12228, N121);
not NOT1 (N12235, N12208);
or OR4 (N12236, N12231, N1837, N9104, N10566);
or OR2 (N12237, N12224, N2855);
nand NAND2 (N12238, N12232, N6369);
xor XOR2 (N12239, N12229, N9781);
nand NAND4 (N12240, N12230, N9503, N10694, N8774);
nand NAND4 (N12241, N12216, N3233, N1917, N9727);
buf BUF1 (N12242, N12239);
buf BUF1 (N12243, N12242);
nand NAND4 (N12244, N12225, N9391, N10196, N1873);
nor NOR2 (N12245, N12244, N2377);
nor NOR2 (N12246, N12238, N8536);
nand NAND2 (N12247, N12240, N47);
buf BUF1 (N12248, N12237);
and AND3 (N12249, N12247, N6986, N9891);
or OR2 (N12250, N12246, N1443);
nor NOR4 (N12251, N12245, N4291, N2841, N11032);
xor XOR2 (N12252, N12243, N10716);
not NOT1 (N12253, N12241);
buf BUF1 (N12254, N12251);
buf BUF1 (N12255, N12234);
not NOT1 (N12256, N12255);
not NOT1 (N12257, N12253);
xor XOR2 (N12258, N12233, N9002);
not NOT1 (N12259, N12258);
nor NOR2 (N12260, N12249, N12017);
xor XOR2 (N12261, N12236, N8616);
or OR3 (N12262, N12259, N7314, N11157);
or OR3 (N12263, N12235, N1325, N1052);
or OR3 (N12264, N12263, N11497, N2362);
and AND3 (N12265, N12262, N10194, N8893);
nor NOR4 (N12266, N12261, N8733, N5268, N5943);
nand NAND2 (N12267, N12252, N9694);
xor XOR2 (N12268, N12266, N5908);
buf BUF1 (N12269, N12248);
nand NAND3 (N12270, N12250, N6888, N4066);
buf BUF1 (N12271, N12268);
xor XOR2 (N12272, N12265, N12105);
not NOT1 (N12273, N12257);
xor XOR2 (N12274, N12272, N4760);
xor XOR2 (N12275, N12270, N381);
or OR2 (N12276, N12256, N9777);
nor NOR2 (N12277, N12264, N10251);
and AND2 (N12278, N12277, N8598);
not NOT1 (N12279, N12278);
nand NAND4 (N12280, N12274, N7675, N5768, N5326);
buf BUF1 (N12281, N12271);
not NOT1 (N12282, N12267);
and AND4 (N12283, N12282, N1608, N9588, N6255);
or OR3 (N12284, N12280, N6866, N8876);
nor NOR3 (N12285, N12279, N5741, N5650);
nor NOR4 (N12286, N12285, N10329, N5282, N7475);
or OR4 (N12287, N12286, N8933, N10911, N10933);
not NOT1 (N12288, N12254);
or OR3 (N12289, N12269, N720, N364);
nand NAND2 (N12290, N12273, N1541);
buf BUF1 (N12291, N12288);
xor XOR2 (N12292, N12290, N10889);
and AND4 (N12293, N12283, N3669, N9797, N1167);
not NOT1 (N12294, N12276);
nor NOR2 (N12295, N12292, N9797);
nand NAND3 (N12296, N12287, N336, N5885);
or OR4 (N12297, N12293, N878, N6048, N1163);
xor XOR2 (N12298, N12275, N3084);
not NOT1 (N12299, N12294);
nor NOR2 (N12300, N12291, N11092);
buf BUF1 (N12301, N12281);
or OR3 (N12302, N12298, N1311, N2009);
nand NAND4 (N12303, N12300, N3526, N7150, N11059);
not NOT1 (N12304, N12302);
or OR3 (N12305, N12299, N2274, N7426);
xor XOR2 (N12306, N12260, N4214);
not NOT1 (N12307, N12301);
or OR3 (N12308, N12297, N5750, N6673);
or OR4 (N12309, N12296, N9567, N1227, N7579);
xor XOR2 (N12310, N12284, N3226);
not NOT1 (N12311, N12304);
buf BUF1 (N12312, N12310);
nand NAND4 (N12313, N12309, N4071, N11213, N5768);
or OR2 (N12314, N12289, N4592);
xor XOR2 (N12315, N12307, N7773);
buf BUF1 (N12316, N12315);
nand NAND2 (N12317, N12295, N7053);
xor XOR2 (N12318, N12314, N5135);
or OR4 (N12319, N12317, N11377, N10927, N515);
nand NAND3 (N12320, N12308, N7920, N8164);
and AND2 (N12321, N12318, N8900);
buf BUF1 (N12322, N12306);
xor XOR2 (N12323, N12320, N9654);
not NOT1 (N12324, N12316);
buf BUF1 (N12325, N12311);
nand NAND3 (N12326, N12322, N10786, N650);
nor NOR4 (N12327, N12321, N10717, N1805, N10658);
nor NOR2 (N12328, N12326, N2970);
buf BUF1 (N12329, N12312);
or OR4 (N12330, N12323, N6303, N3599, N3410);
not NOT1 (N12331, N12319);
not NOT1 (N12332, N12331);
and AND3 (N12333, N12324, N7852, N3683);
nor NOR4 (N12334, N12313, N8599, N510, N12326);
not NOT1 (N12335, N12327);
nor NOR3 (N12336, N12329, N6435, N6680);
nand NAND3 (N12337, N12336, N2260, N6087);
nor NOR2 (N12338, N12305, N7034);
nor NOR4 (N12339, N12328, N10833, N7988, N7975);
buf BUF1 (N12340, N12335);
xor XOR2 (N12341, N12330, N7356);
or OR4 (N12342, N12338, N5580, N8782, N2767);
nor NOR4 (N12343, N12334, N10370, N4759, N11700);
nand NAND3 (N12344, N12332, N847, N10062);
not NOT1 (N12345, N12303);
nand NAND4 (N12346, N12341, N2835, N8277, N5817);
nor NOR2 (N12347, N12342, N8308);
or OR3 (N12348, N12333, N7413, N11740);
and AND4 (N12349, N12343, N8979, N3016, N11709);
not NOT1 (N12350, N12348);
nor NOR4 (N12351, N12337, N6502, N10259, N170);
not NOT1 (N12352, N12349);
or OR3 (N12353, N12325, N2142, N11259);
or OR3 (N12354, N12344, N9278, N5105);
not NOT1 (N12355, N12345);
and AND3 (N12356, N12351, N2502, N7962);
nand NAND3 (N12357, N12346, N6163, N10951);
not NOT1 (N12358, N12356);
nor NOR2 (N12359, N12352, N6390);
nand NAND3 (N12360, N12354, N5254, N3940);
buf BUF1 (N12361, N12357);
nor NOR4 (N12362, N12358, N5733, N1394, N1016);
and AND3 (N12363, N12339, N11947, N12129);
not NOT1 (N12364, N12340);
xor XOR2 (N12365, N12362, N10920);
nor NOR4 (N12366, N12347, N9886, N10141, N11061);
or OR4 (N12367, N12364, N10364, N982, N6126);
xor XOR2 (N12368, N12367, N7308);
not NOT1 (N12369, N12361);
nand NAND2 (N12370, N12368, N7168);
not NOT1 (N12371, N12366);
and AND3 (N12372, N12365, N1769, N4669);
nand NAND2 (N12373, N12355, N8141);
not NOT1 (N12374, N12363);
not NOT1 (N12375, N12370);
nand NAND3 (N12376, N12353, N4352, N3644);
and AND2 (N12377, N12376, N2349);
not NOT1 (N12378, N12375);
xor XOR2 (N12379, N12360, N1554);
nor NOR3 (N12380, N12359, N6758, N3525);
or OR3 (N12381, N12350, N12009, N3279);
xor XOR2 (N12382, N12371, N12099);
nand NAND4 (N12383, N12369, N3700, N7490, N7982);
not NOT1 (N12384, N12383);
and AND3 (N12385, N12379, N280, N11913);
nand NAND3 (N12386, N12373, N9501, N5293);
buf BUF1 (N12387, N12385);
and AND2 (N12388, N12378, N2629);
buf BUF1 (N12389, N12388);
buf BUF1 (N12390, N12387);
buf BUF1 (N12391, N12384);
or OR2 (N12392, N12382, N10968);
not NOT1 (N12393, N12380);
buf BUF1 (N12394, N12374);
or OR2 (N12395, N12393, N9756);
or OR3 (N12396, N12395, N5577, N6720);
not NOT1 (N12397, N12396);
xor XOR2 (N12398, N12390, N3596);
nor NOR2 (N12399, N12377, N9058);
not NOT1 (N12400, N12398);
buf BUF1 (N12401, N12391);
xor XOR2 (N12402, N12394, N1237);
nor NOR4 (N12403, N12399, N7723, N1768, N10651);
nor NOR2 (N12404, N12372, N5573);
and AND2 (N12405, N12401, N11643);
nor NOR2 (N12406, N12397, N1710);
xor XOR2 (N12407, N12402, N7515);
buf BUF1 (N12408, N12403);
not NOT1 (N12409, N12404);
xor XOR2 (N12410, N12392, N4878);
not NOT1 (N12411, N12406);
buf BUF1 (N12412, N12389);
nor NOR2 (N12413, N12408, N2707);
nor NOR2 (N12414, N12381, N1188);
xor XOR2 (N12415, N12413, N12015);
not NOT1 (N12416, N12414);
or OR2 (N12417, N12411, N4123);
or OR2 (N12418, N12405, N5526);
xor XOR2 (N12419, N12418, N7192);
not NOT1 (N12420, N12400);
not NOT1 (N12421, N12417);
xor XOR2 (N12422, N12415, N8681);
nor NOR3 (N12423, N12409, N659, N202);
and AND2 (N12424, N12422, N6871);
nor NOR4 (N12425, N12410, N2825, N7354, N5043);
not NOT1 (N12426, N12421);
not NOT1 (N12427, N12425);
buf BUF1 (N12428, N12386);
buf BUF1 (N12429, N12407);
nand NAND4 (N12430, N12419, N8478, N4903, N8215);
and AND3 (N12431, N12430, N5466, N6649);
not NOT1 (N12432, N12423);
not NOT1 (N12433, N12427);
nand NAND3 (N12434, N12424, N10956, N11406);
or OR2 (N12435, N12412, N11608);
nor NOR3 (N12436, N12429, N6177, N4623);
not NOT1 (N12437, N12426);
not NOT1 (N12438, N12416);
nor NOR3 (N12439, N12438, N9997, N3991);
buf BUF1 (N12440, N12431);
nand NAND2 (N12441, N12432, N7373);
xor XOR2 (N12442, N12433, N764);
or OR4 (N12443, N12437, N5974, N4297, N9316);
buf BUF1 (N12444, N12443);
buf BUF1 (N12445, N12444);
buf BUF1 (N12446, N12439);
or OR4 (N12447, N12446, N5391, N3113, N10482);
or OR2 (N12448, N12435, N951);
buf BUF1 (N12449, N12447);
not NOT1 (N12450, N12441);
buf BUF1 (N12451, N12442);
or OR3 (N12452, N12448, N7107, N4992);
and AND3 (N12453, N12434, N7149, N8563);
xor XOR2 (N12454, N12450, N2330);
and AND2 (N12455, N12436, N8457);
not NOT1 (N12456, N12452);
nand NAND4 (N12457, N12449, N12227, N11135, N11367);
nor NOR4 (N12458, N12440, N7340, N9549, N7597);
nor NOR2 (N12459, N12420, N6707);
xor XOR2 (N12460, N12458, N5480);
xor XOR2 (N12461, N12455, N10980);
not NOT1 (N12462, N12451);
and AND4 (N12463, N12460, N9727, N3121, N904);
nand NAND3 (N12464, N12445, N4665, N6500);
xor XOR2 (N12465, N12459, N3969);
nand NAND2 (N12466, N12464, N8509);
and AND3 (N12467, N12456, N6947, N11563);
nor NOR2 (N12468, N12428, N3217);
or OR3 (N12469, N12468, N9733, N9453);
nor NOR4 (N12470, N12457, N8124, N6002, N1087);
not NOT1 (N12471, N12462);
buf BUF1 (N12472, N12471);
not NOT1 (N12473, N12454);
or OR3 (N12474, N12470, N7230, N3426);
buf BUF1 (N12475, N12463);
or OR3 (N12476, N12465, N12433, N10362);
buf BUF1 (N12477, N12467);
or OR3 (N12478, N12461, N4840, N7913);
not NOT1 (N12479, N12478);
buf BUF1 (N12480, N12479);
buf BUF1 (N12481, N12477);
nor NOR2 (N12482, N12473, N7401);
buf BUF1 (N12483, N12472);
nand NAND3 (N12484, N12476, N9859, N4936);
xor XOR2 (N12485, N12475, N4901);
and AND4 (N12486, N12481, N2266, N3337, N2611);
nand NAND3 (N12487, N12469, N1443, N6075);
xor XOR2 (N12488, N12453, N5919);
nand NAND3 (N12489, N12488, N6008, N9914);
nor NOR2 (N12490, N12487, N5135);
buf BUF1 (N12491, N12489);
xor XOR2 (N12492, N12483, N5395);
xor XOR2 (N12493, N12492, N4244);
nor NOR3 (N12494, N12466, N1984, N10439);
not NOT1 (N12495, N12485);
and AND2 (N12496, N12484, N9606);
not NOT1 (N12497, N12486);
buf BUF1 (N12498, N12496);
not NOT1 (N12499, N12495);
not NOT1 (N12500, N12497);
or OR2 (N12501, N12490, N11261);
nor NOR3 (N12502, N12474, N5360, N4420);
and AND4 (N12503, N12494, N616, N5958, N8345);
not NOT1 (N12504, N12491);
nor NOR3 (N12505, N12504, N5584, N12155);
buf BUF1 (N12506, N12499);
or OR3 (N12507, N12503, N1832, N3834);
nand NAND3 (N12508, N12507, N11408, N4855);
buf BUF1 (N12509, N12500);
nand NAND2 (N12510, N12498, N5436);
nor NOR3 (N12511, N12482, N5291, N8647);
buf BUF1 (N12512, N12509);
or OR2 (N12513, N12502, N11086);
and AND2 (N12514, N12511, N11311);
or OR3 (N12515, N12510, N11417, N10559);
and AND4 (N12516, N12480, N6241, N1715, N9888);
not NOT1 (N12517, N12505);
or OR3 (N12518, N12513, N9290, N1434);
not NOT1 (N12519, N12515);
nand NAND3 (N12520, N12512, N10783, N10636);
or OR4 (N12521, N12501, N11702, N6786, N8795);
nand NAND2 (N12522, N12518, N10849);
or OR3 (N12523, N12506, N5648, N4181);
nand NAND3 (N12524, N12508, N2921, N2777);
and AND3 (N12525, N12520, N1419, N9431);
not NOT1 (N12526, N12522);
nand NAND4 (N12527, N12523, N10096, N4309, N10211);
nand NAND4 (N12528, N12526, N1513, N2245, N10683);
xor XOR2 (N12529, N12519, N4478);
and AND4 (N12530, N12517, N1400, N5638, N6776);
or OR3 (N12531, N12528, N9776, N9301);
nor NOR3 (N12532, N12531, N7275, N10862);
nor NOR4 (N12533, N12514, N6914, N5333, N10968);
and AND4 (N12534, N12532, N2768, N837, N5231);
buf BUF1 (N12535, N12516);
not NOT1 (N12536, N12535);
or OR3 (N12537, N12493, N2734, N7718);
not NOT1 (N12538, N12525);
or OR2 (N12539, N12536, N7463);
not NOT1 (N12540, N12538);
nand NAND3 (N12541, N12537, N4351, N5788);
and AND2 (N12542, N12534, N7974);
nor NOR3 (N12543, N12527, N3091, N11176);
or OR3 (N12544, N12540, N10828, N9606);
nor NOR3 (N12545, N12530, N8733, N2435);
nand NAND4 (N12546, N12541, N11559, N844, N5876);
xor XOR2 (N12547, N12529, N317);
nor NOR2 (N12548, N12539, N8914);
or OR4 (N12549, N12542, N3408, N2073, N2289);
not NOT1 (N12550, N12546);
or OR3 (N12551, N12550, N8153, N10241);
nand NAND4 (N12552, N12521, N8995, N12303, N5012);
buf BUF1 (N12553, N12543);
and AND4 (N12554, N12552, N9279, N10171, N5354);
or OR4 (N12555, N12549, N12255, N1856, N1030);
nor NOR4 (N12556, N12547, N11146, N6721, N11712);
xor XOR2 (N12557, N12553, N11315);
or OR3 (N12558, N12554, N7525, N661);
nand NAND3 (N12559, N12533, N10247, N10321);
not NOT1 (N12560, N12544);
and AND4 (N12561, N12548, N4624, N603, N920);
buf BUF1 (N12562, N12557);
nor NOR4 (N12563, N12545, N734, N11142, N2855);
nand NAND4 (N12564, N12559, N2811, N5681, N2872);
xor XOR2 (N12565, N12562, N11372);
and AND3 (N12566, N12564, N6837, N7474);
nand NAND4 (N12567, N12551, N2703, N6834, N5360);
nand NAND3 (N12568, N12556, N4860, N2606);
or OR2 (N12569, N12566, N8304);
and AND2 (N12570, N12563, N7969);
not NOT1 (N12571, N12560);
or OR4 (N12572, N12570, N10004, N12382, N5427);
and AND2 (N12573, N12565, N473);
xor XOR2 (N12574, N12569, N8948);
buf BUF1 (N12575, N12568);
xor XOR2 (N12576, N12567, N12068);
buf BUF1 (N12577, N12524);
not NOT1 (N12578, N12573);
nand NAND4 (N12579, N12571, N7399, N9583, N9807);
or OR4 (N12580, N12576, N595, N6119, N559);
nor NOR3 (N12581, N12555, N11249, N11621);
xor XOR2 (N12582, N12575, N9491);
not NOT1 (N12583, N12577);
not NOT1 (N12584, N12583);
not NOT1 (N12585, N12579);
or OR4 (N12586, N12572, N11583, N3950, N8396);
nand NAND2 (N12587, N12586, N10710);
xor XOR2 (N12588, N12580, N7833);
nor NOR3 (N12589, N12588, N8892, N5596);
and AND2 (N12590, N12574, N1194);
and AND4 (N12591, N12581, N10997, N1953, N8287);
and AND2 (N12592, N12578, N6811);
not NOT1 (N12593, N12558);
not NOT1 (N12594, N12584);
xor XOR2 (N12595, N12561, N8029);
xor XOR2 (N12596, N12592, N1266);
and AND2 (N12597, N12596, N3911);
and AND2 (N12598, N12594, N6215);
and AND3 (N12599, N12591, N6835, N8371);
buf BUF1 (N12600, N12593);
not NOT1 (N12601, N12587);
nor NOR3 (N12602, N12582, N10377, N8167);
not NOT1 (N12603, N12600);
or OR4 (N12604, N12597, N11133, N10509, N1093);
not NOT1 (N12605, N12604);
not NOT1 (N12606, N12585);
not NOT1 (N12607, N12606);
xor XOR2 (N12608, N12595, N9657);
or OR3 (N12609, N12603, N5589, N7286);
or OR4 (N12610, N12601, N2665, N3070, N11441);
nor NOR2 (N12611, N12608, N1813);
and AND3 (N12612, N12610, N4245, N12229);
not NOT1 (N12613, N12589);
and AND2 (N12614, N12605, N2950);
buf BUF1 (N12615, N12599);
not NOT1 (N12616, N12615);
nor NOR4 (N12617, N12613, N11560, N294, N3412);
nor NOR2 (N12618, N12609, N983);
not NOT1 (N12619, N12602);
not NOT1 (N12620, N12614);
and AND2 (N12621, N12618, N81);
not NOT1 (N12622, N12590);
nand NAND4 (N12623, N12598, N7959, N312, N6104);
or OR2 (N12624, N12616, N9555);
buf BUF1 (N12625, N12607);
xor XOR2 (N12626, N12619, N7647);
or OR3 (N12627, N12625, N10774, N11359);
buf BUF1 (N12628, N12612);
nor NOR4 (N12629, N12628, N9940, N7893, N12542);
nor NOR3 (N12630, N12611, N3018, N11709);
nand NAND2 (N12631, N12623, N6159);
nor NOR2 (N12632, N12617, N5342);
not NOT1 (N12633, N12622);
and AND4 (N12634, N12620, N7140, N4864, N12094);
nand NAND3 (N12635, N12633, N4, N11633);
buf BUF1 (N12636, N12627);
nand NAND4 (N12637, N12635, N6596, N9443, N5019);
not NOT1 (N12638, N12630);
xor XOR2 (N12639, N12631, N7518);
and AND3 (N12640, N12637, N10745, N7929);
nand NAND3 (N12641, N12621, N6382, N2905);
and AND4 (N12642, N12624, N6871, N4036, N1260);
xor XOR2 (N12643, N12626, N8051);
or OR4 (N12644, N12641, N9144, N9081, N986);
and AND4 (N12645, N12642, N2735, N7540, N6039);
nor NOR4 (N12646, N12632, N567, N8932, N4829);
not NOT1 (N12647, N12629);
nand NAND4 (N12648, N12643, N12403, N3111, N1922);
buf BUF1 (N12649, N12646);
nand NAND4 (N12650, N12638, N6787, N11656, N4331);
or OR4 (N12651, N12644, N433, N11196, N10539);
xor XOR2 (N12652, N12639, N3593);
buf BUF1 (N12653, N12645);
and AND2 (N12654, N12651, N3624);
not NOT1 (N12655, N12634);
nor NOR2 (N12656, N12636, N5819);
and AND4 (N12657, N12640, N8600, N4239, N5366);
and AND4 (N12658, N12650, N12344, N7666, N7579);
nand NAND4 (N12659, N12654, N5657, N12244, N6977);
xor XOR2 (N12660, N12658, N6015);
and AND3 (N12661, N12657, N2194, N3824);
and AND4 (N12662, N12655, N5460, N2433, N4948);
not NOT1 (N12663, N12659);
buf BUF1 (N12664, N12660);
not NOT1 (N12665, N12652);
nor NOR2 (N12666, N12649, N5743);
nand NAND2 (N12667, N12663, N3154);
nor NOR4 (N12668, N12656, N1311, N4804, N9703);
xor XOR2 (N12669, N12661, N5432);
and AND4 (N12670, N12668, N3929, N1604, N4840);
nor NOR4 (N12671, N12666, N5153, N1593, N11580);
nand NAND2 (N12672, N12667, N670);
xor XOR2 (N12673, N12669, N12107);
and AND2 (N12674, N12648, N1332);
not NOT1 (N12675, N12664);
buf BUF1 (N12676, N12647);
nor NOR2 (N12677, N12653, N8172);
nor NOR3 (N12678, N12673, N9209, N9202);
and AND2 (N12679, N12675, N7857);
nand NAND3 (N12680, N12676, N131, N2055);
and AND4 (N12681, N12677, N8582, N3312, N3239);
and AND3 (N12682, N12665, N6732, N12480);
or OR4 (N12683, N12670, N12085, N2054, N8294);
or OR3 (N12684, N12678, N10289, N11930);
and AND4 (N12685, N12680, N5920, N3665, N9999);
and AND2 (N12686, N12685, N10460);
nand NAND4 (N12687, N12674, N12231, N3719, N6931);
xor XOR2 (N12688, N12682, N4676);
not NOT1 (N12689, N12671);
not NOT1 (N12690, N12684);
not NOT1 (N12691, N12681);
and AND4 (N12692, N12679, N12173, N3773, N5551);
or OR3 (N12693, N12692, N10633, N3769);
and AND2 (N12694, N12686, N4599);
nand NAND4 (N12695, N12690, N5322, N12655, N6253);
buf BUF1 (N12696, N12693);
xor XOR2 (N12697, N12694, N6596);
buf BUF1 (N12698, N12689);
and AND3 (N12699, N12698, N4384, N2323);
nor NOR2 (N12700, N12696, N5891);
buf BUF1 (N12701, N12697);
or OR4 (N12702, N12691, N7733, N1461, N5892);
nand NAND2 (N12703, N12699, N12007);
buf BUF1 (N12704, N12687);
nor NOR4 (N12705, N12672, N961, N9404, N6950);
or OR4 (N12706, N12662, N12701, N4920, N8607);
or OR3 (N12707, N4808, N1667, N85);
xor XOR2 (N12708, N12706, N5657);
nand NAND4 (N12709, N12683, N829, N2736, N5680);
not NOT1 (N12710, N12700);
buf BUF1 (N12711, N12688);
or OR4 (N12712, N12705, N5536, N9077, N10079);
xor XOR2 (N12713, N12702, N9379);
not NOT1 (N12714, N12710);
nor NOR3 (N12715, N12712, N339, N7117);
and AND3 (N12716, N12715, N10066, N9164);
nand NAND2 (N12717, N12703, N7537);
and AND3 (N12718, N12704, N735, N10027);
nor NOR2 (N12719, N12718, N2178);
not NOT1 (N12720, N12711);
xor XOR2 (N12721, N12713, N2968);
or OR3 (N12722, N12719, N3391, N2365);
or OR4 (N12723, N12716, N10281, N592, N10999);
nand NAND3 (N12724, N12717, N8387, N1433);
or OR2 (N12725, N12714, N2533);
buf BUF1 (N12726, N12721);
nand NAND4 (N12727, N12707, N2124, N8921, N3060);
nand NAND3 (N12728, N12723, N10063, N786);
or OR2 (N12729, N12724, N8869);
or OR2 (N12730, N12728, N8473);
not NOT1 (N12731, N12725);
not NOT1 (N12732, N12730);
xor XOR2 (N12733, N12709, N3367);
nor NOR2 (N12734, N12695, N7440);
buf BUF1 (N12735, N12727);
or OR3 (N12736, N12731, N4555, N7720);
not NOT1 (N12737, N12735);
nor NOR4 (N12738, N12736, N2161, N2144, N7532);
xor XOR2 (N12739, N12732, N4299);
or OR2 (N12740, N12737, N5461);
nand NAND2 (N12741, N12726, N4459);
and AND4 (N12742, N12708, N12114, N1754, N2379);
or OR4 (N12743, N12740, N7906, N11889, N8745);
buf BUF1 (N12744, N12742);
or OR2 (N12745, N12722, N9191);
and AND2 (N12746, N12729, N7721);
buf BUF1 (N12747, N12733);
not NOT1 (N12748, N12734);
or OR2 (N12749, N12744, N7016);
nand NAND4 (N12750, N12741, N2489, N4895, N7733);
and AND3 (N12751, N12746, N9564, N9916);
or OR2 (N12752, N12743, N6533);
buf BUF1 (N12753, N12750);
and AND3 (N12754, N12752, N4486, N6376);
or OR3 (N12755, N12747, N8172, N1078);
not NOT1 (N12756, N12739);
buf BUF1 (N12757, N12756);
not NOT1 (N12758, N12748);
or OR2 (N12759, N12754, N5517);
nor NOR2 (N12760, N12720, N11795);
nand NAND3 (N12761, N12760, N9544, N3814);
not NOT1 (N12762, N12738);
or OR2 (N12763, N12758, N9050);
xor XOR2 (N12764, N12759, N4196);
or OR2 (N12765, N12763, N8798);
and AND4 (N12766, N12764, N2808, N7945, N962);
nor NOR4 (N12767, N12757, N11576, N1557, N11506);
or OR3 (N12768, N12762, N2776, N7278);
nor NOR4 (N12769, N12767, N2822, N9458, N11111);
or OR3 (N12770, N12766, N11342, N9843);
and AND3 (N12771, N12755, N8891, N11602);
or OR4 (N12772, N12751, N10935, N1532, N6047);
and AND4 (N12773, N12761, N3709, N7796, N3924);
xor XOR2 (N12774, N12745, N7859);
nand NAND4 (N12775, N12753, N7755, N690, N6818);
nor NOR3 (N12776, N12749, N5445, N9114);
xor XOR2 (N12777, N12771, N1704);
buf BUF1 (N12778, N12768);
and AND4 (N12779, N12770, N2351, N5723, N6395);
xor XOR2 (N12780, N12769, N1231);
nand NAND3 (N12781, N12780, N5461, N10202);
not NOT1 (N12782, N12779);
and AND4 (N12783, N12777, N8683, N11401, N11521);
buf BUF1 (N12784, N12772);
buf BUF1 (N12785, N12784);
and AND3 (N12786, N12776, N5142, N8125);
or OR2 (N12787, N12786, N10596);
buf BUF1 (N12788, N12783);
nor NOR4 (N12789, N12787, N11853, N7462, N523);
or OR2 (N12790, N12785, N7198);
xor XOR2 (N12791, N12778, N11687);
xor XOR2 (N12792, N12789, N954);
or OR3 (N12793, N12791, N5709, N5591);
buf BUF1 (N12794, N12765);
nand NAND4 (N12795, N12788, N9174, N181, N5573);
xor XOR2 (N12796, N12775, N444);
nand NAND2 (N12797, N12790, N9260);
nand NAND3 (N12798, N12795, N7864, N10924);
xor XOR2 (N12799, N12782, N3461);
and AND3 (N12800, N12794, N6709, N1619);
nor NOR4 (N12801, N12797, N983, N7491, N6464);
xor XOR2 (N12802, N12781, N9323);
or OR4 (N12803, N12800, N9008, N8778, N5373);
not NOT1 (N12804, N12796);
and AND3 (N12805, N12802, N5235, N12300);
or OR4 (N12806, N12804, N11471, N8410, N10644);
not NOT1 (N12807, N12805);
or OR4 (N12808, N12773, N12227, N6159, N7494);
buf BUF1 (N12809, N12793);
not NOT1 (N12810, N12803);
xor XOR2 (N12811, N12806, N2693);
or OR3 (N12812, N12811, N8379, N1181);
or OR3 (N12813, N12807, N3013, N11497);
nand NAND2 (N12814, N12809, N7619);
or OR4 (N12815, N12801, N11811, N9663, N11395);
nand NAND3 (N12816, N12808, N12433, N6379);
buf BUF1 (N12817, N12792);
buf BUF1 (N12818, N12815);
xor XOR2 (N12819, N12798, N4103);
or OR4 (N12820, N12817, N8974, N1012, N10971);
and AND4 (N12821, N12816, N8378, N8956, N9954);
nand NAND4 (N12822, N12814, N375, N7176, N1043);
buf BUF1 (N12823, N12799);
nor NOR4 (N12824, N12818, N4895, N1333, N538);
or OR2 (N12825, N12822, N5239);
or OR4 (N12826, N12774, N11707, N4767, N10568);
xor XOR2 (N12827, N12821, N9280);
not NOT1 (N12828, N12813);
or OR4 (N12829, N12823, N10108, N3109, N3703);
xor XOR2 (N12830, N12825, N3435);
buf BUF1 (N12831, N12824);
and AND3 (N12832, N12827, N12036, N12065);
not NOT1 (N12833, N12812);
and AND2 (N12834, N12819, N10905);
xor XOR2 (N12835, N12828, N5360);
nor NOR2 (N12836, N12810, N11983);
or OR2 (N12837, N12836, N1657);
nor NOR3 (N12838, N12820, N6203, N11677);
nand NAND2 (N12839, N12831, N374);
xor XOR2 (N12840, N12837, N12546);
nor NOR3 (N12841, N12832, N7733, N8222);
nor NOR3 (N12842, N12833, N8455, N6245);
buf BUF1 (N12843, N12835);
and AND4 (N12844, N12834, N5846, N3393, N7563);
xor XOR2 (N12845, N12842, N8727);
buf BUF1 (N12846, N12839);
not NOT1 (N12847, N12838);
not NOT1 (N12848, N12840);
and AND4 (N12849, N12847, N12352, N3343, N11537);
or OR4 (N12850, N12846, N12541, N11586, N10450);
xor XOR2 (N12851, N12830, N2034);
and AND4 (N12852, N12851, N1005, N10574, N2901);
not NOT1 (N12853, N12843);
not NOT1 (N12854, N12841);
buf BUF1 (N12855, N12845);
or OR2 (N12856, N12854, N10033);
xor XOR2 (N12857, N12849, N116);
or OR4 (N12858, N12844, N2213, N10224, N3568);
xor XOR2 (N12859, N12856, N8679);
not NOT1 (N12860, N12857);
nand NAND4 (N12861, N12855, N9791, N1608, N7162);
xor XOR2 (N12862, N12861, N3334);
or OR3 (N12863, N12848, N8166, N12002);
and AND2 (N12864, N12859, N9532);
nand NAND2 (N12865, N12858, N7775);
nor NOR4 (N12866, N12829, N12704, N8547, N10752);
or OR4 (N12867, N12866, N8657, N11110, N5658);
xor XOR2 (N12868, N12862, N4202);
nor NOR4 (N12869, N12867, N10132, N1573, N1777);
not NOT1 (N12870, N12850);
not NOT1 (N12871, N12853);
nor NOR4 (N12872, N12869, N361, N2055, N7868);
or OR3 (N12873, N12826, N12363, N12305);
or OR2 (N12874, N12872, N12484);
xor XOR2 (N12875, N12870, N1886);
not NOT1 (N12876, N12863);
not NOT1 (N12877, N12871);
nand NAND3 (N12878, N12876, N11024, N9890);
not NOT1 (N12879, N12852);
buf BUF1 (N12880, N12877);
and AND4 (N12881, N12880, N10268, N1022, N389);
and AND3 (N12882, N12878, N10548, N9938);
nand NAND3 (N12883, N12882, N11944, N7584);
or OR4 (N12884, N12875, N6997, N7319, N10902);
not NOT1 (N12885, N12881);
and AND4 (N12886, N12884, N7617, N5848, N7804);
xor XOR2 (N12887, N12885, N8658);
nor NOR2 (N12888, N12883, N6645);
nand NAND2 (N12889, N12886, N4252);
buf BUF1 (N12890, N12860);
xor XOR2 (N12891, N12874, N9758);
nand NAND2 (N12892, N12879, N868);
and AND3 (N12893, N12889, N950, N8769);
nand NAND2 (N12894, N12892, N9168);
xor XOR2 (N12895, N12868, N12535);
xor XOR2 (N12896, N12864, N1346);
xor XOR2 (N12897, N12896, N9671);
buf BUF1 (N12898, N12891);
not NOT1 (N12899, N12888);
and AND4 (N12900, N12895, N11783, N5460, N5700);
or OR2 (N12901, N12873, N12174);
not NOT1 (N12902, N12900);
and AND4 (N12903, N12901, N10001, N7765, N10292);
and AND2 (N12904, N12899, N5692);
or OR4 (N12905, N12893, N4564, N5129, N4064);
buf BUF1 (N12906, N12903);
and AND2 (N12907, N12897, N5154);
nor NOR4 (N12908, N12887, N5953, N2470, N4609);
not NOT1 (N12909, N12906);
nand NAND4 (N12910, N12908, N9585, N6374, N5258);
not NOT1 (N12911, N12894);
or OR4 (N12912, N12905, N4753, N7043, N2809);
xor XOR2 (N12913, N12911, N9473);
xor XOR2 (N12914, N12910, N10385);
xor XOR2 (N12915, N12913, N10137);
nand NAND3 (N12916, N12904, N3970, N2169);
xor XOR2 (N12917, N12890, N7409);
xor XOR2 (N12918, N12898, N2183);
nor NOR3 (N12919, N12907, N2611, N1256);
nor NOR2 (N12920, N12865, N2641);
or OR4 (N12921, N12916, N3809, N8689, N12716);
xor XOR2 (N12922, N12921, N6612);
buf BUF1 (N12923, N12920);
buf BUF1 (N12924, N12902);
or OR2 (N12925, N12914, N7378);
not NOT1 (N12926, N12919);
not NOT1 (N12927, N12917);
xor XOR2 (N12928, N12915, N9336);
or OR2 (N12929, N12924, N1555);
nand NAND2 (N12930, N12925, N1786);
nor NOR4 (N12931, N12930, N2931, N1282, N11229);
xor XOR2 (N12932, N12929, N4193);
xor XOR2 (N12933, N12918, N10669);
nor NOR4 (N12934, N12912, N9164, N11559, N4519);
nand NAND3 (N12935, N12909, N6179, N5552);
nor NOR2 (N12936, N12923, N325);
not NOT1 (N12937, N12932);
nor NOR3 (N12938, N12934, N8817, N738);
xor XOR2 (N12939, N12922, N8523);
or OR4 (N12940, N12928, N8754, N12007, N3165);
nand NAND4 (N12941, N12931, N10327, N11929, N10478);
or OR4 (N12942, N12941, N7732, N5766, N4436);
xor XOR2 (N12943, N12926, N5246);
not NOT1 (N12944, N12937);
buf BUF1 (N12945, N12927);
nor NOR4 (N12946, N12939, N104, N10961, N1709);
nand NAND3 (N12947, N12935, N7362, N4339);
buf BUF1 (N12948, N12936);
or OR3 (N12949, N12944, N5234, N11869);
not NOT1 (N12950, N12943);
xor XOR2 (N12951, N12948, N11840);
buf BUF1 (N12952, N12938);
buf BUF1 (N12953, N12949);
or OR3 (N12954, N12953, N12479, N7294);
nor NOR2 (N12955, N12952, N2879);
and AND4 (N12956, N12942, N12919, N10387, N6042);
xor XOR2 (N12957, N12945, N11708);
nor NOR4 (N12958, N12957, N10458, N9171, N6542);
nor NOR3 (N12959, N12951, N11437, N7331);
buf BUF1 (N12960, N12956);
not NOT1 (N12961, N12947);
or OR2 (N12962, N12950, N9183);
not NOT1 (N12963, N12961);
buf BUF1 (N12964, N12933);
not NOT1 (N12965, N12964);
not NOT1 (N12966, N12960);
or OR3 (N12967, N12962, N10900, N2353);
or OR4 (N12968, N12967, N7510, N3531, N12295);
nand NAND2 (N12969, N12966, N159);
buf BUF1 (N12970, N12955);
and AND3 (N12971, N12963, N4667, N7436);
nand NAND2 (N12972, N12940, N837);
xor XOR2 (N12973, N12969, N10414);
xor XOR2 (N12974, N12972, N4335);
nor NOR3 (N12975, N12968, N705, N5594);
buf BUF1 (N12976, N12974);
or OR2 (N12977, N12973, N1257);
buf BUF1 (N12978, N12971);
buf BUF1 (N12979, N12958);
buf BUF1 (N12980, N12959);
not NOT1 (N12981, N12979);
nand NAND4 (N12982, N12975, N2863, N11343, N6672);
and AND4 (N12983, N12976, N8750, N10551, N409);
nand NAND2 (N12984, N12954, N11093);
not NOT1 (N12985, N12981);
or OR4 (N12986, N12977, N2847, N3688, N944);
xor XOR2 (N12987, N12980, N966);
and AND3 (N12988, N12984, N3887, N560);
or OR3 (N12989, N12965, N877, N2049);
and AND4 (N12990, N12988, N4151, N3088, N3631);
and AND2 (N12991, N12986, N4854);
nor NOR3 (N12992, N12991, N56, N7353);
xor XOR2 (N12993, N12946, N12304);
nor NOR3 (N12994, N12982, N10707, N4154);
or OR4 (N12995, N12990, N1682, N4757, N5566);
nand NAND3 (N12996, N12985, N12430, N2907);
nand NAND3 (N12997, N12992, N7301, N4994);
and AND2 (N12998, N12989, N9254);
nor NOR4 (N12999, N12995, N4472, N480, N5454);
or OR4 (N13000, N12994, N7962, N2775, N3503);
not NOT1 (N13001, N13000);
not NOT1 (N13002, N12993);
nor NOR4 (N13003, N13002, N2057, N10795, N3842);
buf BUF1 (N13004, N12987);
not NOT1 (N13005, N12997);
or OR2 (N13006, N13005, N1272);
xor XOR2 (N13007, N12998, N12136);
and AND2 (N13008, N12983, N4141);
xor XOR2 (N13009, N12999, N4817);
nand NAND3 (N13010, N12978, N11972, N4615);
and AND3 (N13011, N13007, N10210, N4563);
nor NOR4 (N13012, N13001, N323, N410, N1724);
xor XOR2 (N13013, N12970, N12902);
or OR4 (N13014, N13008, N1498, N11346, N9626);
nor NOR4 (N13015, N13012, N4964, N8576, N1335);
xor XOR2 (N13016, N13010, N3222);
buf BUF1 (N13017, N13004);
buf BUF1 (N13018, N13014);
xor XOR2 (N13019, N13015, N4253);
and AND3 (N13020, N12996, N2690, N4582);
nor NOR4 (N13021, N13019, N11424, N3378, N11514);
or OR2 (N13022, N13009, N1012);
buf BUF1 (N13023, N13006);
and AND3 (N13024, N13011, N6857, N3268);
and AND2 (N13025, N13003, N12294);
nand NAND2 (N13026, N13022, N8332);
and AND2 (N13027, N13021, N7148);
nand NAND4 (N13028, N13017, N1647, N6746, N1020);
nor NOR2 (N13029, N13025, N7052);
not NOT1 (N13030, N13016);
nor NOR3 (N13031, N13028, N8428, N1204);
xor XOR2 (N13032, N13031, N7942);
nand NAND2 (N13033, N13026, N5346);
and AND2 (N13034, N13030, N9452);
nand NAND2 (N13035, N13023, N1942);
or OR2 (N13036, N13032, N392);
buf BUF1 (N13037, N13013);
xor XOR2 (N13038, N13018, N11573);
and AND2 (N13039, N13038, N11037);
buf BUF1 (N13040, N13033);
nor NOR4 (N13041, N13035, N4777, N12369, N12415);
buf BUF1 (N13042, N13027);
buf BUF1 (N13043, N13037);
or OR3 (N13044, N13040, N1849, N2262);
xor XOR2 (N13045, N13036, N1299);
nand NAND4 (N13046, N13042, N8505, N12294, N9729);
xor XOR2 (N13047, N13029, N6461);
not NOT1 (N13048, N13020);
nor NOR2 (N13049, N13044, N915);
or OR3 (N13050, N13043, N2652, N3245);
nor NOR2 (N13051, N13024, N7901);
xor XOR2 (N13052, N13049, N8249);
nor NOR3 (N13053, N13047, N8165, N3239);
nor NOR3 (N13054, N13052, N8735, N11210);
xor XOR2 (N13055, N13041, N6069);
nor NOR2 (N13056, N13050, N12973);
nor NOR2 (N13057, N13034, N10021);
nand NAND2 (N13058, N13048, N11382);
or OR3 (N13059, N13054, N9801, N13057);
nor NOR4 (N13060, N90, N7008, N5743, N10509);
or OR3 (N13061, N13039, N690, N6604);
xor XOR2 (N13062, N13051, N10416);
buf BUF1 (N13063, N13046);
nand NAND3 (N13064, N13060, N7270, N12298);
and AND4 (N13065, N13053, N6959, N11658, N10457);
nor NOR4 (N13066, N13061, N3846, N4312, N5725);
nor NOR3 (N13067, N13066, N4800, N464);
not NOT1 (N13068, N13058);
not NOT1 (N13069, N13059);
and AND2 (N13070, N13045, N3152);
nand NAND4 (N13071, N13055, N6346, N8374, N333);
xor XOR2 (N13072, N13070, N957);
buf BUF1 (N13073, N13065);
and AND3 (N13074, N13072, N4249, N4112);
or OR3 (N13075, N13073, N10749, N5291);
or OR3 (N13076, N13062, N260, N5941);
or OR4 (N13077, N13064, N5120, N1915, N8769);
nor NOR4 (N13078, N13069, N12410, N8065, N3299);
nand NAND2 (N13079, N13078, N9498);
xor XOR2 (N13080, N13067, N10647);
xor XOR2 (N13081, N13079, N3733);
or OR4 (N13082, N13081, N2363, N10050, N7130);
buf BUF1 (N13083, N13076);
and AND4 (N13084, N13068, N2694, N11755, N12424);
buf BUF1 (N13085, N13071);
buf BUF1 (N13086, N13075);
or OR3 (N13087, N13082, N11756, N7077);
xor XOR2 (N13088, N13087, N7462);
not NOT1 (N13089, N13056);
not NOT1 (N13090, N13063);
nor NOR4 (N13091, N13084, N11092, N12235, N11834);
not NOT1 (N13092, N13089);
not NOT1 (N13093, N13092);
buf BUF1 (N13094, N13088);
xor XOR2 (N13095, N13091, N4478);
nand NAND4 (N13096, N13077, N3883, N116, N5003);
nor NOR2 (N13097, N13096, N12547);
or OR2 (N13098, N13085, N11986);
buf BUF1 (N13099, N13097);
nor NOR3 (N13100, N13093, N2958, N11707);
or OR4 (N13101, N13095, N8879, N10694, N11454);
nor NOR3 (N13102, N13086, N9057, N4553);
or OR2 (N13103, N13102, N11773);
and AND3 (N13104, N13101, N3081, N8076);
xor XOR2 (N13105, N13104, N3146);
xor XOR2 (N13106, N13094, N4340);
and AND2 (N13107, N13098, N4813);
xor XOR2 (N13108, N13099, N633);
xor XOR2 (N13109, N13090, N4883);
nand NAND4 (N13110, N13107, N2883, N401, N3624);
not NOT1 (N13111, N13074);
or OR2 (N13112, N13109, N425);
xor XOR2 (N13113, N13103, N12857);
nor NOR2 (N13114, N13100, N11592);
and AND3 (N13115, N13114, N2225, N6546);
nand NAND4 (N13116, N13111, N3663, N6199, N3476);
xor XOR2 (N13117, N13113, N6382);
buf BUF1 (N13118, N13110);
xor XOR2 (N13119, N13116, N9255);
and AND3 (N13120, N13118, N10451, N7385);
and AND2 (N13121, N13083, N7986);
xor XOR2 (N13122, N13117, N4125);
not NOT1 (N13123, N13119);
and AND2 (N13124, N13105, N5672);
not NOT1 (N13125, N13123);
or OR4 (N13126, N13122, N4377, N4221, N5752);
not NOT1 (N13127, N13121);
buf BUF1 (N13128, N13080);
buf BUF1 (N13129, N13128);
nand NAND4 (N13130, N13127, N6847, N3787, N6870);
not NOT1 (N13131, N13120);
and AND4 (N13132, N13125, N12140, N10762, N5101);
buf BUF1 (N13133, N13106);
nor NOR2 (N13134, N13129, N12778);
nand NAND2 (N13135, N13130, N820);
and AND4 (N13136, N13135, N7090, N274, N9446);
nor NOR3 (N13137, N13108, N5126, N5264);
not NOT1 (N13138, N13136);
and AND3 (N13139, N13133, N10798, N800);
or OR3 (N13140, N13138, N3314, N9537);
nor NOR2 (N13141, N13115, N4892);
or OR4 (N13142, N13139, N13012, N11383, N6128);
or OR3 (N13143, N13112, N7208, N5413);
nor NOR2 (N13144, N13143, N8599);
nor NOR2 (N13145, N13142, N11678);
and AND3 (N13146, N13140, N4125, N10536);
nand NAND4 (N13147, N13134, N3109, N11267, N5228);
nand NAND3 (N13148, N13126, N2802, N9720);
and AND2 (N13149, N13146, N1874);
nand NAND2 (N13150, N13137, N9573);
buf BUF1 (N13151, N13149);
not NOT1 (N13152, N13144);
not NOT1 (N13153, N13141);
and AND4 (N13154, N13153, N5371, N8743, N7196);
not NOT1 (N13155, N13148);
xor XOR2 (N13156, N13132, N6792);
not NOT1 (N13157, N13156);
nor NOR4 (N13158, N13154, N487, N5812, N11541);
nand NAND2 (N13159, N13124, N461);
nor NOR3 (N13160, N13152, N2894, N11840);
and AND2 (N13161, N13159, N9282);
and AND4 (N13162, N13150, N8031, N6140, N6776);
nand NAND2 (N13163, N13162, N12318);
not NOT1 (N13164, N13155);
and AND4 (N13165, N13158, N10937, N8240, N5242);
and AND2 (N13166, N13163, N5447);
or OR2 (N13167, N13157, N257);
xor XOR2 (N13168, N13145, N1888);
nand NAND4 (N13169, N13147, N5551, N9752, N703);
nor NOR3 (N13170, N13165, N11799, N10502);
nand NAND3 (N13171, N13151, N1038, N2154);
and AND2 (N13172, N13167, N10886);
nand NAND2 (N13173, N13170, N4088);
and AND3 (N13174, N13169, N3653, N3362);
nand NAND3 (N13175, N13171, N2153, N4099);
buf BUF1 (N13176, N13160);
buf BUF1 (N13177, N13168);
or OR2 (N13178, N13174, N5284);
not NOT1 (N13179, N13161);
not NOT1 (N13180, N13177);
not NOT1 (N13181, N13175);
xor XOR2 (N13182, N13173, N174);
buf BUF1 (N13183, N13181);
and AND3 (N13184, N13164, N7628, N626);
nor NOR3 (N13185, N13131, N11529, N7030);
nand NAND2 (N13186, N13180, N6683);
nand NAND2 (N13187, N13172, N4352);
or OR4 (N13188, N13186, N327, N6767, N11150);
not NOT1 (N13189, N13187);
xor XOR2 (N13190, N13188, N6912);
nand NAND2 (N13191, N13185, N8449);
not NOT1 (N13192, N13166);
not NOT1 (N13193, N13179);
or OR2 (N13194, N13184, N7620);
or OR2 (N13195, N13190, N10046);
nor NOR4 (N13196, N13191, N7792, N11467, N7532);
nor NOR2 (N13197, N13183, N8239);
nand NAND2 (N13198, N13194, N2930);
or OR4 (N13199, N13189, N8545, N2166, N3506);
buf BUF1 (N13200, N13178);
nor NOR3 (N13201, N13199, N8736, N4638);
xor XOR2 (N13202, N13192, N11531);
or OR4 (N13203, N13176, N4138, N3258, N12680);
buf BUF1 (N13204, N13202);
nor NOR2 (N13205, N13198, N4602);
or OR3 (N13206, N13182, N6400, N6971);
not NOT1 (N13207, N13203);
or OR2 (N13208, N13207, N12747);
buf BUF1 (N13209, N13205);
xor XOR2 (N13210, N13196, N6899);
buf BUF1 (N13211, N13204);
nand NAND2 (N13212, N13209, N2906);
xor XOR2 (N13213, N13210, N1994);
xor XOR2 (N13214, N13193, N10676);
nand NAND3 (N13215, N13208, N2985, N4694);
not NOT1 (N13216, N13214);
nor NOR4 (N13217, N13211, N8783, N11321, N5239);
xor XOR2 (N13218, N13216, N5872);
nor NOR3 (N13219, N13212, N9916, N4398);
not NOT1 (N13220, N13218);
and AND3 (N13221, N13217, N12201, N11302);
xor XOR2 (N13222, N13201, N4511);
not NOT1 (N13223, N13195);
not NOT1 (N13224, N13206);
buf BUF1 (N13225, N13222);
nor NOR3 (N13226, N13223, N7691, N11741);
or OR2 (N13227, N13220, N1287);
nand NAND4 (N13228, N13225, N4871, N9409, N2827);
and AND3 (N13229, N13213, N12714, N5983);
nand NAND3 (N13230, N13215, N1793, N1265);
not NOT1 (N13231, N13227);
nor NOR4 (N13232, N13228, N2816, N10458, N8872);
xor XOR2 (N13233, N13224, N8842);
not NOT1 (N13234, N13233);
xor XOR2 (N13235, N13200, N12312);
xor XOR2 (N13236, N13234, N4752);
nor NOR3 (N13237, N13197, N5568, N11672);
nand NAND3 (N13238, N13221, N10152, N2397);
buf BUF1 (N13239, N13229);
nand NAND2 (N13240, N13235, N7156);
xor XOR2 (N13241, N13240, N10573);
buf BUF1 (N13242, N13239);
not NOT1 (N13243, N13232);
nor NOR3 (N13244, N13238, N238, N3670);
buf BUF1 (N13245, N13219);
xor XOR2 (N13246, N13241, N3060);
not NOT1 (N13247, N13237);
or OR2 (N13248, N13243, N11453);
or OR2 (N13249, N13226, N10142);
buf BUF1 (N13250, N13236);
nand NAND3 (N13251, N13250, N4487, N6293);
or OR4 (N13252, N13230, N9370, N12112, N11823);
xor XOR2 (N13253, N13245, N4935);
or OR2 (N13254, N13251, N4886);
xor XOR2 (N13255, N13246, N1378);
buf BUF1 (N13256, N13244);
or OR2 (N13257, N13247, N9478);
nand NAND3 (N13258, N13257, N4698, N2921);
not NOT1 (N13259, N13248);
and AND3 (N13260, N13231, N7385, N5081);
nand NAND3 (N13261, N13254, N3100, N5136);
not NOT1 (N13262, N13259);
or OR3 (N13263, N13261, N3416, N7527);
buf BUF1 (N13264, N13253);
or OR4 (N13265, N13242, N6695, N4916, N4550);
xor XOR2 (N13266, N13263, N6143);
nor NOR4 (N13267, N13266, N9859, N5498, N10082);
not NOT1 (N13268, N13267);
and AND3 (N13269, N13255, N8806, N8876);
buf BUF1 (N13270, N13262);
and AND2 (N13271, N13258, N5671);
nand NAND2 (N13272, N13269, N7946);
xor XOR2 (N13273, N13265, N6327);
and AND2 (N13274, N13249, N9797);
not NOT1 (N13275, N13252);
nor NOR3 (N13276, N13272, N5899, N4280);
buf BUF1 (N13277, N13260);
xor XOR2 (N13278, N13274, N2658);
nand NAND3 (N13279, N13273, N6730, N1208);
and AND3 (N13280, N13277, N708, N1888);
xor XOR2 (N13281, N13264, N10387);
or OR2 (N13282, N13280, N4760);
and AND3 (N13283, N13271, N10452, N7091);
nand NAND2 (N13284, N13268, N2398);
xor XOR2 (N13285, N13276, N11940);
nor NOR4 (N13286, N13284, N3674, N12283, N8143);
nand NAND4 (N13287, N13270, N12726, N10720, N9038);
nor NOR4 (N13288, N13287, N8343, N1767, N6443);
or OR4 (N13289, N13282, N1682, N12272, N10778);
or OR4 (N13290, N13275, N6714, N1047, N12915);
buf BUF1 (N13291, N13285);
nor NOR3 (N13292, N13281, N7397, N2510);
xor XOR2 (N13293, N13289, N12099);
and AND4 (N13294, N13279, N8648, N9788, N7696);
buf BUF1 (N13295, N13288);
nand NAND3 (N13296, N13292, N512, N9025);
buf BUF1 (N13297, N13256);
buf BUF1 (N13298, N13286);
buf BUF1 (N13299, N13296);
or OR4 (N13300, N13278, N2065, N12099, N9420);
xor XOR2 (N13301, N13298, N3020);
nand NAND2 (N13302, N13295, N2062);
or OR2 (N13303, N13291, N373);
xor XOR2 (N13304, N13303, N9978);
xor XOR2 (N13305, N13299, N2663);
nor NOR4 (N13306, N13304, N3414, N4763, N5476);
buf BUF1 (N13307, N13293);
and AND4 (N13308, N13283, N8003, N10772, N2408);
not NOT1 (N13309, N13290);
and AND4 (N13310, N13302, N12106, N12435, N12273);
buf BUF1 (N13311, N13310);
xor XOR2 (N13312, N13308, N7374);
buf BUF1 (N13313, N13309);
buf BUF1 (N13314, N13301);
and AND4 (N13315, N13297, N4858, N131, N10947);
not NOT1 (N13316, N13306);
or OR4 (N13317, N13314, N4231, N9291, N5689);
not NOT1 (N13318, N13307);
or OR4 (N13319, N13316, N2394, N1641, N6829);
or OR3 (N13320, N13318, N10550, N10315);
nor NOR4 (N13321, N13312, N4476, N6039, N3020);
and AND4 (N13322, N13317, N11445, N8745, N3320);
or OR4 (N13323, N13300, N1806, N1656, N1008);
nand NAND2 (N13324, N13320, N10667);
or OR4 (N13325, N13322, N7698, N5321, N3724);
and AND3 (N13326, N13311, N2364, N10786);
nand NAND2 (N13327, N13325, N9548);
or OR3 (N13328, N13324, N3297, N10653);
xor XOR2 (N13329, N13326, N3498);
nand NAND3 (N13330, N13319, N9000, N12060);
not NOT1 (N13331, N13327);
xor XOR2 (N13332, N13328, N709);
xor XOR2 (N13333, N13305, N12644);
nor NOR2 (N13334, N13333, N2478);
nor NOR4 (N13335, N13330, N10598, N1214, N994);
and AND3 (N13336, N13334, N11371, N9024);
not NOT1 (N13337, N13313);
nor NOR4 (N13338, N13323, N1969, N372, N8573);
nor NOR3 (N13339, N13315, N9915, N6349);
xor XOR2 (N13340, N13331, N8023);
and AND3 (N13341, N13339, N4026, N5748);
nand NAND4 (N13342, N13294, N605, N12979, N5046);
and AND4 (N13343, N13337, N9310, N6865, N7214);
not NOT1 (N13344, N13321);
and AND2 (N13345, N13340, N10570);
buf BUF1 (N13346, N13329);
not NOT1 (N13347, N13336);
nor NOR2 (N13348, N13346, N10088);
and AND3 (N13349, N13344, N10801, N1322);
xor XOR2 (N13350, N13338, N10876);
buf BUF1 (N13351, N13347);
not NOT1 (N13352, N13349);
buf BUF1 (N13353, N13335);
buf BUF1 (N13354, N13351);
and AND4 (N13355, N13332, N11747, N10002, N10464);
nor NOR2 (N13356, N13350, N7564);
nor NOR4 (N13357, N13356, N12185, N5016, N7502);
and AND3 (N13358, N13353, N4285, N437);
xor XOR2 (N13359, N13345, N9482);
nor NOR3 (N13360, N13359, N1127, N2499);
nand NAND3 (N13361, N13358, N5966, N6375);
xor XOR2 (N13362, N13357, N13100);
xor XOR2 (N13363, N13360, N741);
and AND4 (N13364, N13341, N2067, N6570, N10610);
buf BUF1 (N13365, N13361);
nand NAND4 (N13366, N13352, N7557, N2564, N9680);
or OR4 (N13367, N13348, N9139, N8751, N12888);
and AND3 (N13368, N13342, N8591, N216);
nor NOR4 (N13369, N13362, N2850, N5886, N11580);
nor NOR4 (N13370, N13354, N1270, N1787, N11314);
nor NOR2 (N13371, N13369, N1983);
and AND2 (N13372, N13364, N13367);
or OR2 (N13373, N5022, N2008);
nor NOR2 (N13374, N13370, N9804);
xor XOR2 (N13375, N13343, N12217);
nor NOR4 (N13376, N13368, N3296, N1061, N4413);
and AND2 (N13377, N13375, N51);
buf BUF1 (N13378, N13376);
not NOT1 (N13379, N13363);
nand NAND3 (N13380, N13366, N6646, N3470);
not NOT1 (N13381, N13355);
not NOT1 (N13382, N13365);
xor XOR2 (N13383, N13378, N5384);
or OR4 (N13384, N13377, N2476, N2301, N722);
buf BUF1 (N13385, N13381);
or OR4 (N13386, N13379, N7262, N8176, N122);
or OR4 (N13387, N13374, N3524, N5641, N12717);
buf BUF1 (N13388, N13371);
or OR4 (N13389, N13387, N9615, N9092, N4828);
xor XOR2 (N13390, N13386, N8369);
buf BUF1 (N13391, N13384);
buf BUF1 (N13392, N13372);
not NOT1 (N13393, N13383);
buf BUF1 (N13394, N13392);
or OR3 (N13395, N13385, N3504, N101);
nor NOR3 (N13396, N13380, N12751, N295);
and AND4 (N13397, N13395, N3798, N4300, N12074);
nor NOR3 (N13398, N13382, N4872, N6448);
or OR4 (N13399, N13397, N5749, N4054, N9516);
not NOT1 (N13400, N13391);
nor NOR2 (N13401, N13396, N10980);
and AND3 (N13402, N13388, N3311, N6118);
or OR4 (N13403, N13400, N13197, N3662, N5782);
xor XOR2 (N13404, N13403, N1079);
nor NOR2 (N13405, N13404, N7975);
and AND4 (N13406, N13401, N1465, N6900, N12175);
or OR4 (N13407, N13406, N7194, N11450, N1150);
nand NAND2 (N13408, N13393, N574);
buf BUF1 (N13409, N13373);
buf BUF1 (N13410, N13394);
buf BUF1 (N13411, N13409);
not NOT1 (N13412, N13405);
nor NOR4 (N13413, N13412, N1497, N10509, N11149);
nand NAND4 (N13414, N13398, N12850, N4746, N7790);
nor NOR4 (N13415, N13402, N3500, N12139, N7925);
nand NAND3 (N13416, N13413, N749, N2828);
buf BUF1 (N13417, N13390);
nand NAND2 (N13418, N13410, N6742);
nand NAND4 (N13419, N13418, N9194, N8016, N2705);
not NOT1 (N13420, N13417);
nor NOR4 (N13421, N13419, N6176, N10701, N2237);
nand NAND4 (N13422, N13399, N7772, N6030, N4833);
and AND4 (N13423, N13407, N6912, N5831, N10134);
xor XOR2 (N13424, N13389, N11623);
and AND4 (N13425, N13422, N9090, N10467, N8719);
or OR4 (N13426, N13425, N3579, N1657, N4415);
buf BUF1 (N13427, N13414);
buf BUF1 (N13428, N13421);
or OR4 (N13429, N13424, N8388, N331, N8621);
nor NOR3 (N13430, N13428, N2319, N7508);
nand NAND2 (N13431, N13415, N1344);
nand NAND3 (N13432, N13420, N6610, N1595);
not NOT1 (N13433, N13408);
and AND3 (N13434, N13427, N6249, N2948);
nor NOR2 (N13435, N13430, N9534);
nor NOR3 (N13436, N13432, N5824, N6299);
xor XOR2 (N13437, N13411, N10801);
buf BUF1 (N13438, N13434);
or OR4 (N13439, N13426, N3914, N597, N6521);
nand NAND2 (N13440, N13438, N8087);
xor XOR2 (N13441, N13423, N8616);
nor NOR4 (N13442, N13433, N11784, N7738, N6074);
nor NOR4 (N13443, N13439, N2425, N12839, N5885);
xor XOR2 (N13444, N13443, N2415);
buf BUF1 (N13445, N13436);
or OR4 (N13446, N13431, N57, N3914, N3549);
and AND3 (N13447, N13446, N1705, N13417);
xor XOR2 (N13448, N13435, N8878);
not NOT1 (N13449, N13447);
buf BUF1 (N13450, N13444);
nor NOR2 (N13451, N13449, N9186);
and AND2 (N13452, N13441, N10701);
xor XOR2 (N13453, N13440, N2253);
nand NAND3 (N13454, N13437, N7168, N7211);
nor NOR4 (N13455, N13429, N11761, N11723, N7017);
not NOT1 (N13456, N13454);
buf BUF1 (N13457, N13455);
buf BUF1 (N13458, N13450);
and AND4 (N13459, N13457, N12906, N10374, N9818);
or OR3 (N13460, N13452, N323, N8305);
xor XOR2 (N13461, N13456, N5512);
and AND4 (N13462, N13416, N12528, N3517, N5919);
xor XOR2 (N13463, N13448, N7977);
buf BUF1 (N13464, N13458);
nor NOR4 (N13465, N13464, N5211, N11824, N4227);
nor NOR3 (N13466, N13465, N3927, N2229);
or OR2 (N13467, N13453, N7820);
xor XOR2 (N13468, N13442, N11360);
nand NAND4 (N13469, N13463, N4450, N2205, N11285);
xor XOR2 (N13470, N13445, N8596);
and AND2 (N13471, N13470, N2633);
buf BUF1 (N13472, N13466);
and AND2 (N13473, N13461, N8398);
and AND2 (N13474, N13451, N3985);
xor XOR2 (N13475, N13459, N9286);
buf BUF1 (N13476, N13475);
xor XOR2 (N13477, N13471, N3220);
nor NOR4 (N13478, N13469, N3255, N7212, N8881);
buf BUF1 (N13479, N13462);
and AND2 (N13480, N13472, N179);
not NOT1 (N13481, N13479);
nand NAND4 (N13482, N13477, N13200, N13231, N6968);
or OR3 (N13483, N13460, N3720, N11151);
not NOT1 (N13484, N13476);
or OR3 (N13485, N13478, N5740, N5083);
not NOT1 (N13486, N13485);
xor XOR2 (N13487, N13483, N9589);
buf BUF1 (N13488, N13474);
not NOT1 (N13489, N13487);
or OR2 (N13490, N13486, N3766);
xor XOR2 (N13491, N13473, N10757);
nand NAND3 (N13492, N13489, N12266, N13378);
buf BUF1 (N13493, N13482);
not NOT1 (N13494, N13492);
and AND3 (N13495, N13488, N12520, N7747);
not NOT1 (N13496, N13467);
buf BUF1 (N13497, N13480);
or OR2 (N13498, N13496, N8796);
xor XOR2 (N13499, N13491, N7868);
buf BUF1 (N13500, N13495);
not NOT1 (N13501, N13481);
and AND4 (N13502, N13490, N9679, N11162, N3634);
nand NAND3 (N13503, N13497, N10885, N2965);
buf BUF1 (N13504, N13493);
nand NAND2 (N13505, N13503, N2806);
not NOT1 (N13506, N13500);
or OR3 (N13507, N13501, N6136, N10611);
buf BUF1 (N13508, N13499);
buf BUF1 (N13509, N13468);
xor XOR2 (N13510, N13508, N7936);
nor NOR3 (N13511, N13502, N9922, N11305);
xor XOR2 (N13512, N13510, N11252);
nand NAND2 (N13513, N13509, N10878);
buf BUF1 (N13514, N13513);
nor NOR2 (N13515, N13505, N10434);
nor NOR3 (N13516, N13484, N12502, N582);
nand NAND2 (N13517, N13506, N10070);
or OR3 (N13518, N13512, N13152, N10966);
and AND4 (N13519, N13511, N13506, N9515, N6855);
nor NOR3 (N13520, N13494, N9550, N3879);
not NOT1 (N13521, N13498);
nor NOR4 (N13522, N13514, N10763, N4421, N11715);
and AND3 (N13523, N13517, N7649, N10134);
or OR4 (N13524, N13518, N3707, N3335, N6467);
not NOT1 (N13525, N13516);
and AND3 (N13526, N13519, N6660, N5436);
xor XOR2 (N13527, N13521, N4383);
not NOT1 (N13528, N13504);
not NOT1 (N13529, N13527);
buf BUF1 (N13530, N13515);
xor XOR2 (N13531, N13522, N1900);
or OR3 (N13532, N13525, N5939, N8424);
nand NAND2 (N13533, N13530, N11222);
not NOT1 (N13534, N13523);
nor NOR4 (N13535, N13529, N9515, N6639, N8650);
and AND2 (N13536, N13520, N1586);
and AND3 (N13537, N13528, N12167, N1639);
not NOT1 (N13538, N13535);
nor NOR3 (N13539, N13507, N6273, N11328);
nand NAND2 (N13540, N13531, N10633);
xor XOR2 (N13541, N13533, N1785);
nand NAND3 (N13542, N13537, N10310, N12807);
not NOT1 (N13543, N13536);
and AND4 (N13544, N13526, N3710, N7617, N3328);
xor XOR2 (N13545, N13538, N12754);
xor XOR2 (N13546, N13524, N2016);
not NOT1 (N13547, N13546);
nor NOR4 (N13548, N13541, N7679, N4529, N10281);
nand NAND2 (N13549, N13545, N3548);
nand NAND3 (N13550, N13547, N1518, N2628);
and AND2 (N13551, N13540, N8145);
nand NAND3 (N13552, N13542, N13483, N8032);
not NOT1 (N13553, N13550);
nor NOR4 (N13554, N13553, N1285, N1440, N10445);
and AND2 (N13555, N13544, N2368);
not NOT1 (N13556, N13539);
buf BUF1 (N13557, N13552);
and AND4 (N13558, N13557, N13335, N8723, N4348);
buf BUF1 (N13559, N13558);
nand NAND3 (N13560, N13534, N4933, N2142);
and AND3 (N13561, N13559, N3302, N3780);
or OR2 (N13562, N13561, N6623);
buf BUF1 (N13563, N13532);
or OR3 (N13564, N13560, N5172, N7895);
and AND3 (N13565, N13549, N3668, N12839);
nor NOR4 (N13566, N13565, N6420, N642, N6121);
or OR4 (N13567, N13551, N5760, N1675, N7245);
buf BUF1 (N13568, N13564);
or OR2 (N13569, N13548, N12312);
nand NAND3 (N13570, N13566, N6510, N2950);
nand NAND2 (N13571, N13562, N4704);
nor NOR2 (N13572, N13543, N10957);
and AND4 (N13573, N13563, N9297, N2224, N532);
and AND3 (N13574, N13570, N9456, N5471);
xor XOR2 (N13575, N13556, N3954);
xor XOR2 (N13576, N13554, N3526);
nor NOR2 (N13577, N13572, N8914);
not NOT1 (N13578, N13573);
nand NAND3 (N13579, N13575, N12830, N8675);
nand NAND3 (N13580, N13579, N8859, N12902);
and AND2 (N13581, N13555, N12630);
nor NOR2 (N13582, N13578, N2301);
or OR3 (N13583, N13581, N2365, N10486);
not NOT1 (N13584, N13580);
and AND4 (N13585, N13584, N1852, N5461, N7313);
buf BUF1 (N13586, N13582);
or OR3 (N13587, N13568, N2846, N4657);
nor NOR2 (N13588, N13583, N8021);
nand NAND2 (N13589, N13576, N11721);
nor NOR2 (N13590, N13588, N12960);
not NOT1 (N13591, N13585);
and AND4 (N13592, N13586, N1270, N12980, N7592);
buf BUF1 (N13593, N13590);
buf BUF1 (N13594, N13574);
nor NOR2 (N13595, N13589, N4666);
nand NAND2 (N13596, N13591, N4853);
and AND4 (N13597, N13571, N3256, N2927, N8304);
buf BUF1 (N13598, N13569);
or OR2 (N13599, N13598, N1723);
not NOT1 (N13600, N13592);
buf BUF1 (N13601, N13594);
xor XOR2 (N13602, N13587, N12353);
not NOT1 (N13603, N13595);
buf BUF1 (N13604, N13603);
and AND2 (N13605, N13601, N1243);
not NOT1 (N13606, N13593);
or OR4 (N13607, N13597, N2061, N10245, N12892);
xor XOR2 (N13608, N13596, N10746);
nor NOR4 (N13609, N13567, N11658, N7071, N5787);
buf BUF1 (N13610, N13607);
nor NOR4 (N13611, N13605, N9930, N1112, N11060);
buf BUF1 (N13612, N13577);
not NOT1 (N13613, N13608);
and AND4 (N13614, N13599, N11818, N4327, N10078);
and AND3 (N13615, N13610, N7606, N10056);
buf BUF1 (N13616, N13602);
nor NOR2 (N13617, N13604, N1745);
buf BUF1 (N13618, N13616);
nor NOR2 (N13619, N13611, N3619);
nand NAND4 (N13620, N13613, N3678, N13529, N4514);
buf BUF1 (N13621, N13614);
nor NOR4 (N13622, N13600, N2098, N1882, N13266);
not NOT1 (N13623, N13609);
or OR4 (N13624, N13620, N6955, N12460, N8784);
not NOT1 (N13625, N13621);
not NOT1 (N13626, N13617);
and AND3 (N13627, N13624, N7460, N5517);
xor XOR2 (N13628, N13606, N4304);
nor NOR2 (N13629, N13623, N8966);
and AND4 (N13630, N13626, N8036, N10274, N6398);
buf BUF1 (N13631, N13612);
not NOT1 (N13632, N13629);
not NOT1 (N13633, N13615);
and AND3 (N13634, N13628, N9432, N11495);
not NOT1 (N13635, N13622);
buf BUF1 (N13636, N13633);
and AND2 (N13637, N13634, N12382);
nor NOR3 (N13638, N13618, N4818, N2608);
buf BUF1 (N13639, N13638);
not NOT1 (N13640, N13625);
nor NOR4 (N13641, N13637, N6859, N7009, N2602);
xor XOR2 (N13642, N13639, N1377);
nor NOR2 (N13643, N13631, N4531);
and AND3 (N13644, N13641, N11733, N6292);
nor NOR4 (N13645, N13636, N8342, N8904, N9675);
and AND2 (N13646, N13642, N1535);
or OR4 (N13647, N13645, N4729, N7681, N6703);
buf BUF1 (N13648, N13630);
xor XOR2 (N13649, N13644, N2507);
or OR4 (N13650, N13632, N8098, N6274, N7013);
and AND3 (N13651, N13643, N13273, N3341);
nand NAND4 (N13652, N13635, N2468, N949, N3819);
not NOT1 (N13653, N13640);
buf BUF1 (N13654, N13653);
xor XOR2 (N13655, N13619, N3556);
or OR4 (N13656, N13649, N1042, N11231, N3621);
not NOT1 (N13657, N13652);
or OR4 (N13658, N13647, N6250, N7759, N8828);
not NOT1 (N13659, N13651);
and AND4 (N13660, N13656, N10199, N4917, N3809);
and AND3 (N13661, N13659, N4354, N10121);
not NOT1 (N13662, N13658);
nand NAND3 (N13663, N13662, N4460, N11366);
and AND2 (N13664, N13654, N7028);
buf BUF1 (N13665, N13657);
or OR3 (N13666, N13663, N9591, N11921);
not NOT1 (N13667, N13665);
nor NOR4 (N13668, N13661, N7047, N1664, N6909);
nor NOR4 (N13669, N13666, N8416, N12470, N2163);
and AND4 (N13670, N13664, N10029, N240, N11178);
nand NAND3 (N13671, N13668, N2455, N13126);
xor XOR2 (N13672, N13660, N1593);
not NOT1 (N13673, N13650);
or OR4 (N13674, N13673, N1965, N4207, N11708);
or OR4 (N13675, N13667, N4146, N11054, N9702);
nor NOR4 (N13676, N13669, N6407, N11238, N2562);
or OR2 (N13677, N13671, N3179);
buf BUF1 (N13678, N13655);
xor XOR2 (N13679, N13672, N1008);
not NOT1 (N13680, N13646);
and AND4 (N13681, N13627, N4751, N3092, N9823);
buf BUF1 (N13682, N13680);
and AND3 (N13683, N13675, N2481, N12807);
buf BUF1 (N13684, N13677);
xor XOR2 (N13685, N13648, N7343);
nor NOR2 (N13686, N13670, N3712);
buf BUF1 (N13687, N13679);
nor NOR4 (N13688, N13676, N3647, N11516, N681);
xor XOR2 (N13689, N13688, N11757);
and AND4 (N13690, N13674, N11214, N1308, N9297);
nand NAND3 (N13691, N13687, N11403, N6417);
buf BUF1 (N13692, N13691);
and AND4 (N13693, N13686, N11989, N3076, N6854);
or OR2 (N13694, N13690, N1519);
xor XOR2 (N13695, N13678, N10526);
not NOT1 (N13696, N13681);
and AND3 (N13697, N13682, N3372, N4248);
nand NAND2 (N13698, N13697, N9576);
or OR3 (N13699, N13683, N11656, N5306);
not NOT1 (N13700, N13695);
nor NOR3 (N13701, N13696, N5957, N2586);
and AND3 (N13702, N13684, N8538, N9107);
not NOT1 (N13703, N13698);
nor NOR4 (N13704, N13692, N12629, N10644, N10916);
xor XOR2 (N13705, N13704, N9483);
or OR3 (N13706, N13705, N10337, N5848);
or OR2 (N13707, N13701, N7712);
not NOT1 (N13708, N13699);
or OR2 (N13709, N13707, N1913);
nand NAND3 (N13710, N13702, N17, N10174);
or OR2 (N13711, N13693, N2735);
nor NOR2 (N13712, N13700, N4512);
nand NAND3 (N13713, N13685, N12893, N3297);
xor XOR2 (N13714, N13706, N3142);
nor NOR4 (N13715, N13689, N278, N5627, N219);
nor NOR4 (N13716, N13709, N2426, N5889, N8740);
xor XOR2 (N13717, N13694, N3513);
xor XOR2 (N13718, N13716, N3072);
and AND4 (N13719, N13714, N416, N4931, N3950);
buf BUF1 (N13720, N13711);
nand NAND2 (N13721, N13712, N2744);
or OR4 (N13722, N13719, N10095, N1693, N11781);
xor XOR2 (N13723, N13721, N10109);
xor XOR2 (N13724, N13715, N9954);
nand NAND4 (N13725, N13717, N2313, N12935, N4694);
and AND3 (N13726, N13723, N443, N1006);
and AND2 (N13727, N13724, N639);
and AND4 (N13728, N13725, N7850, N2435, N10105);
nor NOR2 (N13729, N13727, N3634);
not NOT1 (N13730, N13729);
nor NOR4 (N13731, N13718, N1325, N6635, N1879);
buf BUF1 (N13732, N13730);
and AND3 (N13733, N13720, N6451, N1478);
and AND2 (N13734, N13703, N7490);
and AND4 (N13735, N13733, N751, N8387, N10757);
not NOT1 (N13736, N13726);
not NOT1 (N13737, N13736);
or OR4 (N13738, N13722, N1998, N3272, N4318);
or OR2 (N13739, N13738, N11600);
or OR3 (N13740, N13732, N13682, N1433);
nor NOR4 (N13741, N13737, N8339, N940, N5147);
buf BUF1 (N13742, N13739);
buf BUF1 (N13743, N13742);
or OR2 (N13744, N13731, N5635);
xor XOR2 (N13745, N13741, N12950);
nand NAND2 (N13746, N13710, N7580);
not NOT1 (N13747, N13744);
nor NOR2 (N13748, N13735, N6923);
nor NOR2 (N13749, N13745, N3377);
or OR2 (N13750, N13713, N4049);
buf BUF1 (N13751, N13750);
xor XOR2 (N13752, N13743, N9937);
nor NOR4 (N13753, N13751, N58, N12348, N6516);
and AND3 (N13754, N13747, N13360, N5283);
xor XOR2 (N13755, N13749, N3254);
nor NOR2 (N13756, N13708, N2418);
or OR2 (N13757, N13752, N5591);
xor XOR2 (N13758, N13728, N8742);
and AND3 (N13759, N13756, N3112, N12410);
nor NOR4 (N13760, N13755, N4758, N11092, N7756);
buf BUF1 (N13761, N13760);
and AND2 (N13762, N13759, N242);
and AND2 (N13763, N13761, N6489);
xor XOR2 (N13764, N13754, N13760);
or OR3 (N13765, N13753, N5155, N1333);
not NOT1 (N13766, N13762);
not NOT1 (N13767, N13758);
buf BUF1 (N13768, N13734);
buf BUF1 (N13769, N13740);
and AND2 (N13770, N13768, N6134);
xor XOR2 (N13771, N13748, N12252);
or OR4 (N13772, N13746, N4576, N1444, N11082);
nand NAND3 (N13773, N13770, N12773, N8958);
buf BUF1 (N13774, N13771);
and AND3 (N13775, N13764, N7283, N7153);
or OR2 (N13776, N13775, N8585);
not NOT1 (N13777, N13776);
nor NOR4 (N13778, N13757, N7234, N1696, N12664);
and AND2 (N13779, N13769, N5942);
nand NAND4 (N13780, N13763, N12213, N12293, N4959);
not NOT1 (N13781, N13777);
nand NAND2 (N13782, N13774, N7197);
and AND3 (N13783, N13780, N5629, N12246);
nor NOR2 (N13784, N13767, N9378);
buf BUF1 (N13785, N13782);
nor NOR3 (N13786, N13766, N2225, N10613);
xor XOR2 (N13787, N13785, N4132);
buf BUF1 (N13788, N13765);
or OR2 (N13789, N13788, N11299);
or OR4 (N13790, N13779, N6700, N7989, N13586);
or OR4 (N13791, N13787, N359, N5465, N557);
xor XOR2 (N13792, N13789, N10856);
nor NOR3 (N13793, N13773, N9117, N5004);
nor NOR4 (N13794, N13783, N4424, N3310, N2863);
nand NAND4 (N13795, N13784, N3066, N9995, N7111);
nor NOR2 (N13796, N13791, N9563);
nor NOR2 (N13797, N13790, N6526);
xor XOR2 (N13798, N13795, N12100);
xor XOR2 (N13799, N13796, N1795);
nand NAND3 (N13800, N13793, N12977, N4241);
xor XOR2 (N13801, N13798, N6057);
nand NAND3 (N13802, N13778, N2220, N8536);
not NOT1 (N13803, N13781);
not NOT1 (N13804, N13772);
xor XOR2 (N13805, N13800, N6614);
nor NOR2 (N13806, N13801, N3255);
buf BUF1 (N13807, N13806);
nor NOR4 (N13808, N13807, N4887, N285, N2952);
buf BUF1 (N13809, N13799);
buf BUF1 (N13810, N13808);
nand NAND3 (N13811, N13803, N11821, N13737);
nand NAND2 (N13812, N13794, N1571);
nor NOR3 (N13813, N13811, N12265, N7608);
nor NOR3 (N13814, N13812, N864, N9500);
nand NAND4 (N13815, N13814, N11736, N7669, N4509);
not NOT1 (N13816, N13805);
nor NOR2 (N13817, N13802, N1287);
nand NAND2 (N13818, N13810, N6599);
xor XOR2 (N13819, N13809, N7260);
nand NAND4 (N13820, N13797, N6787, N9547, N7416);
buf BUF1 (N13821, N13819);
xor XOR2 (N13822, N13818, N1091);
buf BUF1 (N13823, N13816);
xor XOR2 (N13824, N13817, N66);
or OR3 (N13825, N13815, N8841, N888);
and AND3 (N13826, N13823, N7899, N3454);
buf BUF1 (N13827, N13821);
not NOT1 (N13828, N13786);
nor NOR2 (N13829, N13827, N2367);
and AND3 (N13830, N13822, N6421, N3448);
xor XOR2 (N13831, N13804, N9533);
buf BUF1 (N13832, N13829);
xor XOR2 (N13833, N13813, N4268);
xor XOR2 (N13834, N13826, N3603);
and AND3 (N13835, N13825, N13000, N1403);
nor NOR4 (N13836, N13834, N13791, N272, N8294);
nand NAND4 (N13837, N13820, N3015, N2964, N9028);
nand NAND3 (N13838, N13830, N12494, N1585);
nor NOR4 (N13839, N13828, N6092, N5009, N4242);
not NOT1 (N13840, N13831);
nor NOR4 (N13841, N13833, N2817, N11974, N10375);
nand NAND4 (N13842, N13824, N5243, N5461, N4695);
buf BUF1 (N13843, N13842);
and AND3 (N13844, N13838, N12120, N2538);
nor NOR2 (N13845, N13839, N3597);
nor NOR2 (N13846, N13792, N3508);
or OR4 (N13847, N13837, N1129, N4356, N13773);
buf BUF1 (N13848, N13836);
nand NAND3 (N13849, N13847, N6495, N9556);
and AND3 (N13850, N13840, N11653, N5701);
nand NAND2 (N13851, N13841, N12785);
or OR3 (N13852, N13843, N3851, N198);
and AND2 (N13853, N13832, N13294);
or OR2 (N13854, N13851, N8319);
and AND4 (N13855, N13850, N1410, N7507, N5493);
nand NAND3 (N13856, N13854, N1723, N2244);
buf BUF1 (N13857, N13844);
xor XOR2 (N13858, N13849, N7860);
or OR2 (N13859, N13856, N2639);
nand NAND2 (N13860, N13858, N9812);
buf BUF1 (N13861, N13848);
or OR4 (N13862, N13852, N4441, N4230, N5734);
or OR2 (N13863, N13857, N120);
xor XOR2 (N13864, N13862, N5790);
buf BUF1 (N13865, N13864);
nand NAND2 (N13866, N13859, N4326);
buf BUF1 (N13867, N13865);
not NOT1 (N13868, N13860);
nor NOR2 (N13869, N13845, N9353);
buf BUF1 (N13870, N13868);
or OR4 (N13871, N13855, N2607, N404, N13828);
and AND3 (N13872, N13867, N506, N1371);
or OR3 (N13873, N13870, N11855, N6342);
nor NOR3 (N13874, N13871, N724, N12109);
buf BUF1 (N13875, N13866);
not NOT1 (N13876, N13835);
nor NOR2 (N13877, N13875, N12442);
and AND2 (N13878, N13876, N5305);
or OR3 (N13879, N13878, N176, N10899);
not NOT1 (N13880, N13863);
nand NAND2 (N13881, N13877, N2303);
and AND4 (N13882, N13861, N2363, N3045, N5709);
not NOT1 (N13883, N13869);
nand NAND4 (N13884, N13873, N9301, N1664, N4073);
and AND2 (N13885, N13880, N5081);
not NOT1 (N13886, N13879);
not NOT1 (N13887, N13884);
buf BUF1 (N13888, N13881);
xor XOR2 (N13889, N13853, N6849);
xor XOR2 (N13890, N13882, N1409);
xor XOR2 (N13891, N13883, N8476);
xor XOR2 (N13892, N13888, N5213);
not NOT1 (N13893, N13889);
or OR3 (N13894, N13872, N3738, N6408);
buf BUF1 (N13895, N13890);
not NOT1 (N13896, N13846);
not NOT1 (N13897, N13891);
not NOT1 (N13898, N13874);
nor NOR3 (N13899, N13885, N5573, N11303);
or OR4 (N13900, N13895, N11274, N9186, N7355);
not NOT1 (N13901, N13892);
nor NOR3 (N13902, N13886, N3435, N6919);
or OR2 (N13903, N13887, N10472);
and AND4 (N13904, N13894, N3692, N4151, N9474);
not NOT1 (N13905, N13904);
xor XOR2 (N13906, N13896, N13796);
xor XOR2 (N13907, N13899, N10082);
xor XOR2 (N13908, N13900, N11803);
nand NAND4 (N13909, N13903, N11648, N9508, N1537);
and AND2 (N13910, N13893, N2744);
or OR4 (N13911, N13902, N8757, N8549, N10459);
nor NOR3 (N13912, N13898, N13689, N10219);
nand NAND2 (N13913, N13909, N13540);
and AND4 (N13914, N13905, N12615, N9525, N13627);
not NOT1 (N13915, N13913);
xor XOR2 (N13916, N13915, N1267);
not NOT1 (N13917, N13907);
nor NOR3 (N13918, N13917, N7139, N10508);
nor NOR4 (N13919, N13916, N12930, N10233, N33);
nor NOR3 (N13920, N13908, N9448, N5378);
nand NAND4 (N13921, N13914, N6684, N5683, N625);
nor NOR2 (N13922, N13901, N3238);
and AND3 (N13923, N13906, N7797, N9102);
not NOT1 (N13924, N13921);
nand NAND2 (N13925, N13912, N9781);
and AND3 (N13926, N13918, N3925, N12608);
and AND3 (N13927, N13923, N8030, N9745);
not NOT1 (N13928, N13925);
buf BUF1 (N13929, N13919);
nand NAND4 (N13930, N13897, N12496, N13735, N10591);
nor NOR2 (N13931, N13930, N12794);
nor NOR4 (N13932, N13922, N5148, N2394, N8840);
nor NOR2 (N13933, N13924, N9446);
or OR4 (N13934, N13928, N6273, N9557, N9619);
nand NAND2 (N13935, N13920, N6426);
buf BUF1 (N13936, N13910);
nor NOR3 (N13937, N13935, N6412, N575);
and AND4 (N13938, N13933, N5321, N2666, N4909);
not NOT1 (N13939, N13937);
not NOT1 (N13940, N13926);
buf BUF1 (N13941, N13939);
not NOT1 (N13942, N13932);
or OR2 (N13943, N13942, N3007);
xor XOR2 (N13944, N13941, N8400);
not NOT1 (N13945, N13911);
nor NOR3 (N13946, N13945, N6041, N9382);
nor NOR4 (N13947, N13936, N9691, N10393, N12250);
xor XOR2 (N13948, N13929, N10836);
nor NOR4 (N13949, N13946, N10885, N9982, N7116);
nor NOR2 (N13950, N13943, N13001);
not NOT1 (N13951, N13948);
or OR4 (N13952, N13944, N7652, N865, N8579);
nor NOR4 (N13953, N13952, N4323, N8027, N7789);
or OR2 (N13954, N13949, N2709);
nand NAND2 (N13955, N13927, N1162);
and AND2 (N13956, N13955, N2960);
nor NOR2 (N13957, N13956, N4420);
not NOT1 (N13958, N13954);
buf BUF1 (N13959, N13958);
buf BUF1 (N13960, N13931);
or OR2 (N13961, N13938, N2365);
xor XOR2 (N13962, N13951, N8871);
and AND2 (N13963, N13957, N10898);
or OR2 (N13964, N13934, N3025);
or OR4 (N13965, N13947, N3942, N7580, N12751);
xor XOR2 (N13966, N13960, N3375);
not NOT1 (N13967, N13965);
nand NAND3 (N13968, N13959, N3875, N8794);
and AND2 (N13969, N13953, N3548);
nor NOR2 (N13970, N13969, N7856);
not NOT1 (N13971, N13964);
nand NAND2 (N13972, N13962, N2769);
nand NAND4 (N13973, N13972, N12132, N5722, N266);
xor XOR2 (N13974, N13940, N1182);
and AND3 (N13975, N13971, N13647, N8514);
buf BUF1 (N13976, N13975);
nor NOR3 (N13977, N13967, N11403, N1675);
nand NAND2 (N13978, N13973, N7640);
or OR2 (N13979, N13966, N11840);
or OR3 (N13980, N13963, N13879, N7339);
nand NAND4 (N13981, N13968, N5223, N4966, N4283);
and AND4 (N13982, N13974, N2864, N597, N12932);
nor NOR4 (N13983, N13976, N7081, N3927, N724);
buf BUF1 (N13984, N13961);
or OR4 (N13985, N13984, N6215, N6070, N10159);
and AND4 (N13986, N13981, N9617, N12473, N4237);
and AND2 (N13987, N13979, N663);
buf BUF1 (N13988, N13970);
buf BUF1 (N13989, N13988);
nand NAND2 (N13990, N13950, N6090);
buf BUF1 (N13991, N13987);
and AND4 (N13992, N13980, N11548, N1059, N2977);
or OR2 (N13993, N13983, N7860);
and AND4 (N13994, N13992, N4105, N13617, N9249);
nand NAND4 (N13995, N13986, N8849, N4395, N7534);
nand NAND3 (N13996, N13991, N2870, N12723);
xor XOR2 (N13997, N13996, N10734);
buf BUF1 (N13998, N13982);
xor XOR2 (N13999, N13998, N1670);
nand NAND4 (N14000, N13990, N13638, N2016, N9190);
nand NAND3 (N14001, N13978, N1628, N8346);
or OR2 (N14002, N13993, N3645);
or OR3 (N14003, N14000, N8820, N8143);
and AND3 (N14004, N13977, N5154, N8762);
or OR3 (N14005, N13994, N6838, N13365);
or OR3 (N14006, N14005, N10280, N3001);
xor XOR2 (N14007, N13985, N12653);
not NOT1 (N14008, N14007);
or OR4 (N14009, N13997, N8754, N12620, N6644);
nor NOR3 (N14010, N14006, N11766, N1725);
or OR3 (N14011, N14010, N9776, N9432);
not NOT1 (N14012, N14003);
xor XOR2 (N14013, N13995, N4933);
xor XOR2 (N14014, N14001, N5649);
not NOT1 (N14015, N14011);
and AND4 (N14016, N14004, N5453, N13672, N3959);
buf BUF1 (N14017, N14013);
buf BUF1 (N14018, N13989);
xor XOR2 (N14019, N14012, N7847);
nand NAND2 (N14020, N14002, N4464);
or OR4 (N14021, N14009, N11374, N10471, N10226);
or OR4 (N14022, N14021, N6606, N8415, N5654);
or OR3 (N14023, N13999, N10917, N5625);
nor NOR3 (N14024, N14015, N7206, N13192);
xor XOR2 (N14025, N14024, N4356);
nor NOR2 (N14026, N14016, N3454);
not NOT1 (N14027, N14020);
nand NAND4 (N14028, N14017, N11524, N8574, N8921);
not NOT1 (N14029, N14023);
or OR2 (N14030, N14022, N6854);
xor XOR2 (N14031, N14008, N5634);
nand NAND4 (N14032, N14027, N13719, N13730, N7680);
or OR2 (N14033, N14030, N10141);
xor XOR2 (N14034, N14014, N11212);
nand NAND4 (N14035, N14033, N794, N6819, N11997);
or OR3 (N14036, N14018, N1919, N9287);
nor NOR2 (N14037, N14035, N8980);
buf BUF1 (N14038, N14037);
nand NAND3 (N14039, N14029, N9382, N13018);
buf BUF1 (N14040, N14019);
xor XOR2 (N14041, N14040, N13189);
xor XOR2 (N14042, N14041, N5573);
nand NAND3 (N14043, N14026, N13091, N632);
not NOT1 (N14044, N14036);
buf BUF1 (N14045, N14038);
nor NOR3 (N14046, N14042, N9349, N11772);
or OR2 (N14047, N14043, N3234);
nor NOR3 (N14048, N14034, N4275, N11692);
nor NOR2 (N14049, N14048, N13381);
or OR3 (N14050, N14044, N13503, N8658);
and AND4 (N14051, N14032, N2578, N13190, N5096);
xor XOR2 (N14052, N14039, N4463);
and AND2 (N14053, N14046, N1136);
not NOT1 (N14054, N14052);
xor XOR2 (N14055, N14053, N10102);
or OR2 (N14056, N14051, N9681);
xor XOR2 (N14057, N14049, N2110);
buf BUF1 (N14058, N14047);
buf BUF1 (N14059, N14058);
and AND4 (N14060, N14028, N6456, N11393, N3467);
xor XOR2 (N14061, N14055, N11082);
not NOT1 (N14062, N14050);
buf BUF1 (N14063, N14056);
nand NAND3 (N14064, N14060, N1342, N1623);
buf BUF1 (N14065, N14031);
and AND4 (N14066, N14045, N11370, N6903, N11612);
xor XOR2 (N14067, N14062, N7325);
and AND3 (N14068, N14063, N11446, N12568);
buf BUF1 (N14069, N14057);
or OR2 (N14070, N14069, N3507);
or OR2 (N14071, N14065, N11908);
not NOT1 (N14072, N14064);
buf BUF1 (N14073, N14059);
nand NAND3 (N14074, N14071, N10414, N12434);
nor NOR4 (N14075, N14070, N11888, N9208, N6734);
or OR4 (N14076, N14067, N7890, N7875, N2841);
nor NOR4 (N14077, N14068, N11259, N1530, N13500);
and AND4 (N14078, N14075, N1527, N13709, N13278);
nand NAND4 (N14079, N14078, N5642, N12894, N462);
xor XOR2 (N14080, N14079, N7208);
nor NOR4 (N14081, N14066, N56, N4870, N3468);
nand NAND4 (N14082, N14025, N1954, N12568, N7010);
or OR2 (N14083, N14081, N11094);
or OR3 (N14084, N14080, N2625, N7110);
and AND2 (N14085, N14076, N8187);
nor NOR3 (N14086, N14061, N1808, N11538);
or OR4 (N14087, N14072, N12784, N5650, N6729);
nand NAND4 (N14088, N14054, N6457, N6659, N3243);
xor XOR2 (N14089, N14086, N1701);
or OR2 (N14090, N14085, N4750);
nor NOR3 (N14091, N14090, N4182, N2018);
nand NAND3 (N14092, N14083, N12145, N5272);
xor XOR2 (N14093, N14091, N10537);
xor XOR2 (N14094, N14084, N7794);
buf BUF1 (N14095, N14094);
nand NAND4 (N14096, N14077, N8667, N12455, N8507);
not NOT1 (N14097, N14087);
not NOT1 (N14098, N14082);
xor XOR2 (N14099, N14089, N4369);
or OR2 (N14100, N14073, N9911);
nor NOR2 (N14101, N14098, N3980);
xor XOR2 (N14102, N14095, N1400);
or OR3 (N14103, N14074, N10159, N749);
xor XOR2 (N14104, N14102, N10314);
not NOT1 (N14105, N14097);
not NOT1 (N14106, N14088);
not NOT1 (N14107, N14106);
xor XOR2 (N14108, N14099, N1693);
not NOT1 (N14109, N14104);
buf BUF1 (N14110, N14096);
not NOT1 (N14111, N14105);
xor XOR2 (N14112, N14092, N12468);
nor NOR4 (N14113, N14111, N8077, N11203, N775);
buf BUF1 (N14114, N14103);
nand NAND2 (N14115, N14100, N1449);
and AND2 (N14116, N14115, N8965);
and AND2 (N14117, N14093, N442);
or OR3 (N14118, N14113, N5019, N6442);
xor XOR2 (N14119, N14110, N10038);
xor XOR2 (N14120, N14107, N4686);
and AND3 (N14121, N14101, N1792, N7551);
buf BUF1 (N14122, N14112);
nor NOR3 (N14123, N14121, N13702, N13361);
or OR2 (N14124, N14109, N11243);
xor XOR2 (N14125, N14119, N12432);
and AND4 (N14126, N14125, N2516, N4928, N6681);
nand NAND4 (N14127, N14114, N3838, N5749, N10061);
not NOT1 (N14128, N14127);
and AND2 (N14129, N14108, N12539);
nand NAND2 (N14130, N14129, N178);
and AND2 (N14131, N14120, N1014);
nor NOR2 (N14132, N14118, N5332);
nor NOR2 (N14133, N14117, N6573);
or OR3 (N14134, N14116, N3141, N10925);
not NOT1 (N14135, N14124);
xor XOR2 (N14136, N14134, N5789);
and AND4 (N14137, N14123, N1879, N933, N13983);
or OR3 (N14138, N14122, N9646, N2403);
xor XOR2 (N14139, N14137, N7817);
or OR2 (N14140, N14131, N10157);
nor NOR4 (N14141, N14133, N1121, N10819, N1422);
buf BUF1 (N14142, N14126);
not NOT1 (N14143, N14132);
xor XOR2 (N14144, N14135, N12029);
buf BUF1 (N14145, N14138);
or OR2 (N14146, N14139, N12802);
buf BUF1 (N14147, N14136);
not NOT1 (N14148, N14140);
nor NOR3 (N14149, N14147, N23, N2859);
nand NAND4 (N14150, N14143, N7035, N11654, N5344);
buf BUF1 (N14151, N14150);
xor XOR2 (N14152, N14144, N4191);
or OR4 (N14153, N14152, N6582, N2403, N2156);
or OR3 (N14154, N14141, N5053, N4482);
nor NOR4 (N14155, N14153, N11584, N11065, N12178);
buf BUF1 (N14156, N14142);
buf BUF1 (N14157, N14155);
nor NOR4 (N14158, N14154, N10441, N5138, N800);
buf BUF1 (N14159, N14148);
nor NOR4 (N14160, N14157, N11513, N8942, N679);
and AND2 (N14161, N14146, N2728);
not NOT1 (N14162, N14160);
xor XOR2 (N14163, N14159, N4850);
buf BUF1 (N14164, N14149);
buf BUF1 (N14165, N14161);
or OR3 (N14166, N14145, N11670, N5230);
not NOT1 (N14167, N14130);
or OR4 (N14168, N14167, N8642, N1546, N5942);
or OR2 (N14169, N14166, N6808);
or OR2 (N14170, N14158, N10732);
xor XOR2 (N14171, N14170, N2798);
buf BUF1 (N14172, N14163);
xor XOR2 (N14173, N14169, N8376);
nand NAND4 (N14174, N14165, N13164, N2328, N10960);
buf BUF1 (N14175, N14173);
and AND2 (N14176, N14164, N4116);
or OR4 (N14177, N14168, N5513, N5589, N11276);
nor NOR3 (N14178, N14128, N6316, N10191);
nor NOR3 (N14179, N14177, N10844, N3213);
nand NAND2 (N14180, N14179, N2567);
nor NOR4 (N14181, N14174, N9673, N13487, N7591);
nor NOR3 (N14182, N14171, N7561, N7054);
buf BUF1 (N14183, N14176);
or OR2 (N14184, N14172, N469);
nor NOR2 (N14185, N14175, N6768);
nand NAND3 (N14186, N14182, N1750, N7486);
or OR4 (N14187, N14180, N8121, N8587, N13404);
buf BUF1 (N14188, N14181);
nor NOR4 (N14189, N14162, N44, N13601, N11624);
and AND3 (N14190, N14178, N898, N11403);
or OR4 (N14191, N14183, N12189, N5778, N14072);
nand NAND4 (N14192, N14191, N107, N36, N3981);
nor NOR2 (N14193, N14187, N394);
xor XOR2 (N14194, N14156, N5474);
nand NAND2 (N14195, N14189, N913);
nand NAND2 (N14196, N14190, N8117);
not NOT1 (N14197, N14188);
not NOT1 (N14198, N14193);
nand NAND4 (N14199, N14197, N7501, N163, N8730);
nand NAND4 (N14200, N14192, N3255, N8671, N5848);
not NOT1 (N14201, N14198);
not NOT1 (N14202, N14185);
nor NOR3 (N14203, N14195, N11865, N5342);
nor NOR3 (N14204, N14196, N4870, N10696);
not NOT1 (N14205, N14184);
nor NOR4 (N14206, N14199, N9775, N8698, N5228);
and AND4 (N14207, N14206, N531, N2044, N13777);
not NOT1 (N14208, N14205);
and AND4 (N14209, N14200, N4177, N9057, N11703);
nand NAND3 (N14210, N14194, N11582, N12082);
buf BUF1 (N14211, N14210);
buf BUF1 (N14212, N14202);
nand NAND2 (N14213, N14208, N11325);
nand NAND3 (N14214, N14186, N3069, N13117);
buf BUF1 (N14215, N14207);
or OR3 (N14216, N14151, N11371, N11769);
nor NOR3 (N14217, N14214, N10219, N87);
and AND4 (N14218, N14212, N10440, N13517, N5960);
buf BUF1 (N14219, N14204);
buf BUF1 (N14220, N14217);
not NOT1 (N14221, N14220);
or OR3 (N14222, N14216, N12122, N2838);
and AND3 (N14223, N14215, N8366, N2723);
or OR2 (N14224, N14211, N5812);
not NOT1 (N14225, N14209);
or OR2 (N14226, N14219, N1465);
nor NOR2 (N14227, N14225, N6328);
or OR4 (N14228, N14203, N10811, N7477, N810);
buf BUF1 (N14229, N14223);
nand NAND3 (N14230, N14224, N11995, N11841);
or OR2 (N14231, N14218, N10072);
xor XOR2 (N14232, N14227, N111);
nand NAND3 (N14233, N14201, N977, N2321);
nand NAND3 (N14234, N14229, N11338, N4056);
not NOT1 (N14235, N14221);
nand NAND4 (N14236, N14231, N192, N5132, N2414);
not NOT1 (N14237, N14232);
nor NOR3 (N14238, N14236, N840, N8073);
and AND2 (N14239, N14213, N2809);
not NOT1 (N14240, N14238);
or OR2 (N14241, N14222, N12990);
or OR2 (N14242, N14228, N11419);
xor XOR2 (N14243, N14233, N8220);
buf BUF1 (N14244, N14243);
xor XOR2 (N14245, N14234, N8597);
buf BUF1 (N14246, N14237);
or OR3 (N14247, N14235, N461, N4023);
nand NAND2 (N14248, N14226, N8637);
or OR4 (N14249, N14230, N2502, N7478, N7746);
buf BUF1 (N14250, N14242);
and AND4 (N14251, N14240, N12640, N7703, N1796);
xor XOR2 (N14252, N14247, N10563);
not NOT1 (N14253, N14245);
not NOT1 (N14254, N14253);
not NOT1 (N14255, N14250);
buf BUF1 (N14256, N14241);
or OR4 (N14257, N14251, N4261, N9710, N4951);
and AND2 (N14258, N14254, N12572);
nand NAND2 (N14259, N14252, N13091);
and AND2 (N14260, N14255, N919);
xor XOR2 (N14261, N14259, N6784);
and AND2 (N14262, N14246, N14017);
not NOT1 (N14263, N14260);
not NOT1 (N14264, N14248);
nor NOR2 (N14265, N14264, N3155);
xor XOR2 (N14266, N14244, N2242);
buf BUF1 (N14267, N14249);
and AND3 (N14268, N14262, N6102, N145);
nand NAND4 (N14269, N14257, N4531, N2580, N12403);
xor XOR2 (N14270, N14261, N3337);
buf BUF1 (N14271, N14270);
or OR4 (N14272, N14265, N11255, N4711, N7081);
nor NOR2 (N14273, N14272, N4726);
and AND4 (N14274, N14266, N6759, N6609, N2029);
xor XOR2 (N14275, N14239, N879);
and AND2 (N14276, N14256, N9753);
nand NAND2 (N14277, N14276, N12993);
or OR2 (N14278, N14267, N13886);
and AND2 (N14279, N14278, N1171);
buf BUF1 (N14280, N14277);
buf BUF1 (N14281, N14263);
and AND3 (N14282, N14273, N1515, N12806);
not NOT1 (N14283, N14279);
buf BUF1 (N14284, N14282);
nand NAND4 (N14285, N14271, N1460, N1453, N11636);
nor NOR2 (N14286, N14275, N1506);
xor XOR2 (N14287, N14281, N13888);
buf BUF1 (N14288, N14284);
xor XOR2 (N14289, N14269, N5929);
not NOT1 (N14290, N14283);
not NOT1 (N14291, N14280);
not NOT1 (N14292, N14288);
not NOT1 (N14293, N14290);
or OR4 (N14294, N14293, N11908, N9967, N13341);
nand NAND4 (N14295, N14294, N8940, N9740, N8076);
nor NOR3 (N14296, N14287, N2892, N8929);
and AND3 (N14297, N14286, N3534, N11203);
not NOT1 (N14298, N14285);
or OR2 (N14299, N14258, N4749);
or OR3 (N14300, N14298, N2852, N4153);
or OR4 (N14301, N14274, N954, N2608, N12337);
buf BUF1 (N14302, N14301);
xor XOR2 (N14303, N14296, N3656);
and AND3 (N14304, N14292, N9277, N13385);
buf BUF1 (N14305, N14291);
nor NOR2 (N14306, N14297, N12051);
nor NOR3 (N14307, N14304, N8887, N9510);
nand NAND2 (N14308, N14306, N12895);
buf BUF1 (N14309, N14305);
or OR4 (N14310, N14307, N9222, N9287, N13714);
or OR3 (N14311, N14309, N7872, N1604);
not NOT1 (N14312, N14295);
and AND4 (N14313, N14312, N3273, N14119, N9986);
not NOT1 (N14314, N14302);
buf BUF1 (N14315, N14308);
not NOT1 (N14316, N14310);
not NOT1 (N14317, N14315);
and AND3 (N14318, N14311, N3501, N4546);
xor XOR2 (N14319, N14299, N4950);
not NOT1 (N14320, N14316);
buf BUF1 (N14321, N14303);
and AND4 (N14322, N14320, N1550, N10269, N3579);
not NOT1 (N14323, N14268);
and AND3 (N14324, N14300, N2643, N2554);
not NOT1 (N14325, N14319);
not NOT1 (N14326, N14314);
xor XOR2 (N14327, N14289, N1449);
nor NOR2 (N14328, N14313, N3892);
and AND2 (N14329, N14325, N10087);
nor NOR4 (N14330, N14328, N8537, N14069, N1490);
buf BUF1 (N14331, N14324);
not NOT1 (N14332, N14323);
xor XOR2 (N14333, N14318, N4935);
nand NAND4 (N14334, N14329, N3266, N14264, N13144);
xor XOR2 (N14335, N14327, N1247);
not NOT1 (N14336, N14321);
buf BUF1 (N14337, N14331);
xor XOR2 (N14338, N14337, N12941);
or OR4 (N14339, N14322, N1792, N10633, N7247);
or OR3 (N14340, N14326, N11500, N6385);
and AND2 (N14341, N14330, N4287);
buf BUF1 (N14342, N14332);
nand NAND2 (N14343, N14317, N4334);
xor XOR2 (N14344, N14339, N644);
nand NAND4 (N14345, N14333, N3248, N13077, N1291);
xor XOR2 (N14346, N14334, N977);
not NOT1 (N14347, N14342);
nand NAND4 (N14348, N14345, N928, N10989, N9766);
not NOT1 (N14349, N14343);
xor XOR2 (N14350, N14344, N636);
and AND4 (N14351, N14346, N11941, N3655, N11893);
xor XOR2 (N14352, N14351, N7897);
nand NAND3 (N14353, N14349, N5693, N5904);
or OR4 (N14354, N14352, N2234, N880, N7003);
and AND2 (N14355, N14353, N11982);
or OR4 (N14356, N14341, N13638, N8914, N9592);
nor NOR4 (N14357, N14336, N7373, N14107, N2319);
not NOT1 (N14358, N14357);
and AND3 (N14359, N14355, N14082, N4012);
nand NAND3 (N14360, N14340, N10420, N8929);
xor XOR2 (N14361, N14347, N5956);
and AND3 (N14362, N14360, N12536, N10036);
nand NAND3 (N14363, N14361, N10751, N9706);
nand NAND3 (N14364, N14356, N13612, N279);
nand NAND3 (N14365, N14350, N3514, N12292);
nor NOR2 (N14366, N14364, N11354);
buf BUF1 (N14367, N14362);
nor NOR4 (N14368, N14348, N1593, N6661, N11235);
or OR4 (N14369, N14335, N13577, N7023, N6544);
not NOT1 (N14370, N14366);
nand NAND4 (N14371, N14363, N8617, N4224, N9715);
nand NAND2 (N14372, N14338, N8821);
buf BUF1 (N14373, N14370);
buf BUF1 (N14374, N14372);
xor XOR2 (N14375, N14365, N6921);
or OR4 (N14376, N14375, N568, N9422, N6200);
xor XOR2 (N14377, N14354, N12809);
xor XOR2 (N14378, N14377, N12748);
nor NOR3 (N14379, N14358, N3987, N12078);
nand NAND4 (N14380, N14376, N13037, N12463, N13180);
or OR4 (N14381, N14367, N12082, N8107, N13858);
and AND2 (N14382, N14368, N3997);
buf BUF1 (N14383, N14371);
nor NOR3 (N14384, N14383, N5720, N11114);
xor XOR2 (N14385, N14379, N4150);
nand NAND3 (N14386, N14373, N7347, N4088);
not NOT1 (N14387, N14369);
nand NAND4 (N14388, N14378, N4115, N3010, N12378);
not NOT1 (N14389, N14380);
not NOT1 (N14390, N14374);
or OR2 (N14391, N14390, N3601);
buf BUF1 (N14392, N14384);
buf BUF1 (N14393, N14388);
buf BUF1 (N14394, N14382);
or OR3 (N14395, N14394, N7649, N3713);
nor NOR4 (N14396, N14359, N629, N6307, N6676);
buf BUF1 (N14397, N14385);
and AND2 (N14398, N14397, N10707);
and AND2 (N14399, N14391, N4402);
and AND4 (N14400, N14393, N3782, N2094, N13738);
xor XOR2 (N14401, N14398, N3755);
and AND2 (N14402, N14389, N5610);
and AND4 (N14403, N14395, N11292, N2321, N1674);
or OR2 (N14404, N14392, N10366);
nand NAND4 (N14405, N14396, N10710, N3180, N7156);
xor XOR2 (N14406, N14401, N844);
buf BUF1 (N14407, N14403);
and AND3 (N14408, N14399, N11566, N5675);
or OR2 (N14409, N14408, N1283);
not NOT1 (N14410, N14386);
nand NAND3 (N14411, N14410, N7310, N6338);
or OR4 (N14412, N14409, N405, N7656, N13677);
buf BUF1 (N14413, N14381);
or OR4 (N14414, N14402, N1568, N9863, N9586);
xor XOR2 (N14415, N14414, N3633);
or OR2 (N14416, N14387, N13836);
not NOT1 (N14417, N14413);
nand NAND3 (N14418, N14415, N3921, N1488);
nor NOR3 (N14419, N14416, N1390, N2090);
not NOT1 (N14420, N14407);
nand NAND3 (N14421, N14406, N7907, N2508);
or OR3 (N14422, N14405, N12140, N9421);
and AND4 (N14423, N14400, N3366, N9304, N13830);
not NOT1 (N14424, N14417);
xor XOR2 (N14425, N14423, N2823);
or OR3 (N14426, N14412, N6500, N12483);
xor XOR2 (N14427, N14404, N5522);
nand NAND3 (N14428, N14421, N7809, N584);
not NOT1 (N14429, N14422);
xor XOR2 (N14430, N14411, N7091);
and AND2 (N14431, N14420, N3703);
nand NAND4 (N14432, N14431, N6283, N9481, N1179);
and AND4 (N14433, N14426, N6159, N12538, N5536);
or OR4 (N14434, N14432, N2366, N9932, N11902);
or OR2 (N14435, N14419, N8457);
buf BUF1 (N14436, N14425);
and AND4 (N14437, N14436, N7437, N13854, N2113);
nand NAND3 (N14438, N14427, N2227, N9534);
not NOT1 (N14439, N14429);
and AND2 (N14440, N14433, N4145);
and AND2 (N14441, N14434, N13033);
nand NAND2 (N14442, N14435, N13774);
and AND3 (N14443, N14438, N6082, N26);
nor NOR2 (N14444, N14418, N12164);
not NOT1 (N14445, N14442);
xor XOR2 (N14446, N14445, N10513);
or OR4 (N14447, N14439, N7472, N7408, N11554);
nor NOR4 (N14448, N14447, N3914, N4167, N5920);
nor NOR3 (N14449, N14437, N2150, N6520);
not NOT1 (N14450, N14440);
not NOT1 (N14451, N14446);
and AND2 (N14452, N14443, N4349);
nand NAND3 (N14453, N14428, N9270, N10787);
and AND4 (N14454, N14450, N8315, N8000, N12063);
buf BUF1 (N14455, N14453);
or OR4 (N14456, N14449, N4495, N3349, N3663);
and AND4 (N14457, N14441, N1135, N11125, N8842);
nor NOR4 (N14458, N14454, N13061, N393, N9784);
not NOT1 (N14459, N14430);
or OR3 (N14460, N14455, N4926, N7768);
nand NAND2 (N14461, N14451, N118);
nand NAND2 (N14462, N14457, N9993);
xor XOR2 (N14463, N14458, N12321);
xor XOR2 (N14464, N14460, N6566);
nand NAND2 (N14465, N14444, N1905);
or OR2 (N14466, N14461, N14456);
not NOT1 (N14467, N10396);
xor XOR2 (N14468, N14465, N5606);
xor XOR2 (N14469, N14459, N10988);
and AND2 (N14470, N14467, N12131);
xor XOR2 (N14471, N14468, N10740);
and AND4 (N14472, N14452, N215, N6817, N11327);
nand NAND3 (N14473, N14469, N10355, N2007);
and AND2 (N14474, N14448, N12545);
and AND3 (N14475, N14473, N4108, N10526);
nand NAND4 (N14476, N14466, N13886, N2010, N12334);
xor XOR2 (N14477, N14471, N8948);
buf BUF1 (N14478, N14477);
not NOT1 (N14479, N14474);
nor NOR2 (N14480, N14479, N10098);
nand NAND2 (N14481, N14476, N8087);
buf BUF1 (N14482, N14424);
and AND3 (N14483, N14478, N3242, N116);
and AND2 (N14484, N14464, N3936);
not NOT1 (N14485, N14480);
and AND2 (N14486, N14472, N14387);
or OR4 (N14487, N14463, N7072, N3209, N9967);
nand NAND3 (N14488, N14485, N6518, N5764);
not NOT1 (N14489, N14488);
or OR4 (N14490, N14481, N5055, N6325, N4119);
buf BUF1 (N14491, N14475);
and AND4 (N14492, N14470, N481, N6861, N1048);
and AND4 (N14493, N14486, N3644, N12312, N985);
and AND2 (N14494, N14487, N11152);
or OR4 (N14495, N14494, N12124, N12968, N2045);
nand NAND4 (N14496, N14491, N11527, N9830, N4322);
buf BUF1 (N14497, N14496);
xor XOR2 (N14498, N14489, N9820);
and AND2 (N14499, N14484, N9643);
buf BUF1 (N14500, N14498);
not NOT1 (N14501, N14492);
xor XOR2 (N14502, N14497, N548);
nand NAND4 (N14503, N14483, N4000, N2984, N13643);
xor XOR2 (N14504, N14462, N6862);
buf BUF1 (N14505, N14503);
not NOT1 (N14506, N14502);
nor NOR3 (N14507, N14505, N2725, N3504);
and AND2 (N14508, N14493, N9825);
nand NAND4 (N14509, N14490, N13658, N7568, N11978);
buf BUF1 (N14510, N14500);
buf BUF1 (N14511, N14507);
not NOT1 (N14512, N14504);
and AND2 (N14513, N14512, N3173);
xor XOR2 (N14514, N14499, N2784);
buf BUF1 (N14515, N14511);
xor XOR2 (N14516, N14495, N11941);
nand NAND2 (N14517, N14482, N8077);
not NOT1 (N14518, N14516);
nor NOR3 (N14519, N14513, N12958, N12712);
not NOT1 (N14520, N14518);
xor XOR2 (N14521, N14515, N10343);
nand NAND4 (N14522, N14509, N7151, N1386, N897);
nand NAND4 (N14523, N14506, N11437, N200, N13003);
buf BUF1 (N14524, N14522);
or OR3 (N14525, N14519, N10564, N11152);
buf BUF1 (N14526, N14521);
xor XOR2 (N14527, N14525, N12680);
and AND2 (N14528, N14501, N4062);
buf BUF1 (N14529, N14523);
and AND3 (N14530, N14524, N11197, N7490);
buf BUF1 (N14531, N14530);
or OR3 (N14532, N14520, N13769, N6352);
nor NOR4 (N14533, N14532, N11095, N833, N5961);
or OR2 (N14534, N14533, N9356);
buf BUF1 (N14535, N14528);
xor XOR2 (N14536, N14517, N10078);
buf BUF1 (N14537, N14531);
nor NOR3 (N14538, N14537, N5812, N9748);
not NOT1 (N14539, N14529);
nand NAND4 (N14540, N14538, N10949, N8150, N3228);
not NOT1 (N14541, N14508);
not NOT1 (N14542, N14514);
nand NAND4 (N14543, N14534, N14172, N5478, N3986);
not NOT1 (N14544, N14541);
or OR2 (N14545, N14539, N7853);
or OR3 (N14546, N14527, N5305, N8875);
nor NOR4 (N14547, N14510, N7265, N6078, N9885);
buf BUF1 (N14548, N14546);
and AND3 (N14549, N14547, N12184, N8071);
not NOT1 (N14550, N14535);
nor NOR2 (N14551, N14526, N7010);
nor NOR2 (N14552, N14545, N8329);
xor XOR2 (N14553, N14549, N8745);
and AND2 (N14554, N14551, N12364);
buf BUF1 (N14555, N14536);
or OR2 (N14556, N14550, N834);
nand NAND3 (N14557, N14555, N3091, N7837);
buf BUF1 (N14558, N14554);
and AND3 (N14559, N14542, N4015, N12927);
nor NOR2 (N14560, N14540, N14395);
or OR2 (N14561, N14544, N10073);
buf BUF1 (N14562, N14543);
nor NOR3 (N14563, N14560, N5393, N3846);
and AND4 (N14564, N14557, N5213, N10084, N6788);
nor NOR4 (N14565, N14548, N14394, N10584, N1217);
or OR2 (N14566, N14562, N14043);
nand NAND2 (N14567, N14564, N5236);
nor NOR3 (N14568, N14558, N2707, N14439);
xor XOR2 (N14569, N14566, N13280);
nand NAND2 (N14570, N14569, N2149);
and AND3 (N14571, N14563, N3597, N3217);
not NOT1 (N14572, N14556);
not NOT1 (N14573, N14565);
not NOT1 (N14574, N14571);
xor XOR2 (N14575, N14567, N2680);
and AND3 (N14576, N14572, N14324, N8528);
buf BUF1 (N14577, N14574);
nand NAND4 (N14578, N14573, N9507, N1254, N3497);
buf BUF1 (N14579, N14561);
buf BUF1 (N14580, N14579);
or OR2 (N14581, N14578, N3187);
buf BUF1 (N14582, N14559);
nor NOR2 (N14583, N14553, N9802);
not NOT1 (N14584, N14575);
or OR3 (N14585, N14583, N5210, N6280);
nand NAND3 (N14586, N14584, N4549, N5324);
not NOT1 (N14587, N14581);
xor XOR2 (N14588, N14582, N8889);
and AND2 (N14589, N14585, N1413);
or OR2 (N14590, N14589, N226);
not NOT1 (N14591, N14576);
nor NOR3 (N14592, N14577, N251, N3161);
nand NAND4 (N14593, N14580, N5043, N8524, N7706);
buf BUF1 (N14594, N14587);
buf BUF1 (N14595, N14568);
or OR2 (N14596, N14590, N4213);
not NOT1 (N14597, N14586);
xor XOR2 (N14598, N14597, N11863);
buf BUF1 (N14599, N14592);
xor XOR2 (N14600, N14593, N718);
not NOT1 (N14601, N14598);
and AND2 (N14602, N14552, N3262);
buf BUF1 (N14603, N14588);
buf BUF1 (N14604, N14602);
xor XOR2 (N14605, N14600, N5733);
nand NAND3 (N14606, N14603, N1616, N7788);
nand NAND4 (N14607, N14604, N11048, N13716, N1802);
or OR4 (N14608, N14570, N2459, N5711, N1732);
nand NAND3 (N14609, N14596, N14548, N11626);
or OR2 (N14610, N14601, N7068);
or OR2 (N14611, N14591, N6337);
buf BUF1 (N14612, N14594);
not NOT1 (N14613, N14611);
and AND3 (N14614, N14608, N9027, N10679);
and AND4 (N14615, N14605, N11225, N11319, N5204);
or OR2 (N14616, N14606, N1935);
nor NOR3 (N14617, N14607, N10170, N13314);
and AND4 (N14618, N14617, N4377, N7792, N4386);
and AND2 (N14619, N14615, N12884);
not NOT1 (N14620, N14610);
and AND3 (N14621, N14595, N7745, N8338);
nand NAND2 (N14622, N14614, N430);
buf BUF1 (N14623, N14599);
nor NOR3 (N14624, N14620, N5123, N11977);
and AND2 (N14625, N14624, N10271);
or OR4 (N14626, N14622, N8929, N11511, N2008);
buf BUF1 (N14627, N14616);
nor NOR3 (N14628, N14609, N3558, N4632);
and AND4 (N14629, N14626, N3338, N6552, N11403);
nor NOR4 (N14630, N14618, N12401, N3983, N564);
buf BUF1 (N14631, N14630);
buf BUF1 (N14632, N14621);
and AND3 (N14633, N14627, N8124, N13090);
not NOT1 (N14634, N14612);
and AND4 (N14635, N14625, N3486, N1102, N8896);
not NOT1 (N14636, N14628);
or OR4 (N14637, N14632, N12178, N14183, N12929);
not NOT1 (N14638, N14634);
nor NOR2 (N14639, N14633, N6744);
nor NOR2 (N14640, N14636, N8544);
or OR3 (N14641, N14629, N5209, N5131);
or OR2 (N14642, N14640, N5642);
and AND3 (N14643, N14638, N5713, N1859);
nand NAND2 (N14644, N14613, N8545);
xor XOR2 (N14645, N14642, N6563);
not NOT1 (N14646, N14637);
nor NOR4 (N14647, N14646, N2847, N602, N7570);
nand NAND3 (N14648, N14641, N10179, N8192);
xor XOR2 (N14649, N14635, N1197);
not NOT1 (N14650, N14631);
or OR3 (N14651, N14623, N10618, N2267);
or OR2 (N14652, N14643, N12907);
nand NAND2 (N14653, N14648, N5327);
nand NAND4 (N14654, N14644, N3757, N13394, N5202);
buf BUF1 (N14655, N14652);
nor NOR4 (N14656, N14639, N3266, N14379, N7232);
not NOT1 (N14657, N14645);
buf BUF1 (N14658, N14654);
xor XOR2 (N14659, N14651, N6547);
not NOT1 (N14660, N14655);
not NOT1 (N14661, N14650);
not NOT1 (N14662, N14619);
buf BUF1 (N14663, N14649);
buf BUF1 (N14664, N14653);
xor XOR2 (N14665, N14663, N8409);
not NOT1 (N14666, N14647);
buf BUF1 (N14667, N14661);
nor NOR3 (N14668, N14660, N13717, N5426);
buf BUF1 (N14669, N14664);
or OR3 (N14670, N14662, N683, N386);
buf BUF1 (N14671, N14667);
nor NOR4 (N14672, N14659, N5217, N6983, N6831);
or OR2 (N14673, N14671, N620);
nor NOR3 (N14674, N14672, N8784, N5389);
xor XOR2 (N14675, N14666, N5168);
or OR3 (N14676, N14674, N9312, N9616);
nand NAND3 (N14677, N14665, N7763, N7608);
not NOT1 (N14678, N14668);
nor NOR4 (N14679, N14657, N3025, N8679, N14367);
and AND3 (N14680, N14676, N6536, N9714);
buf BUF1 (N14681, N14670);
xor XOR2 (N14682, N14658, N11791);
buf BUF1 (N14683, N14677);
nand NAND2 (N14684, N14656, N11524);
not NOT1 (N14685, N14683);
and AND3 (N14686, N14669, N3302, N8775);
nand NAND3 (N14687, N14679, N14024, N11557);
and AND3 (N14688, N14681, N14084, N4069);
and AND3 (N14689, N14684, N9866, N8987);
buf BUF1 (N14690, N14675);
or OR2 (N14691, N14682, N5267);
not NOT1 (N14692, N14686);
xor XOR2 (N14693, N14673, N12227);
and AND3 (N14694, N14693, N10594, N9306);
xor XOR2 (N14695, N14687, N5106);
nor NOR4 (N14696, N14688, N12108, N9867, N8650);
buf BUF1 (N14697, N14692);
not NOT1 (N14698, N14680);
or OR4 (N14699, N14685, N11165, N6339, N9076);
and AND2 (N14700, N14691, N12894);
xor XOR2 (N14701, N14697, N8720);
and AND4 (N14702, N14696, N12484, N9125, N8564);
xor XOR2 (N14703, N14702, N3469);
or OR4 (N14704, N14698, N4098, N2651, N2847);
nor NOR3 (N14705, N14690, N6056, N6451);
xor XOR2 (N14706, N14704, N11793);
nand NAND2 (N14707, N14703, N9954);
buf BUF1 (N14708, N14700);
nand NAND3 (N14709, N14689, N376, N454);
not NOT1 (N14710, N14701);
xor XOR2 (N14711, N14705, N12420);
buf BUF1 (N14712, N14708);
or OR2 (N14713, N14695, N9375);
not NOT1 (N14714, N14711);
nand NAND3 (N14715, N14694, N1968, N5777);
buf BUF1 (N14716, N14714);
not NOT1 (N14717, N14678);
buf BUF1 (N14718, N14712);
xor XOR2 (N14719, N14699, N5056);
buf BUF1 (N14720, N14709);
xor XOR2 (N14721, N14719, N10503);
nand NAND4 (N14722, N14707, N8638, N11506, N7574);
xor XOR2 (N14723, N14713, N4342);
and AND2 (N14724, N14723, N11614);
xor XOR2 (N14725, N14716, N12681);
or OR3 (N14726, N14722, N14722, N6740);
nand NAND4 (N14727, N14725, N14089, N14273, N12250);
or OR2 (N14728, N14715, N11300);
xor XOR2 (N14729, N14724, N14372);
not NOT1 (N14730, N14728);
and AND3 (N14731, N14726, N1991, N723);
nor NOR3 (N14732, N14710, N3377, N13658);
nor NOR4 (N14733, N14731, N12119, N4924, N10280);
nor NOR2 (N14734, N14733, N13547);
buf BUF1 (N14735, N14717);
and AND4 (N14736, N14706, N6748, N12849, N4208);
or OR2 (N14737, N14721, N3608);
not NOT1 (N14738, N14735);
not NOT1 (N14739, N14732);
not NOT1 (N14740, N14737);
nand NAND4 (N14741, N14736, N11409, N10590, N3316);
xor XOR2 (N14742, N14739, N6014);
and AND4 (N14743, N14718, N927, N13996, N12332);
not NOT1 (N14744, N14720);
xor XOR2 (N14745, N14734, N9480);
not NOT1 (N14746, N14744);
and AND2 (N14747, N14730, N1756);
and AND2 (N14748, N14727, N10489);
xor XOR2 (N14749, N14748, N14649);
or OR3 (N14750, N14745, N1873, N10935);
or OR4 (N14751, N14742, N14734, N1492, N9763);
nand NAND3 (N14752, N14750, N13461, N1675);
nor NOR2 (N14753, N14743, N2716);
buf BUF1 (N14754, N14740);
buf BUF1 (N14755, N14753);
nor NOR3 (N14756, N14751, N7965, N8652);
nor NOR4 (N14757, N14749, N2584, N13775, N3329);
buf BUF1 (N14758, N14741);
nand NAND4 (N14759, N14755, N1787, N410, N7016);
buf BUF1 (N14760, N14752);
buf BUF1 (N14761, N14759);
not NOT1 (N14762, N14760);
buf BUF1 (N14763, N14754);
not NOT1 (N14764, N14761);
not NOT1 (N14765, N14757);
or OR4 (N14766, N14764, N3988, N9711, N7217);
and AND2 (N14767, N14765, N10719);
nor NOR3 (N14768, N14763, N5227, N5583);
not NOT1 (N14769, N14756);
not NOT1 (N14770, N14746);
or OR4 (N14771, N14747, N1437, N12055, N7248);
not NOT1 (N14772, N14771);
buf BUF1 (N14773, N14729);
xor XOR2 (N14774, N14768, N12575);
xor XOR2 (N14775, N14772, N5572);
or OR3 (N14776, N14762, N6190, N11750);
buf BUF1 (N14777, N14775);
nor NOR4 (N14778, N14774, N5041, N252, N12044);
nand NAND2 (N14779, N14770, N11914);
nor NOR4 (N14780, N14758, N9849, N8890, N12389);
not NOT1 (N14781, N14776);
nand NAND2 (N14782, N14779, N12563);
not NOT1 (N14783, N14769);
or OR3 (N14784, N14782, N3971, N14445);
and AND3 (N14785, N14738, N5038, N13000);
nand NAND3 (N14786, N14766, N5587, N6698);
and AND4 (N14787, N14777, N2865, N4991, N9018);
and AND2 (N14788, N14787, N12125);
xor XOR2 (N14789, N14767, N11186);
nand NAND2 (N14790, N14780, N5610);
nand NAND2 (N14791, N14781, N6760);
or OR3 (N14792, N14778, N1551, N4150);
and AND2 (N14793, N14784, N4225);
or OR4 (N14794, N14788, N4988, N2000, N5780);
nand NAND2 (N14795, N14793, N1476);
nand NAND2 (N14796, N14791, N11698);
and AND2 (N14797, N14786, N6998);
buf BUF1 (N14798, N14794);
or OR4 (N14799, N14783, N5600, N8114, N9772);
nor NOR4 (N14800, N14795, N3340, N2392, N2186);
nand NAND3 (N14801, N14785, N9192, N8695);
nor NOR4 (N14802, N14801, N5726, N5711, N12599);
and AND4 (N14803, N14798, N2269, N4996, N10194);
nand NAND2 (N14804, N14789, N13915);
or OR3 (N14805, N14797, N12836, N3289);
xor XOR2 (N14806, N14805, N7713);
not NOT1 (N14807, N14804);
and AND4 (N14808, N14796, N10151, N13803, N1059);
nor NOR2 (N14809, N14790, N5427);
nor NOR3 (N14810, N14806, N7839, N4620);
and AND2 (N14811, N14809, N8345);
and AND2 (N14812, N14792, N2395);
and AND4 (N14813, N14810, N4963, N762, N9623);
nand NAND4 (N14814, N14773, N14698, N1485, N11025);
not NOT1 (N14815, N14799);
nor NOR3 (N14816, N14815, N8215, N6573);
nand NAND3 (N14817, N14814, N1391, N9284);
or OR2 (N14818, N14807, N7989);
buf BUF1 (N14819, N14803);
not NOT1 (N14820, N14813);
nand NAND3 (N14821, N14816, N7265, N10609);
and AND2 (N14822, N14812, N3068);
not NOT1 (N14823, N14817);
nor NOR4 (N14824, N14820, N1198, N247, N6738);
not NOT1 (N14825, N14819);
or OR4 (N14826, N14824, N11827, N12632, N594);
nand NAND4 (N14827, N14802, N1288, N13705, N8357);
not NOT1 (N14828, N14821);
nor NOR4 (N14829, N14808, N7611, N13177, N13849);
and AND4 (N14830, N14823, N5297, N13596, N10474);
not NOT1 (N14831, N14822);
xor XOR2 (N14832, N14825, N11003);
or OR4 (N14833, N14818, N8828, N5527, N1934);
not NOT1 (N14834, N14828);
buf BUF1 (N14835, N14831);
nand NAND4 (N14836, N14833, N5063, N5758, N6405);
not NOT1 (N14837, N14830);
nand NAND3 (N14838, N14835, N4780, N10726);
and AND3 (N14839, N14836, N5586, N2306);
not NOT1 (N14840, N14837);
and AND2 (N14841, N14832, N9161);
not NOT1 (N14842, N14838);
xor XOR2 (N14843, N14839, N6569);
not NOT1 (N14844, N14840);
xor XOR2 (N14845, N14800, N2547);
not NOT1 (N14846, N14845);
not NOT1 (N14847, N14827);
not NOT1 (N14848, N14846);
and AND3 (N14849, N14842, N5687, N5183);
not NOT1 (N14850, N14826);
nor NOR3 (N14851, N14849, N4734, N8550);
xor XOR2 (N14852, N14829, N3709);
or OR3 (N14853, N14850, N5106, N4974);
not NOT1 (N14854, N14853);
not NOT1 (N14855, N14843);
nor NOR3 (N14856, N14841, N12316, N12385);
or OR3 (N14857, N14811, N12093, N10837);
not NOT1 (N14858, N14852);
xor XOR2 (N14859, N14844, N13368);
xor XOR2 (N14860, N14834, N13133);
nor NOR3 (N14861, N14856, N13988, N3481);
or OR2 (N14862, N14857, N10142);
and AND2 (N14863, N14854, N5818);
nand NAND3 (N14864, N14848, N2552, N13740);
not NOT1 (N14865, N14847);
xor XOR2 (N14866, N14858, N10503);
nor NOR4 (N14867, N14851, N278, N1264, N4152);
and AND4 (N14868, N14862, N9790, N7565, N6962);
and AND2 (N14869, N14864, N13096);
buf BUF1 (N14870, N14868);
and AND4 (N14871, N14866, N8293, N952, N4578);
xor XOR2 (N14872, N14870, N2097);
not NOT1 (N14873, N14865);
xor XOR2 (N14874, N14871, N8830);
nor NOR3 (N14875, N14873, N1790, N6239);
nand NAND2 (N14876, N14863, N6650);
and AND4 (N14877, N14869, N10402, N12922, N4056);
nand NAND2 (N14878, N14877, N8832);
not NOT1 (N14879, N14860);
not NOT1 (N14880, N14872);
xor XOR2 (N14881, N14879, N2894);
or OR2 (N14882, N14876, N5073);
and AND4 (N14883, N14882, N10167, N14108, N8062);
nand NAND3 (N14884, N14859, N9076, N523);
not NOT1 (N14885, N14881);
xor XOR2 (N14886, N14875, N12475);
buf BUF1 (N14887, N14861);
or OR4 (N14888, N14855, N4720, N8209, N8090);
xor XOR2 (N14889, N14885, N35);
nand NAND3 (N14890, N14887, N8173, N6999);
xor XOR2 (N14891, N14880, N1978);
not NOT1 (N14892, N14883);
not NOT1 (N14893, N14878);
nor NOR2 (N14894, N14888, N7368);
not NOT1 (N14895, N14889);
nor NOR4 (N14896, N14891, N2979, N8962, N10174);
not NOT1 (N14897, N14893);
nor NOR4 (N14898, N14874, N12457, N2849, N13070);
and AND2 (N14899, N14886, N573);
not NOT1 (N14900, N14897);
and AND3 (N14901, N14896, N6130, N10254);
buf BUF1 (N14902, N14895);
xor XOR2 (N14903, N14884, N5219);
nor NOR3 (N14904, N14890, N51, N13418);
not NOT1 (N14905, N14901);
buf BUF1 (N14906, N14867);
nand NAND4 (N14907, N14898, N12239, N9443, N12073);
or OR4 (N14908, N14903, N11617, N4019, N4591);
not NOT1 (N14909, N14892);
xor XOR2 (N14910, N14909, N9751);
xor XOR2 (N14911, N14905, N7940);
nand NAND2 (N14912, N14907, N11561);
nor NOR3 (N14913, N14902, N6892, N10478);
buf BUF1 (N14914, N14900);
not NOT1 (N14915, N14894);
xor XOR2 (N14916, N14904, N6986);
nand NAND2 (N14917, N14915, N4338);
buf BUF1 (N14918, N14917);
nor NOR4 (N14919, N14908, N10094, N3659, N10519);
buf BUF1 (N14920, N14910);
nand NAND4 (N14921, N14919, N5774, N12503, N10462);
not NOT1 (N14922, N14911);
and AND4 (N14923, N14912, N9562, N12697, N12842);
or OR3 (N14924, N14922, N10686, N2778);
buf BUF1 (N14925, N14924);
buf BUF1 (N14926, N14920);
and AND2 (N14927, N14918, N10610);
not NOT1 (N14928, N14927);
or OR2 (N14929, N14928, N8999);
not NOT1 (N14930, N14925);
not NOT1 (N14931, N14913);
and AND2 (N14932, N14899, N5464);
nand NAND3 (N14933, N14916, N5140, N8486);
nand NAND2 (N14934, N14926, N3472);
buf BUF1 (N14935, N14906);
not NOT1 (N14936, N14934);
nor NOR2 (N14937, N14930, N4346);
nor NOR2 (N14938, N14931, N8056);
buf BUF1 (N14939, N14914);
nor NOR3 (N14940, N14921, N7538, N13701);
not NOT1 (N14941, N14923);
and AND2 (N14942, N14938, N1941);
nor NOR2 (N14943, N14932, N13111);
nand NAND4 (N14944, N14940, N9737, N13165, N1157);
not NOT1 (N14945, N14933);
xor XOR2 (N14946, N14935, N9886);
xor XOR2 (N14947, N14943, N4940);
not NOT1 (N14948, N14936);
and AND2 (N14949, N14941, N6756);
or OR3 (N14950, N14947, N5861, N13483);
buf BUF1 (N14951, N14950);
buf BUF1 (N14952, N14942);
or OR4 (N14953, N14948, N6791, N6957, N2687);
nand NAND3 (N14954, N14951, N3633, N11644);
xor XOR2 (N14955, N14949, N9693);
and AND3 (N14956, N14946, N13612, N10079);
and AND2 (N14957, N14953, N7223);
nor NOR3 (N14958, N14929, N6633, N6389);
and AND3 (N14959, N14939, N14700, N3929);
nand NAND2 (N14960, N14945, N9941);
nand NAND3 (N14961, N14957, N1629, N12545);
or OR3 (N14962, N14959, N3916, N13841);
not NOT1 (N14963, N14961);
nor NOR3 (N14964, N14958, N8857, N2629);
nand NAND3 (N14965, N14964, N13566, N9734);
nor NOR4 (N14966, N14944, N8078, N5581, N1435);
buf BUF1 (N14967, N14965);
buf BUF1 (N14968, N14967);
buf BUF1 (N14969, N14962);
nand NAND2 (N14970, N14969, N895);
xor XOR2 (N14971, N14968, N12159);
not NOT1 (N14972, N14956);
buf BUF1 (N14973, N14954);
or OR4 (N14974, N14972, N13023, N6279, N5572);
nor NOR3 (N14975, N14970, N1689, N11347);
nor NOR3 (N14976, N14974, N6277, N11020);
nand NAND4 (N14977, N14976, N12836, N2846, N8930);
xor XOR2 (N14978, N14966, N4033);
buf BUF1 (N14979, N14960);
or OR2 (N14980, N14973, N5221);
xor XOR2 (N14981, N14979, N6896);
nor NOR4 (N14982, N14963, N3562, N9845, N5191);
xor XOR2 (N14983, N14955, N8410);
or OR2 (N14984, N14975, N8193);
buf BUF1 (N14985, N14978);
xor XOR2 (N14986, N14952, N2482);
not NOT1 (N14987, N14986);
not NOT1 (N14988, N14987);
nand NAND4 (N14989, N14985, N483, N4559, N1783);
xor XOR2 (N14990, N14989, N5612);
not NOT1 (N14991, N14977);
and AND3 (N14992, N14991, N758, N12181);
and AND2 (N14993, N14990, N7109);
or OR4 (N14994, N14983, N448, N2398, N455);
buf BUF1 (N14995, N14981);
nor NOR2 (N14996, N14992, N7507);
or OR3 (N14997, N14937, N8467, N2759);
xor XOR2 (N14998, N14993, N13548);
nand NAND2 (N14999, N14995, N9404);
or OR3 (N15000, N14980, N3503, N1448);
nor NOR4 (N15001, N15000, N7644, N6487, N6543);
nand NAND4 (N15002, N14999, N9444, N11628, N14002);
or OR4 (N15003, N14997, N9063, N9893, N7118);
not NOT1 (N15004, N14998);
and AND2 (N15005, N14994, N2882);
nor NOR2 (N15006, N15002, N14568);
nor NOR3 (N15007, N14996, N9700, N12743);
xor XOR2 (N15008, N14988, N14061);
not NOT1 (N15009, N15004);
not NOT1 (N15010, N15009);
not NOT1 (N15011, N15006);
nand NAND2 (N15012, N15011, N13734);
xor XOR2 (N15013, N15008, N7290);
and AND3 (N15014, N14984, N10675, N7370);
and AND4 (N15015, N15005, N586, N12262, N4976);
xor XOR2 (N15016, N14982, N5431);
and AND2 (N15017, N15010, N1932);
xor XOR2 (N15018, N15017, N2450);
buf BUF1 (N15019, N15014);
and AND4 (N15020, N15015, N14, N1166, N11787);
and AND2 (N15021, N15013, N4533);
buf BUF1 (N15022, N15019);
buf BUF1 (N15023, N15001);
or OR3 (N15024, N15021, N5173, N3065);
buf BUF1 (N15025, N15018);
xor XOR2 (N15026, N15024, N2282);
or OR4 (N15027, N15020, N9536, N12785, N495);
or OR4 (N15028, N15016, N180, N5413, N5950);
or OR3 (N15029, N15012, N3301, N5356);
xor XOR2 (N15030, N15026, N9900);
not NOT1 (N15031, N15029);
buf BUF1 (N15032, N15022);
and AND3 (N15033, N15027, N2685, N12183);
xor XOR2 (N15034, N15028, N9694);
buf BUF1 (N15035, N15007);
nor NOR4 (N15036, N15034, N1814, N12281, N10256);
nand NAND4 (N15037, N15030, N4526, N3853, N10824);
xor XOR2 (N15038, N15033, N14784);
not NOT1 (N15039, N15031);
buf BUF1 (N15040, N15037);
buf BUF1 (N15041, N15003);
xor XOR2 (N15042, N15039, N12575);
and AND4 (N15043, N15040, N10025, N14565, N5831);
xor XOR2 (N15044, N15038, N4093);
or OR4 (N15045, N15023, N5098, N13939, N5738);
not NOT1 (N15046, N15032);
buf BUF1 (N15047, N15044);
or OR2 (N15048, N15047, N10613);
nor NOR3 (N15049, N15045, N14451, N8497);
and AND3 (N15050, N15049, N9450, N5439);
nor NOR4 (N15051, N15041, N5233, N991, N6554);
and AND3 (N15052, N15051, N5584, N4536);
xor XOR2 (N15053, N15050, N6323);
xor XOR2 (N15054, N15035, N8972);
and AND3 (N15055, N15048, N574, N3987);
buf BUF1 (N15056, N15052);
buf BUF1 (N15057, N15056);
and AND4 (N15058, N15046, N399, N6468, N7208);
or OR2 (N15059, N15057, N10286);
and AND3 (N15060, N15053, N13463, N1355);
and AND3 (N15061, N14971, N12880, N3726);
or OR3 (N15062, N15043, N9214, N4139);
xor XOR2 (N15063, N15036, N13889);
nand NAND4 (N15064, N15063, N5345, N14738, N11724);
nor NOR4 (N15065, N15062, N9706, N5723, N11301);
not NOT1 (N15066, N15025);
and AND2 (N15067, N15061, N8691);
or OR2 (N15068, N15060, N7467);
nor NOR2 (N15069, N15065, N11845);
nor NOR3 (N15070, N15058, N621, N12584);
not NOT1 (N15071, N15042);
nor NOR2 (N15072, N15055, N1082);
not NOT1 (N15073, N15066);
xor XOR2 (N15074, N15054, N11824);
or OR4 (N15075, N15069, N2588, N9084, N6361);
nand NAND3 (N15076, N15074, N1149, N13452);
nor NOR3 (N15077, N15076, N6260, N4231);
not NOT1 (N15078, N15064);
nor NOR3 (N15079, N15078, N7051, N2649);
not NOT1 (N15080, N15077);
nand NAND3 (N15081, N15079, N10274, N14787);
not NOT1 (N15082, N15081);
and AND3 (N15083, N15059, N2946, N3913);
not NOT1 (N15084, N15073);
nor NOR3 (N15085, N15072, N301, N3309);
xor XOR2 (N15086, N15068, N7407);
xor XOR2 (N15087, N15070, N6921);
and AND3 (N15088, N15067, N9804, N5541);
not NOT1 (N15089, N15087);
and AND4 (N15090, N15082, N14365, N12012, N1175);
nor NOR4 (N15091, N15089, N1794, N8725, N317);
nand NAND4 (N15092, N15075, N4298, N12647, N9331);
buf BUF1 (N15093, N15092);
buf BUF1 (N15094, N15091);
nand NAND2 (N15095, N15093, N14103);
nor NOR4 (N15096, N15090, N2472, N10780, N13230);
xor XOR2 (N15097, N15086, N3456);
or OR2 (N15098, N15096, N4654);
or OR4 (N15099, N15098, N11030, N11830, N15092);
and AND4 (N15100, N15095, N12072, N1005, N130);
xor XOR2 (N15101, N15088, N793);
or OR2 (N15102, N15084, N15040);
nor NOR2 (N15103, N15071, N3965);
buf BUF1 (N15104, N15080);
buf BUF1 (N15105, N15097);
and AND3 (N15106, N15099, N7043, N3980);
nor NOR4 (N15107, N15102, N14785, N741, N1808);
not NOT1 (N15108, N15105);
xor XOR2 (N15109, N15100, N939);
not NOT1 (N15110, N15101);
xor XOR2 (N15111, N15083, N12675);
buf BUF1 (N15112, N15108);
not NOT1 (N15113, N15109);
not NOT1 (N15114, N15085);
not NOT1 (N15115, N15103);
nand NAND2 (N15116, N15111, N11778);
nor NOR4 (N15117, N15094, N2639, N11125, N2662);
nand NAND4 (N15118, N15107, N14502, N2273, N3640);
nand NAND4 (N15119, N15116, N11340, N1803, N7950);
and AND4 (N15120, N15106, N14435, N1259, N2178);
or OR4 (N15121, N15115, N7976, N2034, N3811);
or OR3 (N15122, N15119, N1347, N2958);
buf BUF1 (N15123, N15121);
not NOT1 (N15124, N15113);
xor XOR2 (N15125, N15114, N12720);
not NOT1 (N15126, N15110);
not NOT1 (N15127, N15122);
xor XOR2 (N15128, N15118, N9632);
or OR4 (N15129, N15104, N5731, N1763, N5027);
nor NOR3 (N15130, N15128, N4656, N4623);
xor XOR2 (N15131, N15129, N10177);
buf BUF1 (N15132, N15120);
nand NAND4 (N15133, N15126, N3623, N10595, N1626);
xor XOR2 (N15134, N15130, N3250);
buf BUF1 (N15135, N15131);
nand NAND2 (N15136, N15117, N3348);
not NOT1 (N15137, N15133);
buf BUF1 (N15138, N15125);
nor NOR4 (N15139, N15138, N6898, N4534, N2376);
buf BUF1 (N15140, N15137);
or OR4 (N15141, N15134, N1990, N12723, N6375);
nand NAND4 (N15142, N15112, N10013, N6295, N12264);
xor XOR2 (N15143, N15127, N10318);
xor XOR2 (N15144, N15132, N1631);
or OR2 (N15145, N15142, N6753);
or OR2 (N15146, N15145, N8983);
xor XOR2 (N15147, N15141, N12303);
xor XOR2 (N15148, N15139, N10414);
nand NAND4 (N15149, N15146, N6236, N14471, N8187);
buf BUF1 (N15150, N15123);
or OR3 (N15151, N15150, N2672, N855);
nor NOR2 (N15152, N15148, N5316);
not NOT1 (N15153, N15144);
or OR4 (N15154, N15136, N12841, N10857, N11635);
and AND2 (N15155, N15143, N13074);
nand NAND4 (N15156, N15140, N1438, N11069, N12534);
or OR2 (N15157, N15149, N11507);
nor NOR3 (N15158, N15152, N4172, N9231);
or OR4 (N15159, N15135, N2472, N10245, N14459);
and AND4 (N15160, N15124, N8796, N11892, N350);
and AND2 (N15161, N15158, N5871);
xor XOR2 (N15162, N15157, N1810);
not NOT1 (N15163, N15147);
not NOT1 (N15164, N15151);
buf BUF1 (N15165, N15155);
or OR4 (N15166, N15154, N10285, N2979, N14684);
not NOT1 (N15167, N15166);
and AND3 (N15168, N15162, N4387, N12928);
nand NAND2 (N15169, N15165, N6458);
and AND2 (N15170, N15164, N14046);
xor XOR2 (N15171, N15161, N3016);
nor NOR2 (N15172, N15167, N1154);
buf BUF1 (N15173, N15153);
and AND3 (N15174, N15156, N14877, N14152);
and AND2 (N15175, N15163, N4346);
and AND4 (N15176, N15169, N13578, N8755, N3905);
buf BUF1 (N15177, N15159);
buf BUF1 (N15178, N15168);
and AND2 (N15179, N15170, N14007);
and AND4 (N15180, N15178, N5842, N6451, N10138);
not NOT1 (N15181, N15160);
nor NOR3 (N15182, N15180, N5076, N11501);
not NOT1 (N15183, N15171);
or OR4 (N15184, N15172, N4329, N7250, N6721);
and AND3 (N15185, N15183, N9312, N7047);
xor XOR2 (N15186, N15175, N3963);
buf BUF1 (N15187, N15179);
nand NAND3 (N15188, N15181, N434, N8928);
not NOT1 (N15189, N15173);
buf BUF1 (N15190, N15174);
xor XOR2 (N15191, N15190, N10679);
and AND4 (N15192, N15177, N3604, N359, N3428);
xor XOR2 (N15193, N15191, N1067);
or OR4 (N15194, N15186, N4224, N8675, N12870);
and AND2 (N15195, N15194, N1556);
xor XOR2 (N15196, N15184, N14859);
nor NOR4 (N15197, N15195, N2974, N14207, N9900);
nand NAND2 (N15198, N15182, N10504);
and AND2 (N15199, N15188, N8280);
or OR3 (N15200, N15196, N10718, N8033);
not NOT1 (N15201, N15185);
nand NAND2 (N15202, N15198, N3523);
xor XOR2 (N15203, N15192, N4037);
nor NOR4 (N15204, N15200, N8125, N5778, N8218);
nand NAND3 (N15205, N15189, N9229, N12981);
not NOT1 (N15206, N15204);
nand NAND2 (N15207, N15197, N6161);
not NOT1 (N15208, N15207);
or OR2 (N15209, N15208, N13599);
buf BUF1 (N15210, N15193);
and AND4 (N15211, N15203, N8655, N10612, N6131);
nand NAND2 (N15212, N15209, N2334);
nor NOR3 (N15213, N15199, N3522, N555);
xor XOR2 (N15214, N15187, N12432);
not NOT1 (N15215, N15205);
xor XOR2 (N15216, N15211, N12983);
xor XOR2 (N15217, N15176, N14615);
or OR4 (N15218, N15215, N11527, N3115, N4439);
nor NOR4 (N15219, N15212, N11883, N4981, N14290);
or OR4 (N15220, N15213, N4529, N6208, N12658);
and AND3 (N15221, N15206, N1812, N3663);
nand NAND3 (N15222, N15221, N932, N1115);
nor NOR3 (N15223, N15219, N7758, N10283);
or OR4 (N15224, N15201, N8410, N5227, N3651);
xor XOR2 (N15225, N15214, N6568);
nor NOR2 (N15226, N15222, N1780);
nor NOR3 (N15227, N15220, N11841, N1186);
and AND4 (N15228, N15227, N3431, N6349, N8980);
nand NAND3 (N15229, N15202, N7064, N13999);
or OR2 (N15230, N15224, N3258);
buf BUF1 (N15231, N15217);
buf BUF1 (N15232, N15223);
not NOT1 (N15233, N15230);
buf BUF1 (N15234, N15210);
or OR3 (N15235, N15216, N13142, N4084);
buf BUF1 (N15236, N15231);
and AND3 (N15237, N15226, N4459, N10857);
or OR3 (N15238, N15237, N2738, N2502);
nand NAND2 (N15239, N15232, N13146);
buf BUF1 (N15240, N15218);
nor NOR4 (N15241, N15228, N1947, N14220, N5127);
and AND3 (N15242, N15240, N8228, N9641);
and AND4 (N15243, N15225, N14027, N277, N4734);
buf BUF1 (N15244, N15233);
or OR4 (N15245, N15239, N13544, N739, N14174);
xor XOR2 (N15246, N15245, N12742);
xor XOR2 (N15247, N15234, N12440);
and AND4 (N15248, N15247, N13578, N13154, N14380);
or OR4 (N15249, N15243, N13351, N657, N1201);
and AND4 (N15250, N15235, N3235, N10664, N1576);
and AND2 (N15251, N15241, N3430);
and AND3 (N15252, N15244, N5918, N14054);
nor NOR2 (N15253, N15238, N10950);
and AND3 (N15254, N15253, N3316, N5684);
buf BUF1 (N15255, N15236);
or OR2 (N15256, N15229, N14232);
and AND3 (N15257, N15256, N5998, N8157);
xor XOR2 (N15258, N15251, N3425);
not NOT1 (N15259, N15246);
buf BUF1 (N15260, N15257);
not NOT1 (N15261, N15250);
nand NAND3 (N15262, N15249, N1784, N2440);
or OR2 (N15263, N15255, N6908);
buf BUF1 (N15264, N15254);
xor XOR2 (N15265, N15252, N2549);
or OR2 (N15266, N15260, N9321);
buf BUF1 (N15267, N15248);
xor XOR2 (N15268, N15261, N9375);
or OR2 (N15269, N15266, N12066);
not NOT1 (N15270, N15267);
nor NOR2 (N15271, N15268, N4075);
or OR3 (N15272, N15242, N1656, N3427);
buf BUF1 (N15273, N15272);
nor NOR2 (N15274, N15262, N9537);
xor XOR2 (N15275, N15265, N8283);
not NOT1 (N15276, N15273);
or OR3 (N15277, N15258, N12732, N3999);
nor NOR4 (N15278, N15259, N11791, N8737, N6888);
xor XOR2 (N15279, N15276, N9573);
and AND4 (N15280, N15274, N12786, N1926, N5589);
xor XOR2 (N15281, N15277, N2219);
buf BUF1 (N15282, N15263);
and AND3 (N15283, N15278, N15087, N1042);
or OR2 (N15284, N15282, N14908);
and AND4 (N15285, N15280, N11438, N14497, N13603);
buf BUF1 (N15286, N15283);
buf BUF1 (N15287, N15270);
xor XOR2 (N15288, N15286, N2851);
and AND4 (N15289, N15279, N11080, N14574, N186);
and AND4 (N15290, N15275, N7155, N5896, N10677);
nand NAND4 (N15291, N15289, N3938, N1316, N8266);
not NOT1 (N15292, N15288);
nand NAND2 (N15293, N15269, N3263);
nand NAND4 (N15294, N15264, N876, N3520, N10384);
nor NOR4 (N15295, N15285, N8017, N8046, N7743);
or OR2 (N15296, N15281, N10319);
buf BUF1 (N15297, N15287);
nor NOR3 (N15298, N15294, N1146, N3704);
nor NOR4 (N15299, N15290, N11502, N9667, N14176);
nor NOR2 (N15300, N15292, N6506);
nor NOR2 (N15301, N15295, N6001);
buf BUF1 (N15302, N15297);
xor XOR2 (N15303, N15271, N13865);
not NOT1 (N15304, N15296);
buf BUF1 (N15305, N15291);
nand NAND3 (N15306, N15298, N1565, N5248);
and AND2 (N15307, N15301, N13457);
and AND2 (N15308, N15303, N2926);
and AND4 (N15309, N15305, N1699, N2219, N4920);
nor NOR2 (N15310, N15302, N8585);
or OR2 (N15311, N15308, N10461);
nor NOR4 (N15312, N15284, N14140, N6128, N5655);
xor XOR2 (N15313, N15311, N13649);
xor XOR2 (N15314, N15312, N3446);
xor XOR2 (N15315, N15310, N3794);
nand NAND2 (N15316, N15307, N12343);
nor NOR2 (N15317, N15314, N3984);
buf BUF1 (N15318, N15299);
buf BUF1 (N15319, N15304);
nor NOR2 (N15320, N15293, N624);
xor XOR2 (N15321, N15317, N5344);
buf BUF1 (N15322, N15316);
and AND4 (N15323, N15306, N1221, N6511, N12017);
not NOT1 (N15324, N15319);
nand NAND4 (N15325, N15323, N8272, N4373, N15316);
buf BUF1 (N15326, N15322);
and AND3 (N15327, N15320, N1356, N8171);
or OR3 (N15328, N15324, N12042, N7707);
or OR3 (N15329, N15300, N12927, N11089);
xor XOR2 (N15330, N15326, N10467);
buf BUF1 (N15331, N15318);
buf BUF1 (N15332, N15313);
nor NOR2 (N15333, N15309, N12766);
and AND2 (N15334, N15331, N1878);
buf BUF1 (N15335, N15333);
not NOT1 (N15336, N15325);
and AND3 (N15337, N15329, N11718, N4854);
buf BUF1 (N15338, N15315);
not NOT1 (N15339, N15321);
nand NAND3 (N15340, N15336, N6789, N2090);
and AND2 (N15341, N15327, N14908);
nor NOR3 (N15342, N15341, N175, N5323);
xor XOR2 (N15343, N15338, N14078);
not NOT1 (N15344, N15328);
xor XOR2 (N15345, N15334, N6476);
and AND4 (N15346, N15343, N12778, N11306, N7866);
xor XOR2 (N15347, N15344, N8013);
nand NAND3 (N15348, N15337, N2450, N5611);
or OR4 (N15349, N15346, N7332, N11447, N8415);
buf BUF1 (N15350, N15348);
or OR2 (N15351, N15335, N6049);
and AND4 (N15352, N15350, N8140, N7539, N13425);
buf BUF1 (N15353, N15351);
nor NOR4 (N15354, N15330, N14034, N13953, N6760);
not NOT1 (N15355, N15340);
nor NOR2 (N15356, N15339, N2996);
or OR2 (N15357, N15354, N13806);
buf BUF1 (N15358, N15342);
nand NAND4 (N15359, N15332, N4716, N13093, N11937);
not NOT1 (N15360, N15355);
nor NOR3 (N15361, N15360, N1120, N11950);
not NOT1 (N15362, N15347);
nor NOR3 (N15363, N15349, N3448, N12316);
and AND3 (N15364, N15359, N5743, N12070);
nor NOR2 (N15365, N15358, N12638);
not NOT1 (N15366, N15345);
and AND4 (N15367, N15356, N10245, N2554, N11204);
not NOT1 (N15368, N15357);
nand NAND4 (N15369, N15368, N1484, N4754, N3924);
not NOT1 (N15370, N15362);
and AND4 (N15371, N15364, N1101, N465, N5619);
or OR2 (N15372, N15365, N10401);
not NOT1 (N15373, N15366);
not NOT1 (N15374, N15367);
nor NOR3 (N15375, N15352, N11917, N6377);
nor NOR3 (N15376, N15373, N7109, N2140);
not NOT1 (N15377, N15372);
or OR2 (N15378, N15353, N12382);
xor XOR2 (N15379, N15371, N10707);
and AND4 (N15380, N15376, N9954, N29, N8067);
xor XOR2 (N15381, N15374, N9615);
buf BUF1 (N15382, N15378);
and AND3 (N15383, N15380, N751, N12848);
buf BUF1 (N15384, N15382);
not NOT1 (N15385, N15377);
nor NOR2 (N15386, N15363, N11933);
nand NAND3 (N15387, N15370, N7927, N11913);
not NOT1 (N15388, N15384);
buf BUF1 (N15389, N15361);
nor NOR2 (N15390, N15375, N9983);
buf BUF1 (N15391, N15385);
nor NOR2 (N15392, N15386, N5668);
and AND2 (N15393, N15388, N4235);
or OR2 (N15394, N15369, N15058);
nand NAND2 (N15395, N15387, N5758);
or OR3 (N15396, N15389, N5344, N2937);
buf BUF1 (N15397, N15394);
xor XOR2 (N15398, N15379, N11501);
or OR3 (N15399, N15396, N13641, N10066);
not NOT1 (N15400, N15383);
or OR4 (N15401, N15391, N3951, N12791, N11225);
buf BUF1 (N15402, N15399);
not NOT1 (N15403, N15392);
xor XOR2 (N15404, N15390, N5345);
nand NAND3 (N15405, N15398, N2895, N14042);
or OR3 (N15406, N15403, N7215, N13663);
or OR2 (N15407, N15401, N2276);
not NOT1 (N15408, N15400);
and AND2 (N15409, N15404, N5820);
buf BUF1 (N15410, N15393);
not NOT1 (N15411, N15397);
and AND3 (N15412, N15410, N12927, N13164);
not NOT1 (N15413, N15406);
nand NAND3 (N15414, N15405, N15272, N13655);
not NOT1 (N15415, N15414);
nor NOR4 (N15416, N15415, N12085, N435, N11501);
buf BUF1 (N15417, N15411);
nor NOR4 (N15418, N15408, N1030, N8824, N7057);
nor NOR4 (N15419, N15412, N7049, N9760, N14985);
and AND4 (N15420, N15395, N12197, N12269, N6842);
xor XOR2 (N15421, N15407, N4918);
not NOT1 (N15422, N15419);
nor NOR4 (N15423, N15402, N14121, N579, N12373);
xor XOR2 (N15424, N15409, N137);
nand NAND4 (N15425, N15381, N6062, N11695, N3431);
nor NOR4 (N15426, N15417, N11872, N12983, N1424);
not NOT1 (N15427, N15420);
not NOT1 (N15428, N15427);
nor NOR2 (N15429, N15413, N2788);
buf BUF1 (N15430, N15424);
nand NAND2 (N15431, N15423, N6276);
xor XOR2 (N15432, N15430, N379);
and AND3 (N15433, N15425, N8071, N3147);
nor NOR2 (N15434, N15421, N14253);
not NOT1 (N15435, N15432);
xor XOR2 (N15436, N15418, N12200);
or OR3 (N15437, N15429, N2784, N3666);
not NOT1 (N15438, N15416);
nor NOR2 (N15439, N15431, N9801);
xor XOR2 (N15440, N15435, N12531);
nand NAND3 (N15441, N15422, N7714, N10892);
buf BUF1 (N15442, N15428);
buf BUF1 (N15443, N15441);
xor XOR2 (N15444, N15443, N12801);
and AND3 (N15445, N15444, N1798, N9717);
nor NOR3 (N15446, N15440, N3397, N83);
or OR4 (N15447, N15433, N3881, N14146, N14234);
buf BUF1 (N15448, N15437);
and AND3 (N15449, N15426, N1545, N8548);
not NOT1 (N15450, N15434);
not NOT1 (N15451, N15445);
nor NOR2 (N15452, N15442, N12347);
nor NOR3 (N15453, N15452, N5597, N1439);
or OR4 (N15454, N15448, N7354, N14671, N5124);
xor XOR2 (N15455, N15436, N11628);
nor NOR3 (N15456, N15453, N3712, N2670);
nor NOR3 (N15457, N15439, N2193, N972);
or OR2 (N15458, N15446, N11230);
and AND3 (N15459, N15455, N12891, N2993);
buf BUF1 (N15460, N15449);
xor XOR2 (N15461, N15450, N10060);
xor XOR2 (N15462, N15438, N15032);
xor XOR2 (N15463, N15454, N6702);
and AND3 (N15464, N15451, N213, N2219);
and AND4 (N15465, N15447, N776, N5348, N14309);
xor XOR2 (N15466, N15461, N4889);
and AND3 (N15467, N15466, N8449, N327);
not NOT1 (N15468, N15467);
and AND2 (N15469, N15462, N1113);
xor XOR2 (N15470, N15458, N10103);
or OR4 (N15471, N15470, N847, N6715, N7663);
nor NOR4 (N15472, N15456, N3759, N2251, N3584);
xor XOR2 (N15473, N15465, N8526);
and AND3 (N15474, N15469, N11253, N11986);
buf BUF1 (N15475, N15474);
or OR4 (N15476, N15468, N4879, N8657, N11695);
nor NOR3 (N15477, N15475, N13233, N10811);
nand NAND2 (N15478, N15457, N6642);
buf BUF1 (N15479, N15473);
xor XOR2 (N15480, N15459, N14417);
xor XOR2 (N15481, N15478, N12137);
nand NAND4 (N15482, N15477, N13007, N5674, N12822);
nand NAND4 (N15483, N15480, N13641, N2917, N13684);
nor NOR3 (N15484, N15472, N3122, N14899);
or OR4 (N15485, N15481, N4489, N13213, N12323);
buf BUF1 (N15486, N15483);
or OR3 (N15487, N15484, N4430, N2673);
nand NAND4 (N15488, N15485, N6230, N897, N10353);
or OR2 (N15489, N15460, N12288);
nand NAND4 (N15490, N15476, N14192, N10111, N571);
nand NAND3 (N15491, N15487, N10169, N5958);
and AND2 (N15492, N15463, N4345);
and AND3 (N15493, N15492, N9617, N8471);
xor XOR2 (N15494, N15491, N6939);
or OR4 (N15495, N15479, N1603, N1035, N8410);
xor XOR2 (N15496, N15495, N1108);
or OR3 (N15497, N15486, N13631, N6588);
or OR2 (N15498, N15496, N15142);
buf BUF1 (N15499, N15488);
nand NAND2 (N15500, N15493, N11103);
buf BUF1 (N15501, N15471);
or OR2 (N15502, N15489, N1068);
not NOT1 (N15503, N15464);
and AND3 (N15504, N15499, N4449, N174);
buf BUF1 (N15505, N15497);
nor NOR3 (N15506, N15501, N6412, N4838);
nand NAND3 (N15507, N15498, N2330, N11297);
xor XOR2 (N15508, N15506, N10971);
xor XOR2 (N15509, N15490, N11144);
nand NAND3 (N15510, N15504, N13835, N12950);
nand NAND4 (N15511, N15482, N7959, N5279, N6503);
and AND3 (N15512, N15502, N1694, N11371);
nand NAND4 (N15513, N15507, N3518, N3430, N1901);
xor XOR2 (N15514, N15509, N126);
or OR4 (N15515, N15512, N14026, N5351, N267);
buf BUF1 (N15516, N15513);
or OR3 (N15517, N15510, N168, N8690);
nor NOR3 (N15518, N15500, N10781, N239);
not NOT1 (N15519, N15514);
and AND2 (N15520, N15503, N3145);
or OR3 (N15521, N15516, N12288, N937);
nand NAND4 (N15522, N15521, N13724, N4378, N1393);
not NOT1 (N15523, N15505);
or OR4 (N15524, N15519, N11662, N14437, N11404);
or OR2 (N15525, N15511, N7249);
and AND3 (N15526, N15517, N8345, N5678);
or OR2 (N15527, N15524, N4042);
nor NOR2 (N15528, N15527, N11677);
or OR4 (N15529, N15515, N14818, N11447, N7723);
xor XOR2 (N15530, N15494, N1861);
nand NAND4 (N15531, N15529, N7446, N2168, N10204);
not NOT1 (N15532, N15520);
or OR4 (N15533, N15531, N2830, N6414, N533);
not NOT1 (N15534, N15518);
xor XOR2 (N15535, N15525, N7445);
and AND2 (N15536, N15530, N10162);
nor NOR4 (N15537, N15533, N10106, N7522, N7078);
nor NOR2 (N15538, N15522, N14570);
not NOT1 (N15539, N15526);
not NOT1 (N15540, N15532);
not NOT1 (N15541, N15536);
or OR2 (N15542, N15538, N2674);
or OR4 (N15543, N15539, N2116, N10762, N14031);
or OR4 (N15544, N15541, N7030, N10089, N14340);
not NOT1 (N15545, N15523);
xor XOR2 (N15546, N15534, N1006);
not NOT1 (N15547, N15537);
buf BUF1 (N15548, N15528);
nor NOR3 (N15549, N15508, N197, N12860);
xor XOR2 (N15550, N15548, N12899);
or OR4 (N15551, N15546, N2200, N5725, N13439);
xor XOR2 (N15552, N15551, N9473);
xor XOR2 (N15553, N15550, N77);
buf BUF1 (N15554, N15549);
buf BUF1 (N15555, N15553);
nand NAND4 (N15556, N15543, N9022, N8572, N14784);
buf BUF1 (N15557, N15535);
or OR2 (N15558, N15556, N10656);
and AND4 (N15559, N15544, N5434, N980, N5425);
xor XOR2 (N15560, N15542, N11659);
and AND4 (N15561, N15554, N11510, N902, N15332);
buf BUF1 (N15562, N15555);
and AND4 (N15563, N15547, N266, N3715, N14852);
and AND2 (N15564, N15560, N6597);
xor XOR2 (N15565, N15561, N11258);
nor NOR3 (N15566, N15552, N14881, N3683);
and AND3 (N15567, N15563, N6141, N1755);
not NOT1 (N15568, N15565);
buf BUF1 (N15569, N15558);
nand NAND2 (N15570, N15564, N15496);
nor NOR4 (N15571, N15559, N3267, N1933, N9952);
and AND3 (N15572, N15569, N6588, N10024);
xor XOR2 (N15573, N15562, N2305);
or OR4 (N15574, N15557, N5849, N1212, N13475);
not NOT1 (N15575, N15574);
nand NAND4 (N15576, N15568, N2905, N7727, N3147);
or OR2 (N15577, N15566, N15037);
nand NAND2 (N15578, N15577, N5501);
nand NAND2 (N15579, N15540, N6281);
nor NOR3 (N15580, N15573, N11817, N11376);
nor NOR4 (N15581, N15576, N5476, N2716, N14641);
xor XOR2 (N15582, N15572, N14470);
nor NOR4 (N15583, N15578, N1429, N2807, N8472);
buf BUF1 (N15584, N15583);
xor XOR2 (N15585, N15567, N11847);
nand NAND4 (N15586, N15585, N10522, N6762, N2419);
nor NOR3 (N15587, N15582, N3743, N6628);
or OR4 (N15588, N15545, N4142, N5618, N8190);
buf BUF1 (N15589, N15586);
or OR4 (N15590, N15570, N11787, N10564, N12435);
xor XOR2 (N15591, N15589, N2182);
xor XOR2 (N15592, N15584, N797);
xor XOR2 (N15593, N15591, N11552);
buf BUF1 (N15594, N15579);
and AND3 (N15595, N15592, N6093, N10195);
buf BUF1 (N15596, N15593);
xor XOR2 (N15597, N15587, N15153);
xor XOR2 (N15598, N15571, N5621);
buf BUF1 (N15599, N15590);
nor NOR4 (N15600, N15599, N2799, N15402, N14611);
and AND4 (N15601, N15581, N5837, N7067, N9390);
or OR4 (N15602, N15595, N13859, N1934, N838);
nand NAND4 (N15603, N15600, N178, N4374, N2362);
buf BUF1 (N15604, N15594);
xor XOR2 (N15605, N15603, N9721);
and AND3 (N15606, N15602, N15038, N11836);
nor NOR4 (N15607, N15606, N5241, N3960, N703);
and AND2 (N15608, N15597, N11747);
nand NAND3 (N15609, N15575, N11920, N9299);
nor NOR3 (N15610, N15609, N11711, N14371);
nor NOR2 (N15611, N15605, N265);
or OR2 (N15612, N15610, N6466);
nand NAND3 (N15613, N15601, N1255, N7124);
xor XOR2 (N15614, N15612, N635);
nor NOR4 (N15615, N15580, N9813, N12581, N7483);
not NOT1 (N15616, N15596);
xor XOR2 (N15617, N15613, N11888);
or OR2 (N15618, N15607, N6808);
and AND4 (N15619, N15608, N10836, N14050, N6193);
and AND3 (N15620, N15618, N9726, N9938);
nand NAND3 (N15621, N15598, N7588, N11956);
not NOT1 (N15622, N15611);
or OR2 (N15623, N15620, N13850);
nand NAND2 (N15624, N15614, N7218);
or OR4 (N15625, N15604, N5700, N15461, N12733);
or OR3 (N15626, N15615, N1846, N9691);
buf BUF1 (N15627, N15617);
and AND2 (N15628, N15626, N10378);
nand NAND4 (N15629, N15628, N1942, N14901, N8178);
xor XOR2 (N15630, N15622, N6510);
or OR2 (N15631, N15630, N218);
and AND3 (N15632, N15627, N3787, N15112);
nor NOR2 (N15633, N15632, N4309);
nand NAND3 (N15634, N15588, N5303, N90);
buf BUF1 (N15635, N15619);
nand NAND4 (N15636, N15635, N10671, N3107, N12333);
nand NAND4 (N15637, N15625, N2985, N5064, N8284);
nor NOR2 (N15638, N15631, N7417);
not NOT1 (N15639, N15637);
or OR2 (N15640, N15633, N3235);
xor XOR2 (N15641, N15624, N7509);
xor XOR2 (N15642, N15640, N15328);
nand NAND2 (N15643, N15641, N3114);
or OR2 (N15644, N15629, N13286);
xor XOR2 (N15645, N15634, N13750);
buf BUF1 (N15646, N15621);
nand NAND4 (N15647, N15646, N7972, N6517, N9632);
or OR3 (N15648, N15623, N8669, N4959);
not NOT1 (N15649, N15636);
not NOT1 (N15650, N15638);
xor XOR2 (N15651, N15650, N1350);
nand NAND3 (N15652, N15648, N8861, N14285);
not NOT1 (N15653, N15643);
not NOT1 (N15654, N15649);
nor NOR3 (N15655, N15653, N8361, N11317);
nor NOR3 (N15656, N15616, N6215, N12882);
not NOT1 (N15657, N15652);
or OR3 (N15658, N15651, N6007, N6386);
and AND2 (N15659, N15654, N5002);
not NOT1 (N15660, N15659);
nand NAND3 (N15661, N15645, N926, N2186);
nor NOR3 (N15662, N15657, N13255, N12105);
buf BUF1 (N15663, N15639);
or OR4 (N15664, N15642, N12932, N9871, N7297);
buf BUF1 (N15665, N15663);
buf BUF1 (N15666, N15661);
not NOT1 (N15667, N15647);
nand NAND2 (N15668, N15660, N11465);
not NOT1 (N15669, N15665);
xor XOR2 (N15670, N15668, N3161);
buf BUF1 (N15671, N15666);
buf BUF1 (N15672, N15671);
xor XOR2 (N15673, N15669, N4598);
xor XOR2 (N15674, N15673, N6284);
nor NOR2 (N15675, N15667, N1538);
buf BUF1 (N15676, N15664);
nor NOR2 (N15677, N15656, N7633);
nand NAND3 (N15678, N15672, N2125, N9996);
not NOT1 (N15679, N15678);
or OR2 (N15680, N15676, N14596);
buf BUF1 (N15681, N15662);
not NOT1 (N15682, N15674);
nor NOR2 (N15683, N15655, N14832);
nor NOR2 (N15684, N15683, N1219);
not NOT1 (N15685, N15679);
xor XOR2 (N15686, N15685, N5866);
xor XOR2 (N15687, N15680, N6446);
nor NOR2 (N15688, N15681, N14403);
buf BUF1 (N15689, N15675);
and AND4 (N15690, N15644, N11917, N4013, N15253);
not NOT1 (N15691, N15688);
nor NOR4 (N15692, N15689, N1421, N9792, N4230);
not NOT1 (N15693, N15687);
xor XOR2 (N15694, N15686, N8687);
nor NOR4 (N15695, N15677, N8109, N14546, N9109);
xor XOR2 (N15696, N15658, N4200);
buf BUF1 (N15697, N15692);
xor XOR2 (N15698, N15695, N2407);
nor NOR3 (N15699, N15694, N10641, N5972);
xor XOR2 (N15700, N15691, N7820);
buf BUF1 (N15701, N15700);
buf BUF1 (N15702, N15684);
buf BUF1 (N15703, N15701);
nor NOR2 (N15704, N15699, N11987);
and AND2 (N15705, N15702, N9114);
nor NOR3 (N15706, N15696, N3954, N8916);
and AND4 (N15707, N15682, N4767, N6993, N477);
buf BUF1 (N15708, N15704);
and AND3 (N15709, N15697, N6096, N2424);
buf BUF1 (N15710, N15690);
not NOT1 (N15711, N15698);
xor XOR2 (N15712, N15709, N2945);
or OR4 (N15713, N15706, N5034, N1346, N5056);
nor NOR3 (N15714, N15713, N11734, N2435);
nand NAND3 (N15715, N15708, N4416, N8045);
buf BUF1 (N15716, N15714);
not NOT1 (N15717, N15712);
xor XOR2 (N15718, N15707, N11482);
xor XOR2 (N15719, N15718, N9040);
buf BUF1 (N15720, N15670);
buf BUF1 (N15721, N15693);
not NOT1 (N15722, N15717);
xor XOR2 (N15723, N15721, N1646);
and AND4 (N15724, N15719, N9821, N4682, N12039);
not NOT1 (N15725, N15720);
nand NAND3 (N15726, N15725, N5575, N6035);
nand NAND3 (N15727, N15724, N13359, N12497);
nor NOR3 (N15728, N15705, N799, N8439);
and AND4 (N15729, N15727, N2811, N12439, N4294);
not NOT1 (N15730, N15703);
or OR4 (N15731, N15722, N101, N5867, N12986);
nand NAND3 (N15732, N15729, N12087, N6532);
not NOT1 (N15733, N15710);
and AND3 (N15734, N15715, N13866, N8099);
nor NOR2 (N15735, N15723, N15523);
xor XOR2 (N15736, N15735, N8837);
and AND4 (N15737, N15734, N8779, N12485, N12767);
xor XOR2 (N15738, N15726, N4482);
xor XOR2 (N15739, N15711, N14528);
nand NAND2 (N15740, N15737, N6123);
nor NOR3 (N15741, N15740, N7954, N11591);
nor NOR2 (N15742, N15716, N3256);
nor NOR2 (N15743, N15741, N4014);
not NOT1 (N15744, N15736);
or OR2 (N15745, N15732, N3448);
not NOT1 (N15746, N15744);
nand NAND3 (N15747, N15743, N2984, N12023);
nand NAND4 (N15748, N15738, N8806, N11968, N10973);
not NOT1 (N15749, N15733);
nand NAND2 (N15750, N15747, N14629);
xor XOR2 (N15751, N15739, N4854);
nand NAND3 (N15752, N15746, N14073, N14368);
buf BUF1 (N15753, N15745);
nor NOR2 (N15754, N15749, N3890);
nand NAND2 (N15755, N15752, N378);
buf BUF1 (N15756, N15750);
or OR4 (N15757, N15742, N12101, N13345, N12000);
and AND4 (N15758, N15753, N10180, N1491, N11784);
and AND2 (N15759, N15758, N13620);
nor NOR3 (N15760, N15728, N2026, N10590);
or OR2 (N15761, N15760, N13416);
and AND3 (N15762, N15757, N883, N9881);
nor NOR2 (N15763, N15748, N11823);
nor NOR2 (N15764, N15754, N9436);
buf BUF1 (N15765, N15764);
and AND4 (N15766, N15763, N2586, N14262, N15208);
not NOT1 (N15767, N15766);
xor XOR2 (N15768, N15762, N7651);
not NOT1 (N15769, N15767);
nor NOR3 (N15770, N15731, N993, N79);
nor NOR3 (N15771, N15769, N4630, N14954);
not NOT1 (N15772, N15771);
nor NOR2 (N15773, N15770, N2183);
nand NAND2 (N15774, N15761, N11195);
not NOT1 (N15775, N15730);
and AND4 (N15776, N15768, N5224, N9687, N13329);
not NOT1 (N15777, N15772);
not NOT1 (N15778, N15756);
xor XOR2 (N15779, N15751, N14120);
nand NAND4 (N15780, N15765, N5073, N9760, N11373);
or OR4 (N15781, N15775, N9367, N9288, N6002);
nand NAND4 (N15782, N15780, N4954, N3939, N5954);
or OR3 (N15783, N15778, N12637, N4146);
xor XOR2 (N15784, N15777, N7796);
nor NOR2 (N15785, N15784, N11870);
or OR2 (N15786, N15755, N10597);
not NOT1 (N15787, N15786);
nand NAND3 (N15788, N15787, N770, N4089);
buf BUF1 (N15789, N15776);
not NOT1 (N15790, N15774);
or OR3 (N15791, N15779, N15696, N2590);
xor XOR2 (N15792, N15782, N924);
buf BUF1 (N15793, N15785);
buf BUF1 (N15794, N15791);
or OR2 (N15795, N15794, N9461);
xor XOR2 (N15796, N15795, N5007);
xor XOR2 (N15797, N15793, N6911);
or OR2 (N15798, N15796, N8395);
and AND4 (N15799, N15781, N4438, N2909, N9131);
xor XOR2 (N15800, N15789, N10791);
or OR4 (N15801, N15800, N2491, N5801, N14937);
nor NOR2 (N15802, N15790, N333);
not NOT1 (N15803, N15801);
xor XOR2 (N15804, N15792, N15488);
not NOT1 (N15805, N15788);
and AND3 (N15806, N15797, N13916, N7494);
buf BUF1 (N15807, N15798);
buf BUF1 (N15808, N15802);
not NOT1 (N15809, N15759);
nor NOR4 (N15810, N15804, N12246, N15218, N7904);
buf BUF1 (N15811, N15783);
nor NOR2 (N15812, N15811, N642);
xor XOR2 (N15813, N15799, N12608);
xor XOR2 (N15814, N15807, N4482);
xor XOR2 (N15815, N15813, N5194);
nand NAND4 (N15816, N15808, N6085, N15586, N8769);
or OR3 (N15817, N15814, N3791, N1832);
not NOT1 (N15818, N15773);
xor XOR2 (N15819, N15817, N9436);
or OR4 (N15820, N15806, N14753, N10307, N9039);
xor XOR2 (N15821, N15820, N14360);
or OR2 (N15822, N15805, N8484);
buf BUF1 (N15823, N15812);
or OR4 (N15824, N15803, N11506, N1866, N3066);
not NOT1 (N15825, N15816);
and AND4 (N15826, N15821, N3042, N1066, N10423);
or OR3 (N15827, N15815, N2224, N2021);
xor XOR2 (N15828, N15818, N9107);
and AND4 (N15829, N15827, N5334, N13381, N6659);
buf BUF1 (N15830, N15819);
not NOT1 (N15831, N15824);
or OR4 (N15832, N15829, N13747, N13705, N10152);
nand NAND3 (N15833, N15823, N14649, N8918);
not NOT1 (N15834, N15830);
or OR2 (N15835, N15809, N7034);
and AND2 (N15836, N15825, N5644);
or OR2 (N15837, N15831, N4021);
or OR4 (N15838, N15837, N5286, N12751, N9686);
or OR3 (N15839, N15822, N13621, N11483);
and AND4 (N15840, N15826, N1856, N1547, N8392);
nand NAND3 (N15841, N15833, N96, N2201);
nor NOR2 (N15842, N15839, N15220);
not NOT1 (N15843, N15835);
buf BUF1 (N15844, N15840);
not NOT1 (N15845, N15843);
nand NAND2 (N15846, N15838, N1454);
nand NAND2 (N15847, N15834, N8155);
buf BUF1 (N15848, N15832);
not NOT1 (N15849, N15848);
nand NAND2 (N15850, N15810, N13456);
nand NAND4 (N15851, N15845, N1845, N9542, N11821);
and AND3 (N15852, N15850, N6733, N11796);
or OR2 (N15853, N15849, N10739);
xor XOR2 (N15854, N15851, N1151);
nor NOR4 (N15855, N15847, N10705, N2365, N5758);
nor NOR3 (N15856, N15828, N4692, N2067);
nand NAND3 (N15857, N15844, N1149, N13965);
buf BUF1 (N15858, N15841);
not NOT1 (N15859, N15854);
xor XOR2 (N15860, N15846, N6838);
or OR2 (N15861, N15860, N4665);
not NOT1 (N15862, N15852);
or OR4 (N15863, N15856, N14285, N6554, N6457);
nand NAND3 (N15864, N15863, N8806, N5994);
xor XOR2 (N15865, N15858, N6654);
nor NOR2 (N15866, N15842, N3299);
nand NAND2 (N15867, N15861, N8252);
xor XOR2 (N15868, N15866, N9534);
or OR3 (N15869, N15836, N14080, N12992);
not NOT1 (N15870, N15868);
xor XOR2 (N15871, N15855, N8563);
nand NAND3 (N15872, N15857, N3864, N528);
nor NOR2 (N15873, N15867, N13083);
xor XOR2 (N15874, N15873, N3802);
nor NOR3 (N15875, N15869, N4146, N6540);
nor NOR2 (N15876, N15865, N14735);
or OR3 (N15877, N15859, N13674, N2341);
and AND2 (N15878, N15872, N222);
nor NOR3 (N15879, N15870, N3276, N15732);
buf BUF1 (N15880, N15877);
nor NOR3 (N15881, N15880, N14219, N9096);
and AND2 (N15882, N15862, N3499);
not NOT1 (N15883, N15871);
nor NOR2 (N15884, N15879, N13683);
xor XOR2 (N15885, N15853, N9580);
nand NAND3 (N15886, N15882, N3479, N8424);
and AND4 (N15887, N15875, N3089, N9528, N589);
xor XOR2 (N15888, N15876, N3573);
buf BUF1 (N15889, N15881);
nor NOR3 (N15890, N15889, N15231, N14330);
nor NOR2 (N15891, N15886, N2023);
and AND2 (N15892, N15874, N10684);
and AND3 (N15893, N15890, N15303, N8994);
or OR2 (N15894, N15887, N5458);
and AND2 (N15895, N15883, N2704);
and AND2 (N15896, N15878, N1959);
buf BUF1 (N15897, N15892);
not NOT1 (N15898, N15896);
xor XOR2 (N15899, N15897, N5828);
nor NOR2 (N15900, N15885, N7780);
buf BUF1 (N15901, N15893);
xor XOR2 (N15902, N15895, N826);
buf BUF1 (N15903, N15901);
xor XOR2 (N15904, N15894, N5595);
xor XOR2 (N15905, N15891, N4357);
nor NOR4 (N15906, N15905, N1032, N3899, N11701);
or OR3 (N15907, N15903, N6826, N2317);
not NOT1 (N15908, N15902);
and AND4 (N15909, N15884, N779, N13321, N14824);
nand NAND3 (N15910, N15888, N9854, N9837);
nand NAND3 (N15911, N15899, N11415, N8966);
nand NAND3 (N15912, N15907, N2975, N6010);
nand NAND3 (N15913, N15906, N3193, N1425);
and AND2 (N15914, N15898, N3638);
and AND4 (N15915, N15908, N2305, N14417, N8006);
not NOT1 (N15916, N15912);
and AND3 (N15917, N15916, N9508, N2448);
nand NAND3 (N15918, N15913, N4428, N12026);
xor XOR2 (N15919, N15909, N15394);
and AND3 (N15920, N15917, N8745, N14358);
or OR3 (N15921, N15900, N12441, N15163);
xor XOR2 (N15922, N15904, N7273);
or OR2 (N15923, N15915, N14232);
not NOT1 (N15924, N15919);
nor NOR4 (N15925, N15923, N13588, N14640, N3687);
nand NAND2 (N15926, N15924, N6412);
not NOT1 (N15927, N15918);
and AND3 (N15928, N15926, N14068, N10759);
and AND4 (N15929, N15911, N8236, N13078, N13249);
xor XOR2 (N15930, N15929, N7901);
buf BUF1 (N15931, N15930);
not NOT1 (N15932, N15914);
or OR3 (N15933, N15910, N6905, N2820);
xor XOR2 (N15934, N15864, N4772);
not NOT1 (N15935, N15922);
xor XOR2 (N15936, N15931, N7735);
and AND3 (N15937, N15921, N7096, N6364);
buf BUF1 (N15938, N15935);
xor XOR2 (N15939, N15920, N12056);
or OR2 (N15940, N15937, N11354);
nor NOR3 (N15941, N15938, N294, N9728);
not NOT1 (N15942, N15934);
nor NOR3 (N15943, N15933, N10624, N9741);
nand NAND4 (N15944, N15928, N3145, N4996, N1124);
nand NAND4 (N15945, N15941, N622, N4516, N4786);
xor XOR2 (N15946, N15942, N3202);
or OR2 (N15947, N15927, N8936);
or OR3 (N15948, N15945, N73, N11301);
nor NOR2 (N15949, N15940, N14868);
nand NAND3 (N15950, N15936, N1488, N7105);
xor XOR2 (N15951, N15944, N5496);
and AND2 (N15952, N15943, N11980);
xor XOR2 (N15953, N15948, N6326);
nor NOR4 (N15954, N15950, N3145, N11099, N11786);
or OR4 (N15955, N15932, N13254, N12352, N7686);
not NOT1 (N15956, N15953);
nand NAND4 (N15957, N15946, N12840, N12657, N14628);
not NOT1 (N15958, N15925);
nor NOR3 (N15959, N15957, N13122, N5403);
nor NOR2 (N15960, N15956, N1691);
nor NOR3 (N15961, N15959, N11852, N13064);
not NOT1 (N15962, N15951);
buf BUF1 (N15963, N15958);
buf BUF1 (N15964, N15960);
nand NAND3 (N15965, N15949, N15304, N2325);
nand NAND4 (N15966, N15952, N13868, N7740, N830);
nand NAND4 (N15967, N15964, N3411, N8907, N5671);
not NOT1 (N15968, N15955);
buf BUF1 (N15969, N15947);
or OR4 (N15970, N15939, N9438, N14274, N10095);
and AND2 (N15971, N15970, N7328);
and AND4 (N15972, N15967, N4819, N1751, N7001);
and AND4 (N15973, N15969, N2188, N173, N8218);
xor XOR2 (N15974, N15973, N3330);
not NOT1 (N15975, N15966);
not NOT1 (N15976, N15972);
or OR2 (N15977, N15976, N13148);
nand NAND4 (N15978, N15954, N4164, N15929, N14314);
buf BUF1 (N15979, N15961);
nand NAND2 (N15980, N15979, N9548);
not NOT1 (N15981, N15977);
nor NOR2 (N15982, N15968, N792);
nor NOR2 (N15983, N15963, N1466);
buf BUF1 (N15984, N15981);
buf BUF1 (N15985, N15962);
buf BUF1 (N15986, N15984);
buf BUF1 (N15987, N15986);
xor XOR2 (N15988, N15971, N7183);
xor XOR2 (N15989, N15985, N82);
not NOT1 (N15990, N15982);
xor XOR2 (N15991, N15965, N5326);
and AND3 (N15992, N15990, N6919, N4849);
nor NOR4 (N15993, N15992, N11275, N8958, N9588);
nand NAND4 (N15994, N15988, N15250, N2928, N6526);
nor NOR4 (N15995, N15991, N12127, N9848, N631);
and AND3 (N15996, N15978, N11716, N13884);
nand NAND3 (N15997, N15996, N4058, N12424);
nor NOR3 (N15998, N15995, N12861, N10368);
xor XOR2 (N15999, N15980, N12869);
buf BUF1 (N16000, N15998);
not NOT1 (N16001, N16000);
nor NOR2 (N16002, N15997, N109);
nor NOR4 (N16003, N15987, N635, N1037, N2929);
or OR3 (N16004, N15993, N12630, N1246);
not NOT1 (N16005, N15989);
not NOT1 (N16006, N15994);
or OR3 (N16007, N16002, N7890, N6464);
and AND4 (N16008, N16006, N10932, N14511, N463);
nand NAND3 (N16009, N15974, N1222, N11051);
and AND2 (N16010, N16004, N9978);
and AND2 (N16011, N16001, N8700);
nand NAND4 (N16012, N16007, N9027, N5374, N11381);
not NOT1 (N16013, N16009);
and AND3 (N16014, N16010, N10123, N10852);
and AND3 (N16015, N15975, N12025, N13728);
and AND3 (N16016, N16015, N4315, N10278);
not NOT1 (N16017, N16008);
nand NAND4 (N16018, N16014, N8558, N12516, N3033);
or OR4 (N16019, N16018, N3305, N12270, N12896);
and AND3 (N16020, N16019, N2150, N12790);
not NOT1 (N16021, N15983);
xor XOR2 (N16022, N16012, N6318);
buf BUF1 (N16023, N15999);
nand NAND2 (N16024, N16021, N12323);
xor XOR2 (N16025, N16013, N10076);
not NOT1 (N16026, N16024);
xor XOR2 (N16027, N16022, N3653);
and AND2 (N16028, N16020, N19);
or OR4 (N16029, N16028, N489, N4382, N2432);
nand NAND3 (N16030, N16023, N7707, N14594);
nand NAND3 (N16031, N16016, N12431, N5483);
xor XOR2 (N16032, N16003, N8567);
xor XOR2 (N16033, N16029, N10636);
buf BUF1 (N16034, N16005);
or OR3 (N16035, N16031, N2027, N16023);
xor XOR2 (N16036, N16011, N7335);
buf BUF1 (N16037, N16026);
nand NAND4 (N16038, N16035, N1522, N15471, N13583);
or OR4 (N16039, N16034, N6765, N3698, N8043);
not NOT1 (N16040, N16039);
or OR3 (N16041, N16038, N8472, N7905);
nand NAND3 (N16042, N16030, N3169, N6661);
and AND4 (N16043, N16042, N11583, N14187, N1667);
nand NAND4 (N16044, N16041, N15590, N12246, N9816);
xor XOR2 (N16045, N16017, N14773);
nor NOR3 (N16046, N16044, N8009, N3778);
nand NAND3 (N16047, N16027, N1068, N7697);
nor NOR2 (N16048, N16043, N486);
nand NAND2 (N16049, N16045, N9650);
xor XOR2 (N16050, N16048, N14127);
nor NOR4 (N16051, N16036, N1086, N12913, N10470);
nor NOR4 (N16052, N16049, N3193, N6911, N14642);
nor NOR2 (N16053, N16025, N9020);
not NOT1 (N16054, N16052);
nor NOR2 (N16055, N16033, N12380);
nor NOR2 (N16056, N16046, N4573);
nand NAND2 (N16057, N16032, N3791);
nor NOR4 (N16058, N16053, N14070, N3782, N59);
nor NOR4 (N16059, N16050, N5560, N13214, N6400);
not NOT1 (N16060, N16057);
xor XOR2 (N16061, N16060, N4111);
not NOT1 (N16062, N16040);
or OR3 (N16063, N16037, N11908, N16036);
xor XOR2 (N16064, N16058, N9840);
not NOT1 (N16065, N16059);
not NOT1 (N16066, N16065);
buf BUF1 (N16067, N16054);
or OR2 (N16068, N16056, N13892);
not NOT1 (N16069, N16047);
not NOT1 (N16070, N16061);
nand NAND2 (N16071, N16064, N9958);
or OR4 (N16072, N16071, N12106, N9491, N4458);
nand NAND4 (N16073, N16070, N9612, N1395, N9258);
nor NOR3 (N16074, N16063, N1337, N7156);
xor XOR2 (N16075, N16072, N3543);
xor XOR2 (N16076, N16075, N9947);
nand NAND2 (N16077, N16062, N8749);
or OR2 (N16078, N16068, N9152);
and AND2 (N16079, N16076, N13141);
not NOT1 (N16080, N16079);
xor XOR2 (N16081, N16067, N11158);
or OR3 (N16082, N16073, N2606, N14535);
or OR4 (N16083, N16077, N2925, N8062, N3826);
or OR2 (N16084, N16081, N6584);
not NOT1 (N16085, N16078);
xor XOR2 (N16086, N16082, N3543);
nor NOR4 (N16087, N16066, N3893, N8238, N15654);
nor NOR2 (N16088, N16051, N524);
nor NOR3 (N16089, N16088, N1800, N15448);
not NOT1 (N16090, N16069);
or OR4 (N16091, N16084, N11487, N15811, N2255);
buf BUF1 (N16092, N16089);
nor NOR2 (N16093, N16083, N12290);
nand NAND3 (N16094, N16090, N13844, N7061);
xor XOR2 (N16095, N16055, N11335);
xor XOR2 (N16096, N16087, N14125);
nor NOR2 (N16097, N16095, N5609);
and AND4 (N16098, N16092, N5133, N5536, N6084);
buf BUF1 (N16099, N16086);
buf BUF1 (N16100, N16099);
xor XOR2 (N16101, N16093, N10116);
and AND2 (N16102, N16074, N4293);
or OR4 (N16103, N16101, N10832, N8495, N12347);
not NOT1 (N16104, N16091);
or OR3 (N16105, N16096, N12903, N1998);
nand NAND3 (N16106, N16097, N9734, N3764);
nand NAND3 (N16107, N16103, N436, N5824);
nand NAND2 (N16108, N16106, N8249);
nor NOR2 (N16109, N16108, N3740);
nand NAND3 (N16110, N16098, N8333, N635);
and AND4 (N16111, N16100, N9724, N15015, N7617);
nor NOR3 (N16112, N16080, N4541, N12954);
xor XOR2 (N16113, N16111, N5916);
not NOT1 (N16114, N16085);
xor XOR2 (N16115, N16114, N7573);
nor NOR4 (N16116, N16110, N12626, N8145, N8756);
and AND4 (N16117, N16107, N9713, N15129, N2542);
not NOT1 (N16118, N16102);
and AND4 (N16119, N16109, N10991, N1540, N11058);
nand NAND4 (N16120, N16119, N2024, N5222, N4235);
nand NAND3 (N16121, N16115, N5307, N12226);
nor NOR4 (N16122, N16112, N10938, N14489, N12517);
not NOT1 (N16123, N16120);
or OR2 (N16124, N16104, N12587);
or OR4 (N16125, N16105, N1011, N6250, N1442);
and AND2 (N16126, N16118, N3733);
not NOT1 (N16127, N16124);
not NOT1 (N16128, N16116);
or OR3 (N16129, N16123, N654, N6014);
nor NOR4 (N16130, N16094, N5154, N5394, N991);
xor XOR2 (N16131, N16113, N9077);
nand NAND4 (N16132, N16121, N9955, N9820, N4704);
or OR4 (N16133, N16129, N10773, N1039, N2042);
and AND4 (N16134, N16132, N9825, N11634, N5520);
or OR4 (N16135, N16134, N8569, N12919, N2852);
nor NOR4 (N16136, N16128, N7427, N11087, N15273);
nand NAND4 (N16137, N16135, N5576, N5796, N13744);
nor NOR2 (N16138, N16117, N14464);
nor NOR4 (N16139, N16127, N14815, N13567, N3353);
nor NOR4 (N16140, N16130, N2562, N16076, N2209);
and AND4 (N16141, N16136, N8009, N15537, N1796);
nand NAND2 (N16142, N16125, N9097);
nand NAND4 (N16143, N16126, N11723, N12797, N5478);
nor NOR4 (N16144, N16140, N15115, N2276, N13218);
and AND2 (N16145, N16122, N4711);
nor NOR2 (N16146, N16143, N9944);
or OR2 (N16147, N16138, N15378);
nand NAND2 (N16148, N16137, N7107);
nor NOR4 (N16149, N16144, N4588, N13438, N9855);
nor NOR3 (N16150, N16148, N10605, N15643);
xor XOR2 (N16151, N16145, N8807);
nor NOR4 (N16152, N16146, N8885, N12210, N15780);
not NOT1 (N16153, N16152);
xor XOR2 (N16154, N16139, N7371);
and AND4 (N16155, N16149, N7546, N2208, N16148);
xor XOR2 (N16156, N16151, N3330);
nor NOR3 (N16157, N16142, N9884, N7693);
and AND2 (N16158, N16155, N1613);
nor NOR2 (N16159, N16157, N2595);
buf BUF1 (N16160, N16156);
nand NAND2 (N16161, N16153, N12911);
or OR2 (N16162, N16131, N10472);
buf BUF1 (N16163, N16150);
and AND4 (N16164, N16141, N14406, N15021, N11916);
not NOT1 (N16165, N16164);
or OR2 (N16166, N16133, N12310);
xor XOR2 (N16167, N16165, N5947);
nor NOR4 (N16168, N16166, N8435, N4458, N5350);
xor XOR2 (N16169, N16167, N16077);
buf BUF1 (N16170, N16161);
xor XOR2 (N16171, N16147, N13642);
or OR3 (N16172, N16168, N9878, N15084);
and AND4 (N16173, N16169, N9133, N4041, N12279);
nand NAND3 (N16174, N16163, N10750, N15427);
nor NOR2 (N16175, N16162, N10086);
or OR4 (N16176, N16172, N8512, N2525, N4763);
and AND4 (N16177, N16159, N6103, N9613, N1315);
nor NOR3 (N16178, N16174, N7537, N1032);
or OR4 (N16179, N16176, N6684, N7001, N10123);
not NOT1 (N16180, N16173);
nor NOR2 (N16181, N16171, N12981);
nor NOR3 (N16182, N16179, N4418, N12158);
or OR3 (N16183, N16175, N6666, N2649);
buf BUF1 (N16184, N16182);
nand NAND2 (N16185, N16154, N14196);
nor NOR3 (N16186, N16160, N3278, N234);
or OR2 (N16187, N16177, N9776);
xor XOR2 (N16188, N16178, N4507);
and AND3 (N16189, N16158, N11452, N14567);
xor XOR2 (N16190, N16180, N7447);
nand NAND2 (N16191, N16184, N7825);
buf BUF1 (N16192, N16188);
not NOT1 (N16193, N16192);
buf BUF1 (N16194, N16181);
and AND4 (N16195, N16185, N15738, N6601, N12279);
nor NOR2 (N16196, N16194, N9212);
or OR2 (N16197, N16195, N197);
buf BUF1 (N16198, N16197);
or OR4 (N16199, N16198, N4287, N9885, N14104);
not NOT1 (N16200, N16187);
buf BUF1 (N16201, N16190);
buf BUF1 (N16202, N16191);
not NOT1 (N16203, N16193);
nor NOR4 (N16204, N16199, N3178, N11802, N8516);
not NOT1 (N16205, N16200);
nor NOR4 (N16206, N16203, N7735, N9467, N8190);
and AND3 (N16207, N16186, N2262, N7126);
and AND3 (N16208, N16201, N14899, N15786);
nor NOR3 (N16209, N16202, N6812, N4694);
nor NOR3 (N16210, N16204, N5026, N8102);
not NOT1 (N16211, N16196);
nor NOR4 (N16212, N16209, N8238, N9278, N1701);
or OR4 (N16213, N16212, N14574, N3359, N12120);
and AND4 (N16214, N16183, N13870, N8788, N5220);
xor XOR2 (N16215, N16210, N4108);
nor NOR4 (N16216, N16206, N9753, N6734, N12670);
or OR4 (N16217, N16207, N4119, N14590, N11169);
buf BUF1 (N16218, N16214);
or OR3 (N16219, N16170, N12219, N12553);
xor XOR2 (N16220, N16211, N13966);
and AND3 (N16221, N16217, N3670, N12921);
and AND3 (N16222, N16218, N11657, N11291);
and AND3 (N16223, N16216, N7019, N2283);
and AND2 (N16224, N16189, N8022);
xor XOR2 (N16225, N16224, N13649);
not NOT1 (N16226, N16222);
nor NOR2 (N16227, N16213, N10090);
xor XOR2 (N16228, N16223, N7228);
and AND3 (N16229, N16227, N13491, N14108);
and AND2 (N16230, N16226, N14443);
or OR3 (N16231, N16230, N1610, N1830);
and AND4 (N16232, N16215, N1461, N3819, N9508);
nand NAND3 (N16233, N16221, N94, N8915);
and AND4 (N16234, N16228, N5173, N5976, N4638);
not NOT1 (N16235, N16205);
not NOT1 (N16236, N16220);
nand NAND3 (N16237, N16229, N12418, N15854);
not NOT1 (N16238, N16234);
or OR3 (N16239, N16208, N13344, N6238);
buf BUF1 (N16240, N16239);
nor NOR2 (N16241, N16235, N4024);
buf BUF1 (N16242, N16237);
and AND3 (N16243, N16242, N2054, N2852);
nand NAND4 (N16244, N16236, N10241, N3014, N3385);
or OR2 (N16245, N16244, N4682);
nor NOR4 (N16246, N16219, N187, N9926, N15262);
and AND3 (N16247, N16240, N1922, N9235);
or OR4 (N16248, N16246, N15356, N3854, N3257);
xor XOR2 (N16249, N16241, N1974);
or OR4 (N16250, N16243, N11426, N2032, N3044);
not NOT1 (N16251, N16248);
nor NOR3 (N16252, N16249, N7087, N5869);
nor NOR2 (N16253, N16245, N6113);
xor XOR2 (N16254, N16250, N15429);
or OR4 (N16255, N16231, N7723, N12436, N1311);
nand NAND3 (N16256, N16225, N5054, N10266);
xor XOR2 (N16257, N16238, N14189);
not NOT1 (N16258, N16257);
not NOT1 (N16259, N16233);
nor NOR4 (N16260, N16252, N4541, N10612, N3168);
xor XOR2 (N16261, N16253, N11412);
xor XOR2 (N16262, N16259, N10902);
and AND4 (N16263, N16251, N1774, N14936, N1545);
not NOT1 (N16264, N16254);
buf BUF1 (N16265, N16258);
not NOT1 (N16266, N16232);
or OR2 (N16267, N16266, N1287);
nand NAND2 (N16268, N16267, N12205);
xor XOR2 (N16269, N16247, N11603);
and AND3 (N16270, N16264, N1277, N16197);
buf BUF1 (N16271, N16269);
nor NOR4 (N16272, N16270, N596, N3144, N10669);
nand NAND2 (N16273, N16265, N13330);
nor NOR2 (N16274, N16263, N2070);
xor XOR2 (N16275, N16261, N5661);
not NOT1 (N16276, N16256);
buf BUF1 (N16277, N16273);
nor NOR4 (N16278, N16260, N9314, N8183, N4758);
nand NAND2 (N16279, N16278, N13675);
nand NAND4 (N16280, N16279, N1472, N8272, N5766);
and AND4 (N16281, N16277, N14138, N13565, N6410);
nand NAND4 (N16282, N16276, N9993, N5551, N2102);
nor NOR3 (N16283, N16272, N2368, N2172);
xor XOR2 (N16284, N16271, N1457);
nand NAND2 (N16285, N16282, N4314);
buf BUF1 (N16286, N16268);
buf BUF1 (N16287, N16255);
nand NAND4 (N16288, N16274, N4579, N4486, N11952);
buf BUF1 (N16289, N16275);
and AND3 (N16290, N16281, N4488, N5894);
or OR4 (N16291, N16288, N601, N2548, N4825);
xor XOR2 (N16292, N16286, N12786);
buf BUF1 (N16293, N16290);
buf BUF1 (N16294, N16289);
and AND3 (N16295, N16283, N1082, N9957);
nand NAND2 (N16296, N16292, N16275);
xor XOR2 (N16297, N16284, N13615);
nor NOR2 (N16298, N16294, N8355);
not NOT1 (N16299, N16298);
xor XOR2 (N16300, N16262, N3342);
not NOT1 (N16301, N16293);
not NOT1 (N16302, N16280);
nor NOR4 (N16303, N16302, N12679, N14400, N5532);
buf BUF1 (N16304, N16296);
or OR3 (N16305, N16304, N984, N987);
and AND4 (N16306, N16287, N2956, N12795, N16282);
buf BUF1 (N16307, N16299);
not NOT1 (N16308, N16305);
nor NOR2 (N16309, N16300, N681);
nor NOR2 (N16310, N16308, N1423);
buf BUF1 (N16311, N16285);
and AND3 (N16312, N16297, N14564, N13449);
buf BUF1 (N16313, N16310);
and AND4 (N16314, N16306, N14996, N12833, N10316);
or OR4 (N16315, N16307, N4817, N7137, N3474);
nor NOR4 (N16316, N16303, N14933, N5691, N6369);
nand NAND2 (N16317, N16309, N9101);
not NOT1 (N16318, N16316);
nor NOR4 (N16319, N16311, N9212, N3652, N9780);
and AND3 (N16320, N16318, N8059, N14912);
not NOT1 (N16321, N16291);
nand NAND3 (N16322, N16315, N6832, N8856);
not NOT1 (N16323, N16301);
or OR3 (N16324, N16322, N3549, N13412);
not NOT1 (N16325, N16324);
xor XOR2 (N16326, N16321, N11097);
buf BUF1 (N16327, N16319);
or OR4 (N16328, N16320, N4213, N2635, N4696);
nor NOR3 (N16329, N16295, N10555, N222);
and AND4 (N16330, N16312, N11117, N7096, N869);
or OR2 (N16331, N16330, N15862);
or OR2 (N16332, N16328, N9760);
and AND4 (N16333, N16314, N9988, N1199, N5765);
buf BUF1 (N16334, N16325);
or OR2 (N16335, N16317, N674);
nor NOR3 (N16336, N16335, N1938, N3890);
and AND4 (N16337, N16313, N15996, N1217, N11651);
nor NOR4 (N16338, N16332, N7065, N941, N6136);
not NOT1 (N16339, N16326);
nor NOR3 (N16340, N16334, N12338, N12304);
nand NAND4 (N16341, N16331, N6170, N4285, N14239);
not NOT1 (N16342, N16337);
or OR3 (N16343, N16336, N4238, N6750);
buf BUF1 (N16344, N16338);
nand NAND3 (N16345, N16327, N7471, N6472);
nor NOR3 (N16346, N16344, N10193, N3598);
and AND2 (N16347, N16339, N12698);
buf BUF1 (N16348, N16346);
xor XOR2 (N16349, N16323, N14060);
buf BUF1 (N16350, N16333);
and AND3 (N16351, N16347, N14592, N9798);
nor NOR4 (N16352, N16351, N13396, N6997, N862);
or OR2 (N16353, N16329, N13900);
nor NOR4 (N16354, N16345, N2996, N2146, N14440);
and AND3 (N16355, N16349, N11719, N4272);
and AND3 (N16356, N16355, N14806, N3287);
xor XOR2 (N16357, N16340, N6911);
not NOT1 (N16358, N16343);
xor XOR2 (N16359, N16348, N5087);
or OR3 (N16360, N16350, N13681, N13476);
nand NAND4 (N16361, N16356, N14416, N3962, N10644);
and AND3 (N16362, N16359, N14339, N5408);
or OR3 (N16363, N16353, N4451, N4941);
not NOT1 (N16364, N16341);
or OR3 (N16365, N16354, N2545, N1458);
and AND4 (N16366, N16363, N7783, N12052, N12949);
not NOT1 (N16367, N16360);
nand NAND3 (N16368, N16342, N2497, N1630);
xor XOR2 (N16369, N16358, N229);
or OR2 (N16370, N16366, N7340);
nand NAND4 (N16371, N16369, N8681, N527, N25);
nand NAND2 (N16372, N16365, N6934);
and AND2 (N16373, N16370, N6464);
nor NOR4 (N16374, N16371, N12716, N12456, N8253);
xor XOR2 (N16375, N16373, N11188);
buf BUF1 (N16376, N16374);
buf BUF1 (N16377, N16375);
not NOT1 (N16378, N16367);
xor XOR2 (N16379, N16362, N2822);
not NOT1 (N16380, N16376);
or OR4 (N16381, N16377, N4303, N6172, N10999);
xor XOR2 (N16382, N16380, N8831);
nor NOR4 (N16383, N16382, N16316, N7074, N7091);
buf BUF1 (N16384, N16379);
or OR2 (N16385, N16378, N9947);
nand NAND2 (N16386, N16381, N8802);
or OR4 (N16387, N16386, N6834, N5507, N4660);
buf BUF1 (N16388, N16383);
not NOT1 (N16389, N16385);
nand NAND4 (N16390, N16361, N5713, N7146, N4037);
buf BUF1 (N16391, N16364);
or OR4 (N16392, N16391, N247, N14033, N10787);
or OR2 (N16393, N16392, N2203);
nor NOR3 (N16394, N16390, N7989, N6992);
or OR3 (N16395, N16372, N12864, N3425);
and AND4 (N16396, N16357, N9616, N4322, N2695);
nor NOR4 (N16397, N16387, N1776, N11471, N3149);
xor XOR2 (N16398, N16388, N10114);
not NOT1 (N16399, N16396);
xor XOR2 (N16400, N16393, N10529);
nor NOR3 (N16401, N16398, N13057, N2741);
nand NAND4 (N16402, N16384, N12999, N6571, N13831);
and AND4 (N16403, N16389, N352, N10396, N5638);
and AND3 (N16404, N16400, N15406, N11304);
not NOT1 (N16405, N16403);
nor NOR3 (N16406, N16394, N8848, N11669);
or OR3 (N16407, N16401, N15336, N4327);
xor XOR2 (N16408, N16368, N14784);
nand NAND2 (N16409, N16397, N4046);
buf BUF1 (N16410, N16402);
xor XOR2 (N16411, N16399, N5197);
and AND3 (N16412, N16410, N11536, N6460);
not NOT1 (N16413, N16405);
or OR3 (N16414, N16395, N10859, N16014);
or OR3 (N16415, N16409, N10344, N9917);
or OR4 (N16416, N16407, N14245, N8161, N14777);
nor NOR4 (N16417, N16404, N13194, N9064, N12956);
nand NAND4 (N16418, N16408, N6584, N5906, N3282);
not NOT1 (N16419, N16406);
xor XOR2 (N16420, N16417, N9045);
nand NAND3 (N16421, N16413, N1777, N14028);
nand NAND3 (N16422, N16420, N11091, N2840);
not NOT1 (N16423, N16415);
or OR2 (N16424, N16423, N15752);
not NOT1 (N16425, N16421);
not NOT1 (N16426, N16352);
or OR4 (N16427, N16411, N5227, N638, N12745);
nand NAND3 (N16428, N16416, N11289, N10724);
xor XOR2 (N16429, N16426, N25);
nand NAND3 (N16430, N16427, N10948, N11354);
xor XOR2 (N16431, N16428, N1405);
or OR4 (N16432, N16412, N3111, N16306, N394);
or OR2 (N16433, N16432, N1716);
nor NOR2 (N16434, N16414, N363);
nor NOR2 (N16435, N16424, N629);
not NOT1 (N16436, N16434);
xor XOR2 (N16437, N16431, N872);
nand NAND4 (N16438, N16435, N10378, N10676, N3019);
buf BUF1 (N16439, N16433);
buf BUF1 (N16440, N16439);
not NOT1 (N16441, N16438);
nor NOR3 (N16442, N16418, N14006, N3895);
buf BUF1 (N16443, N16419);
buf BUF1 (N16444, N16443);
nor NOR3 (N16445, N16440, N13747, N13102);
or OR3 (N16446, N16444, N10585, N11067);
or OR2 (N16447, N16422, N12484);
nand NAND3 (N16448, N16429, N5850, N16110);
or OR2 (N16449, N16448, N4633);
or OR2 (N16450, N16442, N66);
or OR4 (N16451, N16445, N1655, N7428, N15919);
or OR4 (N16452, N16437, N6487, N8806, N6806);
nor NOR2 (N16453, N16430, N2169);
or OR3 (N16454, N16450, N9820, N1870);
nor NOR3 (N16455, N16425, N356, N8095);
or OR4 (N16456, N16451, N1867, N13471, N7245);
or OR4 (N16457, N16454, N8415, N13426, N5620);
or OR2 (N16458, N16455, N10665);
xor XOR2 (N16459, N16447, N8374);
or OR3 (N16460, N16456, N10985, N9464);
not NOT1 (N16461, N16459);
and AND2 (N16462, N16458, N14862);
nor NOR2 (N16463, N16446, N14143);
nand NAND2 (N16464, N16463, N1692);
and AND3 (N16465, N16453, N10241, N10822);
nor NOR4 (N16466, N16449, N16324, N12404, N13702);
buf BUF1 (N16467, N16462);
xor XOR2 (N16468, N16464, N2210);
or OR3 (N16469, N16461, N15786, N2630);
not NOT1 (N16470, N16452);
buf BUF1 (N16471, N16436);
and AND2 (N16472, N16466, N486);
nand NAND3 (N16473, N16457, N12985, N10224);
nor NOR3 (N16474, N16441, N4571, N7939);
and AND2 (N16475, N16465, N16119);
xor XOR2 (N16476, N16470, N8724);
or OR4 (N16477, N16469, N16162, N4459, N7958);
or OR4 (N16478, N16468, N12357, N4492, N9487);
nand NAND4 (N16479, N16475, N5826, N7602, N15897);
xor XOR2 (N16480, N16476, N9776);
not NOT1 (N16481, N16471);
nor NOR3 (N16482, N16460, N14112, N2826);
nand NAND4 (N16483, N16479, N4417, N15082, N6382);
buf BUF1 (N16484, N16474);
nand NAND4 (N16485, N16482, N7824, N2383, N9579);
nor NOR3 (N16486, N16481, N1993, N15179);
not NOT1 (N16487, N16483);
nor NOR4 (N16488, N16478, N2237, N11412, N5149);
or OR3 (N16489, N16486, N15174, N10589);
or OR4 (N16490, N16467, N3155, N6003, N7868);
xor XOR2 (N16491, N16480, N6016);
or OR2 (N16492, N16485, N7016);
and AND3 (N16493, N16477, N8516, N6596);
xor XOR2 (N16494, N16492, N10637);
nand NAND3 (N16495, N16484, N6205, N12298);
nor NOR2 (N16496, N16488, N11059);
or OR3 (N16497, N16490, N4669, N6535);
nand NAND2 (N16498, N16495, N3502);
or OR4 (N16499, N16494, N2925, N7418, N15853);
not NOT1 (N16500, N16473);
nor NOR2 (N16501, N16496, N15489);
nand NAND3 (N16502, N16497, N7295, N1109);
not NOT1 (N16503, N16472);
nor NOR2 (N16504, N16493, N12126);
not NOT1 (N16505, N16503);
not NOT1 (N16506, N16501);
not NOT1 (N16507, N16504);
and AND2 (N16508, N16491, N12033);
not NOT1 (N16509, N16499);
and AND4 (N16510, N16507, N11546, N12538, N13532);
nand NAND2 (N16511, N16500, N15922);
nand NAND4 (N16512, N16487, N12026, N2063, N14959);
or OR4 (N16513, N16509, N2266, N8920, N3118);
nor NOR2 (N16514, N16513, N1765);
xor XOR2 (N16515, N16489, N13252);
buf BUF1 (N16516, N16511);
not NOT1 (N16517, N16516);
or OR4 (N16518, N16508, N5592, N424, N7642);
or OR4 (N16519, N16506, N1968, N13860, N1476);
buf BUF1 (N16520, N16517);
nor NOR2 (N16521, N16502, N5500);
xor XOR2 (N16522, N16510, N6921);
nor NOR2 (N16523, N16514, N13717);
nor NOR2 (N16524, N16519, N11704);
nand NAND2 (N16525, N16515, N12592);
buf BUF1 (N16526, N16521);
buf BUF1 (N16527, N16512);
xor XOR2 (N16528, N16526, N15226);
buf BUF1 (N16529, N16524);
xor XOR2 (N16530, N16505, N14823);
and AND3 (N16531, N16529, N5042, N2612);
or OR4 (N16532, N16522, N12304, N6454, N164);
or OR4 (N16533, N16525, N4378, N4410, N6938);
not NOT1 (N16534, N16523);
buf BUF1 (N16535, N16518);
or OR2 (N16536, N16530, N15236);
or OR3 (N16537, N16520, N10636, N8081);
or OR4 (N16538, N16498, N493, N629, N13335);
buf BUF1 (N16539, N16535);
or OR4 (N16540, N16537, N986, N14635, N3586);
xor XOR2 (N16541, N16531, N4369);
nor NOR2 (N16542, N16539, N12694);
or OR3 (N16543, N16534, N13520, N3745);
not NOT1 (N16544, N16538);
xor XOR2 (N16545, N16541, N4026);
or OR2 (N16546, N16536, N1037);
buf BUF1 (N16547, N16543);
not NOT1 (N16548, N16533);
xor XOR2 (N16549, N16547, N9807);
xor XOR2 (N16550, N16546, N3965);
nand NAND4 (N16551, N16550, N6431, N8272, N13816);
buf BUF1 (N16552, N16548);
xor XOR2 (N16553, N16542, N1207);
and AND2 (N16554, N16532, N4929);
buf BUF1 (N16555, N16527);
buf BUF1 (N16556, N16551);
xor XOR2 (N16557, N16554, N1017);
not NOT1 (N16558, N16555);
not NOT1 (N16559, N16552);
nand NAND2 (N16560, N16559, N13066);
buf BUF1 (N16561, N16528);
buf BUF1 (N16562, N16557);
buf BUF1 (N16563, N16562);
nor NOR4 (N16564, N16553, N4218, N4179, N947);
nand NAND3 (N16565, N16545, N1256, N193);
not NOT1 (N16566, N16556);
xor XOR2 (N16567, N16561, N3517);
not NOT1 (N16568, N16566);
or OR2 (N16569, N16560, N3829);
buf BUF1 (N16570, N16540);
xor XOR2 (N16571, N16570, N4723);
not NOT1 (N16572, N16563);
or OR3 (N16573, N16558, N11818, N12779);
and AND3 (N16574, N16572, N11489, N3237);
and AND3 (N16575, N16573, N12187, N4572);
nand NAND3 (N16576, N16564, N6545, N10285);
or OR2 (N16577, N16576, N10289);
xor XOR2 (N16578, N16568, N1721);
not NOT1 (N16579, N16565);
nor NOR2 (N16580, N16567, N4831);
buf BUF1 (N16581, N16544);
and AND2 (N16582, N16549, N8970);
nand NAND3 (N16583, N16581, N3566, N6043);
not NOT1 (N16584, N16571);
nor NOR2 (N16585, N16577, N2776);
xor XOR2 (N16586, N16585, N5724);
or OR4 (N16587, N16579, N1462, N9112, N4323);
or OR3 (N16588, N16569, N15958, N15584);
xor XOR2 (N16589, N16586, N12865);
and AND2 (N16590, N16574, N15034);
xor XOR2 (N16591, N16590, N5102);
nand NAND3 (N16592, N16587, N13835, N6396);
and AND2 (N16593, N16578, N14872);
or OR4 (N16594, N16582, N850, N5286, N8880);
nand NAND2 (N16595, N16580, N7511);
and AND3 (N16596, N16592, N6140, N3493);
not NOT1 (N16597, N16575);
or OR3 (N16598, N16593, N8274, N13452);
xor XOR2 (N16599, N16594, N6182);
nand NAND4 (N16600, N16589, N2863, N5315, N11044);
xor XOR2 (N16601, N16584, N8366);
nor NOR4 (N16602, N16600, N8935, N14046, N2926);
and AND3 (N16603, N16598, N8103, N10382);
and AND4 (N16604, N16588, N10846, N9523, N13620);
nor NOR4 (N16605, N16595, N860, N6873, N7010);
buf BUF1 (N16606, N16602);
buf BUF1 (N16607, N16591);
or OR4 (N16608, N16599, N3256, N3558, N13118);
nor NOR4 (N16609, N16601, N3957, N595, N4031);
or OR2 (N16610, N16597, N12871);
and AND2 (N16611, N16596, N2971);
nor NOR4 (N16612, N16608, N13588, N14908, N4493);
or OR3 (N16613, N16605, N13266, N11153);
xor XOR2 (N16614, N16603, N6312);
not NOT1 (N16615, N16611);
xor XOR2 (N16616, N16610, N12296);
or OR4 (N16617, N16613, N11875, N13479, N4520);
buf BUF1 (N16618, N16617);
not NOT1 (N16619, N16616);
or OR3 (N16620, N16607, N15171, N10793);
buf BUF1 (N16621, N16604);
and AND4 (N16622, N16618, N13502, N6166, N8111);
nor NOR4 (N16623, N16606, N11168, N10249, N15422);
nor NOR2 (N16624, N16583, N8445);
nand NAND4 (N16625, N16620, N9983, N1068, N1844);
and AND3 (N16626, N16622, N15076, N1613);
nand NAND3 (N16627, N16625, N6439, N11389);
and AND2 (N16628, N16624, N12434);
nor NOR4 (N16629, N16619, N2430, N15904, N15641);
buf BUF1 (N16630, N16629);
not NOT1 (N16631, N16609);
buf BUF1 (N16632, N16615);
and AND2 (N16633, N16631, N3230);
nand NAND2 (N16634, N16626, N4481);
buf BUF1 (N16635, N16614);
and AND3 (N16636, N16621, N3367, N5595);
nand NAND3 (N16637, N16627, N3442, N4548);
not NOT1 (N16638, N16634);
not NOT1 (N16639, N16632);
buf BUF1 (N16640, N16633);
buf BUF1 (N16641, N16640);
not NOT1 (N16642, N16641);
or OR2 (N16643, N16623, N12719);
buf BUF1 (N16644, N16643);
or OR2 (N16645, N16636, N1076);
nor NOR3 (N16646, N16645, N7048, N3011);
not NOT1 (N16647, N16639);
not NOT1 (N16648, N16628);
buf BUF1 (N16649, N16612);
nand NAND2 (N16650, N16648, N1649);
not NOT1 (N16651, N16650);
nor NOR3 (N16652, N16647, N16477, N4373);
nand NAND2 (N16653, N16651, N2357);
buf BUF1 (N16654, N16649);
xor XOR2 (N16655, N16630, N9206);
nor NOR2 (N16656, N16638, N8557);
or OR3 (N16657, N16654, N66, N2759);
xor XOR2 (N16658, N16653, N14627);
buf BUF1 (N16659, N16644);
or OR2 (N16660, N16646, N12810);
xor XOR2 (N16661, N16658, N5314);
and AND2 (N16662, N16637, N11537);
not NOT1 (N16663, N16656);
not NOT1 (N16664, N16635);
not NOT1 (N16665, N16652);
or OR3 (N16666, N16661, N3634, N10330);
and AND3 (N16667, N16655, N12200, N8975);
nor NOR2 (N16668, N16665, N11319);
or OR2 (N16669, N16667, N8373);
nor NOR4 (N16670, N16659, N13961, N2314, N14678);
not NOT1 (N16671, N16670);
not NOT1 (N16672, N16664);
not NOT1 (N16673, N16671);
buf BUF1 (N16674, N16657);
buf BUF1 (N16675, N16668);
xor XOR2 (N16676, N16675, N4565);
xor XOR2 (N16677, N16642, N5013);
not NOT1 (N16678, N16662);
nand NAND4 (N16679, N16663, N11037, N11770, N6478);
nor NOR4 (N16680, N16660, N6608, N781, N8907);
nand NAND3 (N16681, N16678, N15356, N4694);
not NOT1 (N16682, N16681);
nor NOR4 (N16683, N16674, N12756, N12619, N4110);
not NOT1 (N16684, N16680);
xor XOR2 (N16685, N16672, N4553);
or OR4 (N16686, N16669, N15163, N9929, N16406);
buf BUF1 (N16687, N16682);
xor XOR2 (N16688, N16677, N1513);
nor NOR3 (N16689, N16683, N9300, N15259);
nand NAND3 (N16690, N16687, N10061, N9408);
or OR2 (N16691, N16689, N13071);
xor XOR2 (N16692, N16679, N11872);
xor XOR2 (N16693, N16666, N8968);
nand NAND4 (N16694, N16690, N7933, N7250, N1525);
not NOT1 (N16695, N16685);
xor XOR2 (N16696, N16688, N13015);
buf BUF1 (N16697, N16693);
xor XOR2 (N16698, N16676, N15100);
or OR4 (N16699, N16694, N5569, N1069, N6625);
buf BUF1 (N16700, N16699);
buf BUF1 (N16701, N16700);
xor XOR2 (N16702, N16686, N1870);
nand NAND3 (N16703, N16697, N9639, N117);
not NOT1 (N16704, N16692);
or OR4 (N16705, N16673, N6479, N12318, N20);
or OR2 (N16706, N16695, N10246);
nand NAND4 (N16707, N16691, N9222, N12452, N8772);
not NOT1 (N16708, N16684);
and AND4 (N16709, N16707, N10754, N1708, N6794);
xor XOR2 (N16710, N16708, N12756);
nor NOR3 (N16711, N16706, N1816, N4674);
buf BUF1 (N16712, N16705);
buf BUF1 (N16713, N16711);
xor XOR2 (N16714, N16702, N3236);
xor XOR2 (N16715, N16712, N10800);
and AND3 (N16716, N16703, N10961, N3553);
xor XOR2 (N16717, N16713, N1581);
xor XOR2 (N16718, N16715, N3024);
buf BUF1 (N16719, N16696);
nand NAND3 (N16720, N16718, N1583, N14718);
nor NOR2 (N16721, N16710, N4855);
and AND3 (N16722, N16716, N14791, N5488);
xor XOR2 (N16723, N16719, N1171);
not NOT1 (N16724, N16720);
buf BUF1 (N16725, N16723);
or OR3 (N16726, N16701, N13556, N2952);
and AND3 (N16727, N16721, N8755, N10385);
nor NOR3 (N16728, N16727, N14345, N11831);
nor NOR2 (N16729, N16724, N61);
and AND3 (N16730, N16717, N10743, N274);
nand NAND2 (N16731, N16728, N14654);
buf BUF1 (N16732, N16722);
xor XOR2 (N16733, N16731, N8911);
nand NAND2 (N16734, N16732, N11781);
nand NAND4 (N16735, N16730, N2457, N3169, N7074);
buf BUF1 (N16736, N16729);
nand NAND2 (N16737, N16704, N5545);
xor XOR2 (N16738, N16725, N6291);
buf BUF1 (N16739, N16736);
and AND2 (N16740, N16726, N3405);
xor XOR2 (N16741, N16740, N960);
nor NOR2 (N16742, N16738, N9622);
xor XOR2 (N16743, N16733, N857);
nor NOR4 (N16744, N16735, N3998, N12977, N13694);
and AND4 (N16745, N16739, N241, N9420, N4478);
not NOT1 (N16746, N16745);
xor XOR2 (N16747, N16743, N13333);
nand NAND2 (N16748, N16744, N7567);
buf BUF1 (N16749, N16741);
and AND2 (N16750, N16746, N8191);
not NOT1 (N16751, N16714);
or OR2 (N16752, N16751, N12418);
xor XOR2 (N16753, N16750, N12148);
nand NAND3 (N16754, N16742, N7553, N8174);
or OR2 (N16755, N16737, N4734);
buf BUF1 (N16756, N16755);
nor NOR2 (N16757, N16698, N5821);
nand NAND4 (N16758, N16749, N13274, N1446, N6520);
and AND4 (N16759, N16758, N2947, N8525, N11566);
xor XOR2 (N16760, N16747, N10404);
and AND4 (N16761, N16748, N12110, N11802, N6624);
or OR2 (N16762, N16754, N15038);
nand NAND3 (N16763, N16753, N14077, N3778);
buf BUF1 (N16764, N16757);
xor XOR2 (N16765, N16764, N2280);
xor XOR2 (N16766, N16760, N6057);
buf BUF1 (N16767, N16762);
nand NAND2 (N16768, N16767, N13471);
nor NOR4 (N16769, N16752, N13308, N3660, N184);
nor NOR4 (N16770, N16765, N10211, N10532, N14986);
xor XOR2 (N16771, N16769, N5061);
xor XOR2 (N16772, N16756, N1829);
or OR4 (N16773, N16768, N216, N7120, N2230);
nand NAND3 (N16774, N16773, N6137, N3099);
nand NAND2 (N16775, N16774, N202);
or OR2 (N16776, N16772, N74);
xor XOR2 (N16777, N16770, N14182);
nand NAND3 (N16778, N16763, N8293, N2418);
or OR2 (N16779, N16734, N15680);
nor NOR2 (N16780, N16766, N4393);
buf BUF1 (N16781, N16761);
and AND4 (N16782, N16759, N13160, N16049, N4570);
or OR3 (N16783, N16775, N5079, N10709);
buf BUF1 (N16784, N16776);
and AND4 (N16785, N16783, N10680, N7043, N7430);
nand NAND3 (N16786, N16785, N13482, N15125);
and AND2 (N16787, N16778, N15231);
or OR2 (N16788, N16784, N6392);
buf BUF1 (N16789, N16780);
not NOT1 (N16790, N16777);
buf BUF1 (N16791, N16782);
xor XOR2 (N16792, N16790, N13667);
not NOT1 (N16793, N16791);
and AND4 (N16794, N16781, N13010, N16501, N6199);
buf BUF1 (N16795, N16794);
xor XOR2 (N16796, N16786, N6736);
buf BUF1 (N16797, N16789);
buf BUF1 (N16798, N16792);
and AND2 (N16799, N16793, N9833);
nand NAND4 (N16800, N16771, N4689, N12934, N10314);
not NOT1 (N16801, N16709);
nand NAND3 (N16802, N16779, N7511, N11565);
nand NAND2 (N16803, N16798, N3010);
buf BUF1 (N16804, N16795);
or OR4 (N16805, N16802, N15930, N1596, N8756);
nand NAND4 (N16806, N16804, N2351, N6716, N16801);
not NOT1 (N16807, N16669);
buf BUF1 (N16808, N16799);
and AND4 (N16809, N16788, N752, N11876, N951);
nand NAND3 (N16810, N16796, N11686, N6722);
nand NAND4 (N16811, N16787, N7280, N5211, N4350);
buf BUF1 (N16812, N16803);
not NOT1 (N16813, N16812);
and AND2 (N16814, N16808, N408);
xor XOR2 (N16815, N16797, N3482);
xor XOR2 (N16816, N16809, N16144);
nand NAND2 (N16817, N16813, N8376);
nand NAND4 (N16818, N16806, N8167, N731, N469);
nor NOR3 (N16819, N16800, N12230, N14095);
buf BUF1 (N16820, N16817);
nor NOR3 (N16821, N16816, N14386, N6200);
not NOT1 (N16822, N16815);
or OR2 (N16823, N16822, N4521);
buf BUF1 (N16824, N16810);
not NOT1 (N16825, N16820);
xor XOR2 (N16826, N16823, N16485);
or OR4 (N16827, N16821, N4668, N1243, N127);
and AND2 (N16828, N16825, N8512);
not NOT1 (N16829, N16814);
nor NOR4 (N16830, N16811, N6623, N2584, N15507);
or OR3 (N16831, N16828, N8932, N5008);
or OR2 (N16832, N16831, N12475);
and AND2 (N16833, N16824, N12807);
or OR2 (N16834, N16827, N16675);
xor XOR2 (N16835, N16819, N9126);
not NOT1 (N16836, N16826);
not NOT1 (N16837, N16835);
xor XOR2 (N16838, N16807, N14669);
nor NOR4 (N16839, N16818, N671, N1550, N1357);
xor XOR2 (N16840, N16805, N8888);
or OR4 (N16841, N16840, N6140, N2125, N7960);
nand NAND4 (N16842, N16833, N3934, N3183, N16146);
xor XOR2 (N16843, N16838, N12397);
xor XOR2 (N16844, N16842, N7045);
and AND3 (N16845, N16841, N13310, N5239);
nand NAND3 (N16846, N16844, N1292, N10461);
not NOT1 (N16847, N16832);
buf BUF1 (N16848, N16837);
not NOT1 (N16849, N16829);
not NOT1 (N16850, N16830);
nor NOR3 (N16851, N16848, N5635, N8676);
not NOT1 (N16852, N16834);
and AND2 (N16853, N16843, N4641);
or OR2 (N16854, N16847, N8991);
nor NOR2 (N16855, N16839, N16485);
not NOT1 (N16856, N16854);
xor XOR2 (N16857, N16851, N201);
not NOT1 (N16858, N16850);
xor XOR2 (N16859, N16855, N7845);
nand NAND3 (N16860, N16857, N8199, N7981);
nand NAND2 (N16861, N16849, N4493);
nand NAND2 (N16862, N16856, N12820);
nor NOR3 (N16863, N16859, N15185, N8211);
or OR4 (N16864, N16860, N16008, N2439, N1142);
not NOT1 (N16865, N16858);
or OR4 (N16866, N16864, N15718, N11915, N4496);
not NOT1 (N16867, N16846);
buf BUF1 (N16868, N16862);
not NOT1 (N16869, N16865);
nand NAND3 (N16870, N16863, N8212, N9064);
buf BUF1 (N16871, N16861);
or OR4 (N16872, N16836, N6725, N496, N12258);
nand NAND3 (N16873, N16853, N9968, N5720);
xor XOR2 (N16874, N16870, N16580);
xor XOR2 (N16875, N16867, N12938);
nor NOR3 (N16876, N16874, N8450, N12808);
nor NOR2 (N16877, N16873, N13046);
buf BUF1 (N16878, N16868);
buf BUF1 (N16879, N16869);
not NOT1 (N16880, N16877);
nand NAND4 (N16881, N16845, N1696, N14129, N7882);
nor NOR2 (N16882, N16879, N6600);
buf BUF1 (N16883, N16871);
xor XOR2 (N16884, N16875, N15006);
nor NOR4 (N16885, N16884, N15430, N4668, N16072);
not NOT1 (N16886, N16882);
or OR3 (N16887, N16883, N15281, N9322);
xor XOR2 (N16888, N16885, N6675);
nand NAND4 (N16889, N16876, N9916, N7155, N10089);
buf BUF1 (N16890, N16886);
and AND3 (N16891, N16889, N4208, N9348);
and AND2 (N16892, N16852, N3142);
not NOT1 (N16893, N16881);
nand NAND2 (N16894, N16880, N10096);
xor XOR2 (N16895, N16894, N13945);
and AND2 (N16896, N16893, N2667);
xor XOR2 (N16897, N16896, N123);
nor NOR3 (N16898, N16887, N7854, N2553);
buf BUF1 (N16899, N16895);
xor XOR2 (N16900, N16866, N15071);
buf BUF1 (N16901, N16897);
or OR3 (N16902, N16888, N9730, N11829);
nor NOR2 (N16903, N16901, N13239);
or OR3 (N16904, N16878, N13779, N5560);
or OR4 (N16905, N16891, N8705, N12937, N7610);
nor NOR3 (N16906, N16890, N8656, N10577);
and AND4 (N16907, N16892, N7700, N14519, N15486);
or OR3 (N16908, N16899, N12742, N11535);
and AND4 (N16909, N16898, N8560, N14997, N3832);
nor NOR2 (N16910, N16908, N5672);
buf BUF1 (N16911, N16910);
nor NOR3 (N16912, N16906, N5929, N11333);
not NOT1 (N16913, N16903);
and AND3 (N16914, N16907, N10961, N10701);
and AND3 (N16915, N16905, N9033, N11047);
xor XOR2 (N16916, N16872, N2516);
and AND2 (N16917, N16909, N2987);
nor NOR4 (N16918, N16917, N3948, N4790, N11684);
nor NOR4 (N16919, N16915, N5020, N3871, N15795);
or OR2 (N16920, N16914, N13580);
nor NOR2 (N16921, N16911, N15746);
not NOT1 (N16922, N16921);
nor NOR3 (N16923, N16902, N4263, N16514);
nor NOR4 (N16924, N16913, N14899, N5508, N10665);
not NOT1 (N16925, N16912);
xor XOR2 (N16926, N16919, N9342);
buf BUF1 (N16927, N16900);
and AND2 (N16928, N16923, N7455);
nand NAND2 (N16929, N16927, N7494);
nor NOR3 (N16930, N16916, N10714, N6289);
nor NOR2 (N16931, N16925, N5415);
or OR3 (N16932, N16918, N15480, N7265);
buf BUF1 (N16933, N16928);
not NOT1 (N16934, N16920);
nor NOR2 (N16935, N16933, N7758);
xor XOR2 (N16936, N16935, N9868);
not NOT1 (N16937, N16936);
buf BUF1 (N16938, N16904);
nand NAND2 (N16939, N16930, N14843);
nand NAND2 (N16940, N16934, N6431);
or OR3 (N16941, N16940, N107, N6249);
or OR3 (N16942, N16931, N11086, N5685);
buf BUF1 (N16943, N16938);
and AND2 (N16944, N16924, N8256);
nor NOR3 (N16945, N16922, N14128, N16012);
nor NOR3 (N16946, N16942, N1466, N13169);
or OR4 (N16947, N16926, N7400, N11224, N12044);
not NOT1 (N16948, N16932);
or OR4 (N16949, N16948, N10398, N13871, N13997);
and AND4 (N16950, N16937, N11958, N6369, N3268);
xor XOR2 (N16951, N16944, N15171);
or OR3 (N16952, N16945, N3213, N744);
xor XOR2 (N16953, N16950, N5732);
buf BUF1 (N16954, N16953);
nor NOR4 (N16955, N16941, N7540, N3498, N1130);
or OR2 (N16956, N16949, N10154);
buf BUF1 (N16957, N16943);
and AND3 (N16958, N16954, N1189, N5308);
and AND3 (N16959, N16952, N4037, N16900);
not NOT1 (N16960, N16958);
buf BUF1 (N16961, N16947);
and AND2 (N16962, N16946, N12890);
not NOT1 (N16963, N16960);
or OR2 (N16964, N16959, N12474);
buf BUF1 (N16965, N16963);
xor XOR2 (N16966, N16964, N13686);
not NOT1 (N16967, N16929);
and AND2 (N16968, N16951, N9363);
not NOT1 (N16969, N16957);
xor XOR2 (N16970, N16966, N1129);
nand NAND4 (N16971, N16968, N3396, N6283, N15931);
nand NAND4 (N16972, N16962, N3603, N16584, N13653);
xor XOR2 (N16973, N16969, N16823);
xor XOR2 (N16974, N16971, N1969);
nor NOR2 (N16975, N16961, N16361);
and AND4 (N16976, N16970, N14720, N9800, N7652);
not NOT1 (N16977, N16973);
xor XOR2 (N16978, N16939, N7796);
buf BUF1 (N16979, N16977);
buf BUF1 (N16980, N16955);
not NOT1 (N16981, N16965);
and AND3 (N16982, N16967, N7189, N2482);
nor NOR4 (N16983, N16974, N16454, N13382, N8405);
nor NOR4 (N16984, N16982, N123, N774, N2029);
nand NAND3 (N16985, N16981, N1698, N5635);
nor NOR4 (N16986, N16975, N16083, N1350, N9112);
nor NOR4 (N16987, N16984, N2121, N594, N10153);
nor NOR3 (N16988, N16987, N10072, N13516);
not NOT1 (N16989, N16978);
buf BUF1 (N16990, N16986);
buf BUF1 (N16991, N16983);
nand NAND3 (N16992, N16980, N7750, N8778);
or OR2 (N16993, N16979, N15413);
xor XOR2 (N16994, N16972, N5743);
nor NOR2 (N16995, N16956, N897);
and AND3 (N16996, N16990, N5187, N5285);
nor NOR2 (N16997, N16989, N1631);
not NOT1 (N16998, N16993);
nand NAND2 (N16999, N16976, N14472);
or OR2 (N17000, N16985, N11916);
or OR2 (N17001, N17000, N14926);
nor NOR4 (N17002, N16999, N13898, N6814, N8237);
nand NAND2 (N17003, N16998, N16709);
and AND4 (N17004, N16991, N9000, N7878, N13042);
and AND4 (N17005, N16995, N11419, N3512, N6364);
nand NAND3 (N17006, N17002, N14994, N1834);
xor XOR2 (N17007, N16994, N14832);
nor NOR4 (N17008, N16988, N1306, N2910, N9825);
or OR2 (N17009, N16996, N5304);
xor XOR2 (N17010, N17006, N9588);
and AND4 (N17011, N16992, N9686, N202, N11009);
buf BUF1 (N17012, N17007);
buf BUF1 (N17013, N17011);
xor XOR2 (N17014, N17008, N6048);
and AND4 (N17015, N17003, N10515, N3896, N5563);
xor XOR2 (N17016, N16997, N3107);
buf BUF1 (N17017, N17016);
nor NOR4 (N17018, N17004, N7952, N14696, N7750);
buf BUF1 (N17019, N17018);
not NOT1 (N17020, N17001);
nand NAND3 (N17021, N17020, N5563, N6813);
and AND3 (N17022, N17015, N5922, N809);
and AND3 (N17023, N17022, N6143, N5471);
and AND3 (N17024, N17017, N1683, N6328);
and AND3 (N17025, N17023, N9269, N2526);
buf BUF1 (N17026, N17025);
and AND2 (N17027, N17013, N11125);
buf BUF1 (N17028, N17009);
or OR4 (N17029, N17027, N12971, N4400, N16163);
xor XOR2 (N17030, N17005, N16778);
buf BUF1 (N17031, N17029);
nor NOR2 (N17032, N17031, N2509);
or OR4 (N17033, N17014, N10034, N1070, N3107);
or OR4 (N17034, N17012, N10067, N7790, N10385);
or OR2 (N17035, N17026, N8793);
xor XOR2 (N17036, N17035, N13749);
buf BUF1 (N17037, N17010);
nor NOR3 (N17038, N17037, N13782, N9361);
nor NOR3 (N17039, N17030, N16859, N9847);
nor NOR4 (N17040, N17036, N14374, N11607, N3427);
xor XOR2 (N17041, N17040, N14895);
buf BUF1 (N17042, N17033);
buf BUF1 (N17043, N17038);
or OR4 (N17044, N17042, N4484, N11635, N8906);
nor NOR2 (N17045, N17034, N13619);
nand NAND4 (N17046, N17041, N2825, N2763, N15525);
xor XOR2 (N17047, N17028, N5594);
nor NOR4 (N17048, N17046, N16902, N1272, N12275);
not NOT1 (N17049, N17019);
and AND4 (N17050, N17045, N16387, N12899, N4524);
and AND3 (N17051, N17043, N3406, N395);
not NOT1 (N17052, N17032);
or OR2 (N17053, N17051, N9001);
and AND3 (N17054, N17052, N6007, N6953);
or OR2 (N17055, N17047, N4254);
xor XOR2 (N17056, N17039, N5881);
xor XOR2 (N17057, N17021, N1997);
and AND4 (N17058, N17055, N6490, N10836, N8133);
and AND3 (N17059, N17044, N4336, N15257);
nand NAND4 (N17060, N17058, N2376, N16645, N2038);
or OR3 (N17061, N17056, N3965, N4964);
buf BUF1 (N17062, N17050);
xor XOR2 (N17063, N17054, N516);
or OR4 (N17064, N17053, N2525, N15805, N3929);
buf BUF1 (N17065, N17062);
xor XOR2 (N17066, N17048, N3893);
xor XOR2 (N17067, N17063, N13210);
not NOT1 (N17068, N17060);
nor NOR2 (N17069, N17067, N6120);
xor XOR2 (N17070, N17068, N15559);
not NOT1 (N17071, N17069);
nand NAND3 (N17072, N17049, N744, N15777);
buf BUF1 (N17073, N17024);
nor NOR3 (N17074, N17065, N6947, N3266);
or OR2 (N17075, N17073, N11453);
nor NOR2 (N17076, N17071, N2422);
nand NAND4 (N17077, N17066, N12938, N1730, N1950);
nand NAND4 (N17078, N17077, N15942, N14967, N14864);
nand NAND3 (N17079, N17064, N4256, N1569);
nor NOR2 (N17080, N17075, N13502);
xor XOR2 (N17081, N17072, N3953);
not NOT1 (N17082, N17070);
or OR4 (N17083, N17074, N11721, N15493, N2059);
not NOT1 (N17084, N17082);
nor NOR2 (N17085, N17078, N15121);
or OR3 (N17086, N17084, N1367, N3238);
not NOT1 (N17087, N17080);
buf BUF1 (N17088, N17081);
nand NAND3 (N17089, N17086, N13982, N13170);
or OR4 (N17090, N17059, N483, N8386, N16229);
nand NAND4 (N17091, N17088, N16284, N9311, N13739);
not NOT1 (N17092, N17089);
or OR4 (N17093, N17087, N11178, N8952, N12987);
or OR2 (N17094, N17093, N8172);
and AND2 (N17095, N17079, N8511);
buf BUF1 (N17096, N17090);
not NOT1 (N17097, N17094);
nor NOR3 (N17098, N17095, N100, N11743);
buf BUF1 (N17099, N17098);
or OR3 (N17100, N17085, N1913, N9263);
xor XOR2 (N17101, N17092, N16923);
or OR3 (N17102, N17076, N15949, N16803);
not NOT1 (N17103, N17091);
or OR3 (N17104, N17100, N12917, N5573);
or OR3 (N17105, N17103, N13049, N16937);
or OR4 (N17106, N17061, N268, N1899, N6980);
nor NOR4 (N17107, N17104, N4298, N14053, N8635);
nand NAND4 (N17108, N17096, N3200, N8379, N7220);
or OR4 (N17109, N17057, N8198, N4749, N3667);
buf BUF1 (N17110, N17106);
and AND4 (N17111, N17083, N13017, N4421, N2243);
xor XOR2 (N17112, N17108, N5933);
not NOT1 (N17113, N17110);
not NOT1 (N17114, N17102);
buf BUF1 (N17115, N17097);
not NOT1 (N17116, N17111);
or OR3 (N17117, N17112, N1753, N4533);
nand NAND3 (N17118, N17101, N3474, N16695);
nor NOR3 (N17119, N17116, N7231, N3160);
nand NAND2 (N17120, N17109, N287);
nor NOR3 (N17121, N17113, N12019, N6314);
nor NOR4 (N17122, N17121, N12281, N4189, N6512);
and AND2 (N17123, N17107, N6547);
nor NOR3 (N17124, N17119, N15975, N6577);
or OR4 (N17125, N17115, N11060, N15274, N1580);
not NOT1 (N17126, N17114);
and AND4 (N17127, N17105, N11683, N15627, N1421);
xor XOR2 (N17128, N17122, N13363);
nor NOR3 (N17129, N17124, N9676, N16980);
not NOT1 (N17130, N17129);
nand NAND3 (N17131, N17126, N5541, N3326);
and AND4 (N17132, N17120, N5227, N6581, N2097);
nand NAND3 (N17133, N17131, N15300, N12205);
or OR2 (N17134, N17123, N15795);
and AND2 (N17135, N17132, N16116);
and AND2 (N17136, N17127, N14239);
nand NAND2 (N17137, N17125, N15064);
not NOT1 (N17138, N17137);
nand NAND2 (N17139, N17133, N16062);
not NOT1 (N17140, N17128);
and AND3 (N17141, N17138, N14866, N16805);
or OR4 (N17142, N17136, N8050, N12014, N5247);
nand NAND3 (N17143, N17130, N8935, N13001);
and AND3 (N17144, N17099, N5894, N13417);
nand NAND4 (N17145, N17139, N6735, N7815, N14552);
buf BUF1 (N17146, N17117);
not NOT1 (N17147, N17143);
and AND3 (N17148, N17147, N10849, N5033);
nand NAND4 (N17149, N17146, N3583, N5938, N3464);
nor NOR4 (N17150, N17140, N9276, N5928, N9146);
buf BUF1 (N17151, N17148);
nand NAND2 (N17152, N17135, N186);
nor NOR2 (N17153, N17145, N14216);
nor NOR4 (N17154, N17134, N12942, N5517, N11598);
and AND4 (N17155, N17142, N4172, N9524, N2776);
not NOT1 (N17156, N17118);
buf BUF1 (N17157, N17150);
nor NOR3 (N17158, N17157, N13959, N10224);
nand NAND2 (N17159, N17151, N10394);
nand NAND2 (N17160, N17144, N6749);
or OR3 (N17161, N17159, N15452, N14472);
nand NAND4 (N17162, N17161, N1410, N10511, N16552);
xor XOR2 (N17163, N17153, N11183);
xor XOR2 (N17164, N17155, N11948);
nor NOR4 (N17165, N17154, N8308, N13972, N5648);
and AND2 (N17166, N17156, N6288);
and AND3 (N17167, N17152, N9609, N9835);
not NOT1 (N17168, N17166);
xor XOR2 (N17169, N17160, N2463);
not NOT1 (N17170, N17158);
nand NAND4 (N17171, N17165, N6060, N8039, N7551);
nand NAND3 (N17172, N17163, N1981, N201);
not NOT1 (N17173, N17172);
nor NOR2 (N17174, N17171, N9326);
not NOT1 (N17175, N17169);
nor NOR4 (N17176, N17164, N7095, N517, N3635);
and AND4 (N17177, N17149, N11601, N2410, N4056);
and AND2 (N17178, N17167, N4462);
not NOT1 (N17179, N17162);
buf BUF1 (N17180, N17174);
and AND4 (N17181, N17178, N1764, N3747, N10742);
and AND2 (N17182, N17173, N12368);
nand NAND2 (N17183, N17175, N3686);
xor XOR2 (N17184, N17181, N14509);
buf BUF1 (N17185, N17170);
and AND2 (N17186, N17185, N1809);
xor XOR2 (N17187, N17182, N10191);
or OR2 (N17188, N17186, N11062);
and AND4 (N17189, N17188, N2925, N14921, N6076);
buf BUF1 (N17190, N17189);
or OR4 (N17191, N17176, N7743, N6501, N14566);
and AND2 (N17192, N17180, N2247);
not NOT1 (N17193, N17187);
xor XOR2 (N17194, N17168, N11532);
nand NAND3 (N17195, N17184, N1079, N13027);
or OR2 (N17196, N17177, N11252);
and AND2 (N17197, N17141, N12671);
xor XOR2 (N17198, N17179, N2165);
xor XOR2 (N17199, N17190, N16487);
or OR2 (N17200, N17199, N884);
not NOT1 (N17201, N17183);
not NOT1 (N17202, N17200);
or OR2 (N17203, N17195, N16683);
nor NOR4 (N17204, N17191, N13475, N5945, N8574);
or OR4 (N17205, N17196, N10079, N4955, N10047);
xor XOR2 (N17206, N17203, N13720);
or OR2 (N17207, N17192, N7401);
xor XOR2 (N17208, N17202, N3619);
nor NOR4 (N17209, N17201, N8049, N6346, N298);
nor NOR3 (N17210, N17207, N13935, N2255);
nand NAND3 (N17211, N17204, N17065, N13202);
nand NAND3 (N17212, N17206, N2483, N751);
nand NAND2 (N17213, N17193, N10868);
and AND2 (N17214, N17213, N14877);
nand NAND3 (N17215, N17210, N10222, N10303);
nor NOR2 (N17216, N17212, N15556);
not NOT1 (N17217, N17205);
nor NOR2 (N17218, N17197, N14178);
buf BUF1 (N17219, N17211);
or OR2 (N17220, N17194, N5435);
buf BUF1 (N17221, N17208);
xor XOR2 (N17222, N17214, N11969);
nor NOR4 (N17223, N17222, N9305, N6266, N2220);
or OR2 (N17224, N17216, N14304);
not NOT1 (N17225, N17220);
nor NOR2 (N17226, N17221, N8704);
buf BUF1 (N17227, N17218);
nor NOR4 (N17228, N17224, N6820, N9432, N8483);
not NOT1 (N17229, N17209);
nand NAND2 (N17230, N17223, N6139);
nor NOR2 (N17231, N17229, N7293);
nor NOR4 (N17232, N17228, N2579, N9755, N11346);
nand NAND3 (N17233, N17232, N9541, N16218);
xor XOR2 (N17234, N17198, N17123);
or OR2 (N17235, N17233, N16351);
xor XOR2 (N17236, N17230, N13402);
nand NAND3 (N17237, N17227, N12259, N17132);
buf BUF1 (N17238, N17215);
buf BUF1 (N17239, N17225);
and AND2 (N17240, N17237, N5253);
nand NAND3 (N17241, N17240, N3775, N2646);
and AND3 (N17242, N17226, N16825, N6225);
nor NOR3 (N17243, N17219, N7500, N4360);
nor NOR3 (N17244, N17217, N10340, N10641);
xor XOR2 (N17245, N17234, N7455);
and AND2 (N17246, N17243, N4179);
nand NAND3 (N17247, N17246, N3284, N17032);
or OR4 (N17248, N17241, N13637, N7232, N12393);
buf BUF1 (N17249, N17248);
buf BUF1 (N17250, N17242);
nand NAND4 (N17251, N17244, N16487, N5920, N5090);
nand NAND3 (N17252, N17238, N6057, N17240);
nor NOR2 (N17253, N17247, N12202);
not NOT1 (N17254, N17253);
nor NOR4 (N17255, N17252, N15772, N11855, N3288);
nand NAND2 (N17256, N17239, N3735);
or OR4 (N17257, N17236, N13424, N335, N11322);
nand NAND2 (N17258, N17257, N16672);
nand NAND4 (N17259, N17258, N9620, N15688, N2269);
nor NOR2 (N17260, N17245, N1751);
buf BUF1 (N17261, N17254);
or OR2 (N17262, N17235, N11130);
nand NAND2 (N17263, N17249, N15341);
or OR3 (N17264, N17256, N1266, N14088);
buf BUF1 (N17265, N17259);
and AND3 (N17266, N17261, N12189, N11919);
and AND2 (N17267, N17266, N13202);
nand NAND3 (N17268, N17260, N15293, N16044);
or OR3 (N17269, N17250, N12192, N13395);
or OR3 (N17270, N17269, N9088, N885);
nor NOR4 (N17271, N17263, N3896, N5085, N13932);
buf BUF1 (N17272, N17265);
not NOT1 (N17273, N17270);
xor XOR2 (N17274, N17251, N1449);
or OR4 (N17275, N17268, N13790, N6537, N13440);
buf BUF1 (N17276, N17271);
buf BUF1 (N17277, N17267);
not NOT1 (N17278, N17274);
nand NAND4 (N17279, N17273, N1002, N2170, N9035);
xor XOR2 (N17280, N17272, N3023);
or OR2 (N17281, N17275, N15305);
buf BUF1 (N17282, N17279);
and AND4 (N17283, N17264, N9050, N15344, N16041);
nor NOR2 (N17284, N17282, N7437);
and AND3 (N17285, N17278, N4637, N15925);
and AND3 (N17286, N17277, N1044, N2505);
nand NAND3 (N17287, N17283, N11097, N12265);
not NOT1 (N17288, N17287);
buf BUF1 (N17289, N17231);
buf BUF1 (N17290, N17284);
and AND2 (N17291, N17262, N16341);
nor NOR2 (N17292, N17285, N14455);
nand NAND2 (N17293, N17291, N4864);
nand NAND4 (N17294, N17276, N3323, N9303, N13865);
and AND2 (N17295, N17286, N300);
not NOT1 (N17296, N17280);
nor NOR2 (N17297, N17293, N871);
and AND3 (N17298, N17297, N16808, N16657);
nor NOR4 (N17299, N17288, N13222, N16589, N3942);
nand NAND3 (N17300, N17289, N12052, N6427);
nand NAND2 (N17301, N17294, N10389);
xor XOR2 (N17302, N17255, N10472);
nand NAND4 (N17303, N17301, N5358, N13123, N4107);
buf BUF1 (N17304, N17303);
nor NOR4 (N17305, N17296, N11957, N11328, N15687);
nand NAND3 (N17306, N17300, N17089, N5364);
xor XOR2 (N17307, N17299, N438);
nor NOR2 (N17308, N17298, N7047);
buf BUF1 (N17309, N17306);
nand NAND4 (N17310, N17308, N5172, N16489, N8071);
xor XOR2 (N17311, N17305, N13032);
nor NOR2 (N17312, N17309, N8072);
or OR3 (N17313, N17295, N15756, N14470);
nor NOR2 (N17314, N17292, N9284);
and AND4 (N17315, N17313, N11913, N15551, N16850);
xor XOR2 (N17316, N17281, N2096);
nand NAND2 (N17317, N17302, N8054);
nor NOR2 (N17318, N17311, N6801);
and AND4 (N17319, N17316, N2491, N4384, N820);
nor NOR3 (N17320, N17290, N4843, N10427);
and AND4 (N17321, N17312, N16623, N2743, N725);
buf BUF1 (N17322, N17319);
nand NAND3 (N17323, N17307, N15792, N14755);
nand NAND4 (N17324, N17321, N14576, N9281, N13879);
not NOT1 (N17325, N17322);
not NOT1 (N17326, N17310);
buf BUF1 (N17327, N17320);
nor NOR3 (N17328, N17325, N10194, N9364);
buf BUF1 (N17329, N17318);
nor NOR2 (N17330, N17315, N5338);
xor XOR2 (N17331, N17326, N11332);
buf BUF1 (N17332, N17331);
buf BUF1 (N17333, N17330);
and AND2 (N17334, N17328, N6166);
not NOT1 (N17335, N17332);
and AND3 (N17336, N17314, N9284, N12935);
nor NOR4 (N17337, N17335, N12539, N5688, N8289);
or OR2 (N17338, N17333, N14792);
buf BUF1 (N17339, N17329);
nand NAND2 (N17340, N17327, N11484);
not NOT1 (N17341, N17340);
nor NOR3 (N17342, N17341, N16556, N2823);
not NOT1 (N17343, N17324);
nand NAND3 (N17344, N17323, N6371, N12214);
nand NAND3 (N17345, N17339, N5648, N11287);
nor NOR2 (N17346, N17317, N15650);
nand NAND4 (N17347, N17334, N122, N16796, N15139);
not NOT1 (N17348, N17338);
buf BUF1 (N17349, N17343);
buf BUF1 (N17350, N17342);
xor XOR2 (N17351, N17350, N12491);
nor NOR4 (N17352, N17349, N9792, N5685, N9506);
buf BUF1 (N17353, N17347);
and AND2 (N17354, N17348, N3234);
and AND4 (N17355, N17351, N3910, N16249, N8803);
and AND2 (N17356, N17352, N11013);
nand NAND2 (N17357, N17346, N11718);
and AND2 (N17358, N17345, N627);
and AND3 (N17359, N17358, N11457, N15924);
or OR2 (N17360, N17359, N578);
buf BUF1 (N17361, N17354);
not NOT1 (N17362, N17357);
and AND3 (N17363, N17337, N13170, N16703);
and AND4 (N17364, N17353, N14753, N10946, N16183);
buf BUF1 (N17365, N17361);
not NOT1 (N17366, N17362);
not NOT1 (N17367, N17366);
nand NAND2 (N17368, N17367, N2720);
and AND4 (N17369, N17368, N491, N13588, N5960);
and AND3 (N17370, N17369, N6719, N6103);
nor NOR3 (N17371, N17360, N3953, N10004);
and AND2 (N17372, N17355, N8469);
not NOT1 (N17373, N17336);
not NOT1 (N17374, N17371);
and AND4 (N17375, N17304, N2050, N2080, N8352);
or OR2 (N17376, N17372, N9619);
and AND3 (N17377, N17356, N5068, N11606);
buf BUF1 (N17378, N17365);
not NOT1 (N17379, N17378);
buf BUF1 (N17380, N17374);
buf BUF1 (N17381, N17375);
buf BUF1 (N17382, N17344);
nor NOR2 (N17383, N17373, N2433);
nand NAND3 (N17384, N17380, N15250, N4987);
and AND2 (N17385, N17370, N8930);
buf BUF1 (N17386, N17383);
or OR2 (N17387, N17377, N14031);
nor NOR3 (N17388, N17386, N10600, N15744);
or OR3 (N17389, N17364, N8922, N9184);
and AND4 (N17390, N17384, N13184, N15295, N5486);
nor NOR2 (N17391, N17387, N2211);
xor XOR2 (N17392, N17389, N7973);
nand NAND4 (N17393, N17392, N16556, N2116, N9187);
or OR3 (N17394, N17390, N10676, N10028);
not NOT1 (N17395, N17391);
or OR3 (N17396, N17363, N6986, N9429);
or OR3 (N17397, N17385, N3448, N11460);
xor XOR2 (N17398, N17395, N9779);
and AND3 (N17399, N17376, N8991, N6291);
and AND2 (N17400, N17382, N9260);
nor NOR2 (N17401, N17379, N15336);
buf BUF1 (N17402, N17393);
not NOT1 (N17403, N17401);
and AND3 (N17404, N17403, N3234, N16878);
and AND3 (N17405, N17404, N12100, N721);
buf BUF1 (N17406, N17388);
nor NOR3 (N17407, N17405, N17269, N3483);
nand NAND4 (N17408, N17407, N2146, N6335, N6895);
not NOT1 (N17409, N17406);
nor NOR3 (N17410, N17400, N531, N17283);
nor NOR3 (N17411, N17396, N5529, N11982);
or OR2 (N17412, N17409, N8087);
or OR2 (N17413, N17402, N8221);
and AND4 (N17414, N17408, N1184, N6166, N11313);
not NOT1 (N17415, N17398);
buf BUF1 (N17416, N17414);
buf BUF1 (N17417, N17394);
not NOT1 (N17418, N17381);
nor NOR4 (N17419, N17415, N14024, N974, N11668);
or OR2 (N17420, N17412, N11063);
and AND2 (N17421, N17413, N15299);
or OR3 (N17422, N17418, N1521, N16035);
and AND4 (N17423, N17420, N10974, N8374, N9617);
nor NOR2 (N17424, N17422, N13872);
not NOT1 (N17425, N17397);
or OR4 (N17426, N17424, N13940, N4661, N13489);
buf BUF1 (N17427, N17425);
not NOT1 (N17428, N17421);
xor XOR2 (N17429, N17428, N10722);
nor NOR4 (N17430, N17416, N14364, N14270, N13511);
and AND2 (N17431, N17411, N16);
xor XOR2 (N17432, N17426, N2472);
not NOT1 (N17433, N17431);
not NOT1 (N17434, N17429);
and AND2 (N17435, N17432, N5967);
nand NAND4 (N17436, N17419, N8294, N4806, N5169);
or OR3 (N17437, N17430, N4865, N6873);
and AND2 (N17438, N17410, N7452);
not NOT1 (N17439, N17438);
nor NOR3 (N17440, N17433, N14631, N5436);
and AND3 (N17441, N17437, N7317, N7010);
or OR4 (N17442, N17435, N365, N17304, N3123);
nand NAND3 (N17443, N17427, N3310, N2524);
nor NOR4 (N17444, N17443, N1124, N8586, N10964);
nor NOR2 (N17445, N17439, N7244);
or OR4 (N17446, N17445, N12003, N14269, N2711);
xor XOR2 (N17447, N17442, N12120);
nor NOR4 (N17448, N17417, N2379, N725, N11624);
or OR4 (N17449, N17440, N12494, N7286, N5653);
nand NAND2 (N17450, N17449, N110);
or OR3 (N17451, N17448, N11359, N13172);
xor XOR2 (N17452, N17436, N9697);
xor XOR2 (N17453, N17452, N636);
nand NAND3 (N17454, N17446, N16929, N6835);
xor XOR2 (N17455, N17434, N16199);
nor NOR3 (N17456, N17451, N12590, N1240);
xor XOR2 (N17457, N17447, N6894);
nor NOR3 (N17458, N17423, N3345, N12065);
or OR4 (N17459, N17441, N9050, N12633, N3477);
not NOT1 (N17460, N17450);
xor XOR2 (N17461, N17453, N6968);
not NOT1 (N17462, N17444);
or OR3 (N17463, N17399, N13309, N7229);
not NOT1 (N17464, N17458);
not NOT1 (N17465, N17463);
xor XOR2 (N17466, N17459, N1495);
not NOT1 (N17467, N17464);
nor NOR3 (N17468, N17460, N10908, N7502);
nand NAND3 (N17469, N17457, N3632, N4820);
buf BUF1 (N17470, N17456);
nand NAND2 (N17471, N17469, N15736);
and AND4 (N17472, N17454, N9566, N12885, N16560);
nor NOR2 (N17473, N17468, N15650);
not NOT1 (N17474, N17465);
or OR3 (N17475, N17473, N708, N15306);
buf BUF1 (N17476, N17455);
buf BUF1 (N17477, N17471);
or OR4 (N17478, N17467, N6482, N2914, N5796);
or OR3 (N17479, N17474, N10562, N15219);
not NOT1 (N17480, N17479);
buf BUF1 (N17481, N17478);
or OR2 (N17482, N17477, N11454);
xor XOR2 (N17483, N17480, N7093);
not NOT1 (N17484, N17475);
nand NAND3 (N17485, N17482, N6545, N6213);
nand NAND4 (N17486, N17484, N483, N15270, N8818);
xor XOR2 (N17487, N17470, N1540);
buf BUF1 (N17488, N17483);
and AND3 (N17489, N17461, N3447, N6225);
buf BUF1 (N17490, N17488);
and AND3 (N17491, N17462, N16160, N985);
not NOT1 (N17492, N17466);
buf BUF1 (N17493, N17476);
not NOT1 (N17494, N17491);
buf BUF1 (N17495, N17490);
or OR4 (N17496, N17481, N2809, N11409, N16860);
and AND2 (N17497, N17472, N8057);
nand NAND3 (N17498, N17485, N15285, N14834);
and AND2 (N17499, N17486, N13600);
nand NAND4 (N17500, N17489, N8408, N102, N14167);
not NOT1 (N17501, N17500);
not NOT1 (N17502, N17494);
buf BUF1 (N17503, N17496);
nand NAND2 (N17504, N17493, N10540);
or OR2 (N17505, N17499, N2892);
and AND4 (N17506, N17502, N8075, N5507, N12457);
and AND2 (N17507, N17495, N11451);
nor NOR2 (N17508, N17506, N15601);
or OR2 (N17509, N17503, N13847);
buf BUF1 (N17510, N17487);
buf BUF1 (N17511, N17509);
nand NAND2 (N17512, N17507, N8142);
buf BUF1 (N17513, N17508);
xor XOR2 (N17514, N17512, N2078);
nor NOR2 (N17515, N17501, N9743);
and AND3 (N17516, N17510, N7148, N91);
nand NAND4 (N17517, N17511, N321, N7076, N4841);
and AND2 (N17518, N17492, N7608);
and AND4 (N17519, N17518, N4767, N13995, N10852);
xor XOR2 (N17520, N17504, N7785);
nor NOR3 (N17521, N17514, N17446, N16919);
nor NOR3 (N17522, N17520, N35, N16298);
or OR3 (N17523, N17497, N186, N1220);
not NOT1 (N17524, N17521);
nor NOR2 (N17525, N17513, N13043);
and AND4 (N17526, N17524, N4982, N1321, N5150);
and AND2 (N17527, N17515, N6735);
or OR4 (N17528, N17519, N4085, N3509, N10732);
xor XOR2 (N17529, N17523, N12984);
and AND3 (N17530, N17528, N118, N14615);
nand NAND3 (N17531, N17517, N8829, N8421);
and AND2 (N17532, N17498, N16862);
not NOT1 (N17533, N17526);
buf BUF1 (N17534, N17533);
nand NAND4 (N17535, N17534, N12260, N194, N9505);
nor NOR4 (N17536, N17529, N16037, N13192, N3080);
not NOT1 (N17537, N17525);
nand NAND3 (N17538, N17527, N104, N9351);
buf BUF1 (N17539, N17532);
not NOT1 (N17540, N17539);
buf BUF1 (N17541, N17536);
xor XOR2 (N17542, N17531, N5188);
and AND3 (N17543, N17538, N10141, N8385);
and AND4 (N17544, N17541, N15091, N2573, N8457);
not NOT1 (N17545, N17516);
or OR3 (N17546, N17537, N9282, N11760);
and AND4 (N17547, N17535, N15650, N1817, N12216);
nor NOR3 (N17548, N17545, N12806, N5822);
or OR2 (N17549, N17543, N1956);
or OR3 (N17550, N17505, N13793, N13805);
or OR2 (N17551, N17540, N671);
not NOT1 (N17552, N17550);
and AND3 (N17553, N17552, N15272, N10035);
not NOT1 (N17554, N17551);
nor NOR4 (N17555, N17546, N4187, N17379, N16848);
xor XOR2 (N17556, N17547, N14048);
nor NOR2 (N17557, N17555, N7972);
and AND2 (N17558, N17557, N5269);
nand NAND2 (N17559, N17549, N7503);
buf BUF1 (N17560, N17530);
buf BUF1 (N17561, N17560);
not NOT1 (N17562, N17559);
buf BUF1 (N17563, N17544);
or OR2 (N17564, N17563, N11678);
nor NOR4 (N17565, N17564, N5986, N15651, N4505);
and AND3 (N17566, N17553, N13385, N7148);
or OR4 (N17567, N17522, N1935, N16896, N322);
not NOT1 (N17568, N17565);
buf BUF1 (N17569, N17554);
buf BUF1 (N17570, N17569);
nor NOR3 (N17571, N17567, N14534, N14507);
not NOT1 (N17572, N17562);
buf BUF1 (N17573, N17561);
not NOT1 (N17574, N17570);
not NOT1 (N17575, N17566);
and AND3 (N17576, N17571, N3064, N13577);
buf BUF1 (N17577, N17556);
not NOT1 (N17578, N17572);
nand NAND3 (N17579, N17575, N6027, N16965);
nand NAND4 (N17580, N17568, N11608, N12701, N11837);
buf BUF1 (N17581, N17579);
xor XOR2 (N17582, N17558, N6171);
not NOT1 (N17583, N17580);
and AND2 (N17584, N17573, N15648);
buf BUF1 (N17585, N17582);
nand NAND4 (N17586, N17585, N13962, N14955, N16701);
nand NAND4 (N17587, N17542, N16074, N10494, N8280);
nand NAND3 (N17588, N17574, N16902, N12025);
nor NOR4 (N17589, N17586, N12302, N3540, N10297);
not NOT1 (N17590, N17588);
not NOT1 (N17591, N17576);
or OR2 (N17592, N17583, N6121);
or OR2 (N17593, N17590, N8434);
or OR2 (N17594, N17548, N17357);
not NOT1 (N17595, N17589);
nor NOR2 (N17596, N17584, N8772);
nand NAND4 (N17597, N17594, N16633, N6236, N2361);
nor NOR4 (N17598, N17597, N17533, N10904, N10441);
not NOT1 (N17599, N17577);
nor NOR3 (N17600, N17599, N15990, N12180);
xor XOR2 (N17601, N17581, N14409);
nor NOR3 (N17602, N17593, N1400, N17216);
xor XOR2 (N17603, N17591, N16604);
nand NAND4 (N17604, N17596, N3178, N6533, N16900);
and AND4 (N17605, N17602, N10069, N16551, N1655);
not NOT1 (N17606, N17598);
nor NOR2 (N17607, N17600, N2738);
and AND3 (N17608, N17587, N4695, N4445);
buf BUF1 (N17609, N17578);
nor NOR4 (N17610, N17604, N15274, N5686, N15031);
xor XOR2 (N17611, N17606, N1750);
buf BUF1 (N17612, N17609);
buf BUF1 (N17613, N17603);
or OR4 (N17614, N17613, N6571, N6067, N13360);
buf BUF1 (N17615, N17607);
nor NOR3 (N17616, N17608, N8776, N12818);
nand NAND4 (N17617, N17616, N16651, N91, N5378);
not NOT1 (N17618, N17610);
and AND3 (N17619, N17614, N14058, N7447);
nand NAND4 (N17620, N17619, N12851, N551, N3685);
or OR2 (N17621, N17601, N13058);
and AND3 (N17622, N17618, N633, N9585);
or OR3 (N17623, N17617, N6800, N13426);
or OR3 (N17624, N17620, N1834, N14245);
nand NAND3 (N17625, N17622, N4383, N14924);
nand NAND4 (N17626, N17625, N6310, N904, N47);
nor NOR2 (N17627, N17611, N7988);
xor XOR2 (N17628, N17627, N15604);
or OR2 (N17629, N17615, N13079);
buf BUF1 (N17630, N17629);
nand NAND4 (N17631, N17592, N9468, N3640, N2598);
or OR2 (N17632, N17630, N3250);
or OR4 (N17633, N17621, N14221, N12180, N5652);
nand NAND2 (N17634, N17626, N10660);
or OR4 (N17635, N17633, N6310, N1228, N3878);
buf BUF1 (N17636, N17635);
nor NOR2 (N17637, N17632, N12361);
nand NAND3 (N17638, N17624, N553, N7001);
not NOT1 (N17639, N17636);
or OR4 (N17640, N17631, N17261, N15585, N4049);
and AND2 (N17641, N17628, N1039);
not NOT1 (N17642, N17637);
or OR3 (N17643, N17642, N7221, N11581);
not NOT1 (N17644, N17634);
nand NAND3 (N17645, N17641, N1920, N11248);
and AND3 (N17646, N17612, N16020, N2716);
and AND4 (N17647, N17595, N8963, N9000, N5191);
and AND3 (N17648, N17645, N1767, N6539);
or OR3 (N17649, N17605, N7411, N4851);
nor NOR4 (N17650, N17647, N2879, N15581, N15042);
nor NOR4 (N17651, N17650, N500, N10227, N12465);
nand NAND4 (N17652, N17639, N8535, N11658, N10123);
nand NAND4 (N17653, N17646, N4440, N13761, N3550);
nand NAND4 (N17654, N17651, N12168, N980, N4055);
nor NOR2 (N17655, N17638, N16085);
nand NAND3 (N17656, N17655, N8815, N3289);
buf BUF1 (N17657, N17656);
nor NOR2 (N17658, N17657, N11974);
and AND2 (N17659, N17623, N15520);
buf BUF1 (N17660, N17648);
nand NAND4 (N17661, N17660, N3175, N4450, N16018);
nand NAND4 (N17662, N17644, N14000, N6336, N7650);
xor XOR2 (N17663, N17649, N5638);
not NOT1 (N17664, N17662);
and AND3 (N17665, N17664, N3616, N3150);
and AND3 (N17666, N17665, N14188, N3329);
and AND3 (N17667, N17640, N5072, N10435);
not NOT1 (N17668, N17663);
nor NOR3 (N17669, N17659, N3005, N7322);
nor NOR4 (N17670, N17652, N3857, N4367, N8093);
nand NAND4 (N17671, N17670, N9772, N12323, N16898);
and AND4 (N17672, N17643, N13748, N1404, N12766);
buf BUF1 (N17673, N17654);
and AND4 (N17674, N17658, N4397, N8455, N16337);
nor NOR4 (N17675, N17674, N11329, N11810, N16088);
buf BUF1 (N17676, N17666);
or OR4 (N17677, N17671, N3516, N12219, N393);
or OR4 (N17678, N17673, N9141, N16783, N7487);
buf BUF1 (N17679, N17675);
xor XOR2 (N17680, N17667, N13139);
buf BUF1 (N17681, N17680);
and AND4 (N17682, N17653, N15455, N8264, N17597);
nand NAND4 (N17683, N17669, N4631, N7, N7259);
or OR3 (N17684, N17672, N1682, N14009);
xor XOR2 (N17685, N17678, N12568);
not NOT1 (N17686, N17676);
not NOT1 (N17687, N17681);
and AND2 (N17688, N17687, N12690);
or OR2 (N17689, N17661, N206);
xor XOR2 (N17690, N17682, N8310);
buf BUF1 (N17691, N17689);
nand NAND3 (N17692, N17679, N9550, N14435);
nand NAND4 (N17693, N17688, N17053, N11024, N11232);
nor NOR3 (N17694, N17693, N11139, N9077);
nand NAND2 (N17695, N17690, N14916);
or OR4 (N17696, N17683, N5490, N1744, N5591);
or OR2 (N17697, N17692, N9881);
nor NOR2 (N17698, N17691, N12263);
or OR4 (N17699, N17698, N11653, N5342, N10816);
buf BUF1 (N17700, N17699);
or OR4 (N17701, N17694, N13033, N5139, N7507);
or OR2 (N17702, N17677, N17011);
buf BUF1 (N17703, N17695);
nor NOR2 (N17704, N17696, N4213);
buf BUF1 (N17705, N17686);
and AND2 (N17706, N17684, N15416);
or OR4 (N17707, N17702, N16341, N13712, N1739);
buf BUF1 (N17708, N17707);
and AND2 (N17709, N17704, N17436);
nor NOR2 (N17710, N17705, N7821);
and AND2 (N17711, N17706, N14022);
nand NAND2 (N17712, N17710, N13771);
and AND2 (N17713, N17703, N6099);
buf BUF1 (N17714, N17685);
and AND3 (N17715, N17697, N15653, N11518);
nor NOR4 (N17716, N17708, N5651, N13910, N13754);
and AND2 (N17717, N17668, N17668);
buf BUF1 (N17718, N17711);
xor XOR2 (N17719, N17713, N372);
and AND4 (N17720, N17717, N15359, N10618, N14681);
xor XOR2 (N17721, N17719, N6606);
xor XOR2 (N17722, N17721, N12667);
not NOT1 (N17723, N17712);
buf BUF1 (N17724, N17714);
nor NOR4 (N17725, N17709, N248, N14324, N11647);
xor XOR2 (N17726, N17716, N2582);
nand NAND2 (N17727, N17700, N3554);
xor XOR2 (N17728, N17715, N2998);
buf BUF1 (N17729, N17726);
xor XOR2 (N17730, N17724, N15499);
and AND2 (N17731, N17727, N16439);
xor XOR2 (N17732, N17722, N7334);
not NOT1 (N17733, N17731);
or OR3 (N17734, N17720, N16843, N12005);
nand NAND4 (N17735, N17732, N16654, N8081, N17673);
nor NOR3 (N17736, N17730, N15508, N4554);
nand NAND2 (N17737, N17733, N14874);
nand NAND3 (N17738, N17718, N11071, N15426);
and AND4 (N17739, N17734, N7893, N16135, N10001);
not NOT1 (N17740, N17739);
nor NOR3 (N17741, N17729, N13482, N2618);
xor XOR2 (N17742, N17740, N2230);
or OR3 (N17743, N17741, N11568, N11188);
not NOT1 (N17744, N17723);
or OR4 (N17745, N17744, N7813, N11816, N1435);
nand NAND3 (N17746, N17701, N7519, N6128);
or OR2 (N17747, N17745, N5406);
not NOT1 (N17748, N17738);
nor NOR2 (N17749, N17737, N12022);
nand NAND2 (N17750, N17736, N5816);
xor XOR2 (N17751, N17746, N8560);
and AND3 (N17752, N17735, N7741, N2549);
not NOT1 (N17753, N17750);
xor XOR2 (N17754, N17742, N5982);
not NOT1 (N17755, N17728);
and AND2 (N17756, N17753, N2946);
nand NAND3 (N17757, N17751, N17217, N5676);
buf BUF1 (N17758, N17757);
not NOT1 (N17759, N17743);
nand NAND3 (N17760, N17749, N5624, N2045);
xor XOR2 (N17761, N17748, N5611);
or OR3 (N17762, N17752, N17674, N12474);
or OR3 (N17763, N17755, N10818, N6701);
buf BUF1 (N17764, N17758);
and AND4 (N17765, N17747, N14372, N8815, N5370);
and AND2 (N17766, N17759, N10806);
nand NAND2 (N17767, N17764, N6359);
or OR3 (N17768, N17763, N242, N5738);
nor NOR2 (N17769, N17768, N1544);
and AND2 (N17770, N17756, N1815);
xor XOR2 (N17771, N17762, N1637);
nand NAND4 (N17772, N17754, N3590, N1639, N9055);
and AND2 (N17773, N17767, N4342);
and AND3 (N17774, N17771, N13153, N5686);
nand NAND4 (N17775, N17760, N13110, N282, N461);
and AND2 (N17776, N17761, N7710);
buf BUF1 (N17777, N17765);
nor NOR4 (N17778, N17775, N13328, N7501, N2197);
and AND4 (N17779, N17777, N4803, N11743, N6501);
not NOT1 (N17780, N17770);
buf BUF1 (N17781, N17766);
nor NOR3 (N17782, N17725, N7816, N11029);
nor NOR3 (N17783, N17772, N5907, N15542);
or OR3 (N17784, N17780, N9568, N9448);
nor NOR4 (N17785, N17784, N6487, N10516, N8417);
or OR3 (N17786, N17782, N7494, N7913);
or OR3 (N17787, N17783, N4700, N15103);
nor NOR4 (N17788, N17774, N10900, N10266, N10835);
xor XOR2 (N17789, N17773, N615);
buf BUF1 (N17790, N17786);
nor NOR3 (N17791, N17785, N9726, N648);
buf BUF1 (N17792, N17789);
xor XOR2 (N17793, N17788, N14846);
nor NOR4 (N17794, N17779, N7908, N8789, N8007);
nand NAND2 (N17795, N17791, N16929);
nand NAND2 (N17796, N17795, N14034);
xor XOR2 (N17797, N17794, N15869);
and AND2 (N17798, N17797, N5542);
buf BUF1 (N17799, N17769);
xor XOR2 (N17800, N17792, N16204);
buf BUF1 (N17801, N17776);
nand NAND4 (N17802, N17787, N4915, N7323, N8128);
buf BUF1 (N17803, N17799);
xor XOR2 (N17804, N17798, N9799);
buf BUF1 (N17805, N17800);
nand NAND2 (N17806, N17778, N4736);
and AND4 (N17807, N17806, N12607, N5421, N780);
buf BUF1 (N17808, N17807);
buf BUF1 (N17809, N17801);
or OR2 (N17810, N17809, N16023);
nand NAND3 (N17811, N17793, N17315, N11975);
xor XOR2 (N17812, N17781, N4229);
and AND4 (N17813, N17790, N16326, N12976, N10626);
not NOT1 (N17814, N17808);
nand NAND4 (N17815, N17802, N2272, N13203, N7263);
nand NAND3 (N17816, N17811, N1102, N902);
not NOT1 (N17817, N17803);
not NOT1 (N17818, N17814);
nand NAND3 (N17819, N17796, N16100, N12425);
nand NAND2 (N17820, N17816, N3042);
buf BUF1 (N17821, N17804);
not NOT1 (N17822, N17810);
nand NAND4 (N17823, N17815, N2252, N6760, N16443);
nand NAND3 (N17824, N17812, N887, N17235);
buf BUF1 (N17825, N17822);
buf BUF1 (N17826, N17819);
or OR2 (N17827, N17824, N3156);
buf BUF1 (N17828, N17825);
nor NOR2 (N17829, N17827, N5343);
or OR3 (N17830, N17820, N6567, N6480);
xor XOR2 (N17831, N17817, N8725);
nor NOR2 (N17832, N17818, N15170);
or OR3 (N17833, N17826, N9902, N15162);
nor NOR4 (N17834, N17805, N12343, N13033, N1140);
and AND3 (N17835, N17813, N3169, N4813);
nand NAND3 (N17836, N17834, N12742, N3163);
buf BUF1 (N17837, N17831);
and AND2 (N17838, N17828, N15115);
nand NAND3 (N17839, N17821, N7689, N2957);
or OR4 (N17840, N17835, N1208, N9642, N14910);
nor NOR2 (N17841, N17840, N4483);
buf BUF1 (N17842, N17839);
buf BUF1 (N17843, N17842);
or OR2 (N17844, N17830, N17380);
not NOT1 (N17845, N17823);
not NOT1 (N17846, N17837);
buf BUF1 (N17847, N17832);
nor NOR4 (N17848, N17847, N15045, N9957, N2812);
xor XOR2 (N17849, N17848, N3001);
buf BUF1 (N17850, N17829);
or OR3 (N17851, N17843, N5654, N976);
or OR2 (N17852, N17833, N76);
and AND2 (N17853, N17846, N4628);
nand NAND4 (N17854, N17850, N9995, N11635, N16389);
nand NAND2 (N17855, N17845, N8383);
or OR2 (N17856, N17849, N11633);
buf BUF1 (N17857, N17852);
buf BUF1 (N17858, N17844);
and AND2 (N17859, N17854, N4185);
nor NOR2 (N17860, N17858, N6488);
buf BUF1 (N17861, N17859);
nand NAND3 (N17862, N17851, N6989, N15805);
or OR3 (N17863, N17861, N6282, N4674);
buf BUF1 (N17864, N17857);
and AND4 (N17865, N17856, N15781, N2742, N6668);
buf BUF1 (N17866, N17863);
buf BUF1 (N17867, N17838);
and AND2 (N17868, N17836, N4144);
or OR2 (N17869, N17855, N16859);
xor XOR2 (N17870, N17853, N3894);
not NOT1 (N17871, N17866);
xor XOR2 (N17872, N17864, N6873);
xor XOR2 (N17873, N17870, N8731);
nand NAND4 (N17874, N17841, N8273, N11833, N6411);
xor XOR2 (N17875, N17874, N16990);
buf BUF1 (N17876, N17873);
buf BUF1 (N17877, N17875);
and AND2 (N17878, N17876, N9891);
not NOT1 (N17879, N17872);
or OR2 (N17880, N17862, N17248);
or OR2 (N17881, N17865, N4188);
or OR3 (N17882, N17869, N3505, N2000);
not NOT1 (N17883, N17878);
or OR3 (N17884, N17871, N10178, N12047);
not NOT1 (N17885, N17882);
xor XOR2 (N17886, N17881, N5526);
nor NOR2 (N17887, N17886, N1072);
and AND4 (N17888, N17880, N10469, N5096, N1899);
nand NAND2 (N17889, N17884, N14340);
xor XOR2 (N17890, N17868, N9144);
nor NOR3 (N17891, N17883, N14632, N580);
and AND4 (N17892, N17885, N590, N13002, N16777);
not NOT1 (N17893, N17879);
buf BUF1 (N17894, N17888);
and AND4 (N17895, N17893, N15185, N9047, N8129);
or OR3 (N17896, N17890, N7653, N13965);
or OR3 (N17897, N17891, N15913, N14744);
xor XOR2 (N17898, N17889, N10450);
nor NOR2 (N17899, N17896, N16029);
nand NAND4 (N17900, N17897, N11904, N12072, N1558);
nand NAND3 (N17901, N17900, N17825, N14068);
and AND3 (N17902, N17860, N9648, N14424);
buf BUF1 (N17903, N17894);
buf BUF1 (N17904, N17902);
or OR2 (N17905, N17903, N3575);
nor NOR3 (N17906, N17867, N15702, N15934);
nor NOR2 (N17907, N17892, N7307);
and AND2 (N17908, N17898, N17808);
and AND3 (N17909, N17877, N5341, N3129);
nor NOR4 (N17910, N17907, N11741, N16901, N6268);
and AND2 (N17911, N17899, N7070);
and AND2 (N17912, N17906, N3532);
and AND2 (N17913, N17901, N9202);
or OR4 (N17914, N17904, N10823, N15705, N4792);
not NOT1 (N17915, N17909);
nand NAND2 (N17916, N17912, N5335);
not NOT1 (N17917, N17887);
xor XOR2 (N17918, N17908, N12741);
xor XOR2 (N17919, N17918, N11479);
or OR4 (N17920, N17917, N15245, N15790, N7729);
nor NOR3 (N17921, N17910, N5786, N13585);
or OR2 (N17922, N17911, N15207);
and AND4 (N17923, N17922, N3887, N1545, N15373);
nand NAND4 (N17924, N17916, N7030, N2668, N13850);
or OR4 (N17925, N17924, N7302, N1042, N11837);
nand NAND3 (N17926, N17913, N7767, N7202);
not NOT1 (N17927, N17920);
and AND3 (N17928, N17915, N3785, N6926);
buf BUF1 (N17929, N17925);
and AND2 (N17930, N17921, N4659);
nor NOR2 (N17931, N17914, N3389);
nand NAND4 (N17932, N17929, N13125, N11648, N2343);
nor NOR2 (N17933, N17928, N8759);
nor NOR2 (N17934, N17923, N13234);
not NOT1 (N17935, N17930);
buf BUF1 (N17936, N17926);
nor NOR4 (N17937, N17931, N2449, N15793, N3174);
or OR3 (N17938, N17927, N15416, N8416);
nor NOR4 (N17939, N17937, N11405, N16540, N5458);
buf BUF1 (N17940, N17939);
and AND3 (N17941, N17936, N16105, N3102);
buf BUF1 (N17942, N17938);
or OR3 (N17943, N17941, N5605, N17576);
nand NAND4 (N17944, N17933, N2216, N10083, N15965);
or OR2 (N17945, N17895, N3476);
xor XOR2 (N17946, N17919, N283);
nor NOR4 (N17947, N17934, N5465, N7592, N1147);
buf BUF1 (N17948, N17905);
xor XOR2 (N17949, N17943, N8519);
nor NOR2 (N17950, N17932, N16159);
or OR2 (N17951, N17945, N10941);
nand NAND4 (N17952, N17940, N11423, N392, N1592);
and AND2 (N17953, N17935, N4721);
buf BUF1 (N17954, N17952);
and AND3 (N17955, N17949, N11390, N13625);
or OR2 (N17956, N17948, N16429);
and AND2 (N17957, N17954, N4468);
nor NOR2 (N17958, N17946, N7754);
nand NAND3 (N17959, N17958, N10494, N3108);
xor XOR2 (N17960, N17959, N4272);
buf BUF1 (N17961, N17947);
buf BUF1 (N17962, N17957);
or OR2 (N17963, N17960, N13134);
xor XOR2 (N17964, N17953, N6715);
not NOT1 (N17965, N17955);
nand NAND2 (N17966, N17965, N6749);
nand NAND4 (N17967, N17942, N14756, N6642, N11558);
and AND2 (N17968, N17964, N7501);
nor NOR4 (N17969, N17966, N7416, N17495, N15605);
not NOT1 (N17970, N17963);
and AND2 (N17971, N17968, N4);
and AND3 (N17972, N17971, N6448, N17225);
nand NAND3 (N17973, N17956, N623, N16469);
nor NOR4 (N17974, N17950, N17642, N15943, N8205);
not NOT1 (N17975, N17972);
nand NAND4 (N17976, N17970, N16744, N14942, N3804);
xor XOR2 (N17977, N17976, N17772);
not NOT1 (N17978, N17975);
or OR2 (N17979, N17944, N6913);
or OR3 (N17980, N17969, N11236, N14209);
not NOT1 (N17981, N17961);
and AND4 (N17982, N17977, N1091, N5997, N11574);
nand NAND4 (N17983, N17951, N3558, N1261, N11270);
not NOT1 (N17984, N17962);
buf BUF1 (N17985, N17978);
and AND3 (N17986, N17982, N7959, N4243);
buf BUF1 (N17987, N17974);
xor XOR2 (N17988, N17981, N10564);
or OR4 (N17989, N17985, N3482, N10799, N972);
buf BUF1 (N17990, N17967);
or OR3 (N17991, N17979, N14804, N2798);
buf BUF1 (N17992, N17989);
or OR2 (N17993, N17987, N2257);
or OR3 (N17994, N17992, N6360, N5999);
nand NAND2 (N17995, N17980, N5631);
not NOT1 (N17996, N17988);
nand NAND3 (N17997, N17984, N3699, N10388);
or OR2 (N17998, N17986, N11102);
nor NOR3 (N17999, N17983, N16185, N16998);
buf BUF1 (N18000, N17994);
nor NOR3 (N18001, N17995, N9000, N3605);
nand NAND4 (N18002, N18001, N11833, N3127, N2381);
xor XOR2 (N18003, N18002, N17199);
buf BUF1 (N18004, N17997);
or OR2 (N18005, N17998, N16052);
buf BUF1 (N18006, N18000);
xor XOR2 (N18007, N17996, N14442);
xor XOR2 (N18008, N17990, N6909);
nand NAND2 (N18009, N18004, N16165);
not NOT1 (N18010, N17993);
buf BUF1 (N18011, N18010);
nand NAND3 (N18012, N18005, N10862, N17877);
nor NOR3 (N18013, N18006, N17842, N9107);
not NOT1 (N18014, N17999);
or OR2 (N18015, N18011, N15367);
buf BUF1 (N18016, N18015);
or OR4 (N18017, N18007, N12384, N6156, N364);
and AND4 (N18018, N18014, N1515, N5456, N14313);
nand NAND3 (N18019, N18012, N2656, N293);
not NOT1 (N18020, N18018);
nand NAND2 (N18021, N18019, N4328);
nor NOR4 (N18022, N18021, N3658, N6015, N673);
buf BUF1 (N18023, N18017);
buf BUF1 (N18024, N18023);
nand NAND4 (N18025, N18008, N2064, N8981, N3950);
buf BUF1 (N18026, N18022);
nor NOR4 (N18027, N18003, N5139, N10314, N5072);
buf BUF1 (N18028, N18024);
nand NAND2 (N18029, N17973, N5382);
not NOT1 (N18030, N18016);
and AND4 (N18031, N18020, N15963, N15746, N12847);
nand NAND4 (N18032, N18031, N4847, N6060, N7964);
buf BUF1 (N18033, N18028);
nand NAND3 (N18034, N17991, N13936, N9867);
not NOT1 (N18035, N18009);
and AND2 (N18036, N18030, N9765);
xor XOR2 (N18037, N18027, N11120);
not NOT1 (N18038, N18035);
and AND2 (N18039, N18026, N13876);
nor NOR3 (N18040, N18025, N14323, N5645);
and AND2 (N18041, N18013, N4061);
buf BUF1 (N18042, N18041);
nand NAND4 (N18043, N18040, N10280, N17252, N17370);
nor NOR4 (N18044, N18042, N2243, N4875, N8871);
nand NAND2 (N18045, N18033, N12575);
nor NOR3 (N18046, N18029, N13410, N7189);
nor NOR3 (N18047, N18045, N11618, N1021);
nand NAND3 (N18048, N18046, N12470, N6063);
or OR3 (N18049, N18044, N7966, N2702);
nand NAND3 (N18050, N18039, N15769, N5844);
and AND3 (N18051, N18043, N8980, N16401);
not NOT1 (N18052, N18032);
or OR2 (N18053, N18052, N537);
and AND2 (N18054, N18036, N3932);
xor XOR2 (N18055, N18034, N8690);
nor NOR3 (N18056, N18053, N7724, N1724);
and AND2 (N18057, N18037, N10116);
nand NAND2 (N18058, N18038, N11640);
nor NOR3 (N18059, N18047, N11956, N14067);
and AND4 (N18060, N18048, N9778, N4677, N16735);
and AND2 (N18061, N18055, N9985);
nor NOR4 (N18062, N18049, N8943, N5942, N17035);
nor NOR2 (N18063, N18051, N1623);
or OR3 (N18064, N18056, N16050, N16454);
not NOT1 (N18065, N18057);
and AND3 (N18066, N18064, N2253, N1975);
nor NOR4 (N18067, N18059, N10373, N1955, N7023);
buf BUF1 (N18068, N18058);
nor NOR2 (N18069, N18066, N17878);
nor NOR2 (N18070, N18068, N11227);
xor XOR2 (N18071, N18063, N1310);
or OR4 (N18072, N18067, N17544, N5990, N7948);
and AND2 (N18073, N18071, N3129);
xor XOR2 (N18074, N18073, N17029);
xor XOR2 (N18075, N18062, N1091);
xor XOR2 (N18076, N18050, N16257);
and AND2 (N18077, N18060, N12881);
not NOT1 (N18078, N18072);
not NOT1 (N18079, N18065);
xor XOR2 (N18080, N18074, N9591);
and AND3 (N18081, N18080, N9851, N5044);
xor XOR2 (N18082, N18075, N7703);
and AND2 (N18083, N18054, N6129);
nand NAND3 (N18084, N18061, N996, N9330);
or OR3 (N18085, N18081, N7754, N7895);
buf BUF1 (N18086, N18084);
nand NAND3 (N18087, N18085, N15812, N4242);
nor NOR4 (N18088, N18078, N5554, N1701, N17970);
xor XOR2 (N18089, N18076, N8977);
nand NAND4 (N18090, N18077, N6990, N11732, N3136);
and AND3 (N18091, N18088, N6254, N11030);
nand NAND2 (N18092, N18089, N155);
nand NAND3 (N18093, N18086, N10810, N9816);
or OR2 (N18094, N18079, N10194);
or OR2 (N18095, N18069, N634);
or OR3 (N18096, N18094, N13583, N10947);
not NOT1 (N18097, N18083);
xor XOR2 (N18098, N18070, N7723);
xor XOR2 (N18099, N18087, N17692);
not NOT1 (N18100, N18098);
nand NAND4 (N18101, N18099, N9094, N6896, N17630);
buf BUF1 (N18102, N18091);
nor NOR2 (N18103, N18095, N14268);
and AND4 (N18104, N18097, N14174, N869, N9933);
and AND2 (N18105, N18082, N15673);
not NOT1 (N18106, N18093);
not NOT1 (N18107, N18106);
and AND3 (N18108, N18096, N1175, N1053);
not NOT1 (N18109, N18102);
or OR2 (N18110, N18109, N10175);
or OR4 (N18111, N18103, N6026, N11658, N7148);
buf BUF1 (N18112, N18107);
nor NOR4 (N18113, N18105, N7946, N9021, N14292);
xor XOR2 (N18114, N18090, N752);
buf BUF1 (N18115, N18114);
nand NAND3 (N18116, N18104, N17314, N11044);
or OR2 (N18117, N18110, N4927);
or OR2 (N18118, N18116, N440);
or OR2 (N18119, N18112, N5668);
nand NAND3 (N18120, N18115, N13104, N239);
or OR2 (N18121, N18113, N1643);
not NOT1 (N18122, N18121);
nand NAND2 (N18123, N18092, N15225);
xor XOR2 (N18124, N18111, N15568);
and AND2 (N18125, N18117, N16529);
xor XOR2 (N18126, N18118, N14452);
or OR2 (N18127, N18120, N11358);
buf BUF1 (N18128, N18100);
or OR3 (N18129, N18101, N11561, N188);
nor NOR3 (N18130, N18128, N7612, N1768);
and AND4 (N18131, N18124, N16297, N3278, N9852);
buf BUF1 (N18132, N18125);
and AND3 (N18133, N18122, N1290, N11437);
xor XOR2 (N18134, N18126, N13626);
and AND4 (N18135, N18132, N16072, N8582, N17724);
and AND3 (N18136, N18129, N2279, N5197);
and AND3 (N18137, N18135, N8672, N16325);
and AND3 (N18138, N18131, N2625, N4133);
nand NAND2 (N18139, N18137, N11243);
nor NOR2 (N18140, N18123, N1565);
not NOT1 (N18141, N18130);
not NOT1 (N18142, N18133);
buf BUF1 (N18143, N18138);
not NOT1 (N18144, N18142);
nor NOR2 (N18145, N18140, N4441);
xor XOR2 (N18146, N18136, N10779);
nand NAND3 (N18147, N18141, N5466, N7580);
buf BUF1 (N18148, N18144);
nand NAND4 (N18149, N18139, N3303, N2067, N1398);
or OR4 (N18150, N18119, N1377, N3032, N7564);
not NOT1 (N18151, N18150);
not NOT1 (N18152, N18145);
nand NAND4 (N18153, N18147, N2254, N6000, N2747);
xor XOR2 (N18154, N18151, N2561);
xor XOR2 (N18155, N18108, N1957);
xor XOR2 (N18156, N18152, N5815);
and AND4 (N18157, N18143, N16743, N17209, N17969);
buf BUF1 (N18158, N18153);
buf BUF1 (N18159, N18146);
not NOT1 (N18160, N18159);
or OR3 (N18161, N18148, N8379, N7801);
buf BUF1 (N18162, N18157);
not NOT1 (N18163, N18160);
nand NAND2 (N18164, N18127, N13763);
and AND2 (N18165, N18163, N17582);
xor XOR2 (N18166, N18165, N9527);
or OR3 (N18167, N18166, N5895, N1568);
or OR3 (N18168, N18167, N11439, N379);
or OR3 (N18169, N18158, N6825, N16120);
nor NOR2 (N18170, N18154, N377);
or OR4 (N18171, N18134, N259, N8643, N2778);
buf BUF1 (N18172, N18170);
and AND3 (N18173, N18161, N2181, N327);
not NOT1 (N18174, N18156);
nand NAND3 (N18175, N18168, N4973, N896);
xor XOR2 (N18176, N18164, N7957);
buf BUF1 (N18177, N18174);
or OR3 (N18178, N18173, N3938, N16156);
and AND4 (N18179, N18177, N8179, N13537, N3597);
not NOT1 (N18180, N18155);
buf BUF1 (N18181, N18169);
not NOT1 (N18182, N18175);
not NOT1 (N18183, N18178);
or OR2 (N18184, N18176, N15663);
nor NOR2 (N18185, N18184, N11813);
nand NAND3 (N18186, N18183, N11678, N10097);
or OR3 (N18187, N18171, N6796, N11697);
nor NOR2 (N18188, N18179, N5648);
or OR3 (N18189, N18172, N13075, N7313);
nor NOR2 (N18190, N18189, N13744);
and AND2 (N18191, N18186, N9641);
xor XOR2 (N18192, N18182, N4888);
or OR4 (N18193, N18190, N11113, N5363, N17697);
not NOT1 (N18194, N18193);
and AND4 (N18195, N18180, N11983, N996, N17913);
nor NOR3 (N18196, N18185, N5278, N1613);
or OR3 (N18197, N18188, N17475, N8528);
xor XOR2 (N18198, N18196, N16843);
buf BUF1 (N18199, N18198);
nand NAND2 (N18200, N18199, N1785);
not NOT1 (N18201, N18181);
not NOT1 (N18202, N18197);
buf BUF1 (N18203, N18187);
nor NOR2 (N18204, N18194, N16074);
xor XOR2 (N18205, N18203, N13100);
nand NAND2 (N18206, N18162, N5589);
and AND4 (N18207, N18192, N13080, N7592, N9877);
and AND4 (N18208, N18149, N12909, N10967, N12454);
and AND4 (N18209, N18204, N5746, N6297, N17670);
buf BUF1 (N18210, N18207);
or OR4 (N18211, N18208, N15967, N15583, N9639);
not NOT1 (N18212, N18211);
and AND3 (N18213, N18210, N6124, N7811);
and AND2 (N18214, N18201, N9765);
xor XOR2 (N18215, N18214, N14121);
or OR4 (N18216, N18205, N1722, N10916, N10052);
and AND2 (N18217, N18202, N14232);
xor XOR2 (N18218, N18213, N569);
xor XOR2 (N18219, N18195, N11670);
and AND3 (N18220, N18219, N1523, N13325);
and AND2 (N18221, N18206, N6745);
xor XOR2 (N18222, N18215, N11272);
not NOT1 (N18223, N18220);
and AND4 (N18224, N18223, N15845, N4541, N8529);
nor NOR3 (N18225, N18224, N839, N8029);
or OR4 (N18226, N18221, N3694, N8230, N2163);
buf BUF1 (N18227, N18200);
and AND3 (N18228, N18226, N5411, N9320);
and AND3 (N18229, N18225, N11722, N13323);
nand NAND4 (N18230, N18218, N13258, N15663, N4552);
not NOT1 (N18231, N18227);
nand NAND3 (N18232, N18230, N5229, N12320);
nand NAND3 (N18233, N18222, N10130, N10790);
or OR3 (N18234, N18228, N8478, N14672);
or OR4 (N18235, N18231, N6374, N6541, N10139);
xor XOR2 (N18236, N18235, N4447);
nor NOR4 (N18237, N18232, N5592, N13449, N11789);
and AND3 (N18238, N18217, N8389, N14016);
xor XOR2 (N18239, N18234, N10661);
nand NAND4 (N18240, N18236, N10774, N9431, N9793);
and AND2 (N18241, N18237, N17950);
nor NOR2 (N18242, N18209, N15224);
or OR4 (N18243, N18242, N456, N10935, N16359);
nand NAND3 (N18244, N18191, N1164, N6552);
nand NAND4 (N18245, N18229, N7507, N15673, N17618);
not NOT1 (N18246, N18239);
nor NOR4 (N18247, N18245, N11659, N15924, N6657);
not NOT1 (N18248, N18212);
nor NOR2 (N18249, N18238, N447);
and AND4 (N18250, N18216, N11900, N17838, N2751);
buf BUF1 (N18251, N18249);
nor NOR2 (N18252, N18233, N2308);
or OR3 (N18253, N18244, N5552, N4087);
nand NAND4 (N18254, N18250, N5811, N11503, N940);
nand NAND3 (N18255, N18241, N3444, N6128);
buf BUF1 (N18256, N18253);
xor XOR2 (N18257, N18255, N1954);
not NOT1 (N18258, N18251);
not NOT1 (N18259, N18258);
nor NOR3 (N18260, N18247, N14536, N339);
xor XOR2 (N18261, N18240, N10136);
not NOT1 (N18262, N18256);
nor NOR2 (N18263, N18246, N11574);
not NOT1 (N18264, N18257);
nand NAND4 (N18265, N18248, N150, N3540, N9590);
buf BUF1 (N18266, N18262);
and AND2 (N18267, N18265, N9383);
or OR4 (N18268, N18259, N7198, N10016, N1342);
buf BUF1 (N18269, N18267);
xor XOR2 (N18270, N18243, N3211);
xor XOR2 (N18271, N18261, N11921);
or OR2 (N18272, N18260, N4064);
xor XOR2 (N18273, N18252, N3435);
or OR4 (N18274, N18271, N13123, N14948, N10534);
nor NOR4 (N18275, N18263, N18058, N10722, N13232);
not NOT1 (N18276, N18266);
not NOT1 (N18277, N18264);
buf BUF1 (N18278, N18254);
nor NOR4 (N18279, N18277, N13903, N6838, N2549);
not NOT1 (N18280, N18279);
xor XOR2 (N18281, N18270, N12001);
nor NOR3 (N18282, N18280, N6868, N9703);
or OR4 (N18283, N18278, N11853, N17819, N16580);
nand NAND4 (N18284, N18281, N2916, N645, N7624);
not NOT1 (N18285, N18269);
or OR2 (N18286, N18276, N7418);
not NOT1 (N18287, N18268);
not NOT1 (N18288, N18283);
nand NAND2 (N18289, N18284, N9744);
buf BUF1 (N18290, N18287);
nand NAND3 (N18291, N18282, N6358, N5006);
or OR4 (N18292, N18289, N10893, N3874, N313);
nand NAND4 (N18293, N18275, N11549, N3457, N16919);
or OR4 (N18294, N18273, N11492, N7135, N16731);
and AND2 (N18295, N18292, N16671);
and AND3 (N18296, N18285, N1880, N2659);
nor NOR2 (N18297, N18274, N16760);
nor NOR4 (N18298, N18288, N10525, N9000, N8454);
not NOT1 (N18299, N18290);
nand NAND3 (N18300, N18293, N3493, N12991);
and AND3 (N18301, N18299, N7695, N9672);
nor NOR3 (N18302, N18297, N14730, N371);
buf BUF1 (N18303, N18296);
nand NAND4 (N18304, N18294, N12399, N12793, N647);
or OR3 (N18305, N18303, N228, N12455);
nand NAND4 (N18306, N18300, N8588, N3968, N4625);
and AND3 (N18307, N18298, N5086, N390);
or OR3 (N18308, N18302, N11238, N13950);
and AND4 (N18309, N18306, N6600, N9732, N9458);
and AND3 (N18310, N18309, N2352, N14180);
buf BUF1 (N18311, N18286);
xor XOR2 (N18312, N18304, N9371);
not NOT1 (N18313, N18310);
not NOT1 (N18314, N18313);
xor XOR2 (N18315, N18291, N14203);
or OR4 (N18316, N18295, N17921, N927, N12643);
buf BUF1 (N18317, N18314);
xor XOR2 (N18318, N18311, N14346);
nor NOR4 (N18319, N18318, N3239, N9652, N5513);
xor XOR2 (N18320, N18301, N7207);
nor NOR2 (N18321, N18308, N11137);
xor XOR2 (N18322, N18316, N15715);
xor XOR2 (N18323, N18272, N3471);
nor NOR2 (N18324, N18312, N11550);
xor XOR2 (N18325, N18307, N11162);
xor XOR2 (N18326, N18317, N3338);
or OR4 (N18327, N18315, N6705, N5015, N12887);
nand NAND2 (N18328, N18322, N4740);
xor XOR2 (N18329, N18305, N6925);
nand NAND2 (N18330, N18323, N16004);
nor NOR2 (N18331, N18327, N3726);
buf BUF1 (N18332, N18328);
nor NOR2 (N18333, N18324, N16174);
buf BUF1 (N18334, N18320);
nor NOR4 (N18335, N18326, N8579, N1865, N9434);
and AND3 (N18336, N18321, N7988, N466);
buf BUF1 (N18337, N18329);
or OR3 (N18338, N18330, N2212, N17250);
nor NOR2 (N18339, N18337, N8809);
buf BUF1 (N18340, N18339);
not NOT1 (N18341, N18333);
xor XOR2 (N18342, N18340, N5826);
nand NAND2 (N18343, N18334, N16451);
nor NOR3 (N18344, N18338, N1016, N16215);
nor NOR4 (N18345, N18331, N7782, N18328, N11035);
nor NOR4 (N18346, N18335, N5047, N18064, N1642);
not NOT1 (N18347, N18346);
buf BUF1 (N18348, N18347);
buf BUF1 (N18349, N18319);
or OR3 (N18350, N18336, N1189, N14298);
or OR2 (N18351, N18332, N16770);
buf BUF1 (N18352, N18345);
or OR2 (N18353, N18351, N10317);
nand NAND4 (N18354, N18342, N18343, N10742, N17790);
or OR3 (N18355, N10376, N5774, N17414);
nor NOR4 (N18356, N18348, N11120, N5356, N6991);
buf BUF1 (N18357, N18325);
and AND3 (N18358, N18354, N4117, N2035);
nand NAND3 (N18359, N18350, N12456, N16103);
or OR2 (N18360, N18357, N1639);
nand NAND3 (N18361, N18353, N4370, N281);
buf BUF1 (N18362, N18358);
not NOT1 (N18363, N18344);
and AND2 (N18364, N18360, N8869);
xor XOR2 (N18365, N18363, N2517);
buf BUF1 (N18366, N18365);
xor XOR2 (N18367, N18349, N537);
not NOT1 (N18368, N18362);
buf BUF1 (N18369, N18367);
buf BUF1 (N18370, N18368);
nand NAND2 (N18371, N18355, N14112);
nand NAND3 (N18372, N18369, N12244, N15747);
not NOT1 (N18373, N18359);
xor XOR2 (N18374, N18373, N14602);
xor XOR2 (N18375, N18370, N15332);
or OR2 (N18376, N18356, N12831);
xor XOR2 (N18377, N18341, N6796);
not NOT1 (N18378, N18366);
nand NAND3 (N18379, N18376, N17535, N18234);
and AND4 (N18380, N18361, N13557, N16891, N8363);
buf BUF1 (N18381, N18374);
or OR2 (N18382, N18375, N5702);
nand NAND4 (N18383, N18379, N2656, N918, N8337);
nor NOR4 (N18384, N18364, N15998, N15624, N4125);
nor NOR2 (N18385, N18380, N10042);
not NOT1 (N18386, N18381);
not NOT1 (N18387, N18383);
or OR4 (N18388, N18387, N17873, N14680, N7564);
not NOT1 (N18389, N18372);
not NOT1 (N18390, N18382);
or OR2 (N18391, N18388, N7790);
not NOT1 (N18392, N18377);
and AND4 (N18393, N18386, N11840, N4176, N14103);
nor NOR4 (N18394, N18384, N7585, N8591, N4804);
and AND2 (N18395, N18371, N9725);
buf BUF1 (N18396, N18395);
xor XOR2 (N18397, N18352, N5155);
and AND3 (N18398, N18391, N11056, N18265);
xor XOR2 (N18399, N18385, N13411);
not NOT1 (N18400, N18378);
buf BUF1 (N18401, N18393);
xor XOR2 (N18402, N18398, N1332);
not NOT1 (N18403, N18397);
buf BUF1 (N18404, N18396);
xor XOR2 (N18405, N18399, N15659);
and AND4 (N18406, N18389, N13851, N5381, N14225);
nand NAND4 (N18407, N18406, N14440, N9808, N397);
nor NOR2 (N18408, N18404, N10290);
buf BUF1 (N18409, N18403);
not NOT1 (N18410, N18407);
buf BUF1 (N18411, N18400);
or OR4 (N18412, N18390, N7689, N6409, N3738);
and AND2 (N18413, N18394, N16053);
or OR4 (N18414, N18392, N3835, N11122, N6347);
not NOT1 (N18415, N18401);
nor NOR4 (N18416, N18410, N12823, N5497, N12396);
or OR3 (N18417, N18416, N7517, N16940);
xor XOR2 (N18418, N18412, N14339);
and AND4 (N18419, N18408, N4771, N10172, N14046);
nor NOR3 (N18420, N18409, N9220, N16229);
not NOT1 (N18421, N18415);
nor NOR2 (N18422, N18417, N11057);
and AND2 (N18423, N18420, N6481);
nand NAND3 (N18424, N18422, N10754, N2665);
not NOT1 (N18425, N18402);
nor NOR4 (N18426, N18413, N6108, N14052, N12467);
not NOT1 (N18427, N18425);
xor XOR2 (N18428, N18423, N14595);
nor NOR4 (N18429, N18411, N5649, N8603, N14082);
or OR3 (N18430, N18429, N14544, N14191);
nand NAND3 (N18431, N18418, N7539, N12795);
buf BUF1 (N18432, N18419);
buf BUF1 (N18433, N18428);
nand NAND4 (N18434, N18432, N13036, N888, N9204);
and AND2 (N18435, N18421, N4426);
nor NOR4 (N18436, N18414, N18387, N10162, N16781);
not NOT1 (N18437, N18426);
nand NAND3 (N18438, N18434, N9288, N18086);
and AND4 (N18439, N18431, N11375, N583, N16127);
nor NOR4 (N18440, N18436, N906, N13386, N3423);
not NOT1 (N18441, N18405);
and AND4 (N18442, N18424, N9461, N15806, N18068);
or OR2 (N18443, N18433, N5440);
not NOT1 (N18444, N18439);
nor NOR4 (N18445, N18443, N16031, N4027, N16231);
nor NOR2 (N18446, N18440, N2726);
buf BUF1 (N18447, N18445);
nand NAND3 (N18448, N18435, N5416, N1443);
xor XOR2 (N18449, N18447, N17260);
nand NAND4 (N18450, N18441, N2206, N18100, N8985);
nand NAND3 (N18451, N18448, N13362, N7713);
nand NAND3 (N18452, N18446, N8252, N4827);
and AND3 (N18453, N18438, N5373, N7213);
xor XOR2 (N18454, N18451, N17492);
and AND3 (N18455, N18442, N16401, N15882);
or OR3 (N18456, N18430, N15876, N14101);
xor XOR2 (N18457, N18449, N11771);
xor XOR2 (N18458, N18456, N6764);
or OR2 (N18459, N18450, N5929);
nand NAND3 (N18460, N18427, N14337, N15632);
nand NAND3 (N18461, N18454, N14879, N17780);
nand NAND2 (N18462, N18437, N6618);
nor NOR4 (N18463, N18457, N15947, N1952, N2498);
not NOT1 (N18464, N18459);
or OR3 (N18465, N18460, N11398, N14651);
xor XOR2 (N18466, N18461, N16432);
nor NOR3 (N18467, N18453, N8660, N8295);
nand NAND4 (N18468, N18465, N9312, N12435, N14597);
buf BUF1 (N18469, N18467);
nor NOR2 (N18470, N18452, N11505);
not NOT1 (N18471, N18466);
or OR2 (N18472, N18463, N442);
xor XOR2 (N18473, N18472, N17203);
or OR2 (N18474, N18470, N6469);
buf BUF1 (N18475, N18471);
buf BUF1 (N18476, N18462);
xor XOR2 (N18477, N18476, N7077);
nand NAND2 (N18478, N18477, N15439);
or OR4 (N18479, N18464, N11647, N15713, N2848);
or OR2 (N18480, N18444, N5285);
xor XOR2 (N18481, N18458, N10990);
nand NAND4 (N18482, N18468, N15204, N14733, N1383);
not NOT1 (N18483, N18473);
nand NAND3 (N18484, N18475, N11076, N7489);
not NOT1 (N18485, N18482);
and AND4 (N18486, N18469, N12400, N16115, N8843);
and AND3 (N18487, N18474, N10812, N14728);
nor NOR2 (N18488, N18486, N14490);
nor NOR4 (N18489, N18478, N17994, N7993, N4271);
or OR4 (N18490, N18480, N14416, N8861, N13690);
xor XOR2 (N18491, N18479, N16179);
and AND4 (N18492, N18484, N860, N11107, N2372);
not NOT1 (N18493, N18481);
and AND3 (N18494, N18489, N10629, N14403);
xor XOR2 (N18495, N18490, N468);
xor XOR2 (N18496, N18492, N14120);
nor NOR2 (N18497, N18493, N18215);
nand NAND4 (N18498, N18494, N1336, N6623, N16765);
nor NOR3 (N18499, N18495, N639, N14506);
nand NAND3 (N18500, N18483, N10341, N11658);
nand NAND3 (N18501, N18498, N1347, N5482);
nand NAND4 (N18502, N18488, N6140, N11407, N179);
nand NAND2 (N18503, N18502, N8197);
buf BUF1 (N18504, N18503);
and AND3 (N18505, N18491, N16299, N3881);
nor NOR4 (N18506, N18504, N1883, N4850, N16184);
or OR4 (N18507, N18500, N14461, N10245, N14296);
or OR4 (N18508, N18506, N13972, N13958, N4865);
and AND3 (N18509, N18496, N17663, N16670);
and AND2 (N18510, N18501, N8716);
buf BUF1 (N18511, N18507);
buf BUF1 (N18512, N18510);
or OR4 (N18513, N18455, N6510, N8515, N10017);
and AND4 (N18514, N18511, N11611, N2718, N4408);
not NOT1 (N18515, N18512);
not NOT1 (N18516, N18515);
nand NAND2 (N18517, N18497, N11753);
xor XOR2 (N18518, N18505, N9950);
xor XOR2 (N18519, N18509, N4547);
or OR2 (N18520, N18513, N13641);
not NOT1 (N18521, N18499);
buf BUF1 (N18522, N18519);
or OR2 (N18523, N18516, N259);
not NOT1 (N18524, N18517);
buf BUF1 (N18525, N18524);
xor XOR2 (N18526, N18485, N16046);
nand NAND4 (N18527, N18525, N4364, N5832, N4832);
xor XOR2 (N18528, N18508, N13966);
or OR2 (N18529, N18520, N359);
xor XOR2 (N18530, N18518, N18420);
buf BUF1 (N18531, N18526);
and AND4 (N18532, N18527, N78, N12438, N1387);
xor XOR2 (N18533, N18523, N17677);
buf BUF1 (N18534, N18533);
and AND2 (N18535, N18487, N4978);
xor XOR2 (N18536, N18532, N5013);
buf BUF1 (N18537, N18531);
or OR3 (N18538, N18514, N16428, N10232);
buf BUF1 (N18539, N18529);
or OR3 (N18540, N18536, N16672, N5626);
nand NAND4 (N18541, N18535, N2354, N18494, N3123);
nor NOR2 (N18542, N18540, N8965);
or OR3 (N18543, N18522, N14049, N16386);
xor XOR2 (N18544, N18528, N15972);
not NOT1 (N18545, N18541);
buf BUF1 (N18546, N18544);
xor XOR2 (N18547, N18543, N15532);
not NOT1 (N18548, N18539);
not NOT1 (N18549, N18548);
xor XOR2 (N18550, N18538, N3710);
or OR4 (N18551, N18545, N4540, N3962, N7289);
xor XOR2 (N18552, N18530, N4082);
and AND3 (N18553, N18546, N3498, N11884);
and AND4 (N18554, N18551, N12956, N8592, N1155);
nand NAND4 (N18555, N18534, N2534, N18554, N16296);
and AND2 (N18556, N957, N14394);
nand NAND4 (N18557, N18521, N1694, N16932, N4791);
and AND2 (N18558, N18555, N18521);
xor XOR2 (N18559, N18552, N6180);
or OR4 (N18560, N18553, N13175, N6325, N13834);
and AND3 (N18561, N18542, N2974, N14825);
buf BUF1 (N18562, N18557);
not NOT1 (N18563, N18547);
nor NOR2 (N18564, N18560, N4304);
or OR4 (N18565, N18563, N5724, N14664, N8479);
xor XOR2 (N18566, N18556, N9125);
nor NOR3 (N18567, N18549, N12421, N3209);
and AND2 (N18568, N18566, N2493);
xor XOR2 (N18569, N18561, N1219);
not NOT1 (N18570, N18559);
nor NOR3 (N18571, N18550, N9378, N6840);
buf BUF1 (N18572, N18568);
or OR4 (N18573, N18564, N16349, N10503, N716);
and AND3 (N18574, N18558, N4089, N14559);
nand NAND2 (N18575, N18569, N5122);
xor XOR2 (N18576, N18572, N4467);
nor NOR3 (N18577, N18575, N6583, N5387);
xor XOR2 (N18578, N18570, N2867);
not NOT1 (N18579, N18574);
not NOT1 (N18580, N18567);
nor NOR2 (N18581, N18576, N9552);
xor XOR2 (N18582, N18565, N10590);
and AND2 (N18583, N18562, N18260);
xor XOR2 (N18584, N18578, N5077);
nor NOR3 (N18585, N18577, N2929, N14801);
xor XOR2 (N18586, N18571, N11897);
not NOT1 (N18587, N18573);
not NOT1 (N18588, N18585);
buf BUF1 (N18589, N18580);
nor NOR3 (N18590, N18583, N18562, N10300);
buf BUF1 (N18591, N18579);
or OR3 (N18592, N18591, N11365, N10890);
nor NOR4 (N18593, N18584, N10566, N12718, N14901);
or OR4 (N18594, N18587, N9746, N3551, N3174);
xor XOR2 (N18595, N18586, N5000);
and AND3 (N18596, N18594, N5198, N3739);
and AND2 (N18597, N18596, N390);
nand NAND2 (N18598, N18537, N7055);
or OR3 (N18599, N18588, N15764, N6794);
buf BUF1 (N18600, N18581);
or OR3 (N18601, N18595, N17957, N16405);
nand NAND2 (N18602, N18582, N723);
or OR3 (N18603, N18599, N3795, N10050);
xor XOR2 (N18604, N18593, N1335);
not NOT1 (N18605, N18603);
or OR3 (N18606, N18604, N5517, N5832);
xor XOR2 (N18607, N18606, N1273);
buf BUF1 (N18608, N18598);
nor NOR2 (N18609, N18589, N3353);
xor XOR2 (N18610, N18605, N6828);
not NOT1 (N18611, N18602);
or OR2 (N18612, N18597, N4042);
buf BUF1 (N18613, N18609);
buf BUF1 (N18614, N18592);
nand NAND2 (N18615, N18613, N15171);
nand NAND2 (N18616, N18608, N10004);
buf BUF1 (N18617, N18615);
or OR3 (N18618, N18616, N1335, N7435);
and AND4 (N18619, N18618, N2162, N14877, N8605);
buf BUF1 (N18620, N18611);
and AND2 (N18621, N18607, N1618);
nor NOR4 (N18622, N18614, N9882, N10983, N1225);
and AND4 (N18623, N18617, N2617, N10235, N12849);
xor XOR2 (N18624, N18590, N3224);
xor XOR2 (N18625, N18600, N1633);
buf BUF1 (N18626, N18601);
nor NOR4 (N18627, N18624, N3206, N12226, N4562);
or OR2 (N18628, N18620, N18476);
xor XOR2 (N18629, N18622, N17277);
not NOT1 (N18630, N18612);
not NOT1 (N18631, N18627);
and AND4 (N18632, N18621, N16741, N13936, N17298);
nand NAND2 (N18633, N18610, N11013);
xor XOR2 (N18634, N18631, N14166);
and AND3 (N18635, N18633, N6784, N9787);
nand NAND2 (N18636, N18628, N17722);
or OR2 (N18637, N18634, N11102);
or OR3 (N18638, N18630, N6963, N17827);
buf BUF1 (N18639, N18626);
buf BUF1 (N18640, N18619);
buf BUF1 (N18641, N18629);
xor XOR2 (N18642, N18632, N8521);
nor NOR4 (N18643, N18635, N14496, N16006, N9141);
or OR4 (N18644, N18623, N1028, N5418, N4848);
xor XOR2 (N18645, N18638, N5424);
or OR2 (N18646, N18643, N14132);
buf BUF1 (N18647, N18637);
nand NAND2 (N18648, N18641, N10746);
xor XOR2 (N18649, N18636, N10708);
not NOT1 (N18650, N18639);
not NOT1 (N18651, N18647);
or OR2 (N18652, N18649, N1156);
and AND4 (N18653, N18648, N214, N3851, N16113);
or OR2 (N18654, N18646, N13966);
nor NOR3 (N18655, N18640, N3672, N10620);
nor NOR4 (N18656, N18645, N4990, N6516, N17697);
buf BUF1 (N18657, N18644);
nand NAND2 (N18658, N18642, N13688);
nor NOR3 (N18659, N18655, N16620, N15167);
buf BUF1 (N18660, N18658);
and AND4 (N18661, N18653, N1695, N15927, N14220);
nor NOR3 (N18662, N18657, N1859, N15156);
or OR2 (N18663, N18660, N10804);
not NOT1 (N18664, N18651);
xor XOR2 (N18665, N18659, N16844);
or OR2 (N18666, N18656, N1756);
or OR2 (N18667, N18665, N12134);
and AND4 (N18668, N18663, N15149, N12808, N3451);
not NOT1 (N18669, N18662);
xor XOR2 (N18670, N18650, N1439);
and AND4 (N18671, N18668, N13222, N3938, N807);
buf BUF1 (N18672, N18669);
nor NOR2 (N18673, N18670, N3523);
nor NOR2 (N18674, N18666, N9693);
nand NAND2 (N18675, N18664, N2400);
buf BUF1 (N18676, N18675);
or OR3 (N18677, N18676, N14488, N3879);
xor XOR2 (N18678, N18625, N5433);
xor XOR2 (N18679, N18661, N9152);
nand NAND2 (N18680, N18652, N4474);
xor XOR2 (N18681, N18677, N7086);
nor NOR4 (N18682, N18681, N10259, N9565, N15843);
nor NOR4 (N18683, N18667, N9199, N2191, N5190);
buf BUF1 (N18684, N18654);
xor XOR2 (N18685, N18674, N9500);
and AND3 (N18686, N18682, N7743, N13839);
nor NOR4 (N18687, N18684, N1501, N2212, N14829);
buf BUF1 (N18688, N18673);
buf BUF1 (N18689, N18678);
and AND3 (N18690, N18687, N7804, N15929);
xor XOR2 (N18691, N18686, N6283);
or OR4 (N18692, N18685, N1634, N10569, N6711);
nand NAND3 (N18693, N18680, N11245, N15068);
nor NOR2 (N18694, N18679, N11780);
nor NOR2 (N18695, N18683, N11663);
nor NOR3 (N18696, N18692, N14794, N13170);
and AND4 (N18697, N18689, N2489, N5639, N10830);
not NOT1 (N18698, N18672);
buf BUF1 (N18699, N18694);
buf BUF1 (N18700, N18696);
or OR4 (N18701, N18699, N17723, N14184, N10908);
and AND4 (N18702, N18691, N8228, N12901, N13260);
buf BUF1 (N18703, N18700);
nand NAND4 (N18704, N18698, N8345, N18565, N2203);
nor NOR2 (N18705, N18671, N14836);
or OR4 (N18706, N18697, N14256, N15893, N1260);
not NOT1 (N18707, N18702);
nand NAND2 (N18708, N18693, N18231);
nand NAND2 (N18709, N18701, N12005);
or OR2 (N18710, N18709, N2808);
nand NAND2 (N18711, N18704, N13955);
nor NOR2 (N18712, N18706, N14526);
buf BUF1 (N18713, N18688);
buf BUF1 (N18714, N18711);
nand NAND2 (N18715, N18695, N6890);
xor XOR2 (N18716, N18690, N13695);
nand NAND4 (N18717, N18707, N16496, N2933, N12242);
xor XOR2 (N18718, N18716, N2154);
or OR2 (N18719, N18717, N8947);
or OR3 (N18720, N18714, N18697, N3664);
buf BUF1 (N18721, N18719);
buf BUF1 (N18722, N18715);
or OR3 (N18723, N18722, N17516, N7465);
buf BUF1 (N18724, N18721);
nor NOR2 (N18725, N18718, N10354);
buf BUF1 (N18726, N18723);
nand NAND4 (N18727, N18720, N10667, N13229, N14083);
not NOT1 (N18728, N18710);
xor XOR2 (N18729, N18712, N8416);
buf BUF1 (N18730, N18713);
or OR2 (N18731, N18727, N1327);
not NOT1 (N18732, N18725);
nand NAND2 (N18733, N18724, N8199);
xor XOR2 (N18734, N18703, N6348);
nand NAND2 (N18735, N18734, N18426);
nand NAND3 (N18736, N18730, N16969, N9968);
nand NAND4 (N18737, N18708, N11467, N6763, N18633);
nand NAND3 (N18738, N18732, N5864, N2320);
not NOT1 (N18739, N18736);
or OR2 (N18740, N18733, N15351);
nor NOR2 (N18741, N18705, N7536);
not NOT1 (N18742, N18737);
nor NOR4 (N18743, N18728, N12578, N10810, N5385);
nor NOR2 (N18744, N18740, N8672);
xor XOR2 (N18745, N18741, N2093);
or OR3 (N18746, N18735, N1228, N16731);
nor NOR3 (N18747, N18726, N18690, N7860);
or OR3 (N18748, N18745, N16002, N14244);
and AND3 (N18749, N18742, N13011, N16825);
or OR2 (N18750, N18744, N17701);
nor NOR2 (N18751, N18748, N2521);
nand NAND3 (N18752, N18729, N15304, N13659);
nor NOR2 (N18753, N18752, N3344);
xor XOR2 (N18754, N18753, N11535);
or OR2 (N18755, N18754, N3370);
not NOT1 (N18756, N18743);
nand NAND3 (N18757, N18746, N12440, N12394);
xor XOR2 (N18758, N18738, N10351);
and AND4 (N18759, N18757, N17568, N3639, N8535);
buf BUF1 (N18760, N18749);
not NOT1 (N18761, N18760);
or OR3 (N18762, N18761, N4090, N10505);
buf BUF1 (N18763, N18751);
or OR4 (N18764, N18750, N3882, N14247, N14468);
and AND4 (N18765, N18758, N12274, N13269, N9404);
nand NAND3 (N18766, N18755, N16901, N9856);
nor NOR4 (N18767, N18759, N8970, N5990, N9088);
nand NAND2 (N18768, N18763, N2131);
nor NOR2 (N18769, N18739, N14508);
xor XOR2 (N18770, N18747, N17733);
not NOT1 (N18771, N18770);
nand NAND4 (N18772, N18768, N13412, N7812, N2106);
buf BUF1 (N18773, N18766);
nand NAND4 (N18774, N18773, N16943, N13151, N13762);
buf BUF1 (N18775, N18772);
and AND4 (N18776, N18762, N9455, N1238, N15969);
not NOT1 (N18777, N18775);
xor XOR2 (N18778, N18731, N5777);
buf BUF1 (N18779, N18756);
nor NOR3 (N18780, N18765, N8908, N1027);
or OR2 (N18781, N18767, N2540);
nor NOR3 (N18782, N18781, N7903, N9844);
xor XOR2 (N18783, N18769, N9590);
xor XOR2 (N18784, N18777, N12569);
and AND2 (N18785, N18784, N17544);
xor XOR2 (N18786, N18778, N10965);
not NOT1 (N18787, N18786);
xor XOR2 (N18788, N18764, N18473);
buf BUF1 (N18789, N18774);
nand NAND3 (N18790, N18783, N4694, N9291);
not NOT1 (N18791, N18771);
not NOT1 (N18792, N18776);
not NOT1 (N18793, N18790);
nor NOR4 (N18794, N18789, N2524, N17342, N16998);
not NOT1 (N18795, N18780);
buf BUF1 (N18796, N18793);
or OR4 (N18797, N18782, N5745, N12453, N1317);
not NOT1 (N18798, N18791);
or OR4 (N18799, N18785, N1188, N10634, N3371);
nand NAND2 (N18800, N18799, N16053);
buf BUF1 (N18801, N18792);
xor XOR2 (N18802, N18787, N16355);
not NOT1 (N18803, N18794);
nand NAND2 (N18804, N18803, N6357);
xor XOR2 (N18805, N18779, N5815);
or OR3 (N18806, N18800, N11712, N14121);
nor NOR3 (N18807, N18788, N13907, N8181);
and AND3 (N18808, N18796, N9316, N1123);
xor XOR2 (N18809, N18797, N4880);
nand NAND4 (N18810, N18804, N13158, N18122, N9552);
buf BUF1 (N18811, N18806);
buf BUF1 (N18812, N18811);
xor XOR2 (N18813, N18807, N17020);
and AND3 (N18814, N18798, N14033, N12303);
and AND4 (N18815, N18808, N105, N17091, N14878);
xor XOR2 (N18816, N18810, N9917);
buf BUF1 (N18817, N18815);
and AND4 (N18818, N18817, N6778, N8710, N9809);
and AND2 (N18819, N18805, N11090);
or OR2 (N18820, N18814, N10263);
buf BUF1 (N18821, N18813);
xor XOR2 (N18822, N18795, N16111);
or OR2 (N18823, N18819, N18684);
xor XOR2 (N18824, N18820, N18164);
buf BUF1 (N18825, N18802);
xor XOR2 (N18826, N18821, N3380);
nor NOR2 (N18827, N18801, N9711);
buf BUF1 (N18828, N18816);
nor NOR2 (N18829, N18827, N3838);
and AND2 (N18830, N18826, N1321);
or OR3 (N18831, N18823, N10949, N17887);
and AND3 (N18832, N18829, N7840, N8062);
and AND3 (N18833, N18824, N9319, N7555);
nor NOR3 (N18834, N18830, N15188, N17708);
xor XOR2 (N18835, N18812, N7382);
nor NOR2 (N18836, N18834, N416);
or OR3 (N18837, N18828, N14082, N11245);
nand NAND2 (N18838, N18825, N5888);
not NOT1 (N18839, N18809);
buf BUF1 (N18840, N18836);
buf BUF1 (N18841, N18833);
buf BUF1 (N18842, N18832);
nand NAND2 (N18843, N18822, N14728);
xor XOR2 (N18844, N18842, N5782);
not NOT1 (N18845, N18837);
buf BUF1 (N18846, N18838);
buf BUF1 (N18847, N18843);
not NOT1 (N18848, N18844);
nand NAND2 (N18849, N18839, N7422);
xor XOR2 (N18850, N18845, N200);
nand NAND2 (N18851, N18841, N10222);
xor XOR2 (N18852, N18850, N13331);
buf BUF1 (N18853, N18846);
nand NAND4 (N18854, N18851, N5387, N15133, N4185);
or OR2 (N18855, N18835, N3146);
xor XOR2 (N18856, N18852, N16302);
nor NOR3 (N18857, N18840, N13320, N14374);
and AND2 (N18858, N18856, N5672);
xor XOR2 (N18859, N18849, N12213);
xor XOR2 (N18860, N18855, N1471);
xor XOR2 (N18861, N18857, N5791);
not NOT1 (N18862, N18848);
nor NOR2 (N18863, N18858, N210);
xor XOR2 (N18864, N18862, N6183);
nand NAND3 (N18865, N18853, N9145, N12251);
xor XOR2 (N18866, N18863, N1668);
or OR3 (N18867, N18831, N4637, N11219);
buf BUF1 (N18868, N18847);
nor NOR2 (N18869, N18865, N6192);
xor XOR2 (N18870, N18818, N1780);
or OR2 (N18871, N18867, N4649);
nor NOR2 (N18872, N18864, N10537);
or OR3 (N18873, N18854, N2968, N15718);
and AND3 (N18874, N18860, N18271, N7807);
or OR2 (N18875, N18866, N1380);
xor XOR2 (N18876, N18872, N16270);
xor XOR2 (N18877, N18861, N1339);
buf BUF1 (N18878, N18877);
not NOT1 (N18879, N18874);
nand NAND2 (N18880, N18859, N5375);
nand NAND3 (N18881, N18870, N5473, N3456);
or OR2 (N18882, N18871, N9551);
nor NOR2 (N18883, N18881, N6008);
buf BUF1 (N18884, N18878);
or OR2 (N18885, N18884, N6827);
not NOT1 (N18886, N18883);
not NOT1 (N18887, N18869);
nor NOR2 (N18888, N18882, N8156);
buf BUF1 (N18889, N18876);
not NOT1 (N18890, N18873);
buf BUF1 (N18891, N18886);
and AND2 (N18892, N18887, N5350);
nor NOR4 (N18893, N18892, N14403, N10439, N9095);
not NOT1 (N18894, N18879);
or OR3 (N18895, N18880, N13735, N1868);
not NOT1 (N18896, N18889);
not NOT1 (N18897, N18891);
not NOT1 (N18898, N18888);
and AND3 (N18899, N18890, N4277, N13696);
not NOT1 (N18900, N18895);
not NOT1 (N18901, N18894);
not NOT1 (N18902, N18885);
xor XOR2 (N18903, N18896, N12640);
nand NAND2 (N18904, N18868, N6765);
and AND3 (N18905, N18899, N15753, N4208);
nor NOR2 (N18906, N18893, N16337);
and AND4 (N18907, N18906, N8250, N952, N14085);
and AND2 (N18908, N18905, N12314);
nor NOR2 (N18909, N18907, N4155);
or OR2 (N18910, N18900, N18891);
buf BUF1 (N18911, N18903);
buf BUF1 (N18912, N18901);
buf BUF1 (N18913, N18902);
or OR2 (N18914, N18911, N6771);
nand NAND4 (N18915, N18912, N8835, N1598, N4594);
buf BUF1 (N18916, N18913);
not NOT1 (N18917, N18875);
nor NOR3 (N18918, N18904, N5086, N1908);
nor NOR3 (N18919, N18910, N17368, N11223);
buf BUF1 (N18920, N18919);
nor NOR3 (N18921, N18914, N4388, N7234);
not NOT1 (N18922, N18916);
and AND2 (N18923, N18908, N5657);
and AND4 (N18924, N18918, N1094, N8137, N6401);
nor NOR2 (N18925, N18917, N8272);
and AND4 (N18926, N18909, N15632, N11508, N1121);
not NOT1 (N18927, N18915);
or OR4 (N18928, N18897, N3974, N18013, N7215);
nor NOR3 (N18929, N18926, N1553, N14056);
buf BUF1 (N18930, N18920);
not NOT1 (N18931, N18923);
buf BUF1 (N18932, N18898);
nand NAND4 (N18933, N18929, N6401, N5268, N11130);
nor NOR3 (N18934, N18932, N14001, N5814);
xor XOR2 (N18935, N18931, N12805);
nand NAND3 (N18936, N18934, N18337, N1176);
buf BUF1 (N18937, N18922);
nor NOR2 (N18938, N18937, N12228);
buf BUF1 (N18939, N18921);
nand NAND4 (N18940, N18935, N4019, N12609, N15959);
buf BUF1 (N18941, N18933);
nand NAND4 (N18942, N18925, N4003, N10846, N7239);
or OR3 (N18943, N18938, N7025, N9140);
not NOT1 (N18944, N18940);
buf BUF1 (N18945, N18941);
not NOT1 (N18946, N18936);
and AND2 (N18947, N18944, N10696);
not NOT1 (N18948, N18942);
nand NAND2 (N18949, N18945, N5816);
nor NOR3 (N18950, N18943, N16995, N7693);
xor XOR2 (N18951, N18928, N898);
buf BUF1 (N18952, N18950);
nand NAND2 (N18953, N18927, N6365);
nand NAND2 (N18954, N18951, N14374);
buf BUF1 (N18955, N18948);
nor NOR3 (N18956, N18953, N16259, N3201);
buf BUF1 (N18957, N18952);
nand NAND4 (N18958, N18954, N14937, N10265, N9661);
buf BUF1 (N18959, N18957);
nand NAND2 (N18960, N18959, N15131);
not NOT1 (N18961, N18955);
nand NAND3 (N18962, N18949, N724, N15667);
nand NAND4 (N18963, N18956, N4547, N12737, N16824);
or OR3 (N18964, N18930, N14236, N18220);
and AND2 (N18965, N18960, N16687);
nand NAND2 (N18966, N18965, N13413);
xor XOR2 (N18967, N18958, N14889);
not NOT1 (N18968, N18967);
and AND3 (N18969, N18963, N499, N4695);
buf BUF1 (N18970, N18962);
buf BUF1 (N18971, N18961);
xor XOR2 (N18972, N18971, N14974);
nor NOR3 (N18973, N18972, N3413, N3757);
buf BUF1 (N18974, N18964);
nor NOR4 (N18975, N18973, N16787, N13303, N9443);
xor XOR2 (N18976, N18924, N16650);
xor XOR2 (N18977, N18966, N2242);
buf BUF1 (N18978, N18947);
and AND2 (N18979, N18969, N13187);
nand NAND3 (N18980, N18975, N433, N18030);
nor NOR3 (N18981, N18970, N14160, N17198);
or OR3 (N18982, N18974, N13750, N12452);
or OR2 (N18983, N18939, N6796);
nand NAND2 (N18984, N18946, N18033);
buf BUF1 (N18985, N18982);
nor NOR2 (N18986, N18979, N16185);
or OR4 (N18987, N18980, N467, N8576, N14694);
or OR4 (N18988, N18968, N17668, N1307, N6858);
nor NOR3 (N18989, N18976, N10782, N5617);
nor NOR2 (N18990, N18985, N1582);
nor NOR4 (N18991, N18983, N8936, N9015, N6855);
or OR2 (N18992, N18981, N15684);
nor NOR3 (N18993, N18989, N15498, N12085);
not NOT1 (N18994, N18988);
buf BUF1 (N18995, N18978);
nand NAND3 (N18996, N18977, N4726, N6020);
or OR4 (N18997, N18994, N16791, N6642, N10942);
buf BUF1 (N18998, N18984);
not NOT1 (N18999, N18996);
nor NOR4 (N19000, N18990, N12253, N5344, N17202);
not NOT1 (N19001, N18999);
xor XOR2 (N19002, N18995, N12297);
and AND3 (N19003, N18986, N4251, N18771);
nor NOR4 (N19004, N18992, N11817, N9100, N2723);
nand NAND4 (N19005, N18991, N16550, N18760, N8166);
xor XOR2 (N19006, N18987, N6287);
buf BUF1 (N19007, N19002);
nor NOR2 (N19008, N19000, N13034);
and AND3 (N19009, N18997, N3178, N2437);
nor NOR3 (N19010, N18998, N13704, N4562);
or OR3 (N19011, N19007, N14890, N6481);
or OR3 (N19012, N19003, N12077, N9850);
and AND2 (N19013, N19008, N1484);
or OR3 (N19014, N19005, N15615, N5539);
nor NOR3 (N19015, N19014, N7538, N40);
or OR3 (N19016, N19013, N4610, N11671);
or OR3 (N19017, N19006, N2861, N14328);
or OR2 (N19018, N19017, N18846);
or OR2 (N19019, N19004, N18457);
or OR4 (N19020, N18993, N9269, N3849, N16213);
not NOT1 (N19021, N19001);
buf BUF1 (N19022, N19009);
xor XOR2 (N19023, N19015, N2287);
or OR4 (N19024, N19010, N17667, N9204, N13845);
buf BUF1 (N19025, N19020);
buf BUF1 (N19026, N19016);
xor XOR2 (N19027, N19022, N6257);
nand NAND4 (N19028, N19011, N13380, N14028, N6456);
and AND4 (N19029, N19012, N10321, N1540, N408);
xor XOR2 (N19030, N19025, N13148);
nand NAND4 (N19031, N19024, N7668, N7562, N7451);
xor XOR2 (N19032, N19021, N17252);
and AND3 (N19033, N19032, N5694, N7786);
xor XOR2 (N19034, N19018, N6555);
not NOT1 (N19035, N19033);
or OR4 (N19036, N19031, N16075, N9190, N18931);
not NOT1 (N19037, N19030);
nor NOR4 (N19038, N19023, N2301, N18644, N18208);
xor XOR2 (N19039, N19036, N5339);
buf BUF1 (N19040, N19029);
nor NOR2 (N19041, N19039, N4752);
and AND3 (N19042, N19040, N12015, N5492);
and AND2 (N19043, N19034, N6284);
nand NAND3 (N19044, N19037, N6205, N11804);
nand NAND2 (N19045, N19028, N5901);
and AND4 (N19046, N19042, N972, N7482, N5111);
xor XOR2 (N19047, N19043, N5467);
or OR3 (N19048, N19046, N18057, N6384);
or OR4 (N19049, N19027, N7046, N18994, N6376);
nand NAND4 (N19050, N19047, N10137, N17692, N15172);
xor XOR2 (N19051, N19035, N10349);
and AND4 (N19052, N19038, N12295, N13691, N17663);
nand NAND4 (N19053, N19041, N3677, N9124, N10233);
nand NAND3 (N19054, N19049, N3817, N3930);
or OR4 (N19055, N19019, N6425, N16070, N9871);
not NOT1 (N19056, N19052);
xor XOR2 (N19057, N19053, N11056);
buf BUF1 (N19058, N19057);
buf BUF1 (N19059, N19056);
not NOT1 (N19060, N19026);
and AND4 (N19061, N19048, N15714, N190, N8583);
nand NAND3 (N19062, N19059, N9811, N3969);
nand NAND3 (N19063, N19060, N5259, N12651);
not NOT1 (N19064, N19062);
buf BUF1 (N19065, N19055);
not NOT1 (N19066, N19044);
xor XOR2 (N19067, N19065, N17290);
and AND3 (N19068, N19058, N5240, N14630);
buf BUF1 (N19069, N19054);
xor XOR2 (N19070, N19064, N13751);
buf BUF1 (N19071, N19050);
or OR4 (N19072, N19067, N11814, N14701, N7091);
or OR4 (N19073, N19068, N11280, N9709, N7251);
xor XOR2 (N19074, N19071, N16849);
buf BUF1 (N19075, N19070);
not NOT1 (N19076, N19051);
xor XOR2 (N19077, N19061, N235);
not NOT1 (N19078, N19074);
buf BUF1 (N19079, N19066);
xor XOR2 (N19080, N19045, N14279);
not NOT1 (N19081, N19075);
or OR2 (N19082, N19079, N6338);
xor XOR2 (N19083, N19076, N13938);
buf BUF1 (N19084, N19063);
xor XOR2 (N19085, N19073, N12774);
xor XOR2 (N19086, N19080, N16162);
buf BUF1 (N19087, N19084);
not NOT1 (N19088, N19072);
or OR3 (N19089, N19082, N12650, N7146);
nand NAND4 (N19090, N19086, N11477, N17891, N8221);
xor XOR2 (N19091, N19090, N3381);
xor XOR2 (N19092, N19087, N7666);
xor XOR2 (N19093, N19078, N13564);
nand NAND2 (N19094, N19089, N3944);
xor XOR2 (N19095, N19085, N16418);
or OR4 (N19096, N19069, N19057, N2930, N17761);
nor NOR3 (N19097, N19092, N4467, N16003);
or OR4 (N19098, N19096, N14770, N3010, N9527);
or OR4 (N19099, N19094, N552, N7385, N8523);
xor XOR2 (N19100, N19077, N14279);
xor XOR2 (N19101, N19097, N14771);
and AND3 (N19102, N19100, N3428, N16982);
nand NAND3 (N19103, N19102, N16477, N16744);
not NOT1 (N19104, N19103);
or OR4 (N19105, N19081, N17364, N9366, N3740);
nor NOR4 (N19106, N19101, N7486, N8377, N4306);
buf BUF1 (N19107, N19105);
xor XOR2 (N19108, N19083, N18970);
buf BUF1 (N19109, N19099);
nor NOR4 (N19110, N19095, N15666, N13525, N2964);
and AND3 (N19111, N19110, N16956, N12560);
nand NAND2 (N19112, N19106, N4396);
nand NAND4 (N19113, N19093, N8392, N12830, N7865);
or OR2 (N19114, N19111, N15611);
xor XOR2 (N19115, N19114, N4084);
or OR3 (N19116, N19115, N2728, N8644);
nand NAND2 (N19117, N19116, N1634);
nor NOR2 (N19118, N19113, N13209);
or OR3 (N19119, N19118, N9578, N5943);
nor NOR3 (N19120, N19108, N15863, N592);
nand NAND4 (N19121, N19104, N7545, N824, N17063);
xor XOR2 (N19122, N19121, N12889);
nand NAND3 (N19123, N19117, N14929, N8163);
nor NOR3 (N19124, N19119, N13911, N7099);
nand NAND4 (N19125, N19109, N3521, N4508, N3976);
buf BUF1 (N19126, N19122);
buf BUF1 (N19127, N19123);
or OR4 (N19128, N19124, N1918, N5069, N5491);
not NOT1 (N19129, N19128);
nand NAND3 (N19130, N19126, N16499, N14233);
xor XOR2 (N19131, N19127, N16141);
nor NOR4 (N19132, N19098, N18004, N1823, N9278);
nand NAND4 (N19133, N19112, N8381, N17317, N2505);
or OR4 (N19134, N19091, N1255, N1658, N10673);
nor NOR3 (N19135, N19107, N10982, N6594);
nand NAND3 (N19136, N19131, N5906, N13796);
not NOT1 (N19137, N19125);
buf BUF1 (N19138, N19088);
xor XOR2 (N19139, N19133, N886);
not NOT1 (N19140, N19138);
nor NOR2 (N19141, N19136, N14687);
nor NOR2 (N19142, N19137, N16005);
and AND2 (N19143, N19135, N15666);
and AND2 (N19144, N19132, N17195);
xor XOR2 (N19145, N19142, N14001);
or OR3 (N19146, N19145, N5047, N14570);
nand NAND3 (N19147, N19146, N12053, N13134);
buf BUF1 (N19148, N19141);
nor NOR4 (N19149, N19129, N16174, N4045, N1392);
not NOT1 (N19150, N19134);
buf BUF1 (N19151, N19140);
xor XOR2 (N19152, N19149, N13500);
not NOT1 (N19153, N19130);
and AND2 (N19154, N19143, N18469);
or OR3 (N19155, N19154, N6722, N15576);
and AND3 (N19156, N19148, N4255, N1914);
xor XOR2 (N19157, N19139, N11054);
buf BUF1 (N19158, N19152);
nand NAND4 (N19159, N19157, N408, N15557, N15226);
not NOT1 (N19160, N19153);
and AND2 (N19161, N19151, N17067);
nor NOR4 (N19162, N19160, N14025, N16250, N8741);
or OR3 (N19163, N19120, N914, N10216);
nor NOR4 (N19164, N19150, N10768, N2353, N6069);
or OR2 (N19165, N19161, N1713);
not NOT1 (N19166, N19158);
nor NOR2 (N19167, N19166, N18099);
or OR4 (N19168, N19162, N3946, N732, N6887);
not NOT1 (N19169, N19168);
nand NAND4 (N19170, N19159, N1127, N8440, N12827);
nand NAND2 (N19171, N19167, N12156);
not NOT1 (N19172, N19169);
or OR3 (N19173, N19144, N890, N7659);
nand NAND2 (N19174, N19173, N6165);
buf BUF1 (N19175, N19147);
or OR4 (N19176, N19175, N1818, N18132, N8147);
nand NAND3 (N19177, N19170, N8652, N17168);
buf BUF1 (N19178, N19177);
or OR3 (N19179, N19172, N5574, N16505);
and AND2 (N19180, N19163, N1402);
or OR2 (N19181, N19156, N6672);
nand NAND2 (N19182, N19178, N11399);
xor XOR2 (N19183, N19174, N16818);
nor NOR4 (N19184, N19176, N5645, N13017, N5328);
nand NAND3 (N19185, N19164, N17664, N14551);
nand NAND2 (N19186, N19182, N13250);
and AND3 (N19187, N19186, N17928, N12080);
not NOT1 (N19188, N19179);
and AND3 (N19189, N19155, N2526, N1822);
or OR2 (N19190, N19180, N11926);
buf BUF1 (N19191, N19187);
nand NAND3 (N19192, N19183, N10895, N2906);
and AND3 (N19193, N19184, N6318, N15405);
nand NAND4 (N19194, N19165, N17792, N8455, N18068);
buf BUF1 (N19195, N19193);
buf BUF1 (N19196, N19189);
and AND3 (N19197, N19190, N1397, N4880);
xor XOR2 (N19198, N19192, N8277);
or OR2 (N19199, N19197, N19109);
buf BUF1 (N19200, N19199);
xor XOR2 (N19201, N19188, N13472);
xor XOR2 (N19202, N19181, N5322);
nand NAND3 (N19203, N19200, N10423, N10973);
not NOT1 (N19204, N19171);
or OR3 (N19205, N19198, N1948, N7694);
xor XOR2 (N19206, N19202, N15331);
xor XOR2 (N19207, N19203, N13779);
buf BUF1 (N19208, N19204);
and AND3 (N19209, N19194, N18083, N3923);
nand NAND3 (N19210, N19196, N4139, N771);
nor NOR4 (N19211, N19207, N14370, N1377, N14118);
not NOT1 (N19212, N19185);
and AND2 (N19213, N19195, N16207);
nor NOR3 (N19214, N19210, N13564, N12456);
nor NOR3 (N19215, N19209, N10772, N4883);
nor NOR4 (N19216, N19215, N15393, N3651, N12191);
buf BUF1 (N19217, N19213);
nor NOR4 (N19218, N19191, N10606, N18644, N15544);
or OR2 (N19219, N19205, N10288);
nand NAND3 (N19220, N19212, N1657, N8130);
nor NOR3 (N19221, N19208, N14392, N12629);
not NOT1 (N19222, N19219);
and AND4 (N19223, N19222, N8477, N15125, N11013);
buf BUF1 (N19224, N19221);
xor XOR2 (N19225, N19217, N815);
or OR4 (N19226, N19216, N1714, N10496, N5419);
not NOT1 (N19227, N19220);
nand NAND4 (N19228, N19201, N17684, N16684, N18239);
or OR4 (N19229, N19206, N10443, N17365, N1148);
nor NOR3 (N19230, N19225, N124, N18232);
and AND2 (N19231, N19214, N13312);
not NOT1 (N19232, N19231);
not NOT1 (N19233, N19218);
buf BUF1 (N19234, N19229);
not NOT1 (N19235, N19228);
buf BUF1 (N19236, N19230);
and AND3 (N19237, N19235, N7936, N17093);
xor XOR2 (N19238, N19237, N6444);
buf BUF1 (N19239, N19224);
and AND2 (N19240, N19239, N3531);
nand NAND3 (N19241, N19234, N15961, N636);
xor XOR2 (N19242, N19241, N10026);
or OR3 (N19243, N19227, N8637, N9127);
xor XOR2 (N19244, N19232, N18456);
and AND2 (N19245, N19243, N5585);
nor NOR3 (N19246, N19233, N10252, N11608);
nand NAND3 (N19247, N19238, N16286, N102);
buf BUF1 (N19248, N19236);
nor NOR2 (N19249, N19240, N992);
xor XOR2 (N19250, N19223, N869);
nor NOR3 (N19251, N19250, N1667, N17945);
nand NAND4 (N19252, N19249, N6195, N8519, N13801);
and AND3 (N19253, N19247, N11458, N6363);
or OR4 (N19254, N19251, N4361, N5976, N14389);
and AND4 (N19255, N19245, N12432, N6282, N1911);
xor XOR2 (N19256, N19248, N3389);
nand NAND2 (N19257, N19211, N471);
buf BUF1 (N19258, N19253);
xor XOR2 (N19259, N19246, N9623);
or OR4 (N19260, N19255, N14174, N896, N16050);
and AND3 (N19261, N19257, N11504, N18552);
or OR3 (N19262, N19256, N2778, N10030);
not NOT1 (N19263, N19261);
or OR4 (N19264, N19254, N8169, N9033, N1789);
not NOT1 (N19265, N19258);
buf BUF1 (N19266, N19264);
xor XOR2 (N19267, N19263, N9597);
xor XOR2 (N19268, N19265, N17041);
buf BUF1 (N19269, N19244);
or OR3 (N19270, N19262, N11642, N14085);
not NOT1 (N19271, N19268);
or OR4 (N19272, N19269, N12638, N24, N2751);
nor NOR4 (N19273, N19260, N452, N1456, N14327);
or OR2 (N19274, N19242, N8632);
xor XOR2 (N19275, N19271, N8622);
not NOT1 (N19276, N19275);
and AND3 (N19277, N19276, N16707, N5214);
nand NAND2 (N19278, N19273, N7071);
and AND2 (N19279, N19277, N19162);
not NOT1 (N19280, N19266);
buf BUF1 (N19281, N19270);
and AND4 (N19282, N19279, N18484, N2803, N14328);
nor NOR4 (N19283, N19282, N2970, N15614, N5100);
buf BUF1 (N19284, N19252);
buf BUF1 (N19285, N19283);
and AND2 (N19286, N19278, N5657);
nand NAND3 (N19287, N19285, N388, N6261);
nand NAND2 (N19288, N19259, N12303);
nor NOR3 (N19289, N19287, N1664, N15597);
not NOT1 (N19290, N19286);
buf BUF1 (N19291, N19267);
not NOT1 (N19292, N19281);
or OR3 (N19293, N19284, N17021, N1885);
and AND2 (N19294, N19280, N16800);
buf BUF1 (N19295, N19290);
not NOT1 (N19296, N19274);
nor NOR2 (N19297, N19291, N4540);
buf BUF1 (N19298, N19289);
not NOT1 (N19299, N19296);
xor XOR2 (N19300, N19297, N8487);
nand NAND2 (N19301, N19293, N14448);
xor XOR2 (N19302, N19301, N16870);
buf BUF1 (N19303, N19226);
nor NOR3 (N19304, N19294, N16735, N15720);
nand NAND4 (N19305, N19272, N17082, N2137, N8212);
and AND2 (N19306, N19302, N11904);
or OR2 (N19307, N19305, N11308);
not NOT1 (N19308, N19303);
buf BUF1 (N19309, N19300);
or OR3 (N19310, N19306, N8698, N1539);
nor NOR2 (N19311, N19304, N4113);
xor XOR2 (N19312, N19309, N11033);
buf BUF1 (N19313, N19308);
xor XOR2 (N19314, N19310, N16292);
nor NOR2 (N19315, N19299, N5524);
nand NAND4 (N19316, N19292, N14750, N7103, N4687);
buf BUF1 (N19317, N19295);
xor XOR2 (N19318, N19311, N11241);
buf BUF1 (N19319, N19317);
and AND3 (N19320, N19315, N9388, N3271);
buf BUF1 (N19321, N19314);
or OR2 (N19322, N19321, N3787);
or OR2 (N19323, N19318, N15401);
not NOT1 (N19324, N19298);
buf BUF1 (N19325, N19313);
and AND4 (N19326, N19323, N5823, N1472, N11605);
or OR2 (N19327, N19324, N13525);
xor XOR2 (N19328, N19312, N390);
or OR2 (N19329, N19327, N6008);
buf BUF1 (N19330, N19328);
nand NAND3 (N19331, N19307, N3449, N15367);
nor NOR2 (N19332, N19331, N11050);
not NOT1 (N19333, N19288);
xor XOR2 (N19334, N19332, N7956);
xor XOR2 (N19335, N19316, N10715);
not NOT1 (N19336, N19326);
xor XOR2 (N19337, N19322, N3441);
nand NAND4 (N19338, N19333, N9530, N3201, N16798);
xor XOR2 (N19339, N19334, N3170);
or OR3 (N19340, N19337, N19184, N11958);
and AND2 (N19341, N19335, N17565);
not NOT1 (N19342, N19329);
buf BUF1 (N19343, N19319);
nor NOR3 (N19344, N19330, N13631, N17389);
or OR2 (N19345, N19336, N3487);
and AND3 (N19346, N19340, N10741, N15468);
or OR2 (N19347, N19320, N6473);
nand NAND4 (N19348, N19343, N18739, N17621, N3183);
and AND2 (N19349, N19346, N10388);
nand NAND3 (N19350, N19325, N18042, N3647);
and AND3 (N19351, N19342, N2862, N16229);
or OR3 (N19352, N19341, N14198, N12106);
nand NAND2 (N19353, N19344, N5314);
not NOT1 (N19354, N19353);
nand NAND3 (N19355, N19348, N1036, N6891);
and AND2 (N19356, N19350, N8331);
nor NOR4 (N19357, N19339, N11643, N13980, N14167);
nand NAND2 (N19358, N19357, N9821);
xor XOR2 (N19359, N19347, N13455);
nor NOR3 (N19360, N19352, N18806, N1449);
or OR2 (N19361, N19351, N14968);
not NOT1 (N19362, N19338);
buf BUF1 (N19363, N19355);
or OR4 (N19364, N19362, N85, N13400, N17803);
buf BUF1 (N19365, N19364);
not NOT1 (N19366, N19363);
xor XOR2 (N19367, N19349, N12240);
nand NAND2 (N19368, N19354, N4410);
nor NOR3 (N19369, N19366, N7583, N8824);
or OR3 (N19370, N19365, N16853, N8636);
nor NOR2 (N19371, N19369, N17857);
buf BUF1 (N19372, N19370);
nand NAND3 (N19373, N19345, N3258, N3995);
and AND3 (N19374, N19371, N15698, N12340);
nand NAND4 (N19375, N19367, N19042, N16161, N7512);
nand NAND2 (N19376, N19361, N10414);
and AND4 (N19377, N19376, N14707, N16710, N11921);
not NOT1 (N19378, N19368);
nor NOR3 (N19379, N19372, N7947, N14566);
xor XOR2 (N19380, N19377, N1866);
and AND2 (N19381, N19375, N1393);
nand NAND3 (N19382, N19356, N3305, N8854);
not NOT1 (N19383, N19382);
buf BUF1 (N19384, N19360);
xor XOR2 (N19385, N19379, N12922);
and AND4 (N19386, N19385, N1550, N12135, N3379);
buf BUF1 (N19387, N19384);
nor NOR4 (N19388, N19387, N475, N8320, N14770);
nor NOR4 (N19389, N19373, N9823, N9533, N13195);
nor NOR3 (N19390, N19388, N14075, N344);
xor XOR2 (N19391, N19389, N74);
buf BUF1 (N19392, N19383);
or OR3 (N19393, N19390, N15256, N8002);
and AND3 (N19394, N19391, N4200, N2642);
nand NAND4 (N19395, N19378, N18299, N5052, N15645);
nor NOR4 (N19396, N19359, N13436, N13791, N5922);
or OR2 (N19397, N19394, N658);
nand NAND2 (N19398, N19358, N2858);
not NOT1 (N19399, N19392);
and AND4 (N19400, N19396, N16567, N14036, N13182);
xor XOR2 (N19401, N19397, N11611);
nor NOR2 (N19402, N19381, N18078);
or OR4 (N19403, N19398, N2101, N2501, N6559);
and AND2 (N19404, N19399, N16801);
xor XOR2 (N19405, N19402, N1225);
nand NAND3 (N19406, N19401, N6650, N13965);
not NOT1 (N19407, N19405);
buf BUF1 (N19408, N19395);
nand NAND3 (N19409, N19406, N6845, N16139);
xor XOR2 (N19410, N19403, N15463);
or OR2 (N19411, N19380, N17865);
and AND3 (N19412, N19409, N492, N18470);
and AND4 (N19413, N19393, N14577, N19080, N10283);
xor XOR2 (N19414, N19411, N15329);
xor XOR2 (N19415, N19414, N5489);
nand NAND4 (N19416, N19404, N10099, N17624, N14417);
nor NOR4 (N19417, N19415, N8857, N14992, N7989);
and AND4 (N19418, N19400, N10097, N3807, N5632);
nor NOR3 (N19419, N19416, N7483, N6189);
not NOT1 (N19420, N19417);
xor XOR2 (N19421, N19412, N538);
or OR4 (N19422, N19419, N671, N7610, N15790);
not NOT1 (N19423, N19418);
and AND4 (N19424, N19374, N2791, N15679, N18239);
nand NAND4 (N19425, N19421, N13140, N11449, N2323);
not NOT1 (N19426, N19410);
and AND3 (N19427, N19425, N7389, N10643);
xor XOR2 (N19428, N19423, N15718);
nand NAND3 (N19429, N19413, N15354, N14866);
and AND2 (N19430, N19422, N12464);
nor NOR2 (N19431, N19386, N4635);
or OR4 (N19432, N19428, N9019, N13223, N16334);
not NOT1 (N19433, N19426);
nand NAND3 (N19434, N19432, N7705, N6361);
or OR2 (N19435, N19430, N11525);
and AND3 (N19436, N19420, N1987, N12941);
not NOT1 (N19437, N19434);
nor NOR4 (N19438, N19424, N5490, N14921, N10041);
and AND2 (N19439, N19438, N2048);
xor XOR2 (N19440, N19437, N16099);
nor NOR4 (N19441, N19427, N2080, N7249, N6798);
nand NAND4 (N19442, N19433, N3229, N7053, N10727);
nand NAND4 (N19443, N19431, N14655, N12345, N12767);
nand NAND2 (N19444, N19408, N2066);
buf BUF1 (N19445, N19429);
or OR4 (N19446, N19439, N17942, N16489, N13910);
xor XOR2 (N19447, N19445, N7171);
buf BUF1 (N19448, N19436);
nor NOR2 (N19449, N19447, N15107);
nor NOR3 (N19450, N19440, N11535, N14232);
and AND3 (N19451, N19443, N1146, N12892);
nand NAND4 (N19452, N19451, N4369, N13283, N6843);
not NOT1 (N19453, N19442);
and AND4 (N19454, N19435, N942, N4564, N2512);
nor NOR2 (N19455, N19452, N2638);
buf BUF1 (N19456, N19455);
and AND3 (N19457, N19446, N10641, N17292);
not NOT1 (N19458, N19407);
not NOT1 (N19459, N19449);
xor XOR2 (N19460, N19441, N449);
or OR2 (N19461, N19456, N5423);
not NOT1 (N19462, N19458);
buf BUF1 (N19463, N19450);
xor XOR2 (N19464, N19461, N15900);
and AND2 (N19465, N19448, N8245);
not NOT1 (N19466, N19463);
nand NAND4 (N19467, N19462, N3983, N18286, N9998);
buf BUF1 (N19468, N19454);
buf BUF1 (N19469, N19460);
nor NOR4 (N19470, N19453, N15191, N16418, N3731);
or OR4 (N19471, N19466, N6953, N6281, N8939);
nor NOR3 (N19472, N19469, N12658, N1242);
not NOT1 (N19473, N19467);
buf BUF1 (N19474, N19459);
and AND3 (N19475, N19457, N1072, N11525);
buf BUF1 (N19476, N19465);
or OR2 (N19477, N19473, N14462);
not NOT1 (N19478, N19474);
or OR4 (N19479, N19444, N18917, N2590, N13414);
and AND2 (N19480, N19478, N18806);
not NOT1 (N19481, N19475);
or OR3 (N19482, N19476, N10004, N6716);
or OR3 (N19483, N19464, N16850, N9376);
nor NOR2 (N19484, N19480, N1984);
not NOT1 (N19485, N19470);
xor XOR2 (N19486, N19477, N1895);
xor XOR2 (N19487, N19482, N1318);
nor NOR2 (N19488, N19486, N4857);
not NOT1 (N19489, N19484);
nand NAND2 (N19490, N19471, N12253);
and AND2 (N19491, N19468, N12543);
nor NOR2 (N19492, N19479, N16335);
buf BUF1 (N19493, N19492);
and AND3 (N19494, N19472, N13963, N5948);
xor XOR2 (N19495, N19483, N17329);
not NOT1 (N19496, N19485);
not NOT1 (N19497, N19488);
buf BUF1 (N19498, N19496);
xor XOR2 (N19499, N19495, N1365);
nand NAND2 (N19500, N19499, N833);
nand NAND2 (N19501, N19493, N10713);
xor XOR2 (N19502, N19481, N17386);
not NOT1 (N19503, N19487);
not NOT1 (N19504, N19502);
or OR2 (N19505, N19491, N7921);
xor XOR2 (N19506, N19504, N14298);
and AND2 (N19507, N19490, N12977);
not NOT1 (N19508, N19500);
nand NAND4 (N19509, N19501, N3805, N11619, N8705);
not NOT1 (N19510, N19505);
and AND4 (N19511, N19498, N16457, N11409, N17121);
nor NOR3 (N19512, N19510, N19028, N3154);
xor XOR2 (N19513, N19506, N18898);
or OR3 (N19514, N19511, N15491, N2148);
nand NAND3 (N19515, N19509, N2302, N17417);
nor NOR3 (N19516, N19512, N10266, N6668);
or OR3 (N19517, N19513, N4484, N7969);
xor XOR2 (N19518, N19508, N5476);
buf BUF1 (N19519, N19517);
not NOT1 (N19520, N19497);
nor NOR2 (N19521, N19520, N13867);
nor NOR2 (N19522, N19494, N8210);
nor NOR4 (N19523, N19515, N19486, N5645, N5578);
nand NAND4 (N19524, N19521, N9489, N4498, N1169);
nor NOR3 (N19525, N19503, N586, N4098);
buf BUF1 (N19526, N19523);
buf BUF1 (N19527, N19526);
buf BUF1 (N19528, N19518);
not NOT1 (N19529, N19489);
not NOT1 (N19530, N19525);
and AND2 (N19531, N19507, N8921);
buf BUF1 (N19532, N19516);
nand NAND3 (N19533, N19530, N17441, N6993);
xor XOR2 (N19534, N19528, N12433);
or OR4 (N19535, N19519, N1519, N8411, N226);
not NOT1 (N19536, N19529);
nor NOR2 (N19537, N19536, N15417);
buf BUF1 (N19538, N19514);
nor NOR3 (N19539, N19527, N15906, N12564);
not NOT1 (N19540, N19535);
buf BUF1 (N19541, N19534);
and AND2 (N19542, N19533, N17315);
or OR3 (N19543, N19538, N17014, N8018);
nor NOR3 (N19544, N19531, N1740, N4303);
and AND3 (N19545, N19524, N2391, N16938);
or OR4 (N19546, N19544, N16389, N677, N858);
not NOT1 (N19547, N19539);
buf BUF1 (N19548, N19546);
not NOT1 (N19549, N19540);
not NOT1 (N19550, N19549);
not NOT1 (N19551, N19542);
not NOT1 (N19552, N19547);
xor XOR2 (N19553, N19545, N6833);
nand NAND4 (N19554, N19548, N9439, N5366, N18830);
nand NAND3 (N19555, N19543, N9933, N13473);
nand NAND4 (N19556, N19532, N6142, N14409, N18098);
and AND4 (N19557, N19554, N15040, N163, N307);
buf BUF1 (N19558, N19556);
buf BUF1 (N19559, N19552);
nand NAND2 (N19560, N19559, N15008);
buf BUF1 (N19561, N19541);
not NOT1 (N19562, N19555);
xor XOR2 (N19563, N19561, N17241);
not NOT1 (N19564, N19560);
and AND4 (N19565, N19564, N13463, N10788, N13431);
nor NOR3 (N19566, N19563, N5669, N8263);
nand NAND3 (N19567, N19551, N12468, N1186);
and AND4 (N19568, N19557, N9295, N3255, N15033);
xor XOR2 (N19569, N19553, N12543);
and AND3 (N19570, N19569, N1327, N11775);
or OR2 (N19571, N19562, N13026);
or OR3 (N19572, N19550, N18256, N5358);
nor NOR3 (N19573, N19565, N2745, N5374);
or OR2 (N19574, N19573, N6443);
buf BUF1 (N19575, N19568);
not NOT1 (N19576, N19571);
xor XOR2 (N19577, N19576, N12335);
or OR2 (N19578, N19570, N16471);
nor NOR2 (N19579, N19575, N3420);
buf BUF1 (N19580, N19577);
nand NAND2 (N19581, N19579, N1066);
nor NOR3 (N19582, N19572, N386, N14360);
not NOT1 (N19583, N19558);
buf BUF1 (N19584, N19580);
not NOT1 (N19585, N19581);
not NOT1 (N19586, N19578);
buf BUF1 (N19587, N19537);
buf BUF1 (N19588, N19586);
nand NAND4 (N19589, N19522, N11644, N18006, N8881);
buf BUF1 (N19590, N19574);
not NOT1 (N19591, N19588);
nor NOR3 (N19592, N19585, N80, N8635);
not NOT1 (N19593, N19589);
not NOT1 (N19594, N19583);
or OR3 (N19595, N19593, N9381, N10293);
and AND2 (N19596, N19590, N15490);
or OR2 (N19597, N19587, N6172);
buf BUF1 (N19598, N19582);
and AND3 (N19599, N19584, N2451, N8479);
buf BUF1 (N19600, N19596);
nor NOR2 (N19601, N19597, N5552);
or OR2 (N19602, N19595, N4280);
nand NAND4 (N19603, N19566, N80, N8624, N15618);
nor NOR3 (N19604, N19567, N19038, N3335);
nor NOR3 (N19605, N19592, N13843, N7991);
not NOT1 (N19606, N19602);
and AND2 (N19607, N19606, N2708);
nand NAND2 (N19608, N19600, N1751);
buf BUF1 (N19609, N19605);
not NOT1 (N19610, N19603);
not NOT1 (N19611, N19608);
or OR2 (N19612, N19599, N13954);
nand NAND4 (N19613, N19612, N16735, N16189, N9265);
nand NAND3 (N19614, N19604, N18150, N2962);
nor NOR4 (N19615, N19601, N5159, N18307, N12165);
xor XOR2 (N19616, N19611, N2764);
or OR4 (N19617, N19609, N16366, N7440, N4362);
nor NOR3 (N19618, N19617, N43, N398);
nand NAND3 (N19619, N19610, N6604, N18211);
and AND3 (N19620, N19618, N15594, N2817);
buf BUF1 (N19621, N19594);
buf BUF1 (N19622, N19619);
not NOT1 (N19623, N19620);
xor XOR2 (N19624, N19607, N8755);
nor NOR2 (N19625, N19598, N16461);
buf BUF1 (N19626, N19622);
xor XOR2 (N19627, N19613, N14179);
buf BUF1 (N19628, N19591);
buf BUF1 (N19629, N19625);
and AND3 (N19630, N19615, N6744, N12291);
nand NAND3 (N19631, N19624, N7789, N3516);
not NOT1 (N19632, N19623);
and AND2 (N19633, N19627, N5213);
xor XOR2 (N19634, N19630, N4998);
not NOT1 (N19635, N19614);
buf BUF1 (N19636, N19621);
nor NOR3 (N19637, N19628, N2914, N4764);
nand NAND4 (N19638, N19633, N16233, N9589, N14875);
not NOT1 (N19639, N19616);
nor NOR4 (N19640, N19635, N6436, N9529, N15145);
and AND3 (N19641, N19632, N5040, N8291);
xor XOR2 (N19642, N19636, N5709);
and AND4 (N19643, N19639, N11064, N13353, N6257);
xor XOR2 (N19644, N19642, N12177);
buf BUF1 (N19645, N19629);
or OR4 (N19646, N19641, N10362, N16688, N5062);
or OR4 (N19647, N19643, N261, N9323, N5155);
not NOT1 (N19648, N19644);
nor NOR2 (N19649, N19648, N1224);
and AND2 (N19650, N19647, N6799);
or OR3 (N19651, N19640, N659, N3314);
or OR2 (N19652, N19650, N12772);
xor XOR2 (N19653, N19631, N9583);
buf BUF1 (N19654, N19645);
and AND3 (N19655, N19638, N6325, N10130);
or OR3 (N19656, N19654, N758, N19095);
xor XOR2 (N19657, N19651, N8138);
nand NAND4 (N19658, N19655, N11751, N3630, N14423);
and AND3 (N19659, N19658, N12761, N9832);
buf BUF1 (N19660, N19652);
buf BUF1 (N19661, N19634);
and AND4 (N19662, N19626, N18808, N7441, N840);
nand NAND4 (N19663, N19659, N13952, N3237, N3272);
xor XOR2 (N19664, N19653, N8628);
nand NAND3 (N19665, N19656, N7555, N3168);
buf BUF1 (N19666, N19657);
xor XOR2 (N19667, N19637, N9429);
and AND2 (N19668, N19649, N17419);
or OR2 (N19669, N19661, N13968);
nor NOR3 (N19670, N19660, N4572, N5356);
not NOT1 (N19671, N19669);
and AND2 (N19672, N19666, N13678);
nor NOR4 (N19673, N19664, N5201, N6229, N15238);
nor NOR2 (N19674, N19673, N3990);
or OR3 (N19675, N19672, N9625, N4497);
xor XOR2 (N19676, N19665, N15126);
nand NAND3 (N19677, N19674, N16914, N2202);
nand NAND2 (N19678, N19668, N10216);
xor XOR2 (N19679, N19670, N14563);
xor XOR2 (N19680, N19678, N11593);
nor NOR2 (N19681, N19676, N10890);
or OR4 (N19682, N19646, N18418, N132, N15013);
nor NOR3 (N19683, N19681, N4255, N18886);
and AND2 (N19684, N19680, N4793);
nand NAND2 (N19685, N19683, N18560);
buf BUF1 (N19686, N19662);
or OR2 (N19687, N19675, N16494);
nor NOR3 (N19688, N19679, N12245, N9629);
not NOT1 (N19689, N19667);
not NOT1 (N19690, N19671);
nor NOR3 (N19691, N19684, N5886, N5901);
or OR4 (N19692, N19690, N5482, N3530, N17907);
and AND2 (N19693, N19687, N7943);
buf BUF1 (N19694, N19689);
and AND4 (N19695, N19694, N14455, N15607, N9007);
buf BUF1 (N19696, N19691);
buf BUF1 (N19697, N19695);
nand NAND4 (N19698, N19677, N14931, N16009, N7901);
nand NAND2 (N19699, N19696, N14199);
buf BUF1 (N19700, N19663);
buf BUF1 (N19701, N19697);
buf BUF1 (N19702, N19688);
nor NOR2 (N19703, N19682, N8850);
not NOT1 (N19704, N19700);
or OR3 (N19705, N19701, N19190, N18391);
or OR3 (N19706, N19704, N13892, N13833);
and AND2 (N19707, N19702, N16113);
buf BUF1 (N19708, N19703);
nor NOR2 (N19709, N19699, N9812);
buf BUF1 (N19710, N19705);
and AND4 (N19711, N19708, N11153, N7014, N4694);
and AND4 (N19712, N19698, N12213, N14066, N4544);
nand NAND3 (N19713, N19686, N8617, N11999);
buf BUF1 (N19714, N19713);
or OR4 (N19715, N19714, N18662, N5851, N59);
nor NOR3 (N19716, N19707, N13855, N17741);
xor XOR2 (N19717, N19710, N2528);
and AND2 (N19718, N19717, N3926);
or OR4 (N19719, N19693, N16286, N6715, N5369);
nand NAND3 (N19720, N19685, N7398, N12311);
and AND4 (N19721, N19692, N4434, N4306, N12638);
not NOT1 (N19722, N19719);
nand NAND4 (N19723, N19718, N17779, N18333, N16448);
and AND2 (N19724, N19716, N3058);
and AND3 (N19725, N19706, N13830, N17813);
buf BUF1 (N19726, N19720);
nand NAND3 (N19727, N19723, N3206, N16040);
or OR4 (N19728, N19724, N588, N12641, N19284);
and AND4 (N19729, N19715, N15497, N14711, N402);
and AND3 (N19730, N19721, N2034, N17537);
not NOT1 (N19731, N19709);
nor NOR2 (N19732, N19722, N4758);
buf BUF1 (N19733, N19727);
xor XOR2 (N19734, N19732, N10291);
nor NOR2 (N19735, N19725, N14037);
and AND4 (N19736, N19712, N1450, N14795, N12086);
and AND3 (N19737, N19711, N11454, N3665);
nand NAND4 (N19738, N19726, N3839, N14966, N1177);
and AND4 (N19739, N19728, N11689, N7996, N1516);
nor NOR2 (N19740, N19737, N2293);
buf BUF1 (N19741, N19735);
xor XOR2 (N19742, N19730, N9234);
not NOT1 (N19743, N19729);
or OR4 (N19744, N19738, N9732, N3314, N3736);
xor XOR2 (N19745, N19743, N8573);
not NOT1 (N19746, N19741);
xor XOR2 (N19747, N19744, N17846);
xor XOR2 (N19748, N19740, N17142);
or OR2 (N19749, N19742, N10164);
and AND4 (N19750, N19746, N11715, N18482, N9133);
xor XOR2 (N19751, N19748, N18204);
buf BUF1 (N19752, N19751);
xor XOR2 (N19753, N19745, N2760);
or OR2 (N19754, N19752, N10892);
buf BUF1 (N19755, N19747);
nand NAND2 (N19756, N19734, N10274);
and AND3 (N19757, N19731, N4419, N15621);
xor XOR2 (N19758, N19754, N16672);
not NOT1 (N19759, N19755);
not NOT1 (N19760, N19750);
not NOT1 (N19761, N19758);
nor NOR2 (N19762, N19759, N11271);
xor XOR2 (N19763, N19756, N2820);
xor XOR2 (N19764, N19757, N663);
nor NOR2 (N19765, N19733, N5587);
buf BUF1 (N19766, N19763);
not NOT1 (N19767, N19761);
nand NAND2 (N19768, N19765, N5780);
nand NAND4 (N19769, N19736, N7580, N935, N7552);
buf BUF1 (N19770, N19767);
nor NOR2 (N19771, N19753, N13764);
or OR2 (N19772, N19760, N8795);
and AND2 (N19773, N19739, N6278);
xor XOR2 (N19774, N19770, N636);
xor XOR2 (N19775, N19772, N7632);
or OR2 (N19776, N19762, N15714);
not NOT1 (N19777, N19775);
nand NAND3 (N19778, N19773, N8634, N7084);
nand NAND2 (N19779, N19749, N18441);
or OR2 (N19780, N19776, N11945);
nor NOR2 (N19781, N19780, N9064);
xor XOR2 (N19782, N19779, N15322);
nand NAND2 (N19783, N19768, N8612);
and AND4 (N19784, N19782, N3709, N17472, N18342);
buf BUF1 (N19785, N19778);
or OR4 (N19786, N19785, N2939, N3991, N19375);
xor XOR2 (N19787, N19783, N15469);
xor XOR2 (N19788, N19774, N16995);
or OR3 (N19789, N19766, N5202, N7076);
buf BUF1 (N19790, N19764);
nand NAND4 (N19791, N19784, N11435, N10966, N13386);
not NOT1 (N19792, N19787);
buf BUF1 (N19793, N19791);
or OR2 (N19794, N19781, N15156);
xor XOR2 (N19795, N19793, N5551);
buf BUF1 (N19796, N19795);
or OR3 (N19797, N19794, N15068, N13435);
not NOT1 (N19798, N19790);
buf BUF1 (N19799, N19792);
nor NOR4 (N19800, N19786, N17180, N482, N8720);
or OR3 (N19801, N19798, N8257, N3883);
not NOT1 (N19802, N19801);
or OR2 (N19803, N19802, N13429);
and AND4 (N19804, N19769, N3042, N19030, N11518);
and AND3 (N19805, N19800, N19134, N10487);
not NOT1 (N19806, N19789);
buf BUF1 (N19807, N19788);
nor NOR3 (N19808, N19771, N14470, N4882);
nand NAND4 (N19809, N19807, N16335, N10297, N11054);
nor NOR3 (N19810, N19797, N3614, N2914);
xor XOR2 (N19811, N19796, N11013);
nor NOR4 (N19812, N19805, N8396, N8509, N16998);
buf BUF1 (N19813, N19808);
not NOT1 (N19814, N19777);
nor NOR3 (N19815, N19799, N11729, N17884);
and AND3 (N19816, N19814, N7017, N2269);
nor NOR2 (N19817, N19813, N13293);
and AND4 (N19818, N19804, N1368, N18322, N463);
not NOT1 (N19819, N19806);
and AND2 (N19820, N19803, N445);
buf BUF1 (N19821, N19817);
not NOT1 (N19822, N19812);
or OR4 (N19823, N19819, N12807, N6927, N18124);
or OR4 (N19824, N19822, N6761, N10176, N496);
buf BUF1 (N19825, N19810);
xor XOR2 (N19826, N19821, N6275);
or OR4 (N19827, N19816, N14802, N10981, N18709);
and AND3 (N19828, N19824, N9574, N5632);
not NOT1 (N19829, N19809);
nand NAND4 (N19830, N19823, N8308, N358, N9212);
not NOT1 (N19831, N19825);
and AND2 (N19832, N19829, N18563);
xor XOR2 (N19833, N19830, N9804);
xor XOR2 (N19834, N19828, N11580);
or OR4 (N19835, N19827, N3901, N13528, N18057);
nand NAND2 (N19836, N19826, N6314);
buf BUF1 (N19837, N19833);
nor NOR4 (N19838, N19834, N8849, N13980, N8888);
xor XOR2 (N19839, N19832, N15190);
or OR4 (N19840, N19831, N17506, N7467, N1372);
nor NOR4 (N19841, N19836, N7356, N7662, N13602);
buf BUF1 (N19842, N19840);
and AND4 (N19843, N19838, N10624, N8221, N10459);
and AND4 (N19844, N19820, N13141, N8367, N9241);
nor NOR2 (N19845, N19842, N13931);
or OR3 (N19846, N19843, N3677, N885);
nor NOR2 (N19847, N19841, N314);
or OR3 (N19848, N19835, N12724, N10286);
not NOT1 (N19849, N19815);
xor XOR2 (N19850, N19849, N3755);
or OR4 (N19851, N19850, N9636, N17444, N13450);
or OR3 (N19852, N19845, N12843, N8934);
nand NAND4 (N19853, N19818, N6140, N18511, N2423);
and AND2 (N19854, N19848, N2388);
buf BUF1 (N19855, N19854);
xor XOR2 (N19856, N19839, N17563);
or OR4 (N19857, N19846, N10377, N16402, N789);
xor XOR2 (N19858, N19844, N14014);
nor NOR4 (N19859, N19837, N16971, N12849, N2311);
nand NAND3 (N19860, N19855, N8771, N9168);
nor NOR3 (N19861, N19856, N16413, N4092);
and AND2 (N19862, N19852, N2042);
nand NAND4 (N19863, N19853, N16573, N10171, N9235);
and AND2 (N19864, N19847, N15633);
or OR2 (N19865, N19862, N8133);
nand NAND4 (N19866, N19860, N3764, N18612, N12480);
nand NAND3 (N19867, N19865, N19230, N16224);
xor XOR2 (N19868, N19857, N4315);
xor XOR2 (N19869, N19863, N3939);
or OR2 (N19870, N19866, N16902);
and AND4 (N19871, N19861, N10804, N14254, N10194);
not NOT1 (N19872, N19868);
and AND3 (N19873, N19872, N17931, N15637);
xor XOR2 (N19874, N19864, N15894);
not NOT1 (N19875, N19870);
nand NAND2 (N19876, N19851, N10202);
or OR4 (N19877, N19876, N8572, N8163, N7489);
not NOT1 (N19878, N19875);
or OR3 (N19879, N19871, N704, N1745);
buf BUF1 (N19880, N19869);
nor NOR2 (N19881, N19858, N7290);
or OR4 (N19882, N19880, N8823, N4756, N17886);
or OR2 (N19883, N19873, N4895);
or OR4 (N19884, N19867, N1112, N1204, N5445);
xor XOR2 (N19885, N19882, N14031);
buf BUF1 (N19886, N19874);
and AND3 (N19887, N19877, N13103, N5278);
nor NOR2 (N19888, N19884, N12884);
not NOT1 (N19889, N19859);
or OR4 (N19890, N19883, N10677, N15610, N4701);
not NOT1 (N19891, N19886);
buf BUF1 (N19892, N19878);
not NOT1 (N19893, N19890);
not NOT1 (N19894, N19887);
buf BUF1 (N19895, N19888);
and AND4 (N19896, N19893, N2077, N19250, N8342);
or OR2 (N19897, N19881, N18398);
xor XOR2 (N19898, N19891, N17710);
xor XOR2 (N19899, N19896, N3764);
and AND4 (N19900, N19898, N19801, N10065, N4712);
not NOT1 (N19901, N19897);
buf BUF1 (N19902, N19895);
xor XOR2 (N19903, N19811, N3476);
buf BUF1 (N19904, N19889);
buf BUF1 (N19905, N19892);
buf BUF1 (N19906, N19901);
not NOT1 (N19907, N19906);
not NOT1 (N19908, N19904);
or OR3 (N19909, N19885, N16454, N8237);
or OR2 (N19910, N19899, N12048);
and AND2 (N19911, N19910, N3767);
not NOT1 (N19912, N19909);
and AND2 (N19913, N19903, N3536);
nand NAND3 (N19914, N19907, N13877, N10840);
nand NAND2 (N19915, N19914, N17876);
or OR3 (N19916, N19915, N6734, N6032);
and AND3 (N19917, N19905, N6000, N5904);
nor NOR2 (N19918, N19894, N7217);
or OR4 (N19919, N19916, N2679, N5997, N6020);
or OR2 (N19920, N19919, N10982);
buf BUF1 (N19921, N19879);
xor XOR2 (N19922, N19913, N9394);
and AND2 (N19923, N19912, N18859);
or OR2 (N19924, N19920, N2799);
buf BUF1 (N19925, N19908);
not NOT1 (N19926, N19917);
not NOT1 (N19927, N19925);
nand NAND3 (N19928, N19926, N9, N16502);
and AND2 (N19929, N19900, N17198);
or OR4 (N19930, N19918, N2905, N9414, N5000);
nor NOR3 (N19931, N19928, N11026, N1210);
not NOT1 (N19932, N19930);
buf BUF1 (N19933, N19927);
not NOT1 (N19934, N19922);
not NOT1 (N19935, N19929);
not NOT1 (N19936, N19935);
and AND3 (N19937, N19924, N5711, N8335);
and AND2 (N19938, N19932, N13341);
or OR2 (N19939, N19911, N11765);
nand NAND3 (N19940, N19921, N13222, N17900);
not NOT1 (N19941, N19938);
not NOT1 (N19942, N19902);
xor XOR2 (N19943, N19934, N7844);
buf BUF1 (N19944, N19931);
not NOT1 (N19945, N19933);
not NOT1 (N19946, N19939);
and AND2 (N19947, N19936, N10061);
nor NOR2 (N19948, N19937, N6116);
nand NAND3 (N19949, N19923, N14661, N10655);
nand NAND3 (N19950, N19941, N6768, N16393);
nor NOR4 (N19951, N19946, N17279, N16001, N823);
and AND4 (N19952, N19942, N11601, N15513, N9173);
and AND4 (N19953, N19949, N16698, N17932, N19486);
xor XOR2 (N19954, N19952, N2775);
and AND4 (N19955, N19940, N10513, N13076, N16657);
not NOT1 (N19956, N19950);
and AND4 (N19957, N19955, N7153, N15224, N7892);
not NOT1 (N19958, N19957);
or OR2 (N19959, N19951, N17714);
not NOT1 (N19960, N19959);
or OR2 (N19961, N19960, N11125);
and AND3 (N19962, N19947, N4340, N1570);
xor XOR2 (N19963, N19944, N13254);
nor NOR4 (N19964, N19953, N17132, N16164, N9973);
not NOT1 (N19965, N19958);
nand NAND2 (N19966, N19954, N10146);
and AND3 (N19967, N19956, N18289, N8190);
nand NAND3 (N19968, N19967, N6209, N18190);
nand NAND3 (N19969, N19943, N15977, N14656);
xor XOR2 (N19970, N19961, N5461);
nand NAND2 (N19971, N19970, N2754);
buf BUF1 (N19972, N19969);
nor NOR3 (N19973, N19972, N14073, N10967);
nand NAND3 (N19974, N19973, N2915, N9735);
buf BUF1 (N19975, N19971);
nor NOR4 (N19976, N19948, N19502, N7592, N3602);
nor NOR3 (N19977, N19945, N13602, N11862);
or OR4 (N19978, N19976, N10147, N16480, N14650);
buf BUF1 (N19979, N19966);
or OR4 (N19980, N19963, N6326, N2815, N11363);
and AND3 (N19981, N19977, N17427, N9569);
and AND2 (N19982, N19978, N4146);
not NOT1 (N19983, N19975);
buf BUF1 (N19984, N19982);
not NOT1 (N19985, N19968);
nor NOR2 (N19986, N19974, N5823);
or OR4 (N19987, N19980, N9654, N14971, N18209);
or OR3 (N19988, N19964, N2450, N5446);
not NOT1 (N19989, N19983);
nor NOR2 (N19990, N19984, N9160);
buf BUF1 (N19991, N19962);
xor XOR2 (N19992, N19989, N2107);
buf BUF1 (N19993, N19981);
not NOT1 (N19994, N19979);
buf BUF1 (N19995, N19988);
not NOT1 (N19996, N19987);
nand NAND4 (N19997, N19996, N10905, N4876, N4674);
xor XOR2 (N19998, N19965, N12578);
not NOT1 (N19999, N19986);
and AND2 (N20000, N19990, N14517);
or OR3 (N20001, N19997, N2443, N4893);
nand NAND4 (N20002, N19999, N8302, N3246, N2564);
or OR3 (N20003, N19993, N18899, N19922);
nand NAND3 (N20004, N19994, N612, N4127);
xor XOR2 (N20005, N20001, N5979);
or OR3 (N20006, N19991, N12042, N12632);
nor NOR2 (N20007, N20006, N8612);
xor XOR2 (N20008, N19998, N8415);
buf BUF1 (N20009, N20007);
nor NOR3 (N20010, N20003, N5971, N15442);
xor XOR2 (N20011, N19995, N6019);
xor XOR2 (N20012, N19992, N15528);
or OR2 (N20013, N20008, N2497);
buf BUF1 (N20014, N20013);
xor XOR2 (N20015, N20012, N4208);
nand NAND4 (N20016, N20015, N14888, N19974, N12386);
buf BUF1 (N20017, N20000);
buf BUF1 (N20018, N20002);
xor XOR2 (N20019, N20018, N16955);
or OR2 (N20020, N20017, N17097);
or OR3 (N20021, N20019, N6760, N8906);
nor NOR4 (N20022, N20010, N4000, N6915, N15077);
nor NOR2 (N20023, N20022, N8544);
nand NAND2 (N20024, N20014, N5518);
or OR3 (N20025, N19985, N7275, N158);
xor XOR2 (N20026, N20009, N19852);
buf BUF1 (N20027, N20020);
not NOT1 (N20028, N20025);
buf BUF1 (N20029, N20027);
xor XOR2 (N20030, N20026, N6255);
not NOT1 (N20031, N20005);
and AND3 (N20032, N20021, N7693, N17115);
and AND3 (N20033, N20024, N1870, N20010);
nand NAND4 (N20034, N20033, N17226, N15038, N4852);
buf BUF1 (N20035, N20029);
and AND2 (N20036, N20016, N6725);
xor XOR2 (N20037, N20036, N19838);
or OR3 (N20038, N20023, N3135, N6653);
and AND4 (N20039, N20038, N17836, N5298, N16711);
not NOT1 (N20040, N20004);
nand NAND2 (N20041, N20028, N8420);
nor NOR4 (N20042, N20040, N8413, N10739, N10150);
nor NOR2 (N20043, N20037, N18554);
xor XOR2 (N20044, N20032, N6814);
buf BUF1 (N20045, N20011);
nor NOR3 (N20046, N20031, N13668, N7061);
not NOT1 (N20047, N20035);
buf BUF1 (N20048, N20044);
nor NOR4 (N20049, N20046, N13442, N6184, N5042);
and AND4 (N20050, N20043, N9727, N11300, N6473);
xor XOR2 (N20051, N20048, N8732);
nor NOR4 (N20052, N20051, N18108, N8215, N11734);
xor XOR2 (N20053, N20047, N15130);
not NOT1 (N20054, N20041);
nand NAND3 (N20055, N20045, N1063, N11105);
nand NAND4 (N20056, N20030, N1933, N12925, N18975);
xor XOR2 (N20057, N20053, N15922);
and AND2 (N20058, N20054, N3086);
buf BUF1 (N20059, N20049);
or OR3 (N20060, N20042, N3576, N19996);
xor XOR2 (N20061, N20056, N19388);
buf BUF1 (N20062, N20050);
nor NOR3 (N20063, N20058, N1295, N15883);
xor XOR2 (N20064, N20057, N16224);
not NOT1 (N20065, N20055);
nor NOR2 (N20066, N20064, N9923);
not NOT1 (N20067, N20039);
nand NAND4 (N20068, N20059, N19776, N2060, N1977);
or OR4 (N20069, N20062, N18293, N15327, N6709);
xor XOR2 (N20070, N20060, N5225);
buf BUF1 (N20071, N20067);
buf BUF1 (N20072, N20063);
xor XOR2 (N20073, N20070, N8814);
not NOT1 (N20074, N20069);
nand NAND4 (N20075, N20071, N14160, N9832, N16547);
buf BUF1 (N20076, N20075);
and AND3 (N20077, N20066, N5981, N2577);
and AND4 (N20078, N20074, N9189, N5552, N3563);
or OR4 (N20079, N20078, N18585, N3263, N1744);
not NOT1 (N20080, N20061);
not NOT1 (N20081, N20068);
nor NOR2 (N20082, N20072, N6049);
or OR3 (N20083, N20077, N16548, N10585);
or OR4 (N20084, N20081, N3929, N16009, N4814);
or OR3 (N20085, N20083, N10363, N9134);
and AND2 (N20086, N20065, N2297);
nor NOR3 (N20087, N20034, N9458, N18436);
xor XOR2 (N20088, N20076, N3361);
buf BUF1 (N20089, N20087);
buf BUF1 (N20090, N20079);
xor XOR2 (N20091, N20082, N18905);
nor NOR3 (N20092, N20052, N848, N19232);
xor XOR2 (N20093, N20090, N15835);
buf BUF1 (N20094, N20073);
or OR2 (N20095, N20089, N18074);
and AND3 (N20096, N20094, N7872, N567);
or OR2 (N20097, N20088, N1716);
and AND2 (N20098, N20080, N18727);
not NOT1 (N20099, N20098);
and AND3 (N20100, N20099, N3660, N6088);
nor NOR2 (N20101, N20093, N436);
nand NAND2 (N20102, N20101, N18860);
and AND2 (N20103, N20100, N12468);
nor NOR3 (N20104, N20091, N5733, N5222);
and AND4 (N20105, N20097, N9826, N9403, N15548);
or OR2 (N20106, N20102, N10511);
nor NOR3 (N20107, N20104, N2885, N6017);
nor NOR3 (N20108, N20086, N14166, N17428);
and AND2 (N20109, N20084, N19543);
and AND2 (N20110, N20092, N1659);
not NOT1 (N20111, N20103);
buf BUF1 (N20112, N20107);
nor NOR2 (N20113, N20105, N17410);
not NOT1 (N20114, N20113);
or OR2 (N20115, N20109, N19103);
nor NOR2 (N20116, N20106, N10498);
and AND4 (N20117, N20115, N225, N17321, N547);
or OR3 (N20118, N20114, N8127, N16524);
xor XOR2 (N20119, N20095, N13642);
and AND4 (N20120, N20118, N9038, N10573, N14631);
xor XOR2 (N20121, N20117, N16166);
and AND4 (N20122, N20110, N17909, N2893, N1318);
buf BUF1 (N20123, N20108);
nor NOR4 (N20124, N20119, N319, N19822, N10492);
and AND2 (N20125, N20116, N7565);
or OR2 (N20126, N20112, N4402);
xor XOR2 (N20127, N20096, N11397);
and AND2 (N20128, N20127, N16534);
xor XOR2 (N20129, N20122, N15676);
nand NAND2 (N20130, N20126, N309);
not NOT1 (N20131, N20129);
nor NOR4 (N20132, N20125, N6459, N11448, N1392);
nand NAND3 (N20133, N20120, N9987, N10884);
nor NOR2 (N20134, N20111, N8997);
xor XOR2 (N20135, N20131, N2101);
and AND3 (N20136, N20124, N11271, N1221);
or OR4 (N20137, N20130, N8363, N14327, N657);
not NOT1 (N20138, N20137);
nand NAND4 (N20139, N20135, N1692, N14370, N4591);
and AND4 (N20140, N20132, N2803, N1170, N9088);
nand NAND2 (N20141, N20085, N5274);
xor XOR2 (N20142, N20140, N5961);
not NOT1 (N20143, N20139);
and AND4 (N20144, N20141, N4005, N5142, N13846);
nor NOR4 (N20145, N20136, N5177, N8905, N3433);
xor XOR2 (N20146, N20145, N7125);
and AND4 (N20147, N20146, N10275, N12032, N7577);
and AND2 (N20148, N20142, N7931);
buf BUF1 (N20149, N20144);
buf BUF1 (N20150, N20147);
buf BUF1 (N20151, N20134);
or OR4 (N20152, N20138, N11039, N17292, N3506);
xor XOR2 (N20153, N20123, N18603);
nand NAND4 (N20154, N20148, N11610, N6052, N6164);
or OR2 (N20155, N20121, N18405);
not NOT1 (N20156, N20151);
or OR2 (N20157, N20143, N16421);
nand NAND4 (N20158, N20128, N10925, N8565, N15215);
xor XOR2 (N20159, N20152, N13261);
not NOT1 (N20160, N20157);
buf BUF1 (N20161, N20160);
and AND2 (N20162, N20149, N11246);
not NOT1 (N20163, N20156);
or OR2 (N20164, N20162, N5643);
buf BUF1 (N20165, N20155);
nor NOR4 (N20166, N20161, N13967, N4562, N18815);
nor NOR2 (N20167, N20153, N1489);
buf BUF1 (N20168, N20165);
and AND2 (N20169, N20164, N8908);
nand NAND3 (N20170, N20167, N16629, N19396);
not NOT1 (N20171, N20150);
xor XOR2 (N20172, N20171, N161);
xor XOR2 (N20173, N20172, N9866);
xor XOR2 (N20174, N20169, N5429);
or OR3 (N20175, N20158, N17874, N9113);
or OR3 (N20176, N20174, N2803, N6359);
xor XOR2 (N20177, N20175, N16539);
xor XOR2 (N20178, N20133, N18437);
and AND2 (N20179, N20178, N16478);
xor XOR2 (N20180, N20177, N19291);
or OR3 (N20181, N20176, N1130, N18017);
or OR4 (N20182, N20173, N5808, N17244, N725);
buf BUF1 (N20183, N20154);
or OR3 (N20184, N20182, N19730, N11643);
nor NOR2 (N20185, N20181, N344);
and AND3 (N20186, N20183, N14741, N19447);
buf BUF1 (N20187, N20186);
buf BUF1 (N20188, N20179);
xor XOR2 (N20189, N20170, N15809);
not NOT1 (N20190, N20166);
or OR4 (N20191, N20163, N363, N16542, N1627);
nor NOR3 (N20192, N20187, N17055, N16125);
buf BUF1 (N20193, N20180);
not NOT1 (N20194, N20168);
and AND3 (N20195, N20184, N12113, N17412);
nand NAND3 (N20196, N20189, N5939, N19261);
nand NAND2 (N20197, N20190, N6170);
buf BUF1 (N20198, N20193);
not NOT1 (N20199, N20185);
nor NOR4 (N20200, N20197, N8939, N18110, N1341);
nand NAND2 (N20201, N20196, N3320);
nor NOR4 (N20202, N20191, N16299, N4250, N10265);
or OR2 (N20203, N20200, N8769);
nor NOR2 (N20204, N20202, N1212);
nor NOR2 (N20205, N20192, N5395);
not NOT1 (N20206, N20159);
nor NOR4 (N20207, N20195, N14820, N8423, N7981);
and AND4 (N20208, N20207, N10981, N16084, N19836);
buf BUF1 (N20209, N20188);
or OR4 (N20210, N20201, N19297, N15646, N7667);
buf BUF1 (N20211, N20208);
buf BUF1 (N20212, N20199);
buf BUF1 (N20213, N20211);
or OR4 (N20214, N20204, N17701, N8877, N11523);
not NOT1 (N20215, N20209);
nor NOR2 (N20216, N20213, N19666);
buf BUF1 (N20217, N20215);
xor XOR2 (N20218, N20203, N7752);
not NOT1 (N20219, N20194);
xor XOR2 (N20220, N20210, N16060);
nor NOR4 (N20221, N20206, N4885, N3675, N3263);
nor NOR2 (N20222, N20221, N7862);
nand NAND3 (N20223, N20220, N8744, N5235);
not NOT1 (N20224, N20214);
nand NAND3 (N20225, N20216, N2555, N13971);
nand NAND2 (N20226, N20217, N9535);
nor NOR2 (N20227, N20223, N16677);
buf BUF1 (N20228, N20219);
nand NAND4 (N20229, N20225, N18314, N3426, N7150);
nand NAND3 (N20230, N20226, N19441, N19358);
buf BUF1 (N20231, N20198);
and AND4 (N20232, N20231, N19349, N6632, N1543);
nand NAND3 (N20233, N20230, N7844, N846);
xor XOR2 (N20234, N20205, N19044);
nor NOR4 (N20235, N20228, N13575, N16327, N12765);
or OR2 (N20236, N20224, N1326);
nor NOR3 (N20237, N20229, N4215, N13501);
nand NAND2 (N20238, N20232, N6487);
nand NAND3 (N20239, N20222, N10714, N4372);
xor XOR2 (N20240, N20227, N1432);
not NOT1 (N20241, N20237);
xor XOR2 (N20242, N20235, N2092);
xor XOR2 (N20243, N20241, N11377);
buf BUF1 (N20244, N20212);
nand NAND2 (N20245, N20239, N7326);
or OR2 (N20246, N20218, N3022);
not NOT1 (N20247, N20236);
buf BUF1 (N20248, N20243);
or OR4 (N20249, N20248, N19726, N8437, N19841);
or OR4 (N20250, N20249, N9344, N2609, N249);
or OR4 (N20251, N20233, N3840, N10681, N18661);
xor XOR2 (N20252, N20245, N18687);
nor NOR4 (N20253, N20242, N11304, N8584, N13822);
nor NOR3 (N20254, N20251, N3963, N14546);
nand NAND4 (N20255, N20253, N12259, N18480, N6090);
xor XOR2 (N20256, N20250, N17366);
xor XOR2 (N20257, N20234, N3991);
not NOT1 (N20258, N20247);
buf BUF1 (N20259, N20252);
or OR4 (N20260, N20246, N2655, N2461, N15679);
not NOT1 (N20261, N20257);
xor XOR2 (N20262, N20238, N10596);
and AND2 (N20263, N20256, N14658);
xor XOR2 (N20264, N20240, N8683);
or OR2 (N20265, N20255, N16628);
nand NAND3 (N20266, N20263, N13329, N17842);
buf BUF1 (N20267, N20244);
xor XOR2 (N20268, N20258, N11425);
nor NOR4 (N20269, N20264, N16367, N17980, N3551);
or OR3 (N20270, N20260, N13534, N6417);
and AND2 (N20271, N20254, N18275);
xor XOR2 (N20272, N20266, N12333);
and AND3 (N20273, N20268, N20203, N8322);
xor XOR2 (N20274, N20262, N18266);
or OR4 (N20275, N20269, N312, N13972, N1092);
or OR3 (N20276, N20271, N4825, N9495);
nor NOR4 (N20277, N20272, N12933, N18451, N3143);
and AND3 (N20278, N20276, N11209, N9682);
xor XOR2 (N20279, N20273, N13129);
not NOT1 (N20280, N20259);
nor NOR2 (N20281, N20280, N11522);
nor NOR3 (N20282, N20281, N16616, N7052);
nor NOR2 (N20283, N20275, N3674);
or OR2 (N20284, N20274, N7803);
buf BUF1 (N20285, N20277);
or OR2 (N20286, N20261, N14923);
not NOT1 (N20287, N20270);
buf BUF1 (N20288, N20267);
nand NAND3 (N20289, N20265, N4194, N1963);
or OR3 (N20290, N20278, N4869, N4658);
and AND3 (N20291, N20288, N11379, N4630);
nand NAND3 (N20292, N20283, N4831, N15957);
nand NAND3 (N20293, N20284, N7915, N9996);
nor NOR3 (N20294, N20293, N11769, N13097);
not NOT1 (N20295, N20282);
nor NOR4 (N20296, N20286, N1412, N644, N19913);
and AND3 (N20297, N20292, N5639, N6751);
and AND2 (N20298, N20295, N16482);
or OR4 (N20299, N20279, N3000, N17446, N9592);
buf BUF1 (N20300, N20287);
not NOT1 (N20301, N20296);
or OR3 (N20302, N20299, N2870, N3709);
nor NOR4 (N20303, N20294, N10981, N1686, N7893);
buf BUF1 (N20304, N20285);
xor XOR2 (N20305, N20303, N11801);
buf BUF1 (N20306, N20290);
xor XOR2 (N20307, N20302, N10747);
xor XOR2 (N20308, N20306, N4661);
nor NOR2 (N20309, N20307, N6122);
or OR4 (N20310, N20300, N5439, N5858, N10761);
or OR2 (N20311, N20309, N13498);
nand NAND2 (N20312, N20311, N5085);
not NOT1 (N20313, N20289);
buf BUF1 (N20314, N20312);
not NOT1 (N20315, N20298);
buf BUF1 (N20316, N20310);
nor NOR3 (N20317, N20301, N12994, N9476);
or OR2 (N20318, N20314, N10117);
or OR2 (N20319, N20291, N10920);
or OR3 (N20320, N20317, N109, N902);
nor NOR4 (N20321, N20305, N278, N10375, N9138);
and AND3 (N20322, N20320, N7948, N12383);
or OR3 (N20323, N20308, N12586, N9359);
or OR3 (N20324, N20321, N2064, N4079);
and AND3 (N20325, N20318, N17149, N14056);
nor NOR2 (N20326, N20297, N5743);
xor XOR2 (N20327, N20313, N9200);
xor XOR2 (N20328, N20322, N4571);
not NOT1 (N20329, N20323);
nand NAND2 (N20330, N20316, N16950);
not NOT1 (N20331, N20328);
or OR4 (N20332, N20326, N7200, N11548, N15899);
or OR3 (N20333, N20325, N1273, N6789);
xor XOR2 (N20334, N20330, N18907);
buf BUF1 (N20335, N20324);
not NOT1 (N20336, N20335);
nand NAND3 (N20337, N20336, N13504, N19262);
nand NAND3 (N20338, N20319, N19118, N10728);
and AND4 (N20339, N20329, N466, N15766, N16452);
not NOT1 (N20340, N20327);
buf BUF1 (N20341, N20304);
xor XOR2 (N20342, N20332, N5112);
not NOT1 (N20343, N20334);
not NOT1 (N20344, N20342);
xor XOR2 (N20345, N20333, N2727);
buf BUF1 (N20346, N20338);
xor XOR2 (N20347, N20345, N16807);
nor NOR2 (N20348, N20341, N4563);
not NOT1 (N20349, N20339);
not NOT1 (N20350, N20315);
nor NOR2 (N20351, N20350, N136);
or OR4 (N20352, N20346, N7140, N18855, N3403);
and AND2 (N20353, N20352, N17562);
and AND4 (N20354, N20349, N10534, N5718, N4001);
nand NAND4 (N20355, N20347, N17698, N14288, N16724);
nand NAND4 (N20356, N20344, N1744, N13601, N16533);
nor NOR2 (N20357, N20356, N3655);
nand NAND2 (N20358, N20357, N7576);
nor NOR4 (N20359, N20340, N9507, N17493, N11261);
not NOT1 (N20360, N20351);
xor XOR2 (N20361, N20331, N2963);
or OR4 (N20362, N20354, N9469, N11238, N15461);
xor XOR2 (N20363, N20353, N16588);
or OR2 (N20364, N20343, N9735);
nor NOR4 (N20365, N20348, N10488, N15187, N7184);
nor NOR4 (N20366, N20359, N6253, N6800, N12724);
not NOT1 (N20367, N20364);
or OR2 (N20368, N20337, N7514);
and AND2 (N20369, N20365, N15319);
nand NAND4 (N20370, N20367, N3649, N17893, N10498);
xor XOR2 (N20371, N20361, N1217);
nand NAND2 (N20372, N20360, N11959);
nand NAND3 (N20373, N20369, N16711, N19258);
or OR2 (N20374, N20366, N1749);
or OR4 (N20375, N20371, N13641, N15239, N13313);
xor XOR2 (N20376, N20368, N15039);
and AND2 (N20377, N20362, N15903);
not NOT1 (N20378, N20372);
not NOT1 (N20379, N20374);
nor NOR4 (N20380, N20358, N14860, N451, N14581);
nand NAND4 (N20381, N20375, N17191, N2652, N44);
and AND4 (N20382, N20355, N18545, N16484, N2941);
or OR4 (N20383, N20381, N18504, N16513, N4662);
or OR3 (N20384, N20378, N14265, N14071);
not NOT1 (N20385, N20370);
nor NOR4 (N20386, N20363, N7206, N5130, N17126);
or OR2 (N20387, N20384, N15903);
and AND3 (N20388, N20382, N3968, N7903);
not NOT1 (N20389, N20377);
nor NOR4 (N20390, N20376, N14842, N3900, N9555);
and AND4 (N20391, N20383, N11457, N14675, N6652);
nor NOR3 (N20392, N20389, N14541, N12967);
nor NOR4 (N20393, N20385, N12824, N11676, N7824);
nand NAND3 (N20394, N20388, N19530, N20185);
buf BUF1 (N20395, N20380);
nor NOR3 (N20396, N20391, N7983, N14061);
buf BUF1 (N20397, N20387);
and AND3 (N20398, N20396, N17670, N8594);
not NOT1 (N20399, N20397);
or OR4 (N20400, N20393, N11766, N14778, N18970);
buf BUF1 (N20401, N20390);
and AND4 (N20402, N20395, N871, N15918, N12616);
nor NOR3 (N20403, N20373, N19929, N13757);
or OR4 (N20404, N20401, N14350, N154, N565);
buf BUF1 (N20405, N20402);
nor NOR4 (N20406, N20392, N13400, N17682, N16751);
or OR3 (N20407, N20379, N1869, N6847);
buf BUF1 (N20408, N20386);
or OR2 (N20409, N20400, N17467);
not NOT1 (N20410, N20398);
or OR3 (N20411, N20403, N5684, N5620);
or OR3 (N20412, N20404, N12897, N10461);
buf BUF1 (N20413, N20411);
nor NOR4 (N20414, N20406, N15984, N18132, N7214);
nand NAND4 (N20415, N20413, N16544, N5477, N12441);
and AND4 (N20416, N20409, N18780, N14669, N14645);
and AND2 (N20417, N20410, N8171);
not NOT1 (N20418, N20407);
not NOT1 (N20419, N20399);
nor NOR3 (N20420, N20394, N16476, N5737);
not NOT1 (N20421, N20420);
xor XOR2 (N20422, N20414, N4443);
not NOT1 (N20423, N20418);
xor XOR2 (N20424, N20412, N7210);
xor XOR2 (N20425, N20416, N6751);
and AND2 (N20426, N20421, N15988);
xor XOR2 (N20427, N20426, N1891);
buf BUF1 (N20428, N20423);
not NOT1 (N20429, N20422);
nand NAND4 (N20430, N20429, N8028, N8680, N5900);
and AND2 (N20431, N20427, N12783);
and AND2 (N20432, N20431, N18107);
nor NOR3 (N20433, N20432, N6203, N8556);
not NOT1 (N20434, N20415);
or OR2 (N20435, N20433, N677);
buf BUF1 (N20436, N20419);
xor XOR2 (N20437, N20428, N3763);
not NOT1 (N20438, N20424);
buf BUF1 (N20439, N20436);
xor XOR2 (N20440, N20425, N1624);
xor XOR2 (N20441, N20417, N8168);
or OR2 (N20442, N20408, N6192);
not NOT1 (N20443, N20439);
nand NAND4 (N20444, N20441, N18830, N17660, N14912);
and AND4 (N20445, N20405, N14305, N8984, N19076);
buf BUF1 (N20446, N20435);
nor NOR3 (N20447, N20442, N11979, N7327);
buf BUF1 (N20448, N20447);
nor NOR2 (N20449, N20434, N7718);
xor XOR2 (N20450, N20449, N19461);
not NOT1 (N20451, N20440);
buf BUF1 (N20452, N20448);
buf BUF1 (N20453, N20445);
xor XOR2 (N20454, N20450, N10771);
nand NAND2 (N20455, N20437, N13154);
and AND3 (N20456, N20454, N14686, N12271);
or OR4 (N20457, N20446, N3629, N19446, N8995);
buf BUF1 (N20458, N20430);
nand NAND3 (N20459, N20451, N19051, N2211);
nand NAND3 (N20460, N20453, N6545, N4955);
not NOT1 (N20461, N20459);
and AND4 (N20462, N20456, N19149, N11741, N14693);
and AND4 (N20463, N20444, N10492, N3840, N14281);
nand NAND4 (N20464, N20457, N1947, N12231, N12060);
nor NOR3 (N20465, N20463, N1852, N14296);
and AND2 (N20466, N20438, N4452);
nand NAND2 (N20467, N20460, N16055);
buf BUF1 (N20468, N20461);
and AND3 (N20469, N20467, N997, N17101);
or OR3 (N20470, N20458, N15848, N1216);
not NOT1 (N20471, N20464);
not NOT1 (N20472, N20452);
or OR3 (N20473, N20466, N877, N19390);
buf BUF1 (N20474, N20468);
not NOT1 (N20475, N20465);
not NOT1 (N20476, N20469);
buf BUF1 (N20477, N20471);
nor NOR2 (N20478, N20477, N7231);
and AND4 (N20479, N20478, N8424, N11958, N18540);
not NOT1 (N20480, N20473);
nor NOR4 (N20481, N20472, N9329, N18061, N19962);
and AND4 (N20482, N20480, N11250, N20315, N1633);
buf BUF1 (N20483, N20455);
xor XOR2 (N20484, N20475, N19094);
or OR2 (N20485, N20484, N9212);
buf BUF1 (N20486, N20483);
xor XOR2 (N20487, N20482, N6391);
not NOT1 (N20488, N20443);
and AND3 (N20489, N20487, N4273, N5715);
nand NAND3 (N20490, N20479, N13365, N4138);
or OR2 (N20491, N20488, N2855);
xor XOR2 (N20492, N20474, N10828);
buf BUF1 (N20493, N20476);
and AND4 (N20494, N20470, N3688, N15188, N4619);
nand NAND2 (N20495, N20494, N7366);
nor NOR3 (N20496, N20486, N11864, N17301);
nand NAND3 (N20497, N20496, N2240, N13266);
nand NAND3 (N20498, N20491, N10976, N8463);
xor XOR2 (N20499, N20497, N11326);
or OR3 (N20500, N20493, N1970, N17439);
nor NOR2 (N20501, N20490, N17532);
xor XOR2 (N20502, N20500, N18704);
not NOT1 (N20503, N20501);
or OR2 (N20504, N20499, N14063);
not NOT1 (N20505, N20481);
nand NAND2 (N20506, N20498, N10201);
xor XOR2 (N20507, N20492, N1753);
not NOT1 (N20508, N20495);
and AND4 (N20509, N20506, N14709, N16820, N18482);
and AND4 (N20510, N20462, N8733, N19252, N8908);
or OR2 (N20511, N20505, N12225);
xor XOR2 (N20512, N20510, N434);
buf BUF1 (N20513, N20503);
and AND3 (N20514, N20512, N11235, N6555);
xor XOR2 (N20515, N20489, N12970);
not NOT1 (N20516, N20514);
or OR4 (N20517, N20509, N9472, N270, N11507);
nor NOR3 (N20518, N20485, N76, N14687);
nand NAND4 (N20519, N20511, N7387, N18138, N8340);
not NOT1 (N20520, N20519);
xor XOR2 (N20521, N20513, N4899);
and AND3 (N20522, N20520, N7657, N5872);
nand NAND2 (N20523, N20507, N4874);
not NOT1 (N20524, N20517);
and AND3 (N20525, N20502, N4807, N14041);
not NOT1 (N20526, N20521);
nand NAND3 (N20527, N20516, N10793, N2385);
or OR2 (N20528, N20518, N10420);
and AND2 (N20529, N20526, N17451);
not NOT1 (N20530, N20504);
nand NAND3 (N20531, N20525, N17810, N5540);
xor XOR2 (N20532, N20523, N124);
and AND2 (N20533, N20531, N4398);
nand NAND2 (N20534, N20530, N16349);
not NOT1 (N20535, N20515);
nor NOR2 (N20536, N20533, N13255);
and AND4 (N20537, N20527, N15049, N14955, N17966);
nor NOR4 (N20538, N20528, N3102, N18018, N2391);
nand NAND3 (N20539, N20529, N14615, N1362);
not NOT1 (N20540, N20535);
nor NOR3 (N20541, N20537, N9312, N7051);
xor XOR2 (N20542, N20538, N6507);
xor XOR2 (N20543, N20542, N4727);
or OR2 (N20544, N20534, N13260);
nor NOR4 (N20545, N20544, N8574, N13336, N8572);
or OR3 (N20546, N20532, N4250, N6381);
nor NOR2 (N20547, N20524, N14920);
and AND3 (N20548, N20547, N1486, N5055);
not NOT1 (N20549, N20536);
not NOT1 (N20550, N20545);
not NOT1 (N20551, N20543);
and AND4 (N20552, N20540, N13372, N15786, N2804);
buf BUF1 (N20553, N20551);
xor XOR2 (N20554, N20539, N11069);
xor XOR2 (N20555, N20508, N16254);
or OR4 (N20556, N20555, N13364, N7732, N7145);
or OR2 (N20557, N20556, N221);
nand NAND2 (N20558, N20554, N4251);
nor NOR3 (N20559, N20553, N19514, N19039);
nand NAND2 (N20560, N20552, N5094);
nand NAND4 (N20561, N20522, N20136, N14920, N5519);
and AND2 (N20562, N20560, N17842);
nand NAND4 (N20563, N20561, N6149, N18765, N1860);
nand NAND2 (N20564, N20558, N20204);
nor NOR2 (N20565, N20541, N10642);
xor XOR2 (N20566, N20564, N11259);
nand NAND3 (N20567, N20559, N14083, N14510);
nand NAND2 (N20568, N20565, N16739);
nand NAND2 (N20569, N20563, N8708);
and AND3 (N20570, N20546, N19310, N19084);
or OR2 (N20571, N20550, N4011);
and AND2 (N20572, N20548, N18986);
nand NAND2 (N20573, N20568, N6710);
not NOT1 (N20574, N20569);
buf BUF1 (N20575, N20574);
nor NOR3 (N20576, N20575, N6796, N11037);
buf BUF1 (N20577, N20566);
xor XOR2 (N20578, N20577, N18553);
nand NAND2 (N20579, N20571, N11073);
buf BUF1 (N20580, N20573);
nor NOR2 (N20581, N20567, N471);
and AND3 (N20582, N20576, N12912, N7320);
nor NOR4 (N20583, N20582, N9294, N16832, N18151);
xor XOR2 (N20584, N20570, N11222);
xor XOR2 (N20585, N20572, N3524);
nor NOR4 (N20586, N20580, N396, N4495, N17639);
and AND2 (N20587, N20585, N11873);
or OR4 (N20588, N20579, N7334, N3050, N1219);
xor XOR2 (N20589, N20562, N6387);
and AND2 (N20590, N20589, N4457);
and AND2 (N20591, N20590, N2537);
buf BUF1 (N20592, N20584);
or OR2 (N20593, N20578, N146);
xor XOR2 (N20594, N20588, N17477);
xor XOR2 (N20595, N20557, N6621);
nand NAND2 (N20596, N20583, N1189);
not NOT1 (N20597, N20549);
xor XOR2 (N20598, N20592, N8364);
nor NOR4 (N20599, N20591, N312, N9039, N16251);
and AND4 (N20600, N20593, N9231, N17141, N19082);
and AND3 (N20601, N20596, N1213, N16765);
nand NAND4 (N20602, N20581, N6698, N11519, N1258);
and AND3 (N20603, N20587, N6320, N2500);
nor NOR3 (N20604, N20602, N8468, N19660);
not NOT1 (N20605, N20599);
and AND4 (N20606, N20598, N51, N2383, N1564);
not NOT1 (N20607, N20586);
or OR2 (N20608, N20594, N572);
not NOT1 (N20609, N20607);
and AND3 (N20610, N20604, N16944, N2575);
nor NOR4 (N20611, N20595, N14484, N17440, N8070);
xor XOR2 (N20612, N20600, N4648);
nor NOR2 (N20613, N20605, N3737);
or OR2 (N20614, N20613, N7605);
and AND3 (N20615, N20608, N4268, N1395);
not NOT1 (N20616, N20614);
and AND4 (N20617, N20609, N4242, N13147, N19905);
not NOT1 (N20618, N20597);
buf BUF1 (N20619, N20601);
not NOT1 (N20620, N20603);
xor XOR2 (N20621, N20610, N2068);
and AND4 (N20622, N20611, N13803, N12255, N10694);
and AND2 (N20623, N20620, N10015);
nor NOR4 (N20624, N20622, N16768, N658, N723);
buf BUF1 (N20625, N20617);
nand NAND4 (N20626, N20606, N5824, N11357, N13563);
nor NOR2 (N20627, N20625, N12509);
xor XOR2 (N20628, N20627, N10825);
not NOT1 (N20629, N20624);
and AND3 (N20630, N20628, N20569, N3872);
buf BUF1 (N20631, N20621);
not NOT1 (N20632, N20630);
or OR4 (N20633, N20631, N19367, N2617, N1676);
and AND2 (N20634, N20612, N16342);
not NOT1 (N20635, N20623);
buf BUF1 (N20636, N20629);
xor XOR2 (N20637, N20615, N13583);
nand NAND2 (N20638, N20637, N15890);
nand NAND3 (N20639, N20626, N15832, N12831);
buf BUF1 (N20640, N20633);
nand NAND2 (N20641, N20636, N2676);
xor XOR2 (N20642, N20639, N7245);
or OR2 (N20643, N20619, N15215);
nor NOR2 (N20644, N20632, N239);
and AND3 (N20645, N20643, N18000, N3237);
or OR3 (N20646, N20616, N10046, N14178);
not NOT1 (N20647, N20646);
nor NOR2 (N20648, N20638, N5975);
and AND3 (N20649, N20634, N17875, N10263);
nor NOR2 (N20650, N20649, N4618);
or OR3 (N20651, N20650, N1526, N6926);
nand NAND3 (N20652, N20642, N5558, N19192);
not NOT1 (N20653, N20652);
or OR4 (N20654, N20645, N20397, N7526, N3395);
not NOT1 (N20655, N20640);
nand NAND4 (N20656, N20655, N13749, N2105, N17499);
and AND2 (N20657, N20656, N9662);
or OR3 (N20658, N20618, N15198, N12663);
buf BUF1 (N20659, N20635);
nand NAND4 (N20660, N20648, N3663, N16592, N17727);
buf BUF1 (N20661, N20647);
nor NOR4 (N20662, N20641, N11092, N8533, N16562);
not NOT1 (N20663, N20657);
nand NAND2 (N20664, N20651, N6841);
buf BUF1 (N20665, N20658);
or OR2 (N20666, N20661, N11578);
not NOT1 (N20667, N20663);
buf BUF1 (N20668, N20644);
nand NAND2 (N20669, N20654, N2330);
and AND4 (N20670, N20659, N15059, N7085, N14130);
buf BUF1 (N20671, N20669);
and AND3 (N20672, N20662, N1865, N7653);
buf BUF1 (N20673, N20653);
and AND4 (N20674, N20672, N18649, N10201, N12700);
and AND2 (N20675, N20668, N9464);
buf BUF1 (N20676, N20671);
and AND3 (N20677, N20675, N7922, N3959);
or OR3 (N20678, N20677, N2421, N13849);
nand NAND4 (N20679, N20676, N1109, N18084, N19987);
buf BUF1 (N20680, N20679);
nor NOR2 (N20681, N20667, N8861);
and AND2 (N20682, N20665, N1646);
not NOT1 (N20683, N20680);
xor XOR2 (N20684, N20682, N15218);
and AND3 (N20685, N20670, N13344, N3815);
xor XOR2 (N20686, N20660, N8322);
not NOT1 (N20687, N20678);
nand NAND2 (N20688, N20683, N12871);
buf BUF1 (N20689, N20686);
nand NAND4 (N20690, N20687, N14967, N17807, N8609);
not NOT1 (N20691, N20688);
not NOT1 (N20692, N20685);
and AND3 (N20693, N20673, N20342, N320);
buf BUF1 (N20694, N20692);
not NOT1 (N20695, N20681);
and AND3 (N20696, N20690, N3399, N6511);
not NOT1 (N20697, N20666);
not NOT1 (N20698, N20695);
not NOT1 (N20699, N20664);
not NOT1 (N20700, N20689);
nand NAND4 (N20701, N20674, N16678, N6331, N17428);
nor NOR3 (N20702, N20697, N4790, N18703);
or OR4 (N20703, N20694, N334, N694, N6052);
or OR2 (N20704, N20696, N17297);
nand NAND4 (N20705, N20693, N12051, N16019, N20444);
and AND2 (N20706, N20704, N8593);
xor XOR2 (N20707, N20691, N614);
not NOT1 (N20708, N20706);
or OR3 (N20709, N20698, N15373, N11000);
or OR2 (N20710, N20705, N13422);
nand NAND2 (N20711, N20710, N7463);
not NOT1 (N20712, N20702);
xor XOR2 (N20713, N20701, N1557);
nand NAND4 (N20714, N20707, N11726, N7399, N1637);
not NOT1 (N20715, N20700);
or OR4 (N20716, N20712, N14580, N16931, N12668);
not NOT1 (N20717, N20709);
xor XOR2 (N20718, N20699, N3578);
xor XOR2 (N20719, N20711, N12512);
or OR2 (N20720, N20703, N3812);
buf BUF1 (N20721, N20717);
or OR3 (N20722, N20715, N9320, N13734);
nor NOR2 (N20723, N20720, N8526);
xor XOR2 (N20724, N20722, N7916);
nand NAND4 (N20725, N20713, N19147, N19884, N16754);
xor XOR2 (N20726, N20714, N1204);
and AND3 (N20727, N20723, N9373, N4011);
not NOT1 (N20728, N20708);
nor NOR4 (N20729, N20718, N10930, N9362, N4150);
and AND4 (N20730, N20725, N19936, N12150, N6425);
or OR4 (N20731, N20684, N14084, N3536, N8334);
not NOT1 (N20732, N20727);
nor NOR3 (N20733, N20728, N7012, N15729);
and AND4 (N20734, N20731, N15761, N6990, N11175);
nand NAND3 (N20735, N20719, N18052, N12843);
not NOT1 (N20736, N20735);
not NOT1 (N20737, N20726);
and AND4 (N20738, N20737, N13909, N7981, N18484);
xor XOR2 (N20739, N20738, N10366);
xor XOR2 (N20740, N20733, N3040);
nor NOR4 (N20741, N20721, N10195, N4993, N7419);
nor NOR4 (N20742, N20736, N12310, N4716, N10978);
not NOT1 (N20743, N20716);
nor NOR3 (N20744, N20739, N4126, N4971);
xor XOR2 (N20745, N20724, N4414);
xor XOR2 (N20746, N20742, N15226);
xor XOR2 (N20747, N20734, N7336);
buf BUF1 (N20748, N20741);
buf BUF1 (N20749, N20744);
and AND2 (N20750, N20745, N5875);
and AND4 (N20751, N20729, N918, N13541, N14743);
not NOT1 (N20752, N20749);
buf BUF1 (N20753, N20748);
and AND3 (N20754, N20752, N9168, N12130);
and AND4 (N20755, N20750, N1536, N4970, N8802);
not NOT1 (N20756, N20754);
and AND2 (N20757, N20730, N3781);
nand NAND3 (N20758, N20746, N414, N6013);
not NOT1 (N20759, N20740);
xor XOR2 (N20760, N20747, N2355);
and AND3 (N20761, N20759, N5647, N1213);
nand NAND3 (N20762, N20753, N9556, N15563);
xor XOR2 (N20763, N20761, N19606);
nand NAND3 (N20764, N20751, N1982, N973);
or OR4 (N20765, N20743, N5344, N13683, N5849);
buf BUF1 (N20766, N20762);
and AND4 (N20767, N20756, N17348, N17373, N2472);
nor NOR2 (N20768, N20758, N13691);
and AND4 (N20769, N20767, N13349, N20408, N8645);
xor XOR2 (N20770, N20732, N18897);
not NOT1 (N20771, N20766);
nor NOR2 (N20772, N20760, N3402);
nand NAND2 (N20773, N20772, N13747);
buf BUF1 (N20774, N20764);
and AND2 (N20775, N20769, N13411);
nand NAND2 (N20776, N20755, N11640);
xor XOR2 (N20777, N20768, N12246);
not NOT1 (N20778, N20771);
buf BUF1 (N20779, N20765);
or OR4 (N20780, N20773, N12879, N6427, N2092);
or OR3 (N20781, N20777, N14498, N9569);
xor XOR2 (N20782, N20779, N9545);
or OR4 (N20783, N20782, N15784, N9339, N13598);
and AND3 (N20784, N20763, N16693, N13120);
or OR4 (N20785, N20780, N10339, N14577, N4431);
xor XOR2 (N20786, N20776, N13711);
xor XOR2 (N20787, N20781, N12965);
buf BUF1 (N20788, N20783);
or OR3 (N20789, N20775, N16393, N495);
nand NAND3 (N20790, N20786, N5311, N13000);
buf BUF1 (N20791, N20788);
or OR4 (N20792, N20787, N7491, N18946, N11692);
xor XOR2 (N20793, N20757, N11526);
and AND3 (N20794, N20793, N14622, N16817);
nor NOR2 (N20795, N20790, N4459);
xor XOR2 (N20796, N20795, N7015);
nand NAND2 (N20797, N20794, N6975);
nand NAND3 (N20798, N20792, N7933, N14909);
nand NAND3 (N20799, N20785, N7751, N18619);
nand NAND3 (N20800, N20789, N4782, N20789);
nand NAND2 (N20801, N20774, N16020);
nand NAND2 (N20802, N20796, N12677);
nor NOR4 (N20803, N20800, N20750, N656, N3582);
buf BUF1 (N20804, N20784);
nand NAND4 (N20805, N20797, N19910, N17962, N11187);
buf BUF1 (N20806, N20770);
nand NAND3 (N20807, N20778, N1632, N3079);
nand NAND4 (N20808, N20801, N14995, N15501, N9291);
not NOT1 (N20809, N20798);
xor XOR2 (N20810, N20803, N5681);
or OR4 (N20811, N20799, N5943, N3912, N18218);
nand NAND4 (N20812, N20809, N16046, N16039, N1537);
nor NOR3 (N20813, N20811, N20597, N6931);
buf BUF1 (N20814, N20813);
nor NOR2 (N20815, N20791, N13675);
and AND3 (N20816, N20814, N20275, N17694);
xor XOR2 (N20817, N20802, N14790);
nand NAND3 (N20818, N20817, N17322, N20224);
nand NAND2 (N20819, N20805, N4232);
nor NOR4 (N20820, N20807, N6689, N1045, N4475);
not NOT1 (N20821, N20820);
nand NAND3 (N20822, N20818, N10614, N6024);
nand NAND4 (N20823, N20808, N14948, N16538, N9433);
xor XOR2 (N20824, N20819, N12381);
not NOT1 (N20825, N20822);
nand NAND3 (N20826, N20804, N16878, N7630);
nand NAND4 (N20827, N20825, N17135, N5156, N3048);
xor XOR2 (N20828, N20810, N18541);
nor NOR4 (N20829, N20812, N15626, N14141, N7816);
nand NAND2 (N20830, N20828, N288);
nor NOR4 (N20831, N20821, N12148, N8319, N19890);
not NOT1 (N20832, N20830);
or OR3 (N20833, N20829, N16259, N16322);
not NOT1 (N20834, N20832);
not NOT1 (N20835, N20827);
not NOT1 (N20836, N20815);
and AND3 (N20837, N20834, N4188, N4564);
xor XOR2 (N20838, N20836, N17633);
not NOT1 (N20839, N20838);
buf BUF1 (N20840, N20833);
not NOT1 (N20841, N20835);
nand NAND3 (N20842, N20841, N2344, N12352);
nand NAND4 (N20843, N20806, N8642, N18685, N5849);
not NOT1 (N20844, N20831);
xor XOR2 (N20845, N20816, N16268);
xor XOR2 (N20846, N20840, N20514);
not NOT1 (N20847, N20844);
nand NAND4 (N20848, N20823, N9977, N2013, N17877);
not NOT1 (N20849, N20843);
xor XOR2 (N20850, N20837, N18556);
buf BUF1 (N20851, N20842);
and AND4 (N20852, N20826, N20822, N10770, N14048);
or OR2 (N20853, N20839, N12749);
not NOT1 (N20854, N20847);
not NOT1 (N20855, N20853);
buf BUF1 (N20856, N20846);
nor NOR2 (N20857, N20845, N1618);
buf BUF1 (N20858, N20848);
not NOT1 (N20859, N20850);
xor XOR2 (N20860, N20852, N19938);
buf BUF1 (N20861, N20849);
and AND3 (N20862, N20824, N7912, N2551);
buf BUF1 (N20863, N20854);
xor XOR2 (N20864, N20861, N4534);
or OR2 (N20865, N20863, N7776);
buf BUF1 (N20866, N20856);
or OR2 (N20867, N20851, N10106);
not NOT1 (N20868, N20867);
nand NAND4 (N20869, N20862, N13027, N16337, N16431);
not NOT1 (N20870, N20865);
buf BUF1 (N20871, N20859);
nor NOR4 (N20872, N20871, N10294, N12286, N11305);
or OR3 (N20873, N20870, N9470, N9586);
buf BUF1 (N20874, N20864);
nor NOR3 (N20875, N20860, N16715, N6729);
not NOT1 (N20876, N20869);
nor NOR4 (N20877, N20868, N10318, N15268, N3835);
xor XOR2 (N20878, N20858, N9804);
nor NOR2 (N20879, N20872, N14698);
not NOT1 (N20880, N20875);
and AND3 (N20881, N20866, N12958, N7598);
buf BUF1 (N20882, N20855);
xor XOR2 (N20883, N20873, N2206);
nand NAND3 (N20884, N20880, N16996, N10356);
nor NOR4 (N20885, N20877, N1979, N259, N18069);
and AND4 (N20886, N20878, N14786, N571, N13045);
nor NOR3 (N20887, N20857, N19748, N8508);
nor NOR2 (N20888, N20882, N14979);
or OR3 (N20889, N20874, N11780, N17736);
or OR2 (N20890, N20887, N12585);
or OR4 (N20891, N20881, N3293, N11988, N18429);
and AND3 (N20892, N20884, N17887, N8268);
not NOT1 (N20893, N20889);
nor NOR2 (N20894, N20885, N3237);
and AND3 (N20895, N20879, N4211, N16444);
buf BUF1 (N20896, N20894);
xor XOR2 (N20897, N20890, N6337);
and AND4 (N20898, N20876, N14346, N9729, N9034);
nor NOR3 (N20899, N20895, N3390, N889);
or OR2 (N20900, N20897, N10308);
not NOT1 (N20901, N20899);
nand NAND3 (N20902, N20886, N11135, N19174);
and AND3 (N20903, N20901, N5012, N20012);
not NOT1 (N20904, N20893);
and AND2 (N20905, N20883, N18929);
xor XOR2 (N20906, N20888, N19089);
and AND4 (N20907, N20896, N12053, N4664, N2648);
not NOT1 (N20908, N20891);
xor XOR2 (N20909, N20902, N19558);
not NOT1 (N20910, N20908);
xor XOR2 (N20911, N20892, N19700);
and AND3 (N20912, N20903, N3906, N2690);
and AND3 (N20913, N20905, N17049, N7267);
buf BUF1 (N20914, N20911);
not NOT1 (N20915, N20898);
xor XOR2 (N20916, N20906, N12593);
and AND4 (N20917, N20909, N17014, N16072, N4793);
nand NAND2 (N20918, N20915, N17333);
buf BUF1 (N20919, N20900);
nand NAND3 (N20920, N20918, N1321, N11732);
xor XOR2 (N20921, N20912, N3871);
nor NOR3 (N20922, N20920, N15432, N7627);
or OR4 (N20923, N20914, N18420, N5062, N4426);
buf BUF1 (N20924, N20916);
and AND2 (N20925, N20913, N9941);
or OR2 (N20926, N20925, N3333);
not NOT1 (N20927, N20910);
or OR3 (N20928, N20926, N14022, N2971);
and AND3 (N20929, N20922, N8016, N20068);
or OR3 (N20930, N20904, N15860, N7096);
xor XOR2 (N20931, N20919, N8024);
not NOT1 (N20932, N20927);
or OR4 (N20933, N20929, N12780, N15569, N10769);
xor XOR2 (N20934, N20928, N2384);
and AND4 (N20935, N20931, N13237, N2562, N5185);
or OR3 (N20936, N20935, N16577, N420);
buf BUF1 (N20937, N20936);
nand NAND4 (N20938, N20933, N10110, N18950, N3211);
xor XOR2 (N20939, N20917, N8610);
and AND3 (N20940, N20939, N15188, N5258);
nand NAND3 (N20941, N20907, N3866, N16108);
nor NOR4 (N20942, N20924, N2273, N8756, N17428);
nand NAND3 (N20943, N20932, N10945, N3385);
not NOT1 (N20944, N20930);
nand NAND3 (N20945, N20943, N18605, N10744);
buf BUF1 (N20946, N20940);
nor NOR4 (N20947, N20938, N6718, N10520, N20553);
nor NOR3 (N20948, N20947, N12303, N18104);
xor XOR2 (N20949, N20923, N16260);
nor NOR3 (N20950, N20941, N5987, N3068);
or OR3 (N20951, N20942, N20686, N3725);
xor XOR2 (N20952, N20948, N18113);
buf BUF1 (N20953, N20951);
nor NOR3 (N20954, N20952, N9708, N16044);
xor XOR2 (N20955, N20944, N5668);
xor XOR2 (N20956, N20950, N14092);
not NOT1 (N20957, N20934);
nand NAND4 (N20958, N20954, N13387, N7011, N19390);
not NOT1 (N20959, N20946);
not NOT1 (N20960, N20957);
buf BUF1 (N20961, N20937);
not NOT1 (N20962, N20953);
nand NAND2 (N20963, N20961, N6674);
not NOT1 (N20964, N20958);
and AND3 (N20965, N20963, N1634, N13546);
xor XOR2 (N20966, N20962, N11549);
and AND2 (N20967, N20945, N9111);
not NOT1 (N20968, N20956);
buf BUF1 (N20969, N20967);
nor NOR4 (N20970, N20959, N9405, N1523, N452);
or OR2 (N20971, N20949, N12106);
and AND3 (N20972, N20968, N45, N16884);
not NOT1 (N20973, N20921);
and AND2 (N20974, N20966, N16125);
or OR2 (N20975, N20971, N597);
and AND4 (N20976, N20969, N13775, N18736, N8193);
and AND4 (N20977, N20970, N15795, N12754, N6294);
buf BUF1 (N20978, N20965);
and AND4 (N20979, N20972, N16015, N116, N9611);
not NOT1 (N20980, N20979);
nor NOR3 (N20981, N20955, N15223, N3132);
not NOT1 (N20982, N20978);
or OR4 (N20983, N20964, N3479, N17221, N11036);
xor XOR2 (N20984, N20982, N8311);
buf BUF1 (N20985, N20981);
buf BUF1 (N20986, N20984);
or OR4 (N20987, N20975, N4641, N11919, N2848);
nor NOR2 (N20988, N20974, N981);
xor XOR2 (N20989, N20977, N20791);
and AND2 (N20990, N20973, N15494);
nand NAND4 (N20991, N20983, N7567, N3221, N5300);
not NOT1 (N20992, N20988);
nor NOR2 (N20993, N20960, N17604);
buf BUF1 (N20994, N20990);
not NOT1 (N20995, N20991);
buf BUF1 (N20996, N20976);
nand NAND3 (N20997, N20989, N17192, N7874);
nand NAND4 (N20998, N20994, N5591, N12572, N2985);
nor NOR3 (N20999, N20995, N3604, N3476);
buf BUF1 (N21000, N20986);
buf BUF1 (N21001, N20987);
not NOT1 (N21002, N20999);
xor XOR2 (N21003, N21002, N7291);
or OR3 (N21004, N20993, N19350, N15063);
or OR3 (N21005, N20998, N9327, N8408);
xor XOR2 (N21006, N21001, N13214);
buf BUF1 (N21007, N20997);
nor NOR2 (N21008, N21000, N10008);
and AND2 (N21009, N21007, N18348);
and AND3 (N21010, N20992, N9302, N12582);
not NOT1 (N21011, N21006);
nor NOR3 (N21012, N21011, N15574, N15304);
not NOT1 (N21013, N21005);
buf BUF1 (N21014, N21008);
or OR4 (N21015, N20996, N9302, N1586, N2920);
nand NAND3 (N21016, N21013, N11780, N1022);
nor NOR3 (N21017, N21014, N20374, N5684);
xor XOR2 (N21018, N21017, N14958);
buf BUF1 (N21019, N21012);
and AND2 (N21020, N21010, N8153);
nor NOR4 (N21021, N21009, N575, N19140, N13779);
nor NOR2 (N21022, N21018, N2978);
or OR3 (N21023, N21004, N12255, N17580);
nand NAND4 (N21024, N21019, N12730, N14891, N14115);
not NOT1 (N21025, N21003);
xor XOR2 (N21026, N21020, N1252);
nor NOR2 (N21027, N21023, N6211);
nor NOR4 (N21028, N21024, N2198, N20649, N9359);
nand NAND2 (N21029, N20980, N13156);
not NOT1 (N21030, N21028);
buf BUF1 (N21031, N21025);
xor XOR2 (N21032, N21030, N11349);
xor XOR2 (N21033, N21027, N3993);
or OR4 (N21034, N21031, N6414, N1558, N15895);
buf BUF1 (N21035, N21033);
not NOT1 (N21036, N21022);
not NOT1 (N21037, N21034);
not NOT1 (N21038, N21015);
or OR2 (N21039, N21026, N12241);
and AND4 (N21040, N21038, N4831, N1040, N2503);
and AND2 (N21041, N21039, N14424);
buf BUF1 (N21042, N21029);
buf BUF1 (N21043, N21032);
nor NOR4 (N21044, N21035, N12717, N2704, N14519);
nor NOR2 (N21045, N21043, N6852);
and AND4 (N21046, N21036, N9637, N2283, N2828);
or OR4 (N21047, N21045, N4722, N20361, N13381);
or OR2 (N21048, N21016, N4373);
buf BUF1 (N21049, N21042);
nor NOR4 (N21050, N20985, N3636, N18595, N8715);
nand NAND2 (N21051, N21048, N2828);
nand NAND3 (N21052, N21041, N4879, N18423);
and AND4 (N21053, N21047, N20988, N9256, N15195);
or OR4 (N21054, N21021, N2476, N3777, N5397);
or OR3 (N21055, N21052, N13783, N3300);
buf BUF1 (N21056, N21054);
and AND3 (N21057, N21051, N13917, N10489);
buf BUF1 (N21058, N21046);
or OR4 (N21059, N21053, N15015, N1056, N12640);
nand NAND2 (N21060, N21040, N5534);
or OR2 (N21061, N21057, N19657);
nor NOR2 (N21062, N21050, N17071);
or OR3 (N21063, N21037, N16677, N9660);
xor XOR2 (N21064, N21058, N18080);
buf BUF1 (N21065, N21063);
and AND3 (N21066, N21062, N18873, N14275);
buf BUF1 (N21067, N21066);
or OR4 (N21068, N21056, N11692, N3465, N18350);
nand NAND3 (N21069, N21065, N13734, N14394);
buf BUF1 (N21070, N21044);
not NOT1 (N21071, N21055);
xor XOR2 (N21072, N21071, N12624);
xor XOR2 (N21073, N21059, N17832);
or OR2 (N21074, N21049, N9216);
nand NAND4 (N21075, N21061, N11179, N14751, N15977);
and AND4 (N21076, N21072, N5957, N21014, N5641);
nor NOR4 (N21077, N21070, N16179, N11487, N12709);
and AND3 (N21078, N21068, N2125, N16384);
nor NOR4 (N21079, N21076, N19050, N15380, N17875);
xor XOR2 (N21080, N21078, N6887);
not NOT1 (N21081, N21073);
or OR3 (N21082, N21074, N2719, N11232);
nor NOR2 (N21083, N21077, N18149);
and AND4 (N21084, N21081, N20693, N5477, N17659);
and AND3 (N21085, N21080, N6753, N17588);
or OR2 (N21086, N21064, N5323);
and AND3 (N21087, N21069, N11954, N8916);
xor XOR2 (N21088, N21087, N8891);
not NOT1 (N21089, N21086);
nor NOR4 (N21090, N21085, N16863, N3507, N4667);
and AND4 (N21091, N21075, N5441, N8789, N2920);
and AND4 (N21092, N21090, N14249, N3253, N2725);
nor NOR2 (N21093, N21079, N5349);
not NOT1 (N21094, N21091);
nor NOR2 (N21095, N21084, N16232);
nand NAND2 (N21096, N21082, N2898);
buf BUF1 (N21097, N21094);
buf BUF1 (N21098, N21093);
or OR2 (N21099, N21096, N15995);
nand NAND4 (N21100, N21060, N19576, N3614, N10570);
not NOT1 (N21101, N21088);
not NOT1 (N21102, N21100);
xor XOR2 (N21103, N21099, N1025);
and AND3 (N21104, N21103, N4613, N6374);
or OR3 (N21105, N21092, N629, N4043);
nor NOR4 (N21106, N21067, N15977, N15560, N4615);
nor NOR4 (N21107, N21106, N10190, N16324, N3065);
buf BUF1 (N21108, N21102);
xor XOR2 (N21109, N21107, N508);
nand NAND4 (N21110, N21097, N1540, N13207, N2650);
or OR2 (N21111, N21109, N5657);
nand NAND4 (N21112, N21089, N10212, N861, N1637);
or OR3 (N21113, N21105, N7027, N19368);
not NOT1 (N21114, N21110);
and AND2 (N21115, N21108, N16040);
nand NAND4 (N21116, N21101, N2822, N16940, N18019);
and AND3 (N21117, N21104, N7977, N9167);
nor NOR4 (N21118, N21095, N3027, N3384, N2603);
nor NOR3 (N21119, N21098, N17489, N6810);
buf BUF1 (N21120, N21113);
nand NAND2 (N21121, N21116, N13158);
or OR4 (N21122, N21111, N16157, N3154, N19705);
nand NAND2 (N21123, N21122, N8962);
not NOT1 (N21124, N21083);
and AND4 (N21125, N21124, N18973, N11730, N3254);
xor XOR2 (N21126, N21125, N18043);
buf BUF1 (N21127, N21120);
nand NAND3 (N21128, N21118, N11820, N1058);
nor NOR4 (N21129, N21127, N1851, N8619, N15703);
buf BUF1 (N21130, N21129);
or OR4 (N21131, N21128, N11248, N1953, N18774);
nor NOR3 (N21132, N21121, N19668, N18289);
xor XOR2 (N21133, N21117, N8798);
buf BUF1 (N21134, N21130);
xor XOR2 (N21135, N21119, N8890);
nor NOR2 (N21136, N21114, N13279);
and AND2 (N21137, N21131, N13263);
nor NOR4 (N21138, N21115, N3902, N12068, N1953);
not NOT1 (N21139, N21123);
nand NAND2 (N21140, N21139, N10098);
nor NOR2 (N21141, N21132, N20595);
buf BUF1 (N21142, N21137);
buf BUF1 (N21143, N21135);
xor XOR2 (N21144, N21134, N18301);
nand NAND2 (N21145, N21126, N5158);
nor NOR2 (N21146, N21145, N623);
nor NOR4 (N21147, N21136, N3993, N19981, N15885);
and AND3 (N21148, N21147, N18396, N17222);
nand NAND3 (N21149, N21140, N2765, N7520);
nand NAND3 (N21150, N21141, N14827, N8182);
buf BUF1 (N21151, N21142);
xor XOR2 (N21152, N21151, N18645);
buf BUF1 (N21153, N21144);
and AND3 (N21154, N21149, N7889, N5989);
buf BUF1 (N21155, N21146);
nand NAND2 (N21156, N21133, N9495);
and AND4 (N21157, N21153, N12287, N17131, N18203);
not NOT1 (N21158, N21154);
buf BUF1 (N21159, N21152);
buf BUF1 (N21160, N21138);
not NOT1 (N21161, N21157);
nand NAND2 (N21162, N21150, N2461);
and AND2 (N21163, N21159, N20293);
xor XOR2 (N21164, N21163, N5698);
and AND4 (N21165, N21164, N4611, N20459, N6138);
nand NAND3 (N21166, N21155, N13157, N18643);
nand NAND2 (N21167, N21148, N16993);
xor XOR2 (N21168, N21160, N5589);
or OR2 (N21169, N21162, N17559);
nand NAND4 (N21170, N21166, N2254, N14823, N5878);
buf BUF1 (N21171, N21169);
buf BUF1 (N21172, N21158);
and AND2 (N21173, N21172, N17682);
buf BUF1 (N21174, N21161);
xor XOR2 (N21175, N21165, N17246);
nor NOR3 (N21176, N21171, N15592, N13871);
and AND3 (N21177, N21176, N5715, N13146);
nand NAND3 (N21178, N21175, N11608, N2481);
nand NAND4 (N21179, N21156, N6967, N21006, N10270);
nand NAND4 (N21180, N21168, N8138, N20952, N6477);
or OR4 (N21181, N21167, N13052, N3084, N16513);
nor NOR4 (N21182, N21143, N10726, N19397, N6781);
buf BUF1 (N21183, N21181);
buf BUF1 (N21184, N21179);
nand NAND3 (N21185, N21170, N14827, N14331);
and AND2 (N21186, N21180, N17397);
nand NAND4 (N21187, N21112, N4809, N20365, N14473);
xor XOR2 (N21188, N21186, N694);
not NOT1 (N21189, N21185);
xor XOR2 (N21190, N21184, N11050);
xor XOR2 (N21191, N21189, N853);
and AND3 (N21192, N21174, N7834, N13099);
or OR3 (N21193, N21190, N16055, N3963);
xor XOR2 (N21194, N21191, N4186);
not NOT1 (N21195, N21188);
xor XOR2 (N21196, N21183, N11748);
nor NOR2 (N21197, N21182, N5883);
nor NOR2 (N21198, N21193, N16592);
buf BUF1 (N21199, N21178);
nand NAND2 (N21200, N21194, N298);
xor XOR2 (N21201, N21192, N4079);
xor XOR2 (N21202, N21201, N12011);
nor NOR3 (N21203, N21197, N1854, N11565);
not NOT1 (N21204, N21173);
xor XOR2 (N21205, N21199, N2983);
not NOT1 (N21206, N21200);
xor XOR2 (N21207, N21206, N1633);
xor XOR2 (N21208, N21202, N3848);
xor XOR2 (N21209, N21177, N8202);
nand NAND3 (N21210, N21203, N14838, N727);
xor XOR2 (N21211, N21187, N21038);
buf BUF1 (N21212, N21198);
nor NOR3 (N21213, N21210, N7558, N10950);
buf BUF1 (N21214, N21195);
nand NAND4 (N21215, N21211, N20186, N13457, N4710);
xor XOR2 (N21216, N21215, N7482);
and AND4 (N21217, N21214, N5018, N17176, N13869);
and AND4 (N21218, N21196, N4167, N11666, N16922);
nor NOR2 (N21219, N21216, N4421);
buf BUF1 (N21220, N21204);
and AND3 (N21221, N21209, N5670, N10275);
nand NAND4 (N21222, N21208, N1778, N6330, N9249);
nor NOR4 (N21223, N21212, N8307, N20206, N14550);
xor XOR2 (N21224, N21217, N20037);
xor XOR2 (N21225, N21224, N8740);
xor XOR2 (N21226, N21222, N8107);
nor NOR3 (N21227, N21218, N7869, N13541);
buf BUF1 (N21228, N21225);
nand NAND3 (N21229, N21205, N17016, N20667);
nand NAND3 (N21230, N21226, N2203, N5158);
or OR4 (N21231, N21230, N4937, N13898, N18349);
xor XOR2 (N21232, N21229, N8633);
nand NAND4 (N21233, N21228, N11374, N13083, N11273);
or OR4 (N21234, N21232, N15517, N19700, N12907);
or OR4 (N21235, N21221, N19086, N8091, N3245);
and AND2 (N21236, N21234, N2076);
or OR2 (N21237, N21233, N19471);
and AND3 (N21238, N21213, N13434, N12249);
nor NOR2 (N21239, N21231, N9020);
nand NAND3 (N21240, N21237, N15919, N14645);
xor XOR2 (N21241, N21238, N17037);
not NOT1 (N21242, N21236);
and AND2 (N21243, N21223, N12954);
nor NOR3 (N21244, N21240, N5616, N9032);
buf BUF1 (N21245, N21242);
and AND3 (N21246, N21239, N12250, N12292);
not NOT1 (N21247, N21235);
buf BUF1 (N21248, N21241);
buf BUF1 (N21249, N21243);
xor XOR2 (N21250, N21207, N7240);
xor XOR2 (N21251, N21248, N11783);
xor XOR2 (N21252, N21246, N7211);
buf BUF1 (N21253, N21251);
nor NOR4 (N21254, N21247, N17992, N8928, N7375);
not NOT1 (N21255, N21227);
xor XOR2 (N21256, N21252, N11480);
nor NOR3 (N21257, N21250, N13033, N6365);
not NOT1 (N21258, N21249);
xor XOR2 (N21259, N21219, N3649);
xor XOR2 (N21260, N21244, N11204);
buf BUF1 (N21261, N21259);
nor NOR4 (N21262, N21261, N14820, N20291, N13501);
nand NAND2 (N21263, N21260, N15610);
nor NOR3 (N21264, N21220, N18245, N7472);
or OR3 (N21265, N21254, N5618, N15221);
xor XOR2 (N21266, N21256, N9233);
xor XOR2 (N21267, N21258, N19045);
nand NAND2 (N21268, N21265, N18935);
nand NAND2 (N21269, N21253, N8195);
nor NOR4 (N21270, N21255, N18462, N4417, N14455);
nand NAND2 (N21271, N21270, N3978);
buf BUF1 (N21272, N21269);
not NOT1 (N21273, N21264);
nand NAND4 (N21274, N21245, N2849, N13074, N11913);
xor XOR2 (N21275, N21257, N16916);
nand NAND3 (N21276, N21266, N13701, N10425);
nand NAND2 (N21277, N21262, N18907);
nand NAND4 (N21278, N21271, N4048, N17770, N16106);
nor NOR4 (N21279, N21274, N4424, N17833, N2072);
and AND3 (N21280, N21273, N11016, N10744);
or OR4 (N21281, N21279, N18995, N7533, N7596);
nand NAND2 (N21282, N21275, N9647);
buf BUF1 (N21283, N21281);
buf BUF1 (N21284, N21268);
nor NOR2 (N21285, N21280, N17698);
buf BUF1 (N21286, N21278);
and AND4 (N21287, N21286, N20575, N7324, N18848);
not NOT1 (N21288, N21272);
buf BUF1 (N21289, N21283);
buf BUF1 (N21290, N21276);
or OR3 (N21291, N21267, N9582, N15253);
or OR2 (N21292, N21287, N9608);
nand NAND2 (N21293, N21291, N8334);
xor XOR2 (N21294, N21282, N8842);
or OR3 (N21295, N21277, N15508, N17469);
xor XOR2 (N21296, N21295, N12638);
or OR4 (N21297, N21289, N8109, N10934, N1285);
or OR3 (N21298, N21284, N9794, N8750);
nor NOR3 (N21299, N21288, N15295, N5044);
and AND2 (N21300, N21298, N1286);
xor XOR2 (N21301, N21299, N17269);
nand NAND4 (N21302, N21292, N6349, N10100, N18212);
or OR3 (N21303, N21301, N10540, N14237);
nor NOR3 (N21304, N21296, N16180, N10791);
or OR2 (N21305, N21304, N8526);
not NOT1 (N21306, N21285);
xor XOR2 (N21307, N21263, N19575);
nand NAND3 (N21308, N21300, N197, N20552);
or OR2 (N21309, N21303, N3839);
nor NOR2 (N21310, N21305, N18303);
nand NAND4 (N21311, N21302, N15729, N2090, N16885);
and AND2 (N21312, N21294, N16300);
or OR4 (N21313, N21308, N8226, N8706, N4850);
and AND2 (N21314, N21312, N13424);
nand NAND3 (N21315, N21311, N9317, N13812);
not NOT1 (N21316, N21306);
not NOT1 (N21317, N21307);
and AND4 (N21318, N21297, N8417, N19576, N19440);
and AND4 (N21319, N21315, N3951, N20701, N3459);
nor NOR4 (N21320, N21317, N19099, N5605, N20144);
nand NAND2 (N21321, N21316, N3972);
nand NAND4 (N21322, N21318, N16953, N3300, N20086);
or OR2 (N21323, N21310, N20699);
not NOT1 (N21324, N21293);
buf BUF1 (N21325, N21319);
and AND2 (N21326, N21325, N18880);
nor NOR4 (N21327, N21320, N5302, N14893, N15863);
buf BUF1 (N21328, N21290);
nor NOR3 (N21329, N21322, N2755, N2321);
buf BUF1 (N21330, N21326);
not NOT1 (N21331, N21329);
not NOT1 (N21332, N21313);
xor XOR2 (N21333, N21324, N21243);
buf BUF1 (N21334, N21332);
or OR3 (N21335, N21327, N10736, N13278);
or OR2 (N21336, N21335, N7454);
and AND2 (N21337, N21333, N6744);
nand NAND4 (N21338, N21328, N18785, N17723, N1651);
nor NOR2 (N21339, N21337, N14788);
or OR4 (N21340, N21339, N4993, N18705, N14075);
xor XOR2 (N21341, N21309, N13298);
nand NAND4 (N21342, N21338, N15079, N6194, N17919);
nand NAND3 (N21343, N21334, N19925, N5568);
nand NAND4 (N21344, N21331, N9527, N10131, N14900);
buf BUF1 (N21345, N21342);
buf BUF1 (N21346, N21336);
buf BUF1 (N21347, N21344);
or OR3 (N21348, N21340, N9748, N10741);
buf BUF1 (N21349, N21321);
not NOT1 (N21350, N21341);
not NOT1 (N21351, N21345);
nand NAND3 (N21352, N21343, N2328, N17926);
nor NOR3 (N21353, N21349, N2907, N3930);
nor NOR3 (N21354, N21347, N15383, N7972);
and AND3 (N21355, N21330, N6113, N12253);
nand NAND4 (N21356, N21352, N11259, N13272, N16256);
and AND3 (N21357, N21323, N6350, N14421);
nand NAND4 (N21358, N21346, N453, N1746, N17015);
xor XOR2 (N21359, N21348, N7336);
buf BUF1 (N21360, N21359);
nor NOR3 (N21361, N21356, N9776, N3252);
buf BUF1 (N21362, N21354);
nand NAND3 (N21363, N21361, N5754, N4967);
and AND3 (N21364, N21353, N19815, N240);
not NOT1 (N21365, N21314);
nor NOR2 (N21366, N21357, N5713);
or OR2 (N21367, N21355, N11871);
and AND3 (N21368, N21366, N9818, N314);
and AND4 (N21369, N21351, N14843, N9779, N21233);
nand NAND4 (N21370, N21350, N17545, N8014, N16272);
not NOT1 (N21371, N21364);
and AND4 (N21372, N21368, N16778, N6035, N3391);
nand NAND4 (N21373, N21372, N8483, N9814, N10918);
or OR2 (N21374, N21371, N7658);
nor NOR3 (N21375, N21365, N17758, N11601);
or OR2 (N21376, N21374, N20785);
nand NAND4 (N21377, N21375, N20873, N13079, N9545);
or OR2 (N21378, N21376, N744);
not NOT1 (N21379, N21363);
xor XOR2 (N21380, N21378, N11925);
xor XOR2 (N21381, N21360, N6681);
not NOT1 (N21382, N21373);
not NOT1 (N21383, N21382);
and AND3 (N21384, N21369, N13603, N12182);
not NOT1 (N21385, N21358);
not NOT1 (N21386, N21370);
not NOT1 (N21387, N21383);
nor NOR4 (N21388, N21377, N7661, N12546, N2877);
nor NOR4 (N21389, N21385, N1550, N15972, N12423);
xor XOR2 (N21390, N21389, N6976);
xor XOR2 (N21391, N21380, N21148);
xor XOR2 (N21392, N21367, N12370);
xor XOR2 (N21393, N21362, N20247);
and AND4 (N21394, N21390, N11454, N19524, N11421);
or OR3 (N21395, N21391, N11740, N10340);
and AND4 (N21396, N21393, N16482, N16215, N19741);
buf BUF1 (N21397, N21386);
xor XOR2 (N21398, N21395, N1424);
buf BUF1 (N21399, N21381);
buf BUF1 (N21400, N21388);
xor XOR2 (N21401, N21397, N9255);
nand NAND3 (N21402, N21396, N11464, N8014);
buf BUF1 (N21403, N21394);
xor XOR2 (N21404, N21403, N18523);
buf BUF1 (N21405, N21401);
nor NOR4 (N21406, N21398, N20985, N4340, N1598);
xor XOR2 (N21407, N21406, N10536);
nor NOR3 (N21408, N21405, N11137, N2868);
or OR2 (N21409, N21392, N11641);
nor NOR4 (N21410, N21402, N20842, N6708, N9601);
and AND2 (N21411, N21400, N18239);
nand NAND4 (N21412, N21387, N11932, N11029, N13077);
nand NAND3 (N21413, N21399, N16572, N14396);
or OR4 (N21414, N21413, N4500, N18828, N13536);
nand NAND4 (N21415, N21414, N18056, N6465, N6281);
or OR4 (N21416, N21409, N11775, N17941, N793);
buf BUF1 (N21417, N21379);
or OR4 (N21418, N21416, N5550, N4242, N16832);
not NOT1 (N21419, N21412);
nand NAND3 (N21420, N21411, N60, N11665);
nand NAND4 (N21421, N21407, N17771, N18919, N7319);
not NOT1 (N21422, N21408);
xor XOR2 (N21423, N21420, N6436);
nor NOR3 (N21424, N21404, N5649, N1488);
and AND4 (N21425, N21424, N2007, N4791, N12905);
or OR3 (N21426, N21419, N8012, N3326);
nor NOR2 (N21427, N21384, N316);
or OR2 (N21428, N21421, N4552);
or OR3 (N21429, N21418, N20726, N8796);
not NOT1 (N21430, N21417);
nand NAND4 (N21431, N21422, N6123, N20315, N16776);
not NOT1 (N21432, N21415);
and AND4 (N21433, N21430, N15059, N16236, N1042);
or OR2 (N21434, N21431, N15013);
xor XOR2 (N21435, N21429, N20376);
buf BUF1 (N21436, N21433);
buf BUF1 (N21437, N21423);
and AND3 (N21438, N21434, N18697, N15288);
and AND4 (N21439, N21425, N8677, N15167, N14527);
or OR4 (N21440, N21435, N13359, N6024, N20221);
buf BUF1 (N21441, N21428);
and AND3 (N21442, N21432, N143, N18999);
and AND3 (N21443, N21441, N10211, N3491);
xor XOR2 (N21444, N21443, N13039);
not NOT1 (N21445, N21444);
nand NAND2 (N21446, N21445, N12805);
xor XOR2 (N21447, N21442, N1634);
nand NAND4 (N21448, N21438, N1154, N13307, N9774);
and AND2 (N21449, N21439, N7496);
or OR3 (N21450, N21427, N10971, N5568);
nor NOR2 (N21451, N21426, N13242);
and AND2 (N21452, N21450, N7413);
nor NOR3 (N21453, N21451, N20733, N1700);
buf BUF1 (N21454, N21440);
nand NAND3 (N21455, N21437, N15847, N12592);
and AND4 (N21456, N21410, N4185, N70, N9442);
nor NOR4 (N21457, N21453, N5148, N3846, N4659);
or OR2 (N21458, N21447, N10918);
buf BUF1 (N21459, N21446);
and AND3 (N21460, N21457, N15747, N6687);
buf BUF1 (N21461, N21448);
xor XOR2 (N21462, N21436, N19145);
or OR3 (N21463, N21456, N11655, N21143);
xor XOR2 (N21464, N21463, N4368);
buf BUF1 (N21465, N21464);
or OR2 (N21466, N21462, N21090);
not NOT1 (N21467, N21455);
nand NAND4 (N21468, N21454, N15577, N5451, N13083);
buf BUF1 (N21469, N21449);
nand NAND2 (N21470, N21467, N18199);
not NOT1 (N21471, N21458);
and AND4 (N21472, N21460, N17731, N3247, N3655);
buf BUF1 (N21473, N21471);
buf BUF1 (N21474, N21469);
nand NAND4 (N21475, N21474, N708, N18512, N8839);
nor NOR3 (N21476, N21452, N3139, N18809);
and AND2 (N21477, N21466, N5909);
nand NAND4 (N21478, N21461, N877, N11554, N5553);
nand NAND3 (N21479, N21468, N7793, N2444);
or OR3 (N21480, N21476, N5350, N18635);
and AND2 (N21481, N21473, N15442);
and AND3 (N21482, N21478, N1349, N16002);
or OR4 (N21483, N21465, N20989, N9311, N2320);
not NOT1 (N21484, N21479);
buf BUF1 (N21485, N21480);
xor XOR2 (N21486, N21472, N14713);
buf BUF1 (N21487, N21475);
buf BUF1 (N21488, N21484);
nand NAND2 (N21489, N21488, N3917);
nor NOR4 (N21490, N21470, N8114, N468, N16787);
nor NOR4 (N21491, N21485, N3714, N18018, N20751);
not NOT1 (N21492, N21490);
buf BUF1 (N21493, N21491);
or OR4 (N21494, N21492, N8708, N20552, N15209);
and AND3 (N21495, N21493, N6308, N2593);
or OR3 (N21496, N21482, N16497, N740);
nand NAND2 (N21497, N21495, N13220);
xor XOR2 (N21498, N21489, N4610);
and AND2 (N21499, N21483, N18233);
nor NOR2 (N21500, N21496, N8584);
or OR4 (N21501, N21498, N17158, N17763, N17665);
and AND2 (N21502, N21501, N7554);
nor NOR4 (N21503, N21477, N12146, N2292, N1402);
not NOT1 (N21504, N21503);
or OR4 (N21505, N21499, N15944, N13133, N8324);
nand NAND2 (N21506, N21504, N16780);
xor XOR2 (N21507, N21506, N151);
not NOT1 (N21508, N21500);
buf BUF1 (N21509, N21487);
buf BUF1 (N21510, N21508);
buf BUF1 (N21511, N21459);
or OR3 (N21512, N21502, N9142, N14408);
not NOT1 (N21513, N21507);
nor NOR3 (N21514, N21512, N19245, N8053);
xor XOR2 (N21515, N21514, N14182);
xor XOR2 (N21516, N21510, N842);
buf BUF1 (N21517, N21511);
nand NAND3 (N21518, N21513, N15589, N17331);
nor NOR2 (N21519, N21494, N3284);
nor NOR3 (N21520, N21509, N15158, N18302);
nor NOR2 (N21521, N21486, N4419);
nand NAND2 (N21522, N21517, N16870);
nand NAND3 (N21523, N21521, N8080, N13712);
buf BUF1 (N21524, N21522);
xor XOR2 (N21525, N21518, N19620);
and AND2 (N21526, N21523, N14210);
xor XOR2 (N21527, N21497, N5570);
nand NAND4 (N21528, N21519, N5343, N9153, N1398);
xor XOR2 (N21529, N21505, N10068);
buf BUF1 (N21530, N21527);
and AND4 (N21531, N21528, N18232, N9264, N2215);
or OR3 (N21532, N21531, N10399, N665);
buf BUF1 (N21533, N21515);
xor XOR2 (N21534, N21524, N11519);
buf BUF1 (N21535, N21529);
or OR2 (N21536, N21525, N5629);
and AND3 (N21537, N21533, N6954, N18423);
xor XOR2 (N21538, N21481, N1226);
xor XOR2 (N21539, N21535, N459);
nand NAND3 (N21540, N21520, N3193, N2534);
or OR3 (N21541, N21536, N13041, N2240);
nor NOR4 (N21542, N21532, N3242, N13056, N11794);
or OR3 (N21543, N21534, N15171, N14907);
or OR4 (N21544, N21537, N9863, N14729, N1607);
nand NAND3 (N21545, N21538, N17881, N2064);
not NOT1 (N21546, N21541);
and AND2 (N21547, N21530, N9333);
not NOT1 (N21548, N21539);
xor XOR2 (N21549, N21526, N11554);
not NOT1 (N21550, N21546);
xor XOR2 (N21551, N21544, N14216);
nand NAND4 (N21552, N21547, N12252, N15577, N13700);
or OR4 (N21553, N21551, N7771, N10153, N10596);
xor XOR2 (N21554, N21549, N13613);
or OR3 (N21555, N21552, N17738, N17046);
nor NOR2 (N21556, N21516, N17778);
nor NOR2 (N21557, N21550, N3952);
or OR4 (N21558, N21542, N13651, N20137, N20053);
nand NAND3 (N21559, N21554, N11390, N10625);
not NOT1 (N21560, N21556);
nor NOR2 (N21561, N21558, N864);
buf BUF1 (N21562, N21540);
or OR3 (N21563, N21557, N15755, N9352);
or OR4 (N21564, N21562, N11078, N10157, N641);
nand NAND2 (N21565, N21560, N1977);
buf BUF1 (N21566, N21553);
nand NAND3 (N21567, N21566, N14430, N1522);
nor NOR2 (N21568, N21545, N4770);
buf BUF1 (N21569, N21563);
nand NAND3 (N21570, N21543, N629, N7931);
xor XOR2 (N21571, N21555, N8851);
nand NAND2 (N21572, N21569, N10989);
not NOT1 (N21573, N21561);
not NOT1 (N21574, N21573);
nand NAND2 (N21575, N21564, N820);
or OR3 (N21576, N21565, N11124, N15787);
nor NOR3 (N21577, N21571, N12046, N8025);
and AND2 (N21578, N21574, N17343);
or OR4 (N21579, N21572, N17356, N2596, N19079);
nand NAND2 (N21580, N21567, N9210);
and AND4 (N21581, N21575, N5554, N5405, N14061);
nand NAND3 (N21582, N21570, N5824, N13777);
nor NOR2 (N21583, N21579, N2772);
and AND3 (N21584, N21578, N13860, N19403);
not NOT1 (N21585, N21568);
xor XOR2 (N21586, N21577, N838);
or OR4 (N21587, N21559, N9231, N2905, N3053);
not NOT1 (N21588, N21583);
nand NAND2 (N21589, N21584, N14300);
or OR3 (N21590, N21586, N12583, N3374);
or OR2 (N21591, N21587, N13812);
buf BUF1 (N21592, N21590);
nand NAND2 (N21593, N21576, N20015);
or OR4 (N21594, N21582, N2849, N1510, N1968);
and AND4 (N21595, N21588, N15621, N16158, N12197);
nand NAND4 (N21596, N21593, N8818, N13167, N2473);
buf BUF1 (N21597, N21585);
buf BUF1 (N21598, N21581);
nor NOR3 (N21599, N21597, N5908, N7735);
buf BUF1 (N21600, N21596);
nor NOR3 (N21601, N21591, N10857, N1207);
xor XOR2 (N21602, N21594, N2499);
buf BUF1 (N21603, N21592);
or OR3 (N21604, N21603, N13529, N6484);
or OR4 (N21605, N21589, N3810, N8408, N4993);
not NOT1 (N21606, N21600);
or OR4 (N21607, N21605, N17753, N11660, N4038);
and AND4 (N21608, N21602, N1720, N17754, N4357);
nand NAND3 (N21609, N21601, N15222, N2784);
and AND2 (N21610, N21607, N16178);
buf BUF1 (N21611, N21598);
nand NAND3 (N21612, N21610, N3953, N17891);
buf BUF1 (N21613, N21611);
and AND4 (N21614, N21604, N11623, N5699, N19409);
xor XOR2 (N21615, N21548, N2012);
not NOT1 (N21616, N21615);
or OR3 (N21617, N21616, N3919, N5985);
not NOT1 (N21618, N21608);
nand NAND3 (N21619, N21618, N8461, N18247);
nor NOR4 (N21620, N21580, N16378, N19993, N20877);
buf BUF1 (N21621, N21612);
not NOT1 (N21622, N21606);
xor XOR2 (N21623, N21622, N15201);
not NOT1 (N21624, N21620);
nand NAND2 (N21625, N21614, N15521);
nand NAND2 (N21626, N21619, N17673);
buf BUF1 (N21627, N21624);
not NOT1 (N21628, N21599);
nand NAND2 (N21629, N21623, N15849);
nor NOR4 (N21630, N21625, N7999, N15470, N1181);
and AND3 (N21631, N21630, N21484, N9350);
and AND3 (N21632, N21628, N21541, N10552);
xor XOR2 (N21633, N21632, N19179);
buf BUF1 (N21634, N21627);
not NOT1 (N21635, N21633);
or OR3 (N21636, N21609, N18035, N14117);
or OR2 (N21637, N21595, N16985);
buf BUF1 (N21638, N21634);
nor NOR2 (N21639, N21635, N7080);
xor XOR2 (N21640, N21631, N413);
nand NAND4 (N21641, N21621, N10859, N11687, N1812);
or OR2 (N21642, N21640, N4114);
nand NAND2 (N21643, N21617, N3210);
nor NOR3 (N21644, N21641, N19303, N15116);
and AND4 (N21645, N21626, N15530, N1877, N1389);
or OR4 (N21646, N21639, N5166, N6294, N18301);
or OR3 (N21647, N21637, N6789, N21589);
and AND4 (N21648, N21646, N19618, N5620, N18139);
or OR4 (N21649, N21643, N1259, N12384, N12755);
or OR3 (N21650, N21644, N19360, N16982);
buf BUF1 (N21651, N21649);
nand NAND4 (N21652, N21629, N4549, N16842, N17130);
nand NAND4 (N21653, N21652, N21233, N675, N18657);
nand NAND2 (N21654, N21645, N17829);
not NOT1 (N21655, N21651);
nand NAND4 (N21656, N21655, N9303, N21014, N15651);
nand NAND4 (N21657, N21648, N13064, N20044, N7058);
buf BUF1 (N21658, N21613);
nor NOR2 (N21659, N21658, N18082);
and AND3 (N21660, N21657, N13123, N8164);
xor XOR2 (N21661, N21647, N2550);
buf BUF1 (N21662, N21661);
nand NAND4 (N21663, N21659, N7311, N2331, N8799);
buf BUF1 (N21664, N21650);
or OR4 (N21665, N21662, N4044, N19106, N19910);
buf BUF1 (N21666, N21638);
nand NAND3 (N21667, N21656, N1629, N11305);
or OR4 (N21668, N21667, N538, N19940, N1014);
nand NAND4 (N21669, N21664, N13124, N3173, N866);
and AND4 (N21670, N21653, N13690, N16797, N5814);
buf BUF1 (N21671, N21666);
or OR3 (N21672, N21660, N15783, N1691);
not NOT1 (N21673, N21663);
buf BUF1 (N21674, N21668);
and AND3 (N21675, N21642, N3828, N9425);
or OR3 (N21676, N21674, N1255, N7584);
xor XOR2 (N21677, N21675, N13410);
not NOT1 (N21678, N21669);
not NOT1 (N21679, N21672);
and AND2 (N21680, N21654, N620);
nor NOR3 (N21681, N21636, N8917, N11889);
nor NOR3 (N21682, N21677, N7037, N1506);
or OR2 (N21683, N21676, N19607);
buf BUF1 (N21684, N21671);
nor NOR3 (N21685, N21678, N8601, N14597);
not NOT1 (N21686, N21665);
and AND2 (N21687, N21684, N11815);
xor XOR2 (N21688, N21680, N20217);
nor NOR3 (N21689, N21683, N2428, N8660);
not NOT1 (N21690, N21681);
not NOT1 (N21691, N21670);
nor NOR2 (N21692, N21673, N3741);
and AND4 (N21693, N21692, N8157, N12743, N5505);
not NOT1 (N21694, N21691);
and AND4 (N21695, N21690, N8652, N19651, N15514);
xor XOR2 (N21696, N21682, N11686);
or OR3 (N21697, N21685, N13134, N16740);
not NOT1 (N21698, N21693);
nor NOR2 (N21699, N21694, N17919);
or OR2 (N21700, N21688, N18554);
not NOT1 (N21701, N21689);
buf BUF1 (N21702, N21701);
nand NAND2 (N21703, N21687, N5543);
not NOT1 (N21704, N21686);
or OR3 (N21705, N21700, N20546, N4668);
not NOT1 (N21706, N21705);
buf BUF1 (N21707, N21706);
xor XOR2 (N21708, N21704, N14754);
xor XOR2 (N21709, N21697, N12853);
nor NOR2 (N21710, N21703, N4581);
or OR2 (N21711, N21708, N5752);
or OR2 (N21712, N21698, N2868);
buf BUF1 (N21713, N21699);
xor XOR2 (N21714, N21713, N9914);
or OR4 (N21715, N21696, N1452, N12599, N13901);
buf BUF1 (N21716, N21707);
and AND2 (N21717, N21709, N20252);
nand NAND4 (N21718, N21717, N16739, N16838, N3632);
nand NAND3 (N21719, N21715, N13674, N5671);
not NOT1 (N21720, N21712);
nand NAND3 (N21721, N21695, N13164, N15285);
nand NAND3 (N21722, N21679, N4480, N19947);
not NOT1 (N21723, N21722);
xor XOR2 (N21724, N21721, N20888);
nand NAND2 (N21725, N21702, N10718);
and AND2 (N21726, N21714, N15768);
not NOT1 (N21727, N21720);
and AND2 (N21728, N21727, N3204);
and AND2 (N21729, N21710, N3494);
or OR3 (N21730, N21723, N861, N10815);
buf BUF1 (N21731, N21719);
nor NOR2 (N21732, N21725, N16100);
nand NAND4 (N21733, N21718, N12561, N9090, N18195);
not NOT1 (N21734, N21724);
xor XOR2 (N21735, N21730, N19576);
xor XOR2 (N21736, N21716, N12482);
or OR2 (N21737, N21731, N19455);
nor NOR4 (N21738, N21728, N18345, N7368, N18121);
nand NAND3 (N21739, N21726, N15239, N543);
or OR3 (N21740, N21737, N4708, N2537);
or OR4 (N21741, N21740, N15548, N20078, N8103);
or OR2 (N21742, N21735, N6272);
and AND2 (N21743, N21732, N8934);
or OR2 (N21744, N21736, N18757);
or OR3 (N21745, N21742, N17285, N20850);
xor XOR2 (N21746, N21738, N19799);
nor NOR3 (N21747, N21739, N1407, N21028);
nand NAND2 (N21748, N21734, N16863);
not NOT1 (N21749, N21748);
nor NOR2 (N21750, N21747, N6104);
nand NAND4 (N21751, N21746, N15055, N16358, N15183);
xor XOR2 (N21752, N21729, N12158);
or OR4 (N21753, N21750, N6277, N15442, N16857);
nor NOR3 (N21754, N21749, N11159, N17948);
xor XOR2 (N21755, N21744, N13549);
xor XOR2 (N21756, N21711, N17761);
buf BUF1 (N21757, N21751);
and AND4 (N21758, N21756, N1488, N16712, N19458);
nor NOR2 (N21759, N21741, N19145);
and AND3 (N21760, N21752, N592, N7080);
nor NOR2 (N21761, N21733, N5583);
xor XOR2 (N21762, N21758, N7168);
buf BUF1 (N21763, N21754);
not NOT1 (N21764, N21759);
or OR2 (N21765, N21753, N12330);
or OR4 (N21766, N21743, N19389, N9656, N3993);
nand NAND3 (N21767, N21760, N7140, N13449);
nand NAND3 (N21768, N21755, N14049, N20584);
nor NOR4 (N21769, N21763, N14328, N3356, N16758);
or OR3 (N21770, N21767, N10769, N6862);
nand NAND2 (N21771, N21745, N21460);
not NOT1 (N21772, N21765);
not NOT1 (N21773, N21772);
buf BUF1 (N21774, N21773);
or OR2 (N21775, N21774, N847);
or OR4 (N21776, N21769, N13552, N6165, N4662);
nand NAND3 (N21777, N21771, N21719, N194);
nor NOR3 (N21778, N21762, N8692, N20919);
not NOT1 (N21779, N21778);
nor NOR2 (N21780, N21777, N799);
nor NOR4 (N21781, N21770, N11756, N10310, N377);
and AND4 (N21782, N21781, N20415, N10527, N13350);
xor XOR2 (N21783, N21780, N6825);
xor XOR2 (N21784, N21779, N11345);
nand NAND3 (N21785, N21764, N6073, N1417);
or OR2 (N21786, N21784, N364);
not NOT1 (N21787, N21766);
not NOT1 (N21788, N21783);
and AND4 (N21789, N21788, N19167, N18140, N18975);
not NOT1 (N21790, N21786);
and AND2 (N21791, N21776, N16549);
nor NOR3 (N21792, N21789, N5969, N8091);
xor XOR2 (N21793, N21785, N15224);
nor NOR3 (N21794, N21775, N14190, N12798);
nor NOR2 (N21795, N21787, N1308);
nor NOR3 (N21796, N21791, N17137, N8002);
xor XOR2 (N21797, N21794, N4484);
xor XOR2 (N21798, N21761, N18697);
and AND3 (N21799, N21797, N10371, N20471);
buf BUF1 (N21800, N21782);
or OR2 (N21801, N21757, N4445);
buf BUF1 (N21802, N21793);
nor NOR3 (N21803, N21768, N11730, N4150);
nor NOR2 (N21804, N21803, N7948);
xor XOR2 (N21805, N21798, N3640);
nand NAND3 (N21806, N21801, N2979, N12524);
nor NOR4 (N21807, N21800, N17470, N11701, N17326);
not NOT1 (N21808, N21807);
buf BUF1 (N21809, N21805);
nand NAND2 (N21810, N21790, N16140);
and AND2 (N21811, N21804, N8240);
not NOT1 (N21812, N21810);
not NOT1 (N21813, N21811);
or OR2 (N21814, N21796, N7923);
nor NOR2 (N21815, N21806, N19811);
and AND2 (N21816, N21813, N20341);
buf BUF1 (N21817, N21802);
nor NOR3 (N21818, N21799, N3580, N19414);
not NOT1 (N21819, N21816);
nor NOR3 (N21820, N21819, N15988, N15799);
not NOT1 (N21821, N21795);
not NOT1 (N21822, N21817);
buf BUF1 (N21823, N21812);
nor NOR2 (N21824, N21792, N5496);
nand NAND2 (N21825, N21814, N14617);
nor NOR4 (N21826, N21824, N2234, N5100, N20802);
or OR3 (N21827, N21820, N1551, N18697);
nor NOR2 (N21828, N21822, N5202);
nand NAND3 (N21829, N21823, N203, N5515);
or OR2 (N21830, N21818, N6269);
and AND4 (N21831, N21829, N17040, N7014, N15143);
buf BUF1 (N21832, N21826);
nand NAND4 (N21833, N21827, N3297, N3242, N12705);
nand NAND3 (N21834, N21821, N9258, N14575);
not NOT1 (N21835, N21834);
and AND3 (N21836, N21828, N6045, N14801);
or OR3 (N21837, N21815, N14226, N19681);
buf BUF1 (N21838, N21830);
and AND3 (N21839, N21825, N17790, N15613);
buf BUF1 (N21840, N21808);
nand NAND4 (N21841, N21838, N3868, N11847, N17755);
buf BUF1 (N21842, N21809);
nand NAND4 (N21843, N21833, N15565, N18889, N19007);
xor XOR2 (N21844, N21841, N20708);
xor XOR2 (N21845, N21836, N20148);
not NOT1 (N21846, N21835);
or OR2 (N21847, N21844, N15513);
nor NOR3 (N21848, N21837, N17792, N14835);
xor XOR2 (N21849, N21842, N19075);
and AND2 (N21850, N21831, N15455);
or OR4 (N21851, N21849, N11763, N18135, N16865);
not NOT1 (N21852, N21840);
buf BUF1 (N21853, N21847);
nor NOR2 (N21854, N21848, N1602);
xor XOR2 (N21855, N21839, N15551);
or OR2 (N21856, N21843, N4212);
and AND2 (N21857, N21850, N10167);
and AND3 (N21858, N21854, N14898, N5717);
not NOT1 (N21859, N21855);
buf BUF1 (N21860, N21857);
xor XOR2 (N21861, N21858, N2550);
and AND4 (N21862, N21860, N3064, N1142, N13336);
not NOT1 (N21863, N21851);
or OR4 (N21864, N21853, N870, N9945, N17885);
xor XOR2 (N21865, N21856, N11291);
and AND3 (N21866, N21859, N5651, N3292);
nand NAND4 (N21867, N21861, N14536, N10712, N14369);
nand NAND2 (N21868, N21845, N8726);
xor XOR2 (N21869, N21864, N9645);
nand NAND2 (N21870, N21862, N1708);
not NOT1 (N21871, N21870);
or OR4 (N21872, N21865, N2510, N20180, N9673);
or OR4 (N21873, N21832, N10302, N14858, N21034);
nand NAND4 (N21874, N21872, N12418, N11277, N3460);
and AND2 (N21875, N21846, N6245);
buf BUF1 (N21876, N21869);
nand NAND3 (N21877, N21868, N14582, N17359);
not NOT1 (N21878, N21863);
buf BUF1 (N21879, N21867);
xor XOR2 (N21880, N21876, N9777);
and AND4 (N21881, N21878, N15456, N21613, N8711);
nor NOR3 (N21882, N21873, N3404, N13694);
nand NAND2 (N21883, N21881, N1802);
nand NAND2 (N21884, N21882, N4206);
xor XOR2 (N21885, N21875, N13241);
xor XOR2 (N21886, N21880, N3133);
nand NAND4 (N21887, N21884, N16758, N9910, N2189);
and AND3 (N21888, N21885, N17614, N18418);
buf BUF1 (N21889, N21887);
xor XOR2 (N21890, N21889, N16054);
xor XOR2 (N21891, N21871, N20656);
or OR2 (N21892, N21886, N4904);
and AND3 (N21893, N21852, N16819, N2943);
and AND3 (N21894, N21890, N13925, N11460);
and AND4 (N21895, N21866, N1988, N9592, N8433);
or OR4 (N21896, N21894, N16152, N15122, N13390);
xor XOR2 (N21897, N21891, N14963);
or OR3 (N21898, N21896, N13513, N17044);
or OR4 (N21899, N21879, N10414, N6358, N17698);
and AND2 (N21900, N21897, N10780);
xor XOR2 (N21901, N21888, N9619);
buf BUF1 (N21902, N21893);
nand NAND4 (N21903, N21899, N4908, N6419, N14072);
nor NOR4 (N21904, N21874, N11743, N10701, N5768);
not NOT1 (N21905, N21877);
nor NOR2 (N21906, N21901, N17665);
xor XOR2 (N21907, N21883, N4416);
not NOT1 (N21908, N21903);
and AND2 (N21909, N21902, N17163);
buf BUF1 (N21910, N21907);
not NOT1 (N21911, N21909);
nor NOR4 (N21912, N21895, N6048, N15541, N18324);
not NOT1 (N21913, N21911);
and AND3 (N21914, N21906, N21017, N3583);
not NOT1 (N21915, N21913);
nand NAND3 (N21916, N21912, N578, N3001);
nor NOR2 (N21917, N21904, N21311);
nand NAND2 (N21918, N21915, N5666);
or OR4 (N21919, N21905, N19712, N13413, N1949);
nand NAND4 (N21920, N21914, N6950, N13053, N3704);
nor NOR3 (N21921, N21916, N21152, N20382);
buf BUF1 (N21922, N21900);
not NOT1 (N21923, N21908);
xor XOR2 (N21924, N21921, N2106);
or OR3 (N21925, N21924, N9096, N13378);
xor XOR2 (N21926, N21920, N18100);
nand NAND2 (N21927, N21925, N4240);
nor NOR3 (N21928, N21923, N8459, N1692);
not NOT1 (N21929, N21910);
nand NAND4 (N21930, N21917, N13408, N6978, N11983);
nor NOR2 (N21931, N21926, N17326);
not NOT1 (N21932, N21930);
xor XOR2 (N21933, N21918, N7574);
buf BUF1 (N21934, N21933);
or OR4 (N21935, N21929, N1805, N20048, N12852);
buf BUF1 (N21936, N21934);
buf BUF1 (N21937, N21935);
or OR3 (N21938, N21892, N6196, N782);
not NOT1 (N21939, N21919);
buf BUF1 (N21940, N21938);
nand NAND3 (N21941, N21936, N17955, N15867);
xor XOR2 (N21942, N21931, N11819);
buf BUF1 (N21943, N21942);
nand NAND4 (N21944, N21940, N15974, N4373, N6044);
and AND2 (N21945, N21927, N21594);
xor XOR2 (N21946, N21928, N13436);
nand NAND3 (N21947, N21945, N12379, N1474);
nand NAND3 (N21948, N21947, N1996, N8724);
and AND4 (N21949, N21941, N13733, N6475, N163);
nand NAND3 (N21950, N21939, N8565, N14607);
nand NAND2 (N21951, N21950, N9206);
buf BUF1 (N21952, N21946);
buf BUF1 (N21953, N21943);
nand NAND4 (N21954, N21953, N3095, N21799, N21715);
nor NOR3 (N21955, N21951, N8440, N3470);
buf BUF1 (N21956, N21954);
or OR4 (N21957, N21937, N73, N12147, N3051);
buf BUF1 (N21958, N21949);
and AND4 (N21959, N21955, N11697, N7404, N12436);
nor NOR2 (N21960, N21922, N3979);
or OR3 (N21961, N21944, N15083, N20366);
buf BUF1 (N21962, N21960);
not NOT1 (N21963, N21932);
buf BUF1 (N21964, N21963);
not NOT1 (N21965, N21964);
nor NOR3 (N21966, N21958, N986, N2679);
nand NAND4 (N21967, N21952, N4754, N7528, N10878);
and AND4 (N21968, N21948, N18499, N12976, N6337);
and AND3 (N21969, N21959, N8905, N2839);
buf BUF1 (N21970, N21966);
not NOT1 (N21971, N21969);
or OR4 (N21972, N21962, N16212, N9317, N16731);
xor XOR2 (N21973, N21898, N16995);
not NOT1 (N21974, N21956);
buf BUF1 (N21975, N21971);
not NOT1 (N21976, N21957);
nor NOR2 (N21977, N21975, N4726);
or OR2 (N21978, N21968, N3726);
nor NOR3 (N21979, N21965, N21087, N6013);
not NOT1 (N21980, N21979);
nand NAND2 (N21981, N21973, N10139);
nand NAND2 (N21982, N21976, N7470);
nand NAND3 (N21983, N21977, N11253, N21550);
xor XOR2 (N21984, N21972, N4656);
or OR2 (N21985, N21982, N275);
not NOT1 (N21986, N21970);
nor NOR3 (N21987, N21978, N3056, N7624);
and AND2 (N21988, N21974, N13678);
nor NOR3 (N21989, N21986, N20198, N16243);
or OR2 (N21990, N21984, N11154);
and AND3 (N21991, N21988, N15854, N14948);
nand NAND4 (N21992, N21991, N10827, N11526, N786);
nand NAND3 (N21993, N21989, N4903, N11940);
nor NOR2 (N21994, N21993, N4692);
or OR4 (N21995, N21967, N3232, N15499, N5600);
nand NAND3 (N21996, N21994, N1450, N13724);
buf BUF1 (N21997, N21990);
nand NAND4 (N21998, N21997, N18542, N10602, N13139);
nor NOR3 (N21999, N21980, N19065, N20326);
and AND2 (N22000, N21981, N6081);
not NOT1 (N22001, N21995);
buf BUF1 (N22002, N21987);
nor NOR3 (N22003, N22001, N17251, N6665);
buf BUF1 (N22004, N21961);
nand NAND4 (N22005, N22000, N6079, N1190, N8795);
not NOT1 (N22006, N21985);
nor NOR3 (N22007, N21996, N12316, N18469);
nor NOR2 (N22008, N22003, N4600);
nand NAND2 (N22009, N21992, N15341);
nand NAND3 (N22010, N21999, N8117, N7205);
buf BUF1 (N22011, N22008);
buf BUF1 (N22012, N22009);
and AND4 (N22013, N22010, N11989, N20853, N13618);
or OR2 (N22014, N22012, N19545);
nor NOR2 (N22015, N22013, N5376);
not NOT1 (N22016, N22011);
buf BUF1 (N22017, N21983);
and AND2 (N22018, N22006, N19254);
or OR4 (N22019, N22015, N93, N19676, N11567);
nand NAND3 (N22020, N22007, N1419, N2854);
buf BUF1 (N22021, N22002);
not NOT1 (N22022, N22020);
not NOT1 (N22023, N22017);
or OR3 (N22024, N22014, N4055, N3089);
buf BUF1 (N22025, N22018);
nor NOR4 (N22026, N22022, N9563, N6068, N5829);
and AND2 (N22027, N22025, N21701);
not NOT1 (N22028, N22016);
and AND4 (N22029, N22019, N8259, N8875, N5655);
nor NOR3 (N22030, N22026, N18157, N531);
xor XOR2 (N22031, N22024, N13834);
nor NOR3 (N22032, N22021, N12402, N6644);
nand NAND4 (N22033, N22028, N9102, N11359, N13876);
or OR4 (N22034, N22023, N5992, N5641, N3831);
nor NOR2 (N22035, N22033, N11730);
not NOT1 (N22036, N22030);
nor NOR2 (N22037, N22032, N18403);
nand NAND4 (N22038, N22004, N17802, N4463, N19807);
buf BUF1 (N22039, N22029);
xor XOR2 (N22040, N22039, N20333);
nor NOR4 (N22041, N22037, N18885, N6092, N11109);
and AND4 (N22042, N22041, N5285, N19802, N11139);
buf BUF1 (N22043, N22038);
xor XOR2 (N22044, N22005, N972);
or OR3 (N22045, N22031, N6869, N7244);
nor NOR2 (N22046, N22027, N212);
nand NAND3 (N22047, N22034, N3530, N4906);
nand NAND4 (N22048, N22042, N6134, N12291, N12240);
nand NAND4 (N22049, N22043, N9325, N9709, N21996);
or OR2 (N22050, N22044, N12550);
and AND2 (N22051, N22047, N12993);
nor NOR2 (N22052, N21998, N11545);
and AND4 (N22053, N22040, N6037, N10121, N4540);
and AND3 (N22054, N22052, N3647, N15120);
buf BUF1 (N22055, N22035);
nand NAND4 (N22056, N22046, N6641, N19362, N14295);
not NOT1 (N22057, N22051);
xor XOR2 (N22058, N22056, N14588);
and AND3 (N22059, N22049, N4560, N16806);
xor XOR2 (N22060, N22045, N16165);
nand NAND2 (N22061, N22059, N7154);
and AND3 (N22062, N22053, N16978, N18426);
and AND2 (N22063, N22057, N1853);
buf BUF1 (N22064, N22050);
xor XOR2 (N22065, N22064, N2594);
or OR2 (N22066, N22055, N11002);
nand NAND4 (N22067, N22062, N17695, N17936, N1051);
xor XOR2 (N22068, N22063, N13062);
nor NOR2 (N22069, N22067, N8186);
buf BUF1 (N22070, N22068);
and AND4 (N22071, N22054, N5719, N19378, N5338);
xor XOR2 (N22072, N22066, N17398);
not NOT1 (N22073, N22036);
nor NOR2 (N22074, N22070, N3092);
and AND3 (N22075, N22073, N16615, N3941);
not NOT1 (N22076, N22060);
not NOT1 (N22077, N22071);
nand NAND3 (N22078, N22077, N5575, N16778);
and AND2 (N22079, N22072, N20476);
nor NOR3 (N22080, N22078, N19931, N4399);
nor NOR2 (N22081, N22075, N14611);
buf BUF1 (N22082, N22081);
or OR3 (N22083, N22080, N2330, N18779);
buf BUF1 (N22084, N22065);
or OR4 (N22085, N22061, N3495, N8031, N238);
or OR4 (N22086, N22079, N8783, N20112, N2485);
nor NOR3 (N22087, N22074, N16486, N14604);
nor NOR4 (N22088, N22086, N14820, N17398, N17008);
nor NOR4 (N22089, N22058, N42, N16802, N11221);
and AND2 (N22090, N22089, N18924);
buf BUF1 (N22091, N22076);
or OR4 (N22092, N22083, N2464, N8486, N8683);
nand NAND3 (N22093, N22088, N17886, N10);
or OR4 (N22094, N22092, N9630, N14129, N15896);
buf BUF1 (N22095, N22093);
or OR3 (N22096, N22085, N15810, N14135);
nor NOR4 (N22097, N22082, N10169, N15600, N15390);
and AND3 (N22098, N22090, N16647, N17749);
or OR4 (N22099, N22069, N12734, N13616, N7766);
not NOT1 (N22100, N22096);
buf BUF1 (N22101, N22099);
or OR3 (N22102, N22097, N8640, N11303);
or OR2 (N22103, N22095, N9781);
buf BUF1 (N22104, N22084);
or OR2 (N22105, N22102, N896);
nor NOR4 (N22106, N22104, N9527, N3829, N3278);
xor XOR2 (N22107, N22087, N2954);
nor NOR3 (N22108, N22106, N13902, N12120);
or OR4 (N22109, N22091, N1817, N20287, N5227);
or OR4 (N22110, N22101, N18627, N3123, N2203);
xor XOR2 (N22111, N22048, N2681);
and AND4 (N22112, N22110, N10825, N16002, N21609);
and AND4 (N22113, N22098, N17946, N15082, N2352);
buf BUF1 (N22114, N22113);
nor NOR4 (N22115, N22109, N5110, N6368, N17658);
buf BUF1 (N22116, N22108);
nand NAND2 (N22117, N22116, N94);
nor NOR2 (N22118, N22107, N16786);
and AND2 (N22119, N22100, N5820);
buf BUF1 (N22120, N22112);
nand NAND4 (N22121, N22111, N11903, N6797, N20516);
nand NAND4 (N22122, N22094, N16149, N3264, N7168);
nor NOR4 (N22123, N22115, N10927, N6207, N8138);
buf BUF1 (N22124, N22105);
nand NAND2 (N22125, N22117, N8288);
nor NOR3 (N22126, N22121, N2336, N9692);
or OR3 (N22127, N22120, N12021, N15029);
buf BUF1 (N22128, N22126);
xor XOR2 (N22129, N22128, N12067);
xor XOR2 (N22130, N22125, N6836);
xor XOR2 (N22131, N22130, N582);
nand NAND3 (N22132, N22131, N1520, N20181);
nand NAND4 (N22133, N22122, N6941, N21182, N17460);
and AND3 (N22134, N22133, N5147, N17414);
or OR2 (N22135, N22134, N8317);
or OR4 (N22136, N22114, N12552, N6776, N20142);
xor XOR2 (N22137, N22123, N10380);
not NOT1 (N22138, N22129);
not NOT1 (N22139, N22132);
and AND3 (N22140, N22135, N16713, N14363);
not NOT1 (N22141, N22138);
not NOT1 (N22142, N22137);
nor NOR2 (N22143, N22118, N16764);
nand NAND3 (N22144, N22136, N4284, N2501);
buf BUF1 (N22145, N22103);
nor NOR4 (N22146, N22141, N3030, N13073, N8343);
or OR4 (N22147, N22143, N1011, N7578, N14226);
or OR4 (N22148, N22127, N10123, N3621, N2392);
nand NAND3 (N22149, N22140, N6065, N3975);
nor NOR3 (N22150, N22149, N9609, N9249);
or OR4 (N22151, N22124, N7119, N21385, N16400);
not NOT1 (N22152, N22119);
nor NOR3 (N22153, N22144, N121, N2195);
not NOT1 (N22154, N22142);
and AND4 (N22155, N22147, N17735, N14826, N1029);
and AND2 (N22156, N22148, N21865);
xor XOR2 (N22157, N22151, N9771);
nand NAND2 (N22158, N22152, N576);
or OR3 (N22159, N22155, N22129, N7538);
not NOT1 (N22160, N22154);
not NOT1 (N22161, N22153);
or OR2 (N22162, N22161, N5941);
or OR2 (N22163, N22159, N8493);
nor NOR3 (N22164, N22160, N565, N16183);
nor NOR3 (N22165, N22162, N7303, N16720);
nor NOR4 (N22166, N22145, N13040, N8533, N19101);
and AND2 (N22167, N22146, N16362);
buf BUF1 (N22168, N22163);
and AND4 (N22169, N22158, N8264, N14659, N8233);
nand NAND2 (N22170, N22167, N20911);
and AND2 (N22171, N22165, N431);
nand NAND4 (N22172, N22150, N13426, N12238, N21168);
buf BUF1 (N22173, N22156);
nor NOR2 (N22174, N22170, N9115);
and AND3 (N22175, N22157, N133, N14777);
xor XOR2 (N22176, N22173, N19187);
xor XOR2 (N22177, N22172, N12104);
not NOT1 (N22178, N22139);
xor XOR2 (N22179, N22171, N5552);
or OR4 (N22180, N22174, N13821, N17258, N15833);
not NOT1 (N22181, N22180);
and AND3 (N22182, N22178, N16732, N17284);
buf BUF1 (N22183, N22182);
or OR2 (N22184, N22179, N13878);
not NOT1 (N22185, N22166);
xor XOR2 (N22186, N22181, N10967);
buf BUF1 (N22187, N22164);
buf BUF1 (N22188, N22176);
and AND3 (N22189, N22183, N165, N3121);
xor XOR2 (N22190, N22175, N20770);
not NOT1 (N22191, N22185);
and AND4 (N22192, N22187, N11134, N20611, N13299);
buf BUF1 (N22193, N22168);
nand NAND4 (N22194, N22186, N16053, N5292, N13462);
nand NAND3 (N22195, N22184, N10228, N20081);
xor XOR2 (N22196, N22177, N18238);
buf BUF1 (N22197, N22193);
and AND2 (N22198, N22192, N7570);
or OR4 (N22199, N22189, N19308, N18124, N5849);
nor NOR4 (N22200, N22195, N15073, N11286, N8608);
and AND4 (N22201, N22169, N16809, N9955, N19707);
and AND3 (N22202, N22198, N3482, N17845);
not NOT1 (N22203, N22201);
nand NAND4 (N22204, N22203, N13608, N16230, N4969);
nor NOR4 (N22205, N22194, N12136, N20273, N1690);
nand NAND2 (N22206, N22196, N11065);
not NOT1 (N22207, N22206);
nor NOR2 (N22208, N22204, N8976);
xor XOR2 (N22209, N22199, N5711);
not NOT1 (N22210, N22197);
xor XOR2 (N22211, N22205, N20847);
nand NAND4 (N22212, N22202, N15057, N12239, N21020);
xor XOR2 (N22213, N22209, N17123);
nand NAND2 (N22214, N22207, N18478);
xor XOR2 (N22215, N22208, N13394);
buf BUF1 (N22216, N22214);
nand NAND3 (N22217, N22216, N17499, N21491);
not NOT1 (N22218, N22213);
or OR4 (N22219, N22188, N14603, N20740, N5594);
nor NOR4 (N22220, N22215, N16230, N20415, N15210);
or OR3 (N22221, N22212, N8637, N6020);
and AND2 (N22222, N22210, N6999);
and AND4 (N22223, N22190, N17581, N21324, N1472);
nand NAND4 (N22224, N22221, N18959, N2969, N8273);
not NOT1 (N22225, N22200);
buf BUF1 (N22226, N22223);
nand NAND2 (N22227, N22218, N8483);
buf BUF1 (N22228, N22191);
nor NOR4 (N22229, N22227, N3326, N15985, N674);
buf BUF1 (N22230, N22228);
nor NOR3 (N22231, N22225, N1768, N7557);
buf BUF1 (N22232, N22226);
not NOT1 (N22233, N22231);
nand NAND3 (N22234, N22220, N15898, N6568);
not NOT1 (N22235, N22233);
buf BUF1 (N22236, N22224);
nand NAND2 (N22237, N22217, N3290);
xor XOR2 (N22238, N22237, N14563);
buf BUF1 (N22239, N22229);
nand NAND3 (N22240, N22238, N2339, N11683);
xor XOR2 (N22241, N22232, N11736);
nor NOR4 (N22242, N22236, N9670, N7771, N4810);
buf BUF1 (N22243, N22242);
or OR3 (N22244, N22219, N13040, N15688);
buf BUF1 (N22245, N22222);
nor NOR3 (N22246, N22240, N3966, N12813);
or OR3 (N22247, N22230, N2010, N3242);
or OR4 (N22248, N22247, N20967, N17333, N18018);
or OR2 (N22249, N22245, N9274);
nor NOR3 (N22250, N22241, N9100, N5148);
nand NAND2 (N22251, N22246, N17641);
not NOT1 (N22252, N22249);
xor XOR2 (N22253, N22252, N15129);
or OR3 (N22254, N22253, N21561, N3913);
or OR2 (N22255, N22211, N21546);
not NOT1 (N22256, N22250);
nand NAND4 (N22257, N22251, N9837, N3144, N14061);
nand NAND4 (N22258, N22243, N11012, N2270, N13517);
not NOT1 (N22259, N22257);
nand NAND3 (N22260, N22239, N11627, N12659);
or OR3 (N22261, N22244, N17015, N3369);
xor XOR2 (N22262, N22256, N166);
or OR2 (N22263, N22258, N13705);
buf BUF1 (N22264, N22261);
xor XOR2 (N22265, N22263, N19696);
and AND2 (N22266, N22248, N864);
nand NAND3 (N22267, N22254, N5917, N9860);
buf BUF1 (N22268, N22265);
and AND2 (N22269, N22268, N13488);
not NOT1 (N22270, N22255);
nand NAND2 (N22271, N22260, N17677);
or OR2 (N22272, N22269, N21567);
xor XOR2 (N22273, N22259, N8652);
xor XOR2 (N22274, N22272, N1394);
xor XOR2 (N22275, N22271, N11702);
and AND4 (N22276, N22274, N14483, N16010, N7244);
buf BUF1 (N22277, N22234);
not NOT1 (N22278, N22266);
nand NAND3 (N22279, N22276, N21089, N13327);
buf BUF1 (N22280, N22279);
or OR2 (N22281, N22275, N4753);
nor NOR4 (N22282, N22262, N5793, N3004, N3312);
not NOT1 (N22283, N22280);
xor XOR2 (N22284, N22264, N2052);
not NOT1 (N22285, N22278);
buf BUF1 (N22286, N22277);
and AND3 (N22287, N22281, N3578, N22241);
or OR4 (N22288, N22282, N1970, N7078, N7940);
xor XOR2 (N22289, N22267, N3237);
xor XOR2 (N22290, N22284, N1126);
nand NAND3 (N22291, N22287, N13580, N12573);
and AND2 (N22292, N22283, N4433);
not NOT1 (N22293, N22286);
and AND3 (N22294, N22235, N2563, N14734);
buf BUF1 (N22295, N22293);
buf BUF1 (N22296, N22288);
nor NOR2 (N22297, N22285, N16782);
and AND2 (N22298, N22295, N21469);
not NOT1 (N22299, N22296);
buf BUF1 (N22300, N22289);
not NOT1 (N22301, N22290);
or OR3 (N22302, N22300, N5184, N9051);
nor NOR2 (N22303, N22273, N14295);
not NOT1 (N22304, N22303);
or OR4 (N22305, N22304, N17902, N18022, N299);
nand NAND4 (N22306, N22299, N12677, N17018, N6131);
not NOT1 (N22307, N22301);
and AND3 (N22308, N22305, N13448, N19126);
nand NAND3 (N22309, N22292, N16530, N15703);
xor XOR2 (N22310, N22298, N4722);
nand NAND4 (N22311, N22291, N15448, N21319, N13047);
and AND3 (N22312, N22297, N4919, N10718);
nor NOR3 (N22313, N22306, N19405, N12204);
and AND2 (N22314, N22307, N5794);
and AND4 (N22315, N22302, N6985, N16877, N7569);
not NOT1 (N22316, N22314);
buf BUF1 (N22317, N22315);
nor NOR2 (N22318, N22294, N10730);
or OR4 (N22319, N22311, N16937, N21467, N20639);
xor XOR2 (N22320, N22316, N22125);
nand NAND4 (N22321, N22318, N19622, N16055, N419);
and AND4 (N22322, N22313, N4738, N16783, N5339);
buf BUF1 (N22323, N22309);
or OR3 (N22324, N22270, N19040, N13058);
and AND4 (N22325, N22321, N11881, N2790, N19054);
buf BUF1 (N22326, N22324);
not NOT1 (N22327, N22308);
nand NAND4 (N22328, N22325, N21743, N983, N14257);
xor XOR2 (N22329, N22312, N3108);
or OR4 (N22330, N22319, N16618, N17779, N1080);
nand NAND4 (N22331, N22330, N19203, N3311, N20013);
xor XOR2 (N22332, N22328, N18780);
nor NOR4 (N22333, N22317, N432, N21401, N8603);
not NOT1 (N22334, N22322);
buf BUF1 (N22335, N22331);
nor NOR2 (N22336, N22323, N16185);
buf BUF1 (N22337, N22334);
nand NAND2 (N22338, N22320, N997);
not NOT1 (N22339, N22337);
not NOT1 (N22340, N22335);
not NOT1 (N22341, N22332);
not NOT1 (N22342, N22338);
buf BUF1 (N22343, N22327);
buf BUF1 (N22344, N22342);
not NOT1 (N22345, N22333);
nor NOR2 (N22346, N22336, N14292);
xor XOR2 (N22347, N22346, N7734);
xor XOR2 (N22348, N22329, N17705);
xor XOR2 (N22349, N22345, N18190);
nand NAND3 (N22350, N22344, N10503, N9032);
not NOT1 (N22351, N22343);
nor NOR2 (N22352, N22340, N22216);
xor XOR2 (N22353, N22326, N19153);
nor NOR2 (N22354, N22347, N13355);
or OR2 (N22355, N22354, N13353);
xor XOR2 (N22356, N22350, N10968);
nor NOR3 (N22357, N22339, N9714, N2076);
buf BUF1 (N22358, N22356);
or OR2 (N22359, N22349, N460);
nand NAND4 (N22360, N22358, N15027, N3218, N5909);
not NOT1 (N22361, N22360);
buf BUF1 (N22362, N22348);
or OR4 (N22363, N22310, N17355, N14036, N833);
nand NAND3 (N22364, N22357, N221, N12044);
or OR2 (N22365, N22353, N12219);
nor NOR2 (N22366, N22352, N18036);
nor NOR4 (N22367, N22351, N18548, N18974, N20467);
xor XOR2 (N22368, N22361, N14019);
buf BUF1 (N22369, N22367);
not NOT1 (N22370, N22365);
buf BUF1 (N22371, N22363);
and AND4 (N22372, N22370, N17586, N15367, N6322);
and AND3 (N22373, N22362, N3718, N5683);
or OR3 (N22374, N22369, N19778, N2945);
not NOT1 (N22375, N22364);
not NOT1 (N22376, N22372);
xor XOR2 (N22377, N22373, N3155);
and AND4 (N22378, N22359, N8446, N8491, N13635);
buf BUF1 (N22379, N22371);
not NOT1 (N22380, N22375);
xor XOR2 (N22381, N22376, N18456);
not NOT1 (N22382, N22341);
nor NOR2 (N22383, N22381, N6503);
or OR4 (N22384, N22379, N15047, N4413, N12189);
nand NAND3 (N22385, N22380, N6795, N21324);
not NOT1 (N22386, N22382);
or OR3 (N22387, N22385, N20772, N14132);
buf BUF1 (N22388, N22374);
nor NOR3 (N22389, N22387, N14696, N8650);
and AND2 (N22390, N22368, N1620);
xor XOR2 (N22391, N22366, N4065);
nand NAND4 (N22392, N22389, N21319, N21573, N2029);
and AND4 (N22393, N22383, N11550, N2429, N13757);
nor NOR3 (N22394, N22386, N14463, N5298);
and AND2 (N22395, N22378, N3563);
not NOT1 (N22396, N22391);
nor NOR3 (N22397, N22355, N22114, N21544);
and AND4 (N22398, N22377, N2090, N5400, N19131);
buf BUF1 (N22399, N22393);
not NOT1 (N22400, N22395);
nor NOR4 (N22401, N22397, N9864, N4210, N4917);
or OR3 (N22402, N22401, N14656, N17116);
and AND2 (N22403, N22402, N9682);
or OR4 (N22404, N22388, N18263, N1406, N16657);
xor XOR2 (N22405, N22404, N5862);
xor XOR2 (N22406, N22398, N2490);
and AND4 (N22407, N22400, N19351, N22221, N18936);
xor XOR2 (N22408, N22390, N4447);
not NOT1 (N22409, N22405);
xor XOR2 (N22410, N22394, N50);
not NOT1 (N22411, N22399);
buf BUF1 (N22412, N22411);
or OR3 (N22413, N22406, N21829, N8927);
xor XOR2 (N22414, N22408, N21119);
nor NOR3 (N22415, N22412, N10718, N15724);
nand NAND3 (N22416, N22415, N9808, N6230);
and AND2 (N22417, N22413, N19044);
not NOT1 (N22418, N22416);
or OR3 (N22419, N22392, N13202, N12447);
nand NAND2 (N22420, N22419, N254);
and AND2 (N22421, N22396, N5362);
and AND4 (N22422, N22407, N10297, N20791, N4241);
not NOT1 (N22423, N22418);
not NOT1 (N22424, N22422);
nand NAND4 (N22425, N22410, N20754, N17798, N13464);
nor NOR2 (N22426, N22423, N13259);
nand NAND4 (N22427, N22409, N14406, N20325, N16050);
not NOT1 (N22428, N22417);
xor XOR2 (N22429, N22414, N6817);
and AND2 (N22430, N22403, N5582);
xor XOR2 (N22431, N22424, N10774);
and AND4 (N22432, N22426, N15136, N10379, N10668);
xor XOR2 (N22433, N22431, N11228);
buf BUF1 (N22434, N22384);
buf BUF1 (N22435, N22429);
nor NOR4 (N22436, N22434, N22306, N21489, N17799);
nor NOR2 (N22437, N22425, N15065);
nor NOR4 (N22438, N22427, N1801, N1026, N6613);
and AND4 (N22439, N22432, N3798, N19684, N3749);
nand NAND4 (N22440, N22437, N13547, N2779, N11802);
xor XOR2 (N22441, N22430, N10647);
nor NOR3 (N22442, N22439, N4881, N7207);
and AND2 (N22443, N22428, N17780);
buf BUF1 (N22444, N22420);
nand NAND3 (N22445, N22440, N11205, N1926);
or OR4 (N22446, N22433, N4410, N19008, N17474);
not NOT1 (N22447, N22444);
buf BUF1 (N22448, N22421);
nor NOR2 (N22449, N22443, N8320);
not NOT1 (N22450, N22442);
nand NAND3 (N22451, N22450, N5263, N10885);
xor XOR2 (N22452, N22447, N14571);
nor NOR4 (N22453, N22438, N4477, N19647, N1266);
nand NAND3 (N22454, N22446, N18423, N8713);
nor NOR3 (N22455, N22454, N12890, N18591);
not NOT1 (N22456, N22452);
buf BUF1 (N22457, N22448);
buf BUF1 (N22458, N22449);
buf BUF1 (N22459, N22457);
and AND4 (N22460, N22455, N15192, N16608, N4026);
not NOT1 (N22461, N22435);
xor XOR2 (N22462, N22445, N6229);
and AND4 (N22463, N22453, N19306, N9671, N11700);
nand NAND3 (N22464, N22451, N20724, N4955);
or OR2 (N22465, N22464, N19465);
buf BUF1 (N22466, N22460);
or OR2 (N22467, N22459, N16165);
xor XOR2 (N22468, N22462, N18949);
nor NOR4 (N22469, N22468, N3053, N16057, N19389);
nor NOR3 (N22470, N22463, N15864, N1987);
buf BUF1 (N22471, N22441);
nor NOR3 (N22472, N22465, N21138, N15141);
or OR4 (N22473, N22470, N3178, N21756, N8679);
nor NOR3 (N22474, N22458, N16867, N9280);
buf BUF1 (N22475, N22474);
nor NOR4 (N22476, N22436, N2495, N8666, N8262);
or OR3 (N22477, N22475, N8628, N8063);
or OR3 (N22478, N22466, N2433, N10380);
xor XOR2 (N22479, N22478, N16414);
xor XOR2 (N22480, N22476, N9466);
and AND2 (N22481, N22469, N75);
nand NAND2 (N22482, N22467, N18186);
xor XOR2 (N22483, N22480, N21590);
not NOT1 (N22484, N22472);
not NOT1 (N22485, N22483);
nand NAND2 (N22486, N22473, N6401);
xor XOR2 (N22487, N22481, N5823);
buf BUF1 (N22488, N22471);
or OR4 (N22489, N22484, N19926, N8734, N17374);
nor NOR2 (N22490, N22488, N21184);
or OR3 (N22491, N22456, N15147, N11900);
nor NOR2 (N22492, N22486, N7943);
or OR2 (N22493, N22487, N7878);
not NOT1 (N22494, N22493);
nor NOR2 (N22495, N22477, N2877);
nand NAND2 (N22496, N22495, N15241);
and AND4 (N22497, N22490, N13275, N2973, N3396);
or OR4 (N22498, N22494, N18633, N4927, N21307);
nor NOR3 (N22499, N22491, N3486, N1680);
nor NOR2 (N22500, N22489, N20384);
nand NAND3 (N22501, N22500, N3762, N14239);
nand NAND3 (N22502, N22461, N19441, N5595);
nor NOR2 (N22503, N22498, N11012);
not NOT1 (N22504, N22479);
xor XOR2 (N22505, N22499, N9301);
not NOT1 (N22506, N22501);
xor XOR2 (N22507, N22502, N16883);
nand NAND4 (N22508, N22482, N288, N4285, N20516);
and AND3 (N22509, N22496, N10354, N1750);
nor NOR2 (N22510, N22508, N21754);
buf BUF1 (N22511, N22509);
buf BUF1 (N22512, N22492);
not NOT1 (N22513, N22512);
nor NOR4 (N22514, N22485, N10313, N8871, N20161);
and AND3 (N22515, N22513, N5739, N5754);
or OR4 (N22516, N22504, N21576, N11759, N20275);
nor NOR3 (N22517, N22497, N1687, N13683);
and AND4 (N22518, N22507, N15496, N15692, N12052);
and AND4 (N22519, N22517, N19948, N18279, N8188);
and AND3 (N22520, N22516, N22151, N4700);
nand NAND3 (N22521, N22505, N19094, N2915);
nor NOR3 (N22522, N22519, N209, N19523);
nor NOR4 (N22523, N22518, N3522, N4468, N10969);
nand NAND4 (N22524, N22523, N14189, N5358, N10171);
not NOT1 (N22525, N22503);
nand NAND3 (N22526, N22520, N16441, N10752);
xor XOR2 (N22527, N22521, N334);
nand NAND2 (N22528, N22525, N18066);
and AND4 (N22529, N22510, N18311, N14593, N8243);
buf BUF1 (N22530, N22527);
nand NAND3 (N22531, N22529, N5689, N6009);
or OR2 (N22532, N22531, N4435);
buf BUF1 (N22533, N22515);
nor NOR4 (N22534, N22506, N10488, N11983, N11738);
nand NAND4 (N22535, N22533, N18046, N14, N18437);
xor XOR2 (N22536, N22526, N18949);
and AND3 (N22537, N22536, N20596, N6983);
nor NOR3 (N22538, N22514, N9455, N19117);
or OR4 (N22539, N22524, N9364, N20701, N15865);
not NOT1 (N22540, N22530);
nor NOR4 (N22541, N22538, N4650, N3720, N13606);
not NOT1 (N22542, N22532);
nand NAND4 (N22543, N22522, N21997, N13695, N4435);
or OR2 (N22544, N22534, N11346);
and AND4 (N22545, N22540, N7790, N10620, N22487);
not NOT1 (N22546, N22537);
or OR4 (N22547, N22546, N4774, N16680, N3825);
or OR4 (N22548, N22528, N11828, N21458, N12847);
xor XOR2 (N22549, N22541, N13083);
and AND2 (N22550, N22542, N1519);
or OR2 (N22551, N22544, N7777);
or OR2 (N22552, N22551, N13894);
nor NOR3 (N22553, N22552, N2655, N12542);
buf BUF1 (N22554, N22539);
nor NOR3 (N22555, N22553, N9235, N13383);
and AND2 (N22556, N22543, N11992);
or OR2 (N22557, N22548, N6873);
nand NAND2 (N22558, N22550, N7678);
nand NAND2 (N22559, N22547, N19681);
buf BUF1 (N22560, N22511);
nor NOR4 (N22561, N22556, N3508, N5472, N4460);
and AND2 (N22562, N22549, N3255);
nand NAND2 (N22563, N22557, N18047);
buf BUF1 (N22564, N22561);
nand NAND2 (N22565, N22555, N2934);
and AND3 (N22566, N22563, N19050, N9767);
not NOT1 (N22567, N22559);
xor XOR2 (N22568, N22558, N1110);
or OR3 (N22569, N22565, N2131, N17755);
nand NAND3 (N22570, N22569, N16364, N3301);
not NOT1 (N22571, N22564);
or OR4 (N22572, N22568, N1806, N4573, N11390);
nor NOR2 (N22573, N22554, N17057);
not NOT1 (N22574, N22560);
nor NOR2 (N22575, N22574, N17736);
and AND2 (N22576, N22567, N13718);
and AND3 (N22577, N22566, N9562, N12755);
xor XOR2 (N22578, N22545, N6858);
xor XOR2 (N22579, N22577, N19092);
nand NAND3 (N22580, N22570, N20189, N16021);
and AND4 (N22581, N22535, N20966, N7547, N11914);
and AND2 (N22582, N22572, N11662);
xor XOR2 (N22583, N22576, N3660);
and AND2 (N22584, N22562, N6385);
nand NAND3 (N22585, N22584, N10691, N10379);
xor XOR2 (N22586, N22573, N11523);
or OR2 (N22587, N22585, N17639);
xor XOR2 (N22588, N22583, N12815);
and AND4 (N22589, N22571, N1421, N2496, N17515);
xor XOR2 (N22590, N22589, N10702);
not NOT1 (N22591, N22582);
xor XOR2 (N22592, N22588, N19583);
xor XOR2 (N22593, N22592, N558);
not NOT1 (N22594, N22578);
xor XOR2 (N22595, N22580, N8145);
or OR4 (N22596, N22590, N20454, N8097, N7047);
or OR4 (N22597, N22587, N20679, N21951, N21112);
nor NOR4 (N22598, N22594, N21418, N17069, N1598);
nand NAND4 (N22599, N22597, N13743, N4297, N5155);
not NOT1 (N22600, N22593);
nand NAND4 (N22601, N22599, N22287, N6504, N7129);
and AND2 (N22602, N22600, N14880);
and AND4 (N22603, N22579, N5723, N10866, N16915);
nand NAND3 (N22604, N22603, N16556, N8341);
and AND3 (N22605, N22586, N6045, N32);
nor NOR2 (N22606, N22596, N16533);
or OR4 (N22607, N22602, N1626, N22043, N16889);
xor XOR2 (N22608, N22591, N15076);
buf BUF1 (N22609, N22606);
nor NOR2 (N22610, N22605, N1000);
buf BUF1 (N22611, N22595);
nor NOR3 (N22612, N22601, N3443, N6662);
buf BUF1 (N22613, N22581);
nand NAND3 (N22614, N22612, N1696, N15016);
buf BUF1 (N22615, N22575);
nor NOR4 (N22616, N22609, N3065, N1673, N9866);
and AND4 (N22617, N22616, N135, N18833, N14377);
nor NOR2 (N22618, N22617, N7093);
buf BUF1 (N22619, N22618);
nor NOR3 (N22620, N22615, N22256, N2583);
buf BUF1 (N22621, N22611);
nand NAND3 (N22622, N22598, N7849, N15309);
nand NAND4 (N22623, N22619, N20254, N18388, N16773);
or OR2 (N22624, N22623, N9815);
not NOT1 (N22625, N22622);
or OR4 (N22626, N22620, N11937, N15457, N9812);
not NOT1 (N22627, N22610);
and AND4 (N22628, N22608, N22120, N10392, N9467);
not NOT1 (N22629, N22621);
or OR2 (N22630, N22627, N16300);
and AND3 (N22631, N22624, N22121, N678);
and AND4 (N22632, N22604, N2295, N10126, N7391);
nand NAND3 (N22633, N22629, N4422, N18585);
xor XOR2 (N22634, N22607, N833);
or OR2 (N22635, N22614, N9147);
xor XOR2 (N22636, N22613, N430);
or OR4 (N22637, N22632, N21833, N14588, N5554);
not NOT1 (N22638, N22628);
xor XOR2 (N22639, N22625, N13459);
or OR3 (N22640, N22634, N12276, N5380);
nor NOR2 (N22641, N22630, N22381);
nand NAND4 (N22642, N22640, N5644, N6535, N13726);
nand NAND2 (N22643, N22642, N10374);
not NOT1 (N22644, N22626);
not NOT1 (N22645, N22633);
and AND2 (N22646, N22636, N1161);
not NOT1 (N22647, N22645);
buf BUF1 (N22648, N22631);
nand NAND3 (N22649, N22647, N2973, N6789);
nor NOR4 (N22650, N22641, N19849, N4427, N7267);
xor XOR2 (N22651, N22638, N14804);
nand NAND4 (N22652, N22643, N12276, N15899, N17131);
or OR4 (N22653, N22646, N22121, N21401, N22355);
xor XOR2 (N22654, N22650, N13415);
xor XOR2 (N22655, N22651, N6628);
not NOT1 (N22656, N22649);
buf BUF1 (N22657, N22655);
xor XOR2 (N22658, N22637, N14313);
not NOT1 (N22659, N22654);
not NOT1 (N22660, N22657);
and AND3 (N22661, N22648, N4356, N20355);
or OR4 (N22662, N22658, N14354, N17558, N5426);
and AND4 (N22663, N22644, N17302, N22125, N21958);
nor NOR4 (N22664, N22652, N8809, N1155, N2429);
xor XOR2 (N22665, N22635, N16563);
nand NAND3 (N22666, N22656, N2486, N7433);
buf BUF1 (N22667, N22659);
buf BUF1 (N22668, N22639);
xor XOR2 (N22669, N22661, N1622);
xor XOR2 (N22670, N22669, N7015);
nand NAND2 (N22671, N22663, N18368);
xor XOR2 (N22672, N22660, N11663);
xor XOR2 (N22673, N22662, N8717);
nand NAND4 (N22674, N22653, N3195, N20370, N2196);
not NOT1 (N22675, N22671);
and AND2 (N22676, N22674, N11862);
nor NOR4 (N22677, N22676, N2921, N9104, N6946);
and AND2 (N22678, N22664, N755);
not NOT1 (N22679, N22673);
not NOT1 (N22680, N22667);
nand NAND3 (N22681, N22672, N19365, N3550);
nand NAND3 (N22682, N22679, N6890, N6988);
not NOT1 (N22683, N22681);
nand NAND4 (N22684, N22665, N3730, N12372, N4212);
and AND2 (N22685, N22684, N12762);
not NOT1 (N22686, N22683);
buf BUF1 (N22687, N22668);
and AND2 (N22688, N22678, N20564);
nand NAND3 (N22689, N22675, N6918, N12433);
not NOT1 (N22690, N22686);
and AND2 (N22691, N22680, N14027);
buf BUF1 (N22692, N22689);
nor NOR2 (N22693, N22691, N1964);
xor XOR2 (N22694, N22677, N15577);
nand NAND2 (N22695, N22682, N6133);
nor NOR2 (N22696, N22692, N10684);
nand NAND3 (N22697, N22687, N14380, N17956);
xor XOR2 (N22698, N22690, N12760);
and AND3 (N22699, N22698, N9913, N7761);
nor NOR2 (N22700, N22693, N10515);
not NOT1 (N22701, N22696);
or OR3 (N22702, N22666, N18595, N12514);
nand NAND3 (N22703, N22699, N9891, N3498);
xor XOR2 (N22704, N22685, N15037);
nand NAND3 (N22705, N22703, N13337, N7507);
not NOT1 (N22706, N22702);
nand NAND4 (N22707, N22694, N17792, N20159, N11006);
buf BUF1 (N22708, N22695);
buf BUF1 (N22709, N22708);
nor NOR2 (N22710, N22709, N15729);
or OR4 (N22711, N22710, N76, N8230, N16241);
or OR4 (N22712, N22697, N22308, N6117, N13218);
nand NAND3 (N22713, N22670, N18394, N4864);
nand NAND3 (N22714, N22704, N1170, N2454);
not NOT1 (N22715, N22706);
or OR2 (N22716, N22715, N20627);
not NOT1 (N22717, N22688);
buf BUF1 (N22718, N22712);
xor XOR2 (N22719, N22700, N2173);
not NOT1 (N22720, N22717);
or OR3 (N22721, N22713, N6953, N17841);
not NOT1 (N22722, N22705);
not NOT1 (N22723, N22719);
xor XOR2 (N22724, N22711, N17861);
not NOT1 (N22725, N22722);
xor XOR2 (N22726, N22725, N18181);
and AND4 (N22727, N22723, N21692, N11120, N15119);
not NOT1 (N22728, N22718);
buf BUF1 (N22729, N22714);
and AND3 (N22730, N22701, N18358, N4183);
or OR4 (N22731, N22727, N13304, N19803, N17429);
and AND4 (N22732, N22724, N6941, N21376, N12296);
buf BUF1 (N22733, N22707);
or OR2 (N22734, N22732, N10303);
buf BUF1 (N22735, N22730);
nand NAND2 (N22736, N22731, N2324);
buf BUF1 (N22737, N22729);
nor NOR4 (N22738, N22733, N18544, N43, N8039);
nand NAND2 (N22739, N22721, N6914);
xor XOR2 (N22740, N22728, N16261);
and AND3 (N22741, N22734, N2129, N16813);
or OR4 (N22742, N22738, N5569, N3672, N19088);
xor XOR2 (N22743, N22737, N9733);
nand NAND2 (N22744, N22743, N6088);
not NOT1 (N22745, N22740);
buf BUF1 (N22746, N22716);
and AND3 (N22747, N22746, N6499, N7525);
nor NOR3 (N22748, N22744, N21557, N8923);
not NOT1 (N22749, N22742);
or OR4 (N22750, N22720, N20881, N21007, N16640);
nor NOR2 (N22751, N22741, N14886);
and AND4 (N22752, N22747, N14741, N14655, N8750);
nor NOR3 (N22753, N22749, N15471, N15668);
and AND4 (N22754, N22753, N20158, N1664, N10392);
buf BUF1 (N22755, N22726);
and AND2 (N22756, N22739, N20366);
nor NOR2 (N22757, N22736, N9205);
or OR3 (N22758, N22750, N9501, N11942);
or OR3 (N22759, N22751, N18239, N66);
nand NAND3 (N22760, N22754, N22636, N22283);
or OR3 (N22761, N22759, N21242, N7309);
buf BUF1 (N22762, N22761);
buf BUF1 (N22763, N22748);
or OR2 (N22764, N22752, N2084);
nor NOR3 (N22765, N22758, N520, N15717);
nor NOR3 (N22766, N22756, N16695, N9744);
and AND4 (N22767, N22760, N9094, N9855, N15904);
buf BUF1 (N22768, N22755);
and AND2 (N22769, N22768, N19171);
buf BUF1 (N22770, N22764);
nand NAND2 (N22771, N22762, N16865);
xor XOR2 (N22772, N22745, N2388);
not NOT1 (N22773, N22767);
or OR2 (N22774, N22765, N9189);
nor NOR3 (N22775, N22774, N5510, N4913);
not NOT1 (N22776, N22766);
not NOT1 (N22777, N22771);
or OR4 (N22778, N22735, N15674, N7921, N9435);
or OR3 (N22779, N22769, N9092, N14041);
nand NAND2 (N22780, N22772, N8085);
or OR4 (N22781, N22763, N3146, N3181, N8906);
or OR4 (N22782, N22773, N15422, N5062, N22389);
xor XOR2 (N22783, N22757, N5756);
and AND4 (N22784, N22782, N11300, N10605, N16188);
buf BUF1 (N22785, N22770);
buf BUF1 (N22786, N22783);
nor NOR2 (N22787, N22778, N20273);
buf BUF1 (N22788, N22777);
nand NAND4 (N22789, N22779, N3278, N5850, N18236);
and AND2 (N22790, N22789, N3797);
or OR2 (N22791, N22787, N2817);
xor XOR2 (N22792, N22776, N17550);
nor NOR3 (N22793, N22786, N6673, N348);
not NOT1 (N22794, N22790);
buf BUF1 (N22795, N22791);
and AND4 (N22796, N22793, N17819, N14692, N627);
or OR3 (N22797, N22796, N7565, N18969);
not NOT1 (N22798, N22784);
and AND4 (N22799, N22792, N15164, N12961, N4149);
and AND3 (N22800, N22780, N2425, N272);
buf BUF1 (N22801, N22785);
buf BUF1 (N22802, N22800);
nand NAND2 (N22803, N22798, N14290);
not NOT1 (N22804, N22788);
and AND3 (N22805, N22804, N732, N17832);
nor NOR3 (N22806, N22775, N17224, N11247);
nor NOR4 (N22807, N22806, N5685, N8543, N12503);
nand NAND3 (N22808, N22807, N3275, N3832);
nand NAND3 (N22809, N22801, N3257, N13118);
xor XOR2 (N22810, N22809, N20495);
or OR3 (N22811, N22799, N14941, N10456);
or OR3 (N22812, N22803, N15484, N9763);
xor XOR2 (N22813, N22795, N22235);
nor NOR3 (N22814, N22811, N14490, N17865);
not NOT1 (N22815, N22805);
not NOT1 (N22816, N22781);
or OR2 (N22817, N22813, N17872);
not NOT1 (N22818, N22815);
nor NOR3 (N22819, N22818, N8367, N22418);
nand NAND4 (N22820, N22819, N16682, N13500, N13788);
not NOT1 (N22821, N22814);
and AND2 (N22822, N22812, N18120);
nand NAND2 (N22823, N22817, N3555);
nand NAND4 (N22824, N22823, N22171, N14923, N13219);
or OR3 (N22825, N22816, N17744, N20080);
nand NAND2 (N22826, N22808, N16560);
and AND3 (N22827, N22810, N7410, N18363);
nor NOR2 (N22828, N22825, N2575);
nand NAND4 (N22829, N22822, N17477, N20916, N16783);
nor NOR3 (N22830, N22824, N15403, N15935);
or OR2 (N22831, N22821, N131);
and AND4 (N22832, N22831, N13477, N10614, N2975);
xor XOR2 (N22833, N22830, N10050);
or OR3 (N22834, N22797, N9408, N9984);
xor XOR2 (N22835, N22802, N5642);
nor NOR2 (N22836, N22834, N5031);
and AND2 (N22837, N22820, N16996);
buf BUF1 (N22838, N22829);
xor XOR2 (N22839, N22835, N1393);
not NOT1 (N22840, N22833);
or OR2 (N22841, N22828, N6079);
not NOT1 (N22842, N22837);
xor XOR2 (N22843, N22838, N10346);
nor NOR3 (N22844, N22832, N4057, N4092);
xor XOR2 (N22845, N22840, N21813);
buf BUF1 (N22846, N22843);
nand NAND4 (N22847, N22846, N16137, N5109, N17978);
or OR3 (N22848, N22839, N16821, N1998);
or OR2 (N22849, N22827, N6673);
nor NOR3 (N22850, N22842, N14832, N15190);
nand NAND2 (N22851, N22850, N19770);
xor XOR2 (N22852, N22845, N7050);
not NOT1 (N22853, N22826);
or OR4 (N22854, N22844, N13789, N12267, N19182);
buf BUF1 (N22855, N22849);
nor NOR3 (N22856, N22848, N15499, N10158);
nand NAND2 (N22857, N22853, N2958);
or OR3 (N22858, N22855, N3983, N16279);
not NOT1 (N22859, N22841);
not NOT1 (N22860, N22852);
nor NOR4 (N22861, N22847, N13786, N22108, N19179);
xor XOR2 (N22862, N22859, N6106);
buf BUF1 (N22863, N22862);
not NOT1 (N22864, N22856);
xor XOR2 (N22865, N22860, N16411);
nor NOR4 (N22866, N22858, N6199, N5736, N5837);
buf BUF1 (N22867, N22865);
not NOT1 (N22868, N22861);
buf BUF1 (N22869, N22866);
nor NOR3 (N22870, N22857, N22730, N8780);
xor XOR2 (N22871, N22851, N17871);
xor XOR2 (N22872, N22868, N16011);
or OR4 (N22873, N22872, N14715, N8783, N19975);
or OR2 (N22874, N22867, N18709);
and AND3 (N22875, N22869, N21726, N2732);
xor XOR2 (N22876, N22836, N11920);
not NOT1 (N22877, N22863);
and AND2 (N22878, N22870, N2408);
nand NAND3 (N22879, N22854, N10409, N20929);
nor NOR3 (N22880, N22871, N9195, N3595);
xor XOR2 (N22881, N22875, N9704);
nand NAND4 (N22882, N22794, N17612, N17373, N20656);
buf BUF1 (N22883, N22880);
or OR4 (N22884, N22876, N1533, N12642, N7941);
and AND3 (N22885, N22883, N22710, N20129);
nand NAND3 (N22886, N22881, N22373, N17360);
nand NAND2 (N22887, N22877, N19950);
nand NAND2 (N22888, N22886, N9116);
nand NAND4 (N22889, N22879, N10837, N6684, N19097);
xor XOR2 (N22890, N22873, N16287);
nand NAND2 (N22891, N22888, N12163);
or OR3 (N22892, N22885, N16831, N13751);
xor XOR2 (N22893, N22864, N5751);
xor XOR2 (N22894, N22882, N16976);
nand NAND3 (N22895, N22890, N15184, N16208);
not NOT1 (N22896, N22887);
buf BUF1 (N22897, N22895);
not NOT1 (N22898, N22874);
xor XOR2 (N22899, N22896, N19236);
nor NOR4 (N22900, N22884, N11297, N6873, N17199);
xor XOR2 (N22901, N22900, N9610);
nor NOR4 (N22902, N22901, N13247, N21805, N14245);
not NOT1 (N22903, N22889);
nand NAND3 (N22904, N22897, N9952, N15284);
xor XOR2 (N22905, N22891, N4136);
nand NAND4 (N22906, N22898, N18395, N17638, N22623);
not NOT1 (N22907, N22899);
and AND2 (N22908, N22907, N17467);
buf BUF1 (N22909, N22906);
buf BUF1 (N22910, N22905);
and AND4 (N22911, N22902, N10866, N9886, N18019);
xor XOR2 (N22912, N22904, N15431);
or OR2 (N22913, N22892, N4712);
nor NOR3 (N22914, N22913, N9861, N7707);
xor XOR2 (N22915, N22894, N8394);
not NOT1 (N22916, N22911);
not NOT1 (N22917, N22916);
nand NAND3 (N22918, N22914, N1414, N19953);
not NOT1 (N22919, N22893);
not NOT1 (N22920, N22909);
nor NOR4 (N22921, N22915, N9728, N7390, N16275);
or OR4 (N22922, N22878, N10279, N13326, N10174);
buf BUF1 (N22923, N22922);
not NOT1 (N22924, N22910);
not NOT1 (N22925, N22924);
buf BUF1 (N22926, N22925);
or OR4 (N22927, N22926, N7689, N2126, N12293);
not NOT1 (N22928, N22923);
and AND3 (N22929, N22921, N1209, N12016);
xor XOR2 (N22930, N22929, N7567);
buf BUF1 (N22931, N22928);
and AND2 (N22932, N22918, N10324);
or OR3 (N22933, N22920, N17176, N22197);
xor XOR2 (N22934, N22927, N2034);
xor XOR2 (N22935, N22932, N22075);
or OR4 (N22936, N22917, N21541, N2255, N16998);
and AND4 (N22937, N22934, N22286, N5273, N1883);
buf BUF1 (N22938, N22903);
and AND2 (N22939, N22937, N5401);
nand NAND2 (N22940, N22931, N19837);
xor XOR2 (N22941, N22939, N19831);
or OR3 (N22942, N22930, N17758, N18307);
buf BUF1 (N22943, N22935);
buf BUF1 (N22944, N22938);
and AND3 (N22945, N22936, N20761, N20587);
and AND3 (N22946, N22933, N18309, N22208);
and AND2 (N22947, N22908, N129);
nand NAND4 (N22948, N22945, N5801, N5179, N13738);
nand NAND2 (N22949, N22942, N22355);
buf BUF1 (N22950, N22912);
buf BUF1 (N22951, N22941);
or OR3 (N22952, N22947, N15226, N12158);
buf BUF1 (N22953, N22951);
xor XOR2 (N22954, N22949, N17767);
nand NAND2 (N22955, N22950, N11121);
nand NAND4 (N22956, N22953, N6899, N20985, N7455);
and AND4 (N22957, N22943, N171, N13828, N18480);
xor XOR2 (N22958, N22952, N17194);
buf BUF1 (N22959, N22957);
or OR3 (N22960, N22944, N18632, N14987);
xor XOR2 (N22961, N22958, N14690);
not NOT1 (N22962, N22961);
or OR3 (N22963, N22959, N4258, N16636);
nand NAND2 (N22964, N22960, N18181);
nor NOR4 (N22965, N22948, N6682, N1379, N15327);
nand NAND2 (N22966, N22963, N12105);
nor NOR4 (N22967, N22964, N10220, N17876, N14198);
buf BUF1 (N22968, N22966);
nor NOR4 (N22969, N22968, N4695, N15303, N6336);
buf BUF1 (N22970, N22965);
not NOT1 (N22971, N22954);
and AND3 (N22972, N22946, N4867, N3422);
not NOT1 (N22973, N22940);
nor NOR3 (N22974, N22973, N13707, N12112);
nor NOR2 (N22975, N22967, N18887);
nor NOR2 (N22976, N22972, N12597);
nand NAND3 (N22977, N22974, N17277, N19214);
not NOT1 (N22978, N22975);
not NOT1 (N22979, N22956);
nand NAND4 (N22980, N22962, N13733, N12813, N6297);
or OR4 (N22981, N22919, N10560, N20750, N14417);
nand NAND4 (N22982, N22981, N21823, N12216, N20966);
or OR4 (N22983, N22977, N19240, N18501, N6252);
or OR3 (N22984, N22955, N8513, N18110);
xor XOR2 (N22985, N22984, N22217);
nand NAND3 (N22986, N22979, N16965, N22633);
nor NOR3 (N22987, N22971, N1532, N11299);
and AND3 (N22988, N22985, N4907, N1126);
or OR3 (N22989, N22982, N1733, N14805);
not NOT1 (N22990, N22986);
xor XOR2 (N22991, N22969, N8125);
nor NOR4 (N22992, N22989, N1549, N16871, N7815);
or OR3 (N22993, N22987, N18103, N12114);
and AND4 (N22994, N22970, N5938, N7203, N7691);
nor NOR3 (N22995, N22988, N20147, N13552);
not NOT1 (N22996, N22992);
xor XOR2 (N22997, N22995, N14450);
nor NOR3 (N22998, N22997, N17392, N7167);
xor XOR2 (N22999, N22993, N16001);
buf BUF1 (N23000, N22990);
and AND3 (N23001, N22994, N5452, N4743);
xor XOR2 (N23002, N22999, N20153);
or OR2 (N23003, N22996, N545);
nor NOR4 (N23004, N22976, N7180, N15570, N19044);
nor NOR4 (N23005, N23001, N9448, N22829, N7751);
nor NOR3 (N23006, N23005, N17084, N5896);
not NOT1 (N23007, N22978);
xor XOR2 (N23008, N22991, N21096);
nand NAND3 (N23009, N23007, N7530, N2142);
and AND4 (N23010, N23002, N8272, N12501, N21073);
not NOT1 (N23011, N23006);
and AND2 (N23012, N23003, N20506);
not NOT1 (N23013, N23011);
buf BUF1 (N23014, N23012);
not NOT1 (N23015, N23004);
not NOT1 (N23016, N23008);
and AND3 (N23017, N23000, N6762, N16940);
nand NAND4 (N23018, N22998, N6760, N19664, N20324);
and AND2 (N23019, N22983, N6319);
and AND4 (N23020, N23017, N19747, N8348, N21082);
or OR3 (N23021, N23014, N2415, N7054);
nor NOR4 (N23022, N23020, N17690, N12656, N17308);
and AND2 (N23023, N23021, N13553);
nand NAND4 (N23024, N23015, N11416, N21900, N18937);
nor NOR4 (N23025, N23023, N14675, N21217, N8413);
xor XOR2 (N23026, N23018, N1995);
nor NOR2 (N23027, N23010, N5581);
nor NOR3 (N23028, N23025, N8092, N3384);
nor NOR2 (N23029, N23027, N18434);
buf BUF1 (N23030, N22980);
and AND2 (N23031, N23022, N22116);
not NOT1 (N23032, N23028);
buf BUF1 (N23033, N23031);
nand NAND4 (N23034, N23024, N21867, N16681, N6319);
or OR3 (N23035, N23016, N2654, N12035);
or OR3 (N23036, N23034, N3226, N1307);
nand NAND2 (N23037, N23030, N20785);
nand NAND3 (N23038, N23036, N22140, N12517);
buf BUF1 (N23039, N23029);
buf BUF1 (N23040, N23033);
or OR2 (N23041, N23037, N3008);
not NOT1 (N23042, N23041);
and AND4 (N23043, N23019, N14852, N11881, N6305);
not NOT1 (N23044, N23009);
nand NAND2 (N23045, N23044, N586);
xor XOR2 (N23046, N23026, N19998);
nand NAND4 (N23047, N23040, N20936, N5130, N22589);
not NOT1 (N23048, N23042);
or OR3 (N23049, N23013, N5295, N21427);
xor XOR2 (N23050, N23039, N10768);
and AND3 (N23051, N23045, N22036, N2784);
not NOT1 (N23052, N23049);
not NOT1 (N23053, N23035);
xor XOR2 (N23054, N23032, N15971);
buf BUF1 (N23055, N23050);
xor XOR2 (N23056, N23053, N16556);
buf BUF1 (N23057, N23043);
nand NAND2 (N23058, N23051, N14968);
or OR4 (N23059, N23047, N17502, N12772, N6668);
nor NOR3 (N23060, N23059, N21417, N10745);
and AND3 (N23061, N23048, N18472, N15282);
nor NOR3 (N23062, N23056, N14733, N9515);
nor NOR2 (N23063, N23062, N12951);
or OR3 (N23064, N23055, N12063, N8440);
and AND2 (N23065, N23054, N1693);
and AND2 (N23066, N23052, N17565);
nand NAND2 (N23067, N23038, N3027);
buf BUF1 (N23068, N23060);
nand NAND3 (N23069, N23065, N22396, N11161);
or OR4 (N23070, N23066, N19504, N17078, N11646);
nor NOR4 (N23071, N23068, N11235, N5828, N135);
and AND4 (N23072, N23061, N5814, N3509, N8950);
or OR3 (N23073, N23046, N16448, N12400);
not NOT1 (N23074, N23070);
nand NAND3 (N23075, N23072, N835, N11002);
nand NAND2 (N23076, N23074, N21855);
nor NOR4 (N23077, N23075, N5076, N6711, N1695);
xor XOR2 (N23078, N23057, N10287);
nand NAND2 (N23079, N23064, N5668);
xor XOR2 (N23080, N23079, N21354);
nand NAND4 (N23081, N23076, N2539, N10534, N15813);
buf BUF1 (N23082, N23058);
not NOT1 (N23083, N23077);
not NOT1 (N23084, N23080);
not NOT1 (N23085, N23084);
nand NAND3 (N23086, N23073, N13507, N8433);
or OR2 (N23087, N23082, N22392);
or OR2 (N23088, N23067, N11923);
or OR2 (N23089, N23078, N2376);
xor XOR2 (N23090, N23087, N17316);
buf BUF1 (N23091, N23063);
nor NOR4 (N23092, N23071, N22046, N2973, N19288);
buf BUF1 (N23093, N23083);
nor NOR3 (N23094, N23086, N5433, N9885);
nand NAND4 (N23095, N23093, N1274, N22295, N11334);
or OR4 (N23096, N23091, N22499, N13882, N15986);
nand NAND4 (N23097, N23096, N13138, N16503, N16227);
or OR4 (N23098, N23085, N4154, N965, N11215);
or OR2 (N23099, N23097, N18887);
xor XOR2 (N23100, N23069, N15334);
or OR4 (N23101, N23099, N9973, N7488, N11389);
or OR2 (N23102, N23081, N14715);
or OR4 (N23103, N23094, N9015, N13798, N11248);
nor NOR4 (N23104, N23098, N21853, N15574, N1537);
nand NAND3 (N23105, N23090, N11951, N561);
not NOT1 (N23106, N23102);
xor XOR2 (N23107, N23103, N11952);
or OR2 (N23108, N23089, N17002);
not NOT1 (N23109, N23105);
not NOT1 (N23110, N23107);
or OR2 (N23111, N23108, N17032);
and AND2 (N23112, N23092, N21527);
and AND2 (N23113, N23104, N1860);
not NOT1 (N23114, N23100);
and AND4 (N23115, N23095, N7201, N4953, N12684);
buf BUF1 (N23116, N23114);
or OR4 (N23117, N23109, N12956, N5763, N20525);
buf BUF1 (N23118, N23117);
not NOT1 (N23119, N23113);
xor XOR2 (N23120, N23106, N6798);
nor NOR2 (N23121, N23112, N6585);
or OR3 (N23122, N23118, N17920, N16553);
buf BUF1 (N23123, N23115);
not NOT1 (N23124, N23101);
or OR3 (N23125, N23123, N12033, N14479);
not NOT1 (N23126, N23122);
not NOT1 (N23127, N23125);
not NOT1 (N23128, N23110);
or OR2 (N23129, N23119, N6197);
nor NOR2 (N23130, N23120, N126);
nor NOR3 (N23131, N23127, N11836, N925);
or OR4 (N23132, N23126, N14257, N2054, N19272);
or OR4 (N23133, N23128, N6991, N7377, N1034);
buf BUF1 (N23134, N23121);
nor NOR3 (N23135, N23130, N15545, N5628);
not NOT1 (N23136, N23133);
nor NOR3 (N23137, N23134, N10433, N19783);
nor NOR2 (N23138, N23088, N3078);
nor NOR3 (N23139, N23116, N5893, N15122);
nor NOR2 (N23140, N23138, N5247);
nand NAND4 (N23141, N23137, N1925, N18081, N7577);
not NOT1 (N23142, N23141);
and AND2 (N23143, N23131, N22826);
nor NOR3 (N23144, N23140, N12761, N12154);
xor XOR2 (N23145, N23142, N10809);
not NOT1 (N23146, N23129);
xor XOR2 (N23147, N23143, N4879);
nand NAND3 (N23148, N23135, N6411, N16561);
or OR4 (N23149, N23111, N15149, N3750, N15267);
buf BUF1 (N23150, N23148);
xor XOR2 (N23151, N23136, N20233);
and AND2 (N23152, N23132, N4354);
and AND3 (N23153, N23151, N18439, N7769);
nor NOR4 (N23154, N23153, N16176, N98, N21352);
nor NOR2 (N23155, N23124, N21732);
nand NAND3 (N23156, N23152, N9568, N3994);
or OR2 (N23157, N23156, N12454);
buf BUF1 (N23158, N23147);
and AND2 (N23159, N23145, N21880);
nor NOR2 (N23160, N23157, N12455);
nand NAND4 (N23161, N23146, N6669, N12961, N22863);
and AND2 (N23162, N23144, N9279);
or OR2 (N23163, N23155, N4592);
not NOT1 (N23164, N23149);
xor XOR2 (N23165, N23164, N5308);
buf BUF1 (N23166, N23165);
buf BUF1 (N23167, N23159);
and AND3 (N23168, N23167, N11554, N10529);
or OR2 (N23169, N23168, N17470);
buf BUF1 (N23170, N23169);
or OR3 (N23171, N23161, N18233, N22603);
xor XOR2 (N23172, N23163, N7281);
not NOT1 (N23173, N23139);
buf BUF1 (N23174, N23150);
not NOT1 (N23175, N23160);
nand NAND4 (N23176, N23174, N9737, N3121, N11953);
or OR3 (N23177, N23171, N20176, N331);
nand NAND3 (N23178, N23173, N9663, N15408);
not NOT1 (N23179, N23158);
nor NOR4 (N23180, N23154, N17762, N5539, N15117);
nand NAND4 (N23181, N23176, N13400, N11994, N10414);
not NOT1 (N23182, N23180);
or OR2 (N23183, N23182, N8159);
and AND2 (N23184, N23177, N23034);
nand NAND3 (N23185, N23181, N3199, N18612);
or OR4 (N23186, N23170, N17577, N1711, N15489);
not NOT1 (N23187, N23185);
nand NAND4 (N23188, N23183, N23077, N17609, N6243);
and AND3 (N23189, N23178, N2604, N11614);
not NOT1 (N23190, N23189);
nor NOR4 (N23191, N23162, N22108, N9041, N23188);
nor NOR4 (N23192, N20778, N22626, N1660, N11311);
xor XOR2 (N23193, N23166, N19588);
nor NOR2 (N23194, N23191, N21132);
not NOT1 (N23195, N23194);
nor NOR3 (N23196, N23187, N19795, N7194);
or OR2 (N23197, N23196, N6401);
buf BUF1 (N23198, N23179);
or OR2 (N23199, N23184, N2760);
nand NAND4 (N23200, N23175, N13895, N11184, N10993);
nand NAND4 (N23201, N23193, N4364, N22726, N13555);
buf BUF1 (N23202, N23186);
or OR2 (N23203, N23190, N10721);
xor XOR2 (N23204, N23197, N937);
not NOT1 (N23205, N23199);
buf BUF1 (N23206, N23205);
and AND4 (N23207, N23206, N13810, N20994, N5070);
or OR3 (N23208, N23172, N16433, N20078);
nand NAND3 (N23209, N23200, N13778, N500);
xor XOR2 (N23210, N23203, N932);
not NOT1 (N23211, N23192);
and AND2 (N23212, N23209, N212);
nand NAND4 (N23213, N23195, N19738, N963, N1191);
or OR3 (N23214, N23210, N13001, N23065);
or OR3 (N23215, N23212, N13614, N14609);
or OR3 (N23216, N23215, N10008, N3408);
buf BUF1 (N23217, N23211);
and AND4 (N23218, N23202, N11087, N11390, N6253);
nor NOR4 (N23219, N23214, N5263, N16940, N6810);
nor NOR3 (N23220, N23198, N6836, N15522);
or OR2 (N23221, N23213, N12872);
not NOT1 (N23222, N23216);
and AND3 (N23223, N23222, N2517, N20266);
or OR3 (N23224, N23207, N20927, N13938);
not NOT1 (N23225, N23201);
buf BUF1 (N23226, N23224);
or OR4 (N23227, N23220, N517, N10647, N16080);
buf BUF1 (N23228, N23208);
not NOT1 (N23229, N23223);
or OR2 (N23230, N23228, N22701);
nor NOR3 (N23231, N23219, N13556, N4275);
nor NOR4 (N23232, N23229, N12576, N2447, N19594);
buf BUF1 (N23233, N23225);
and AND3 (N23234, N23218, N9472, N4910);
buf BUF1 (N23235, N23233);
and AND2 (N23236, N23232, N14808);
xor XOR2 (N23237, N23236, N10373);
and AND4 (N23238, N23204, N9383, N12204, N16447);
buf BUF1 (N23239, N23231);
not NOT1 (N23240, N23238);
or OR2 (N23241, N23230, N823);
xor XOR2 (N23242, N23240, N10137);
nor NOR4 (N23243, N23234, N14376, N1611, N2138);
and AND2 (N23244, N23221, N11982);
buf BUF1 (N23245, N23226);
buf BUF1 (N23246, N23244);
xor XOR2 (N23247, N23235, N8575);
nor NOR3 (N23248, N23217, N17348, N12674);
xor XOR2 (N23249, N23245, N7162);
buf BUF1 (N23250, N23248);
xor XOR2 (N23251, N23241, N22565);
or OR4 (N23252, N23251, N18676, N11178, N22905);
not NOT1 (N23253, N23249);
not NOT1 (N23254, N23243);
nand NAND4 (N23255, N23247, N11144, N4121, N4327);
buf BUF1 (N23256, N23252);
or OR3 (N23257, N23227, N19405, N6118);
xor XOR2 (N23258, N23237, N5295);
nor NOR2 (N23259, N23242, N15716);
nand NAND3 (N23260, N23239, N16808, N6023);
not NOT1 (N23261, N23250);
nand NAND4 (N23262, N23259, N21140, N14103, N5421);
buf BUF1 (N23263, N23246);
not NOT1 (N23264, N23258);
nand NAND4 (N23265, N23256, N289, N15641, N18735);
nor NOR2 (N23266, N23263, N17939);
buf BUF1 (N23267, N23264);
and AND4 (N23268, N23266, N12688, N18527, N14041);
xor XOR2 (N23269, N23257, N10291);
nor NOR4 (N23270, N23265, N653, N1271, N14454);
not NOT1 (N23271, N23267);
nand NAND3 (N23272, N23254, N9492, N19070);
nand NAND3 (N23273, N23269, N2103, N9740);
or OR3 (N23274, N23272, N10878, N21712);
not NOT1 (N23275, N23261);
nor NOR3 (N23276, N23255, N14722, N13921);
nor NOR3 (N23277, N23276, N22694, N20901);
buf BUF1 (N23278, N23260);
xor XOR2 (N23279, N23270, N6311);
nand NAND4 (N23280, N23273, N3319, N4614, N1938);
buf BUF1 (N23281, N23271);
buf BUF1 (N23282, N23253);
buf BUF1 (N23283, N23262);
buf BUF1 (N23284, N23281);
not NOT1 (N23285, N23282);
and AND2 (N23286, N23277, N9109);
xor XOR2 (N23287, N23275, N22755);
nor NOR2 (N23288, N23287, N1249);
buf BUF1 (N23289, N23286);
xor XOR2 (N23290, N23284, N11939);
buf BUF1 (N23291, N23283);
nor NOR4 (N23292, N23289, N20922, N21010, N15623);
not NOT1 (N23293, N23279);
buf BUF1 (N23294, N23288);
not NOT1 (N23295, N23292);
and AND4 (N23296, N23268, N22087, N14148, N6056);
nand NAND4 (N23297, N23280, N19509, N21448, N21252);
buf BUF1 (N23298, N23291);
or OR3 (N23299, N23290, N14379, N8059);
not NOT1 (N23300, N23294);
nand NAND2 (N23301, N23295, N5653);
nor NOR3 (N23302, N23293, N21623, N5646);
nor NOR4 (N23303, N23302, N13592, N8684, N10689);
nand NAND4 (N23304, N23297, N17901, N2489, N9343);
and AND4 (N23305, N23296, N20904, N21558, N1705);
nand NAND2 (N23306, N23278, N10427);
not NOT1 (N23307, N23301);
not NOT1 (N23308, N23300);
nor NOR2 (N23309, N23304, N1985);
buf BUF1 (N23310, N23306);
and AND3 (N23311, N23303, N1245, N4596);
and AND3 (N23312, N23285, N1236, N19438);
not NOT1 (N23313, N23274);
xor XOR2 (N23314, N23310, N13722);
not NOT1 (N23315, N23298);
xor XOR2 (N23316, N23311, N2001);
nor NOR4 (N23317, N23312, N13021, N7057, N6066);
or OR4 (N23318, N23313, N14700, N7704, N10791);
not NOT1 (N23319, N23308);
not NOT1 (N23320, N23305);
not NOT1 (N23321, N23307);
nand NAND3 (N23322, N23321, N10031, N8524);
nand NAND4 (N23323, N23320, N14729, N22641, N11657);
xor XOR2 (N23324, N23316, N22794);
or OR3 (N23325, N23314, N21836, N2929);
not NOT1 (N23326, N23299);
buf BUF1 (N23327, N23318);
not NOT1 (N23328, N23317);
and AND2 (N23329, N23315, N20923);
buf BUF1 (N23330, N23329);
and AND3 (N23331, N23319, N5431, N2243);
not NOT1 (N23332, N23323);
nor NOR3 (N23333, N23309, N1546, N21911);
not NOT1 (N23334, N23327);
nand NAND3 (N23335, N23325, N3495, N6354);
nand NAND3 (N23336, N23328, N15245, N5351);
xor XOR2 (N23337, N23322, N17815);
nand NAND4 (N23338, N23336, N9068, N18949, N14324);
xor XOR2 (N23339, N23331, N23251);
or OR3 (N23340, N23326, N20302, N22285);
nor NOR2 (N23341, N23338, N9960);
nor NOR4 (N23342, N23340, N4762, N3325, N1877);
not NOT1 (N23343, N23324);
and AND4 (N23344, N23337, N22769, N20619, N15127);
nand NAND3 (N23345, N23341, N21975, N16257);
nor NOR3 (N23346, N23330, N16010, N13272);
or OR3 (N23347, N23335, N14812, N18292);
buf BUF1 (N23348, N23339);
or OR4 (N23349, N23344, N14745, N20946, N14431);
not NOT1 (N23350, N23348);
not NOT1 (N23351, N23333);
xor XOR2 (N23352, N23342, N12311);
or OR2 (N23353, N23332, N16696);
nand NAND3 (N23354, N23352, N22816, N6768);
buf BUF1 (N23355, N23343);
xor XOR2 (N23356, N23345, N12058);
nand NAND3 (N23357, N23346, N8015, N12048);
buf BUF1 (N23358, N23355);
nor NOR2 (N23359, N23357, N21262);
nor NOR2 (N23360, N23347, N11736);
xor XOR2 (N23361, N23360, N18557);
buf BUF1 (N23362, N23351);
xor XOR2 (N23363, N23359, N5332);
not NOT1 (N23364, N23356);
buf BUF1 (N23365, N23349);
nand NAND4 (N23366, N23350, N4079, N2886, N934);
nand NAND3 (N23367, N23365, N17405, N6094);
nand NAND3 (N23368, N23354, N1585, N2327);
nor NOR2 (N23369, N23367, N16221);
xor XOR2 (N23370, N23366, N20155);
nand NAND3 (N23371, N23364, N12483, N4791);
nor NOR4 (N23372, N23353, N15971, N8347, N21492);
xor XOR2 (N23373, N23372, N8130);
and AND2 (N23374, N23368, N13419);
nand NAND2 (N23375, N23334, N16117);
not NOT1 (N23376, N23370);
nand NAND2 (N23377, N23376, N20938);
nor NOR2 (N23378, N23374, N826);
xor XOR2 (N23379, N23361, N22222);
and AND4 (N23380, N23362, N12398, N11339, N3774);
or OR4 (N23381, N23380, N12919, N19300, N9149);
and AND3 (N23382, N23377, N8522, N14062);
nand NAND2 (N23383, N23382, N4310);
or OR2 (N23384, N23371, N3924);
nand NAND2 (N23385, N23358, N18975);
nor NOR3 (N23386, N23373, N191, N18788);
nand NAND4 (N23387, N23383, N22165, N13022, N23122);
buf BUF1 (N23388, N23379);
nor NOR3 (N23389, N23363, N22824, N22280);
not NOT1 (N23390, N23385);
nand NAND2 (N23391, N23381, N16466);
nand NAND3 (N23392, N23390, N9894, N98);
buf BUF1 (N23393, N23384);
not NOT1 (N23394, N23388);
xor XOR2 (N23395, N23378, N17785);
not NOT1 (N23396, N23369);
or OR2 (N23397, N23391, N19266);
and AND2 (N23398, N23389, N11386);
or OR3 (N23399, N23398, N10805, N17192);
or OR2 (N23400, N23393, N900);
nand NAND4 (N23401, N23399, N19665, N20250, N6520);
nor NOR4 (N23402, N23392, N3395, N1629, N2680);
nor NOR4 (N23403, N23394, N4048, N6944, N22846);
nor NOR3 (N23404, N23396, N19892, N3257);
nand NAND3 (N23405, N23402, N275, N13832);
or OR3 (N23406, N23401, N13519, N13154);
nor NOR2 (N23407, N23404, N8479);
xor XOR2 (N23408, N23403, N21446);
or OR2 (N23409, N23397, N1710);
buf BUF1 (N23410, N23387);
nor NOR3 (N23411, N23375, N16956, N9678);
and AND3 (N23412, N23407, N14927, N4140);
nor NOR2 (N23413, N23411, N4757);
not NOT1 (N23414, N23412);
not NOT1 (N23415, N23413);
and AND2 (N23416, N23386, N10247);
nor NOR3 (N23417, N23406, N19900, N1391);
nand NAND3 (N23418, N23417, N19214, N21032);
and AND4 (N23419, N23410, N22914, N5861, N2658);
xor XOR2 (N23420, N23395, N9254);
nor NOR2 (N23421, N23420, N22965);
nand NAND4 (N23422, N23418, N6319, N22955, N17202);
or OR2 (N23423, N23408, N5681);
not NOT1 (N23424, N23422);
xor XOR2 (N23425, N23409, N23050);
or OR2 (N23426, N23425, N6949);
not NOT1 (N23427, N23416);
buf BUF1 (N23428, N23426);
xor XOR2 (N23429, N23400, N5343);
buf BUF1 (N23430, N23415);
nor NOR2 (N23431, N23424, N8744);
buf BUF1 (N23432, N23431);
buf BUF1 (N23433, N23432);
nand NAND2 (N23434, N23405, N7957);
or OR4 (N23435, N23421, N2805, N3082, N10331);
nand NAND4 (N23436, N23428, N20484, N9938, N1512);
xor XOR2 (N23437, N23419, N21475);
xor XOR2 (N23438, N23430, N5963);
nor NOR3 (N23439, N23437, N12201, N11854);
buf BUF1 (N23440, N23414);
nand NAND4 (N23441, N23436, N16679, N8379, N9225);
and AND2 (N23442, N23440, N15204);
nor NOR4 (N23443, N23439, N18109, N12873, N20943);
or OR4 (N23444, N23434, N3180, N21164, N7836);
nand NAND4 (N23445, N23433, N12093, N14675, N3154);
and AND3 (N23446, N23438, N16888, N22213);
not NOT1 (N23447, N23445);
xor XOR2 (N23448, N23444, N21060);
xor XOR2 (N23449, N23423, N10295);
buf BUF1 (N23450, N23427);
xor XOR2 (N23451, N23446, N11521);
xor XOR2 (N23452, N23450, N5182);
xor XOR2 (N23453, N23442, N7750);
xor XOR2 (N23454, N23453, N2312);
or OR2 (N23455, N23447, N14693);
nand NAND2 (N23456, N23451, N3682);
nor NOR4 (N23457, N23443, N22780, N21495, N10221);
xor XOR2 (N23458, N23456, N2655);
not NOT1 (N23459, N23452);
nand NAND2 (N23460, N23435, N7913);
and AND3 (N23461, N23448, N14985, N17228);
not NOT1 (N23462, N23449);
nor NOR2 (N23463, N23455, N20487);
buf BUF1 (N23464, N23441);
nor NOR4 (N23465, N23463, N21077, N3902, N55);
nor NOR4 (N23466, N23459, N15365, N23384, N13242);
xor XOR2 (N23467, N23465, N1809);
not NOT1 (N23468, N23462);
nand NAND2 (N23469, N23460, N11072);
not NOT1 (N23470, N23458);
nand NAND2 (N23471, N23454, N22054);
not NOT1 (N23472, N23467);
nor NOR4 (N23473, N23466, N3845, N12797, N18311);
not NOT1 (N23474, N23472);
xor XOR2 (N23475, N23457, N21175);
buf BUF1 (N23476, N23473);
xor XOR2 (N23477, N23476, N8012);
xor XOR2 (N23478, N23464, N7270);
not NOT1 (N23479, N23429);
and AND4 (N23480, N23469, N15940, N9220, N22855);
xor XOR2 (N23481, N23475, N3452);
and AND4 (N23482, N23481, N686, N13428, N3261);
xor XOR2 (N23483, N23479, N22296);
and AND4 (N23484, N23468, N12888, N13403, N16186);
not NOT1 (N23485, N23484);
or OR4 (N23486, N23485, N2367, N13275, N5767);
not NOT1 (N23487, N23480);
buf BUF1 (N23488, N23487);
nand NAND3 (N23489, N23477, N7805, N8536);
nand NAND2 (N23490, N23470, N18172);
xor XOR2 (N23491, N23488, N9558);
not NOT1 (N23492, N23478);
buf BUF1 (N23493, N23483);
nor NOR3 (N23494, N23486, N16090, N16031);
and AND3 (N23495, N23474, N14162, N2769);
not NOT1 (N23496, N23492);
nand NAND3 (N23497, N23495, N12191, N9349);
nor NOR2 (N23498, N23496, N18553);
nor NOR3 (N23499, N23494, N14765, N6496);
buf BUF1 (N23500, N23482);
buf BUF1 (N23501, N23489);
or OR2 (N23502, N23497, N11183);
nand NAND2 (N23503, N23461, N1393);
and AND2 (N23504, N23499, N22656);
buf BUF1 (N23505, N23501);
buf BUF1 (N23506, N23493);
and AND4 (N23507, N23503, N23128, N10946, N10087);
nand NAND4 (N23508, N23471, N22628, N10575, N9617);
nor NOR2 (N23509, N23507, N21503);
not NOT1 (N23510, N23509);
nor NOR2 (N23511, N23506, N1360);
or OR3 (N23512, N23502, N5798, N486);
buf BUF1 (N23513, N23490);
and AND2 (N23514, N23508, N935);
not NOT1 (N23515, N23498);
xor XOR2 (N23516, N23514, N8999);
or OR2 (N23517, N23491, N9941);
nor NOR3 (N23518, N23504, N17673, N6035);
nand NAND3 (N23519, N23513, N18714, N7706);
buf BUF1 (N23520, N23511);
xor XOR2 (N23521, N23520, N22519);
not NOT1 (N23522, N23512);
xor XOR2 (N23523, N23516, N22431);
or OR2 (N23524, N23523, N5050);
or OR2 (N23525, N23515, N4035);
buf BUF1 (N23526, N23518);
nor NOR2 (N23527, N23526, N22730);
buf BUF1 (N23528, N23505);
xor XOR2 (N23529, N23500, N14958);
not NOT1 (N23530, N23524);
nor NOR2 (N23531, N23521, N13371);
and AND2 (N23532, N23530, N963);
xor XOR2 (N23533, N23531, N6068);
not NOT1 (N23534, N23517);
buf BUF1 (N23535, N23534);
nand NAND2 (N23536, N23533, N1528);
or OR2 (N23537, N23528, N4550);
and AND4 (N23538, N23510, N12543, N615, N540);
xor XOR2 (N23539, N23538, N22798);
not NOT1 (N23540, N23536);
or OR4 (N23541, N23535, N11621, N18500, N17213);
nor NOR2 (N23542, N23541, N23374);
nor NOR2 (N23543, N23542, N17328);
or OR3 (N23544, N23525, N10634, N22560);
or OR3 (N23545, N23519, N23039, N8556);
buf BUF1 (N23546, N23539);
nand NAND2 (N23547, N23537, N5285);
nor NOR3 (N23548, N23547, N7617, N18037);
or OR4 (N23549, N23529, N4238, N4549, N6574);
nor NOR3 (N23550, N23532, N4712, N2161);
nor NOR3 (N23551, N23540, N4748, N1347);
and AND2 (N23552, N23546, N12374);
nor NOR4 (N23553, N23544, N23006, N3098, N1148);
nand NAND3 (N23554, N23550, N3050, N18236);
nand NAND2 (N23555, N23545, N14751);
nor NOR3 (N23556, N23549, N1622, N10116);
not NOT1 (N23557, N23556);
and AND4 (N23558, N23554, N17315, N22028, N19740);
and AND3 (N23559, N23553, N18889, N2246);
nand NAND3 (N23560, N23522, N16998, N16655);
not NOT1 (N23561, N23551);
buf BUF1 (N23562, N23561);
nand NAND4 (N23563, N23543, N4977, N19261, N9047);
nand NAND2 (N23564, N23559, N8608);
xor XOR2 (N23565, N23548, N16431);
xor XOR2 (N23566, N23562, N18139);
nor NOR4 (N23567, N23552, N14729, N18987, N2805);
or OR3 (N23568, N23558, N11915, N7113);
nand NAND3 (N23569, N23564, N20799, N21645);
nand NAND3 (N23570, N23563, N6000, N14143);
and AND3 (N23571, N23566, N3813, N22840);
buf BUF1 (N23572, N23570);
nor NOR2 (N23573, N23569, N5343);
buf BUF1 (N23574, N23560);
not NOT1 (N23575, N23527);
or OR2 (N23576, N23568, N3196);
buf BUF1 (N23577, N23557);
nor NOR3 (N23578, N23577, N18401, N2783);
xor XOR2 (N23579, N23578, N414);
xor XOR2 (N23580, N23579, N7267);
nor NOR4 (N23581, N23565, N18283, N7386, N11534);
nor NOR3 (N23582, N23574, N11044, N3636);
nor NOR2 (N23583, N23581, N6378);
nand NAND3 (N23584, N23555, N5045, N2752);
buf BUF1 (N23585, N23583);
and AND2 (N23586, N23573, N17651);
and AND3 (N23587, N23584, N9488, N22322);
nand NAND2 (N23588, N23572, N23517);
nand NAND3 (N23589, N23567, N20578, N21733);
or OR3 (N23590, N23580, N19886, N14714);
nor NOR3 (N23591, N23582, N16118, N3531);
nand NAND3 (N23592, N23575, N15479, N13420);
not NOT1 (N23593, N23571);
xor XOR2 (N23594, N23593, N13873);
not NOT1 (N23595, N23591);
nor NOR4 (N23596, N23587, N18820, N19320, N1549);
and AND2 (N23597, N23590, N400);
or OR3 (N23598, N23597, N15113, N13597);
nand NAND4 (N23599, N23598, N18945, N14386, N15734);
buf BUF1 (N23600, N23599);
and AND2 (N23601, N23594, N9734);
buf BUF1 (N23602, N23592);
nor NOR2 (N23603, N23585, N12871);
not NOT1 (N23604, N23596);
buf BUF1 (N23605, N23595);
and AND4 (N23606, N23604, N1706, N16755, N12669);
or OR4 (N23607, N23606, N17325, N4231, N18841);
nor NOR2 (N23608, N23605, N12171);
or OR2 (N23609, N23602, N13140);
xor XOR2 (N23610, N23601, N15090);
not NOT1 (N23611, N23610);
not NOT1 (N23612, N23576);
and AND2 (N23613, N23609, N19855);
or OR2 (N23614, N23612, N7447);
or OR2 (N23615, N23611, N9822);
nand NAND4 (N23616, N23603, N4633, N12811, N13035);
or OR2 (N23617, N23586, N2340);
not NOT1 (N23618, N23607);
and AND3 (N23619, N23615, N1529, N17588);
xor XOR2 (N23620, N23618, N21056);
and AND3 (N23621, N23617, N23607, N13057);
not NOT1 (N23622, N23613);
and AND4 (N23623, N23621, N13417, N23586, N15176);
or OR4 (N23624, N23623, N4232, N16984, N5733);
and AND4 (N23625, N23588, N4758, N14687, N18651);
buf BUF1 (N23626, N23614);
nand NAND2 (N23627, N23608, N5438);
not NOT1 (N23628, N23589);
not NOT1 (N23629, N23625);
or OR2 (N23630, N23619, N20397);
nor NOR2 (N23631, N23626, N3792);
not NOT1 (N23632, N23620);
nor NOR3 (N23633, N23631, N6790, N17261);
and AND4 (N23634, N23630, N1894, N3468, N11198);
xor XOR2 (N23635, N23600, N8117);
not NOT1 (N23636, N23627);
and AND3 (N23637, N23616, N19572, N16823);
and AND2 (N23638, N23632, N19928);
or OR2 (N23639, N23636, N506);
not NOT1 (N23640, N23635);
and AND3 (N23641, N23637, N20266, N19005);
not NOT1 (N23642, N23633);
not NOT1 (N23643, N23629);
xor XOR2 (N23644, N23628, N20734);
and AND2 (N23645, N23624, N8060);
buf BUF1 (N23646, N23622);
xor XOR2 (N23647, N23638, N23404);
buf BUF1 (N23648, N23647);
buf BUF1 (N23649, N23634);
xor XOR2 (N23650, N23639, N7043);
nor NOR3 (N23651, N23642, N7080, N12553);
or OR4 (N23652, N23643, N23355, N18302, N1607);
or OR4 (N23653, N23651, N18842, N16416, N16512);
not NOT1 (N23654, N23652);
and AND3 (N23655, N23641, N15814, N21851);
buf BUF1 (N23656, N23644);
and AND3 (N23657, N23646, N845, N11351);
nor NOR2 (N23658, N23653, N17066);
nand NAND3 (N23659, N23650, N21842, N8614);
not NOT1 (N23660, N23656);
or OR4 (N23661, N23654, N23098, N13692, N17723);
nand NAND4 (N23662, N23658, N11699, N609, N9393);
buf BUF1 (N23663, N23657);
not NOT1 (N23664, N23645);
nor NOR4 (N23665, N23640, N1019, N20618, N23491);
buf BUF1 (N23666, N23660);
not NOT1 (N23667, N23649);
or OR3 (N23668, N23664, N6365, N4398);
buf BUF1 (N23669, N23666);
buf BUF1 (N23670, N23661);
nor NOR3 (N23671, N23665, N16812, N22987);
xor XOR2 (N23672, N23648, N23405);
or OR4 (N23673, N23670, N13043, N2688, N6142);
not NOT1 (N23674, N23671);
nor NOR2 (N23675, N23662, N23365);
nor NOR2 (N23676, N23674, N9925);
or OR3 (N23677, N23655, N12540, N13266);
not NOT1 (N23678, N23669);
not NOT1 (N23679, N23675);
xor XOR2 (N23680, N23679, N16601);
or OR2 (N23681, N23667, N19849);
not NOT1 (N23682, N23680);
not NOT1 (N23683, N23673);
xor XOR2 (N23684, N23682, N22251);
or OR2 (N23685, N23659, N4302);
and AND2 (N23686, N23663, N15396);
nor NOR4 (N23687, N23678, N19334, N22268, N12599);
xor XOR2 (N23688, N23681, N1861);
or OR4 (N23689, N23672, N19709, N20356, N12771);
not NOT1 (N23690, N23685);
not NOT1 (N23691, N23690);
xor XOR2 (N23692, N23677, N14879);
xor XOR2 (N23693, N23687, N8502);
nor NOR2 (N23694, N23676, N21261);
nand NAND3 (N23695, N23683, N3634, N20902);
xor XOR2 (N23696, N23688, N11465);
not NOT1 (N23697, N23689);
not NOT1 (N23698, N23696);
or OR3 (N23699, N23692, N23658, N18311);
or OR4 (N23700, N23684, N11043, N17720, N20630);
xor XOR2 (N23701, N23693, N3465);
nor NOR4 (N23702, N23694, N8070, N14053, N7432);
xor XOR2 (N23703, N23686, N20312);
buf BUF1 (N23704, N23668);
buf BUF1 (N23705, N23704);
nor NOR3 (N23706, N23699, N22629, N10915);
or OR4 (N23707, N23706, N5713, N1728, N4020);
nand NAND2 (N23708, N23702, N14143);
and AND3 (N23709, N23695, N11423, N4743);
or OR3 (N23710, N23703, N1642, N21769);
nor NOR3 (N23711, N23691, N22124, N21236);
and AND4 (N23712, N23701, N23295, N7714, N6837);
buf BUF1 (N23713, N23700);
and AND4 (N23714, N23711, N6059, N11335, N21589);
xor XOR2 (N23715, N23713, N5678);
or OR3 (N23716, N23708, N21322, N6984);
nor NOR2 (N23717, N23716, N13445);
nor NOR3 (N23718, N23697, N16318, N18823);
xor XOR2 (N23719, N23709, N2155);
buf BUF1 (N23720, N23714);
xor XOR2 (N23721, N23707, N17235);
buf BUF1 (N23722, N23712);
buf BUF1 (N23723, N23721);
or OR3 (N23724, N23715, N12809, N12032);
and AND4 (N23725, N23718, N21801, N21955, N15774);
or OR3 (N23726, N23724, N11039, N11336);
or OR3 (N23727, N23726, N8467, N3653);
nor NOR3 (N23728, N23705, N17330, N1994);
nand NAND3 (N23729, N23727, N17957, N20295);
not NOT1 (N23730, N23723);
or OR2 (N23731, N23725, N13661);
nand NAND4 (N23732, N23730, N15904, N9359, N22349);
and AND3 (N23733, N23729, N4938, N21760);
nand NAND2 (N23734, N23720, N11546);
buf BUF1 (N23735, N23733);
and AND2 (N23736, N23710, N2228);
not NOT1 (N23737, N23731);
and AND3 (N23738, N23728, N1857, N18001);
nor NOR4 (N23739, N23698, N14190, N840, N7236);
nor NOR2 (N23740, N23719, N4733);
or OR3 (N23741, N23732, N8118, N19452);
buf BUF1 (N23742, N23737);
or OR2 (N23743, N23735, N22379);
buf BUF1 (N23744, N23722);
and AND3 (N23745, N23741, N9898, N16248);
nor NOR3 (N23746, N23739, N10454, N4926);
buf BUF1 (N23747, N23738);
nand NAND3 (N23748, N23746, N9047, N220);
buf BUF1 (N23749, N23742);
buf BUF1 (N23750, N23740);
nand NAND4 (N23751, N23736, N3182, N16554, N16361);
nand NAND2 (N23752, N23743, N6065);
nor NOR3 (N23753, N23748, N13891, N18178);
buf BUF1 (N23754, N23751);
or OR4 (N23755, N23749, N23403, N5381, N7057);
nor NOR3 (N23756, N23753, N12332, N23058);
nand NAND4 (N23757, N23744, N13737, N11893, N6454);
nand NAND3 (N23758, N23750, N11987, N6708);
xor XOR2 (N23759, N23752, N20873);
buf BUF1 (N23760, N23747);
and AND2 (N23761, N23758, N3932);
nor NOR2 (N23762, N23759, N6204);
xor XOR2 (N23763, N23761, N1712);
nor NOR4 (N23764, N23754, N21367, N18606, N1587);
nor NOR4 (N23765, N23756, N22693, N15310, N15702);
not NOT1 (N23766, N23755);
nand NAND2 (N23767, N23734, N13822);
and AND2 (N23768, N23764, N3178);
buf BUF1 (N23769, N23757);
xor XOR2 (N23770, N23763, N23323);
buf BUF1 (N23771, N23760);
xor XOR2 (N23772, N23762, N6751);
nand NAND3 (N23773, N23772, N7431, N20206);
and AND2 (N23774, N23745, N16065);
or OR4 (N23775, N23768, N8605, N21915, N22176);
nor NOR3 (N23776, N23771, N22565, N4686);
not NOT1 (N23777, N23770);
and AND4 (N23778, N23774, N23174, N265, N20623);
and AND4 (N23779, N23778, N13582, N11517, N272);
buf BUF1 (N23780, N23776);
nor NOR4 (N23781, N23765, N7273, N15564, N17864);
buf BUF1 (N23782, N23780);
or OR4 (N23783, N23777, N9394, N19811, N5406);
and AND2 (N23784, N23766, N18134);
buf BUF1 (N23785, N23767);
buf BUF1 (N23786, N23783);
not NOT1 (N23787, N23781);
or OR4 (N23788, N23769, N18116, N17049, N10854);
buf BUF1 (N23789, N23773);
and AND2 (N23790, N23786, N11358);
buf BUF1 (N23791, N23787);
nor NOR2 (N23792, N23784, N15290);
xor XOR2 (N23793, N23792, N13326);
or OR2 (N23794, N23790, N5627);
not NOT1 (N23795, N23785);
buf BUF1 (N23796, N23789);
nor NOR4 (N23797, N23796, N16151, N1650, N3390);
and AND4 (N23798, N23788, N22374, N15316, N5504);
xor XOR2 (N23799, N23717, N204);
xor XOR2 (N23800, N23794, N16389);
nand NAND4 (N23801, N23798, N20250, N3287, N13990);
nor NOR2 (N23802, N23779, N21865);
buf BUF1 (N23803, N23775);
or OR4 (N23804, N23802, N7738, N13748, N1914);
nand NAND3 (N23805, N23799, N17414, N8176);
xor XOR2 (N23806, N23793, N6680);
nor NOR4 (N23807, N23801, N17278, N5991, N14365);
or OR3 (N23808, N23804, N17366, N2374);
and AND3 (N23809, N23800, N17961, N1552);
not NOT1 (N23810, N23807);
nor NOR4 (N23811, N23810, N9608, N1232, N15843);
buf BUF1 (N23812, N23808);
buf BUF1 (N23813, N23791);
nor NOR3 (N23814, N23803, N5199, N11199);
buf BUF1 (N23815, N23814);
buf BUF1 (N23816, N23795);
not NOT1 (N23817, N23813);
or OR4 (N23818, N23806, N22150, N4935, N18297);
nor NOR3 (N23819, N23817, N11718, N6760);
and AND4 (N23820, N23805, N9232, N17467, N15673);
buf BUF1 (N23821, N23819);
and AND3 (N23822, N23811, N15486, N3823);
nor NOR3 (N23823, N23822, N4397, N23075);
buf BUF1 (N23824, N23820);
nand NAND2 (N23825, N23824, N6731);
or OR3 (N23826, N23815, N1964, N393);
nor NOR4 (N23827, N23797, N5857, N9683, N16791);
or OR4 (N23828, N23825, N15631, N8751, N19038);
or OR4 (N23829, N23826, N5594, N9405, N15293);
xor XOR2 (N23830, N23828, N19646);
nor NOR2 (N23831, N23782, N5413);
buf BUF1 (N23832, N23809);
nor NOR3 (N23833, N23823, N11826, N20148);
and AND3 (N23834, N23818, N19818, N11284);
nor NOR2 (N23835, N23829, N4670);
nor NOR4 (N23836, N23821, N5488, N11871, N11662);
xor XOR2 (N23837, N23835, N502);
nor NOR2 (N23838, N23816, N11209);
and AND4 (N23839, N23827, N10386, N19574, N4653);
nor NOR2 (N23840, N23830, N8266);
or OR4 (N23841, N23833, N7433, N2665, N9357);
buf BUF1 (N23842, N23840);
or OR3 (N23843, N23831, N12733, N15301);
nor NOR2 (N23844, N23841, N594);
and AND3 (N23845, N23842, N7648, N13569);
or OR2 (N23846, N23832, N23048);
buf BUF1 (N23847, N23843);
nand NAND2 (N23848, N23837, N12846);
and AND3 (N23849, N23812, N15637, N5774);
nand NAND3 (N23850, N23847, N7937, N8610);
xor XOR2 (N23851, N23846, N23329);
xor XOR2 (N23852, N23839, N5727);
nor NOR4 (N23853, N23848, N8051, N16185, N18458);
nand NAND4 (N23854, N23852, N10688, N761, N4555);
or OR3 (N23855, N23836, N23259, N3126);
xor XOR2 (N23856, N23845, N18298);
not NOT1 (N23857, N23853);
not NOT1 (N23858, N23851);
nor NOR3 (N23859, N23834, N5772, N12805);
or OR2 (N23860, N23857, N23557);
buf BUF1 (N23861, N23838);
nor NOR2 (N23862, N23860, N4989);
and AND3 (N23863, N23855, N6288, N4722);
xor XOR2 (N23864, N23861, N14033);
and AND4 (N23865, N23844, N10525, N17563, N12100);
and AND3 (N23866, N23859, N463, N17976);
nor NOR4 (N23867, N23865, N12121, N3656, N5368);
not NOT1 (N23868, N23858);
nand NAND3 (N23869, N23864, N6556, N15464);
nor NOR3 (N23870, N23854, N14387, N16891);
xor XOR2 (N23871, N23869, N17399);
and AND4 (N23872, N23870, N9255, N17614, N19265);
buf BUF1 (N23873, N23871);
buf BUF1 (N23874, N23872);
or OR2 (N23875, N23866, N12780);
or OR2 (N23876, N23856, N9385);
nor NOR2 (N23877, N23867, N5460);
not NOT1 (N23878, N23876);
and AND3 (N23879, N23878, N8625, N13533);
nand NAND2 (N23880, N23873, N4935);
buf BUF1 (N23881, N23879);
nor NOR3 (N23882, N23875, N17086, N4145);
or OR4 (N23883, N23863, N18963, N88, N20578);
or OR4 (N23884, N23881, N13249, N1731, N19976);
xor XOR2 (N23885, N23868, N13990);
nor NOR3 (N23886, N23885, N19057, N7169);
buf BUF1 (N23887, N23877);
xor XOR2 (N23888, N23880, N18528);
xor XOR2 (N23889, N23887, N10117);
or OR3 (N23890, N23886, N11367, N8793);
or OR4 (N23891, N23882, N7904, N5672, N19403);
and AND2 (N23892, N23884, N14725);
nand NAND4 (N23893, N23889, N1423, N848, N15458);
nor NOR2 (N23894, N23892, N13235);
xor XOR2 (N23895, N23849, N5489);
nand NAND4 (N23896, N23895, N21186, N2036, N20507);
and AND3 (N23897, N23883, N9735, N11504);
not NOT1 (N23898, N23874);
and AND4 (N23899, N23862, N21287, N23796, N23535);
not NOT1 (N23900, N23893);
nand NAND2 (N23901, N23891, N17488);
nand NAND4 (N23902, N23890, N12716, N21288, N12096);
or OR2 (N23903, N23888, N2137);
not NOT1 (N23904, N23901);
nand NAND2 (N23905, N23894, N13135);
nand NAND3 (N23906, N23899, N4923, N13237);
not NOT1 (N23907, N23903);
nand NAND3 (N23908, N23850, N22133, N2329);
not NOT1 (N23909, N23902);
or OR3 (N23910, N23908, N15817, N11783);
and AND4 (N23911, N23907, N9100, N2541, N11496);
buf BUF1 (N23912, N23904);
nor NOR4 (N23913, N23906, N8549, N15547, N19468);
and AND2 (N23914, N23912, N2291);
nand NAND2 (N23915, N23897, N12091);
buf BUF1 (N23916, N23905);
xor XOR2 (N23917, N23915, N3168);
xor XOR2 (N23918, N23911, N12798);
and AND2 (N23919, N23916, N17038);
nor NOR3 (N23920, N23909, N18400, N21558);
and AND2 (N23921, N23920, N846);
and AND3 (N23922, N23896, N22316, N10192);
buf BUF1 (N23923, N23914);
and AND4 (N23924, N23921, N7404, N23439, N21536);
nor NOR4 (N23925, N23913, N14545, N2926, N14694);
xor XOR2 (N23926, N23918, N13470);
xor XOR2 (N23927, N23924, N8804);
and AND2 (N23928, N23917, N18264);
and AND2 (N23929, N23928, N4563);
not NOT1 (N23930, N23929);
buf BUF1 (N23931, N23910);
nand NAND3 (N23932, N23898, N1746, N22912);
or OR4 (N23933, N23925, N16471, N23562, N846);
or OR2 (N23934, N23922, N10431);
not NOT1 (N23935, N23932);
xor XOR2 (N23936, N23927, N17937);
buf BUF1 (N23937, N23935);
not NOT1 (N23938, N23934);
xor XOR2 (N23939, N23936, N556);
nand NAND4 (N23940, N23937, N16996, N1047, N20288);
not NOT1 (N23941, N23940);
and AND4 (N23942, N23931, N3410, N2889, N320);
and AND2 (N23943, N23941, N8504);
not NOT1 (N23944, N23942);
and AND2 (N23945, N23944, N22504);
nor NOR2 (N23946, N23938, N11695);
nor NOR3 (N23947, N23943, N10758, N7899);
and AND2 (N23948, N23946, N3281);
xor XOR2 (N23949, N23945, N11905);
nor NOR3 (N23950, N23900, N19356, N17556);
buf BUF1 (N23951, N23926);
xor XOR2 (N23952, N23933, N21602);
and AND3 (N23953, N23923, N10703, N20702);
nor NOR4 (N23954, N23952, N891, N21561, N6119);
nand NAND2 (N23955, N23948, N3265);
not NOT1 (N23956, N23953);
xor XOR2 (N23957, N23919, N5170);
buf BUF1 (N23958, N23947);
not NOT1 (N23959, N23956);
or OR3 (N23960, N23950, N9700, N6283);
or OR3 (N23961, N23951, N10586, N5320);
buf BUF1 (N23962, N23930);
buf BUF1 (N23963, N23954);
and AND4 (N23964, N23961, N2049, N20068, N269);
nand NAND3 (N23965, N23959, N19602, N20825);
xor XOR2 (N23966, N23962, N15408);
nor NOR2 (N23967, N23966, N23495);
buf BUF1 (N23968, N23967);
and AND3 (N23969, N23964, N5990, N2192);
nand NAND2 (N23970, N23968, N22827);
not NOT1 (N23971, N23970);
nand NAND4 (N23972, N23965, N3008, N14291, N1940);
buf BUF1 (N23973, N23957);
not NOT1 (N23974, N23960);
nor NOR4 (N23975, N23972, N12912, N16855, N10490);
xor XOR2 (N23976, N23973, N18500);
and AND4 (N23977, N23974, N18078, N17731, N12815);
and AND2 (N23978, N23963, N8972);
nor NOR4 (N23979, N23976, N9059, N23345, N18058);
buf BUF1 (N23980, N23958);
nor NOR4 (N23981, N23971, N23291, N12420, N17376);
buf BUF1 (N23982, N23955);
or OR2 (N23983, N23969, N23653);
and AND4 (N23984, N23980, N1295, N16852, N19127);
nand NAND4 (N23985, N23982, N16063, N13354, N17407);
not NOT1 (N23986, N23984);
xor XOR2 (N23987, N23975, N13904);
xor XOR2 (N23988, N23983, N5816);
or OR4 (N23989, N23987, N16235, N2010, N17870);
nand NAND3 (N23990, N23949, N6878, N6093);
nand NAND2 (N23991, N23979, N5398);
nand NAND4 (N23992, N23990, N9945, N11116, N19658);
and AND3 (N23993, N23977, N20215, N7913);
not NOT1 (N23994, N23981);
not NOT1 (N23995, N23939);
nand NAND4 (N23996, N23986, N11720, N23305, N10895);
not NOT1 (N23997, N23995);
xor XOR2 (N23998, N23993, N17933);
or OR2 (N23999, N23991, N15799);
xor XOR2 (N24000, N23994, N6338);
xor XOR2 (N24001, N23999, N13686);
buf BUF1 (N24002, N23978);
nand NAND4 (N24003, N23998, N14864, N22110, N6073);
and AND2 (N24004, N24002, N19971);
buf BUF1 (N24005, N24004);
and AND4 (N24006, N23992, N14183, N18232, N10599);
nand NAND2 (N24007, N24003, N7416);
or OR2 (N24008, N24001, N16899);
and AND2 (N24009, N23989, N13932);
or OR2 (N24010, N23985, N1257);
or OR4 (N24011, N24009, N3023, N9277, N14457);
or OR2 (N24012, N24000, N7518);
or OR3 (N24013, N24005, N10976, N13127);
xor XOR2 (N24014, N23996, N6637);
and AND3 (N24015, N24006, N4676, N519);
or OR4 (N24016, N24008, N1189, N10809, N23396);
nor NOR3 (N24017, N23988, N4152, N12571);
and AND2 (N24018, N24010, N14187);
xor XOR2 (N24019, N24017, N12999);
and AND3 (N24020, N23997, N1320, N106);
and AND2 (N24021, N24014, N23254);
buf BUF1 (N24022, N24018);
xor XOR2 (N24023, N24007, N4364);
buf BUF1 (N24024, N24015);
nor NOR3 (N24025, N24024, N4810, N6306);
nand NAND4 (N24026, N24023, N10960, N10852, N16029);
nor NOR4 (N24027, N24019, N11810, N12026, N9840);
and AND4 (N24028, N24016, N21411, N1588, N3922);
buf BUF1 (N24029, N24021);
nor NOR2 (N24030, N24013, N20071);
not NOT1 (N24031, N24025);
xor XOR2 (N24032, N24012, N609);
buf BUF1 (N24033, N24031);
or OR3 (N24034, N24029, N5466, N23971);
or OR2 (N24035, N24032, N2549);
nor NOR4 (N24036, N24028, N12533, N16623, N8612);
and AND2 (N24037, N24027, N11169);
nand NAND2 (N24038, N24036, N13864);
xor XOR2 (N24039, N24020, N2396);
and AND4 (N24040, N24011, N7389, N2892, N14039);
buf BUF1 (N24041, N24026);
nand NAND2 (N24042, N24038, N2784);
not NOT1 (N24043, N24035);
buf BUF1 (N24044, N24042);
buf BUF1 (N24045, N24030);
or OR4 (N24046, N24034, N15907, N7541, N12569);
buf BUF1 (N24047, N24039);
buf BUF1 (N24048, N24037);
and AND3 (N24049, N24046, N9165, N6563);
buf BUF1 (N24050, N24022);
and AND4 (N24051, N24049, N18243, N5847, N2613);
buf BUF1 (N24052, N24043);
or OR4 (N24053, N24050, N22930, N12939, N18469);
nor NOR4 (N24054, N24053, N11608, N1534, N22065);
nor NOR4 (N24055, N24041, N9506, N16599, N6518);
xor XOR2 (N24056, N24033, N2489);
nand NAND3 (N24057, N24056, N11596, N12758);
buf BUF1 (N24058, N24047);
and AND4 (N24059, N24054, N4638, N15411, N8331);
nor NOR2 (N24060, N24040, N14777);
not NOT1 (N24061, N24057);
nor NOR3 (N24062, N24060, N9851, N8988);
and AND4 (N24063, N24058, N12961, N409, N6696);
not NOT1 (N24064, N24048);
buf BUF1 (N24065, N24051);
not NOT1 (N24066, N24065);
or OR4 (N24067, N24044, N16203, N139, N6391);
nand NAND2 (N24068, N24067, N12413);
not NOT1 (N24069, N24052);
xor XOR2 (N24070, N24045, N12039);
and AND2 (N24071, N24055, N8195);
xor XOR2 (N24072, N24069, N16713);
or OR2 (N24073, N24061, N7842);
nand NAND2 (N24074, N24064, N654);
or OR4 (N24075, N24071, N17082, N1571, N16032);
buf BUF1 (N24076, N24068);
and AND2 (N24077, N24074, N13297);
buf BUF1 (N24078, N24073);
nor NOR2 (N24079, N24078, N16452);
nand NAND3 (N24080, N24062, N17744, N21365);
nor NOR4 (N24081, N24066, N5101, N1647, N20710);
and AND4 (N24082, N24075, N716, N23334, N2921);
nand NAND3 (N24083, N24076, N9710, N9675);
nand NAND4 (N24084, N24079, N14936, N13152, N11951);
nand NAND2 (N24085, N24063, N23407);
nand NAND2 (N24086, N24084, N10608);
nand NAND2 (N24087, N24081, N8064);
nor NOR4 (N24088, N24070, N3564, N17783, N14067);
xor XOR2 (N24089, N24077, N12851);
nand NAND2 (N24090, N24083, N2532);
and AND2 (N24091, N24085, N11778);
nand NAND3 (N24092, N24059, N23965, N112);
buf BUF1 (N24093, N24092);
nand NAND3 (N24094, N24080, N15739, N2463);
or OR4 (N24095, N24087, N12525, N22440, N8461);
buf BUF1 (N24096, N24091);
or OR2 (N24097, N24089, N3223);
and AND4 (N24098, N24072, N21514, N4658, N3579);
xor XOR2 (N24099, N24090, N15315);
buf BUF1 (N24100, N24096);
and AND3 (N24101, N24095, N4212, N2465);
or OR2 (N24102, N24094, N13912);
buf BUF1 (N24103, N24093);
nand NAND4 (N24104, N24086, N19373, N22274, N11420);
xor XOR2 (N24105, N24082, N11160);
and AND2 (N24106, N24102, N21418);
not NOT1 (N24107, N24097);
or OR3 (N24108, N24101, N14768, N16652);
buf BUF1 (N24109, N24099);
or OR3 (N24110, N24107, N3518, N4098);
xor XOR2 (N24111, N24109, N21692);
nand NAND3 (N24112, N24088, N23824, N6090);
buf BUF1 (N24113, N24111);
nor NOR4 (N24114, N24108, N7082, N7319, N7822);
xor XOR2 (N24115, N24112, N19353);
not NOT1 (N24116, N24110);
and AND4 (N24117, N24104, N19342, N999, N4202);
buf BUF1 (N24118, N24115);
xor XOR2 (N24119, N24106, N10810);
or OR3 (N24120, N24098, N23449, N6143);
buf BUF1 (N24121, N24100);
or OR3 (N24122, N24113, N10213, N23136);
nand NAND4 (N24123, N24118, N5786, N11001, N2579);
or OR3 (N24124, N24123, N15108, N9307);
nand NAND2 (N24125, N24117, N1041);
xor XOR2 (N24126, N24103, N17389);
or OR2 (N24127, N24114, N8290);
or OR3 (N24128, N24127, N10547, N2415);
buf BUF1 (N24129, N24116);
not NOT1 (N24130, N24125);
xor XOR2 (N24131, N24105, N21298);
nand NAND2 (N24132, N24128, N10967);
not NOT1 (N24133, N24124);
not NOT1 (N24134, N24133);
nor NOR2 (N24135, N24126, N831);
not NOT1 (N24136, N24121);
or OR3 (N24137, N24129, N22025, N22702);
and AND4 (N24138, N24132, N21704, N7339, N20238);
nand NAND4 (N24139, N24137, N16714, N3171, N14809);
buf BUF1 (N24140, N24134);
nor NOR2 (N24141, N24138, N895);
not NOT1 (N24142, N24130);
not NOT1 (N24143, N24122);
not NOT1 (N24144, N24131);
buf BUF1 (N24145, N24143);
not NOT1 (N24146, N24120);
nand NAND2 (N24147, N24119, N3449);
nor NOR3 (N24148, N24140, N8985, N11376);
xor XOR2 (N24149, N24135, N20455);
xor XOR2 (N24150, N24146, N10477);
buf BUF1 (N24151, N24144);
xor XOR2 (N24152, N24141, N2064);
nand NAND4 (N24153, N24139, N16507, N6476, N10281);
and AND2 (N24154, N24147, N3294);
and AND4 (N24155, N24136, N2591, N23628, N14144);
buf BUF1 (N24156, N24153);
and AND2 (N24157, N24151, N19434);
not NOT1 (N24158, N24148);
buf BUF1 (N24159, N24150);
not NOT1 (N24160, N24155);
xor XOR2 (N24161, N24157, N4405);
nor NOR4 (N24162, N24158, N12858, N16082, N8565);
or OR4 (N24163, N24154, N16629, N15360, N23664);
buf BUF1 (N24164, N24152);
or OR3 (N24165, N24145, N14400, N13084);
or OR3 (N24166, N24156, N21167, N22771);
xor XOR2 (N24167, N24149, N12550);
xor XOR2 (N24168, N24164, N16161);
nand NAND4 (N24169, N24167, N9035, N10454, N21856);
not NOT1 (N24170, N24162);
nor NOR3 (N24171, N24169, N13148, N9584);
buf BUF1 (N24172, N24166);
nand NAND4 (N24173, N24170, N1797, N6097, N718);
xor XOR2 (N24174, N24142, N14278);
nor NOR3 (N24175, N24159, N6718, N3920);
buf BUF1 (N24176, N24168);
buf BUF1 (N24177, N24160);
nand NAND2 (N24178, N24165, N10402);
and AND3 (N24179, N24176, N20559, N11931);
nor NOR4 (N24180, N24178, N8640, N252, N20757);
or OR2 (N24181, N24177, N23893);
nand NAND2 (N24182, N24175, N23318);
nand NAND2 (N24183, N24179, N22831);
buf BUF1 (N24184, N24163);
xor XOR2 (N24185, N24183, N16484);
not NOT1 (N24186, N24182);
not NOT1 (N24187, N24180);
buf BUF1 (N24188, N24185);
xor XOR2 (N24189, N24186, N8010);
buf BUF1 (N24190, N24184);
buf BUF1 (N24191, N24181);
not NOT1 (N24192, N24173);
nor NOR3 (N24193, N24189, N1847, N18356);
and AND2 (N24194, N24193, N7707);
nand NAND2 (N24195, N24172, N12677);
nor NOR4 (N24196, N24161, N8788, N6800, N4376);
buf BUF1 (N24197, N24195);
xor XOR2 (N24198, N24192, N12839);
nor NOR2 (N24199, N24174, N13920);
buf BUF1 (N24200, N24187);
not NOT1 (N24201, N24198);
nand NAND3 (N24202, N24196, N15308, N14948);
nand NAND2 (N24203, N24171, N860);
nor NOR4 (N24204, N24202, N17342, N3712, N14656);
or OR2 (N24205, N24201, N6964);
buf BUF1 (N24206, N24190);
nor NOR2 (N24207, N24194, N9384);
not NOT1 (N24208, N24207);
buf BUF1 (N24209, N24197);
not NOT1 (N24210, N24191);
xor XOR2 (N24211, N24188, N8895);
buf BUF1 (N24212, N24206);
buf BUF1 (N24213, N24203);
and AND3 (N24214, N24204, N21898, N24141);
buf BUF1 (N24215, N24210);
buf BUF1 (N24216, N24209);
buf BUF1 (N24217, N24212);
and AND2 (N24218, N24215, N17269);
or OR2 (N24219, N24211, N7538);
not NOT1 (N24220, N24205);
and AND4 (N24221, N24208, N15510, N10791, N20477);
nand NAND3 (N24222, N24221, N9789, N17818);
not NOT1 (N24223, N24199);
and AND4 (N24224, N24213, N9746, N16349, N335);
nor NOR2 (N24225, N24222, N7272);
xor XOR2 (N24226, N24200, N15690);
nor NOR4 (N24227, N24214, N814, N10154, N14850);
xor XOR2 (N24228, N24226, N10600);
nand NAND4 (N24229, N24228, N2903, N20890, N9197);
not NOT1 (N24230, N24220);
buf BUF1 (N24231, N24227);
buf BUF1 (N24232, N24218);
and AND2 (N24233, N24230, N12230);
not NOT1 (N24234, N24233);
and AND3 (N24235, N24219, N3645, N18851);
or OR3 (N24236, N24234, N10137, N15861);
not NOT1 (N24237, N24231);
buf BUF1 (N24238, N24217);
not NOT1 (N24239, N24224);
not NOT1 (N24240, N24216);
not NOT1 (N24241, N24238);
nand NAND3 (N24242, N24235, N5199, N6177);
xor XOR2 (N24243, N24223, N10185);
nand NAND4 (N24244, N24243, N9569, N2862, N16616);
nand NAND3 (N24245, N24244, N1511, N11027);
or OR3 (N24246, N24232, N10590, N17732);
xor XOR2 (N24247, N24240, N10423);
not NOT1 (N24248, N24237);
buf BUF1 (N24249, N24242);
xor XOR2 (N24250, N24239, N991);
and AND4 (N24251, N24248, N21705, N373, N5153);
buf BUF1 (N24252, N24241);
buf BUF1 (N24253, N24250);
buf BUF1 (N24254, N24246);
nand NAND3 (N24255, N24252, N6943, N7669);
nand NAND2 (N24256, N24225, N23936);
xor XOR2 (N24257, N24245, N18863);
nand NAND2 (N24258, N24247, N9744);
xor XOR2 (N24259, N24236, N20534);
not NOT1 (N24260, N24257);
or OR2 (N24261, N24229, N8623);
not NOT1 (N24262, N24261);
nand NAND2 (N24263, N24260, N11222);
buf BUF1 (N24264, N24258);
not NOT1 (N24265, N24256);
nor NOR3 (N24266, N24255, N3737, N4598);
and AND4 (N24267, N24266, N19578, N20840, N10807);
nand NAND4 (N24268, N24249, N6378, N24075, N9766);
xor XOR2 (N24269, N24259, N12134);
or OR4 (N24270, N24269, N6749, N11893, N20371);
nand NAND2 (N24271, N24251, N10697);
not NOT1 (N24272, N24263);
or OR4 (N24273, N24253, N7081, N3357, N87);
nand NAND3 (N24274, N24262, N11211, N23052);
not NOT1 (N24275, N24268);
and AND4 (N24276, N24270, N10002, N11544, N21767);
buf BUF1 (N24277, N24274);
xor XOR2 (N24278, N24267, N22128);
xor XOR2 (N24279, N24275, N21808);
and AND4 (N24280, N24264, N6909, N14385, N14938);
buf BUF1 (N24281, N24278);
or OR3 (N24282, N24279, N1608, N22621);
or OR4 (N24283, N24277, N12865, N13357, N13764);
xor XOR2 (N24284, N24282, N16490);
or OR3 (N24285, N24273, N5739, N17009);
xor XOR2 (N24286, N24280, N17690);
and AND4 (N24287, N24283, N2719, N16462, N5574);
and AND4 (N24288, N24271, N22033, N7598, N7587);
nand NAND2 (N24289, N24265, N13140);
or OR3 (N24290, N24287, N9896, N4632);
not NOT1 (N24291, N24281);
or OR2 (N24292, N24289, N9215);
xor XOR2 (N24293, N24284, N4043);
not NOT1 (N24294, N24293);
nand NAND2 (N24295, N24294, N20626);
xor XOR2 (N24296, N24272, N18386);
not NOT1 (N24297, N24296);
buf BUF1 (N24298, N24288);
and AND3 (N24299, N24285, N141, N10856);
xor XOR2 (N24300, N24286, N10891);
xor XOR2 (N24301, N24254, N9025);
not NOT1 (N24302, N24299);
nor NOR3 (N24303, N24276, N24093, N3008);
nand NAND4 (N24304, N24290, N15265, N3788, N13981);
nand NAND3 (N24305, N24304, N5352, N15438);
nand NAND3 (N24306, N24292, N15824, N14582);
buf BUF1 (N24307, N24295);
buf BUF1 (N24308, N24307);
xor XOR2 (N24309, N24308, N12021);
buf BUF1 (N24310, N24302);
buf BUF1 (N24311, N24306);
nand NAND3 (N24312, N24310, N11323, N17775);
nor NOR3 (N24313, N24303, N21590, N22598);
or OR2 (N24314, N24301, N21101);
not NOT1 (N24315, N24291);
xor XOR2 (N24316, N24313, N5782);
nand NAND4 (N24317, N24315, N18791, N23804, N22736);
buf BUF1 (N24318, N24317);
and AND4 (N24319, N24312, N19252, N9971, N10417);
xor XOR2 (N24320, N24297, N381);
xor XOR2 (N24321, N24316, N22316);
or OR2 (N24322, N24311, N21543);
xor XOR2 (N24323, N24322, N15024);
xor XOR2 (N24324, N24319, N11398);
nand NAND4 (N24325, N24320, N18413, N19529, N659);
not NOT1 (N24326, N24318);
or OR4 (N24327, N24321, N19622, N18674, N8532);
not NOT1 (N24328, N24324);
and AND3 (N24329, N24326, N19005, N4778);
xor XOR2 (N24330, N24298, N14432);
or OR3 (N24331, N24328, N10447, N6465);
nand NAND2 (N24332, N24323, N22801);
buf BUF1 (N24333, N24329);
xor XOR2 (N24334, N24331, N17555);
and AND3 (N24335, N24305, N9107, N11904);
nor NOR2 (N24336, N24332, N24044);
nand NAND3 (N24337, N24335, N4673, N12594);
buf BUF1 (N24338, N24309);
or OR2 (N24339, N24327, N4421);
or OR2 (N24340, N24336, N14454);
xor XOR2 (N24341, N24333, N22878);
buf BUF1 (N24342, N24339);
xor XOR2 (N24343, N24341, N13708);
and AND2 (N24344, N24337, N10591);
buf BUF1 (N24345, N24325);
and AND2 (N24346, N24340, N5392);
nand NAND3 (N24347, N24338, N12135, N971);
xor XOR2 (N24348, N24300, N17957);
buf BUF1 (N24349, N24330);
and AND2 (N24350, N24345, N6114);
or OR4 (N24351, N24343, N14901, N7671, N337);
and AND4 (N24352, N24314, N14637, N173, N14777);
not NOT1 (N24353, N24334);
or OR3 (N24354, N24350, N6588, N8394);
buf BUF1 (N24355, N24353);
nor NOR4 (N24356, N24342, N18841, N13227, N22015);
and AND3 (N24357, N24356, N16015, N6427);
not NOT1 (N24358, N24346);
not NOT1 (N24359, N24354);
xor XOR2 (N24360, N24358, N13544);
not NOT1 (N24361, N24355);
buf BUF1 (N24362, N24352);
nand NAND3 (N24363, N24362, N14058, N10579);
nand NAND4 (N24364, N24351, N5847, N17241, N15882);
nor NOR4 (N24365, N24347, N12421, N23632, N9368);
buf BUF1 (N24366, N24348);
and AND2 (N24367, N24359, N2547);
and AND3 (N24368, N24357, N5487, N2552);
or OR4 (N24369, N24361, N15582, N11168, N5271);
xor XOR2 (N24370, N24349, N7153);
xor XOR2 (N24371, N24365, N12148);
buf BUF1 (N24372, N24363);
nand NAND4 (N24373, N24369, N9668, N16950, N13663);
nand NAND4 (N24374, N24360, N4293, N6231, N2476);
nor NOR4 (N24375, N24371, N17370, N22732, N8959);
buf BUF1 (N24376, N24366);
or OR4 (N24377, N24374, N10522, N4679, N1008);
not NOT1 (N24378, N24376);
not NOT1 (N24379, N24377);
buf BUF1 (N24380, N24370);
nand NAND4 (N24381, N24373, N470, N252, N14560);
and AND3 (N24382, N24375, N574, N12645);
nor NOR2 (N24383, N24380, N4493);
buf BUF1 (N24384, N24368);
not NOT1 (N24385, N24382);
nand NAND2 (N24386, N24379, N1020);
and AND2 (N24387, N24378, N1195);
xor XOR2 (N24388, N24372, N20665);
nand NAND3 (N24389, N24364, N4224, N21923);
nor NOR3 (N24390, N24344, N6968, N4601);
nand NAND3 (N24391, N24383, N23926, N5759);
nor NOR4 (N24392, N24390, N15569, N11457, N16550);
and AND3 (N24393, N24388, N6217, N22332);
nand NAND4 (N24394, N24392, N23729, N10156, N11818);
nor NOR3 (N24395, N24384, N8976, N23860);
nor NOR3 (N24396, N24381, N18147, N6089);
nor NOR2 (N24397, N24391, N10718);
xor XOR2 (N24398, N24387, N15968);
and AND2 (N24399, N24385, N22356);
nand NAND3 (N24400, N24399, N6015, N13545);
nand NAND2 (N24401, N24397, N22099);
not NOT1 (N24402, N24396);
nor NOR3 (N24403, N24401, N21684, N17626);
xor XOR2 (N24404, N24389, N3127);
and AND3 (N24405, N24404, N1750, N7833);
buf BUF1 (N24406, N24367);
nand NAND4 (N24407, N24402, N14487, N16305, N9587);
or OR2 (N24408, N24386, N10960);
buf BUF1 (N24409, N24400);
nand NAND3 (N24410, N24403, N5619, N5137);
not NOT1 (N24411, N24393);
or OR4 (N24412, N24405, N553, N10346, N18202);
and AND4 (N24413, N24412, N12425, N22068, N1484);
nand NAND4 (N24414, N24411, N17458, N16555, N7889);
nand NAND3 (N24415, N24408, N11470, N20027);
buf BUF1 (N24416, N24394);
not NOT1 (N24417, N24410);
xor XOR2 (N24418, N24409, N23862);
nor NOR3 (N24419, N24416, N12798, N4530);
and AND3 (N24420, N24415, N11954, N6576);
nand NAND4 (N24421, N24418, N19783, N7178, N14484);
nand NAND2 (N24422, N24413, N6658);
xor XOR2 (N24423, N24420, N21093);
nor NOR4 (N24424, N24419, N18498, N3956, N3483);
nor NOR3 (N24425, N24414, N10056, N7651);
buf BUF1 (N24426, N24407);
or OR3 (N24427, N24417, N1280, N10890);
not NOT1 (N24428, N24398);
nor NOR3 (N24429, N24395, N23243, N7035);
buf BUF1 (N24430, N24422);
xor XOR2 (N24431, N24424, N13511);
or OR2 (N24432, N24421, N14619);
and AND2 (N24433, N24423, N8781);
and AND2 (N24434, N24428, N10860);
not NOT1 (N24435, N24426);
nor NOR3 (N24436, N24429, N17834, N11134);
nor NOR2 (N24437, N24433, N10853);
not NOT1 (N24438, N24435);
and AND3 (N24439, N24434, N7705, N24175);
nor NOR3 (N24440, N24437, N15220, N5548);
not NOT1 (N24441, N24438);
or OR4 (N24442, N24440, N15607, N5963, N19765);
or OR2 (N24443, N24442, N19612);
or OR2 (N24444, N24427, N5145);
buf BUF1 (N24445, N24444);
not NOT1 (N24446, N24443);
buf BUF1 (N24447, N24425);
or OR4 (N24448, N24446, N6977, N18976, N2824);
not NOT1 (N24449, N24441);
nor NOR3 (N24450, N24439, N2431, N22362);
buf BUF1 (N24451, N24432);
and AND3 (N24452, N24447, N9505, N6891);
not NOT1 (N24453, N24431);
and AND4 (N24454, N24451, N23958, N8430, N23053);
nor NOR2 (N24455, N24454, N19278);
nand NAND3 (N24456, N24406, N20038, N2365);
or OR2 (N24457, N24448, N4700);
nor NOR4 (N24458, N24456, N5588, N8423, N6471);
buf BUF1 (N24459, N24449);
not NOT1 (N24460, N24459);
buf BUF1 (N24461, N24430);
buf BUF1 (N24462, N24460);
nand NAND3 (N24463, N24452, N14527, N572);
buf BUF1 (N24464, N24450);
nor NOR4 (N24465, N24445, N2294, N9530, N275);
and AND3 (N24466, N24461, N21632, N22015);
nand NAND4 (N24467, N24462, N15742, N6068, N7612);
xor XOR2 (N24468, N24464, N13588);
not NOT1 (N24469, N24467);
xor XOR2 (N24470, N24455, N20222);
or OR3 (N24471, N24463, N12818, N14789);
not NOT1 (N24472, N24457);
or OR3 (N24473, N24436, N22469, N23540);
xor XOR2 (N24474, N24469, N22474);
or OR2 (N24475, N24466, N55);
buf BUF1 (N24476, N24458);
not NOT1 (N24477, N24465);
buf BUF1 (N24478, N24472);
buf BUF1 (N24479, N24474);
or OR4 (N24480, N24473, N6765, N16400, N9836);
nor NOR2 (N24481, N24478, N11524);
buf BUF1 (N24482, N24470);
not NOT1 (N24483, N24468);
and AND2 (N24484, N24479, N11544);
and AND4 (N24485, N24471, N21368, N12983, N3387);
not NOT1 (N24486, N24453);
not NOT1 (N24487, N24475);
or OR3 (N24488, N24480, N9142, N21219);
xor XOR2 (N24489, N24484, N11754);
buf BUF1 (N24490, N24483);
nor NOR3 (N24491, N24482, N8302, N6579);
not NOT1 (N24492, N24486);
xor XOR2 (N24493, N24485, N4326);
nand NAND4 (N24494, N24492, N24202, N23383, N8062);
buf BUF1 (N24495, N24490);
or OR3 (N24496, N24481, N7276, N10539);
buf BUF1 (N24497, N24488);
not NOT1 (N24498, N24494);
and AND3 (N24499, N24491, N8284, N18339);
or OR3 (N24500, N24476, N20356, N1329);
nor NOR4 (N24501, N24497, N8378, N4914, N8947);
nor NOR2 (N24502, N24496, N22172);
buf BUF1 (N24503, N24489);
xor XOR2 (N24504, N24503, N14235);
nor NOR4 (N24505, N24499, N5854, N10789, N18885);
xor XOR2 (N24506, N24493, N1169);
nor NOR2 (N24507, N24487, N24376);
xor XOR2 (N24508, N24498, N12043);
or OR4 (N24509, N24495, N6952, N11478, N21604);
buf BUF1 (N24510, N24502);
xor XOR2 (N24511, N24500, N23290);
and AND2 (N24512, N24504, N19468);
and AND4 (N24513, N24505, N24135, N13121, N3636);
nor NOR3 (N24514, N24477, N8454, N13173);
not NOT1 (N24515, N24509);
nor NOR2 (N24516, N24501, N7727);
nand NAND4 (N24517, N24510, N15471, N8485, N16383);
nor NOR3 (N24518, N24512, N20397, N11630);
or OR3 (N24519, N24516, N898, N11391);
not NOT1 (N24520, N24513);
nand NAND4 (N24521, N24515, N24492, N20641, N12920);
nor NOR3 (N24522, N24517, N8416, N7838);
nor NOR3 (N24523, N24514, N11799, N170);
and AND4 (N24524, N24520, N12899, N22358, N7506);
and AND2 (N24525, N24506, N571);
nand NAND4 (N24526, N24523, N14210, N21727, N6811);
or OR2 (N24527, N24511, N4699);
or OR2 (N24528, N24521, N24400);
not NOT1 (N24529, N24524);
nand NAND4 (N24530, N24527, N6093, N23980, N17070);
or OR4 (N24531, N24525, N7798, N6224, N7026);
not NOT1 (N24532, N24518);
not NOT1 (N24533, N24528);
not NOT1 (N24534, N24531);
not NOT1 (N24535, N24532);
nand NAND4 (N24536, N24535, N6148, N1512, N5874);
nor NOR3 (N24537, N24533, N159, N8608);
nor NOR3 (N24538, N24530, N7795, N16875);
or OR3 (N24539, N24529, N22147, N13765);
not NOT1 (N24540, N24508);
xor XOR2 (N24541, N24537, N16140);
not NOT1 (N24542, N24538);
or OR3 (N24543, N24519, N1486, N9271);
not NOT1 (N24544, N24542);
and AND2 (N24545, N24536, N19259);
not NOT1 (N24546, N24541);
xor XOR2 (N24547, N24540, N20021);
xor XOR2 (N24548, N24526, N12229);
not NOT1 (N24549, N24544);
and AND4 (N24550, N24539, N8532, N14579, N3182);
buf BUF1 (N24551, N24507);
buf BUF1 (N24552, N24545);
buf BUF1 (N24553, N24546);
nor NOR4 (N24554, N24534, N6716, N3569, N2758);
nand NAND2 (N24555, N24550, N13387);
nand NAND3 (N24556, N24522, N950, N10292);
nor NOR4 (N24557, N24548, N17846, N11849, N3455);
nand NAND4 (N24558, N24543, N20341, N23372, N7224);
nor NOR4 (N24559, N24557, N7919, N15950, N9524);
or OR4 (N24560, N24555, N14905, N13953, N15619);
nand NAND4 (N24561, N24559, N5985, N23885, N17837);
and AND4 (N24562, N24551, N2170, N8154, N8328);
nor NOR4 (N24563, N24552, N14601, N16532, N14885);
not NOT1 (N24564, N24553);
nand NAND3 (N24565, N24562, N5689, N9859);
not NOT1 (N24566, N24554);
buf BUF1 (N24567, N24566);
nor NOR4 (N24568, N24564, N10805, N2797, N4770);
nand NAND4 (N24569, N24567, N24362, N9358, N11167);
xor XOR2 (N24570, N24561, N18910);
and AND2 (N24571, N24563, N17693);
nor NOR3 (N24572, N24560, N6154, N1597);
and AND4 (N24573, N24568, N9989, N4218, N9353);
xor XOR2 (N24574, N24570, N6803);
buf BUF1 (N24575, N24571);
and AND3 (N24576, N24549, N2096, N9132);
nor NOR2 (N24577, N24575, N9755);
or OR2 (N24578, N24573, N10611);
nor NOR3 (N24579, N24578, N4148, N9352);
or OR2 (N24580, N24574, N5876);
or OR3 (N24581, N24572, N19870, N20953);
buf BUF1 (N24582, N24576);
not NOT1 (N24583, N24569);
or OR2 (N24584, N24565, N251);
nand NAND4 (N24585, N24558, N11098, N23219, N7503);
buf BUF1 (N24586, N24585);
nand NAND3 (N24587, N24547, N3390, N12045);
nand NAND4 (N24588, N24586, N1589, N6212, N15600);
xor XOR2 (N24589, N24581, N2597);
or OR4 (N24590, N24589, N20346, N9648, N11826);
xor XOR2 (N24591, N24556, N16683);
or OR4 (N24592, N24590, N10132, N20079, N20142);
nor NOR3 (N24593, N24584, N19498, N15650);
not NOT1 (N24594, N24580);
and AND4 (N24595, N24592, N9068, N6101, N24454);
buf BUF1 (N24596, N24593);
nand NAND4 (N24597, N24577, N15496, N16497, N14589);
nor NOR2 (N24598, N24579, N13817);
and AND2 (N24599, N24591, N3867);
buf BUF1 (N24600, N24588);
buf BUF1 (N24601, N24600);
buf BUF1 (N24602, N24587);
buf BUF1 (N24603, N24596);
xor XOR2 (N24604, N24599, N1722);
nand NAND4 (N24605, N24603, N9869, N6665, N3697);
xor XOR2 (N24606, N24597, N12135);
nor NOR2 (N24607, N24605, N18751);
nand NAND3 (N24608, N24606, N2446, N12804);
or OR2 (N24609, N24598, N9633);
not NOT1 (N24610, N24582);
nand NAND4 (N24611, N24604, N5736, N13739, N17783);
nor NOR2 (N24612, N24583, N1312);
xor XOR2 (N24613, N24602, N10112);
xor XOR2 (N24614, N24594, N274);
and AND3 (N24615, N24595, N20237, N22491);
or OR2 (N24616, N24601, N23881);
nand NAND4 (N24617, N24610, N17704, N15862, N22907);
nand NAND3 (N24618, N24611, N12175, N12039);
nor NOR3 (N24619, N24613, N18594, N23423);
nor NOR2 (N24620, N24607, N19738);
buf BUF1 (N24621, N24617);
xor XOR2 (N24622, N24618, N6474);
and AND2 (N24623, N24622, N10989);
buf BUF1 (N24624, N24608);
and AND4 (N24625, N24614, N5492, N14358, N15363);
not NOT1 (N24626, N24615);
xor XOR2 (N24627, N24621, N9674);
or OR2 (N24628, N24627, N22866);
or OR2 (N24629, N24619, N22585);
nand NAND3 (N24630, N24626, N9547, N20941);
not NOT1 (N24631, N24612);
and AND4 (N24632, N24623, N1064, N16240, N1061);
and AND4 (N24633, N24616, N11065, N308, N2539);
or OR4 (N24634, N24633, N14396, N16645, N3119);
buf BUF1 (N24635, N24609);
nor NOR2 (N24636, N24632, N22510);
and AND2 (N24637, N24631, N14897);
or OR3 (N24638, N24630, N19397, N18898);
or OR2 (N24639, N24624, N24369);
not NOT1 (N24640, N24637);
nor NOR3 (N24641, N24635, N252, N6313);
or OR4 (N24642, N24638, N15199, N528, N21529);
buf BUF1 (N24643, N24641);
nand NAND2 (N24644, N24636, N13154);
nor NOR4 (N24645, N24644, N19564, N15742, N13525);
nor NOR2 (N24646, N24628, N17026);
not NOT1 (N24647, N24629);
xor XOR2 (N24648, N24643, N1226);
or OR3 (N24649, N24645, N3131, N8786);
nor NOR2 (N24650, N24620, N16725);
xor XOR2 (N24651, N24625, N4189);
buf BUF1 (N24652, N24634);
nand NAND2 (N24653, N24652, N11259);
xor XOR2 (N24654, N24650, N12355);
nand NAND3 (N24655, N24649, N10044, N16235);
xor XOR2 (N24656, N24640, N8326);
not NOT1 (N24657, N24639);
nand NAND3 (N24658, N24648, N11954, N6499);
buf BUF1 (N24659, N24651);
nand NAND2 (N24660, N24646, N24197);
nor NOR3 (N24661, N24655, N21494, N8097);
nand NAND4 (N24662, N24660, N24137, N21805, N19304);
buf BUF1 (N24663, N24654);
xor XOR2 (N24664, N24656, N418);
and AND3 (N24665, N24663, N5580, N18083);
nand NAND2 (N24666, N24653, N23996);
and AND3 (N24667, N24664, N1372, N3978);
buf BUF1 (N24668, N24667);
nor NOR4 (N24669, N24662, N18256, N13434, N20356);
nor NOR2 (N24670, N24642, N3807);
not NOT1 (N24671, N24669);
not NOT1 (N24672, N24658);
or OR2 (N24673, N24670, N17629);
nor NOR2 (N24674, N24657, N22852);
not NOT1 (N24675, N24661);
not NOT1 (N24676, N24666);
nor NOR2 (N24677, N24668, N1005);
nor NOR4 (N24678, N24674, N8981, N17554, N18236);
nor NOR2 (N24679, N24647, N1536);
xor XOR2 (N24680, N24675, N14473);
or OR3 (N24681, N24672, N19993, N20478);
not NOT1 (N24682, N24665);
nand NAND4 (N24683, N24676, N22378, N20838, N16160);
buf BUF1 (N24684, N24682);
nor NOR4 (N24685, N24671, N414, N17522, N11578);
not NOT1 (N24686, N24673);
nand NAND4 (N24687, N24683, N7997, N14357, N12222);
nor NOR3 (N24688, N24680, N2437, N23492);
nand NAND2 (N24689, N24684, N6262);
xor XOR2 (N24690, N24677, N1248);
xor XOR2 (N24691, N24686, N11709);
not NOT1 (N24692, N24690);
nand NAND2 (N24693, N24691, N20178);
buf BUF1 (N24694, N24689);
nor NOR3 (N24695, N24681, N22511, N9979);
and AND4 (N24696, N24687, N8111, N15609, N7639);
and AND3 (N24697, N24696, N18330, N21488);
buf BUF1 (N24698, N24693);
xor XOR2 (N24699, N24694, N7786);
nor NOR3 (N24700, N24692, N17595, N16222);
nand NAND3 (N24701, N24697, N1503, N1825);
or OR2 (N24702, N24700, N18099);
and AND3 (N24703, N24698, N24501, N21441);
buf BUF1 (N24704, N24679);
nand NAND4 (N24705, N24695, N14646, N503, N10017);
nor NOR4 (N24706, N24699, N9121, N7354, N20766);
nor NOR2 (N24707, N24678, N23782);
nand NAND3 (N24708, N24659, N5755, N18987);
and AND2 (N24709, N24704, N5212);
nor NOR4 (N24710, N24688, N13426, N5681, N14396);
buf BUF1 (N24711, N24708);
or OR2 (N24712, N24707, N13616);
xor XOR2 (N24713, N24711, N4462);
nand NAND4 (N24714, N24685, N5060, N14362, N3744);
nand NAND3 (N24715, N24712, N1529, N9440);
nor NOR4 (N24716, N24709, N24600, N1755, N5915);
xor XOR2 (N24717, N24705, N17194);
nor NOR2 (N24718, N24702, N3910);
or OR3 (N24719, N24710, N8723, N2243);
buf BUF1 (N24720, N24703);
or OR4 (N24721, N24701, N14125, N24579, N7191);
xor XOR2 (N24722, N24717, N3017);
and AND3 (N24723, N24716, N8947, N7742);
and AND4 (N24724, N24706, N1894, N2844, N21592);
and AND3 (N24725, N24722, N14777, N8904);
xor XOR2 (N24726, N24713, N21766);
and AND4 (N24727, N24720, N3342, N9026, N13691);
nand NAND3 (N24728, N24726, N17473, N21519);
not NOT1 (N24729, N24727);
nand NAND2 (N24730, N24729, N19298);
xor XOR2 (N24731, N24721, N6352);
not NOT1 (N24732, N24725);
buf BUF1 (N24733, N24723);
not NOT1 (N24734, N24715);
nand NAND3 (N24735, N24718, N18287, N9894);
not NOT1 (N24736, N24719);
buf BUF1 (N24737, N24731);
nand NAND2 (N24738, N24728, N7746);
nor NOR4 (N24739, N24734, N20384, N1138, N12177);
xor XOR2 (N24740, N24736, N7064);
xor XOR2 (N24741, N24740, N19014);
buf BUF1 (N24742, N24714);
nor NOR2 (N24743, N24730, N23454);
xor XOR2 (N24744, N24732, N428);
not NOT1 (N24745, N24739);
not NOT1 (N24746, N24733);
nand NAND4 (N24747, N24742, N14811, N20502, N10585);
and AND2 (N24748, N24744, N884);
nand NAND2 (N24749, N24747, N15904);
and AND3 (N24750, N24738, N21923, N21964);
xor XOR2 (N24751, N24748, N695);
or OR4 (N24752, N24750, N20103, N4941, N23010);
buf BUF1 (N24753, N24746);
xor XOR2 (N24754, N24735, N6924);
buf BUF1 (N24755, N24752);
xor XOR2 (N24756, N24724, N15529);
buf BUF1 (N24757, N24756);
xor XOR2 (N24758, N24755, N1434);
not NOT1 (N24759, N24743);
or OR4 (N24760, N24757, N23903, N15683, N19647);
and AND2 (N24761, N24741, N24417);
xor XOR2 (N24762, N24753, N24616);
nor NOR3 (N24763, N24737, N4036, N12019);
xor XOR2 (N24764, N24751, N13860);
not NOT1 (N24765, N24760);
nor NOR3 (N24766, N24764, N2421, N13198);
nor NOR2 (N24767, N24745, N20524);
nor NOR2 (N24768, N24762, N14268);
and AND3 (N24769, N24754, N21758, N9404);
buf BUF1 (N24770, N24765);
buf BUF1 (N24771, N24766);
and AND3 (N24772, N24763, N937, N18423);
or OR4 (N24773, N24770, N7874, N13194, N15593);
and AND4 (N24774, N24758, N14331, N12069, N17247);
nand NAND2 (N24775, N24761, N3012);
nor NOR3 (N24776, N24772, N17503, N19010);
nand NAND2 (N24777, N24749, N2192);
nand NAND4 (N24778, N24759, N21490, N12480, N5020);
nor NOR3 (N24779, N24771, N14008, N10585);
not NOT1 (N24780, N24768);
or OR4 (N24781, N24775, N20627, N8620, N23837);
nor NOR4 (N24782, N24777, N14408, N22305, N21403);
or OR2 (N24783, N24778, N18889);
and AND2 (N24784, N24781, N22023);
not NOT1 (N24785, N24773);
not NOT1 (N24786, N24769);
buf BUF1 (N24787, N24782);
xor XOR2 (N24788, N24780, N2740);
and AND4 (N24789, N24788, N9076, N17947, N7287);
xor XOR2 (N24790, N24787, N24327);
xor XOR2 (N24791, N24784, N7404);
buf BUF1 (N24792, N24783);
and AND2 (N24793, N24774, N6431);
or OR3 (N24794, N24785, N5633, N11061);
xor XOR2 (N24795, N24791, N7855);
nand NAND4 (N24796, N24779, N18007, N11818, N1489);
or OR4 (N24797, N24790, N9639, N2421, N23697);
nand NAND3 (N24798, N24792, N6320, N10709);
xor XOR2 (N24799, N24796, N17149);
buf BUF1 (N24800, N24793);
not NOT1 (N24801, N24800);
or OR4 (N24802, N24799, N12787, N8125, N10809);
buf BUF1 (N24803, N24798);
or OR2 (N24804, N24795, N900);
not NOT1 (N24805, N24794);
nand NAND2 (N24806, N24803, N24644);
xor XOR2 (N24807, N24786, N6969);
nand NAND2 (N24808, N24805, N22927);
or OR2 (N24809, N24801, N21098);
and AND4 (N24810, N24808, N8733, N13208, N2659);
not NOT1 (N24811, N24789);
and AND3 (N24812, N24802, N8682, N15795);
buf BUF1 (N24813, N24812);
or OR4 (N24814, N24813, N6129, N7280, N17742);
nor NOR2 (N24815, N24809, N13807);
not NOT1 (N24816, N24814);
nor NOR2 (N24817, N24767, N23879);
nor NOR2 (N24818, N24811, N6277);
not NOT1 (N24819, N24817);
xor XOR2 (N24820, N24815, N9172);
buf BUF1 (N24821, N24818);
not NOT1 (N24822, N24810);
and AND3 (N24823, N24820, N4577, N4341);
nor NOR4 (N24824, N24819, N1019, N22518, N17581);
nor NOR2 (N24825, N24823, N20693);
not NOT1 (N24826, N24776);
nand NAND4 (N24827, N24807, N14613, N314, N8888);
or OR3 (N24828, N24816, N2005, N2158);
or OR3 (N24829, N24827, N3993, N5958);
or OR4 (N24830, N24804, N11667, N6082, N13038);
xor XOR2 (N24831, N24824, N645);
not NOT1 (N24832, N24822);
not NOT1 (N24833, N24830);
buf BUF1 (N24834, N24828);
buf BUF1 (N24835, N24832);
not NOT1 (N24836, N24826);
buf BUF1 (N24837, N24821);
nor NOR4 (N24838, N24829, N4953, N21067, N15816);
nor NOR3 (N24839, N24837, N23451, N4539);
xor XOR2 (N24840, N24839, N9846);
xor XOR2 (N24841, N24831, N12482);
xor XOR2 (N24842, N24838, N4034);
buf BUF1 (N24843, N24835);
and AND3 (N24844, N24833, N10676, N12689);
or OR4 (N24845, N24841, N13811, N17041, N24654);
not NOT1 (N24846, N24836);
and AND4 (N24847, N24844, N15211, N13543, N22401);
nor NOR4 (N24848, N24825, N7297, N10420, N4580);
nand NAND4 (N24849, N24847, N8065, N18398, N23355);
nor NOR3 (N24850, N24843, N15856, N18562);
xor XOR2 (N24851, N24849, N18705);
and AND4 (N24852, N24834, N18521, N3265, N15331);
buf BUF1 (N24853, N24840);
buf BUF1 (N24854, N24848);
nand NAND3 (N24855, N24853, N4270, N21845);
nor NOR2 (N24856, N24797, N18436);
buf BUF1 (N24857, N24855);
not NOT1 (N24858, N24850);
and AND2 (N24859, N24842, N13725);
xor XOR2 (N24860, N24858, N5022);
not NOT1 (N24861, N24859);
nand NAND3 (N24862, N24861, N12449, N6810);
or OR4 (N24863, N24806, N4455, N12809, N4884);
xor XOR2 (N24864, N24845, N15558);
nand NAND3 (N24865, N24860, N7281, N4451);
not NOT1 (N24866, N24856);
nor NOR3 (N24867, N24857, N12097, N20732);
xor XOR2 (N24868, N24865, N1369);
nor NOR3 (N24869, N24852, N13307, N11514);
xor XOR2 (N24870, N24863, N20415);
xor XOR2 (N24871, N24869, N9235);
nand NAND2 (N24872, N24870, N13079);
nand NAND4 (N24873, N24866, N19233, N20597, N16939);
or OR4 (N24874, N24868, N2199, N11530, N22586);
xor XOR2 (N24875, N24854, N2624);
and AND4 (N24876, N24851, N4326, N493, N21360);
not NOT1 (N24877, N24872);
buf BUF1 (N24878, N24871);
xor XOR2 (N24879, N24873, N2899);
xor XOR2 (N24880, N24874, N19989);
xor XOR2 (N24881, N24880, N9935);
buf BUF1 (N24882, N24862);
nand NAND2 (N24883, N24879, N7938);
nor NOR3 (N24884, N24876, N6263, N18402);
and AND3 (N24885, N24884, N12107, N6164);
or OR4 (N24886, N24875, N15223, N19386, N8293);
buf BUF1 (N24887, N24877);
or OR3 (N24888, N24882, N21544, N21576);
nor NOR4 (N24889, N24886, N12536, N5472, N24006);
or OR3 (N24890, N24864, N11661, N12551);
or OR2 (N24891, N24887, N22013);
nand NAND2 (N24892, N24890, N2987);
not NOT1 (N24893, N24881);
and AND3 (N24894, N24883, N9407, N19226);
nand NAND3 (N24895, N24892, N3410, N8851);
nor NOR2 (N24896, N24878, N18582);
xor XOR2 (N24897, N24894, N7557);
xor XOR2 (N24898, N24846, N2793);
not NOT1 (N24899, N24895);
xor XOR2 (N24900, N24891, N8549);
nand NAND2 (N24901, N24898, N14582);
and AND2 (N24902, N24885, N13706);
buf BUF1 (N24903, N24900);
xor XOR2 (N24904, N24867, N24093);
not NOT1 (N24905, N24902);
nand NAND3 (N24906, N24904, N1172, N4294);
buf BUF1 (N24907, N24889);
xor XOR2 (N24908, N24905, N21607);
xor XOR2 (N24909, N24901, N984);
not NOT1 (N24910, N24888);
or OR4 (N24911, N24897, N6486, N19304, N15668);
and AND4 (N24912, N24906, N23613, N6242, N10673);
xor XOR2 (N24913, N24896, N5659);
nor NOR2 (N24914, N24908, N4866);
buf BUF1 (N24915, N24893);
nand NAND3 (N24916, N24914, N18067, N17751);
xor XOR2 (N24917, N24915, N18914);
and AND4 (N24918, N24912, N4258, N23730, N18835);
nor NOR4 (N24919, N24909, N7723, N14516, N13154);
or OR2 (N24920, N24913, N8439);
or OR2 (N24921, N24920, N24160);
buf BUF1 (N24922, N24903);
buf BUF1 (N24923, N24922);
nor NOR2 (N24924, N24921, N14802);
or OR3 (N24925, N24918, N4423, N15365);
nor NOR2 (N24926, N24907, N14359);
buf BUF1 (N24927, N24919);
xor XOR2 (N24928, N24927, N5358);
nor NOR4 (N24929, N24916, N558, N2390, N356);
nand NAND2 (N24930, N24917, N2293);
xor XOR2 (N24931, N24911, N18838);
nand NAND4 (N24932, N24929, N9007, N9322, N4285);
and AND4 (N24933, N24931, N18124, N13937, N9221);
not NOT1 (N24934, N24899);
and AND2 (N24935, N24930, N2167);
nand NAND2 (N24936, N24910, N1017);
nand NAND3 (N24937, N24928, N17168, N1540);
or OR2 (N24938, N24933, N14773);
and AND3 (N24939, N24923, N20682, N19989);
buf BUF1 (N24940, N24937);
or OR4 (N24941, N24935, N12105, N21964, N10315);
not NOT1 (N24942, N24924);
xor XOR2 (N24943, N24932, N6209);
or OR4 (N24944, N24939, N9109, N11328, N14975);
buf BUF1 (N24945, N24925);
or OR4 (N24946, N24938, N6504, N10431, N13257);
or OR4 (N24947, N24942, N2864, N16509, N23238);
nor NOR3 (N24948, N24940, N751, N11821);
nor NOR3 (N24949, N24947, N22034, N16517);
not NOT1 (N24950, N24946);
nor NOR2 (N24951, N24936, N1452);
buf BUF1 (N24952, N24926);
nand NAND2 (N24953, N24948, N18960);
nor NOR2 (N24954, N24951, N24110);
buf BUF1 (N24955, N24943);
xor XOR2 (N24956, N24955, N20406);
or OR4 (N24957, N24956, N365, N11400, N11638);
buf BUF1 (N24958, N24952);
buf BUF1 (N24959, N24941);
and AND4 (N24960, N24949, N958, N23773, N19934);
buf BUF1 (N24961, N24934);
buf BUF1 (N24962, N24944);
nand NAND3 (N24963, N24958, N9418, N21331);
xor XOR2 (N24964, N24963, N5136);
nand NAND4 (N24965, N24950, N7530, N7638, N8454);
buf BUF1 (N24966, N24954);
or OR3 (N24967, N24961, N15932, N13986);
xor XOR2 (N24968, N24967, N4359);
not NOT1 (N24969, N24959);
nand NAND2 (N24970, N24957, N17297);
buf BUF1 (N24971, N24962);
xor XOR2 (N24972, N24971, N18251);
xor XOR2 (N24973, N24966, N2862);
xor XOR2 (N24974, N24965, N20214);
buf BUF1 (N24975, N24972);
nand NAND4 (N24976, N24968, N20105, N14605, N12230);
not NOT1 (N24977, N24975);
or OR2 (N24978, N24960, N5269);
and AND4 (N24979, N24964, N10776, N17335, N14122);
nor NOR3 (N24980, N24976, N12338, N3492);
nand NAND4 (N24981, N24973, N14736, N1518, N9);
buf BUF1 (N24982, N24978);
or OR3 (N24983, N24982, N3289, N18411);
nand NAND2 (N24984, N24980, N18386);
nor NOR2 (N24985, N24984, N10606);
nor NOR3 (N24986, N24981, N20007, N16854);
buf BUF1 (N24987, N24986);
buf BUF1 (N24988, N24953);
xor XOR2 (N24989, N24969, N170);
not NOT1 (N24990, N24974);
nor NOR4 (N24991, N24977, N18712, N10340, N3151);
nor NOR4 (N24992, N24945, N20333, N16256, N2058);
not NOT1 (N24993, N24979);
nor NOR3 (N24994, N24985, N3375, N14320);
buf BUF1 (N24995, N24990);
xor XOR2 (N24996, N24991, N21614);
nand NAND4 (N24997, N24988, N5529, N14612, N18229);
not NOT1 (N24998, N24993);
nand NAND2 (N24999, N24992, N20628);
nor NOR2 (N25000, N24997, N4598);
not NOT1 (N25001, N24999);
and AND2 (N25002, N24996, N7726);
nand NAND3 (N25003, N24998, N1096, N18326);
nand NAND2 (N25004, N24970, N17753);
xor XOR2 (N25005, N25001, N12049);
or OR3 (N25006, N25002, N903, N7245);
not NOT1 (N25007, N25000);
xor XOR2 (N25008, N25005, N18794);
xor XOR2 (N25009, N24994, N5219);
xor XOR2 (N25010, N24989, N14860);
or OR2 (N25011, N25003, N18854);
xor XOR2 (N25012, N24983, N8378);
buf BUF1 (N25013, N24995);
buf BUF1 (N25014, N25010);
and AND4 (N25015, N25007, N24604, N7566, N18316);
nand NAND2 (N25016, N24987, N217);
nor NOR2 (N25017, N25014, N12602);
and AND2 (N25018, N25004, N16644);
or OR4 (N25019, N25012, N12727, N5928, N24082);
xor XOR2 (N25020, N25013, N8780);
nand NAND4 (N25021, N25006, N19464, N13506, N2301);
or OR2 (N25022, N25009, N11308);
not NOT1 (N25023, N25021);
xor XOR2 (N25024, N25022, N20458);
nor NOR4 (N25025, N25019, N18174, N21365, N23291);
buf BUF1 (N25026, N25023);
nand NAND3 (N25027, N25018, N17280, N8783);
buf BUF1 (N25028, N25017);
buf BUF1 (N25029, N25024);
nor NOR3 (N25030, N25029, N11215, N1329);
buf BUF1 (N25031, N25027);
xor XOR2 (N25032, N25030, N21965);
nand NAND4 (N25033, N25008, N8838, N2574, N3050);
and AND3 (N25034, N25025, N959, N3610);
nor NOR2 (N25035, N25026, N15047);
or OR3 (N25036, N25028, N19107, N17120);
and AND2 (N25037, N25020, N21609);
buf BUF1 (N25038, N25033);
and AND4 (N25039, N25038, N4443, N18922, N16786);
buf BUF1 (N25040, N25011);
buf BUF1 (N25041, N25035);
nand NAND3 (N25042, N25040, N18833, N21746);
or OR2 (N25043, N25032, N64);
nor NOR4 (N25044, N25039, N24890, N4738, N12796);
or OR4 (N25045, N25016, N15027, N17016, N14049);
and AND3 (N25046, N25036, N18400, N15574);
and AND3 (N25047, N25031, N20508, N15613);
buf BUF1 (N25048, N25046);
or OR2 (N25049, N25043, N23639);
nor NOR4 (N25050, N25045, N3440, N512, N24870);
buf BUF1 (N25051, N25037);
buf BUF1 (N25052, N25048);
not NOT1 (N25053, N25044);
not NOT1 (N25054, N25053);
xor XOR2 (N25055, N25052, N22054);
not NOT1 (N25056, N25041);
not NOT1 (N25057, N25054);
nand NAND4 (N25058, N25056, N5355, N12611, N24788);
and AND3 (N25059, N25051, N21894, N12922);
nand NAND3 (N25060, N25050, N9621, N1339);
nor NOR2 (N25061, N25057, N10570);
xor XOR2 (N25062, N25059, N20741);
and AND4 (N25063, N25034, N9079, N3509, N20877);
nor NOR2 (N25064, N25061, N20043);
or OR4 (N25065, N25042, N21807, N2074, N21132);
or OR2 (N25066, N25063, N6702);
not NOT1 (N25067, N25065);
buf BUF1 (N25068, N25067);
xor XOR2 (N25069, N25068, N17829);
not NOT1 (N25070, N25062);
or OR4 (N25071, N25049, N13974, N5077, N48);
nor NOR3 (N25072, N25060, N11592, N14377);
or OR2 (N25073, N25047, N4831);
nor NOR3 (N25074, N25064, N2134, N3866);
xor XOR2 (N25075, N25058, N12499);
xor XOR2 (N25076, N25066, N13462);
not NOT1 (N25077, N25070);
xor XOR2 (N25078, N25075, N5704);
or OR4 (N25079, N25072, N1737, N20980, N19915);
not NOT1 (N25080, N25079);
xor XOR2 (N25081, N25073, N21547);
and AND2 (N25082, N25081, N496);
buf BUF1 (N25083, N25071);
nand NAND3 (N25084, N25078, N819, N19243);
nor NOR2 (N25085, N25015, N24512);
not NOT1 (N25086, N25083);
nor NOR4 (N25087, N25085, N15882, N24029, N22278);
nor NOR4 (N25088, N25055, N12292, N2425, N2173);
not NOT1 (N25089, N25077);
and AND3 (N25090, N25082, N16536, N526);
xor XOR2 (N25091, N25086, N12701);
and AND2 (N25092, N25090, N8814);
xor XOR2 (N25093, N25076, N3870);
xor XOR2 (N25094, N25080, N22211);
nand NAND2 (N25095, N25091, N20989);
or OR4 (N25096, N25087, N20559, N1991, N4730);
and AND4 (N25097, N25093, N1230, N12964, N14665);
buf BUF1 (N25098, N25096);
or OR3 (N25099, N25094, N5721, N22797);
buf BUF1 (N25100, N25099);
nor NOR4 (N25101, N25097, N5984, N22781, N21815);
nor NOR3 (N25102, N25100, N16422, N8761);
nand NAND3 (N25103, N25092, N6558, N2201);
not NOT1 (N25104, N25095);
buf BUF1 (N25105, N25103);
and AND2 (N25106, N25098, N22591);
xor XOR2 (N25107, N25102, N8454);
and AND4 (N25108, N25104, N9549, N19572, N4245);
or OR3 (N25109, N25107, N13346, N18367);
and AND3 (N25110, N25105, N7524, N1869);
not NOT1 (N25111, N25084);
buf BUF1 (N25112, N25074);
nand NAND3 (N25113, N25109, N2003, N790);
buf BUF1 (N25114, N25106);
xor XOR2 (N25115, N25110, N12983);
not NOT1 (N25116, N25111);
not NOT1 (N25117, N25088);
not NOT1 (N25118, N25117);
and AND3 (N25119, N25118, N18701, N12933);
nand NAND4 (N25120, N25108, N4274, N4865, N5077);
not NOT1 (N25121, N25115);
not NOT1 (N25122, N25114);
nor NOR2 (N25123, N25122, N5091);
nor NOR3 (N25124, N25112, N5655, N22564);
and AND3 (N25125, N25120, N14422, N10944);
nand NAND4 (N25126, N25113, N13436, N21969, N11271);
not NOT1 (N25127, N25125);
xor XOR2 (N25128, N25123, N17274);
xor XOR2 (N25129, N25069, N23158);
and AND4 (N25130, N25128, N21543, N17030, N14429);
not NOT1 (N25131, N25101);
not NOT1 (N25132, N25127);
and AND4 (N25133, N25130, N11609, N13596, N21819);
nor NOR3 (N25134, N25126, N18840, N8822);
or OR3 (N25135, N25089, N21414, N9726);
buf BUF1 (N25136, N25124);
nor NOR3 (N25137, N25132, N16117, N19501);
xor XOR2 (N25138, N25136, N14134);
nand NAND3 (N25139, N25134, N24414, N12770);
xor XOR2 (N25140, N25121, N7485);
buf BUF1 (N25141, N25129);
and AND3 (N25142, N25137, N16964, N21898);
not NOT1 (N25143, N25119);
nor NOR2 (N25144, N25142, N5618);
not NOT1 (N25145, N25141);
nand NAND4 (N25146, N25140, N1141, N23453, N11686);
nor NOR3 (N25147, N25143, N10688, N20886);
nor NOR2 (N25148, N25116, N5819);
nor NOR4 (N25149, N25133, N19147, N313, N6055);
nor NOR2 (N25150, N25135, N22067);
nand NAND4 (N25151, N25150, N10217, N6556, N23801);
nor NOR3 (N25152, N25147, N20938, N20076);
xor XOR2 (N25153, N25146, N12422);
nor NOR2 (N25154, N25151, N5766);
xor XOR2 (N25155, N25152, N6291);
not NOT1 (N25156, N25155);
or OR4 (N25157, N25138, N8264, N18294, N20590);
xor XOR2 (N25158, N25154, N25057);
or OR2 (N25159, N25145, N20902);
and AND4 (N25160, N25149, N8178, N2389, N2278);
and AND3 (N25161, N25131, N20316, N24758);
nor NOR2 (N25162, N25139, N24686);
or OR4 (N25163, N25161, N24549, N24782, N14815);
buf BUF1 (N25164, N25153);
nand NAND3 (N25165, N25148, N4490, N25163);
buf BUF1 (N25166, N17652);
not NOT1 (N25167, N25144);
or OR2 (N25168, N25156, N10975);
not NOT1 (N25169, N25160);
buf BUF1 (N25170, N25167);
not NOT1 (N25171, N25166);
and AND2 (N25172, N25159, N9991);
xor XOR2 (N25173, N25165, N18193);
nand NAND4 (N25174, N25158, N20699, N14869, N18491);
nand NAND3 (N25175, N25168, N7174, N12096);
buf BUF1 (N25176, N25169);
nor NOR2 (N25177, N25170, N11631);
nor NOR3 (N25178, N25176, N11896, N10161);
not NOT1 (N25179, N25173);
nand NAND4 (N25180, N25172, N6273, N9585, N3200);
and AND4 (N25181, N25174, N10105, N9997, N19763);
or OR2 (N25182, N25175, N10472);
nand NAND4 (N25183, N25157, N17711, N3096, N12311);
buf BUF1 (N25184, N25171);
nor NOR3 (N25185, N25162, N2949, N19601);
and AND2 (N25186, N25179, N554);
nand NAND2 (N25187, N25180, N9553);
not NOT1 (N25188, N25187);
nand NAND2 (N25189, N25188, N17637);
not NOT1 (N25190, N25189);
nand NAND3 (N25191, N25177, N7798, N5159);
not NOT1 (N25192, N25186);
nand NAND3 (N25193, N25182, N675, N18459);
nor NOR3 (N25194, N25192, N17471, N22103);
and AND4 (N25195, N25191, N13024, N3444, N189);
or OR4 (N25196, N25194, N807, N22547, N13036);
not NOT1 (N25197, N25196);
and AND3 (N25198, N25178, N12423, N2008);
xor XOR2 (N25199, N25183, N13697);
and AND2 (N25200, N25197, N5363);
nand NAND4 (N25201, N25198, N24360, N1940, N4518);
and AND4 (N25202, N25199, N10835, N9481, N1366);
nand NAND3 (N25203, N25202, N18911, N832);
or OR2 (N25204, N25164, N5985);
buf BUF1 (N25205, N25184);
nand NAND3 (N25206, N25205, N888, N23297);
and AND2 (N25207, N25200, N22057);
buf BUF1 (N25208, N25207);
nand NAND4 (N25209, N25206, N6995, N23624, N16848);
nor NOR4 (N25210, N25190, N21250, N6816, N5329);
not NOT1 (N25211, N25210);
and AND3 (N25212, N25193, N11080, N5534);
and AND4 (N25213, N25203, N17401, N11224, N3541);
nor NOR4 (N25214, N25195, N22197, N2631, N13020);
not NOT1 (N25215, N25185);
nor NOR4 (N25216, N25208, N15670, N1385, N9605);
buf BUF1 (N25217, N25211);
and AND4 (N25218, N25214, N18777, N10648, N10408);
buf BUF1 (N25219, N25201);
xor XOR2 (N25220, N25181, N10641);
and AND2 (N25221, N25216, N20027);
or OR2 (N25222, N25215, N21552);
nand NAND2 (N25223, N25209, N18353);
not NOT1 (N25224, N25219);
nor NOR2 (N25225, N25223, N5799);
xor XOR2 (N25226, N25212, N15074);
xor XOR2 (N25227, N25222, N3345);
xor XOR2 (N25228, N25220, N5517);
nand NAND3 (N25229, N25221, N20111, N2703);
and AND4 (N25230, N25228, N15477, N24940, N17010);
nand NAND4 (N25231, N25224, N10383, N16015, N20619);
buf BUF1 (N25232, N25213);
or OR4 (N25233, N25229, N5793, N9572, N22497);
not NOT1 (N25234, N25204);
xor XOR2 (N25235, N25232, N8549);
xor XOR2 (N25236, N25231, N12620);
or OR4 (N25237, N25235, N22092, N22346, N10356);
xor XOR2 (N25238, N25234, N18563);
nor NOR4 (N25239, N25233, N6789, N17198, N24034);
nand NAND4 (N25240, N25238, N25238, N17473, N12885);
buf BUF1 (N25241, N25227);
buf BUF1 (N25242, N25225);
xor XOR2 (N25243, N25241, N4745);
or OR4 (N25244, N25240, N14463, N13807, N11014);
nor NOR4 (N25245, N25226, N7279, N12938, N21280);
and AND4 (N25246, N25239, N15967, N11689, N7159);
or OR4 (N25247, N25230, N12790, N21054, N24347);
and AND2 (N25248, N25236, N4082);
nor NOR2 (N25249, N25218, N1440);
not NOT1 (N25250, N25249);
not NOT1 (N25251, N25217);
nor NOR3 (N25252, N25243, N24319, N16286);
xor XOR2 (N25253, N25251, N18894);
not NOT1 (N25254, N25237);
and AND4 (N25255, N25247, N5363, N1033, N7681);
or OR3 (N25256, N25250, N14387, N9972);
buf BUF1 (N25257, N25253);
buf BUF1 (N25258, N25255);
buf BUF1 (N25259, N25246);
xor XOR2 (N25260, N25248, N5083);
and AND4 (N25261, N25257, N10895, N16975, N11956);
and AND4 (N25262, N25260, N11373, N18155, N14275);
nand NAND3 (N25263, N25254, N13428, N8189);
buf BUF1 (N25264, N25242);
nand NAND2 (N25265, N25264, N17289);
not NOT1 (N25266, N25262);
not NOT1 (N25267, N25265);
nand NAND3 (N25268, N25252, N7727, N20166);
and AND3 (N25269, N25245, N14232, N17114);
nand NAND3 (N25270, N25244, N5552, N193);
nor NOR4 (N25271, N25268, N14738, N775, N21169);
nor NOR3 (N25272, N25271, N13259, N5411);
not NOT1 (N25273, N25270);
not NOT1 (N25274, N25261);
nand NAND2 (N25275, N25258, N15071);
nand NAND2 (N25276, N25263, N20877);
nor NOR4 (N25277, N25275, N14583, N13333, N13825);
nor NOR3 (N25278, N25274, N18753, N11895);
buf BUF1 (N25279, N25277);
nor NOR3 (N25280, N25266, N20831, N8833);
or OR2 (N25281, N25273, N3351);
or OR4 (N25282, N25267, N8572, N16523, N24935);
nor NOR4 (N25283, N25259, N24002, N4054, N18950);
nand NAND3 (N25284, N25276, N7828, N3618);
nand NAND3 (N25285, N25280, N7979, N21720);
nand NAND4 (N25286, N25279, N21457, N24981, N9784);
or OR2 (N25287, N25281, N23494);
nor NOR4 (N25288, N25283, N10009, N16090, N10743);
and AND3 (N25289, N25288, N14280, N13658);
not NOT1 (N25290, N25285);
xor XOR2 (N25291, N25278, N638);
or OR2 (N25292, N25287, N491);
nor NOR2 (N25293, N25282, N8705);
not NOT1 (N25294, N25293);
and AND4 (N25295, N25269, N22397, N3986, N7503);
xor XOR2 (N25296, N25291, N20523);
nor NOR3 (N25297, N25290, N20018, N14886);
nand NAND2 (N25298, N25256, N16446);
nor NOR3 (N25299, N25298, N17097, N21852);
nor NOR4 (N25300, N25297, N24567, N4968, N7569);
buf BUF1 (N25301, N25299);
nand NAND4 (N25302, N25286, N24244, N1780, N24212);
nand NAND4 (N25303, N25272, N16184, N23474, N23262);
and AND3 (N25304, N25302, N10503, N12348);
nand NAND3 (N25305, N25300, N22131, N5084);
nor NOR3 (N25306, N25292, N7937, N7564);
xor XOR2 (N25307, N25295, N21330);
nor NOR3 (N25308, N25303, N20378, N3300);
nor NOR4 (N25309, N25284, N5870, N23100, N10230);
nand NAND4 (N25310, N25308, N12758, N15210, N23628);
nor NOR2 (N25311, N25301, N25131);
nand NAND4 (N25312, N25294, N7895, N10806, N9326);
nand NAND2 (N25313, N25309, N4609);
buf BUF1 (N25314, N25289);
nor NOR4 (N25315, N25314, N410, N16731, N21797);
not NOT1 (N25316, N25296);
xor XOR2 (N25317, N25315, N15215);
xor XOR2 (N25318, N25312, N19704);
not NOT1 (N25319, N25311);
nand NAND3 (N25320, N25319, N5102, N18654);
buf BUF1 (N25321, N25310);
nor NOR2 (N25322, N25313, N16202);
or OR2 (N25323, N25322, N1360);
not NOT1 (N25324, N25318);
xor XOR2 (N25325, N25307, N8647);
or OR4 (N25326, N25321, N24489, N9123, N15780);
or OR2 (N25327, N25306, N22231);
nand NAND4 (N25328, N25316, N15863, N9482, N25029);
and AND4 (N25329, N25317, N21281, N5662, N3339);
and AND4 (N25330, N25329, N14909, N6648, N3560);
nor NOR3 (N25331, N25328, N15739, N12592);
buf BUF1 (N25332, N25326);
buf BUF1 (N25333, N25305);
or OR4 (N25334, N25333, N10240, N20433, N20884);
xor XOR2 (N25335, N25330, N7777);
xor XOR2 (N25336, N25335, N22830);
and AND4 (N25337, N25334, N7029, N3600, N20906);
buf BUF1 (N25338, N25324);
nand NAND4 (N25339, N25337, N12828, N13244, N7847);
and AND3 (N25340, N25336, N17228, N2302);
not NOT1 (N25341, N25332);
nand NAND3 (N25342, N25327, N751, N7);
and AND2 (N25343, N25325, N15403);
xor XOR2 (N25344, N25331, N5239);
nor NOR4 (N25345, N25339, N11452, N13555, N7399);
xor XOR2 (N25346, N25343, N10963);
nand NAND4 (N25347, N25338, N8830, N9507, N21175);
nand NAND2 (N25348, N25346, N13753);
nand NAND4 (N25349, N25342, N1909, N4033, N5733);
or OR3 (N25350, N25320, N4852, N22128);
or OR3 (N25351, N25323, N4423, N14357);
not NOT1 (N25352, N25345);
buf BUF1 (N25353, N25348);
buf BUF1 (N25354, N25351);
not NOT1 (N25355, N25349);
or OR4 (N25356, N25341, N8462, N13680, N23164);
and AND2 (N25357, N25344, N17177);
and AND4 (N25358, N25354, N10935, N10904, N2843);
nand NAND4 (N25359, N25356, N21885, N10408, N23512);
or OR4 (N25360, N25358, N24177, N14978, N21080);
xor XOR2 (N25361, N25352, N18957);
nor NOR3 (N25362, N25355, N962, N18063);
buf BUF1 (N25363, N25362);
or OR4 (N25364, N25359, N1959, N18030, N2621);
nor NOR3 (N25365, N25304, N3713, N16398);
and AND2 (N25366, N25347, N10663);
xor XOR2 (N25367, N25365, N14192);
not NOT1 (N25368, N25350);
nor NOR3 (N25369, N25366, N10769, N17495);
and AND2 (N25370, N25367, N843);
and AND3 (N25371, N25361, N15862, N761);
buf BUF1 (N25372, N25369);
buf BUF1 (N25373, N25370);
nor NOR4 (N25374, N25353, N3101, N1078, N18281);
and AND2 (N25375, N25371, N12348);
nand NAND2 (N25376, N25363, N6747);
not NOT1 (N25377, N25375);
not NOT1 (N25378, N25376);
nor NOR4 (N25379, N25372, N7229, N12373, N10172);
or OR3 (N25380, N25360, N4049, N2278);
xor XOR2 (N25381, N25374, N13256);
nor NOR2 (N25382, N25379, N18439);
nand NAND3 (N25383, N25381, N7814, N6169);
xor XOR2 (N25384, N25357, N24481);
or OR4 (N25385, N25340, N7864, N15127, N8264);
or OR4 (N25386, N25368, N6838, N1255, N10564);
not NOT1 (N25387, N25383);
nor NOR4 (N25388, N25380, N8017, N8007, N14626);
nor NOR4 (N25389, N25382, N4040, N20288, N12309);
nand NAND4 (N25390, N25389, N22286, N6383, N16056);
not NOT1 (N25391, N25377);
xor XOR2 (N25392, N25384, N16098);
xor XOR2 (N25393, N25390, N17656);
not NOT1 (N25394, N25387);
not NOT1 (N25395, N25393);
xor XOR2 (N25396, N25394, N3433);
buf BUF1 (N25397, N25391);
nor NOR2 (N25398, N25385, N24508);
not NOT1 (N25399, N25398);
nand NAND4 (N25400, N25396, N17114, N15092, N3981);
buf BUF1 (N25401, N25378);
buf BUF1 (N25402, N25395);
and AND2 (N25403, N25401, N7346);
buf BUF1 (N25404, N25397);
nor NOR4 (N25405, N25388, N16906, N23667, N5309);
nor NOR3 (N25406, N25405, N14248, N20479);
and AND4 (N25407, N25400, N19081, N7487, N20673);
nor NOR3 (N25408, N25402, N15818, N7737);
buf BUF1 (N25409, N25404);
nand NAND2 (N25410, N25407, N10308);
and AND4 (N25411, N25373, N16400, N16107, N4029);
xor XOR2 (N25412, N25386, N22347);
not NOT1 (N25413, N25403);
and AND3 (N25414, N25411, N247, N10600);
buf BUF1 (N25415, N25408);
xor XOR2 (N25416, N25364, N20888);
buf BUF1 (N25417, N25409);
nand NAND3 (N25418, N25392, N19659, N25228);
or OR4 (N25419, N25415, N5320, N20181, N4257);
nand NAND3 (N25420, N25406, N6663, N3666);
nor NOR3 (N25421, N25419, N22601, N4922);
nand NAND3 (N25422, N25416, N7711, N18936);
not NOT1 (N25423, N25418);
nand NAND3 (N25424, N25421, N21317, N6449);
xor XOR2 (N25425, N25420, N7782);
not NOT1 (N25426, N25412);
or OR4 (N25427, N25422, N10511, N16255, N16646);
nor NOR2 (N25428, N25423, N19405);
not NOT1 (N25429, N25428);
nor NOR2 (N25430, N25426, N8950);
not NOT1 (N25431, N25417);
nor NOR3 (N25432, N25431, N1443, N18384);
buf BUF1 (N25433, N25430);
nand NAND3 (N25434, N25414, N1216, N20634);
not NOT1 (N25435, N25432);
and AND3 (N25436, N25410, N2273, N25232);
xor XOR2 (N25437, N25424, N20365);
xor XOR2 (N25438, N25433, N4083);
buf BUF1 (N25439, N25434);
xor XOR2 (N25440, N25399, N3777);
xor XOR2 (N25441, N25436, N19577);
nand NAND3 (N25442, N25425, N2612, N22021);
nor NOR4 (N25443, N25438, N19467, N1308, N16052);
or OR3 (N25444, N25441, N6945, N17876);
or OR3 (N25445, N25439, N3990, N24190);
and AND4 (N25446, N25437, N10699, N787, N15873);
xor XOR2 (N25447, N25435, N11032);
buf BUF1 (N25448, N25442);
and AND2 (N25449, N25448, N7565);
xor XOR2 (N25450, N25427, N19123);
or OR3 (N25451, N25449, N20384, N20071);
not NOT1 (N25452, N25450);
buf BUF1 (N25453, N25440);
not NOT1 (N25454, N25453);
and AND3 (N25455, N25452, N1928, N11512);
nor NOR2 (N25456, N25445, N11004);
xor XOR2 (N25457, N25455, N10202);
nor NOR2 (N25458, N25446, N1113);
or OR3 (N25459, N25429, N23108, N1004);
nor NOR2 (N25460, N25458, N22401);
not NOT1 (N25461, N25447);
and AND4 (N25462, N25459, N6379, N5637, N10318);
and AND2 (N25463, N25461, N17857);
xor XOR2 (N25464, N25451, N1041);
nand NAND4 (N25465, N25456, N17939, N3144, N12939);
buf BUF1 (N25466, N25444);
buf BUF1 (N25467, N25457);
and AND4 (N25468, N25462, N21775, N1891, N115);
xor XOR2 (N25469, N25443, N8997);
nor NOR2 (N25470, N25464, N9372);
nand NAND4 (N25471, N25466, N16670, N20966, N23901);
xor XOR2 (N25472, N25463, N9786);
nand NAND4 (N25473, N25465, N23607, N853, N7145);
nand NAND3 (N25474, N25469, N21966, N20709);
or OR4 (N25475, N25471, N11828, N17411, N6973);
nand NAND2 (N25476, N25468, N9771);
xor XOR2 (N25477, N25413, N23343);
or OR4 (N25478, N25454, N24358, N21142, N11714);
and AND3 (N25479, N25472, N19476, N8346);
or OR4 (N25480, N25460, N19848, N9696, N24641);
buf BUF1 (N25481, N25479);
not NOT1 (N25482, N25478);
and AND3 (N25483, N25475, N10309, N9268);
xor XOR2 (N25484, N25467, N2055);
or OR2 (N25485, N25483, N19974);
xor XOR2 (N25486, N25476, N17610);
nand NAND3 (N25487, N25480, N18248, N9947);
nand NAND3 (N25488, N25473, N21446, N20737);
or OR4 (N25489, N25474, N4893, N4299, N8230);
or OR3 (N25490, N25488, N2012, N9126);
nor NOR2 (N25491, N25477, N9030);
or OR3 (N25492, N25489, N13874, N22040);
and AND4 (N25493, N25491, N5681, N21412, N259);
nor NOR3 (N25494, N25492, N12510, N24636);
xor XOR2 (N25495, N25470, N7933);
or OR3 (N25496, N25490, N20267, N2650);
xor XOR2 (N25497, N25495, N9394);
and AND3 (N25498, N25494, N1, N17429);
or OR2 (N25499, N25485, N5389);
xor XOR2 (N25500, N25493, N15978);
nor NOR4 (N25501, N25500, N25499, N3177, N14862);
nand NAND2 (N25502, N1821, N23662);
nor NOR3 (N25503, N25496, N15577, N673);
or OR2 (N25504, N25486, N11220);
or OR3 (N25505, N25502, N25485, N12351);
buf BUF1 (N25506, N25503);
and AND4 (N25507, N25506, N25483, N8630, N10638);
not NOT1 (N25508, N25487);
nand NAND4 (N25509, N25481, N11117, N9321, N16935);
not NOT1 (N25510, N25482);
nand NAND2 (N25511, N25509, N11721);
or OR3 (N25512, N25501, N6368, N15400);
nand NAND3 (N25513, N25498, N14022, N2929);
nand NAND3 (N25514, N25511, N13801, N3760);
xor XOR2 (N25515, N25512, N6451);
or OR3 (N25516, N25513, N8780, N15378);
and AND3 (N25517, N25497, N8219, N8346);
xor XOR2 (N25518, N25504, N18772);
nand NAND3 (N25519, N25484, N5070, N3696);
and AND3 (N25520, N25516, N14918, N18319);
xor XOR2 (N25521, N25505, N4798);
buf BUF1 (N25522, N25518);
nand NAND2 (N25523, N25520, N1790);
and AND4 (N25524, N25523, N15868, N16653, N14832);
not NOT1 (N25525, N25508);
or OR4 (N25526, N25521, N2139, N21229, N16614);
nand NAND2 (N25527, N25522, N3761);
nand NAND4 (N25528, N25515, N3621, N23430, N11041);
or OR3 (N25529, N25526, N13379, N15988);
xor XOR2 (N25530, N25510, N4543);
nand NAND2 (N25531, N25517, N13142);
or OR3 (N25532, N25530, N10881, N8840);
xor XOR2 (N25533, N25528, N15106);
nor NOR2 (N25534, N25507, N8015);
buf BUF1 (N25535, N25534);
nor NOR3 (N25536, N25525, N4136, N11102);
and AND4 (N25537, N25535, N22289, N12131, N16938);
or OR2 (N25538, N25531, N15363);
nand NAND2 (N25539, N25532, N23078);
buf BUF1 (N25540, N25514);
nor NOR2 (N25541, N25537, N23719);
buf BUF1 (N25542, N25519);
not NOT1 (N25543, N25538);
not NOT1 (N25544, N25543);
nor NOR3 (N25545, N25539, N12870, N6820);
nor NOR2 (N25546, N25540, N6225);
or OR3 (N25547, N25536, N16999, N4193);
and AND2 (N25548, N25527, N15459);
xor XOR2 (N25549, N25524, N13481);
nor NOR3 (N25550, N25548, N23892, N19870);
not NOT1 (N25551, N25547);
and AND3 (N25552, N25549, N3483, N13224);
buf BUF1 (N25553, N25545);
and AND2 (N25554, N25546, N12117);
or OR2 (N25555, N25552, N3551);
and AND4 (N25556, N25533, N15648, N21521, N5768);
nor NOR2 (N25557, N25553, N5070);
buf BUF1 (N25558, N25555);
nand NAND3 (N25559, N25557, N1432, N4491);
xor XOR2 (N25560, N25554, N3971);
nand NAND3 (N25561, N25556, N8154, N4224);
xor XOR2 (N25562, N25551, N15492);
not NOT1 (N25563, N25550);
nand NAND4 (N25564, N25559, N260, N16962, N4367);
or OR2 (N25565, N25544, N3372);
or OR2 (N25566, N25563, N4543);
nand NAND4 (N25567, N25542, N21653, N3978, N14397);
or OR3 (N25568, N25561, N11589, N12575);
xor XOR2 (N25569, N25541, N12193);
buf BUF1 (N25570, N25558);
or OR4 (N25571, N25568, N963, N164, N18973);
not NOT1 (N25572, N25565);
buf BUF1 (N25573, N25569);
not NOT1 (N25574, N25572);
nor NOR2 (N25575, N25571, N2106);
nor NOR2 (N25576, N25566, N25513);
nor NOR3 (N25577, N25529, N3492, N4644);
buf BUF1 (N25578, N25575);
xor XOR2 (N25579, N25562, N20829);
xor XOR2 (N25580, N25577, N1844);
nor NOR2 (N25581, N25564, N25190);
xor XOR2 (N25582, N25560, N17146);
xor XOR2 (N25583, N25576, N21160);
not NOT1 (N25584, N25582);
or OR3 (N25585, N25581, N985, N8143);
nor NOR2 (N25586, N25579, N1692);
xor XOR2 (N25587, N25573, N5741);
or OR3 (N25588, N25584, N20704, N6814);
nand NAND3 (N25589, N25567, N17573, N24474);
nand NAND3 (N25590, N25589, N25307, N10487);
or OR4 (N25591, N25586, N11060, N4495, N17598);
nand NAND3 (N25592, N25570, N20424, N12149);
and AND2 (N25593, N25588, N14026);
not NOT1 (N25594, N25574);
nor NOR3 (N25595, N25585, N24301, N19285);
or OR2 (N25596, N25595, N7100);
or OR3 (N25597, N25592, N5971, N12462);
xor XOR2 (N25598, N25597, N19381);
and AND4 (N25599, N25587, N11020, N855, N7958);
not NOT1 (N25600, N25598);
and AND3 (N25601, N25583, N13454, N2227);
and AND4 (N25602, N25578, N16555, N21770, N11621);
xor XOR2 (N25603, N25596, N4994);
nor NOR4 (N25604, N25594, N11522, N6456, N11713);
and AND2 (N25605, N25599, N12781);
xor XOR2 (N25606, N25580, N14487);
nor NOR2 (N25607, N25604, N10819);
nand NAND3 (N25608, N25603, N11040, N13041);
nand NAND2 (N25609, N25605, N21734);
buf BUF1 (N25610, N25600);
not NOT1 (N25611, N25602);
buf BUF1 (N25612, N25609);
xor XOR2 (N25613, N25601, N22176);
buf BUF1 (N25614, N25610);
nand NAND2 (N25615, N25608, N3665);
xor XOR2 (N25616, N25611, N23414);
not NOT1 (N25617, N25591);
xor XOR2 (N25618, N25606, N18351);
buf BUF1 (N25619, N25607);
buf BUF1 (N25620, N25619);
buf BUF1 (N25621, N25614);
nand NAND4 (N25622, N25618, N17505, N9710, N19243);
nor NOR2 (N25623, N25613, N5537);
endmodule