// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23;

output N3013,N3018,N3006,N3009,N3016,N3008,N3014,N3022,N3015,N3023;

xor XOR2 (N24, N18, N4);
nor NOR4 (N25, N1, N5, N9, N18);
or OR4 (N26, N10, N15, N14, N13);
buf BUF1 (N27, N12);
or OR3 (N28, N22, N5, N4);
or OR2 (N29, N18, N20);
nor NOR2 (N30, N22, N20);
nor NOR4 (N31, N7, N2, N22, N13);
or OR4 (N32, N19, N5, N15, N8);
buf BUF1 (N33, N29);
nand NAND2 (N34, N15, N29);
nor NOR4 (N35, N30, N27, N16, N22);
nor NOR4 (N36, N3, N12, N12, N8);
nor NOR2 (N37, N24, N20);
nor NOR3 (N38, N37, N30, N25);
and AND4 (N39, N33, N14, N29, N4);
nand NAND2 (N40, N13, N7);
not NOT1 (N41, N34);
xor XOR2 (N42, N32, N41);
or OR3 (N43, N41, N27, N10);
and AND2 (N44, N38, N39);
not NOT1 (N45, N20);
and AND3 (N46, N26, N41, N16);
xor XOR2 (N47, N42, N16);
not NOT1 (N48, N40);
nor NOR3 (N49, N28, N46, N36);
not NOT1 (N50, N9);
xor XOR2 (N51, N34, N23);
not NOT1 (N52, N45);
xor XOR2 (N53, N51, N3);
not NOT1 (N54, N44);
nor NOR4 (N55, N48, N33, N26, N35);
not NOT1 (N56, N21);
xor XOR2 (N57, N55, N1);
and AND3 (N58, N52, N24, N16);
buf BUF1 (N59, N54);
buf BUF1 (N60, N53);
xor XOR2 (N61, N49, N6);
buf BUF1 (N62, N59);
buf BUF1 (N63, N50);
not NOT1 (N64, N43);
or OR2 (N65, N47, N33);
or OR2 (N66, N57, N36);
nor NOR3 (N67, N61, N48, N29);
nand NAND2 (N68, N56, N26);
or OR2 (N69, N64, N27);
nor NOR2 (N70, N65, N62);
or OR3 (N71, N32, N54, N22);
not NOT1 (N72, N69);
or OR4 (N73, N68, N33, N32, N6);
nor NOR2 (N74, N58, N23);
xor XOR2 (N75, N73, N67);
nor NOR2 (N76, N60, N34);
or OR3 (N77, N37, N43, N46);
and AND2 (N78, N63, N12);
and AND2 (N79, N71, N23);
buf BUF1 (N80, N76);
and AND3 (N81, N70, N7, N23);
buf BUF1 (N82, N72);
nor NOR3 (N83, N31, N78, N54);
nand NAND4 (N84, N65, N13, N28, N77);
buf BUF1 (N85, N40);
and AND4 (N86, N85, N5, N49, N78);
nor NOR4 (N87, N75, N14, N78, N19);
and AND4 (N88, N83, N41, N37, N31);
nor NOR4 (N89, N80, N80, N30, N62);
buf BUF1 (N90, N82);
not NOT1 (N91, N87);
or OR2 (N92, N79, N70);
not NOT1 (N93, N89);
or OR2 (N94, N74, N65);
nand NAND2 (N95, N91, N88);
nand NAND3 (N96, N75, N18, N74);
or OR3 (N97, N96, N11, N30);
nor NOR2 (N98, N81, N43);
nand NAND2 (N99, N94, N10);
nor NOR4 (N100, N95, N94, N48, N28);
and AND3 (N101, N100, N61, N57);
or OR2 (N102, N98, N89);
and AND3 (N103, N90, N1, N84);
and AND3 (N104, N101, N10, N24);
buf BUF1 (N105, N68);
not NOT1 (N106, N105);
nand NAND4 (N107, N92, N79, N80, N55);
and AND4 (N108, N102, N32, N35, N97);
buf BUF1 (N109, N61);
xor XOR2 (N110, N93, N37);
or OR2 (N111, N110, N37);
and AND4 (N112, N104, N37, N21, N61);
xor XOR2 (N113, N66, N95);
and AND4 (N114, N86, N42, N73, N89);
xor XOR2 (N115, N113, N85);
buf BUF1 (N116, N107);
and AND2 (N117, N108, N67);
or OR2 (N118, N115, N101);
and AND3 (N119, N103, N33, N42);
buf BUF1 (N120, N99);
and AND2 (N121, N119, N17);
nor NOR3 (N122, N106, N70, N33);
not NOT1 (N123, N118);
not NOT1 (N124, N121);
nor NOR3 (N125, N120, N33, N35);
buf BUF1 (N126, N125);
buf BUF1 (N127, N112);
nand NAND4 (N128, N111, N118, N77, N121);
and AND3 (N129, N126, N109, N103);
buf BUF1 (N130, N97);
xor XOR2 (N131, N128, N112);
xor XOR2 (N132, N130, N33);
not NOT1 (N133, N123);
nor NOR2 (N134, N129, N29);
nand NAND4 (N135, N124, N40, N12, N16);
nand NAND4 (N136, N131, N98, N67, N27);
nor NOR2 (N137, N114, N32);
not NOT1 (N138, N127);
buf BUF1 (N139, N116);
and AND2 (N140, N132, N39);
xor XOR2 (N141, N135, N26);
and AND3 (N142, N137, N66, N128);
nor NOR4 (N143, N133, N122, N114, N109);
or OR2 (N144, N121, N70);
not NOT1 (N145, N139);
not NOT1 (N146, N141);
xor XOR2 (N147, N136, N5);
and AND2 (N148, N117, N142);
or OR2 (N149, N131, N132);
or OR4 (N150, N147, N124, N31, N26);
buf BUF1 (N151, N146);
xor XOR2 (N152, N143, N89);
buf BUF1 (N153, N150);
not NOT1 (N154, N153);
and AND2 (N155, N144, N134);
not NOT1 (N156, N114);
nand NAND2 (N157, N156, N6);
or OR3 (N158, N138, N125, N149);
nand NAND3 (N159, N36, N7, N74);
nor NOR3 (N160, N157, N70, N40);
and AND2 (N161, N140, N121);
xor XOR2 (N162, N145, N99);
buf BUF1 (N163, N158);
or OR4 (N164, N159, N93, N66, N112);
and AND4 (N165, N148, N90, N59, N105);
nor NOR4 (N166, N163, N9, N68, N139);
buf BUF1 (N167, N160);
or OR2 (N168, N161, N60);
not NOT1 (N169, N165);
nand NAND3 (N170, N164, N89, N153);
or OR3 (N171, N151, N143, N91);
nand NAND4 (N172, N170, N19, N96, N170);
or OR3 (N173, N152, N165, N46);
nand NAND3 (N174, N172, N132, N77);
nor NOR4 (N175, N171, N100, N107, N29);
nand NAND3 (N176, N167, N105, N13);
buf BUF1 (N177, N168);
buf BUF1 (N178, N169);
or OR3 (N179, N173, N12, N35);
buf BUF1 (N180, N175);
buf BUF1 (N181, N179);
xor XOR2 (N182, N155, N62);
xor XOR2 (N183, N154, N61);
buf BUF1 (N184, N183);
or OR2 (N185, N181, N23);
xor XOR2 (N186, N166, N108);
nor NOR4 (N187, N177, N73, N81, N141);
or OR2 (N188, N178, N177);
or OR2 (N189, N162, N50);
nor NOR2 (N190, N185, N146);
nand NAND2 (N191, N190, N60);
nand NAND2 (N192, N186, N164);
buf BUF1 (N193, N174);
or OR3 (N194, N191, N32, N181);
xor XOR2 (N195, N182, N49);
or OR4 (N196, N176, N176, N50, N148);
nand NAND3 (N197, N195, N145, N59);
nor NOR2 (N198, N196, N175);
not NOT1 (N199, N197);
xor XOR2 (N200, N193, N199);
or OR4 (N201, N128, N31, N103, N55);
xor XOR2 (N202, N194, N33);
and AND2 (N203, N198, N45);
xor XOR2 (N204, N180, N12);
buf BUF1 (N205, N204);
buf BUF1 (N206, N184);
or OR3 (N207, N202, N186, N112);
not NOT1 (N208, N187);
nor NOR3 (N209, N208, N170, N65);
and AND3 (N210, N189, N174, N182);
and AND3 (N211, N205, N37, N139);
not NOT1 (N212, N210);
buf BUF1 (N213, N192);
nand NAND2 (N214, N200, N208);
or OR3 (N215, N212, N46, N102);
or OR3 (N216, N215, N109, N83);
or OR3 (N217, N216, N191, N91);
and AND4 (N218, N214, N77, N168, N209);
or OR2 (N219, N193, N59);
nand NAND2 (N220, N201, N164);
not NOT1 (N221, N220);
and AND4 (N222, N206, N20, N81, N105);
and AND3 (N223, N217, N159, N26);
not NOT1 (N224, N221);
nand NAND2 (N225, N219, N203);
xor XOR2 (N226, N173, N166);
xor XOR2 (N227, N218, N20);
and AND2 (N228, N207, N51);
not NOT1 (N229, N211);
buf BUF1 (N230, N227);
buf BUF1 (N231, N213);
or OR4 (N232, N231, N41, N149, N75);
xor XOR2 (N233, N228, N75);
xor XOR2 (N234, N229, N179);
nand NAND2 (N235, N233, N15);
nor NOR3 (N236, N230, N162, N79);
and AND3 (N237, N222, N73, N59);
xor XOR2 (N238, N236, N201);
and AND4 (N239, N232, N113, N39, N33);
nand NAND3 (N240, N224, N36, N117);
xor XOR2 (N241, N225, N223);
buf BUF1 (N242, N95);
and AND4 (N243, N234, N23, N119, N85);
not NOT1 (N244, N242);
xor XOR2 (N245, N240, N130);
not NOT1 (N246, N226);
or OR4 (N247, N245, N205, N240, N104);
buf BUF1 (N248, N247);
buf BUF1 (N249, N248);
buf BUF1 (N250, N235);
and AND3 (N251, N246, N44, N62);
or OR2 (N252, N251, N168);
buf BUF1 (N253, N249);
xor XOR2 (N254, N239, N157);
nor NOR2 (N255, N243, N26);
and AND3 (N256, N237, N141, N30);
and AND4 (N257, N244, N39, N142, N100);
buf BUF1 (N258, N252);
nor NOR4 (N259, N250, N140, N70, N183);
nor NOR2 (N260, N238, N145);
not NOT1 (N261, N253);
nor NOR4 (N262, N259, N182, N214, N85);
buf BUF1 (N263, N241);
or OR3 (N264, N260, N199, N105);
xor XOR2 (N265, N256, N121);
and AND2 (N266, N261, N76);
nor NOR2 (N267, N262, N185);
or OR4 (N268, N264, N70, N124, N128);
buf BUF1 (N269, N258);
nor NOR4 (N270, N254, N239, N231, N11);
or OR4 (N271, N268, N36, N233, N42);
or OR3 (N272, N265, N233, N179);
nor NOR2 (N273, N257, N21);
buf BUF1 (N274, N269);
buf BUF1 (N275, N266);
and AND2 (N276, N271, N226);
nand NAND2 (N277, N270, N222);
or OR4 (N278, N276, N212, N62, N223);
and AND2 (N279, N188, N84);
nor NOR2 (N280, N279, N214);
xor XOR2 (N281, N263, N167);
and AND2 (N282, N275, N49);
nor NOR3 (N283, N281, N24, N137);
or OR3 (N284, N267, N115, N195);
or OR4 (N285, N278, N43, N41, N62);
nor NOR2 (N286, N273, N246);
not NOT1 (N287, N274);
xor XOR2 (N288, N282, N77);
and AND2 (N289, N285, N67);
or OR3 (N290, N288, N167, N11);
nor NOR3 (N291, N284, N109, N70);
nor NOR3 (N292, N286, N164, N74);
nand NAND4 (N293, N291, N142, N162, N111);
or OR3 (N294, N293, N145, N218);
xor XOR2 (N295, N290, N27);
xor XOR2 (N296, N287, N192);
buf BUF1 (N297, N296);
xor XOR2 (N298, N295, N76);
nand NAND3 (N299, N255, N89, N234);
nand NAND2 (N300, N292, N169);
not NOT1 (N301, N272);
nor NOR2 (N302, N289, N202);
or OR2 (N303, N298, N151);
nor NOR4 (N304, N300, N30, N28, N25);
and AND2 (N305, N302, N78);
xor XOR2 (N306, N303, N238);
nand NAND4 (N307, N277, N143, N19, N94);
buf BUF1 (N308, N306);
not NOT1 (N309, N308);
xor XOR2 (N310, N283, N130);
and AND4 (N311, N310, N250, N226, N203);
and AND2 (N312, N297, N260);
nor NOR3 (N313, N299, N138, N184);
buf BUF1 (N314, N294);
nor NOR2 (N315, N304, N155);
nor NOR2 (N316, N307, N252);
xor XOR2 (N317, N316, N157);
or OR3 (N318, N315, N282, N53);
nand NAND4 (N319, N301, N308, N184, N151);
xor XOR2 (N320, N319, N37);
or OR3 (N321, N312, N279, N231);
not NOT1 (N322, N314);
and AND3 (N323, N322, N33, N311);
nand NAND4 (N324, N74, N318, N123, N257);
nand NAND4 (N325, N176, N71, N136, N224);
or OR4 (N326, N320, N122, N222, N113);
and AND4 (N327, N323, N129, N134, N285);
nor NOR4 (N328, N280, N92, N305, N149);
nor NOR4 (N329, N266, N327, N40, N215);
buf BUF1 (N330, N115);
or OR4 (N331, N324, N260, N88, N3);
buf BUF1 (N332, N317);
and AND4 (N333, N309, N91, N230, N5);
not NOT1 (N334, N313);
nand NAND3 (N335, N325, N163, N311);
nor NOR2 (N336, N334, N27);
or OR4 (N337, N328, N151, N69, N271);
nand NAND3 (N338, N332, N259, N317);
or OR4 (N339, N330, N305, N5, N327);
not NOT1 (N340, N336);
or OR4 (N341, N335, N84, N312, N137);
buf BUF1 (N342, N331);
nand NAND4 (N343, N341, N247, N222, N172);
and AND3 (N344, N342, N285, N71);
or OR3 (N345, N339, N3, N239);
and AND4 (N346, N321, N63, N139, N160);
buf BUF1 (N347, N343);
nor NOR4 (N348, N337, N298, N214, N249);
nor NOR3 (N349, N333, N26, N82);
and AND2 (N350, N348, N296);
and AND4 (N351, N350, N96, N106, N221);
xor XOR2 (N352, N344, N89);
or OR2 (N353, N340, N31);
xor XOR2 (N354, N346, N200);
and AND4 (N355, N347, N95, N170, N41);
not NOT1 (N356, N352);
nand NAND4 (N357, N353, N256, N195, N130);
not NOT1 (N358, N326);
not NOT1 (N359, N329);
or OR3 (N360, N355, N154, N104);
nor NOR2 (N361, N360, N308);
nor NOR2 (N362, N354, N97);
not NOT1 (N363, N362);
nor NOR3 (N364, N357, N306, N197);
and AND2 (N365, N349, N340);
or OR2 (N366, N338, N160);
buf BUF1 (N367, N351);
or OR3 (N368, N356, N233, N219);
buf BUF1 (N369, N367);
or OR2 (N370, N363, N359);
nor NOR4 (N371, N225, N40, N142, N259);
nor NOR4 (N372, N364, N316, N128, N350);
or OR3 (N373, N345, N166, N92);
buf BUF1 (N374, N368);
nand NAND2 (N375, N374, N37);
not NOT1 (N376, N370);
nand NAND2 (N377, N366, N179);
nand NAND2 (N378, N373, N37);
nor NOR3 (N379, N372, N235, N179);
nand NAND3 (N380, N377, N73, N59);
xor XOR2 (N381, N379, N86);
nor NOR2 (N382, N378, N294);
xor XOR2 (N383, N365, N285);
buf BUF1 (N384, N381);
xor XOR2 (N385, N358, N262);
not NOT1 (N386, N384);
or OR2 (N387, N380, N324);
buf BUF1 (N388, N385);
xor XOR2 (N389, N371, N36);
buf BUF1 (N390, N375);
and AND3 (N391, N369, N34, N222);
nor NOR3 (N392, N383, N108, N347);
nand NAND2 (N393, N389, N217);
not NOT1 (N394, N386);
not NOT1 (N395, N393);
not NOT1 (N396, N376);
not NOT1 (N397, N391);
buf BUF1 (N398, N395);
xor XOR2 (N399, N382, N102);
nor NOR3 (N400, N388, N161, N14);
xor XOR2 (N401, N398, N158);
and AND4 (N402, N390, N290, N345, N1);
not NOT1 (N403, N392);
or OR3 (N404, N399, N198, N374);
xor XOR2 (N405, N361, N220);
nand NAND4 (N406, N396, N41, N274, N322);
not NOT1 (N407, N404);
nand NAND2 (N408, N400, N135);
or OR3 (N409, N408, N83, N28);
and AND2 (N410, N402, N374);
not NOT1 (N411, N387);
not NOT1 (N412, N403);
nor NOR4 (N413, N411, N346, N14, N110);
not NOT1 (N414, N412);
not NOT1 (N415, N401);
buf BUF1 (N416, N407);
not NOT1 (N417, N397);
nand NAND4 (N418, N410, N286, N143, N138);
nand NAND3 (N419, N405, N347, N87);
nor NOR4 (N420, N406, N67, N280, N315);
or OR3 (N421, N413, N95, N278);
or OR4 (N422, N421, N200, N405, N260);
not NOT1 (N423, N418);
buf BUF1 (N424, N420);
nor NOR3 (N425, N394, N315, N42);
nand NAND3 (N426, N415, N395, N289);
not NOT1 (N427, N416);
nand NAND4 (N428, N426, N129, N236, N297);
and AND4 (N429, N422, N423, N190, N332);
xor XOR2 (N430, N396, N209);
nand NAND4 (N431, N425, N336, N8, N166);
or OR2 (N432, N427, N190);
or OR3 (N433, N424, N412, N144);
buf BUF1 (N434, N429);
not NOT1 (N435, N433);
not NOT1 (N436, N419);
not NOT1 (N437, N436);
xor XOR2 (N438, N409, N118);
nor NOR3 (N439, N435, N297, N213);
xor XOR2 (N440, N430, N349);
not NOT1 (N441, N437);
buf BUF1 (N442, N428);
xor XOR2 (N443, N432, N4);
xor XOR2 (N444, N443, N21);
buf BUF1 (N445, N441);
nand NAND4 (N446, N444, N190, N153, N420);
or OR3 (N447, N440, N261, N54);
and AND4 (N448, N434, N181, N414, N3);
xor XOR2 (N449, N275, N132);
xor XOR2 (N450, N442, N114);
buf BUF1 (N451, N450);
nor NOR2 (N452, N439, N407);
or OR2 (N453, N451, N110);
xor XOR2 (N454, N453, N314);
nand NAND4 (N455, N417, N200, N32, N197);
xor XOR2 (N456, N445, N403);
not NOT1 (N457, N431);
or OR3 (N458, N456, N368, N438);
not NOT1 (N459, N52);
buf BUF1 (N460, N449);
xor XOR2 (N461, N457, N231);
and AND2 (N462, N458, N131);
xor XOR2 (N463, N447, N117);
buf BUF1 (N464, N448);
not NOT1 (N465, N461);
nor NOR3 (N466, N462, N293, N156);
and AND2 (N467, N460, N465);
nand NAND4 (N468, N213, N243, N47, N45);
or OR2 (N469, N454, N126);
nor NOR3 (N470, N455, N159, N329);
buf BUF1 (N471, N466);
or OR2 (N472, N471, N125);
nand NAND4 (N473, N446, N385, N50, N394);
nor NOR3 (N474, N452, N347, N90);
xor XOR2 (N475, N464, N222);
buf BUF1 (N476, N463);
nor NOR3 (N477, N475, N225, N457);
nand NAND3 (N478, N476, N350, N292);
buf BUF1 (N479, N467);
xor XOR2 (N480, N468, N450);
and AND3 (N481, N469, N168, N371);
nor NOR2 (N482, N459, N120);
xor XOR2 (N483, N474, N51);
or OR4 (N484, N483, N190, N157, N483);
and AND2 (N485, N482, N138);
xor XOR2 (N486, N477, N452);
xor XOR2 (N487, N473, N232);
xor XOR2 (N488, N470, N114);
nor NOR2 (N489, N472, N103);
buf BUF1 (N490, N478);
buf BUF1 (N491, N480);
nand NAND4 (N492, N488, N168, N469, N372);
nor NOR4 (N493, N489, N56, N425, N464);
or OR3 (N494, N485, N135, N9);
xor XOR2 (N495, N481, N328);
and AND3 (N496, N492, N378, N315);
nor NOR3 (N497, N496, N276, N91);
buf BUF1 (N498, N479);
or OR3 (N499, N486, N99, N469);
nand NAND3 (N500, N487, N103, N446);
xor XOR2 (N501, N497, N313);
not NOT1 (N502, N498);
or OR2 (N503, N484, N205);
not NOT1 (N504, N501);
nor NOR2 (N505, N499, N39);
or OR2 (N506, N500, N229);
not NOT1 (N507, N503);
buf BUF1 (N508, N493);
buf BUF1 (N509, N506);
or OR3 (N510, N494, N477, N205);
or OR2 (N511, N495, N79);
nand NAND3 (N512, N510, N85, N229);
nand NAND2 (N513, N511, N509);
not NOT1 (N514, N2);
buf BUF1 (N515, N504);
buf BUF1 (N516, N515);
buf BUF1 (N517, N490);
not NOT1 (N518, N517);
or OR3 (N519, N512, N141, N427);
and AND4 (N520, N505, N332, N446, N19);
and AND3 (N521, N507, N39, N170);
or OR4 (N522, N520, N430, N257, N484);
nor NOR4 (N523, N519, N31, N100, N116);
nand NAND2 (N524, N502, N450);
xor XOR2 (N525, N508, N477);
nand NAND3 (N526, N514, N203, N292);
nor NOR3 (N527, N491, N36, N429);
xor XOR2 (N528, N518, N267);
xor XOR2 (N529, N528, N397);
nor NOR2 (N530, N524, N320);
or OR3 (N531, N522, N321, N498);
nor NOR2 (N532, N530, N63);
nand NAND3 (N533, N525, N464, N110);
and AND4 (N534, N513, N157, N49, N300);
xor XOR2 (N535, N527, N528);
not NOT1 (N536, N529);
nor NOR2 (N537, N535, N39);
not NOT1 (N538, N533);
nand NAND4 (N539, N526, N336, N438, N162);
xor XOR2 (N540, N538, N309);
nor NOR2 (N541, N536, N49);
xor XOR2 (N542, N523, N217);
nor NOR4 (N543, N521, N344, N185, N51);
xor XOR2 (N544, N516, N413);
not NOT1 (N545, N539);
not NOT1 (N546, N540);
not NOT1 (N547, N542);
xor XOR2 (N548, N531, N456);
and AND4 (N549, N537, N84, N147, N333);
nand NAND2 (N550, N543, N100);
xor XOR2 (N551, N532, N385);
and AND2 (N552, N541, N395);
xor XOR2 (N553, N552, N471);
xor XOR2 (N554, N553, N313);
buf BUF1 (N555, N534);
nor NOR2 (N556, N555, N384);
and AND4 (N557, N554, N98, N33, N38);
or OR4 (N558, N549, N206, N292, N371);
and AND2 (N559, N544, N493);
not NOT1 (N560, N546);
xor XOR2 (N561, N551, N304);
buf BUF1 (N562, N557);
or OR4 (N563, N556, N535, N419, N298);
nand NAND3 (N564, N561, N195, N480);
nand NAND2 (N565, N560, N39);
or OR3 (N566, N548, N524, N503);
and AND4 (N567, N562, N470, N549, N74);
nor NOR2 (N568, N550, N178);
not NOT1 (N569, N558);
buf BUF1 (N570, N545);
or OR3 (N571, N567, N191, N7);
and AND2 (N572, N563, N331);
nand NAND2 (N573, N569, N170);
not NOT1 (N574, N559);
not NOT1 (N575, N547);
buf BUF1 (N576, N574);
or OR3 (N577, N568, N566, N39);
nor NOR2 (N578, N216, N222);
buf BUF1 (N579, N570);
and AND2 (N580, N565, N429);
xor XOR2 (N581, N575, N9);
and AND4 (N582, N572, N215, N560, N223);
not NOT1 (N583, N577);
not NOT1 (N584, N583);
buf BUF1 (N585, N582);
or OR2 (N586, N576, N508);
and AND3 (N587, N571, N413, N41);
buf BUF1 (N588, N580);
buf BUF1 (N589, N584);
nand NAND3 (N590, N589, N505, N524);
or OR2 (N591, N585, N41);
or OR2 (N592, N564, N290);
and AND3 (N593, N591, N248, N323);
or OR2 (N594, N586, N216);
not NOT1 (N595, N588);
not NOT1 (N596, N587);
or OR4 (N597, N573, N393, N296, N418);
nor NOR3 (N598, N579, N427, N390);
xor XOR2 (N599, N595, N231);
buf BUF1 (N600, N596);
and AND2 (N601, N593, N443);
buf BUF1 (N602, N581);
and AND4 (N603, N600, N230, N180, N2);
and AND3 (N604, N601, N283, N100);
or OR3 (N605, N599, N361, N229);
nor NOR2 (N606, N603, N82);
xor XOR2 (N607, N602, N250);
xor XOR2 (N608, N578, N280);
not NOT1 (N609, N604);
or OR3 (N610, N590, N461, N410);
buf BUF1 (N611, N609);
xor XOR2 (N612, N606, N157);
and AND3 (N613, N607, N161, N185);
or OR3 (N614, N613, N480, N33);
and AND2 (N615, N610, N44);
or OR4 (N616, N597, N479, N336, N361);
nor NOR4 (N617, N611, N55, N359, N552);
not NOT1 (N618, N608);
nor NOR2 (N619, N592, N543);
or OR3 (N620, N615, N449, N333);
not NOT1 (N621, N619);
xor XOR2 (N622, N594, N285);
nor NOR3 (N623, N620, N292, N614);
or OR3 (N624, N272, N473, N493);
nor NOR4 (N625, N623, N403, N608, N398);
or OR3 (N626, N624, N17, N559);
buf BUF1 (N627, N621);
nor NOR2 (N628, N616, N573);
nand NAND3 (N629, N628, N506, N424);
nor NOR2 (N630, N612, N87);
not NOT1 (N631, N625);
nor NOR3 (N632, N631, N601, N125);
nor NOR2 (N633, N598, N379);
xor XOR2 (N634, N622, N19);
buf BUF1 (N635, N605);
nor NOR4 (N636, N630, N614, N466, N464);
and AND4 (N637, N618, N317, N253, N340);
or OR2 (N638, N627, N143);
nor NOR3 (N639, N638, N251, N312);
not NOT1 (N640, N626);
buf BUF1 (N641, N617);
nand NAND4 (N642, N635, N234, N554, N170);
nor NOR3 (N643, N634, N382, N33);
or OR4 (N644, N642, N455, N640, N558);
buf BUF1 (N645, N167);
buf BUF1 (N646, N636);
nor NOR2 (N647, N639, N115);
nor NOR4 (N648, N632, N346, N130, N375);
or OR3 (N649, N647, N599, N571);
nand NAND2 (N650, N649, N57);
and AND4 (N651, N643, N8, N76, N610);
nand NAND4 (N652, N644, N287, N359, N284);
nor NOR4 (N653, N646, N547, N442, N24);
not NOT1 (N654, N648);
nor NOR3 (N655, N633, N394, N480);
or OR4 (N656, N641, N442, N32, N497);
buf BUF1 (N657, N656);
and AND4 (N658, N653, N531, N621, N33);
or OR2 (N659, N637, N194);
nor NOR4 (N660, N645, N580, N308, N57);
nor NOR4 (N661, N660, N604, N450, N268);
buf BUF1 (N662, N657);
not NOT1 (N663, N651);
or OR3 (N664, N650, N152, N58);
xor XOR2 (N665, N664, N541);
buf BUF1 (N666, N659);
or OR4 (N667, N658, N308, N399, N162);
and AND2 (N668, N661, N150);
xor XOR2 (N669, N629, N159);
or OR2 (N670, N654, N115);
not NOT1 (N671, N665);
not NOT1 (N672, N667);
and AND3 (N673, N666, N264, N404);
not NOT1 (N674, N655);
buf BUF1 (N675, N668);
buf BUF1 (N676, N674);
or OR2 (N677, N671, N285);
xor XOR2 (N678, N662, N320);
or OR3 (N679, N652, N118, N209);
not NOT1 (N680, N679);
nand NAND3 (N681, N672, N255, N630);
buf BUF1 (N682, N663);
not NOT1 (N683, N675);
xor XOR2 (N684, N673, N637);
or OR4 (N685, N683, N463, N650, N630);
not NOT1 (N686, N680);
nand NAND2 (N687, N678, N218);
nor NOR4 (N688, N670, N213, N141, N71);
buf BUF1 (N689, N685);
buf BUF1 (N690, N688);
or OR2 (N691, N669, N561);
and AND4 (N692, N691, N230, N531, N436);
xor XOR2 (N693, N677, N51);
xor XOR2 (N694, N681, N152);
nor NOR2 (N695, N694, N529);
and AND3 (N696, N676, N676, N291);
nand NAND2 (N697, N684, N362);
nand NAND2 (N698, N690, N667);
not NOT1 (N699, N698);
or OR2 (N700, N699, N690);
buf BUF1 (N701, N700);
xor XOR2 (N702, N686, N661);
buf BUF1 (N703, N692);
and AND4 (N704, N693, N448, N88, N47);
and AND3 (N705, N697, N347, N510);
or OR2 (N706, N695, N256);
buf BUF1 (N707, N703);
nor NOR2 (N708, N705, N122);
not NOT1 (N709, N708);
nand NAND4 (N710, N696, N248, N600, N172);
buf BUF1 (N711, N710);
nor NOR3 (N712, N682, N704, N627);
nand NAND2 (N713, N468, N482);
not NOT1 (N714, N713);
not NOT1 (N715, N712);
and AND4 (N716, N714, N590, N377, N21);
not NOT1 (N717, N711);
nand NAND3 (N718, N687, N564, N464);
xor XOR2 (N719, N702, N317);
nor NOR4 (N720, N707, N202, N552, N682);
or OR4 (N721, N709, N226, N39, N553);
xor XOR2 (N722, N720, N161);
xor XOR2 (N723, N715, N513);
and AND3 (N724, N723, N636, N481);
or OR3 (N725, N724, N195, N150);
buf BUF1 (N726, N716);
nand NAND2 (N727, N722, N483);
or OR4 (N728, N689, N617, N439, N188);
not NOT1 (N729, N717);
and AND4 (N730, N726, N319, N145, N406);
nand NAND2 (N731, N721, N277);
or OR4 (N732, N718, N515, N708, N90);
nand NAND2 (N733, N731, N607);
not NOT1 (N734, N732);
buf BUF1 (N735, N701);
buf BUF1 (N736, N728);
nand NAND3 (N737, N719, N234, N668);
and AND4 (N738, N729, N556, N347, N178);
or OR4 (N739, N727, N381, N17, N192);
nand NAND2 (N740, N736, N509);
not NOT1 (N741, N739);
nor NOR3 (N742, N737, N318, N300);
or OR3 (N743, N738, N305, N257);
not NOT1 (N744, N730);
nor NOR4 (N745, N741, N438, N368, N332);
not NOT1 (N746, N745);
or OR3 (N747, N706, N20, N122);
nand NAND2 (N748, N743, N282);
not NOT1 (N749, N748);
not NOT1 (N750, N740);
buf BUF1 (N751, N733);
not NOT1 (N752, N746);
xor XOR2 (N753, N751, N667);
buf BUF1 (N754, N744);
nand NAND3 (N755, N735, N69, N390);
not NOT1 (N756, N749);
buf BUF1 (N757, N725);
nor NOR3 (N758, N755, N154, N186);
or OR2 (N759, N756, N629);
or OR2 (N760, N757, N390);
and AND2 (N761, N747, N213);
buf BUF1 (N762, N758);
nand NAND2 (N763, N750, N478);
and AND3 (N764, N760, N86, N89);
nor NOR4 (N765, N759, N205, N116, N2);
not NOT1 (N766, N754);
not NOT1 (N767, N734);
or OR3 (N768, N763, N697, N370);
nand NAND2 (N769, N768, N596);
or OR4 (N770, N753, N59, N236, N16);
and AND4 (N771, N767, N540, N78, N630);
not NOT1 (N772, N742);
buf BUF1 (N773, N752);
not NOT1 (N774, N769);
or OR4 (N775, N761, N420, N411, N680);
or OR2 (N776, N773, N248);
buf BUF1 (N777, N774);
and AND3 (N778, N775, N634, N31);
xor XOR2 (N779, N776, N391);
or OR2 (N780, N764, N253);
nand NAND4 (N781, N779, N621, N512, N499);
xor XOR2 (N782, N780, N330);
and AND3 (N783, N772, N333, N342);
or OR4 (N784, N777, N778, N250, N242);
xor XOR2 (N785, N182, N554);
not NOT1 (N786, N771);
nor NOR4 (N787, N781, N180, N199, N120);
buf BUF1 (N788, N762);
nor NOR3 (N789, N765, N434, N283);
and AND2 (N790, N783, N97);
not NOT1 (N791, N787);
nor NOR4 (N792, N785, N228, N388, N571);
and AND3 (N793, N792, N275, N253);
buf BUF1 (N794, N791);
or OR2 (N795, N788, N487);
or OR3 (N796, N790, N622, N734);
buf BUF1 (N797, N782);
nor NOR3 (N798, N766, N365, N98);
not NOT1 (N799, N770);
xor XOR2 (N800, N789, N95);
or OR2 (N801, N798, N176);
nand NAND4 (N802, N795, N269, N658, N322);
and AND4 (N803, N801, N410, N318, N3);
nand NAND3 (N804, N799, N362, N730);
not NOT1 (N805, N804);
and AND4 (N806, N786, N394, N154, N107);
and AND4 (N807, N793, N674, N705, N318);
not NOT1 (N808, N807);
nand NAND3 (N809, N794, N736, N380);
or OR2 (N810, N806, N430);
xor XOR2 (N811, N808, N304);
xor XOR2 (N812, N796, N58);
nand NAND2 (N813, N805, N765);
xor XOR2 (N814, N797, N227);
nand NAND2 (N815, N812, N433);
and AND3 (N816, N811, N517, N45);
xor XOR2 (N817, N815, N130);
nor NOR3 (N818, N802, N665, N574);
or OR3 (N819, N800, N738, N522);
and AND4 (N820, N810, N507, N49, N99);
and AND4 (N821, N820, N423, N163, N772);
xor XOR2 (N822, N809, N38);
not NOT1 (N823, N784);
and AND4 (N824, N821, N578, N55, N357);
and AND3 (N825, N813, N439, N778);
nand NAND4 (N826, N819, N588, N130, N735);
nor NOR2 (N827, N825, N156);
or OR4 (N828, N827, N474, N309, N171);
nor NOR4 (N829, N803, N372, N316, N64);
not NOT1 (N830, N823);
buf BUF1 (N831, N828);
buf BUF1 (N832, N830);
and AND4 (N833, N817, N581, N28, N225);
nor NOR3 (N834, N831, N181, N32);
xor XOR2 (N835, N829, N748);
xor XOR2 (N836, N834, N28);
and AND2 (N837, N826, N736);
xor XOR2 (N838, N835, N432);
nand NAND2 (N839, N832, N419);
nor NOR4 (N840, N838, N111, N178, N375);
and AND2 (N841, N824, N662);
and AND3 (N842, N814, N19, N588);
xor XOR2 (N843, N842, N342);
nand NAND2 (N844, N818, N475);
and AND3 (N845, N837, N192, N401);
or OR3 (N846, N816, N546, N128);
or OR3 (N847, N846, N393, N708);
not NOT1 (N848, N843);
nand NAND2 (N849, N840, N845);
xor XOR2 (N850, N592, N804);
xor XOR2 (N851, N850, N647);
and AND4 (N852, N822, N468, N790, N368);
not NOT1 (N853, N833);
and AND4 (N854, N852, N664, N63, N296);
and AND2 (N855, N851, N145);
or OR4 (N856, N844, N119, N117, N741);
or OR3 (N857, N847, N621, N614);
nand NAND2 (N858, N857, N598);
and AND3 (N859, N849, N737, N251);
xor XOR2 (N860, N854, N252);
not NOT1 (N861, N841);
nor NOR4 (N862, N848, N571, N410, N696);
or OR3 (N863, N855, N621, N373);
or OR2 (N864, N861, N187);
nand NAND3 (N865, N839, N759, N321);
xor XOR2 (N866, N836, N500);
buf BUF1 (N867, N864);
nand NAND2 (N868, N859, N783);
xor XOR2 (N869, N862, N490);
nand NAND3 (N870, N860, N638, N356);
or OR3 (N871, N869, N404, N484);
buf BUF1 (N872, N871);
nand NAND4 (N873, N863, N278, N607, N31);
buf BUF1 (N874, N870);
xor XOR2 (N875, N867, N577);
not NOT1 (N876, N858);
nand NAND3 (N877, N853, N274, N621);
or OR3 (N878, N868, N238, N147);
xor XOR2 (N879, N876, N132);
nor NOR2 (N880, N875, N763);
and AND3 (N881, N866, N611, N269);
not NOT1 (N882, N856);
xor XOR2 (N883, N879, N446);
or OR3 (N884, N883, N576, N491);
buf BUF1 (N885, N881);
or OR4 (N886, N882, N716, N743, N350);
or OR4 (N887, N886, N479, N571, N464);
buf BUF1 (N888, N884);
nand NAND2 (N889, N888, N25);
xor XOR2 (N890, N877, N786);
buf BUF1 (N891, N889);
not NOT1 (N892, N872);
not NOT1 (N893, N887);
xor XOR2 (N894, N885, N42);
nand NAND4 (N895, N894, N536, N516, N247);
or OR3 (N896, N880, N458, N166);
or OR4 (N897, N874, N547, N2, N709);
nand NAND4 (N898, N892, N536, N524, N425);
buf BUF1 (N899, N893);
and AND2 (N900, N890, N887);
nor NOR2 (N901, N900, N293);
xor XOR2 (N902, N865, N271);
or OR4 (N903, N895, N440, N849, N617);
and AND4 (N904, N891, N507, N772, N514);
or OR3 (N905, N902, N403, N811);
not NOT1 (N906, N873);
and AND2 (N907, N898, N762);
nor NOR4 (N908, N897, N701, N174, N791);
xor XOR2 (N909, N907, N527);
and AND3 (N910, N896, N381, N289);
and AND2 (N911, N903, N227);
xor XOR2 (N912, N910, N374);
buf BUF1 (N913, N901);
nor NOR3 (N914, N912, N512, N469);
or OR4 (N915, N908, N80, N229, N32);
nor NOR2 (N916, N878, N268);
xor XOR2 (N917, N906, N28);
nand NAND2 (N918, N911, N867);
xor XOR2 (N919, N917, N595);
and AND4 (N920, N918, N536, N185, N477);
not NOT1 (N921, N913);
and AND3 (N922, N904, N336, N666);
nand NAND2 (N923, N920, N764);
xor XOR2 (N924, N909, N16);
not NOT1 (N925, N923);
buf BUF1 (N926, N916);
or OR4 (N927, N921, N63, N175, N893);
and AND4 (N928, N924, N410, N635, N279);
or OR2 (N929, N926, N313);
xor XOR2 (N930, N915, N812);
xor XOR2 (N931, N899, N863);
not NOT1 (N932, N930);
buf BUF1 (N933, N929);
nor NOR2 (N934, N925, N610);
nand NAND3 (N935, N919, N873, N620);
and AND2 (N936, N905, N20);
nor NOR4 (N937, N932, N556, N677, N547);
xor XOR2 (N938, N933, N220);
and AND2 (N939, N928, N575);
or OR3 (N940, N938, N858, N741);
or OR3 (N941, N927, N526, N865);
not NOT1 (N942, N941);
xor XOR2 (N943, N936, N871);
buf BUF1 (N944, N922);
xor XOR2 (N945, N914, N147);
nand NAND4 (N946, N942, N41, N492, N165);
nand NAND4 (N947, N931, N327, N147, N391);
nor NOR2 (N948, N940, N258);
or OR2 (N949, N934, N483);
and AND2 (N950, N946, N488);
and AND2 (N951, N948, N504);
not NOT1 (N952, N939);
buf BUF1 (N953, N944);
nand NAND4 (N954, N952, N164, N655, N72);
nand NAND2 (N955, N951, N311);
buf BUF1 (N956, N945);
or OR4 (N957, N956, N194, N219, N885);
buf BUF1 (N958, N955);
nor NOR3 (N959, N937, N52, N800);
not NOT1 (N960, N958);
nand NAND4 (N961, N935, N75, N511, N685);
nand NAND4 (N962, N961, N953, N488, N842);
or OR3 (N963, N304, N637, N207);
not NOT1 (N964, N962);
nor NOR3 (N965, N957, N956, N500);
nor NOR2 (N966, N943, N498);
nand NAND2 (N967, N959, N584);
nor NOR3 (N968, N967, N712, N660);
or OR4 (N969, N964, N63, N331, N586);
buf BUF1 (N970, N949);
or OR2 (N971, N969, N553);
nand NAND4 (N972, N971, N450, N396, N717);
xor XOR2 (N973, N960, N605);
buf BUF1 (N974, N954);
buf BUF1 (N975, N966);
buf BUF1 (N976, N947);
nand NAND2 (N977, N963, N64);
not NOT1 (N978, N975);
and AND4 (N979, N965, N847, N595, N969);
xor XOR2 (N980, N972, N753);
buf BUF1 (N981, N970);
nand NAND3 (N982, N977, N302, N241);
nor NOR4 (N983, N979, N529, N921, N638);
buf BUF1 (N984, N981);
nor NOR3 (N985, N982, N340, N138);
nand NAND4 (N986, N980, N832, N61, N247);
nor NOR2 (N987, N950, N64);
nor NOR2 (N988, N984, N464);
not NOT1 (N989, N968);
or OR4 (N990, N986, N765, N772, N870);
xor XOR2 (N991, N976, N875);
buf BUF1 (N992, N974);
nand NAND4 (N993, N985, N397, N561, N381);
xor XOR2 (N994, N989, N47);
and AND4 (N995, N978, N407, N153, N864);
or OR3 (N996, N987, N382, N947);
nor NOR2 (N997, N994, N470);
not NOT1 (N998, N996);
and AND2 (N999, N973, N921);
buf BUF1 (N1000, N998);
and AND2 (N1001, N992, N992);
nand NAND4 (N1002, N995, N185, N299, N508);
buf BUF1 (N1003, N1001);
nand NAND2 (N1004, N993, N871);
xor XOR2 (N1005, N991, N145);
nand NAND4 (N1006, N1002, N828, N843, N966);
not NOT1 (N1007, N1005);
nor NOR3 (N1008, N990, N313, N296);
or OR4 (N1009, N997, N637, N466, N502);
nand NAND2 (N1010, N983, N748);
buf BUF1 (N1011, N1010);
not NOT1 (N1012, N1011);
buf BUF1 (N1013, N1006);
or OR3 (N1014, N1000, N58, N319);
xor XOR2 (N1015, N1009, N908);
buf BUF1 (N1016, N1013);
and AND4 (N1017, N1003, N261, N549, N185);
nor NOR4 (N1018, N999, N740, N997, N564);
xor XOR2 (N1019, N1017, N972);
xor XOR2 (N1020, N1007, N306);
xor XOR2 (N1021, N1008, N440);
and AND2 (N1022, N1004, N731);
xor XOR2 (N1023, N1012, N339);
not NOT1 (N1024, N1014);
nand NAND4 (N1025, N988, N582, N372, N655);
nand NAND3 (N1026, N1023, N525, N380);
nor NOR4 (N1027, N1015, N71, N1018, N53);
nor NOR3 (N1028, N1006, N903, N678);
buf BUF1 (N1029, N1026);
not NOT1 (N1030, N1024);
and AND2 (N1031, N1029, N400);
nand NAND3 (N1032, N1030, N378, N1030);
buf BUF1 (N1033, N1025);
buf BUF1 (N1034, N1020);
not NOT1 (N1035, N1019);
buf BUF1 (N1036, N1035);
nor NOR2 (N1037, N1036, N891);
xor XOR2 (N1038, N1028, N918);
nor NOR2 (N1039, N1022, N543);
nand NAND4 (N1040, N1039, N871, N573, N346);
buf BUF1 (N1041, N1034);
nand NAND3 (N1042, N1041, N267, N69);
nand NAND4 (N1043, N1016, N1021, N425, N226);
xor XOR2 (N1044, N693, N961);
or OR4 (N1045, N1042, N880, N586, N507);
xor XOR2 (N1046, N1033, N250);
xor XOR2 (N1047, N1044, N669);
or OR3 (N1048, N1046, N599, N236);
not NOT1 (N1049, N1038);
or OR4 (N1050, N1047, N458, N628, N406);
not NOT1 (N1051, N1045);
nand NAND3 (N1052, N1032, N142, N365);
not NOT1 (N1053, N1031);
not NOT1 (N1054, N1053);
buf BUF1 (N1055, N1043);
nand NAND2 (N1056, N1055, N557);
or OR2 (N1057, N1048, N150);
or OR4 (N1058, N1049, N157, N581, N706);
not NOT1 (N1059, N1054);
buf BUF1 (N1060, N1058);
or OR2 (N1061, N1027, N706);
and AND3 (N1062, N1037, N433, N670);
not NOT1 (N1063, N1060);
not NOT1 (N1064, N1059);
buf BUF1 (N1065, N1051);
nor NOR3 (N1066, N1040, N785, N941);
and AND4 (N1067, N1050, N255, N202, N646);
not NOT1 (N1068, N1066);
buf BUF1 (N1069, N1056);
buf BUF1 (N1070, N1052);
nand NAND3 (N1071, N1057, N1045, N985);
or OR2 (N1072, N1062, N116);
and AND2 (N1073, N1072, N406);
not NOT1 (N1074, N1063);
nor NOR4 (N1075, N1067, N634, N610, N106);
nor NOR2 (N1076, N1075, N468);
and AND4 (N1077, N1073, N163, N506, N477);
nor NOR2 (N1078, N1076, N557);
buf BUF1 (N1079, N1065);
not NOT1 (N1080, N1068);
or OR4 (N1081, N1074, N1072, N448, N1035);
and AND3 (N1082, N1061, N865, N271);
not NOT1 (N1083, N1078);
nand NAND2 (N1084, N1083, N204);
not NOT1 (N1085, N1070);
nor NOR4 (N1086, N1077, N956, N1020, N264);
nor NOR4 (N1087, N1064, N637, N671, N338);
and AND2 (N1088, N1082, N1042);
buf BUF1 (N1089, N1086);
not NOT1 (N1090, N1081);
xor XOR2 (N1091, N1089, N45);
and AND4 (N1092, N1071, N591, N58, N328);
buf BUF1 (N1093, N1080);
nor NOR2 (N1094, N1092, N177);
buf BUF1 (N1095, N1087);
xor XOR2 (N1096, N1094, N604);
xor XOR2 (N1097, N1090, N403);
nand NAND4 (N1098, N1088, N236, N277, N278);
and AND4 (N1099, N1093, N554, N839, N550);
nand NAND2 (N1100, N1095, N50);
and AND2 (N1101, N1099, N977);
and AND4 (N1102, N1079, N1011, N879, N1079);
xor XOR2 (N1103, N1098, N248);
nor NOR3 (N1104, N1069, N358, N149);
nor NOR2 (N1105, N1085, N372);
or OR2 (N1106, N1100, N931);
nor NOR4 (N1107, N1104, N668, N197, N919);
not NOT1 (N1108, N1102);
xor XOR2 (N1109, N1106, N238);
not NOT1 (N1110, N1084);
xor XOR2 (N1111, N1091, N275);
nand NAND4 (N1112, N1109, N308, N809, N208);
not NOT1 (N1113, N1097);
xor XOR2 (N1114, N1110, N1068);
buf BUF1 (N1115, N1108);
xor XOR2 (N1116, N1115, N722);
buf BUF1 (N1117, N1105);
buf BUF1 (N1118, N1111);
not NOT1 (N1119, N1112);
xor XOR2 (N1120, N1117, N820);
and AND4 (N1121, N1120, N528, N1015, N971);
not NOT1 (N1122, N1116);
buf BUF1 (N1123, N1118);
or OR3 (N1124, N1096, N1020, N429);
xor XOR2 (N1125, N1122, N917);
not NOT1 (N1126, N1121);
xor XOR2 (N1127, N1103, N766);
and AND2 (N1128, N1125, N1007);
nand NAND4 (N1129, N1113, N1078, N921, N949);
not NOT1 (N1130, N1123);
buf BUF1 (N1131, N1119);
nor NOR3 (N1132, N1126, N924, N932);
buf BUF1 (N1133, N1107);
xor XOR2 (N1134, N1132, N628);
or OR4 (N1135, N1131, N158, N12, N768);
or OR2 (N1136, N1128, N1088);
not NOT1 (N1137, N1124);
xor XOR2 (N1138, N1134, N133);
xor XOR2 (N1139, N1127, N825);
nand NAND4 (N1140, N1114, N136, N363, N814);
nor NOR4 (N1141, N1133, N458, N669, N858);
nor NOR3 (N1142, N1135, N406, N541);
nor NOR4 (N1143, N1137, N25, N30, N611);
not NOT1 (N1144, N1130);
nand NAND2 (N1145, N1141, N833);
or OR4 (N1146, N1143, N312, N840, N356);
nor NOR2 (N1147, N1136, N396);
not NOT1 (N1148, N1145);
nand NAND4 (N1149, N1146, N1100, N788, N859);
and AND3 (N1150, N1147, N963, N1145);
not NOT1 (N1151, N1129);
and AND4 (N1152, N1144, N155, N1041, N394);
not NOT1 (N1153, N1150);
xor XOR2 (N1154, N1149, N153);
nor NOR4 (N1155, N1151, N478, N27, N928);
or OR4 (N1156, N1153, N663, N203, N905);
nand NAND4 (N1157, N1154, N840, N350, N361);
nand NAND3 (N1158, N1152, N388, N507);
xor XOR2 (N1159, N1148, N996);
nand NAND2 (N1160, N1142, N425);
not NOT1 (N1161, N1155);
xor XOR2 (N1162, N1140, N49);
xor XOR2 (N1163, N1157, N975);
and AND3 (N1164, N1101, N602, N1056);
nand NAND4 (N1165, N1158, N775, N638, N1064);
xor XOR2 (N1166, N1165, N377);
xor XOR2 (N1167, N1138, N1073);
and AND2 (N1168, N1159, N146);
nand NAND4 (N1169, N1156, N58, N522, N247);
and AND3 (N1170, N1163, N369, N471);
or OR4 (N1171, N1170, N1114, N768, N221);
not NOT1 (N1172, N1171);
buf BUF1 (N1173, N1172);
not NOT1 (N1174, N1164);
xor XOR2 (N1175, N1169, N699);
and AND3 (N1176, N1167, N6, N453);
not NOT1 (N1177, N1166);
xor XOR2 (N1178, N1177, N94);
nor NOR2 (N1179, N1175, N666);
nor NOR3 (N1180, N1162, N308, N21);
buf BUF1 (N1181, N1179);
xor XOR2 (N1182, N1180, N216);
nor NOR4 (N1183, N1139, N942, N202, N892);
nand NAND3 (N1184, N1174, N475, N1149);
or OR2 (N1185, N1168, N42);
not NOT1 (N1186, N1183);
buf BUF1 (N1187, N1178);
nor NOR4 (N1188, N1176, N190, N297, N496);
not NOT1 (N1189, N1188);
buf BUF1 (N1190, N1182);
or OR3 (N1191, N1190, N960, N374);
nand NAND4 (N1192, N1173, N1189, N228, N1086);
and AND4 (N1193, N67, N755, N278, N695);
not NOT1 (N1194, N1187);
and AND4 (N1195, N1194, N136, N942, N1103);
nand NAND2 (N1196, N1193, N826);
nand NAND2 (N1197, N1160, N155);
or OR3 (N1198, N1186, N619, N888);
nor NOR2 (N1199, N1195, N382);
xor XOR2 (N1200, N1196, N358);
nor NOR3 (N1201, N1185, N359, N1096);
buf BUF1 (N1202, N1197);
buf BUF1 (N1203, N1200);
or OR3 (N1204, N1184, N786, N385);
xor XOR2 (N1205, N1192, N617);
nand NAND4 (N1206, N1205, N446, N1066, N576);
not NOT1 (N1207, N1202);
not NOT1 (N1208, N1201);
not NOT1 (N1209, N1206);
buf BUF1 (N1210, N1209);
or OR2 (N1211, N1199, N1123);
and AND2 (N1212, N1161, N465);
xor XOR2 (N1213, N1207, N565);
not NOT1 (N1214, N1191);
and AND3 (N1215, N1213, N1177, N373);
not NOT1 (N1216, N1214);
nor NOR2 (N1217, N1216, N802);
or OR2 (N1218, N1212, N761);
nor NOR3 (N1219, N1181, N463, N536);
buf BUF1 (N1220, N1211);
nor NOR3 (N1221, N1204, N692, N167);
or OR2 (N1222, N1220, N746);
and AND4 (N1223, N1221, N889, N715, N637);
buf BUF1 (N1224, N1198);
and AND2 (N1225, N1224, N783);
nand NAND4 (N1226, N1225, N555, N789, N570);
or OR2 (N1227, N1210, N313);
nor NOR4 (N1228, N1223, N320, N481, N1057);
and AND4 (N1229, N1226, N266, N795, N1143);
buf BUF1 (N1230, N1222);
and AND4 (N1231, N1215, N353, N637, N602);
not NOT1 (N1232, N1227);
not NOT1 (N1233, N1229);
and AND4 (N1234, N1219, N975, N93, N1133);
nor NOR3 (N1235, N1233, N643, N896);
or OR3 (N1236, N1230, N764, N1235);
nand NAND3 (N1237, N1092, N1184, N347);
and AND4 (N1238, N1217, N454, N832, N570);
or OR3 (N1239, N1236, N221, N1164);
nor NOR3 (N1240, N1234, N61, N1054);
and AND2 (N1241, N1203, N259);
not NOT1 (N1242, N1240);
xor XOR2 (N1243, N1208, N94);
nand NAND3 (N1244, N1232, N1088, N1171);
nor NOR4 (N1245, N1231, N1084, N1170, N735);
nor NOR2 (N1246, N1218, N1070);
or OR3 (N1247, N1238, N870, N432);
not NOT1 (N1248, N1245);
and AND4 (N1249, N1237, N36, N965, N783);
nor NOR2 (N1250, N1239, N21);
nand NAND4 (N1251, N1228, N858, N764, N1076);
or OR4 (N1252, N1242, N694, N185, N1119);
or OR2 (N1253, N1243, N861);
xor XOR2 (N1254, N1253, N1098);
not NOT1 (N1255, N1252);
and AND4 (N1256, N1254, N926, N1043, N391);
or OR4 (N1257, N1255, N202, N654, N25);
buf BUF1 (N1258, N1248);
buf BUF1 (N1259, N1244);
or OR4 (N1260, N1256, N581, N611, N551);
nor NOR2 (N1261, N1241, N216);
or OR2 (N1262, N1249, N1186);
and AND3 (N1263, N1258, N409, N833);
buf BUF1 (N1264, N1246);
not NOT1 (N1265, N1262);
nor NOR4 (N1266, N1259, N380, N399, N864);
xor XOR2 (N1267, N1251, N493);
nand NAND3 (N1268, N1267, N1159, N790);
not NOT1 (N1269, N1247);
nor NOR2 (N1270, N1263, N623);
nand NAND3 (N1271, N1261, N439, N1019);
nand NAND2 (N1272, N1269, N725);
not NOT1 (N1273, N1250);
nand NAND3 (N1274, N1272, N357, N218);
buf BUF1 (N1275, N1271);
nand NAND2 (N1276, N1275, N730);
and AND3 (N1277, N1266, N577, N777);
buf BUF1 (N1278, N1276);
or OR3 (N1279, N1264, N175, N1180);
nand NAND2 (N1280, N1265, N977);
xor XOR2 (N1281, N1268, N1052);
nand NAND4 (N1282, N1274, N1145, N296, N1022);
xor XOR2 (N1283, N1278, N637);
or OR2 (N1284, N1280, N536);
xor XOR2 (N1285, N1284, N972);
xor XOR2 (N1286, N1257, N855);
or OR3 (N1287, N1281, N908, N646);
or OR3 (N1288, N1285, N241, N1013);
nand NAND4 (N1289, N1287, N620, N287, N1039);
buf BUF1 (N1290, N1288);
nand NAND3 (N1291, N1273, N205, N1003);
not NOT1 (N1292, N1270);
buf BUF1 (N1293, N1283);
not NOT1 (N1294, N1282);
nand NAND2 (N1295, N1294, N961);
buf BUF1 (N1296, N1279);
buf BUF1 (N1297, N1286);
nor NOR2 (N1298, N1289, N403);
nand NAND3 (N1299, N1277, N1234, N1195);
nand NAND3 (N1300, N1296, N392, N490);
nand NAND2 (N1301, N1300, N829);
and AND2 (N1302, N1297, N756);
or OR2 (N1303, N1293, N1045);
nand NAND2 (N1304, N1299, N1225);
nand NAND3 (N1305, N1292, N468, N529);
nand NAND3 (N1306, N1298, N298, N1112);
nor NOR4 (N1307, N1290, N919, N1067, N1020);
nand NAND2 (N1308, N1302, N684);
xor XOR2 (N1309, N1304, N574);
nor NOR2 (N1310, N1307, N658);
buf BUF1 (N1311, N1295);
nand NAND2 (N1312, N1303, N74);
nand NAND3 (N1313, N1312, N856, N230);
nand NAND2 (N1314, N1309, N397);
buf BUF1 (N1315, N1314);
and AND4 (N1316, N1310, N929, N611, N72);
and AND4 (N1317, N1301, N275, N971, N221);
not NOT1 (N1318, N1308);
buf BUF1 (N1319, N1305);
nand NAND4 (N1320, N1319, N173, N488, N849);
not NOT1 (N1321, N1320);
nor NOR3 (N1322, N1317, N364, N1103);
buf BUF1 (N1323, N1318);
or OR3 (N1324, N1260, N189, N526);
nor NOR2 (N1325, N1315, N434);
and AND3 (N1326, N1311, N1318, N416);
nand NAND4 (N1327, N1291, N66, N854, N1249);
or OR2 (N1328, N1323, N35);
buf BUF1 (N1329, N1328);
not NOT1 (N1330, N1313);
xor XOR2 (N1331, N1326, N179);
nor NOR2 (N1332, N1316, N49);
buf BUF1 (N1333, N1321);
nor NOR3 (N1334, N1329, N376, N648);
and AND2 (N1335, N1332, N439);
xor XOR2 (N1336, N1334, N1067);
xor XOR2 (N1337, N1324, N470);
nand NAND4 (N1338, N1325, N527, N539, N1189);
nor NOR4 (N1339, N1330, N295, N260, N381);
not NOT1 (N1340, N1336);
and AND2 (N1341, N1335, N569);
nor NOR4 (N1342, N1331, N1324, N207, N41);
and AND4 (N1343, N1322, N173, N157, N513);
not NOT1 (N1344, N1339);
nor NOR3 (N1345, N1333, N745, N323);
or OR2 (N1346, N1327, N1082);
nand NAND2 (N1347, N1342, N529);
nor NOR2 (N1348, N1337, N251);
nor NOR4 (N1349, N1341, N1082, N427, N999);
buf BUF1 (N1350, N1340);
and AND3 (N1351, N1306, N57, N103);
nand NAND3 (N1352, N1350, N918, N509);
xor XOR2 (N1353, N1345, N929);
buf BUF1 (N1354, N1348);
buf BUF1 (N1355, N1338);
xor XOR2 (N1356, N1352, N775);
nor NOR4 (N1357, N1354, N38, N529, N566);
nor NOR2 (N1358, N1356, N469);
nor NOR3 (N1359, N1358, N780, N749);
not NOT1 (N1360, N1357);
nand NAND3 (N1361, N1355, N690, N1154);
buf BUF1 (N1362, N1346);
or OR3 (N1363, N1360, N852, N255);
or OR4 (N1364, N1359, N264, N479, N289);
not NOT1 (N1365, N1364);
buf BUF1 (N1366, N1347);
and AND4 (N1367, N1353, N179, N1182, N401);
nor NOR3 (N1368, N1362, N788, N636);
nor NOR3 (N1369, N1361, N627, N278);
and AND2 (N1370, N1343, N621);
nand NAND4 (N1371, N1370, N559, N1035, N16);
not NOT1 (N1372, N1365);
xor XOR2 (N1373, N1351, N51);
not NOT1 (N1374, N1367);
not NOT1 (N1375, N1374);
not NOT1 (N1376, N1369);
nand NAND3 (N1377, N1373, N1321, N1148);
nor NOR4 (N1378, N1377, N247, N88, N730);
buf BUF1 (N1379, N1371);
xor XOR2 (N1380, N1372, N760);
xor XOR2 (N1381, N1368, N509);
not NOT1 (N1382, N1366);
nor NOR2 (N1383, N1363, N928);
not NOT1 (N1384, N1381);
xor XOR2 (N1385, N1375, N624);
not NOT1 (N1386, N1378);
and AND3 (N1387, N1384, N1110, N733);
buf BUF1 (N1388, N1380);
nor NOR2 (N1389, N1385, N832);
and AND4 (N1390, N1388, N246, N668, N360);
xor XOR2 (N1391, N1344, N400);
nor NOR2 (N1392, N1349, N614);
xor XOR2 (N1393, N1387, N826);
or OR3 (N1394, N1392, N467, N557);
and AND4 (N1395, N1383, N1082, N1164, N942);
xor XOR2 (N1396, N1390, N552);
or OR2 (N1397, N1395, N227);
and AND4 (N1398, N1394, N1348, N842, N204);
nor NOR2 (N1399, N1393, N1023);
buf BUF1 (N1400, N1382);
nand NAND3 (N1401, N1391, N1000, N219);
xor XOR2 (N1402, N1376, N984);
and AND3 (N1403, N1401, N1318, N732);
xor XOR2 (N1404, N1389, N343);
buf BUF1 (N1405, N1386);
xor XOR2 (N1406, N1404, N1284);
not NOT1 (N1407, N1400);
buf BUF1 (N1408, N1398);
buf BUF1 (N1409, N1397);
buf BUF1 (N1410, N1396);
xor XOR2 (N1411, N1409, N569);
or OR4 (N1412, N1407, N755, N559, N509);
nand NAND3 (N1413, N1408, N430, N1185);
or OR3 (N1414, N1412, N1286, N522);
buf BUF1 (N1415, N1414);
buf BUF1 (N1416, N1405);
not NOT1 (N1417, N1379);
xor XOR2 (N1418, N1413, N930);
xor XOR2 (N1419, N1410, N1321);
and AND2 (N1420, N1411, N620);
not NOT1 (N1421, N1417);
buf BUF1 (N1422, N1402);
or OR4 (N1423, N1418, N824, N436, N831);
xor XOR2 (N1424, N1419, N146);
xor XOR2 (N1425, N1406, N1037);
and AND4 (N1426, N1421, N1033, N1135, N604);
buf BUF1 (N1427, N1420);
and AND2 (N1428, N1423, N557);
nor NOR4 (N1429, N1426, N1161, N70, N1091);
or OR4 (N1430, N1424, N1243, N542, N530);
and AND2 (N1431, N1416, N1251);
nand NAND4 (N1432, N1427, N502, N89, N983);
xor XOR2 (N1433, N1432, N895);
and AND2 (N1434, N1422, N100);
nor NOR4 (N1435, N1399, N545, N479, N1102);
not NOT1 (N1436, N1425);
nor NOR2 (N1437, N1415, N854);
xor XOR2 (N1438, N1434, N791);
not NOT1 (N1439, N1428);
nand NAND2 (N1440, N1435, N106);
xor XOR2 (N1441, N1433, N179);
xor XOR2 (N1442, N1439, N320);
nand NAND2 (N1443, N1430, N99);
not NOT1 (N1444, N1442);
xor XOR2 (N1445, N1429, N1043);
and AND2 (N1446, N1445, N1140);
xor XOR2 (N1447, N1441, N1401);
and AND2 (N1448, N1437, N1149);
not NOT1 (N1449, N1431);
xor XOR2 (N1450, N1403, N714);
buf BUF1 (N1451, N1438);
not NOT1 (N1452, N1440);
or OR2 (N1453, N1451, N1081);
buf BUF1 (N1454, N1448);
or OR4 (N1455, N1453, N808, N857, N1082);
buf BUF1 (N1456, N1446);
nand NAND4 (N1457, N1452, N752, N191, N964);
not NOT1 (N1458, N1436);
nand NAND3 (N1459, N1458, N498, N865);
buf BUF1 (N1460, N1443);
buf BUF1 (N1461, N1447);
not NOT1 (N1462, N1457);
and AND4 (N1463, N1461, N1320, N510, N597);
or OR4 (N1464, N1450, N1073, N1099, N1203);
buf BUF1 (N1465, N1444);
nand NAND4 (N1466, N1454, N369, N928, N775);
nand NAND3 (N1467, N1459, N96, N498);
nand NAND3 (N1468, N1467, N1459, N685);
xor XOR2 (N1469, N1464, N1375);
nand NAND3 (N1470, N1460, N137, N981);
xor XOR2 (N1471, N1470, N981);
xor XOR2 (N1472, N1463, N175);
and AND4 (N1473, N1472, N1288, N672, N1391);
and AND3 (N1474, N1456, N1320, N1054);
nor NOR3 (N1475, N1462, N570, N1266);
not NOT1 (N1476, N1471);
and AND4 (N1477, N1474, N294, N1346, N748);
xor XOR2 (N1478, N1465, N648);
and AND2 (N1479, N1469, N1459);
nand NAND2 (N1480, N1475, N392);
or OR2 (N1481, N1455, N1278);
and AND4 (N1482, N1466, N1063, N734, N1281);
not NOT1 (N1483, N1476);
nor NOR3 (N1484, N1483, N1249, N867);
xor XOR2 (N1485, N1480, N783);
xor XOR2 (N1486, N1478, N352);
not NOT1 (N1487, N1468);
nor NOR4 (N1488, N1473, N775, N158, N984);
or OR4 (N1489, N1481, N368, N893, N1294);
xor XOR2 (N1490, N1486, N1296);
and AND4 (N1491, N1489, N1349, N82, N1137);
nand NAND3 (N1492, N1482, N436, N630);
or OR2 (N1493, N1491, N1168);
nand NAND2 (N1494, N1488, N1117);
xor XOR2 (N1495, N1449, N407);
or OR2 (N1496, N1479, N1394);
or OR4 (N1497, N1496, N541, N318, N1066);
and AND2 (N1498, N1487, N1067);
not NOT1 (N1499, N1498);
or OR4 (N1500, N1495, N103, N254, N656);
nor NOR4 (N1501, N1493, N433, N758, N735);
not NOT1 (N1502, N1497);
nand NAND4 (N1503, N1485, N451, N1413, N134);
xor XOR2 (N1504, N1484, N1089);
not NOT1 (N1505, N1477);
nand NAND3 (N1506, N1500, N687, N297);
buf BUF1 (N1507, N1502);
nor NOR4 (N1508, N1506, N879, N1071, N33);
nand NAND3 (N1509, N1505, N926, N1093);
or OR3 (N1510, N1490, N1019, N928);
not NOT1 (N1511, N1501);
and AND2 (N1512, N1507, N512);
nor NOR3 (N1513, N1504, N1076, N695);
xor XOR2 (N1514, N1494, N886);
and AND2 (N1515, N1514, N716);
or OR3 (N1516, N1515, N896, N606);
nor NOR3 (N1517, N1499, N247, N269);
and AND4 (N1518, N1511, N142, N1474, N1090);
nand NAND2 (N1519, N1509, N106);
not NOT1 (N1520, N1513);
and AND2 (N1521, N1518, N50);
nor NOR4 (N1522, N1521, N543, N561, N1090);
nand NAND4 (N1523, N1516, N68, N408, N1153);
or OR4 (N1524, N1520, N1178, N819, N19);
or OR3 (N1525, N1523, N721, N797);
not NOT1 (N1526, N1525);
and AND2 (N1527, N1508, N1163);
nor NOR4 (N1528, N1522, N946, N608, N477);
xor XOR2 (N1529, N1517, N523);
or OR4 (N1530, N1524, N1263, N178, N1140);
or OR2 (N1531, N1492, N423);
xor XOR2 (N1532, N1503, N445);
nand NAND3 (N1533, N1531, N1454, N1296);
or OR3 (N1534, N1528, N794, N1143);
xor XOR2 (N1535, N1533, N1520);
buf BUF1 (N1536, N1527);
and AND4 (N1537, N1534, N664, N1499, N1134);
buf BUF1 (N1538, N1510);
xor XOR2 (N1539, N1530, N9);
or OR3 (N1540, N1538, N952, N971);
nand NAND3 (N1541, N1529, N768, N1438);
xor XOR2 (N1542, N1526, N1321);
and AND3 (N1543, N1537, N1444, N1449);
or OR4 (N1544, N1542, N1142, N1261, N438);
xor XOR2 (N1545, N1532, N445);
or OR4 (N1546, N1544, N891, N651, N1408);
not NOT1 (N1547, N1519);
buf BUF1 (N1548, N1543);
or OR4 (N1549, N1548, N1087, N1181, N568);
not NOT1 (N1550, N1536);
not NOT1 (N1551, N1546);
not NOT1 (N1552, N1551);
buf BUF1 (N1553, N1545);
buf BUF1 (N1554, N1540);
or OR2 (N1555, N1552, N1382);
nand NAND2 (N1556, N1554, N1215);
xor XOR2 (N1557, N1539, N448);
nor NOR3 (N1558, N1556, N1167, N690);
and AND4 (N1559, N1555, N794, N775, N1039);
nor NOR4 (N1560, N1541, N451, N258, N1455);
nor NOR2 (N1561, N1512, N751);
nor NOR4 (N1562, N1558, N660, N1411, N122);
not NOT1 (N1563, N1535);
not NOT1 (N1564, N1557);
or OR3 (N1565, N1563, N1479, N825);
or OR4 (N1566, N1562, N233, N928, N1400);
nor NOR4 (N1567, N1553, N1146, N1107, N40);
not NOT1 (N1568, N1559);
nor NOR4 (N1569, N1550, N851, N901, N597);
nor NOR2 (N1570, N1560, N650);
nor NOR3 (N1571, N1564, N1218, N97);
nand NAND3 (N1572, N1547, N1290, N1416);
nor NOR4 (N1573, N1572, N1139, N987, N392);
nand NAND3 (N1574, N1566, N1518, N1301);
buf BUF1 (N1575, N1573);
nor NOR3 (N1576, N1575, N220, N752);
buf BUF1 (N1577, N1571);
nand NAND4 (N1578, N1569, N1073, N320, N419);
nor NOR4 (N1579, N1549, N163, N1468, N792);
and AND2 (N1580, N1567, N579);
and AND2 (N1581, N1578, N1028);
nor NOR4 (N1582, N1579, N1339, N879, N1326);
nand NAND4 (N1583, N1577, N704, N859, N1157);
and AND2 (N1584, N1568, N379);
xor XOR2 (N1585, N1584, N856);
xor XOR2 (N1586, N1580, N310);
or OR2 (N1587, N1561, N1510);
xor XOR2 (N1588, N1587, N708);
xor XOR2 (N1589, N1574, N1445);
xor XOR2 (N1590, N1583, N1265);
buf BUF1 (N1591, N1576);
not NOT1 (N1592, N1581);
or OR4 (N1593, N1570, N356, N121, N73);
or OR3 (N1594, N1588, N176, N1193);
nand NAND2 (N1595, N1582, N1245);
not NOT1 (N1596, N1585);
or OR3 (N1597, N1593, N753, N960);
nor NOR4 (N1598, N1592, N571, N1519, N1037);
or OR2 (N1599, N1591, N1420);
or OR3 (N1600, N1590, N1111, N9);
and AND3 (N1601, N1586, N23, N1216);
and AND4 (N1602, N1589, N125, N1134, N1024);
and AND4 (N1603, N1602, N740, N728, N390);
and AND3 (N1604, N1603, N952, N1154);
nand NAND2 (N1605, N1595, N1366);
and AND3 (N1606, N1596, N63, N1368);
nand NAND2 (N1607, N1604, N701);
not NOT1 (N1608, N1594);
nor NOR3 (N1609, N1600, N101, N1267);
buf BUF1 (N1610, N1565);
and AND4 (N1611, N1605, N682, N69, N72);
buf BUF1 (N1612, N1608);
or OR2 (N1613, N1601, N1480);
nor NOR3 (N1614, N1597, N1203, N878);
nor NOR3 (N1615, N1612, N304, N668);
nor NOR4 (N1616, N1614, N638, N556, N1162);
or OR3 (N1617, N1598, N914, N1583);
nor NOR3 (N1618, N1616, N1003, N1256);
buf BUF1 (N1619, N1615);
and AND3 (N1620, N1611, N1076, N757);
buf BUF1 (N1621, N1617);
xor XOR2 (N1622, N1618, N1565);
xor XOR2 (N1623, N1609, N1322);
not NOT1 (N1624, N1622);
not NOT1 (N1625, N1621);
nand NAND4 (N1626, N1607, N959, N670, N410);
not NOT1 (N1627, N1620);
or OR4 (N1628, N1623, N1156, N377, N926);
nand NAND3 (N1629, N1613, N1073, N1365);
xor XOR2 (N1630, N1629, N513);
nand NAND3 (N1631, N1610, N463, N1069);
buf BUF1 (N1632, N1619);
buf BUF1 (N1633, N1632);
or OR2 (N1634, N1599, N491);
nand NAND3 (N1635, N1633, N995, N308);
nand NAND4 (N1636, N1626, N1545, N1355, N358);
nor NOR3 (N1637, N1625, N1498, N708);
buf BUF1 (N1638, N1635);
or OR3 (N1639, N1627, N690, N1176);
nand NAND4 (N1640, N1634, N831, N925, N766);
xor XOR2 (N1641, N1631, N1053);
nand NAND4 (N1642, N1641, N1355, N1404, N1144);
nand NAND2 (N1643, N1637, N800);
nor NOR2 (N1644, N1640, N968);
or OR4 (N1645, N1636, N781, N116, N1351);
or OR3 (N1646, N1639, N1584, N1472);
nor NOR4 (N1647, N1624, N585, N287, N1008);
or OR4 (N1648, N1642, N1252, N1504, N731);
not NOT1 (N1649, N1645);
xor XOR2 (N1650, N1647, N1434);
xor XOR2 (N1651, N1649, N713);
and AND4 (N1652, N1648, N1041, N1241, N348);
or OR4 (N1653, N1650, N988, N1503, N1267);
not NOT1 (N1654, N1630);
not NOT1 (N1655, N1652);
and AND3 (N1656, N1606, N487, N706);
or OR3 (N1657, N1654, N1458, N1309);
and AND2 (N1658, N1653, N534);
not NOT1 (N1659, N1655);
nand NAND2 (N1660, N1658, N1623);
nor NOR3 (N1661, N1659, N577, N1354);
xor XOR2 (N1662, N1644, N177);
nand NAND4 (N1663, N1638, N1558, N1496, N1337);
nor NOR2 (N1664, N1628, N262);
xor XOR2 (N1665, N1656, N422);
not NOT1 (N1666, N1661);
and AND4 (N1667, N1643, N256, N1318, N704);
nand NAND4 (N1668, N1665, N541, N1317, N1235);
buf BUF1 (N1669, N1663);
buf BUF1 (N1670, N1660);
xor XOR2 (N1671, N1668, N1476);
nand NAND4 (N1672, N1670, N1303, N418, N414);
or OR4 (N1673, N1671, N1573, N260, N1588);
xor XOR2 (N1674, N1657, N426);
buf BUF1 (N1675, N1672);
xor XOR2 (N1676, N1646, N94);
and AND2 (N1677, N1666, N999);
buf BUF1 (N1678, N1673);
nand NAND4 (N1679, N1678, N132, N1067, N634);
xor XOR2 (N1680, N1664, N827);
nor NOR4 (N1681, N1680, N1033, N1163, N1600);
xor XOR2 (N1682, N1667, N629);
and AND2 (N1683, N1681, N460);
not NOT1 (N1684, N1683);
nand NAND2 (N1685, N1662, N1291);
or OR3 (N1686, N1685, N604, N1369);
not NOT1 (N1687, N1684);
nand NAND3 (N1688, N1651, N1184, N571);
nand NAND2 (N1689, N1688, N1434);
nor NOR2 (N1690, N1679, N848);
xor XOR2 (N1691, N1669, N1406);
and AND4 (N1692, N1676, N1474, N1361, N392);
or OR4 (N1693, N1674, N786, N1360, N1190);
buf BUF1 (N1694, N1690);
buf BUF1 (N1695, N1691);
nand NAND4 (N1696, N1689, N789, N815, N1419);
nor NOR4 (N1697, N1695, N1273, N1576, N1528);
buf BUF1 (N1698, N1694);
not NOT1 (N1699, N1682);
xor XOR2 (N1700, N1686, N1111);
nor NOR4 (N1701, N1697, N519, N1699, N389);
nor NOR3 (N1702, N899, N1308, N458);
nand NAND4 (N1703, N1677, N1133, N90, N1076);
or OR2 (N1704, N1687, N882);
buf BUF1 (N1705, N1692);
nand NAND3 (N1706, N1675, N1197, N924);
xor XOR2 (N1707, N1698, N171);
nor NOR3 (N1708, N1702, N633, N408);
nor NOR3 (N1709, N1704, N1440, N1686);
nand NAND2 (N1710, N1701, N1485);
and AND2 (N1711, N1696, N561);
and AND3 (N1712, N1711, N1334, N702);
not NOT1 (N1713, N1705);
and AND3 (N1714, N1693, N1519, N1145);
or OR3 (N1715, N1700, N1388, N742);
xor XOR2 (N1716, N1712, N234);
not NOT1 (N1717, N1715);
xor XOR2 (N1718, N1717, N716);
not NOT1 (N1719, N1703);
xor XOR2 (N1720, N1707, N1205);
buf BUF1 (N1721, N1710);
nor NOR2 (N1722, N1721, N360);
or OR3 (N1723, N1716, N906, N48);
not NOT1 (N1724, N1723);
nand NAND3 (N1725, N1713, N808, N1146);
nand NAND4 (N1726, N1722, N1040, N91, N296);
nand NAND2 (N1727, N1726, N121);
not NOT1 (N1728, N1718);
nor NOR4 (N1729, N1709, N706, N151, N1562);
nand NAND2 (N1730, N1708, N910);
buf BUF1 (N1731, N1725);
xor XOR2 (N1732, N1720, N1199);
xor XOR2 (N1733, N1706, N1682);
buf BUF1 (N1734, N1729);
xor XOR2 (N1735, N1733, N657);
and AND3 (N1736, N1719, N1580, N8);
and AND3 (N1737, N1735, N367, N1087);
nand NAND4 (N1738, N1727, N745, N794, N1036);
nand NAND4 (N1739, N1732, N205, N1088, N1496);
and AND4 (N1740, N1728, N1605, N726, N146);
nor NOR2 (N1741, N1731, N237);
or OR3 (N1742, N1734, N863, N7);
buf BUF1 (N1743, N1739);
and AND2 (N1744, N1737, N88);
or OR4 (N1745, N1740, N1178, N167, N1567);
nor NOR3 (N1746, N1744, N1051, N300);
and AND2 (N1747, N1730, N1049);
xor XOR2 (N1748, N1742, N869);
nand NAND3 (N1749, N1724, N283, N448);
xor XOR2 (N1750, N1714, N993);
or OR2 (N1751, N1750, N95);
or OR4 (N1752, N1736, N1024, N1679, N1684);
and AND4 (N1753, N1743, N1049, N1744, N1188);
or OR3 (N1754, N1738, N538, N50);
or OR4 (N1755, N1745, N1211, N1504, N967);
not NOT1 (N1756, N1741);
buf BUF1 (N1757, N1751);
xor XOR2 (N1758, N1752, N1209);
nand NAND4 (N1759, N1756, N509, N130, N229);
and AND2 (N1760, N1759, N236);
nand NAND2 (N1761, N1755, N916);
or OR3 (N1762, N1757, N1464, N683);
nand NAND2 (N1763, N1754, N1589);
not NOT1 (N1764, N1753);
buf BUF1 (N1765, N1762);
buf BUF1 (N1766, N1763);
or OR2 (N1767, N1765, N22);
not NOT1 (N1768, N1764);
and AND2 (N1769, N1761, N1126);
or OR4 (N1770, N1758, N1679, N135, N90);
not NOT1 (N1771, N1770);
nor NOR3 (N1772, N1749, N273, N653);
xor XOR2 (N1773, N1767, N860);
not NOT1 (N1774, N1747);
buf BUF1 (N1775, N1773);
or OR4 (N1776, N1775, N1430, N1082, N238);
nor NOR3 (N1777, N1772, N436, N462);
buf BUF1 (N1778, N1776);
nor NOR4 (N1779, N1778, N615, N963, N774);
nand NAND4 (N1780, N1768, N1369, N1705, N776);
or OR2 (N1781, N1774, N621);
buf BUF1 (N1782, N1779);
not NOT1 (N1783, N1781);
and AND3 (N1784, N1769, N1589, N1420);
nand NAND2 (N1785, N1766, N759);
buf BUF1 (N1786, N1785);
and AND2 (N1787, N1786, N1625);
nor NOR3 (N1788, N1748, N868, N623);
and AND2 (N1789, N1787, N859);
or OR3 (N1790, N1783, N1480, N250);
nand NAND2 (N1791, N1784, N1653);
and AND4 (N1792, N1771, N619, N857, N1416);
or OR3 (N1793, N1791, N1518, N1586);
nor NOR3 (N1794, N1790, N1614, N650);
nor NOR4 (N1795, N1746, N1699, N995, N1414);
or OR3 (N1796, N1782, N770, N929);
not NOT1 (N1797, N1792);
xor XOR2 (N1798, N1795, N92);
and AND2 (N1799, N1797, N208);
not NOT1 (N1800, N1777);
nand NAND2 (N1801, N1794, N861);
and AND2 (N1802, N1780, N1707);
and AND4 (N1803, N1789, N1004, N1202, N407);
nor NOR2 (N1804, N1803, N697);
and AND3 (N1805, N1788, N586, N438);
and AND4 (N1806, N1804, N1276, N1144, N1359);
and AND3 (N1807, N1760, N409, N609);
not NOT1 (N1808, N1807);
not NOT1 (N1809, N1802);
and AND2 (N1810, N1801, N81);
and AND4 (N1811, N1810, N1080, N929, N1513);
and AND2 (N1812, N1806, N642);
not NOT1 (N1813, N1808);
nand NAND3 (N1814, N1798, N1650, N1163);
xor XOR2 (N1815, N1800, N970);
nor NOR3 (N1816, N1793, N743, N270);
not NOT1 (N1817, N1815);
and AND2 (N1818, N1814, N309);
not NOT1 (N1819, N1809);
and AND3 (N1820, N1799, N1028, N36);
nand NAND4 (N1821, N1813, N675, N758, N302);
xor XOR2 (N1822, N1796, N112);
xor XOR2 (N1823, N1819, N204);
not NOT1 (N1824, N1812);
and AND4 (N1825, N1818, N138, N1694, N1749);
nand NAND2 (N1826, N1822, N338);
and AND4 (N1827, N1821, N978, N731, N1225);
or OR4 (N1828, N1825, N293, N1394, N530);
or OR2 (N1829, N1823, N679);
not NOT1 (N1830, N1811);
nor NOR2 (N1831, N1830, N1161);
and AND3 (N1832, N1828, N1489, N985);
buf BUF1 (N1833, N1827);
or OR4 (N1834, N1817, N140, N816, N1142);
not NOT1 (N1835, N1816);
nor NOR3 (N1836, N1826, N1102, N574);
and AND3 (N1837, N1836, N1222, N1364);
nor NOR3 (N1838, N1837, N911, N1517);
buf BUF1 (N1839, N1838);
nor NOR3 (N1840, N1835, N1518, N334);
or OR4 (N1841, N1840, N142, N134, N1133);
not NOT1 (N1842, N1832);
buf BUF1 (N1843, N1842);
xor XOR2 (N1844, N1833, N1326);
and AND2 (N1845, N1805, N280);
nor NOR3 (N1846, N1845, N1747, N638);
xor XOR2 (N1847, N1824, N754);
buf BUF1 (N1848, N1831);
not NOT1 (N1849, N1820);
not NOT1 (N1850, N1848);
buf BUF1 (N1851, N1843);
buf BUF1 (N1852, N1846);
nand NAND2 (N1853, N1844, N1191);
nor NOR3 (N1854, N1850, N582, N694);
nor NOR4 (N1855, N1829, N98, N4, N792);
or OR4 (N1856, N1839, N1239, N1373, N241);
buf BUF1 (N1857, N1852);
buf BUF1 (N1858, N1855);
nor NOR2 (N1859, N1841, N873);
buf BUF1 (N1860, N1853);
nor NOR2 (N1861, N1854, N691);
xor XOR2 (N1862, N1861, N1284);
xor XOR2 (N1863, N1862, N538);
or OR2 (N1864, N1856, N1518);
and AND2 (N1865, N1859, N27);
and AND4 (N1866, N1858, N74, N1546, N410);
and AND2 (N1867, N1849, N1716);
not NOT1 (N1868, N1866);
or OR3 (N1869, N1864, N8, N1400);
nand NAND4 (N1870, N1863, N260, N908, N1751);
buf BUF1 (N1871, N1868);
buf BUF1 (N1872, N1860);
nor NOR3 (N1873, N1851, N1027, N28);
nor NOR4 (N1874, N1869, N791, N1385, N288);
and AND4 (N1875, N1834, N1197, N923, N1494);
nor NOR4 (N1876, N1865, N380, N1085, N119);
nor NOR3 (N1877, N1867, N1699, N1081);
xor XOR2 (N1878, N1871, N147);
nand NAND4 (N1879, N1872, N1639, N307, N1202);
or OR4 (N1880, N1873, N957, N938, N1876);
xor XOR2 (N1881, N33, N1853);
buf BUF1 (N1882, N1874);
buf BUF1 (N1883, N1879);
and AND2 (N1884, N1882, N1186);
buf BUF1 (N1885, N1857);
or OR3 (N1886, N1885, N1787, N828);
nor NOR4 (N1887, N1847, N1875, N374, N1175);
xor XOR2 (N1888, N651, N1660);
and AND3 (N1889, N1880, N1723, N1527);
nand NAND4 (N1890, N1886, N538, N1485, N383);
xor XOR2 (N1891, N1870, N881);
or OR3 (N1892, N1881, N149, N1619);
nand NAND4 (N1893, N1888, N1760, N1643, N453);
or OR4 (N1894, N1893, N1463, N1467, N1414);
buf BUF1 (N1895, N1878);
xor XOR2 (N1896, N1892, N535);
buf BUF1 (N1897, N1890);
or OR4 (N1898, N1883, N1868, N705, N461);
or OR3 (N1899, N1884, N1139, N285);
buf BUF1 (N1900, N1889);
not NOT1 (N1901, N1895);
and AND3 (N1902, N1894, N618, N1507);
not NOT1 (N1903, N1877);
nor NOR4 (N1904, N1887, N980, N1, N1029);
not NOT1 (N1905, N1899);
or OR4 (N1906, N1891, N234, N478, N37);
nor NOR3 (N1907, N1905, N310, N931);
and AND4 (N1908, N1902, N1130, N1454, N1551);
nand NAND3 (N1909, N1908, N650, N1443);
not NOT1 (N1910, N1900);
nor NOR4 (N1911, N1901, N1124, N218, N1710);
nor NOR2 (N1912, N1896, N1012);
not NOT1 (N1913, N1903);
not NOT1 (N1914, N1906);
nor NOR3 (N1915, N1911, N403, N297);
not NOT1 (N1916, N1914);
not NOT1 (N1917, N1915);
or OR4 (N1918, N1916, N982, N783, N1553);
xor XOR2 (N1919, N1904, N1368);
or OR3 (N1920, N1898, N119, N584);
not NOT1 (N1921, N1909);
buf BUF1 (N1922, N1897);
xor XOR2 (N1923, N1918, N1016);
and AND4 (N1924, N1912, N1539, N1418, N680);
and AND4 (N1925, N1924, N169, N141, N1309);
nor NOR3 (N1926, N1921, N1698, N742);
nand NAND2 (N1927, N1925, N1655);
not NOT1 (N1928, N1922);
xor XOR2 (N1929, N1927, N747);
nand NAND3 (N1930, N1929, N667, N1485);
xor XOR2 (N1931, N1917, N1398);
buf BUF1 (N1932, N1931);
nand NAND2 (N1933, N1920, N1876);
nor NOR3 (N1934, N1930, N1871, N141);
buf BUF1 (N1935, N1933);
buf BUF1 (N1936, N1932);
and AND4 (N1937, N1936, N1750, N456, N683);
buf BUF1 (N1938, N1923);
xor XOR2 (N1939, N1910, N767);
buf BUF1 (N1940, N1938);
not NOT1 (N1941, N1926);
and AND4 (N1942, N1928, N308, N1098, N183);
xor XOR2 (N1943, N1939, N1599);
or OR4 (N1944, N1934, N201, N1597, N1242);
not NOT1 (N1945, N1913);
xor XOR2 (N1946, N1919, N336);
buf BUF1 (N1947, N1907);
or OR3 (N1948, N1942, N1595, N1688);
not NOT1 (N1949, N1947);
and AND3 (N1950, N1949, N865, N90);
buf BUF1 (N1951, N1948);
not NOT1 (N1952, N1946);
nor NOR4 (N1953, N1944, N1794, N975, N1212);
buf BUF1 (N1954, N1950);
or OR4 (N1955, N1953, N900, N1660, N778);
nand NAND3 (N1956, N1940, N236, N819);
or OR4 (N1957, N1951, N1910, N1666, N1797);
not NOT1 (N1958, N1943);
nor NOR2 (N1959, N1937, N1514);
not NOT1 (N1960, N1956);
nand NAND3 (N1961, N1941, N1036, N1800);
buf BUF1 (N1962, N1960);
buf BUF1 (N1963, N1959);
or OR2 (N1964, N1955, N449);
nand NAND4 (N1965, N1954, N825, N1262, N402);
or OR4 (N1966, N1958, N1068, N75, N776);
nand NAND4 (N1967, N1965, N266, N1551, N1741);
and AND2 (N1968, N1935, N734);
buf BUF1 (N1969, N1964);
and AND2 (N1970, N1966, N15);
xor XOR2 (N1971, N1968, N1356);
nand NAND4 (N1972, N1945, N1379, N1897, N659);
and AND2 (N1973, N1962, N1826);
xor XOR2 (N1974, N1972, N203);
nor NOR4 (N1975, N1957, N957, N1401, N360);
buf BUF1 (N1976, N1967);
and AND2 (N1977, N1963, N466);
xor XOR2 (N1978, N1974, N1946);
buf BUF1 (N1979, N1971);
or OR3 (N1980, N1978, N1404, N1859);
and AND2 (N1981, N1976, N276);
xor XOR2 (N1982, N1979, N851);
buf BUF1 (N1983, N1961);
nor NOR3 (N1984, N1983, N1193, N1835);
xor XOR2 (N1985, N1973, N989);
nand NAND2 (N1986, N1982, N214);
or OR3 (N1987, N1969, N1766, N690);
not NOT1 (N1988, N1986);
not NOT1 (N1989, N1984);
nand NAND2 (N1990, N1980, N1141);
nand NAND4 (N1991, N1981, N587, N966, N1420);
not NOT1 (N1992, N1985);
xor XOR2 (N1993, N1987, N533);
xor XOR2 (N1994, N1991, N607);
nand NAND4 (N1995, N1988, N295, N460, N1306);
buf BUF1 (N1996, N1977);
nor NOR3 (N1997, N1990, N1450, N1483);
and AND4 (N1998, N1975, N3, N1564, N433);
nand NAND3 (N1999, N1970, N314, N223);
or OR4 (N2000, N1996, N1404, N1078, N1765);
and AND3 (N2001, N1998, N283, N1479);
nand NAND3 (N2002, N2000, N1365, N630);
and AND2 (N2003, N1989, N1472);
xor XOR2 (N2004, N1952, N1133);
and AND2 (N2005, N1999, N732);
or OR2 (N2006, N1993, N263);
xor XOR2 (N2007, N1994, N1651);
and AND2 (N2008, N1997, N36);
nor NOR2 (N2009, N1995, N351);
nor NOR2 (N2010, N1992, N854);
nor NOR4 (N2011, N2001, N1577, N1676, N1438);
and AND2 (N2012, N2011, N1688);
nand NAND3 (N2013, N2005, N1992, N1140);
not NOT1 (N2014, N2004);
not NOT1 (N2015, N2002);
not NOT1 (N2016, N2013);
and AND2 (N2017, N2008, N617);
or OR2 (N2018, N2010, N1855);
and AND4 (N2019, N2006, N1953, N946, N1756);
or OR2 (N2020, N2019, N750);
not NOT1 (N2021, N2003);
not NOT1 (N2022, N2016);
not NOT1 (N2023, N2014);
and AND2 (N2024, N2023, N539);
or OR2 (N2025, N2018, N80);
not NOT1 (N2026, N2015);
and AND3 (N2027, N2024, N1354, N886);
nand NAND2 (N2028, N2026, N100);
or OR2 (N2029, N2012, N556);
xor XOR2 (N2030, N2025, N99);
or OR2 (N2031, N2022, N1152);
xor XOR2 (N2032, N2029, N157);
xor XOR2 (N2033, N2031, N1508);
xor XOR2 (N2034, N2028, N1173);
nor NOR3 (N2035, N2030, N1958, N1026);
nor NOR2 (N2036, N2007, N1688);
xor XOR2 (N2037, N2027, N1048);
and AND4 (N2038, N2032, N1488, N1898, N156);
buf BUF1 (N2039, N2036);
xor XOR2 (N2040, N2038, N1815);
nand NAND2 (N2041, N2009, N1847);
and AND3 (N2042, N2041, N934, N722);
xor XOR2 (N2043, N2037, N1066);
buf BUF1 (N2044, N2021);
buf BUF1 (N2045, N2034);
or OR4 (N2046, N2043, N1597, N1478, N1825);
nand NAND3 (N2047, N2044, N747, N823);
xor XOR2 (N2048, N2047, N1882);
or OR4 (N2049, N2039, N634, N1408, N742);
not NOT1 (N2050, N2049);
nor NOR3 (N2051, N2048, N1903, N389);
and AND3 (N2052, N2050, N1355, N34);
not NOT1 (N2053, N2045);
buf BUF1 (N2054, N2033);
and AND2 (N2055, N2054, N1659);
and AND4 (N2056, N2052, N1501, N849, N127);
nor NOR4 (N2057, N2035, N1268, N662, N1652);
nor NOR2 (N2058, N2053, N1844);
and AND3 (N2059, N2058, N661, N29);
not NOT1 (N2060, N2017);
or OR3 (N2061, N2055, N1329, N1109);
nand NAND4 (N2062, N2020, N1562, N1249, N861);
buf BUF1 (N2063, N2056);
buf BUF1 (N2064, N2042);
or OR2 (N2065, N2046, N1643);
or OR2 (N2066, N2040, N1592);
not NOT1 (N2067, N2061);
or OR4 (N2068, N2060, N2050, N224, N1389);
xor XOR2 (N2069, N2068, N1902);
not NOT1 (N2070, N2051);
not NOT1 (N2071, N2059);
nand NAND2 (N2072, N2067, N1970);
nand NAND2 (N2073, N2066, N1539);
not NOT1 (N2074, N2065);
and AND3 (N2075, N2064, N897, N1639);
buf BUF1 (N2076, N2072);
nand NAND3 (N2077, N2063, N50, N66);
buf BUF1 (N2078, N2062);
nor NOR3 (N2079, N2074, N1191, N1470);
nand NAND4 (N2080, N2069, N1143, N386, N619);
nor NOR2 (N2081, N2071, N215);
nand NAND3 (N2082, N2057, N576, N7);
nand NAND3 (N2083, N2076, N688, N1819);
not NOT1 (N2084, N2080);
not NOT1 (N2085, N2079);
buf BUF1 (N2086, N2081);
xor XOR2 (N2087, N2075, N869);
xor XOR2 (N2088, N2082, N1849);
buf BUF1 (N2089, N2087);
buf BUF1 (N2090, N2070);
and AND3 (N2091, N2085, N1070, N1492);
or OR3 (N2092, N2088, N201, N561);
and AND4 (N2093, N2089, N940, N497, N1773);
nor NOR3 (N2094, N2091, N1197, N752);
nor NOR4 (N2095, N2077, N927, N491, N1147);
xor XOR2 (N2096, N2095, N810);
not NOT1 (N2097, N2086);
nor NOR3 (N2098, N2092, N21, N745);
nor NOR3 (N2099, N2078, N1556, N671);
and AND2 (N2100, N2084, N1009);
xor XOR2 (N2101, N2097, N1367);
nand NAND4 (N2102, N2098, N1474, N1259, N908);
buf BUF1 (N2103, N2102);
and AND3 (N2104, N2103, N1359, N1437);
nor NOR3 (N2105, N2073, N1299, N1449);
nand NAND3 (N2106, N2096, N830, N2044);
or OR4 (N2107, N2094, N1089, N935, N661);
nand NAND3 (N2108, N2093, N1297, N286);
buf BUF1 (N2109, N2101);
or OR2 (N2110, N2104, N563);
xor XOR2 (N2111, N2110, N1347);
buf BUF1 (N2112, N2090);
nand NAND3 (N2113, N2083, N529, N1498);
nor NOR2 (N2114, N2108, N19);
xor XOR2 (N2115, N2114, N1564);
not NOT1 (N2116, N2099);
xor XOR2 (N2117, N2116, N1388);
buf BUF1 (N2118, N2100);
nand NAND3 (N2119, N2109, N666, N2090);
xor XOR2 (N2120, N2119, N1400);
nor NOR4 (N2121, N2107, N1945, N1538, N763);
and AND3 (N2122, N2115, N1721, N1852);
buf BUF1 (N2123, N2106);
buf BUF1 (N2124, N2122);
buf BUF1 (N2125, N2112);
nand NAND4 (N2126, N2125, N1162, N1726, N927);
xor XOR2 (N2127, N2111, N1476);
or OR2 (N2128, N2117, N2006);
nand NAND4 (N2129, N2124, N1846, N898, N493);
xor XOR2 (N2130, N2127, N1639);
nand NAND4 (N2131, N2118, N1267, N367, N906);
nor NOR3 (N2132, N2123, N1575, N816);
nor NOR3 (N2133, N2120, N1431, N1378);
xor XOR2 (N2134, N2133, N280);
not NOT1 (N2135, N2131);
buf BUF1 (N2136, N2128);
nor NOR3 (N2137, N2135, N1898, N2028);
or OR4 (N2138, N2130, N193, N2109, N1944);
not NOT1 (N2139, N2126);
nor NOR3 (N2140, N2105, N1069, N1912);
buf BUF1 (N2141, N2132);
buf BUF1 (N2142, N2113);
and AND2 (N2143, N2136, N189);
xor XOR2 (N2144, N2143, N2105);
and AND3 (N2145, N2144, N1582, N229);
or OR4 (N2146, N2141, N980, N501, N966);
nand NAND4 (N2147, N2139, N1852, N1795, N725);
buf BUF1 (N2148, N2140);
not NOT1 (N2149, N2148);
or OR3 (N2150, N2142, N590, N199);
and AND3 (N2151, N2150, N804, N813);
nor NOR2 (N2152, N2138, N1923);
and AND2 (N2153, N2129, N1982);
not NOT1 (N2154, N2149);
nor NOR4 (N2155, N2154, N1081, N1498, N1302);
or OR3 (N2156, N2155, N1937, N610);
nand NAND3 (N2157, N2147, N761, N902);
not NOT1 (N2158, N2121);
and AND3 (N2159, N2137, N465, N1919);
xor XOR2 (N2160, N2151, N660);
xor XOR2 (N2161, N2158, N959);
and AND4 (N2162, N2145, N745, N1436, N1367);
nand NAND2 (N2163, N2156, N1820);
or OR2 (N2164, N2162, N451);
not NOT1 (N2165, N2160);
not NOT1 (N2166, N2157);
and AND2 (N2167, N2164, N1552);
nand NAND3 (N2168, N2146, N557, N132);
buf BUF1 (N2169, N2168);
buf BUF1 (N2170, N2165);
and AND3 (N2171, N2169, N1124, N264);
nor NOR4 (N2172, N2152, N1992, N750, N1638);
and AND4 (N2173, N2153, N266, N1919, N889);
and AND2 (N2174, N2172, N1736);
or OR4 (N2175, N2163, N721, N889, N428);
or OR3 (N2176, N2159, N1770, N333);
nand NAND3 (N2177, N2174, N2022, N380);
buf BUF1 (N2178, N2173);
buf BUF1 (N2179, N2175);
nor NOR2 (N2180, N2166, N860);
nand NAND3 (N2181, N2170, N2107, N2041);
nand NAND4 (N2182, N2176, N146, N1859, N1545);
xor XOR2 (N2183, N2171, N1149);
nor NOR4 (N2184, N2167, N137, N792, N371);
nor NOR3 (N2185, N2161, N88, N1405);
nand NAND2 (N2186, N2183, N424);
nor NOR3 (N2187, N2181, N1096, N511);
buf BUF1 (N2188, N2185);
nor NOR2 (N2189, N2182, N739);
and AND4 (N2190, N2177, N887, N13, N1617);
and AND4 (N2191, N2189, N1833, N2066, N597);
nor NOR3 (N2192, N2188, N753, N2178);
not NOT1 (N2193, N882);
nor NOR4 (N2194, N2191, N2106, N1929, N1513);
and AND2 (N2195, N2194, N1965);
and AND3 (N2196, N2192, N745, N1889);
buf BUF1 (N2197, N2196);
or OR2 (N2198, N2186, N895);
or OR4 (N2199, N2190, N783, N357, N1000);
nor NOR2 (N2200, N2193, N2148);
or OR4 (N2201, N2200, N893, N1660, N1061);
and AND3 (N2202, N2184, N594, N1614);
and AND3 (N2203, N2180, N1047, N2036);
or OR4 (N2204, N2202, N376, N268, N2094);
or OR2 (N2205, N2198, N2050);
buf BUF1 (N2206, N2204);
and AND2 (N2207, N2187, N1432);
nor NOR2 (N2208, N2134, N774);
xor XOR2 (N2209, N2201, N2081);
or OR2 (N2210, N2197, N352);
nor NOR4 (N2211, N2209, N1705, N1866, N1823);
not NOT1 (N2212, N2207);
buf BUF1 (N2213, N2203);
nand NAND2 (N2214, N2208, N1173);
or OR4 (N2215, N2199, N1649, N122, N500);
xor XOR2 (N2216, N2211, N400);
and AND3 (N2217, N2210, N1892, N2047);
xor XOR2 (N2218, N2215, N2046);
nand NAND4 (N2219, N2218, N1455, N1527, N1208);
or OR2 (N2220, N2179, N170);
nand NAND3 (N2221, N2216, N352, N1957);
not NOT1 (N2222, N2220);
and AND3 (N2223, N2214, N54, N911);
and AND3 (N2224, N2217, N519, N871);
nor NOR4 (N2225, N2213, N518, N493, N1796);
buf BUF1 (N2226, N2205);
xor XOR2 (N2227, N2221, N66);
and AND4 (N2228, N2219, N539, N1406, N1251);
or OR4 (N2229, N2224, N863, N190, N923);
or OR2 (N2230, N2222, N1794);
nand NAND4 (N2231, N2227, N863, N190, N1362);
xor XOR2 (N2232, N2195, N1802);
not NOT1 (N2233, N2206);
nand NAND3 (N2234, N2231, N184, N67);
or OR3 (N2235, N2230, N553, N252);
buf BUF1 (N2236, N2226);
and AND3 (N2237, N2232, N1092, N1937);
and AND2 (N2238, N2228, N1596);
or OR3 (N2239, N2234, N187, N769);
nand NAND3 (N2240, N2239, N782, N41);
and AND4 (N2241, N2225, N959, N1960, N875);
nand NAND4 (N2242, N2235, N1779, N1623, N2103);
not NOT1 (N2243, N2242);
buf BUF1 (N2244, N2223);
xor XOR2 (N2245, N2241, N2106);
or OR2 (N2246, N2233, N1874);
or OR2 (N2247, N2243, N381);
xor XOR2 (N2248, N2238, N501);
or OR4 (N2249, N2248, N634, N1368, N1596);
nand NAND2 (N2250, N2237, N1104);
xor XOR2 (N2251, N2244, N1659);
not NOT1 (N2252, N2229);
not NOT1 (N2253, N2240);
nor NOR4 (N2254, N2249, N2021, N1251, N1041);
nand NAND4 (N2255, N2247, N309, N169, N1449);
nand NAND2 (N2256, N2246, N2149);
and AND2 (N2257, N2236, N2037);
nand NAND4 (N2258, N2245, N1552, N2171, N23);
or OR3 (N2259, N2212, N1730, N600);
nand NAND4 (N2260, N2257, N1865, N776, N889);
xor XOR2 (N2261, N2259, N1127);
buf BUF1 (N2262, N2254);
or OR3 (N2263, N2262, N2038, N1375);
and AND4 (N2264, N2252, N1389, N58, N964);
nor NOR2 (N2265, N2258, N1574);
and AND4 (N2266, N2261, N1132, N927, N1642);
xor XOR2 (N2267, N2250, N2044);
xor XOR2 (N2268, N2263, N1271);
nor NOR3 (N2269, N2266, N2195, N693);
nand NAND4 (N2270, N2253, N2136, N1529, N772);
nand NAND2 (N2271, N2255, N247);
nor NOR3 (N2272, N2268, N52, N2184);
or OR4 (N2273, N2269, N2232, N1850, N937);
nor NOR2 (N2274, N2272, N1574);
not NOT1 (N2275, N2256);
buf BUF1 (N2276, N2260);
and AND4 (N2277, N2265, N2190, N388, N1091);
xor XOR2 (N2278, N2275, N532);
buf BUF1 (N2279, N2276);
nor NOR2 (N2280, N2277, N1701);
or OR3 (N2281, N2271, N1471, N187);
nor NOR4 (N2282, N2278, N871, N446, N862);
not NOT1 (N2283, N2274);
xor XOR2 (N2284, N2281, N356);
nor NOR2 (N2285, N2270, N2086);
and AND4 (N2286, N2279, N2092, N1265, N14);
xor XOR2 (N2287, N2284, N1398);
and AND3 (N2288, N2287, N231, N464);
buf BUF1 (N2289, N2286);
nand NAND2 (N2290, N2267, N1797);
and AND4 (N2291, N2282, N47, N1251, N2150);
not NOT1 (N2292, N2283);
or OR3 (N2293, N2285, N2161, N729);
or OR3 (N2294, N2291, N2221, N1923);
or OR3 (N2295, N2251, N1997, N1709);
nor NOR3 (N2296, N2280, N1426, N1075);
not NOT1 (N2297, N2292);
and AND3 (N2298, N2293, N752, N1699);
xor XOR2 (N2299, N2295, N87);
nand NAND4 (N2300, N2298, N633, N668, N1584);
xor XOR2 (N2301, N2290, N1400);
and AND3 (N2302, N2289, N1036, N2150);
not NOT1 (N2303, N2296);
buf BUF1 (N2304, N2273);
not NOT1 (N2305, N2288);
nor NOR4 (N2306, N2297, N50, N244, N1771);
or OR3 (N2307, N2305, N532, N1766);
nand NAND3 (N2308, N2264, N255, N578);
nor NOR3 (N2309, N2299, N1700, N1097);
xor XOR2 (N2310, N2303, N856);
nand NAND4 (N2311, N2302, N1866, N120, N1708);
xor XOR2 (N2312, N2309, N2015);
nand NAND4 (N2313, N2308, N714, N2043, N498);
xor XOR2 (N2314, N2313, N1769);
xor XOR2 (N2315, N2304, N1157);
nor NOR4 (N2316, N2314, N1140, N2130, N367);
not NOT1 (N2317, N2311);
not NOT1 (N2318, N2317);
nand NAND4 (N2319, N2294, N391, N1456, N595);
nand NAND4 (N2320, N2306, N2137, N2298, N1310);
nor NOR2 (N2321, N2320, N2111);
and AND3 (N2322, N2321, N974, N552);
and AND2 (N2323, N2318, N109);
or OR4 (N2324, N2323, N344, N1428, N387);
nand NAND3 (N2325, N2322, N526, N114);
xor XOR2 (N2326, N2300, N360);
buf BUF1 (N2327, N2326);
nor NOR2 (N2328, N2310, N763);
xor XOR2 (N2329, N2319, N105);
or OR2 (N2330, N2327, N539);
nand NAND4 (N2331, N2329, N2179, N1737, N1262);
or OR4 (N2332, N2325, N923, N1279, N1486);
and AND2 (N2333, N2301, N1076);
and AND3 (N2334, N2315, N48, N132);
not NOT1 (N2335, N2307);
or OR2 (N2336, N2324, N945);
or OR4 (N2337, N2316, N563, N382, N1530);
and AND3 (N2338, N2337, N1998, N1583);
not NOT1 (N2339, N2333);
and AND2 (N2340, N2312, N1405);
or OR3 (N2341, N2334, N842, N395);
buf BUF1 (N2342, N2339);
nor NOR2 (N2343, N2338, N1031);
buf BUF1 (N2344, N2340);
nand NAND2 (N2345, N2344, N1684);
nand NAND2 (N2346, N2331, N1709);
not NOT1 (N2347, N2345);
xor XOR2 (N2348, N2346, N776);
or OR3 (N2349, N2342, N1950, N867);
not NOT1 (N2350, N2330);
xor XOR2 (N2351, N2343, N1303);
not NOT1 (N2352, N2348);
xor XOR2 (N2353, N2350, N1295);
buf BUF1 (N2354, N2347);
or OR3 (N2355, N2351, N978, N1102);
buf BUF1 (N2356, N2355);
buf BUF1 (N2357, N2352);
buf BUF1 (N2358, N2335);
or OR2 (N2359, N2356, N1510);
buf BUF1 (N2360, N2341);
or OR4 (N2361, N2354, N1272, N1134, N685);
and AND4 (N2362, N2361, N62, N1423, N299);
and AND2 (N2363, N2360, N1683);
nor NOR3 (N2364, N2336, N1897, N2069);
or OR2 (N2365, N2359, N1570);
not NOT1 (N2366, N2353);
buf BUF1 (N2367, N2365);
or OR3 (N2368, N2357, N99, N1112);
or OR4 (N2369, N2367, N2125, N897, N1632);
nand NAND2 (N2370, N2363, N1364);
buf BUF1 (N2371, N2370);
xor XOR2 (N2372, N2358, N1679);
and AND2 (N2373, N2364, N313);
nor NOR4 (N2374, N2349, N754, N1554, N349);
xor XOR2 (N2375, N2368, N893);
and AND4 (N2376, N2374, N140, N2122, N321);
and AND4 (N2377, N2369, N1707, N150, N1552);
and AND4 (N2378, N2372, N2283, N2344, N133);
buf BUF1 (N2379, N2375);
not NOT1 (N2380, N2376);
not NOT1 (N2381, N2371);
nor NOR2 (N2382, N2373, N1514);
or OR2 (N2383, N2362, N633);
nor NOR3 (N2384, N2328, N1212, N1456);
nor NOR3 (N2385, N2332, N1983, N1667);
nor NOR2 (N2386, N2381, N526);
not NOT1 (N2387, N2383);
not NOT1 (N2388, N2379);
xor XOR2 (N2389, N2386, N1301);
buf BUF1 (N2390, N2380);
nor NOR3 (N2391, N2389, N2220, N393);
buf BUF1 (N2392, N2391);
not NOT1 (N2393, N2385);
nor NOR2 (N2394, N2387, N1438);
buf BUF1 (N2395, N2378);
nand NAND4 (N2396, N2377, N1719, N488, N679);
xor XOR2 (N2397, N2382, N1542);
buf BUF1 (N2398, N2394);
nand NAND2 (N2399, N2384, N1502);
not NOT1 (N2400, N2393);
nand NAND2 (N2401, N2397, N553);
or OR3 (N2402, N2400, N2286, N1929);
xor XOR2 (N2403, N2401, N815);
and AND4 (N2404, N2388, N565, N881, N898);
buf BUF1 (N2405, N2395);
and AND2 (N2406, N2399, N421);
or OR4 (N2407, N2396, N748, N1207, N1712);
nand NAND3 (N2408, N2398, N1977, N1248);
nand NAND3 (N2409, N2405, N945, N1526);
not NOT1 (N2410, N2390);
and AND4 (N2411, N2408, N1641, N744, N1255);
nor NOR4 (N2412, N2411, N983, N881, N1947);
and AND4 (N2413, N2404, N2179, N755, N52);
and AND3 (N2414, N2392, N1019, N2347);
buf BUF1 (N2415, N2410);
nand NAND2 (N2416, N2414, N1443);
xor XOR2 (N2417, N2412, N1751);
not NOT1 (N2418, N2402);
not NOT1 (N2419, N2366);
or OR4 (N2420, N2418, N1611, N1392, N2060);
not NOT1 (N2421, N2419);
or OR3 (N2422, N2420, N351, N780);
or OR4 (N2423, N2421, N2281, N1658, N158);
buf BUF1 (N2424, N2406);
buf BUF1 (N2425, N2424);
xor XOR2 (N2426, N2407, N1815);
nand NAND2 (N2427, N2409, N2007);
buf BUF1 (N2428, N2403);
and AND2 (N2429, N2415, N1027);
not NOT1 (N2430, N2417);
buf BUF1 (N2431, N2422);
nor NOR3 (N2432, N2431, N653, N234);
nor NOR2 (N2433, N2428, N1419);
nand NAND3 (N2434, N2413, N59, N2328);
buf BUF1 (N2435, N2432);
nand NAND3 (N2436, N2427, N1301, N1933);
nand NAND2 (N2437, N2426, N1431);
xor XOR2 (N2438, N2430, N1506);
not NOT1 (N2439, N2429);
nor NOR3 (N2440, N2434, N479, N1675);
or OR3 (N2441, N2416, N590, N888);
buf BUF1 (N2442, N2433);
and AND3 (N2443, N2435, N2216, N179);
nor NOR2 (N2444, N2423, N2059);
nand NAND4 (N2445, N2440, N2299, N1867, N188);
nor NOR2 (N2446, N2425, N1911);
buf BUF1 (N2447, N2436);
nor NOR2 (N2448, N2437, N1750);
or OR2 (N2449, N2443, N718);
nand NAND2 (N2450, N2446, N1457);
xor XOR2 (N2451, N2447, N2292);
xor XOR2 (N2452, N2442, N496);
nand NAND3 (N2453, N2448, N1632, N1728);
xor XOR2 (N2454, N2453, N329);
and AND4 (N2455, N2451, N1149, N477, N698);
xor XOR2 (N2456, N2449, N1655);
xor XOR2 (N2457, N2444, N964);
or OR2 (N2458, N2439, N92);
xor XOR2 (N2459, N2458, N2076);
not NOT1 (N2460, N2456);
buf BUF1 (N2461, N2452);
and AND3 (N2462, N2445, N1618, N361);
nor NOR3 (N2463, N2462, N558, N1353);
buf BUF1 (N2464, N2450);
nand NAND4 (N2465, N2454, N359, N2290, N1073);
nor NOR4 (N2466, N2457, N380, N1071, N447);
nand NAND3 (N2467, N2463, N2014, N585);
xor XOR2 (N2468, N2438, N460);
not NOT1 (N2469, N2466);
xor XOR2 (N2470, N2468, N954);
xor XOR2 (N2471, N2464, N988);
not NOT1 (N2472, N2459);
nor NOR4 (N2473, N2461, N395, N1136, N225);
nor NOR2 (N2474, N2455, N993);
not NOT1 (N2475, N2460);
not NOT1 (N2476, N2465);
and AND2 (N2477, N2441, N508);
buf BUF1 (N2478, N2475);
nor NOR2 (N2479, N2470, N693);
and AND4 (N2480, N2477, N1501, N693, N1456);
xor XOR2 (N2481, N2469, N1557);
buf BUF1 (N2482, N2478);
buf BUF1 (N2483, N2482);
buf BUF1 (N2484, N2476);
and AND4 (N2485, N2474, N1755, N465, N878);
buf BUF1 (N2486, N2471);
not NOT1 (N2487, N2479);
and AND2 (N2488, N2484, N656);
nand NAND2 (N2489, N2486, N1828);
buf BUF1 (N2490, N2472);
and AND3 (N2491, N2488, N1266, N1163);
buf BUF1 (N2492, N2483);
buf BUF1 (N2493, N2481);
xor XOR2 (N2494, N2485, N375);
and AND3 (N2495, N2487, N1381, N1766);
xor XOR2 (N2496, N2467, N275);
nor NOR4 (N2497, N2492, N1217, N2227, N1218);
xor XOR2 (N2498, N2480, N1659);
and AND2 (N2499, N2494, N688);
nor NOR4 (N2500, N2491, N924, N43, N575);
not NOT1 (N2501, N2495);
and AND2 (N2502, N2499, N2380);
buf BUF1 (N2503, N2498);
or OR3 (N2504, N2501, N474, N1981);
not NOT1 (N2505, N2503);
nand NAND3 (N2506, N2497, N1577, N2263);
not NOT1 (N2507, N2505);
and AND3 (N2508, N2490, N1739, N77);
and AND2 (N2509, N2504, N1847);
buf BUF1 (N2510, N2473);
nor NOR4 (N2511, N2508, N2093, N765, N2411);
nor NOR2 (N2512, N2496, N1219);
nand NAND2 (N2513, N2507, N1165);
nor NOR2 (N2514, N2489, N1474);
nand NAND4 (N2515, N2502, N2137, N535, N2465);
xor XOR2 (N2516, N2513, N2309);
buf BUF1 (N2517, N2500);
xor XOR2 (N2518, N2509, N2432);
xor XOR2 (N2519, N2515, N573);
nand NAND4 (N2520, N2518, N2119, N1934, N2132);
buf BUF1 (N2521, N2506);
nor NOR3 (N2522, N2510, N990, N1096);
and AND4 (N2523, N2493, N361, N1907, N2407);
buf BUF1 (N2524, N2520);
xor XOR2 (N2525, N2512, N46);
nor NOR3 (N2526, N2517, N2033, N2156);
nor NOR2 (N2527, N2523, N1394);
not NOT1 (N2528, N2527);
and AND4 (N2529, N2516, N789, N527, N510);
xor XOR2 (N2530, N2511, N2161);
and AND4 (N2531, N2514, N1357, N2502, N1030);
nor NOR4 (N2532, N2524, N1783, N196, N2001);
nand NAND4 (N2533, N2531, N1012, N280, N1405);
nand NAND3 (N2534, N2525, N982, N2459);
nor NOR2 (N2535, N2533, N2124);
not NOT1 (N2536, N2522);
xor XOR2 (N2537, N2529, N843);
nand NAND4 (N2538, N2534, N380, N640, N1636);
nand NAND2 (N2539, N2536, N1275);
nand NAND2 (N2540, N2530, N1333);
xor XOR2 (N2541, N2538, N2187);
or OR3 (N2542, N2521, N810, N1299);
xor XOR2 (N2543, N2541, N1362);
or OR3 (N2544, N2519, N1274, N523);
nor NOR3 (N2545, N2544, N839, N997);
buf BUF1 (N2546, N2545);
buf BUF1 (N2547, N2537);
buf BUF1 (N2548, N2547);
nand NAND4 (N2549, N2542, N2207, N1144, N2201);
buf BUF1 (N2550, N2543);
buf BUF1 (N2551, N2535);
nor NOR3 (N2552, N2540, N1144, N1126);
not NOT1 (N2553, N2532);
and AND3 (N2554, N2528, N1029, N1353);
nor NOR4 (N2555, N2553, N156, N400, N2291);
buf BUF1 (N2556, N2526);
or OR4 (N2557, N2548, N642, N664, N1744);
not NOT1 (N2558, N2539);
or OR3 (N2559, N2554, N2214, N2166);
nor NOR4 (N2560, N2559, N684, N1563, N337);
nand NAND4 (N2561, N2546, N2321, N2462, N2218);
nor NOR2 (N2562, N2560, N1424);
nand NAND2 (N2563, N2555, N1121);
and AND2 (N2564, N2561, N1447);
nor NOR3 (N2565, N2563, N279, N2479);
buf BUF1 (N2566, N2550);
or OR2 (N2567, N2564, N681);
nor NOR2 (N2568, N2549, N275);
not NOT1 (N2569, N2557);
not NOT1 (N2570, N2569);
and AND2 (N2571, N2552, N269);
or OR3 (N2572, N2565, N1364, N2427);
not NOT1 (N2573, N2572);
xor XOR2 (N2574, N2556, N1486);
and AND3 (N2575, N2574, N542, N953);
buf BUF1 (N2576, N2562);
not NOT1 (N2577, N2566);
xor XOR2 (N2578, N2567, N402);
and AND4 (N2579, N2577, N2546, N523, N859);
or OR3 (N2580, N2575, N63, N1324);
nor NOR4 (N2581, N2570, N2052, N2018, N2260);
nand NAND3 (N2582, N2578, N200, N1734);
and AND2 (N2583, N2579, N1306);
nor NOR3 (N2584, N2583, N571, N519);
and AND3 (N2585, N2573, N1343, N532);
nand NAND3 (N2586, N2558, N1291, N2219);
not NOT1 (N2587, N2586);
nand NAND2 (N2588, N2576, N672);
nand NAND2 (N2589, N2581, N1381);
and AND2 (N2590, N2585, N451);
xor XOR2 (N2591, N2582, N1104);
or OR3 (N2592, N2580, N935, N1542);
nand NAND3 (N2593, N2592, N1513, N629);
or OR4 (N2594, N2591, N2489, N810, N56);
buf BUF1 (N2595, N2590);
nand NAND4 (N2596, N2593, N678, N395, N385);
xor XOR2 (N2597, N2589, N1804);
nor NOR4 (N2598, N2596, N979, N377, N269);
buf BUF1 (N2599, N2597);
nand NAND4 (N2600, N2584, N417, N1835, N715);
nor NOR2 (N2601, N2594, N2262);
not NOT1 (N2602, N2599);
buf BUF1 (N2603, N2600);
and AND2 (N2604, N2587, N641);
or OR3 (N2605, N2602, N714, N2541);
and AND3 (N2606, N2605, N367, N1719);
or OR3 (N2607, N2551, N2342, N1713);
nand NAND2 (N2608, N2571, N628);
and AND3 (N2609, N2598, N791, N1531);
nor NOR2 (N2610, N2603, N638);
buf BUF1 (N2611, N2609);
nand NAND2 (N2612, N2604, N1824);
nand NAND3 (N2613, N2601, N59, N369);
not NOT1 (N2614, N2595);
buf BUF1 (N2615, N2612);
nor NOR3 (N2616, N2568, N2066, N1560);
and AND3 (N2617, N2616, N1621, N1001);
or OR2 (N2618, N2606, N1862);
nand NAND2 (N2619, N2617, N1938);
or OR3 (N2620, N2618, N1967, N2281);
not NOT1 (N2621, N2608);
xor XOR2 (N2622, N2619, N1175);
xor XOR2 (N2623, N2613, N2442);
and AND3 (N2624, N2621, N2159, N2056);
nand NAND4 (N2625, N2611, N921, N2308, N2241);
buf BUF1 (N2626, N2623);
buf BUF1 (N2627, N2615);
nand NAND4 (N2628, N2625, N457, N183, N480);
and AND3 (N2629, N2628, N2628, N1518);
or OR3 (N2630, N2588, N33, N1859);
and AND2 (N2631, N2624, N1839);
not NOT1 (N2632, N2631);
buf BUF1 (N2633, N2614);
buf BUF1 (N2634, N2622);
xor XOR2 (N2635, N2627, N1401);
or OR4 (N2636, N2626, N639, N2096, N1415);
buf BUF1 (N2637, N2620);
xor XOR2 (N2638, N2633, N1304);
buf BUF1 (N2639, N2607);
nor NOR4 (N2640, N2636, N1279, N844, N401);
nand NAND2 (N2641, N2632, N28);
nand NAND3 (N2642, N2610, N1153, N1970);
nor NOR3 (N2643, N2641, N2202, N888);
nor NOR2 (N2644, N2635, N2396);
and AND2 (N2645, N2639, N164);
not NOT1 (N2646, N2644);
nand NAND2 (N2647, N2640, N448);
and AND3 (N2648, N2634, N1086, N1272);
nor NOR2 (N2649, N2638, N546);
not NOT1 (N2650, N2642);
nand NAND2 (N2651, N2649, N1589);
nand NAND3 (N2652, N2646, N1226, N406);
xor XOR2 (N2653, N2652, N1408);
and AND4 (N2654, N2645, N1353, N374, N348);
nand NAND4 (N2655, N2650, N2506, N1240, N1963);
nand NAND2 (N2656, N2654, N560);
and AND2 (N2657, N2647, N518);
or OR3 (N2658, N2657, N735, N1416);
and AND2 (N2659, N2648, N1451);
nand NAND3 (N2660, N2655, N526, N1833);
buf BUF1 (N2661, N2629);
not NOT1 (N2662, N2661);
and AND2 (N2663, N2651, N662);
xor XOR2 (N2664, N2643, N86);
xor XOR2 (N2665, N2664, N1036);
nor NOR3 (N2666, N2653, N1439, N2061);
and AND3 (N2667, N2659, N2605, N360);
and AND2 (N2668, N2665, N2667);
buf BUF1 (N2669, N2362);
or OR3 (N2670, N2663, N1698, N2641);
or OR2 (N2671, N2669, N761);
not NOT1 (N2672, N2666);
nand NAND3 (N2673, N2637, N717, N2476);
or OR2 (N2674, N2660, N2605);
or OR2 (N2675, N2630, N1558);
and AND4 (N2676, N2658, N2673, N2180, N271);
not NOT1 (N2677, N782);
nor NOR3 (N2678, N2668, N509, N323);
nand NAND3 (N2679, N2674, N502, N2092);
nand NAND2 (N2680, N2670, N1834);
xor XOR2 (N2681, N2676, N1032);
nand NAND2 (N2682, N2662, N583);
not NOT1 (N2683, N2656);
nor NOR3 (N2684, N2679, N1713, N1480);
not NOT1 (N2685, N2683);
and AND2 (N2686, N2677, N1452);
xor XOR2 (N2687, N2678, N1109);
buf BUF1 (N2688, N2675);
xor XOR2 (N2689, N2671, N711);
nand NAND4 (N2690, N2685, N1963, N1437, N2099);
and AND2 (N2691, N2688, N1909);
or OR4 (N2692, N2681, N1274, N768, N2344);
xor XOR2 (N2693, N2672, N2618);
or OR3 (N2694, N2687, N1895, N750);
not NOT1 (N2695, N2689);
nor NOR2 (N2696, N2693, N813);
nor NOR3 (N2697, N2694, N1144, N2481);
not NOT1 (N2698, N2686);
or OR4 (N2699, N2698, N2098, N1315, N616);
not NOT1 (N2700, N2691);
xor XOR2 (N2701, N2680, N2002);
nor NOR2 (N2702, N2700, N1681);
or OR2 (N2703, N2692, N2564);
and AND4 (N2704, N2684, N2003, N1017, N2564);
nor NOR4 (N2705, N2690, N180, N2646, N2388);
nand NAND2 (N2706, N2703, N1019);
xor XOR2 (N2707, N2705, N2391);
or OR4 (N2708, N2707, N499, N1232, N2011);
nand NAND2 (N2709, N2704, N2094);
xor XOR2 (N2710, N2702, N2042);
or OR4 (N2711, N2709, N1591, N2424, N2547);
and AND2 (N2712, N2697, N1750);
buf BUF1 (N2713, N2699);
and AND2 (N2714, N2712, N923);
xor XOR2 (N2715, N2711, N1474);
xor XOR2 (N2716, N2715, N1052);
and AND2 (N2717, N2710, N1649);
and AND4 (N2718, N2701, N497, N2515, N1789);
nor NOR2 (N2719, N2713, N1396);
not NOT1 (N2720, N2682);
buf BUF1 (N2721, N2706);
buf BUF1 (N2722, N2719);
buf BUF1 (N2723, N2695);
not NOT1 (N2724, N2716);
not NOT1 (N2725, N2718);
or OR4 (N2726, N2721, N2564, N2574, N1445);
nand NAND2 (N2727, N2714, N1927);
buf BUF1 (N2728, N2708);
nand NAND4 (N2729, N2720, N259, N2401, N1489);
not NOT1 (N2730, N2729);
nand NAND4 (N2731, N2696, N673, N1918, N1562);
and AND4 (N2732, N2726, N83, N45, N1894);
nand NAND2 (N2733, N2717, N765);
nand NAND3 (N2734, N2731, N1258, N1394);
not NOT1 (N2735, N2724);
or OR2 (N2736, N2722, N1563);
nand NAND3 (N2737, N2730, N2485, N1695);
not NOT1 (N2738, N2735);
buf BUF1 (N2739, N2723);
nor NOR4 (N2740, N2727, N1103, N2309, N2039);
xor XOR2 (N2741, N2738, N2031);
nor NOR2 (N2742, N2740, N1868);
and AND3 (N2743, N2733, N1700, N667);
or OR2 (N2744, N2736, N1006);
nand NAND3 (N2745, N2744, N2739, N2479);
or OR2 (N2746, N1711, N757);
nand NAND4 (N2747, N2745, N2374, N1811, N463);
nand NAND4 (N2748, N2746, N1036, N1962, N2301);
xor XOR2 (N2749, N2725, N1184);
and AND4 (N2750, N2737, N541, N1037, N2144);
or OR4 (N2751, N2728, N1952, N338, N2673);
not NOT1 (N2752, N2751);
nand NAND4 (N2753, N2732, N1311, N403, N2537);
nor NOR4 (N2754, N2753, N1624, N410, N670);
or OR2 (N2755, N2741, N2025);
and AND3 (N2756, N2742, N2501, N700);
nor NOR4 (N2757, N2747, N78, N1054, N2133);
buf BUF1 (N2758, N2756);
xor XOR2 (N2759, N2755, N305);
and AND2 (N2760, N2759, N1817);
nor NOR3 (N2761, N2754, N2282, N1883);
or OR4 (N2762, N2750, N2418, N630, N1329);
nor NOR2 (N2763, N2762, N1703);
buf BUF1 (N2764, N2734);
or OR4 (N2765, N2763, N121, N1230, N2343);
not NOT1 (N2766, N2761);
or OR4 (N2767, N2758, N1502, N2480, N2683);
and AND2 (N2768, N2765, N670);
buf BUF1 (N2769, N2766);
or OR2 (N2770, N2760, N1728);
buf BUF1 (N2771, N2757);
nor NOR4 (N2772, N2770, N467, N2409, N1085);
nand NAND3 (N2773, N2772, N762, N2498);
nor NOR2 (N2774, N2749, N1766);
xor XOR2 (N2775, N2774, N1946);
xor XOR2 (N2776, N2768, N2355);
nor NOR3 (N2777, N2764, N350, N2452);
xor XOR2 (N2778, N2771, N775);
buf BUF1 (N2779, N2743);
buf BUF1 (N2780, N2769);
nor NOR4 (N2781, N2776, N945, N526, N412);
buf BUF1 (N2782, N2752);
nand NAND4 (N2783, N2775, N1274, N1252, N2205);
buf BUF1 (N2784, N2748);
and AND2 (N2785, N2782, N1633);
or OR4 (N2786, N2785, N1260, N858, N1248);
buf BUF1 (N2787, N2786);
or OR4 (N2788, N2780, N27, N176, N1566);
nor NOR2 (N2789, N2779, N1700);
nor NOR3 (N2790, N2778, N239, N2335);
nand NAND4 (N2791, N2787, N871, N44, N1565);
buf BUF1 (N2792, N2791);
or OR2 (N2793, N2790, N2132);
or OR4 (N2794, N2789, N710, N1304, N389);
nor NOR2 (N2795, N2794, N2225);
or OR3 (N2796, N2792, N997, N1413);
and AND4 (N2797, N2773, N853, N792, N1830);
not NOT1 (N2798, N2793);
and AND2 (N2799, N2784, N2788);
or OR4 (N2800, N196, N807, N783, N1675);
or OR4 (N2801, N2796, N2490, N98, N2780);
and AND4 (N2802, N2781, N1215, N2344, N1176);
nor NOR2 (N2803, N2800, N700);
nand NAND4 (N2804, N2798, N2181, N612, N637);
nor NOR4 (N2805, N2801, N1435, N1423, N2790);
or OR2 (N2806, N2777, N2288);
nor NOR4 (N2807, N2803, N1985, N2355, N919);
nand NAND2 (N2808, N2795, N188);
not NOT1 (N2809, N2767);
nand NAND4 (N2810, N2799, N1975, N2292, N2502);
xor XOR2 (N2811, N2783, N2564);
buf BUF1 (N2812, N2797);
xor XOR2 (N2813, N2806, N2375);
xor XOR2 (N2814, N2813, N883);
nand NAND4 (N2815, N2804, N1011, N884, N505);
xor XOR2 (N2816, N2811, N1363);
or OR2 (N2817, N2812, N2399);
not NOT1 (N2818, N2815);
not NOT1 (N2819, N2818);
nor NOR2 (N2820, N2810, N2049);
buf BUF1 (N2821, N2814);
nor NOR4 (N2822, N2807, N1490, N2806, N2126);
or OR3 (N2823, N2821, N2103, N2821);
buf BUF1 (N2824, N2819);
and AND3 (N2825, N2824, N711, N1804);
xor XOR2 (N2826, N2820, N518);
nor NOR2 (N2827, N2802, N496);
xor XOR2 (N2828, N2826, N2489);
or OR3 (N2829, N2809, N951, N2489);
nand NAND2 (N2830, N2829, N77);
nor NOR2 (N2831, N2823, N392);
nand NAND3 (N2832, N2822, N944, N2192);
nand NAND4 (N2833, N2828, N1561, N1408, N2639);
and AND3 (N2834, N2830, N431, N1919);
xor XOR2 (N2835, N2833, N1107);
nor NOR4 (N2836, N2831, N1051, N1425, N718);
buf BUF1 (N2837, N2832);
or OR3 (N2838, N2836, N120, N167);
nand NAND2 (N2839, N2837, N1571);
buf BUF1 (N2840, N2808);
xor XOR2 (N2841, N2827, N2812);
nor NOR4 (N2842, N2838, N2253, N2012, N749);
nor NOR3 (N2843, N2825, N1966, N157);
not NOT1 (N2844, N2842);
nand NAND2 (N2845, N2817, N813);
buf BUF1 (N2846, N2816);
nor NOR3 (N2847, N2846, N2807, N2821);
nand NAND2 (N2848, N2847, N1271);
and AND3 (N2849, N2841, N447, N672);
buf BUF1 (N2850, N2834);
nor NOR2 (N2851, N2849, N1699);
xor XOR2 (N2852, N2840, N380);
buf BUF1 (N2853, N2843);
buf BUF1 (N2854, N2850);
nor NOR2 (N2855, N2839, N2763);
xor XOR2 (N2856, N2835, N218);
not NOT1 (N2857, N2851);
buf BUF1 (N2858, N2845);
nor NOR2 (N2859, N2848, N1619);
or OR4 (N2860, N2858, N2466, N2255, N68);
not NOT1 (N2861, N2852);
buf BUF1 (N2862, N2857);
xor XOR2 (N2863, N2860, N421);
buf BUF1 (N2864, N2844);
not NOT1 (N2865, N2864);
and AND3 (N2866, N2862, N1554, N1284);
and AND4 (N2867, N2853, N2838, N901, N254);
and AND4 (N2868, N2854, N1139, N1824, N935);
and AND2 (N2869, N2805, N2542);
nand NAND4 (N2870, N2856, N1504, N2230, N783);
buf BUF1 (N2871, N2859);
nor NOR4 (N2872, N2867, N1490, N2526, N2488);
and AND3 (N2873, N2868, N1893, N1479);
and AND4 (N2874, N2865, N1640, N2678, N1487);
xor XOR2 (N2875, N2866, N2219);
nand NAND2 (N2876, N2869, N1866);
nor NOR2 (N2877, N2863, N513);
and AND3 (N2878, N2872, N1086, N1862);
nor NOR2 (N2879, N2870, N1159);
buf BUF1 (N2880, N2874);
buf BUF1 (N2881, N2878);
nor NOR3 (N2882, N2875, N1601, N1053);
nand NAND4 (N2883, N2880, N615, N1134, N9);
and AND4 (N2884, N2883, N712, N2293, N1101);
nand NAND3 (N2885, N2882, N1807, N2179);
or OR4 (N2886, N2877, N2076, N181, N876);
buf BUF1 (N2887, N2885);
buf BUF1 (N2888, N2879);
buf BUF1 (N2889, N2871);
nor NOR4 (N2890, N2888, N2666, N1022, N955);
nand NAND2 (N2891, N2887, N1789);
xor XOR2 (N2892, N2876, N1321);
nand NAND2 (N2893, N2861, N1196);
xor XOR2 (N2894, N2881, N703);
nor NOR2 (N2895, N2855, N911);
nand NAND3 (N2896, N2894, N2851, N505);
nor NOR4 (N2897, N2895, N1391, N2276, N1304);
nand NAND2 (N2898, N2873, N2007);
buf BUF1 (N2899, N2892);
buf BUF1 (N2900, N2890);
or OR4 (N2901, N2884, N1259, N2193, N1679);
nand NAND4 (N2902, N2900, N1195, N615, N2068);
xor XOR2 (N2903, N2899, N2440);
or OR3 (N2904, N2898, N1207, N2682);
xor XOR2 (N2905, N2901, N2566);
or OR3 (N2906, N2891, N1085, N924);
nand NAND4 (N2907, N2889, N1813, N533, N903);
buf BUF1 (N2908, N2902);
buf BUF1 (N2909, N2908);
xor XOR2 (N2910, N2904, N2019);
buf BUF1 (N2911, N2896);
and AND2 (N2912, N2897, N1957);
or OR2 (N2913, N2907, N2074);
nor NOR3 (N2914, N2909, N1926, N1640);
or OR3 (N2915, N2906, N2103, N1959);
xor XOR2 (N2916, N2912, N2767);
nor NOR4 (N2917, N2886, N111, N1119, N427);
nor NOR4 (N2918, N2893, N1937, N1898, N2869);
or OR3 (N2919, N2916, N1604, N2395);
nor NOR4 (N2920, N2915, N1918, N2698, N1938);
or OR4 (N2921, N2917, N2629, N861, N2531);
buf BUF1 (N2922, N2910);
nor NOR4 (N2923, N2921, N305, N1856, N517);
buf BUF1 (N2924, N2919);
nor NOR2 (N2925, N2911, N1859);
xor XOR2 (N2926, N2925, N1151);
and AND2 (N2927, N2903, N577);
or OR3 (N2928, N2914, N191, N2486);
not NOT1 (N2929, N2922);
nor NOR2 (N2930, N2923, N2434);
or OR4 (N2931, N2930, N83, N944, N876);
nor NOR4 (N2932, N2929, N1414, N328, N1657);
or OR3 (N2933, N2927, N1657, N2689);
not NOT1 (N2934, N2918);
not NOT1 (N2935, N2933);
and AND4 (N2936, N2934, N304, N105, N2095);
xor XOR2 (N2937, N2935, N2887);
or OR4 (N2938, N2905, N677, N1723, N2164);
not NOT1 (N2939, N2938);
nor NOR3 (N2940, N2939, N1998, N2680);
not NOT1 (N2941, N2940);
or OR2 (N2942, N2924, N1070);
xor XOR2 (N2943, N2913, N1274);
or OR3 (N2944, N2936, N723, N1716);
nor NOR2 (N2945, N2944, N1443);
buf BUF1 (N2946, N2943);
nor NOR3 (N2947, N2945, N1527, N2123);
nand NAND2 (N2948, N2931, N2261);
xor XOR2 (N2949, N2928, N1794);
xor XOR2 (N2950, N2932, N1239);
nand NAND4 (N2951, N2937, N437, N226, N2591);
nor NOR3 (N2952, N2950, N1825, N2279);
nand NAND3 (N2953, N2920, N597, N1999);
nand NAND2 (N2954, N2946, N1324);
xor XOR2 (N2955, N2947, N1429);
or OR3 (N2956, N2926, N956, N1565);
or OR3 (N2957, N2952, N2133, N1775);
xor XOR2 (N2958, N2942, N193);
buf BUF1 (N2959, N2953);
buf BUF1 (N2960, N2959);
buf BUF1 (N2961, N2949);
buf BUF1 (N2962, N2954);
and AND2 (N2963, N2956, N2008);
nor NOR3 (N2964, N2948, N2125, N1655);
and AND4 (N2965, N2964, N1677, N2114, N1830);
xor XOR2 (N2966, N2963, N808);
xor XOR2 (N2967, N2962, N1314);
buf BUF1 (N2968, N2955);
nor NOR3 (N2969, N2965, N2769, N679);
xor XOR2 (N2970, N2958, N812);
nor NOR2 (N2971, N2966, N1896);
not NOT1 (N2972, N2951);
and AND2 (N2973, N2957, N351);
or OR3 (N2974, N2972, N1991, N1103);
not NOT1 (N2975, N2960);
and AND3 (N2976, N2968, N934, N699);
buf BUF1 (N2977, N2976);
and AND4 (N2978, N2967, N2947, N471, N1837);
xor XOR2 (N2979, N2961, N1818);
nor NOR4 (N2980, N2974, N1454, N2647, N1882);
or OR4 (N2981, N2979, N1879, N2648, N2673);
nand NAND3 (N2982, N2971, N1422, N611);
or OR2 (N2983, N2982, N1258);
nand NAND3 (N2984, N2983, N2473, N1687);
or OR2 (N2985, N2970, N2274);
nand NAND3 (N2986, N2980, N1371, N116);
or OR4 (N2987, N2969, N2228, N348, N1011);
nand NAND4 (N2988, N2975, N1225, N1443, N2583);
nor NOR3 (N2989, N2941, N983, N2728);
buf BUF1 (N2990, N2981);
nand NAND4 (N2991, N2985, N1609, N1615, N874);
or OR2 (N2992, N2978, N2593);
xor XOR2 (N2993, N2984, N158);
nand NAND3 (N2994, N2977, N2438, N1977);
nand NAND3 (N2995, N2986, N1722, N1430);
nand NAND2 (N2996, N2988, N439);
and AND2 (N2997, N2994, N2643);
buf BUF1 (N2998, N2989);
buf BUF1 (N2999, N2993);
nand NAND4 (N3000, N2990, N56, N1742, N297);
or OR3 (N3001, N2987, N2810, N1985);
xor XOR2 (N3002, N3001, N541);
and AND3 (N3003, N2999, N1729, N1999);
nor NOR2 (N3004, N3000, N577);
not NOT1 (N3005, N2992);
nor NOR4 (N3006, N2991, N2433, N1503, N2600);
xor XOR2 (N3007, N3002, N2289);
nand NAND4 (N3008, N3004, N53, N2066, N1942);
or OR2 (N3009, N3005, N2430);
buf BUF1 (N3010, N2997);
not NOT1 (N3011, N3007);
nor NOR2 (N3012, N3003, N727);
or OR3 (N3013, N3010, N856, N1969);
or OR2 (N3014, N2973, N591);
buf BUF1 (N3015, N2998);
not NOT1 (N3016, N3012);
xor XOR2 (N3017, N2996, N1390);
nand NAND2 (N3018, N2995, N2263);
nor NOR2 (N3019, N3011, N2466);
and AND2 (N3020, N3019, N2482);
or OR4 (N3021, N3017, N1031, N2496, N378);
xor XOR2 (N3022, N3020, N1754);
xor XOR2 (N3023, N3021, N1870);
endmodule