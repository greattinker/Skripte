// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19;

output N4015,N4014,N4009,N4016,N4000,N4007,N4018,N4011,N3997,N4019;

xor XOR2 (N20, N5, N15);
nand NAND2 (N21, N12, N13);
xor XOR2 (N22, N14, N5);
nand NAND2 (N23, N17, N3);
buf BUF1 (N24, N22);
nand NAND4 (N25, N8, N17, N13, N20);
not NOT1 (N26, N7);
and AND3 (N27, N6, N7, N21);
or OR4 (N28, N16, N12, N13, N3);
xor XOR2 (N29, N11, N28);
or OR3 (N30, N28, N19, N6);
buf BUF1 (N31, N27);
and AND2 (N32, N21, N8);
xor XOR2 (N33, N15, N6);
nor NOR2 (N34, N5, N25);
nor NOR3 (N35, N6, N12, N1);
buf BUF1 (N36, N29);
or OR3 (N37, N30, N3, N23);
or OR4 (N38, N13, N29, N5, N29);
xor XOR2 (N39, N26, N26);
or OR3 (N40, N36, N34, N21);
and AND4 (N41, N24, N39, N18, N9);
nor NOR2 (N42, N39, N41);
xor XOR2 (N43, N11, N26);
and AND3 (N44, N18, N4, N11);
not NOT1 (N45, N42);
not NOT1 (N46, N38);
or OR2 (N47, N32, N25);
not NOT1 (N48, N47);
nand NAND3 (N49, N45, N20, N48);
nand NAND4 (N50, N31, N10, N7, N48);
not NOT1 (N51, N34);
nor NOR2 (N52, N33, N4);
buf BUF1 (N53, N43);
nand NAND3 (N54, N46, N45, N6);
buf BUF1 (N55, N51);
buf BUF1 (N56, N35);
buf BUF1 (N57, N37);
or OR3 (N58, N50, N33, N29);
or OR2 (N59, N49, N47);
or OR4 (N60, N58, N21, N26, N36);
and AND2 (N61, N44, N22);
buf BUF1 (N62, N61);
nor NOR4 (N63, N54, N48, N50, N20);
buf BUF1 (N64, N55);
nand NAND2 (N65, N60, N55);
not NOT1 (N66, N65);
xor XOR2 (N67, N56, N6);
nor NOR2 (N68, N62, N33);
or OR4 (N69, N57, N36, N26, N31);
nand NAND2 (N70, N66, N35);
nand NAND4 (N71, N67, N22, N43, N19);
nand NAND3 (N72, N59, N48, N54);
not NOT1 (N73, N40);
or OR3 (N74, N63, N37, N10);
not NOT1 (N75, N52);
or OR4 (N76, N75, N19, N1, N11);
or OR4 (N77, N76, N10, N43, N20);
and AND4 (N78, N74, N21, N66, N38);
nor NOR4 (N79, N73, N47, N32, N77);
and AND3 (N80, N18, N21, N20);
nand NAND2 (N81, N72, N3);
or OR2 (N82, N64, N65);
nand NAND4 (N83, N70, N73, N17, N23);
or OR3 (N84, N81, N59, N61);
and AND2 (N85, N68, N52);
nand NAND2 (N86, N79, N23);
buf BUF1 (N87, N82);
nor NOR3 (N88, N87, N12, N43);
not NOT1 (N89, N86);
nor NOR4 (N90, N80, N44, N74, N30);
or OR3 (N91, N78, N9, N27);
not NOT1 (N92, N91);
nor NOR2 (N93, N53, N46);
or OR2 (N94, N69, N57);
buf BUF1 (N95, N90);
xor XOR2 (N96, N93, N87);
nor NOR2 (N97, N85, N27);
nand NAND2 (N98, N96, N88);
not NOT1 (N99, N33);
or OR3 (N100, N84, N20, N5);
nor NOR3 (N101, N92, N55, N39);
nor NOR3 (N102, N71, N53, N53);
not NOT1 (N103, N89);
and AND3 (N104, N94, N82, N27);
and AND3 (N105, N101, N60, N76);
nor NOR2 (N106, N83, N54);
or OR2 (N107, N99, N63);
and AND4 (N108, N95, N15, N48, N103);
nor NOR4 (N109, N2, N15, N10, N58);
nor NOR2 (N110, N108, N77);
xor XOR2 (N111, N106, N83);
nor NOR2 (N112, N104, N79);
xor XOR2 (N113, N111, N47);
xor XOR2 (N114, N97, N54);
not NOT1 (N115, N109);
buf BUF1 (N116, N105);
nor NOR2 (N117, N116, N62);
xor XOR2 (N118, N117, N21);
buf BUF1 (N119, N100);
and AND3 (N120, N98, N94, N64);
and AND3 (N121, N110, N101, N1);
or OR2 (N122, N102, N34);
and AND2 (N123, N120, N48);
not NOT1 (N124, N123);
buf BUF1 (N125, N122);
nand NAND3 (N126, N114, N95, N52);
and AND4 (N127, N112, N92, N113, N109);
or OR3 (N128, N73, N29, N88);
xor XOR2 (N129, N121, N18);
and AND4 (N130, N128, N86, N99, N110);
nand NAND2 (N131, N107, N49);
nor NOR2 (N132, N127, N31);
xor XOR2 (N133, N118, N102);
and AND3 (N134, N132, N123, N35);
buf BUF1 (N135, N130);
nand NAND2 (N136, N125, N87);
or OR4 (N137, N133, N26, N54, N18);
nand NAND2 (N138, N126, N62);
and AND2 (N139, N137, N63);
and AND3 (N140, N135, N139, N40);
not NOT1 (N141, N80);
not NOT1 (N142, N115);
buf BUF1 (N143, N131);
xor XOR2 (N144, N119, N89);
buf BUF1 (N145, N124);
not NOT1 (N146, N145);
nor NOR4 (N147, N134, N25, N66, N12);
nor NOR2 (N148, N136, N115);
and AND2 (N149, N144, N89);
nand NAND3 (N150, N138, N149, N97);
or OR3 (N151, N127, N19, N116);
or OR3 (N152, N141, N139, N8);
not NOT1 (N153, N143);
not NOT1 (N154, N129);
and AND3 (N155, N146, N86, N26);
xor XOR2 (N156, N153, N112);
not NOT1 (N157, N155);
buf BUF1 (N158, N154);
or OR2 (N159, N152, N150);
nor NOR4 (N160, N5, N37, N28, N91);
buf BUF1 (N161, N140);
not NOT1 (N162, N160);
buf BUF1 (N163, N142);
nor NOR3 (N164, N162, N162, N134);
or OR2 (N165, N147, N2);
nand NAND3 (N166, N163, N65, N17);
or OR2 (N167, N156, N9);
nand NAND4 (N168, N148, N92, N103, N97);
nor NOR4 (N169, N158, N136, N45, N124);
and AND4 (N170, N165, N54, N139, N47);
not NOT1 (N171, N167);
xor XOR2 (N172, N171, N29);
and AND2 (N173, N151, N35);
xor XOR2 (N174, N157, N22);
nand NAND4 (N175, N166, N9, N24, N152);
xor XOR2 (N176, N173, N140);
buf BUF1 (N177, N174);
buf BUF1 (N178, N159);
or OR2 (N179, N172, N98);
not NOT1 (N180, N170);
buf BUF1 (N181, N164);
buf BUF1 (N182, N180);
buf BUF1 (N183, N177);
xor XOR2 (N184, N183, N31);
buf BUF1 (N185, N182);
or OR4 (N186, N168, N117, N8, N62);
nand NAND2 (N187, N176, N116);
not NOT1 (N188, N179);
not NOT1 (N189, N161);
nor NOR4 (N190, N189, N145, N101, N40);
nor NOR2 (N191, N184, N89);
nand NAND3 (N192, N178, N52, N152);
nand NAND2 (N193, N188, N164);
and AND3 (N194, N187, N105, N124);
nor NOR2 (N195, N192, N126);
and AND3 (N196, N186, N49, N67);
xor XOR2 (N197, N196, N99);
nand NAND2 (N198, N195, N137);
and AND3 (N199, N175, N42, N154);
nand NAND4 (N200, N185, N153, N178, N178);
and AND2 (N201, N169, N147);
or OR3 (N202, N181, N90, N1);
xor XOR2 (N203, N200, N85);
nand NAND3 (N204, N191, N164, N78);
and AND3 (N205, N202, N182, N136);
nor NOR4 (N206, N201, N104, N119, N55);
or OR3 (N207, N204, N203, N118);
xor XOR2 (N208, N8, N53);
xor XOR2 (N209, N198, N123);
or OR4 (N210, N206, N121, N206, N164);
nor NOR3 (N211, N199, N180, N14);
not NOT1 (N212, N190);
nand NAND3 (N213, N205, N200, N4);
xor XOR2 (N214, N193, N128);
nor NOR4 (N215, N208, N93, N74, N180);
nand NAND3 (N216, N212, N84, N183);
xor XOR2 (N217, N194, N142);
and AND2 (N218, N211, N170);
not NOT1 (N219, N215);
and AND3 (N220, N210, N65, N165);
and AND2 (N221, N213, N185);
xor XOR2 (N222, N197, N99);
xor XOR2 (N223, N218, N79);
nor NOR4 (N224, N207, N215, N190, N54);
nand NAND3 (N225, N224, N51, N3);
nor NOR4 (N226, N209, N183, N199, N29);
xor XOR2 (N227, N223, N138);
nor NOR2 (N228, N219, N169);
nand NAND3 (N229, N217, N31, N128);
and AND2 (N230, N228, N77);
nand NAND4 (N231, N225, N160, N40, N178);
buf BUF1 (N232, N229);
nand NAND3 (N233, N222, N177, N12);
and AND3 (N234, N221, N176, N53);
and AND3 (N235, N234, N5, N7);
not NOT1 (N236, N227);
and AND2 (N237, N230, N99);
nor NOR3 (N238, N237, N23, N16);
not NOT1 (N239, N232);
or OR3 (N240, N233, N20, N199);
or OR3 (N241, N226, N203, N187);
buf BUF1 (N242, N238);
or OR3 (N243, N236, N236, N15);
and AND4 (N244, N216, N179, N232, N152);
not NOT1 (N245, N241);
nand NAND2 (N246, N240, N23);
and AND4 (N247, N246, N185, N188, N130);
not NOT1 (N248, N243);
or OR4 (N249, N242, N156, N112, N47);
not NOT1 (N250, N231);
nand NAND3 (N251, N249, N81, N109);
nand NAND3 (N252, N235, N118, N181);
and AND3 (N253, N244, N165, N24);
not NOT1 (N254, N252);
nand NAND2 (N255, N239, N176);
not NOT1 (N256, N214);
or OR2 (N257, N248, N44);
not NOT1 (N258, N245);
not NOT1 (N259, N220);
or OR4 (N260, N251, N248, N82, N192);
nor NOR3 (N261, N247, N147, N123);
and AND4 (N262, N261, N158, N131, N18);
and AND3 (N263, N256, N79, N159);
nand NAND4 (N264, N250, N130, N67, N194);
buf BUF1 (N265, N255);
nand NAND3 (N266, N257, N76, N232);
nand NAND4 (N267, N263, N219, N193, N31);
nor NOR3 (N268, N253, N44, N129);
not NOT1 (N269, N266);
and AND4 (N270, N264, N13, N90, N55);
nor NOR4 (N271, N265, N216, N74, N179);
not NOT1 (N272, N269);
or OR2 (N273, N262, N184);
or OR3 (N274, N254, N40, N82);
buf BUF1 (N275, N258);
not NOT1 (N276, N259);
nand NAND4 (N277, N274, N60, N254, N48);
buf BUF1 (N278, N277);
not NOT1 (N279, N268);
not NOT1 (N280, N278);
nand NAND3 (N281, N280, N260, N127);
or OR4 (N282, N153, N159, N277, N127);
nor NOR2 (N283, N276, N199);
nand NAND2 (N284, N273, N136);
nand NAND4 (N285, N275, N56, N256, N91);
not NOT1 (N286, N285);
nor NOR4 (N287, N281, N207, N151, N187);
xor XOR2 (N288, N272, N287);
nor NOR3 (N289, N243, N254, N2);
and AND2 (N290, N289, N283);
or OR3 (N291, N277, N167, N141);
and AND3 (N292, N286, N214, N275);
or OR4 (N293, N267, N23, N63, N234);
buf BUF1 (N294, N284);
buf BUF1 (N295, N282);
buf BUF1 (N296, N271);
nor NOR2 (N297, N291, N164);
nor NOR2 (N298, N293, N118);
not NOT1 (N299, N279);
or OR4 (N300, N290, N207, N126, N185);
buf BUF1 (N301, N295);
and AND3 (N302, N294, N212, N57);
buf BUF1 (N303, N302);
nand NAND4 (N304, N270, N91, N270, N204);
nand NAND2 (N305, N299, N293);
buf BUF1 (N306, N298);
buf BUF1 (N307, N303);
nand NAND2 (N308, N292, N2);
xor XOR2 (N309, N300, N90);
and AND3 (N310, N288, N89, N131);
and AND4 (N311, N297, N126, N136, N171);
nand NAND3 (N312, N308, N268, N137);
nand NAND2 (N313, N304, N144);
nand NAND3 (N314, N296, N310, N37);
or OR4 (N315, N37, N74, N139, N234);
not NOT1 (N316, N312);
nand NAND4 (N317, N313, N171, N35, N103);
or OR3 (N318, N301, N151, N105);
nor NOR3 (N319, N318, N200, N211);
buf BUF1 (N320, N314);
not NOT1 (N321, N320);
and AND3 (N322, N309, N178, N292);
nand NAND4 (N323, N321, N119, N128, N202);
buf BUF1 (N324, N317);
nand NAND3 (N325, N323, N161, N36);
and AND3 (N326, N305, N269, N301);
and AND3 (N327, N311, N321, N137);
or OR3 (N328, N307, N291, N59);
nor NOR2 (N329, N319, N311);
nand NAND3 (N330, N326, N146, N92);
not NOT1 (N331, N315);
nor NOR2 (N332, N328, N233);
nand NAND3 (N333, N316, N272, N98);
nor NOR4 (N334, N332, N134, N176, N218);
nand NAND3 (N335, N324, N208, N60);
not NOT1 (N336, N322);
xor XOR2 (N337, N329, N221);
or OR4 (N338, N333, N212, N307, N130);
or OR2 (N339, N325, N273);
nor NOR3 (N340, N337, N178, N32);
nand NAND3 (N341, N327, N232, N322);
nand NAND2 (N342, N335, N118);
or OR3 (N343, N306, N187, N55);
or OR4 (N344, N343, N50, N335, N322);
nor NOR3 (N345, N339, N250, N4);
xor XOR2 (N346, N344, N139);
nand NAND4 (N347, N346, N244, N86, N91);
or OR2 (N348, N336, N151);
not NOT1 (N349, N348);
or OR4 (N350, N334, N226, N189, N335);
xor XOR2 (N351, N347, N340);
or OR4 (N352, N71, N186, N34, N110);
nor NOR4 (N353, N352, N81, N328, N204);
xor XOR2 (N354, N342, N289);
and AND2 (N355, N354, N302);
not NOT1 (N356, N350);
xor XOR2 (N357, N355, N50);
nor NOR4 (N358, N330, N95, N210, N113);
buf BUF1 (N359, N345);
or OR3 (N360, N356, N217, N51);
or OR4 (N361, N338, N134, N41, N189);
xor XOR2 (N362, N349, N326);
nor NOR2 (N363, N358, N185);
not NOT1 (N364, N361);
not NOT1 (N365, N362);
or OR4 (N366, N353, N110, N285, N180);
xor XOR2 (N367, N365, N2);
xor XOR2 (N368, N357, N195);
or OR2 (N369, N341, N81);
buf BUF1 (N370, N369);
xor XOR2 (N371, N364, N100);
or OR3 (N372, N371, N295, N360);
or OR4 (N373, N11, N232, N120, N239);
and AND3 (N374, N366, N50, N82);
or OR2 (N375, N363, N60);
xor XOR2 (N376, N359, N57);
nand NAND2 (N377, N351, N141);
or OR2 (N378, N377, N142);
and AND3 (N379, N372, N212, N250);
or OR4 (N380, N379, N134, N306, N111);
buf BUF1 (N381, N376);
nand NAND4 (N382, N378, N230, N297, N343);
xor XOR2 (N383, N375, N52);
xor XOR2 (N384, N331, N196);
xor XOR2 (N385, N384, N243);
or OR2 (N386, N370, N315);
or OR3 (N387, N386, N37, N135);
buf BUF1 (N388, N381);
not NOT1 (N389, N367);
or OR3 (N390, N387, N62, N101);
xor XOR2 (N391, N374, N237);
not NOT1 (N392, N382);
or OR2 (N393, N390, N357);
nand NAND3 (N394, N393, N2, N58);
and AND2 (N395, N380, N199);
buf BUF1 (N396, N373);
not NOT1 (N397, N383);
not NOT1 (N398, N397);
buf BUF1 (N399, N385);
or OR4 (N400, N398, N23, N249, N85);
not NOT1 (N401, N396);
nor NOR2 (N402, N391, N127);
buf BUF1 (N403, N388);
and AND4 (N404, N401, N331, N342, N28);
or OR2 (N405, N394, N385);
xor XOR2 (N406, N368, N251);
not NOT1 (N407, N403);
xor XOR2 (N408, N404, N72);
nor NOR3 (N409, N402, N292, N50);
or OR2 (N410, N405, N337);
or OR4 (N411, N408, N308, N278, N160);
or OR4 (N412, N389, N348, N249, N360);
nand NAND2 (N413, N407, N2);
and AND4 (N414, N410, N305, N178, N175);
buf BUF1 (N415, N395);
or OR4 (N416, N415, N123, N410, N95);
or OR2 (N417, N409, N107);
and AND4 (N418, N392, N96, N401, N173);
nand NAND2 (N419, N417, N304);
xor XOR2 (N420, N412, N238);
and AND3 (N421, N400, N366, N384);
nor NOR2 (N422, N406, N274);
xor XOR2 (N423, N420, N272);
nor NOR4 (N424, N416, N163, N146, N156);
xor XOR2 (N425, N413, N157);
nor NOR4 (N426, N424, N323, N235, N197);
nor NOR4 (N427, N411, N45, N252, N29);
or OR3 (N428, N421, N11, N101);
not NOT1 (N429, N418);
buf BUF1 (N430, N427);
and AND4 (N431, N399, N28, N365, N82);
xor XOR2 (N432, N430, N224);
not NOT1 (N433, N425);
or OR2 (N434, N428, N239);
xor XOR2 (N435, N434, N410);
nand NAND4 (N436, N426, N63, N130, N192);
xor XOR2 (N437, N432, N431);
and AND2 (N438, N86, N376);
or OR4 (N439, N438, N116, N229, N436);
nand NAND2 (N440, N3, N188);
buf BUF1 (N441, N414);
not NOT1 (N442, N435);
xor XOR2 (N443, N439, N19);
nor NOR3 (N444, N437, N187, N106);
and AND2 (N445, N443, N393);
or OR4 (N446, N422, N118, N325, N269);
xor XOR2 (N447, N419, N401);
nor NOR2 (N448, N441, N340);
and AND2 (N449, N423, N368);
or OR2 (N450, N444, N385);
or OR4 (N451, N429, N384, N307, N416);
xor XOR2 (N452, N447, N385);
and AND3 (N453, N452, N274, N435);
and AND4 (N454, N451, N219, N47, N335);
nor NOR3 (N455, N445, N181, N88);
xor XOR2 (N456, N449, N6);
nand NAND2 (N457, N453, N219);
buf BUF1 (N458, N457);
not NOT1 (N459, N440);
not NOT1 (N460, N442);
and AND3 (N461, N454, N179, N129);
not NOT1 (N462, N460);
or OR2 (N463, N462, N221);
nand NAND2 (N464, N459, N386);
nor NOR2 (N465, N463, N23);
and AND2 (N466, N446, N391);
nor NOR4 (N467, N433, N290, N465, N371);
nor NOR4 (N468, N363, N406, N200, N69);
and AND2 (N469, N448, N350);
nor NOR4 (N470, N455, N69, N425, N36);
not NOT1 (N471, N469);
or OR4 (N472, N450, N75, N373, N248);
and AND3 (N473, N456, N139, N422);
or OR2 (N474, N464, N292);
not NOT1 (N475, N467);
nor NOR3 (N476, N458, N416, N360);
buf BUF1 (N477, N476);
or OR3 (N478, N472, N45, N9);
buf BUF1 (N479, N461);
buf BUF1 (N480, N474);
not NOT1 (N481, N471);
and AND2 (N482, N481, N2);
xor XOR2 (N483, N475, N377);
nor NOR3 (N484, N479, N400, N132);
or OR4 (N485, N480, N262, N295, N155);
and AND2 (N486, N478, N187);
and AND4 (N487, N485, N70, N220, N58);
not NOT1 (N488, N477);
and AND2 (N489, N488, N35);
or OR2 (N490, N470, N295);
nand NAND2 (N491, N484, N322);
not NOT1 (N492, N468);
not NOT1 (N493, N482);
and AND4 (N494, N466, N59, N438, N412);
or OR4 (N495, N492, N459, N359, N374);
not NOT1 (N496, N489);
or OR4 (N497, N493, N23, N392, N226);
xor XOR2 (N498, N491, N123);
nor NOR4 (N499, N487, N282, N179, N330);
buf BUF1 (N500, N483);
buf BUF1 (N501, N499);
not NOT1 (N502, N495);
or OR3 (N503, N501, N167, N44);
xor XOR2 (N504, N497, N286);
buf BUF1 (N505, N502);
nand NAND3 (N506, N498, N399, N229);
buf BUF1 (N507, N490);
nor NOR4 (N508, N507, N199, N62, N278);
nand NAND2 (N509, N504, N264);
or OR4 (N510, N486, N354, N435, N257);
buf BUF1 (N511, N509);
buf BUF1 (N512, N494);
not NOT1 (N513, N510);
nor NOR2 (N514, N506, N275);
not NOT1 (N515, N473);
and AND2 (N516, N508, N511);
or OR3 (N517, N63, N141, N155);
not NOT1 (N518, N512);
buf BUF1 (N519, N516);
nor NOR4 (N520, N519, N341, N454, N255);
or OR4 (N521, N505, N315, N120, N344);
and AND2 (N522, N521, N485);
nor NOR4 (N523, N517, N243, N67, N79);
or OR3 (N524, N503, N251, N349);
buf BUF1 (N525, N523);
or OR3 (N526, N514, N362, N191);
nor NOR3 (N527, N513, N29, N25);
xor XOR2 (N528, N496, N61);
nand NAND3 (N529, N520, N388, N57);
nand NAND4 (N530, N528, N451, N519, N453);
nand NAND2 (N531, N527, N461);
or OR2 (N532, N515, N37);
and AND2 (N533, N531, N296);
and AND3 (N534, N524, N241, N504);
and AND3 (N535, N522, N191, N6);
nand NAND3 (N536, N500, N248, N435);
and AND2 (N537, N530, N356);
nor NOR2 (N538, N536, N309);
or OR3 (N539, N529, N455, N177);
or OR2 (N540, N533, N104);
not NOT1 (N541, N518);
nor NOR3 (N542, N541, N62, N49);
nand NAND4 (N543, N537, N174, N43, N171);
buf BUF1 (N544, N540);
buf BUF1 (N545, N538);
not NOT1 (N546, N543);
nor NOR3 (N547, N544, N441, N456);
or OR2 (N548, N534, N130);
nor NOR4 (N549, N535, N140, N148, N302);
and AND2 (N550, N526, N21);
or OR3 (N551, N548, N322, N171);
buf BUF1 (N552, N550);
nand NAND2 (N553, N549, N217);
buf BUF1 (N554, N545);
xor XOR2 (N555, N525, N370);
not NOT1 (N556, N553);
xor XOR2 (N557, N546, N255);
xor XOR2 (N558, N547, N198);
and AND4 (N559, N558, N266, N262, N391);
nand NAND4 (N560, N555, N318, N261, N505);
buf BUF1 (N561, N532);
not NOT1 (N562, N557);
or OR3 (N563, N554, N240, N330);
or OR4 (N564, N551, N525, N136, N346);
and AND2 (N565, N562, N450);
buf BUF1 (N566, N552);
not NOT1 (N567, N556);
buf BUF1 (N568, N539);
not NOT1 (N569, N560);
nand NAND3 (N570, N569, N479, N491);
and AND2 (N571, N564, N349);
or OR4 (N572, N570, N454, N174, N37);
nor NOR3 (N573, N559, N439, N23);
buf BUF1 (N574, N571);
xor XOR2 (N575, N561, N170);
nor NOR4 (N576, N572, N510, N248, N287);
xor XOR2 (N577, N574, N96);
nor NOR4 (N578, N577, N511, N24, N311);
xor XOR2 (N579, N542, N382);
and AND4 (N580, N568, N482, N25, N55);
not NOT1 (N581, N580);
buf BUF1 (N582, N573);
nand NAND3 (N583, N581, N554, N348);
not NOT1 (N584, N575);
nor NOR2 (N585, N563, N380);
xor XOR2 (N586, N566, N516);
or OR4 (N587, N579, N54, N12, N214);
not NOT1 (N588, N567);
not NOT1 (N589, N565);
xor XOR2 (N590, N578, N307);
buf BUF1 (N591, N589);
or OR3 (N592, N591, N557, N104);
or OR4 (N593, N587, N329, N186, N29);
xor XOR2 (N594, N590, N554);
buf BUF1 (N595, N592);
xor XOR2 (N596, N585, N418);
xor XOR2 (N597, N584, N501);
or OR2 (N598, N597, N248);
or OR4 (N599, N595, N16, N477, N361);
nand NAND4 (N600, N588, N118, N480, N431);
or OR3 (N601, N598, N109, N209);
not NOT1 (N602, N583);
and AND3 (N603, N582, N169, N446);
and AND2 (N604, N594, N364);
nor NOR4 (N605, N602, N136, N549, N171);
xor XOR2 (N606, N586, N483);
and AND4 (N607, N599, N516, N389, N181);
nor NOR4 (N608, N607, N85, N303, N409);
or OR3 (N609, N604, N278, N47);
and AND2 (N610, N601, N315);
nand NAND3 (N611, N609, N597, N36);
nor NOR2 (N612, N608, N355);
not NOT1 (N613, N603);
or OR2 (N614, N610, N554);
nand NAND4 (N615, N611, N493, N513, N249);
not NOT1 (N616, N593);
or OR2 (N617, N605, N41);
nand NAND4 (N618, N576, N128, N255, N302);
and AND2 (N619, N617, N516);
or OR2 (N620, N615, N365);
and AND3 (N621, N600, N55, N586);
nor NOR3 (N622, N606, N587, N17);
or OR2 (N623, N616, N372);
xor XOR2 (N624, N619, N505);
or OR3 (N625, N612, N553, N494);
not NOT1 (N626, N623);
nand NAND4 (N627, N624, N318, N333, N412);
not NOT1 (N628, N622);
nor NOR2 (N629, N618, N551);
or OR4 (N630, N629, N582, N130, N237);
and AND4 (N631, N626, N346, N517, N188);
or OR4 (N632, N621, N86, N141, N537);
nand NAND3 (N633, N632, N432, N174);
not NOT1 (N634, N614);
not NOT1 (N635, N625);
nand NAND4 (N636, N620, N454, N248, N450);
xor XOR2 (N637, N631, N558);
nand NAND4 (N638, N633, N81, N30, N180);
nor NOR4 (N639, N630, N411, N448, N561);
nand NAND3 (N640, N636, N480, N525);
nor NOR3 (N641, N635, N438, N633);
xor XOR2 (N642, N627, N404);
buf BUF1 (N643, N637);
xor XOR2 (N644, N642, N259);
nor NOR3 (N645, N596, N404, N431);
nor NOR3 (N646, N644, N25, N144);
nand NAND2 (N647, N646, N279);
xor XOR2 (N648, N613, N618);
and AND2 (N649, N638, N118);
not NOT1 (N650, N648);
xor XOR2 (N651, N649, N333);
nor NOR2 (N652, N628, N75);
nand NAND2 (N653, N639, N127);
nand NAND4 (N654, N643, N325, N585, N320);
xor XOR2 (N655, N645, N602);
xor XOR2 (N656, N654, N108);
nand NAND2 (N657, N634, N468);
and AND2 (N658, N647, N568);
nor NOR3 (N659, N641, N431, N283);
not NOT1 (N660, N657);
nand NAND4 (N661, N650, N606, N215, N117);
or OR3 (N662, N655, N65, N520);
not NOT1 (N663, N640);
buf BUF1 (N664, N663);
nor NOR4 (N665, N656, N590, N547, N378);
buf BUF1 (N666, N651);
nor NOR4 (N667, N665, N311, N204, N393);
nand NAND3 (N668, N658, N474, N331);
not NOT1 (N669, N664);
and AND4 (N670, N652, N67, N553, N15);
not NOT1 (N671, N653);
or OR4 (N672, N659, N507, N664, N297);
not NOT1 (N673, N667);
buf BUF1 (N674, N670);
nor NOR3 (N675, N662, N543, N368);
xor XOR2 (N676, N671, N427);
nor NOR3 (N677, N669, N119, N366);
nand NAND3 (N678, N666, N286, N296);
not NOT1 (N679, N674);
and AND4 (N680, N668, N129, N131, N16);
or OR2 (N681, N677, N318);
buf BUF1 (N682, N680);
nor NOR2 (N683, N676, N533);
and AND3 (N684, N679, N386, N644);
xor XOR2 (N685, N682, N596);
xor XOR2 (N686, N673, N646);
not NOT1 (N687, N660);
or OR3 (N688, N672, N562, N132);
xor XOR2 (N689, N685, N582);
not NOT1 (N690, N678);
and AND2 (N691, N683, N532);
nor NOR4 (N692, N688, N160, N386, N578);
or OR3 (N693, N691, N142, N93);
xor XOR2 (N694, N693, N509);
and AND4 (N695, N689, N181, N310, N666);
buf BUF1 (N696, N690);
xor XOR2 (N697, N695, N125);
xor XOR2 (N698, N686, N289);
buf BUF1 (N699, N696);
nor NOR2 (N700, N694, N565);
nor NOR4 (N701, N699, N193, N343, N125);
not NOT1 (N702, N687);
buf BUF1 (N703, N692);
nand NAND2 (N704, N675, N105);
and AND4 (N705, N684, N381, N688, N138);
nor NOR2 (N706, N698, N611);
xor XOR2 (N707, N703, N580);
and AND3 (N708, N706, N497, N56);
nand NAND3 (N709, N705, N327, N282);
nor NOR2 (N710, N697, N598);
not NOT1 (N711, N704);
not NOT1 (N712, N700);
xor XOR2 (N713, N701, N116);
buf BUF1 (N714, N707);
nor NOR2 (N715, N713, N464);
nor NOR3 (N716, N715, N25, N294);
or OR3 (N717, N661, N677, N280);
and AND2 (N718, N714, N553);
xor XOR2 (N719, N708, N252);
and AND3 (N720, N710, N164, N521);
xor XOR2 (N721, N709, N636);
nor NOR2 (N722, N717, N607);
and AND2 (N723, N722, N182);
nor NOR3 (N724, N719, N551, N435);
and AND2 (N725, N718, N360);
buf BUF1 (N726, N723);
nand NAND2 (N727, N681, N660);
nor NOR2 (N728, N721, N522);
or OR4 (N729, N711, N664, N310, N646);
not NOT1 (N730, N725);
not NOT1 (N731, N724);
and AND3 (N732, N731, N335, N291);
xor XOR2 (N733, N728, N291);
and AND4 (N734, N729, N430, N511, N260);
nor NOR2 (N735, N732, N425);
buf BUF1 (N736, N734);
nor NOR3 (N737, N730, N87, N325);
not NOT1 (N738, N735);
or OR4 (N739, N733, N325, N36, N48);
and AND2 (N740, N736, N489);
nand NAND4 (N741, N727, N667, N276, N68);
not NOT1 (N742, N716);
or OR4 (N743, N739, N131, N531, N260);
or OR2 (N744, N712, N63);
buf BUF1 (N745, N702);
buf BUF1 (N746, N743);
not NOT1 (N747, N738);
or OR4 (N748, N747, N98, N562, N201);
buf BUF1 (N749, N748);
not NOT1 (N750, N740);
nand NAND3 (N751, N749, N258, N309);
nand NAND2 (N752, N720, N644);
or OR2 (N753, N752, N169);
nand NAND3 (N754, N751, N738, N103);
buf BUF1 (N755, N750);
nor NOR2 (N756, N741, N314);
buf BUF1 (N757, N744);
buf BUF1 (N758, N755);
buf BUF1 (N759, N757);
and AND2 (N760, N745, N538);
nand NAND3 (N761, N758, N214, N120);
and AND3 (N762, N726, N557, N751);
and AND3 (N763, N737, N684, N317);
and AND2 (N764, N753, N175);
xor XOR2 (N765, N763, N430);
not NOT1 (N766, N759);
xor XOR2 (N767, N761, N759);
not NOT1 (N768, N760);
buf BUF1 (N769, N762);
or OR2 (N770, N746, N45);
and AND3 (N771, N742, N447, N205);
or OR2 (N772, N769, N31);
nand NAND3 (N773, N765, N484, N261);
nor NOR4 (N774, N768, N64, N506, N737);
not NOT1 (N775, N772);
nand NAND4 (N776, N774, N570, N560, N171);
not NOT1 (N777, N770);
not NOT1 (N778, N764);
nand NAND3 (N779, N771, N661, N270);
not NOT1 (N780, N754);
buf BUF1 (N781, N773);
nand NAND3 (N782, N778, N603, N494);
buf BUF1 (N783, N767);
not NOT1 (N784, N756);
nand NAND4 (N785, N777, N320, N522, N286);
not NOT1 (N786, N779);
or OR2 (N787, N783, N311);
xor XOR2 (N788, N775, N309);
and AND2 (N789, N776, N403);
xor XOR2 (N790, N786, N290);
not NOT1 (N791, N766);
and AND2 (N792, N791, N56);
nand NAND4 (N793, N787, N132, N750, N451);
not NOT1 (N794, N780);
xor XOR2 (N795, N784, N614);
or OR3 (N796, N781, N574, N223);
xor XOR2 (N797, N792, N710);
buf BUF1 (N798, N795);
xor XOR2 (N799, N798, N475);
not NOT1 (N800, N797);
and AND4 (N801, N794, N269, N373, N580);
not NOT1 (N802, N796);
and AND4 (N803, N785, N591, N209, N110);
buf BUF1 (N804, N801);
nand NAND3 (N805, N803, N695, N496);
not NOT1 (N806, N799);
and AND3 (N807, N806, N499, N620);
or OR3 (N808, N782, N518, N398);
xor XOR2 (N809, N808, N417);
not NOT1 (N810, N790);
or OR2 (N811, N789, N300);
and AND4 (N812, N809, N465, N138, N494);
xor XOR2 (N813, N812, N368);
or OR2 (N814, N813, N663);
nand NAND3 (N815, N814, N374, N448);
buf BUF1 (N816, N810);
xor XOR2 (N817, N804, N178);
nand NAND2 (N818, N800, N627);
nor NOR4 (N819, N818, N31, N655, N625);
not NOT1 (N820, N807);
xor XOR2 (N821, N811, N551);
and AND4 (N822, N821, N388, N53, N304);
nor NOR2 (N823, N817, N603);
not NOT1 (N824, N788);
or OR2 (N825, N805, N200);
nand NAND3 (N826, N823, N105, N343);
and AND3 (N827, N822, N84, N665);
or OR4 (N828, N820, N798, N65, N427);
or OR2 (N829, N828, N634);
and AND3 (N830, N827, N689, N715);
or OR2 (N831, N802, N803);
or OR2 (N832, N825, N469);
not NOT1 (N833, N829);
nand NAND2 (N834, N826, N140);
or OR2 (N835, N816, N687);
not NOT1 (N836, N834);
or OR3 (N837, N830, N188, N777);
and AND2 (N838, N824, N329);
buf BUF1 (N839, N832);
nand NAND2 (N840, N815, N544);
nor NOR2 (N841, N836, N687);
xor XOR2 (N842, N837, N633);
buf BUF1 (N843, N840);
buf BUF1 (N844, N831);
buf BUF1 (N845, N839);
or OR3 (N846, N844, N315, N85);
not NOT1 (N847, N833);
buf BUF1 (N848, N819);
buf BUF1 (N849, N845);
buf BUF1 (N850, N838);
and AND3 (N851, N850, N342, N601);
not NOT1 (N852, N846);
not NOT1 (N853, N851);
xor XOR2 (N854, N848, N785);
or OR4 (N855, N847, N608, N352, N596);
buf BUF1 (N856, N854);
nand NAND2 (N857, N852, N424);
buf BUF1 (N858, N857);
nand NAND3 (N859, N858, N119, N567);
xor XOR2 (N860, N849, N791);
buf BUF1 (N861, N855);
nand NAND3 (N862, N842, N80, N521);
buf BUF1 (N863, N860);
xor XOR2 (N864, N856, N20);
xor XOR2 (N865, N853, N340);
and AND2 (N866, N865, N742);
nand NAND2 (N867, N835, N505);
nand NAND4 (N868, N843, N49, N617, N94);
nand NAND2 (N869, N861, N118);
nor NOR2 (N870, N864, N434);
and AND2 (N871, N841, N300);
nor NOR4 (N872, N870, N711, N549, N200);
xor XOR2 (N873, N793, N368);
nand NAND2 (N874, N862, N75);
xor XOR2 (N875, N863, N553);
buf BUF1 (N876, N866);
buf BUF1 (N877, N876);
nand NAND4 (N878, N869, N650, N454, N208);
buf BUF1 (N879, N872);
not NOT1 (N880, N868);
buf BUF1 (N881, N874);
buf BUF1 (N882, N880);
or OR4 (N883, N875, N260, N858, N698);
nor NOR4 (N884, N859, N160, N471, N826);
nand NAND2 (N885, N877, N82);
xor XOR2 (N886, N882, N683);
and AND2 (N887, N867, N210);
and AND2 (N888, N886, N871);
nand NAND3 (N889, N99, N692, N113);
or OR2 (N890, N878, N571);
nor NOR2 (N891, N884, N827);
xor XOR2 (N892, N873, N520);
xor XOR2 (N893, N885, N595);
buf BUF1 (N894, N883);
nor NOR4 (N895, N890, N130, N452, N523);
and AND2 (N896, N888, N654);
xor XOR2 (N897, N894, N84);
not NOT1 (N898, N896);
xor XOR2 (N899, N889, N108);
not NOT1 (N900, N892);
nor NOR3 (N901, N900, N50, N77);
nand NAND2 (N902, N898, N363);
buf BUF1 (N903, N902);
buf BUF1 (N904, N897);
nor NOR2 (N905, N904, N542);
buf BUF1 (N906, N899);
or OR2 (N907, N879, N549);
nand NAND2 (N908, N901, N300);
or OR4 (N909, N895, N844, N631, N54);
nor NOR3 (N910, N906, N251, N847);
xor XOR2 (N911, N910, N431);
nand NAND2 (N912, N903, N477);
xor XOR2 (N913, N909, N827);
or OR4 (N914, N893, N24, N793, N686);
and AND4 (N915, N905, N536, N72, N262);
nor NOR4 (N916, N881, N322, N888, N303);
nor NOR4 (N917, N912, N88, N889, N805);
buf BUF1 (N918, N914);
or OR3 (N919, N891, N326, N194);
or OR3 (N920, N918, N850, N310);
or OR4 (N921, N911, N485, N270, N612);
and AND4 (N922, N913, N267, N722, N48);
xor XOR2 (N923, N907, N237);
nand NAND2 (N924, N916, N309);
nor NOR4 (N925, N917, N399, N615, N665);
xor XOR2 (N926, N919, N627);
or OR2 (N927, N915, N123);
or OR2 (N928, N925, N234);
buf BUF1 (N929, N927);
and AND4 (N930, N887, N644, N76, N416);
or OR3 (N931, N920, N625, N360);
xor XOR2 (N932, N908, N129);
not NOT1 (N933, N928);
buf BUF1 (N934, N930);
nand NAND4 (N935, N921, N553, N574, N599);
not NOT1 (N936, N924);
nand NAND2 (N937, N922, N398);
or OR3 (N938, N937, N272, N251);
nor NOR3 (N939, N933, N120, N597);
nand NAND3 (N940, N931, N106, N97);
not NOT1 (N941, N934);
not NOT1 (N942, N940);
or OR3 (N943, N935, N328, N678);
nand NAND4 (N944, N938, N355, N705, N240);
buf BUF1 (N945, N926);
buf BUF1 (N946, N945);
or OR3 (N947, N929, N723, N638);
or OR2 (N948, N923, N580);
xor XOR2 (N949, N948, N470);
buf BUF1 (N950, N936);
and AND3 (N951, N947, N713, N383);
or OR2 (N952, N932, N442);
and AND3 (N953, N946, N344, N735);
or OR2 (N954, N941, N594);
not NOT1 (N955, N944);
and AND2 (N956, N954, N626);
and AND2 (N957, N956, N693);
xor XOR2 (N958, N951, N154);
nand NAND2 (N959, N942, N880);
nor NOR4 (N960, N943, N847, N801, N41);
xor XOR2 (N961, N953, N401);
nand NAND2 (N962, N955, N917);
nor NOR3 (N963, N952, N870, N587);
nor NOR2 (N964, N939, N334);
nand NAND4 (N965, N964, N244, N711, N225);
or OR4 (N966, N958, N942, N752, N200);
buf BUF1 (N967, N962);
buf BUF1 (N968, N960);
buf BUF1 (N969, N968);
and AND3 (N970, N949, N854, N569);
buf BUF1 (N971, N961);
or OR2 (N972, N965, N195);
or OR3 (N973, N959, N604, N806);
buf BUF1 (N974, N970);
not NOT1 (N975, N973);
nand NAND3 (N976, N967, N251, N319);
and AND3 (N977, N975, N19, N522);
and AND2 (N978, N976, N504);
xor XOR2 (N979, N978, N562);
buf BUF1 (N980, N974);
xor XOR2 (N981, N963, N638);
buf BUF1 (N982, N950);
and AND2 (N983, N971, N204);
not NOT1 (N984, N972);
and AND4 (N985, N957, N492, N52, N327);
xor XOR2 (N986, N980, N305);
or OR3 (N987, N984, N620, N702);
nand NAND4 (N988, N987, N75, N590, N312);
and AND3 (N989, N985, N723, N893);
not NOT1 (N990, N977);
and AND4 (N991, N983, N14, N292, N883);
not NOT1 (N992, N981);
nand NAND3 (N993, N982, N250, N587);
or OR3 (N994, N979, N69, N2);
buf BUF1 (N995, N986);
nand NAND4 (N996, N991, N328, N566, N222);
nand NAND3 (N997, N988, N770, N411);
xor XOR2 (N998, N992, N799);
xor XOR2 (N999, N966, N818);
xor XOR2 (N1000, N998, N485);
buf BUF1 (N1001, N1000);
or OR2 (N1002, N997, N969);
and AND4 (N1003, N594, N766, N475, N689);
buf BUF1 (N1004, N999);
xor XOR2 (N1005, N993, N155);
or OR4 (N1006, N1004, N627, N88, N948);
and AND2 (N1007, N989, N714);
nor NOR2 (N1008, N1005, N896);
nor NOR3 (N1009, N995, N328, N864);
or OR2 (N1010, N1007, N1008);
buf BUF1 (N1011, N805);
and AND2 (N1012, N996, N574);
nor NOR4 (N1013, N1010, N870, N440, N463);
or OR4 (N1014, N1006, N791, N267, N997);
nand NAND2 (N1015, N1002, N692);
not NOT1 (N1016, N1001);
xor XOR2 (N1017, N1013, N328);
not NOT1 (N1018, N1012);
buf BUF1 (N1019, N1011);
not NOT1 (N1020, N1018);
nand NAND3 (N1021, N1015, N857, N892);
not NOT1 (N1022, N1016);
not NOT1 (N1023, N990);
nor NOR3 (N1024, N1021, N322, N248);
or OR2 (N1025, N1017, N68);
xor XOR2 (N1026, N1019, N232);
nor NOR2 (N1027, N1025, N498);
buf BUF1 (N1028, N1020);
not NOT1 (N1029, N1003);
and AND4 (N1030, N1022, N458, N110, N465);
and AND2 (N1031, N1028, N628);
and AND4 (N1032, N1026, N1021, N71, N407);
and AND4 (N1033, N1032, N313, N550, N974);
or OR2 (N1034, N1027, N394);
or OR4 (N1035, N1034, N170, N470, N94);
nor NOR3 (N1036, N1030, N719, N873);
buf BUF1 (N1037, N994);
or OR4 (N1038, N1023, N846, N903, N614);
nor NOR3 (N1039, N1024, N80, N392);
not NOT1 (N1040, N1031);
buf BUF1 (N1041, N1036);
or OR2 (N1042, N1014, N1011);
nand NAND4 (N1043, N1037, N434, N142, N242);
buf BUF1 (N1044, N1043);
nand NAND2 (N1045, N1029, N251);
nor NOR2 (N1046, N1045, N464);
and AND4 (N1047, N1041, N73, N656, N547);
nor NOR4 (N1048, N1047, N960, N489, N490);
or OR4 (N1049, N1039, N581, N405, N10);
nor NOR3 (N1050, N1035, N560, N758);
not NOT1 (N1051, N1049);
nand NAND3 (N1052, N1044, N470, N397);
nand NAND3 (N1053, N1050, N460, N23);
xor XOR2 (N1054, N1042, N799);
not NOT1 (N1055, N1009);
and AND3 (N1056, N1051, N792, N884);
xor XOR2 (N1057, N1048, N598);
and AND2 (N1058, N1055, N533);
buf BUF1 (N1059, N1058);
not NOT1 (N1060, N1033);
and AND2 (N1061, N1054, N543);
and AND2 (N1062, N1057, N602);
xor XOR2 (N1063, N1052, N111);
buf BUF1 (N1064, N1056);
not NOT1 (N1065, N1053);
and AND3 (N1066, N1046, N325, N222);
nand NAND4 (N1067, N1065, N720, N117, N889);
nor NOR4 (N1068, N1066, N357, N751, N622);
xor XOR2 (N1069, N1063, N505);
xor XOR2 (N1070, N1064, N360);
or OR3 (N1071, N1060, N730, N378);
buf BUF1 (N1072, N1040);
xor XOR2 (N1073, N1070, N1003);
and AND3 (N1074, N1059, N684, N333);
nor NOR4 (N1075, N1062, N479, N359, N234);
not NOT1 (N1076, N1072);
not NOT1 (N1077, N1068);
or OR2 (N1078, N1073, N947);
buf BUF1 (N1079, N1077);
xor XOR2 (N1080, N1078, N28);
xor XOR2 (N1081, N1061, N790);
and AND4 (N1082, N1069, N1070, N987, N1029);
or OR4 (N1083, N1067, N401, N384, N228);
or OR2 (N1084, N1083, N320);
xor XOR2 (N1085, N1075, N991);
xor XOR2 (N1086, N1081, N654);
and AND2 (N1087, N1085, N149);
or OR3 (N1088, N1071, N117, N36);
and AND4 (N1089, N1086, N580, N148, N844);
nor NOR3 (N1090, N1082, N162, N776);
buf BUF1 (N1091, N1087);
not NOT1 (N1092, N1089);
xor XOR2 (N1093, N1092, N490);
and AND2 (N1094, N1076, N222);
not NOT1 (N1095, N1038);
nor NOR3 (N1096, N1095, N620, N88);
nand NAND4 (N1097, N1079, N972, N397, N1017);
nand NAND3 (N1098, N1094, N337, N161);
or OR4 (N1099, N1093, N166, N526, N505);
nand NAND3 (N1100, N1096, N268, N405);
buf BUF1 (N1101, N1099);
buf BUF1 (N1102, N1074);
nand NAND4 (N1103, N1080, N15, N785, N146);
not NOT1 (N1104, N1101);
xor XOR2 (N1105, N1102, N387);
not NOT1 (N1106, N1105);
or OR2 (N1107, N1100, N964);
or OR2 (N1108, N1090, N441);
or OR4 (N1109, N1091, N677, N615, N55);
xor XOR2 (N1110, N1084, N1044);
or OR2 (N1111, N1104, N990);
and AND2 (N1112, N1108, N793);
or OR4 (N1113, N1106, N899, N770, N969);
and AND3 (N1114, N1111, N895, N1081);
nor NOR4 (N1115, N1097, N969, N1069, N1108);
not NOT1 (N1116, N1110);
not NOT1 (N1117, N1115);
buf BUF1 (N1118, N1113);
buf BUF1 (N1119, N1118);
and AND3 (N1120, N1107, N222, N774);
buf BUF1 (N1121, N1088);
and AND4 (N1122, N1120, N185, N874, N255);
nor NOR2 (N1123, N1112, N753);
nand NAND3 (N1124, N1119, N547, N807);
or OR3 (N1125, N1116, N652, N346);
xor XOR2 (N1126, N1103, N377);
xor XOR2 (N1127, N1123, N833);
nand NAND2 (N1128, N1125, N684);
and AND4 (N1129, N1117, N1053, N761, N583);
or OR2 (N1130, N1126, N915);
nor NOR4 (N1131, N1128, N593, N921, N1023);
nand NAND2 (N1132, N1129, N785);
or OR4 (N1133, N1131, N532, N825, N873);
and AND3 (N1134, N1098, N564, N281);
and AND4 (N1135, N1130, N868, N834, N1031);
buf BUF1 (N1136, N1133);
xor XOR2 (N1137, N1121, N962);
nand NAND3 (N1138, N1136, N540, N285);
or OR4 (N1139, N1132, N336, N970, N247);
nand NAND2 (N1140, N1134, N930);
nand NAND3 (N1141, N1114, N274, N321);
buf BUF1 (N1142, N1109);
or OR2 (N1143, N1124, N870);
nand NAND3 (N1144, N1141, N657, N906);
not NOT1 (N1145, N1140);
not NOT1 (N1146, N1138);
nor NOR2 (N1147, N1145, N1075);
not NOT1 (N1148, N1144);
buf BUF1 (N1149, N1135);
nand NAND3 (N1150, N1127, N421, N981);
and AND2 (N1151, N1149, N68);
and AND2 (N1152, N1151, N473);
xor XOR2 (N1153, N1150, N1045);
and AND4 (N1154, N1142, N1082, N543, N1011);
and AND2 (N1155, N1148, N201);
not NOT1 (N1156, N1137);
nand NAND3 (N1157, N1156, N560, N857);
and AND4 (N1158, N1152, N902, N530, N841);
nor NOR3 (N1159, N1146, N928, N81);
nand NAND2 (N1160, N1147, N607);
xor XOR2 (N1161, N1155, N1074);
not NOT1 (N1162, N1153);
buf BUF1 (N1163, N1162);
not NOT1 (N1164, N1157);
nand NAND2 (N1165, N1158, N405);
buf BUF1 (N1166, N1165);
not NOT1 (N1167, N1166);
not NOT1 (N1168, N1164);
nor NOR3 (N1169, N1154, N548, N472);
not NOT1 (N1170, N1167);
buf BUF1 (N1171, N1160);
nand NAND2 (N1172, N1139, N755);
nor NOR4 (N1173, N1172, N1063, N98, N354);
nor NOR2 (N1174, N1122, N120);
not NOT1 (N1175, N1163);
buf BUF1 (N1176, N1171);
xor XOR2 (N1177, N1168, N1043);
buf BUF1 (N1178, N1174);
nand NAND3 (N1179, N1176, N837, N1014);
xor XOR2 (N1180, N1173, N3);
not NOT1 (N1181, N1178);
and AND3 (N1182, N1170, N362, N856);
not NOT1 (N1183, N1159);
buf BUF1 (N1184, N1161);
buf BUF1 (N1185, N1177);
not NOT1 (N1186, N1143);
nand NAND2 (N1187, N1181, N573);
or OR3 (N1188, N1180, N440, N768);
nand NAND2 (N1189, N1186, N572);
xor XOR2 (N1190, N1179, N237);
and AND4 (N1191, N1189, N22, N1106, N797);
nand NAND3 (N1192, N1190, N905, N115);
nor NOR2 (N1193, N1182, N956);
and AND2 (N1194, N1193, N609);
buf BUF1 (N1195, N1187);
buf BUF1 (N1196, N1194);
or OR2 (N1197, N1191, N1125);
buf BUF1 (N1198, N1188);
xor XOR2 (N1199, N1185, N694);
buf BUF1 (N1200, N1198);
buf BUF1 (N1201, N1199);
and AND3 (N1202, N1169, N756, N820);
xor XOR2 (N1203, N1192, N370);
not NOT1 (N1204, N1195);
xor XOR2 (N1205, N1197, N948);
buf BUF1 (N1206, N1201);
xor XOR2 (N1207, N1205, N253);
nor NOR4 (N1208, N1202, N817, N796, N1098);
xor XOR2 (N1209, N1196, N45);
buf BUF1 (N1210, N1207);
nor NOR2 (N1211, N1204, N1087);
xor XOR2 (N1212, N1206, N578);
or OR4 (N1213, N1203, N974, N700, N111);
or OR3 (N1214, N1212, N814, N1195);
nor NOR4 (N1215, N1208, N732, N980, N912);
and AND4 (N1216, N1175, N939, N155, N246);
or OR2 (N1217, N1215, N686);
and AND4 (N1218, N1184, N285, N1058, N869);
nand NAND2 (N1219, N1210, N1013);
nor NOR2 (N1220, N1213, N96);
nor NOR2 (N1221, N1214, N340);
buf BUF1 (N1222, N1220);
not NOT1 (N1223, N1218);
buf BUF1 (N1224, N1216);
nor NOR4 (N1225, N1223, N1152, N128, N538);
and AND4 (N1226, N1200, N608, N1022, N96);
not NOT1 (N1227, N1221);
xor XOR2 (N1228, N1219, N884);
not NOT1 (N1229, N1226);
nor NOR2 (N1230, N1209, N468);
nand NAND2 (N1231, N1224, N232);
nor NOR4 (N1232, N1225, N732, N518, N1046);
nand NAND4 (N1233, N1227, N1064, N627, N251);
or OR2 (N1234, N1217, N1132);
or OR4 (N1235, N1232, N91, N47, N164);
xor XOR2 (N1236, N1231, N987);
nand NAND4 (N1237, N1183, N632, N1099, N248);
nand NAND4 (N1238, N1222, N1122, N481, N1168);
not NOT1 (N1239, N1230);
and AND3 (N1240, N1228, N1238, N437);
nor NOR2 (N1241, N2, N348);
xor XOR2 (N1242, N1237, N306);
xor XOR2 (N1243, N1233, N49);
nand NAND2 (N1244, N1242, N47);
buf BUF1 (N1245, N1239);
or OR2 (N1246, N1240, N673);
and AND2 (N1247, N1236, N227);
nor NOR3 (N1248, N1245, N297, N818);
or OR2 (N1249, N1211, N594);
or OR2 (N1250, N1246, N715);
buf BUF1 (N1251, N1243);
and AND3 (N1252, N1234, N260, N249);
or OR3 (N1253, N1241, N327, N630);
nand NAND3 (N1254, N1250, N1047, N305);
nand NAND3 (N1255, N1244, N1207, N859);
buf BUF1 (N1256, N1251);
nand NAND2 (N1257, N1253, N743);
nand NAND4 (N1258, N1249, N17, N1213, N629);
xor XOR2 (N1259, N1256, N1000);
xor XOR2 (N1260, N1247, N834);
buf BUF1 (N1261, N1257);
xor XOR2 (N1262, N1229, N7);
buf BUF1 (N1263, N1261);
not NOT1 (N1264, N1262);
nand NAND2 (N1265, N1260, N139);
and AND3 (N1266, N1248, N929, N605);
and AND4 (N1267, N1264, N114, N48, N725);
or OR4 (N1268, N1255, N366, N862, N983);
xor XOR2 (N1269, N1258, N523);
nand NAND4 (N1270, N1263, N49, N401, N933);
nor NOR4 (N1271, N1252, N152, N1196, N975);
and AND3 (N1272, N1265, N782, N1186);
buf BUF1 (N1273, N1259);
not NOT1 (N1274, N1268);
and AND3 (N1275, N1267, N298, N382);
not NOT1 (N1276, N1270);
nor NOR4 (N1277, N1235, N1090, N919, N939);
or OR4 (N1278, N1266, N1273, N1143, N472);
not NOT1 (N1279, N137);
xor XOR2 (N1280, N1278, N1249);
or OR2 (N1281, N1271, N940);
buf BUF1 (N1282, N1254);
not NOT1 (N1283, N1276);
buf BUF1 (N1284, N1281);
and AND2 (N1285, N1274, N788);
or OR3 (N1286, N1285, N126, N627);
and AND2 (N1287, N1272, N776);
not NOT1 (N1288, N1282);
nand NAND4 (N1289, N1280, N119, N503, N293);
xor XOR2 (N1290, N1289, N1211);
nor NOR3 (N1291, N1287, N1226, N425);
or OR2 (N1292, N1286, N551);
not NOT1 (N1293, N1288);
nand NAND3 (N1294, N1279, N212, N839);
buf BUF1 (N1295, N1293);
and AND2 (N1296, N1295, N152);
or OR4 (N1297, N1269, N582, N807, N1258);
not NOT1 (N1298, N1292);
nand NAND2 (N1299, N1277, N1213);
nor NOR3 (N1300, N1298, N586, N1275);
xor XOR2 (N1301, N1187, N146);
not NOT1 (N1302, N1290);
nand NAND2 (N1303, N1291, N1126);
xor XOR2 (N1304, N1303, N983);
nand NAND3 (N1305, N1283, N269, N547);
not NOT1 (N1306, N1300);
nand NAND3 (N1307, N1306, N918, N1256);
not NOT1 (N1308, N1302);
and AND2 (N1309, N1301, N150);
not NOT1 (N1310, N1307);
not NOT1 (N1311, N1299);
or OR3 (N1312, N1311, N255, N798);
and AND4 (N1313, N1309, N1236, N1001, N1146);
buf BUF1 (N1314, N1304);
nand NAND4 (N1315, N1297, N601, N33, N870);
buf BUF1 (N1316, N1310);
nor NOR3 (N1317, N1296, N817, N269);
xor XOR2 (N1318, N1314, N500);
xor XOR2 (N1319, N1313, N241);
not NOT1 (N1320, N1317);
xor XOR2 (N1321, N1312, N558);
not NOT1 (N1322, N1318);
and AND4 (N1323, N1305, N1247, N489, N326);
xor XOR2 (N1324, N1315, N1305);
and AND2 (N1325, N1308, N685);
buf BUF1 (N1326, N1316);
and AND4 (N1327, N1321, N970, N151, N712);
not NOT1 (N1328, N1325);
buf BUF1 (N1329, N1284);
and AND3 (N1330, N1294, N1046, N841);
not NOT1 (N1331, N1327);
not NOT1 (N1332, N1322);
nor NOR4 (N1333, N1319, N193, N1057, N845);
nand NAND3 (N1334, N1330, N1075, N385);
not NOT1 (N1335, N1332);
or OR4 (N1336, N1320, N338, N1110, N1032);
xor XOR2 (N1337, N1328, N827);
nand NAND2 (N1338, N1337, N922);
xor XOR2 (N1339, N1329, N1004);
nor NOR4 (N1340, N1335, N346, N744, N1290);
xor XOR2 (N1341, N1340, N1020);
and AND4 (N1342, N1339, N654, N1281, N809);
and AND4 (N1343, N1326, N1279, N988, N664);
not NOT1 (N1344, N1341);
buf BUF1 (N1345, N1343);
xor XOR2 (N1346, N1333, N68);
xor XOR2 (N1347, N1338, N728);
or OR2 (N1348, N1346, N909);
and AND3 (N1349, N1336, N849, N1081);
buf BUF1 (N1350, N1344);
nor NOR2 (N1351, N1349, N513);
nor NOR4 (N1352, N1347, N1164, N266, N956);
or OR3 (N1353, N1342, N284, N1183);
not NOT1 (N1354, N1334);
buf BUF1 (N1355, N1324);
xor XOR2 (N1356, N1353, N995);
buf BUF1 (N1357, N1350);
buf BUF1 (N1358, N1355);
xor XOR2 (N1359, N1348, N385);
nand NAND4 (N1360, N1357, N714, N1079, N787);
or OR4 (N1361, N1331, N590, N617, N1135);
nand NAND2 (N1362, N1354, N12);
nor NOR2 (N1363, N1356, N763);
xor XOR2 (N1364, N1359, N298);
not NOT1 (N1365, N1361);
or OR2 (N1366, N1345, N740);
xor XOR2 (N1367, N1360, N822);
or OR2 (N1368, N1363, N1070);
and AND3 (N1369, N1367, N480, N957);
or OR3 (N1370, N1368, N1259, N22);
not NOT1 (N1371, N1370);
nand NAND2 (N1372, N1358, N1119);
nand NAND3 (N1373, N1365, N704, N135);
not NOT1 (N1374, N1352);
and AND3 (N1375, N1351, N961, N1097);
nand NAND4 (N1376, N1375, N58, N242, N1231);
or OR4 (N1377, N1369, N404, N682, N1072);
and AND3 (N1378, N1364, N1208, N1336);
nor NOR4 (N1379, N1378, N568, N395, N814);
buf BUF1 (N1380, N1371);
nor NOR3 (N1381, N1323, N179, N807);
buf BUF1 (N1382, N1376);
or OR2 (N1383, N1373, N180);
xor XOR2 (N1384, N1377, N583);
nor NOR4 (N1385, N1379, N68, N204, N903);
or OR2 (N1386, N1381, N371);
buf BUF1 (N1387, N1386);
not NOT1 (N1388, N1372);
buf BUF1 (N1389, N1385);
and AND4 (N1390, N1380, N102, N576, N1319);
nor NOR4 (N1391, N1382, N279, N280, N16);
xor XOR2 (N1392, N1391, N828);
nand NAND3 (N1393, N1383, N758, N957);
not NOT1 (N1394, N1362);
not NOT1 (N1395, N1390);
not NOT1 (N1396, N1388);
not NOT1 (N1397, N1393);
xor XOR2 (N1398, N1396, N236);
nor NOR3 (N1399, N1384, N570, N75);
and AND2 (N1400, N1374, N1369);
buf BUF1 (N1401, N1392);
not NOT1 (N1402, N1395);
xor XOR2 (N1403, N1387, N890);
nor NOR2 (N1404, N1399, N882);
buf BUF1 (N1405, N1404);
buf BUF1 (N1406, N1405);
or OR4 (N1407, N1402, N1102, N1210, N854);
not NOT1 (N1408, N1394);
buf BUF1 (N1409, N1397);
or OR3 (N1410, N1398, N452, N151);
and AND3 (N1411, N1400, N289, N619);
and AND4 (N1412, N1408, N157, N1249, N1317);
xor XOR2 (N1413, N1366, N121);
buf BUF1 (N1414, N1413);
and AND2 (N1415, N1389, N263);
nor NOR2 (N1416, N1415, N1070);
xor XOR2 (N1417, N1409, N459);
nand NAND4 (N1418, N1414, N1181, N629, N958);
or OR3 (N1419, N1401, N916, N1401);
nor NOR3 (N1420, N1419, N839, N1332);
buf BUF1 (N1421, N1411);
not NOT1 (N1422, N1416);
nor NOR3 (N1423, N1417, N148, N1238);
nand NAND3 (N1424, N1422, N910, N440);
not NOT1 (N1425, N1423);
nor NOR3 (N1426, N1406, N473, N816);
xor XOR2 (N1427, N1425, N1257);
nand NAND2 (N1428, N1410, N153);
and AND3 (N1429, N1428, N1158, N554);
and AND2 (N1430, N1429, N241);
not NOT1 (N1431, N1403);
nand NAND4 (N1432, N1420, N764, N686, N941);
not NOT1 (N1433, N1418);
nor NOR2 (N1434, N1432, N1170);
or OR4 (N1435, N1421, N1224, N357, N153);
not NOT1 (N1436, N1424);
and AND2 (N1437, N1435, N789);
or OR4 (N1438, N1430, N333, N200, N894);
buf BUF1 (N1439, N1438);
xor XOR2 (N1440, N1439, N948);
nand NAND2 (N1441, N1426, N770);
not NOT1 (N1442, N1440);
nor NOR4 (N1443, N1433, N747, N982, N1029);
xor XOR2 (N1444, N1431, N418);
or OR3 (N1445, N1412, N98, N527);
and AND3 (N1446, N1441, N255, N337);
or OR3 (N1447, N1407, N412, N641);
and AND3 (N1448, N1434, N524, N459);
nand NAND2 (N1449, N1442, N228);
nor NOR3 (N1450, N1444, N463, N1188);
and AND4 (N1451, N1443, N464, N4, N686);
or OR2 (N1452, N1446, N789);
nor NOR3 (N1453, N1447, N1360, N151);
not NOT1 (N1454, N1453);
or OR2 (N1455, N1452, N308);
or OR2 (N1456, N1436, N186);
and AND2 (N1457, N1456, N183);
not NOT1 (N1458, N1451);
nand NAND3 (N1459, N1437, N370, N185);
nor NOR2 (N1460, N1427, N1077);
or OR4 (N1461, N1457, N1396, N444, N1221);
nor NOR3 (N1462, N1455, N706, N1083);
or OR3 (N1463, N1460, N321, N1041);
nor NOR3 (N1464, N1449, N406, N745);
or OR2 (N1465, N1458, N1211);
xor XOR2 (N1466, N1450, N919);
and AND4 (N1467, N1466, N1234, N20, N1432);
nand NAND2 (N1468, N1448, N1403);
nand NAND4 (N1469, N1463, N1358, N1138, N288);
not NOT1 (N1470, N1461);
nor NOR3 (N1471, N1468, N682, N1246);
and AND3 (N1472, N1454, N785, N1213);
or OR4 (N1473, N1445, N203, N1067, N1315);
nand NAND2 (N1474, N1459, N1023);
nand NAND2 (N1475, N1472, N1347);
buf BUF1 (N1476, N1464);
xor XOR2 (N1477, N1469, N577);
not NOT1 (N1478, N1477);
nand NAND2 (N1479, N1473, N1019);
not NOT1 (N1480, N1470);
xor XOR2 (N1481, N1474, N515);
or OR2 (N1482, N1479, N484);
and AND3 (N1483, N1478, N679, N158);
buf BUF1 (N1484, N1481);
and AND3 (N1485, N1465, N54, N639);
nand NAND2 (N1486, N1475, N198);
nor NOR3 (N1487, N1482, N578, N541);
buf BUF1 (N1488, N1467);
buf BUF1 (N1489, N1485);
and AND2 (N1490, N1487, N370);
xor XOR2 (N1491, N1476, N415);
or OR4 (N1492, N1484, N1231, N269, N600);
or OR2 (N1493, N1471, N503);
buf BUF1 (N1494, N1491);
buf BUF1 (N1495, N1492);
and AND3 (N1496, N1488, N875, N1202);
buf BUF1 (N1497, N1489);
and AND2 (N1498, N1493, N294);
not NOT1 (N1499, N1495);
buf BUF1 (N1500, N1498);
not NOT1 (N1501, N1462);
nor NOR4 (N1502, N1500, N559, N789, N392);
or OR4 (N1503, N1499, N539, N858, N1444);
nand NAND4 (N1504, N1501, N286, N820, N666);
and AND4 (N1505, N1504, N1256, N8, N353);
xor XOR2 (N1506, N1503, N1278);
buf BUF1 (N1507, N1483);
or OR3 (N1508, N1490, N396, N757);
xor XOR2 (N1509, N1497, N201);
xor XOR2 (N1510, N1480, N1417);
or OR3 (N1511, N1496, N953, N148);
nand NAND2 (N1512, N1508, N54);
nand NAND4 (N1513, N1510, N1499, N256, N470);
and AND3 (N1514, N1513, N1285, N1513);
not NOT1 (N1515, N1494);
buf BUF1 (N1516, N1509);
and AND4 (N1517, N1516, N927, N120, N975);
nor NOR2 (N1518, N1486, N219);
nand NAND3 (N1519, N1505, N706, N1378);
not NOT1 (N1520, N1507);
not NOT1 (N1521, N1514);
nor NOR2 (N1522, N1511, N287);
and AND2 (N1523, N1520, N137);
or OR2 (N1524, N1512, N99);
or OR4 (N1525, N1515, N1236, N609, N720);
not NOT1 (N1526, N1525);
and AND3 (N1527, N1506, N954, N1187);
buf BUF1 (N1528, N1502);
buf BUF1 (N1529, N1526);
nor NOR3 (N1530, N1518, N1323, N756);
and AND4 (N1531, N1528, N740, N681, N1511);
buf BUF1 (N1532, N1529);
buf BUF1 (N1533, N1521);
xor XOR2 (N1534, N1533, N748);
nor NOR3 (N1535, N1532, N1075, N1201);
and AND2 (N1536, N1523, N1236);
nor NOR3 (N1537, N1519, N1154, N1128);
and AND2 (N1538, N1536, N416);
or OR3 (N1539, N1531, N817, N952);
nand NAND2 (N1540, N1524, N817);
or OR4 (N1541, N1527, N1423, N1322, N1472);
nand NAND2 (N1542, N1522, N510);
not NOT1 (N1543, N1540);
or OR4 (N1544, N1534, N178, N733, N1110);
not NOT1 (N1545, N1542);
nand NAND3 (N1546, N1530, N160, N1395);
not NOT1 (N1547, N1546);
not NOT1 (N1548, N1537);
nand NAND3 (N1549, N1539, N1297, N212);
nor NOR4 (N1550, N1541, N894, N174, N951);
nand NAND4 (N1551, N1538, N1509, N1113, N160);
nor NOR3 (N1552, N1517, N262, N1456);
xor XOR2 (N1553, N1552, N186);
or OR2 (N1554, N1545, N1208);
nand NAND2 (N1555, N1549, N1082);
not NOT1 (N1556, N1551);
buf BUF1 (N1557, N1554);
not NOT1 (N1558, N1557);
buf BUF1 (N1559, N1547);
nor NOR2 (N1560, N1550, N717);
buf BUF1 (N1561, N1544);
and AND2 (N1562, N1548, N1538);
nor NOR4 (N1563, N1543, N831, N126, N1453);
and AND3 (N1564, N1556, N668, N1303);
nand NAND4 (N1565, N1553, N1295, N855, N488);
and AND2 (N1566, N1563, N261);
nand NAND2 (N1567, N1566, N67);
not NOT1 (N1568, N1535);
and AND3 (N1569, N1561, N710, N1233);
nand NAND3 (N1570, N1564, N630, N1304);
buf BUF1 (N1571, N1562);
xor XOR2 (N1572, N1569, N1401);
or OR4 (N1573, N1567, N1272, N1280, N1391);
nand NAND4 (N1574, N1571, N208, N65, N797);
not NOT1 (N1575, N1568);
xor XOR2 (N1576, N1555, N727);
nand NAND4 (N1577, N1574, N418, N191, N161);
or OR4 (N1578, N1565, N845, N951, N1348);
xor XOR2 (N1579, N1577, N377);
xor XOR2 (N1580, N1576, N676);
nor NOR3 (N1581, N1572, N1286, N837);
nand NAND3 (N1582, N1581, N550, N32);
not NOT1 (N1583, N1578);
nor NOR4 (N1584, N1570, N1279, N500, N1532);
or OR3 (N1585, N1560, N212, N481);
or OR4 (N1586, N1583, N541, N163, N830);
or OR4 (N1587, N1585, N1207, N748, N844);
and AND3 (N1588, N1575, N1392, N510);
nand NAND2 (N1589, N1573, N1060);
nand NAND2 (N1590, N1589, N221);
nor NOR2 (N1591, N1558, N1235);
nor NOR4 (N1592, N1580, N173, N484, N960);
or OR2 (N1593, N1584, N944);
or OR4 (N1594, N1591, N335, N723, N1491);
and AND4 (N1595, N1593, N451, N588, N1355);
nor NOR4 (N1596, N1590, N1176, N442, N82);
xor XOR2 (N1597, N1587, N1457);
and AND3 (N1598, N1596, N1409, N1204);
nand NAND4 (N1599, N1598, N1124, N1590, N1125);
nand NAND2 (N1600, N1592, N1450);
and AND4 (N1601, N1597, N1085, N323, N943);
nor NOR4 (N1602, N1594, N855, N1452, N709);
not NOT1 (N1603, N1595);
or OR2 (N1604, N1599, N1479);
and AND4 (N1605, N1579, N1579, N108, N1139);
nor NOR2 (N1606, N1586, N933);
or OR4 (N1607, N1600, N457, N1418, N545);
buf BUF1 (N1608, N1602);
or OR4 (N1609, N1606, N1005, N75, N509);
or OR4 (N1610, N1582, N1462, N1277, N899);
buf BUF1 (N1611, N1610);
buf BUF1 (N1612, N1605);
buf BUF1 (N1613, N1588);
or OR2 (N1614, N1613, N925);
not NOT1 (N1615, N1607);
xor XOR2 (N1616, N1614, N846);
not NOT1 (N1617, N1611);
nor NOR2 (N1618, N1612, N1069);
and AND4 (N1619, N1608, N1144, N475, N214);
not NOT1 (N1620, N1604);
nand NAND4 (N1621, N1618, N1164, N656, N406);
and AND4 (N1622, N1621, N1083, N769, N827);
and AND2 (N1623, N1559, N347);
nand NAND3 (N1624, N1615, N849, N331);
not NOT1 (N1625, N1601);
xor XOR2 (N1626, N1623, N902);
and AND3 (N1627, N1620, N215, N357);
and AND3 (N1628, N1619, N742, N733);
or OR3 (N1629, N1624, N405, N458);
and AND2 (N1630, N1616, N487);
xor XOR2 (N1631, N1609, N48);
buf BUF1 (N1632, N1631);
buf BUF1 (N1633, N1625);
xor XOR2 (N1634, N1627, N135);
or OR3 (N1635, N1630, N227, N96);
and AND2 (N1636, N1626, N340);
nand NAND2 (N1637, N1617, N1051);
and AND2 (N1638, N1634, N139);
buf BUF1 (N1639, N1637);
not NOT1 (N1640, N1638);
xor XOR2 (N1641, N1628, N1342);
nand NAND4 (N1642, N1633, N187, N522, N128);
not NOT1 (N1643, N1629);
xor XOR2 (N1644, N1642, N1003);
xor XOR2 (N1645, N1641, N547);
buf BUF1 (N1646, N1635);
or OR3 (N1647, N1644, N69, N328);
nand NAND4 (N1648, N1639, N299, N1413, N1530);
not NOT1 (N1649, N1636);
or OR4 (N1650, N1646, N560, N665, N1385);
nor NOR4 (N1651, N1645, N918, N1142, N201);
not NOT1 (N1652, N1647);
not NOT1 (N1653, N1643);
and AND2 (N1654, N1652, N941);
and AND3 (N1655, N1650, N717, N1249);
and AND3 (N1656, N1648, N538, N1334);
nand NAND4 (N1657, N1651, N694, N1350, N109);
nand NAND3 (N1658, N1649, N336, N1319);
not NOT1 (N1659, N1632);
and AND2 (N1660, N1657, N324);
not NOT1 (N1661, N1655);
xor XOR2 (N1662, N1622, N918);
nor NOR2 (N1663, N1659, N456);
xor XOR2 (N1664, N1662, N249);
and AND2 (N1665, N1663, N1232);
or OR2 (N1666, N1654, N570);
or OR2 (N1667, N1664, N1392);
buf BUF1 (N1668, N1640);
not NOT1 (N1669, N1653);
not NOT1 (N1670, N1660);
xor XOR2 (N1671, N1656, N601);
buf BUF1 (N1672, N1668);
nor NOR3 (N1673, N1672, N1078, N805);
or OR4 (N1674, N1669, N229, N1132, N113);
and AND4 (N1675, N1658, N1256, N1618, N1127);
xor XOR2 (N1676, N1661, N973);
or OR3 (N1677, N1674, N793, N547);
nor NOR3 (N1678, N1677, N468, N174);
nand NAND4 (N1679, N1667, N1546, N148, N637);
not NOT1 (N1680, N1603);
xor XOR2 (N1681, N1670, N850);
nor NOR4 (N1682, N1676, N949, N1122, N1290);
or OR3 (N1683, N1671, N440, N1196);
buf BUF1 (N1684, N1666);
or OR4 (N1685, N1683, N722, N1518, N366);
not NOT1 (N1686, N1675);
nand NAND4 (N1687, N1686, N529, N1387, N871);
nand NAND2 (N1688, N1684, N1506);
and AND3 (N1689, N1679, N1168, N1376);
or OR3 (N1690, N1678, N410, N1513);
or OR4 (N1691, N1690, N1617, N1284, N144);
xor XOR2 (N1692, N1680, N383);
not NOT1 (N1693, N1691);
or OR4 (N1694, N1665, N756, N212, N904);
and AND4 (N1695, N1693, N411, N968, N1461);
or OR4 (N1696, N1685, N389, N784, N1413);
and AND2 (N1697, N1688, N1480);
xor XOR2 (N1698, N1694, N1486);
buf BUF1 (N1699, N1687);
nor NOR2 (N1700, N1689, N1111);
buf BUF1 (N1701, N1697);
nor NOR3 (N1702, N1681, N1011, N270);
nand NAND3 (N1703, N1673, N804, N1535);
buf BUF1 (N1704, N1682);
nor NOR3 (N1705, N1696, N1653, N1383);
not NOT1 (N1706, N1698);
xor XOR2 (N1707, N1704, N1367);
or OR4 (N1708, N1695, N549, N315, N1414);
nor NOR4 (N1709, N1702, N1369, N321, N377);
nor NOR4 (N1710, N1709, N435, N734, N242);
or OR3 (N1711, N1708, N1360, N620);
or OR3 (N1712, N1706, N69, N722);
not NOT1 (N1713, N1710);
and AND3 (N1714, N1711, N442, N1240);
and AND3 (N1715, N1703, N1381, N1615);
buf BUF1 (N1716, N1712);
buf BUF1 (N1717, N1714);
not NOT1 (N1718, N1701);
not NOT1 (N1719, N1715);
and AND2 (N1720, N1692, N470);
and AND4 (N1721, N1707, N651, N839, N354);
and AND4 (N1722, N1716, N51, N1521, N377);
buf BUF1 (N1723, N1719);
buf BUF1 (N1724, N1705);
not NOT1 (N1725, N1722);
not NOT1 (N1726, N1700);
nand NAND2 (N1727, N1718, N882);
buf BUF1 (N1728, N1720);
not NOT1 (N1729, N1723);
or OR3 (N1730, N1721, N1009, N1536);
xor XOR2 (N1731, N1727, N302);
or OR4 (N1732, N1725, N701, N1264, N216);
and AND4 (N1733, N1731, N205, N739, N1261);
xor XOR2 (N1734, N1717, N643);
nand NAND3 (N1735, N1733, N130, N1097);
buf BUF1 (N1736, N1732);
xor XOR2 (N1737, N1728, N497);
and AND3 (N1738, N1730, N418, N1212);
and AND3 (N1739, N1736, N764, N908);
nand NAND2 (N1740, N1724, N970);
nor NOR3 (N1741, N1699, N163, N1505);
and AND2 (N1742, N1737, N879);
buf BUF1 (N1743, N1738);
xor XOR2 (N1744, N1734, N1528);
xor XOR2 (N1745, N1742, N1242);
and AND3 (N1746, N1745, N1640, N1629);
nand NAND2 (N1747, N1726, N1680);
not NOT1 (N1748, N1747);
and AND3 (N1749, N1746, N1076, N1489);
nand NAND4 (N1750, N1729, N1661, N897, N41);
nand NAND2 (N1751, N1740, N10);
not NOT1 (N1752, N1713);
and AND2 (N1753, N1739, N1462);
nor NOR4 (N1754, N1749, N1685, N1376, N1447);
nand NAND2 (N1755, N1743, N913);
nor NOR2 (N1756, N1741, N1737);
nor NOR4 (N1757, N1752, N1014, N220, N566);
nand NAND4 (N1758, N1757, N335, N1196, N1069);
not NOT1 (N1759, N1748);
nand NAND4 (N1760, N1750, N682, N1099, N788);
or OR2 (N1761, N1758, N788);
xor XOR2 (N1762, N1755, N1614);
or OR2 (N1763, N1735, N1173);
nand NAND4 (N1764, N1763, N347, N985, N170);
or OR2 (N1765, N1764, N1638);
nor NOR3 (N1766, N1756, N417, N1205);
not NOT1 (N1767, N1765);
or OR4 (N1768, N1766, N1716, N963, N159);
not NOT1 (N1769, N1751);
xor XOR2 (N1770, N1768, N327);
nand NAND3 (N1771, N1767, N1298, N253);
or OR3 (N1772, N1753, N1312, N1468);
buf BUF1 (N1773, N1759);
nand NAND4 (N1774, N1771, N1445, N1026, N1488);
nand NAND2 (N1775, N1744, N887);
nor NOR2 (N1776, N1775, N1599);
nor NOR3 (N1777, N1772, N1746, N988);
nor NOR4 (N1778, N1776, N1471, N626, N1581);
or OR3 (N1779, N1754, N1074, N605);
and AND4 (N1780, N1773, N587, N350, N1501);
or OR3 (N1781, N1774, N612, N1470);
and AND3 (N1782, N1780, N839, N489);
xor XOR2 (N1783, N1762, N1515);
or OR2 (N1784, N1769, N74);
and AND3 (N1785, N1781, N1476, N999);
nand NAND4 (N1786, N1761, N262, N289, N1208);
buf BUF1 (N1787, N1782);
buf BUF1 (N1788, N1779);
not NOT1 (N1789, N1784);
nor NOR3 (N1790, N1770, N404, N1669);
nand NAND2 (N1791, N1785, N1029);
nand NAND3 (N1792, N1778, N142, N822);
nor NOR4 (N1793, N1790, N277, N176, N454);
and AND2 (N1794, N1760, N1790);
or OR3 (N1795, N1783, N981, N1257);
and AND2 (N1796, N1793, N1320);
buf BUF1 (N1797, N1777);
nor NOR3 (N1798, N1787, N1748, N1365);
buf BUF1 (N1799, N1792);
nor NOR4 (N1800, N1786, N909, N289, N1701);
and AND3 (N1801, N1794, N1065, N1206);
and AND4 (N1802, N1800, N5, N1503, N993);
or OR2 (N1803, N1798, N92);
or OR2 (N1804, N1788, N1305);
xor XOR2 (N1805, N1803, N1648);
nor NOR4 (N1806, N1796, N1586, N1340, N1519);
nor NOR4 (N1807, N1805, N1742, N1040, N838);
nand NAND2 (N1808, N1806, N535);
buf BUF1 (N1809, N1797);
and AND2 (N1810, N1804, N1307);
buf BUF1 (N1811, N1789);
and AND3 (N1812, N1809, N231, N1558);
xor XOR2 (N1813, N1799, N192);
not NOT1 (N1814, N1813);
or OR3 (N1815, N1807, N400, N1175);
buf BUF1 (N1816, N1802);
nand NAND3 (N1817, N1814, N1587, N185);
buf BUF1 (N1818, N1815);
not NOT1 (N1819, N1808);
buf BUF1 (N1820, N1810);
xor XOR2 (N1821, N1817, N1742);
nor NOR3 (N1822, N1811, N1477, N22);
buf BUF1 (N1823, N1819);
buf BUF1 (N1824, N1820);
or OR4 (N1825, N1801, N149, N1171, N1190);
nand NAND2 (N1826, N1816, N1210);
or OR2 (N1827, N1826, N783);
not NOT1 (N1828, N1824);
and AND3 (N1829, N1795, N786, N100);
not NOT1 (N1830, N1821);
nand NAND3 (N1831, N1812, N103, N896);
not NOT1 (N1832, N1822);
or OR3 (N1833, N1791, N1105, N902);
nand NAND3 (N1834, N1833, N403, N818);
not NOT1 (N1835, N1818);
not NOT1 (N1836, N1827);
and AND4 (N1837, N1825, N961, N1053, N821);
xor XOR2 (N1838, N1835, N1017);
or OR4 (N1839, N1832, N866, N369, N1025);
nor NOR4 (N1840, N1837, N952, N1535, N603);
or OR2 (N1841, N1828, N1560);
buf BUF1 (N1842, N1840);
nand NAND3 (N1843, N1836, N1250, N1330);
nor NOR2 (N1844, N1831, N419);
and AND3 (N1845, N1843, N1464, N435);
nand NAND3 (N1846, N1838, N1836, N98);
nand NAND4 (N1847, N1845, N1711, N1806, N478);
nor NOR2 (N1848, N1839, N548);
nor NOR3 (N1849, N1844, N1680, N1336);
not NOT1 (N1850, N1834);
xor XOR2 (N1851, N1848, N449);
not NOT1 (N1852, N1842);
nand NAND4 (N1853, N1850, N1350, N790, N461);
buf BUF1 (N1854, N1830);
or OR3 (N1855, N1841, N1212, N1351);
nand NAND4 (N1856, N1853, N960, N1343, N1220);
buf BUF1 (N1857, N1854);
nand NAND2 (N1858, N1829, N1180);
and AND4 (N1859, N1852, N1543, N1396, N351);
or OR4 (N1860, N1859, N320, N715, N1415);
and AND3 (N1861, N1856, N775, N830);
nor NOR4 (N1862, N1860, N1472, N1104, N1801);
xor XOR2 (N1863, N1857, N338);
nand NAND2 (N1864, N1855, N1723);
and AND4 (N1865, N1849, N729, N1266, N1728);
buf BUF1 (N1866, N1861);
not NOT1 (N1867, N1858);
xor XOR2 (N1868, N1823, N435);
xor XOR2 (N1869, N1865, N1368);
xor XOR2 (N1870, N1868, N1066);
buf BUF1 (N1871, N1870);
nand NAND3 (N1872, N1862, N212, N1635);
buf BUF1 (N1873, N1847);
or OR3 (N1874, N1846, N1352, N1785);
xor XOR2 (N1875, N1867, N684);
nand NAND2 (N1876, N1864, N429);
nand NAND2 (N1877, N1869, N806);
buf BUF1 (N1878, N1863);
nand NAND4 (N1879, N1866, N1755, N1324, N959);
buf BUF1 (N1880, N1872);
nor NOR2 (N1881, N1880, N810);
or OR3 (N1882, N1874, N779, N747);
and AND2 (N1883, N1882, N1070);
or OR4 (N1884, N1879, N1232, N699, N1381);
nor NOR3 (N1885, N1851, N1348, N962);
buf BUF1 (N1886, N1884);
xor XOR2 (N1887, N1876, N702);
buf BUF1 (N1888, N1878);
nor NOR4 (N1889, N1875, N1696, N141, N1727);
nand NAND2 (N1890, N1889, N766);
buf BUF1 (N1891, N1887);
nor NOR4 (N1892, N1890, N1509, N1809, N481);
nand NAND2 (N1893, N1883, N257);
buf BUF1 (N1894, N1886);
nor NOR2 (N1895, N1888, N1313);
or OR3 (N1896, N1881, N63, N460);
not NOT1 (N1897, N1885);
nand NAND3 (N1898, N1877, N895, N1423);
nand NAND4 (N1899, N1871, N349, N523, N956);
and AND2 (N1900, N1897, N1025);
nand NAND2 (N1901, N1898, N1045);
nand NAND4 (N1902, N1891, N600, N227, N391);
and AND2 (N1903, N1900, N525);
nand NAND4 (N1904, N1895, N1083, N1183, N1490);
nor NOR4 (N1905, N1894, N1898, N260, N826);
or OR3 (N1906, N1892, N279, N1109);
or OR4 (N1907, N1902, N1717, N1422, N891);
xor XOR2 (N1908, N1906, N719);
nand NAND4 (N1909, N1893, N291, N775, N798);
or OR2 (N1910, N1903, N505);
xor XOR2 (N1911, N1904, N1476);
or OR3 (N1912, N1911, N12, N1852);
nand NAND4 (N1913, N1912, N772, N900, N1470);
nand NAND3 (N1914, N1899, N527, N1659);
xor XOR2 (N1915, N1905, N252);
xor XOR2 (N1916, N1908, N1645);
not NOT1 (N1917, N1914);
nand NAND2 (N1918, N1913, N1484);
not NOT1 (N1919, N1873);
and AND2 (N1920, N1916, N650);
nor NOR2 (N1921, N1917, N1095);
or OR2 (N1922, N1920, N1607);
nor NOR4 (N1923, N1919, N1713, N1327, N315);
nand NAND4 (N1924, N1896, N999, N1165, N326);
nor NOR4 (N1925, N1924, N462, N1075, N1530);
or OR4 (N1926, N1901, N1129, N49, N1732);
or OR3 (N1927, N1921, N1764, N1191);
xor XOR2 (N1928, N1925, N419);
and AND4 (N1929, N1922, N1808, N1739, N375);
and AND4 (N1930, N1929, N199, N1059, N762);
and AND2 (N1931, N1926, N1334);
or OR3 (N1932, N1923, N1810, N213);
nor NOR2 (N1933, N1930, N558);
not NOT1 (N1934, N1931);
xor XOR2 (N1935, N1910, N1378);
not NOT1 (N1936, N1933);
not NOT1 (N1937, N1932);
buf BUF1 (N1938, N1935);
or OR4 (N1939, N1936, N236, N1460, N1411);
buf BUF1 (N1940, N1927);
not NOT1 (N1941, N1939);
nand NAND2 (N1942, N1937, N305);
xor XOR2 (N1943, N1907, N776);
buf BUF1 (N1944, N1915);
xor XOR2 (N1945, N1938, N1731);
not NOT1 (N1946, N1934);
nand NAND2 (N1947, N1940, N670);
and AND3 (N1948, N1945, N509, N996);
or OR4 (N1949, N1943, N1028, N1721, N561);
buf BUF1 (N1950, N1909);
and AND2 (N1951, N1918, N1194);
and AND3 (N1952, N1951, N1036, N1427);
and AND2 (N1953, N1952, N1834);
and AND4 (N1954, N1949, N41, N211, N806);
not NOT1 (N1955, N1941);
and AND4 (N1956, N1947, N1167, N250, N568);
nor NOR4 (N1957, N1956, N165, N1150, N866);
and AND4 (N1958, N1946, N1092, N1430, N1263);
or OR2 (N1959, N1954, N376);
nor NOR3 (N1960, N1944, N1697, N1942);
and AND4 (N1961, N52, N479, N737, N1688);
or OR3 (N1962, N1959, N641, N1524);
buf BUF1 (N1963, N1960);
or OR4 (N1964, N1955, N1700, N1129, N388);
xor XOR2 (N1965, N1958, N236);
or OR2 (N1966, N1948, N70);
and AND4 (N1967, N1964, N111, N1793, N1011);
not NOT1 (N1968, N1967);
xor XOR2 (N1969, N1950, N557);
or OR4 (N1970, N1968, N1764, N812, N1537);
xor XOR2 (N1971, N1966, N1001);
or OR2 (N1972, N1963, N1069);
and AND2 (N1973, N1969, N939);
nor NOR2 (N1974, N1953, N300);
and AND4 (N1975, N1957, N730, N507, N1531);
xor XOR2 (N1976, N1965, N1096);
nor NOR4 (N1977, N1970, N1478, N1143, N479);
not NOT1 (N1978, N1977);
not NOT1 (N1979, N1973);
xor XOR2 (N1980, N1979, N1957);
nor NOR3 (N1981, N1962, N14, N976);
and AND3 (N1982, N1975, N1592, N842);
nand NAND3 (N1983, N1981, N1726, N1126);
not NOT1 (N1984, N1928);
not NOT1 (N1985, N1984);
nor NOR2 (N1986, N1971, N932);
and AND2 (N1987, N1982, N851);
not NOT1 (N1988, N1974);
nor NOR2 (N1989, N1983, N1253);
nor NOR2 (N1990, N1980, N1351);
and AND3 (N1991, N1990, N1746, N1291);
nand NAND4 (N1992, N1986, N312, N36, N1535);
nand NAND4 (N1993, N1988, N488, N1233, N906);
or OR4 (N1994, N1972, N1783, N1867, N720);
buf BUF1 (N1995, N1976);
or OR3 (N1996, N1993, N142, N182);
nand NAND2 (N1997, N1995, N1038);
nor NOR3 (N1998, N1987, N166, N210);
or OR3 (N1999, N1991, N422, N1304);
not NOT1 (N2000, N1999);
xor XOR2 (N2001, N1994, N1045);
nand NAND3 (N2002, N1996, N1268, N1579);
or OR2 (N2003, N1997, N200);
xor XOR2 (N2004, N2001, N1957);
not NOT1 (N2005, N1992);
xor XOR2 (N2006, N1985, N666);
nor NOR2 (N2007, N2000, N1580);
not NOT1 (N2008, N2005);
nor NOR3 (N2009, N2008, N1980, N1963);
nor NOR2 (N2010, N2006, N1126);
and AND2 (N2011, N1978, N1136);
nand NAND2 (N2012, N2010, N1922);
and AND3 (N2013, N2002, N473, N67);
xor XOR2 (N2014, N1989, N880);
or OR3 (N2015, N2012, N198, N1477);
buf BUF1 (N2016, N1998);
xor XOR2 (N2017, N2011, N1290);
nand NAND2 (N2018, N2007, N1649);
not NOT1 (N2019, N2018);
not NOT1 (N2020, N2009);
or OR3 (N2021, N2019, N709, N845);
not NOT1 (N2022, N2016);
xor XOR2 (N2023, N1961, N1591);
and AND3 (N2024, N2015, N88, N757);
nor NOR2 (N2025, N2023, N523);
and AND3 (N2026, N2025, N464, N644);
xor XOR2 (N2027, N2020, N1560);
or OR4 (N2028, N2014, N1634, N1281, N1503);
xor XOR2 (N2029, N2013, N573);
nor NOR4 (N2030, N2028, N1847, N745, N551);
and AND3 (N2031, N2017, N1546, N1275);
and AND2 (N2032, N2027, N450);
not NOT1 (N2033, N2026);
nand NAND3 (N2034, N2033, N1823, N678);
buf BUF1 (N2035, N2021);
not NOT1 (N2036, N2031);
and AND3 (N2037, N2004, N125, N1700);
not NOT1 (N2038, N2022);
or OR4 (N2039, N2036, N103, N836, N1712);
buf BUF1 (N2040, N2039);
nand NAND4 (N2041, N2040, N290, N676, N1778);
xor XOR2 (N2042, N2029, N1925);
and AND2 (N2043, N2035, N34);
buf BUF1 (N2044, N2041);
and AND2 (N2045, N2044, N315);
not NOT1 (N2046, N2042);
nand NAND3 (N2047, N2003, N1570, N184);
or OR4 (N2048, N2043, N799, N1971, N918);
or OR4 (N2049, N2046, N1049, N1576, N1567);
buf BUF1 (N2050, N2037);
xor XOR2 (N2051, N2049, N1389);
not NOT1 (N2052, N2024);
not NOT1 (N2053, N2051);
xor XOR2 (N2054, N2032, N528);
nor NOR3 (N2055, N2052, N431, N866);
and AND3 (N2056, N2054, N1177, N2051);
or OR3 (N2057, N2055, N1678, N580);
not NOT1 (N2058, N2047);
not NOT1 (N2059, N2058);
nor NOR2 (N2060, N2045, N833);
not NOT1 (N2061, N2048);
buf BUF1 (N2062, N2056);
nand NAND3 (N2063, N2034, N1540, N1571);
xor XOR2 (N2064, N2059, N568);
not NOT1 (N2065, N2064);
and AND2 (N2066, N2065, N553);
buf BUF1 (N2067, N2063);
and AND4 (N2068, N2060, N1087, N874, N1385);
xor XOR2 (N2069, N2061, N1355);
not NOT1 (N2070, N2050);
nand NAND3 (N2071, N2067, N965, N1122);
xor XOR2 (N2072, N2062, N353);
or OR2 (N2073, N2070, N812);
or OR2 (N2074, N2057, N618);
nand NAND4 (N2075, N2073, N927, N2062, N2006);
buf BUF1 (N2076, N2030);
nor NOR4 (N2077, N2053, N1974, N1022, N211);
nand NAND3 (N2078, N2071, N439, N263);
nor NOR3 (N2079, N2075, N227, N659);
and AND3 (N2080, N2077, N1495, N921);
and AND3 (N2081, N2078, N1691, N1088);
not NOT1 (N2082, N2038);
not NOT1 (N2083, N2074);
and AND3 (N2084, N2083, N1135, N1494);
and AND4 (N2085, N2080, N1949, N1284, N1082);
or OR3 (N2086, N2085, N1685, N1028);
nor NOR4 (N2087, N2072, N1028, N1944, N293);
xor XOR2 (N2088, N2082, N1202);
buf BUF1 (N2089, N2084);
nand NAND2 (N2090, N2089, N1805);
nand NAND2 (N2091, N2081, N2030);
or OR4 (N2092, N2090, N1698, N1825, N1552);
not NOT1 (N2093, N2069);
not NOT1 (N2094, N2088);
xor XOR2 (N2095, N2068, N282);
nand NAND4 (N2096, N2076, N1936, N909, N1600);
buf BUF1 (N2097, N2086);
xor XOR2 (N2098, N2095, N1781);
and AND2 (N2099, N2097, N596);
nor NOR4 (N2100, N2096, N1767, N1071, N916);
nor NOR3 (N2101, N2098, N423, N504);
not NOT1 (N2102, N2087);
xor XOR2 (N2103, N2101, N1898);
and AND4 (N2104, N2094, N1119, N1465, N572);
and AND4 (N2105, N2091, N535, N1218, N10);
not NOT1 (N2106, N2099);
and AND2 (N2107, N2066, N1267);
or OR2 (N2108, N2103, N1130);
or OR4 (N2109, N2104, N1764, N392, N72);
buf BUF1 (N2110, N2106);
and AND3 (N2111, N2092, N689, N1838);
nand NAND2 (N2112, N2093, N104);
and AND2 (N2113, N2108, N890);
buf BUF1 (N2114, N2105);
nand NAND3 (N2115, N2102, N222, N1900);
nor NOR4 (N2116, N2113, N1856, N235, N16);
not NOT1 (N2117, N2107);
nand NAND3 (N2118, N2079, N151, N1717);
xor XOR2 (N2119, N2115, N1083);
buf BUF1 (N2120, N2114);
not NOT1 (N2121, N2100);
nor NOR3 (N2122, N2121, N2066, N565);
xor XOR2 (N2123, N2110, N1805);
not NOT1 (N2124, N2117);
nand NAND3 (N2125, N2111, N1910, N1818);
nand NAND2 (N2126, N2109, N1067);
nor NOR2 (N2127, N2116, N1040);
nor NOR4 (N2128, N2120, N304, N1173, N78);
nand NAND3 (N2129, N2123, N1893, N1052);
not NOT1 (N2130, N2124);
nand NAND3 (N2131, N2127, N484, N1124);
or OR2 (N2132, N2112, N1701);
or OR4 (N2133, N2129, N440, N627, N1056);
xor XOR2 (N2134, N2133, N1576);
not NOT1 (N2135, N2122);
nor NOR3 (N2136, N2119, N683, N147);
nor NOR4 (N2137, N2128, N332, N585, N2007);
nor NOR3 (N2138, N2125, N765, N147);
nor NOR3 (N2139, N2131, N597, N1362);
nor NOR3 (N2140, N2130, N1540, N376);
nand NAND2 (N2141, N2118, N1158);
and AND3 (N2142, N2139, N2040, N1514);
not NOT1 (N2143, N2132);
or OR2 (N2144, N2143, N1012);
buf BUF1 (N2145, N2126);
not NOT1 (N2146, N2145);
nand NAND2 (N2147, N2134, N1157);
and AND2 (N2148, N2135, N1723);
nor NOR3 (N2149, N2137, N84, N1418);
and AND2 (N2150, N2142, N1752);
not NOT1 (N2151, N2138);
nor NOR3 (N2152, N2141, N990, N2001);
nor NOR4 (N2153, N2146, N1904, N1153, N1526);
not NOT1 (N2154, N2150);
not NOT1 (N2155, N2147);
and AND4 (N2156, N2148, N1288, N1300, N1453);
or OR2 (N2157, N2155, N1037);
and AND3 (N2158, N2136, N1616, N2071);
and AND4 (N2159, N2152, N267, N563, N1188);
nor NOR4 (N2160, N2153, N396, N1497, N1564);
not NOT1 (N2161, N2160);
nand NAND4 (N2162, N2157, N319, N1134, N1032);
buf BUF1 (N2163, N2144);
and AND3 (N2164, N2149, N875, N1012);
buf BUF1 (N2165, N2154);
nor NOR2 (N2166, N2158, N344);
buf BUF1 (N2167, N2162);
xor XOR2 (N2168, N2151, N1572);
buf BUF1 (N2169, N2167);
and AND2 (N2170, N2165, N873);
or OR3 (N2171, N2161, N637, N951);
not NOT1 (N2172, N2164);
nand NAND2 (N2173, N2172, N993);
nor NOR3 (N2174, N2171, N442, N1856);
not NOT1 (N2175, N2174);
or OR4 (N2176, N2175, N417, N227, N2035);
and AND3 (N2177, N2168, N777, N1589);
xor XOR2 (N2178, N2166, N1047);
not NOT1 (N2179, N2140);
nand NAND2 (N2180, N2159, N1771);
and AND4 (N2181, N2179, N1021, N1408, N1103);
or OR2 (N2182, N2176, N492);
and AND3 (N2183, N2177, N1484, N873);
nand NAND2 (N2184, N2169, N774);
buf BUF1 (N2185, N2178);
not NOT1 (N2186, N2182);
nand NAND3 (N2187, N2185, N156, N1859);
buf BUF1 (N2188, N2183);
nand NAND3 (N2189, N2181, N809, N34);
or OR3 (N2190, N2163, N1362, N454);
nand NAND2 (N2191, N2190, N716);
buf BUF1 (N2192, N2187);
nand NAND4 (N2193, N2170, N668, N1579, N528);
buf BUF1 (N2194, N2191);
buf BUF1 (N2195, N2194);
nand NAND3 (N2196, N2180, N147, N613);
xor XOR2 (N2197, N2156, N1838);
not NOT1 (N2198, N2195);
buf BUF1 (N2199, N2193);
not NOT1 (N2200, N2199);
nand NAND3 (N2201, N2198, N362, N910);
not NOT1 (N2202, N2184);
not NOT1 (N2203, N2189);
or OR3 (N2204, N2186, N2045, N1180);
xor XOR2 (N2205, N2204, N433);
or OR4 (N2206, N2188, N1781, N1794, N2039);
buf BUF1 (N2207, N2201);
nor NOR3 (N2208, N2203, N1214, N1447);
or OR2 (N2209, N2192, N931);
xor XOR2 (N2210, N2173, N1500);
and AND3 (N2211, N2208, N1200, N1596);
xor XOR2 (N2212, N2205, N457);
buf BUF1 (N2213, N2212);
not NOT1 (N2214, N2202);
nor NOR2 (N2215, N2209, N1356);
xor XOR2 (N2216, N2206, N1177);
not NOT1 (N2217, N2196);
nor NOR4 (N2218, N2216, N1165, N1552, N1370);
xor XOR2 (N2219, N2215, N2162);
buf BUF1 (N2220, N2197);
or OR3 (N2221, N2200, N490, N707);
and AND2 (N2222, N2207, N1621);
xor XOR2 (N2223, N2211, N1882);
nand NAND3 (N2224, N2218, N1646, N1806);
xor XOR2 (N2225, N2219, N300);
or OR4 (N2226, N2221, N341, N1244, N2113);
or OR2 (N2227, N2217, N1509);
nor NOR3 (N2228, N2227, N1375, N1064);
xor XOR2 (N2229, N2222, N2214);
and AND2 (N2230, N56, N148);
nor NOR4 (N2231, N2220, N381, N234, N1144);
buf BUF1 (N2232, N2228);
buf BUF1 (N2233, N2225);
nor NOR3 (N2234, N2210, N727, N340);
nand NAND3 (N2235, N2226, N1346, N1092);
and AND2 (N2236, N2234, N1620);
and AND2 (N2237, N2235, N979);
nand NAND4 (N2238, N2232, N521, N993, N1572);
xor XOR2 (N2239, N2230, N1334);
nand NAND2 (N2240, N2237, N175);
and AND3 (N2241, N2223, N1118, N1059);
or OR2 (N2242, N2238, N1190);
or OR4 (N2243, N2241, N292, N1213, N2212);
xor XOR2 (N2244, N2213, N69);
nand NAND3 (N2245, N2239, N2040, N804);
xor XOR2 (N2246, N2242, N1676);
or OR2 (N2247, N2246, N285);
or OR2 (N2248, N2240, N1552);
not NOT1 (N2249, N2243);
xor XOR2 (N2250, N2224, N628);
xor XOR2 (N2251, N2229, N1895);
buf BUF1 (N2252, N2247);
and AND2 (N2253, N2251, N1020);
nor NOR2 (N2254, N2253, N1238);
and AND2 (N2255, N2254, N1017);
nand NAND3 (N2256, N2252, N742, N1584);
not NOT1 (N2257, N2245);
not NOT1 (N2258, N2231);
and AND3 (N2259, N2257, N2063, N633);
xor XOR2 (N2260, N2250, N1897);
and AND3 (N2261, N2260, N2212, N2057);
not NOT1 (N2262, N2244);
not NOT1 (N2263, N2261);
buf BUF1 (N2264, N2263);
not NOT1 (N2265, N2258);
xor XOR2 (N2266, N2249, N715);
and AND2 (N2267, N2266, N1519);
nand NAND2 (N2268, N2233, N1419);
xor XOR2 (N2269, N2259, N1415);
and AND4 (N2270, N2264, N1022, N1172, N1252);
or OR2 (N2271, N2268, N2242);
nor NOR2 (N2272, N2255, N518);
nand NAND4 (N2273, N2267, N2063, N1041, N614);
not NOT1 (N2274, N2272);
or OR4 (N2275, N2256, N266, N1195, N406);
buf BUF1 (N2276, N2262);
or OR3 (N2277, N2275, N1085, N1782);
xor XOR2 (N2278, N2265, N1287);
and AND3 (N2279, N2276, N1738, N2071);
or OR3 (N2280, N2269, N2112, N228);
buf BUF1 (N2281, N2273);
buf BUF1 (N2282, N2278);
nor NOR2 (N2283, N2277, N1939);
and AND3 (N2284, N2280, N1934, N512);
nand NAND4 (N2285, N2281, N1545, N1706, N2198);
nor NOR2 (N2286, N2279, N1022);
nor NOR4 (N2287, N2270, N2115, N1104, N273);
nor NOR3 (N2288, N2286, N1943, N698);
not NOT1 (N2289, N2285);
not NOT1 (N2290, N2274);
or OR4 (N2291, N2283, N1995, N1593, N1782);
and AND2 (N2292, N2287, N1734);
or OR2 (N2293, N2288, N1387);
and AND2 (N2294, N2248, N2073);
xor XOR2 (N2295, N2284, N1450);
and AND4 (N2296, N2236, N1214, N1915, N2247);
buf BUF1 (N2297, N2289);
or OR3 (N2298, N2290, N170, N2029);
nand NAND3 (N2299, N2293, N695, N159);
xor XOR2 (N2300, N2299, N2177);
and AND4 (N2301, N2296, N522, N342, N1328);
and AND2 (N2302, N2294, N1947);
xor XOR2 (N2303, N2291, N497);
xor XOR2 (N2304, N2282, N1934);
or OR2 (N2305, N2297, N1543);
not NOT1 (N2306, N2301);
and AND4 (N2307, N2292, N1240, N1910, N1958);
or OR4 (N2308, N2295, N2084, N872, N1081);
xor XOR2 (N2309, N2308, N1088);
not NOT1 (N2310, N2302);
xor XOR2 (N2311, N2305, N836);
buf BUF1 (N2312, N2310);
and AND4 (N2313, N2300, N2136, N1713, N944);
nor NOR3 (N2314, N2306, N1030, N1667);
nand NAND4 (N2315, N2311, N979, N93, N235);
or OR2 (N2316, N2307, N2016);
and AND2 (N2317, N2313, N2091);
nand NAND4 (N2318, N2304, N328, N2174, N1118);
or OR4 (N2319, N2314, N948, N1105, N629);
xor XOR2 (N2320, N2316, N388);
xor XOR2 (N2321, N2309, N892);
and AND3 (N2322, N2303, N765, N421);
nand NAND4 (N2323, N2321, N2197, N1542, N440);
nand NAND2 (N2324, N2315, N2290);
not NOT1 (N2325, N2323);
buf BUF1 (N2326, N2271);
nand NAND4 (N2327, N2320, N257, N2114, N2111);
and AND2 (N2328, N2322, N542);
nand NAND4 (N2329, N2328, N669, N1238, N1327);
buf BUF1 (N2330, N2318);
buf BUF1 (N2331, N2330);
xor XOR2 (N2332, N2325, N1564);
and AND2 (N2333, N2317, N407);
nand NAND3 (N2334, N2332, N264, N1895);
and AND3 (N2335, N2298, N926, N1356);
not NOT1 (N2336, N2326);
not NOT1 (N2337, N2331);
buf BUF1 (N2338, N2333);
buf BUF1 (N2339, N2327);
or OR3 (N2340, N2324, N1024, N337);
or OR2 (N2341, N2339, N1924);
xor XOR2 (N2342, N2340, N1405);
buf BUF1 (N2343, N2334);
nand NAND4 (N2344, N2343, N1777, N1559, N618);
not NOT1 (N2345, N2338);
nand NAND4 (N2346, N2336, N2334, N1808, N2328);
nand NAND2 (N2347, N2312, N673);
and AND4 (N2348, N2344, N1713, N1768, N2009);
not NOT1 (N2349, N2329);
or OR2 (N2350, N2341, N407);
nor NOR3 (N2351, N2350, N2063, N411);
buf BUF1 (N2352, N2342);
buf BUF1 (N2353, N2347);
and AND4 (N2354, N2348, N684, N2085, N1757);
xor XOR2 (N2355, N2346, N1301);
and AND2 (N2356, N2355, N981);
and AND4 (N2357, N2354, N2319, N432, N1974);
and AND4 (N2358, N2298, N904, N1995, N643);
xor XOR2 (N2359, N2345, N686);
xor XOR2 (N2360, N2351, N1697);
buf BUF1 (N2361, N2360);
or OR4 (N2362, N2349, N2044, N516, N111);
buf BUF1 (N2363, N2362);
nor NOR3 (N2364, N2335, N1368, N2296);
nor NOR2 (N2365, N2361, N757);
nor NOR3 (N2366, N2364, N778, N276);
buf BUF1 (N2367, N2363);
buf BUF1 (N2368, N2358);
and AND2 (N2369, N2337, N397);
and AND4 (N2370, N2365, N1793, N138, N1871);
or OR2 (N2371, N2367, N1914);
buf BUF1 (N2372, N2368);
buf BUF1 (N2373, N2357);
buf BUF1 (N2374, N2373);
buf BUF1 (N2375, N2370);
nand NAND4 (N2376, N2366, N1958, N209, N358);
and AND2 (N2377, N2375, N1929);
not NOT1 (N2378, N2377);
and AND3 (N2379, N2371, N2192, N1412);
and AND2 (N2380, N2352, N2138);
nand NAND2 (N2381, N2372, N44);
nand NAND3 (N2382, N2353, N1923, N2169);
nand NAND4 (N2383, N2376, N2197, N978, N1570);
nand NAND2 (N2384, N2378, N1825);
not NOT1 (N2385, N2369);
or OR3 (N2386, N2379, N2295, N1967);
or OR3 (N2387, N2386, N1341, N1872);
and AND4 (N2388, N2380, N1000, N511, N2159);
nand NAND2 (N2389, N2382, N2117);
nor NOR4 (N2390, N2381, N1612, N1344, N1138);
not NOT1 (N2391, N2374);
not NOT1 (N2392, N2385);
and AND4 (N2393, N2391, N1773, N824, N913);
not NOT1 (N2394, N2389);
not NOT1 (N2395, N2390);
or OR2 (N2396, N2356, N2200);
not NOT1 (N2397, N2395);
not NOT1 (N2398, N2393);
or OR2 (N2399, N2388, N2108);
not NOT1 (N2400, N2396);
nand NAND3 (N2401, N2399, N1754, N250);
nor NOR3 (N2402, N2392, N687, N268);
nand NAND2 (N2403, N2398, N439);
buf BUF1 (N2404, N2394);
not NOT1 (N2405, N2384);
nor NOR2 (N2406, N2405, N2125);
nand NAND4 (N2407, N2387, N538, N468, N1125);
and AND3 (N2408, N2402, N1456, N2256);
buf BUF1 (N2409, N2403);
nor NOR4 (N2410, N2359, N1697, N1929, N279);
nor NOR2 (N2411, N2410, N563);
nand NAND2 (N2412, N2404, N219);
nand NAND4 (N2413, N2383, N1674, N1031, N1991);
or OR4 (N2414, N2401, N2276, N391, N2260);
not NOT1 (N2415, N2407);
not NOT1 (N2416, N2411);
nor NOR4 (N2417, N2406, N1910, N1069, N1023);
and AND3 (N2418, N2412, N2002, N2059);
nor NOR3 (N2419, N2414, N1980, N1322);
nand NAND2 (N2420, N2415, N403);
nor NOR2 (N2421, N2416, N1556);
and AND3 (N2422, N2413, N1536, N1927);
not NOT1 (N2423, N2418);
and AND4 (N2424, N2409, N1808, N2105, N29);
xor XOR2 (N2425, N2422, N2305);
and AND4 (N2426, N2420, N1114, N863, N2199);
nor NOR3 (N2427, N2426, N2277, N1665);
buf BUF1 (N2428, N2427);
or OR2 (N2429, N2419, N425);
nand NAND4 (N2430, N2408, N338, N2278, N2318);
or OR4 (N2431, N2429, N1416, N2203, N2000);
xor XOR2 (N2432, N2417, N1101);
not NOT1 (N2433, N2425);
nand NAND4 (N2434, N2428, N2290, N245, N1934);
nand NAND4 (N2435, N2397, N596, N35, N274);
nand NAND2 (N2436, N2430, N1325);
not NOT1 (N2437, N2400);
nand NAND4 (N2438, N2435, N651, N1083, N1042);
buf BUF1 (N2439, N2431);
xor XOR2 (N2440, N2424, N24);
xor XOR2 (N2441, N2432, N384);
buf BUF1 (N2442, N2439);
buf BUF1 (N2443, N2434);
and AND2 (N2444, N2436, N2353);
buf BUF1 (N2445, N2438);
nand NAND2 (N2446, N2437, N1307);
or OR3 (N2447, N2441, N2010, N84);
or OR2 (N2448, N2423, N2128);
buf BUF1 (N2449, N2443);
not NOT1 (N2450, N2440);
nor NOR4 (N2451, N2448, N1921, N2320, N1919);
nand NAND2 (N2452, N2450, N1271);
or OR2 (N2453, N2433, N965);
not NOT1 (N2454, N2449);
buf BUF1 (N2455, N2421);
xor XOR2 (N2456, N2453, N1662);
buf BUF1 (N2457, N2452);
and AND2 (N2458, N2447, N2288);
buf BUF1 (N2459, N2444);
nor NOR3 (N2460, N2458, N1724, N930);
not NOT1 (N2461, N2455);
nand NAND3 (N2462, N2451, N221, N2198);
not NOT1 (N2463, N2460);
not NOT1 (N2464, N2446);
nor NOR3 (N2465, N2457, N1332, N1486);
nor NOR3 (N2466, N2465, N2160, N1883);
buf BUF1 (N2467, N2466);
nand NAND3 (N2468, N2464, N702, N1766);
or OR2 (N2469, N2454, N410);
not NOT1 (N2470, N2445);
buf BUF1 (N2471, N2456);
xor XOR2 (N2472, N2461, N1209);
buf BUF1 (N2473, N2471);
and AND3 (N2474, N2467, N1446, N1300);
and AND2 (N2475, N2462, N2098);
and AND3 (N2476, N2442, N1320, N1895);
nor NOR2 (N2477, N2468, N205);
xor XOR2 (N2478, N2476, N1606);
and AND3 (N2479, N2459, N959, N740);
buf BUF1 (N2480, N2475);
not NOT1 (N2481, N2472);
xor XOR2 (N2482, N2477, N2029);
xor XOR2 (N2483, N2469, N2218);
nand NAND3 (N2484, N2474, N274, N1265);
buf BUF1 (N2485, N2483);
nand NAND2 (N2486, N2478, N2317);
buf BUF1 (N2487, N2480);
and AND3 (N2488, N2470, N1470, N223);
not NOT1 (N2489, N2479);
nand NAND3 (N2490, N2484, N948, N69);
not NOT1 (N2491, N2473);
or OR2 (N2492, N2482, N1218);
and AND2 (N2493, N2489, N1563);
nand NAND2 (N2494, N2491, N1412);
nor NOR3 (N2495, N2481, N603, N2341);
not NOT1 (N2496, N2490);
not NOT1 (N2497, N2493);
nor NOR2 (N2498, N2486, N2286);
nand NAND3 (N2499, N2492, N2050, N2174);
or OR2 (N2500, N2488, N1765);
or OR2 (N2501, N2500, N1004);
and AND4 (N2502, N2499, N481, N746, N1001);
nand NAND2 (N2503, N2463, N551);
and AND2 (N2504, N2502, N2106);
or OR4 (N2505, N2498, N1570, N2422, N676);
or OR2 (N2506, N2505, N1337);
buf BUF1 (N2507, N2497);
nand NAND4 (N2508, N2495, N1475, N1896, N220);
nand NAND4 (N2509, N2496, N466, N1811, N1950);
nand NAND3 (N2510, N2506, N967, N2426);
buf BUF1 (N2511, N2487);
and AND3 (N2512, N2510, N1368, N1885);
not NOT1 (N2513, N2485);
xor XOR2 (N2514, N2513, N242);
buf BUF1 (N2515, N2501);
and AND3 (N2516, N2515, N101, N1968);
or OR3 (N2517, N2503, N1255, N1923);
buf BUF1 (N2518, N2507);
nand NAND2 (N2519, N2516, N979);
not NOT1 (N2520, N2509);
xor XOR2 (N2521, N2520, N477);
or OR3 (N2522, N2514, N1760, N1056);
xor XOR2 (N2523, N2518, N502);
or OR2 (N2524, N2494, N1325);
nor NOR4 (N2525, N2512, N386, N1538, N195);
buf BUF1 (N2526, N2511);
nand NAND2 (N2527, N2524, N1158);
nand NAND4 (N2528, N2525, N646, N936, N491);
nor NOR3 (N2529, N2508, N1683, N2207);
not NOT1 (N2530, N2517);
not NOT1 (N2531, N2519);
nor NOR4 (N2532, N2521, N1430, N192, N2300);
buf BUF1 (N2533, N2527);
nor NOR3 (N2534, N2526, N641, N411);
not NOT1 (N2535, N2532);
xor XOR2 (N2536, N2529, N2444);
and AND2 (N2537, N2536, N2259);
and AND3 (N2538, N2522, N2257, N1355);
or OR4 (N2539, N2530, N1241, N2387, N2108);
nand NAND3 (N2540, N2531, N547, N1588);
or OR4 (N2541, N2528, N1392, N481, N1125);
buf BUF1 (N2542, N2541);
nand NAND3 (N2543, N2540, N1768, N744);
or OR3 (N2544, N2542, N359, N1390);
buf BUF1 (N2545, N2537);
or OR4 (N2546, N2543, N99, N1753, N263);
not NOT1 (N2547, N2538);
buf BUF1 (N2548, N2535);
nor NOR3 (N2549, N2545, N2481, N1245);
buf BUF1 (N2550, N2533);
or OR3 (N2551, N2549, N418, N1886);
nor NOR2 (N2552, N2546, N2168);
or OR4 (N2553, N2523, N10, N912, N1735);
nand NAND2 (N2554, N2547, N247);
not NOT1 (N2555, N2539);
nor NOR4 (N2556, N2551, N1579, N2539, N2030);
nand NAND3 (N2557, N2534, N1381, N630);
nor NOR4 (N2558, N2544, N1363, N158, N1813);
nor NOR3 (N2559, N2552, N2512, N1545);
buf BUF1 (N2560, N2548);
and AND4 (N2561, N2560, N1976, N2493, N1380);
and AND4 (N2562, N2504, N1545, N983, N767);
buf BUF1 (N2563, N2561);
buf BUF1 (N2564, N2563);
xor XOR2 (N2565, N2558, N2045);
xor XOR2 (N2566, N2557, N1286);
and AND4 (N2567, N2555, N1903, N1276, N602);
not NOT1 (N2568, N2559);
buf BUF1 (N2569, N2568);
nand NAND2 (N2570, N2550, N413);
nor NOR4 (N2571, N2566, N344, N2310, N1245);
nor NOR2 (N2572, N2564, N1894);
nand NAND2 (N2573, N2554, N582);
or OR2 (N2574, N2565, N1790);
nand NAND2 (N2575, N2574, N2477);
buf BUF1 (N2576, N2553);
buf BUF1 (N2577, N2572);
buf BUF1 (N2578, N2577);
nor NOR2 (N2579, N2569, N1911);
and AND3 (N2580, N2562, N689, N2371);
buf BUF1 (N2581, N2576);
xor XOR2 (N2582, N2580, N512);
nand NAND3 (N2583, N2556, N1132, N108);
and AND3 (N2584, N2571, N1128, N677);
not NOT1 (N2585, N2578);
nor NOR3 (N2586, N2575, N528, N1792);
and AND2 (N2587, N2584, N1138);
or OR4 (N2588, N2586, N777, N1580, N1043);
buf BUF1 (N2589, N2573);
or OR3 (N2590, N2589, N1738, N2135);
xor XOR2 (N2591, N2587, N1510);
or OR2 (N2592, N2582, N1416);
nor NOR3 (N2593, N2588, N360, N738);
nand NAND2 (N2594, N2592, N1111);
xor XOR2 (N2595, N2583, N2231);
and AND3 (N2596, N2570, N954, N547);
or OR2 (N2597, N2595, N334);
and AND2 (N2598, N2567, N1799);
and AND4 (N2599, N2591, N209, N1451, N2387);
buf BUF1 (N2600, N2597);
and AND4 (N2601, N2590, N2107, N2308, N1176);
nand NAND3 (N2602, N2581, N2382, N1628);
nor NOR3 (N2603, N2600, N1692, N1142);
nand NAND3 (N2604, N2594, N1483, N1587);
buf BUF1 (N2605, N2593);
xor XOR2 (N2606, N2598, N192);
buf BUF1 (N2607, N2596);
or OR3 (N2608, N2604, N31, N1212);
nor NOR4 (N2609, N2599, N1872, N1496, N1453);
nand NAND4 (N2610, N2605, N1302, N1428, N738);
nand NAND2 (N2611, N2601, N958);
nor NOR2 (N2612, N2608, N844);
buf BUF1 (N2613, N2607);
or OR2 (N2614, N2613, N2267);
buf BUF1 (N2615, N2611);
buf BUF1 (N2616, N2606);
and AND4 (N2617, N2610, N1684, N1865, N1526);
or OR2 (N2618, N2579, N298);
or OR3 (N2619, N2614, N2530, N1660);
nand NAND4 (N2620, N2612, N428, N1785, N1102);
buf BUF1 (N2621, N2603);
buf BUF1 (N2622, N2618);
or OR2 (N2623, N2585, N2254);
nand NAND4 (N2624, N2615, N530, N684, N2301);
nor NOR2 (N2625, N2621, N980);
nor NOR4 (N2626, N2624, N1197, N1409, N2028);
buf BUF1 (N2627, N2622);
buf BUF1 (N2628, N2609);
nand NAND2 (N2629, N2616, N999);
buf BUF1 (N2630, N2619);
not NOT1 (N2631, N2626);
or OR2 (N2632, N2630, N1245);
and AND4 (N2633, N2625, N1558, N2312, N260);
nand NAND3 (N2634, N2602, N1526, N1052);
buf BUF1 (N2635, N2631);
nand NAND4 (N2636, N2620, N1167, N1710, N2513);
or OR3 (N2637, N2634, N2594, N807);
nand NAND4 (N2638, N2617, N1686, N2373, N1595);
buf BUF1 (N2639, N2638);
or OR2 (N2640, N2636, N60);
or OR4 (N2641, N2635, N1921, N1034, N2328);
and AND4 (N2642, N2627, N1748, N1483, N1102);
and AND2 (N2643, N2640, N188);
or OR2 (N2644, N2643, N86);
not NOT1 (N2645, N2623);
nor NOR3 (N2646, N2644, N2293, N2605);
nor NOR3 (N2647, N2646, N1603, N263);
nor NOR3 (N2648, N2639, N1614, N31);
or OR2 (N2649, N2632, N95);
and AND4 (N2650, N2628, N1780, N1072, N1733);
or OR2 (N2651, N2645, N2608);
not NOT1 (N2652, N2649);
xor XOR2 (N2653, N2651, N915);
buf BUF1 (N2654, N2652);
or OR2 (N2655, N2654, N1431);
and AND3 (N2656, N2629, N2139, N2206);
not NOT1 (N2657, N2641);
nor NOR4 (N2658, N2657, N1257, N194, N1744);
or OR3 (N2659, N2637, N1468, N487);
xor XOR2 (N2660, N2647, N1956);
not NOT1 (N2661, N2650);
and AND3 (N2662, N2661, N1145, N2142);
nand NAND3 (N2663, N2658, N1468, N1733);
not NOT1 (N2664, N2660);
buf BUF1 (N2665, N2663);
nor NOR3 (N2666, N2656, N2189, N2317);
not NOT1 (N2667, N2655);
or OR2 (N2668, N2666, N2021);
not NOT1 (N2669, N2662);
buf BUF1 (N2670, N2665);
or OR2 (N2671, N2633, N1796);
and AND2 (N2672, N2664, N671);
or OR3 (N2673, N2669, N535, N1913);
nand NAND4 (N2674, N2673, N94, N1422, N532);
buf BUF1 (N2675, N2672);
nand NAND2 (N2676, N2671, N2183);
xor XOR2 (N2677, N2648, N301);
xor XOR2 (N2678, N2675, N946);
not NOT1 (N2679, N2670);
or OR3 (N2680, N2678, N1188, N899);
buf BUF1 (N2681, N2674);
nor NOR4 (N2682, N2668, N1986, N2597, N1720);
buf BUF1 (N2683, N2659);
or OR3 (N2684, N2679, N1948, N2577);
not NOT1 (N2685, N2684);
buf BUF1 (N2686, N2642);
nor NOR2 (N2687, N2682, N2644);
not NOT1 (N2688, N2686);
or OR3 (N2689, N2677, N594, N682);
buf BUF1 (N2690, N2687);
and AND3 (N2691, N2676, N1194, N1284);
buf BUF1 (N2692, N2653);
or OR2 (N2693, N2692, N768);
or OR4 (N2694, N2688, N2687, N2249, N2021);
and AND2 (N2695, N2693, N1567);
or OR4 (N2696, N2691, N920, N808, N2450);
nor NOR3 (N2697, N2680, N1001, N723);
not NOT1 (N2698, N2690);
not NOT1 (N2699, N2689);
or OR3 (N2700, N2694, N1293, N427);
and AND4 (N2701, N2683, N1549, N199, N191);
nand NAND4 (N2702, N2681, N2535, N2552, N1671);
xor XOR2 (N2703, N2702, N1915);
buf BUF1 (N2704, N2685);
and AND2 (N2705, N2704, N2336);
buf BUF1 (N2706, N2697);
nor NOR4 (N2707, N2705, N204, N1463, N398);
not NOT1 (N2708, N2707);
xor XOR2 (N2709, N2698, N2537);
xor XOR2 (N2710, N2708, N1456);
nand NAND2 (N2711, N2667, N871);
nor NOR3 (N2712, N2695, N1752, N2247);
and AND2 (N2713, N2711, N1103);
xor XOR2 (N2714, N2699, N592);
nand NAND3 (N2715, N2710, N1904, N1631);
and AND3 (N2716, N2712, N1214, N1926);
buf BUF1 (N2717, N2700);
or OR3 (N2718, N2715, N2221, N2053);
buf BUF1 (N2719, N2696);
xor XOR2 (N2720, N2716, N2537);
buf BUF1 (N2721, N2720);
not NOT1 (N2722, N2717);
nand NAND4 (N2723, N2714, N502, N720, N860);
nand NAND4 (N2724, N2713, N1731, N801, N1457);
buf BUF1 (N2725, N2706);
nor NOR2 (N2726, N2701, N92);
nor NOR3 (N2727, N2709, N2284, N1467);
nor NOR2 (N2728, N2724, N1171);
buf BUF1 (N2729, N2728);
nor NOR3 (N2730, N2721, N2027, N2301);
xor XOR2 (N2731, N2725, N1406);
or OR3 (N2732, N2718, N42, N2417);
nand NAND3 (N2733, N2731, N879, N2693);
not NOT1 (N2734, N2729);
buf BUF1 (N2735, N2719);
buf BUF1 (N2736, N2730);
nor NOR2 (N2737, N2727, N2355);
buf BUF1 (N2738, N2722);
not NOT1 (N2739, N2703);
xor XOR2 (N2740, N2723, N1287);
buf BUF1 (N2741, N2738);
not NOT1 (N2742, N2735);
nand NAND2 (N2743, N2726, N2549);
not NOT1 (N2744, N2737);
xor XOR2 (N2745, N2733, N127);
xor XOR2 (N2746, N2736, N467);
xor XOR2 (N2747, N2740, N2135);
buf BUF1 (N2748, N2732);
buf BUF1 (N2749, N2734);
xor XOR2 (N2750, N2747, N2452);
not NOT1 (N2751, N2742);
buf BUF1 (N2752, N2743);
buf BUF1 (N2753, N2751);
buf BUF1 (N2754, N2741);
not NOT1 (N2755, N2749);
and AND3 (N2756, N2754, N1564, N2753);
xor XOR2 (N2757, N2590, N598);
xor XOR2 (N2758, N2744, N978);
xor XOR2 (N2759, N2755, N1766);
not NOT1 (N2760, N2748);
and AND2 (N2761, N2750, N2027);
or OR3 (N2762, N2760, N404, N406);
and AND2 (N2763, N2746, N2014);
not NOT1 (N2764, N2745);
and AND4 (N2765, N2762, N2449, N701, N1532);
nor NOR2 (N2766, N2757, N656);
xor XOR2 (N2767, N2759, N1834);
or OR3 (N2768, N2767, N1103, N1759);
and AND3 (N2769, N2766, N453, N1627);
nor NOR2 (N2770, N2756, N1409);
buf BUF1 (N2771, N2763);
not NOT1 (N2772, N2761);
and AND3 (N2773, N2752, N1584, N438);
and AND3 (N2774, N2773, N2159, N596);
nand NAND4 (N2775, N2769, N231, N2247, N1531);
buf BUF1 (N2776, N2758);
and AND4 (N2777, N2771, N1448, N2049, N2528);
not NOT1 (N2778, N2777);
buf BUF1 (N2779, N2765);
and AND2 (N2780, N2770, N2379);
or OR2 (N2781, N2739, N2157);
nand NAND2 (N2782, N2778, N1295);
not NOT1 (N2783, N2775);
nor NOR2 (N2784, N2774, N1449);
nand NAND4 (N2785, N2764, N177, N359, N538);
or OR4 (N2786, N2785, N8, N1935, N892);
and AND4 (N2787, N2776, N1460, N1301, N1368);
nor NOR2 (N2788, N2782, N2538);
buf BUF1 (N2789, N2779);
xor XOR2 (N2790, N2780, N2046);
xor XOR2 (N2791, N2784, N2511);
buf BUF1 (N2792, N2781);
buf BUF1 (N2793, N2789);
buf BUF1 (N2794, N2791);
and AND3 (N2795, N2768, N1491, N309);
or OR3 (N2796, N2794, N857, N529);
nand NAND2 (N2797, N2792, N1978);
or OR4 (N2798, N2787, N667, N41, N1);
not NOT1 (N2799, N2772);
buf BUF1 (N2800, N2799);
or OR3 (N2801, N2800, N50, N496);
nor NOR4 (N2802, N2795, N2313, N1446, N1402);
nand NAND3 (N2803, N2802, N1783, N1454);
not NOT1 (N2804, N2788);
nor NOR2 (N2805, N2801, N1241);
nor NOR2 (N2806, N2803, N1911);
nand NAND3 (N2807, N2783, N2463, N1450);
nor NOR3 (N2808, N2806, N1062, N539);
nand NAND4 (N2809, N2808, N773, N990, N1517);
buf BUF1 (N2810, N2796);
not NOT1 (N2811, N2793);
buf BUF1 (N2812, N2810);
not NOT1 (N2813, N2811);
or OR4 (N2814, N2797, N1324, N1813, N875);
not NOT1 (N2815, N2807);
or OR4 (N2816, N2790, N1341, N1483, N1657);
and AND2 (N2817, N2812, N1865);
and AND2 (N2818, N2798, N1842);
nor NOR3 (N2819, N2805, N1233, N2293);
or OR3 (N2820, N2819, N2384, N2212);
nand NAND2 (N2821, N2786, N2553);
nor NOR3 (N2822, N2821, N1764, N2810);
or OR4 (N2823, N2813, N2648, N2026, N195);
nor NOR4 (N2824, N2817, N2607, N58, N1164);
or OR3 (N2825, N2809, N1146, N1476);
xor XOR2 (N2826, N2814, N1047);
not NOT1 (N2827, N2804);
nor NOR4 (N2828, N2824, N2450, N2231, N1343);
xor XOR2 (N2829, N2823, N178);
buf BUF1 (N2830, N2829);
or OR2 (N2831, N2827, N2278);
not NOT1 (N2832, N2826);
xor XOR2 (N2833, N2825, N913);
and AND4 (N2834, N2831, N156, N1403, N1224);
buf BUF1 (N2835, N2832);
nand NAND3 (N2836, N2828, N1430, N1905);
or OR3 (N2837, N2833, N2502, N308);
buf BUF1 (N2838, N2816);
nor NOR3 (N2839, N2834, N1640, N1646);
or OR3 (N2840, N2818, N1970, N1142);
nand NAND2 (N2841, N2815, N487);
nand NAND3 (N2842, N2838, N2154, N1330);
and AND2 (N2843, N2839, N2002);
nand NAND2 (N2844, N2836, N2577);
nand NAND2 (N2845, N2822, N1019);
buf BUF1 (N2846, N2820);
xor XOR2 (N2847, N2835, N1675);
not NOT1 (N2848, N2844);
or OR4 (N2849, N2841, N1331, N147, N1471);
not NOT1 (N2850, N2837);
nand NAND4 (N2851, N2847, N139, N1002, N1932);
or OR4 (N2852, N2849, N614, N1298, N1426);
nand NAND4 (N2853, N2840, N440, N2363, N810);
not NOT1 (N2854, N2846);
buf BUF1 (N2855, N2852);
nor NOR3 (N2856, N2851, N1612, N2344);
nor NOR2 (N2857, N2853, N2605);
nor NOR4 (N2858, N2845, N2204, N1195, N943);
or OR3 (N2859, N2854, N2440, N1426);
or OR4 (N2860, N2850, N2747, N2457, N1717);
nor NOR3 (N2861, N2855, N231, N2353);
buf BUF1 (N2862, N2858);
and AND4 (N2863, N2862, N2283, N1985, N2587);
or OR3 (N2864, N2848, N1719, N1637);
nor NOR2 (N2865, N2843, N2790);
nand NAND4 (N2866, N2860, N183, N2022, N447);
nor NOR2 (N2867, N2857, N527);
nor NOR3 (N2868, N2867, N174, N936);
xor XOR2 (N2869, N2861, N600);
nor NOR4 (N2870, N2868, N641, N494, N2275);
buf BUF1 (N2871, N2863);
or OR3 (N2872, N2869, N7, N1263);
nand NAND2 (N2873, N2842, N2806);
buf BUF1 (N2874, N2859);
nand NAND4 (N2875, N2865, N1031, N1749, N126);
or OR4 (N2876, N2871, N397, N1450, N1360);
or OR2 (N2877, N2830, N20);
nor NOR4 (N2878, N2872, N1019, N776, N301);
and AND4 (N2879, N2864, N662, N2162, N2712);
nor NOR2 (N2880, N2856, N2470);
buf BUF1 (N2881, N2873);
nor NOR3 (N2882, N2879, N2094, N1194);
nor NOR2 (N2883, N2876, N2818);
nor NOR3 (N2884, N2866, N17, N1237);
or OR3 (N2885, N2884, N2630, N549);
nand NAND3 (N2886, N2875, N1693, N181);
buf BUF1 (N2887, N2882);
and AND4 (N2888, N2881, N808, N1023, N795);
not NOT1 (N2889, N2887);
nor NOR2 (N2890, N2888, N1980);
nand NAND2 (N2891, N2877, N184);
and AND3 (N2892, N2880, N87, N1676);
xor XOR2 (N2893, N2891, N1590);
and AND2 (N2894, N2878, N2823);
nand NAND3 (N2895, N2892, N2694, N2779);
nand NAND2 (N2896, N2894, N1220);
not NOT1 (N2897, N2896);
and AND3 (N2898, N2893, N570, N2714);
xor XOR2 (N2899, N2890, N1213);
or OR4 (N2900, N2897, N539, N1818, N1069);
not NOT1 (N2901, N2874);
not NOT1 (N2902, N2900);
buf BUF1 (N2903, N2889);
nand NAND4 (N2904, N2898, N1174, N292, N662);
nand NAND2 (N2905, N2870, N2830);
nor NOR2 (N2906, N2886, N1918);
nor NOR3 (N2907, N2904, N364, N305);
nor NOR3 (N2908, N2907, N2498, N2691);
buf BUF1 (N2909, N2899);
not NOT1 (N2910, N2903);
nand NAND3 (N2911, N2883, N2113, N2786);
nor NOR3 (N2912, N2885, N951, N690);
buf BUF1 (N2913, N2895);
buf BUF1 (N2914, N2910);
nor NOR3 (N2915, N2913, N2712, N2885);
not NOT1 (N2916, N2909);
buf BUF1 (N2917, N2914);
not NOT1 (N2918, N2908);
and AND4 (N2919, N2905, N1524, N2412, N835);
nand NAND3 (N2920, N2919, N35, N1537);
or OR3 (N2921, N2920, N1182, N680);
xor XOR2 (N2922, N2916, N750);
and AND3 (N2923, N2912, N1691, N2007);
xor XOR2 (N2924, N2917, N1840);
not NOT1 (N2925, N2922);
not NOT1 (N2926, N2906);
buf BUF1 (N2927, N2925);
buf BUF1 (N2928, N2923);
xor XOR2 (N2929, N2926, N474);
or OR4 (N2930, N2927, N2723, N2558, N341);
or OR3 (N2931, N2915, N2380, N1625);
and AND2 (N2932, N2930, N1125);
nor NOR3 (N2933, N2928, N2801, N1136);
nor NOR3 (N2934, N2918, N2172, N184);
nor NOR2 (N2935, N2932, N1161);
nand NAND3 (N2936, N2921, N619, N1549);
or OR3 (N2937, N2911, N1642, N2932);
nor NOR3 (N2938, N2902, N2596, N2451);
xor XOR2 (N2939, N2937, N1282);
nor NOR2 (N2940, N2931, N890);
and AND4 (N2941, N2935, N1839, N2248, N2331);
or OR2 (N2942, N2901, N2218);
nor NOR2 (N2943, N2929, N458);
or OR4 (N2944, N2933, N2822, N2409, N2345);
nor NOR3 (N2945, N2924, N2473, N2771);
xor XOR2 (N2946, N2936, N919);
nor NOR2 (N2947, N2939, N946);
xor XOR2 (N2948, N2942, N313);
not NOT1 (N2949, N2946);
or OR3 (N2950, N2940, N2251, N558);
buf BUF1 (N2951, N2943);
nor NOR4 (N2952, N2950, N2582, N556, N137);
buf BUF1 (N2953, N2951);
buf BUF1 (N2954, N2941);
nor NOR3 (N2955, N2934, N2461, N500);
not NOT1 (N2956, N2953);
and AND3 (N2957, N2952, N431, N1999);
nand NAND2 (N2958, N2948, N375);
and AND4 (N2959, N2958, N797, N1374, N1317);
buf BUF1 (N2960, N2957);
not NOT1 (N2961, N2944);
xor XOR2 (N2962, N2938, N2043);
nor NOR3 (N2963, N2960, N891, N2864);
or OR2 (N2964, N2961, N1189);
buf BUF1 (N2965, N2962);
nand NAND3 (N2966, N2954, N20, N1591);
nor NOR4 (N2967, N2956, N2331, N2907, N783);
and AND4 (N2968, N2964, N784, N1556, N1245);
nor NOR4 (N2969, N2965, N1538, N2792, N1505);
nand NAND2 (N2970, N2945, N1679);
xor XOR2 (N2971, N2968, N2375);
nand NAND2 (N2972, N2971, N305);
not NOT1 (N2973, N2966);
not NOT1 (N2974, N2963);
nor NOR3 (N2975, N2955, N261, N2722);
or OR3 (N2976, N2947, N982, N1466);
buf BUF1 (N2977, N2974);
or OR2 (N2978, N2972, N2028);
not NOT1 (N2979, N2975);
nand NAND3 (N2980, N2976, N76, N2043);
not NOT1 (N2981, N2973);
and AND4 (N2982, N2967, N1480, N1281, N2560);
nor NOR3 (N2983, N2949, N1947, N1299);
not NOT1 (N2984, N2981);
buf BUF1 (N2985, N2959);
nor NOR2 (N2986, N2977, N1633);
or OR4 (N2987, N2983, N1870, N1429, N1702);
and AND2 (N2988, N2979, N1161);
nand NAND3 (N2989, N2984, N2528, N78);
or OR4 (N2990, N2986, N872, N1607, N948);
or OR3 (N2991, N2990, N1085, N1091);
and AND3 (N2992, N2985, N1386, N721);
nand NAND4 (N2993, N2987, N2391, N1314, N1675);
buf BUF1 (N2994, N2980);
or OR3 (N2995, N2978, N2870, N1089);
nor NOR2 (N2996, N2970, N1358);
and AND4 (N2997, N2995, N2474, N148, N1504);
or OR3 (N2998, N2988, N1720, N2585);
xor XOR2 (N2999, N2996, N2823);
nand NAND3 (N3000, N2997, N682, N696);
not NOT1 (N3001, N2991);
nor NOR3 (N3002, N2969, N307, N245);
and AND3 (N3003, N2998, N1678, N1546);
or OR3 (N3004, N2989, N1039, N1598);
buf BUF1 (N3005, N2993);
not NOT1 (N3006, N2999);
nor NOR4 (N3007, N2982, N566, N438, N2458);
and AND2 (N3008, N3007, N2309);
nand NAND4 (N3009, N3006, N358, N1850, N1081);
buf BUF1 (N3010, N3005);
and AND2 (N3011, N3008, N1409);
not NOT1 (N3012, N3003);
nand NAND2 (N3013, N3010, N1884);
nor NOR4 (N3014, N3002, N795, N2757, N557);
nor NOR4 (N3015, N3001, N1575, N509, N1999);
not NOT1 (N3016, N3000);
and AND3 (N3017, N3015, N2745, N294);
not NOT1 (N3018, N3009);
xor XOR2 (N3019, N3013, N1817);
and AND4 (N3020, N3014, N1482, N250, N2248);
and AND3 (N3021, N3011, N51, N737);
xor XOR2 (N3022, N3020, N654);
or OR2 (N3023, N3016, N285);
buf BUF1 (N3024, N3019);
nand NAND2 (N3025, N3021, N2287);
not NOT1 (N3026, N2992);
not NOT1 (N3027, N3022);
buf BUF1 (N3028, N3027);
or OR2 (N3029, N3024, N99);
not NOT1 (N3030, N3018);
not NOT1 (N3031, N3026);
and AND4 (N3032, N3004, N1083, N2728, N2829);
nand NAND3 (N3033, N3029, N1522, N636);
buf BUF1 (N3034, N3033);
buf BUF1 (N3035, N3030);
nor NOR4 (N3036, N2994, N404, N2215, N2222);
buf BUF1 (N3037, N3034);
buf BUF1 (N3038, N3035);
nand NAND2 (N3039, N3017, N1068);
xor XOR2 (N3040, N3012, N1323);
xor XOR2 (N3041, N3025, N2864);
xor XOR2 (N3042, N3037, N634);
buf BUF1 (N3043, N3036);
or OR4 (N3044, N3032, N443, N495, N1953);
nand NAND2 (N3045, N3038, N1954);
nor NOR4 (N3046, N3031, N703, N1321, N2775);
buf BUF1 (N3047, N3023);
not NOT1 (N3048, N3046);
xor XOR2 (N3049, N3044, N973);
buf BUF1 (N3050, N3040);
not NOT1 (N3051, N3041);
and AND4 (N3052, N3042, N55, N675, N1081);
xor XOR2 (N3053, N3043, N1288);
or OR2 (N3054, N3047, N2485);
or OR3 (N3055, N3052, N2795, N2654);
nand NAND4 (N3056, N3045, N717, N2160, N1502);
and AND2 (N3057, N3054, N133);
not NOT1 (N3058, N3049);
or OR4 (N3059, N3056, N1688, N2189, N2075);
nand NAND2 (N3060, N3048, N458);
not NOT1 (N3061, N3051);
and AND3 (N3062, N3050, N320, N2203);
buf BUF1 (N3063, N3060);
not NOT1 (N3064, N3062);
xor XOR2 (N3065, N3061, N2164);
xor XOR2 (N3066, N3057, N2846);
and AND2 (N3067, N3028, N689);
nor NOR2 (N3068, N3055, N1674);
and AND4 (N3069, N3067, N2092, N1493, N270);
and AND4 (N3070, N3069, N1808, N972, N1484);
xor XOR2 (N3071, N3065, N2429);
xor XOR2 (N3072, N3039, N2846);
nand NAND2 (N3073, N3066, N332);
xor XOR2 (N3074, N3071, N1971);
nand NAND4 (N3075, N3068, N3039, N1274, N2456);
xor XOR2 (N3076, N3074, N2651);
buf BUF1 (N3077, N3058);
or OR2 (N3078, N3053, N2331);
nand NAND3 (N3079, N3059, N1685, N2805);
xor XOR2 (N3080, N3079, N275);
nand NAND4 (N3081, N3076, N1764, N441, N2372);
or OR2 (N3082, N3075, N628);
or OR2 (N3083, N3073, N932);
or OR3 (N3084, N3077, N2282, N2713);
not NOT1 (N3085, N3063);
xor XOR2 (N3086, N3078, N1983);
buf BUF1 (N3087, N3080);
nand NAND3 (N3088, N3086, N263, N339);
xor XOR2 (N3089, N3083, N1898);
buf BUF1 (N3090, N3088);
or OR3 (N3091, N3072, N1765, N1584);
nand NAND2 (N3092, N3085, N273);
not NOT1 (N3093, N3084);
nand NAND2 (N3094, N3064, N1928);
not NOT1 (N3095, N3070);
not NOT1 (N3096, N3092);
xor XOR2 (N3097, N3095, N2081);
not NOT1 (N3098, N3081);
xor XOR2 (N3099, N3094, N119);
nand NAND2 (N3100, N3096, N1577);
buf BUF1 (N3101, N3091);
and AND2 (N3102, N3093, N47);
not NOT1 (N3103, N3102);
and AND2 (N3104, N3101, N181);
and AND3 (N3105, N3097, N2108, N2128);
nor NOR4 (N3106, N3104, N2353, N1255, N2679);
not NOT1 (N3107, N3103);
buf BUF1 (N3108, N3100);
xor XOR2 (N3109, N3106, N1592);
buf BUF1 (N3110, N3109);
xor XOR2 (N3111, N3105, N1796);
and AND2 (N3112, N3099, N527);
buf BUF1 (N3113, N3090);
buf BUF1 (N3114, N3108);
and AND3 (N3115, N3112, N2972, N2905);
nor NOR3 (N3116, N3114, N672, N1187);
xor XOR2 (N3117, N3113, N1582);
and AND4 (N3118, N3082, N2147, N110, N1084);
not NOT1 (N3119, N3089);
and AND3 (N3120, N3107, N291, N667);
or OR3 (N3121, N3111, N1058, N2329);
or OR3 (N3122, N3121, N2055, N2199);
buf BUF1 (N3123, N3118);
nor NOR2 (N3124, N3120, N204);
not NOT1 (N3125, N3116);
or OR4 (N3126, N3124, N2910, N1060, N2985);
not NOT1 (N3127, N3115);
and AND4 (N3128, N3125, N2099, N2863, N99);
xor XOR2 (N3129, N3123, N1648);
and AND3 (N3130, N3087, N239, N1962);
or OR2 (N3131, N3126, N1636);
nor NOR2 (N3132, N3122, N29);
buf BUF1 (N3133, N3127);
not NOT1 (N3134, N3133);
nor NOR3 (N3135, N3098, N2232, N2100);
nand NAND4 (N3136, N3135, N633, N2249, N2983);
nand NAND3 (N3137, N3136, N1568, N2642);
and AND2 (N3138, N3119, N1704);
or OR2 (N3139, N3130, N1918);
xor XOR2 (N3140, N3138, N2093);
buf BUF1 (N3141, N3131);
nand NAND2 (N3142, N3140, N218);
not NOT1 (N3143, N3129);
nor NOR4 (N3144, N3132, N975, N3084, N1655);
buf BUF1 (N3145, N3141);
xor XOR2 (N3146, N3110, N1982);
nor NOR3 (N3147, N3145, N1193, N2979);
or OR4 (N3148, N3147, N2604, N1074, N3007);
and AND4 (N3149, N3137, N807, N2092, N392);
xor XOR2 (N3150, N3149, N2967);
not NOT1 (N3151, N3146);
not NOT1 (N3152, N3143);
not NOT1 (N3153, N3152);
not NOT1 (N3154, N3150);
nor NOR4 (N3155, N3148, N1639, N2394, N476);
nor NOR2 (N3156, N3155, N1949);
or OR3 (N3157, N3117, N2300, N2297);
not NOT1 (N3158, N3142);
not NOT1 (N3159, N3158);
not NOT1 (N3160, N3154);
nor NOR4 (N3161, N3128, N428, N1140, N2273);
nand NAND2 (N3162, N3153, N2177);
nand NAND4 (N3163, N3162, N928, N1451, N614);
and AND4 (N3164, N3159, N662, N1119, N1344);
or OR3 (N3165, N3139, N503, N1603);
not NOT1 (N3166, N3163);
not NOT1 (N3167, N3164);
and AND2 (N3168, N3156, N760);
not NOT1 (N3169, N3144);
not NOT1 (N3170, N3151);
or OR3 (N3171, N3160, N939, N1922);
nand NAND3 (N3172, N3157, N753, N255);
nand NAND2 (N3173, N3168, N844);
nand NAND2 (N3174, N3170, N1668);
buf BUF1 (N3175, N3167);
not NOT1 (N3176, N3161);
xor XOR2 (N3177, N3173, N3114);
buf BUF1 (N3178, N3177);
buf BUF1 (N3179, N3171);
nor NOR2 (N3180, N3166, N1455);
nand NAND4 (N3181, N3178, N246, N1600, N582);
or OR3 (N3182, N3134, N3025, N2962);
nor NOR2 (N3183, N3182, N2255);
xor XOR2 (N3184, N3183, N167);
buf BUF1 (N3185, N3174);
not NOT1 (N3186, N3176);
nor NOR3 (N3187, N3181, N915, N1187);
xor XOR2 (N3188, N3180, N835);
nor NOR3 (N3189, N3187, N1188, N1451);
and AND3 (N3190, N3188, N1819, N2754);
or OR3 (N3191, N3172, N1516, N1245);
xor XOR2 (N3192, N3165, N1756);
buf BUF1 (N3193, N3175);
xor XOR2 (N3194, N3189, N1774);
buf BUF1 (N3195, N3184);
not NOT1 (N3196, N3193);
nand NAND4 (N3197, N3186, N1735, N2364, N2492);
and AND3 (N3198, N3185, N41, N2621);
xor XOR2 (N3199, N3191, N1894);
or OR3 (N3200, N3192, N1302, N793);
buf BUF1 (N3201, N3190);
buf BUF1 (N3202, N3198);
nand NAND4 (N3203, N3200, N1748, N722, N2001);
or OR4 (N3204, N3196, N30, N1782, N3177);
and AND4 (N3205, N3203, N1149, N2918, N2857);
xor XOR2 (N3206, N3195, N2521);
and AND4 (N3207, N3199, N1583, N214, N2743);
buf BUF1 (N3208, N3197);
nor NOR2 (N3209, N3169, N1832);
and AND3 (N3210, N3205, N2341, N1942);
xor XOR2 (N3211, N3204, N1455);
nand NAND4 (N3212, N3206, N74, N1953, N2773);
xor XOR2 (N3213, N3212, N2910);
nor NOR2 (N3214, N3194, N1134);
nor NOR4 (N3215, N3209, N1462, N2118, N1150);
nor NOR2 (N3216, N3214, N2760);
xor XOR2 (N3217, N3216, N2419);
not NOT1 (N3218, N3201);
xor XOR2 (N3219, N3215, N3204);
or OR4 (N3220, N3218, N2118, N121, N2679);
nor NOR4 (N3221, N3217, N1530, N2934, N36);
not NOT1 (N3222, N3213);
nor NOR3 (N3223, N3208, N1458, N427);
nor NOR2 (N3224, N3207, N1557);
nor NOR3 (N3225, N3219, N39, N1119);
nand NAND3 (N3226, N3211, N1390, N2537);
not NOT1 (N3227, N3222);
nor NOR4 (N3228, N3210, N2969, N653, N3224);
nor NOR4 (N3229, N1812, N1489, N2554, N2840);
nand NAND3 (N3230, N3223, N581, N1874);
and AND2 (N3231, N3230, N72);
not NOT1 (N3232, N3179);
and AND2 (N3233, N3220, N1943);
not NOT1 (N3234, N3202);
nand NAND3 (N3235, N3228, N924, N2839);
nand NAND3 (N3236, N3235, N846, N1984);
xor XOR2 (N3237, N3234, N1322);
nand NAND2 (N3238, N3231, N2808);
buf BUF1 (N3239, N3233);
not NOT1 (N3240, N3225);
and AND3 (N3241, N3240, N2374, N493);
buf BUF1 (N3242, N3227);
xor XOR2 (N3243, N3238, N2858);
and AND2 (N3244, N3241, N1006);
and AND3 (N3245, N3229, N2153, N1739);
not NOT1 (N3246, N3237);
not NOT1 (N3247, N3226);
xor XOR2 (N3248, N3244, N1281);
or OR2 (N3249, N3239, N2971);
nor NOR3 (N3250, N3221, N2655, N3006);
xor XOR2 (N3251, N3247, N2899);
nor NOR3 (N3252, N3249, N2598, N445);
nor NOR4 (N3253, N3250, N2, N1245, N3199);
nor NOR3 (N3254, N3253, N1550, N2683);
xor XOR2 (N3255, N3248, N2100);
not NOT1 (N3256, N3246);
nand NAND4 (N3257, N3243, N350, N1715, N3086);
and AND4 (N3258, N3252, N945, N961, N1859);
nor NOR2 (N3259, N3236, N953);
and AND2 (N3260, N3256, N2389);
nand NAND4 (N3261, N3258, N1497, N1148, N1640);
buf BUF1 (N3262, N3242);
and AND3 (N3263, N3260, N748, N2102);
xor XOR2 (N3264, N3259, N395);
nor NOR2 (N3265, N3263, N677);
not NOT1 (N3266, N3251);
xor XOR2 (N3267, N3265, N721);
and AND2 (N3268, N3261, N771);
or OR4 (N3269, N3268, N75, N1193, N839);
or OR3 (N3270, N3257, N2469, N497);
not NOT1 (N3271, N3232);
or OR2 (N3272, N3245, N1302);
not NOT1 (N3273, N3266);
and AND3 (N3274, N3269, N1539, N674);
nor NOR4 (N3275, N3274, N352, N1689, N802);
or OR3 (N3276, N3270, N2079, N1954);
or OR4 (N3277, N3276, N1210, N1938, N194);
or OR4 (N3278, N3273, N956, N1115, N2936);
and AND4 (N3279, N3271, N1303, N1181, N1614);
nand NAND3 (N3280, N3262, N1044, N2040);
or OR3 (N3281, N3267, N1844, N1964);
xor XOR2 (N3282, N3254, N2281);
xor XOR2 (N3283, N3281, N3106);
nand NAND2 (N3284, N3278, N2141);
not NOT1 (N3285, N3282);
nand NAND3 (N3286, N3272, N1814, N3192);
not NOT1 (N3287, N3264);
or OR2 (N3288, N3255, N1136);
nor NOR2 (N3289, N3287, N645);
not NOT1 (N3290, N3286);
nand NAND2 (N3291, N3280, N2168);
not NOT1 (N3292, N3291);
xor XOR2 (N3293, N3285, N1240);
and AND4 (N3294, N3279, N1751, N2222, N648);
nand NAND2 (N3295, N3294, N2491);
or OR3 (N3296, N3277, N1236, N1440);
buf BUF1 (N3297, N3290);
xor XOR2 (N3298, N3296, N1703);
or OR3 (N3299, N3289, N2715, N1957);
and AND2 (N3300, N3275, N1215);
and AND2 (N3301, N3298, N2204);
nor NOR3 (N3302, N3293, N2408, N1951);
xor XOR2 (N3303, N3292, N280);
xor XOR2 (N3304, N3302, N85);
and AND4 (N3305, N3303, N2799, N2219, N2565);
xor XOR2 (N3306, N3299, N141);
or OR2 (N3307, N3295, N329);
and AND4 (N3308, N3306, N2636, N1693, N2898);
or OR2 (N3309, N3300, N1094);
nand NAND3 (N3310, N3284, N3095, N2022);
buf BUF1 (N3311, N3304);
buf BUF1 (N3312, N3301);
and AND3 (N3313, N3309, N2840, N1336);
and AND4 (N3314, N3307, N1598, N2659, N301);
xor XOR2 (N3315, N3305, N176);
nor NOR3 (N3316, N3297, N2109, N1268);
nor NOR3 (N3317, N3312, N1991, N1269);
nor NOR2 (N3318, N3317, N2842);
xor XOR2 (N3319, N3314, N1616);
not NOT1 (N3320, N3315);
buf BUF1 (N3321, N3311);
not NOT1 (N3322, N3320);
nor NOR3 (N3323, N3310, N1550, N2326);
xor XOR2 (N3324, N3323, N756);
or OR3 (N3325, N3316, N3311, N758);
buf BUF1 (N3326, N3313);
or OR4 (N3327, N3325, N2559, N2416, N1157);
buf BUF1 (N3328, N3319);
nand NAND2 (N3329, N3308, N1165);
not NOT1 (N3330, N3322);
nor NOR3 (N3331, N3326, N3044, N420);
xor XOR2 (N3332, N3321, N1043);
and AND3 (N3333, N3330, N1426, N2701);
and AND4 (N3334, N3331, N840, N1383, N2994);
xor XOR2 (N3335, N3283, N1840);
xor XOR2 (N3336, N3288, N2759);
buf BUF1 (N3337, N3318);
or OR3 (N3338, N3334, N2854, N331);
xor XOR2 (N3339, N3333, N2135);
buf BUF1 (N3340, N3337);
and AND4 (N3341, N3329, N962, N1823, N924);
nor NOR3 (N3342, N3341, N2481, N1868);
nand NAND4 (N3343, N3338, N2122, N1050, N1663);
or OR4 (N3344, N3339, N1908, N1885, N1677);
or OR2 (N3345, N3342, N714);
or OR4 (N3346, N3340, N3284, N2773, N2556);
or OR2 (N3347, N3324, N517);
or OR3 (N3348, N3335, N884, N364);
not NOT1 (N3349, N3343);
not NOT1 (N3350, N3347);
nand NAND4 (N3351, N3328, N3157, N853, N1896);
not NOT1 (N3352, N3351);
nand NAND2 (N3353, N3336, N3007);
not NOT1 (N3354, N3346);
or OR4 (N3355, N3349, N490, N3173, N1529);
nor NOR3 (N3356, N3350, N358, N814);
and AND3 (N3357, N3348, N27, N723);
xor XOR2 (N3358, N3352, N455);
nor NOR2 (N3359, N3356, N8);
not NOT1 (N3360, N3344);
or OR4 (N3361, N3358, N553, N2335, N203);
buf BUF1 (N3362, N3332);
buf BUF1 (N3363, N3355);
and AND4 (N3364, N3361, N78, N1876, N388);
xor XOR2 (N3365, N3364, N2729);
or OR2 (N3366, N3345, N2087);
xor XOR2 (N3367, N3354, N790);
not NOT1 (N3368, N3366);
buf BUF1 (N3369, N3359);
and AND2 (N3370, N3369, N3006);
or OR2 (N3371, N3353, N2545);
and AND3 (N3372, N3362, N3021, N2113);
and AND2 (N3373, N3371, N3012);
or OR4 (N3374, N3357, N906, N937, N2794);
nor NOR4 (N3375, N3372, N1000, N2893, N2166);
or OR2 (N3376, N3373, N603);
nor NOR4 (N3377, N3360, N1454, N1912, N717);
or OR4 (N3378, N3365, N1881, N2036, N3265);
or OR4 (N3379, N3375, N2913, N1717, N1008);
nor NOR2 (N3380, N3368, N453);
nor NOR4 (N3381, N3370, N2918, N3113, N46);
or OR4 (N3382, N3376, N186, N2687, N2067);
nand NAND2 (N3383, N3378, N705);
xor XOR2 (N3384, N3380, N133);
nand NAND2 (N3385, N3383, N2029);
nor NOR2 (N3386, N3384, N2303);
not NOT1 (N3387, N3363);
or OR2 (N3388, N3327, N2200);
buf BUF1 (N3389, N3381);
xor XOR2 (N3390, N3388, N2194);
nand NAND4 (N3391, N3382, N881, N302, N1737);
nor NOR4 (N3392, N3391, N2321, N3370, N1611);
not NOT1 (N3393, N3386);
or OR2 (N3394, N3377, N2591);
buf BUF1 (N3395, N3374);
buf BUF1 (N3396, N3367);
nor NOR2 (N3397, N3396, N2916);
xor XOR2 (N3398, N3390, N260);
xor XOR2 (N3399, N3379, N2755);
and AND3 (N3400, N3393, N3045, N1522);
or OR3 (N3401, N3397, N2466, N2116);
buf BUF1 (N3402, N3395);
nand NAND3 (N3403, N3399, N1608, N3012);
not NOT1 (N3404, N3398);
nand NAND3 (N3405, N3403, N1898, N1860);
not NOT1 (N3406, N3402);
or OR3 (N3407, N3389, N2049, N183);
not NOT1 (N3408, N3407);
xor XOR2 (N3409, N3408, N3092);
xor XOR2 (N3410, N3401, N2365);
not NOT1 (N3411, N3387);
or OR4 (N3412, N3409, N630, N3284, N633);
or OR4 (N3413, N3404, N1036, N329, N3348);
nand NAND4 (N3414, N3411, N1013, N3319, N1873);
xor XOR2 (N3415, N3414, N2552);
nor NOR2 (N3416, N3392, N2242);
and AND3 (N3417, N3410, N2274, N2137);
buf BUF1 (N3418, N3416);
xor XOR2 (N3419, N3412, N1058);
not NOT1 (N3420, N3385);
xor XOR2 (N3421, N3417, N1526);
xor XOR2 (N3422, N3400, N3022);
or OR4 (N3423, N3418, N1863, N1399, N3217);
nand NAND4 (N3424, N3420, N2524, N1477, N3378);
nor NOR2 (N3425, N3394, N3071);
or OR2 (N3426, N3413, N1398);
xor XOR2 (N3427, N3421, N105);
xor XOR2 (N3428, N3422, N2699);
nor NOR2 (N3429, N3423, N871);
buf BUF1 (N3430, N3424);
xor XOR2 (N3431, N3405, N975);
and AND2 (N3432, N3415, N2011);
not NOT1 (N3433, N3432);
buf BUF1 (N3434, N3430);
or OR4 (N3435, N3434, N1092, N2957, N380);
and AND2 (N3436, N3429, N1794);
or OR2 (N3437, N3436, N365);
buf BUF1 (N3438, N3427);
buf BUF1 (N3439, N3435);
or OR3 (N3440, N3428, N3295, N2715);
nand NAND4 (N3441, N3425, N1233, N3242, N1381);
nand NAND3 (N3442, N3441, N2707, N3279);
nor NOR4 (N3443, N3440, N1304, N2507, N1261);
buf BUF1 (N3444, N3426);
not NOT1 (N3445, N3442);
buf BUF1 (N3446, N3438);
nand NAND2 (N3447, N3431, N3120);
buf BUF1 (N3448, N3419);
nor NOR3 (N3449, N3445, N874, N2250);
not NOT1 (N3450, N3437);
buf BUF1 (N3451, N3443);
not NOT1 (N3452, N3449);
or OR2 (N3453, N3447, N2752);
or OR3 (N3454, N3452, N1266, N3184);
xor XOR2 (N3455, N3406, N2064);
and AND4 (N3456, N3439, N2093, N149, N3351);
and AND3 (N3457, N3455, N79, N1336);
nor NOR4 (N3458, N3453, N3034, N170, N2267);
and AND3 (N3459, N3457, N88, N1552);
nor NOR2 (N3460, N3444, N2467);
buf BUF1 (N3461, N3433);
and AND4 (N3462, N3458, N2359, N2587, N109);
not NOT1 (N3463, N3460);
xor XOR2 (N3464, N3462, N596);
buf BUF1 (N3465, N3446);
xor XOR2 (N3466, N3454, N941);
and AND3 (N3467, N3451, N2666, N1429);
nor NOR2 (N3468, N3459, N1738);
not NOT1 (N3469, N3466);
buf BUF1 (N3470, N3467);
not NOT1 (N3471, N3468);
nand NAND3 (N3472, N3456, N2701, N2305);
nand NAND2 (N3473, N3472, N102);
not NOT1 (N3474, N3473);
not NOT1 (N3475, N3450);
nand NAND4 (N3476, N3461, N1988, N1794, N2363);
or OR2 (N3477, N3474, N948);
xor XOR2 (N3478, N3471, N2703);
not NOT1 (N3479, N3476);
nor NOR4 (N3480, N3470, N1522, N1512, N2321);
buf BUF1 (N3481, N3469);
not NOT1 (N3482, N3475);
xor XOR2 (N3483, N3464, N3118);
and AND3 (N3484, N3479, N1426, N2917);
nor NOR2 (N3485, N3463, N1302);
nor NOR2 (N3486, N3484, N2368);
nor NOR2 (N3487, N3482, N953);
buf BUF1 (N3488, N3465);
nor NOR2 (N3489, N3483, N209);
nor NOR4 (N3490, N3477, N3160, N1459, N2999);
buf BUF1 (N3491, N3489);
not NOT1 (N3492, N3481);
nor NOR4 (N3493, N3486, N1149, N930, N731);
or OR4 (N3494, N3491, N2678, N3024, N3023);
and AND3 (N3495, N3487, N1650, N72);
and AND2 (N3496, N3494, N1487);
nor NOR3 (N3497, N3493, N1309, N184);
nand NAND2 (N3498, N3497, N1100);
nor NOR2 (N3499, N3448, N1520);
xor XOR2 (N3500, N3490, N2368);
nor NOR3 (N3501, N3499, N559, N3458);
nand NAND3 (N3502, N3501, N1557, N1842);
not NOT1 (N3503, N3478);
nand NAND4 (N3504, N3480, N2991, N3001, N1177);
nand NAND2 (N3505, N3485, N1098);
nor NOR4 (N3506, N3492, N922, N1505, N2827);
buf BUF1 (N3507, N3505);
nand NAND3 (N3508, N3502, N1420, N2774);
nor NOR2 (N3509, N3508, N2948);
buf BUF1 (N3510, N3498);
xor XOR2 (N3511, N3503, N2930);
nand NAND2 (N3512, N3495, N2950);
and AND2 (N3513, N3506, N1418);
nor NOR2 (N3514, N3511, N1225);
nor NOR2 (N3515, N3504, N131);
not NOT1 (N3516, N3513);
or OR3 (N3517, N3510, N3161, N2018);
not NOT1 (N3518, N3516);
nand NAND2 (N3519, N3507, N591);
buf BUF1 (N3520, N3519);
not NOT1 (N3521, N3515);
or OR4 (N3522, N3520, N1614, N1438, N108);
buf BUF1 (N3523, N3509);
not NOT1 (N3524, N3517);
nor NOR3 (N3525, N3514, N25, N2133);
nand NAND2 (N3526, N3518, N1190);
nor NOR3 (N3527, N3526, N1183, N837);
xor XOR2 (N3528, N3512, N2187);
xor XOR2 (N3529, N3523, N3173);
nand NAND3 (N3530, N3529, N1503, N2789);
and AND3 (N3531, N3527, N2355, N834);
buf BUF1 (N3532, N3500);
buf BUF1 (N3533, N3522);
or OR2 (N3534, N3528, N1107);
xor XOR2 (N3535, N3524, N1513);
nand NAND3 (N3536, N3530, N1834, N2784);
buf BUF1 (N3537, N3525);
nor NOR4 (N3538, N3531, N684, N1981, N60);
xor XOR2 (N3539, N3521, N188);
xor XOR2 (N3540, N3537, N2895);
nor NOR2 (N3541, N3540, N2528);
nor NOR3 (N3542, N3539, N1305, N1023);
buf BUF1 (N3543, N3496);
buf BUF1 (N3544, N3534);
xor XOR2 (N3545, N3541, N655);
and AND4 (N3546, N3536, N1696, N1458, N2736);
and AND4 (N3547, N3533, N1566, N716, N3480);
nand NAND2 (N3548, N3547, N513);
buf BUF1 (N3549, N3535);
and AND2 (N3550, N3546, N3429);
buf BUF1 (N3551, N3548);
not NOT1 (N3552, N3543);
nor NOR4 (N3553, N3532, N2111, N2402, N3183);
nor NOR4 (N3554, N3552, N1935, N994, N310);
buf BUF1 (N3555, N3549);
and AND2 (N3556, N3553, N2680);
xor XOR2 (N3557, N3488, N3260);
nand NAND4 (N3558, N3550, N3087, N3128, N2662);
or OR2 (N3559, N3554, N2871);
xor XOR2 (N3560, N3559, N532);
buf BUF1 (N3561, N3544);
nor NOR4 (N3562, N3555, N1766, N627, N1423);
nor NOR4 (N3563, N3557, N1832, N870, N952);
nand NAND2 (N3564, N3556, N411);
not NOT1 (N3565, N3562);
nor NOR2 (N3566, N3561, N104);
not NOT1 (N3567, N3551);
or OR3 (N3568, N3545, N3517, N1542);
nor NOR3 (N3569, N3538, N2796, N1911);
or OR3 (N3570, N3567, N1166, N2318);
and AND4 (N3571, N3558, N2081, N1724, N2581);
buf BUF1 (N3572, N3570);
nor NOR3 (N3573, N3572, N1660, N2521);
buf BUF1 (N3574, N3568);
buf BUF1 (N3575, N3542);
xor XOR2 (N3576, N3564, N424);
nand NAND3 (N3577, N3565, N701, N2180);
nor NOR4 (N3578, N3566, N284, N3452, N2301);
nor NOR2 (N3579, N3575, N2750);
nor NOR3 (N3580, N3569, N1555, N1238);
buf BUF1 (N3581, N3577);
xor XOR2 (N3582, N3573, N1838);
not NOT1 (N3583, N3574);
and AND2 (N3584, N3578, N1592);
not NOT1 (N3585, N3582);
xor XOR2 (N3586, N3560, N2494);
not NOT1 (N3587, N3583);
or OR3 (N3588, N3580, N12, N2164);
or OR4 (N3589, N3571, N1113, N164, N2722);
not NOT1 (N3590, N3581);
nor NOR3 (N3591, N3563, N3238, N1004);
nor NOR4 (N3592, N3589, N449, N1973, N3378);
buf BUF1 (N3593, N3592);
not NOT1 (N3594, N3590);
or OR4 (N3595, N3579, N152, N1944, N1058);
xor XOR2 (N3596, N3591, N2052);
nand NAND2 (N3597, N3595, N2163);
or OR4 (N3598, N3594, N2141, N2396, N724);
not NOT1 (N3599, N3598);
or OR3 (N3600, N3596, N1018, N1148);
or OR4 (N3601, N3585, N2239, N225, N3152);
or OR3 (N3602, N3600, N1717, N1638);
xor XOR2 (N3603, N3597, N2049);
and AND4 (N3604, N3584, N1474, N658, N3599);
xor XOR2 (N3605, N1053, N3298);
not NOT1 (N3606, N3601);
or OR4 (N3607, N3586, N1964, N661, N16);
nand NAND3 (N3608, N3587, N1513, N1859);
and AND3 (N3609, N3593, N1653, N1181);
or OR2 (N3610, N3609, N1124);
nor NOR3 (N3611, N3602, N2380, N323);
buf BUF1 (N3612, N3607);
and AND3 (N3613, N3611, N1122, N2065);
xor XOR2 (N3614, N3588, N2440);
nand NAND3 (N3615, N3603, N720, N2577);
nor NOR2 (N3616, N3613, N2770);
and AND2 (N3617, N3614, N3509);
and AND3 (N3618, N3606, N2412, N1252);
nor NOR4 (N3619, N3612, N44, N3287, N31);
not NOT1 (N3620, N3615);
or OR4 (N3621, N3605, N1506, N2365, N1221);
not NOT1 (N3622, N3617);
nor NOR4 (N3623, N3619, N2547, N1343, N3267);
not NOT1 (N3624, N3610);
xor XOR2 (N3625, N3620, N3492);
and AND2 (N3626, N3576, N155);
buf BUF1 (N3627, N3604);
xor XOR2 (N3628, N3627, N3522);
xor XOR2 (N3629, N3618, N1312);
not NOT1 (N3630, N3621);
not NOT1 (N3631, N3608);
buf BUF1 (N3632, N3624);
or OR3 (N3633, N3626, N2361, N1106);
or OR2 (N3634, N3633, N3376);
nand NAND3 (N3635, N3632, N3030, N2864);
nor NOR4 (N3636, N3628, N677, N499, N1923);
xor XOR2 (N3637, N3629, N3619);
not NOT1 (N3638, N3616);
and AND3 (N3639, N3638, N1548, N2751);
nand NAND3 (N3640, N3631, N2289, N1615);
xor XOR2 (N3641, N3637, N104);
or OR4 (N3642, N3635, N2958, N1674, N1753);
xor XOR2 (N3643, N3641, N643);
xor XOR2 (N3644, N3639, N2653);
buf BUF1 (N3645, N3642);
xor XOR2 (N3646, N3623, N535);
buf BUF1 (N3647, N3634);
or OR2 (N3648, N3643, N3440);
and AND4 (N3649, N3645, N526, N496, N392);
buf BUF1 (N3650, N3625);
not NOT1 (N3651, N3650);
nor NOR3 (N3652, N3647, N1448, N2551);
or OR2 (N3653, N3640, N1648);
and AND3 (N3654, N3651, N2744, N3222);
nand NAND2 (N3655, N3653, N2046);
and AND4 (N3656, N3649, N2952, N2077, N909);
or OR2 (N3657, N3655, N260);
nand NAND2 (N3658, N3636, N1876);
not NOT1 (N3659, N3658);
and AND3 (N3660, N3652, N2168, N1590);
xor XOR2 (N3661, N3659, N1575);
nor NOR3 (N3662, N3654, N1319, N7);
xor XOR2 (N3663, N3656, N3196);
or OR4 (N3664, N3662, N1829, N188, N1029);
nor NOR4 (N3665, N3646, N1548, N474, N2181);
nand NAND2 (N3666, N3661, N734);
and AND2 (N3667, N3665, N1771);
not NOT1 (N3668, N3664);
xor XOR2 (N3669, N3660, N3434);
buf BUF1 (N3670, N3657);
buf BUF1 (N3671, N3644);
xor XOR2 (N3672, N3648, N3481);
not NOT1 (N3673, N3663);
and AND3 (N3674, N3670, N1073, N3443);
and AND3 (N3675, N3630, N2850, N1261);
nor NOR3 (N3676, N3671, N583, N882);
not NOT1 (N3677, N3666);
buf BUF1 (N3678, N3675);
nand NAND3 (N3679, N3674, N914, N1511);
not NOT1 (N3680, N3673);
xor XOR2 (N3681, N3668, N82);
xor XOR2 (N3682, N3672, N414);
nand NAND4 (N3683, N3679, N3543, N2395, N963);
xor XOR2 (N3684, N3622, N2642);
nand NAND4 (N3685, N3678, N1778, N1903, N3127);
or OR2 (N3686, N3676, N522);
buf BUF1 (N3687, N3685);
and AND3 (N3688, N3669, N612, N3323);
buf BUF1 (N3689, N3680);
buf BUF1 (N3690, N3681);
or OR4 (N3691, N3686, N1984, N1014, N3666);
or OR3 (N3692, N3688, N1513, N2236);
nand NAND2 (N3693, N3667, N1580);
not NOT1 (N3694, N3691);
nor NOR4 (N3695, N3692, N3042, N1643, N316);
not NOT1 (N3696, N3684);
buf BUF1 (N3697, N3689);
nor NOR4 (N3698, N3687, N1528, N3106, N759);
and AND2 (N3699, N3690, N880);
and AND3 (N3700, N3683, N161, N2454);
not NOT1 (N3701, N3700);
nor NOR4 (N3702, N3695, N2056, N2996, N779);
buf BUF1 (N3703, N3698);
nor NOR3 (N3704, N3696, N1161, N157);
or OR4 (N3705, N3702, N2650, N3296, N728);
or OR2 (N3706, N3705, N2638);
nor NOR2 (N3707, N3706, N3064);
buf BUF1 (N3708, N3682);
not NOT1 (N3709, N3707);
not NOT1 (N3710, N3701);
or OR2 (N3711, N3697, N2512);
or OR4 (N3712, N3708, N2706, N1014, N1931);
and AND3 (N3713, N3703, N3495, N2342);
nand NAND2 (N3714, N3677, N703);
nand NAND2 (N3715, N3709, N990);
not NOT1 (N3716, N3711);
or OR2 (N3717, N3713, N2844);
nor NOR3 (N3718, N3712, N88, N3662);
buf BUF1 (N3719, N3704);
nor NOR4 (N3720, N3693, N2750, N1040, N3532);
not NOT1 (N3721, N3719);
nor NOR4 (N3722, N3721, N927, N3512, N2321);
nor NOR4 (N3723, N3714, N1647, N3631, N1213);
nor NOR2 (N3724, N3722, N3688);
buf BUF1 (N3725, N3723);
nor NOR3 (N3726, N3715, N2016, N156);
xor XOR2 (N3727, N3718, N276);
nand NAND2 (N3728, N3727, N1558);
nand NAND4 (N3729, N3726, N2380, N2798, N166);
nand NAND2 (N3730, N3694, N3186);
xor XOR2 (N3731, N3717, N1106);
buf BUF1 (N3732, N3730);
buf BUF1 (N3733, N3724);
and AND4 (N3734, N3725, N809, N2703, N3568);
and AND2 (N3735, N3734, N484);
not NOT1 (N3736, N3699);
or OR4 (N3737, N3732, N2030, N3246, N1014);
xor XOR2 (N3738, N3728, N3290);
or OR3 (N3739, N3737, N2966, N3625);
nor NOR4 (N3740, N3720, N2419, N2567, N1946);
xor XOR2 (N3741, N3735, N503);
and AND4 (N3742, N3710, N1301, N2191, N1453);
or OR2 (N3743, N3739, N1353);
not NOT1 (N3744, N3741);
xor XOR2 (N3745, N3740, N431);
nand NAND2 (N3746, N3745, N2647);
or OR2 (N3747, N3731, N531);
not NOT1 (N3748, N3738);
and AND4 (N3749, N3733, N2129, N2149, N243);
nand NAND3 (N3750, N3748, N2084, N2723);
xor XOR2 (N3751, N3746, N3701);
nand NAND4 (N3752, N3729, N1175, N1906, N3589);
not NOT1 (N3753, N3749);
not NOT1 (N3754, N3747);
not NOT1 (N3755, N3753);
not NOT1 (N3756, N3743);
nor NOR3 (N3757, N3736, N3625, N805);
nor NOR3 (N3758, N3757, N1469, N361);
xor XOR2 (N3759, N3755, N86);
nor NOR4 (N3760, N3752, N1, N3589, N272);
not NOT1 (N3761, N3751);
nand NAND3 (N3762, N3759, N113, N499);
not NOT1 (N3763, N3758);
nor NOR4 (N3764, N3744, N2375, N1431, N3130);
nor NOR3 (N3765, N3742, N475, N3361);
and AND2 (N3766, N3764, N1443);
buf BUF1 (N3767, N3754);
xor XOR2 (N3768, N3750, N3137);
buf BUF1 (N3769, N3766);
not NOT1 (N3770, N3762);
and AND4 (N3771, N3760, N3020, N1413, N3435);
and AND2 (N3772, N3767, N801);
buf BUF1 (N3773, N3765);
nand NAND3 (N3774, N3763, N505, N817);
buf BUF1 (N3775, N3756);
buf BUF1 (N3776, N3770);
and AND4 (N3777, N3775, N3096, N2514, N2963);
and AND3 (N3778, N3777, N2183, N3649);
nand NAND3 (N3779, N3778, N3280, N24);
not NOT1 (N3780, N3774);
not NOT1 (N3781, N3769);
nor NOR3 (N3782, N3771, N2735, N1016);
nand NAND4 (N3783, N3780, N1299, N1028, N2311);
and AND4 (N3784, N3776, N1898, N1390, N2280);
xor XOR2 (N3785, N3783, N1811);
nor NOR3 (N3786, N3782, N484, N2192);
nand NAND2 (N3787, N3716, N3060);
buf BUF1 (N3788, N3772);
and AND2 (N3789, N3784, N711);
or OR3 (N3790, N3785, N1681, N1346);
not NOT1 (N3791, N3781);
xor XOR2 (N3792, N3761, N1861);
xor XOR2 (N3793, N3789, N1801);
nand NAND4 (N3794, N3792, N751, N2563, N6);
nor NOR2 (N3795, N3773, N1809);
and AND4 (N3796, N3794, N1290, N2741, N425);
xor XOR2 (N3797, N3795, N1411);
or OR4 (N3798, N3790, N1791, N1630, N2043);
nor NOR4 (N3799, N3793, N2318, N1636, N672);
and AND3 (N3800, N3796, N390, N1204);
and AND2 (N3801, N3799, N1724);
xor XOR2 (N3802, N3786, N1815);
or OR2 (N3803, N3797, N523);
or OR2 (N3804, N3779, N3424);
nand NAND4 (N3805, N3791, N3246, N987, N428);
xor XOR2 (N3806, N3787, N1083);
and AND4 (N3807, N3800, N2479, N1317, N3101);
buf BUF1 (N3808, N3768);
buf BUF1 (N3809, N3788);
buf BUF1 (N3810, N3809);
nor NOR4 (N3811, N3803, N1825, N2740, N2993);
nand NAND2 (N3812, N3804, N3171);
or OR4 (N3813, N3812, N3794, N2818, N175);
buf BUF1 (N3814, N3798);
and AND4 (N3815, N3805, N664, N1124, N2191);
not NOT1 (N3816, N3802);
nand NAND2 (N3817, N3813, N203);
and AND3 (N3818, N3801, N1106, N420);
nand NAND2 (N3819, N3817, N830);
and AND3 (N3820, N3807, N1143, N2985);
and AND4 (N3821, N3814, N1717, N1008, N3594);
buf BUF1 (N3822, N3821);
nand NAND2 (N3823, N3808, N3455);
not NOT1 (N3824, N3819);
xor XOR2 (N3825, N3810, N2547);
not NOT1 (N3826, N3806);
buf BUF1 (N3827, N3820);
buf BUF1 (N3828, N3823);
nand NAND4 (N3829, N3825, N3329, N1979, N3137);
nor NOR4 (N3830, N3827, N960, N2909, N312);
buf BUF1 (N3831, N3818);
buf BUF1 (N3832, N3826);
and AND2 (N3833, N3822, N2131);
and AND4 (N3834, N3811, N2562, N694, N3307);
buf BUF1 (N3835, N3834);
and AND2 (N3836, N3816, N517);
and AND4 (N3837, N3828, N228, N7, N559);
or OR3 (N3838, N3835, N2555, N152);
nor NOR3 (N3839, N3838, N2345, N1468);
nand NAND3 (N3840, N3837, N643, N3730);
and AND2 (N3841, N3832, N2181);
and AND2 (N3842, N3836, N2588);
nand NAND4 (N3843, N3840, N961, N1413, N1554);
or OR4 (N3844, N3841, N14, N2163, N654);
buf BUF1 (N3845, N3842);
nand NAND3 (N3846, N3815, N1349, N3208);
nor NOR4 (N3847, N3844, N2285, N1982, N1074);
nor NOR4 (N3848, N3847, N996, N321, N3111);
nand NAND3 (N3849, N3839, N2831, N518);
xor XOR2 (N3850, N3833, N500);
nand NAND3 (N3851, N3850, N1653, N699);
and AND4 (N3852, N3846, N1900, N399, N3304);
nor NOR3 (N3853, N3830, N720, N2553);
and AND4 (N3854, N3845, N1203, N1505, N3363);
or OR3 (N3855, N3852, N2630, N1790);
not NOT1 (N3856, N3851);
and AND3 (N3857, N3829, N2028, N209);
not NOT1 (N3858, N3854);
buf BUF1 (N3859, N3849);
xor XOR2 (N3860, N3843, N1542);
xor XOR2 (N3861, N3859, N2192);
nor NOR2 (N3862, N3848, N2267);
or OR2 (N3863, N3857, N2995);
nand NAND4 (N3864, N3861, N977, N2714, N3250);
buf BUF1 (N3865, N3853);
and AND2 (N3866, N3860, N316);
buf BUF1 (N3867, N3865);
buf BUF1 (N3868, N3831);
nor NOR4 (N3869, N3866, N1957, N213, N2150);
and AND2 (N3870, N3867, N1796);
nand NAND3 (N3871, N3824, N3509, N425);
buf BUF1 (N3872, N3863);
nand NAND4 (N3873, N3871, N2271, N3047, N1330);
or OR3 (N3874, N3864, N1764, N525);
nand NAND4 (N3875, N3862, N2859, N3282, N1701);
not NOT1 (N3876, N3872);
nor NOR4 (N3877, N3856, N3874, N849, N141);
and AND2 (N3878, N466, N921);
xor XOR2 (N3879, N3855, N3570);
buf BUF1 (N3880, N3868);
and AND4 (N3881, N3858, N2715, N3487, N1267);
xor XOR2 (N3882, N3875, N3799);
and AND4 (N3883, N3880, N934, N76, N1699);
buf BUF1 (N3884, N3879);
xor XOR2 (N3885, N3876, N25);
and AND4 (N3886, N3878, N2220, N3256, N235);
not NOT1 (N3887, N3873);
and AND3 (N3888, N3881, N2002, N3484);
nor NOR4 (N3889, N3882, N228, N2493, N1320);
nor NOR3 (N3890, N3888, N1494, N2983);
or OR4 (N3891, N3885, N524, N1823, N602);
buf BUF1 (N3892, N3890);
not NOT1 (N3893, N3886);
xor XOR2 (N3894, N3884, N1523);
nand NAND2 (N3895, N3889, N2473);
buf BUF1 (N3896, N3870);
or OR3 (N3897, N3883, N3811, N516);
and AND2 (N3898, N3869, N2085);
nor NOR4 (N3899, N3897, N641, N3508, N3035);
nand NAND2 (N3900, N3877, N2861);
not NOT1 (N3901, N3887);
buf BUF1 (N3902, N3896);
nor NOR4 (N3903, N3902, N2967, N1024, N2292);
or OR4 (N3904, N3895, N1982, N1180, N849);
buf BUF1 (N3905, N3894);
nand NAND3 (N3906, N3891, N1429, N2338);
and AND4 (N3907, N3900, N3227, N1627, N3522);
not NOT1 (N3908, N3905);
or OR3 (N3909, N3907, N2826, N793);
nor NOR4 (N3910, N3892, N3471, N305, N1462);
nor NOR2 (N3911, N3908, N3892);
nand NAND3 (N3912, N3910, N946, N1856);
buf BUF1 (N3913, N3898);
nor NOR3 (N3914, N3893, N1894, N14);
or OR3 (N3915, N3913, N1219, N1003);
not NOT1 (N3916, N3903);
nand NAND2 (N3917, N3899, N3073);
not NOT1 (N3918, N3904);
and AND2 (N3919, N3915, N2129);
nor NOR4 (N3920, N3918, N1099, N2875, N963);
nor NOR2 (N3921, N3919, N313);
or OR2 (N3922, N3917, N3165);
xor XOR2 (N3923, N3922, N2072);
buf BUF1 (N3924, N3916);
buf BUF1 (N3925, N3906);
nor NOR2 (N3926, N3911, N1657);
nor NOR2 (N3927, N3901, N2277);
buf BUF1 (N3928, N3921);
xor XOR2 (N3929, N3920, N1481);
and AND3 (N3930, N3926, N2523, N906);
xor XOR2 (N3931, N3909, N3784);
or OR2 (N3932, N3928, N2557);
or OR2 (N3933, N3925, N1193);
or OR2 (N3934, N3931, N1805);
not NOT1 (N3935, N3932);
buf BUF1 (N3936, N3933);
xor XOR2 (N3937, N3924, N2968);
nor NOR3 (N3938, N3930, N3842, N1811);
xor XOR2 (N3939, N3936, N723);
or OR2 (N3940, N3938, N2872);
nand NAND4 (N3941, N3940, N929, N3360, N863);
not NOT1 (N3942, N3927);
nand NAND3 (N3943, N3935, N220, N585);
or OR4 (N3944, N3929, N2217, N3216, N165);
buf BUF1 (N3945, N3937);
nand NAND4 (N3946, N3941, N832, N1391, N2044);
or OR4 (N3947, N3923, N2785, N2455, N195);
and AND2 (N3948, N3946, N3137);
buf BUF1 (N3949, N3945);
or OR2 (N3950, N3944, N2517);
nor NOR4 (N3951, N3914, N2972, N831, N3106);
or OR4 (N3952, N3950, N2463, N1140, N551);
nand NAND3 (N3953, N3912, N345, N3814);
nand NAND3 (N3954, N3934, N644, N3556);
and AND2 (N3955, N3952, N3584);
not NOT1 (N3956, N3947);
nand NAND2 (N3957, N3943, N3181);
xor XOR2 (N3958, N3951, N3525);
not NOT1 (N3959, N3948);
buf BUF1 (N3960, N3957);
xor XOR2 (N3961, N3956, N1833);
not NOT1 (N3962, N3955);
nand NAND3 (N3963, N3939, N959, N1772);
nand NAND2 (N3964, N3942, N769);
nand NAND2 (N3965, N3953, N1941);
nor NOR2 (N3966, N3964, N3126);
or OR4 (N3967, N3959, N2736, N1779, N1916);
nor NOR4 (N3968, N3963, N3673, N1008, N137);
or OR3 (N3969, N3966, N27, N1113);
or OR4 (N3970, N3958, N252, N1952, N1483);
not NOT1 (N3971, N3960);
and AND2 (N3972, N3967, N3675);
xor XOR2 (N3973, N3961, N3606);
nand NAND3 (N3974, N3971, N293, N3350);
or OR3 (N3975, N3949, N1719, N2440);
nand NAND3 (N3976, N3974, N2964, N3784);
xor XOR2 (N3977, N3972, N1981);
and AND3 (N3978, N3977, N3487, N2854);
not NOT1 (N3979, N3970);
and AND3 (N3980, N3975, N2929, N1012);
or OR4 (N3981, N3973, N2344, N3173, N1540);
and AND2 (N3982, N3954, N1879);
buf BUF1 (N3983, N3978);
nand NAND2 (N3984, N3976, N1532);
nand NAND3 (N3985, N3968, N1291, N616);
not NOT1 (N3986, N3980);
nor NOR3 (N3987, N3962, N3377, N3663);
not NOT1 (N3988, N3984);
buf BUF1 (N3989, N3979);
and AND3 (N3990, N3988, N2555, N1865);
not NOT1 (N3991, N3982);
and AND2 (N3992, N3990, N1827);
or OR2 (N3993, N3991, N3778);
nor NOR3 (N3994, N3992, N3683, N2743);
or OR2 (N3995, N3983, N131);
nand NAND3 (N3996, N3969, N1890, N613);
not NOT1 (N3997, N3987);
nand NAND4 (N3998, N3985, N1564, N3804, N2641);
nand NAND4 (N3999, N3996, N828, N2055, N3046);
nor NOR2 (N4000, N3981, N3437);
and AND2 (N4001, N3995, N1664);
xor XOR2 (N4002, N4001, N780);
not NOT1 (N4003, N4002);
xor XOR2 (N4004, N3965, N2131);
xor XOR2 (N4005, N4003, N2150);
and AND3 (N4006, N3998, N278, N3793);
not NOT1 (N4007, N3986);
buf BUF1 (N4008, N3993);
nor NOR4 (N4009, N3989, N207, N1418, N2753);
nor NOR2 (N4010, N4005, N2898);
buf BUF1 (N4011, N4008);
nor NOR3 (N4012, N3999, N1380, N2629);
not NOT1 (N4013, N4010);
nor NOR3 (N4014, N4012, N3893, N3178);
buf BUF1 (N4015, N4004);
nand NAND4 (N4016, N4006, N1776, N815, N89);
and AND2 (N4017, N4013, N1192);
or OR4 (N4018, N4017, N542, N1182, N3216);
or OR3 (N4019, N3994, N2212, N2499);
endmodule