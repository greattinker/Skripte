// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16;

output N25602,N25613,N25610,N25589,N25615,N25612,N25607,N25614,N25611,N25616;

not NOT1 (N17, N8);
nand NAND3 (N18, N10, N12, N12);
xor XOR2 (N19, N14, N8);
and AND2 (N20, N8, N18);
or OR3 (N21, N20, N14, N4);
and AND2 (N22, N1, N7);
not NOT1 (N23, N4);
nand NAND2 (N24, N5, N23);
nor NOR4 (N25, N21, N20, N21, N21);
nor NOR3 (N26, N22, N5, N22);
not NOT1 (N27, N14);
buf BUF1 (N28, N9);
and AND3 (N29, N20, N5, N2);
or OR4 (N30, N3, N29, N6, N6);
and AND2 (N31, N14, N11);
or OR3 (N32, N9, N11, N19);
buf BUF1 (N33, N17);
or OR4 (N34, N18, N5, N6, N28);
not NOT1 (N35, N25);
and AND2 (N36, N30, N11);
or OR2 (N37, N36, N19);
or OR2 (N38, N6, N12);
and AND3 (N39, N26, N21, N11);
and AND2 (N40, N39, N32);
nand NAND4 (N41, N18, N25, N29, N22);
not NOT1 (N42, N31);
nand NAND2 (N43, N33, N19);
and AND2 (N44, N38, N10);
nand NAND4 (N45, N35, N23, N40, N43);
not NOT1 (N46, N35);
xor XOR2 (N47, N4, N8);
nand NAND4 (N48, N37, N3, N33, N18);
not NOT1 (N49, N27);
xor XOR2 (N50, N45, N29);
and AND2 (N51, N50, N42);
nand NAND3 (N52, N45, N41, N38);
and AND2 (N53, N9, N43);
and AND2 (N54, N44, N43);
and AND3 (N55, N47, N1, N22);
xor XOR2 (N56, N34, N20);
and AND4 (N57, N46, N35, N28, N46);
buf BUF1 (N58, N51);
nor NOR3 (N59, N58, N11, N20);
or OR3 (N60, N54, N32, N32);
or OR3 (N61, N56, N39, N31);
buf BUF1 (N62, N55);
buf BUF1 (N63, N49);
buf BUF1 (N64, N53);
nand NAND4 (N65, N59, N18, N16, N64);
nor NOR3 (N66, N13, N8, N41);
not NOT1 (N67, N61);
nand NAND2 (N68, N65, N43);
xor XOR2 (N69, N48, N4);
and AND2 (N70, N60, N10);
and AND4 (N71, N66, N66, N7, N69);
and AND3 (N72, N60, N63, N49);
xor XOR2 (N73, N7, N65);
nor NOR3 (N74, N73, N56, N22);
xor XOR2 (N75, N74, N49);
nand NAND2 (N76, N52, N33);
nor NOR3 (N77, N68, N40, N16);
nor NOR2 (N78, N57, N50);
xor XOR2 (N79, N76, N15);
or OR3 (N80, N70, N17, N33);
not NOT1 (N81, N79);
and AND3 (N82, N62, N74, N75);
or OR3 (N83, N29, N78, N16);
nor NOR3 (N84, N52, N64, N54);
buf BUF1 (N85, N84);
not NOT1 (N86, N71);
nand NAND3 (N87, N80, N64, N3);
not NOT1 (N88, N85);
xor XOR2 (N89, N88, N24);
buf BUF1 (N90, N86);
xor XOR2 (N91, N56, N42);
nor NOR2 (N92, N83, N30);
not NOT1 (N93, N81);
buf BUF1 (N94, N92);
nor NOR4 (N95, N94, N25, N7, N86);
not NOT1 (N96, N87);
nand NAND4 (N97, N91, N1, N69, N85);
and AND2 (N98, N93, N77);
nand NAND2 (N99, N77, N59);
nor NOR3 (N100, N90, N59, N82);
xor XOR2 (N101, N10, N19);
and AND4 (N102, N67, N7, N99, N76);
not NOT1 (N103, N8);
nand NAND2 (N104, N96, N3);
buf BUF1 (N105, N103);
nand NAND4 (N106, N101, N66, N50, N56);
not NOT1 (N107, N104);
and AND3 (N108, N106, N81, N42);
nand NAND4 (N109, N105, N17, N23, N106);
or OR4 (N110, N98, N66, N99, N35);
xor XOR2 (N111, N102, N64);
and AND4 (N112, N108, N27, N75, N8);
buf BUF1 (N113, N110);
xor XOR2 (N114, N72, N109);
and AND4 (N115, N75, N25, N18, N4);
nand NAND3 (N116, N114, N52, N15);
nor NOR3 (N117, N113, N3, N40);
xor XOR2 (N118, N97, N7);
or OR4 (N119, N117, N117, N9, N64);
nor NOR3 (N120, N107, N9, N15);
and AND4 (N121, N95, N88, N120, N52);
buf BUF1 (N122, N112);
buf BUF1 (N123, N97);
not NOT1 (N124, N118);
buf BUF1 (N125, N119);
nor NOR4 (N126, N116, N82, N107, N18);
or OR2 (N127, N122, N39);
or OR3 (N128, N115, N96, N49);
or OR2 (N129, N111, N17);
and AND4 (N130, N125, N66, N83, N82);
and AND4 (N131, N130, N70, N17, N94);
nor NOR2 (N132, N123, N124);
or OR4 (N133, N8, N10, N38, N76);
or OR4 (N134, N129, N78, N22, N85);
not NOT1 (N135, N121);
nor NOR2 (N136, N127, N128);
xor XOR2 (N137, N136, N91);
not NOT1 (N138, N69);
nand NAND2 (N139, N131, N57);
buf BUF1 (N140, N100);
nor NOR2 (N141, N133, N51);
and AND2 (N142, N135, N103);
nand NAND2 (N143, N139, N85);
nand NAND2 (N144, N143, N88);
nand NAND4 (N145, N138, N114, N138, N69);
xor XOR2 (N146, N132, N95);
nand NAND4 (N147, N89, N100, N65, N60);
or OR2 (N148, N147, N20);
and AND4 (N149, N140, N23, N77, N22);
xor XOR2 (N150, N148, N109);
nor NOR3 (N151, N144, N142, N4);
buf BUF1 (N152, N125);
nor NOR4 (N153, N149, N144, N103, N66);
xor XOR2 (N154, N137, N2);
buf BUF1 (N155, N153);
nor NOR2 (N156, N151, N27);
xor XOR2 (N157, N145, N150);
xor XOR2 (N158, N1, N48);
xor XOR2 (N159, N158, N155);
or OR3 (N160, N49, N123, N13);
and AND4 (N161, N156, N32, N61, N134);
xor XOR2 (N162, N116, N117);
or OR4 (N163, N141, N24, N120, N159);
nand NAND4 (N164, N38, N12, N10, N110);
nor NOR4 (N165, N126, N75, N39, N58);
not NOT1 (N166, N160);
or OR3 (N167, N146, N166, N67);
or OR3 (N168, N23, N140, N123);
or OR2 (N169, N165, N5);
xor XOR2 (N170, N163, N73);
xor XOR2 (N171, N157, N48);
xor XOR2 (N172, N162, N7);
not NOT1 (N173, N161);
nand NAND3 (N174, N172, N82, N72);
buf BUF1 (N175, N167);
and AND2 (N176, N164, N103);
nor NOR4 (N177, N173, N133, N14, N24);
nand NAND2 (N178, N171, N7);
not NOT1 (N179, N174);
and AND2 (N180, N152, N76);
nor NOR4 (N181, N177, N56, N95, N23);
and AND2 (N182, N175, N68);
not NOT1 (N183, N178);
buf BUF1 (N184, N176);
buf BUF1 (N185, N180);
xor XOR2 (N186, N179, N112);
or OR3 (N187, N154, N92, N72);
not NOT1 (N188, N182);
and AND3 (N189, N168, N57, N51);
not NOT1 (N190, N185);
xor XOR2 (N191, N184, N170);
nor NOR2 (N192, N173, N32);
not NOT1 (N193, N191);
xor XOR2 (N194, N181, N187);
nor NOR2 (N195, N192, N192);
or OR2 (N196, N34, N87);
nor NOR2 (N197, N189, N137);
and AND2 (N198, N186, N169);
and AND3 (N199, N101, N136, N89);
not NOT1 (N200, N190);
or OR4 (N201, N194, N33, N39, N110);
nand NAND2 (N202, N201, N192);
nor NOR4 (N203, N196, N113, N165, N72);
nand NAND3 (N204, N195, N124, N199);
buf BUF1 (N205, N10);
nor NOR3 (N206, N197, N170, N92);
nand NAND2 (N207, N183, N133);
xor XOR2 (N208, N204, N27);
not NOT1 (N209, N202);
nand NAND4 (N210, N193, N30, N143, N169);
buf BUF1 (N211, N209);
nand NAND4 (N212, N206, N101, N80, N183);
and AND2 (N213, N203, N126);
buf BUF1 (N214, N207);
and AND3 (N215, N200, N133, N187);
buf BUF1 (N216, N211);
and AND4 (N217, N210, N168, N62, N137);
xor XOR2 (N218, N214, N190);
nand NAND3 (N219, N208, N152, N5);
nor NOR3 (N220, N188, N133, N128);
nor NOR2 (N221, N205, N131);
buf BUF1 (N222, N220);
xor XOR2 (N223, N215, N96);
nand NAND3 (N224, N219, N75, N177);
and AND2 (N225, N224, N164);
nor NOR3 (N226, N218, N194, N70);
nand NAND2 (N227, N223, N137);
buf BUF1 (N228, N226);
not NOT1 (N229, N216);
buf BUF1 (N230, N217);
not NOT1 (N231, N230);
nand NAND2 (N232, N222, N84);
buf BUF1 (N233, N232);
or OR3 (N234, N221, N75, N17);
buf BUF1 (N235, N234);
or OR2 (N236, N213, N77);
not NOT1 (N237, N212);
xor XOR2 (N238, N229, N174);
xor XOR2 (N239, N228, N220);
nand NAND2 (N240, N236, N125);
nor NOR3 (N241, N235, N8, N186);
nand NAND4 (N242, N198, N239, N21, N58);
nor NOR3 (N243, N99, N118, N234);
xor XOR2 (N244, N233, N58);
buf BUF1 (N245, N240);
or OR2 (N246, N238, N232);
xor XOR2 (N247, N225, N169);
or OR3 (N248, N227, N11, N3);
buf BUF1 (N249, N242);
or OR3 (N250, N243, N129, N69);
or OR2 (N251, N248, N171);
or OR3 (N252, N237, N43, N209);
and AND4 (N253, N252, N247, N216, N12);
nor NOR4 (N254, N149, N42, N4, N83);
nor NOR3 (N255, N246, N200, N79);
buf BUF1 (N256, N255);
buf BUF1 (N257, N250);
or OR3 (N258, N249, N97, N178);
buf BUF1 (N259, N244);
not NOT1 (N260, N259);
nand NAND3 (N261, N253, N124, N248);
not NOT1 (N262, N258);
buf BUF1 (N263, N254);
or OR2 (N264, N263, N238);
or OR2 (N265, N260, N145);
xor XOR2 (N266, N245, N208);
and AND4 (N267, N266, N85, N165, N197);
and AND4 (N268, N267, N161, N184, N106);
and AND4 (N269, N261, N27, N7, N82);
xor XOR2 (N270, N264, N62);
xor XOR2 (N271, N270, N226);
buf BUF1 (N272, N265);
xor XOR2 (N273, N271, N80);
and AND4 (N274, N269, N248, N262, N13);
or OR3 (N275, N25, N158, N264);
xor XOR2 (N276, N256, N36);
or OR2 (N277, N241, N31);
nor NOR4 (N278, N277, N113, N234, N212);
and AND3 (N279, N274, N179, N40);
xor XOR2 (N280, N231, N212);
not NOT1 (N281, N257);
buf BUF1 (N282, N278);
buf BUF1 (N283, N280);
not NOT1 (N284, N251);
nor NOR2 (N285, N281, N163);
nand NAND2 (N286, N279, N262);
not NOT1 (N287, N285);
or OR2 (N288, N282, N77);
xor XOR2 (N289, N275, N109);
xor XOR2 (N290, N286, N162);
and AND3 (N291, N273, N106, N102);
not NOT1 (N292, N287);
nand NAND2 (N293, N272, N212);
or OR2 (N294, N276, N134);
buf BUF1 (N295, N288);
nand NAND3 (N296, N284, N98, N37);
buf BUF1 (N297, N283);
nand NAND4 (N298, N292, N219, N31, N128);
and AND3 (N299, N295, N12, N169);
xor XOR2 (N300, N296, N67);
or OR2 (N301, N268, N156);
not NOT1 (N302, N300);
not NOT1 (N303, N302);
not NOT1 (N304, N303);
nor NOR3 (N305, N297, N75, N148);
not NOT1 (N306, N304);
or OR3 (N307, N298, N192, N102);
nand NAND3 (N308, N306, N31, N12);
not NOT1 (N309, N293);
not NOT1 (N310, N301);
or OR4 (N311, N294, N139, N33, N305);
nor NOR3 (N312, N110, N205, N120);
xor XOR2 (N313, N311, N241);
buf BUF1 (N314, N309);
nand NAND4 (N315, N313, N299, N143, N159);
nand NAND2 (N316, N6, N245);
nand NAND4 (N317, N290, N285, N32, N256);
nor NOR4 (N318, N316, N171, N267, N149);
xor XOR2 (N319, N317, N259);
not NOT1 (N320, N310);
nor NOR2 (N321, N312, N34);
or OR4 (N322, N307, N85, N75, N260);
and AND3 (N323, N291, N253, N255);
not NOT1 (N324, N319);
nand NAND2 (N325, N315, N174);
or OR4 (N326, N320, N292, N221, N274);
not NOT1 (N327, N308);
xor XOR2 (N328, N289, N303);
nor NOR2 (N329, N321, N237);
nor NOR3 (N330, N323, N75, N67);
and AND2 (N331, N322, N43);
not NOT1 (N332, N318);
or OR3 (N333, N325, N303, N228);
nor NOR3 (N334, N324, N216, N25);
not NOT1 (N335, N329);
nand NAND4 (N336, N330, N17, N204, N89);
nor NOR3 (N337, N326, N37, N56);
and AND3 (N338, N334, N327, N48);
or OR4 (N339, N273, N10, N283, N219);
or OR2 (N340, N314, N117);
or OR2 (N341, N332, N182);
not NOT1 (N342, N338);
or OR4 (N343, N337, N58, N36, N337);
and AND4 (N344, N342, N245, N201, N115);
and AND3 (N345, N331, N103, N159);
xor XOR2 (N346, N341, N210);
nand NAND3 (N347, N344, N230, N117);
buf BUF1 (N348, N347);
or OR3 (N349, N336, N197, N314);
or OR2 (N350, N333, N283);
not NOT1 (N351, N346);
nand NAND4 (N352, N328, N313, N50, N123);
nand NAND4 (N353, N351, N159, N8, N272);
buf BUF1 (N354, N340);
nand NAND3 (N355, N350, N185, N339);
and AND2 (N356, N175, N75);
nand NAND4 (N357, N355, N108, N293, N46);
not NOT1 (N358, N335);
xor XOR2 (N359, N352, N257);
not NOT1 (N360, N345);
or OR4 (N361, N354, N230, N312, N240);
and AND3 (N362, N343, N121, N313);
xor XOR2 (N363, N359, N335);
not NOT1 (N364, N360);
or OR2 (N365, N362, N97);
not NOT1 (N366, N361);
nand NAND4 (N367, N357, N311, N135, N323);
not NOT1 (N368, N353);
nor NOR3 (N369, N368, N67, N166);
or OR3 (N370, N358, N302, N43);
nand NAND2 (N371, N366, N237);
nor NOR2 (N372, N364, N161);
buf BUF1 (N373, N371);
nand NAND3 (N374, N372, N6, N259);
not NOT1 (N375, N367);
nor NOR3 (N376, N363, N111, N297);
xor XOR2 (N377, N365, N292);
nand NAND4 (N378, N376, N346, N323, N234);
buf BUF1 (N379, N356);
nand NAND2 (N380, N379, N80);
xor XOR2 (N381, N349, N22);
xor XOR2 (N382, N377, N346);
not NOT1 (N383, N380);
or OR4 (N384, N375, N339, N186, N74);
buf BUF1 (N385, N370);
nor NOR4 (N386, N381, N140, N24, N209);
not NOT1 (N387, N384);
or OR4 (N388, N374, N265, N211, N305);
buf BUF1 (N389, N373);
nand NAND3 (N390, N383, N111, N231);
xor XOR2 (N391, N378, N302);
or OR2 (N392, N386, N305);
and AND4 (N393, N348, N265, N352, N101);
and AND4 (N394, N392, N98, N84, N138);
or OR2 (N395, N387, N303);
not NOT1 (N396, N390);
or OR2 (N397, N388, N367);
or OR2 (N398, N397, N149);
xor XOR2 (N399, N382, N74);
or OR4 (N400, N393, N139, N362, N349);
nor NOR4 (N401, N389, N60, N353, N149);
and AND2 (N402, N369, N148);
not NOT1 (N403, N385);
xor XOR2 (N404, N403, N322);
nor NOR2 (N405, N394, N209);
and AND2 (N406, N404, N17);
buf BUF1 (N407, N400);
xor XOR2 (N408, N396, N190);
buf BUF1 (N409, N398);
or OR3 (N410, N407, N266, N336);
xor XOR2 (N411, N401, N289);
buf BUF1 (N412, N411);
or OR2 (N413, N391, N76);
buf BUF1 (N414, N406);
not NOT1 (N415, N408);
nor NOR3 (N416, N412, N214, N184);
not NOT1 (N417, N410);
or OR3 (N418, N414, N224, N10);
nand NAND3 (N419, N416, N268, N46);
xor XOR2 (N420, N402, N63);
not NOT1 (N421, N420);
nor NOR4 (N422, N418, N199, N286, N171);
buf BUF1 (N423, N405);
not NOT1 (N424, N419);
and AND3 (N425, N417, N343, N28);
xor XOR2 (N426, N395, N394);
and AND2 (N427, N424, N333);
nand NAND3 (N428, N409, N240, N189);
buf BUF1 (N429, N415);
nand NAND4 (N430, N425, N375, N115, N424);
or OR2 (N431, N430, N201);
not NOT1 (N432, N429);
and AND3 (N433, N426, N79, N392);
nand NAND2 (N434, N422, N159);
nor NOR2 (N435, N399, N208);
nand NAND3 (N436, N432, N293, N205);
xor XOR2 (N437, N431, N69);
buf BUF1 (N438, N428);
not NOT1 (N439, N423);
buf BUF1 (N440, N434);
nand NAND4 (N441, N413, N302, N58, N206);
nand NAND2 (N442, N433, N423);
nor NOR3 (N443, N436, N279, N94);
or OR4 (N444, N438, N42, N284, N402);
not NOT1 (N445, N443);
nor NOR3 (N446, N427, N246, N425);
or OR3 (N447, N442, N177, N362);
not NOT1 (N448, N437);
nor NOR2 (N449, N444, N37);
buf BUF1 (N450, N447);
and AND3 (N451, N440, N245, N239);
buf BUF1 (N452, N448);
xor XOR2 (N453, N435, N389);
nand NAND2 (N454, N446, N193);
nor NOR2 (N455, N452, N353);
or OR3 (N456, N451, N34, N321);
xor XOR2 (N457, N455, N347);
buf BUF1 (N458, N456);
not NOT1 (N459, N450);
not NOT1 (N460, N457);
buf BUF1 (N461, N458);
and AND3 (N462, N454, N65, N377);
nand NAND4 (N463, N460, N33, N312, N378);
buf BUF1 (N464, N421);
not NOT1 (N465, N463);
nor NOR3 (N466, N462, N202, N62);
or OR2 (N467, N465, N275);
buf BUF1 (N468, N441);
nand NAND3 (N469, N466, N257, N423);
xor XOR2 (N470, N469, N272);
nand NAND4 (N471, N449, N292, N267, N389);
or OR4 (N472, N445, N146, N169, N390);
nand NAND3 (N473, N471, N192, N226);
nand NAND3 (N474, N473, N83, N142);
xor XOR2 (N475, N464, N307);
buf BUF1 (N476, N459);
buf BUF1 (N477, N461);
nand NAND2 (N478, N472, N430);
nand NAND3 (N479, N477, N18, N371);
nor NOR4 (N480, N475, N168, N97, N276);
or OR2 (N481, N476, N81);
nand NAND4 (N482, N480, N195, N30, N451);
nor NOR4 (N483, N467, N227, N383, N216);
and AND2 (N484, N479, N65);
nor NOR4 (N485, N484, N477, N167, N166);
not NOT1 (N486, N481);
or OR4 (N487, N483, N177, N46, N440);
or OR2 (N488, N485, N185);
xor XOR2 (N489, N474, N357);
nor NOR4 (N490, N482, N284, N353, N6);
or OR3 (N491, N453, N397, N386);
buf BUF1 (N492, N468);
not NOT1 (N493, N470);
or OR3 (N494, N490, N74, N163);
and AND2 (N495, N492, N20);
xor XOR2 (N496, N495, N439);
buf BUF1 (N497, N379);
and AND3 (N498, N478, N160, N66);
nand NAND2 (N499, N498, N87);
xor XOR2 (N500, N499, N25);
and AND3 (N501, N486, N470, N391);
buf BUF1 (N502, N500);
nor NOR4 (N503, N488, N74, N297, N140);
nand NAND3 (N504, N489, N280, N110);
and AND3 (N505, N502, N334, N495);
nor NOR4 (N506, N503, N259, N435, N359);
nand NAND4 (N507, N505, N486, N239, N95);
xor XOR2 (N508, N496, N145);
or OR3 (N509, N507, N210, N179);
or OR2 (N510, N493, N23);
buf BUF1 (N511, N491);
or OR4 (N512, N501, N423, N305, N161);
xor XOR2 (N513, N506, N22);
or OR4 (N514, N511, N342, N504, N277);
not NOT1 (N515, N245);
or OR4 (N516, N510, N131, N346, N9);
buf BUF1 (N517, N513);
and AND3 (N518, N487, N360, N291);
or OR3 (N519, N515, N326, N206);
and AND2 (N520, N494, N273);
and AND4 (N521, N518, N176, N417, N193);
xor XOR2 (N522, N517, N230);
buf BUF1 (N523, N497);
nand NAND4 (N524, N512, N64, N99, N365);
buf BUF1 (N525, N522);
not NOT1 (N526, N514);
and AND3 (N527, N526, N195, N11);
or OR4 (N528, N516, N73, N255, N96);
xor XOR2 (N529, N524, N43);
and AND4 (N530, N509, N429, N489, N489);
or OR4 (N531, N527, N230, N72, N388);
xor XOR2 (N532, N523, N357);
and AND3 (N533, N532, N227, N359);
and AND3 (N534, N525, N454, N188);
xor XOR2 (N535, N528, N64);
nand NAND2 (N536, N520, N317);
or OR4 (N537, N535, N400, N226, N351);
and AND2 (N538, N521, N190);
or OR2 (N539, N508, N478);
nand NAND4 (N540, N534, N313, N446, N49);
not NOT1 (N541, N537);
or OR2 (N542, N538, N299);
nor NOR4 (N543, N519, N111, N154, N413);
and AND3 (N544, N536, N35, N9);
and AND4 (N545, N529, N514, N297, N542);
or OR2 (N546, N2, N24);
and AND2 (N547, N545, N167);
nand NAND2 (N548, N546, N387);
nor NOR3 (N549, N539, N307, N542);
nor NOR2 (N550, N548, N366);
nand NAND2 (N551, N550, N243);
and AND2 (N552, N551, N490);
not NOT1 (N553, N543);
not NOT1 (N554, N544);
nor NOR4 (N555, N554, N84, N423, N36);
nand NAND3 (N556, N555, N162, N327);
nand NAND4 (N557, N553, N182, N484, N488);
nand NAND3 (N558, N533, N417, N499);
xor XOR2 (N559, N552, N159);
not NOT1 (N560, N558);
or OR4 (N561, N556, N102, N428, N139);
not NOT1 (N562, N560);
and AND2 (N563, N561, N292);
or OR3 (N564, N540, N367, N282);
nor NOR2 (N565, N530, N494);
nor NOR2 (N566, N562, N250);
or OR2 (N567, N549, N17);
nand NAND2 (N568, N566, N449);
xor XOR2 (N569, N567, N261);
and AND4 (N570, N564, N29, N311, N2);
and AND2 (N571, N563, N268);
not NOT1 (N572, N559);
nand NAND4 (N573, N571, N203, N403, N216);
nand NAND2 (N574, N557, N329);
nand NAND2 (N575, N565, N57);
or OR2 (N576, N569, N71);
not NOT1 (N577, N547);
xor XOR2 (N578, N577, N137);
buf BUF1 (N579, N575);
xor XOR2 (N580, N568, N306);
nor NOR4 (N581, N570, N188, N446, N76);
buf BUF1 (N582, N580);
and AND3 (N583, N582, N528, N145);
or OR4 (N584, N579, N128, N508, N368);
xor XOR2 (N585, N541, N559);
nand NAND4 (N586, N574, N59, N496, N428);
not NOT1 (N587, N576);
nor NOR3 (N588, N583, N391, N78);
buf BUF1 (N589, N581);
or OR2 (N590, N578, N520);
not NOT1 (N591, N587);
not NOT1 (N592, N584);
xor XOR2 (N593, N585, N276);
buf BUF1 (N594, N589);
and AND4 (N595, N591, N526, N426, N213);
nor NOR3 (N596, N573, N370, N246);
not NOT1 (N597, N572);
nor NOR3 (N598, N588, N402, N502);
or OR3 (N599, N597, N267, N481);
nand NAND4 (N600, N531, N280, N126, N571);
buf BUF1 (N601, N600);
nor NOR3 (N602, N593, N491, N486);
nor NOR4 (N603, N592, N146, N323, N332);
nand NAND4 (N604, N602, N413, N53, N560);
or OR3 (N605, N599, N430, N357);
nand NAND2 (N606, N590, N433);
buf BUF1 (N607, N601);
buf BUF1 (N608, N604);
or OR3 (N609, N605, N590, N54);
or OR2 (N610, N598, N183);
not NOT1 (N611, N610);
xor XOR2 (N612, N596, N239);
not NOT1 (N613, N609);
nor NOR4 (N614, N586, N95, N90, N339);
nand NAND3 (N615, N606, N319, N137);
not NOT1 (N616, N612);
not NOT1 (N617, N607);
xor XOR2 (N618, N594, N388);
xor XOR2 (N619, N613, N133);
buf BUF1 (N620, N616);
not NOT1 (N621, N617);
nand NAND2 (N622, N620, N362);
or OR4 (N623, N621, N514, N81, N270);
not NOT1 (N624, N603);
buf BUF1 (N625, N614);
not NOT1 (N626, N608);
not NOT1 (N627, N625);
xor XOR2 (N628, N624, N445);
or OR2 (N629, N611, N358);
not NOT1 (N630, N595);
and AND4 (N631, N619, N115, N478, N608);
nand NAND4 (N632, N623, N378, N44, N334);
buf BUF1 (N633, N629);
buf BUF1 (N634, N615);
nor NOR3 (N635, N633, N142, N59);
nand NAND2 (N636, N622, N223);
buf BUF1 (N637, N632);
xor XOR2 (N638, N630, N620);
nor NOR3 (N639, N636, N577, N477);
xor XOR2 (N640, N627, N27);
not NOT1 (N641, N639);
buf BUF1 (N642, N634);
not NOT1 (N643, N641);
not NOT1 (N644, N631);
not NOT1 (N645, N637);
or OR3 (N646, N640, N421, N114);
nor NOR2 (N647, N638, N373);
and AND2 (N648, N628, N317);
buf BUF1 (N649, N635);
and AND3 (N650, N626, N7, N552);
nor NOR4 (N651, N648, N252, N58, N252);
not NOT1 (N652, N645);
not NOT1 (N653, N647);
xor XOR2 (N654, N653, N610);
xor XOR2 (N655, N651, N218);
and AND4 (N656, N654, N8, N106, N496);
not NOT1 (N657, N650);
xor XOR2 (N658, N618, N311);
nand NAND3 (N659, N642, N540, N106);
buf BUF1 (N660, N644);
xor XOR2 (N661, N646, N445);
nor NOR4 (N662, N655, N326, N27, N416);
or OR3 (N663, N659, N344, N551);
nor NOR4 (N664, N662, N401, N644, N175);
and AND4 (N665, N660, N233, N470, N589);
buf BUF1 (N666, N665);
not NOT1 (N667, N666);
not NOT1 (N668, N657);
or OR4 (N669, N664, N347, N337, N436);
and AND2 (N670, N652, N491);
or OR3 (N671, N670, N471, N209);
nor NOR3 (N672, N649, N183, N195);
or OR4 (N673, N656, N65, N302, N301);
not NOT1 (N674, N669);
nor NOR2 (N675, N663, N453);
and AND4 (N676, N668, N446, N501, N489);
buf BUF1 (N677, N667);
buf BUF1 (N678, N672);
or OR2 (N679, N674, N131);
or OR2 (N680, N676, N269);
not NOT1 (N681, N643);
nand NAND2 (N682, N675, N220);
or OR4 (N683, N671, N679, N32, N335);
nor NOR2 (N684, N107, N101);
and AND2 (N685, N661, N358);
xor XOR2 (N686, N677, N630);
or OR3 (N687, N684, N353, N240);
and AND4 (N688, N681, N318, N258, N637);
nor NOR2 (N689, N682, N35);
not NOT1 (N690, N678);
xor XOR2 (N691, N683, N20);
and AND4 (N692, N685, N561, N639, N38);
nor NOR3 (N693, N688, N571, N584);
or OR2 (N694, N658, N325);
nand NAND4 (N695, N694, N462, N102, N12);
or OR3 (N696, N673, N256, N158);
not NOT1 (N697, N696);
nand NAND3 (N698, N697, N298, N307);
nand NAND3 (N699, N691, N199, N352);
xor XOR2 (N700, N692, N486);
buf BUF1 (N701, N687);
buf BUF1 (N702, N699);
xor XOR2 (N703, N700, N624);
not NOT1 (N704, N702);
nor NOR3 (N705, N703, N398, N54);
xor XOR2 (N706, N686, N531);
nor NOR4 (N707, N695, N161, N675, N584);
nand NAND2 (N708, N707, N654);
nor NOR2 (N709, N701, N287);
xor XOR2 (N710, N705, N272);
not NOT1 (N711, N680);
and AND3 (N712, N710, N354, N645);
nor NOR2 (N713, N689, N637);
not NOT1 (N714, N711);
or OR3 (N715, N706, N633, N335);
buf BUF1 (N716, N715);
or OR4 (N717, N708, N198, N649, N475);
nor NOR4 (N718, N712, N413, N251, N663);
nand NAND4 (N719, N704, N591, N205, N578);
or OR3 (N720, N709, N25, N287);
or OR3 (N721, N718, N564, N120);
nand NAND2 (N722, N717, N342);
and AND2 (N723, N720, N440);
and AND4 (N724, N722, N676, N596, N328);
buf BUF1 (N725, N724);
nand NAND2 (N726, N713, N558);
buf BUF1 (N727, N714);
and AND3 (N728, N719, N680, N723);
xor XOR2 (N729, N539, N593);
buf BUF1 (N730, N690);
and AND2 (N731, N725, N331);
or OR4 (N732, N731, N703, N365, N123);
or OR4 (N733, N727, N698, N675, N243);
or OR2 (N734, N147, N548);
and AND3 (N735, N728, N409, N279);
xor XOR2 (N736, N733, N13);
buf BUF1 (N737, N721);
nand NAND3 (N738, N732, N36, N683);
buf BUF1 (N739, N726);
nand NAND4 (N740, N734, N621, N197, N83);
and AND4 (N741, N716, N500, N233, N601);
or OR4 (N742, N741, N449, N451, N706);
buf BUF1 (N743, N693);
not NOT1 (N744, N742);
xor XOR2 (N745, N744, N318);
not NOT1 (N746, N740);
nor NOR4 (N747, N743, N551, N514, N590);
nand NAND2 (N748, N738, N136);
and AND3 (N749, N730, N555, N131);
nor NOR3 (N750, N729, N501, N122);
buf BUF1 (N751, N737);
xor XOR2 (N752, N739, N568);
or OR3 (N753, N748, N285, N332);
nand NAND3 (N754, N745, N449, N28);
xor XOR2 (N755, N749, N706);
or OR4 (N756, N755, N413, N226, N89);
nor NOR3 (N757, N750, N329, N27);
nor NOR2 (N758, N753, N609);
buf BUF1 (N759, N752);
xor XOR2 (N760, N751, N114);
and AND4 (N761, N754, N759, N186, N312);
not NOT1 (N762, N458);
not NOT1 (N763, N762);
nor NOR3 (N764, N736, N11, N456);
nand NAND3 (N765, N758, N358, N264);
buf BUF1 (N766, N760);
xor XOR2 (N767, N747, N461);
nor NOR2 (N768, N757, N270);
or OR2 (N769, N765, N617);
or OR2 (N770, N763, N227);
xor XOR2 (N771, N770, N380);
and AND3 (N772, N768, N564, N285);
or OR4 (N773, N756, N357, N175, N731);
buf BUF1 (N774, N735);
not NOT1 (N775, N774);
or OR3 (N776, N773, N249, N46);
or OR4 (N777, N775, N24, N212, N67);
nand NAND2 (N778, N766, N316);
nor NOR2 (N779, N772, N310);
buf BUF1 (N780, N764);
or OR4 (N781, N777, N681, N682, N575);
and AND4 (N782, N769, N668, N276, N582);
and AND2 (N783, N780, N231);
buf BUF1 (N784, N761);
or OR2 (N785, N776, N250);
and AND3 (N786, N778, N568, N297);
xor XOR2 (N787, N784, N5);
xor XOR2 (N788, N783, N353);
not NOT1 (N789, N788);
and AND2 (N790, N789, N319);
nand NAND3 (N791, N781, N391, N14);
or OR3 (N792, N782, N602, N302);
nor NOR4 (N793, N790, N320, N234, N386);
nor NOR4 (N794, N767, N438, N271, N84);
buf BUF1 (N795, N792);
buf BUF1 (N796, N779);
not NOT1 (N797, N791);
not NOT1 (N798, N746);
xor XOR2 (N799, N771, N327);
and AND3 (N800, N796, N727, N61);
xor XOR2 (N801, N797, N113);
or OR4 (N802, N793, N570, N254, N499);
or OR2 (N803, N802, N378);
or OR3 (N804, N803, N342, N86);
nand NAND4 (N805, N798, N665, N284, N17);
xor XOR2 (N806, N804, N508);
nand NAND4 (N807, N785, N626, N94, N564);
or OR2 (N808, N805, N323);
nor NOR3 (N809, N806, N304, N790);
and AND4 (N810, N795, N759, N103, N171);
xor XOR2 (N811, N807, N160);
nand NAND2 (N812, N810, N349);
xor XOR2 (N813, N801, N494);
not NOT1 (N814, N808);
or OR4 (N815, N800, N601, N683, N314);
or OR3 (N816, N815, N489, N6);
buf BUF1 (N817, N787);
buf BUF1 (N818, N786);
and AND3 (N819, N813, N293, N27);
and AND2 (N820, N809, N742);
buf BUF1 (N821, N818);
xor XOR2 (N822, N794, N122);
nand NAND3 (N823, N819, N724, N555);
xor XOR2 (N824, N814, N181);
nor NOR3 (N825, N799, N777, N737);
buf BUF1 (N826, N816);
nand NAND3 (N827, N826, N61, N196);
nor NOR2 (N828, N821, N496);
and AND4 (N829, N824, N18, N769, N739);
or OR4 (N830, N822, N443, N588, N233);
nand NAND4 (N831, N812, N714, N226, N27);
nand NAND3 (N832, N820, N88, N233);
not NOT1 (N833, N831);
not NOT1 (N834, N811);
or OR3 (N835, N827, N256, N435);
not NOT1 (N836, N834);
nand NAND2 (N837, N832, N457);
or OR3 (N838, N830, N505, N106);
not NOT1 (N839, N837);
buf BUF1 (N840, N823);
and AND2 (N841, N829, N109);
and AND4 (N842, N841, N796, N177, N293);
and AND3 (N843, N825, N476, N114);
or OR4 (N844, N838, N419, N379, N491);
nand NAND3 (N845, N833, N316, N563);
and AND4 (N846, N844, N734, N196, N832);
and AND4 (N847, N835, N63, N100, N500);
xor XOR2 (N848, N836, N144);
not NOT1 (N849, N843);
not NOT1 (N850, N842);
and AND2 (N851, N828, N672);
or OR2 (N852, N851, N709);
or OR2 (N853, N839, N182);
buf BUF1 (N854, N846);
not NOT1 (N855, N854);
nand NAND4 (N856, N847, N214, N666, N221);
and AND4 (N857, N856, N354, N734, N592);
buf BUF1 (N858, N817);
not NOT1 (N859, N852);
xor XOR2 (N860, N859, N432);
nor NOR2 (N861, N860, N684);
buf BUF1 (N862, N855);
not NOT1 (N863, N858);
xor XOR2 (N864, N863, N712);
nand NAND3 (N865, N840, N386, N754);
xor XOR2 (N866, N861, N291);
nor NOR2 (N867, N857, N58);
nand NAND4 (N868, N849, N342, N471, N858);
xor XOR2 (N869, N848, N82);
nor NOR4 (N870, N866, N73, N775, N792);
and AND4 (N871, N867, N566, N36, N208);
xor XOR2 (N872, N868, N342);
and AND4 (N873, N872, N788, N756, N213);
xor XOR2 (N874, N862, N90);
nor NOR4 (N875, N853, N492, N7, N125);
and AND3 (N876, N870, N251, N539);
not NOT1 (N877, N871);
and AND4 (N878, N869, N421, N491, N225);
and AND4 (N879, N875, N576, N809, N280);
or OR3 (N880, N873, N24, N598);
nor NOR3 (N881, N876, N560, N623);
nor NOR4 (N882, N877, N809, N26, N837);
or OR3 (N883, N864, N428, N369);
nand NAND2 (N884, N845, N759);
xor XOR2 (N885, N879, N504);
and AND4 (N886, N885, N126, N819, N52);
nor NOR3 (N887, N883, N396, N150);
and AND4 (N888, N886, N125, N106, N873);
nor NOR2 (N889, N878, N585);
nand NAND4 (N890, N865, N457, N874, N529);
and AND4 (N891, N277, N828, N157, N407);
nor NOR4 (N892, N881, N311, N132, N244);
nor NOR2 (N893, N882, N162);
not NOT1 (N894, N891);
nand NAND3 (N895, N890, N651, N63);
nor NOR2 (N896, N850, N149);
not NOT1 (N897, N884);
and AND2 (N898, N897, N111);
and AND3 (N899, N889, N274, N226);
nand NAND2 (N900, N887, N489);
xor XOR2 (N901, N900, N161);
and AND3 (N902, N895, N329, N429);
nor NOR3 (N903, N902, N142, N826);
buf BUF1 (N904, N898);
xor XOR2 (N905, N903, N824);
and AND2 (N906, N888, N418);
nor NOR3 (N907, N904, N687, N21);
nor NOR3 (N908, N907, N589, N171);
nand NAND3 (N909, N899, N843, N68);
not NOT1 (N910, N880);
nand NAND2 (N911, N894, N367);
and AND4 (N912, N892, N486, N748, N485);
or OR2 (N913, N896, N863);
nor NOR3 (N914, N913, N212, N560);
or OR4 (N915, N893, N789, N126, N266);
nand NAND2 (N916, N914, N300);
nand NAND2 (N917, N912, N636);
nor NOR4 (N918, N906, N811, N817, N246);
or OR3 (N919, N908, N529, N380);
or OR2 (N920, N918, N130);
and AND3 (N921, N910, N578, N377);
not NOT1 (N922, N916);
nand NAND3 (N923, N911, N918, N405);
not NOT1 (N924, N905);
buf BUF1 (N925, N921);
nor NOR3 (N926, N909, N274, N61);
not NOT1 (N927, N925);
nand NAND3 (N928, N922, N46, N458);
nand NAND3 (N929, N928, N83, N153);
not NOT1 (N930, N915);
or OR3 (N931, N926, N637, N807);
xor XOR2 (N932, N927, N520);
buf BUF1 (N933, N929);
buf BUF1 (N934, N932);
and AND2 (N935, N934, N756);
and AND4 (N936, N919, N812, N788, N440);
nor NOR3 (N937, N935, N296, N265);
and AND2 (N938, N924, N792);
not NOT1 (N939, N901);
nor NOR2 (N940, N923, N428);
not NOT1 (N941, N938);
and AND2 (N942, N930, N22);
nor NOR4 (N943, N933, N262, N936, N810);
xor XOR2 (N944, N503, N869);
or OR4 (N945, N944, N426, N829, N163);
and AND3 (N946, N943, N471, N409);
nor NOR3 (N947, N939, N652, N762);
buf BUF1 (N948, N917);
nor NOR3 (N949, N931, N432, N650);
buf BUF1 (N950, N948);
buf BUF1 (N951, N950);
or OR3 (N952, N946, N519, N230);
and AND4 (N953, N937, N538, N285, N655);
buf BUF1 (N954, N941);
nand NAND4 (N955, N942, N380, N60, N810);
not NOT1 (N956, N940);
xor XOR2 (N957, N945, N579);
nor NOR2 (N958, N953, N303);
buf BUF1 (N959, N951);
nand NAND3 (N960, N957, N942, N636);
or OR3 (N961, N958, N789, N617);
xor XOR2 (N962, N949, N765);
xor XOR2 (N963, N955, N648);
or OR2 (N964, N961, N693);
or OR3 (N965, N920, N301, N324);
and AND2 (N966, N954, N59);
xor XOR2 (N967, N960, N109);
nor NOR4 (N968, N967, N264, N489, N958);
and AND2 (N969, N965, N55);
not NOT1 (N970, N956);
buf BUF1 (N971, N969);
buf BUF1 (N972, N952);
buf BUF1 (N973, N962);
or OR2 (N974, N947, N65);
nand NAND3 (N975, N972, N161, N10);
or OR3 (N976, N964, N798, N928);
nand NAND4 (N977, N976, N711, N212, N664);
buf BUF1 (N978, N975);
or OR4 (N979, N970, N181, N696, N426);
buf BUF1 (N980, N977);
not NOT1 (N981, N980);
nor NOR4 (N982, N979, N278, N716, N2);
nor NOR2 (N983, N981, N75);
buf BUF1 (N984, N983);
or OR2 (N985, N974, N635);
nor NOR2 (N986, N963, N69);
buf BUF1 (N987, N973);
buf BUF1 (N988, N987);
and AND2 (N989, N984, N725);
nand NAND2 (N990, N989, N694);
buf BUF1 (N991, N986);
nor NOR3 (N992, N978, N960, N551);
not NOT1 (N993, N966);
nand NAND2 (N994, N990, N51);
and AND4 (N995, N992, N242, N959, N170);
and AND3 (N996, N761, N774, N460);
not NOT1 (N997, N991);
buf BUF1 (N998, N988);
xor XOR2 (N999, N995, N814);
nand NAND3 (N1000, N985, N294, N751);
xor XOR2 (N1001, N994, N855);
nor NOR4 (N1002, N1000, N636, N463, N217);
and AND4 (N1003, N993, N817, N746, N387);
not NOT1 (N1004, N982);
or OR2 (N1005, N968, N886);
xor XOR2 (N1006, N1005, N538);
and AND2 (N1007, N971, N438);
or OR3 (N1008, N1002, N688, N1006);
nor NOR3 (N1009, N556, N152, N379);
nor NOR3 (N1010, N997, N580, N843);
or OR4 (N1011, N999, N365, N239, N98);
not NOT1 (N1012, N1010);
or OR4 (N1013, N998, N193, N754, N461);
nor NOR4 (N1014, N1008, N95, N666, N21);
xor XOR2 (N1015, N1013, N801);
nor NOR3 (N1016, N1003, N213, N889);
nand NAND4 (N1017, N1012, N56, N522, N758);
nor NOR2 (N1018, N1009, N423);
nor NOR3 (N1019, N1015, N629, N156);
or OR4 (N1020, N1014, N317, N349, N956);
nand NAND4 (N1021, N1019, N816, N831, N282);
xor XOR2 (N1022, N996, N915);
nand NAND4 (N1023, N1017, N1009, N362, N244);
not NOT1 (N1024, N1022);
nor NOR3 (N1025, N1016, N796, N574);
or OR2 (N1026, N1021, N47);
or OR3 (N1027, N1001, N672, N686);
nor NOR3 (N1028, N1023, N81, N448);
or OR3 (N1029, N1025, N658, N995);
and AND2 (N1030, N1029, N584);
nor NOR4 (N1031, N1027, N1015, N402, N304);
nor NOR3 (N1032, N1024, N114, N961);
nor NOR4 (N1033, N1020, N196, N783, N602);
and AND2 (N1034, N1028, N486);
buf BUF1 (N1035, N1007);
nand NAND4 (N1036, N1004, N688, N156, N546);
nand NAND3 (N1037, N1011, N536, N835);
xor XOR2 (N1038, N1034, N717);
buf BUF1 (N1039, N1031);
nor NOR3 (N1040, N1033, N460, N971);
not NOT1 (N1041, N1040);
xor XOR2 (N1042, N1026, N794);
xor XOR2 (N1043, N1018, N379);
buf BUF1 (N1044, N1030);
xor XOR2 (N1045, N1037, N1038);
nand NAND3 (N1046, N340, N682, N782);
or OR2 (N1047, N1045, N863);
buf BUF1 (N1048, N1041);
nor NOR3 (N1049, N1046, N803, N130);
xor XOR2 (N1050, N1032, N842);
not NOT1 (N1051, N1049);
and AND2 (N1052, N1048, N428);
or OR2 (N1053, N1035, N526);
not NOT1 (N1054, N1051);
nand NAND3 (N1055, N1043, N537, N678);
and AND2 (N1056, N1044, N922);
nand NAND2 (N1057, N1053, N768);
nand NAND3 (N1058, N1036, N473, N1030);
xor XOR2 (N1059, N1039, N116);
nand NAND2 (N1060, N1058, N362);
not NOT1 (N1061, N1060);
xor XOR2 (N1062, N1052, N129);
not NOT1 (N1063, N1050);
xor XOR2 (N1064, N1055, N114);
nor NOR3 (N1065, N1054, N420, N368);
or OR2 (N1066, N1057, N488);
not NOT1 (N1067, N1066);
nand NAND4 (N1068, N1065, N168, N895, N1064);
or OR4 (N1069, N59, N584, N486, N1025);
xor XOR2 (N1070, N1069, N797);
nand NAND4 (N1071, N1059, N672, N850, N254);
nor NOR4 (N1072, N1056, N298, N541, N170);
and AND4 (N1073, N1062, N326, N288, N108);
buf BUF1 (N1074, N1067);
not NOT1 (N1075, N1070);
xor XOR2 (N1076, N1075, N734);
and AND2 (N1077, N1047, N1040);
xor XOR2 (N1078, N1071, N3);
nand NAND4 (N1079, N1077, N745, N172, N1036);
nand NAND4 (N1080, N1072, N309, N872, N38);
not NOT1 (N1081, N1068);
nor NOR4 (N1082, N1074, N918, N1073, N604);
buf BUF1 (N1083, N536);
xor XOR2 (N1084, N1061, N395);
not NOT1 (N1085, N1076);
or OR2 (N1086, N1042, N791);
xor XOR2 (N1087, N1085, N1045);
or OR3 (N1088, N1086, N869, N905);
not NOT1 (N1089, N1078);
nor NOR4 (N1090, N1089, N841, N256, N803);
not NOT1 (N1091, N1090);
buf BUF1 (N1092, N1083);
or OR3 (N1093, N1084, N1069, N759);
buf BUF1 (N1094, N1092);
buf BUF1 (N1095, N1082);
xor XOR2 (N1096, N1063, N98);
not NOT1 (N1097, N1080);
not NOT1 (N1098, N1088);
or OR4 (N1099, N1093, N949, N182, N1036);
nand NAND3 (N1100, N1097, N591, N366);
nor NOR3 (N1101, N1091, N140, N764);
nor NOR2 (N1102, N1087, N1006);
nor NOR3 (N1103, N1096, N307, N534);
nor NOR2 (N1104, N1100, N346);
buf BUF1 (N1105, N1081);
not NOT1 (N1106, N1105);
not NOT1 (N1107, N1102);
nor NOR2 (N1108, N1104, N853);
buf BUF1 (N1109, N1103);
buf BUF1 (N1110, N1107);
not NOT1 (N1111, N1098);
not NOT1 (N1112, N1111);
nor NOR2 (N1113, N1106, N614);
buf BUF1 (N1114, N1099);
and AND4 (N1115, N1113, N758, N408, N997);
nor NOR3 (N1116, N1094, N543, N993);
buf BUF1 (N1117, N1110);
or OR2 (N1118, N1116, N627);
or OR2 (N1119, N1114, N413);
xor XOR2 (N1120, N1115, N1056);
and AND2 (N1121, N1120, N394);
or OR4 (N1122, N1119, N422, N639, N61);
xor XOR2 (N1123, N1118, N258);
xor XOR2 (N1124, N1121, N962);
xor XOR2 (N1125, N1079, N594);
or OR2 (N1126, N1112, N492);
and AND3 (N1127, N1109, N25, N708);
not NOT1 (N1128, N1127);
or OR3 (N1129, N1123, N916, N900);
xor XOR2 (N1130, N1124, N1055);
nand NAND4 (N1131, N1095, N333, N1023, N106);
and AND3 (N1132, N1125, N712, N542);
nor NOR4 (N1133, N1126, N401, N1103, N862);
buf BUF1 (N1134, N1130);
and AND2 (N1135, N1108, N522);
not NOT1 (N1136, N1117);
xor XOR2 (N1137, N1133, N1067);
xor XOR2 (N1138, N1122, N166);
buf BUF1 (N1139, N1134);
or OR4 (N1140, N1135, N724, N639, N330);
xor XOR2 (N1141, N1140, N584);
not NOT1 (N1142, N1138);
nor NOR3 (N1143, N1132, N1002, N798);
or OR2 (N1144, N1128, N169);
and AND3 (N1145, N1141, N160, N801);
nand NAND3 (N1146, N1145, N308, N216);
xor XOR2 (N1147, N1142, N1079);
nor NOR2 (N1148, N1136, N346);
nor NOR4 (N1149, N1147, N1064, N271, N786);
nor NOR2 (N1150, N1149, N64);
or OR3 (N1151, N1131, N155, N1046);
nand NAND4 (N1152, N1139, N25, N294, N727);
not NOT1 (N1153, N1152);
and AND3 (N1154, N1146, N498, N272);
and AND3 (N1155, N1144, N64, N1107);
nor NOR4 (N1156, N1148, N1150, N856, N162);
and AND2 (N1157, N989, N287);
xor XOR2 (N1158, N1129, N674);
nor NOR4 (N1159, N1156, N327, N881, N703);
buf BUF1 (N1160, N1158);
and AND4 (N1161, N1155, N1134, N239, N416);
nor NOR2 (N1162, N1160, N179);
buf BUF1 (N1163, N1159);
nand NAND2 (N1164, N1101, N379);
buf BUF1 (N1165, N1161);
nand NAND2 (N1166, N1157, N824);
buf BUF1 (N1167, N1143);
nand NAND2 (N1168, N1151, N529);
nor NOR2 (N1169, N1162, N668);
nor NOR2 (N1170, N1154, N345);
nand NAND4 (N1171, N1167, N66, N83, N531);
nand NAND2 (N1172, N1170, N1127);
xor XOR2 (N1173, N1171, N749);
xor XOR2 (N1174, N1153, N539);
not NOT1 (N1175, N1164);
xor XOR2 (N1176, N1175, N950);
xor XOR2 (N1177, N1172, N505);
not NOT1 (N1178, N1168);
and AND4 (N1179, N1169, N356, N707, N846);
nand NAND4 (N1180, N1173, N369, N620, N10);
not NOT1 (N1181, N1177);
nor NOR3 (N1182, N1181, N146, N384);
nand NAND2 (N1183, N1163, N149);
and AND4 (N1184, N1165, N23, N996, N257);
buf BUF1 (N1185, N1137);
buf BUF1 (N1186, N1179);
or OR4 (N1187, N1180, N87, N610, N302);
buf BUF1 (N1188, N1178);
nand NAND2 (N1189, N1188, N816);
xor XOR2 (N1190, N1174, N330);
not NOT1 (N1191, N1176);
buf BUF1 (N1192, N1184);
and AND4 (N1193, N1186, N970, N927, N927);
buf BUF1 (N1194, N1192);
not NOT1 (N1195, N1194);
or OR4 (N1196, N1193, N783, N858, N720);
nand NAND3 (N1197, N1185, N815, N807);
and AND2 (N1198, N1187, N883);
or OR4 (N1199, N1166, N852, N287, N811);
xor XOR2 (N1200, N1190, N400);
or OR2 (N1201, N1200, N709);
or OR2 (N1202, N1198, N1116);
or OR3 (N1203, N1201, N232, N473);
nand NAND3 (N1204, N1182, N329, N527);
buf BUF1 (N1205, N1191);
or OR4 (N1206, N1196, N1194, N1196, N608);
nand NAND2 (N1207, N1202, N180);
nand NAND2 (N1208, N1206, N1054);
buf BUF1 (N1209, N1199);
xor XOR2 (N1210, N1209, N35);
and AND3 (N1211, N1207, N370, N905);
buf BUF1 (N1212, N1208);
buf BUF1 (N1213, N1205);
buf BUF1 (N1214, N1203);
nor NOR4 (N1215, N1213, N280, N912, N745);
and AND3 (N1216, N1197, N384, N427);
or OR2 (N1217, N1189, N151);
and AND4 (N1218, N1212, N541, N110, N334);
nor NOR3 (N1219, N1216, N750, N54);
buf BUF1 (N1220, N1204);
and AND2 (N1221, N1211, N164);
nor NOR3 (N1222, N1218, N82, N316);
xor XOR2 (N1223, N1195, N586);
not NOT1 (N1224, N1219);
not NOT1 (N1225, N1210);
or OR2 (N1226, N1225, N1225);
nand NAND4 (N1227, N1217, N894, N172, N317);
buf BUF1 (N1228, N1220);
xor XOR2 (N1229, N1227, N710);
nand NAND4 (N1230, N1224, N1040, N386, N1031);
nand NAND3 (N1231, N1221, N283, N110);
or OR4 (N1232, N1228, N1150, N219, N935);
xor XOR2 (N1233, N1230, N782);
buf BUF1 (N1234, N1222);
xor XOR2 (N1235, N1229, N942);
and AND3 (N1236, N1183, N272, N270);
or OR4 (N1237, N1215, N964, N1035, N697);
and AND3 (N1238, N1232, N436, N161);
nand NAND2 (N1239, N1233, N1030);
and AND2 (N1240, N1236, N50);
buf BUF1 (N1241, N1235);
or OR3 (N1242, N1231, N229, N107);
not NOT1 (N1243, N1242);
buf BUF1 (N1244, N1237);
xor XOR2 (N1245, N1243, N1005);
xor XOR2 (N1246, N1245, N1207);
or OR2 (N1247, N1223, N1185);
not NOT1 (N1248, N1241);
nor NOR2 (N1249, N1226, N154);
not NOT1 (N1250, N1239);
or OR2 (N1251, N1244, N893);
and AND4 (N1252, N1248, N1142, N494, N458);
nand NAND3 (N1253, N1234, N739, N284);
buf BUF1 (N1254, N1252);
not NOT1 (N1255, N1250);
not NOT1 (N1256, N1255);
and AND2 (N1257, N1246, N245);
nand NAND2 (N1258, N1214, N766);
and AND3 (N1259, N1258, N454, N922);
not NOT1 (N1260, N1238);
nand NAND4 (N1261, N1240, N449, N116, N1100);
nand NAND3 (N1262, N1259, N1249, N1237);
xor XOR2 (N1263, N864, N348);
buf BUF1 (N1264, N1253);
nand NAND2 (N1265, N1257, N1226);
and AND4 (N1266, N1261, N667, N753, N724);
xor XOR2 (N1267, N1265, N347);
xor XOR2 (N1268, N1254, N8);
and AND3 (N1269, N1264, N8, N964);
or OR4 (N1270, N1262, N744, N315, N710);
nor NOR3 (N1271, N1247, N1074, N403);
buf BUF1 (N1272, N1260);
nand NAND4 (N1273, N1256, N250, N1203, N1268);
nand NAND3 (N1274, N589, N387, N863);
nand NAND2 (N1275, N1267, N759);
nand NAND2 (N1276, N1271, N43);
nor NOR2 (N1277, N1273, N343);
xor XOR2 (N1278, N1270, N939);
nor NOR2 (N1279, N1263, N67);
nor NOR3 (N1280, N1278, N151, N556);
or OR2 (N1281, N1277, N1177);
buf BUF1 (N1282, N1275);
xor XOR2 (N1283, N1280, N65);
xor XOR2 (N1284, N1282, N1282);
and AND4 (N1285, N1272, N993, N343, N1154);
and AND3 (N1286, N1251, N1070, N960);
buf BUF1 (N1287, N1274);
xor XOR2 (N1288, N1269, N680);
not NOT1 (N1289, N1286);
buf BUF1 (N1290, N1288);
xor XOR2 (N1291, N1281, N907);
buf BUF1 (N1292, N1291);
not NOT1 (N1293, N1287);
xor XOR2 (N1294, N1292, N1288);
xor XOR2 (N1295, N1279, N463);
buf BUF1 (N1296, N1276);
or OR4 (N1297, N1289, N558, N1243, N324);
nand NAND3 (N1298, N1283, N1008, N889);
buf BUF1 (N1299, N1295);
nor NOR4 (N1300, N1293, N328, N116, N810);
nor NOR2 (N1301, N1297, N521);
nor NOR2 (N1302, N1284, N574);
nor NOR3 (N1303, N1298, N203, N122);
or OR3 (N1304, N1299, N1082, N280);
buf BUF1 (N1305, N1294);
not NOT1 (N1306, N1290);
nor NOR2 (N1307, N1301, N703);
buf BUF1 (N1308, N1307);
and AND3 (N1309, N1308, N129, N707);
xor XOR2 (N1310, N1304, N307);
nand NAND3 (N1311, N1305, N516, N1055);
not NOT1 (N1312, N1311);
or OR4 (N1313, N1303, N1193, N252, N1237);
or OR4 (N1314, N1302, N1248, N1173, N517);
or OR2 (N1315, N1309, N1258);
nand NAND3 (N1316, N1312, N399, N481);
nand NAND2 (N1317, N1314, N259);
xor XOR2 (N1318, N1285, N995);
buf BUF1 (N1319, N1266);
and AND3 (N1320, N1317, N432, N1070);
and AND4 (N1321, N1300, N65, N360, N70);
nand NAND4 (N1322, N1310, N362, N1198, N138);
and AND2 (N1323, N1306, N326);
and AND4 (N1324, N1296, N590, N588, N461);
and AND4 (N1325, N1323, N592, N1324, N208);
nand NAND4 (N1326, N602, N1319, N363, N314);
and AND4 (N1327, N674, N487, N489, N513);
not NOT1 (N1328, N1320);
nand NAND2 (N1329, N1326, N994);
not NOT1 (N1330, N1321);
nand NAND3 (N1331, N1325, N769, N1009);
nor NOR2 (N1332, N1330, N840);
and AND3 (N1333, N1316, N1020, N1296);
and AND4 (N1334, N1318, N175, N688, N756);
and AND3 (N1335, N1313, N15, N1053);
xor XOR2 (N1336, N1331, N624);
nor NOR4 (N1337, N1335, N172, N256, N1120);
nand NAND2 (N1338, N1333, N1147);
xor XOR2 (N1339, N1336, N65);
or OR3 (N1340, N1327, N1326, N688);
nand NAND4 (N1341, N1338, N1053, N321, N1272);
and AND2 (N1342, N1337, N66);
xor XOR2 (N1343, N1332, N979);
xor XOR2 (N1344, N1343, N66);
buf BUF1 (N1345, N1322);
or OR2 (N1346, N1334, N178);
buf BUF1 (N1347, N1344);
not NOT1 (N1348, N1329);
nor NOR3 (N1349, N1341, N1244, N113);
nor NOR4 (N1350, N1328, N1327, N402, N509);
nand NAND4 (N1351, N1339, N861, N484, N1134);
and AND4 (N1352, N1346, N1302, N347, N1098);
not NOT1 (N1353, N1315);
buf BUF1 (N1354, N1353);
nor NOR4 (N1355, N1354, N1328, N610, N1218);
xor XOR2 (N1356, N1340, N976);
buf BUF1 (N1357, N1356);
not NOT1 (N1358, N1351);
or OR3 (N1359, N1348, N239, N353);
buf BUF1 (N1360, N1359);
nand NAND3 (N1361, N1360, N1288, N478);
nor NOR2 (N1362, N1357, N853);
or OR3 (N1363, N1358, N135, N1270);
or OR4 (N1364, N1352, N558, N1094, N491);
or OR4 (N1365, N1355, N875, N417, N1131);
buf BUF1 (N1366, N1361);
nor NOR4 (N1367, N1362, N606, N633, N510);
nand NAND3 (N1368, N1366, N256, N420);
and AND3 (N1369, N1367, N735, N693);
not NOT1 (N1370, N1342);
nand NAND2 (N1371, N1370, N846);
and AND3 (N1372, N1368, N142, N658);
not NOT1 (N1373, N1369);
and AND4 (N1374, N1373, N131, N1130, N1039);
not NOT1 (N1375, N1364);
not NOT1 (N1376, N1349);
or OR2 (N1377, N1347, N311);
not NOT1 (N1378, N1350);
or OR4 (N1379, N1372, N1219, N597, N55);
nand NAND4 (N1380, N1371, N686, N1073, N1242);
buf BUF1 (N1381, N1376);
nand NAND2 (N1382, N1378, N1129);
xor XOR2 (N1383, N1379, N940);
and AND3 (N1384, N1381, N867, N1080);
xor XOR2 (N1385, N1345, N1240);
nand NAND2 (N1386, N1374, N740);
buf BUF1 (N1387, N1377);
not NOT1 (N1388, N1363);
nor NOR2 (N1389, N1385, N542);
or OR4 (N1390, N1386, N676, N500, N168);
not NOT1 (N1391, N1365);
buf BUF1 (N1392, N1387);
nor NOR3 (N1393, N1391, N1342, N150);
xor XOR2 (N1394, N1390, N385);
or OR3 (N1395, N1392, N844, N719);
nand NAND4 (N1396, N1382, N1295, N826, N152);
or OR3 (N1397, N1394, N27, N970);
xor XOR2 (N1398, N1393, N371);
nand NAND4 (N1399, N1398, N912, N750, N249);
xor XOR2 (N1400, N1375, N562);
nand NAND2 (N1401, N1400, N9);
not NOT1 (N1402, N1395);
not NOT1 (N1403, N1380);
nor NOR3 (N1404, N1401, N1268, N1388);
not NOT1 (N1405, N573);
and AND2 (N1406, N1402, N49);
and AND2 (N1407, N1397, N1285);
nor NOR4 (N1408, N1383, N914, N1370, N855);
or OR2 (N1409, N1403, N338);
buf BUF1 (N1410, N1409);
and AND2 (N1411, N1399, N540);
xor XOR2 (N1412, N1410, N786);
nand NAND2 (N1413, N1396, N489);
and AND4 (N1414, N1384, N510, N1222, N462);
xor XOR2 (N1415, N1413, N335);
buf BUF1 (N1416, N1389);
xor XOR2 (N1417, N1405, N948);
and AND2 (N1418, N1412, N886);
and AND2 (N1419, N1404, N931);
buf BUF1 (N1420, N1406);
nand NAND2 (N1421, N1414, N155);
xor XOR2 (N1422, N1421, N118);
not NOT1 (N1423, N1418);
not NOT1 (N1424, N1422);
and AND4 (N1425, N1407, N359, N1021, N900);
buf BUF1 (N1426, N1423);
and AND2 (N1427, N1424, N239);
and AND3 (N1428, N1426, N64, N1370);
or OR2 (N1429, N1417, N1409);
and AND4 (N1430, N1415, N497, N773, N500);
nand NAND4 (N1431, N1427, N817, N965, N484);
nand NAND2 (N1432, N1428, N949);
buf BUF1 (N1433, N1419);
buf BUF1 (N1434, N1432);
nor NOR3 (N1435, N1408, N939, N294);
xor XOR2 (N1436, N1416, N517);
not NOT1 (N1437, N1411);
not NOT1 (N1438, N1435);
xor XOR2 (N1439, N1437, N711);
nand NAND3 (N1440, N1433, N628, N936);
or OR2 (N1441, N1431, N1061);
and AND3 (N1442, N1439, N70, N153);
nand NAND2 (N1443, N1438, N272);
not NOT1 (N1444, N1434);
not NOT1 (N1445, N1420);
or OR3 (N1446, N1425, N268, N1343);
nor NOR4 (N1447, N1443, N280, N825, N993);
or OR4 (N1448, N1447, N969, N1110, N287);
or OR4 (N1449, N1429, N1310, N1135, N1174);
or OR4 (N1450, N1442, N925, N323, N1047);
and AND2 (N1451, N1436, N1145);
and AND3 (N1452, N1445, N84, N70);
xor XOR2 (N1453, N1449, N746);
nor NOR2 (N1454, N1448, N1273);
nand NAND2 (N1455, N1430, N159);
xor XOR2 (N1456, N1444, N783);
buf BUF1 (N1457, N1446);
nand NAND4 (N1458, N1456, N890, N901, N378);
nor NOR3 (N1459, N1451, N762, N554);
and AND3 (N1460, N1455, N97, N499);
not NOT1 (N1461, N1454);
nor NOR2 (N1462, N1440, N787);
xor XOR2 (N1463, N1457, N1234);
buf BUF1 (N1464, N1452);
and AND3 (N1465, N1463, N476, N405);
xor XOR2 (N1466, N1450, N90);
nor NOR3 (N1467, N1466, N176, N754);
nor NOR2 (N1468, N1465, N523);
and AND4 (N1469, N1462, N112, N625, N1248);
buf BUF1 (N1470, N1441);
nor NOR2 (N1471, N1453, N1230);
xor XOR2 (N1472, N1460, N722);
or OR4 (N1473, N1469, N1187, N231, N772);
buf BUF1 (N1474, N1459);
and AND2 (N1475, N1467, N1228);
not NOT1 (N1476, N1473);
and AND4 (N1477, N1468, N1217, N74, N780);
not NOT1 (N1478, N1464);
nand NAND3 (N1479, N1476, N334, N225);
nand NAND2 (N1480, N1458, N441);
buf BUF1 (N1481, N1480);
and AND4 (N1482, N1475, N327, N94, N1315);
nor NOR4 (N1483, N1482, N669, N832, N1134);
and AND4 (N1484, N1472, N222, N924, N789);
buf BUF1 (N1485, N1470);
nand NAND4 (N1486, N1478, N859, N1153, N1023);
or OR4 (N1487, N1477, N381, N1061, N1257);
nor NOR4 (N1488, N1461, N681, N21, N3);
or OR4 (N1489, N1479, N283, N430, N850);
xor XOR2 (N1490, N1471, N322);
xor XOR2 (N1491, N1486, N911);
buf BUF1 (N1492, N1490);
nand NAND3 (N1493, N1484, N1006, N836);
buf BUF1 (N1494, N1485);
not NOT1 (N1495, N1474);
or OR4 (N1496, N1491, N1009, N1450, N1309);
buf BUF1 (N1497, N1481);
or OR4 (N1498, N1493, N1255, N650, N655);
xor XOR2 (N1499, N1487, N1441);
or OR2 (N1500, N1483, N635);
not NOT1 (N1501, N1496);
or OR4 (N1502, N1488, N765, N360, N957);
or OR3 (N1503, N1499, N353, N1247);
nand NAND4 (N1504, N1500, N1088, N737, N766);
xor XOR2 (N1505, N1489, N1046);
and AND4 (N1506, N1503, N890, N66, N335);
buf BUF1 (N1507, N1497);
nor NOR3 (N1508, N1507, N515, N785);
not NOT1 (N1509, N1501);
nor NOR4 (N1510, N1508, N749, N319, N133);
nor NOR2 (N1511, N1506, N163);
or OR3 (N1512, N1505, N648, N1331);
not NOT1 (N1513, N1492);
nor NOR3 (N1514, N1511, N239, N1042);
nor NOR2 (N1515, N1510, N473);
xor XOR2 (N1516, N1515, N501);
nand NAND2 (N1517, N1498, N498);
buf BUF1 (N1518, N1502);
xor XOR2 (N1519, N1518, N1227);
or OR3 (N1520, N1516, N1263, N566);
and AND4 (N1521, N1514, N151, N1212, N198);
buf BUF1 (N1522, N1512);
or OR3 (N1523, N1520, N1027, N613);
nor NOR2 (N1524, N1494, N1109);
xor XOR2 (N1525, N1523, N1188);
buf BUF1 (N1526, N1513);
not NOT1 (N1527, N1526);
buf BUF1 (N1528, N1504);
not NOT1 (N1529, N1522);
nor NOR4 (N1530, N1509, N844, N234, N1474);
and AND2 (N1531, N1530, N1158);
not NOT1 (N1532, N1495);
not NOT1 (N1533, N1527);
and AND4 (N1534, N1528, N629, N182, N292);
nand NAND3 (N1535, N1529, N377, N749);
buf BUF1 (N1536, N1525);
buf BUF1 (N1537, N1517);
buf BUF1 (N1538, N1536);
or OR4 (N1539, N1524, N199, N1518, N1176);
nor NOR4 (N1540, N1538, N885, N977, N1427);
buf BUF1 (N1541, N1537);
or OR2 (N1542, N1540, N879);
xor XOR2 (N1543, N1521, N1239);
nand NAND3 (N1544, N1542, N731, N497);
xor XOR2 (N1545, N1534, N703);
and AND3 (N1546, N1531, N1300, N1071);
not NOT1 (N1547, N1545);
buf BUF1 (N1548, N1543);
and AND4 (N1549, N1548, N586, N602, N1513);
nand NAND4 (N1550, N1533, N991, N308, N1492);
xor XOR2 (N1551, N1519, N1511);
xor XOR2 (N1552, N1535, N486);
and AND4 (N1553, N1544, N84, N1087, N722);
and AND4 (N1554, N1549, N1343, N1201, N595);
not NOT1 (N1555, N1532);
not NOT1 (N1556, N1541);
nor NOR2 (N1557, N1551, N208);
buf BUF1 (N1558, N1547);
or OR4 (N1559, N1550, N287, N79, N1555);
or OR2 (N1560, N1206, N1272);
or OR2 (N1561, N1554, N666);
nand NAND2 (N1562, N1539, N331);
nand NAND3 (N1563, N1561, N714, N1393);
and AND2 (N1564, N1558, N1135);
nor NOR4 (N1565, N1552, N640, N441, N1006);
nor NOR3 (N1566, N1564, N1182, N1365);
buf BUF1 (N1567, N1559);
or OR3 (N1568, N1565, N800, N1453);
and AND2 (N1569, N1562, N1491);
xor XOR2 (N1570, N1568, N583);
not NOT1 (N1571, N1566);
buf BUF1 (N1572, N1569);
or OR2 (N1573, N1560, N1300);
and AND4 (N1574, N1573, N879, N785, N668);
and AND2 (N1575, N1574, N912);
or OR2 (N1576, N1572, N1510);
nand NAND3 (N1577, N1571, N1040, N784);
not NOT1 (N1578, N1575);
nor NOR2 (N1579, N1553, N1020);
nand NAND3 (N1580, N1579, N478, N1091);
buf BUF1 (N1581, N1546);
nand NAND2 (N1582, N1557, N1518);
or OR4 (N1583, N1556, N1122, N1287, N533);
xor XOR2 (N1584, N1581, N133);
not NOT1 (N1585, N1582);
or OR3 (N1586, N1577, N1554, N1544);
or OR2 (N1587, N1576, N1177);
buf BUF1 (N1588, N1583);
nand NAND3 (N1589, N1584, N1424, N1403);
and AND2 (N1590, N1563, N603);
nand NAND3 (N1591, N1586, N146, N436);
not NOT1 (N1592, N1578);
or OR4 (N1593, N1570, N1273, N1400, N1378);
nor NOR2 (N1594, N1580, N1068);
and AND2 (N1595, N1594, N136);
nand NAND2 (N1596, N1588, N1529);
xor XOR2 (N1597, N1589, N1528);
buf BUF1 (N1598, N1597);
nor NOR3 (N1599, N1585, N795, N1328);
or OR4 (N1600, N1595, N832, N1106, N261);
nor NOR3 (N1601, N1590, N441, N1273);
xor XOR2 (N1602, N1598, N1507);
nor NOR2 (N1603, N1592, N623);
and AND2 (N1604, N1601, N190);
and AND4 (N1605, N1596, N614, N17, N1509);
buf BUF1 (N1606, N1593);
not NOT1 (N1607, N1604);
not NOT1 (N1608, N1606);
and AND4 (N1609, N1605, N252, N857, N586);
buf BUF1 (N1610, N1600);
nand NAND2 (N1611, N1610, N327);
nor NOR2 (N1612, N1587, N1538);
nor NOR4 (N1613, N1612, N1226, N755, N1335);
not NOT1 (N1614, N1599);
or OR2 (N1615, N1609, N1052);
not NOT1 (N1616, N1607);
and AND4 (N1617, N1603, N1553, N948, N1497);
nand NAND2 (N1618, N1608, N1550);
buf BUF1 (N1619, N1591);
and AND3 (N1620, N1618, N1447, N812);
buf BUF1 (N1621, N1615);
xor XOR2 (N1622, N1602, N1071);
nand NAND3 (N1623, N1613, N1030, N476);
or OR4 (N1624, N1567, N1417, N1335, N746);
nor NOR3 (N1625, N1616, N872, N1505);
buf BUF1 (N1626, N1621);
nor NOR2 (N1627, N1625, N1230);
xor XOR2 (N1628, N1614, N1126);
xor XOR2 (N1629, N1626, N1273);
xor XOR2 (N1630, N1627, N432);
nor NOR2 (N1631, N1622, N206);
and AND3 (N1632, N1611, N158, N423);
or OR3 (N1633, N1628, N43, N157);
or OR3 (N1634, N1624, N128, N1626);
not NOT1 (N1635, N1620);
buf BUF1 (N1636, N1633);
nor NOR3 (N1637, N1631, N1459, N805);
nor NOR3 (N1638, N1617, N762, N969);
not NOT1 (N1639, N1637);
or OR2 (N1640, N1632, N582);
nand NAND2 (N1641, N1634, N342);
buf BUF1 (N1642, N1639);
not NOT1 (N1643, N1638);
or OR3 (N1644, N1619, N747, N1589);
buf BUF1 (N1645, N1641);
buf BUF1 (N1646, N1630);
nand NAND4 (N1647, N1642, N250, N1356, N1232);
not NOT1 (N1648, N1643);
xor XOR2 (N1649, N1644, N1090);
nand NAND3 (N1650, N1646, N74, N1106);
not NOT1 (N1651, N1649);
buf BUF1 (N1652, N1645);
nor NOR3 (N1653, N1651, N1495, N821);
buf BUF1 (N1654, N1652);
xor XOR2 (N1655, N1629, N1245);
and AND3 (N1656, N1655, N672, N1068);
or OR4 (N1657, N1656, N413, N941, N191);
nand NAND3 (N1658, N1657, N1230, N719);
or OR3 (N1659, N1640, N965, N322);
and AND4 (N1660, N1647, N1567, N719, N1507);
buf BUF1 (N1661, N1659);
nand NAND4 (N1662, N1653, N390, N139, N1647);
nor NOR3 (N1663, N1661, N435, N1104);
or OR3 (N1664, N1662, N1275, N91);
buf BUF1 (N1665, N1648);
nor NOR4 (N1666, N1623, N809, N793, N1221);
nor NOR4 (N1667, N1665, N496, N944, N1493);
xor XOR2 (N1668, N1666, N1122);
or OR4 (N1669, N1636, N900, N1585, N708);
and AND2 (N1670, N1650, N470);
nand NAND4 (N1671, N1658, N20, N438, N201);
and AND4 (N1672, N1654, N1180, N358, N1600);
buf BUF1 (N1673, N1670);
nor NOR4 (N1674, N1672, N401, N481, N449);
not NOT1 (N1675, N1673);
not NOT1 (N1676, N1671);
buf BUF1 (N1677, N1676);
and AND2 (N1678, N1675, N247);
or OR3 (N1679, N1667, N796, N1110);
nand NAND4 (N1680, N1674, N1345, N1403, N1174);
nor NOR4 (N1681, N1663, N186, N1126, N1234);
and AND4 (N1682, N1678, N1240, N779, N184);
nor NOR3 (N1683, N1682, N768, N41);
or OR4 (N1684, N1668, N795, N546, N1408);
not NOT1 (N1685, N1680);
nand NAND2 (N1686, N1664, N572);
or OR3 (N1687, N1679, N642, N337);
and AND4 (N1688, N1685, N1106, N535, N1162);
xor XOR2 (N1689, N1688, N44);
nand NAND2 (N1690, N1677, N483);
not NOT1 (N1691, N1635);
not NOT1 (N1692, N1690);
buf BUF1 (N1693, N1660);
nor NOR2 (N1694, N1689, N160);
nor NOR2 (N1695, N1684, N569);
nor NOR4 (N1696, N1683, N1131, N405, N706);
xor XOR2 (N1697, N1687, N683);
nand NAND3 (N1698, N1694, N736, N1653);
buf BUF1 (N1699, N1691);
xor XOR2 (N1700, N1699, N147);
nand NAND3 (N1701, N1695, N921, N146);
not NOT1 (N1702, N1681);
or OR3 (N1703, N1692, N1165, N935);
or OR2 (N1704, N1669, N221);
xor XOR2 (N1705, N1698, N1093);
xor XOR2 (N1706, N1693, N704);
buf BUF1 (N1707, N1701);
not NOT1 (N1708, N1704);
and AND4 (N1709, N1703, N840, N1278, N1002);
not NOT1 (N1710, N1708);
and AND3 (N1711, N1696, N419, N922);
not NOT1 (N1712, N1711);
nor NOR4 (N1713, N1707, N405, N347, N1086);
and AND2 (N1714, N1706, N1637);
and AND4 (N1715, N1709, N1173, N1526, N289);
buf BUF1 (N1716, N1686);
not NOT1 (N1717, N1702);
or OR2 (N1718, N1716, N496);
or OR2 (N1719, N1714, N111);
and AND4 (N1720, N1715, N834, N923, N72);
and AND3 (N1721, N1710, N524, N140);
and AND2 (N1722, N1720, N1425);
nand NAND2 (N1723, N1705, N300);
and AND2 (N1724, N1712, N1209);
or OR3 (N1725, N1721, N1520, N415);
not NOT1 (N1726, N1718);
or OR3 (N1727, N1717, N1388, N1028);
not NOT1 (N1728, N1726);
xor XOR2 (N1729, N1723, N1633);
or OR3 (N1730, N1719, N315, N1290);
and AND4 (N1731, N1724, N1652, N437, N1347);
nand NAND3 (N1732, N1725, N842, N1721);
buf BUF1 (N1733, N1697);
and AND4 (N1734, N1731, N713, N1642, N111);
nor NOR4 (N1735, N1700, N952, N4, N1034);
or OR2 (N1736, N1733, N1030);
nor NOR3 (N1737, N1730, N1336, N92);
nand NAND2 (N1738, N1727, N487);
and AND3 (N1739, N1737, N945, N1556);
and AND3 (N1740, N1729, N1204, N683);
not NOT1 (N1741, N1740);
or OR4 (N1742, N1728, N478, N1255, N971);
nor NOR4 (N1743, N1739, N1437, N1652, N1094);
nand NAND3 (N1744, N1738, N1002, N1533);
not NOT1 (N1745, N1743);
and AND2 (N1746, N1741, N566);
and AND2 (N1747, N1735, N1071);
nor NOR2 (N1748, N1742, N1295);
and AND2 (N1749, N1736, N379);
nor NOR2 (N1750, N1744, N1560);
or OR4 (N1751, N1745, N668, N1652, N1473);
xor XOR2 (N1752, N1751, N1147);
nor NOR3 (N1753, N1750, N1115, N395);
xor XOR2 (N1754, N1734, N423);
nor NOR2 (N1755, N1753, N802);
or OR3 (N1756, N1748, N1005, N321);
buf BUF1 (N1757, N1732);
and AND4 (N1758, N1746, N1253, N1579, N1276);
and AND2 (N1759, N1747, N993);
buf BUF1 (N1760, N1749);
nand NAND3 (N1761, N1759, N1159, N844);
buf BUF1 (N1762, N1755);
or OR2 (N1763, N1722, N1526);
or OR3 (N1764, N1761, N220, N597);
not NOT1 (N1765, N1763);
or OR4 (N1766, N1754, N795, N211, N1621);
nand NAND3 (N1767, N1762, N1691, N379);
xor XOR2 (N1768, N1764, N184);
not NOT1 (N1769, N1760);
or OR3 (N1770, N1767, N748, N379);
not NOT1 (N1771, N1765);
and AND3 (N1772, N1756, N1708, N1136);
xor XOR2 (N1773, N1770, N1695);
and AND2 (N1774, N1713, N372);
nand NAND2 (N1775, N1773, N665);
not NOT1 (N1776, N1757);
xor XOR2 (N1777, N1775, N1123);
nand NAND2 (N1778, N1777, N1103);
buf BUF1 (N1779, N1776);
or OR2 (N1780, N1779, N840);
and AND4 (N1781, N1768, N1706, N424, N970);
nor NOR4 (N1782, N1774, N1023, N1573, N1335);
nand NAND4 (N1783, N1778, N288, N1073, N1462);
not NOT1 (N1784, N1772);
or OR2 (N1785, N1769, N1591);
not NOT1 (N1786, N1783);
not NOT1 (N1787, N1771);
buf BUF1 (N1788, N1780);
and AND3 (N1789, N1752, N1764, N674);
and AND4 (N1790, N1758, N1616, N1686, N1071);
nor NOR2 (N1791, N1786, N876);
not NOT1 (N1792, N1788);
not NOT1 (N1793, N1781);
not NOT1 (N1794, N1792);
xor XOR2 (N1795, N1791, N1549);
xor XOR2 (N1796, N1782, N1728);
nor NOR2 (N1797, N1784, N174);
nand NAND4 (N1798, N1794, N1459, N546, N645);
buf BUF1 (N1799, N1790);
xor XOR2 (N1800, N1785, N64);
nor NOR4 (N1801, N1800, N508, N1251, N1767);
xor XOR2 (N1802, N1793, N28);
xor XOR2 (N1803, N1789, N74);
not NOT1 (N1804, N1801);
xor XOR2 (N1805, N1796, N852);
xor XOR2 (N1806, N1803, N1704);
and AND3 (N1807, N1804, N333, N1013);
nor NOR2 (N1808, N1806, N1738);
buf BUF1 (N1809, N1802);
xor XOR2 (N1810, N1766, N619);
not NOT1 (N1811, N1807);
nand NAND3 (N1812, N1798, N1635, N1355);
xor XOR2 (N1813, N1810, N584);
xor XOR2 (N1814, N1811, N920);
not NOT1 (N1815, N1809);
buf BUF1 (N1816, N1799);
and AND4 (N1817, N1812, N320, N1758, N782);
not NOT1 (N1818, N1817);
buf BUF1 (N1819, N1815);
and AND4 (N1820, N1797, N1272, N339, N60);
not NOT1 (N1821, N1820);
buf BUF1 (N1822, N1816);
nor NOR3 (N1823, N1813, N996, N1495);
nor NOR4 (N1824, N1819, N1044, N523, N522);
nor NOR4 (N1825, N1787, N1773, N23, N348);
nor NOR4 (N1826, N1805, N793, N732, N405);
nand NAND2 (N1827, N1825, N1478);
nand NAND4 (N1828, N1826, N1184, N470, N536);
xor XOR2 (N1829, N1823, N1493);
xor XOR2 (N1830, N1822, N1419);
and AND3 (N1831, N1830, N284, N574);
not NOT1 (N1832, N1808);
and AND4 (N1833, N1832, N1061, N1059, N520);
and AND3 (N1834, N1828, N869, N596);
nand NAND2 (N1835, N1821, N967);
buf BUF1 (N1836, N1795);
buf BUF1 (N1837, N1824);
nor NOR2 (N1838, N1833, N160);
or OR3 (N1839, N1835, N1529, N144);
buf BUF1 (N1840, N1834);
xor XOR2 (N1841, N1831, N797);
or OR2 (N1842, N1827, N1554);
nor NOR2 (N1843, N1840, N803);
not NOT1 (N1844, N1837);
nor NOR4 (N1845, N1829, N427, N1599, N1119);
xor XOR2 (N1846, N1842, N976);
or OR2 (N1847, N1843, N1205);
nor NOR2 (N1848, N1839, N188);
or OR2 (N1849, N1841, N1205);
not NOT1 (N1850, N1818);
not NOT1 (N1851, N1838);
and AND2 (N1852, N1814, N245);
buf BUF1 (N1853, N1846);
nor NOR4 (N1854, N1849, N1265, N866, N1171);
buf BUF1 (N1855, N1850);
nand NAND2 (N1856, N1847, N146);
not NOT1 (N1857, N1836);
xor XOR2 (N1858, N1852, N169);
nand NAND2 (N1859, N1845, N1610);
xor XOR2 (N1860, N1858, N1205);
and AND2 (N1861, N1856, N843);
not NOT1 (N1862, N1848);
not NOT1 (N1863, N1860);
and AND3 (N1864, N1853, N1423, N1079);
not NOT1 (N1865, N1863);
or OR3 (N1866, N1862, N1310, N383);
xor XOR2 (N1867, N1865, N1373);
xor XOR2 (N1868, N1867, N244);
nand NAND2 (N1869, N1861, N763);
nor NOR3 (N1870, N1864, N68, N1398);
nand NAND4 (N1871, N1869, N362, N1377, N308);
nor NOR3 (N1872, N1855, N1741, N352);
buf BUF1 (N1873, N1844);
not NOT1 (N1874, N1868);
xor XOR2 (N1875, N1873, N791);
and AND2 (N1876, N1854, N1153);
xor XOR2 (N1877, N1870, N669);
and AND2 (N1878, N1876, N231);
nand NAND2 (N1879, N1866, N40);
nand NAND4 (N1880, N1872, N271, N1415, N291);
nor NOR3 (N1881, N1880, N95, N1542);
buf BUF1 (N1882, N1857);
nand NAND2 (N1883, N1878, N1635);
nor NOR3 (N1884, N1871, N1876, N964);
nor NOR3 (N1885, N1882, N1414, N270);
nor NOR3 (N1886, N1875, N1413, N464);
or OR3 (N1887, N1885, N523, N467);
nor NOR4 (N1888, N1874, N518, N1220, N1391);
xor XOR2 (N1889, N1879, N1166);
or OR4 (N1890, N1859, N1293, N71, N1183);
not NOT1 (N1891, N1887);
xor XOR2 (N1892, N1888, N1718);
or OR4 (N1893, N1886, N290, N522, N352);
nor NOR4 (N1894, N1893, N1358, N263, N1032);
and AND3 (N1895, N1881, N1496, N1722);
not NOT1 (N1896, N1884);
buf BUF1 (N1897, N1894);
buf BUF1 (N1898, N1877);
and AND2 (N1899, N1895, N1175);
nand NAND3 (N1900, N1891, N1740, N458);
or OR2 (N1901, N1900, N677);
and AND3 (N1902, N1899, N1898, N684);
not NOT1 (N1903, N1444);
nor NOR3 (N1904, N1902, N748, N412);
or OR4 (N1905, N1904, N626, N511, N624);
not NOT1 (N1906, N1883);
nor NOR2 (N1907, N1851, N1154);
xor XOR2 (N1908, N1901, N231);
nand NAND4 (N1909, N1896, N457, N1403, N303);
or OR2 (N1910, N1906, N27);
nand NAND2 (N1911, N1905, N1789);
or OR3 (N1912, N1892, N831, N1452);
or OR2 (N1913, N1889, N602);
xor XOR2 (N1914, N1909, N1421);
xor XOR2 (N1915, N1911, N1564);
or OR3 (N1916, N1910, N765, N1469);
or OR2 (N1917, N1912, N1317);
or OR2 (N1918, N1908, N869);
and AND2 (N1919, N1897, N807);
nand NAND2 (N1920, N1917, N642);
nand NAND4 (N1921, N1907, N1740, N400, N343);
not NOT1 (N1922, N1918);
and AND4 (N1923, N1921, N596, N1117, N1061);
xor XOR2 (N1924, N1923, N250);
or OR3 (N1925, N1890, N14, N1886);
nand NAND2 (N1926, N1922, N162);
nor NOR3 (N1927, N1915, N835, N947);
or OR2 (N1928, N1920, N1820);
buf BUF1 (N1929, N1924);
nor NOR4 (N1930, N1916, N1316, N1644, N496);
buf BUF1 (N1931, N1903);
not NOT1 (N1932, N1927);
nand NAND3 (N1933, N1926, N737, N153);
or OR2 (N1934, N1928, N1661);
nor NOR3 (N1935, N1934, N1047, N546);
not NOT1 (N1936, N1919);
nand NAND3 (N1937, N1935, N1469, N1613);
and AND3 (N1938, N1929, N527, N118);
or OR3 (N1939, N1932, N1769, N1574);
buf BUF1 (N1940, N1913);
and AND4 (N1941, N1931, N1552, N1289, N1635);
buf BUF1 (N1942, N1933);
nor NOR4 (N1943, N1939, N1324, N1054, N115);
and AND3 (N1944, N1941, N822, N1291);
buf BUF1 (N1945, N1944);
and AND2 (N1946, N1930, N748);
not NOT1 (N1947, N1936);
nor NOR4 (N1948, N1938, N1838, N1456, N338);
xor XOR2 (N1949, N1947, N591);
nor NOR4 (N1950, N1945, N217, N476, N38);
buf BUF1 (N1951, N1948);
and AND2 (N1952, N1937, N612);
not NOT1 (N1953, N1914);
not NOT1 (N1954, N1925);
not NOT1 (N1955, N1951);
nor NOR3 (N1956, N1942, N9, N659);
nor NOR2 (N1957, N1946, N96);
nor NOR3 (N1958, N1957, N1661, N1143);
nand NAND3 (N1959, N1950, N494, N1795);
nand NAND3 (N1960, N1949, N1368, N737);
buf BUF1 (N1961, N1960);
nand NAND2 (N1962, N1956, N1850);
xor XOR2 (N1963, N1952, N809);
or OR2 (N1964, N1943, N1732);
or OR3 (N1965, N1954, N1209, N1783);
nand NAND4 (N1966, N1961, N494, N1387, N979);
and AND4 (N1967, N1963, N1513, N1035, N1210);
not NOT1 (N1968, N1965);
buf BUF1 (N1969, N1964);
nand NAND3 (N1970, N1953, N1059, N1236);
buf BUF1 (N1971, N1962);
not NOT1 (N1972, N1968);
or OR2 (N1973, N1955, N1710);
and AND2 (N1974, N1959, N194);
or OR3 (N1975, N1967, N787, N805);
not NOT1 (N1976, N1970);
not NOT1 (N1977, N1940);
or OR4 (N1978, N1971, N407, N694, N1022);
nand NAND3 (N1979, N1958, N1082, N75);
xor XOR2 (N1980, N1974, N1346);
or OR4 (N1981, N1979, N1890, N1572, N834);
nand NAND2 (N1982, N1981, N1521);
xor XOR2 (N1983, N1982, N251);
or OR2 (N1984, N1980, N1872);
and AND3 (N1985, N1973, N1872, N886);
or OR4 (N1986, N1972, N695, N1551, N1631);
buf BUF1 (N1987, N1986);
xor XOR2 (N1988, N1975, N669);
nand NAND2 (N1989, N1977, N1818);
or OR4 (N1990, N1984, N1720, N596, N1681);
buf BUF1 (N1991, N1985);
buf BUF1 (N1992, N1991);
nand NAND2 (N1993, N1988, N1779);
xor XOR2 (N1994, N1976, N1885);
nand NAND4 (N1995, N1989, N1109, N1547, N1752);
xor XOR2 (N1996, N1990, N1899);
xor XOR2 (N1997, N1969, N1913);
buf BUF1 (N1998, N1997);
buf BUF1 (N1999, N1987);
or OR2 (N2000, N1992, N619);
xor XOR2 (N2001, N1998, N505);
nand NAND2 (N2002, N2001, N954);
not NOT1 (N2003, N1995);
not NOT1 (N2004, N1999);
and AND3 (N2005, N2003, N175, N706);
buf BUF1 (N2006, N2005);
or OR3 (N2007, N1978, N1055, N385);
and AND3 (N2008, N2006, N1511, N810);
not NOT1 (N2009, N2007);
and AND3 (N2010, N2009, N509, N383);
nand NAND4 (N2011, N1994, N1156, N960, N133);
nand NAND2 (N2012, N2010, N549);
and AND4 (N2013, N2004, N567, N172, N1438);
and AND4 (N2014, N2012, N1235, N311, N120);
xor XOR2 (N2015, N2013, N327);
and AND3 (N2016, N2015, N1528, N1703);
not NOT1 (N2017, N1996);
nand NAND2 (N2018, N2008, N117);
nand NAND3 (N2019, N1993, N877, N1715);
and AND4 (N2020, N2002, N1431, N1545, N471);
buf BUF1 (N2021, N2019);
xor XOR2 (N2022, N2011, N624);
buf BUF1 (N2023, N2020);
not NOT1 (N2024, N2014);
xor XOR2 (N2025, N1966, N1893);
nand NAND2 (N2026, N2016, N45);
xor XOR2 (N2027, N1983, N1942);
or OR3 (N2028, N2021, N848, N152);
xor XOR2 (N2029, N2022, N242);
and AND4 (N2030, N2017, N1814, N750, N1818);
buf BUF1 (N2031, N2024);
nor NOR2 (N2032, N2018, N1725);
not NOT1 (N2033, N2030);
nor NOR2 (N2034, N2029, N324);
and AND3 (N2035, N2026, N1543, N1927);
nand NAND4 (N2036, N2023, N444, N1766, N1715);
buf BUF1 (N2037, N2031);
xor XOR2 (N2038, N2027, N1743);
and AND2 (N2039, N2025, N693);
nand NAND4 (N2040, N2038, N191, N1328, N682);
and AND3 (N2041, N2035, N1408, N1623);
not NOT1 (N2042, N2028);
not NOT1 (N2043, N2039);
buf BUF1 (N2044, N2041);
xor XOR2 (N2045, N2043, N1253);
buf BUF1 (N2046, N2045);
or OR2 (N2047, N2034, N346);
buf BUF1 (N2048, N2040);
nand NAND4 (N2049, N2032, N690, N1466, N31);
nor NOR3 (N2050, N2048, N764, N14);
or OR4 (N2051, N2042, N1605, N1028, N1058);
not NOT1 (N2052, N2049);
xor XOR2 (N2053, N2046, N692);
buf BUF1 (N2054, N2037);
xor XOR2 (N2055, N2033, N1533);
buf BUF1 (N2056, N2054);
or OR3 (N2057, N2056, N1122, N1309);
nand NAND4 (N2058, N2057, N566, N624, N173);
nand NAND3 (N2059, N2055, N1176, N522);
nand NAND3 (N2060, N2059, N1101, N684);
xor XOR2 (N2061, N2060, N1195);
buf BUF1 (N2062, N2051);
and AND3 (N2063, N2044, N585, N728);
xor XOR2 (N2064, N2050, N1310);
xor XOR2 (N2065, N2058, N1808);
xor XOR2 (N2066, N2036, N1383);
and AND3 (N2067, N2063, N66, N1022);
nor NOR2 (N2068, N2066, N286);
and AND4 (N2069, N2062, N910, N1851, N467);
or OR4 (N2070, N2068, N31, N748, N1128);
and AND4 (N2071, N2070, N1416, N1396, N1573);
not NOT1 (N2072, N2065);
buf BUF1 (N2073, N2072);
nor NOR4 (N2074, N2069, N1917, N2000, N565);
or OR3 (N2075, N1536, N2034, N1131);
xor XOR2 (N2076, N2075, N545);
nand NAND4 (N2077, N2061, N197, N871, N1016);
or OR2 (N2078, N2052, N1902);
xor XOR2 (N2079, N2076, N229);
and AND3 (N2080, N2074, N1631, N2004);
not NOT1 (N2081, N2078);
nand NAND2 (N2082, N2064, N1503);
xor XOR2 (N2083, N2081, N197);
xor XOR2 (N2084, N2071, N671);
buf BUF1 (N2085, N2079);
and AND2 (N2086, N2077, N1163);
xor XOR2 (N2087, N2073, N1841);
nor NOR4 (N2088, N2080, N1164, N780, N134);
not NOT1 (N2089, N2047);
buf BUF1 (N2090, N2087);
buf BUF1 (N2091, N2090);
or OR2 (N2092, N2088, N722);
nand NAND3 (N2093, N2089, N889, N464);
nand NAND4 (N2094, N2085, N745, N808, N936);
nand NAND4 (N2095, N2092, N1588, N1401, N1149);
xor XOR2 (N2096, N2095, N1197);
nand NAND2 (N2097, N2093, N1072);
nor NOR2 (N2098, N2083, N932);
nor NOR3 (N2099, N2098, N1847, N187);
and AND3 (N2100, N2082, N1970, N461);
nand NAND2 (N2101, N2091, N1149);
buf BUF1 (N2102, N2097);
xor XOR2 (N2103, N2096, N972);
and AND2 (N2104, N2053, N895);
xor XOR2 (N2105, N2102, N372);
nand NAND4 (N2106, N2067, N938, N1794, N1239);
or OR2 (N2107, N2094, N131);
or OR2 (N2108, N2101, N953);
nor NOR2 (N2109, N2105, N668);
or OR3 (N2110, N2099, N1319, N280);
not NOT1 (N2111, N2109);
xor XOR2 (N2112, N2110, N485);
and AND4 (N2113, N2106, N982, N1179, N637);
nand NAND3 (N2114, N2100, N1379, N1143);
and AND4 (N2115, N2084, N978, N1491, N1491);
not NOT1 (N2116, N2103);
or OR3 (N2117, N2104, N49, N1334);
and AND4 (N2118, N2111, N1019, N1214, N239);
nor NOR4 (N2119, N2116, N1175, N1998, N1223);
xor XOR2 (N2120, N2115, N494);
nand NAND2 (N2121, N2086, N740);
xor XOR2 (N2122, N2119, N2109);
nor NOR3 (N2123, N2118, N427, N872);
or OR2 (N2124, N2120, N352);
and AND3 (N2125, N2122, N1179, N1411);
nor NOR2 (N2126, N2124, N295);
nand NAND3 (N2127, N2123, N1203, N1677);
buf BUF1 (N2128, N2127);
nand NAND4 (N2129, N2117, N1705, N1369, N1377);
buf BUF1 (N2130, N2112);
nor NOR3 (N2131, N2107, N954, N484);
and AND3 (N2132, N2114, N697, N609);
buf BUF1 (N2133, N2125);
not NOT1 (N2134, N2132);
or OR3 (N2135, N2134, N694, N177);
xor XOR2 (N2136, N2121, N316);
not NOT1 (N2137, N2131);
buf BUF1 (N2138, N2137);
nor NOR2 (N2139, N2136, N1102);
or OR3 (N2140, N2126, N1504, N876);
nand NAND3 (N2141, N2135, N1783, N1203);
and AND2 (N2142, N2141, N1151);
and AND3 (N2143, N2139, N899, N1107);
xor XOR2 (N2144, N2142, N531);
nor NOR2 (N2145, N2133, N1241);
buf BUF1 (N2146, N2128);
not NOT1 (N2147, N2130);
and AND3 (N2148, N2146, N846, N1818);
and AND4 (N2149, N2147, N1081, N2053, N754);
or OR4 (N2150, N2145, N1553, N1443, N545);
buf BUF1 (N2151, N2113);
xor XOR2 (N2152, N2148, N1077);
or OR3 (N2153, N2129, N1485, N1101);
or OR3 (N2154, N2153, N424, N1256);
or OR4 (N2155, N2150, N1115, N1676, N1651);
or OR3 (N2156, N2151, N225, N892);
and AND3 (N2157, N2154, N1466, N2085);
and AND2 (N2158, N2155, N1360);
nand NAND3 (N2159, N2138, N1148, N133);
xor XOR2 (N2160, N2159, N1618);
buf BUF1 (N2161, N2140);
xor XOR2 (N2162, N2157, N924);
and AND2 (N2163, N2144, N1807);
and AND3 (N2164, N2161, N840, N1642);
nor NOR3 (N2165, N2143, N1935, N2059);
nand NAND4 (N2166, N2160, N764, N1176, N936);
nand NAND4 (N2167, N2166, N1001, N2103, N487);
buf BUF1 (N2168, N2162);
xor XOR2 (N2169, N2165, N650);
buf BUF1 (N2170, N2163);
and AND3 (N2171, N2152, N787, N353);
nor NOR3 (N2172, N2169, N1712, N1903);
buf BUF1 (N2173, N2168);
nor NOR3 (N2174, N2167, N1648, N167);
buf BUF1 (N2175, N2164);
or OR2 (N2176, N2108, N1098);
xor XOR2 (N2177, N2175, N894);
nand NAND2 (N2178, N2158, N630);
nand NAND3 (N2179, N2149, N833, N1527);
nand NAND2 (N2180, N2172, N1935);
not NOT1 (N2181, N2179);
buf BUF1 (N2182, N2170);
nand NAND4 (N2183, N2182, N2129, N1012, N2123);
or OR3 (N2184, N2178, N1141, N128);
nand NAND2 (N2185, N2171, N1709);
nor NOR4 (N2186, N2173, N2071, N2131, N140);
and AND2 (N2187, N2176, N1996);
not NOT1 (N2188, N2187);
buf BUF1 (N2189, N2185);
or OR3 (N2190, N2188, N1194, N977);
buf BUF1 (N2191, N2190);
and AND4 (N2192, N2184, N858, N154, N1216);
not NOT1 (N2193, N2186);
buf BUF1 (N2194, N2189);
xor XOR2 (N2195, N2181, N2065);
nor NOR4 (N2196, N2192, N660, N791, N1964);
buf BUF1 (N2197, N2194);
xor XOR2 (N2198, N2156, N1144);
not NOT1 (N2199, N2198);
nor NOR2 (N2200, N2199, N1504);
buf BUF1 (N2201, N2195);
nand NAND3 (N2202, N2196, N1316, N740);
nand NAND4 (N2203, N2200, N362, N1598, N2140);
buf BUF1 (N2204, N2177);
not NOT1 (N2205, N2204);
buf BUF1 (N2206, N2197);
and AND3 (N2207, N2201, N1794, N1417);
buf BUF1 (N2208, N2174);
and AND2 (N2209, N2183, N512);
nor NOR4 (N2210, N2206, N210, N147, N2055);
or OR3 (N2211, N2193, N389, N1503);
buf BUF1 (N2212, N2211);
nor NOR3 (N2213, N2191, N274, N714);
not NOT1 (N2214, N2207);
and AND2 (N2215, N2212, N803);
and AND2 (N2216, N2213, N161);
and AND2 (N2217, N2208, N1082);
nor NOR2 (N2218, N2209, N573);
and AND2 (N2219, N2215, N1149);
not NOT1 (N2220, N2219);
and AND2 (N2221, N2205, N2127);
not NOT1 (N2222, N2203);
nor NOR2 (N2223, N2222, N794);
xor XOR2 (N2224, N2202, N44);
or OR3 (N2225, N2217, N324, N1325);
xor XOR2 (N2226, N2216, N1557);
xor XOR2 (N2227, N2223, N309);
nand NAND4 (N2228, N2220, N299, N369, N1508);
buf BUF1 (N2229, N2180);
and AND4 (N2230, N2229, N1087, N644, N380);
not NOT1 (N2231, N2230);
xor XOR2 (N2232, N2224, N609);
and AND4 (N2233, N2221, N848, N1876, N2108);
nor NOR3 (N2234, N2227, N1774, N474);
nand NAND2 (N2235, N2214, N375);
and AND4 (N2236, N2234, N1847, N1482, N856);
and AND4 (N2237, N2218, N1110, N400, N550);
nor NOR2 (N2238, N2235, N5);
nand NAND2 (N2239, N2238, N2237);
nor NOR4 (N2240, N1977, N979, N67, N1136);
or OR3 (N2241, N2239, N997, N1679);
nand NAND2 (N2242, N2228, N36);
buf BUF1 (N2243, N2241);
not NOT1 (N2244, N2236);
buf BUF1 (N2245, N2225);
buf BUF1 (N2246, N2244);
and AND2 (N2247, N2226, N775);
and AND2 (N2248, N2247, N284);
nand NAND2 (N2249, N2242, N1935);
buf BUF1 (N2250, N2210);
or OR3 (N2251, N2246, N140, N1463);
buf BUF1 (N2252, N2243);
nand NAND3 (N2253, N2240, N2070, N2212);
not NOT1 (N2254, N2251);
and AND2 (N2255, N2250, N1866);
xor XOR2 (N2256, N2231, N1336);
buf BUF1 (N2257, N2248);
or OR4 (N2258, N2254, N443, N390, N1734);
nor NOR4 (N2259, N2233, N51, N2131, N803);
not NOT1 (N2260, N2252);
or OR4 (N2261, N2253, N1208, N2234, N454);
xor XOR2 (N2262, N2261, N286);
xor XOR2 (N2263, N2258, N1586);
nand NAND2 (N2264, N2232, N1027);
nor NOR4 (N2265, N2260, N2117, N399, N1983);
and AND3 (N2266, N2249, N344, N932);
or OR3 (N2267, N2263, N1048, N528);
nand NAND2 (N2268, N2255, N1120);
buf BUF1 (N2269, N2259);
nand NAND2 (N2270, N2266, N806);
buf BUF1 (N2271, N2270);
buf BUF1 (N2272, N2265);
not NOT1 (N2273, N2272);
xor XOR2 (N2274, N2273, N948);
and AND3 (N2275, N2257, N1953, N1564);
buf BUF1 (N2276, N2264);
buf BUF1 (N2277, N2269);
nor NOR2 (N2278, N2245, N61);
not NOT1 (N2279, N2262);
or OR2 (N2280, N2274, N753);
buf BUF1 (N2281, N2268);
or OR2 (N2282, N2267, N1969);
nand NAND4 (N2283, N2271, N2170, N582, N151);
nor NOR3 (N2284, N2283, N703, N1261);
or OR3 (N2285, N2275, N1547, N176);
buf BUF1 (N2286, N2284);
not NOT1 (N2287, N2285);
and AND2 (N2288, N2279, N522);
buf BUF1 (N2289, N2278);
or OR3 (N2290, N2281, N386, N2111);
and AND3 (N2291, N2286, N1364, N1480);
buf BUF1 (N2292, N2282);
and AND3 (N2293, N2289, N1013, N1290);
or OR2 (N2294, N2256, N1805);
not NOT1 (N2295, N2277);
nor NOR2 (N2296, N2280, N1441);
or OR3 (N2297, N2287, N2208, N495);
not NOT1 (N2298, N2276);
buf BUF1 (N2299, N2290);
or OR4 (N2300, N2299, N946, N1281, N599);
and AND3 (N2301, N2296, N242, N329);
nor NOR2 (N2302, N2293, N2099);
nand NAND4 (N2303, N2300, N313, N633, N303);
or OR2 (N2304, N2297, N2284);
buf BUF1 (N2305, N2304);
not NOT1 (N2306, N2295);
or OR3 (N2307, N2292, N796, N2279);
or OR2 (N2308, N2303, N872);
not NOT1 (N2309, N2302);
not NOT1 (N2310, N2291);
nor NOR4 (N2311, N2294, N1717, N1225, N808);
nand NAND2 (N2312, N2306, N362);
or OR3 (N2313, N2309, N1948, N382);
not NOT1 (N2314, N2288);
and AND4 (N2315, N2310, N462, N1452, N931);
or OR3 (N2316, N2305, N1516, N674);
nand NAND3 (N2317, N2312, N190, N1686);
buf BUF1 (N2318, N2308);
and AND2 (N2319, N2298, N17);
xor XOR2 (N2320, N2313, N1742);
nor NOR4 (N2321, N2315, N381, N1252, N1620);
xor XOR2 (N2322, N2320, N1578);
buf BUF1 (N2323, N2307);
xor XOR2 (N2324, N2301, N191);
nand NAND3 (N2325, N2316, N560, N2315);
xor XOR2 (N2326, N2322, N2305);
not NOT1 (N2327, N2324);
xor XOR2 (N2328, N2323, N1907);
nor NOR3 (N2329, N2321, N1131, N2050);
and AND4 (N2330, N2328, N1636, N1346, N1119);
not NOT1 (N2331, N2325);
buf BUF1 (N2332, N2327);
buf BUF1 (N2333, N2332);
xor XOR2 (N2334, N2319, N1732);
not NOT1 (N2335, N2329);
xor XOR2 (N2336, N2318, N1607);
xor XOR2 (N2337, N2333, N1774);
buf BUF1 (N2338, N2337);
xor XOR2 (N2339, N2334, N667);
nor NOR4 (N2340, N2326, N1992, N922, N893);
and AND3 (N2341, N2330, N943, N1809);
not NOT1 (N2342, N2335);
not NOT1 (N2343, N2331);
nand NAND2 (N2344, N2311, N991);
nor NOR4 (N2345, N2342, N551, N504, N1399);
xor XOR2 (N2346, N2345, N1354);
or OR4 (N2347, N2314, N1419, N1098, N2022);
nor NOR2 (N2348, N2317, N1527);
not NOT1 (N2349, N2347);
and AND2 (N2350, N2340, N2203);
nand NAND2 (N2351, N2336, N338);
xor XOR2 (N2352, N2344, N340);
nand NAND4 (N2353, N2352, N1099, N1062, N320);
or OR3 (N2354, N2346, N527, N1655);
buf BUF1 (N2355, N2343);
nand NAND4 (N2356, N2341, N147, N1059, N1243);
buf BUF1 (N2357, N2350);
or OR3 (N2358, N2339, N370, N1973);
nor NOR2 (N2359, N2358, N1577);
and AND4 (N2360, N2351, N1166, N157, N312);
xor XOR2 (N2361, N2349, N1483);
xor XOR2 (N2362, N2359, N1864);
xor XOR2 (N2363, N2338, N1521);
xor XOR2 (N2364, N2361, N2040);
and AND4 (N2365, N2353, N491, N1728, N155);
buf BUF1 (N2366, N2348);
or OR2 (N2367, N2357, N1304);
or OR4 (N2368, N2362, N1285, N1448, N1530);
buf BUF1 (N2369, N2360);
and AND4 (N2370, N2368, N2018, N1796, N91);
buf BUF1 (N2371, N2366);
nand NAND2 (N2372, N2363, N718);
and AND2 (N2373, N2370, N921);
not NOT1 (N2374, N2365);
and AND2 (N2375, N2374, N1567);
nand NAND2 (N2376, N2372, N1708);
and AND3 (N2377, N2375, N166, N16);
not NOT1 (N2378, N2355);
nor NOR4 (N2379, N2364, N579, N1388, N1718);
nor NOR4 (N2380, N2367, N357, N972, N1188);
or OR2 (N2381, N2354, N1663);
nor NOR2 (N2382, N2379, N17);
and AND2 (N2383, N2380, N1302);
nand NAND4 (N2384, N2381, N148, N265, N829);
xor XOR2 (N2385, N2369, N2247);
and AND4 (N2386, N2382, N1080, N346, N1995);
nor NOR3 (N2387, N2356, N1238, N479);
nand NAND4 (N2388, N2387, N324, N389, N2035);
buf BUF1 (N2389, N2373);
xor XOR2 (N2390, N2388, N343);
buf BUF1 (N2391, N2389);
buf BUF1 (N2392, N2391);
nor NOR2 (N2393, N2390, N108);
xor XOR2 (N2394, N2392, N1116);
buf BUF1 (N2395, N2383);
buf BUF1 (N2396, N2376);
and AND4 (N2397, N2395, N2129, N416, N597);
nor NOR3 (N2398, N2371, N932, N889);
xor XOR2 (N2399, N2385, N463);
not NOT1 (N2400, N2394);
nand NAND4 (N2401, N2384, N1484, N1984, N1211);
nor NOR2 (N2402, N2377, N1488);
nand NAND2 (N2403, N2393, N1254);
xor XOR2 (N2404, N2396, N1213);
nor NOR3 (N2405, N2386, N1781, N1595);
xor XOR2 (N2406, N2402, N1550);
or OR2 (N2407, N2398, N1871);
xor XOR2 (N2408, N2406, N218);
nor NOR3 (N2409, N2397, N1480, N240);
nor NOR4 (N2410, N2404, N1772, N777, N1495);
buf BUF1 (N2411, N2401);
or OR2 (N2412, N2403, N742);
and AND4 (N2413, N2409, N2110, N1949, N1353);
xor XOR2 (N2414, N2407, N2364);
nand NAND4 (N2415, N2412, N718, N1919, N816);
buf BUF1 (N2416, N2400);
buf BUF1 (N2417, N2416);
xor XOR2 (N2418, N2410, N124);
nand NAND4 (N2419, N2408, N562, N567, N724);
nand NAND4 (N2420, N2411, N1713, N491, N1900);
or OR2 (N2421, N2399, N824);
nand NAND2 (N2422, N2421, N235);
nand NAND2 (N2423, N2415, N2257);
xor XOR2 (N2424, N2414, N906);
nand NAND4 (N2425, N2418, N1861, N626, N2392);
and AND4 (N2426, N2424, N21, N1518, N1953);
nor NOR3 (N2427, N2413, N31, N2337);
buf BUF1 (N2428, N2425);
or OR3 (N2429, N2422, N72, N227);
or OR2 (N2430, N2378, N360);
and AND4 (N2431, N2423, N363, N2327, N1531);
nand NAND4 (N2432, N2426, N231, N1307, N730);
buf BUF1 (N2433, N2432);
or OR3 (N2434, N2433, N1085, N481);
or OR4 (N2435, N2417, N759, N1349, N793);
nand NAND4 (N2436, N2431, N1776, N1357, N556);
or OR2 (N2437, N2427, N671);
or OR3 (N2438, N2434, N695, N334);
or OR2 (N2439, N2430, N468);
nor NOR3 (N2440, N2420, N1904, N83);
or OR4 (N2441, N2439, N1142, N926, N555);
xor XOR2 (N2442, N2435, N381);
buf BUF1 (N2443, N2437);
nor NOR4 (N2444, N2419, N2346, N691, N796);
nand NAND4 (N2445, N2440, N1181, N701, N1469);
buf BUF1 (N2446, N2444);
or OR4 (N2447, N2405, N1407, N1444, N1713);
nor NOR3 (N2448, N2447, N974, N236);
xor XOR2 (N2449, N2448, N1357);
not NOT1 (N2450, N2429);
nand NAND4 (N2451, N2428, N1193, N39, N1813);
or OR2 (N2452, N2436, N2190);
or OR4 (N2453, N2445, N2168, N881, N359);
buf BUF1 (N2454, N2452);
nor NOR3 (N2455, N2449, N1289, N448);
or OR2 (N2456, N2438, N12);
not NOT1 (N2457, N2455);
nor NOR4 (N2458, N2441, N877, N629, N371);
buf BUF1 (N2459, N2458);
nor NOR2 (N2460, N2454, N1244);
nand NAND2 (N2461, N2453, N419);
nor NOR2 (N2462, N2443, N634);
and AND4 (N2463, N2461, N2455, N2454, N1861);
xor XOR2 (N2464, N2442, N457);
not NOT1 (N2465, N2459);
nand NAND3 (N2466, N2462, N1059, N2213);
or OR4 (N2467, N2456, N2171, N2110, N1271);
nor NOR3 (N2468, N2446, N1294, N626);
nand NAND3 (N2469, N2463, N2149, N788);
nand NAND3 (N2470, N2469, N1598, N2273);
xor XOR2 (N2471, N2467, N1838);
nor NOR4 (N2472, N2464, N1411, N1148, N338);
not NOT1 (N2473, N2451);
and AND3 (N2474, N2468, N276, N2473);
or OR2 (N2475, N2252, N169);
not NOT1 (N2476, N2470);
nand NAND3 (N2477, N2471, N878, N411);
and AND2 (N2478, N2457, N509);
not NOT1 (N2479, N2475);
nor NOR4 (N2480, N2450, N950, N500, N461);
not NOT1 (N2481, N2478);
and AND2 (N2482, N2481, N1645);
and AND3 (N2483, N2465, N502, N725);
nor NOR4 (N2484, N2479, N1070, N1781, N1728);
or OR4 (N2485, N2480, N1187, N2339, N60);
and AND2 (N2486, N2476, N601);
nor NOR3 (N2487, N2460, N1930, N803);
buf BUF1 (N2488, N2466);
or OR4 (N2489, N2485, N1071, N1171, N2037);
buf BUF1 (N2490, N2486);
nor NOR4 (N2491, N2477, N2431, N1398, N1665);
not NOT1 (N2492, N2490);
buf BUF1 (N2493, N2491);
not NOT1 (N2494, N2482);
or OR4 (N2495, N2484, N2472, N364, N1281);
xor XOR2 (N2496, N2490, N1970);
or OR2 (N2497, N2496, N239);
and AND4 (N2498, N2487, N274, N598, N791);
not NOT1 (N2499, N2498);
xor XOR2 (N2500, N2499, N2444);
xor XOR2 (N2501, N2500, N485);
nand NAND3 (N2502, N2501, N389, N365);
nor NOR4 (N2503, N2483, N2492, N104, N2199);
or OR4 (N2504, N1205, N2253, N135, N405);
xor XOR2 (N2505, N2504, N1154);
and AND4 (N2506, N2493, N2019, N815, N1359);
buf BUF1 (N2507, N2474);
nor NOR3 (N2508, N2497, N801, N738);
xor XOR2 (N2509, N2508, N1195);
not NOT1 (N2510, N2489);
xor XOR2 (N2511, N2506, N1254);
nor NOR2 (N2512, N2507, N2021);
not NOT1 (N2513, N2511);
nor NOR4 (N2514, N2503, N402, N13, N351);
or OR2 (N2515, N2512, N1381);
nand NAND2 (N2516, N2505, N1361);
buf BUF1 (N2517, N2513);
buf BUF1 (N2518, N2515);
buf BUF1 (N2519, N2510);
buf BUF1 (N2520, N2517);
nor NOR2 (N2521, N2509, N954);
buf BUF1 (N2522, N2495);
xor XOR2 (N2523, N2516, N720);
nand NAND3 (N2524, N2494, N504, N2083);
buf BUF1 (N2525, N2520);
nor NOR4 (N2526, N2488, N708, N1875, N420);
not NOT1 (N2527, N2502);
and AND2 (N2528, N2527, N2206);
and AND4 (N2529, N2525, N437, N315, N1322);
or OR4 (N2530, N2526, N955, N272, N660);
buf BUF1 (N2531, N2524);
and AND4 (N2532, N2514, N316, N2166, N889);
or OR4 (N2533, N2532, N1132, N1518, N2167);
buf BUF1 (N2534, N2519);
buf BUF1 (N2535, N2528);
nand NAND2 (N2536, N2530, N2371);
or OR2 (N2537, N2535, N1532);
buf BUF1 (N2538, N2529);
not NOT1 (N2539, N2523);
not NOT1 (N2540, N2536);
and AND4 (N2541, N2522, N2230, N2034, N1042);
not NOT1 (N2542, N2541);
nor NOR2 (N2543, N2537, N481);
and AND2 (N2544, N2531, N1311);
xor XOR2 (N2545, N2538, N703);
and AND3 (N2546, N2540, N545, N1418);
not NOT1 (N2547, N2534);
xor XOR2 (N2548, N2544, N85);
nand NAND4 (N2549, N2548, N1511, N1889, N1671);
and AND2 (N2550, N2549, N1029);
xor XOR2 (N2551, N2518, N2533);
xor XOR2 (N2552, N2316, N1414);
or OR4 (N2553, N2545, N739, N1607, N1838);
nand NAND4 (N2554, N2552, N1257, N527, N1539);
and AND2 (N2555, N2542, N2515);
or OR2 (N2556, N2553, N155);
or OR3 (N2557, N2556, N2346, N1023);
and AND4 (N2558, N2539, N842, N1443, N2474);
or OR2 (N2559, N2546, N394);
nand NAND4 (N2560, N2551, N1804, N1314, N51);
nand NAND3 (N2561, N2554, N746, N1585);
nor NOR2 (N2562, N2543, N1282);
or OR2 (N2563, N2547, N2506);
and AND3 (N2564, N2557, N2356, N1442);
not NOT1 (N2565, N2561);
nand NAND3 (N2566, N2564, N1681, N749);
or OR3 (N2567, N2566, N2085, N1772);
not NOT1 (N2568, N2563);
not NOT1 (N2569, N2559);
xor XOR2 (N2570, N2568, N1727);
xor XOR2 (N2571, N2555, N2097);
xor XOR2 (N2572, N2571, N759);
buf BUF1 (N2573, N2565);
nand NAND2 (N2574, N2567, N1695);
or OR4 (N2575, N2573, N2193, N582, N1668);
nand NAND2 (N2576, N2572, N1856);
buf BUF1 (N2577, N2562);
and AND2 (N2578, N2570, N190);
nand NAND2 (N2579, N2576, N1784);
or OR3 (N2580, N2577, N1616, N1315);
and AND4 (N2581, N2575, N768, N1882, N2404);
or OR4 (N2582, N2560, N1983, N1383, N1576);
and AND4 (N2583, N2550, N1569, N1787, N1683);
nor NOR3 (N2584, N2580, N20, N143);
and AND3 (N2585, N2579, N2264, N1079);
not NOT1 (N2586, N2583);
and AND4 (N2587, N2585, N2426, N1318, N616);
xor XOR2 (N2588, N2578, N1210);
buf BUF1 (N2589, N2586);
xor XOR2 (N2590, N2558, N2400);
and AND4 (N2591, N2574, N1462, N532, N2171);
buf BUF1 (N2592, N2591);
nor NOR3 (N2593, N2589, N1882, N878);
not NOT1 (N2594, N2588);
or OR4 (N2595, N2581, N234, N107, N1463);
not NOT1 (N2596, N2594);
and AND3 (N2597, N2569, N2267, N286);
and AND2 (N2598, N2596, N941);
nor NOR4 (N2599, N2521, N943, N943, N398);
and AND3 (N2600, N2599, N1739, N434);
not NOT1 (N2601, N2590);
or OR2 (N2602, N2592, N780);
or OR2 (N2603, N2593, N1973);
xor XOR2 (N2604, N2598, N1383);
nor NOR4 (N2605, N2587, N2307, N2073, N1352);
not NOT1 (N2606, N2595);
or OR2 (N2607, N2601, N2227);
not NOT1 (N2608, N2604);
or OR2 (N2609, N2597, N188);
xor XOR2 (N2610, N2609, N1563);
or OR4 (N2611, N2610, N1693, N689, N771);
xor XOR2 (N2612, N2605, N1850);
nor NOR4 (N2613, N2606, N2518, N812, N1065);
or OR2 (N2614, N2611, N2101);
xor XOR2 (N2615, N2600, N215);
and AND3 (N2616, N2613, N54, N2515);
not NOT1 (N2617, N2614);
and AND3 (N2618, N2602, N1277, N2466);
nand NAND3 (N2619, N2618, N727, N2554);
not NOT1 (N2620, N2619);
nor NOR3 (N2621, N2615, N1300, N2280);
nand NAND3 (N2622, N2620, N824, N2219);
nand NAND2 (N2623, N2621, N1458);
not NOT1 (N2624, N2622);
and AND2 (N2625, N2623, N2377);
xor XOR2 (N2626, N2607, N590);
or OR2 (N2627, N2616, N2305);
buf BUF1 (N2628, N2584);
or OR3 (N2629, N2612, N254, N1558);
buf BUF1 (N2630, N2624);
and AND4 (N2631, N2617, N724, N2300, N1575);
nor NOR4 (N2632, N2626, N65, N2110, N1477);
and AND2 (N2633, N2625, N198);
buf BUF1 (N2634, N2627);
nor NOR4 (N2635, N2603, N2004, N1779, N1885);
and AND4 (N2636, N2628, N1679, N1939, N1995);
buf BUF1 (N2637, N2630);
buf BUF1 (N2638, N2637);
nand NAND3 (N2639, N2635, N1192, N823);
and AND2 (N2640, N2633, N1811);
and AND4 (N2641, N2608, N432, N2374, N2096);
or OR2 (N2642, N2640, N2045);
nor NOR3 (N2643, N2639, N329, N547);
and AND3 (N2644, N2629, N151, N1770);
nand NAND3 (N2645, N2641, N181, N2010);
xor XOR2 (N2646, N2642, N1682);
xor XOR2 (N2647, N2634, N512);
xor XOR2 (N2648, N2647, N1900);
nand NAND4 (N2649, N2646, N2312, N1972, N123);
xor XOR2 (N2650, N2649, N2344);
or OR3 (N2651, N2632, N1552, N1076);
or OR2 (N2652, N2651, N1560);
nor NOR3 (N2653, N2638, N1740, N1728);
or OR3 (N2654, N2631, N913, N2632);
or OR2 (N2655, N2643, N183);
nand NAND4 (N2656, N2582, N29, N931, N1916);
and AND3 (N2657, N2644, N1758, N884);
and AND4 (N2658, N2657, N1929, N2050, N1493);
not NOT1 (N2659, N2636);
not NOT1 (N2660, N2656);
or OR2 (N2661, N2660, N2122);
or OR4 (N2662, N2645, N2303, N1372, N1364);
not NOT1 (N2663, N2654);
nor NOR2 (N2664, N2652, N1761);
and AND4 (N2665, N2658, N2471, N300, N1384);
nor NOR2 (N2666, N2662, N2360);
nor NOR2 (N2667, N2666, N7);
not NOT1 (N2668, N2667);
and AND4 (N2669, N2663, N2366, N352, N1052);
buf BUF1 (N2670, N2669);
or OR4 (N2671, N2655, N1474, N105, N2221);
nor NOR2 (N2672, N2648, N102);
not NOT1 (N2673, N2659);
nand NAND2 (N2674, N2668, N1132);
buf BUF1 (N2675, N2664);
or OR4 (N2676, N2670, N445, N1741, N642);
and AND4 (N2677, N2673, N2440, N897, N1149);
xor XOR2 (N2678, N2671, N1330);
xor XOR2 (N2679, N2678, N1832);
or OR3 (N2680, N2665, N1095, N418);
nand NAND3 (N2681, N2677, N2153, N1214);
and AND4 (N2682, N2674, N772, N142, N1168);
or OR2 (N2683, N2681, N2364);
nand NAND3 (N2684, N2672, N2274, N1676);
or OR4 (N2685, N2653, N746, N1436, N389);
nand NAND2 (N2686, N2683, N2207);
or OR3 (N2687, N2675, N662, N835);
xor XOR2 (N2688, N2650, N1080);
buf BUF1 (N2689, N2687);
xor XOR2 (N2690, N2689, N608);
buf BUF1 (N2691, N2686);
xor XOR2 (N2692, N2688, N192);
nor NOR2 (N2693, N2684, N589);
or OR2 (N2694, N2676, N1931);
xor XOR2 (N2695, N2690, N1369);
or OR3 (N2696, N2694, N2082, N934);
or OR2 (N2697, N2693, N277);
or OR2 (N2698, N2661, N2559);
nand NAND3 (N2699, N2691, N593, N2320);
buf BUF1 (N2700, N2699);
buf BUF1 (N2701, N2685);
xor XOR2 (N2702, N2698, N1618);
nand NAND4 (N2703, N2700, N1376, N229, N1520);
nor NOR4 (N2704, N2682, N2603, N669, N2243);
nand NAND2 (N2705, N2679, N895);
nor NOR4 (N2706, N2704, N1787, N2007, N1057);
nor NOR4 (N2707, N2706, N257, N1641, N2368);
not NOT1 (N2708, N2680);
xor XOR2 (N2709, N2701, N815);
buf BUF1 (N2710, N2696);
buf BUF1 (N2711, N2702);
nor NOR2 (N2712, N2709, N409);
buf BUF1 (N2713, N2705);
nand NAND2 (N2714, N2697, N830);
nand NAND2 (N2715, N2707, N287);
not NOT1 (N2716, N2710);
buf BUF1 (N2717, N2715);
not NOT1 (N2718, N2713);
nand NAND3 (N2719, N2712, N1069, N2428);
xor XOR2 (N2720, N2703, N1095);
buf BUF1 (N2721, N2716);
not NOT1 (N2722, N2719);
and AND4 (N2723, N2711, N730, N1004, N1540);
nor NOR4 (N2724, N2717, N2079, N333, N81);
nand NAND2 (N2725, N2718, N567);
or OR4 (N2726, N2723, N1113, N2593, N2028);
and AND2 (N2727, N2725, N1828);
nor NOR2 (N2728, N2720, N930);
nand NAND4 (N2729, N2728, N1554, N2413, N2676);
or OR2 (N2730, N2722, N2257);
or OR2 (N2731, N2726, N876);
buf BUF1 (N2732, N2714);
and AND2 (N2733, N2730, N292);
nand NAND2 (N2734, N2724, N883);
or OR3 (N2735, N2695, N878, N792);
nand NAND3 (N2736, N2735, N136, N1898);
nor NOR3 (N2737, N2721, N2165, N673);
not NOT1 (N2738, N2736);
xor XOR2 (N2739, N2738, N2454);
not NOT1 (N2740, N2737);
not NOT1 (N2741, N2729);
and AND3 (N2742, N2731, N1167, N964);
and AND2 (N2743, N2741, N273);
nor NOR2 (N2744, N2708, N921);
or OR3 (N2745, N2732, N1393, N1620);
nand NAND4 (N2746, N2692, N1614, N2655, N1844);
buf BUF1 (N2747, N2746);
xor XOR2 (N2748, N2747, N758);
nor NOR2 (N2749, N2727, N1632);
not NOT1 (N2750, N2740);
nor NOR3 (N2751, N2734, N656, N1802);
not NOT1 (N2752, N2744);
xor XOR2 (N2753, N2733, N307);
buf BUF1 (N2754, N2750);
xor XOR2 (N2755, N2751, N554);
xor XOR2 (N2756, N2745, N2106);
nor NOR2 (N2757, N2753, N2722);
buf BUF1 (N2758, N2755);
or OR4 (N2759, N2752, N1528, N1132, N2494);
or OR3 (N2760, N2748, N1461, N983);
nor NOR4 (N2761, N2739, N103, N2311, N125);
nor NOR2 (N2762, N2754, N636);
or OR4 (N2763, N2749, N824, N1285, N711);
buf BUF1 (N2764, N2761);
not NOT1 (N2765, N2760);
nand NAND2 (N2766, N2763, N1319);
xor XOR2 (N2767, N2742, N2691);
not NOT1 (N2768, N2765);
buf BUF1 (N2769, N2743);
xor XOR2 (N2770, N2757, N1225);
and AND4 (N2771, N2767, N1562, N610, N2111);
nand NAND2 (N2772, N2768, N1356);
buf BUF1 (N2773, N2758);
buf BUF1 (N2774, N2769);
xor XOR2 (N2775, N2772, N2556);
or OR4 (N2776, N2775, N385, N838, N623);
buf BUF1 (N2777, N2756);
or OR4 (N2778, N2759, N2275, N2517, N2265);
or OR2 (N2779, N2762, N2358);
not NOT1 (N2780, N2777);
not NOT1 (N2781, N2774);
nor NOR4 (N2782, N2773, N892, N504, N193);
xor XOR2 (N2783, N2764, N1178);
xor XOR2 (N2784, N2766, N255);
nor NOR3 (N2785, N2779, N2206, N1018);
not NOT1 (N2786, N2785);
nand NAND3 (N2787, N2780, N2214, N810);
xor XOR2 (N2788, N2783, N494);
xor XOR2 (N2789, N2770, N2143);
not NOT1 (N2790, N2789);
not NOT1 (N2791, N2788);
not NOT1 (N2792, N2790);
nor NOR4 (N2793, N2778, N457, N932, N33);
and AND3 (N2794, N2782, N1064, N2467);
xor XOR2 (N2795, N2794, N2750);
buf BUF1 (N2796, N2784);
nor NOR3 (N2797, N2795, N2206, N1078);
not NOT1 (N2798, N2791);
nand NAND4 (N2799, N2798, N2112, N1402, N339);
xor XOR2 (N2800, N2787, N2199);
buf BUF1 (N2801, N2793);
nor NOR4 (N2802, N2801, N531, N1545, N1540);
nand NAND3 (N2803, N2786, N1750, N144);
nand NAND3 (N2804, N2800, N2284, N2223);
not NOT1 (N2805, N2796);
nor NOR2 (N2806, N2797, N1520);
nor NOR3 (N2807, N2806, N761, N1724);
buf BUF1 (N2808, N2802);
not NOT1 (N2809, N2804);
not NOT1 (N2810, N2771);
not NOT1 (N2811, N2805);
and AND4 (N2812, N2803, N714, N1610, N1785);
xor XOR2 (N2813, N2808, N1676);
not NOT1 (N2814, N2781);
nand NAND2 (N2815, N2810, N184);
nand NAND3 (N2816, N2809, N1509, N2089);
and AND2 (N2817, N2816, N2702);
or OR4 (N2818, N2813, N1965, N949, N569);
or OR2 (N2819, N2799, N75);
not NOT1 (N2820, N2814);
nor NOR2 (N2821, N2776, N865);
nor NOR4 (N2822, N2807, N1794, N1983, N1075);
buf BUF1 (N2823, N2819);
not NOT1 (N2824, N2811);
or OR3 (N2825, N2822, N657, N2103);
and AND3 (N2826, N2817, N1307, N2217);
or OR3 (N2827, N2824, N2395, N1784);
xor XOR2 (N2828, N2818, N1283);
xor XOR2 (N2829, N2826, N725);
xor XOR2 (N2830, N2823, N1453);
buf BUF1 (N2831, N2827);
not NOT1 (N2832, N2821);
xor XOR2 (N2833, N2832, N579);
nand NAND3 (N2834, N2815, N2384, N834);
and AND2 (N2835, N2825, N2045);
nand NAND3 (N2836, N2829, N1436, N1064);
xor XOR2 (N2837, N2830, N2364);
nor NOR4 (N2838, N2820, N1920, N472, N1006);
and AND2 (N2839, N2837, N2163);
nor NOR2 (N2840, N2834, N2537);
or OR3 (N2841, N2812, N883, N374);
xor XOR2 (N2842, N2839, N1227);
and AND3 (N2843, N2792, N2360, N429);
not NOT1 (N2844, N2835);
nand NAND3 (N2845, N2828, N939, N1758);
nand NAND3 (N2846, N2843, N228, N862);
nand NAND4 (N2847, N2836, N1964, N2311, N462);
and AND2 (N2848, N2833, N2320);
buf BUF1 (N2849, N2831);
nand NAND2 (N2850, N2840, N2588);
nor NOR2 (N2851, N2845, N2514);
not NOT1 (N2852, N2850);
xor XOR2 (N2853, N2851, N1962);
nand NAND4 (N2854, N2838, N1559, N1123, N1165);
nor NOR4 (N2855, N2847, N2794, N1769, N274);
buf BUF1 (N2856, N2852);
nand NAND3 (N2857, N2848, N89, N748);
and AND3 (N2858, N2849, N2000, N1180);
and AND4 (N2859, N2844, N1017, N557, N2073);
nand NAND2 (N2860, N2855, N2675);
xor XOR2 (N2861, N2856, N1121);
xor XOR2 (N2862, N2846, N2445);
not NOT1 (N2863, N2861);
nand NAND2 (N2864, N2860, N2650);
xor XOR2 (N2865, N2859, N770);
nor NOR3 (N2866, N2857, N431, N1663);
or OR4 (N2867, N2866, N1905, N617, N2367);
xor XOR2 (N2868, N2854, N2550);
nand NAND2 (N2869, N2858, N665);
nand NAND4 (N2870, N2853, N423, N203, N2209);
not NOT1 (N2871, N2863);
not NOT1 (N2872, N2869);
or OR3 (N2873, N2867, N266, N2455);
xor XOR2 (N2874, N2842, N2272);
buf BUF1 (N2875, N2862);
buf BUF1 (N2876, N2872);
nor NOR4 (N2877, N2871, N614, N243, N1573);
and AND4 (N2878, N2864, N95, N316, N2460);
or OR3 (N2879, N2868, N2826, N1919);
not NOT1 (N2880, N2841);
xor XOR2 (N2881, N2877, N2199);
buf BUF1 (N2882, N2880);
not NOT1 (N2883, N2870);
nand NAND4 (N2884, N2883, N1710, N420, N2222);
buf BUF1 (N2885, N2881);
xor XOR2 (N2886, N2882, N1451);
nor NOR2 (N2887, N2865, N2500);
nand NAND3 (N2888, N2878, N985, N1784);
buf BUF1 (N2889, N2886);
not NOT1 (N2890, N2873);
not NOT1 (N2891, N2885);
xor XOR2 (N2892, N2879, N2586);
or OR4 (N2893, N2888, N1298, N680, N2617);
and AND2 (N2894, N2890, N2038);
not NOT1 (N2895, N2875);
nand NAND3 (N2896, N2894, N651, N658);
or OR3 (N2897, N2874, N2280, N961);
nand NAND2 (N2898, N2896, N125);
nor NOR3 (N2899, N2889, N2742, N1371);
nor NOR4 (N2900, N2891, N2072, N1660, N2596);
buf BUF1 (N2901, N2893);
nor NOR3 (N2902, N2900, N1253, N1279);
buf BUF1 (N2903, N2902);
xor XOR2 (N2904, N2884, N328);
not NOT1 (N2905, N2903);
and AND3 (N2906, N2887, N2205, N496);
or OR2 (N2907, N2898, N1024);
xor XOR2 (N2908, N2897, N2433);
buf BUF1 (N2909, N2895);
xor XOR2 (N2910, N2907, N2633);
nand NAND4 (N2911, N2876, N669, N2689, N1935);
nor NOR4 (N2912, N2899, N1568, N2193, N2887);
buf BUF1 (N2913, N2911);
nand NAND3 (N2914, N2909, N1352, N2568);
buf BUF1 (N2915, N2910);
nor NOR4 (N2916, N2913, N638, N1673, N2421);
not NOT1 (N2917, N2904);
nand NAND4 (N2918, N2901, N938, N1665, N1905);
and AND4 (N2919, N2905, N889, N510, N1712);
and AND2 (N2920, N2906, N576);
nand NAND4 (N2921, N2912, N1532, N2082, N1838);
buf BUF1 (N2922, N2915);
nor NOR3 (N2923, N2892, N1433, N2325);
and AND3 (N2924, N2916, N1676, N2118);
nor NOR2 (N2925, N2917, N671);
nor NOR2 (N2926, N2922, N1717);
xor XOR2 (N2927, N2908, N2885);
not NOT1 (N2928, N2919);
nand NAND4 (N2929, N2921, N2300, N1271, N2166);
and AND3 (N2930, N2920, N1987, N886);
or OR4 (N2931, N2929, N2091, N1399, N15);
xor XOR2 (N2932, N2918, N1248);
not NOT1 (N2933, N2931);
or OR4 (N2934, N2925, N1423, N2704, N87);
not NOT1 (N2935, N2930);
nand NAND2 (N2936, N2934, N2618);
buf BUF1 (N2937, N2927);
buf BUF1 (N2938, N2932);
xor XOR2 (N2939, N2933, N1022);
buf BUF1 (N2940, N2914);
buf BUF1 (N2941, N2936);
or OR3 (N2942, N2941, N2423, N982);
nand NAND3 (N2943, N2939, N2128, N164);
buf BUF1 (N2944, N2942);
and AND3 (N2945, N2940, N1146, N1269);
not NOT1 (N2946, N2935);
or OR4 (N2947, N2945, N2840, N1065, N1925);
xor XOR2 (N2948, N2924, N1979);
nor NOR4 (N2949, N2943, N1951, N280, N983);
and AND2 (N2950, N2926, N2447);
nor NOR4 (N2951, N2928, N1890, N1071, N2576);
or OR2 (N2952, N2923, N279);
nor NOR2 (N2953, N2950, N2543);
not NOT1 (N2954, N2949);
buf BUF1 (N2955, N2937);
or OR4 (N2956, N2955, N388, N1350, N1825);
buf BUF1 (N2957, N2954);
nor NOR4 (N2958, N2953, N452, N1163, N2206);
nor NOR2 (N2959, N2938, N4);
xor XOR2 (N2960, N2959, N1359);
and AND2 (N2961, N2956, N2440);
or OR3 (N2962, N2951, N381, N2121);
or OR2 (N2963, N2948, N615);
xor XOR2 (N2964, N2957, N1571);
nor NOR3 (N2965, N2944, N1415, N1949);
nor NOR3 (N2966, N2962, N354, N1214);
nand NAND2 (N2967, N2952, N2059);
xor XOR2 (N2968, N2965, N1749);
nor NOR2 (N2969, N2947, N1302);
nor NOR2 (N2970, N2960, N260);
not NOT1 (N2971, N2968);
nor NOR3 (N2972, N2958, N1283, N1296);
nor NOR4 (N2973, N2969, N2047, N550, N2837);
nand NAND3 (N2974, N2971, N2708, N701);
not NOT1 (N2975, N2967);
nor NOR4 (N2976, N2975, N1953, N379, N1725);
not NOT1 (N2977, N2974);
or OR4 (N2978, N2964, N1512, N2846, N2579);
nor NOR2 (N2979, N2978, N828);
not NOT1 (N2980, N2972);
and AND2 (N2981, N2970, N2327);
xor XOR2 (N2982, N2966, N1590);
or OR3 (N2983, N2980, N2287, N232);
nor NOR4 (N2984, N2983, N2952, N1894, N2084);
not NOT1 (N2985, N2973);
nor NOR4 (N2986, N2979, N2184, N875, N1195);
or OR3 (N2987, N2961, N709, N602);
and AND3 (N2988, N2986, N966, N1934);
and AND3 (N2989, N2987, N1643, N1239);
and AND3 (N2990, N2989, N2383, N1156);
nand NAND4 (N2991, N2982, N2128, N2100, N1069);
nor NOR4 (N2992, N2985, N1567, N1259, N2909);
or OR4 (N2993, N2981, N184, N924, N649);
nor NOR4 (N2994, N2992, N1932, N1980, N1492);
nor NOR2 (N2995, N2946, N2526);
nor NOR2 (N2996, N2990, N810);
or OR3 (N2997, N2976, N855, N69);
not NOT1 (N2998, N2994);
nand NAND4 (N2999, N2963, N1739, N1060, N2174);
and AND2 (N3000, N2997, N587);
xor XOR2 (N3001, N2977, N1642);
or OR4 (N3002, N2996, N535, N270, N1460);
not NOT1 (N3003, N2991);
and AND4 (N3004, N3001, N780, N750, N820);
nand NAND2 (N3005, N2993, N431);
xor XOR2 (N3006, N3005, N2090);
and AND4 (N3007, N3002, N1829, N1740, N2572);
xor XOR2 (N3008, N2988, N199);
not NOT1 (N3009, N2995);
or OR4 (N3010, N3006, N2363, N2454, N2985);
buf BUF1 (N3011, N3000);
buf BUF1 (N3012, N3011);
or OR3 (N3013, N3007, N867, N963);
xor XOR2 (N3014, N3008, N2177);
nand NAND4 (N3015, N3010, N942, N1906, N2306);
and AND2 (N3016, N2998, N697);
or OR4 (N3017, N3013, N790, N943, N759);
or OR3 (N3018, N3016, N2639, N538);
buf BUF1 (N3019, N3003);
nand NAND2 (N3020, N2984, N2234);
nor NOR3 (N3021, N2999, N539, N354);
not NOT1 (N3022, N3018);
not NOT1 (N3023, N3014);
not NOT1 (N3024, N3020);
nor NOR2 (N3025, N3009, N2573);
and AND3 (N3026, N3004, N1822, N1805);
buf BUF1 (N3027, N3017);
xor XOR2 (N3028, N3012, N331);
xor XOR2 (N3029, N3023, N2938);
nand NAND3 (N3030, N3026, N584, N1624);
xor XOR2 (N3031, N3028, N1280);
or OR2 (N3032, N3029, N2028);
not NOT1 (N3033, N3027);
and AND3 (N3034, N3019, N1774, N140);
nand NAND2 (N3035, N3033, N1004);
nor NOR4 (N3036, N3022, N537, N2047, N218);
nand NAND3 (N3037, N3015, N953, N2711);
xor XOR2 (N3038, N3025, N2239);
and AND2 (N3039, N3021, N1109);
or OR3 (N3040, N3024, N2752, N254);
xor XOR2 (N3041, N3039, N1095);
nor NOR2 (N3042, N3034, N1253);
and AND4 (N3043, N3038, N1898, N1986, N708);
xor XOR2 (N3044, N3041, N2995);
and AND2 (N3045, N3040, N753);
not NOT1 (N3046, N3036);
or OR2 (N3047, N3031, N1248);
nand NAND3 (N3048, N3035, N1072, N2654);
not NOT1 (N3049, N3037);
xor XOR2 (N3050, N3032, N1582);
nor NOR2 (N3051, N3030, N2825);
and AND4 (N3052, N3048, N1550, N1873, N2616);
or OR2 (N3053, N3052, N882);
xor XOR2 (N3054, N3046, N2937);
nor NOR3 (N3055, N3049, N2017, N798);
buf BUF1 (N3056, N3042);
and AND2 (N3057, N3043, N394);
nor NOR3 (N3058, N3050, N2017, N168);
or OR2 (N3059, N3051, N831);
not NOT1 (N3060, N3045);
nand NAND4 (N3061, N3059, N1106, N1417, N13);
or OR3 (N3062, N3055, N1610, N729);
or OR4 (N3063, N3044, N972, N564, N1925);
or OR3 (N3064, N3063, N1480, N575);
or OR4 (N3065, N3062, N1574, N268, N672);
nand NAND4 (N3066, N3065, N1966, N454, N1334);
not NOT1 (N3067, N3058);
or OR2 (N3068, N3061, N1822);
nand NAND3 (N3069, N3066, N1717, N1756);
nor NOR4 (N3070, N3057, N2304, N1437, N2819);
buf BUF1 (N3071, N3067);
not NOT1 (N3072, N3068);
nor NOR3 (N3073, N3054, N1939, N1305);
buf BUF1 (N3074, N3047);
buf BUF1 (N3075, N3071);
or OR4 (N3076, N3064, N2839, N2725, N43);
not NOT1 (N3077, N3070);
not NOT1 (N3078, N3076);
buf BUF1 (N3079, N3074);
or OR4 (N3080, N3069, N1244, N2638, N2781);
buf BUF1 (N3081, N3079);
nand NAND2 (N3082, N3056, N2089);
or OR3 (N3083, N3081, N2046, N2829);
nand NAND2 (N3084, N3075, N276);
buf BUF1 (N3085, N3060);
and AND2 (N3086, N3078, N939);
and AND2 (N3087, N3086, N2486);
or OR3 (N3088, N3082, N1092, N2003);
nor NOR4 (N3089, N3080, N26, N1457, N580);
buf BUF1 (N3090, N3089);
nor NOR4 (N3091, N3073, N1201, N1659, N1923);
not NOT1 (N3092, N3087);
not NOT1 (N3093, N3053);
xor XOR2 (N3094, N3084, N531);
nor NOR3 (N3095, N3085, N1392, N15);
nand NAND4 (N3096, N3091, N2257, N3062, N639);
buf BUF1 (N3097, N3072);
not NOT1 (N3098, N3096);
not NOT1 (N3099, N3095);
not NOT1 (N3100, N3090);
and AND2 (N3101, N3083, N2308);
xor XOR2 (N3102, N3097, N2475);
buf BUF1 (N3103, N3094);
nor NOR3 (N3104, N3092, N498, N2474);
nor NOR2 (N3105, N3103, N1487);
or OR3 (N3106, N3100, N114, N752);
nor NOR4 (N3107, N3093, N590, N1734, N1013);
or OR2 (N3108, N3098, N2205);
nor NOR4 (N3109, N3077, N2197, N81, N187);
nor NOR2 (N3110, N3107, N2779);
or OR4 (N3111, N3109, N2528, N2826, N795);
nand NAND3 (N3112, N3110, N266, N3058);
xor XOR2 (N3113, N3101, N2083);
not NOT1 (N3114, N3088);
xor XOR2 (N3115, N3112, N2270);
xor XOR2 (N3116, N3111, N420);
nor NOR3 (N3117, N3104, N2972, N497);
or OR4 (N3118, N3117, N2803, N868, N3094);
and AND4 (N3119, N3113, N1202, N1901, N1562);
nor NOR4 (N3120, N3105, N1327, N371, N2278);
nor NOR3 (N3121, N3106, N1902, N2272);
buf BUF1 (N3122, N3116);
xor XOR2 (N3123, N3121, N2981);
buf BUF1 (N3124, N3114);
nor NOR3 (N3125, N3115, N2976, N537);
or OR3 (N3126, N3125, N2792, N1470);
nand NAND4 (N3127, N3118, N712, N1874, N1211);
buf BUF1 (N3128, N3108);
or OR2 (N3129, N3127, N451);
nor NOR2 (N3130, N3099, N1190);
nor NOR2 (N3131, N3124, N667);
xor XOR2 (N3132, N3129, N2938);
and AND4 (N3133, N3128, N1101, N2631, N2675);
nand NAND2 (N3134, N3120, N719);
or OR4 (N3135, N3122, N2156, N422, N659);
not NOT1 (N3136, N3126);
and AND2 (N3137, N3135, N2643);
nor NOR4 (N3138, N3130, N340, N191, N194);
and AND2 (N3139, N3137, N1548);
and AND2 (N3140, N3133, N474);
not NOT1 (N3141, N3102);
not NOT1 (N3142, N3132);
and AND3 (N3143, N3140, N1157, N2641);
xor XOR2 (N3144, N3136, N1234);
not NOT1 (N3145, N3141);
and AND2 (N3146, N3119, N1806);
buf BUF1 (N3147, N3146);
xor XOR2 (N3148, N3144, N754);
or OR4 (N3149, N3139, N1630, N1297, N1985);
and AND3 (N3150, N3131, N356, N3114);
nor NOR3 (N3151, N3138, N731, N444);
nor NOR3 (N3152, N3143, N904, N1054);
nand NAND2 (N3153, N3123, N1161);
or OR3 (N3154, N3134, N291, N118);
nor NOR4 (N3155, N3154, N1073, N29, N1472);
xor XOR2 (N3156, N3142, N212);
nor NOR3 (N3157, N3153, N1654, N905);
xor XOR2 (N3158, N3152, N566);
not NOT1 (N3159, N3145);
not NOT1 (N3160, N3148);
or OR4 (N3161, N3160, N1962, N2334, N1642);
and AND3 (N3162, N3150, N1675, N842);
or OR2 (N3163, N3156, N2695);
not NOT1 (N3164, N3161);
or OR2 (N3165, N3155, N2602);
xor XOR2 (N3166, N3164, N2012);
or OR2 (N3167, N3158, N2663);
or OR4 (N3168, N3147, N1568, N2689, N225);
nor NOR4 (N3169, N3167, N1493, N2375, N486);
nand NAND4 (N3170, N3163, N2873, N2776, N2104);
buf BUF1 (N3171, N3165);
nor NOR2 (N3172, N3171, N390);
not NOT1 (N3173, N3159);
not NOT1 (N3174, N3151);
and AND4 (N3175, N3173, N2774, N2563, N708);
xor XOR2 (N3176, N3149, N3138);
nor NOR2 (N3177, N3157, N498);
not NOT1 (N3178, N3172);
nor NOR2 (N3179, N3169, N122);
not NOT1 (N3180, N3168);
xor XOR2 (N3181, N3174, N3177);
and AND3 (N3182, N397, N861, N557);
not NOT1 (N3183, N3176);
nor NOR4 (N3184, N3182, N1305, N8, N1680);
nand NAND3 (N3185, N3181, N1832, N1707);
and AND3 (N3186, N3170, N3048, N1002);
buf BUF1 (N3187, N3183);
buf BUF1 (N3188, N3178);
not NOT1 (N3189, N3180);
and AND4 (N3190, N3166, N866, N2564, N949);
nor NOR3 (N3191, N3186, N366, N109);
nor NOR3 (N3192, N3188, N1341, N994);
nand NAND3 (N3193, N3189, N1939, N1753);
nand NAND4 (N3194, N3162, N2738, N2831, N99);
and AND3 (N3195, N3187, N583, N1257);
and AND3 (N3196, N3192, N577, N3048);
nand NAND2 (N3197, N3175, N171);
buf BUF1 (N3198, N3185);
or OR4 (N3199, N3195, N1307, N1948, N1343);
xor XOR2 (N3200, N3190, N41);
and AND2 (N3201, N3191, N1925);
xor XOR2 (N3202, N3197, N3031);
nand NAND3 (N3203, N3184, N1735, N367);
or OR2 (N3204, N3194, N891);
and AND3 (N3205, N3203, N1151, N749);
not NOT1 (N3206, N3193);
and AND2 (N3207, N3206, N28);
not NOT1 (N3208, N3205);
or OR2 (N3209, N3202, N1004);
not NOT1 (N3210, N3200);
or OR3 (N3211, N3208, N2514, N1612);
nand NAND3 (N3212, N3201, N1682, N1753);
nor NOR2 (N3213, N3199, N2785);
xor XOR2 (N3214, N3213, N711);
not NOT1 (N3215, N3196);
xor XOR2 (N3216, N3210, N2580);
nor NOR4 (N3217, N3211, N1020, N1454, N1151);
not NOT1 (N3218, N3216);
or OR2 (N3219, N3212, N2827);
and AND3 (N3220, N3217, N1245, N2547);
or OR2 (N3221, N3214, N202);
xor XOR2 (N3222, N3179, N2506);
not NOT1 (N3223, N3222);
buf BUF1 (N3224, N3204);
not NOT1 (N3225, N3207);
buf BUF1 (N3226, N3224);
not NOT1 (N3227, N3221);
nor NOR2 (N3228, N3226, N1035);
buf BUF1 (N3229, N3225);
not NOT1 (N3230, N3220);
nand NAND4 (N3231, N3228, N14, N1656, N218);
and AND4 (N3232, N3219, N594, N2232, N2437);
not NOT1 (N3233, N3230);
and AND3 (N3234, N3218, N2537, N2213);
buf BUF1 (N3235, N3234);
nand NAND3 (N3236, N3198, N285, N566);
xor XOR2 (N3237, N3229, N529);
or OR4 (N3238, N3209, N1679, N2390, N2475);
nand NAND2 (N3239, N3238, N1919);
buf BUF1 (N3240, N3236);
xor XOR2 (N3241, N3239, N2094);
nor NOR3 (N3242, N3241, N1208, N494);
nor NOR4 (N3243, N3227, N587, N649, N2806);
and AND2 (N3244, N3242, N2017);
not NOT1 (N3245, N3233);
and AND3 (N3246, N3240, N2368, N2377);
not NOT1 (N3247, N3237);
buf BUF1 (N3248, N3232);
nand NAND4 (N3249, N3245, N2562, N2553, N183);
and AND3 (N3250, N3235, N1662, N1954);
nor NOR3 (N3251, N3243, N761, N125);
nand NAND3 (N3252, N3251, N2402, N1526);
and AND4 (N3253, N3248, N115, N2876, N2042);
or OR4 (N3254, N3244, N613, N1974, N3126);
and AND4 (N3255, N3249, N2777, N187, N900);
not NOT1 (N3256, N3231);
nor NOR2 (N3257, N3255, N853);
buf BUF1 (N3258, N3254);
buf BUF1 (N3259, N3258);
or OR4 (N3260, N3215, N3166, N1828, N2901);
or OR4 (N3261, N3252, N1738, N1986, N2464);
and AND3 (N3262, N3223, N2247, N57);
buf BUF1 (N3263, N3260);
nor NOR3 (N3264, N3263, N1480, N740);
or OR3 (N3265, N3262, N1603, N2792);
and AND2 (N3266, N3265, N2258);
or OR2 (N3267, N3259, N2863);
or OR3 (N3268, N3267, N1774, N39);
buf BUF1 (N3269, N3247);
nor NOR3 (N3270, N3246, N763, N3256);
and AND4 (N3271, N2187, N442, N1226, N142);
buf BUF1 (N3272, N3261);
xor XOR2 (N3273, N3257, N201);
or OR3 (N3274, N3253, N1843, N863);
xor XOR2 (N3275, N3264, N738);
and AND3 (N3276, N3270, N872, N2208);
buf BUF1 (N3277, N3271);
or OR3 (N3278, N3250, N403, N1036);
xor XOR2 (N3279, N3268, N2510);
and AND4 (N3280, N3276, N3011, N399, N1293);
or OR3 (N3281, N3279, N2411, N3145);
and AND2 (N3282, N3272, N1538);
buf BUF1 (N3283, N3278);
buf BUF1 (N3284, N3280);
not NOT1 (N3285, N3283);
and AND3 (N3286, N3269, N445, N2);
nor NOR4 (N3287, N3282, N553, N2550, N3211);
nor NOR3 (N3288, N3286, N1877, N1926);
and AND3 (N3289, N3287, N1064, N1428);
nand NAND2 (N3290, N3277, N3209);
or OR2 (N3291, N3288, N2187);
xor XOR2 (N3292, N3274, N1170);
nor NOR3 (N3293, N3285, N3065, N422);
not NOT1 (N3294, N3291);
nor NOR2 (N3295, N3281, N1201);
or OR3 (N3296, N3289, N1205, N3038);
nand NAND4 (N3297, N3275, N1907, N2664, N2562);
nand NAND2 (N3298, N3292, N2663);
buf BUF1 (N3299, N3296);
not NOT1 (N3300, N3266);
buf BUF1 (N3301, N3297);
or OR4 (N3302, N3300, N1860, N2245, N3012);
xor XOR2 (N3303, N3295, N30);
or OR3 (N3304, N3302, N3169, N436);
buf BUF1 (N3305, N3304);
not NOT1 (N3306, N3294);
buf BUF1 (N3307, N3303);
nor NOR2 (N3308, N3299, N2646);
buf BUF1 (N3309, N3306);
xor XOR2 (N3310, N3307, N1186);
nor NOR3 (N3311, N3309, N718, N793);
not NOT1 (N3312, N3284);
xor XOR2 (N3313, N3298, N1075);
not NOT1 (N3314, N3293);
nand NAND2 (N3315, N3313, N363);
nand NAND3 (N3316, N3308, N1190, N3141);
xor XOR2 (N3317, N3316, N1723);
or OR4 (N3318, N3273, N1828, N1593, N2052);
buf BUF1 (N3319, N3317);
or OR4 (N3320, N3315, N799, N244, N3278);
xor XOR2 (N3321, N3290, N1583);
nor NOR3 (N3322, N3305, N1421, N39);
nor NOR3 (N3323, N3322, N294, N2007);
not NOT1 (N3324, N3311);
or OR4 (N3325, N3318, N1800, N1394, N488);
buf BUF1 (N3326, N3310);
buf BUF1 (N3327, N3320);
xor XOR2 (N3328, N3319, N593);
not NOT1 (N3329, N3321);
buf BUF1 (N3330, N3323);
and AND4 (N3331, N3330, N232, N2051, N191);
and AND2 (N3332, N3326, N940);
and AND2 (N3333, N3312, N2407);
not NOT1 (N3334, N3327);
nor NOR3 (N3335, N3328, N2071, N2063);
not NOT1 (N3336, N3335);
xor XOR2 (N3337, N3314, N2906);
xor XOR2 (N3338, N3324, N730);
xor XOR2 (N3339, N3301, N1095);
xor XOR2 (N3340, N3337, N2622);
xor XOR2 (N3341, N3331, N2526);
or OR2 (N3342, N3333, N1267);
and AND2 (N3343, N3332, N884);
nand NAND2 (N3344, N3343, N1791);
nand NAND3 (N3345, N3339, N367, N1999);
nor NOR3 (N3346, N3344, N2301, N2114);
or OR4 (N3347, N3340, N2422, N3336, N619);
nand NAND4 (N3348, N1131, N1552, N374, N2752);
nor NOR2 (N3349, N3329, N1923);
not NOT1 (N3350, N3334);
or OR2 (N3351, N3347, N375);
nor NOR3 (N3352, N3346, N1998, N1079);
buf BUF1 (N3353, N3338);
and AND3 (N3354, N3345, N549, N1860);
nand NAND4 (N3355, N3354, N2932, N2030, N646);
or OR2 (N3356, N3348, N1522);
buf BUF1 (N3357, N3325);
nor NOR3 (N3358, N3356, N14, N1661);
nand NAND2 (N3359, N3351, N16);
and AND2 (N3360, N3350, N2838);
nor NOR2 (N3361, N3342, N2637);
nor NOR2 (N3362, N3341, N1884);
and AND3 (N3363, N3353, N51, N1123);
nor NOR4 (N3364, N3359, N201, N3209, N506);
not NOT1 (N3365, N3352);
and AND3 (N3366, N3362, N3193, N1683);
nor NOR4 (N3367, N3357, N3189, N2461, N1464);
xor XOR2 (N3368, N3358, N2344);
nor NOR2 (N3369, N3368, N1268);
nand NAND4 (N3370, N3367, N180, N2316, N3029);
and AND2 (N3371, N3349, N2670);
or OR4 (N3372, N3366, N1725, N2934, N484);
buf BUF1 (N3373, N3355);
nor NOR4 (N3374, N3370, N948, N607, N573);
nand NAND2 (N3375, N3365, N1922);
xor XOR2 (N3376, N3371, N1041);
or OR3 (N3377, N3360, N2192, N1337);
nand NAND3 (N3378, N3375, N674, N355);
xor XOR2 (N3379, N3372, N3033);
and AND3 (N3380, N3377, N2321, N2965);
not NOT1 (N3381, N3380);
buf BUF1 (N3382, N3363);
and AND4 (N3383, N3381, N1713, N2352, N599);
nand NAND2 (N3384, N3361, N1411);
and AND3 (N3385, N3379, N217, N895);
xor XOR2 (N3386, N3376, N2060);
and AND4 (N3387, N3373, N2197, N721, N426);
nand NAND3 (N3388, N3382, N3046, N2451);
nand NAND4 (N3389, N3386, N788, N1982, N1298);
nand NAND2 (N3390, N3385, N1396);
nand NAND3 (N3391, N3384, N1047, N2396);
nand NAND2 (N3392, N3383, N1072);
not NOT1 (N3393, N3378);
or OR4 (N3394, N3364, N3045, N2015, N1674);
nand NAND2 (N3395, N3392, N2632);
not NOT1 (N3396, N3374);
nand NAND4 (N3397, N3388, N740, N393, N3158);
nand NAND2 (N3398, N3391, N2488);
xor XOR2 (N3399, N3393, N1161);
nand NAND3 (N3400, N3387, N1205, N1693);
buf BUF1 (N3401, N3400);
or OR3 (N3402, N3397, N1355, N2128);
xor XOR2 (N3403, N3399, N2428);
xor XOR2 (N3404, N3395, N1863);
nor NOR2 (N3405, N3394, N965);
and AND2 (N3406, N3402, N3022);
buf BUF1 (N3407, N3369);
nand NAND2 (N3408, N3389, N2751);
buf BUF1 (N3409, N3398);
nand NAND4 (N3410, N3408, N3246, N3370, N3354);
and AND3 (N3411, N3404, N2024, N3026);
nor NOR2 (N3412, N3403, N2627);
nor NOR4 (N3413, N3406, N763, N2985, N698);
nand NAND4 (N3414, N3411, N2331, N1756, N2496);
nand NAND2 (N3415, N3401, N2270);
nor NOR3 (N3416, N3413, N489, N1534);
nor NOR2 (N3417, N3414, N1518);
nand NAND2 (N3418, N3407, N2957);
xor XOR2 (N3419, N3418, N1508);
and AND3 (N3420, N3419, N3010, N3225);
nor NOR4 (N3421, N3417, N811, N3108, N3242);
buf BUF1 (N3422, N3412);
nor NOR4 (N3423, N3409, N617, N2449, N2306);
buf BUF1 (N3424, N3396);
or OR2 (N3425, N3410, N2493);
not NOT1 (N3426, N3423);
nand NAND2 (N3427, N3405, N3206);
not NOT1 (N3428, N3416);
nand NAND2 (N3429, N3424, N698);
not NOT1 (N3430, N3420);
nor NOR3 (N3431, N3390, N1111, N2536);
buf BUF1 (N3432, N3431);
and AND3 (N3433, N3422, N2428, N2948);
buf BUF1 (N3434, N3428);
nand NAND4 (N3435, N3430, N699, N3296, N3381);
and AND4 (N3436, N3415, N2920, N133, N1093);
and AND2 (N3437, N3435, N561);
nor NOR4 (N3438, N3427, N1407, N439, N2346);
xor XOR2 (N3439, N3429, N2551);
nand NAND3 (N3440, N3426, N1216, N1608);
buf BUF1 (N3441, N3425);
buf BUF1 (N3442, N3437);
nor NOR3 (N3443, N3434, N2189, N836);
or OR3 (N3444, N3443, N173, N48);
buf BUF1 (N3445, N3436);
nand NAND2 (N3446, N3441, N1521);
nor NOR2 (N3447, N3440, N3446);
or OR2 (N3448, N1735, N1758);
and AND3 (N3449, N3448, N2651, N268);
nor NOR4 (N3450, N3447, N2083, N3366, N3083);
not NOT1 (N3451, N3433);
xor XOR2 (N3452, N3438, N103);
xor XOR2 (N3453, N3444, N2839);
not NOT1 (N3454, N3452);
buf BUF1 (N3455, N3454);
nand NAND2 (N3456, N3451, N594);
buf BUF1 (N3457, N3456);
nand NAND2 (N3458, N3453, N3031);
or OR2 (N3459, N3421, N1255);
nor NOR2 (N3460, N3432, N3076);
nand NAND4 (N3461, N3458, N965, N825, N1729);
buf BUF1 (N3462, N3459);
xor XOR2 (N3463, N3445, N578);
nand NAND2 (N3464, N3461, N709);
nor NOR4 (N3465, N3450, N779, N2240, N395);
nor NOR3 (N3466, N3465, N227, N1717);
not NOT1 (N3467, N3463);
xor XOR2 (N3468, N3466, N559);
nor NOR3 (N3469, N3464, N2768, N1795);
or OR2 (N3470, N3469, N2331);
xor XOR2 (N3471, N3455, N1883);
nor NOR2 (N3472, N3470, N874);
or OR3 (N3473, N3472, N884, N1242);
xor XOR2 (N3474, N3462, N519);
or OR2 (N3475, N3471, N591);
nand NAND4 (N3476, N3474, N1647, N56, N1086);
buf BUF1 (N3477, N3468);
xor XOR2 (N3478, N3467, N2308);
xor XOR2 (N3479, N3478, N1933);
nor NOR4 (N3480, N3460, N1647, N477, N1624);
or OR3 (N3481, N3479, N1718, N1133);
or OR3 (N3482, N3449, N2427, N314);
nand NAND3 (N3483, N3473, N1460, N1922);
and AND3 (N3484, N3483, N1171, N878);
nand NAND2 (N3485, N3439, N248);
and AND4 (N3486, N3477, N1470, N1688, N2123);
and AND4 (N3487, N3482, N1132, N1032, N513);
not NOT1 (N3488, N3486);
nor NOR4 (N3489, N3480, N2549, N590, N2552);
and AND3 (N3490, N3488, N3392, N868);
not NOT1 (N3491, N3476);
not NOT1 (N3492, N3457);
buf BUF1 (N3493, N3491);
buf BUF1 (N3494, N3475);
buf BUF1 (N3495, N3492);
or OR2 (N3496, N3484, N1007);
and AND4 (N3497, N3496, N1797, N2693, N728);
not NOT1 (N3498, N3490);
nor NOR2 (N3499, N3489, N796);
buf BUF1 (N3500, N3487);
and AND2 (N3501, N3485, N2980);
nor NOR3 (N3502, N3494, N2794, N2476);
buf BUF1 (N3503, N3501);
not NOT1 (N3504, N3481);
buf BUF1 (N3505, N3498);
and AND4 (N3506, N3504, N883, N2993, N2700);
buf BUF1 (N3507, N3503);
not NOT1 (N3508, N3500);
buf BUF1 (N3509, N3502);
not NOT1 (N3510, N3507);
and AND4 (N3511, N3497, N2134, N1020, N62);
xor XOR2 (N3512, N3442, N1975);
buf BUF1 (N3513, N3510);
and AND4 (N3514, N3512, N160, N2939, N2782);
buf BUF1 (N3515, N3506);
and AND3 (N3516, N3513, N3304, N3394);
nor NOR4 (N3517, N3505, N619, N1478, N2075);
buf BUF1 (N3518, N3493);
and AND4 (N3519, N3516, N2339, N2246, N2427);
nor NOR3 (N3520, N3509, N1224, N224);
nor NOR4 (N3521, N3508, N1097, N11, N22);
nor NOR3 (N3522, N3518, N59, N2205);
xor XOR2 (N3523, N3499, N2397);
or OR2 (N3524, N3523, N1096);
and AND3 (N3525, N3514, N364, N1356);
not NOT1 (N3526, N3517);
nor NOR3 (N3527, N3495, N1482, N2160);
xor XOR2 (N3528, N3519, N1176);
buf BUF1 (N3529, N3524);
not NOT1 (N3530, N3525);
nand NAND3 (N3531, N3530, N1589, N911);
and AND2 (N3532, N3515, N2475);
and AND3 (N3533, N3531, N2690, N979);
nor NOR4 (N3534, N3528, N1691, N389, N1661);
not NOT1 (N3535, N3527);
not NOT1 (N3536, N3511);
buf BUF1 (N3537, N3536);
nand NAND2 (N3538, N3529, N1999);
and AND4 (N3539, N3537, N3505, N3458, N2626);
not NOT1 (N3540, N3533);
xor XOR2 (N3541, N3520, N297);
and AND2 (N3542, N3540, N2217);
not NOT1 (N3543, N3532);
not NOT1 (N3544, N3526);
and AND3 (N3545, N3542, N3095, N3016);
xor XOR2 (N3546, N3539, N2626);
xor XOR2 (N3547, N3538, N3394);
or OR3 (N3548, N3543, N1223, N616);
not NOT1 (N3549, N3534);
buf BUF1 (N3550, N3548);
buf BUF1 (N3551, N3545);
or OR4 (N3552, N3550, N1069, N248, N1267);
nor NOR2 (N3553, N3522, N2123);
nor NOR2 (N3554, N3546, N608);
xor XOR2 (N3555, N3553, N2264);
nand NAND3 (N3556, N3521, N1371, N1685);
and AND2 (N3557, N3551, N2633);
xor XOR2 (N3558, N3535, N717);
or OR3 (N3559, N3541, N3233, N632);
nand NAND3 (N3560, N3557, N331, N2765);
nand NAND2 (N3561, N3558, N2109);
xor XOR2 (N3562, N3549, N1925);
buf BUF1 (N3563, N3556);
and AND3 (N3564, N3547, N2705, N2648);
buf BUF1 (N3565, N3552);
nor NOR2 (N3566, N3561, N2216);
xor XOR2 (N3567, N3544, N980);
xor XOR2 (N3568, N3565, N2087);
xor XOR2 (N3569, N3554, N2619);
nor NOR4 (N3570, N3564, N3111, N1287, N579);
nand NAND4 (N3571, N3566, N937, N1486, N159);
and AND3 (N3572, N3562, N1293, N3125);
nand NAND2 (N3573, N3559, N1921);
and AND4 (N3574, N3572, N419, N1270, N1393);
xor XOR2 (N3575, N3570, N764);
xor XOR2 (N3576, N3575, N2588);
nor NOR2 (N3577, N3571, N2363);
not NOT1 (N3578, N3568);
xor XOR2 (N3579, N3560, N861);
nand NAND3 (N3580, N3569, N3056, N650);
and AND3 (N3581, N3577, N3496, N2717);
xor XOR2 (N3582, N3555, N7);
xor XOR2 (N3583, N3579, N593);
and AND4 (N3584, N3582, N970, N518, N1696);
buf BUF1 (N3585, N3581);
and AND3 (N3586, N3573, N1380, N2075);
nor NOR2 (N3587, N3585, N752);
not NOT1 (N3588, N3583);
and AND3 (N3589, N3580, N2806, N2974);
and AND3 (N3590, N3589, N521, N1482);
and AND4 (N3591, N3588, N1117, N2428, N2126);
not NOT1 (N3592, N3563);
and AND4 (N3593, N3584, N3388, N40, N556);
buf BUF1 (N3594, N3593);
buf BUF1 (N3595, N3592);
nand NAND4 (N3596, N3594, N3198, N1784, N729);
or OR4 (N3597, N3576, N1432, N1510, N831);
nor NOR4 (N3598, N3591, N749, N3396, N459);
xor XOR2 (N3599, N3586, N198);
and AND4 (N3600, N3599, N2416, N1446, N2520);
not NOT1 (N3601, N3598);
or OR2 (N3602, N3597, N876);
or OR2 (N3603, N3590, N2611);
not NOT1 (N3604, N3567);
xor XOR2 (N3605, N3574, N136);
nor NOR3 (N3606, N3604, N21, N3320);
and AND3 (N3607, N3602, N1367, N2243);
or OR4 (N3608, N3600, N3522, N2379, N1354);
nor NOR4 (N3609, N3608, N98, N3179, N3245);
nor NOR3 (N3610, N3595, N2051, N1992);
nand NAND2 (N3611, N3609, N242);
buf BUF1 (N3612, N3603);
xor XOR2 (N3613, N3610, N2039);
and AND3 (N3614, N3578, N1866, N416);
nor NOR3 (N3615, N3601, N3138, N1612);
nor NOR3 (N3616, N3605, N2199, N1978);
or OR2 (N3617, N3596, N2097);
xor XOR2 (N3618, N3606, N2263);
buf BUF1 (N3619, N3612);
nand NAND3 (N3620, N3617, N43, N2508);
and AND3 (N3621, N3611, N476, N1900);
nand NAND2 (N3622, N3620, N1916);
xor XOR2 (N3623, N3607, N1418);
or OR2 (N3624, N3623, N596);
not NOT1 (N3625, N3619);
xor XOR2 (N3626, N3614, N2957);
nor NOR2 (N3627, N3621, N3114);
or OR4 (N3628, N3624, N601, N1926, N1962);
xor XOR2 (N3629, N3613, N3464);
not NOT1 (N3630, N3629);
nor NOR2 (N3631, N3616, N1843);
nor NOR3 (N3632, N3626, N839, N1875);
buf BUF1 (N3633, N3632);
xor XOR2 (N3634, N3628, N1432);
nand NAND3 (N3635, N3627, N1863, N2134);
and AND3 (N3636, N3631, N3017, N2472);
nand NAND2 (N3637, N3625, N1459);
nor NOR2 (N3638, N3636, N1531);
nor NOR4 (N3639, N3633, N1173, N1017, N2107);
xor XOR2 (N3640, N3637, N3225);
not NOT1 (N3641, N3640);
nor NOR3 (N3642, N3641, N3477, N2065);
nand NAND4 (N3643, N3630, N840, N642, N568);
xor XOR2 (N3644, N3642, N2739);
nor NOR3 (N3645, N3638, N3126, N1629);
nor NOR4 (N3646, N3639, N3640, N3257, N224);
nor NOR3 (N3647, N3643, N413, N3317);
and AND3 (N3648, N3622, N567, N699);
and AND2 (N3649, N3644, N460);
nand NAND3 (N3650, N3645, N740, N906);
buf BUF1 (N3651, N3634);
and AND4 (N3652, N3649, N2218, N3402, N2037);
nor NOR4 (N3653, N3615, N2383, N320, N2764);
xor XOR2 (N3654, N3653, N1231);
xor XOR2 (N3655, N3635, N90);
nor NOR2 (N3656, N3655, N525);
nor NOR3 (N3657, N3646, N3323, N1703);
xor XOR2 (N3658, N3652, N2777);
not NOT1 (N3659, N3648);
or OR2 (N3660, N3656, N1835);
xor XOR2 (N3661, N3658, N1692);
or OR4 (N3662, N3587, N3068, N540, N413);
nand NAND4 (N3663, N3618, N1516, N3581, N1788);
nand NAND3 (N3664, N3651, N1722, N1941);
buf BUF1 (N3665, N3657);
nand NAND2 (N3666, N3664, N3575);
or OR3 (N3667, N3647, N276, N1154);
nand NAND2 (N3668, N3660, N1269);
nor NOR4 (N3669, N3663, N1618, N1316, N2478);
nand NAND2 (N3670, N3669, N1632);
nand NAND4 (N3671, N3665, N3177, N3414, N2640);
and AND4 (N3672, N3659, N1324, N3204, N611);
not NOT1 (N3673, N3668);
and AND3 (N3674, N3654, N1293, N2259);
not NOT1 (N3675, N3650);
buf BUF1 (N3676, N3667);
nand NAND2 (N3677, N3675, N2835);
or OR2 (N3678, N3674, N3299);
and AND4 (N3679, N3662, N2818, N1016, N1653);
and AND3 (N3680, N3671, N3523, N3081);
nor NOR3 (N3681, N3678, N3479, N2333);
buf BUF1 (N3682, N3679);
nor NOR2 (N3683, N3666, N1471);
or OR4 (N3684, N3676, N1244, N2274, N2735);
not NOT1 (N3685, N3680);
or OR4 (N3686, N3685, N1021, N727, N2412);
nor NOR2 (N3687, N3683, N1222);
not NOT1 (N3688, N3673);
not NOT1 (N3689, N3686);
buf BUF1 (N3690, N3684);
and AND3 (N3691, N3682, N2591, N384);
nor NOR4 (N3692, N3691, N2887, N2669, N874);
not NOT1 (N3693, N3690);
or OR2 (N3694, N3677, N3228);
not NOT1 (N3695, N3670);
nor NOR2 (N3696, N3688, N1413);
and AND3 (N3697, N3672, N2307, N2580);
buf BUF1 (N3698, N3693);
nand NAND3 (N3699, N3687, N1010, N2142);
and AND3 (N3700, N3695, N75, N3248);
and AND2 (N3701, N3696, N334);
and AND4 (N3702, N3661, N962, N1431, N132);
buf BUF1 (N3703, N3681);
nor NOR2 (N3704, N3697, N652);
nor NOR3 (N3705, N3704, N1040, N1321);
buf BUF1 (N3706, N3700);
not NOT1 (N3707, N3701);
nand NAND3 (N3708, N3698, N523, N3064);
nand NAND4 (N3709, N3702, N616, N1324, N1702);
not NOT1 (N3710, N3694);
nand NAND2 (N3711, N3689, N2644);
or OR3 (N3712, N3703, N3046, N2659);
nand NAND3 (N3713, N3712, N1379, N2631);
nor NOR3 (N3714, N3708, N426, N281);
not NOT1 (N3715, N3706);
not NOT1 (N3716, N3710);
or OR4 (N3717, N3715, N619, N1778, N577);
nand NAND4 (N3718, N3705, N1558, N1312, N465);
and AND3 (N3719, N3716, N2284, N3623);
or OR3 (N3720, N3699, N1533, N1128);
nand NAND4 (N3721, N3717, N312, N1672, N230);
buf BUF1 (N3722, N3707);
xor XOR2 (N3723, N3718, N268);
and AND3 (N3724, N3723, N3100, N2981);
buf BUF1 (N3725, N3721);
buf BUF1 (N3726, N3719);
xor XOR2 (N3727, N3714, N608);
or OR3 (N3728, N3727, N2657, N2050);
nand NAND4 (N3729, N3726, N3001, N2016, N2195);
or OR4 (N3730, N3720, N706, N1371, N1806);
nor NOR2 (N3731, N3709, N746);
not NOT1 (N3732, N3728);
nand NAND4 (N3733, N3732, N2635, N1616, N3632);
buf BUF1 (N3734, N3692);
and AND4 (N3735, N3722, N2454, N2275, N2146);
nor NOR3 (N3736, N3735, N312, N2050);
or OR2 (N3737, N3729, N2450);
nor NOR2 (N3738, N3713, N911);
xor XOR2 (N3739, N3737, N1026);
and AND3 (N3740, N3730, N122, N3228);
nand NAND3 (N3741, N3734, N2665, N3153);
or OR4 (N3742, N3739, N1757, N3028, N3359);
and AND2 (N3743, N3725, N2985);
or OR2 (N3744, N3740, N998);
nand NAND2 (N3745, N3733, N178);
buf BUF1 (N3746, N3743);
and AND2 (N3747, N3742, N2451);
xor XOR2 (N3748, N3745, N3608);
not NOT1 (N3749, N3711);
xor XOR2 (N3750, N3731, N2489);
and AND4 (N3751, N3744, N1557, N3013, N3278);
nor NOR2 (N3752, N3736, N3373);
nor NOR3 (N3753, N3749, N1155, N3406);
nor NOR2 (N3754, N3724, N3318);
and AND2 (N3755, N3750, N1218);
or OR4 (N3756, N3753, N3724, N2872, N1338);
or OR3 (N3757, N3755, N1232, N3236);
xor XOR2 (N3758, N3748, N3468);
nor NOR4 (N3759, N3758, N653, N903, N1257);
nor NOR4 (N3760, N3756, N264, N2666, N2558);
nor NOR2 (N3761, N3752, N2662);
nor NOR4 (N3762, N3754, N442, N1331, N590);
or OR4 (N3763, N3762, N3689, N3528, N771);
nand NAND3 (N3764, N3759, N1367, N1441);
not NOT1 (N3765, N3763);
buf BUF1 (N3766, N3747);
xor XOR2 (N3767, N3765, N2371);
xor XOR2 (N3768, N3746, N114);
and AND4 (N3769, N3761, N3472, N126, N1261);
nand NAND3 (N3770, N3764, N3058, N107);
buf BUF1 (N3771, N3760);
and AND2 (N3772, N3770, N3248);
xor XOR2 (N3773, N3741, N2817);
xor XOR2 (N3774, N3767, N1004);
nand NAND3 (N3775, N3768, N1554, N1790);
and AND2 (N3776, N3772, N3012);
and AND2 (N3777, N3738, N1106);
xor XOR2 (N3778, N3751, N2337);
or OR2 (N3779, N3771, N2511);
or OR2 (N3780, N3779, N3276);
xor XOR2 (N3781, N3757, N1581);
not NOT1 (N3782, N3774);
xor XOR2 (N3783, N3780, N3704);
nand NAND4 (N3784, N3776, N2968, N3417, N2655);
xor XOR2 (N3785, N3782, N1702);
nand NAND2 (N3786, N3775, N433);
buf BUF1 (N3787, N3766);
buf BUF1 (N3788, N3787);
nand NAND2 (N3789, N3784, N2279);
not NOT1 (N3790, N3786);
not NOT1 (N3791, N3781);
and AND2 (N3792, N3778, N546);
buf BUF1 (N3793, N3788);
and AND4 (N3794, N3785, N1308, N2214, N637);
nor NOR4 (N3795, N3769, N1554, N3365, N1975);
nor NOR2 (N3796, N3790, N1022);
buf BUF1 (N3797, N3789);
nand NAND3 (N3798, N3796, N3389, N2029);
or OR2 (N3799, N3777, N1330);
buf BUF1 (N3800, N3792);
buf BUF1 (N3801, N3793);
nor NOR3 (N3802, N3797, N1577, N2388);
xor XOR2 (N3803, N3798, N651);
xor XOR2 (N3804, N3773, N1084);
nor NOR4 (N3805, N3801, N2456, N703, N343);
or OR4 (N3806, N3805, N787, N1492, N982);
nand NAND4 (N3807, N3794, N2952, N3279, N2454);
not NOT1 (N3808, N3800);
buf BUF1 (N3809, N3802);
buf BUF1 (N3810, N3809);
nand NAND2 (N3811, N3808, N2635);
not NOT1 (N3812, N3791);
or OR4 (N3813, N3811, N854, N1310, N2629);
nand NAND3 (N3814, N3812, N3139, N3129);
xor XOR2 (N3815, N3795, N2251);
nand NAND3 (N3816, N3799, N1656, N1153);
or OR2 (N3817, N3783, N637);
buf BUF1 (N3818, N3804);
xor XOR2 (N3819, N3815, N3557);
and AND3 (N3820, N3819, N1895, N1764);
nor NOR2 (N3821, N3814, N1617);
buf BUF1 (N3822, N3817);
xor XOR2 (N3823, N3803, N928);
not NOT1 (N3824, N3810);
not NOT1 (N3825, N3821);
xor XOR2 (N3826, N3820, N1977);
nand NAND2 (N3827, N3824, N1700);
and AND3 (N3828, N3807, N1225, N432);
not NOT1 (N3829, N3826);
not NOT1 (N3830, N3818);
or OR2 (N3831, N3806, N2370);
or OR4 (N3832, N3828, N1876, N1520, N169);
nor NOR3 (N3833, N3831, N2112, N3232);
buf BUF1 (N3834, N3830);
nor NOR4 (N3835, N3833, N2718, N2930, N2718);
and AND3 (N3836, N3823, N3045, N2720);
not NOT1 (N3837, N3827);
nor NOR3 (N3838, N3832, N2132, N1981);
and AND2 (N3839, N3825, N1979);
not NOT1 (N3840, N3829);
and AND4 (N3841, N3837, N1595, N163, N3378);
nand NAND3 (N3842, N3841, N3277, N1160);
not NOT1 (N3843, N3840);
and AND4 (N3844, N3834, N1407, N2327, N2057);
and AND2 (N3845, N3816, N1260);
nor NOR2 (N3846, N3813, N2464);
xor XOR2 (N3847, N3838, N1645);
xor XOR2 (N3848, N3822, N292);
xor XOR2 (N3849, N3843, N3407);
and AND3 (N3850, N3844, N319, N268);
nand NAND2 (N3851, N3839, N2781);
buf BUF1 (N3852, N3845);
nand NAND3 (N3853, N3847, N2863, N1948);
nand NAND4 (N3854, N3852, N819, N3391, N3583);
and AND2 (N3855, N3848, N1951);
nor NOR3 (N3856, N3855, N2849, N3256);
xor XOR2 (N3857, N3849, N1916);
and AND2 (N3858, N3850, N2014);
buf BUF1 (N3859, N3854);
buf BUF1 (N3860, N3846);
or OR2 (N3861, N3856, N2481);
and AND3 (N3862, N3859, N3422, N3281);
not NOT1 (N3863, N3861);
nor NOR2 (N3864, N3853, N2046);
buf BUF1 (N3865, N3835);
not NOT1 (N3866, N3842);
not NOT1 (N3867, N3863);
not NOT1 (N3868, N3860);
buf BUF1 (N3869, N3862);
nand NAND4 (N3870, N3864, N1359, N1983, N1947);
nor NOR2 (N3871, N3857, N3374);
and AND4 (N3872, N3858, N1594, N660, N318);
nand NAND4 (N3873, N3867, N3205, N513, N143);
buf BUF1 (N3874, N3866);
xor XOR2 (N3875, N3873, N2827);
nor NOR3 (N3876, N3869, N2809, N490);
nand NAND2 (N3877, N3870, N1566);
nand NAND3 (N3878, N3872, N886, N3286);
and AND3 (N3879, N3865, N2074, N68);
buf BUF1 (N3880, N3874);
not NOT1 (N3881, N3879);
nor NOR4 (N3882, N3868, N145, N2027, N2755);
and AND4 (N3883, N3851, N1870, N472, N1560);
not NOT1 (N3884, N3881);
or OR3 (N3885, N3875, N43, N1789);
or OR2 (N3886, N3877, N241);
or OR3 (N3887, N3878, N1324, N1222);
not NOT1 (N3888, N3871);
nand NAND4 (N3889, N3880, N3333, N1608, N1816);
and AND2 (N3890, N3884, N3786);
buf BUF1 (N3891, N3888);
and AND2 (N3892, N3885, N2519);
nand NAND4 (N3893, N3836, N2865, N2777, N1552);
buf BUF1 (N3894, N3889);
or OR3 (N3895, N3886, N1520, N2444);
xor XOR2 (N3896, N3894, N992);
nor NOR3 (N3897, N3882, N268, N467);
nor NOR4 (N3898, N3891, N773, N2457, N206);
nand NAND4 (N3899, N3876, N1342, N3400, N730);
or OR3 (N3900, N3887, N1168, N3705);
xor XOR2 (N3901, N3893, N1912);
nand NAND3 (N3902, N3890, N2692, N2703);
and AND4 (N3903, N3901, N202, N1814, N2936);
nand NAND3 (N3904, N3892, N1508, N3620);
buf BUF1 (N3905, N3900);
not NOT1 (N3906, N3905);
nor NOR2 (N3907, N3896, N2185);
xor XOR2 (N3908, N3899, N2654);
nor NOR4 (N3909, N3897, N2526, N3094, N3112);
xor XOR2 (N3910, N3883, N1222);
not NOT1 (N3911, N3904);
or OR3 (N3912, N3898, N2566, N1182);
buf BUF1 (N3913, N3903);
buf BUF1 (N3914, N3895);
xor XOR2 (N3915, N3911, N3317);
and AND3 (N3916, N3915, N2420, N3000);
and AND4 (N3917, N3913, N2030, N1721, N393);
buf BUF1 (N3918, N3916);
nand NAND4 (N3919, N3909, N3194, N2659, N1756);
nor NOR4 (N3920, N3908, N1272, N1891, N2857);
not NOT1 (N3921, N3919);
nand NAND3 (N3922, N3920, N2085, N1403);
and AND4 (N3923, N3922, N1268, N2456, N3476);
and AND2 (N3924, N3906, N1339);
nand NAND4 (N3925, N3924, N401, N3263, N3806);
not NOT1 (N3926, N3917);
nor NOR4 (N3927, N3918, N1237, N1370, N3817);
nor NOR3 (N3928, N3902, N143, N3007);
or OR3 (N3929, N3914, N3000, N77);
nand NAND2 (N3930, N3907, N339);
buf BUF1 (N3931, N3927);
and AND3 (N3932, N3926, N1523, N2200);
or OR4 (N3933, N3928, N2813, N2436, N1815);
or OR3 (N3934, N3929, N1235, N1614);
not NOT1 (N3935, N3912);
xor XOR2 (N3936, N3931, N1669);
buf BUF1 (N3937, N3932);
xor XOR2 (N3938, N3935, N3118);
and AND2 (N3939, N3937, N3596);
buf BUF1 (N3940, N3921);
or OR3 (N3941, N3933, N142, N173);
or OR3 (N3942, N3930, N296, N3630);
not NOT1 (N3943, N3936);
not NOT1 (N3944, N3938);
nand NAND3 (N3945, N3923, N395, N2121);
and AND2 (N3946, N3945, N3063);
and AND2 (N3947, N3944, N3336);
buf BUF1 (N3948, N3934);
xor XOR2 (N3949, N3941, N840);
nand NAND4 (N3950, N3948, N3145, N2365, N3242);
xor XOR2 (N3951, N3943, N1617);
nor NOR4 (N3952, N3951, N2802, N1484, N3192);
buf BUF1 (N3953, N3910);
nand NAND3 (N3954, N3925, N3098, N2327);
nor NOR3 (N3955, N3940, N256, N3843);
nor NOR4 (N3956, N3953, N1967, N3866, N2755);
buf BUF1 (N3957, N3954);
not NOT1 (N3958, N3952);
nand NAND2 (N3959, N3946, N3487);
not NOT1 (N3960, N3950);
nor NOR4 (N3961, N3958, N1476, N3500, N2315);
buf BUF1 (N3962, N3960);
not NOT1 (N3963, N3947);
nor NOR3 (N3964, N3939, N2281, N1357);
buf BUF1 (N3965, N3962);
nor NOR2 (N3966, N3942, N94);
buf BUF1 (N3967, N3966);
xor XOR2 (N3968, N3949, N834);
buf BUF1 (N3969, N3968);
xor XOR2 (N3970, N3957, N1553);
not NOT1 (N3971, N3970);
not NOT1 (N3972, N3956);
or OR4 (N3973, N3972, N403, N3641, N938);
and AND4 (N3974, N3967, N2099, N924, N2115);
nand NAND2 (N3975, N3971, N183);
buf BUF1 (N3976, N3963);
and AND2 (N3977, N3965, N3398);
buf BUF1 (N3978, N3969);
not NOT1 (N3979, N3975);
xor XOR2 (N3980, N3977, N2954);
buf BUF1 (N3981, N3964);
nand NAND4 (N3982, N3961, N1831, N2024, N2557);
and AND3 (N3983, N3955, N52, N1897);
nand NAND4 (N3984, N3959, N1616, N3231, N749);
not NOT1 (N3985, N3981);
or OR4 (N3986, N3983, N178, N3780, N2483);
nor NOR3 (N3987, N3978, N3103, N3659);
buf BUF1 (N3988, N3980);
nand NAND4 (N3989, N3986, N3462, N307, N2857);
not NOT1 (N3990, N3982);
xor XOR2 (N3991, N3989, N3967);
and AND2 (N3992, N3987, N1036);
or OR2 (N3993, N3988, N3169);
nor NOR4 (N3994, N3973, N1591, N318, N3579);
or OR3 (N3995, N3976, N1502, N3603);
xor XOR2 (N3996, N3991, N2531);
nor NOR3 (N3997, N3974, N3305, N691);
and AND3 (N3998, N3993, N2183, N2391);
not NOT1 (N3999, N3984);
buf BUF1 (N4000, N3994);
nand NAND2 (N4001, N3979, N1414);
or OR3 (N4002, N4000, N1915, N723);
nand NAND4 (N4003, N3998, N422, N3254, N2761);
buf BUF1 (N4004, N3999);
nand NAND3 (N4005, N3995, N1729, N1717);
or OR4 (N4006, N4004, N80, N541, N2095);
xor XOR2 (N4007, N3996, N2507);
or OR2 (N4008, N4001, N436);
buf BUF1 (N4009, N4007);
and AND2 (N4010, N4008, N58);
buf BUF1 (N4011, N3985);
not NOT1 (N4012, N4003);
nand NAND3 (N4013, N4011, N1293, N769);
xor XOR2 (N4014, N4013, N3443);
buf BUF1 (N4015, N4009);
nor NOR2 (N4016, N4010, N1927);
and AND2 (N4017, N4006, N3192);
and AND4 (N4018, N4015, N3400, N2030, N2498);
buf BUF1 (N4019, N4014);
xor XOR2 (N4020, N4019, N848);
xor XOR2 (N4021, N4016, N795);
or OR4 (N4022, N3990, N2336, N2928, N2850);
xor XOR2 (N4023, N4012, N1754);
not NOT1 (N4024, N3997);
buf BUF1 (N4025, N4018);
xor XOR2 (N4026, N4021, N426);
xor XOR2 (N4027, N4026, N3103);
not NOT1 (N4028, N4022);
not NOT1 (N4029, N4002);
not NOT1 (N4030, N4025);
not NOT1 (N4031, N3992);
and AND4 (N4032, N4031, N378, N3874, N1985);
nand NAND3 (N4033, N4020, N1708, N2409);
not NOT1 (N4034, N4024);
not NOT1 (N4035, N4017);
not NOT1 (N4036, N4035);
nand NAND4 (N4037, N4005, N1095, N2742, N2458);
buf BUF1 (N4038, N4027);
nor NOR2 (N4039, N4032, N381);
or OR2 (N4040, N4030, N1958);
nand NAND3 (N4041, N4039, N497, N1508);
and AND4 (N4042, N4034, N2438, N2431, N2395);
and AND3 (N4043, N4033, N236, N2268);
nand NAND3 (N4044, N4028, N255, N2404);
nand NAND4 (N4045, N4040, N2992, N3354, N1095);
nor NOR2 (N4046, N4042, N2291);
and AND4 (N4047, N4044, N3654, N273, N1584);
buf BUF1 (N4048, N4043);
buf BUF1 (N4049, N4041);
and AND4 (N4050, N4047, N2232, N2116, N1639);
buf BUF1 (N4051, N4046);
nor NOR2 (N4052, N4029, N3466);
buf BUF1 (N4053, N4038);
buf BUF1 (N4054, N4051);
not NOT1 (N4055, N4023);
nand NAND2 (N4056, N4050, N3614);
not NOT1 (N4057, N4054);
buf BUF1 (N4058, N4057);
not NOT1 (N4059, N4049);
not NOT1 (N4060, N4045);
and AND4 (N4061, N4059, N2673, N1188, N3355);
buf BUF1 (N4062, N4053);
buf BUF1 (N4063, N4037);
and AND2 (N4064, N4048, N3153);
not NOT1 (N4065, N4036);
nor NOR3 (N4066, N4060, N3169, N2658);
buf BUF1 (N4067, N4065);
xor XOR2 (N4068, N4058, N330);
xor XOR2 (N4069, N4055, N2530);
and AND3 (N4070, N4056, N4008, N3485);
buf BUF1 (N4071, N4068);
nor NOR2 (N4072, N4070, N46);
and AND3 (N4073, N4062, N1552, N1497);
and AND3 (N4074, N4073, N1610, N2766);
buf BUF1 (N4075, N4063);
xor XOR2 (N4076, N4071, N1813);
nor NOR3 (N4077, N4061, N853, N1919);
and AND2 (N4078, N4074, N2336);
not NOT1 (N4079, N4064);
xor XOR2 (N4080, N4078, N1421);
and AND4 (N4081, N4079, N1352, N3079, N402);
and AND3 (N4082, N4076, N1704, N2636);
not NOT1 (N4083, N4072);
nand NAND3 (N4084, N4066, N4073, N2208);
or OR4 (N4085, N4082, N2307, N2653, N615);
or OR2 (N4086, N4085, N3772);
and AND3 (N4087, N4086, N2014, N4004);
not NOT1 (N4088, N4081);
and AND2 (N4089, N4077, N2467);
xor XOR2 (N4090, N4075, N575);
nor NOR3 (N4091, N4052, N232, N743);
xor XOR2 (N4092, N4080, N3597);
nand NAND4 (N4093, N4090, N3278, N322, N2290);
not NOT1 (N4094, N4067);
nor NOR4 (N4095, N4088, N3437, N3156, N3772);
or OR3 (N4096, N4094, N3484, N1879);
xor XOR2 (N4097, N4084, N327);
nand NAND2 (N4098, N4089, N2895);
nor NOR3 (N4099, N4095, N3217, N2578);
nand NAND2 (N4100, N4093, N2872);
xor XOR2 (N4101, N4092, N2352);
not NOT1 (N4102, N4096);
and AND3 (N4103, N4069, N2611, N171);
nand NAND4 (N4104, N4083, N450, N1045, N362);
nand NAND3 (N4105, N4098, N191, N3776);
nor NOR2 (N4106, N4087, N3073);
nand NAND2 (N4107, N4097, N2997);
nor NOR4 (N4108, N4105, N259, N2712, N3992);
xor XOR2 (N4109, N4102, N44);
not NOT1 (N4110, N4106);
and AND3 (N4111, N4099, N3110, N1409);
buf BUF1 (N4112, N4110);
not NOT1 (N4113, N4103);
buf BUF1 (N4114, N4113);
not NOT1 (N4115, N4111);
xor XOR2 (N4116, N4112, N2896);
nor NOR2 (N4117, N4114, N955);
or OR2 (N4118, N4101, N2961);
xor XOR2 (N4119, N4109, N3397);
and AND2 (N4120, N4108, N1290);
buf BUF1 (N4121, N4107);
or OR2 (N4122, N4115, N2272);
buf BUF1 (N4123, N4119);
nand NAND2 (N4124, N4122, N3912);
not NOT1 (N4125, N4116);
and AND2 (N4126, N4091, N3029);
nand NAND4 (N4127, N4118, N2630, N2826, N1343);
and AND4 (N4128, N4100, N1600, N3899, N592);
nand NAND2 (N4129, N4124, N1869);
buf BUF1 (N4130, N4123);
and AND2 (N4131, N4129, N3607);
nor NOR4 (N4132, N4121, N2206, N1676, N1233);
or OR4 (N4133, N4117, N1892, N2204, N106);
or OR3 (N4134, N4127, N2682, N2349);
or OR2 (N4135, N4131, N1438);
not NOT1 (N4136, N4126);
or OR4 (N4137, N4130, N2726, N425, N3572);
buf BUF1 (N4138, N4135);
or OR4 (N4139, N4138, N3994, N3835, N770);
or OR4 (N4140, N4137, N2204, N1203, N1612);
nand NAND3 (N4141, N4104, N2446, N3870);
xor XOR2 (N4142, N4134, N185);
buf BUF1 (N4143, N4128);
xor XOR2 (N4144, N4120, N1039);
buf BUF1 (N4145, N4139);
nor NOR2 (N4146, N4132, N1854);
and AND3 (N4147, N4144, N1503, N2417);
nand NAND3 (N4148, N4136, N3130, N2612);
nand NAND2 (N4149, N4145, N1868);
not NOT1 (N4150, N4143);
xor XOR2 (N4151, N4142, N434);
buf BUF1 (N4152, N4150);
nand NAND2 (N4153, N4140, N3517);
not NOT1 (N4154, N4141);
and AND4 (N4155, N4151, N571, N1826, N2111);
xor XOR2 (N4156, N4146, N1354);
not NOT1 (N4157, N4148);
not NOT1 (N4158, N4149);
nand NAND3 (N4159, N4158, N993, N3086);
buf BUF1 (N4160, N4125);
nand NAND3 (N4161, N4155, N1863, N2776);
or OR2 (N4162, N4160, N957);
and AND2 (N4163, N4159, N4113);
not NOT1 (N4164, N4154);
not NOT1 (N4165, N4163);
nor NOR3 (N4166, N4147, N3745, N2102);
or OR2 (N4167, N4156, N3221);
xor XOR2 (N4168, N4162, N686);
buf BUF1 (N4169, N4165);
or OR4 (N4170, N4164, N46, N1779, N1062);
xor XOR2 (N4171, N4168, N2927);
buf BUF1 (N4172, N4166);
nor NOR2 (N4173, N4152, N3716);
nor NOR4 (N4174, N4167, N3852, N3428, N663);
xor XOR2 (N4175, N4161, N1782);
and AND4 (N4176, N4174, N775, N210, N863);
buf BUF1 (N4177, N4176);
or OR4 (N4178, N4172, N2798, N2165, N810);
nor NOR3 (N4179, N4171, N3309, N1423);
not NOT1 (N4180, N4169);
nor NOR4 (N4181, N4133, N756, N2995, N3670);
xor XOR2 (N4182, N4153, N2381);
or OR2 (N4183, N4177, N3522);
not NOT1 (N4184, N4182);
xor XOR2 (N4185, N4157, N477);
nand NAND4 (N4186, N4178, N2666, N2932, N635);
nand NAND4 (N4187, N4180, N2816, N1484, N3985);
xor XOR2 (N4188, N4183, N1503);
buf BUF1 (N4189, N4185);
and AND3 (N4190, N4170, N2745, N1763);
buf BUF1 (N4191, N4187);
nor NOR2 (N4192, N4189, N30);
or OR2 (N4193, N4191, N2983);
nor NOR3 (N4194, N4186, N1741, N3639);
and AND2 (N4195, N4173, N2849);
nor NOR3 (N4196, N4190, N242, N989);
buf BUF1 (N4197, N4195);
and AND2 (N4198, N4196, N1826);
nand NAND3 (N4199, N4179, N1684, N1757);
or OR3 (N4200, N4184, N1162, N1755);
nand NAND4 (N4201, N4198, N4190, N3319, N1049);
xor XOR2 (N4202, N4200, N1104);
buf BUF1 (N4203, N4199);
nor NOR4 (N4204, N4188, N3563, N2930, N2672);
nand NAND3 (N4205, N4175, N2265, N2279);
or OR3 (N4206, N4202, N2165, N2293);
nor NOR4 (N4207, N4204, N2924, N247, N3173);
xor XOR2 (N4208, N4193, N3087);
and AND2 (N4209, N4206, N619);
and AND4 (N4210, N4207, N135, N2259, N1205);
buf BUF1 (N4211, N4201);
buf BUF1 (N4212, N4209);
and AND2 (N4213, N4211, N2327);
and AND3 (N4214, N4197, N1067, N3763);
nor NOR4 (N4215, N4208, N98, N2742, N4070);
buf BUF1 (N4216, N4205);
and AND2 (N4217, N4210, N3704);
or OR4 (N4218, N4194, N2877, N543, N3049);
and AND2 (N4219, N4214, N1019);
nand NAND2 (N4220, N4216, N3725);
buf BUF1 (N4221, N4212);
nor NOR2 (N4222, N4192, N1233);
or OR2 (N4223, N4181, N777);
nor NOR3 (N4224, N4220, N1679, N3737);
xor XOR2 (N4225, N4203, N3596);
buf BUF1 (N4226, N4223);
not NOT1 (N4227, N4218);
nor NOR2 (N4228, N4221, N417);
and AND3 (N4229, N4226, N3450, N1361);
nor NOR2 (N4230, N4225, N4067);
xor XOR2 (N4231, N4215, N1462);
buf BUF1 (N4232, N4228);
nor NOR3 (N4233, N4227, N564, N231);
xor XOR2 (N4234, N4224, N1153);
nor NOR2 (N4235, N4219, N463);
nor NOR4 (N4236, N4213, N2780, N2113, N2899);
nor NOR3 (N4237, N4234, N1517, N1883);
xor XOR2 (N4238, N4236, N846);
nor NOR4 (N4239, N4237, N1411, N543, N2588);
buf BUF1 (N4240, N4230);
and AND4 (N4241, N4235, N2674, N1193, N3659);
and AND4 (N4242, N4239, N886, N729, N3444);
not NOT1 (N4243, N4229);
and AND4 (N4244, N4231, N289, N2422, N3367);
and AND4 (N4245, N4233, N3806, N2570, N3578);
nor NOR4 (N4246, N4241, N439, N920, N2900);
not NOT1 (N4247, N4240);
nor NOR3 (N4248, N4245, N3768, N1910);
buf BUF1 (N4249, N4242);
xor XOR2 (N4250, N4232, N3593);
and AND2 (N4251, N4238, N3998);
nor NOR4 (N4252, N4249, N1091, N1570, N1637);
and AND3 (N4253, N4252, N790, N965);
xor XOR2 (N4254, N4253, N3017);
nor NOR2 (N4255, N4248, N3855);
buf BUF1 (N4256, N4217);
not NOT1 (N4257, N4244);
xor XOR2 (N4258, N4251, N2076);
not NOT1 (N4259, N4222);
nor NOR3 (N4260, N4257, N4000, N2432);
and AND4 (N4261, N4250, N1240, N3423, N1623);
nand NAND2 (N4262, N4255, N1895);
nor NOR4 (N4263, N4261, N2901, N3906, N3614);
nand NAND2 (N4264, N4254, N4036);
or OR4 (N4265, N4258, N406, N2100, N1239);
and AND4 (N4266, N4243, N4137, N793, N4222);
and AND2 (N4267, N4246, N2952);
buf BUF1 (N4268, N4264);
or OR2 (N4269, N4256, N1732);
not NOT1 (N4270, N4259);
or OR2 (N4271, N4266, N2709);
not NOT1 (N4272, N4271);
and AND2 (N4273, N4260, N2327);
not NOT1 (N4274, N4268);
and AND3 (N4275, N4265, N2800, N168);
not NOT1 (N4276, N4269);
not NOT1 (N4277, N4272);
or OR3 (N4278, N4274, N3172, N4036);
not NOT1 (N4279, N4275);
or OR2 (N4280, N4276, N3286);
nand NAND2 (N4281, N4263, N1330);
nand NAND3 (N4282, N4270, N162, N1466);
nand NAND2 (N4283, N4267, N2567);
nand NAND2 (N4284, N4247, N3984);
buf BUF1 (N4285, N4281);
nor NOR4 (N4286, N4279, N282, N3934, N2472);
not NOT1 (N4287, N4286);
buf BUF1 (N4288, N4285);
xor XOR2 (N4289, N4283, N3945);
not NOT1 (N4290, N4280);
nand NAND3 (N4291, N4289, N1678, N1246);
nor NOR4 (N4292, N4287, N1875, N1424, N4199);
nor NOR2 (N4293, N4282, N1634);
buf BUF1 (N4294, N4292);
nor NOR3 (N4295, N4294, N586, N2646);
nand NAND2 (N4296, N4288, N2316);
buf BUF1 (N4297, N4295);
xor XOR2 (N4298, N4290, N1209);
nor NOR2 (N4299, N4291, N3408);
nor NOR3 (N4300, N4296, N4103, N3265);
and AND2 (N4301, N4293, N393);
not NOT1 (N4302, N4273);
or OR4 (N4303, N4301, N1300, N593, N2560);
or OR4 (N4304, N4278, N3243, N3773, N3777);
and AND2 (N4305, N4298, N2175);
nand NAND4 (N4306, N4299, N392, N4015, N1844);
xor XOR2 (N4307, N4300, N1172);
not NOT1 (N4308, N4262);
nor NOR3 (N4309, N4307, N1198, N2251);
nand NAND2 (N4310, N4302, N3428);
buf BUF1 (N4311, N4297);
or OR4 (N4312, N4303, N1228, N2006, N824);
not NOT1 (N4313, N4305);
not NOT1 (N4314, N4313);
and AND4 (N4315, N4310, N44, N1272, N1021);
nand NAND3 (N4316, N4284, N3800, N1026);
not NOT1 (N4317, N4316);
buf BUF1 (N4318, N4312);
buf BUF1 (N4319, N4318);
buf BUF1 (N4320, N4277);
not NOT1 (N4321, N4304);
xor XOR2 (N4322, N4306, N4281);
or OR2 (N4323, N4311, N1669);
not NOT1 (N4324, N4315);
nor NOR2 (N4325, N4317, N908);
buf BUF1 (N4326, N4324);
nand NAND2 (N4327, N4325, N696);
not NOT1 (N4328, N4314);
xor XOR2 (N4329, N4328, N2181);
buf BUF1 (N4330, N4308);
and AND4 (N4331, N4329, N3817, N4017, N2422);
xor XOR2 (N4332, N4321, N3322);
nor NOR4 (N4333, N4320, N743, N813, N2390);
or OR2 (N4334, N4332, N2828);
nand NAND4 (N4335, N4322, N245, N4319, N2167);
xor XOR2 (N4336, N1504, N4327);
and AND3 (N4337, N2265, N2083, N322);
buf BUF1 (N4338, N4331);
buf BUF1 (N4339, N4309);
nand NAND2 (N4340, N4330, N2087);
not NOT1 (N4341, N4338);
buf BUF1 (N4342, N4334);
not NOT1 (N4343, N4342);
nand NAND4 (N4344, N4323, N1132, N636, N523);
buf BUF1 (N4345, N4340);
nand NAND3 (N4346, N4336, N2772, N2056);
or OR4 (N4347, N4335, N2545, N1810, N3122);
buf BUF1 (N4348, N4346);
and AND3 (N4349, N4339, N302, N3241);
nor NOR3 (N4350, N4347, N3968, N1063);
xor XOR2 (N4351, N4350, N4036);
buf BUF1 (N4352, N4348);
or OR3 (N4353, N4337, N237, N224);
not NOT1 (N4354, N4341);
xor XOR2 (N4355, N4326, N532);
nand NAND2 (N4356, N4353, N1959);
nand NAND2 (N4357, N4354, N2397);
and AND2 (N4358, N4352, N2462);
xor XOR2 (N4359, N4356, N1542);
not NOT1 (N4360, N4344);
xor XOR2 (N4361, N4351, N3337);
and AND2 (N4362, N4358, N2143);
nand NAND2 (N4363, N4349, N1135);
nand NAND3 (N4364, N4357, N3354, N1901);
nand NAND3 (N4365, N4345, N3569, N839);
or OR4 (N4366, N4362, N3772, N2485, N1855);
nor NOR4 (N4367, N4365, N2800, N1740, N2442);
buf BUF1 (N4368, N4364);
nand NAND2 (N4369, N4359, N1965);
xor XOR2 (N4370, N4361, N2875);
xor XOR2 (N4371, N4360, N1183);
not NOT1 (N4372, N4369);
and AND2 (N4373, N4333, N2319);
or OR3 (N4374, N4366, N2421, N809);
not NOT1 (N4375, N4355);
buf BUF1 (N4376, N4367);
nand NAND4 (N4377, N4368, N233, N4332, N1370);
not NOT1 (N4378, N4375);
buf BUF1 (N4379, N4363);
nor NOR4 (N4380, N4372, N149, N1825, N4171);
xor XOR2 (N4381, N4370, N3752);
buf BUF1 (N4382, N4376);
or OR4 (N4383, N4374, N272, N737, N2229);
xor XOR2 (N4384, N4371, N72);
not NOT1 (N4385, N4380);
not NOT1 (N4386, N4382);
and AND3 (N4387, N4379, N3466, N495);
xor XOR2 (N4388, N4373, N2269);
nand NAND4 (N4389, N4377, N4313, N356, N2216);
not NOT1 (N4390, N4387);
or OR2 (N4391, N4386, N4384);
xor XOR2 (N4392, N3886, N1730);
and AND4 (N4393, N4343, N2062, N2317, N873);
or OR4 (N4394, N4389, N1976, N1609, N792);
and AND4 (N4395, N4385, N367, N2821, N4249);
and AND4 (N4396, N4392, N1775, N3533, N2179);
xor XOR2 (N4397, N4390, N3971);
buf BUF1 (N4398, N4388);
not NOT1 (N4399, N4393);
xor XOR2 (N4400, N4378, N1189);
buf BUF1 (N4401, N4395);
or OR4 (N4402, N4396, N1870, N3919, N2735);
xor XOR2 (N4403, N4399, N3432);
xor XOR2 (N4404, N4394, N761);
nand NAND2 (N4405, N4400, N1621);
and AND3 (N4406, N4383, N484, N576);
buf BUF1 (N4407, N4381);
nor NOR4 (N4408, N4397, N736, N1571, N127);
buf BUF1 (N4409, N4391);
xor XOR2 (N4410, N4409, N1827);
buf BUF1 (N4411, N4406);
buf BUF1 (N4412, N4405);
nand NAND3 (N4413, N4408, N838, N2925);
nand NAND3 (N4414, N4402, N2143, N4392);
nor NOR2 (N4415, N4401, N3572);
nor NOR3 (N4416, N4403, N1456, N411);
not NOT1 (N4417, N4411);
or OR4 (N4418, N4407, N1213, N557, N582);
or OR2 (N4419, N4414, N3602);
buf BUF1 (N4420, N4410);
or OR4 (N4421, N4417, N275, N4139, N1438);
not NOT1 (N4422, N4419);
nand NAND3 (N4423, N4398, N807, N3669);
nand NAND3 (N4424, N4418, N1344, N3749);
nand NAND2 (N4425, N4412, N577);
not NOT1 (N4426, N4425);
and AND4 (N4427, N4426, N1313, N2627, N4166);
nand NAND3 (N4428, N4424, N3491, N752);
xor XOR2 (N4429, N4422, N2449);
or OR4 (N4430, N4415, N1100, N4288, N1885);
not NOT1 (N4431, N4423);
nand NAND2 (N4432, N4430, N242);
not NOT1 (N4433, N4404);
not NOT1 (N4434, N4433);
and AND3 (N4435, N4421, N116, N2068);
nand NAND4 (N4436, N4434, N846, N2556, N3076);
or OR2 (N4437, N4432, N1303);
nor NOR4 (N4438, N4436, N3125, N2112, N733);
not NOT1 (N4439, N4413);
or OR2 (N4440, N4416, N323);
buf BUF1 (N4441, N4437);
not NOT1 (N4442, N4429);
nand NAND2 (N4443, N4438, N4146);
xor XOR2 (N4444, N4431, N2045);
nand NAND4 (N4445, N4428, N3126, N3977, N4073);
xor XOR2 (N4446, N4443, N4063);
nand NAND4 (N4447, N4420, N2090, N2354, N3351);
and AND2 (N4448, N4445, N2928);
buf BUF1 (N4449, N4435);
buf BUF1 (N4450, N4427);
or OR3 (N4451, N4448, N2553, N752);
xor XOR2 (N4452, N4441, N1118);
nand NAND2 (N4453, N4452, N2226);
xor XOR2 (N4454, N4453, N4059);
nand NAND4 (N4455, N4442, N1176, N394, N113);
or OR4 (N4456, N4447, N2827, N3890, N1564);
buf BUF1 (N4457, N4454);
nor NOR3 (N4458, N4444, N3134, N3890);
nand NAND2 (N4459, N4456, N3331);
buf BUF1 (N4460, N4458);
and AND4 (N4461, N4439, N1255, N384, N2742);
xor XOR2 (N4462, N4461, N3861);
and AND4 (N4463, N4451, N3207, N4343, N2605);
and AND3 (N4464, N4440, N4274, N3963);
buf BUF1 (N4465, N4449);
nor NOR4 (N4466, N4457, N3290, N1942, N2399);
buf BUF1 (N4467, N4465);
nand NAND4 (N4468, N4450, N2493, N2035, N4079);
nand NAND4 (N4469, N4468, N1664, N1335, N3174);
nand NAND2 (N4470, N4466, N3224);
xor XOR2 (N4471, N4446, N1099);
and AND2 (N4472, N4459, N1009);
xor XOR2 (N4473, N4467, N556);
buf BUF1 (N4474, N4460);
nor NOR4 (N4475, N4471, N1749, N558, N709);
buf BUF1 (N4476, N4475);
not NOT1 (N4477, N4455);
not NOT1 (N4478, N4469);
and AND3 (N4479, N4476, N2292, N1838);
or OR3 (N4480, N4473, N383, N326);
nor NOR3 (N4481, N4470, N3714, N1873);
and AND4 (N4482, N4480, N1747, N4233, N4224);
and AND3 (N4483, N4479, N1758, N729);
nor NOR4 (N4484, N4464, N2329, N4478, N1285);
and AND4 (N4485, N774, N3669, N1639, N55);
not NOT1 (N4486, N4483);
nand NAND2 (N4487, N4486, N4059);
nor NOR3 (N4488, N4474, N359, N2899);
nor NOR2 (N4489, N4481, N3180);
xor XOR2 (N4490, N4484, N1936);
nor NOR2 (N4491, N4488, N173);
buf BUF1 (N4492, N4485);
or OR3 (N4493, N4491, N3634, N1961);
not NOT1 (N4494, N4492);
xor XOR2 (N4495, N4482, N2420);
buf BUF1 (N4496, N4489);
not NOT1 (N4497, N4493);
and AND4 (N4498, N4495, N1097, N1804, N1741);
or OR2 (N4499, N4494, N3139);
nor NOR4 (N4500, N4477, N2639, N2695, N886);
buf BUF1 (N4501, N4500);
nand NAND4 (N4502, N4497, N4112, N1923, N1002);
nand NAND4 (N4503, N4502, N720, N4436, N846);
nand NAND4 (N4504, N4496, N2534, N2610, N913);
buf BUF1 (N4505, N4503);
xor XOR2 (N4506, N4462, N687);
xor XOR2 (N4507, N4463, N1993);
buf BUF1 (N4508, N4498);
nand NAND3 (N4509, N4501, N2754, N1477);
and AND3 (N4510, N4472, N3227, N3868);
nand NAND4 (N4511, N4506, N1920, N2357, N3467);
buf BUF1 (N4512, N4511);
nor NOR2 (N4513, N4509, N1179);
or OR4 (N4514, N4508, N3360, N2589, N2272);
not NOT1 (N4515, N4505);
not NOT1 (N4516, N4487);
buf BUF1 (N4517, N4504);
nor NOR4 (N4518, N4513, N3818, N2566, N3451);
xor XOR2 (N4519, N4510, N4035);
nand NAND3 (N4520, N4507, N2227, N3693);
not NOT1 (N4521, N4517);
or OR4 (N4522, N4512, N2322, N4519, N191);
and AND3 (N4523, N2862, N2651, N4364);
or OR3 (N4524, N4520, N3186, N2888);
or OR3 (N4525, N4524, N4143, N345);
not NOT1 (N4526, N4518);
buf BUF1 (N4527, N4521);
or OR3 (N4528, N4522, N1290, N3871);
buf BUF1 (N4529, N4523);
nor NOR3 (N4530, N4514, N1627, N2457);
not NOT1 (N4531, N4516);
nor NOR2 (N4532, N4525, N1546);
or OR2 (N4533, N4529, N136);
nor NOR4 (N4534, N4533, N377, N3712, N3850);
nand NAND2 (N4535, N4534, N4340);
buf BUF1 (N4536, N4532);
or OR4 (N4537, N4499, N1622, N1586, N727);
or OR4 (N4538, N4528, N2532, N230, N238);
and AND2 (N4539, N4536, N1527);
nand NAND3 (N4540, N4530, N2173, N4054);
or OR2 (N4541, N4526, N2623);
or OR4 (N4542, N4540, N3624, N2379, N3672);
nor NOR2 (N4543, N4537, N2190);
nor NOR3 (N4544, N4542, N2273, N2616);
xor XOR2 (N4545, N4535, N248);
nand NAND4 (N4546, N4541, N1797, N1892, N1346);
buf BUF1 (N4547, N4538);
nor NOR3 (N4548, N4544, N3640, N3977);
nand NAND4 (N4549, N4546, N123, N20, N4195);
buf BUF1 (N4550, N4547);
buf BUF1 (N4551, N4550);
buf BUF1 (N4552, N4551);
xor XOR2 (N4553, N4515, N2453);
or OR4 (N4554, N4490, N718, N1381, N2599);
nor NOR4 (N4555, N4527, N4190, N3145, N4035);
buf BUF1 (N4556, N4545);
and AND2 (N4557, N4554, N729);
nor NOR3 (N4558, N4549, N574, N81);
buf BUF1 (N4559, N4558);
not NOT1 (N4560, N4555);
xor XOR2 (N4561, N4560, N1486);
or OR2 (N4562, N4531, N2321);
nor NOR2 (N4563, N4539, N1619);
nor NOR2 (N4564, N4561, N2416);
or OR3 (N4565, N4548, N4548, N1317);
and AND4 (N4566, N4564, N3244, N4253, N2188);
not NOT1 (N4567, N4559);
or OR2 (N4568, N4553, N3996);
nor NOR3 (N4569, N4567, N3531, N2084);
or OR3 (N4570, N4569, N873, N3617);
buf BUF1 (N4571, N4568);
buf BUF1 (N4572, N4562);
not NOT1 (N4573, N4571);
xor XOR2 (N4574, N4543, N3097);
and AND2 (N4575, N4557, N956);
xor XOR2 (N4576, N4563, N2175);
and AND3 (N4577, N4556, N2152, N2411);
xor XOR2 (N4578, N4570, N2550);
or OR4 (N4579, N4574, N3126, N4425, N2701);
or OR2 (N4580, N4565, N3168);
nor NOR2 (N4581, N4580, N1778);
nand NAND2 (N4582, N4566, N4497);
or OR4 (N4583, N4578, N368, N2793, N1056);
not NOT1 (N4584, N4576);
nand NAND4 (N4585, N4573, N1467, N3501, N2934);
nand NAND2 (N4586, N4572, N4437);
buf BUF1 (N4587, N4577);
buf BUF1 (N4588, N4552);
xor XOR2 (N4589, N4575, N1015);
buf BUF1 (N4590, N4586);
and AND2 (N4591, N4579, N4468);
not NOT1 (N4592, N4591);
not NOT1 (N4593, N4588);
buf BUF1 (N4594, N4590);
xor XOR2 (N4595, N4585, N290);
nor NOR3 (N4596, N4584, N3395, N1796);
and AND3 (N4597, N4582, N3462, N4409);
not NOT1 (N4598, N4581);
nand NAND3 (N4599, N4589, N3765, N4539);
or OR4 (N4600, N4587, N2763, N3273, N661);
xor XOR2 (N4601, N4598, N1458);
nand NAND2 (N4602, N4593, N2461);
or OR2 (N4603, N4583, N4185);
xor XOR2 (N4604, N4602, N268);
and AND3 (N4605, N4594, N1403, N1451);
and AND3 (N4606, N4605, N2621, N4326);
xor XOR2 (N4607, N4596, N3297);
not NOT1 (N4608, N4592);
xor XOR2 (N4609, N4604, N577);
nor NOR2 (N4610, N4603, N672);
and AND3 (N4611, N4601, N3623, N3178);
not NOT1 (N4612, N4606);
not NOT1 (N4613, N4600);
and AND3 (N4614, N4597, N2154, N3693);
nand NAND4 (N4615, N4609, N1175, N1670, N1150);
not NOT1 (N4616, N4614);
buf BUF1 (N4617, N4599);
and AND3 (N4618, N4610, N3995, N483);
nand NAND3 (N4619, N4595, N3523, N3743);
and AND2 (N4620, N4613, N3277);
nor NOR4 (N4621, N4615, N926, N4172, N4304);
nor NOR3 (N4622, N4607, N4488, N95);
nor NOR3 (N4623, N4617, N748, N2484);
nor NOR3 (N4624, N4621, N4166, N4082);
buf BUF1 (N4625, N4623);
or OR3 (N4626, N4616, N3316, N182);
xor XOR2 (N4627, N4625, N4234);
nand NAND4 (N4628, N4624, N2289, N1329, N1959);
xor XOR2 (N4629, N4612, N1825);
and AND3 (N4630, N4620, N2826, N1882);
or OR3 (N4631, N4608, N2866, N1215);
not NOT1 (N4632, N4626);
and AND2 (N4633, N4628, N534);
and AND4 (N4634, N4629, N3922, N336, N3939);
nand NAND4 (N4635, N4631, N2675, N3022, N1775);
and AND3 (N4636, N4611, N4277, N3576);
or OR4 (N4637, N4627, N1004, N4017, N3422);
and AND4 (N4638, N4634, N2136, N4147, N327);
xor XOR2 (N4639, N4630, N3470);
and AND3 (N4640, N4635, N2545, N558);
not NOT1 (N4641, N4638);
nand NAND2 (N4642, N4633, N3835);
nor NOR4 (N4643, N4619, N3749, N2235, N1898);
nor NOR4 (N4644, N4618, N1593, N392, N2023);
xor XOR2 (N4645, N4636, N1724);
or OR3 (N4646, N4632, N1324, N3489);
or OR2 (N4647, N4637, N4356);
or OR3 (N4648, N4647, N714, N4398);
buf BUF1 (N4649, N4640);
or OR4 (N4650, N4642, N4134, N3702, N2752);
or OR2 (N4651, N4641, N706);
not NOT1 (N4652, N4648);
not NOT1 (N4653, N4650);
buf BUF1 (N4654, N4652);
not NOT1 (N4655, N4643);
buf BUF1 (N4656, N4654);
not NOT1 (N4657, N4651);
not NOT1 (N4658, N4644);
xor XOR2 (N4659, N4657, N1254);
and AND2 (N4660, N4649, N3474);
xor XOR2 (N4661, N4653, N1965);
buf BUF1 (N4662, N4660);
buf BUF1 (N4663, N4639);
or OR4 (N4664, N4655, N1100, N425, N2413);
or OR2 (N4665, N4656, N1229);
nor NOR4 (N4666, N4662, N3584, N2489, N1680);
or OR4 (N4667, N4664, N741, N1315, N404);
buf BUF1 (N4668, N4667);
not NOT1 (N4669, N4665);
not NOT1 (N4670, N4658);
nor NOR3 (N4671, N4663, N1792, N2108);
buf BUF1 (N4672, N4659);
nand NAND4 (N4673, N4622, N1490, N4563, N4138);
and AND3 (N4674, N4668, N2053, N503);
nand NAND3 (N4675, N4672, N3829, N2431);
buf BUF1 (N4676, N4666);
not NOT1 (N4677, N4645);
buf BUF1 (N4678, N4675);
and AND2 (N4679, N4677, N3550);
not NOT1 (N4680, N4679);
buf BUF1 (N4681, N4678);
or OR2 (N4682, N4661, N2027);
not NOT1 (N4683, N4676);
or OR3 (N4684, N4683, N3366, N1802);
nand NAND2 (N4685, N4673, N2042);
buf BUF1 (N4686, N4684);
xor XOR2 (N4687, N4669, N1363);
xor XOR2 (N4688, N4687, N4453);
or OR4 (N4689, N4685, N4574, N468, N560);
and AND2 (N4690, N4670, N1059);
nand NAND3 (N4691, N4686, N988, N3255);
or OR2 (N4692, N4680, N1552);
buf BUF1 (N4693, N4674);
xor XOR2 (N4694, N4692, N494);
not NOT1 (N4695, N4688);
buf BUF1 (N4696, N4689);
nand NAND3 (N4697, N4681, N4555, N3687);
buf BUF1 (N4698, N4694);
or OR3 (N4699, N4697, N3879, N2718);
xor XOR2 (N4700, N4682, N73);
buf BUF1 (N4701, N4698);
nand NAND3 (N4702, N4701, N2502, N3188);
buf BUF1 (N4703, N4690);
and AND4 (N4704, N4695, N1416, N3851, N3423);
or OR3 (N4705, N4704, N2085, N4552);
xor XOR2 (N4706, N4691, N2702);
nand NAND4 (N4707, N4646, N3394, N1799, N4345);
nor NOR3 (N4708, N4700, N2206, N2775);
not NOT1 (N4709, N4702);
nor NOR2 (N4710, N4703, N1850);
buf BUF1 (N4711, N4709);
not NOT1 (N4712, N4705);
nor NOR2 (N4713, N4707, N4187);
xor XOR2 (N4714, N4712, N4199);
and AND2 (N4715, N4699, N2323);
buf BUF1 (N4716, N4671);
and AND4 (N4717, N4696, N3589, N3098, N2005);
xor XOR2 (N4718, N4717, N3223);
and AND4 (N4719, N4711, N3047, N1014, N1813);
xor XOR2 (N4720, N4708, N4574);
or OR3 (N4721, N4720, N3204, N3839);
or OR3 (N4722, N4718, N2607, N4373);
buf BUF1 (N4723, N4719);
or OR4 (N4724, N4706, N4113, N1331, N2427);
buf BUF1 (N4725, N4716);
not NOT1 (N4726, N4724);
xor XOR2 (N4727, N4725, N2618);
buf BUF1 (N4728, N4722);
xor XOR2 (N4729, N4727, N2423);
xor XOR2 (N4730, N4710, N2408);
and AND4 (N4731, N4714, N2444, N1195, N3783);
nand NAND2 (N4732, N4723, N4563);
or OR2 (N4733, N4693, N799);
not NOT1 (N4734, N4726);
buf BUF1 (N4735, N4715);
xor XOR2 (N4736, N4733, N3376);
nand NAND3 (N4737, N4734, N4022, N1335);
or OR3 (N4738, N4728, N3821, N3264);
xor XOR2 (N4739, N4738, N2471);
nand NAND3 (N4740, N4713, N159, N2638);
nand NAND4 (N4741, N4735, N1416, N1093, N1642);
buf BUF1 (N4742, N4737);
not NOT1 (N4743, N4731);
xor XOR2 (N4744, N4742, N3830);
xor XOR2 (N4745, N4730, N1455);
or OR2 (N4746, N4729, N2788);
not NOT1 (N4747, N4740);
buf BUF1 (N4748, N4741);
and AND4 (N4749, N4721, N4418, N4110, N716);
xor XOR2 (N4750, N4748, N4215);
xor XOR2 (N4751, N4750, N3248);
not NOT1 (N4752, N4749);
nor NOR4 (N4753, N4751, N1395, N839, N1975);
nand NAND3 (N4754, N4752, N1544, N2669);
nor NOR2 (N4755, N4754, N3460);
buf BUF1 (N4756, N4736);
not NOT1 (N4757, N4739);
and AND2 (N4758, N4755, N1602);
or OR4 (N4759, N4732, N4249, N3695, N1468);
or OR3 (N4760, N4743, N4396, N3538);
or OR3 (N4761, N4745, N1007, N1421);
xor XOR2 (N4762, N4747, N1879);
nor NOR4 (N4763, N4744, N4311, N608, N3659);
and AND4 (N4764, N4759, N2767, N2797, N2146);
nand NAND3 (N4765, N4763, N3508, N2400);
buf BUF1 (N4766, N4753);
nor NOR3 (N4767, N4765, N49, N2910);
nand NAND2 (N4768, N4758, N2684);
nand NAND2 (N4769, N4768, N3818);
nor NOR4 (N4770, N4761, N4520, N1731, N3514);
xor XOR2 (N4771, N4760, N2067);
not NOT1 (N4772, N4769);
nor NOR3 (N4773, N4756, N4522, N1653);
nor NOR2 (N4774, N4764, N4424);
nand NAND4 (N4775, N4746, N3203, N4493, N3585);
nand NAND2 (N4776, N4766, N883);
not NOT1 (N4777, N4776);
not NOT1 (N4778, N4775);
or OR3 (N4779, N4762, N1021, N4253);
nor NOR2 (N4780, N4778, N747);
nor NOR4 (N4781, N4773, N3474, N380, N4065);
xor XOR2 (N4782, N4767, N547);
and AND2 (N4783, N4772, N3096);
or OR4 (N4784, N4781, N3053, N3892, N3996);
buf BUF1 (N4785, N4770);
not NOT1 (N4786, N4771);
not NOT1 (N4787, N4783);
not NOT1 (N4788, N4757);
nand NAND2 (N4789, N4788, N2909);
nand NAND3 (N4790, N4787, N2121, N3872);
xor XOR2 (N4791, N4779, N3731);
and AND4 (N4792, N4774, N2724, N2561, N4617);
xor XOR2 (N4793, N4789, N3537);
not NOT1 (N4794, N4793);
nand NAND2 (N4795, N4790, N3508);
xor XOR2 (N4796, N4786, N1141);
xor XOR2 (N4797, N4785, N4184);
xor XOR2 (N4798, N4777, N4556);
or OR2 (N4799, N4784, N1569);
or OR2 (N4800, N4780, N1771);
not NOT1 (N4801, N4791);
or OR4 (N4802, N4782, N70, N2947, N2930);
or OR3 (N4803, N4802, N2836, N4545);
nand NAND2 (N4804, N4797, N2060);
nand NAND4 (N4805, N4798, N3544, N1139, N1706);
nor NOR2 (N4806, N4800, N3379);
nor NOR4 (N4807, N4803, N4043, N2066, N2604);
xor XOR2 (N4808, N4796, N3178);
and AND3 (N4809, N4795, N3735, N3822);
or OR4 (N4810, N4809, N3452, N638, N4396);
buf BUF1 (N4811, N4807);
or OR3 (N4812, N4808, N2411, N158);
not NOT1 (N4813, N4804);
xor XOR2 (N4814, N4811, N1391);
not NOT1 (N4815, N4801);
not NOT1 (N4816, N4799);
xor XOR2 (N4817, N4814, N645);
nand NAND2 (N4818, N4812, N1749);
nand NAND3 (N4819, N4792, N849, N4656);
buf BUF1 (N4820, N4819);
xor XOR2 (N4821, N4820, N1973);
or OR4 (N4822, N4813, N3983, N774, N4637);
xor XOR2 (N4823, N4817, N4499);
xor XOR2 (N4824, N4805, N376);
nor NOR4 (N4825, N4815, N2224, N4364, N736);
and AND4 (N4826, N4823, N3419, N1547, N4034);
or OR3 (N4827, N4810, N121, N1879);
not NOT1 (N4828, N4824);
nand NAND2 (N4829, N4794, N431);
xor XOR2 (N4830, N4829, N2674);
buf BUF1 (N4831, N4825);
buf BUF1 (N4832, N4826);
buf BUF1 (N4833, N4830);
nand NAND3 (N4834, N4831, N1622, N291);
and AND2 (N4835, N4834, N22);
nand NAND2 (N4836, N4818, N3552);
and AND2 (N4837, N4806, N521);
or OR3 (N4838, N4837, N3929, N2542);
xor XOR2 (N4839, N4838, N3365);
or OR4 (N4840, N4822, N1909, N1552, N2835);
or OR3 (N4841, N4821, N4297, N99);
nor NOR4 (N4842, N4839, N3940, N3900, N4085);
buf BUF1 (N4843, N4836);
nor NOR3 (N4844, N4843, N1485, N336);
not NOT1 (N4845, N4840);
or OR4 (N4846, N4845, N2372, N889, N92);
nand NAND4 (N4847, N4832, N3779, N1480, N1300);
or OR2 (N4848, N4827, N3584);
and AND4 (N4849, N4846, N2517, N2612, N2221);
and AND3 (N4850, N4842, N1152, N1290);
and AND4 (N4851, N4850, N3734, N3530, N3284);
or OR3 (N4852, N4848, N943, N3274);
or OR2 (N4853, N4849, N2063);
xor XOR2 (N4854, N4835, N2841);
or OR4 (N4855, N4853, N3562, N2641, N378);
nand NAND2 (N4856, N4855, N112);
not NOT1 (N4857, N4854);
or OR4 (N4858, N4856, N4281, N4178, N4332);
and AND4 (N4859, N4841, N927, N4451, N3844);
nand NAND3 (N4860, N4833, N3316, N197);
buf BUF1 (N4861, N4847);
or OR3 (N4862, N4860, N1025, N947);
xor XOR2 (N4863, N4852, N1310);
not NOT1 (N4864, N4844);
and AND4 (N4865, N4862, N1263, N1419, N4691);
nor NOR3 (N4866, N4859, N3336, N2516);
buf BUF1 (N4867, N4866);
not NOT1 (N4868, N4863);
nor NOR4 (N4869, N4865, N3603, N3294, N1541);
xor XOR2 (N4870, N4868, N4771);
nor NOR2 (N4871, N4864, N1205);
and AND2 (N4872, N4867, N1499);
or OR3 (N4873, N4816, N4079, N258);
not NOT1 (N4874, N4872);
and AND4 (N4875, N4858, N1407, N3253, N1435);
or OR4 (N4876, N4871, N2507, N972, N1182);
and AND3 (N4877, N4874, N175, N3210);
and AND3 (N4878, N4876, N1913, N402);
and AND3 (N4879, N4869, N2783, N2592);
nand NAND3 (N4880, N4878, N1499, N3646);
buf BUF1 (N4881, N4828);
or OR2 (N4882, N4873, N4363);
not NOT1 (N4883, N4861);
xor XOR2 (N4884, N4870, N3284);
and AND4 (N4885, N4877, N2225, N2643, N3246);
buf BUF1 (N4886, N4851);
buf BUF1 (N4887, N4880);
xor XOR2 (N4888, N4882, N3885);
nand NAND2 (N4889, N4881, N3635);
and AND4 (N4890, N4885, N856, N1609, N3931);
or OR3 (N4891, N4875, N1136, N3284);
buf BUF1 (N4892, N4890);
buf BUF1 (N4893, N4889);
nor NOR2 (N4894, N4892, N4811);
or OR3 (N4895, N4883, N1116, N3665);
nor NOR4 (N4896, N4887, N983, N3427, N2487);
xor XOR2 (N4897, N4886, N3978);
and AND3 (N4898, N4896, N247, N1411);
nand NAND4 (N4899, N4893, N4377, N364, N4600);
not NOT1 (N4900, N4897);
not NOT1 (N4901, N4899);
xor XOR2 (N4902, N4857, N3857);
not NOT1 (N4903, N4891);
or OR3 (N4904, N4901, N2253, N2960);
not NOT1 (N4905, N4879);
nor NOR2 (N4906, N4895, N2278);
and AND4 (N4907, N4906, N3455, N1224, N287);
xor XOR2 (N4908, N4900, N2753);
buf BUF1 (N4909, N4898);
nand NAND4 (N4910, N4894, N4345, N2568, N2784);
nand NAND2 (N4911, N4908, N4868);
buf BUF1 (N4912, N4911);
nor NOR4 (N4913, N4884, N565, N4308, N879);
nand NAND2 (N4914, N4913, N608);
not NOT1 (N4915, N4903);
nor NOR2 (N4916, N4888, N662);
or OR3 (N4917, N4907, N4503, N927);
not NOT1 (N4918, N4910);
or OR4 (N4919, N4918, N2281, N4142, N3650);
xor XOR2 (N4920, N4905, N3695);
nand NAND2 (N4921, N4919, N4404);
nor NOR4 (N4922, N4909, N3014, N2320, N1176);
or OR4 (N4923, N4912, N2224, N2550, N2556);
xor XOR2 (N4924, N4916, N4448);
nor NOR2 (N4925, N4922, N724);
xor XOR2 (N4926, N4924, N2099);
xor XOR2 (N4927, N4902, N1561);
or OR4 (N4928, N4915, N4826, N4182, N4922);
nand NAND4 (N4929, N4926, N534, N4011, N976);
and AND3 (N4930, N4928, N157, N4059);
or OR2 (N4931, N4917, N4524);
buf BUF1 (N4932, N4923);
not NOT1 (N4933, N4927);
nand NAND4 (N4934, N4904, N4617, N845, N370);
xor XOR2 (N4935, N4930, N4190);
nor NOR2 (N4936, N4929, N1943);
or OR3 (N4937, N4934, N3009, N1557);
not NOT1 (N4938, N4920);
or OR3 (N4939, N4914, N3032, N384);
or OR3 (N4940, N4921, N286, N4637);
or OR2 (N4941, N4939, N4513);
buf BUF1 (N4942, N4940);
nand NAND3 (N4943, N4931, N1322, N443);
xor XOR2 (N4944, N4935, N1766);
nand NAND2 (N4945, N4933, N2581);
and AND4 (N4946, N4938, N3217, N4222, N4697);
nor NOR3 (N4947, N4943, N1922, N2392);
nand NAND3 (N4948, N4925, N1392, N3844);
not NOT1 (N4949, N4941);
or OR2 (N4950, N4936, N1622);
xor XOR2 (N4951, N4942, N172);
and AND4 (N4952, N4951, N3728, N2155, N4360);
or OR4 (N4953, N4944, N705, N1246, N2883);
nand NAND4 (N4954, N4952, N1308, N4778, N4607);
buf BUF1 (N4955, N4950);
nor NOR4 (N4956, N4946, N1267, N866, N2948);
xor XOR2 (N4957, N4945, N3625);
xor XOR2 (N4958, N4956, N4675);
nor NOR4 (N4959, N4948, N4620, N1289, N3234);
nor NOR4 (N4960, N4949, N4718, N4596, N2733);
xor XOR2 (N4961, N4960, N3468);
nor NOR2 (N4962, N4959, N4333);
or OR4 (N4963, N4954, N1143, N3449, N4554);
and AND4 (N4964, N4958, N627, N1999, N2605);
xor XOR2 (N4965, N4932, N959);
nor NOR3 (N4966, N4961, N1566, N1197);
or OR4 (N4967, N4955, N2424, N4758, N3519);
nor NOR4 (N4968, N4962, N4117, N1134, N3745);
not NOT1 (N4969, N4968);
or OR2 (N4970, N4965, N2088);
or OR2 (N4971, N4969, N2722);
and AND2 (N4972, N4966, N901);
nor NOR3 (N4973, N4967, N3182, N468);
xor XOR2 (N4974, N4973, N2273);
buf BUF1 (N4975, N4937);
xor XOR2 (N4976, N4974, N3007);
nand NAND2 (N4977, N4953, N972);
or OR2 (N4978, N4964, N3124);
or OR3 (N4979, N4970, N2087, N754);
nor NOR4 (N4980, N4975, N4962, N2846, N3398);
not NOT1 (N4981, N4957);
nor NOR4 (N4982, N4977, N2773, N3913, N380);
and AND3 (N4983, N4982, N1285, N1669);
not NOT1 (N4984, N4978);
nor NOR3 (N4985, N4979, N4914, N4893);
and AND2 (N4986, N4963, N4543);
not NOT1 (N4987, N4985);
and AND4 (N4988, N4971, N4753, N4795, N655);
and AND4 (N4989, N4983, N4570, N4645, N1545);
not NOT1 (N4990, N4947);
nand NAND4 (N4991, N4981, N4793, N3366, N2724);
buf BUF1 (N4992, N4976);
not NOT1 (N4993, N4984);
or OR2 (N4994, N4989, N383);
and AND4 (N4995, N4980, N777, N78, N3144);
nand NAND3 (N4996, N4987, N431, N735);
or OR4 (N4997, N4972, N375, N4977, N1244);
and AND3 (N4998, N4986, N1166, N776);
and AND2 (N4999, N4990, N1963);
nor NOR4 (N5000, N4993, N2885, N2207, N2285);
not NOT1 (N5001, N4997);
nand NAND3 (N5002, N4988, N4451, N3172);
and AND2 (N5003, N4996, N4815);
nor NOR2 (N5004, N4994, N2128);
xor XOR2 (N5005, N5000, N2421);
and AND3 (N5006, N4999, N4979, N3444);
xor XOR2 (N5007, N5002, N2539);
or OR3 (N5008, N4992, N3530, N1691);
not NOT1 (N5009, N5004);
nand NAND2 (N5010, N5001, N2780);
and AND4 (N5011, N4991, N622, N806, N1047);
or OR4 (N5012, N5006, N3664, N3860, N4587);
not NOT1 (N5013, N5003);
nand NAND4 (N5014, N5008, N387, N1679, N3329);
buf BUF1 (N5015, N5005);
and AND3 (N5016, N5011, N808, N1788);
not NOT1 (N5017, N5010);
not NOT1 (N5018, N5016);
buf BUF1 (N5019, N5013);
or OR2 (N5020, N5009, N3024);
nand NAND3 (N5021, N5014, N3870, N4153);
xor XOR2 (N5022, N4998, N1135);
and AND2 (N5023, N5018, N4254);
nor NOR2 (N5024, N5015, N3042);
nor NOR3 (N5025, N5021, N1657, N4154);
nor NOR3 (N5026, N5019, N2566, N1070);
nor NOR3 (N5027, N5022, N5014, N473);
or OR3 (N5028, N5023, N2683, N3849);
nand NAND4 (N5029, N5028, N1849, N454, N3515);
xor XOR2 (N5030, N5012, N4224);
or OR3 (N5031, N5029, N1686, N913);
not NOT1 (N5032, N5020);
and AND3 (N5033, N4995, N1234, N1049);
nand NAND3 (N5034, N5030, N339, N2764);
buf BUF1 (N5035, N5017);
or OR2 (N5036, N5031, N3537);
not NOT1 (N5037, N5032);
not NOT1 (N5038, N5036);
buf BUF1 (N5039, N5026);
nand NAND2 (N5040, N5037, N346);
not NOT1 (N5041, N5038);
buf BUF1 (N5042, N5041);
buf BUF1 (N5043, N5039);
not NOT1 (N5044, N5027);
nand NAND3 (N5045, N5025, N1022, N2695);
or OR4 (N5046, N5035, N4908, N4928, N4263);
nand NAND3 (N5047, N5007, N355, N4334);
xor XOR2 (N5048, N5033, N1467);
xor XOR2 (N5049, N5045, N3445);
not NOT1 (N5050, N5042);
xor XOR2 (N5051, N5048, N4141);
buf BUF1 (N5052, N5051);
or OR3 (N5053, N5050, N364, N2955);
and AND2 (N5054, N5024, N4598);
and AND3 (N5055, N5046, N4822, N2087);
xor XOR2 (N5056, N5054, N1052);
xor XOR2 (N5057, N5049, N4089);
nor NOR3 (N5058, N5056, N1540, N3617);
and AND2 (N5059, N5052, N1814);
xor XOR2 (N5060, N5059, N2628);
buf BUF1 (N5061, N5058);
nand NAND4 (N5062, N5053, N3071, N4050, N3403);
nor NOR3 (N5063, N5044, N3580, N5);
buf BUF1 (N5064, N5055);
not NOT1 (N5065, N5062);
not NOT1 (N5066, N5064);
nor NOR2 (N5067, N5043, N2473);
buf BUF1 (N5068, N5065);
or OR4 (N5069, N5047, N1864, N1725, N61);
and AND4 (N5070, N5068, N1561, N3129, N4640);
xor XOR2 (N5071, N5069, N3890);
nor NOR3 (N5072, N5070, N4518, N4121);
nor NOR3 (N5073, N5060, N4631, N1910);
xor XOR2 (N5074, N5040, N541);
or OR2 (N5075, N5034, N3693);
nor NOR3 (N5076, N5066, N1614, N4031);
or OR4 (N5077, N5057, N5007, N889, N2394);
nand NAND4 (N5078, N5072, N4488, N4112, N4853);
xor XOR2 (N5079, N5078, N1824);
nor NOR2 (N5080, N5074, N3730);
nand NAND2 (N5081, N5076, N2622);
or OR3 (N5082, N5080, N2648, N1469);
nand NAND4 (N5083, N5081, N4332, N4898, N1066);
buf BUF1 (N5084, N5082);
buf BUF1 (N5085, N5067);
and AND4 (N5086, N5075, N696, N3960, N2670);
buf BUF1 (N5087, N5079);
not NOT1 (N5088, N5077);
and AND2 (N5089, N5083, N4951);
buf BUF1 (N5090, N5063);
and AND4 (N5091, N5088, N2224, N4089, N1625);
not NOT1 (N5092, N5089);
nor NOR2 (N5093, N5084, N3173);
xor XOR2 (N5094, N5061, N447);
buf BUF1 (N5095, N5090);
nand NAND3 (N5096, N5086, N3852, N4523);
nand NAND3 (N5097, N5093, N4828, N4233);
or OR2 (N5098, N5073, N2450);
buf BUF1 (N5099, N5085);
or OR3 (N5100, N5071, N1368, N2110);
and AND4 (N5101, N5100, N1293, N1937, N847);
buf BUF1 (N5102, N5096);
nand NAND3 (N5103, N5101, N3777, N3439);
or OR3 (N5104, N5097, N2479, N133);
nor NOR4 (N5105, N5095, N3467, N4628, N3111);
and AND4 (N5106, N5105, N1311, N2443, N3509);
buf BUF1 (N5107, N5087);
buf BUF1 (N5108, N5099);
not NOT1 (N5109, N5098);
buf BUF1 (N5110, N5103);
nand NAND2 (N5111, N5092, N493);
or OR2 (N5112, N5111, N501);
xor XOR2 (N5113, N5110, N1530);
xor XOR2 (N5114, N5104, N2487);
and AND4 (N5115, N5109, N1479, N1787, N2709);
not NOT1 (N5116, N5106);
nand NAND3 (N5117, N5102, N2706, N841);
buf BUF1 (N5118, N5115);
or OR4 (N5119, N5112, N3324, N1623, N5095);
not NOT1 (N5120, N5091);
xor XOR2 (N5121, N5120, N3577);
buf BUF1 (N5122, N5119);
and AND2 (N5123, N5108, N172);
nor NOR4 (N5124, N5123, N4528, N4537, N4706);
not NOT1 (N5125, N5107);
xor XOR2 (N5126, N5117, N507);
not NOT1 (N5127, N5126);
nor NOR4 (N5128, N5116, N2017, N3989, N1735);
buf BUF1 (N5129, N5127);
buf BUF1 (N5130, N5121);
not NOT1 (N5131, N5128);
xor XOR2 (N5132, N5094, N5009);
xor XOR2 (N5133, N5130, N1625);
nor NOR4 (N5134, N5133, N2235, N2662, N1107);
buf BUF1 (N5135, N5125);
and AND3 (N5136, N5118, N5071, N734);
and AND4 (N5137, N5136, N1282, N4903, N41);
nand NAND2 (N5138, N5132, N2398);
not NOT1 (N5139, N5134);
nand NAND4 (N5140, N5114, N2375, N4864, N4191);
xor XOR2 (N5141, N5135, N1116);
and AND3 (N5142, N5141, N1965, N621);
not NOT1 (N5143, N5142);
buf BUF1 (N5144, N5138);
not NOT1 (N5145, N5144);
or OR4 (N5146, N5124, N20, N3875, N2992);
not NOT1 (N5147, N5131);
nand NAND3 (N5148, N5143, N798, N3724);
and AND4 (N5149, N5148, N1063, N4606, N1994);
or OR3 (N5150, N5129, N4507, N2434);
nand NAND4 (N5151, N5150, N3066, N2057, N1607);
nor NOR3 (N5152, N5140, N3249, N5132);
nand NAND3 (N5153, N5146, N3153, N562);
or OR4 (N5154, N5149, N1950, N3376, N3811);
or OR4 (N5155, N5113, N626, N4713, N1271);
nand NAND4 (N5156, N5139, N3077, N4691, N4683);
not NOT1 (N5157, N5154);
nor NOR3 (N5158, N5137, N797, N2297);
nand NAND4 (N5159, N5155, N3134, N3799, N5047);
xor XOR2 (N5160, N5159, N1519);
and AND3 (N5161, N5122, N1084, N686);
or OR2 (N5162, N5151, N2056);
xor XOR2 (N5163, N5158, N3401);
and AND4 (N5164, N5162, N2067, N750, N4082);
buf BUF1 (N5165, N5164);
nand NAND4 (N5166, N5165, N928, N3367, N1785);
not NOT1 (N5167, N5156);
nand NAND2 (N5168, N5153, N4445);
buf BUF1 (N5169, N5163);
buf BUF1 (N5170, N5166);
nor NOR4 (N5171, N5157, N195, N3106, N530);
xor XOR2 (N5172, N5171, N3421);
and AND2 (N5173, N5145, N492);
xor XOR2 (N5174, N5152, N4105);
not NOT1 (N5175, N5167);
or OR4 (N5176, N5175, N1887, N3666, N2849);
nor NOR4 (N5177, N5170, N5172, N1626, N1151);
and AND3 (N5178, N3019, N2203, N640);
buf BUF1 (N5179, N5160);
not NOT1 (N5180, N5179);
nor NOR4 (N5181, N5178, N621, N3805, N4003);
not NOT1 (N5182, N5176);
xor XOR2 (N5183, N5177, N4322);
and AND3 (N5184, N5180, N205, N2830);
not NOT1 (N5185, N5183);
buf BUF1 (N5186, N5182);
nor NOR2 (N5187, N5168, N4261);
nor NOR2 (N5188, N5181, N942);
and AND3 (N5189, N5186, N4626, N3093);
nor NOR4 (N5190, N5187, N3352, N4654, N4287);
or OR2 (N5191, N5185, N2856);
buf BUF1 (N5192, N5161);
or OR2 (N5193, N5147, N2626);
and AND4 (N5194, N5174, N556, N5156, N3633);
xor XOR2 (N5195, N5190, N1281);
or OR4 (N5196, N5189, N2479, N788, N909);
nor NOR3 (N5197, N5193, N1108, N178);
nor NOR4 (N5198, N5197, N3469, N4773, N1789);
xor XOR2 (N5199, N5195, N4288);
or OR3 (N5200, N5192, N507, N1497);
xor XOR2 (N5201, N5198, N4900);
buf BUF1 (N5202, N5194);
nor NOR2 (N5203, N5173, N1912);
not NOT1 (N5204, N5191);
nor NOR3 (N5205, N5184, N4023, N3567);
nor NOR3 (N5206, N5205, N984, N4563);
and AND3 (N5207, N5201, N3331, N1907);
xor XOR2 (N5208, N5207, N3294);
nand NAND4 (N5209, N5200, N1646, N4921, N3392);
and AND3 (N5210, N5202, N456, N4775);
nand NAND3 (N5211, N5199, N1439, N297);
nand NAND4 (N5212, N5188, N1028, N2391, N1764);
nand NAND4 (N5213, N5203, N5012, N1910, N5210);
buf BUF1 (N5214, N379);
or OR2 (N5215, N5206, N2548);
and AND2 (N5216, N5204, N977);
and AND4 (N5217, N5212, N1121, N1003, N3164);
not NOT1 (N5218, N5196);
buf BUF1 (N5219, N5214);
not NOT1 (N5220, N5219);
buf BUF1 (N5221, N5208);
and AND4 (N5222, N5216, N606, N3870, N1770);
not NOT1 (N5223, N5221);
nor NOR2 (N5224, N5169, N3942);
nand NAND3 (N5225, N5209, N5125, N724);
buf BUF1 (N5226, N5225);
or OR3 (N5227, N5222, N1415, N1758);
nand NAND2 (N5228, N5218, N3552);
not NOT1 (N5229, N5217);
nor NOR3 (N5230, N5226, N2911, N4730);
xor XOR2 (N5231, N5223, N1233);
xor XOR2 (N5232, N5228, N358);
nor NOR4 (N5233, N5229, N2322, N1181, N1236);
not NOT1 (N5234, N5220);
and AND4 (N5235, N5213, N4544, N1650, N341);
xor XOR2 (N5236, N5234, N4347);
nor NOR4 (N5237, N5231, N5163, N281, N5048);
or OR3 (N5238, N5232, N365, N2427);
or OR3 (N5239, N5236, N143, N2702);
xor XOR2 (N5240, N5235, N3167);
nor NOR4 (N5241, N5224, N1654, N4346, N4726);
not NOT1 (N5242, N5233);
nor NOR3 (N5243, N5227, N3833, N3946);
or OR4 (N5244, N5237, N4646, N3677, N4094);
buf BUF1 (N5245, N5211);
not NOT1 (N5246, N5244);
not NOT1 (N5247, N5241);
buf BUF1 (N5248, N5246);
and AND4 (N5249, N5215, N1323, N4459, N1174);
or OR3 (N5250, N5247, N861, N105);
nor NOR4 (N5251, N5250, N4741, N3049, N3727);
xor XOR2 (N5252, N5239, N3121);
or OR2 (N5253, N5248, N72);
nand NAND2 (N5254, N5249, N1362);
xor XOR2 (N5255, N5245, N2216);
not NOT1 (N5256, N5251);
nor NOR4 (N5257, N5252, N4978, N2816, N2136);
xor XOR2 (N5258, N5256, N5078);
or OR4 (N5259, N5258, N1333, N4029, N3142);
or OR3 (N5260, N5243, N492, N1205);
xor XOR2 (N5261, N5253, N4024);
nor NOR4 (N5262, N5257, N3944, N1664, N1603);
xor XOR2 (N5263, N5230, N2200);
nor NOR4 (N5264, N5259, N3169, N3768, N591);
nand NAND4 (N5265, N5238, N4219, N1130, N2397);
or OR4 (N5266, N5254, N4839, N746, N5199);
buf BUF1 (N5267, N5260);
nor NOR2 (N5268, N5262, N4725);
and AND3 (N5269, N5242, N3080, N4930);
nand NAND3 (N5270, N5263, N2963, N5223);
nor NOR4 (N5271, N5266, N2502, N3025, N3164);
buf BUF1 (N5272, N5240);
not NOT1 (N5273, N5255);
or OR3 (N5274, N5269, N3644, N418);
or OR2 (N5275, N5265, N1588);
nor NOR4 (N5276, N5275, N4863, N1602, N3439);
nor NOR2 (N5277, N5274, N2646);
or OR2 (N5278, N5264, N3780);
nand NAND3 (N5279, N5278, N3621, N3770);
nand NAND4 (N5280, N5261, N2744, N3372, N2717);
buf BUF1 (N5281, N5276);
not NOT1 (N5282, N5270);
nand NAND4 (N5283, N5267, N4054, N4119, N491);
nor NOR3 (N5284, N5271, N2478, N3947);
nor NOR3 (N5285, N5268, N2219, N2581);
buf BUF1 (N5286, N5285);
or OR2 (N5287, N5280, N1989);
and AND3 (N5288, N5287, N409, N1346);
or OR4 (N5289, N5283, N2822, N1698, N3567);
nand NAND3 (N5290, N5284, N4685, N2074);
not NOT1 (N5291, N5281);
buf BUF1 (N5292, N5290);
nand NAND3 (N5293, N5286, N1807, N573);
nor NOR4 (N5294, N5288, N4412, N3647, N2448);
and AND3 (N5295, N5293, N4981, N4676);
not NOT1 (N5296, N5273);
and AND3 (N5297, N5277, N3318, N1326);
nand NAND3 (N5298, N5279, N1884, N3536);
or OR4 (N5299, N5298, N2225, N4395, N420);
or OR3 (N5300, N5299, N4022, N1641);
nand NAND2 (N5301, N5282, N2895);
and AND3 (N5302, N5292, N2782, N2707);
nor NOR3 (N5303, N5300, N4841, N3987);
and AND4 (N5304, N5294, N4205, N4871, N4202);
xor XOR2 (N5305, N5302, N4125);
not NOT1 (N5306, N5304);
or OR3 (N5307, N5306, N1053, N34);
nand NAND4 (N5308, N5296, N470, N185, N577);
xor XOR2 (N5309, N5289, N1879);
nand NAND4 (N5310, N5303, N4068, N5017, N1033);
xor XOR2 (N5311, N5272, N3858);
buf BUF1 (N5312, N5311);
nor NOR2 (N5313, N5291, N476);
or OR4 (N5314, N5295, N1424, N2834, N2510);
or OR2 (N5315, N5301, N2142);
nand NAND2 (N5316, N5310, N1183);
xor XOR2 (N5317, N5308, N2521);
xor XOR2 (N5318, N5314, N5062);
buf BUF1 (N5319, N5297);
or OR3 (N5320, N5315, N3398, N1481);
not NOT1 (N5321, N5316);
nor NOR2 (N5322, N5313, N4596);
and AND4 (N5323, N5321, N2498, N315, N1402);
and AND2 (N5324, N5318, N1163);
nand NAND4 (N5325, N5320, N2107, N4907, N355);
or OR2 (N5326, N5309, N1802);
or OR2 (N5327, N5312, N1015);
buf BUF1 (N5328, N5317);
nand NAND4 (N5329, N5307, N4813, N281, N1195);
or OR2 (N5330, N5326, N383);
nor NOR2 (N5331, N5322, N3434);
and AND4 (N5332, N5319, N1369, N4145, N2203);
or OR2 (N5333, N5329, N1538);
xor XOR2 (N5334, N5332, N1700);
not NOT1 (N5335, N5305);
xor XOR2 (N5336, N5327, N4863);
or OR4 (N5337, N5331, N5075, N4891, N3630);
xor XOR2 (N5338, N5336, N5157);
nor NOR4 (N5339, N5337, N1149, N2228, N4923);
xor XOR2 (N5340, N5325, N623);
or OR4 (N5341, N5330, N2513, N2680, N35);
xor XOR2 (N5342, N5335, N1363);
buf BUF1 (N5343, N5338);
xor XOR2 (N5344, N5323, N4353);
xor XOR2 (N5345, N5328, N1724);
not NOT1 (N5346, N5340);
not NOT1 (N5347, N5324);
buf BUF1 (N5348, N5347);
buf BUF1 (N5349, N5334);
nor NOR3 (N5350, N5333, N3908, N3082);
nand NAND2 (N5351, N5341, N5208);
or OR4 (N5352, N5346, N3819, N4554, N2106);
not NOT1 (N5353, N5339);
or OR3 (N5354, N5348, N1615, N2683);
or OR4 (N5355, N5345, N2722, N5052, N3414);
xor XOR2 (N5356, N5353, N3080);
nor NOR2 (N5357, N5355, N4608);
and AND4 (N5358, N5354, N1322, N1149, N2011);
or OR3 (N5359, N5357, N4083, N718);
xor XOR2 (N5360, N5349, N616);
or OR3 (N5361, N5359, N4267, N5107);
xor XOR2 (N5362, N5351, N4662);
nor NOR4 (N5363, N5361, N596, N3200, N3469);
xor XOR2 (N5364, N5362, N616);
buf BUF1 (N5365, N5358);
xor XOR2 (N5366, N5342, N5052);
or OR2 (N5367, N5344, N1152);
nor NOR4 (N5368, N5366, N4708, N2397, N4165);
nor NOR2 (N5369, N5363, N4131);
nor NOR4 (N5370, N5360, N275, N3868, N1446);
and AND4 (N5371, N5352, N1147, N553, N3753);
and AND2 (N5372, N5368, N4594);
buf BUF1 (N5373, N5371);
nand NAND2 (N5374, N5356, N36);
or OR4 (N5375, N5350, N4280, N3235, N1100);
not NOT1 (N5376, N5374);
buf BUF1 (N5377, N5365);
and AND4 (N5378, N5367, N2038, N3447, N3971);
nor NOR3 (N5379, N5378, N1235, N357);
nand NAND4 (N5380, N5370, N3343, N196, N739);
nand NAND3 (N5381, N5364, N3337, N5082);
xor XOR2 (N5382, N5343, N3818);
buf BUF1 (N5383, N5377);
buf BUF1 (N5384, N5381);
not NOT1 (N5385, N5384);
nand NAND2 (N5386, N5369, N364);
buf BUF1 (N5387, N5380);
and AND4 (N5388, N5379, N3080, N168, N2772);
nor NOR2 (N5389, N5386, N4683);
nand NAND3 (N5390, N5389, N1640, N1669);
nand NAND3 (N5391, N5372, N2096, N5223);
nand NAND3 (N5392, N5391, N4748, N879);
nand NAND4 (N5393, N5373, N3868, N5105, N4634);
nor NOR2 (N5394, N5392, N3091);
xor XOR2 (N5395, N5393, N3108);
nand NAND4 (N5396, N5385, N3440, N4478, N3626);
nor NOR2 (N5397, N5383, N3988);
and AND4 (N5398, N5396, N4160, N566, N2917);
not NOT1 (N5399, N5397);
and AND4 (N5400, N5382, N1072, N1875, N2614);
buf BUF1 (N5401, N5375);
or OR4 (N5402, N5401, N3916, N285, N2527);
nor NOR3 (N5403, N5402, N2660, N2255);
or OR2 (N5404, N5376, N5046);
or OR2 (N5405, N5398, N4495);
and AND2 (N5406, N5404, N3198);
not NOT1 (N5407, N5403);
and AND2 (N5408, N5390, N3388);
not NOT1 (N5409, N5394);
buf BUF1 (N5410, N5405);
not NOT1 (N5411, N5409);
nor NOR3 (N5412, N5406, N5305, N2278);
buf BUF1 (N5413, N5412);
not NOT1 (N5414, N5399);
xor XOR2 (N5415, N5408, N403);
buf BUF1 (N5416, N5395);
or OR2 (N5417, N5407, N3397);
and AND3 (N5418, N5417, N2865, N536);
or OR3 (N5419, N5400, N5276, N1073);
not NOT1 (N5420, N5414);
nor NOR4 (N5421, N5416, N3190, N1216, N3694);
nor NOR3 (N5422, N5420, N2496, N5015);
or OR4 (N5423, N5411, N1905, N3102, N850);
not NOT1 (N5424, N5422);
nand NAND4 (N5425, N5424, N1671, N4387, N2330);
or OR2 (N5426, N5419, N444);
not NOT1 (N5427, N5426);
buf BUF1 (N5428, N5413);
nand NAND4 (N5429, N5387, N2996, N3560, N602);
or OR4 (N5430, N5421, N3052, N4299, N848);
not NOT1 (N5431, N5423);
nand NAND2 (N5432, N5429, N5087);
nand NAND4 (N5433, N5432, N4320, N129, N212);
or OR2 (N5434, N5427, N4366);
or OR3 (N5435, N5431, N1178, N833);
and AND4 (N5436, N5410, N4113, N1741, N2034);
or OR3 (N5437, N5415, N1610, N2836);
and AND2 (N5438, N5388, N947);
not NOT1 (N5439, N5435);
and AND2 (N5440, N5428, N3852);
nand NAND3 (N5441, N5438, N918, N2224);
buf BUF1 (N5442, N5430);
buf BUF1 (N5443, N5442);
not NOT1 (N5444, N5425);
and AND2 (N5445, N5444, N2545);
not NOT1 (N5446, N5434);
nor NOR2 (N5447, N5439, N93);
not NOT1 (N5448, N5447);
nand NAND3 (N5449, N5433, N2682, N1619);
and AND3 (N5450, N5445, N4703, N3658);
buf BUF1 (N5451, N5440);
buf BUF1 (N5452, N5446);
nor NOR2 (N5453, N5443, N44);
not NOT1 (N5454, N5437);
nor NOR3 (N5455, N5452, N1053, N5242);
or OR4 (N5456, N5455, N410, N3526, N2819);
or OR4 (N5457, N5418, N4366, N2512, N3700);
and AND4 (N5458, N5457, N3570, N5191, N4925);
nor NOR3 (N5459, N5453, N4076, N2497);
and AND3 (N5460, N5436, N1045, N2808);
or OR3 (N5461, N5460, N5042, N4957);
nor NOR3 (N5462, N5449, N4084, N1038);
xor XOR2 (N5463, N5454, N3956);
xor XOR2 (N5464, N5459, N1584);
nand NAND4 (N5465, N5458, N2717, N3271, N4407);
and AND2 (N5466, N5451, N2330);
or OR4 (N5467, N5441, N3440, N464, N580);
and AND4 (N5468, N5448, N1206, N4559, N2704);
and AND4 (N5469, N5464, N3766, N2376, N1257);
and AND4 (N5470, N5462, N3346, N5424, N2414);
xor XOR2 (N5471, N5463, N4427);
xor XOR2 (N5472, N5466, N2416);
nor NOR2 (N5473, N5465, N1185);
or OR3 (N5474, N5469, N2218, N1427);
buf BUF1 (N5475, N5468);
nand NAND2 (N5476, N5474, N5236);
nor NOR3 (N5477, N5471, N5427, N732);
and AND3 (N5478, N5467, N3418, N2758);
or OR3 (N5479, N5478, N2930, N1996);
buf BUF1 (N5480, N5450);
not NOT1 (N5481, N5473);
xor XOR2 (N5482, N5476, N1545);
xor XOR2 (N5483, N5477, N1919);
buf BUF1 (N5484, N5475);
nor NOR4 (N5485, N5470, N3568, N9, N603);
buf BUF1 (N5486, N5480);
not NOT1 (N5487, N5484);
xor XOR2 (N5488, N5482, N4652);
nor NOR2 (N5489, N5479, N92);
nand NAND2 (N5490, N5456, N1861);
xor XOR2 (N5491, N5486, N3474);
xor XOR2 (N5492, N5483, N4034);
not NOT1 (N5493, N5461);
buf BUF1 (N5494, N5487);
xor XOR2 (N5495, N5485, N5038);
and AND3 (N5496, N5489, N405, N3126);
buf BUF1 (N5497, N5493);
not NOT1 (N5498, N5494);
and AND4 (N5499, N5495, N2887, N2428, N1989);
not NOT1 (N5500, N5488);
or OR3 (N5501, N5481, N692, N1571);
nor NOR3 (N5502, N5498, N1925, N3365);
or OR2 (N5503, N5490, N4183);
and AND4 (N5504, N5502, N915, N4814, N4689);
or OR2 (N5505, N5497, N5171);
buf BUF1 (N5506, N5505);
xor XOR2 (N5507, N5499, N2846);
or OR4 (N5508, N5472, N4463, N5324, N128);
not NOT1 (N5509, N5504);
nor NOR4 (N5510, N5500, N4434, N4286, N4440);
buf BUF1 (N5511, N5492);
buf BUF1 (N5512, N5503);
nand NAND3 (N5513, N5491, N2438, N2808);
nand NAND3 (N5514, N5506, N599, N4238);
nor NOR3 (N5515, N5501, N3177, N4567);
nor NOR2 (N5516, N5513, N1842);
and AND2 (N5517, N5511, N3504);
nor NOR4 (N5518, N5496, N4826, N889, N1542);
nand NAND3 (N5519, N5508, N1585, N3684);
xor XOR2 (N5520, N5510, N5402);
not NOT1 (N5521, N5520);
and AND3 (N5522, N5514, N3015, N3546);
xor XOR2 (N5523, N5515, N507);
or OR2 (N5524, N5509, N2788);
and AND2 (N5525, N5512, N4930);
or OR3 (N5526, N5518, N4176, N2165);
nor NOR2 (N5527, N5522, N1935);
nor NOR2 (N5528, N5525, N49);
nand NAND2 (N5529, N5519, N3352);
buf BUF1 (N5530, N5526);
xor XOR2 (N5531, N5524, N3398);
and AND2 (N5532, N5523, N4830);
xor XOR2 (N5533, N5507, N2300);
and AND4 (N5534, N5528, N707, N126, N4952);
buf BUF1 (N5535, N5532);
nand NAND2 (N5536, N5533, N781);
and AND2 (N5537, N5536, N3844);
and AND3 (N5538, N5535, N2765, N4340);
buf BUF1 (N5539, N5516);
xor XOR2 (N5540, N5537, N2043);
or OR3 (N5541, N5530, N2445, N2600);
xor XOR2 (N5542, N5539, N1083);
or OR4 (N5543, N5531, N1872, N3322, N1199);
not NOT1 (N5544, N5521);
buf BUF1 (N5545, N5542);
xor XOR2 (N5546, N5541, N3505);
buf BUF1 (N5547, N5544);
buf BUF1 (N5548, N5540);
and AND2 (N5549, N5543, N1733);
xor XOR2 (N5550, N5529, N3215);
nor NOR2 (N5551, N5527, N1095);
or OR2 (N5552, N5545, N5180);
not NOT1 (N5553, N5551);
buf BUF1 (N5554, N5552);
buf BUF1 (N5555, N5538);
not NOT1 (N5556, N5549);
and AND4 (N5557, N5556, N4003, N4425, N1617);
buf BUF1 (N5558, N5557);
nor NOR4 (N5559, N5554, N1569, N3492, N60);
or OR3 (N5560, N5534, N2422, N2545);
or OR3 (N5561, N5548, N4703, N2146);
nand NAND2 (N5562, N5546, N921);
not NOT1 (N5563, N5547);
xor XOR2 (N5564, N5559, N3007);
or OR2 (N5565, N5555, N4293);
or OR2 (N5566, N5560, N5005);
and AND2 (N5567, N5565, N5543);
or OR3 (N5568, N5566, N3718, N1189);
or OR3 (N5569, N5562, N4543, N5175);
and AND3 (N5570, N5564, N1577, N38);
nand NAND4 (N5571, N5558, N4368, N4993, N3681);
not NOT1 (N5572, N5561);
xor XOR2 (N5573, N5517, N664);
not NOT1 (N5574, N5553);
nor NOR3 (N5575, N5567, N592, N4088);
buf BUF1 (N5576, N5569);
xor XOR2 (N5577, N5572, N1477);
xor XOR2 (N5578, N5576, N4227);
or OR2 (N5579, N5563, N303);
xor XOR2 (N5580, N5578, N2);
buf BUF1 (N5581, N5577);
and AND4 (N5582, N5579, N994, N4142, N221);
xor XOR2 (N5583, N5575, N2460);
xor XOR2 (N5584, N5580, N1029);
or OR3 (N5585, N5568, N1992, N4947);
not NOT1 (N5586, N5584);
nor NOR4 (N5587, N5586, N291, N3670, N3219);
not NOT1 (N5588, N5550);
xor XOR2 (N5589, N5574, N3592);
and AND4 (N5590, N5573, N1422, N1819, N3760);
xor XOR2 (N5591, N5571, N2889);
nor NOR2 (N5592, N5589, N5484);
nor NOR2 (N5593, N5591, N3265);
not NOT1 (N5594, N5585);
nand NAND2 (N5595, N5581, N5356);
and AND3 (N5596, N5593, N273, N3413);
and AND4 (N5597, N5595, N4333, N1396, N435);
not NOT1 (N5598, N5590);
nor NOR4 (N5599, N5596, N4645, N5450, N2855);
or OR4 (N5600, N5597, N4697, N2867, N2353);
nand NAND2 (N5601, N5570, N4402);
nand NAND4 (N5602, N5582, N405, N4655, N377);
and AND3 (N5603, N5600, N5520, N1346);
buf BUF1 (N5604, N5602);
and AND3 (N5605, N5599, N3211, N3052);
buf BUF1 (N5606, N5604);
buf BUF1 (N5607, N5606);
and AND3 (N5608, N5588, N3936, N3938);
and AND3 (N5609, N5607, N3435, N270);
or OR2 (N5610, N5609, N841);
nand NAND2 (N5611, N5583, N5161);
nand NAND3 (N5612, N5592, N5508, N4215);
nand NAND2 (N5613, N5610, N768);
nor NOR3 (N5614, N5587, N891, N3676);
not NOT1 (N5615, N5605);
nand NAND3 (N5616, N5613, N5217, N5449);
nor NOR3 (N5617, N5594, N4040, N1869);
xor XOR2 (N5618, N5616, N1518);
nand NAND4 (N5619, N5603, N3746, N969, N313);
and AND3 (N5620, N5601, N1150, N2210);
buf BUF1 (N5621, N5611);
and AND3 (N5622, N5608, N3081, N4912);
xor XOR2 (N5623, N5621, N1915);
xor XOR2 (N5624, N5612, N5316);
xor XOR2 (N5625, N5622, N4301);
nor NOR2 (N5626, N5614, N4601);
xor XOR2 (N5627, N5623, N404);
nor NOR3 (N5628, N5615, N3540, N3123);
or OR2 (N5629, N5626, N3000);
nand NAND3 (N5630, N5624, N3991, N3732);
nor NOR4 (N5631, N5630, N4127, N4516, N1775);
and AND4 (N5632, N5625, N4372, N3503, N3187);
nor NOR4 (N5633, N5629, N848, N5620, N220);
nand NAND3 (N5634, N1873, N3981, N1462);
and AND3 (N5635, N5633, N2175, N4032);
xor XOR2 (N5636, N5631, N2437);
and AND2 (N5637, N5619, N3212);
nand NAND2 (N5638, N5627, N2628);
nor NOR3 (N5639, N5637, N2632, N1425);
or OR4 (N5640, N5638, N4481, N5172, N444);
not NOT1 (N5641, N5635);
buf BUF1 (N5642, N5617);
xor XOR2 (N5643, N5618, N2580);
nor NOR3 (N5644, N5636, N911, N4399);
or OR2 (N5645, N5644, N3871);
and AND3 (N5646, N5632, N2013, N1263);
or OR3 (N5647, N5640, N1155, N854);
not NOT1 (N5648, N5639);
nand NAND2 (N5649, N5648, N1617);
nand NAND4 (N5650, N5641, N3699, N5300, N1034);
not NOT1 (N5651, N5634);
nand NAND3 (N5652, N5651, N1365, N2133);
not NOT1 (N5653, N5647);
or OR4 (N5654, N5652, N4630, N1249, N3613);
nor NOR3 (N5655, N5653, N3385, N2937);
nor NOR4 (N5656, N5655, N1769, N1910, N517);
or OR4 (N5657, N5645, N4124, N5598, N706);
and AND2 (N5658, N5470, N1691);
nor NOR3 (N5659, N5643, N3041, N2482);
or OR3 (N5660, N5658, N2918, N2672);
and AND4 (N5661, N5642, N462, N2175, N701);
buf BUF1 (N5662, N5659);
buf BUF1 (N5663, N5661);
and AND2 (N5664, N5650, N900);
nand NAND4 (N5665, N5657, N2776, N2481, N4077);
xor XOR2 (N5666, N5649, N120);
xor XOR2 (N5667, N5656, N2768);
or OR4 (N5668, N5628, N1389, N2637, N941);
nor NOR2 (N5669, N5665, N1784);
not NOT1 (N5670, N5663);
nor NOR3 (N5671, N5646, N762, N538);
buf BUF1 (N5672, N5669);
not NOT1 (N5673, N5668);
not NOT1 (N5674, N5662);
not NOT1 (N5675, N5660);
buf BUF1 (N5676, N5671);
nor NOR2 (N5677, N5675, N551);
and AND2 (N5678, N5676, N4595);
nand NAND3 (N5679, N5672, N2572, N2505);
nor NOR3 (N5680, N5673, N207, N856);
and AND3 (N5681, N5666, N5307, N5343);
buf BUF1 (N5682, N5678);
or OR3 (N5683, N5670, N4503, N3901);
buf BUF1 (N5684, N5667);
nand NAND3 (N5685, N5677, N2598, N5272);
or OR3 (N5686, N5680, N2246, N2613);
buf BUF1 (N5687, N5674);
nand NAND3 (N5688, N5687, N2732, N5343);
and AND4 (N5689, N5681, N3607, N5677, N3376);
not NOT1 (N5690, N5684);
xor XOR2 (N5691, N5689, N466);
xor XOR2 (N5692, N5654, N4973);
nand NAND2 (N5693, N5692, N5129);
nand NAND4 (N5694, N5679, N2154, N593, N5614);
nor NOR2 (N5695, N5694, N2215);
nor NOR2 (N5696, N5693, N4203);
nor NOR3 (N5697, N5683, N1399, N4623);
nand NAND2 (N5698, N5686, N5593);
xor XOR2 (N5699, N5685, N4111);
nand NAND3 (N5700, N5688, N567, N3845);
or OR2 (N5701, N5699, N3712);
and AND2 (N5702, N5696, N3852);
xor XOR2 (N5703, N5691, N72);
nor NOR2 (N5704, N5702, N4604);
nand NAND2 (N5705, N5697, N3696);
buf BUF1 (N5706, N5682);
nor NOR3 (N5707, N5706, N801, N4458);
not NOT1 (N5708, N5703);
nand NAND2 (N5709, N5707, N2990);
not NOT1 (N5710, N5695);
not NOT1 (N5711, N5709);
not NOT1 (N5712, N5700);
nor NOR2 (N5713, N5711, N718);
not NOT1 (N5714, N5664);
or OR3 (N5715, N5690, N1173, N1464);
or OR3 (N5716, N5714, N2511, N1897);
nand NAND4 (N5717, N5712, N4127, N5418, N331);
nand NAND4 (N5718, N5698, N3197, N80, N5550);
and AND2 (N5719, N5710, N4784);
not NOT1 (N5720, N5717);
xor XOR2 (N5721, N5705, N4746);
nor NOR3 (N5722, N5721, N5284, N5407);
nand NAND2 (N5723, N5718, N611);
or OR3 (N5724, N5719, N5125, N2181);
or OR2 (N5725, N5723, N1634);
not NOT1 (N5726, N5722);
and AND3 (N5727, N5725, N2493, N24);
or OR3 (N5728, N5726, N5072, N4952);
xor XOR2 (N5729, N5728, N4407);
or OR4 (N5730, N5729, N3582, N2806, N1562);
and AND4 (N5731, N5708, N3258, N5075, N1553);
nor NOR2 (N5732, N5715, N1874);
xor XOR2 (N5733, N5727, N577);
nor NOR4 (N5734, N5724, N3005, N1377, N4749);
xor XOR2 (N5735, N5713, N3768);
and AND4 (N5736, N5701, N5371, N407, N5301);
nor NOR4 (N5737, N5716, N272, N5477, N1988);
and AND2 (N5738, N5736, N2614);
nand NAND2 (N5739, N5737, N1879);
and AND2 (N5740, N5732, N3954);
and AND3 (N5741, N5731, N17, N4957);
nor NOR4 (N5742, N5733, N5274, N1869, N3497);
and AND2 (N5743, N5740, N3146);
xor XOR2 (N5744, N5720, N5700);
xor XOR2 (N5745, N5739, N90);
not NOT1 (N5746, N5741);
not NOT1 (N5747, N5704);
xor XOR2 (N5748, N5745, N4596);
nor NOR2 (N5749, N5735, N1733);
nand NAND4 (N5750, N5747, N1960, N4743, N535);
nor NOR2 (N5751, N5734, N2795);
or OR2 (N5752, N5750, N4851);
nor NOR2 (N5753, N5751, N789);
nand NAND4 (N5754, N5749, N328, N5678, N3582);
xor XOR2 (N5755, N5748, N5750);
xor XOR2 (N5756, N5746, N5524);
or OR2 (N5757, N5756, N1462);
nor NOR4 (N5758, N5752, N1861, N743, N3975);
buf BUF1 (N5759, N5744);
and AND2 (N5760, N5755, N2193);
nor NOR2 (N5761, N5738, N2531);
nand NAND2 (N5762, N5754, N5500);
nand NAND2 (N5763, N5758, N2756);
xor XOR2 (N5764, N5762, N2988);
and AND3 (N5765, N5761, N3246, N4954);
or OR4 (N5766, N5764, N1621, N3293, N1941);
and AND4 (N5767, N5743, N5711, N4497, N5447);
xor XOR2 (N5768, N5742, N3494);
buf BUF1 (N5769, N5753);
or OR2 (N5770, N5757, N4089);
nor NOR4 (N5771, N5766, N4154, N2513, N4397);
and AND2 (N5772, N5759, N3127);
or OR4 (N5773, N5769, N615, N675, N5603);
not NOT1 (N5774, N5760);
nor NOR4 (N5775, N5763, N324, N2244, N2065);
nand NAND4 (N5776, N5730, N5430, N5397, N1624);
and AND4 (N5777, N5776, N971, N1242, N1193);
nand NAND3 (N5778, N5770, N1299, N3333);
nand NAND2 (N5779, N5778, N4509);
buf BUF1 (N5780, N5765);
not NOT1 (N5781, N5779);
xor XOR2 (N5782, N5767, N183);
xor XOR2 (N5783, N5777, N1235);
nand NAND3 (N5784, N5774, N3220, N346);
nor NOR3 (N5785, N5771, N2780, N5159);
xor XOR2 (N5786, N5773, N2598);
xor XOR2 (N5787, N5783, N5343);
not NOT1 (N5788, N5780);
buf BUF1 (N5789, N5782);
and AND3 (N5790, N5785, N279, N192);
xor XOR2 (N5791, N5786, N758);
xor XOR2 (N5792, N5772, N2351);
nand NAND2 (N5793, N5775, N5685);
xor XOR2 (N5794, N5793, N599);
buf BUF1 (N5795, N5794);
and AND3 (N5796, N5790, N3786, N4575);
buf BUF1 (N5797, N5784);
buf BUF1 (N5798, N5796);
buf BUF1 (N5799, N5798);
and AND2 (N5800, N5799, N3607);
or OR4 (N5801, N5795, N4599, N5727, N4442);
xor XOR2 (N5802, N5791, N617);
nor NOR3 (N5803, N5797, N3344, N3485);
not NOT1 (N5804, N5788);
nor NOR2 (N5805, N5781, N5026);
or OR2 (N5806, N5800, N2017);
not NOT1 (N5807, N5768);
buf BUF1 (N5808, N5803);
xor XOR2 (N5809, N5808, N2880);
not NOT1 (N5810, N5792);
buf BUF1 (N5811, N5789);
nor NOR2 (N5812, N5802, N4455);
xor XOR2 (N5813, N5787, N1022);
xor XOR2 (N5814, N5804, N261);
or OR2 (N5815, N5812, N4999);
or OR3 (N5816, N5809, N5388, N3048);
nor NOR4 (N5817, N5807, N4536, N3768, N731);
and AND3 (N5818, N5813, N2857, N4416);
and AND3 (N5819, N5817, N4744, N5035);
nand NAND3 (N5820, N5810, N2037, N3001);
nor NOR2 (N5821, N5811, N2560);
or OR4 (N5822, N5820, N3307, N3356, N4713);
buf BUF1 (N5823, N5816);
nand NAND3 (N5824, N5806, N4528, N626);
nand NAND3 (N5825, N5815, N1572, N1139);
nor NOR3 (N5826, N5821, N5363, N3157);
nand NAND3 (N5827, N5801, N200, N3862);
nor NOR4 (N5828, N5825, N756, N3490, N3670);
and AND2 (N5829, N5823, N3800);
or OR4 (N5830, N5824, N1087, N5129, N115);
xor XOR2 (N5831, N5826, N1656);
buf BUF1 (N5832, N5805);
buf BUF1 (N5833, N5830);
not NOT1 (N5834, N5833);
or OR4 (N5835, N5829, N5375, N1035, N2624);
nor NOR2 (N5836, N5834, N3315);
and AND3 (N5837, N5828, N4910, N2545);
nor NOR2 (N5838, N5822, N5032);
and AND3 (N5839, N5838, N5117, N4624);
buf BUF1 (N5840, N5839);
and AND3 (N5841, N5819, N1726, N1369);
or OR2 (N5842, N5840, N601);
xor XOR2 (N5843, N5837, N2816);
xor XOR2 (N5844, N5842, N3752);
nor NOR4 (N5845, N5814, N4581, N5137, N3299);
or OR2 (N5846, N5835, N1691);
xor XOR2 (N5847, N5844, N4748);
xor XOR2 (N5848, N5818, N2996);
not NOT1 (N5849, N5847);
not NOT1 (N5850, N5831);
nor NOR3 (N5851, N5841, N1981, N4125);
nor NOR2 (N5852, N5836, N2000);
and AND3 (N5853, N5827, N3947, N1402);
and AND4 (N5854, N5850, N1334, N5406, N5131);
xor XOR2 (N5855, N5845, N1852);
or OR2 (N5856, N5854, N5229);
nand NAND2 (N5857, N5853, N621);
and AND3 (N5858, N5851, N3708, N2939);
or OR3 (N5859, N5858, N5235, N5468);
nand NAND2 (N5860, N5859, N4319);
nand NAND2 (N5861, N5860, N1693);
or OR3 (N5862, N5852, N3098, N3531);
xor XOR2 (N5863, N5849, N4911);
buf BUF1 (N5864, N5861);
nand NAND3 (N5865, N5848, N2916, N3952);
nand NAND4 (N5866, N5865, N5181, N194, N2738);
buf BUF1 (N5867, N5855);
and AND4 (N5868, N5857, N3213, N2789, N4145);
nor NOR4 (N5869, N5864, N1712, N615, N4786);
buf BUF1 (N5870, N5866);
nor NOR2 (N5871, N5846, N4773);
not NOT1 (N5872, N5868);
nor NOR3 (N5873, N5870, N5090, N3283);
xor XOR2 (N5874, N5856, N1612);
not NOT1 (N5875, N5871);
nor NOR2 (N5876, N5867, N5325);
nor NOR3 (N5877, N5873, N3294, N2366);
xor XOR2 (N5878, N5876, N3883);
or OR3 (N5879, N5832, N4039, N5578);
or OR4 (N5880, N5843, N2863, N5414, N5648);
nand NAND2 (N5881, N5863, N3307);
or OR2 (N5882, N5880, N2061);
buf BUF1 (N5883, N5869);
or OR3 (N5884, N5878, N3204, N3670);
buf BUF1 (N5885, N5875);
and AND2 (N5886, N5884, N2890);
and AND2 (N5887, N5882, N3025);
not NOT1 (N5888, N5877);
not NOT1 (N5889, N5883);
and AND2 (N5890, N5887, N1145);
and AND2 (N5891, N5888, N2947);
xor XOR2 (N5892, N5879, N2670);
nand NAND3 (N5893, N5881, N2041, N1501);
or OR3 (N5894, N5889, N3991, N5704);
and AND3 (N5895, N5892, N4623, N5334);
nand NAND2 (N5896, N5886, N4289);
xor XOR2 (N5897, N5885, N1764);
nand NAND4 (N5898, N5894, N4602, N4833, N5115);
xor XOR2 (N5899, N5874, N4841);
nand NAND2 (N5900, N5896, N2087);
buf BUF1 (N5901, N5900);
or OR2 (N5902, N5893, N3519);
or OR4 (N5903, N5901, N1866, N3704, N5091);
xor XOR2 (N5904, N5902, N386);
nand NAND4 (N5905, N5899, N1252, N2489, N2858);
buf BUF1 (N5906, N5862);
nor NOR4 (N5907, N5895, N5464, N4312, N763);
and AND2 (N5908, N5907, N3960);
xor XOR2 (N5909, N5906, N2538);
nor NOR4 (N5910, N5897, N4627, N3700, N2994);
or OR4 (N5911, N5898, N4616, N2070, N2005);
buf BUF1 (N5912, N5872);
nor NOR2 (N5913, N5910, N4906);
nor NOR3 (N5914, N5890, N782, N3353);
xor XOR2 (N5915, N5903, N433);
and AND3 (N5916, N5914, N4233, N3711);
buf BUF1 (N5917, N5891);
buf BUF1 (N5918, N5908);
buf BUF1 (N5919, N5917);
buf BUF1 (N5920, N5905);
xor XOR2 (N5921, N5915, N1075);
and AND3 (N5922, N5918, N2275, N5870);
nand NAND3 (N5923, N5919, N4031, N3834);
nor NOR4 (N5924, N5904, N3742, N92, N5177);
not NOT1 (N5925, N5909);
xor XOR2 (N5926, N5913, N2411);
and AND4 (N5927, N5920, N3367, N2164, N5585);
buf BUF1 (N5928, N5921);
buf BUF1 (N5929, N5922);
and AND4 (N5930, N5929, N1771, N4761, N12);
buf BUF1 (N5931, N5927);
buf BUF1 (N5932, N5912);
nor NOR2 (N5933, N5932, N4526);
not NOT1 (N5934, N5911);
and AND3 (N5935, N5928, N4164, N5121);
buf BUF1 (N5936, N5924);
nand NAND3 (N5937, N5933, N3050, N3379);
or OR4 (N5938, N5935, N1340, N3939, N5125);
buf BUF1 (N5939, N5938);
not NOT1 (N5940, N5934);
or OR2 (N5941, N5939, N3718);
buf BUF1 (N5942, N5916);
xor XOR2 (N5943, N5925, N5636);
xor XOR2 (N5944, N5923, N4720);
nor NOR3 (N5945, N5931, N5668, N4468);
and AND3 (N5946, N5937, N2079, N2279);
buf BUF1 (N5947, N5940);
or OR3 (N5948, N5945, N527, N185);
buf BUF1 (N5949, N5926);
and AND4 (N5950, N5949, N2743, N5131, N4);
and AND2 (N5951, N5936, N5609);
nand NAND2 (N5952, N5930, N5231);
not NOT1 (N5953, N5947);
or OR2 (N5954, N5951, N1412);
buf BUF1 (N5955, N5954);
nand NAND3 (N5956, N5942, N2193, N2775);
buf BUF1 (N5957, N5943);
or OR3 (N5958, N5950, N3603, N4279);
and AND2 (N5959, N5941, N504);
buf BUF1 (N5960, N5959);
or OR2 (N5961, N5955, N4009);
or OR3 (N5962, N5952, N5379, N4073);
not NOT1 (N5963, N5961);
or OR2 (N5964, N5960, N1127);
buf BUF1 (N5965, N5958);
nor NOR3 (N5966, N5953, N4767, N323);
xor XOR2 (N5967, N5964, N2327);
nor NOR3 (N5968, N5946, N3640, N606);
buf BUF1 (N5969, N5963);
or OR2 (N5970, N5969, N5793);
nor NOR3 (N5971, N5965, N209, N5319);
and AND2 (N5972, N5957, N727);
nand NAND3 (N5973, N5962, N3039, N3071);
buf BUF1 (N5974, N5967);
and AND3 (N5975, N5973, N5888, N1420);
not NOT1 (N5976, N5974);
nand NAND2 (N5977, N5975, N205);
nand NAND2 (N5978, N5948, N3755);
not NOT1 (N5979, N5970);
and AND2 (N5980, N5971, N4761);
nor NOR3 (N5981, N5968, N384, N1228);
xor XOR2 (N5982, N5978, N5800);
or OR4 (N5983, N5944, N173, N2872, N2270);
buf BUF1 (N5984, N5956);
xor XOR2 (N5985, N5980, N3616);
not NOT1 (N5986, N5977);
or OR3 (N5987, N5985, N332, N963);
xor XOR2 (N5988, N5979, N1271);
buf BUF1 (N5989, N5966);
or OR2 (N5990, N5988, N1374);
not NOT1 (N5991, N5987);
nor NOR3 (N5992, N5989, N4604, N3819);
or OR3 (N5993, N5976, N5625, N2256);
nand NAND3 (N5994, N5986, N5699, N5754);
nand NAND4 (N5995, N5981, N5903, N934, N3911);
or OR4 (N5996, N5994, N4882, N601, N2076);
or OR2 (N5997, N5984, N2708);
not NOT1 (N5998, N5991);
xor XOR2 (N5999, N5993, N393);
xor XOR2 (N6000, N5972, N3883);
nand NAND2 (N6001, N5990, N3565);
buf BUF1 (N6002, N6000);
nor NOR2 (N6003, N6001, N4328);
nor NOR4 (N6004, N5995, N1457, N4149, N3341);
xor XOR2 (N6005, N5998, N4277);
and AND2 (N6006, N5983, N1542);
and AND2 (N6007, N6003, N5118);
xor XOR2 (N6008, N5996, N5411);
or OR2 (N6009, N6007, N2260);
buf BUF1 (N6010, N6005);
not NOT1 (N6011, N6010);
and AND3 (N6012, N6011, N2207, N5894);
nor NOR4 (N6013, N6006, N2933, N5851, N5673);
or OR2 (N6014, N5999, N3242);
not NOT1 (N6015, N6009);
nand NAND4 (N6016, N6004, N1006, N2889, N3900);
and AND2 (N6017, N6015, N2401);
nor NOR4 (N6018, N5997, N929, N2185, N4310);
nand NAND3 (N6019, N6014, N184, N1867);
or OR2 (N6020, N6012, N1982);
buf BUF1 (N6021, N5992);
or OR2 (N6022, N6019, N109);
not NOT1 (N6023, N6002);
or OR3 (N6024, N6016, N2970, N1940);
and AND2 (N6025, N6021, N106);
nand NAND3 (N6026, N6023, N499, N5968);
and AND2 (N6027, N6018, N2686);
nand NAND2 (N6028, N5982, N2845);
not NOT1 (N6029, N6020);
and AND2 (N6030, N6008, N5458);
and AND2 (N6031, N6027, N5284);
nand NAND2 (N6032, N6031, N5416);
buf BUF1 (N6033, N6032);
not NOT1 (N6034, N6026);
or OR4 (N6035, N6034, N4749, N5288, N4916);
not NOT1 (N6036, N6022);
not NOT1 (N6037, N6025);
or OR4 (N6038, N6036, N190, N4997, N3740);
xor XOR2 (N6039, N6029, N5824);
nand NAND3 (N6040, N6039, N5888, N3865);
xor XOR2 (N6041, N6035, N4820);
nand NAND2 (N6042, N6028, N5132);
xor XOR2 (N6043, N6024, N1712);
xor XOR2 (N6044, N6041, N2215);
buf BUF1 (N6045, N6013);
and AND3 (N6046, N6033, N2166, N3853);
and AND4 (N6047, N6030, N4079, N1260, N5876);
buf BUF1 (N6048, N6045);
buf BUF1 (N6049, N6043);
or OR4 (N6050, N6040, N3389, N2917, N1895);
buf BUF1 (N6051, N6038);
nor NOR3 (N6052, N6047, N4587, N5727);
xor XOR2 (N6053, N6046, N5580);
nor NOR4 (N6054, N6017, N2666, N2870, N4530);
buf BUF1 (N6055, N6037);
buf BUF1 (N6056, N6049);
buf BUF1 (N6057, N6055);
buf BUF1 (N6058, N6052);
not NOT1 (N6059, N6057);
nor NOR4 (N6060, N6044, N2814, N3116, N308);
xor XOR2 (N6061, N6053, N4558);
not NOT1 (N6062, N6060);
buf BUF1 (N6063, N6051);
nor NOR2 (N6064, N6054, N1981);
not NOT1 (N6065, N6059);
and AND4 (N6066, N6056, N3155, N2220, N4418);
xor XOR2 (N6067, N6050, N5718);
buf BUF1 (N6068, N6042);
xor XOR2 (N6069, N6063, N5138);
buf BUF1 (N6070, N6069);
not NOT1 (N6071, N6048);
buf BUF1 (N6072, N6061);
nand NAND3 (N6073, N6058, N5347, N889);
or OR3 (N6074, N6071, N2933, N5144);
not NOT1 (N6075, N6062);
nand NAND2 (N6076, N6072, N3134);
xor XOR2 (N6077, N6064, N679);
or OR3 (N6078, N6067, N5343, N4939);
or OR4 (N6079, N6065, N810, N5061, N2073);
xor XOR2 (N6080, N6073, N2569);
nor NOR3 (N6081, N6074, N5106, N3627);
xor XOR2 (N6082, N6070, N2974);
xor XOR2 (N6083, N6077, N5266);
or OR3 (N6084, N6066, N3136, N404);
nor NOR3 (N6085, N6082, N1825, N4161);
or OR2 (N6086, N6085, N1269);
buf BUF1 (N6087, N6083);
or OR3 (N6088, N6079, N5418, N2475);
xor XOR2 (N6089, N6080, N4144);
or OR2 (N6090, N6068, N1570);
or OR4 (N6091, N6081, N180, N1616, N1048);
nand NAND3 (N6092, N6075, N1821, N3992);
xor XOR2 (N6093, N6091, N3981);
not NOT1 (N6094, N6093);
not NOT1 (N6095, N6084);
or OR3 (N6096, N6078, N5865, N5725);
xor XOR2 (N6097, N6092, N1765);
nand NAND4 (N6098, N6087, N5010, N1847, N4113);
not NOT1 (N6099, N6088);
xor XOR2 (N6100, N6096, N5046);
and AND3 (N6101, N6100, N12, N112);
nor NOR4 (N6102, N6094, N5229, N5016, N1080);
and AND4 (N6103, N6095, N1765, N1445, N1734);
buf BUF1 (N6104, N6101);
or OR2 (N6105, N6099, N5126);
nand NAND3 (N6106, N6089, N701, N5512);
and AND3 (N6107, N6098, N350, N1625);
nand NAND3 (N6108, N6076, N550, N1737);
xor XOR2 (N6109, N6108, N4471);
nor NOR2 (N6110, N6105, N1067);
nand NAND2 (N6111, N6110, N3539);
or OR3 (N6112, N6109, N3990, N3597);
buf BUF1 (N6113, N6107);
not NOT1 (N6114, N6090);
or OR3 (N6115, N6104, N1351, N1156);
or OR3 (N6116, N6114, N2598, N2924);
or OR4 (N6117, N6106, N2719, N2795, N3126);
or OR3 (N6118, N6111, N3913, N2510);
buf BUF1 (N6119, N6118);
buf BUF1 (N6120, N6113);
xor XOR2 (N6121, N6115, N1794);
or OR4 (N6122, N6103, N916, N1668, N4409);
buf BUF1 (N6123, N6086);
or OR4 (N6124, N6119, N341, N1016, N5950);
buf BUF1 (N6125, N6124);
xor XOR2 (N6126, N6122, N5459);
buf BUF1 (N6127, N6121);
buf BUF1 (N6128, N6097);
nand NAND3 (N6129, N6123, N2009, N5445);
nor NOR2 (N6130, N6117, N1398);
and AND2 (N6131, N6129, N3549);
xor XOR2 (N6132, N6120, N4205);
not NOT1 (N6133, N6132);
nor NOR2 (N6134, N6131, N4192);
buf BUF1 (N6135, N6128);
not NOT1 (N6136, N6102);
or OR3 (N6137, N6135, N4312, N1836);
and AND4 (N6138, N6137, N2099, N2876, N1798);
xor XOR2 (N6139, N6136, N380);
and AND3 (N6140, N6130, N2334, N1260);
not NOT1 (N6141, N6139);
nand NAND3 (N6142, N6134, N1995, N2589);
not NOT1 (N6143, N6126);
buf BUF1 (N6144, N6141);
buf BUF1 (N6145, N6127);
xor XOR2 (N6146, N6125, N2101);
not NOT1 (N6147, N6143);
buf BUF1 (N6148, N6116);
or OR2 (N6149, N6146, N2627);
nor NOR3 (N6150, N6144, N5028, N1383);
buf BUF1 (N6151, N6149);
nor NOR4 (N6152, N6138, N4679, N6107, N4595);
xor XOR2 (N6153, N6148, N2493);
not NOT1 (N6154, N6133);
nor NOR4 (N6155, N6140, N4344, N505, N4729);
not NOT1 (N6156, N6154);
buf BUF1 (N6157, N6152);
not NOT1 (N6158, N6156);
or OR3 (N6159, N6145, N3963, N2036);
not NOT1 (N6160, N6112);
buf BUF1 (N6161, N6160);
or OR3 (N6162, N6155, N554, N5210);
xor XOR2 (N6163, N6162, N794);
and AND2 (N6164, N6151, N2395);
not NOT1 (N6165, N6163);
not NOT1 (N6166, N6142);
not NOT1 (N6167, N6147);
and AND4 (N6168, N6164, N5853, N4086, N944);
nand NAND3 (N6169, N6167, N4167, N5276);
buf BUF1 (N6170, N6159);
buf BUF1 (N6171, N6168);
buf BUF1 (N6172, N6153);
not NOT1 (N6173, N6161);
or OR4 (N6174, N6158, N2999, N1771, N2694);
nor NOR2 (N6175, N6166, N3756);
nor NOR4 (N6176, N6157, N5832, N3280, N75);
or OR2 (N6177, N6165, N1432);
nand NAND2 (N6178, N6177, N5702);
xor XOR2 (N6179, N6178, N368);
buf BUF1 (N6180, N6174);
xor XOR2 (N6181, N6169, N5611);
buf BUF1 (N6182, N6150);
not NOT1 (N6183, N6181);
xor XOR2 (N6184, N6175, N157);
or OR4 (N6185, N6180, N1222, N1789, N4543);
and AND3 (N6186, N6171, N170, N3324);
xor XOR2 (N6187, N6186, N3041);
not NOT1 (N6188, N6170);
and AND3 (N6189, N6176, N4162, N3717);
xor XOR2 (N6190, N6185, N2096);
nand NAND4 (N6191, N6187, N5834, N4365, N3749);
nand NAND2 (N6192, N6190, N3393);
and AND3 (N6193, N6189, N1196, N4218);
buf BUF1 (N6194, N6193);
nor NOR3 (N6195, N6194, N5285, N428);
xor XOR2 (N6196, N6183, N1651);
xor XOR2 (N6197, N6188, N124);
not NOT1 (N6198, N6192);
and AND2 (N6199, N6172, N4080);
xor XOR2 (N6200, N6179, N2310);
or OR3 (N6201, N6200, N3966, N3377);
or OR3 (N6202, N6182, N5818, N1301);
nor NOR4 (N6203, N6184, N3215, N4501, N4262);
nor NOR3 (N6204, N6197, N654, N4202);
nor NOR2 (N6205, N6202, N3309);
and AND3 (N6206, N6191, N4887, N1886);
nor NOR3 (N6207, N6206, N6018, N3372);
nand NAND3 (N6208, N6207, N4721, N3361);
nand NAND2 (N6209, N6201, N6116);
xor XOR2 (N6210, N6203, N4689);
not NOT1 (N6211, N6204);
and AND2 (N6212, N6173, N3297);
and AND3 (N6213, N6199, N2615, N1571);
buf BUF1 (N6214, N6195);
nand NAND4 (N6215, N6211, N3664, N5520, N3977);
not NOT1 (N6216, N6198);
nand NAND2 (N6217, N6196, N3654);
nor NOR2 (N6218, N6216, N3394);
buf BUF1 (N6219, N6208);
and AND4 (N6220, N6215, N2896, N5470, N4571);
xor XOR2 (N6221, N6212, N3377);
xor XOR2 (N6222, N6210, N3733);
xor XOR2 (N6223, N6217, N4122);
and AND3 (N6224, N6222, N110, N5845);
xor XOR2 (N6225, N6220, N72);
or OR4 (N6226, N6213, N4683, N3688, N5913);
or OR2 (N6227, N6224, N3875);
not NOT1 (N6228, N6225);
buf BUF1 (N6229, N6219);
nand NAND3 (N6230, N6221, N3814, N6086);
nand NAND4 (N6231, N6214, N3881, N1379, N2350);
or OR4 (N6232, N6223, N3449, N5523, N961);
nand NAND2 (N6233, N6229, N5693);
and AND2 (N6234, N6232, N5550);
xor XOR2 (N6235, N6218, N397);
nor NOR3 (N6236, N6235, N3821, N5667);
xor XOR2 (N6237, N6233, N4008);
and AND3 (N6238, N6230, N1550, N4223);
nor NOR2 (N6239, N6227, N3964);
and AND2 (N6240, N6228, N4091);
buf BUF1 (N6241, N6234);
nor NOR4 (N6242, N6241, N1295, N4424, N2702);
nand NAND2 (N6243, N6236, N3383);
not NOT1 (N6244, N6239);
or OR3 (N6245, N6231, N1446, N5951);
xor XOR2 (N6246, N6242, N3577);
or OR2 (N6247, N6243, N5062);
nand NAND3 (N6248, N6244, N934, N2843);
xor XOR2 (N6249, N6247, N1360);
nor NOR2 (N6250, N6226, N607);
not NOT1 (N6251, N6249);
nor NOR2 (N6252, N6251, N4615);
nor NOR3 (N6253, N6205, N4830, N1797);
nor NOR4 (N6254, N6253, N1989, N5087, N5387);
or OR2 (N6255, N6246, N5324);
xor XOR2 (N6256, N6238, N1957);
not NOT1 (N6257, N6250);
and AND4 (N6258, N6252, N5146, N5547, N3866);
xor XOR2 (N6259, N6254, N1692);
not NOT1 (N6260, N6240);
xor XOR2 (N6261, N6248, N6259);
or OR2 (N6262, N4691, N2219);
nand NAND3 (N6263, N6237, N1370, N5624);
not NOT1 (N6264, N6258);
or OR2 (N6265, N6261, N6020);
or OR3 (N6266, N6245, N1754, N4423);
nor NOR3 (N6267, N6263, N2005, N3374);
or OR2 (N6268, N6256, N5119);
nand NAND2 (N6269, N6260, N829);
and AND3 (N6270, N6257, N3899, N725);
buf BUF1 (N6271, N6265);
or OR2 (N6272, N6262, N2372);
buf BUF1 (N6273, N6255);
nand NAND2 (N6274, N6269, N3284);
nor NOR4 (N6275, N6271, N5325, N3547, N3335);
xor XOR2 (N6276, N6264, N4673);
nor NOR3 (N6277, N6266, N4580, N5926);
xor XOR2 (N6278, N6273, N1343);
nor NOR2 (N6279, N6274, N2544);
buf BUF1 (N6280, N6276);
nand NAND4 (N6281, N6270, N3525, N3556, N684);
buf BUF1 (N6282, N6267);
nor NOR2 (N6283, N6275, N928);
xor XOR2 (N6284, N6209, N1023);
xor XOR2 (N6285, N6272, N6111);
and AND3 (N6286, N6279, N5211, N2790);
and AND2 (N6287, N6268, N5084);
xor XOR2 (N6288, N6283, N5870);
xor XOR2 (N6289, N6285, N5181);
not NOT1 (N6290, N6277);
xor XOR2 (N6291, N6286, N3397);
nand NAND2 (N6292, N6291, N4688);
nand NAND2 (N6293, N6290, N2961);
xor XOR2 (N6294, N6284, N2622);
and AND3 (N6295, N6287, N1542, N981);
nand NAND2 (N6296, N6289, N4376);
nor NOR3 (N6297, N6282, N1117, N3138);
xor XOR2 (N6298, N6280, N6064);
or OR2 (N6299, N6281, N2258);
nor NOR2 (N6300, N6288, N4561);
not NOT1 (N6301, N6292);
xor XOR2 (N6302, N6278, N3364);
not NOT1 (N6303, N6295);
not NOT1 (N6304, N6302);
xor XOR2 (N6305, N6301, N6046);
and AND4 (N6306, N6305, N2384, N4202, N1896);
and AND2 (N6307, N6298, N3576);
not NOT1 (N6308, N6297);
nor NOR4 (N6309, N6294, N863, N6159, N671);
nor NOR4 (N6310, N6304, N3698, N4551, N1906);
buf BUF1 (N6311, N6306);
nor NOR3 (N6312, N6303, N5438, N6253);
not NOT1 (N6313, N6307);
or OR2 (N6314, N6309, N3579);
or OR4 (N6315, N6296, N6310, N1808, N3305);
nand NAND4 (N6316, N540, N1271, N872, N607);
xor XOR2 (N6317, N6300, N3428);
nor NOR2 (N6318, N6311, N165);
or OR4 (N6319, N6315, N3177, N4492, N3939);
or OR3 (N6320, N6293, N3376, N4784);
and AND4 (N6321, N6319, N1236, N2668, N4661);
nor NOR2 (N6322, N6313, N4074);
nor NOR4 (N6323, N6312, N5331, N5910, N5439);
nand NAND4 (N6324, N6321, N6049, N2744, N2760);
not NOT1 (N6325, N6314);
xor XOR2 (N6326, N6323, N3856);
not NOT1 (N6327, N6322);
buf BUF1 (N6328, N6320);
not NOT1 (N6329, N6325);
and AND3 (N6330, N6329, N736, N383);
not NOT1 (N6331, N6326);
buf BUF1 (N6332, N6318);
not NOT1 (N6333, N6316);
xor XOR2 (N6334, N6299, N1493);
not NOT1 (N6335, N6317);
nor NOR3 (N6336, N6328, N3791, N4968);
nand NAND3 (N6337, N6333, N1645, N3468);
nand NAND2 (N6338, N6334, N1361);
and AND3 (N6339, N6337, N228, N2054);
and AND2 (N6340, N6331, N1599);
not NOT1 (N6341, N6330);
not NOT1 (N6342, N6341);
nand NAND3 (N6343, N6342, N86, N2900);
buf BUF1 (N6344, N6340);
nand NAND3 (N6345, N6324, N2051, N3710);
buf BUF1 (N6346, N6308);
buf BUF1 (N6347, N6344);
nand NAND4 (N6348, N6339, N2974, N3480, N493);
buf BUF1 (N6349, N6336);
not NOT1 (N6350, N6332);
nor NOR3 (N6351, N6327, N1722, N257);
buf BUF1 (N6352, N6338);
xor XOR2 (N6353, N6335, N6011);
nor NOR2 (N6354, N6343, N789);
buf BUF1 (N6355, N6350);
not NOT1 (N6356, N6349);
not NOT1 (N6357, N6353);
nor NOR2 (N6358, N6354, N6276);
xor XOR2 (N6359, N6352, N1020);
nand NAND3 (N6360, N6351, N5097, N3938);
and AND4 (N6361, N6347, N4749, N1776, N2273);
xor XOR2 (N6362, N6358, N1789);
nand NAND4 (N6363, N6360, N3100, N4563, N5374);
xor XOR2 (N6364, N6355, N3467);
buf BUF1 (N6365, N6357);
or OR2 (N6366, N6345, N6050);
nor NOR2 (N6367, N6359, N2857);
not NOT1 (N6368, N6367);
nand NAND2 (N6369, N6348, N1145);
buf BUF1 (N6370, N6369);
nor NOR4 (N6371, N6356, N3051, N1708, N3312);
nand NAND3 (N6372, N6361, N1884, N5699);
xor XOR2 (N6373, N6366, N5197);
xor XOR2 (N6374, N6372, N1629);
xor XOR2 (N6375, N6362, N5634);
nor NOR3 (N6376, N6364, N2892, N3488);
nand NAND2 (N6377, N6363, N745);
xor XOR2 (N6378, N6373, N5686);
or OR2 (N6379, N6374, N895);
buf BUF1 (N6380, N6365);
and AND3 (N6381, N6379, N5860, N844);
or OR4 (N6382, N6376, N3278, N1030, N1632);
nand NAND2 (N6383, N6378, N3794);
not NOT1 (N6384, N6375);
buf BUF1 (N6385, N6383);
buf BUF1 (N6386, N6381);
or OR2 (N6387, N6384, N439);
not NOT1 (N6388, N6380);
or OR3 (N6389, N6385, N4689, N1752);
not NOT1 (N6390, N6389);
nor NOR3 (N6391, N6368, N587, N3346);
and AND4 (N6392, N6390, N985, N4604, N977);
not NOT1 (N6393, N6392);
xor XOR2 (N6394, N6387, N4454);
nor NOR4 (N6395, N6388, N3444, N690, N4841);
nand NAND3 (N6396, N6346, N3154, N5781);
buf BUF1 (N6397, N6394);
and AND2 (N6398, N6382, N4559);
or OR4 (N6399, N6398, N4401, N4598, N1778);
not NOT1 (N6400, N6377);
nor NOR4 (N6401, N6386, N2974, N5081, N812);
or OR4 (N6402, N6371, N513, N3451, N1614);
xor XOR2 (N6403, N6395, N3508);
xor XOR2 (N6404, N6401, N2471);
xor XOR2 (N6405, N6396, N1132);
buf BUF1 (N6406, N6393);
or OR3 (N6407, N6405, N772, N5649);
and AND3 (N6408, N6403, N1420, N3080);
and AND4 (N6409, N6399, N2202, N3175, N89);
or OR3 (N6410, N6391, N4775, N806);
nor NOR4 (N6411, N6406, N95, N4787, N2605);
buf BUF1 (N6412, N6410);
buf BUF1 (N6413, N6407);
or OR2 (N6414, N6397, N5697);
xor XOR2 (N6415, N6409, N1039);
nand NAND3 (N6416, N6404, N4959, N2643);
xor XOR2 (N6417, N6413, N4892);
not NOT1 (N6418, N6400);
xor XOR2 (N6419, N6411, N1206);
not NOT1 (N6420, N6416);
nor NOR4 (N6421, N6418, N569, N5747, N3318);
and AND2 (N6422, N6408, N5924);
buf BUF1 (N6423, N6421);
or OR2 (N6424, N6412, N4641);
nor NOR3 (N6425, N6417, N931, N2880);
nor NOR4 (N6426, N6414, N3878, N1309, N2526);
nor NOR2 (N6427, N6420, N3264);
nand NAND2 (N6428, N6425, N4309);
or OR3 (N6429, N6427, N2933, N1872);
not NOT1 (N6430, N6423);
xor XOR2 (N6431, N6422, N5540);
buf BUF1 (N6432, N6430);
not NOT1 (N6433, N6426);
or OR4 (N6434, N6428, N5831, N2910, N1003);
buf BUF1 (N6435, N6429);
nor NOR3 (N6436, N6433, N71, N426);
or OR4 (N6437, N6432, N3936, N5451, N3330);
not NOT1 (N6438, N6424);
buf BUF1 (N6439, N6437);
nor NOR3 (N6440, N6434, N5131, N3396);
nand NAND2 (N6441, N6438, N4510);
nand NAND3 (N6442, N6370, N5695, N1595);
not NOT1 (N6443, N6439);
nand NAND4 (N6444, N6442, N5038, N5219, N198);
buf BUF1 (N6445, N6419);
xor XOR2 (N6446, N6435, N388);
not NOT1 (N6447, N6436);
nand NAND3 (N6448, N6447, N1304, N1700);
or OR3 (N6449, N6415, N2729, N4911);
nand NAND4 (N6450, N6444, N2116, N1844, N6022);
nand NAND2 (N6451, N6440, N6207);
nor NOR2 (N6452, N6451, N3563);
nand NAND3 (N6453, N6402, N4493, N4222);
xor XOR2 (N6454, N6441, N3586);
and AND4 (N6455, N6431, N5392, N6439, N1601);
nor NOR3 (N6456, N6443, N324, N5367);
and AND4 (N6457, N6454, N2973, N774, N4218);
not NOT1 (N6458, N6448);
and AND2 (N6459, N6457, N1012);
not NOT1 (N6460, N6449);
and AND4 (N6461, N6452, N4718, N1137, N2822);
nand NAND4 (N6462, N6445, N1230, N2186, N1646);
or OR4 (N6463, N6459, N1885, N3534, N5225);
or OR2 (N6464, N6446, N6034);
nor NOR2 (N6465, N6453, N2822);
not NOT1 (N6466, N6456);
buf BUF1 (N6467, N6464);
not NOT1 (N6468, N6463);
not NOT1 (N6469, N6466);
buf BUF1 (N6470, N6467);
nand NAND3 (N6471, N6470, N5856, N5796);
nor NOR2 (N6472, N6461, N432);
not NOT1 (N6473, N6462);
or OR4 (N6474, N6469, N4922, N5573, N5173);
not NOT1 (N6475, N6458);
and AND2 (N6476, N6475, N4017);
not NOT1 (N6477, N6473);
or OR2 (N6478, N6460, N5638);
nor NOR2 (N6479, N6455, N2782);
nor NOR3 (N6480, N6474, N1751, N5572);
nand NAND2 (N6481, N6479, N4182);
nand NAND3 (N6482, N6478, N6076, N1252);
and AND3 (N6483, N6481, N1657, N3892);
not NOT1 (N6484, N6476);
buf BUF1 (N6485, N6482);
not NOT1 (N6486, N6450);
nand NAND4 (N6487, N6472, N4767, N5770, N419);
or OR3 (N6488, N6465, N1220, N3998);
nand NAND4 (N6489, N6477, N2468, N1041, N426);
nor NOR3 (N6490, N6483, N3171, N4785);
nor NOR3 (N6491, N6471, N5949, N3908);
nand NAND3 (N6492, N6480, N6328, N564);
not NOT1 (N6493, N6488);
and AND4 (N6494, N6468, N4561, N4550, N5610);
and AND2 (N6495, N6484, N226);
nand NAND4 (N6496, N6490, N3249, N4928, N2001);
buf BUF1 (N6497, N6486);
nand NAND4 (N6498, N6497, N4781, N1893, N1733);
xor XOR2 (N6499, N6489, N5640);
buf BUF1 (N6500, N6496);
xor XOR2 (N6501, N6493, N595);
buf BUF1 (N6502, N6495);
or OR3 (N6503, N6494, N2158, N3477);
buf BUF1 (N6504, N6500);
and AND4 (N6505, N6504, N2205, N2507, N5129);
or OR4 (N6506, N6505, N1593, N5053, N2429);
nand NAND4 (N6507, N6501, N962, N3546, N3396);
and AND3 (N6508, N6506, N3985, N217);
not NOT1 (N6509, N6485);
not NOT1 (N6510, N6508);
nor NOR4 (N6511, N6491, N4407, N699, N4348);
nand NAND3 (N6512, N6492, N2656, N5331);
and AND4 (N6513, N6509, N5649, N3572, N2821);
buf BUF1 (N6514, N6510);
buf BUF1 (N6515, N6513);
and AND4 (N6516, N6498, N4910, N2053, N2394);
nor NOR2 (N6517, N6511, N3509);
buf BUF1 (N6518, N6512);
nor NOR4 (N6519, N6507, N1493, N3364, N1609);
and AND4 (N6520, N6518, N4737, N2273, N4751);
not NOT1 (N6521, N6515);
nor NOR4 (N6522, N6487, N360, N946, N5688);
xor XOR2 (N6523, N6503, N871);
buf BUF1 (N6524, N6523);
nand NAND3 (N6525, N6502, N6065, N2576);
not NOT1 (N6526, N6524);
or OR3 (N6527, N6522, N2, N2807);
xor XOR2 (N6528, N6499, N4668);
nand NAND2 (N6529, N6526, N6240);
nor NOR4 (N6530, N6519, N2795, N2024, N5108);
not NOT1 (N6531, N6527);
xor XOR2 (N6532, N6516, N4934);
not NOT1 (N6533, N6525);
and AND4 (N6534, N6514, N4928, N1083, N6358);
nand NAND4 (N6535, N6530, N1464, N573, N1593);
not NOT1 (N6536, N6529);
nand NAND2 (N6537, N6534, N5429);
nand NAND4 (N6538, N6528, N750, N2732, N5959);
nor NOR3 (N6539, N6538, N6284, N152);
not NOT1 (N6540, N6533);
nor NOR3 (N6541, N6531, N194, N6359);
buf BUF1 (N6542, N6520);
or OR2 (N6543, N6535, N2866);
xor XOR2 (N6544, N6517, N4116);
nor NOR4 (N6545, N6536, N3381, N3618, N3453);
and AND3 (N6546, N6542, N917, N4456);
and AND3 (N6547, N6540, N1290, N1163);
nor NOR4 (N6548, N6545, N5380, N3989, N632);
nand NAND4 (N6549, N6548, N3796, N2888, N5064);
not NOT1 (N6550, N6544);
not NOT1 (N6551, N6550);
nand NAND4 (N6552, N6547, N1439, N2041, N1833);
or OR2 (N6553, N6543, N5727);
nor NOR3 (N6554, N6537, N3476, N6224);
or OR2 (N6555, N6521, N3200);
buf BUF1 (N6556, N6555);
or OR4 (N6557, N6541, N1691, N1919, N3168);
buf BUF1 (N6558, N6553);
nand NAND3 (N6559, N6539, N5622, N1245);
and AND3 (N6560, N6556, N6371, N2394);
nor NOR2 (N6561, N6557, N4400);
xor XOR2 (N6562, N6561, N4457);
buf BUF1 (N6563, N6560);
not NOT1 (N6564, N6549);
not NOT1 (N6565, N6563);
and AND3 (N6566, N6546, N1851, N3091);
xor XOR2 (N6567, N6566, N4484);
nand NAND3 (N6568, N6564, N690, N1683);
xor XOR2 (N6569, N6551, N1435);
and AND3 (N6570, N6532, N5958, N3515);
or OR2 (N6571, N6569, N4692);
or OR3 (N6572, N6565, N784, N2908);
nand NAND3 (N6573, N6571, N4447, N2646);
not NOT1 (N6574, N6558);
and AND2 (N6575, N6552, N4934);
not NOT1 (N6576, N6559);
not NOT1 (N6577, N6568);
nand NAND4 (N6578, N6573, N430, N5212, N173);
xor XOR2 (N6579, N6577, N5130);
buf BUF1 (N6580, N6576);
xor XOR2 (N6581, N6575, N2308);
or OR2 (N6582, N6578, N3883);
buf BUF1 (N6583, N6580);
or OR4 (N6584, N6567, N2029, N1204, N4436);
or OR4 (N6585, N6581, N1505, N2798, N4357);
xor XOR2 (N6586, N6574, N1472);
not NOT1 (N6587, N6583);
xor XOR2 (N6588, N6585, N6096);
nand NAND2 (N6589, N6570, N3519);
xor XOR2 (N6590, N6562, N4989);
nand NAND2 (N6591, N6582, N6522);
and AND2 (N6592, N6590, N6449);
xor XOR2 (N6593, N6579, N696);
nand NAND2 (N6594, N6587, N5928);
and AND2 (N6595, N6588, N2293);
not NOT1 (N6596, N6592);
nand NAND2 (N6597, N6593, N2073);
nor NOR4 (N6598, N6589, N5764, N4275, N5672);
or OR2 (N6599, N6572, N2605);
buf BUF1 (N6600, N6554);
not NOT1 (N6601, N6584);
buf BUF1 (N6602, N6594);
or OR4 (N6603, N6597, N192, N1483, N6372);
and AND4 (N6604, N6591, N5755, N882, N6298);
or OR4 (N6605, N6596, N1688, N2198, N4443);
not NOT1 (N6606, N6604);
or OR4 (N6607, N6606, N2356, N5313, N1112);
nand NAND2 (N6608, N6603, N3565);
xor XOR2 (N6609, N6602, N354);
buf BUF1 (N6610, N6607);
nor NOR4 (N6611, N6608, N5019, N5676, N3299);
xor XOR2 (N6612, N6595, N4992);
xor XOR2 (N6613, N6586, N777);
and AND3 (N6614, N6612, N1044, N1704);
xor XOR2 (N6615, N6611, N5704);
nor NOR2 (N6616, N6599, N4035);
xor XOR2 (N6617, N6614, N6469);
buf BUF1 (N6618, N6613);
buf BUF1 (N6619, N6610);
not NOT1 (N6620, N6616);
xor XOR2 (N6621, N6615, N2645);
or OR3 (N6622, N6600, N3205, N1925);
nand NAND3 (N6623, N6617, N6512, N4163);
or OR2 (N6624, N6623, N2585);
and AND3 (N6625, N6598, N2655, N777);
buf BUF1 (N6626, N6624);
buf BUF1 (N6627, N6618);
not NOT1 (N6628, N6601);
nand NAND4 (N6629, N6625, N6380, N3757, N6037);
buf BUF1 (N6630, N6628);
xor XOR2 (N6631, N6627, N4825);
nor NOR2 (N6632, N6631, N3535);
nand NAND4 (N6633, N6620, N870, N4875, N5609);
nand NAND3 (N6634, N6632, N6085, N4353);
and AND2 (N6635, N6630, N5442);
buf BUF1 (N6636, N6633);
nor NOR4 (N6637, N6636, N3679, N828, N5741);
and AND2 (N6638, N6621, N3767);
and AND3 (N6639, N6634, N4339, N6356);
nand NAND2 (N6640, N6638, N2885);
nand NAND2 (N6641, N6629, N6615);
or OR2 (N6642, N6641, N6199);
xor XOR2 (N6643, N6622, N5373);
xor XOR2 (N6644, N6643, N2356);
nor NOR2 (N6645, N6644, N85);
not NOT1 (N6646, N6635);
buf BUF1 (N6647, N6609);
not NOT1 (N6648, N6646);
nor NOR4 (N6649, N6605, N3428, N534, N4519);
nand NAND3 (N6650, N6648, N2900, N3738);
xor XOR2 (N6651, N6637, N1764);
not NOT1 (N6652, N6649);
not NOT1 (N6653, N6642);
xor XOR2 (N6654, N6619, N5208);
buf BUF1 (N6655, N6654);
and AND3 (N6656, N6653, N2889, N2793);
nor NOR2 (N6657, N6639, N2152);
buf BUF1 (N6658, N6657);
not NOT1 (N6659, N6650);
xor XOR2 (N6660, N6626, N195);
or OR4 (N6661, N6660, N6337, N2708, N4788);
and AND2 (N6662, N6655, N2328);
or OR4 (N6663, N6651, N6537, N1429, N454);
or OR4 (N6664, N6647, N5822, N3025, N6337);
nand NAND3 (N6665, N6661, N311, N505);
nor NOR3 (N6666, N6665, N3066, N3636);
nor NOR2 (N6667, N6656, N3254);
xor XOR2 (N6668, N6659, N3097);
xor XOR2 (N6669, N6640, N3380);
nor NOR3 (N6670, N6663, N690, N2781);
not NOT1 (N6671, N6664);
xor XOR2 (N6672, N6667, N2892);
buf BUF1 (N6673, N6666);
xor XOR2 (N6674, N6669, N3398);
and AND2 (N6675, N6652, N4914);
or OR3 (N6676, N6674, N169, N6093);
buf BUF1 (N6677, N6662);
and AND2 (N6678, N6671, N2312);
nand NAND4 (N6679, N6672, N443, N695, N2727);
xor XOR2 (N6680, N6658, N4545);
nor NOR3 (N6681, N6668, N5070, N1244);
nand NAND2 (N6682, N6675, N3009);
buf BUF1 (N6683, N6678);
not NOT1 (N6684, N6681);
nand NAND4 (N6685, N6670, N537, N1401, N159);
xor XOR2 (N6686, N6684, N3083);
nor NOR3 (N6687, N6677, N300, N1621);
nor NOR2 (N6688, N6682, N6347);
or OR2 (N6689, N6683, N4299);
xor XOR2 (N6690, N6686, N4371);
and AND4 (N6691, N6676, N3446, N3753, N5242);
not NOT1 (N6692, N6691);
nor NOR2 (N6693, N6680, N2868);
not NOT1 (N6694, N6687);
and AND2 (N6695, N6679, N2007);
not NOT1 (N6696, N6692);
nand NAND3 (N6697, N6694, N2406, N696);
or OR4 (N6698, N6688, N5637, N6569, N1384);
nand NAND3 (N6699, N6698, N5213, N5050);
xor XOR2 (N6700, N6673, N4010);
and AND3 (N6701, N6685, N697, N4098);
nor NOR2 (N6702, N6690, N488);
buf BUF1 (N6703, N6702);
not NOT1 (N6704, N6695);
nand NAND4 (N6705, N6704, N2954, N4434, N302);
or OR2 (N6706, N6696, N2230);
buf BUF1 (N6707, N6645);
or OR2 (N6708, N6701, N1935);
nand NAND4 (N6709, N6699, N6234, N1412, N5833);
and AND4 (N6710, N6689, N1613, N225, N2997);
not NOT1 (N6711, N6710);
nor NOR2 (N6712, N6700, N970);
buf BUF1 (N6713, N6707);
xor XOR2 (N6714, N6708, N5237);
nand NAND3 (N6715, N6713, N6689, N1727);
or OR3 (N6716, N6697, N1184, N242);
nor NOR3 (N6717, N6703, N2763, N591);
not NOT1 (N6718, N6693);
buf BUF1 (N6719, N6715);
or OR2 (N6720, N6714, N345);
nand NAND2 (N6721, N6720, N6635);
nor NOR4 (N6722, N6706, N3244, N1762, N3996);
or OR4 (N6723, N6709, N4211, N1812, N3640);
nand NAND2 (N6724, N6711, N4480);
or OR3 (N6725, N6722, N770, N276);
and AND4 (N6726, N6718, N5686, N1976, N5132);
not NOT1 (N6727, N6712);
and AND3 (N6728, N6721, N4116, N6343);
and AND3 (N6729, N6725, N2410, N6153);
xor XOR2 (N6730, N6728, N4927);
not NOT1 (N6731, N6719);
nand NAND2 (N6732, N6723, N2734);
xor XOR2 (N6733, N6727, N1528);
xor XOR2 (N6734, N6731, N802);
not NOT1 (N6735, N6729);
xor XOR2 (N6736, N6726, N4912);
buf BUF1 (N6737, N6716);
nor NOR3 (N6738, N6732, N3483, N6210);
buf BUF1 (N6739, N6705);
nand NAND2 (N6740, N6736, N1847);
buf BUF1 (N6741, N6738);
xor XOR2 (N6742, N6717, N86);
buf BUF1 (N6743, N6735);
nor NOR3 (N6744, N6741, N3126, N3919);
and AND4 (N6745, N6730, N712, N913, N351);
xor XOR2 (N6746, N6742, N1316);
nor NOR3 (N6747, N6734, N3438, N2151);
and AND2 (N6748, N6746, N2772);
or OR4 (N6749, N6724, N5534, N238, N6188);
nand NAND3 (N6750, N6745, N2557, N2912);
or OR2 (N6751, N6740, N1712);
xor XOR2 (N6752, N6744, N4417);
nor NOR2 (N6753, N6752, N3078);
nor NOR2 (N6754, N6751, N3293);
buf BUF1 (N6755, N6737);
not NOT1 (N6756, N6750);
xor XOR2 (N6757, N6749, N6507);
nand NAND4 (N6758, N6747, N1708, N1823, N1300);
buf BUF1 (N6759, N6756);
xor XOR2 (N6760, N6753, N1602);
and AND3 (N6761, N6754, N4677, N3348);
not NOT1 (N6762, N6758);
nor NOR2 (N6763, N6748, N5513);
nand NAND4 (N6764, N6743, N4015, N3430, N6246);
nand NAND2 (N6765, N6762, N125);
buf BUF1 (N6766, N6739);
or OR3 (N6767, N6761, N2490, N5507);
not NOT1 (N6768, N6765);
xor XOR2 (N6769, N6766, N387);
nand NAND4 (N6770, N6768, N6717, N5651, N2434);
nand NAND2 (N6771, N6733, N2793);
and AND3 (N6772, N6755, N2589, N4254);
and AND3 (N6773, N6771, N4568, N5479);
and AND3 (N6774, N6772, N4788, N1674);
not NOT1 (N6775, N6767);
and AND4 (N6776, N6763, N1289, N5319, N6419);
buf BUF1 (N6777, N6773);
or OR3 (N6778, N6759, N301, N6104);
nor NOR2 (N6779, N6769, N4781);
or OR3 (N6780, N6770, N5718, N5558);
nor NOR3 (N6781, N6775, N6139, N4976);
nand NAND3 (N6782, N6777, N726, N3559);
nand NAND2 (N6783, N6760, N1436);
nor NOR4 (N6784, N6764, N6089, N3557, N3554);
nand NAND3 (N6785, N6784, N4826, N4634);
or OR3 (N6786, N6774, N294, N3057);
nand NAND4 (N6787, N6785, N3719, N5686, N4674);
or OR4 (N6788, N6782, N2109, N5611, N2812);
nand NAND3 (N6789, N6783, N6203, N3389);
and AND2 (N6790, N6789, N4374);
nand NAND2 (N6791, N6776, N1290);
or OR2 (N6792, N6780, N2883);
buf BUF1 (N6793, N6791);
buf BUF1 (N6794, N6786);
or OR2 (N6795, N6787, N2873);
nor NOR2 (N6796, N6795, N6227);
not NOT1 (N6797, N6788);
and AND3 (N6798, N6778, N1455, N3028);
nand NAND4 (N6799, N6796, N5401, N3508, N830);
nand NAND4 (N6800, N6797, N1398, N3370, N5919);
nand NAND4 (N6801, N6757, N2539, N4294, N4659);
and AND4 (N6802, N6800, N5381, N2212, N5355);
buf BUF1 (N6803, N6801);
xor XOR2 (N6804, N6792, N1029);
nand NAND3 (N6805, N6803, N1040, N6514);
nand NAND4 (N6806, N6798, N6105, N3616, N6277);
buf BUF1 (N6807, N6799);
and AND3 (N6808, N6802, N2349, N4843);
or OR3 (N6809, N6781, N760, N247);
xor XOR2 (N6810, N6808, N2473);
nand NAND4 (N6811, N6806, N2205, N6449, N1631);
nand NAND3 (N6812, N6811, N4640, N6178);
buf BUF1 (N6813, N6779);
nand NAND4 (N6814, N6810, N4832, N5520, N4869);
or OR2 (N6815, N6813, N236);
xor XOR2 (N6816, N6805, N10);
nor NOR3 (N6817, N6815, N3896, N6330);
not NOT1 (N6818, N6793);
nor NOR2 (N6819, N6818, N1215);
nor NOR3 (N6820, N6809, N3916, N6609);
nand NAND3 (N6821, N6804, N5197, N2901);
or OR3 (N6822, N6807, N31, N1910);
nor NOR4 (N6823, N6812, N1668, N1245, N3292);
nand NAND4 (N6824, N6821, N3443, N6268, N5262);
buf BUF1 (N6825, N6820);
buf BUF1 (N6826, N6814);
or OR2 (N6827, N6819, N6664);
xor XOR2 (N6828, N6794, N5696);
xor XOR2 (N6829, N6790, N3130);
nor NOR4 (N6830, N6829, N3712, N3329, N3725);
nand NAND4 (N6831, N6822, N6376, N835, N6537);
nand NAND3 (N6832, N6830, N5418, N1736);
xor XOR2 (N6833, N6832, N4295);
or OR3 (N6834, N6816, N4993, N704);
nand NAND4 (N6835, N6825, N2920, N804, N4088);
or OR4 (N6836, N6823, N3072, N5689, N2015);
nand NAND2 (N6837, N6834, N1053);
or OR3 (N6838, N6817, N6449, N1074);
buf BUF1 (N6839, N6833);
nand NAND3 (N6840, N6824, N6640, N534);
nor NOR4 (N6841, N6837, N4892, N2426, N2222);
not NOT1 (N6842, N6835);
buf BUF1 (N6843, N6838);
xor XOR2 (N6844, N6840, N219);
nor NOR4 (N6845, N6827, N6390, N5999, N2130);
nor NOR3 (N6846, N6836, N5648, N3288);
and AND3 (N6847, N6843, N4872, N6060);
and AND3 (N6848, N6826, N3181, N6636);
not NOT1 (N6849, N6846);
not NOT1 (N6850, N6845);
xor XOR2 (N6851, N6841, N4251);
not NOT1 (N6852, N6831);
not NOT1 (N6853, N6847);
and AND3 (N6854, N6852, N1474, N4589);
and AND3 (N6855, N6844, N1160, N186);
xor XOR2 (N6856, N6839, N5206);
not NOT1 (N6857, N6851);
xor XOR2 (N6858, N6853, N1045);
nand NAND3 (N6859, N6850, N1382, N3066);
buf BUF1 (N6860, N6859);
buf BUF1 (N6861, N6857);
buf BUF1 (N6862, N6860);
and AND2 (N6863, N6858, N3774);
nand NAND4 (N6864, N6842, N6034, N2441, N2205);
or OR3 (N6865, N6854, N663, N1995);
buf BUF1 (N6866, N6863);
and AND3 (N6867, N6849, N1724, N5900);
or OR2 (N6868, N6856, N1797);
or OR4 (N6869, N6862, N2709, N6784, N1606);
and AND3 (N6870, N6861, N555, N2558);
nand NAND4 (N6871, N6868, N5356, N2565, N601);
nor NOR3 (N6872, N6865, N6261, N2095);
not NOT1 (N6873, N6855);
xor XOR2 (N6874, N6871, N721);
nand NAND2 (N6875, N6869, N2993);
and AND3 (N6876, N6874, N936, N696);
not NOT1 (N6877, N6867);
not NOT1 (N6878, N6875);
xor XOR2 (N6879, N6848, N1957);
not NOT1 (N6880, N6879);
xor XOR2 (N6881, N6870, N4604);
nand NAND2 (N6882, N6880, N6564);
nand NAND4 (N6883, N6828, N1524, N4353, N3520);
xor XOR2 (N6884, N6876, N3672);
nand NAND4 (N6885, N6882, N5987, N2648, N2533);
nor NOR3 (N6886, N6878, N3219, N4659);
buf BUF1 (N6887, N6864);
xor XOR2 (N6888, N6877, N3937);
xor XOR2 (N6889, N6887, N4485);
or OR4 (N6890, N6889, N6134, N5271, N5877);
and AND2 (N6891, N6890, N2181);
xor XOR2 (N6892, N6881, N1883);
not NOT1 (N6893, N6873);
nor NOR2 (N6894, N6892, N1966);
nand NAND2 (N6895, N6893, N5206);
and AND4 (N6896, N6894, N2317, N5477, N4778);
not NOT1 (N6897, N6884);
nor NOR3 (N6898, N6897, N3875, N3965);
or OR3 (N6899, N6872, N1480, N5973);
nor NOR2 (N6900, N6866, N4472);
or OR2 (N6901, N6896, N621);
buf BUF1 (N6902, N6895);
or OR4 (N6903, N6898, N6268, N545, N1751);
buf BUF1 (N6904, N6886);
nand NAND4 (N6905, N6902, N1907, N609, N2446);
not NOT1 (N6906, N6901);
nor NOR4 (N6907, N6906, N4232, N2152, N49);
xor XOR2 (N6908, N6883, N5279);
buf BUF1 (N6909, N6891);
or OR2 (N6910, N6905, N3255);
not NOT1 (N6911, N6904);
nor NOR4 (N6912, N6909, N4452, N236, N352);
buf BUF1 (N6913, N6910);
or OR3 (N6914, N6912, N6113, N3261);
or OR3 (N6915, N6900, N4275, N4762);
or OR3 (N6916, N6908, N841, N2656);
and AND4 (N6917, N6899, N1539, N4498, N3725);
nand NAND2 (N6918, N6888, N1734);
and AND4 (N6919, N6913, N1165, N3889, N678);
xor XOR2 (N6920, N6915, N882);
nand NAND4 (N6921, N6920, N6267, N509, N1040);
xor XOR2 (N6922, N6885, N5892);
and AND2 (N6923, N6922, N2655);
nor NOR4 (N6924, N6907, N5299, N5335, N1712);
not NOT1 (N6925, N6903);
nor NOR3 (N6926, N6925, N6912, N3663);
nand NAND3 (N6927, N6914, N1552, N6584);
not NOT1 (N6928, N6917);
nor NOR2 (N6929, N6911, N1351);
or OR2 (N6930, N6928, N5445);
and AND3 (N6931, N6926, N497, N3026);
buf BUF1 (N6932, N6924);
buf BUF1 (N6933, N6923);
and AND2 (N6934, N6921, N3316);
and AND3 (N6935, N6916, N3131, N6897);
xor XOR2 (N6936, N6929, N3411);
not NOT1 (N6937, N6927);
buf BUF1 (N6938, N6935);
xor XOR2 (N6939, N6930, N6692);
buf BUF1 (N6940, N6931);
nor NOR3 (N6941, N6934, N4708, N5162);
and AND3 (N6942, N6933, N6334, N4088);
nor NOR3 (N6943, N6936, N3667, N6547);
nand NAND3 (N6944, N6940, N774, N6905);
xor XOR2 (N6945, N6942, N6012);
and AND3 (N6946, N6937, N6188, N642);
nor NOR4 (N6947, N6946, N5919, N5516, N244);
buf BUF1 (N6948, N6947);
nor NOR3 (N6949, N6919, N6450, N5464);
not NOT1 (N6950, N6938);
or OR4 (N6951, N6932, N4187, N4505, N5301);
or OR3 (N6952, N6944, N1791, N1743);
xor XOR2 (N6953, N6941, N2124);
buf BUF1 (N6954, N6950);
nand NAND3 (N6955, N6954, N6903, N936);
and AND2 (N6956, N6918, N635);
nor NOR4 (N6957, N6952, N5669, N2203, N357);
xor XOR2 (N6958, N6945, N126);
nand NAND3 (N6959, N6949, N4728, N532);
nand NAND4 (N6960, N6959, N1130, N5904, N1159);
nor NOR2 (N6961, N6956, N5809);
xor XOR2 (N6962, N6958, N5812);
nand NAND2 (N6963, N6943, N403);
buf BUF1 (N6964, N6961);
buf BUF1 (N6965, N6960);
nand NAND2 (N6966, N6965, N6175);
buf BUF1 (N6967, N6951);
nor NOR3 (N6968, N6962, N3936, N3812);
nor NOR2 (N6969, N6939, N1366);
or OR4 (N6970, N6964, N5193, N3403, N5710);
xor XOR2 (N6971, N6955, N132);
nand NAND4 (N6972, N6967, N2079, N5579, N1673);
or OR4 (N6973, N6963, N4000, N3224, N5398);
not NOT1 (N6974, N6968);
nand NAND4 (N6975, N6971, N449, N3738, N4637);
buf BUF1 (N6976, N6969);
nand NAND3 (N6977, N6974, N3457, N6111);
not NOT1 (N6978, N6966);
or OR4 (N6979, N6957, N4411, N1040, N2074);
buf BUF1 (N6980, N6970);
buf BUF1 (N6981, N6948);
or OR2 (N6982, N6953, N1978);
xor XOR2 (N6983, N6982, N540);
buf BUF1 (N6984, N6983);
nand NAND2 (N6985, N6976, N2680);
and AND2 (N6986, N6984, N1105);
or OR3 (N6987, N6980, N1283, N3412);
buf BUF1 (N6988, N6985);
nand NAND2 (N6989, N6975, N3693);
nor NOR3 (N6990, N6979, N5696, N2475);
xor XOR2 (N6991, N6986, N6743);
xor XOR2 (N6992, N6978, N4059);
and AND2 (N6993, N6977, N1012);
and AND4 (N6994, N6992, N3702, N5994, N3814);
xor XOR2 (N6995, N6990, N495);
not NOT1 (N6996, N6973);
nand NAND4 (N6997, N6989, N2074, N5425, N5857);
nand NAND4 (N6998, N6996, N6368, N2631, N4337);
buf BUF1 (N6999, N6981);
nor NOR4 (N7000, N6997, N5472, N733, N1526);
and AND4 (N7001, N6987, N85, N965, N5458);
xor XOR2 (N7002, N6993, N2849);
nor NOR3 (N7003, N6988, N6562, N773);
nor NOR3 (N7004, N6998, N4492, N777);
nand NAND3 (N7005, N6972, N1842, N3577);
and AND2 (N7006, N7004, N2591);
nand NAND4 (N7007, N7000, N6825, N6599, N3535);
buf BUF1 (N7008, N6995);
and AND2 (N7009, N7007, N1868);
not NOT1 (N7010, N7001);
buf BUF1 (N7011, N6999);
nor NOR4 (N7012, N7008, N6512, N4241, N6838);
and AND3 (N7013, N7010, N3548, N4441);
and AND4 (N7014, N7013, N4154, N5420, N977);
xor XOR2 (N7015, N7005, N968);
xor XOR2 (N7016, N7006, N1964);
xor XOR2 (N7017, N7002, N6460);
and AND4 (N7018, N7011, N2877, N4762, N3966);
nand NAND4 (N7019, N6994, N1160, N186, N1646);
xor XOR2 (N7020, N7017, N2731);
nor NOR3 (N7021, N7018, N6692, N324);
not NOT1 (N7022, N7019);
xor XOR2 (N7023, N7014, N806);
xor XOR2 (N7024, N6991, N4477);
or OR4 (N7025, N7023, N2290, N4475, N6821);
nor NOR2 (N7026, N7022, N4737);
not NOT1 (N7027, N7015);
nor NOR4 (N7028, N7025, N6207, N384, N4358);
nand NAND4 (N7029, N7020, N4320, N4139, N3116);
or OR2 (N7030, N7029, N6662);
nor NOR2 (N7031, N7003, N6358);
nand NAND4 (N7032, N7012, N4358, N2876, N1090);
or OR3 (N7033, N7024, N1295, N4941);
not NOT1 (N7034, N7026);
xor XOR2 (N7035, N7021, N1483);
or OR3 (N7036, N7009, N904, N5266);
nand NAND4 (N7037, N7016, N4854, N5924, N4266);
and AND4 (N7038, N7032, N6912, N5256, N1476);
or OR2 (N7039, N7030, N187);
nor NOR4 (N7040, N7028, N2378, N5627, N1848);
or OR2 (N7041, N7035, N2845);
nor NOR4 (N7042, N7034, N1719, N4884, N2510);
xor XOR2 (N7043, N7027, N6352);
nor NOR2 (N7044, N7043, N7035);
and AND2 (N7045, N7041, N5005);
buf BUF1 (N7046, N7045);
not NOT1 (N7047, N7040);
or OR3 (N7048, N7033, N2817, N1341);
buf BUF1 (N7049, N7037);
or OR2 (N7050, N7046, N6983);
xor XOR2 (N7051, N7031, N2580);
and AND4 (N7052, N7050, N5770, N2314, N2838);
and AND4 (N7053, N7049, N1792, N5399, N5824);
xor XOR2 (N7054, N7042, N2097);
not NOT1 (N7055, N7054);
not NOT1 (N7056, N7051);
buf BUF1 (N7057, N7053);
nor NOR2 (N7058, N7044, N4517);
nand NAND4 (N7059, N7038, N4354, N1047, N2838);
nand NAND4 (N7060, N7048, N1329, N4562, N853);
nor NOR4 (N7061, N7059, N5421, N6166, N1071);
xor XOR2 (N7062, N7057, N6339);
buf BUF1 (N7063, N7062);
buf BUF1 (N7064, N7056);
not NOT1 (N7065, N7060);
xor XOR2 (N7066, N7064, N1612);
or OR4 (N7067, N7055, N1665, N3673, N383);
buf BUF1 (N7068, N7039);
nor NOR4 (N7069, N7061, N2113, N2606, N2078);
not NOT1 (N7070, N7067);
or OR4 (N7071, N7070, N2980, N3999, N701);
nor NOR4 (N7072, N7071, N4599, N2095, N5942);
and AND2 (N7073, N7065, N3067);
xor XOR2 (N7074, N7058, N4081);
nor NOR2 (N7075, N7036, N3453);
buf BUF1 (N7076, N7047);
buf BUF1 (N7077, N7063);
xor XOR2 (N7078, N7052, N1607);
buf BUF1 (N7079, N7076);
xor XOR2 (N7080, N7069, N1165);
buf BUF1 (N7081, N7079);
nand NAND4 (N7082, N7078, N4867, N5785, N3740);
nor NOR4 (N7083, N7073, N4215, N25, N4539);
nand NAND2 (N7084, N7072, N1553);
nand NAND4 (N7085, N7074, N4970, N4246, N41);
nand NAND4 (N7086, N7085, N3848, N5277, N1775);
nor NOR3 (N7087, N7086, N4709, N2892);
nor NOR2 (N7088, N7075, N1451);
not NOT1 (N7089, N7066);
buf BUF1 (N7090, N7088);
buf BUF1 (N7091, N7087);
nand NAND3 (N7092, N7080, N6614, N4357);
not NOT1 (N7093, N7092);
xor XOR2 (N7094, N7068, N3612);
nand NAND3 (N7095, N7081, N4140, N875);
not NOT1 (N7096, N7094);
nand NAND3 (N7097, N7084, N3683, N1703);
and AND2 (N7098, N7089, N4829);
xor XOR2 (N7099, N7082, N2656);
buf BUF1 (N7100, N7097);
nor NOR4 (N7101, N7095, N3656, N3245, N1413);
nor NOR4 (N7102, N7091, N2223, N2643, N1810);
nor NOR2 (N7103, N7098, N2502);
and AND4 (N7104, N7093, N1495, N1800, N2763);
not NOT1 (N7105, N7096);
not NOT1 (N7106, N7083);
and AND2 (N7107, N7103, N72);
buf BUF1 (N7108, N7106);
and AND4 (N7109, N7090, N6586, N6368, N6731);
nand NAND4 (N7110, N7105, N6790, N5877, N6251);
not NOT1 (N7111, N7107);
or OR3 (N7112, N7104, N1983, N2429);
xor XOR2 (N7113, N7102, N2630);
not NOT1 (N7114, N7109);
not NOT1 (N7115, N7113);
nor NOR3 (N7116, N7114, N5354, N1984);
nor NOR4 (N7117, N7115, N3506, N4916, N5690);
nand NAND2 (N7118, N7117, N3004);
not NOT1 (N7119, N7101);
nor NOR3 (N7120, N7108, N4055, N2777);
and AND3 (N7121, N7110, N3768, N522);
nand NAND2 (N7122, N7116, N5888);
nand NAND4 (N7123, N7120, N887, N1593, N2917);
buf BUF1 (N7124, N7099);
not NOT1 (N7125, N7118);
or OR2 (N7126, N7123, N5350);
and AND4 (N7127, N7126, N4476, N2740, N5646);
or OR4 (N7128, N7112, N4598, N876, N4704);
nor NOR3 (N7129, N7127, N6746, N3967);
nand NAND4 (N7130, N7128, N3531, N304, N5282);
and AND3 (N7131, N7119, N6061, N4224);
not NOT1 (N7132, N7125);
xor XOR2 (N7133, N7100, N1416);
or OR4 (N7134, N7121, N5408, N5666, N3106);
and AND2 (N7135, N7122, N753);
and AND2 (N7136, N7077, N1605);
xor XOR2 (N7137, N7131, N15);
not NOT1 (N7138, N7134);
buf BUF1 (N7139, N7135);
nand NAND3 (N7140, N7133, N3862, N6843);
and AND2 (N7141, N7124, N1288);
buf BUF1 (N7142, N7136);
and AND2 (N7143, N7139, N6367);
buf BUF1 (N7144, N7141);
not NOT1 (N7145, N7111);
buf BUF1 (N7146, N7137);
nand NAND4 (N7147, N7132, N3243, N445, N3658);
or OR3 (N7148, N7144, N3757, N6263);
buf BUF1 (N7149, N7143);
nor NOR3 (N7150, N7142, N3674, N5775);
and AND2 (N7151, N7145, N5396);
nand NAND3 (N7152, N7150, N1610, N389);
xor XOR2 (N7153, N7152, N6656);
nor NOR2 (N7154, N7148, N6891);
not NOT1 (N7155, N7140);
nor NOR2 (N7156, N7151, N4682);
xor XOR2 (N7157, N7149, N4112);
and AND3 (N7158, N7146, N16, N4038);
xor XOR2 (N7159, N7153, N6273);
nor NOR3 (N7160, N7129, N4683, N321);
buf BUF1 (N7161, N7155);
not NOT1 (N7162, N7161);
nand NAND4 (N7163, N7160, N3640, N173, N1163);
and AND4 (N7164, N7163, N4527, N5659, N4939);
buf BUF1 (N7165, N7162);
and AND4 (N7166, N7147, N1127, N3018, N4386);
xor XOR2 (N7167, N7165, N4019);
or OR4 (N7168, N7158, N50, N5059, N4032);
not NOT1 (N7169, N7130);
and AND2 (N7170, N7166, N1702);
nand NAND3 (N7171, N7159, N1837, N6349);
nor NOR3 (N7172, N7157, N4635, N3619);
nor NOR2 (N7173, N7167, N3510);
xor XOR2 (N7174, N7164, N6258);
nor NOR3 (N7175, N7174, N3817, N6313);
or OR3 (N7176, N7154, N6353, N3391);
not NOT1 (N7177, N7169);
nand NAND2 (N7178, N7171, N824);
nand NAND4 (N7179, N7177, N2316, N2575, N5735);
and AND4 (N7180, N7172, N6681, N1552, N3369);
xor XOR2 (N7181, N7175, N4737);
nand NAND3 (N7182, N7178, N1259, N6879);
nor NOR3 (N7183, N7180, N7040, N4843);
xor XOR2 (N7184, N7183, N213);
nand NAND4 (N7185, N7179, N6190, N4138, N4997);
xor XOR2 (N7186, N7185, N3429);
not NOT1 (N7187, N7182);
nor NOR3 (N7188, N7168, N1474, N1894);
not NOT1 (N7189, N7138);
not NOT1 (N7190, N7170);
nand NAND3 (N7191, N7186, N849, N1166);
buf BUF1 (N7192, N7191);
and AND4 (N7193, N7188, N3941, N5331, N6593);
and AND3 (N7194, N7184, N3355, N1850);
nor NOR2 (N7195, N7181, N4588);
buf BUF1 (N7196, N7194);
nor NOR2 (N7197, N7187, N5396);
and AND3 (N7198, N7173, N3887, N3543);
nand NAND4 (N7199, N7189, N5563, N6119, N2136);
not NOT1 (N7200, N7198);
nand NAND2 (N7201, N7192, N2797);
nand NAND3 (N7202, N7199, N2151, N4206);
nor NOR3 (N7203, N7193, N6944, N275);
nor NOR3 (N7204, N7196, N3150, N5389);
and AND4 (N7205, N7190, N3581, N5610, N1411);
not NOT1 (N7206, N7203);
nand NAND4 (N7207, N7197, N5931, N1982, N926);
not NOT1 (N7208, N7204);
or OR4 (N7209, N7206, N32, N3697, N6007);
nand NAND2 (N7210, N7200, N4170);
xor XOR2 (N7211, N7195, N6892);
nor NOR3 (N7212, N7201, N4699, N6330);
not NOT1 (N7213, N7210);
not NOT1 (N7214, N7209);
nand NAND2 (N7215, N7176, N2057);
nor NOR4 (N7216, N7213, N842, N1761, N590);
or OR4 (N7217, N7215, N234, N4312, N6995);
and AND2 (N7218, N7216, N1233);
buf BUF1 (N7219, N7212);
or OR3 (N7220, N7214, N336, N1108);
nand NAND2 (N7221, N7202, N3114);
or OR2 (N7222, N7217, N3452);
not NOT1 (N7223, N7222);
buf BUF1 (N7224, N7205);
xor XOR2 (N7225, N7224, N5407);
buf BUF1 (N7226, N7220);
nand NAND4 (N7227, N7218, N3404, N6643, N3578);
nor NOR3 (N7228, N7223, N4841, N4501);
not NOT1 (N7229, N7221);
nand NAND3 (N7230, N7156, N886, N3521);
not NOT1 (N7231, N7227);
buf BUF1 (N7232, N7225);
nor NOR3 (N7233, N7226, N603, N66);
not NOT1 (N7234, N7211);
xor XOR2 (N7235, N7219, N1020);
not NOT1 (N7236, N7231);
not NOT1 (N7237, N7230);
and AND2 (N7238, N7229, N1157);
xor XOR2 (N7239, N7235, N6946);
nor NOR4 (N7240, N7234, N2733, N852, N4567);
nand NAND4 (N7241, N7232, N3253, N4291, N6402);
nand NAND2 (N7242, N7207, N951);
buf BUF1 (N7243, N7228);
nand NAND2 (N7244, N7233, N4064);
or OR4 (N7245, N7244, N6336, N1863, N189);
nand NAND2 (N7246, N7241, N1993);
not NOT1 (N7247, N7239);
nor NOR4 (N7248, N7247, N1811, N6401, N4942);
buf BUF1 (N7249, N7238);
or OR2 (N7250, N7242, N6162);
or OR4 (N7251, N7245, N2003, N1714, N512);
nor NOR4 (N7252, N7248, N5748, N5261, N959);
or OR3 (N7253, N7237, N5376, N6937);
or OR4 (N7254, N7253, N4731, N5285, N4873);
xor XOR2 (N7255, N7254, N891);
buf BUF1 (N7256, N7251);
not NOT1 (N7257, N7246);
nand NAND2 (N7258, N7236, N830);
nor NOR4 (N7259, N7258, N6361, N1339, N4565);
not NOT1 (N7260, N7255);
or OR2 (N7261, N7240, N7046);
and AND4 (N7262, N7252, N2798, N5155, N4475);
nor NOR2 (N7263, N7257, N1345);
xor XOR2 (N7264, N7262, N2411);
xor XOR2 (N7265, N7263, N171);
xor XOR2 (N7266, N7259, N1800);
nor NOR2 (N7267, N7208, N3142);
and AND4 (N7268, N7250, N3855, N6941, N5021);
buf BUF1 (N7269, N7256);
xor XOR2 (N7270, N7267, N3406);
or OR3 (N7271, N7269, N1903, N1771);
nand NAND4 (N7272, N7270, N3614, N6930, N1933);
or OR3 (N7273, N7260, N1776, N1840);
xor XOR2 (N7274, N7272, N314);
or OR3 (N7275, N7271, N4758, N986);
and AND4 (N7276, N7264, N6984, N5352, N3672);
nor NOR3 (N7277, N7261, N4228, N3646);
or OR4 (N7278, N7265, N5864, N4044, N2307);
or OR2 (N7279, N7277, N5523);
nor NOR2 (N7280, N7275, N1487);
buf BUF1 (N7281, N7274);
or OR3 (N7282, N7278, N2303, N6138);
xor XOR2 (N7283, N7280, N782);
buf BUF1 (N7284, N7279);
xor XOR2 (N7285, N7281, N7146);
nor NOR4 (N7286, N7284, N6507, N1073, N2476);
nand NAND4 (N7287, N7243, N4689, N2149, N5466);
not NOT1 (N7288, N7266);
nor NOR3 (N7289, N7287, N2338, N1767);
not NOT1 (N7290, N7286);
not NOT1 (N7291, N7249);
not NOT1 (N7292, N7290);
nand NAND3 (N7293, N7291, N4571, N4146);
xor XOR2 (N7294, N7292, N3393);
buf BUF1 (N7295, N7294);
nand NAND3 (N7296, N7289, N3156, N3397);
or OR2 (N7297, N7296, N3765);
nand NAND2 (N7298, N7282, N3738);
nand NAND4 (N7299, N7298, N1475, N456, N7205);
not NOT1 (N7300, N7297);
xor XOR2 (N7301, N7276, N714);
xor XOR2 (N7302, N7300, N4248);
or OR4 (N7303, N7293, N4343, N4250, N6417);
not NOT1 (N7304, N7303);
xor XOR2 (N7305, N7304, N7176);
buf BUF1 (N7306, N7285);
buf BUF1 (N7307, N7288);
nor NOR3 (N7308, N7307, N2130, N2285);
and AND2 (N7309, N7273, N1009);
and AND3 (N7310, N7268, N4261, N3862);
nor NOR3 (N7311, N7295, N2222, N4137);
nor NOR3 (N7312, N7305, N3194, N433);
or OR4 (N7313, N7302, N3427, N5965, N2098);
xor XOR2 (N7314, N7308, N6718);
and AND3 (N7315, N7312, N2496, N4359);
buf BUF1 (N7316, N7310);
buf BUF1 (N7317, N7314);
buf BUF1 (N7318, N7309);
buf BUF1 (N7319, N7283);
and AND3 (N7320, N7306, N3267, N7242);
and AND4 (N7321, N7313, N598, N5403, N5538);
buf BUF1 (N7322, N7315);
nand NAND3 (N7323, N7299, N6065, N5888);
and AND3 (N7324, N7319, N3586, N6168);
not NOT1 (N7325, N7311);
buf BUF1 (N7326, N7322);
nor NOR2 (N7327, N7324, N2882);
xor XOR2 (N7328, N7323, N6055);
nor NOR3 (N7329, N7320, N1895, N787);
nand NAND3 (N7330, N7317, N2849, N3062);
nor NOR2 (N7331, N7316, N428);
and AND3 (N7332, N7327, N3957, N200);
nor NOR4 (N7333, N7321, N4739, N5896, N4139);
nor NOR3 (N7334, N7328, N6635, N1368);
buf BUF1 (N7335, N7333);
or OR2 (N7336, N7332, N1550);
not NOT1 (N7337, N7334);
not NOT1 (N7338, N7318);
or OR4 (N7339, N7330, N6121, N5794, N4087);
not NOT1 (N7340, N7338);
xor XOR2 (N7341, N7325, N5466);
buf BUF1 (N7342, N7301);
and AND3 (N7343, N7329, N611, N4932);
xor XOR2 (N7344, N7340, N6989);
and AND4 (N7345, N7336, N2677, N4296, N5900);
nand NAND3 (N7346, N7337, N2199, N7292);
nor NOR4 (N7347, N7339, N2236, N1670, N6821);
nor NOR3 (N7348, N7345, N1602, N712);
xor XOR2 (N7349, N7346, N3484);
and AND2 (N7350, N7326, N5987);
buf BUF1 (N7351, N7335);
not NOT1 (N7352, N7347);
nand NAND4 (N7353, N7348, N8, N1436, N1119);
not NOT1 (N7354, N7331);
and AND3 (N7355, N7349, N1597, N6581);
or OR2 (N7356, N7351, N1971);
or OR4 (N7357, N7341, N7129, N673, N580);
xor XOR2 (N7358, N7353, N6767);
nand NAND3 (N7359, N7357, N6872, N3051);
or OR2 (N7360, N7344, N4827);
buf BUF1 (N7361, N7343);
not NOT1 (N7362, N7360);
buf BUF1 (N7363, N7361);
and AND4 (N7364, N7363, N34, N4120, N3510);
nor NOR4 (N7365, N7352, N5722, N7302, N227);
nand NAND2 (N7366, N7358, N7140);
buf BUF1 (N7367, N7350);
nand NAND2 (N7368, N7342, N3538);
or OR2 (N7369, N7356, N686);
buf BUF1 (N7370, N7354);
nor NOR4 (N7371, N7364, N2918, N2064, N3065);
nor NOR2 (N7372, N7369, N7129);
nand NAND4 (N7373, N7359, N7220, N6624, N3508);
buf BUF1 (N7374, N7371);
buf BUF1 (N7375, N7373);
or OR4 (N7376, N7367, N1428, N2767, N2845);
xor XOR2 (N7377, N7370, N1361);
nor NOR3 (N7378, N7365, N5355, N2669);
and AND3 (N7379, N7376, N796, N6580);
buf BUF1 (N7380, N7374);
and AND2 (N7381, N7379, N6619);
or OR4 (N7382, N7381, N6145, N6091, N4683);
not NOT1 (N7383, N7378);
nand NAND4 (N7384, N7383, N3892, N5298, N4506);
buf BUF1 (N7385, N7380);
nor NOR3 (N7386, N7366, N3865, N3342);
nand NAND3 (N7387, N7382, N2014, N3456);
not NOT1 (N7388, N7368);
or OR2 (N7389, N7372, N7178);
nor NOR3 (N7390, N7387, N3157, N3365);
not NOT1 (N7391, N7386);
buf BUF1 (N7392, N7375);
buf BUF1 (N7393, N7385);
and AND3 (N7394, N7384, N2923, N5795);
buf BUF1 (N7395, N7388);
nand NAND3 (N7396, N7391, N583, N3853);
xor XOR2 (N7397, N7377, N6727);
nor NOR4 (N7398, N7393, N830, N305, N2944);
or OR2 (N7399, N7398, N1590);
and AND4 (N7400, N7392, N1569, N3379, N738);
nand NAND3 (N7401, N7362, N7001, N2391);
buf BUF1 (N7402, N7390);
xor XOR2 (N7403, N7400, N6700);
buf BUF1 (N7404, N7401);
not NOT1 (N7405, N7395);
nand NAND4 (N7406, N7389, N239, N36, N5248);
and AND3 (N7407, N7404, N573, N353);
not NOT1 (N7408, N7402);
nor NOR3 (N7409, N7407, N2574, N4789);
xor XOR2 (N7410, N7406, N664);
nor NOR4 (N7411, N7410, N6749, N7346, N3178);
buf BUF1 (N7412, N7409);
nor NOR2 (N7413, N7397, N5035);
or OR4 (N7414, N7408, N4313, N2405, N6588);
and AND3 (N7415, N7394, N4647, N4615);
and AND4 (N7416, N7414, N554, N6422, N7405);
buf BUF1 (N7417, N5125);
xor XOR2 (N7418, N7416, N1437);
xor XOR2 (N7419, N7418, N7008);
not NOT1 (N7420, N7417);
and AND2 (N7421, N7396, N2929);
buf BUF1 (N7422, N7403);
nand NAND2 (N7423, N7420, N2257);
nor NOR2 (N7424, N7422, N5219);
buf BUF1 (N7425, N7355);
not NOT1 (N7426, N7399);
buf BUF1 (N7427, N7424);
xor XOR2 (N7428, N7419, N6986);
or OR2 (N7429, N7427, N2074);
xor XOR2 (N7430, N7423, N1766);
and AND3 (N7431, N7429, N1780, N3687);
and AND2 (N7432, N7421, N5465);
and AND4 (N7433, N7426, N5003, N6409, N2804);
not NOT1 (N7434, N7425);
and AND2 (N7435, N7412, N3945);
and AND2 (N7436, N7434, N5031);
buf BUF1 (N7437, N7415);
or OR4 (N7438, N7436, N5525, N2974, N4066);
nand NAND3 (N7439, N7431, N1138, N1776);
xor XOR2 (N7440, N7430, N160);
nor NOR4 (N7441, N7411, N667, N2993, N525);
nand NAND2 (N7442, N7433, N6998);
and AND4 (N7443, N7439, N4953, N1169, N4354);
buf BUF1 (N7444, N7438);
nor NOR4 (N7445, N7443, N6842, N2913, N371);
buf BUF1 (N7446, N7442);
buf BUF1 (N7447, N7437);
or OR2 (N7448, N7444, N3778);
nand NAND2 (N7449, N7435, N1194);
nor NOR2 (N7450, N7413, N4679);
and AND3 (N7451, N7450, N7346, N832);
not NOT1 (N7452, N7446);
nor NOR3 (N7453, N7447, N6568, N468);
nand NAND3 (N7454, N7451, N5359, N2419);
and AND4 (N7455, N7440, N1161, N1437, N3731);
not NOT1 (N7456, N7445);
not NOT1 (N7457, N7454);
xor XOR2 (N7458, N7448, N1493);
xor XOR2 (N7459, N7449, N1676);
xor XOR2 (N7460, N7441, N4929);
xor XOR2 (N7461, N7458, N4651);
and AND3 (N7462, N7452, N2907, N523);
nand NAND2 (N7463, N7459, N3470);
nor NOR2 (N7464, N7432, N57);
or OR4 (N7465, N7463, N219, N1950, N1383);
and AND4 (N7466, N7464, N253, N6163, N7188);
and AND3 (N7467, N7428, N3318, N677);
xor XOR2 (N7468, N7456, N6009);
xor XOR2 (N7469, N7461, N5632);
xor XOR2 (N7470, N7453, N5246);
not NOT1 (N7471, N7455);
or OR3 (N7472, N7468, N6558, N3223);
or OR4 (N7473, N7465, N509, N5311, N549);
or OR3 (N7474, N7470, N3441, N7173);
not NOT1 (N7475, N7469);
xor XOR2 (N7476, N7457, N1366);
xor XOR2 (N7477, N7462, N5568);
not NOT1 (N7478, N7473);
or OR3 (N7479, N7466, N2521, N6773);
nor NOR4 (N7480, N7467, N3803, N2962, N357);
buf BUF1 (N7481, N7460);
and AND4 (N7482, N7481, N2636, N4523, N277);
not NOT1 (N7483, N7475);
nand NAND2 (N7484, N7471, N3268);
nand NAND4 (N7485, N7477, N474, N3918, N2117);
or OR2 (N7486, N7483, N3738);
and AND3 (N7487, N7486, N5801, N3462);
and AND4 (N7488, N7484, N882, N4579, N4472);
xor XOR2 (N7489, N7474, N5591);
xor XOR2 (N7490, N7489, N2064);
nand NAND4 (N7491, N7488, N3723, N3127, N2600);
nor NOR4 (N7492, N7480, N614, N274, N7028);
xor XOR2 (N7493, N7491, N1692);
nor NOR3 (N7494, N7492, N2704, N3863);
nand NAND3 (N7495, N7485, N4490, N2770);
or OR4 (N7496, N7495, N2175, N5969, N732);
nor NOR3 (N7497, N7496, N3889, N5722);
nand NAND4 (N7498, N7472, N1972, N5342, N4797);
not NOT1 (N7499, N7487);
nand NAND2 (N7500, N7482, N2066);
and AND4 (N7501, N7499, N600, N4510, N1803);
and AND3 (N7502, N7494, N2503, N5539);
not NOT1 (N7503, N7502);
or OR3 (N7504, N7493, N5457, N1223);
buf BUF1 (N7505, N7479);
or OR4 (N7506, N7497, N1998, N7446, N5659);
buf BUF1 (N7507, N7504);
nand NAND2 (N7508, N7476, N1083);
or OR2 (N7509, N7508, N974);
or OR3 (N7510, N7500, N3147, N3611);
nor NOR4 (N7511, N7498, N2185, N1173, N5881);
nor NOR4 (N7512, N7509, N7385, N7031, N2687);
nor NOR3 (N7513, N7478, N3051, N3471);
nand NAND4 (N7514, N7513, N1838, N6059, N3438);
buf BUF1 (N7515, N7503);
buf BUF1 (N7516, N7505);
nand NAND2 (N7517, N7501, N4020);
xor XOR2 (N7518, N7506, N4673);
not NOT1 (N7519, N7517);
or OR3 (N7520, N7507, N5468, N4230);
xor XOR2 (N7521, N7514, N6832);
nand NAND3 (N7522, N7510, N2934, N4807);
nand NAND4 (N7523, N7522, N3558, N1323, N1462);
nor NOR4 (N7524, N7518, N1962, N6758, N5247);
or OR2 (N7525, N7520, N2163);
nand NAND4 (N7526, N7512, N1854, N2600, N105);
nand NAND2 (N7527, N7516, N846);
nor NOR3 (N7528, N7523, N6672, N4487);
nand NAND4 (N7529, N7519, N6325, N3252, N3051);
nand NAND2 (N7530, N7515, N5402);
buf BUF1 (N7531, N7526);
not NOT1 (N7532, N7530);
buf BUF1 (N7533, N7524);
nand NAND4 (N7534, N7532, N6051, N2583, N6091);
buf BUF1 (N7535, N7527);
buf BUF1 (N7536, N7531);
nand NAND4 (N7537, N7534, N5425, N478, N3526);
nor NOR3 (N7538, N7525, N4011, N201);
buf BUF1 (N7539, N7521);
nand NAND2 (N7540, N7529, N2292);
and AND4 (N7541, N7528, N3407, N7397, N6697);
xor XOR2 (N7542, N7536, N5725);
or OR2 (N7543, N7541, N5205);
buf BUF1 (N7544, N7535);
or OR3 (N7545, N7537, N1874, N1597);
not NOT1 (N7546, N7533);
not NOT1 (N7547, N7544);
and AND3 (N7548, N7539, N3079, N5343);
nand NAND3 (N7549, N7545, N4544, N3118);
nor NOR2 (N7550, N7542, N2376);
not NOT1 (N7551, N7546);
not NOT1 (N7552, N7511);
not NOT1 (N7553, N7549);
buf BUF1 (N7554, N7547);
not NOT1 (N7555, N7554);
or OR3 (N7556, N7490, N2619, N3756);
nor NOR2 (N7557, N7553, N3261);
and AND3 (N7558, N7550, N6097, N2051);
xor XOR2 (N7559, N7558, N2176);
buf BUF1 (N7560, N7559);
buf BUF1 (N7561, N7548);
buf BUF1 (N7562, N7557);
nand NAND4 (N7563, N7562, N4912, N5550, N3950);
not NOT1 (N7564, N7560);
not NOT1 (N7565, N7543);
or OR2 (N7566, N7563, N7245);
xor XOR2 (N7567, N7552, N1342);
xor XOR2 (N7568, N7538, N102);
xor XOR2 (N7569, N7565, N4755);
nand NAND4 (N7570, N7556, N4469, N3685, N4296);
or OR2 (N7571, N7570, N6178);
xor XOR2 (N7572, N7568, N3360);
xor XOR2 (N7573, N7572, N1002);
buf BUF1 (N7574, N7540);
not NOT1 (N7575, N7551);
nor NOR3 (N7576, N7567, N6277, N3403);
xor XOR2 (N7577, N7575, N6312);
or OR2 (N7578, N7571, N5395);
not NOT1 (N7579, N7574);
not NOT1 (N7580, N7577);
and AND4 (N7581, N7569, N3884, N2015, N6287);
buf BUF1 (N7582, N7581);
or OR3 (N7583, N7561, N606, N2701);
nand NAND2 (N7584, N7579, N6551);
not NOT1 (N7585, N7580);
nor NOR2 (N7586, N7576, N3410);
buf BUF1 (N7587, N7566);
and AND4 (N7588, N7587, N3561, N3699, N7245);
buf BUF1 (N7589, N7578);
nor NOR4 (N7590, N7555, N5252, N7408, N3136);
nand NAND2 (N7591, N7590, N4306);
nand NAND2 (N7592, N7591, N3);
not NOT1 (N7593, N7564);
xor XOR2 (N7594, N7573, N284);
not NOT1 (N7595, N7594);
nand NAND4 (N7596, N7595, N1441, N889, N894);
not NOT1 (N7597, N7585);
nand NAND4 (N7598, N7597, N6634, N3583, N5911);
or OR3 (N7599, N7592, N4720, N2501);
or OR2 (N7600, N7599, N3976);
or OR4 (N7601, N7600, N7306, N5578, N7274);
nand NAND4 (N7602, N7586, N5303, N5815, N7320);
or OR4 (N7603, N7602, N7264, N3589, N628);
xor XOR2 (N7604, N7584, N6307);
buf BUF1 (N7605, N7604);
or OR3 (N7606, N7582, N657, N1277);
nor NOR4 (N7607, N7606, N3965, N6883, N4160);
or OR3 (N7608, N7598, N199, N4994);
or OR3 (N7609, N7608, N4286, N150);
xor XOR2 (N7610, N7609, N2176);
or OR2 (N7611, N7593, N689);
buf BUF1 (N7612, N7605);
nand NAND2 (N7613, N7601, N50);
nand NAND2 (N7614, N7596, N989);
or OR3 (N7615, N7614, N2664, N2507);
nand NAND3 (N7616, N7613, N3601, N3938);
or OR2 (N7617, N7616, N3559);
and AND4 (N7618, N7607, N4945, N3829, N609);
and AND3 (N7619, N7589, N1822, N3523);
xor XOR2 (N7620, N7583, N1196);
or OR3 (N7621, N7612, N6258, N2801);
nand NAND3 (N7622, N7603, N7124, N5455);
and AND2 (N7623, N7610, N561);
and AND4 (N7624, N7617, N5598, N767, N2509);
nor NOR2 (N7625, N7623, N2641);
or OR4 (N7626, N7619, N721, N5859, N5907);
xor XOR2 (N7627, N7622, N1215);
and AND2 (N7628, N7615, N531);
xor XOR2 (N7629, N7621, N5076);
xor XOR2 (N7630, N7588, N5979);
nor NOR4 (N7631, N7620, N4741, N6979, N6084);
not NOT1 (N7632, N7630);
or OR2 (N7633, N7628, N2829);
and AND3 (N7634, N7611, N548, N1997);
buf BUF1 (N7635, N7625);
and AND4 (N7636, N7635, N5000, N3762, N6391);
buf BUF1 (N7637, N7626);
buf BUF1 (N7638, N7618);
xor XOR2 (N7639, N7632, N941);
xor XOR2 (N7640, N7629, N2586);
not NOT1 (N7641, N7627);
and AND3 (N7642, N7636, N2829, N4899);
or OR4 (N7643, N7637, N5032, N6117, N5913);
nor NOR3 (N7644, N7638, N3829, N992);
not NOT1 (N7645, N7624);
xor XOR2 (N7646, N7631, N7259);
not NOT1 (N7647, N7634);
nor NOR2 (N7648, N7633, N7148);
nand NAND3 (N7649, N7639, N5165, N5447);
not NOT1 (N7650, N7644);
xor XOR2 (N7651, N7648, N207);
not NOT1 (N7652, N7645);
nand NAND4 (N7653, N7652, N3335, N7184, N4765);
nor NOR4 (N7654, N7650, N1832, N1380, N2154);
xor XOR2 (N7655, N7651, N986);
and AND4 (N7656, N7641, N2675, N188, N2887);
buf BUF1 (N7657, N7654);
nor NOR4 (N7658, N7653, N1647, N4307, N6340);
or OR4 (N7659, N7656, N2271, N867, N196);
nor NOR3 (N7660, N7643, N1353, N666);
nand NAND4 (N7661, N7660, N5476, N94, N612);
or OR3 (N7662, N7646, N7596, N4336);
nand NAND4 (N7663, N7661, N384, N7657, N3521);
xor XOR2 (N7664, N1912, N5321);
buf BUF1 (N7665, N7647);
or OR3 (N7666, N7665, N7236, N5736);
or OR4 (N7667, N7655, N4081, N2596, N4531);
nand NAND2 (N7668, N7663, N6661);
nand NAND4 (N7669, N7649, N611, N7645, N4925);
not NOT1 (N7670, N7669);
and AND2 (N7671, N7670, N2702);
nor NOR3 (N7672, N7642, N7163, N7307);
nor NOR2 (N7673, N7666, N5718);
nand NAND4 (N7674, N7668, N4278, N2774, N571);
not NOT1 (N7675, N7659);
or OR2 (N7676, N7675, N7545);
nand NAND3 (N7677, N7674, N6695, N5397);
and AND4 (N7678, N7673, N2733, N6086, N5663);
and AND2 (N7679, N7678, N1767);
nor NOR4 (N7680, N7640, N7604, N5510, N2384);
buf BUF1 (N7681, N7671);
or OR3 (N7682, N7672, N3071, N7508);
and AND2 (N7683, N7667, N7430);
nor NOR3 (N7684, N7658, N6586, N3497);
xor XOR2 (N7685, N7662, N4027);
buf BUF1 (N7686, N7683);
and AND2 (N7687, N7679, N4881);
nor NOR4 (N7688, N7685, N6081, N5146, N184);
not NOT1 (N7689, N7684);
nand NAND2 (N7690, N7689, N2320);
or OR2 (N7691, N7690, N4520);
not NOT1 (N7692, N7682);
and AND3 (N7693, N7692, N1427, N6878);
nor NOR2 (N7694, N7686, N6869);
nand NAND2 (N7695, N7677, N1569);
nand NAND2 (N7696, N7694, N7216);
xor XOR2 (N7697, N7681, N3636);
nor NOR4 (N7698, N7676, N1236, N5201, N330);
nor NOR3 (N7699, N7688, N420, N4517);
nand NAND3 (N7700, N7680, N6157, N646);
and AND2 (N7701, N7696, N6693);
and AND4 (N7702, N7695, N1982, N2624, N5616);
nor NOR3 (N7703, N7699, N5686, N2133);
not NOT1 (N7704, N7700);
not NOT1 (N7705, N7697);
or OR3 (N7706, N7687, N5560, N2630);
xor XOR2 (N7707, N7706, N1095);
buf BUF1 (N7708, N7691);
or OR2 (N7709, N7704, N5254);
xor XOR2 (N7710, N7701, N4731);
and AND2 (N7711, N7702, N5226);
not NOT1 (N7712, N7698);
buf BUF1 (N7713, N7709);
xor XOR2 (N7714, N7664, N3532);
not NOT1 (N7715, N7714);
buf BUF1 (N7716, N7710);
or OR2 (N7717, N7716, N5399);
nor NOR3 (N7718, N7708, N3409, N14);
and AND3 (N7719, N7707, N84, N4764);
and AND3 (N7720, N7719, N6962, N4122);
buf BUF1 (N7721, N7718);
nor NOR3 (N7722, N7720, N5587, N7350);
xor XOR2 (N7723, N7713, N993);
nor NOR2 (N7724, N7693, N4851);
or OR2 (N7725, N7723, N4938);
buf BUF1 (N7726, N7705);
buf BUF1 (N7727, N7726);
nand NAND4 (N7728, N7727, N7349, N3249, N281);
xor XOR2 (N7729, N7725, N4943);
buf BUF1 (N7730, N7703);
and AND4 (N7731, N7724, N6194, N597, N1078);
and AND4 (N7732, N7717, N1879, N4812, N1636);
nand NAND3 (N7733, N7729, N6010, N579);
and AND2 (N7734, N7733, N4935);
or OR2 (N7735, N7722, N6533);
buf BUF1 (N7736, N7735);
and AND2 (N7737, N7728, N5465);
xor XOR2 (N7738, N7715, N3924);
nor NOR4 (N7739, N7731, N7380, N3086, N2178);
buf BUF1 (N7740, N7721);
xor XOR2 (N7741, N7711, N823);
buf BUF1 (N7742, N7734);
nor NOR4 (N7743, N7739, N2666, N1968, N3741);
or OR2 (N7744, N7732, N2657);
not NOT1 (N7745, N7712);
and AND4 (N7746, N7743, N3067, N3583, N3131);
nor NOR2 (N7747, N7740, N34);
nor NOR4 (N7748, N7741, N1762, N6180, N4690);
nor NOR4 (N7749, N7737, N6840, N5476, N1571);
nand NAND3 (N7750, N7742, N6362, N5451);
nor NOR3 (N7751, N7748, N5538, N1630);
nand NAND2 (N7752, N7744, N2213);
nand NAND3 (N7753, N7747, N3948, N5232);
nand NAND4 (N7754, N7752, N1695, N809, N4594);
or OR3 (N7755, N7749, N5444, N4325);
nor NOR3 (N7756, N7754, N4110, N4696);
xor XOR2 (N7757, N7746, N2665);
not NOT1 (N7758, N7750);
xor XOR2 (N7759, N7730, N5585);
or OR2 (N7760, N7759, N3600);
nand NAND4 (N7761, N7736, N1210, N2548, N5265);
xor XOR2 (N7762, N7761, N1292);
nor NOR2 (N7763, N7762, N6662);
nor NOR3 (N7764, N7751, N105, N1993);
xor XOR2 (N7765, N7755, N6528);
buf BUF1 (N7766, N7760);
or OR2 (N7767, N7758, N4916);
nor NOR4 (N7768, N7738, N6348, N2519, N3902);
nor NOR3 (N7769, N7768, N4066, N1467);
and AND3 (N7770, N7763, N7748, N1214);
buf BUF1 (N7771, N7753);
and AND4 (N7772, N7770, N774, N153, N552);
nor NOR4 (N7773, N7772, N674, N974, N4509);
not NOT1 (N7774, N7767);
not NOT1 (N7775, N7766);
buf BUF1 (N7776, N7775);
xor XOR2 (N7777, N7757, N7004);
buf BUF1 (N7778, N7764);
not NOT1 (N7779, N7745);
and AND3 (N7780, N7773, N3749, N3313);
or OR4 (N7781, N7780, N679, N3026, N2796);
buf BUF1 (N7782, N7779);
buf BUF1 (N7783, N7756);
or OR3 (N7784, N7777, N4721, N2432);
and AND3 (N7785, N7769, N221, N702);
buf BUF1 (N7786, N7778);
nand NAND4 (N7787, N7782, N4357, N1111, N1416);
or OR3 (N7788, N7785, N2095, N1256);
buf BUF1 (N7789, N7781);
not NOT1 (N7790, N7788);
and AND3 (N7791, N7765, N2403, N5584);
nor NOR2 (N7792, N7776, N6963);
nor NOR4 (N7793, N7783, N3751, N6606, N2866);
or OR2 (N7794, N7789, N223);
or OR2 (N7795, N7771, N6499);
nor NOR2 (N7796, N7784, N6807);
not NOT1 (N7797, N7795);
nor NOR3 (N7798, N7792, N1603, N4289);
not NOT1 (N7799, N7791);
and AND2 (N7800, N7798, N6368);
or OR3 (N7801, N7787, N6609, N363);
nor NOR3 (N7802, N7794, N4105, N2573);
buf BUF1 (N7803, N7790);
and AND4 (N7804, N7796, N7154, N3172, N3311);
nor NOR4 (N7805, N7793, N4670, N3751, N1172);
buf BUF1 (N7806, N7804);
or OR4 (N7807, N7801, N621, N4329, N4257);
or OR4 (N7808, N7799, N6537, N1882, N5945);
nor NOR4 (N7809, N7803, N3649, N7267, N7573);
and AND4 (N7810, N7805, N4745, N5655, N5060);
or OR3 (N7811, N7806, N5897, N5324);
nand NAND3 (N7812, N7811, N6307, N543);
nand NAND4 (N7813, N7802, N730, N3110, N6700);
not NOT1 (N7814, N7807);
nand NAND3 (N7815, N7786, N6929, N4564);
buf BUF1 (N7816, N7812);
buf BUF1 (N7817, N7809);
and AND2 (N7818, N7815, N889);
xor XOR2 (N7819, N7814, N4012);
and AND3 (N7820, N7810, N6748, N7110);
xor XOR2 (N7821, N7819, N4436);
and AND2 (N7822, N7818, N7354);
and AND3 (N7823, N7813, N887, N2528);
nand NAND4 (N7824, N7823, N3322, N7052, N2508);
not NOT1 (N7825, N7824);
buf BUF1 (N7826, N7774);
nor NOR2 (N7827, N7821, N4666);
or OR2 (N7828, N7816, N7370);
nor NOR4 (N7829, N7808, N3058, N6936, N879);
buf BUF1 (N7830, N7829);
nor NOR3 (N7831, N7822, N5734, N2758);
not NOT1 (N7832, N7830);
and AND4 (N7833, N7820, N6757, N2135, N5247);
or OR2 (N7834, N7825, N852);
buf BUF1 (N7835, N7834);
not NOT1 (N7836, N7827);
and AND2 (N7837, N7800, N6560);
xor XOR2 (N7838, N7817, N7327);
not NOT1 (N7839, N7837);
nor NOR2 (N7840, N7836, N1034);
not NOT1 (N7841, N7831);
and AND2 (N7842, N7833, N1782);
or OR3 (N7843, N7839, N5567, N6547);
and AND4 (N7844, N7842, N4303, N7191, N1440);
xor XOR2 (N7845, N7832, N6308);
nand NAND2 (N7846, N7835, N350);
nor NOR2 (N7847, N7845, N5408);
xor XOR2 (N7848, N7840, N1862);
nand NAND2 (N7849, N7843, N7307);
nor NOR4 (N7850, N7847, N6865, N1643, N7782);
not NOT1 (N7851, N7841);
xor XOR2 (N7852, N7851, N2828);
or OR2 (N7853, N7849, N417);
nor NOR2 (N7854, N7844, N5388);
and AND2 (N7855, N7846, N2623);
nand NAND3 (N7856, N7826, N2497, N515);
not NOT1 (N7857, N7797);
and AND3 (N7858, N7850, N6315, N807);
or OR4 (N7859, N7858, N2141, N2243, N6290);
not NOT1 (N7860, N7852);
and AND2 (N7861, N7860, N6684);
not NOT1 (N7862, N7838);
and AND2 (N7863, N7857, N1526);
and AND2 (N7864, N7853, N5831);
xor XOR2 (N7865, N7848, N7694);
xor XOR2 (N7866, N7855, N6140);
nor NOR3 (N7867, N7859, N650, N7079);
nor NOR3 (N7868, N7867, N4476, N1182);
not NOT1 (N7869, N7862);
not NOT1 (N7870, N7864);
or OR4 (N7871, N7868, N3016, N2313, N880);
xor XOR2 (N7872, N7866, N5191);
buf BUF1 (N7873, N7869);
nor NOR4 (N7874, N7828, N2598, N1614, N7098);
not NOT1 (N7875, N7871);
or OR2 (N7876, N7863, N976);
and AND2 (N7877, N7854, N277);
xor XOR2 (N7878, N7856, N7039);
nor NOR4 (N7879, N7870, N2209, N4033, N5971);
buf BUF1 (N7880, N7874);
buf BUF1 (N7881, N7879);
and AND4 (N7882, N7880, N2339, N3262, N7869);
buf BUF1 (N7883, N7872);
or OR3 (N7884, N7882, N242, N627);
buf BUF1 (N7885, N7876);
buf BUF1 (N7886, N7878);
and AND2 (N7887, N7884, N289);
nor NOR4 (N7888, N7875, N1988, N3899, N4617);
and AND2 (N7889, N7877, N4994);
nand NAND2 (N7890, N7888, N4716);
nor NOR2 (N7891, N7887, N7331);
nor NOR3 (N7892, N7890, N1632, N5100);
not NOT1 (N7893, N7886);
buf BUF1 (N7894, N7892);
xor XOR2 (N7895, N7881, N3456);
not NOT1 (N7896, N7885);
or OR3 (N7897, N7865, N6597, N7312);
nand NAND2 (N7898, N7895, N3578);
and AND2 (N7899, N7896, N657);
or OR3 (N7900, N7893, N2506, N6308);
xor XOR2 (N7901, N7898, N6010);
or OR2 (N7902, N7873, N5005);
buf BUF1 (N7903, N7861);
nand NAND4 (N7904, N7901, N1900, N2666, N2026);
buf BUF1 (N7905, N7883);
or OR2 (N7906, N7894, N2962);
buf BUF1 (N7907, N7899);
buf BUF1 (N7908, N7902);
nor NOR3 (N7909, N7891, N6345, N4543);
buf BUF1 (N7910, N7903);
nand NAND2 (N7911, N7897, N1401);
buf BUF1 (N7912, N7911);
not NOT1 (N7913, N7910);
not NOT1 (N7914, N7909);
nor NOR4 (N7915, N7912, N6929, N5569, N3488);
not NOT1 (N7916, N7914);
nand NAND3 (N7917, N7913, N7791, N4028);
and AND3 (N7918, N7906, N2356, N6308);
not NOT1 (N7919, N7918);
xor XOR2 (N7920, N7908, N1098);
nor NOR2 (N7921, N7904, N5145);
nand NAND3 (N7922, N7907, N4391, N3362);
or OR2 (N7923, N7905, N6905);
buf BUF1 (N7924, N7922);
and AND4 (N7925, N7917, N613, N5385, N7785);
nor NOR4 (N7926, N7900, N5519, N4160, N6568);
and AND2 (N7927, N7889, N4066);
or OR4 (N7928, N7920, N1172, N2257, N6029);
xor XOR2 (N7929, N7915, N235);
buf BUF1 (N7930, N7929);
xor XOR2 (N7931, N7926, N5800);
or OR3 (N7932, N7930, N105, N1156);
buf BUF1 (N7933, N7932);
buf BUF1 (N7934, N7923);
or OR3 (N7935, N7928, N1018, N2561);
nor NOR4 (N7936, N7934, N4849, N406, N7129);
not NOT1 (N7937, N7935);
and AND4 (N7938, N7933, N3013, N1604, N325);
nand NAND3 (N7939, N7921, N3371, N5646);
and AND3 (N7940, N7925, N6240, N4727);
nor NOR4 (N7941, N7924, N4346, N7309, N5827);
not NOT1 (N7942, N7939);
buf BUF1 (N7943, N7938);
not NOT1 (N7944, N7943);
not NOT1 (N7945, N7916);
and AND4 (N7946, N7937, N1475, N2480, N5271);
nor NOR3 (N7947, N7945, N5993, N5293);
or OR2 (N7948, N7946, N7170);
xor XOR2 (N7949, N7936, N897);
and AND3 (N7950, N7948, N6471, N5074);
nor NOR4 (N7951, N7941, N2846, N5883, N4785);
and AND3 (N7952, N7950, N4396, N1128);
or OR3 (N7953, N7947, N5080, N3552);
buf BUF1 (N7954, N7951);
nor NOR2 (N7955, N7942, N7279);
nand NAND2 (N7956, N7949, N438);
nor NOR4 (N7957, N7919, N281, N2326, N3502);
buf BUF1 (N7958, N7955);
or OR4 (N7959, N7927, N4933, N3061, N5418);
buf BUF1 (N7960, N7953);
or OR2 (N7961, N7957, N4554);
or OR2 (N7962, N7952, N7800);
nor NOR2 (N7963, N7956, N6964);
xor XOR2 (N7964, N7940, N1661);
or OR2 (N7965, N7958, N3404);
xor XOR2 (N7966, N7962, N1164);
nand NAND3 (N7967, N7965, N353, N712);
or OR3 (N7968, N7954, N2423, N930);
nor NOR2 (N7969, N7960, N674);
buf BUF1 (N7970, N7969);
or OR3 (N7971, N7967, N3985, N7754);
or OR3 (N7972, N7931, N4066, N6407);
xor XOR2 (N7973, N7964, N162);
or OR4 (N7974, N7966, N7298, N2505, N7356);
nand NAND4 (N7975, N7970, N4884, N646, N643);
and AND3 (N7976, N7944, N4240, N5702);
buf BUF1 (N7977, N7968);
not NOT1 (N7978, N7977);
not NOT1 (N7979, N7959);
buf BUF1 (N7980, N7971);
xor XOR2 (N7981, N7974, N2551);
or OR2 (N7982, N7980, N7796);
or OR4 (N7983, N7961, N1809, N3709, N1818);
not NOT1 (N7984, N7978);
not NOT1 (N7985, N7983);
buf BUF1 (N7986, N7973);
or OR3 (N7987, N7984, N1189, N4253);
buf BUF1 (N7988, N7987);
not NOT1 (N7989, N7963);
nor NOR4 (N7990, N7975, N1874, N4592, N7053);
xor XOR2 (N7991, N7988, N7022);
and AND4 (N7992, N7990, N7873, N349, N4332);
and AND3 (N7993, N7991, N5732, N6214);
not NOT1 (N7994, N7986);
buf BUF1 (N7995, N7981);
xor XOR2 (N7996, N7972, N6087);
nand NAND4 (N7997, N7995, N1415, N6837, N7744);
xor XOR2 (N7998, N7976, N5027);
and AND4 (N7999, N7996, N6775, N5865, N4687);
and AND3 (N8000, N7999, N2030, N6783);
xor XOR2 (N8001, N7992, N660);
xor XOR2 (N8002, N7979, N6415);
nand NAND3 (N8003, N7997, N2543, N5701);
nand NAND4 (N8004, N8003, N3572, N4012, N5687);
buf BUF1 (N8005, N8002);
nor NOR2 (N8006, N7989, N7434);
buf BUF1 (N8007, N8006);
nor NOR4 (N8008, N8000, N1741, N5266, N7255);
buf BUF1 (N8009, N7982);
xor XOR2 (N8010, N7994, N5498);
not NOT1 (N8011, N7993);
xor XOR2 (N8012, N8008, N7268);
buf BUF1 (N8013, N8001);
not NOT1 (N8014, N8007);
and AND2 (N8015, N8011, N805);
xor XOR2 (N8016, N8005, N5470);
and AND2 (N8017, N8004, N1812);
xor XOR2 (N8018, N8010, N4161);
nor NOR3 (N8019, N8014, N3875, N2653);
xor XOR2 (N8020, N8017, N1005);
buf BUF1 (N8021, N8009);
or OR4 (N8022, N8012, N7460, N2767, N5295);
nor NOR4 (N8023, N8019, N6319, N7155, N692);
xor XOR2 (N8024, N8020, N3495);
xor XOR2 (N8025, N7998, N1470);
nand NAND3 (N8026, N8023, N610, N781);
or OR2 (N8027, N8026, N2927);
xor XOR2 (N8028, N8024, N3485);
xor XOR2 (N8029, N8021, N1365);
nand NAND2 (N8030, N8013, N3857);
buf BUF1 (N8031, N8022);
and AND3 (N8032, N8018, N4945, N3078);
buf BUF1 (N8033, N8032);
not NOT1 (N8034, N8033);
xor XOR2 (N8035, N8016, N3590);
and AND2 (N8036, N8025, N4545);
xor XOR2 (N8037, N8029, N4005);
or OR3 (N8038, N8036, N4493, N1706);
not NOT1 (N8039, N8031);
buf BUF1 (N8040, N8030);
nand NAND3 (N8041, N8028, N104, N4871);
or OR4 (N8042, N8027, N7728, N7350, N1285);
not NOT1 (N8043, N8015);
not NOT1 (N8044, N8042);
nor NOR3 (N8045, N8037, N3353, N547);
buf BUF1 (N8046, N7985);
buf BUF1 (N8047, N8035);
and AND4 (N8048, N8039, N7281, N2127, N4148);
buf BUF1 (N8049, N8043);
not NOT1 (N8050, N8047);
nand NAND2 (N8051, N8049, N2179);
nand NAND2 (N8052, N8034, N4470);
not NOT1 (N8053, N8046);
not NOT1 (N8054, N8044);
or OR4 (N8055, N8048, N5210, N2621, N7090);
and AND3 (N8056, N8053, N4060, N6364);
xor XOR2 (N8057, N8056, N4823);
or OR4 (N8058, N8051, N6738, N1609, N891);
nor NOR2 (N8059, N8038, N548);
and AND4 (N8060, N8052, N3454, N3278, N5179);
nand NAND3 (N8061, N8054, N6544, N6926);
and AND3 (N8062, N8050, N202, N5568);
nor NOR4 (N8063, N8061, N3344, N4339, N952);
not NOT1 (N8064, N8045);
buf BUF1 (N8065, N8040);
nand NAND2 (N8066, N8055, N6638);
not NOT1 (N8067, N8059);
not NOT1 (N8068, N8064);
nor NOR2 (N8069, N8060, N3397);
and AND4 (N8070, N8067, N2104, N6164, N5304);
not NOT1 (N8071, N8069);
and AND2 (N8072, N8062, N6841);
nand NAND2 (N8073, N8072, N1538);
buf BUF1 (N8074, N8073);
buf BUF1 (N8075, N8071);
nor NOR3 (N8076, N8070, N2996, N8034);
buf BUF1 (N8077, N8068);
or OR4 (N8078, N8065, N5732, N6158, N2048);
nor NOR4 (N8079, N8057, N648, N6259, N6712);
nor NOR3 (N8080, N8077, N975, N1110);
buf BUF1 (N8081, N8075);
and AND3 (N8082, N8066, N3162, N3106);
xor XOR2 (N8083, N8078, N7241);
nor NOR2 (N8084, N8081, N4379);
and AND4 (N8085, N8041, N717, N1696, N5541);
nor NOR3 (N8086, N8074, N2931, N1001);
or OR3 (N8087, N8082, N7054, N5075);
or OR4 (N8088, N8080, N1081, N4980, N1418);
and AND2 (N8089, N8058, N3873);
or OR4 (N8090, N8087, N2040, N871, N7803);
nor NOR2 (N8091, N8063, N3916);
or OR4 (N8092, N8089, N7542, N2001, N1337);
buf BUF1 (N8093, N8091);
nand NAND3 (N8094, N8088, N4392, N2168);
and AND2 (N8095, N8085, N3251);
and AND4 (N8096, N8084, N4887, N5059, N6421);
and AND3 (N8097, N8093, N4434, N8006);
not NOT1 (N8098, N8097);
buf BUF1 (N8099, N8090);
buf BUF1 (N8100, N8076);
or OR4 (N8101, N8094, N2773, N7838, N3018);
xor XOR2 (N8102, N8101, N1583);
buf BUF1 (N8103, N8092);
not NOT1 (N8104, N8102);
buf BUF1 (N8105, N8103);
xor XOR2 (N8106, N8083, N972);
buf BUF1 (N8107, N8100);
nand NAND4 (N8108, N8086, N4201, N7967, N1088);
buf BUF1 (N8109, N8108);
buf BUF1 (N8110, N8079);
buf BUF1 (N8111, N8107);
and AND4 (N8112, N8111, N5944, N2275, N530);
not NOT1 (N8113, N8095);
or OR2 (N8114, N8104, N7265);
nor NOR3 (N8115, N8106, N7823, N475);
or OR4 (N8116, N8113, N6969, N596, N3039);
not NOT1 (N8117, N8114);
buf BUF1 (N8118, N8105);
or OR4 (N8119, N8099, N5258, N5438, N2410);
buf BUF1 (N8120, N8109);
or OR4 (N8121, N8112, N5576, N5209, N2640);
nor NOR3 (N8122, N8119, N7591, N1431);
not NOT1 (N8123, N8121);
xor XOR2 (N8124, N8115, N843);
nand NAND4 (N8125, N8124, N3996, N622, N5582);
xor XOR2 (N8126, N8125, N7396);
nor NOR4 (N8127, N8110, N4098, N2043, N2730);
nand NAND4 (N8128, N8123, N6880, N6625, N4969);
nand NAND2 (N8129, N8128, N6392);
buf BUF1 (N8130, N8116);
or OR4 (N8131, N8129, N1414, N99, N3907);
nand NAND3 (N8132, N8127, N5232, N736);
not NOT1 (N8133, N8131);
not NOT1 (N8134, N8133);
and AND2 (N8135, N8134, N3283);
xor XOR2 (N8136, N8132, N6190);
not NOT1 (N8137, N8096);
nand NAND2 (N8138, N8136, N7246);
xor XOR2 (N8139, N8130, N2947);
nor NOR2 (N8140, N8118, N5642);
or OR2 (N8141, N8126, N2943);
and AND2 (N8142, N8122, N6474);
nand NAND4 (N8143, N8098, N3765, N3094, N5950);
or OR3 (N8144, N8137, N4191, N2045);
xor XOR2 (N8145, N8142, N7167);
not NOT1 (N8146, N8138);
xor XOR2 (N8147, N8140, N2950);
and AND4 (N8148, N8147, N5000, N2859, N482);
nand NAND2 (N8149, N8117, N6152);
or OR3 (N8150, N8135, N2586, N3268);
xor XOR2 (N8151, N8150, N7752);
and AND2 (N8152, N8151, N4013);
buf BUF1 (N8153, N8120);
or OR4 (N8154, N8145, N1806, N7357, N3656);
or OR4 (N8155, N8148, N2637, N5814, N3115);
xor XOR2 (N8156, N8141, N1814);
buf BUF1 (N8157, N8154);
or OR3 (N8158, N8139, N266, N3421);
and AND4 (N8159, N8149, N7896, N5353, N2948);
buf BUF1 (N8160, N8159);
nand NAND4 (N8161, N8146, N6414, N1942, N1876);
not NOT1 (N8162, N8152);
xor XOR2 (N8163, N8144, N8077);
not NOT1 (N8164, N8157);
buf BUF1 (N8165, N8155);
buf BUF1 (N8166, N8143);
buf BUF1 (N8167, N8162);
xor XOR2 (N8168, N8160, N3023);
or OR2 (N8169, N8168, N2925);
xor XOR2 (N8170, N8169, N1644);
nor NOR2 (N8171, N8170, N4381);
nand NAND2 (N8172, N8164, N7301);
xor XOR2 (N8173, N8161, N4334);
xor XOR2 (N8174, N8163, N7764);
not NOT1 (N8175, N8153);
xor XOR2 (N8176, N8166, N1108);
xor XOR2 (N8177, N8174, N7571);
nor NOR4 (N8178, N8175, N3095, N5046, N3486);
not NOT1 (N8179, N8176);
or OR4 (N8180, N8156, N1266, N6221, N5161);
xor XOR2 (N8181, N8171, N6639);
not NOT1 (N8182, N8167);
and AND4 (N8183, N8179, N4811, N318, N2608);
not NOT1 (N8184, N8180);
not NOT1 (N8185, N8183);
not NOT1 (N8186, N8172);
and AND4 (N8187, N8182, N600, N133, N3769);
nand NAND2 (N8188, N8187, N4103);
buf BUF1 (N8189, N8184);
nor NOR2 (N8190, N8173, N7933);
and AND3 (N8191, N8178, N1470, N6496);
xor XOR2 (N8192, N8181, N2331);
or OR4 (N8193, N8186, N766, N4059, N7711);
buf BUF1 (N8194, N8188);
not NOT1 (N8195, N8165);
nand NAND3 (N8196, N8195, N719, N7474);
buf BUF1 (N8197, N8189);
buf BUF1 (N8198, N8177);
nor NOR4 (N8199, N8198, N7958, N212, N5591);
or OR3 (N8200, N8190, N3865, N3425);
nor NOR3 (N8201, N8199, N686, N1424);
nand NAND4 (N8202, N8201, N2606, N6895, N7435);
buf BUF1 (N8203, N8158);
nand NAND2 (N8204, N8193, N5804);
xor XOR2 (N8205, N8196, N1072);
nor NOR3 (N8206, N8185, N3272, N3634);
and AND4 (N8207, N8191, N4249, N1398, N1670);
nand NAND4 (N8208, N8197, N7055, N6012, N7855);
or OR3 (N8209, N8192, N1795, N4634);
xor XOR2 (N8210, N8204, N2304);
or OR4 (N8211, N8194, N1341, N2401, N7444);
nor NOR3 (N8212, N8209, N3643, N2696);
xor XOR2 (N8213, N8203, N5325);
nand NAND4 (N8214, N8211, N3597, N5193, N2958);
nor NOR2 (N8215, N8208, N3048);
or OR2 (N8216, N8213, N5269);
nand NAND4 (N8217, N8210, N1488, N1598, N6497);
nor NOR4 (N8218, N8215, N321, N3853, N3097);
or OR3 (N8219, N8207, N7797, N7200);
and AND3 (N8220, N8212, N7047, N3060);
and AND2 (N8221, N8216, N4293);
buf BUF1 (N8222, N8200);
buf BUF1 (N8223, N8206);
or OR4 (N8224, N8205, N2356, N3643, N7681);
or OR2 (N8225, N8219, N7582);
and AND3 (N8226, N8217, N1002, N5366);
nand NAND2 (N8227, N8224, N6603);
nand NAND4 (N8228, N8218, N7629, N5780, N7787);
not NOT1 (N8229, N8225);
not NOT1 (N8230, N8220);
nand NAND2 (N8231, N8221, N2448);
nand NAND2 (N8232, N8230, N2957);
not NOT1 (N8233, N8214);
or OR4 (N8234, N8223, N1857, N6487, N3449);
and AND3 (N8235, N8227, N1172, N692);
nand NAND4 (N8236, N8226, N3505, N4195, N8159);
or OR3 (N8237, N8232, N6665, N5633);
and AND2 (N8238, N8237, N2606);
nand NAND4 (N8239, N8229, N7655, N2550, N3578);
not NOT1 (N8240, N8222);
or OR3 (N8241, N8238, N4520, N4269);
nand NAND3 (N8242, N8202, N8198, N481);
nand NAND3 (N8243, N8233, N2984, N3790);
buf BUF1 (N8244, N8239);
buf BUF1 (N8245, N8234);
xor XOR2 (N8246, N8243, N7806);
buf BUF1 (N8247, N8241);
nor NOR2 (N8248, N8235, N4257);
xor XOR2 (N8249, N8242, N2433);
xor XOR2 (N8250, N8248, N152);
not NOT1 (N8251, N8240);
nor NOR4 (N8252, N8244, N4556, N2744, N6105);
not NOT1 (N8253, N8245);
and AND2 (N8254, N8247, N7086);
not NOT1 (N8255, N8246);
or OR3 (N8256, N8250, N7833, N3757);
buf BUF1 (N8257, N8256);
buf BUF1 (N8258, N8254);
xor XOR2 (N8259, N8255, N1107);
not NOT1 (N8260, N8249);
and AND3 (N8261, N8258, N4954, N1974);
not NOT1 (N8262, N8252);
xor XOR2 (N8263, N8262, N5270);
and AND4 (N8264, N8231, N7266, N1814, N83);
nand NAND4 (N8265, N8259, N7491, N13, N5386);
nor NOR4 (N8266, N8253, N6575, N1859, N7041);
and AND4 (N8267, N8263, N8205, N4818, N4068);
nand NAND4 (N8268, N8261, N3687, N1127, N513);
or OR2 (N8269, N8228, N3088);
nor NOR4 (N8270, N8266, N7227, N5270, N7722);
buf BUF1 (N8271, N8264);
nand NAND2 (N8272, N8268, N2578);
not NOT1 (N8273, N8271);
nor NOR3 (N8274, N8270, N1913, N880);
and AND2 (N8275, N8274, N971);
not NOT1 (N8276, N8251);
buf BUF1 (N8277, N8260);
xor XOR2 (N8278, N8236, N4833);
buf BUF1 (N8279, N8267);
not NOT1 (N8280, N8273);
or OR3 (N8281, N8280, N2809, N6592);
and AND2 (N8282, N8276, N3850);
buf BUF1 (N8283, N8279);
xor XOR2 (N8284, N8277, N6140);
and AND3 (N8285, N8269, N3601, N7438);
or OR2 (N8286, N8283, N7566);
nor NOR3 (N8287, N8281, N4746, N4754);
xor XOR2 (N8288, N8278, N5401);
and AND2 (N8289, N8272, N210);
buf BUF1 (N8290, N8287);
nor NOR4 (N8291, N8286, N1572, N8011, N1897);
xor XOR2 (N8292, N8290, N4220);
not NOT1 (N8293, N8275);
or OR3 (N8294, N8282, N8185, N3009);
buf BUF1 (N8295, N8294);
nand NAND4 (N8296, N8293, N808, N1124, N568);
not NOT1 (N8297, N8257);
nor NOR4 (N8298, N8289, N5931, N6858, N5629);
and AND2 (N8299, N8295, N2646);
xor XOR2 (N8300, N8299, N1275);
nand NAND3 (N8301, N8292, N1553, N7633);
buf BUF1 (N8302, N8291);
and AND4 (N8303, N8284, N5928, N6687, N7330);
nand NAND4 (N8304, N8301, N2240, N8135, N2829);
nor NOR3 (N8305, N8300, N4814, N4408);
buf BUF1 (N8306, N8285);
nand NAND2 (N8307, N8297, N433);
nor NOR2 (N8308, N8307, N1868);
nand NAND3 (N8309, N8288, N6917, N6232);
buf BUF1 (N8310, N8296);
buf BUF1 (N8311, N8309);
buf BUF1 (N8312, N8265);
buf BUF1 (N8313, N8303);
or OR2 (N8314, N8306, N2462);
nor NOR2 (N8315, N8310, N2331);
xor XOR2 (N8316, N8302, N3596);
nand NAND3 (N8317, N8312, N6198, N964);
not NOT1 (N8318, N8313);
and AND3 (N8319, N8308, N593, N6592);
not NOT1 (N8320, N8319);
nand NAND2 (N8321, N8316, N440);
nand NAND4 (N8322, N8305, N5207, N2216, N6602);
or OR4 (N8323, N8298, N7117, N6575, N46);
nand NAND3 (N8324, N8314, N6246, N8045);
and AND3 (N8325, N8315, N7873, N96);
nand NAND4 (N8326, N8324, N2582, N4632, N1103);
not NOT1 (N8327, N8323);
and AND2 (N8328, N8318, N2187);
nand NAND3 (N8329, N8322, N6571, N3256);
and AND4 (N8330, N8325, N5929, N6380, N1112);
or OR3 (N8331, N8317, N4324, N2441);
xor XOR2 (N8332, N8321, N4797);
xor XOR2 (N8333, N8328, N5703);
and AND4 (N8334, N8332, N6770, N4950, N1899);
or OR4 (N8335, N8334, N5726, N247, N7424);
buf BUF1 (N8336, N8326);
and AND2 (N8337, N8327, N4321);
xor XOR2 (N8338, N8311, N1231);
nand NAND3 (N8339, N8335, N809, N3086);
not NOT1 (N8340, N8331);
or OR4 (N8341, N8333, N1536, N2074, N148);
or OR3 (N8342, N8339, N5599, N5848);
buf BUF1 (N8343, N8320);
buf BUF1 (N8344, N8340);
or OR3 (N8345, N8336, N4354, N5978);
nor NOR4 (N8346, N8345, N4064, N2645, N6261);
nand NAND3 (N8347, N8329, N4495, N3255);
nor NOR4 (N8348, N8342, N5398, N6789, N7111);
buf BUF1 (N8349, N8348);
and AND3 (N8350, N8341, N6058, N1373);
buf BUF1 (N8351, N8350);
buf BUF1 (N8352, N8349);
nor NOR2 (N8353, N8304, N4260);
not NOT1 (N8354, N8353);
nand NAND3 (N8355, N8344, N6128, N378);
nor NOR3 (N8356, N8347, N4572, N7072);
or OR4 (N8357, N8354, N3059, N3828, N1236);
not NOT1 (N8358, N8346);
not NOT1 (N8359, N8343);
nand NAND2 (N8360, N8338, N6389);
nor NOR4 (N8361, N8351, N282, N3586, N3570);
and AND4 (N8362, N8330, N6299, N4708, N2049);
nand NAND4 (N8363, N8362, N2621, N2911, N6191);
xor XOR2 (N8364, N8359, N7189);
and AND2 (N8365, N8357, N998);
not NOT1 (N8366, N8358);
and AND2 (N8367, N8356, N2537);
or OR4 (N8368, N8352, N1888, N2081, N3925);
xor XOR2 (N8369, N8368, N2896);
not NOT1 (N8370, N8361);
xor XOR2 (N8371, N8363, N2018);
nor NOR4 (N8372, N8366, N2407, N4985, N166);
xor XOR2 (N8373, N8367, N7469);
and AND4 (N8374, N8337, N6363, N6802, N3817);
and AND3 (N8375, N8365, N5103, N2539);
and AND3 (N8376, N8370, N8309, N2926);
xor XOR2 (N8377, N8372, N6579);
nand NAND3 (N8378, N8369, N1544, N7375);
nor NOR4 (N8379, N8364, N5730, N2398, N3301);
buf BUF1 (N8380, N8374);
nor NOR3 (N8381, N8380, N3704, N1551);
buf BUF1 (N8382, N8371);
and AND2 (N8383, N8355, N7757);
not NOT1 (N8384, N8383);
or OR3 (N8385, N8384, N6909, N1856);
not NOT1 (N8386, N8378);
xor XOR2 (N8387, N8379, N227);
nor NOR2 (N8388, N8377, N341);
and AND4 (N8389, N8382, N8103, N5402, N5714);
and AND3 (N8390, N8376, N3, N2083);
nand NAND2 (N8391, N8385, N6251);
buf BUF1 (N8392, N8375);
xor XOR2 (N8393, N8373, N8134);
and AND4 (N8394, N8389, N594, N5541, N1467);
buf BUF1 (N8395, N8381);
nor NOR3 (N8396, N8387, N8260, N4227);
nand NAND2 (N8397, N8386, N7634);
nand NAND2 (N8398, N8393, N2759);
nor NOR2 (N8399, N8390, N6422);
not NOT1 (N8400, N8391);
not NOT1 (N8401, N8396);
not NOT1 (N8402, N8397);
nand NAND4 (N8403, N8388, N576, N5177, N4235);
buf BUF1 (N8404, N8403);
nand NAND2 (N8405, N8400, N5991);
or OR3 (N8406, N8394, N3069, N4371);
nor NOR2 (N8407, N8399, N6341);
and AND2 (N8408, N8406, N2163);
not NOT1 (N8409, N8360);
and AND3 (N8410, N8404, N3349, N2489);
not NOT1 (N8411, N8392);
nor NOR3 (N8412, N8402, N5986, N4893);
xor XOR2 (N8413, N8395, N2468);
and AND4 (N8414, N8410, N3231, N4023, N159);
and AND2 (N8415, N8414, N6538);
and AND4 (N8416, N8415, N5623, N8367, N107);
nor NOR4 (N8417, N8405, N6588, N5826, N2478);
nor NOR2 (N8418, N8398, N2540);
nor NOR4 (N8419, N8418, N2626, N5087, N6030);
nor NOR3 (N8420, N8408, N4331, N4281);
xor XOR2 (N8421, N8420, N5410);
not NOT1 (N8422, N8421);
nand NAND2 (N8423, N8419, N3058);
nor NOR2 (N8424, N8417, N2948);
or OR4 (N8425, N8416, N5610, N7246, N7973);
xor XOR2 (N8426, N8407, N4774);
nor NOR4 (N8427, N8424, N2850, N2363, N5780);
buf BUF1 (N8428, N8401);
not NOT1 (N8429, N8413);
or OR4 (N8430, N8426, N3117, N3739, N3796);
not NOT1 (N8431, N8412);
buf BUF1 (N8432, N8427);
nor NOR2 (N8433, N8411, N14);
nand NAND3 (N8434, N8433, N2449, N2751);
and AND3 (N8435, N8434, N2820, N5282);
or OR3 (N8436, N8423, N5998, N528);
nand NAND2 (N8437, N8409, N2283);
buf BUF1 (N8438, N8436);
nor NOR4 (N8439, N8435, N5558, N1654, N4699);
not NOT1 (N8440, N8425);
nand NAND4 (N8441, N8437, N1045, N2149, N4690);
nor NOR2 (N8442, N8439, N5422);
or OR3 (N8443, N8429, N6466, N5672);
nand NAND3 (N8444, N8430, N4550, N472);
and AND3 (N8445, N8438, N6433, N4519);
not NOT1 (N8446, N8443);
not NOT1 (N8447, N8442);
nand NAND4 (N8448, N8431, N3984, N7161, N3427);
not NOT1 (N8449, N8447);
or OR3 (N8450, N8444, N794, N2964);
not NOT1 (N8451, N8448);
not NOT1 (N8452, N8451);
xor XOR2 (N8453, N8422, N923);
or OR2 (N8454, N8432, N6967);
nand NAND4 (N8455, N8453, N7647, N6127, N467);
xor XOR2 (N8456, N8450, N4472);
and AND3 (N8457, N8441, N3062, N5719);
nand NAND2 (N8458, N8457, N2718);
nand NAND2 (N8459, N8456, N1393);
nand NAND3 (N8460, N8454, N989, N1358);
and AND3 (N8461, N8458, N3517, N4656);
buf BUF1 (N8462, N8428);
buf BUF1 (N8463, N8445);
xor XOR2 (N8464, N8440, N3619);
buf BUF1 (N8465, N8460);
xor XOR2 (N8466, N8459, N4874);
and AND2 (N8467, N8466, N5495);
nand NAND3 (N8468, N8463, N4323, N4348);
nand NAND4 (N8469, N8462, N1652, N4587, N1187);
and AND4 (N8470, N8461, N6144, N3903, N5390);
nand NAND4 (N8471, N8464, N767, N5728, N4836);
buf BUF1 (N8472, N8470);
or OR2 (N8473, N8449, N1774);
and AND2 (N8474, N8465, N2740);
and AND2 (N8475, N8469, N5062);
nand NAND4 (N8476, N8446, N5625, N1714, N5823);
or OR3 (N8477, N8476, N6775, N6684);
or OR3 (N8478, N8467, N3827, N444);
nand NAND4 (N8479, N8473, N6633, N6011, N7086);
buf BUF1 (N8480, N8479);
and AND4 (N8481, N8477, N5018, N6198, N7544);
nand NAND3 (N8482, N8468, N7162, N248);
or OR3 (N8483, N8471, N6701, N7805);
nor NOR3 (N8484, N8455, N4732, N8298);
or OR4 (N8485, N8452, N3104, N4719, N1802);
or OR2 (N8486, N8485, N138);
nor NOR2 (N8487, N8474, N5849);
not NOT1 (N8488, N8484);
not NOT1 (N8489, N8481);
nor NOR3 (N8490, N8489, N1852, N289);
or OR2 (N8491, N8478, N5694);
nor NOR3 (N8492, N8475, N5760, N364);
nor NOR4 (N8493, N8480, N6808, N1420, N2450);
xor XOR2 (N8494, N8492, N2717);
nand NAND2 (N8495, N8490, N7527);
and AND3 (N8496, N8494, N6925, N4144);
not NOT1 (N8497, N8483);
or OR3 (N8498, N8472, N4564, N2485);
not NOT1 (N8499, N8482);
nor NOR3 (N8500, N8491, N171, N5687);
or OR2 (N8501, N8499, N5898);
nor NOR2 (N8502, N8501, N5193);
buf BUF1 (N8503, N8496);
nor NOR2 (N8504, N8503, N6920);
not NOT1 (N8505, N8498);
nand NAND2 (N8506, N8487, N1963);
xor XOR2 (N8507, N8500, N2216);
nand NAND2 (N8508, N8497, N3452);
xor XOR2 (N8509, N8495, N5822);
xor XOR2 (N8510, N8507, N5757);
not NOT1 (N8511, N8488);
nor NOR4 (N8512, N8504, N3698, N2514, N7);
and AND4 (N8513, N8508, N7355, N4851, N5216);
or OR2 (N8514, N8512, N1723);
and AND3 (N8515, N8493, N1580, N6362);
or OR4 (N8516, N8506, N6515, N2063, N4859);
nand NAND2 (N8517, N8513, N3468);
buf BUF1 (N8518, N8514);
or OR2 (N8519, N8518, N2944);
xor XOR2 (N8520, N8511, N7090);
and AND3 (N8521, N8516, N4375, N3378);
or OR3 (N8522, N8520, N4047, N3890);
nand NAND3 (N8523, N8519, N7639, N1783);
not NOT1 (N8524, N8486);
or OR4 (N8525, N8521, N2817, N4436, N7797);
xor XOR2 (N8526, N8517, N6091);
xor XOR2 (N8527, N8524, N6878);
nand NAND3 (N8528, N8510, N3540, N4232);
nand NAND2 (N8529, N8509, N1233);
not NOT1 (N8530, N8529);
and AND4 (N8531, N8505, N3151, N3024, N5579);
nand NAND4 (N8532, N8526, N6035, N5011, N2720);
and AND3 (N8533, N8528, N6578, N4998);
nand NAND4 (N8534, N8530, N7222, N3983, N648);
nor NOR4 (N8535, N8502, N6715, N4401, N5903);
buf BUF1 (N8536, N8532);
xor XOR2 (N8537, N8522, N3496);
or OR3 (N8538, N8515, N8529, N5343);
buf BUF1 (N8539, N8537);
nor NOR4 (N8540, N8536, N3254, N1019, N3188);
buf BUF1 (N8541, N8527);
nand NAND3 (N8542, N8538, N7953, N3201);
buf BUF1 (N8543, N8534);
not NOT1 (N8544, N8543);
xor XOR2 (N8545, N8544, N8429);
xor XOR2 (N8546, N8525, N5932);
not NOT1 (N8547, N8539);
or OR2 (N8548, N8535, N2916);
buf BUF1 (N8549, N8541);
and AND3 (N8550, N8549, N7919, N7359);
buf BUF1 (N8551, N8546);
or OR4 (N8552, N8547, N4285, N1720, N7576);
nand NAND3 (N8553, N8523, N293, N6929);
nand NAND3 (N8554, N8531, N5664, N5335);
and AND4 (N8555, N8533, N7926, N1528, N7322);
not NOT1 (N8556, N8548);
and AND4 (N8557, N8555, N7630, N7296, N5903);
xor XOR2 (N8558, N8540, N6592);
nand NAND3 (N8559, N8550, N6464, N442);
nor NOR2 (N8560, N8542, N5936);
buf BUF1 (N8561, N8559);
or OR2 (N8562, N8545, N1453);
nand NAND3 (N8563, N8561, N1732, N2727);
not NOT1 (N8564, N8563);
xor XOR2 (N8565, N8564, N3495);
and AND2 (N8566, N8565, N213);
nand NAND4 (N8567, N8558, N5836, N7116, N5950);
or OR2 (N8568, N8554, N1292);
not NOT1 (N8569, N8557);
or OR3 (N8570, N8552, N214, N2689);
and AND3 (N8571, N8568, N7898, N4674);
or OR3 (N8572, N8562, N2647, N4605);
and AND4 (N8573, N8556, N3270, N485, N3744);
not NOT1 (N8574, N8567);
or OR2 (N8575, N8560, N1263);
not NOT1 (N8576, N8575);
xor XOR2 (N8577, N8573, N6832);
nand NAND2 (N8578, N8571, N7823);
not NOT1 (N8579, N8551);
and AND4 (N8580, N8579, N3248, N5101, N2262);
buf BUF1 (N8581, N8576);
or OR2 (N8582, N8580, N5367);
and AND2 (N8583, N8566, N4755);
not NOT1 (N8584, N8570);
nor NOR3 (N8585, N8581, N1386, N3853);
xor XOR2 (N8586, N8577, N6722);
buf BUF1 (N8587, N8574);
or OR3 (N8588, N8553, N2603, N4800);
or OR4 (N8589, N8585, N5292, N2339, N7535);
nor NOR2 (N8590, N8588, N1009);
nand NAND3 (N8591, N8584, N8179, N265);
not NOT1 (N8592, N8582);
buf BUF1 (N8593, N8586);
buf BUF1 (N8594, N8593);
or OR4 (N8595, N8572, N2181, N1721, N5777);
buf BUF1 (N8596, N8594);
xor XOR2 (N8597, N8578, N2747);
or OR3 (N8598, N8591, N710, N8301);
buf BUF1 (N8599, N8597);
or OR4 (N8600, N8599, N312, N554, N6279);
not NOT1 (N8601, N8595);
buf BUF1 (N8602, N8587);
nor NOR4 (N8603, N8601, N4569, N6102, N543);
or OR2 (N8604, N8603, N4335);
not NOT1 (N8605, N8569);
and AND3 (N8606, N8590, N4482, N6213);
and AND2 (N8607, N8592, N7254);
and AND2 (N8608, N8600, N2311);
nor NOR2 (N8609, N8602, N6649);
nand NAND4 (N8610, N8596, N6665, N5487, N4628);
buf BUF1 (N8611, N8606);
buf BUF1 (N8612, N8604);
xor XOR2 (N8613, N8612, N5152);
xor XOR2 (N8614, N8583, N4180);
nor NOR2 (N8615, N8613, N546);
nand NAND2 (N8616, N8608, N7766);
or OR2 (N8617, N8605, N8103);
nand NAND2 (N8618, N8615, N7453);
or OR3 (N8619, N8589, N6945, N241);
or OR3 (N8620, N8609, N3674, N5884);
or OR2 (N8621, N8617, N5451);
not NOT1 (N8622, N8616);
nand NAND3 (N8623, N8614, N6589, N1191);
and AND2 (N8624, N8611, N8488);
not NOT1 (N8625, N8622);
buf BUF1 (N8626, N8619);
nand NAND2 (N8627, N8607, N1752);
not NOT1 (N8628, N8610);
and AND2 (N8629, N8620, N4445);
and AND2 (N8630, N8625, N7484);
nand NAND4 (N8631, N8598, N2445, N4389, N5364);
nor NOR2 (N8632, N8631, N22);
buf BUF1 (N8633, N8624);
nor NOR3 (N8634, N8627, N8557, N5719);
nor NOR4 (N8635, N8626, N5033, N5206, N2436);
or OR4 (N8636, N8633, N581, N2723, N2602);
not NOT1 (N8637, N8636);
nand NAND3 (N8638, N8632, N3129, N2186);
or OR2 (N8639, N8634, N6005);
or OR2 (N8640, N8630, N6804);
not NOT1 (N8641, N8621);
nor NOR4 (N8642, N8623, N6593, N3236, N5128);
nand NAND2 (N8643, N8635, N7477);
and AND4 (N8644, N8618, N4756, N8379, N6571);
and AND3 (N8645, N8641, N8209, N133);
buf BUF1 (N8646, N8629);
not NOT1 (N8647, N8628);
and AND2 (N8648, N8647, N8531);
xor XOR2 (N8649, N8638, N1627);
xor XOR2 (N8650, N8639, N8481);
buf BUF1 (N8651, N8642);
nor NOR4 (N8652, N8650, N4092, N3867, N60);
nand NAND2 (N8653, N8645, N8364);
or OR4 (N8654, N8646, N4001, N986, N621);
not NOT1 (N8655, N8653);
nor NOR2 (N8656, N8651, N1329);
xor XOR2 (N8657, N8644, N3828);
nand NAND3 (N8658, N8656, N5088, N7524);
and AND4 (N8659, N8649, N5455, N4068, N615);
nor NOR4 (N8660, N8659, N1440, N2119, N5190);
nor NOR2 (N8661, N8657, N4265);
and AND4 (N8662, N8637, N4244, N6576, N6030);
not NOT1 (N8663, N8661);
xor XOR2 (N8664, N8652, N1167);
buf BUF1 (N8665, N8654);
nor NOR3 (N8666, N8643, N3738, N630);
xor XOR2 (N8667, N8663, N3046);
buf BUF1 (N8668, N8667);
and AND2 (N8669, N8655, N5724);
and AND2 (N8670, N8648, N3454);
and AND2 (N8671, N8662, N319);
not NOT1 (N8672, N8658);
nand NAND2 (N8673, N8665, N4829);
and AND4 (N8674, N8669, N6220, N4081, N1341);
nand NAND3 (N8675, N8674, N214, N1463);
nand NAND4 (N8676, N8664, N5725, N5297, N7267);
nor NOR4 (N8677, N8640, N7113, N2951, N5121);
nor NOR4 (N8678, N8671, N2320, N5948, N7602);
or OR2 (N8679, N8676, N232);
or OR2 (N8680, N8660, N536);
nor NOR3 (N8681, N8672, N7749, N2007);
or OR2 (N8682, N8675, N7046);
buf BUF1 (N8683, N8682);
nand NAND3 (N8684, N8668, N6494, N6096);
and AND3 (N8685, N8673, N7266, N844);
buf BUF1 (N8686, N8684);
nand NAND4 (N8687, N8678, N3820, N3756, N8190);
and AND2 (N8688, N8679, N4104);
xor XOR2 (N8689, N8685, N8091);
xor XOR2 (N8690, N8670, N2559);
or OR4 (N8691, N8689, N4359, N1199, N2271);
nand NAND2 (N8692, N8691, N68);
or OR2 (N8693, N8666, N4063);
buf BUF1 (N8694, N8692);
not NOT1 (N8695, N8681);
nand NAND3 (N8696, N8690, N20, N6951);
xor XOR2 (N8697, N8687, N3220);
nand NAND2 (N8698, N8694, N3139);
nand NAND4 (N8699, N8680, N3064, N7076, N8003);
nand NAND2 (N8700, N8677, N559);
buf BUF1 (N8701, N8697);
and AND2 (N8702, N8696, N6438);
or OR3 (N8703, N8700, N3116, N115);
or OR2 (N8704, N8693, N1421);
nand NAND3 (N8705, N8686, N8481, N5329);
nand NAND3 (N8706, N8698, N5455, N7686);
and AND2 (N8707, N8695, N3786);
or OR2 (N8708, N8683, N2035);
and AND4 (N8709, N8705, N1017, N537, N7772);
not NOT1 (N8710, N8702);
buf BUF1 (N8711, N8706);
or OR3 (N8712, N8709, N2599, N2777);
or OR2 (N8713, N8710, N3814);
and AND3 (N8714, N8707, N6730, N422);
and AND2 (N8715, N8688, N6196);
and AND4 (N8716, N8701, N3030, N5546, N5373);
or OR4 (N8717, N8716, N7647, N3592, N1588);
and AND2 (N8718, N8711, N3958);
and AND3 (N8719, N8718, N1966, N5589);
buf BUF1 (N8720, N8708);
or OR2 (N8721, N8715, N6429);
and AND3 (N8722, N8721, N6253, N6631);
and AND4 (N8723, N8699, N6312, N6850, N6638);
not NOT1 (N8724, N8719);
xor XOR2 (N8725, N8712, N1329);
and AND3 (N8726, N8722, N1920, N771);
nand NAND2 (N8727, N8703, N5931);
and AND3 (N8728, N8714, N139, N8459);
and AND4 (N8729, N8713, N6873, N1181, N4463);
xor XOR2 (N8730, N8727, N8080);
nand NAND2 (N8731, N8720, N4809);
xor XOR2 (N8732, N8729, N379);
or OR3 (N8733, N8726, N5667, N3314);
not NOT1 (N8734, N8724);
and AND4 (N8735, N8717, N7630, N3539, N1930);
xor XOR2 (N8736, N8732, N2159);
and AND2 (N8737, N8731, N6299);
or OR3 (N8738, N8728, N1485, N4617);
nor NOR3 (N8739, N8723, N4187, N1028);
nor NOR2 (N8740, N8725, N8239);
nand NAND3 (N8741, N8737, N4134, N4843);
or OR3 (N8742, N8734, N1553, N5524);
nand NAND3 (N8743, N8735, N2669, N5791);
or OR2 (N8744, N8733, N8582);
nand NAND4 (N8745, N8740, N8483, N2, N4843);
not NOT1 (N8746, N8704);
buf BUF1 (N8747, N8744);
nand NAND3 (N8748, N8742, N2343, N2826);
buf BUF1 (N8749, N8738);
and AND2 (N8750, N8730, N1720);
buf BUF1 (N8751, N8739);
and AND3 (N8752, N8747, N5498, N7240);
xor XOR2 (N8753, N8745, N5354);
nand NAND4 (N8754, N8753, N3103, N5548, N1970);
and AND4 (N8755, N8746, N5858, N5397, N7949);
not NOT1 (N8756, N8754);
buf BUF1 (N8757, N8749);
xor XOR2 (N8758, N8751, N441);
nand NAND2 (N8759, N8750, N2595);
and AND2 (N8760, N8756, N7167);
xor XOR2 (N8761, N8748, N3220);
not NOT1 (N8762, N8736);
or OR4 (N8763, N8755, N427, N6134, N6132);
nand NAND3 (N8764, N8759, N2829, N840);
buf BUF1 (N8765, N8764);
not NOT1 (N8766, N8743);
or OR3 (N8767, N8763, N3785, N8513);
or OR2 (N8768, N8761, N2509);
or OR3 (N8769, N8768, N8369, N6224);
nand NAND3 (N8770, N8752, N3079, N8082);
buf BUF1 (N8771, N8765);
nor NOR3 (N8772, N8758, N2607, N1151);
nand NAND2 (N8773, N8757, N6102);
not NOT1 (N8774, N8769);
xor XOR2 (N8775, N8773, N7239);
buf BUF1 (N8776, N8762);
xor XOR2 (N8777, N8774, N3794);
not NOT1 (N8778, N8760);
xor XOR2 (N8779, N8776, N5496);
not NOT1 (N8780, N8741);
xor XOR2 (N8781, N8780, N1519);
nand NAND2 (N8782, N8778, N3565);
not NOT1 (N8783, N8771);
xor XOR2 (N8784, N8782, N5358);
and AND2 (N8785, N8783, N2328);
and AND3 (N8786, N8770, N1589, N1090);
buf BUF1 (N8787, N8767);
nor NOR4 (N8788, N8787, N1472, N1219, N8046);
buf BUF1 (N8789, N8784);
not NOT1 (N8790, N8781);
not NOT1 (N8791, N8785);
xor XOR2 (N8792, N8790, N7577);
xor XOR2 (N8793, N8772, N2128);
nor NOR3 (N8794, N8793, N1918, N8511);
or OR2 (N8795, N8779, N819);
not NOT1 (N8796, N8786);
xor XOR2 (N8797, N8792, N6753);
or OR2 (N8798, N8795, N14);
buf BUF1 (N8799, N8789);
buf BUF1 (N8800, N8775);
buf BUF1 (N8801, N8777);
nor NOR4 (N8802, N8797, N3924, N7764, N5701);
buf BUF1 (N8803, N8788);
nor NOR4 (N8804, N8794, N6094, N2030, N4007);
nand NAND3 (N8805, N8804, N2541, N7173);
nand NAND4 (N8806, N8800, N3996, N6728, N3169);
nand NAND3 (N8807, N8803, N4839, N1888);
xor XOR2 (N8808, N8799, N1064);
buf BUF1 (N8809, N8807);
and AND4 (N8810, N8809, N2496, N4180, N6286);
nand NAND4 (N8811, N8805, N8412, N7348, N5403);
not NOT1 (N8812, N8766);
nand NAND2 (N8813, N8798, N43);
xor XOR2 (N8814, N8796, N1370);
and AND4 (N8815, N8813, N3152, N3275, N3144);
nand NAND4 (N8816, N8802, N981, N2556, N8611);
and AND4 (N8817, N8810, N1004, N1954, N2205);
xor XOR2 (N8818, N8812, N298);
xor XOR2 (N8819, N8815, N2741);
or OR4 (N8820, N8791, N1037, N7545, N3117);
xor XOR2 (N8821, N8816, N1016);
nand NAND3 (N8822, N8817, N4507, N2865);
nand NAND3 (N8823, N8818, N4637, N4269);
or OR2 (N8824, N8821, N4183);
buf BUF1 (N8825, N8806);
and AND2 (N8826, N8824, N4755);
nand NAND3 (N8827, N8808, N7381, N2150);
xor XOR2 (N8828, N8801, N4736);
nor NOR2 (N8829, N8825, N8433);
xor XOR2 (N8830, N8819, N472);
nor NOR2 (N8831, N8823, N6184);
xor XOR2 (N8832, N8811, N5728);
nand NAND3 (N8833, N8826, N372, N5437);
and AND3 (N8834, N8830, N7295, N3748);
and AND2 (N8835, N8829, N2304);
buf BUF1 (N8836, N8835);
or OR2 (N8837, N8833, N2582);
buf BUF1 (N8838, N8828);
not NOT1 (N8839, N8836);
and AND4 (N8840, N8827, N4149, N2599, N3322);
nor NOR2 (N8841, N8832, N4063);
xor XOR2 (N8842, N8814, N6799);
or OR4 (N8843, N8820, N3370, N5165, N7470);
and AND2 (N8844, N8842, N5416);
or OR3 (N8845, N8838, N59, N355);
nor NOR4 (N8846, N8822, N1716, N1790, N6157);
or OR2 (N8847, N8844, N2022);
not NOT1 (N8848, N8845);
xor XOR2 (N8849, N8847, N7470);
buf BUF1 (N8850, N8831);
and AND4 (N8851, N8837, N6162, N4132, N6805);
and AND3 (N8852, N8841, N5971, N8810);
buf BUF1 (N8853, N8849);
and AND2 (N8854, N8853, N7414);
not NOT1 (N8855, N8850);
or OR4 (N8856, N8839, N830, N6548, N6297);
and AND3 (N8857, N8846, N2670, N7512);
xor XOR2 (N8858, N8840, N200);
or OR3 (N8859, N8843, N6040, N7772);
xor XOR2 (N8860, N8858, N5569);
buf BUF1 (N8861, N8834);
or OR3 (N8862, N8851, N7807, N1554);
and AND4 (N8863, N8854, N1143, N1256, N7850);
nor NOR2 (N8864, N8855, N2292);
nor NOR2 (N8865, N8859, N1545);
buf BUF1 (N8866, N8852);
not NOT1 (N8867, N8848);
not NOT1 (N8868, N8863);
xor XOR2 (N8869, N8867, N6807);
xor XOR2 (N8870, N8869, N2861);
xor XOR2 (N8871, N8857, N7140);
or OR3 (N8872, N8864, N5973, N6869);
not NOT1 (N8873, N8861);
xor XOR2 (N8874, N8872, N1924);
nor NOR3 (N8875, N8871, N4133, N7547);
not NOT1 (N8876, N8868);
nand NAND4 (N8877, N8856, N2817, N1812, N4117);
nand NAND4 (N8878, N8874, N5485, N3743, N6293);
nand NAND3 (N8879, N8876, N7101, N5742);
and AND2 (N8880, N8862, N8675);
buf BUF1 (N8881, N8877);
xor XOR2 (N8882, N8860, N240);
not NOT1 (N8883, N8880);
buf BUF1 (N8884, N8866);
not NOT1 (N8885, N8870);
nand NAND4 (N8886, N8875, N7156, N1356, N8663);
nand NAND4 (N8887, N8873, N8683, N3611, N2005);
nand NAND4 (N8888, N8882, N5576, N6296, N811);
xor XOR2 (N8889, N8885, N6485);
xor XOR2 (N8890, N8888, N3048);
or OR2 (N8891, N8884, N2623);
not NOT1 (N8892, N8883);
xor XOR2 (N8893, N8879, N2125);
buf BUF1 (N8894, N8887);
or OR4 (N8895, N8892, N4820, N1661, N4573);
nand NAND3 (N8896, N8895, N238, N2982);
xor XOR2 (N8897, N8886, N1766);
or OR2 (N8898, N8881, N238);
and AND4 (N8899, N8878, N6507, N2003, N8041);
nor NOR4 (N8900, N8890, N7501, N4250, N3508);
buf BUF1 (N8901, N8865);
nand NAND2 (N8902, N8894, N8166);
not NOT1 (N8903, N8889);
and AND3 (N8904, N8901, N3506, N4789);
xor XOR2 (N8905, N8896, N8610);
or OR2 (N8906, N8899, N7265);
not NOT1 (N8907, N8898);
or OR4 (N8908, N8897, N7857, N6347, N5814);
nand NAND3 (N8909, N8891, N3687, N5385);
not NOT1 (N8910, N8907);
nor NOR3 (N8911, N8902, N4280, N3755);
nand NAND4 (N8912, N8911, N5641, N3144, N3330);
nand NAND2 (N8913, N8906, N7454);
or OR4 (N8914, N8908, N6376, N3397, N16);
or OR2 (N8915, N8900, N1746);
xor XOR2 (N8916, N8915, N124);
or OR3 (N8917, N8914, N1356, N2490);
nor NOR4 (N8918, N8909, N2993, N7697, N1884);
or OR3 (N8919, N8917, N6022, N7633);
not NOT1 (N8920, N8904);
or OR2 (N8921, N8903, N519);
nor NOR4 (N8922, N8920, N3798, N5279, N5950);
nand NAND2 (N8923, N8893, N7144);
xor XOR2 (N8924, N8916, N5784);
or OR2 (N8925, N8918, N7222);
xor XOR2 (N8926, N8913, N4402);
not NOT1 (N8927, N8921);
and AND3 (N8928, N8927, N4788, N2408);
or OR4 (N8929, N8923, N6114, N154, N3523);
not NOT1 (N8930, N8924);
and AND2 (N8931, N8929, N583);
nand NAND4 (N8932, N8930, N727, N5640, N8313);
and AND3 (N8933, N8928, N384, N6509);
nor NOR3 (N8934, N8912, N6968, N6724);
buf BUF1 (N8935, N8925);
or OR3 (N8936, N8910, N5235, N2408);
not NOT1 (N8937, N8919);
and AND2 (N8938, N8934, N2948);
xor XOR2 (N8939, N8922, N7215);
nand NAND2 (N8940, N8936, N646);
buf BUF1 (N8941, N8933);
xor XOR2 (N8942, N8941, N4897);
buf BUF1 (N8943, N8932);
xor XOR2 (N8944, N8935, N1518);
nor NOR4 (N8945, N8937, N8581, N6774, N435);
or OR3 (N8946, N8905, N5584, N7282);
nor NOR4 (N8947, N8944, N8648, N2026, N3676);
not NOT1 (N8948, N8926);
nand NAND2 (N8949, N8940, N1277);
nand NAND3 (N8950, N8949, N3356, N8097);
buf BUF1 (N8951, N8942);
buf BUF1 (N8952, N8943);
and AND3 (N8953, N8952, N4507, N8165);
not NOT1 (N8954, N8946);
xor XOR2 (N8955, N8954, N6387);
nor NOR2 (N8956, N8950, N8540);
nor NOR3 (N8957, N8931, N6516, N6452);
nor NOR4 (N8958, N8945, N5408, N6297, N7497);
nand NAND3 (N8959, N8958, N6600, N3421);
buf BUF1 (N8960, N8957);
buf BUF1 (N8961, N8953);
or OR2 (N8962, N8938, N4219);
and AND2 (N8963, N8947, N1621);
nor NOR2 (N8964, N8955, N5356);
and AND3 (N8965, N8964, N5017, N372);
nand NAND3 (N8966, N8962, N4816, N7933);
nand NAND2 (N8967, N8939, N2779);
not NOT1 (N8968, N8961);
nand NAND3 (N8969, N8948, N3036, N4090);
xor XOR2 (N8970, N8967, N2138);
nor NOR2 (N8971, N8968, N8075);
xor XOR2 (N8972, N8966, N8747);
buf BUF1 (N8973, N8963);
nand NAND2 (N8974, N8973, N8016);
xor XOR2 (N8975, N8972, N8843);
nor NOR4 (N8976, N8959, N2486, N4755, N445);
and AND3 (N8977, N8975, N1111, N6267);
xor XOR2 (N8978, N8976, N2700);
or OR2 (N8979, N8960, N2911);
not NOT1 (N8980, N8965);
not NOT1 (N8981, N8951);
buf BUF1 (N8982, N8978);
not NOT1 (N8983, N8979);
nand NAND3 (N8984, N8980, N314, N4476);
nor NOR2 (N8985, N8981, N4593);
or OR4 (N8986, N8969, N1653, N7422, N4293);
and AND2 (N8987, N8984, N8276);
buf BUF1 (N8988, N8982);
nor NOR2 (N8989, N8974, N1696);
xor XOR2 (N8990, N8987, N1218);
not NOT1 (N8991, N8988);
not NOT1 (N8992, N8971);
not NOT1 (N8993, N8985);
and AND3 (N8994, N8989, N6226, N8213);
nand NAND4 (N8995, N8956, N5999, N359, N5604);
nand NAND3 (N8996, N8983, N3647, N2542);
nand NAND3 (N8997, N8991, N6336, N2772);
nand NAND2 (N8998, N8996, N3053);
buf BUF1 (N8999, N8986);
nand NAND3 (N9000, N8994, N2994, N2279);
and AND2 (N9001, N8997, N3179);
and AND3 (N9002, N9001, N6500, N4012);
nor NOR4 (N9003, N8993, N3495, N4771, N2453);
not NOT1 (N9004, N8992);
buf BUF1 (N9005, N8990);
nor NOR2 (N9006, N8999, N5685);
or OR3 (N9007, N8977, N4301, N4175);
not NOT1 (N9008, N9005);
nor NOR3 (N9009, N9008, N5874, N2817);
xor XOR2 (N9010, N9006, N6532);
xor XOR2 (N9011, N9004, N1347);
nor NOR4 (N9012, N8970, N5122, N1242, N8368);
and AND2 (N9013, N9010, N2151);
nand NAND4 (N9014, N9011, N8570, N6594, N3898);
buf BUF1 (N9015, N9007);
xor XOR2 (N9016, N9002, N3477);
and AND4 (N9017, N9016, N6300, N3608, N3506);
nand NAND4 (N9018, N8995, N8626, N7409, N6603);
xor XOR2 (N9019, N9012, N4822);
nor NOR4 (N9020, N9013, N8046, N1745, N6207);
not NOT1 (N9021, N9003);
nand NAND2 (N9022, N8998, N8976);
xor XOR2 (N9023, N9014, N355);
or OR3 (N9024, N9022, N7253, N1703);
buf BUF1 (N9025, N9024);
or OR4 (N9026, N9019, N8677, N7566, N1826);
xor XOR2 (N9027, N9023, N5614);
or OR3 (N9028, N9025, N8881, N1148);
nor NOR4 (N9029, N9000, N1019, N5269, N3197);
xor XOR2 (N9030, N9026, N5502);
buf BUF1 (N9031, N9021);
or OR4 (N9032, N9027, N3808, N882, N6799);
or OR3 (N9033, N9018, N7812, N5939);
nor NOR4 (N9034, N9009, N7634, N8724, N4447);
nor NOR2 (N9035, N9029, N6758);
not NOT1 (N9036, N9017);
or OR3 (N9037, N9030, N1801, N3024);
and AND4 (N9038, N9020, N422, N3809, N2842);
xor XOR2 (N9039, N9035, N375);
nor NOR4 (N9040, N9034, N1265, N7417, N623);
not NOT1 (N9041, N9033);
xor XOR2 (N9042, N9028, N681);
or OR3 (N9043, N9032, N5305, N2204);
nand NAND2 (N9044, N9015, N6230);
xor XOR2 (N9045, N9037, N2416);
not NOT1 (N9046, N9043);
not NOT1 (N9047, N9041);
and AND2 (N9048, N9039, N8458);
and AND4 (N9049, N9036, N2631, N26, N5757);
nand NAND4 (N9050, N9044, N8696, N1298, N5367);
not NOT1 (N9051, N9040);
not NOT1 (N9052, N9046);
or OR2 (N9053, N9049, N2933);
nand NAND3 (N9054, N9042, N6263, N1185);
buf BUF1 (N9055, N9047);
nor NOR2 (N9056, N9031, N6818);
not NOT1 (N9057, N9054);
and AND3 (N9058, N9057, N8040, N125);
nand NAND3 (N9059, N9058, N977, N5807);
nand NAND2 (N9060, N9038, N1870);
xor XOR2 (N9061, N9045, N1110);
and AND3 (N9062, N9060, N1119, N5801);
buf BUF1 (N9063, N9056);
or OR2 (N9064, N9063, N7376);
and AND4 (N9065, N9062, N6446, N980, N3112);
and AND2 (N9066, N9051, N4649);
not NOT1 (N9067, N9052);
or OR2 (N9068, N9048, N7272);
not NOT1 (N9069, N9067);
or OR2 (N9070, N9064, N5277);
or OR2 (N9071, N9061, N2618);
nor NOR3 (N9072, N9069, N1635, N6599);
or OR4 (N9073, N9050, N6085, N1553, N5067);
buf BUF1 (N9074, N9066);
xor XOR2 (N9075, N9072, N4577);
buf BUF1 (N9076, N9073);
or OR2 (N9077, N9070, N7492);
or OR3 (N9078, N9074, N1164, N7018);
buf BUF1 (N9079, N9075);
or OR3 (N9080, N9059, N1828, N7740);
xor XOR2 (N9081, N9079, N5659);
xor XOR2 (N9082, N9081, N3982);
or OR3 (N9083, N9068, N7212, N8249);
not NOT1 (N9084, N9078);
nor NOR3 (N9085, N9077, N8026, N807);
nand NAND2 (N9086, N9071, N5952);
nor NOR3 (N9087, N9085, N3282, N7343);
or OR4 (N9088, N9083, N6589, N8778, N8406);
nor NOR2 (N9089, N9055, N4035);
and AND4 (N9090, N9065, N7189, N5310, N7260);
xor XOR2 (N9091, N9090, N1451);
xor XOR2 (N9092, N9087, N1432);
nand NAND4 (N9093, N9080, N8542, N1867, N2099);
not NOT1 (N9094, N9053);
not NOT1 (N9095, N9076);
or OR4 (N9096, N9088, N572, N7670, N7217);
nor NOR4 (N9097, N9084, N7102, N8392, N3236);
not NOT1 (N9098, N9092);
buf BUF1 (N9099, N9091);
nand NAND3 (N9100, N9096, N7196, N2447);
buf BUF1 (N9101, N9086);
xor XOR2 (N9102, N9101, N4657);
nand NAND3 (N9103, N9089, N2845, N1190);
not NOT1 (N9104, N9100);
xor XOR2 (N9105, N9094, N877);
or OR2 (N9106, N9099, N3911);
not NOT1 (N9107, N9105);
not NOT1 (N9108, N9093);
xor XOR2 (N9109, N9082, N2033);
or OR2 (N9110, N9103, N7028);
buf BUF1 (N9111, N9109);
buf BUF1 (N9112, N9111);
and AND4 (N9113, N9107, N2583, N8104, N4490);
buf BUF1 (N9114, N9098);
or OR3 (N9115, N9104, N4086, N5048);
xor XOR2 (N9116, N9115, N4764);
and AND3 (N9117, N9112, N4756, N8735);
or OR4 (N9118, N9117, N7943, N8346, N8403);
xor XOR2 (N9119, N9106, N1717);
buf BUF1 (N9120, N9114);
buf BUF1 (N9121, N9116);
and AND4 (N9122, N9118, N4688, N7083, N5742);
not NOT1 (N9123, N9108);
buf BUF1 (N9124, N9119);
buf BUF1 (N9125, N9102);
nor NOR3 (N9126, N9121, N7372, N8344);
or OR4 (N9127, N9124, N3304, N4162, N4045);
nand NAND3 (N9128, N9127, N4376, N3937);
buf BUF1 (N9129, N9123);
xor XOR2 (N9130, N9110, N8113);
xor XOR2 (N9131, N9130, N8292);
not NOT1 (N9132, N9120);
not NOT1 (N9133, N9113);
and AND4 (N9134, N9133, N1589, N2990, N2952);
not NOT1 (N9135, N9128);
nand NAND2 (N9136, N9131, N538);
nand NAND2 (N9137, N9097, N4553);
and AND2 (N9138, N9134, N9104);
and AND3 (N9139, N9122, N3135, N8884);
and AND3 (N9140, N9139, N1840, N1438);
nand NAND3 (N9141, N9129, N6767, N7894);
and AND4 (N9142, N9141, N6253, N2059, N215);
xor XOR2 (N9143, N9136, N4883);
or OR2 (N9144, N9137, N4337);
buf BUF1 (N9145, N9140);
nor NOR4 (N9146, N9142, N6965, N4892, N4562);
nor NOR2 (N9147, N9143, N944);
xor XOR2 (N9148, N9146, N8735);
and AND2 (N9149, N9135, N5232);
or OR3 (N9150, N9125, N3054, N8280);
nor NOR4 (N9151, N9144, N5671, N7932, N8465);
nand NAND2 (N9152, N9147, N8293);
or OR3 (N9153, N9151, N7648, N19);
not NOT1 (N9154, N9132);
buf BUF1 (N9155, N9138);
and AND4 (N9156, N9095, N3107, N7588, N3298);
and AND4 (N9157, N9154, N6009, N8684, N4014);
and AND2 (N9158, N9157, N7537);
nor NOR2 (N9159, N9150, N7704);
nor NOR2 (N9160, N9159, N693);
not NOT1 (N9161, N9156);
xor XOR2 (N9162, N9126, N8521);
nor NOR3 (N9163, N9148, N985, N1882);
nand NAND2 (N9164, N9155, N4218);
nor NOR4 (N9165, N9158, N8152, N3446, N7931);
and AND2 (N9166, N9152, N413);
nor NOR2 (N9167, N9164, N5101);
nor NOR4 (N9168, N9162, N7833, N4312, N3047);
xor XOR2 (N9169, N9145, N48);
and AND4 (N9170, N9149, N4157, N7148, N2777);
not NOT1 (N9171, N9160);
xor XOR2 (N9172, N9161, N7391);
not NOT1 (N9173, N9172);
and AND4 (N9174, N9173, N7483, N1834, N9172);
nand NAND4 (N9175, N9167, N3670, N7361, N619);
not NOT1 (N9176, N9174);
not NOT1 (N9177, N9163);
xor XOR2 (N9178, N9176, N3626);
nand NAND3 (N9179, N9168, N2607, N4391);
buf BUF1 (N9180, N9171);
nand NAND3 (N9181, N9166, N999, N5672);
or OR4 (N9182, N9170, N5441, N8620, N5670);
not NOT1 (N9183, N9169);
nor NOR4 (N9184, N9177, N534, N1680, N300);
and AND4 (N9185, N9183, N6426, N3977, N4836);
and AND2 (N9186, N9182, N4764);
and AND2 (N9187, N9179, N4763);
and AND2 (N9188, N9165, N7567);
buf BUF1 (N9189, N9188);
nor NOR4 (N9190, N9186, N5464, N1513, N9071);
xor XOR2 (N9191, N9175, N432);
nor NOR3 (N9192, N9189, N2332, N5268);
buf BUF1 (N9193, N9185);
nor NOR2 (N9194, N9190, N3724);
xor XOR2 (N9195, N9178, N6665);
nor NOR4 (N9196, N9191, N266, N5478, N1920);
and AND3 (N9197, N9184, N3814, N596);
and AND3 (N9198, N9180, N2580, N8600);
not NOT1 (N9199, N9194);
nand NAND4 (N9200, N9187, N8568, N3778, N532);
xor XOR2 (N9201, N9199, N6548);
not NOT1 (N9202, N9198);
nor NOR3 (N9203, N9193, N6151, N5404);
nor NOR2 (N9204, N9196, N5533);
buf BUF1 (N9205, N9201);
or OR4 (N9206, N9181, N1984, N6366, N4416);
not NOT1 (N9207, N9195);
buf BUF1 (N9208, N9200);
buf BUF1 (N9209, N9202);
xor XOR2 (N9210, N9205, N2568);
buf BUF1 (N9211, N9210);
xor XOR2 (N9212, N9153, N6839);
buf BUF1 (N9213, N9197);
xor XOR2 (N9214, N9209, N5682);
nor NOR3 (N9215, N9206, N9118, N9167);
or OR2 (N9216, N9213, N3294);
or OR4 (N9217, N9214, N5530, N2033, N2245);
and AND4 (N9218, N9192, N1543, N6129, N7877);
or OR4 (N9219, N9218, N6641, N6499, N7474);
buf BUF1 (N9220, N9212);
not NOT1 (N9221, N9204);
and AND2 (N9222, N9203, N3331);
not NOT1 (N9223, N9219);
nand NAND3 (N9224, N9207, N4921, N7377);
and AND2 (N9225, N9222, N3703);
nor NOR3 (N9226, N9224, N7653, N6569);
xor XOR2 (N9227, N9221, N533);
xor XOR2 (N9228, N9225, N7632);
nand NAND3 (N9229, N9227, N60, N2623);
buf BUF1 (N9230, N9211);
nand NAND3 (N9231, N9229, N3511, N5239);
buf BUF1 (N9232, N9220);
or OR2 (N9233, N9223, N3731);
xor XOR2 (N9234, N9215, N8843);
and AND2 (N9235, N9208, N3397);
not NOT1 (N9236, N9233);
nand NAND3 (N9237, N9235, N879, N7419);
and AND4 (N9238, N9236, N9015, N4034, N7140);
xor XOR2 (N9239, N9232, N7045);
or OR4 (N9240, N9234, N4646, N767, N2761);
nand NAND3 (N9241, N9239, N4959, N5777);
buf BUF1 (N9242, N9226);
xor XOR2 (N9243, N9241, N725);
nand NAND2 (N9244, N9216, N7854);
not NOT1 (N9245, N9237);
and AND3 (N9246, N9230, N5483, N6299);
nor NOR3 (N9247, N9217, N5491, N202);
not NOT1 (N9248, N9238);
buf BUF1 (N9249, N9231);
not NOT1 (N9250, N9249);
not NOT1 (N9251, N9246);
not NOT1 (N9252, N9244);
buf BUF1 (N9253, N9245);
or OR4 (N9254, N9250, N7289, N6912, N15);
buf BUF1 (N9255, N9251);
buf BUF1 (N9256, N9254);
or OR4 (N9257, N9255, N2452, N4248, N1910);
xor XOR2 (N9258, N9228, N8461);
or OR4 (N9259, N9247, N3873, N8470, N5457);
nor NOR4 (N9260, N9258, N5654, N3553, N8695);
and AND4 (N9261, N9259, N4614, N6210, N3298);
nor NOR3 (N9262, N9261, N1363, N3943);
nor NOR4 (N9263, N9243, N7754, N6286, N1009);
not NOT1 (N9264, N9260);
nand NAND2 (N9265, N9242, N4844);
or OR2 (N9266, N9262, N2189);
buf BUF1 (N9267, N9253);
xor XOR2 (N9268, N9248, N1905);
nand NAND4 (N9269, N9257, N4800, N2253, N7658);
nor NOR3 (N9270, N9267, N4783, N4954);
nor NOR4 (N9271, N9240, N4720, N7236, N6641);
or OR3 (N9272, N9268, N2748, N3972);
and AND3 (N9273, N9271, N3636, N7323);
or OR3 (N9274, N9263, N5661, N57);
or OR2 (N9275, N9266, N5169);
buf BUF1 (N9276, N9256);
and AND3 (N9277, N9275, N4658, N8664);
nand NAND3 (N9278, N9272, N8453, N3881);
not NOT1 (N9279, N9273);
and AND4 (N9280, N9278, N3083, N5614, N4142);
buf BUF1 (N9281, N9270);
nor NOR3 (N9282, N9276, N2232, N2450);
buf BUF1 (N9283, N9252);
nand NAND4 (N9284, N9282, N3218, N6373, N6595);
or OR3 (N9285, N9279, N6619, N3250);
nand NAND4 (N9286, N9264, N1339, N1933, N2892);
or OR2 (N9287, N9284, N4416);
nor NOR4 (N9288, N9285, N6796, N5804, N8207);
nor NOR2 (N9289, N9274, N2946);
buf BUF1 (N9290, N9288);
buf BUF1 (N9291, N9290);
nand NAND2 (N9292, N9265, N6834);
or OR3 (N9293, N9287, N4455, N7090);
xor XOR2 (N9294, N9286, N5895);
nor NOR2 (N9295, N9280, N7468);
nand NAND2 (N9296, N9295, N5445);
nand NAND3 (N9297, N9281, N5286, N8974);
xor XOR2 (N9298, N9293, N3234);
nand NAND3 (N9299, N9283, N54, N7576);
nand NAND2 (N9300, N9291, N8724);
or OR3 (N9301, N9294, N1530, N4469);
xor XOR2 (N9302, N9277, N1007);
nand NAND3 (N9303, N9296, N965, N6153);
and AND4 (N9304, N9303, N948, N1494, N6548);
not NOT1 (N9305, N9289);
xor XOR2 (N9306, N9292, N1958);
not NOT1 (N9307, N9304);
or OR3 (N9308, N9297, N7037, N4692);
xor XOR2 (N9309, N9269, N1089);
xor XOR2 (N9310, N9302, N5865);
xor XOR2 (N9311, N9307, N3137);
buf BUF1 (N9312, N9299);
not NOT1 (N9313, N9300);
nand NAND4 (N9314, N9309, N1330, N68, N2298);
nor NOR4 (N9315, N9305, N5115, N8388, N7769);
nor NOR2 (N9316, N9313, N959);
nand NAND2 (N9317, N9308, N9041);
nor NOR4 (N9318, N9301, N3666, N3214, N9175);
not NOT1 (N9319, N9317);
buf BUF1 (N9320, N9316);
not NOT1 (N9321, N9318);
nor NOR4 (N9322, N9321, N1796, N8248, N2617);
and AND3 (N9323, N9314, N9303, N6508);
nor NOR4 (N9324, N9320, N1854, N419, N2399);
and AND2 (N9325, N9298, N2070);
xor XOR2 (N9326, N9322, N7431);
and AND2 (N9327, N9326, N8186);
nand NAND4 (N9328, N9324, N5553, N9148, N751);
nand NAND3 (N9329, N9325, N3909, N1107);
buf BUF1 (N9330, N9312);
and AND4 (N9331, N9319, N5576, N50, N1035);
or OR4 (N9332, N9331, N2260, N7809, N686);
buf BUF1 (N9333, N9332);
xor XOR2 (N9334, N9327, N1482);
nor NOR2 (N9335, N9333, N576);
nor NOR4 (N9336, N9315, N8116, N516, N7441);
and AND4 (N9337, N9336, N4587, N6588, N7441);
xor XOR2 (N9338, N9310, N8983);
buf BUF1 (N9339, N9334);
nand NAND4 (N9340, N9311, N4434, N2417, N6429);
nand NAND4 (N9341, N9337, N7398, N1259, N3947);
nor NOR3 (N9342, N9306, N9044, N7561);
and AND4 (N9343, N9330, N4950, N2587, N7436);
xor XOR2 (N9344, N9341, N1120);
xor XOR2 (N9345, N9340, N6106);
nand NAND2 (N9346, N9345, N8046);
xor XOR2 (N9347, N9335, N4941);
buf BUF1 (N9348, N9339);
nor NOR2 (N9349, N9348, N3577);
xor XOR2 (N9350, N9342, N4573);
and AND3 (N9351, N9329, N1073, N8574);
buf BUF1 (N9352, N9344);
nor NOR3 (N9353, N9351, N1745, N4253);
or OR2 (N9354, N9346, N2094);
or OR2 (N9355, N9347, N7662);
buf BUF1 (N9356, N9328);
nand NAND3 (N9357, N9338, N1784, N4573);
and AND3 (N9358, N9355, N6736, N4268);
xor XOR2 (N9359, N9353, N3133);
nand NAND3 (N9360, N9350, N4706, N7449);
xor XOR2 (N9361, N9349, N964);
nand NAND2 (N9362, N9360, N8341);
not NOT1 (N9363, N9343);
xor XOR2 (N9364, N9352, N3466);
nor NOR3 (N9365, N9358, N3011, N8614);
xor XOR2 (N9366, N9323, N1518);
nand NAND3 (N9367, N9364, N2572, N5709);
xor XOR2 (N9368, N9361, N1186);
or OR3 (N9369, N9363, N8801, N1703);
nor NOR2 (N9370, N9354, N2501);
or OR2 (N9371, N9357, N3514);
and AND4 (N9372, N9356, N3673, N3628, N6088);
not NOT1 (N9373, N9365);
nand NAND2 (N9374, N9359, N202);
nand NAND2 (N9375, N9370, N9187);
nand NAND4 (N9376, N9374, N6953, N3517, N2416);
not NOT1 (N9377, N9369);
nand NAND4 (N9378, N9377, N6425, N3236, N5364);
not NOT1 (N9379, N9371);
not NOT1 (N9380, N9372);
not NOT1 (N9381, N9362);
xor XOR2 (N9382, N9367, N6250);
or OR4 (N9383, N9378, N2233, N6164, N8002);
and AND2 (N9384, N9381, N5430);
nor NOR4 (N9385, N9368, N5321, N2641, N3888);
nand NAND2 (N9386, N9384, N1665);
not NOT1 (N9387, N9386);
nand NAND2 (N9388, N9376, N2592);
and AND3 (N9389, N9373, N2764, N2076);
nor NOR2 (N9390, N9379, N8939);
nor NOR4 (N9391, N9387, N5463, N8769, N7711);
or OR3 (N9392, N9375, N6106, N3384);
buf BUF1 (N9393, N9391);
and AND2 (N9394, N9385, N4950);
not NOT1 (N9395, N9393);
buf BUF1 (N9396, N9392);
not NOT1 (N9397, N9394);
xor XOR2 (N9398, N9390, N3781);
xor XOR2 (N9399, N9397, N2974);
not NOT1 (N9400, N9380);
nand NAND3 (N9401, N9395, N2520, N5062);
xor XOR2 (N9402, N9396, N9070);
xor XOR2 (N9403, N9366, N7587);
or OR2 (N9404, N9403, N1920);
not NOT1 (N9405, N9401);
nor NOR3 (N9406, N9389, N2261, N701);
not NOT1 (N9407, N9400);
not NOT1 (N9408, N9405);
not NOT1 (N9409, N9398);
not NOT1 (N9410, N9409);
or OR3 (N9411, N9408, N2992, N888);
and AND4 (N9412, N9407, N4684, N7569, N1497);
not NOT1 (N9413, N9412);
nor NOR4 (N9414, N9410, N2814, N598, N7254);
xor XOR2 (N9415, N9399, N3738);
or OR4 (N9416, N9402, N3114, N5379, N6852);
nor NOR4 (N9417, N9406, N7956, N5142, N4728);
xor XOR2 (N9418, N9383, N4691);
and AND4 (N9419, N9382, N3893, N724, N153);
and AND4 (N9420, N9388, N3930, N237, N4341);
buf BUF1 (N9421, N9420);
and AND3 (N9422, N9421, N4005, N8374);
and AND4 (N9423, N9422, N7009, N891, N1208);
buf BUF1 (N9424, N9415);
and AND4 (N9425, N9411, N2801, N6702, N4430);
not NOT1 (N9426, N9423);
or OR2 (N9427, N9419, N825);
xor XOR2 (N9428, N9427, N2299);
xor XOR2 (N9429, N9424, N5519);
and AND3 (N9430, N9413, N7995, N6538);
not NOT1 (N9431, N9417);
buf BUF1 (N9432, N9418);
nor NOR2 (N9433, N9404, N8964);
nand NAND2 (N9434, N9414, N7089);
buf BUF1 (N9435, N9429);
nand NAND2 (N9436, N9430, N1400);
or OR3 (N9437, N9431, N6026, N8803);
nand NAND3 (N9438, N9425, N3981, N1568);
and AND4 (N9439, N9432, N2273, N4960, N1651);
buf BUF1 (N9440, N9428);
or OR3 (N9441, N9434, N4856, N4670);
buf BUF1 (N9442, N9426);
not NOT1 (N9443, N9437);
buf BUF1 (N9444, N9436);
or OR2 (N9445, N9444, N6572);
buf BUF1 (N9446, N9416);
xor XOR2 (N9447, N9442, N2260);
nand NAND3 (N9448, N9446, N1760, N3057);
nor NOR2 (N9449, N9439, N6942);
xor XOR2 (N9450, N9435, N6977);
nand NAND2 (N9451, N9450, N5726);
buf BUF1 (N9452, N9443);
not NOT1 (N9453, N9440);
nand NAND4 (N9454, N9447, N6656, N795, N9059);
and AND4 (N9455, N9433, N8504, N2013, N384);
nand NAND4 (N9456, N9438, N9224, N8259, N2213);
xor XOR2 (N9457, N9455, N239);
buf BUF1 (N9458, N9454);
not NOT1 (N9459, N9448);
and AND4 (N9460, N9458, N4565, N8207, N8754);
nor NOR4 (N9461, N9460, N5017, N928, N2698);
nand NAND3 (N9462, N9451, N7908, N2621);
not NOT1 (N9463, N9441);
or OR3 (N9464, N9457, N1798, N495);
or OR3 (N9465, N9463, N605, N7292);
not NOT1 (N9466, N9462);
and AND2 (N9467, N9449, N5833);
buf BUF1 (N9468, N9464);
buf BUF1 (N9469, N9453);
or OR4 (N9470, N9456, N4648, N6280, N2572);
nand NAND4 (N9471, N9452, N6535, N5773, N42);
buf BUF1 (N9472, N9468);
not NOT1 (N9473, N9465);
nor NOR2 (N9474, N9461, N5812);
and AND3 (N9475, N9445, N691, N5940);
and AND2 (N9476, N9467, N9099);
nor NOR2 (N9477, N9472, N5824);
not NOT1 (N9478, N9473);
buf BUF1 (N9479, N9476);
or OR2 (N9480, N9471, N4365);
and AND3 (N9481, N9477, N2153, N4377);
xor XOR2 (N9482, N9469, N4157);
nand NAND4 (N9483, N9480, N3716, N8048, N3882);
and AND2 (N9484, N9475, N9261);
and AND4 (N9485, N9479, N1717, N2831, N5131);
not NOT1 (N9486, N9470);
or OR2 (N9487, N9485, N8192);
not NOT1 (N9488, N9484);
or OR3 (N9489, N9459, N6472, N2409);
buf BUF1 (N9490, N9474);
nand NAND3 (N9491, N9478, N1000, N3869);
nor NOR4 (N9492, N9481, N4854, N8463, N6367);
xor XOR2 (N9493, N9482, N7016);
nand NAND4 (N9494, N9488, N2366, N292, N6418);
nor NOR4 (N9495, N9486, N7759, N5534, N1543);
nand NAND3 (N9496, N9494, N2159, N942);
not NOT1 (N9497, N9483);
buf BUF1 (N9498, N9487);
nand NAND3 (N9499, N9496, N1835, N6923);
xor XOR2 (N9500, N9497, N8603);
xor XOR2 (N9501, N9489, N7823);
and AND2 (N9502, N9491, N5253);
and AND4 (N9503, N9502, N7687, N2697, N6776);
or OR3 (N9504, N9495, N284, N6221);
buf BUF1 (N9505, N9498);
and AND3 (N9506, N9493, N8859, N6867);
xor XOR2 (N9507, N9490, N375);
xor XOR2 (N9508, N9505, N4119);
xor XOR2 (N9509, N9499, N7838);
nand NAND3 (N9510, N9501, N8411, N7391);
nand NAND4 (N9511, N9509, N4160, N5399, N4235);
nor NOR3 (N9512, N9466, N9036, N2082);
nor NOR4 (N9513, N9507, N9336, N6242, N9117);
nor NOR2 (N9514, N9513, N1343);
xor XOR2 (N9515, N9504, N8496);
or OR4 (N9516, N9508, N6805, N5142, N1145);
xor XOR2 (N9517, N9500, N1590);
or OR3 (N9518, N9514, N4482, N7611);
nor NOR4 (N9519, N9511, N7817, N7667, N6523);
or OR2 (N9520, N9519, N6900);
or OR3 (N9521, N9515, N2356, N9071);
nor NOR3 (N9522, N9512, N4607, N8380);
buf BUF1 (N9523, N9492);
nand NAND2 (N9524, N9503, N2310);
nand NAND4 (N9525, N9521, N5553, N7416, N395);
xor XOR2 (N9526, N9510, N7266);
nor NOR2 (N9527, N9516, N4923);
xor XOR2 (N9528, N9518, N1931);
xor XOR2 (N9529, N9522, N3360);
or OR3 (N9530, N9526, N5325, N5713);
nor NOR2 (N9531, N9530, N3251);
nor NOR4 (N9532, N9517, N5665, N4628, N1004);
buf BUF1 (N9533, N9532);
and AND4 (N9534, N9533, N5167, N8376, N3368);
or OR4 (N9535, N9524, N2543, N8069, N5341);
xor XOR2 (N9536, N9525, N3916);
or OR4 (N9537, N9506, N6010, N1756, N3393);
not NOT1 (N9538, N9536);
nand NAND2 (N9539, N9520, N3777);
buf BUF1 (N9540, N9534);
nand NAND2 (N9541, N9535, N1449);
and AND3 (N9542, N9538, N5150, N1483);
nor NOR2 (N9543, N9528, N5939);
and AND2 (N9544, N9527, N8780);
nand NAND2 (N9545, N9540, N5710);
xor XOR2 (N9546, N9537, N1262);
xor XOR2 (N9547, N9531, N3369);
and AND3 (N9548, N9539, N1184, N796);
buf BUF1 (N9549, N9529);
buf BUF1 (N9550, N9523);
xor XOR2 (N9551, N9542, N6835);
nand NAND2 (N9552, N9549, N831);
nor NOR4 (N9553, N9545, N2419, N7047, N2484);
buf BUF1 (N9554, N9551);
nor NOR3 (N9555, N9553, N8373, N573);
buf BUF1 (N9556, N9555);
xor XOR2 (N9557, N9546, N3055);
xor XOR2 (N9558, N9543, N860);
xor XOR2 (N9559, N9548, N7504);
nand NAND4 (N9560, N9552, N8246, N2619, N3957);
nand NAND2 (N9561, N9558, N4514);
not NOT1 (N9562, N9544);
xor XOR2 (N9563, N9559, N8827);
not NOT1 (N9564, N9550);
or OR3 (N9565, N9561, N6426, N8776);
buf BUF1 (N9566, N9563);
not NOT1 (N9567, N9547);
or OR4 (N9568, N9562, N6741, N8966, N5029);
or OR2 (N9569, N9564, N1000);
nor NOR2 (N9570, N9565, N9103);
not NOT1 (N9571, N9557);
not NOT1 (N9572, N9570);
and AND2 (N9573, N9541, N2032);
not NOT1 (N9574, N9569);
xor XOR2 (N9575, N9571, N5902);
nand NAND3 (N9576, N9566, N1023, N4068);
and AND3 (N9577, N9574, N3160, N2811);
nor NOR3 (N9578, N9577, N665, N3661);
nor NOR3 (N9579, N9556, N7306, N1471);
nor NOR3 (N9580, N9576, N21, N3345);
xor XOR2 (N9581, N9560, N7053);
nor NOR4 (N9582, N9581, N6105, N1109, N5533);
buf BUF1 (N9583, N9579);
nand NAND3 (N9584, N9578, N290, N2567);
and AND3 (N9585, N9582, N7692, N5673);
xor XOR2 (N9586, N9575, N3992);
nor NOR2 (N9587, N9585, N8959);
xor XOR2 (N9588, N9567, N7012);
and AND3 (N9589, N9572, N6760, N1482);
nand NAND3 (N9590, N9573, N1731, N5845);
or OR2 (N9591, N9554, N916);
nor NOR3 (N9592, N9568, N8304, N9488);
nand NAND3 (N9593, N9592, N8058, N7066);
xor XOR2 (N9594, N9593, N1699);
or OR3 (N9595, N9583, N2542, N2300);
buf BUF1 (N9596, N9595);
nand NAND4 (N9597, N9580, N5207, N5074, N2786);
not NOT1 (N9598, N9597);
nor NOR2 (N9599, N9594, N7863);
not NOT1 (N9600, N9588);
nor NOR4 (N9601, N9598, N2743, N7998, N5753);
and AND4 (N9602, N9586, N2165, N4189, N2018);
not NOT1 (N9603, N9599);
not NOT1 (N9604, N9584);
nand NAND4 (N9605, N9587, N3317, N206, N8205);
buf BUF1 (N9606, N9604);
xor XOR2 (N9607, N9589, N2296);
not NOT1 (N9608, N9602);
buf BUF1 (N9609, N9605);
nor NOR4 (N9610, N9596, N4361, N1761, N3828);
not NOT1 (N9611, N9608);
and AND4 (N9612, N9601, N6538, N1361, N298);
or OR3 (N9613, N9591, N3572, N4711);
and AND2 (N9614, N9606, N2460);
or OR4 (N9615, N9611, N517, N7783, N3324);
or OR3 (N9616, N9607, N5572, N3827);
xor XOR2 (N9617, N9609, N238);
buf BUF1 (N9618, N9616);
not NOT1 (N9619, N9612);
xor XOR2 (N9620, N9590, N2470);
not NOT1 (N9621, N9619);
nand NAND4 (N9622, N9615, N7175, N6339, N4472);
buf BUF1 (N9623, N9621);
xor XOR2 (N9624, N9618, N7948);
or OR2 (N9625, N9600, N2644);
not NOT1 (N9626, N9603);
buf BUF1 (N9627, N9617);
nor NOR2 (N9628, N9623, N5533);
nand NAND3 (N9629, N9626, N274, N1385);
buf BUF1 (N9630, N9624);
buf BUF1 (N9631, N9630);
or OR2 (N9632, N9631, N3810);
nand NAND4 (N9633, N9620, N4032, N7773, N8640);
nand NAND4 (N9634, N9625, N5248, N4559, N5931);
and AND2 (N9635, N9629, N7338);
or OR4 (N9636, N9634, N4051, N7126, N2662);
buf BUF1 (N9637, N9613);
nand NAND2 (N9638, N9610, N4061);
not NOT1 (N9639, N9638);
and AND4 (N9640, N9636, N4014, N6670, N7730);
not NOT1 (N9641, N9640);
nand NAND2 (N9642, N9614, N271);
not NOT1 (N9643, N9635);
nand NAND3 (N9644, N9633, N5627, N2291);
nor NOR4 (N9645, N9637, N5356, N7464, N7896);
buf BUF1 (N9646, N9639);
nand NAND4 (N9647, N9632, N839, N7140, N4075);
buf BUF1 (N9648, N9646);
or OR3 (N9649, N9628, N6974, N780);
not NOT1 (N9650, N9644);
buf BUF1 (N9651, N9650);
and AND4 (N9652, N9648, N2563, N5676, N7541);
not NOT1 (N9653, N9622);
xor XOR2 (N9654, N9642, N4722);
nand NAND2 (N9655, N9653, N8796);
buf BUF1 (N9656, N9651);
not NOT1 (N9657, N9647);
nand NAND4 (N9658, N9654, N4041, N3508, N2128);
buf BUF1 (N9659, N9641);
nor NOR2 (N9660, N9643, N3166);
or OR3 (N9661, N9660, N2219, N3289);
not NOT1 (N9662, N9657);
nand NAND4 (N9663, N9661, N501, N3028, N4767);
not NOT1 (N9664, N9652);
buf BUF1 (N9665, N9649);
and AND4 (N9666, N9662, N2569, N7333, N2179);
nor NOR3 (N9667, N9655, N9052, N7024);
nand NAND4 (N9668, N9627, N2873, N3296, N6832);
buf BUF1 (N9669, N9663);
nand NAND3 (N9670, N9669, N5771, N1316);
not NOT1 (N9671, N9667);
not NOT1 (N9672, N9670);
nor NOR4 (N9673, N9645, N8555, N7026, N7177);
and AND2 (N9674, N9668, N3415);
nor NOR2 (N9675, N9659, N3054);
or OR2 (N9676, N9664, N7033);
xor XOR2 (N9677, N9673, N3043);
not NOT1 (N9678, N9665);
not NOT1 (N9679, N9677);
not NOT1 (N9680, N9671);
nor NOR4 (N9681, N9672, N7282, N3547, N5246);
nand NAND3 (N9682, N9658, N614, N6698);
xor XOR2 (N9683, N9679, N243);
or OR2 (N9684, N9656, N3804);
and AND4 (N9685, N9666, N2258, N5741, N693);
not NOT1 (N9686, N9684);
not NOT1 (N9687, N9686);
nor NOR3 (N9688, N9687, N632, N2234);
and AND3 (N9689, N9685, N673, N4766);
nor NOR4 (N9690, N9682, N1381, N1823, N3497);
xor XOR2 (N9691, N9678, N209);
not NOT1 (N9692, N9691);
nor NOR4 (N9693, N9692, N342, N2234, N1972);
buf BUF1 (N9694, N9681);
not NOT1 (N9695, N9674);
xor XOR2 (N9696, N9688, N2793);
or OR3 (N9697, N9695, N5515, N5019);
or OR2 (N9698, N9694, N7947);
and AND4 (N9699, N9697, N8968, N332, N7788);
nand NAND3 (N9700, N9693, N3457, N1310);
nand NAND2 (N9701, N9675, N3529);
or OR3 (N9702, N9690, N367, N5332);
or OR4 (N9703, N9696, N9219, N876, N4619);
buf BUF1 (N9704, N9701);
nor NOR3 (N9705, N9676, N3906, N6964);
nand NAND2 (N9706, N9703, N5321);
and AND2 (N9707, N9680, N6385);
not NOT1 (N9708, N9705);
or OR3 (N9709, N9689, N2005, N972);
not NOT1 (N9710, N9704);
and AND3 (N9711, N9707, N231, N3971);
not NOT1 (N9712, N9700);
or OR3 (N9713, N9712, N1547, N3268);
not NOT1 (N9714, N9698);
or OR4 (N9715, N9714, N6255, N6270, N3636);
buf BUF1 (N9716, N9713);
and AND3 (N9717, N9683, N2861, N8063);
not NOT1 (N9718, N9715);
xor XOR2 (N9719, N9699, N727);
xor XOR2 (N9720, N9708, N8817);
or OR2 (N9721, N9711, N4169);
nor NOR4 (N9722, N9717, N2557, N6460, N3624);
nor NOR2 (N9723, N9710, N5497);
and AND4 (N9724, N9716, N8936, N469, N924);
not NOT1 (N9725, N9718);
not NOT1 (N9726, N9722);
nor NOR2 (N9727, N9725, N5546);
or OR3 (N9728, N9721, N602, N7436);
or OR2 (N9729, N9727, N378);
xor XOR2 (N9730, N9724, N5287);
or OR3 (N9731, N9720, N4373, N4200);
buf BUF1 (N9732, N9729);
nor NOR4 (N9733, N9706, N3835, N8439, N8924);
buf BUF1 (N9734, N9730);
and AND4 (N9735, N9702, N8811, N2150, N907);
xor XOR2 (N9736, N9734, N9259);
and AND3 (N9737, N9731, N4312, N4834);
buf BUF1 (N9738, N9735);
buf BUF1 (N9739, N9728);
buf BUF1 (N9740, N9709);
not NOT1 (N9741, N9736);
xor XOR2 (N9742, N9726, N632);
nand NAND4 (N9743, N9740, N3636, N7171, N2823);
not NOT1 (N9744, N9733);
or OR4 (N9745, N9737, N5613, N9623, N9693);
nor NOR3 (N9746, N9723, N2327, N4594);
nand NAND3 (N9747, N9732, N7090, N1638);
nor NOR3 (N9748, N9747, N521, N7382);
and AND2 (N9749, N9746, N1068);
not NOT1 (N9750, N9749);
nand NAND4 (N9751, N9738, N9443, N5756, N9541);
or OR3 (N9752, N9741, N8547, N7888);
not NOT1 (N9753, N9745);
and AND3 (N9754, N9742, N1651, N8197);
not NOT1 (N9755, N9753);
nand NAND4 (N9756, N9748, N4523, N790, N962);
and AND4 (N9757, N9750, N3830, N9734, N9419);
nor NOR2 (N9758, N9754, N8139);
nand NAND3 (N9759, N9744, N1278, N484);
buf BUF1 (N9760, N9743);
nor NOR3 (N9761, N9719, N8486, N8093);
not NOT1 (N9762, N9755);
not NOT1 (N9763, N9739);
xor XOR2 (N9764, N9761, N3156);
xor XOR2 (N9765, N9764, N7702);
and AND3 (N9766, N9757, N6070, N9532);
xor XOR2 (N9767, N9759, N8692);
not NOT1 (N9768, N9766);
nor NOR4 (N9769, N9756, N1722, N8781, N2025);
buf BUF1 (N9770, N9760);
nand NAND3 (N9771, N9751, N8770, N837);
buf BUF1 (N9772, N9770);
or OR3 (N9773, N9762, N7659, N2590);
not NOT1 (N9774, N9752);
nor NOR3 (N9775, N9772, N856, N7968);
and AND3 (N9776, N9767, N9543, N4011);
buf BUF1 (N9777, N9758);
buf BUF1 (N9778, N9765);
xor XOR2 (N9779, N9774, N7250);
nand NAND2 (N9780, N9778, N480);
and AND4 (N9781, N9771, N9441, N4524, N6770);
buf BUF1 (N9782, N9779);
nor NOR4 (N9783, N9776, N8439, N6485, N1472);
xor XOR2 (N9784, N9763, N7942);
and AND2 (N9785, N9782, N4139);
nor NOR2 (N9786, N9773, N8658);
xor XOR2 (N9787, N9781, N7997);
and AND4 (N9788, N9775, N3548, N1963, N8751);
xor XOR2 (N9789, N9788, N1317);
not NOT1 (N9790, N9780);
xor XOR2 (N9791, N9789, N4488);
not NOT1 (N9792, N9791);
xor XOR2 (N9793, N9787, N5641);
buf BUF1 (N9794, N9786);
nand NAND3 (N9795, N9784, N8468, N8903);
or OR3 (N9796, N9785, N2528, N8830);
or OR2 (N9797, N9769, N4561);
or OR3 (N9798, N9783, N7783, N7409);
and AND4 (N9799, N9792, N8411, N3656, N9510);
buf BUF1 (N9800, N9798);
xor XOR2 (N9801, N9796, N1644);
xor XOR2 (N9802, N9777, N427);
or OR3 (N9803, N9768, N9527, N44);
buf BUF1 (N9804, N9799);
nor NOR2 (N9805, N9790, N113);
nor NOR3 (N9806, N9797, N1044, N1378);
not NOT1 (N9807, N9805);
and AND4 (N9808, N9803, N4339, N858, N340);
not NOT1 (N9809, N9794);
nor NOR4 (N9810, N9801, N3748, N2958, N5985);
nand NAND4 (N9811, N9795, N695, N1812, N7937);
nand NAND4 (N9812, N9808, N5243, N9770, N3821);
or OR2 (N9813, N9810, N3969);
or OR2 (N9814, N9807, N8770);
nand NAND4 (N9815, N9804, N7777, N9346, N5669);
nand NAND4 (N9816, N9814, N7859, N2854, N2102);
not NOT1 (N9817, N9813);
xor XOR2 (N9818, N9811, N5167);
nor NOR2 (N9819, N9809, N3316);
or OR3 (N9820, N9800, N9737, N5675);
or OR2 (N9821, N9819, N9729);
buf BUF1 (N9822, N9816);
nor NOR4 (N9823, N9817, N1230, N5381, N1003);
xor XOR2 (N9824, N9815, N6612);
buf BUF1 (N9825, N9806);
and AND4 (N9826, N9823, N700, N2847, N6152);
and AND2 (N9827, N9825, N5486);
not NOT1 (N9828, N9827);
nand NAND4 (N9829, N9820, N7708, N8599, N2494);
nand NAND3 (N9830, N9821, N2703, N876);
or OR2 (N9831, N9793, N4506);
not NOT1 (N9832, N9826);
not NOT1 (N9833, N9818);
buf BUF1 (N9834, N9802);
nor NOR3 (N9835, N9831, N5151, N9644);
xor XOR2 (N9836, N9828, N7611);
nor NOR3 (N9837, N9834, N5522, N4135);
not NOT1 (N9838, N9822);
and AND3 (N9839, N9830, N6620, N2539);
and AND3 (N9840, N9837, N4718, N2371);
not NOT1 (N9841, N9824);
xor XOR2 (N9842, N9833, N8114);
xor XOR2 (N9843, N9829, N9183);
xor XOR2 (N9844, N9832, N9282);
xor XOR2 (N9845, N9812, N7859);
not NOT1 (N9846, N9841);
and AND2 (N9847, N9846, N6176);
nand NAND3 (N9848, N9847, N8972, N687);
or OR2 (N9849, N9839, N5164);
and AND3 (N9850, N9848, N729, N8707);
nand NAND4 (N9851, N9842, N8337, N2605, N5325);
nand NAND3 (N9852, N9844, N9151, N5265);
and AND4 (N9853, N9835, N6139, N6502, N7491);
xor XOR2 (N9854, N9845, N8861);
nor NOR3 (N9855, N9854, N2068, N9508);
or OR2 (N9856, N9850, N3289);
and AND4 (N9857, N9855, N7196, N1554, N672);
not NOT1 (N9858, N9857);
nand NAND3 (N9859, N9858, N4499, N123);
xor XOR2 (N9860, N9859, N6884);
not NOT1 (N9861, N9840);
not NOT1 (N9862, N9852);
not NOT1 (N9863, N9861);
nand NAND4 (N9864, N9856, N7667, N5864, N3080);
nor NOR2 (N9865, N9862, N3981);
xor XOR2 (N9866, N9860, N3996);
nand NAND3 (N9867, N9838, N1518, N211);
not NOT1 (N9868, N9836);
nor NOR4 (N9869, N9865, N6267, N7941, N2166);
nor NOR3 (N9870, N9867, N8300, N5625);
xor XOR2 (N9871, N9869, N4019);
or OR2 (N9872, N9851, N7788);
and AND3 (N9873, N9871, N81, N7231);
or OR4 (N9874, N9863, N171, N2017, N2595);
buf BUF1 (N9875, N9843);
not NOT1 (N9876, N9870);
nand NAND4 (N9877, N9868, N3393, N2597, N3121);
buf BUF1 (N9878, N9874);
nand NAND3 (N9879, N9875, N3939, N5632);
xor XOR2 (N9880, N9849, N3805);
xor XOR2 (N9881, N9873, N9471);
and AND3 (N9882, N9876, N4948, N7935);
buf BUF1 (N9883, N9880);
xor XOR2 (N9884, N9853, N8296);
or OR2 (N9885, N9872, N9583);
or OR4 (N9886, N9879, N2039, N4377, N9244);
and AND2 (N9887, N9886, N7981);
or OR4 (N9888, N9866, N7083, N5586, N365);
xor XOR2 (N9889, N9864, N2256);
nor NOR4 (N9890, N9882, N58, N7346, N7394);
not NOT1 (N9891, N9878);
xor XOR2 (N9892, N9885, N1891);
not NOT1 (N9893, N9892);
or OR3 (N9894, N9887, N6495, N6263);
or OR2 (N9895, N9881, N5875);
nor NOR2 (N9896, N9888, N2551);
nor NOR4 (N9897, N9889, N6561, N4172, N2547);
nand NAND3 (N9898, N9884, N2426, N3023);
buf BUF1 (N9899, N9898);
or OR4 (N9900, N9896, N9761, N5668, N9328);
not NOT1 (N9901, N9883);
not NOT1 (N9902, N9890);
and AND4 (N9903, N9894, N5728, N5013, N506);
not NOT1 (N9904, N9891);
xor XOR2 (N9905, N9899, N7875);
not NOT1 (N9906, N9903);
nand NAND4 (N9907, N9904, N6111, N8491, N2517);
nand NAND3 (N9908, N9902, N3428, N1813);
nand NAND3 (N9909, N9906, N4473, N5389);
buf BUF1 (N9910, N9905);
not NOT1 (N9911, N9908);
xor XOR2 (N9912, N9910, N2455);
nand NAND3 (N9913, N9909, N7799, N4997);
nor NOR4 (N9914, N9913, N3734, N1982, N1739);
nor NOR4 (N9915, N9907, N73, N4217, N9077);
xor XOR2 (N9916, N9877, N5433);
not NOT1 (N9917, N9911);
buf BUF1 (N9918, N9897);
not NOT1 (N9919, N9916);
and AND2 (N9920, N9917, N6007);
not NOT1 (N9921, N9900);
or OR2 (N9922, N9920, N5069);
nand NAND2 (N9923, N9893, N1868);
buf BUF1 (N9924, N9901);
buf BUF1 (N9925, N9924);
xor XOR2 (N9926, N9923, N2227);
and AND2 (N9927, N9925, N4370);
not NOT1 (N9928, N9912);
and AND2 (N9929, N9915, N9357);
nand NAND3 (N9930, N9929, N6329, N6053);
and AND2 (N9931, N9919, N6050);
xor XOR2 (N9932, N9931, N5810);
xor XOR2 (N9933, N9927, N9919);
xor XOR2 (N9934, N9918, N7306);
buf BUF1 (N9935, N9922);
xor XOR2 (N9936, N9926, N4071);
and AND3 (N9937, N9932, N5264, N2165);
nor NOR2 (N9938, N9930, N8132);
nand NAND2 (N9939, N9934, N1781);
buf BUF1 (N9940, N9921);
nor NOR4 (N9941, N9895, N9393, N4658, N947);
nor NOR2 (N9942, N9935, N8957);
nor NOR3 (N9943, N9938, N1465, N7395);
buf BUF1 (N9944, N9933);
not NOT1 (N9945, N9936);
not NOT1 (N9946, N9944);
nand NAND4 (N9947, N9937, N5712, N5602, N3957);
buf BUF1 (N9948, N9943);
buf BUF1 (N9949, N9946);
buf BUF1 (N9950, N9942);
not NOT1 (N9951, N9950);
and AND3 (N9952, N9940, N9267, N6356);
buf BUF1 (N9953, N9948);
nand NAND2 (N9954, N9947, N2852);
xor XOR2 (N9955, N9953, N6621);
nand NAND4 (N9956, N9941, N2656, N4997, N1580);
nor NOR3 (N9957, N9945, N129, N7687);
nand NAND4 (N9958, N9939, N7287, N6330, N6183);
nor NOR3 (N9959, N9954, N4507, N4116);
buf BUF1 (N9960, N9952);
not NOT1 (N9961, N9960);
not NOT1 (N9962, N9951);
nand NAND4 (N9963, N9962, N4766, N5505, N786);
xor XOR2 (N9964, N9957, N930);
or OR2 (N9965, N9961, N6315);
and AND3 (N9966, N9959, N9146, N8330);
xor XOR2 (N9967, N9914, N241);
buf BUF1 (N9968, N9955);
or OR4 (N9969, N9967, N7266, N5357, N7542);
xor XOR2 (N9970, N9966, N4649);
nand NAND4 (N9971, N9965, N6472, N2103, N4610);
or OR4 (N9972, N9963, N4784, N7472, N6389);
nand NAND3 (N9973, N9949, N3575, N584);
not NOT1 (N9974, N9973);
nor NOR2 (N9975, N9956, N6608);
buf BUF1 (N9976, N9964);
nor NOR3 (N9977, N9928, N7188, N1966);
not NOT1 (N9978, N9971);
buf BUF1 (N9979, N9970);
nand NAND2 (N9980, N9976, N8553);
and AND3 (N9981, N9975, N7789, N4337);
or OR4 (N9982, N9969, N5290, N6928, N4716);
nand NAND3 (N9983, N9978, N6319, N2044);
and AND2 (N9984, N9977, N4174);
xor XOR2 (N9985, N9980, N3748);
not NOT1 (N9986, N9981);
xor XOR2 (N9987, N9958, N8541);
and AND4 (N9988, N9972, N443, N9294, N9466);
and AND2 (N9989, N9986, N1931);
nor NOR3 (N9990, N9983, N6530, N6899);
or OR3 (N9991, N9974, N5771, N8362);
buf BUF1 (N9992, N9987);
nand NAND4 (N9993, N9989, N7390, N3679, N6042);
not NOT1 (N9994, N9982);
nand NAND3 (N9995, N9994, N4189, N504);
nor NOR2 (N9996, N9984, N7390);
xor XOR2 (N9997, N9979, N8969);
xor XOR2 (N9998, N9985, N4661);
and AND3 (N9999, N9991, N1200, N459);
buf BUF1 (N10000, N9996);
not NOT1 (N10001, N9992);
xor XOR2 (N10002, N9993, N3172);
nor NOR2 (N10003, N9990, N4383);
or OR3 (N10004, N9988, N8887, N8455);
or OR3 (N10005, N9968, N494, N2003);
not NOT1 (N10006, N10000);
buf BUF1 (N10007, N9995);
not NOT1 (N10008, N10001);
nand NAND3 (N10009, N10003, N8964, N7814);
nand NAND2 (N10010, N9999, N2111);
buf BUF1 (N10011, N10009);
and AND2 (N10012, N10008, N5928);
not NOT1 (N10013, N10011);
nand NAND4 (N10014, N10013, N4103, N3086, N3625);
and AND2 (N10015, N10010, N6391);
and AND3 (N10016, N10012, N7966, N7318);
and AND4 (N10017, N10006, N8063, N2788, N7779);
nor NOR3 (N10018, N10014, N8075, N8586);
nand NAND4 (N10019, N10007, N6029, N3198, N2998);
not NOT1 (N10020, N10017);
or OR4 (N10021, N10005, N3181, N9635, N9428);
and AND4 (N10022, N10002, N5096, N3002, N457);
not NOT1 (N10023, N10020);
nand NAND4 (N10024, N10019, N62, N5459, N5748);
nor NOR4 (N10025, N10004, N1400, N8531, N8746);
and AND2 (N10026, N10021, N7568);
and AND3 (N10027, N10015, N4629, N177);
not NOT1 (N10028, N10016);
buf BUF1 (N10029, N10024);
nand NAND3 (N10030, N10022, N8351, N8973);
buf BUF1 (N10031, N10028);
nand NAND2 (N10032, N10026, N5257);
and AND4 (N10033, N9998, N6760, N9979, N6208);
nand NAND4 (N10034, N10030, N5744, N5655, N3857);
or OR4 (N10035, N10027, N73, N5597, N7482);
xor XOR2 (N10036, N10023, N4437);
not NOT1 (N10037, N10025);
and AND3 (N10038, N10033, N7648, N1006);
or OR4 (N10039, N10029, N8502, N9287, N4494);
nor NOR3 (N10040, N10018, N2981, N4177);
nor NOR3 (N10041, N10035, N7630, N753);
or OR2 (N10042, N10040, N9359);
and AND3 (N10043, N10039, N2405, N7910);
not NOT1 (N10044, N10043);
nor NOR4 (N10045, N9997, N6872, N7020, N5546);
or OR4 (N10046, N10034, N372, N6746, N1859);
or OR2 (N10047, N10032, N6270);
not NOT1 (N10048, N10031);
and AND2 (N10049, N10044, N9351);
nor NOR3 (N10050, N10036, N9978, N513);
and AND2 (N10051, N10049, N5865);
not NOT1 (N10052, N10038);
xor XOR2 (N10053, N10050, N5052);
xor XOR2 (N10054, N10053, N8246);
not NOT1 (N10055, N10046);
and AND2 (N10056, N10042, N9576);
xor XOR2 (N10057, N10055, N2103);
buf BUF1 (N10058, N10047);
and AND2 (N10059, N10054, N9189);
or OR4 (N10060, N10048, N1451, N6, N9428);
nor NOR3 (N10061, N10060, N9681, N5188);
nor NOR3 (N10062, N10057, N5217, N2659);
or OR3 (N10063, N10056, N6086, N2534);
and AND3 (N10064, N10052, N8199, N8832);
nand NAND3 (N10065, N10063, N3155, N5313);
buf BUF1 (N10066, N10061);
buf BUF1 (N10067, N10064);
xor XOR2 (N10068, N10051, N9271);
not NOT1 (N10069, N10066);
and AND4 (N10070, N10045, N4379, N8374, N5071);
xor XOR2 (N10071, N10041, N2596);
nand NAND4 (N10072, N10062, N3497, N6414, N7690);
xor XOR2 (N10073, N10068, N7924);
nand NAND2 (N10074, N10065, N4936);
buf BUF1 (N10075, N10073);
buf BUF1 (N10076, N10070);
not NOT1 (N10077, N10075);
not NOT1 (N10078, N10067);
nor NOR4 (N10079, N10037, N6533, N9792, N9323);
or OR3 (N10080, N10078, N7766, N5448);
xor XOR2 (N10081, N10072, N5757);
nand NAND3 (N10082, N10079, N4668, N3924);
buf BUF1 (N10083, N10082);
buf BUF1 (N10084, N10058);
nor NOR4 (N10085, N10077, N3299, N948, N2742);
and AND4 (N10086, N10084, N1638, N302, N7509);
nand NAND2 (N10087, N10059, N5227);
nor NOR4 (N10088, N10087, N10061, N8832, N8948);
not NOT1 (N10089, N10076);
and AND2 (N10090, N10086, N8123);
and AND3 (N10091, N10074, N7709, N2724);
not NOT1 (N10092, N10071);
not NOT1 (N10093, N10089);
buf BUF1 (N10094, N10083);
not NOT1 (N10095, N10093);
nand NAND3 (N10096, N10069, N8729, N1841);
not NOT1 (N10097, N10092);
and AND4 (N10098, N10080, N6129, N409, N9323);
nor NOR4 (N10099, N10096, N8100, N3287, N7622);
nor NOR2 (N10100, N10091, N6786);
nor NOR4 (N10101, N10094, N7299, N9920, N958);
or OR2 (N10102, N10097, N6596);
nand NAND3 (N10103, N10101, N5116, N4707);
nand NAND2 (N10104, N10095, N4685);
xor XOR2 (N10105, N10085, N880);
nand NAND4 (N10106, N10090, N6496, N2020, N8281);
buf BUF1 (N10107, N10104);
buf BUF1 (N10108, N10099);
xor XOR2 (N10109, N10098, N7221);
xor XOR2 (N10110, N10081, N4655);
buf BUF1 (N10111, N10109);
xor XOR2 (N10112, N10107, N9013);
buf BUF1 (N10113, N10100);
nand NAND2 (N10114, N10111, N4018);
nor NOR4 (N10115, N10112, N4807, N3212, N3947);
not NOT1 (N10116, N10110);
nand NAND4 (N10117, N10105, N6919, N7133, N4488);
nand NAND3 (N10118, N10115, N5969, N828);
nor NOR3 (N10119, N10113, N6491, N3716);
not NOT1 (N10120, N10116);
nand NAND3 (N10121, N10120, N4643, N871);
nor NOR3 (N10122, N10118, N6378, N3708);
or OR4 (N10123, N10103, N4597, N8205, N3814);
xor XOR2 (N10124, N10123, N5303);
buf BUF1 (N10125, N10124);
and AND4 (N10126, N10125, N5993, N3050, N7449);
nor NOR3 (N10127, N10106, N7016, N6605);
nand NAND4 (N10128, N10127, N9706, N8373, N9841);
or OR4 (N10129, N10117, N9230, N51, N7793);
or OR4 (N10130, N10122, N5742, N3247, N8814);
and AND4 (N10131, N10129, N6476, N8171, N1904);
nor NOR2 (N10132, N10114, N6648);
nor NOR4 (N10133, N10119, N8570, N1443, N3179);
not NOT1 (N10134, N10130);
or OR2 (N10135, N10102, N3671);
nor NOR2 (N10136, N10128, N4030);
or OR3 (N10137, N10134, N7428, N623);
nand NAND4 (N10138, N10137, N9132, N2182, N3669);
and AND4 (N10139, N10121, N935, N5860, N9293);
nand NAND3 (N10140, N10126, N6078, N2182);
xor XOR2 (N10141, N10138, N3347);
buf BUF1 (N10142, N10108);
xor XOR2 (N10143, N10132, N5096);
or OR3 (N10144, N10088, N21, N6928);
xor XOR2 (N10145, N10144, N8225);
xor XOR2 (N10146, N10139, N4142);
or OR2 (N10147, N10141, N3771);
or OR4 (N10148, N10147, N6867, N38, N4115);
nand NAND3 (N10149, N10136, N4125, N6232);
nand NAND2 (N10150, N10148, N990);
nor NOR4 (N10151, N10142, N9132, N6460, N6393);
nor NOR4 (N10152, N10131, N5346, N4001, N9117);
or OR3 (N10153, N10140, N9323, N3367);
nand NAND3 (N10154, N10133, N3919, N4989);
not NOT1 (N10155, N10150);
not NOT1 (N10156, N10152);
nand NAND4 (N10157, N10151, N9662, N4597, N3207);
nor NOR3 (N10158, N10154, N7838, N4865);
nor NOR3 (N10159, N10143, N7047, N4259);
and AND3 (N10160, N10153, N5725, N253);
xor XOR2 (N10161, N10135, N8681);
not NOT1 (N10162, N10157);
and AND2 (N10163, N10161, N8458);
xor XOR2 (N10164, N10149, N249);
buf BUF1 (N10165, N10158);
xor XOR2 (N10166, N10164, N593);
not NOT1 (N10167, N10156);
xor XOR2 (N10168, N10165, N5121);
or OR4 (N10169, N10163, N10034, N6069, N4780);
nor NOR2 (N10170, N10146, N3424);
xor XOR2 (N10171, N10167, N8169);
buf BUF1 (N10172, N10159);
not NOT1 (N10173, N10145);
or OR3 (N10174, N10168, N6826, N7186);
not NOT1 (N10175, N10166);
nand NAND3 (N10176, N10175, N5559, N1318);
nor NOR3 (N10177, N10160, N4866, N2880);
nand NAND2 (N10178, N10169, N34);
or OR4 (N10179, N10155, N9640, N7688, N9945);
xor XOR2 (N10180, N10177, N3858);
nand NAND4 (N10181, N10173, N5179, N3475, N3857);
not NOT1 (N10182, N10179);
nand NAND4 (N10183, N10170, N6302, N683, N6346);
not NOT1 (N10184, N10181);
buf BUF1 (N10185, N10174);
nand NAND4 (N10186, N10182, N1771, N9124, N6505);
not NOT1 (N10187, N10162);
or OR2 (N10188, N10186, N3039);
or OR2 (N10189, N10176, N10042);
buf BUF1 (N10190, N10172);
or OR4 (N10191, N10190, N9416, N3616, N85);
and AND4 (N10192, N10185, N10055, N5469, N7853);
and AND2 (N10193, N10188, N8543);
and AND3 (N10194, N10183, N3005, N6946);
not NOT1 (N10195, N10193);
nand NAND4 (N10196, N10187, N563, N2723, N8207);
not NOT1 (N10197, N10191);
xor XOR2 (N10198, N10196, N9631);
and AND2 (N10199, N10194, N772);
nor NOR4 (N10200, N10189, N1320, N9035, N5714);
and AND2 (N10201, N10195, N6834);
nor NOR4 (N10202, N10198, N1044, N5485, N6182);
nor NOR4 (N10203, N10171, N7784, N4583, N5245);
or OR2 (N10204, N10178, N1737);
and AND3 (N10205, N10202, N5454, N10192);
nand NAND2 (N10206, N6670, N7714);
xor XOR2 (N10207, N10180, N9862);
nand NAND2 (N10208, N10205, N3074);
buf BUF1 (N10209, N10184);
and AND4 (N10210, N10199, N2289, N5897, N9290);
nor NOR3 (N10211, N10203, N5879, N7311);
not NOT1 (N10212, N10208);
nor NOR4 (N10213, N10212, N3184, N7945, N3948);
nor NOR2 (N10214, N10201, N5431);
or OR4 (N10215, N10204, N8881, N9532, N6651);
nand NAND3 (N10216, N10213, N6450, N8317);
nand NAND3 (N10217, N10215, N1016, N9578);
nor NOR4 (N10218, N10206, N5802, N3302, N6464);
not NOT1 (N10219, N10197);
nor NOR2 (N10220, N10217, N3480);
not NOT1 (N10221, N10214);
or OR3 (N10222, N10218, N2210, N4677);
and AND2 (N10223, N10222, N7893);
not NOT1 (N10224, N10223);
nor NOR2 (N10225, N10224, N6109);
or OR2 (N10226, N10207, N3334);
buf BUF1 (N10227, N10221);
or OR3 (N10228, N10227, N710, N10123);
nor NOR3 (N10229, N10209, N589, N3065);
nand NAND2 (N10230, N10200, N766);
and AND4 (N10231, N10211, N6959, N215, N5642);
nand NAND4 (N10232, N10230, N3315, N2604, N341);
not NOT1 (N10233, N10220);
nand NAND3 (N10234, N10225, N9780, N4087);
not NOT1 (N10235, N10232);
buf BUF1 (N10236, N10233);
buf BUF1 (N10237, N10231);
buf BUF1 (N10238, N10235);
and AND2 (N10239, N10236, N8153);
nand NAND3 (N10240, N10229, N7863, N3859);
nand NAND2 (N10241, N10239, N8206);
nand NAND4 (N10242, N10228, N4756, N4764, N2448);
nor NOR3 (N10243, N10241, N6731, N4330);
and AND3 (N10244, N10240, N3058, N2745);
xor XOR2 (N10245, N10234, N1373);
nand NAND4 (N10246, N10243, N1897, N5071, N2892);
or OR2 (N10247, N10216, N739);
not NOT1 (N10248, N10242);
or OR2 (N10249, N10248, N3172);
buf BUF1 (N10250, N10238);
nand NAND4 (N10251, N10210, N5440, N1980, N6928);
and AND4 (N10252, N10251, N9101, N4596, N8035);
or OR2 (N10253, N10249, N10192);
not NOT1 (N10254, N10237);
xor XOR2 (N10255, N10246, N6607);
xor XOR2 (N10256, N10253, N3188);
buf BUF1 (N10257, N10219);
or OR3 (N10258, N10244, N3410, N3207);
or OR4 (N10259, N10254, N9966, N3902, N1843);
or OR4 (N10260, N10247, N611, N8363, N4696);
or OR4 (N10261, N10250, N7887, N4716, N493);
and AND2 (N10262, N10258, N1025);
not NOT1 (N10263, N10257);
and AND3 (N10264, N10259, N60, N1213);
and AND2 (N10265, N10260, N7571);
xor XOR2 (N10266, N10245, N4304);
xor XOR2 (N10267, N10264, N4854);
or OR3 (N10268, N10252, N3570, N9453);
not NOT1 (N10269, N10261);
and AND3 (N10270, N10267, N3115, N8388);
buf BUF1 (N10271, N10255);
nor NOR4 (N10272, N10263, N25, N1973, N3823);
nor NOR2 (N10273, N10265, N6952);
buf BUF1 (N10274, N10256);
or OR4 (N10275, N10262, N2788, N8856, N7514);
nor NOR4 (N10276, N10273, N5642, N10076, N3933);
nor NOR3 (N10277, N10272, N10019, N40);
nor NOR4 (N10278, N10277, N1127, N10088, N1320);
or OR4 (N10279, N10271, N3338, N3021, N8859);
buf BUF1 (N10280, N10268);
nand NAND2 (N10281, N10274, N554);
buf BUF1 (N10282, N10269);
xor XOR2 (N10283, N10278, N6612);
nor NOR4 (N10284, N10270, N1507, N636, N3929);
not NOT1 (N10285, N10266);
buf BUF1 (N10286, N10282);
not NOT1 (N10287, N10285);
nand NAND3 (N10288, N10280, N9732, N6059);
xor XOR2 (N10289, N10287, N4805);
nor NOR3 (N10290, N10283, N1788, N7072);
not NOT1 (N10291, N10276);
or OR3 (N10292, N10279, N7667, N3104);
and AND3 (N10293, N10290, N9136, N3148);
and AND3 (N10294, N10281, N6102, N4824);
and AND3 (N10295, N10284, N1061, N7738);
and AND4 (N10296, N10286, N1395, N8558, N1316);
not NOT1 (N10297, N10292);
nand NAND2 (N10298, N10297, N7439);
nand NAND4 (N10299, N10293, N1148, N2451, N8383);
xor XOR2 (N10300, N10294, N7497);
buf BUF1 (N10301, N10298);
not NOT1 (N10302, N10226);
nand NAND2 (N10303, N10275, N1627);
nand NAND2 (N10304, N10301, N1454);
nand NAND2 (N10305, N10299, N6766);
xor XOR2 (N10306, N10305, N444);
or OR4 (N10307, N10288, N2576, N4555, N7203);
and AND3 (N10308, N10302, N5746, N723);
nand NAND3 (N10309, N10289, N1985, N1673);
buf BUF1 (N10310, N10307);
not NOT1 (N10311, N10310);
nor NOR2 (N10312, N10311, N7831);
nor NOR4 (N10313, N10291, N9550, N2020, N4574);
buf BUF1 (N10314, N10296);
not NOT1 (N10315, N10314);
xor XOR2 (N10316, N10306, N8867);
and AND2 (N10317, N10303, N6049);
xor XOR2 (N10318, N10312, N6937);
and AND4 (N10319, N10318, N4132, N8571, N1710);
buf BUF1 (N10320, N10308);
nor NOR4 (N10321, N10319, N9153, N6643, N8837);
nand NAND2 (N10322, N10315, N650);
buf BUF1 (N10323, N10320);
nor NOR3 (N10324, N10321, N10162, N1096);
not NOT1 (N10325, N10300);
buf BUF1 (N10326, N10323);
buf BUF1 (N10327, N10316);
nor NOR4 (N10328, N10322, N618, N4579, N1799);
xor XOR2 (N10329, N10325, N9916);
or OR4 (N10330, N10317, N3911, N4308, N6510);
not NOT1 (N10331, N10328);
nand NAND2 (N10332, N10304, N226);
nor NOR4 (N10333, N10330, N701, N8284, N453);
buf BUF1 (N10334, N10329);
not NOT1 (N10335, N10334);
nor NOR4 (N10336, N10332, N6494, N4312, N7390);
or OR4 (N10337, N10327, N184, N3796, N5184);
xor XOR2 (N10338, N10295, N5253);
not NOT1 (N10339, N10333);
nor NOR3 (N10340, N10324, N6563, N9435);
nor NOR4 (N10341, N10331, N2651, N5334, N429);
or OR2 (N10342, N10337, N2449);
xor XOR2 (N10343, N10341, N9440);
not NOT1 (N10344, N10336);
buf BUF1 (N10345, N10340);
xor XOR2 (N10346, N10344, N3400);
and AND4 (N10347, N10313, N8534, N6433, N7941);
not NOT1 (N10348, N10346);
buf BUF1 (N10349, N10335);
not NOT1 (N10350, N10339);
xor XOR2 (N10351, N10350, N5571);
or OR3 (N10352, N10345, N3924, N4544);
buf BUF1 (N10353, N10347);
nor NOR2 (N10354, N10352, N5952);
nand NAND3 (N10355, N10342, N4134, N9327);
buf BUF1 (N10356, N10343);
or OR4 (N10357, N10326, N7236, N7168, N7924);
and AND2 (N10358, N10348, N6681);
nand NAND3 (N10359, N10358, N3834, N9878);
nor NOR4 (N10360, N10349, N6263, N4666, N7165);
not NOT1 (N10361, N10360);
buf BUF1 (N10362, N10357);
nand NAND4 (N10363, N10351, N7441, N9586, N9597);
nor NOR4 (N10364, N10354, N4940, N2769, N2796);
and AND3 (N10365, N10338, N4385, N3149);
nand NAND4 (N10366, N10359, N632, N8615, N4880);
xor XOR2 (N10367, N10309, N5704);
and AND4 (N10368, N10356, N1950, N2435, N7669);
nor NOR4 (N10369, N10367, N9137, N9592, N4245);
and AND3 (N10370, N10364, N3014, N3168);
and AND3 (N10371, N10362, N3683, N142);
nor NOR3 (N10372, N10353, N1645, N218);
nand NAND3 (N10373, N10363, N4105, N3423);
or OR2 (N10374, N10368, N4550);
or OR3 (N10375, N10373, N2384, N1738);
or OR4 (N10376, N10355, N6206, N7287, N2312);
or OR2 (N10377, N10371, N7330);
nand NAND4 (N10378, N10377, N5944, N9424, N2405);
buf BUF1 (N10379, N10361);
and AND2 (N10380, N10376, N1926);
not NOT1 (N10381, N10372);
and AND4 (N10382, N10366, N1360, N4220, N7864);
nand NAND4 (N10383, N10374, N4976, N4996, N6531);
nor NOR3 (N10384, N10383, N6093, N7761);
xor XOR2 (N10385, N10375, N1272);
nor NOR3 (N10386, N10381, N3170, N8226);
nand NAND2 (N10387, N10386, N8097);
not NOT1 (N10388, N10380);
or OR3 (N10389, N10370, N7451, N6552);
nand NAND4 (N10390, N10389, N4330, N4779, N8741);
or OR3 (N10391, N10378, N7836, N3883);
xor XOR2 (N10392, N10388, N5410);
xor XOR2 (N10393, N10365, N6);
xor XOR2 (N10394, N10392, N1116);
or OR3 (N10395, N10391, N6292, N9908);
or OR4 (N10396, N10390, N3117, N815, N2264);
buf BUF1 (N10397, N10369);
nand NAND2 (N10398, N10397, N740);
xor XOR2 (N10399, N10398, N3948);
xor XOR2 (N10400, N10387, N9295);
not NOT1 (N10401, N10385);
xor XOR2 (N10402, N10399, N9777);
or OR2 (N10403, N10401, N7722);
nand NAND4 (N10404, N10384, N517, N303, N4198);
nor NOR3 (N10405, N10404, N5118, N3018);
not NOT1 (N10406, N10393);
and AND2 (N10407, N10403, N841);
buf BUF1 (N10408, N10394);
not NOT1 (N10409, N10400);
buf BUF1 (N10410, N10382);
xor XOR2 (N10411, N10406, N4095);
or OR4 (N10412, N10379, N5417, N5177, N8856);
nor NOR2 (N10413, N10395, N9157);
or OR2 (N10414, N10411, N650);
not NOT1 (N10415, N10409);
nor NOR2 (N10416, N10405, N5132);
or OR4 (N10417, N10402, N9501, N5910, N3841);
not NOT1 (N10418, N10414);
buf BUF1 (N10419, N10407);
nand NAND4 (N10420, N10419, N3942, N4788, N7033);
xor XOR2 (N10421, N10410, N3515);
and AND2 (N10422, N10418, N8402);
and AND3 (N10423, N10412, N9445, N6865);
or OR4 (N10424, N10423, N7221, N8531, N7903);
nor NOR3 (N10425, N10422, N4950, N4940);
xor XOR2 (N10426, N10421, N4545);
and AND2 (N10427, N10408, N5598);
nand NAND2 (N10428, N10416, N6616);
xor XOR2 (N10429, N10415, N7708);
buf BUF1 (N10430, N10424);
buf BUF1 (N10431, N10426);
not NOT1 (N10432, N10431);
and AND4 (N10433, N10428, N6190, N8294, N6447);
not NOT1 (N10434, N10430);
and AND3 (N10435, N10396, N10002, N2035);
and AND3 (N10436, N10433, N5904, N9968);
and AND3 (N10437, N10434, N7965, N3586);
not NOT1 (N10438, N10413);
nand NAND2 (N10439, N10420, N8339);
xor XOR2 (N10440, N10429, N5755);
buf BUF1 (N10441, N10437);
nor NOR2 (N10442, N10439, N3048);
buf BUF1 (N10443, N10425);
nand NAND3 (N10444, N10443, N10189, N7112);
and AND3 (N10445, N10427, N8770, N7537);
buf BUF1 (N10446, N10435);
and AND3 (N10447, N10446, N1336, N5639);
or OR4 (N10448, N10442, N10032, N10267, N2857);
buf BUF1 (N10449, N10432);
and AND4 (N10450, N10417, N4830, N6191, N4257);
nor NOR2 (N10451, N10448, N1095);
nand NAND4 (N10452, N10436, N6445, N609, N2680);
not NOT1 (N10453, N10452);
nor NOR2 (N10454, N10447, N5492);
xor XOR2 (N10455, N10450, N6318);
or OR2 (N10456, N10455, N1884);
nor NOR4 (N10457, N10445, N6524, N5312, N3731);
xor XOR2 (N10458, N10444, N10413);
xor XOR2 (N10459, N10451, N4642);
xor XOR2 (N10460, N10449, N3721);
nand NAND4 (N10461, N10457, N10186, N6254, N2336);
buf BUF1 (N10462, N10453);
not NOT1 (N10463, N10458);
xor XOR2 (N10464, N10441, N3565);
or OR2 (N10465, N10454, N5694);
nand NAND2 (N10466, N10463, N5112);
and AND2 (N10467, N10466, N6480);
buf BUF1 (N10468, N10464);
nand NAND4 (N10469, N10461, N558, N569, N1757);
or OR4 (N10470, N10460, N8738, N48, N6305);
nor NOR3 (N10471, N10467, N972, N7881);
xor XOR2 (N10472, N10465, N3680);
xor XOR2 (N10473, N10470, N5425);
and AND3 (N10474, N10472, N8863, N8340);
not NOT1 (N10475, N10473);
nor NOR2 (N10476, N10462, N1587);
nand NAND4 (N10477, N10459, N2519, N2952, N7476);
nor NOR3 (N10478, N10469, N10240, N8716);
nor NOR2 (N10479, N10438, N8070);
or OR2 (N10480, N10471, N397);
buf BUF1 (N10481, N10476);
buf BUF1 (N10482, N10440);
nor NOR3 (N10483, N10468, N1750, N3530);
buf BUF1 (N10484, N10478);
nand NAND3 (N10485, N10475, N4853, N6525);
or OR2 (N10486, N10477, N5817);
nor NOR4 (N10487, N10479, N2963, N8582, N2157);
not NOT1 (N10488, N10484);
buf BUF1 (N10489, N10481);
buf BUF1 (N10490, N10485);
xor XOR2 (N10491, N10474, N4701);
xor XOR2 (N10492, N10456, N2798);
and AND4 (N10493, N10491, N9917, N3043, N7490);
not NOT1 (N10494, N10480);
not NOT1 (N10495, N10490);
or OR3 (N10496, N10483, N6293, N6372);
and AND2 (N10497, N10496, N5371);
not NOT1 (N10498, N10486);
xor XOR2 (N10499, N10482, N6198);
nor NOR2 (N10500, N10499, N2676);
not NOT1 (N10501, N10497);
nor NOR2 (N10502, N10493, N8620);
nand NAND2 (N10503, N10500, N5908);
nor NOR2 (N10504, N10492, N6601);
and AND2 (N10505, N10488, N2089);
not NOT1 (N10506, N10505);
xor XOR2 (N10507, N10502, N3982);
nor NOR3 (N10508, N10489, N4038, N2482);
or OR4 (N10509, N10503, N9193, N298, N1346);
not NOT1 (N10510, N10504);
or OR2 (N10511, N10495, N7530);
buf BUF1 (N10512, N10509);
buf BUF1 (N10513, N10494);
nor NOR4 (N10514, N10487, N5985, N4964, N4086);
xor XOR2 (N10515, N10511, N1958);
nor NOR3 (N10516, N10507, N1980, N5920);
not NOT1 (N10517, N10510);
and AND3 (N10518, N10517, N3343, N6212);
not NOT1 (N10519, N10506);
buf BUF1 (N10520, N10519);
xor XOR2 (N10521, N10516, N5874);
nand NAND3 (N10522, N10508, N8199, N8326);
or OR3 (N10523, N10515, N5590, N3049);
buf BUF1 (N10524, N10513);
nand NAND3 (N10525, N10514, N4352, N6067);
and AND3 (N10526, N10512, N10316, N5419);
nand NAND4 (N10527, N10522, N7477, N10032, N7284);
or OR3 (N10528, N10521, N1391, N10057);
buf BUF1 (N10529, N10520);
and AND2 (N10530, N10498, N3244);
nand NAND3 (N10531, N10528, N8516, N935);
buf BUF1 (N10532, N10526);
nand NAND3 (N10533, N10529, N4758, N10142);
buf BUF1 (N10534, N10518);
nor NOR3 (N10535, N10532, N2231, N7474);
xor XOR2 (N10536, N10525, N4386);
buf BUF1 (N10537, N10523);
and AND3 (N10538, N10536, N5864, N4334);
nand NAND3 (N10539, N10524, N8246, N6260);
and AND3 (N10540, N10539, N7277, N3093);
not NOT1 (N10541, N10538);
not NOT1 (N10542, N10541);
or OR3 (N10543, N10540, N3889, N9274);
nor NOR4 (N10544, N10501, N6839, N959, N1023);
nand NAND4 (N10545, N10544, N2427, N9069, N3836);
nand NAND3 (N10546, N10543, N4359, N334);
xor XOR2 (N10547, N10531, N1395);
nand NAND4 (N10548, N10547, N2817, N2572, N6427);
and AND3 (N10549, N10534, N6378, N6824);
not NOT1 (N10550, N10527);
nor NOR4 (N10551, N10535, N3879, N5174, N6411);
buf BUF1 (N10552, N10551);
not NOT1 (N10553, N10552);
and AND3 (N10554, N10537, N6528, N5296);
buf BUF1 (N10555, N10546);
not NOT1 (N10556, N10553);
buf BUF1 (N10557, N10554);
or OR2 (N10558, N10555, N8752);
nand NAND2 (N10559, N10542, N249);
nand NAND3 (N10560, N10548, N3452, N4015);
buf BUF1 (N10561, N10556);
not NOT1 (N10562, N10557);
and AND2 (N10563, N10559, N2811);
buf BUF1 (N10564, N10549);
buf BUF1 (N10565, N10530);
not NOT1 (N10566, N10565);
xor XOR2 (N10567, N10564, N9826);
or OR3 (N10568, N10550, N5652, N8953);
xor XOR2 (N10569, N10567, N9830);
nand NAND2 (N10570, N10568, N6155);
or OR4 (N10571, N10570, N7805, N2485, N4902);
nor NOR3 (N10572, N10562, N1578, N1264);
and AND3 (N10573, N10566, N1697, N9461);
or OR4 (N10574, N10560, N10013, N3278, N3862);
xor XOR2 (N10575, N10558, N7391);
or OR4 (N10576, N10545, N4795, N9822, N2320);
nor NOR4 (N10577, N10575, N5402, N8687, N9448);
and AND4 (N10578, N10574, N9540, N233, N3950);
xor XOR2 (N10579, N10576, N2841);
nor NOR3 (N10580, N10572, N7090, N3882);
nand NAND3 (N10581, N10563, N7870, N3876);
buf BUF1 (N10582, N10579);
xor XOR2 (N10583, N10580, N5001);
and AND4 (N10584, N10571, N9139, N3646, N8910);
xor XOR2 (N10585, N10561, N6749);
not NOT1 (N10586, N10578);
xor XOR2 (N10587, N10584, N10379);
xor XOR2 (N10588, N10581, N331);
nor NOR2 (N10589, N10587, N3634);
not NOT1 (N10590, N10569);
buf BUF1 (N10591, N10589);
and AND2 (N10592, N10573, N6865);
nand NAND2 (N10593, N10582, N2168);
or OR3 (N10594, N10585, N1021, N10478);
nand NAND2 (N10595, N10591, N392);
and AND3 (N10596, N10583, N8502, N8682);
nor NOR4 (N10597, N10596, N1754, N5555, N8132);
buf BUF1 (N10598, N10588);
nor NOR3 (N10599, N10592, N4225, N472);
buf BUF1 (N10600, N10586);
and AND3 (N10601, N10593, N8034, N4981);
nand NAND2 (N10602, N10597, N361);
or OR3 (N10603, N10533, N2650, N1494);
nand NAND4 (N10604, N10599, N9092, N8196, N9224);
nand NAND3 (N10605, N10595, N1359, N2845);
nand NAND3 (N10606, N10605, N3554, N3971);
and AND4 (N10607, N10594, N3300, N4657, N801);
nor NOR3 (N10608, N10604, N7907, N5489);
nor NOR4 (N10609, N10598, N628, N10118, N3333);
buf BUF1 (N10610, N10609);
not NOT1 (N10611, N10608);
and AND2 (N10612, N10600, N3287);
and AND2 (N10613, N10602, N3856);
and AND3 (N10614, N10611, N6873, N8088);
and AND4 (N10615, N10601, N7246, N6453, N834);
xor XOR2 (N10616, N10612, N2935);
buf BUF1 (N10617, N10614);
nor NOR2 (N10618, N10606, N5086);
not NOT1 (N10619, N10603);
nand NAND4 (N10620, N10610, N3820, N7691, N9060);
xor XOR2 (N10621, N10620, N7952);
buf BUF1 (N10622, N10577);
not NOT1 (N10623, N10622);
nor NOR4 (N10624, N10615, N9845, N7706, N3788);
nor NOR3 (N10625, N10624, N2712, N485);
not NOT1 (N10626, N10619);
nor NOR2 (N10627, N10616, N2448);
or OR4 (N10628, N10607, N5486, N8384, N3921);
and AND4 (N10629, N10621, N5361, N7522, N7573);
buf BUF1 (N10630, N10618);
nor NOR3 (N10631, N10617, N9105, N1799);
or OR3 (N10632, N10627, N4911, N3189);
xor XOR2 (N10633, N10625, N2293);
nor NOR2 (N10634, N10613, N2857);
xor XOR2 (N10635, N10626, N8922);
xor XOR2 (N10636, N10623, N6598);
nor NOR3 (N10637, N10635, N3504, N3370);
nor NOR4 (N10638, N10636, N7121, N4700, N3713);
not NOT1 (N10639, N10638);
xor XOR2 (N10640, N10634, N278);
xor XOR2 (N10641, N10628, N5202);
nor NOR4 (N10642, N10632, N711, N2388, N761);
nor NOR4 (N10643, N10641, N6683, N8559, N6652);
nor NOR2 (N10644, N10629, N3457);
xor XOR2 (N10645, N10630, N3574);
not NOT1 (N10646, N10642);
xor XOR2 (N10647, N10646, N9665);
or OR3 (N10648, N10647, N5371, N4551);
nand NAND4 (N10649, N10640, N10529, N798, N3942);
xor XOR2 (N10650, N10649, N431);
or OR3 (N10651, N10639, N2886, N638);
buf BUF1 (N10652, N10643);
and AND2 (N10653, N10633, N3906);
not NOT1 (N10654, N10651);
not NOT1 (N10655, N10654);
xor XOR2 (N10656, N10653, N9234);
and AND3 (N10657, N10637, N9634, N2449);
and AND3 (N10658, N10631, N8840, N4934);
not NOT1 (N10659, N10655);
and AND3 (N10660, N10644, N1632, N4081);
nor NOR4 (N10661, N10659, N10389, N3689, N9351);
not NOT1 (N10662, N10656);
and AND2 (N10663, N10650, N9841);
or OR4 (N10664, N10660, N5475, N1475, N5032);
nor NOR4 (N10665, N10661, N1501, N2491, N3880);
nor NOR2 (N10666, N10648, N1443);
nor NOR4 (N10667, N10657, N2968, N9531, N9252);
nor NOR4 (N10668, N10645, N8397, N1556, N4225);
or OR4 (N10669, N10662, N3398, N4860, N2157);
nor NOR2 (N10670, N10658, N9997);
not NOT1 (N10671, N10668);
and AND2 (N10672, N10663, N5885);
not NOT1 (N10673, N10671);
buf BUF1 (N10674, N10664);
nor NOR2 (N10675, N10665, N6681);
and AND4 (N10676, N10669, N990, N7305, N7471);
nor NOR3 (N10677, N10590, N9237, N7971);
buf BUF1 (N10678, N10666);
buf BUF1 (N10679, N10670);
xor XOR2 (N10680, N10673, N6428);
buf BUF1 (N10681, N10675);
not NOT1 (N10682, N10667);
nor NOR2 (N10683, N10676, N3603);
not NOT1 (N10684, N10677);
nor NOR4 (N10685, N10678, N10223, N9725, N7580);
or OR2 (N10686, N10680, N2281);
buf BUF1 (N10687, N10684);
buf BUF1 (N10688, N10686);
and AND4 (N10689, N10683, N8723, N4415, N9279);
nand NAND2 (N10690, N10689, N1161);
nor NOR3 (N10691, N10674, N5122, N737);
buf BUF1 (N10692, N10679);
xor XOR2 (N10693, N10691, N1424);
xor XOR2 (N10694, N10682, N2900);
nand NAND4 (N10695, N10681, N1115, N8914, N9017);
and AND3 (N10696, N10693, N6500, N7347);
nand NAND4 (N10697, N10672, N6496, N8644, N2942);
nand NAND2 (N10698, N10687, N8253);
or OR2 (N10699, N10692, N7557);
or OR3 (N10700, N10697, N42, N3928);
xor XOR2 (N10701, N10694, N4225);
not NOT1 (N10702, N10690);
buf BUF1 (N10703, N10702);
and AND3 (N10704, N10652, N10549, N8307);
not NOT1 (N10705, N10700);
and AND2 (N10706, N10703, N140);
buf BUF1 (N10707, N10698);
nand NAND2 (N10708, N10706, N411);
nor NOR3 (N10709, N10696, N1152, N10616);
not NOT1 (N10710, N10695);
not NOT1 (N10711, N10699);
xor XOR2 (N10712, N10688, N477);
buf BUF1 (N10713, N10712);
or OR2 (N10714, N10710, N5514);
nand NAND2 (N10715, N10685, N1644);
and AND2 (N10716, N10715, N7047);
xor XOR2 (N10717, N10714, N7808);
and AND2 (N10718, N10708, N541);
buf BUF1 (N10719, N10716);
and AND2 (N10720, N10717, N6452);
or OR3 (N10721, N10707, N723, N3379);
xor XOR2 (N10722, N10705, N1330);
xor XOR2 (N10723, N10704, N4726);
or OR2 (N10724, N10720, N3768);
nor NOR4 (N10725, N10711, N3128, N10640, N7971);
not NOT1 (N10726, N10719);
nand NAND2 (N10727, N10718, N6488);
or OR2 (N10728, N10727, N7059);
or OR3 (N10729, N10721, N2523, N3860);
nor NOR3 (N10730, N10722, N6487, N8391);
xor XOR2 (N10731, N10724, N706);
nor NOR2 (N10732, N10728, N5656);
nor NOR2 (N10733, N10725, N3385);
xor XOR2 (N10734, N10709, N8565);
nor NOR3 (N10735, N10733, N7109, N431);
nor NOR4 (N10736, N10713, N1359, N6773, N4461);
xor XOR2 (N10737, N10731, N503);
xor XOR2 (N10738, N10730, N456);
and AND3 (N10739, N10732, N9259, N8143);
nor NOR4 (N10740, N10738, N9459, N7219, N6956);
buf BUF1 (N10741, N10701);
xor XOR2 (N10742, N10741, N9293);
and AND3 (N10743, N10734, N4920, N3887);
and AND3 (N10744, N10729, N5011, N3241);
not NOT1 (N10745, N10726);
nand NAND4 (N10746, N10743, N8136, N9957, N3985);
buf BUF1 (N10747, N10740);
nor NOR4 (N10748, N10736, N9492, N8579, N4744);
nand NAND2 (N10749, N10739, N2294);
nand NAND2 (N10750, N10723, N7725);
and AND4 (N10751, N10742, N2405, N260, N2415);
not NOT1 (N10752, N10749);
or OR2 (N10753, N10737, N6754);
and AND2 (N10754, N10752, N6698);
xor XOR2 (N10755, N10746, N3342);
and AND4 (N10756, N10753, N5594, N8514, N10415);
xor XOR2 (N10757, N10755, N10572);
nand NAND3 (N10758, N10757, N9617, N10551);
and AND2 (N10759, N10750, N9856);
xor XOR2 (N10760, N10747, N4121);
or OR4 (N10761, N10745, N2478, N3465, N690);
and AND3 (N10762, N10758, N4430, N4180);
or OR4 (N10763, N10762, N4038, N5803, N9133);
nor NOR3 (N10764, N10763, N3649, N6425);
or OR4 (N10765, N10748, N5458, N10094, N6700);
nor NOR4 (N10766, N10756, N9790, N8842, N5701);
and AND4 (N10767, N10754, N6614, N7572, N3751);
not NOT1 (N10768, N10765);
nor NOR3 (N10769, N10735, N228, N1555);
and AND4 (N10770, N10751, N9406, N9609, N8555);
and AND3 (N10771, N10770, N5750, N2611);
or OR4 (N10772, N10759, N3661, N10457, N3944);
and AND3 (N10773, N10769, N7121, N5737);
nand NAND4 (N10774, N10761, N7461, N4738, N10471);
and AND4 (N10775, N10767, N3031, N7257, N6890);
nor NOR2 (N10776, N10764, N10096);
not NOT1 (N10777, N10766);
nor NOR2 (N10778, N10772, N511);
xor XOR2 (N10779, N10744, N6162);
or OR2 (N10780, N10773, N6058);
or OR2 (N10781, N10771, N7334);
nor NOR4 (N10782, N10781, N1932, N9091, N8683);
not NOT1 (N10783, N10768);
not NOT1 (N10784, N10779);
and AND4 (N10785, N10774, N10245, N9505, N4001);
nand NAND2 (N10786, N10783, N3036);
buf BUF1 (N10787, N10760);
xor XOR2 (N10788, N10776, N4120);
and AND3 (N10789, N10786, N5676, N7646);
or OR4 (N10790, N10780, N6233, N2190, N341);
and AND4 (N10791, N10784, N7031, N974, N5075);
nor NOR2 (N10792, N10777, N2785);
buf BUF1 (N10793, N10785);
buf BUF1 (N10794, N10775);
or OR2 (N10795, N10787, N8152);
and AND3 (N10796, N10788, N4967, N1320);
nor NOR4 (N10797, N10778, N4561, N3958, N646);
and AND3 (N10798, N10791, N8099, N3419);
buf BUF1 (N10799, N10794);
xor XOR2 (N10800, N10792, N1364);
nand NAND4 (N10801, N10793, N8279, N8817, N7409);
not NOT1 (N10802, N10797);
and AND4 (N10803, N10800, N5244, N10079, N8825);
or OR4 (N10804, N10799, N9027, N2183, N587);
and AND3 (N10805, N10801, N2003, N10335);
and AND4 (N10806, N10782, N10645, N2367, N214);
nor NOR4 (N10807, N10790, N2847, N10556, N3434);
nor NOR4 (N10808, N10798, N10794, N2457, N5);
and AND2 (N10809, N10806, N1450);
and AND4 (N10810, N10803, N193, N3801, N892);
buf BUF1 (N10811, N10804);
and AND2 (N10812, N10789, N8326);
and AND2 (N10813, N10811, N2911);
not NOT1 (N10814, N10812);
not NOT1 (N10815, N10813);
nand NAND2 (N10816, N10814, N1317);
nand NAND4 (N10817, N10815, N9054, N10637, N2233);
nand NAND2 (N10818, N10805, N7557);
nand NAND3 (N10819, N10809, N6889, N10697);
or OR4 (N10820, N10819, N4649, N8020, N10431);
xor XOR2 (N10821, N10796, N7085);
nor NOR3 (N10822, N10808, N6628, N10814);
nor NOR4 (N10823, N10807, N6475, N10664, N8937);
or OR3 (N10824, N10817, N1632, N5121);
nand NAND4 (N10825, N10823, N4349, N10283, N2555);
nor NOR3 (N10826, N10795, N2123, N2472);
nor NOR2 (N10827, N10826, N5488);
or OR3 (N10828, N10816, N8402, N8642);
buf BUF1 (N10829, N10810);
and AND3 (N10830, N10827, N1174, N4613);
buf BUF1 (N10831, N10825);
nor NOR2 (N10832, N10830, N2203);
nor NOR3 (N10833, N10821, N2818, N2391);
not NOT1 (N10834, N10824);
xor XOR2 (N10835, N10833, N8983);
not NOT1 (N10836, N10828);
buf BUF1 (N10837, N10822);
and AND2 (N10838, N10820, N418);
buf BUF1 (N10839, N10837);
nor NOR3 (N10840, N10832, N5831, N7173);
xor XOR2 (N10841, N10840, N5353);
nor NOR4 (N10842, N10836, N9537, N3046, N3489);
nor NOR2 (N10843, N10802, N6595);
or OR4 (N10844, N10829, N293, N7891, N8280);
not NOT1 (N10845, N10839);
nand NAND2 (N10846, N10845, N10284);
nor NOR3 (N10847, N10843, N5, N8189);
nor NOR2 (N10848, N10831, N3046);
buf BUF1 (N10849, N10834);
nand NAND4 (N10850, N10838, N4832, N10357, N10057);
not NOT1 (N10851, N10846);
nand NAND4 (N10852, N10835, N8182, N5858, N6979);
xor XOR2 (N10853, N10847, N1924);
nand NAND3 (N10854, N10842, N2702, N304);
nand NAND2 (N10855, N10850, N4821);
nand NAND4 (N10856, N10851, N10590, N10703, N2365);
not NOT1 (N10857, N10853);
nor NOR2 (N10858, N10844, N1488);
not NOT1 (N10859, N10858);
nand NAND2 (N10860, N10857, N10573);
nor NOR4 (N10861, N10848, N4316, N5564, N9642);
or OR4 (N10862, N10841, N10134, N1051, N881);
and AND3 (N10863, N10856, N3933, N7474);
nor NOR2 (N10864, N10854, N2204);
not NOT1 (N10865, N10818);
buf BUF1 (N10866, N10855);
and AND3 (N10867, N10852, N7592, N5992);
nand NAND2 (N10868, N10860, N10045);
xor XOR2 (N10869, N10861, N2224);
and AND4 (N10870, N10862, N4899, N3636, N2393);
nand NAND3 (N10871, N10865, N3989, N3610);
and AND4 (N10872, N10870, N7253, N650, N639);
and AND2 (N10873, N10863, N6416);
not NOT1 (N10874, N10872);
xor XOR2 (N10875, N10869, N7811);
not NOT1 (N10876, N10864);
or OR4 (N10877, N10871, N4910, N4743, N9322);
xor XOR2 (N10878, N10875, N586);
xor XOR2 (N10879, N10866, N5831);
nor NOR4 (N10880, N10873, N9739, N9977, N4999);
xor XOR2 (N10881, N10879, N10149);
nor NOR3 (N10882, N10874, N5749, N5247);
or OR2 (N10883, N10876, N8493);
nand NAND2 (N10884, N10849, N2435);
and AND3 (N10885, N10884, N8862, N9172);
buf BUF1 (N10886, N10859);
not NOT1 (N10887, N10883);
or OR2 (N10888, N10868, N10379);
nor NOR4 (N10889, N10885, N1758, N5474, N8352);
buf BUF1 (N10890, N10881);
or OR4 (N10891, N10877, N6028, N1119, N7751);
buf BUF1 (N10892, N10886);
xor XOR2 (N10893, N10880, N1675);
buf BUF1 (N10894, N10878);
nand NAND3 (N10895, N10891, N4044, N9381);
nand NAND4 (N10896, N10882, N9523, N3237, N9109);
or OR4 (N10897, N10893, N2992, N865, N1196);
and AND3 (N10898, N10894, N2230, N6789);
nand NAND2 (N10899, N10867, N7006);
xor XOR2 (N10900, N10889, N7882);
nand NAND4 (N10901, N10887, N2458, N5743, N8351);
and AND2 (N10902, N10888, N2025);
or OR2 (N10903, N10900, N2922);
not NOT1 (N10904, N10902);
not NOT1 (N10905, N10899);
not NOT1 (N10906, N10896);
nand NAND4 (N10907, N10903, N8472, N5543, N2630);
not NOT1 (N10908, N10895);
and AND2 (N10909, N10908, N4723);
xor XOR2 (N10910, N10897, N4410);
buf BUF1 (N10911, N10898);
and AND2 (N10912, N10905, N9741);
or OR2 (N10913, N10892, N4983);
or OR4 (N10914, N10912, N979, N141, N2161);
and AND4 (N10915, N10890, N5199, N6455, N9019);
nor NOR2 (N10916, N10907, N5036);
and AND2 (N10917, N10906, N2076);
not NOT1 (N10918, N10911);
nor NOR3 (N10919, N10918, N3972, N3933);
and AND2 (N10920, N10915, N3168);
nor NOR4 (N10921, N10913, N6604, N8609, N1107);
and AND3 (N10922, N10909, N8677, N6771);
xor XOR2 (N10923, N10914, N3897);
or OR3 (N10924, N10921, N6838, N1949);
and AND4 (N10925, N10901, N438, N6409, N7314);
buf BUF1 (N10926, N10925);
nand NAND3 (N10927, N10922, N5769, N2098);
or OR2 (N10928, N10920, N10655);
nand NAND2 (N10929, N10916, N469);
or OR2 (N10930, N10917, N6861);
xor XOR2 (N10931, N10926, N1749);
and AND2 (N10932, N10910, N8350);
or OR4 (N10933, N10930, N8595, N8396, N4592);
buf BUF1 (N10934, N10924);
nor NOR3 (N10935, N10932, N412, N7058);
and AND3 (N10936, N10919, N8086, N3135);
xor XOR2 (N10937, N10931, N6336);
and AND4 (N10938, N10904, N4660, N2357, N6154);
or OR4 (N10939, N10935, N7889, N5685, N4486);
nand NAND2 (N10940, N10923, N6922);
nand NAND2 (N10941, N10934, N5946);
and AND3 (N10942, N10933, N8095, N9231);
buf BUF1 (N10943, N10936);
nand NAND4 (N10944, N10943, N10534, N3248, N5976);
nand NAND2 (N10945, N10944, N3536);
nand NAND3 (N10946, N10929, N7030, N10943);
and AND2 (N10947, N10940, N10326);
nor NOR3 (N10948, N10939, N7403, N10897);
xor XOR2 (N10949, N10941, N3817);
nor NOR2 (N10950, N10928, N2565);
buf BUF1 (N10951, N10927);
buf BUF1 (N10952, N10950);
and AND4 (N10953, N10946, N1916, N8249, N3095);
buf BUF1 (N10954, N10948);
buf BUF1 (N10955, N10937);
not NOT1 (N10956, N10951);
not NOT1 (N10957, N10947);
nor NOR4 (N10958, N10956, N10200, N8328, N4031);
not NOT1 (N10959, N10945);
and AND3 (N10960, N10942, N7294, N5726);
xor XOR2 (N10961, N10954, N1669);
buf BUF1 (N10962, N10961);
not NOT1 (N10963, N10959);
or OR4 (N10964, N10953, N8266, N2666, N6160);
and AND3 (N10965, N10960, N1851, N4422);
or OR2 (N10966, N10949, N2802);
nand NAND4 (N10967, N10957, N9630, N2832, N1893);
buf BUF1 (N10968, N10955);
or OR3 (N10969, N10967, N6711, N6194);
or OR4 (N10970, N10965, N5247, N10839, N3002);
xor XOR2 (N10971, N10970, N3189);
nand NAND2 (N10972, N10952, N7002);
xor XOR2 (N10973, N10972, N1019);
or OR3 (N10974, N10963, N9541, N1700);
and AND3 (N10975, N10958, N8350, N5817);
xor XOR2 (N10976, N10969, N9688);
buf BUF1 (N10977, N10976);
nor NOR4 (N10978, N10968, N9033, N8986, N5376);
or OR4 (N10979, N10962, N3194, N8327, N1167);
or OR3 (N10980, N10974, N655, N1356);
not NOT1 (N10981, N10977);
or OR2 (N10982, N10980, N7606);
nand NAND4 (N10983, N10938, N3234, N10632, N1959);
and AND4 (N10984, N10973, N1069, N8057, N1131);
xor XOR2 (N10985, N10981, N4570);
nand NAND3 (N10986, N10975, N10652, N5259);
nand NAND3 (N10987, N10966, N2624, N4413);
buf BUF1 (N10988, N10985);
nor NOR2 (N10989, N10987, N9211);
xor XOR2 (N10990, N10971, N5771);
nor NOR3 (N10991, N10990, N9199, N573);
not NOT1 (N10992, N10979);
nor NOR2 (N10993, N10984, N9286);
and AND4 (N10994, N10991, N8097, N251, N7853);
not NOT1 (N10995, N10994);
and AND3 (N10996, N10986, N5696, N6107);
nor NOR3 (N10997, N10988, N6467, N7576);
nand NAND4 (N10998, N10996, N4329, N1173, N5898);
or OR4 (N10999, N10978, N6017, N350, N1479);
xor XOR2 (N11000, N10992, N7091);
xor XOR2 (N11001, N10999, N767);
not NOT1 (N11002, N11001);
xor XOR2 (N11003, N10997, N6961);
buf BUF1 (N11004, N11003);
and AND2 (N11005, N10998, N2608);
and AND4 (N11006, N10964, N2506, N5468, N9454);
and AND4 (N11007, N10983, N7545, N10541, N7472);
not NOT1 (N11008, N10982);
nand NAND2 (N11009, N11006, N1755);
or OR4 (N11010, N11004, N3445, N9735, N7593);
buf BUF1 (N11011, N10993);
nor NOR3 (N11012, N11007, N10797, N1603);
nand NAND3 (N11013, N10995, N903, N7842);
buf BUF1 (N11014, N11005);
and AND3 (N11015, N11002, N8511, N2047);
and AND3 (N11016, N11011, N10706, N2633);
and AND2 (N11017, N11009, N6024);
buf BUF1 (N11018, N11017);
buf BUF1 (N11019, N11012);
not NOT1 (N11020, N11015);
xor XOR2 (N11021, N11013, N4497);
buf BUF1 (N11022, N11018);
xor XOR2 (N11023, N11008, N2192);
buf BUF1 (N11024, N11021);
or OR2 (N11025, N10989, N10810);
xor XOR2 (N11026, N11024, N4888);
not NOT1 (N11027, N11023);
nand NAND2 (N11028, N11019, N4258);
and AND3 (N11029, N11010, N1248, N7538);
not NOT1 (N11030, N11028);
nand NAND2 (N11031, N11014, N475);
buf BUF1 (N11032, N11000);
and AND2 (N11033, N11022, N6388);
nor NOR3 (N11034, N11030, N1433, N7581);
and AND4 (N11035, N11025, N5991, N9490, N3771);
xor XOR2 (N11036, N11016, N5073);
not NOT1 (N11037, N11029);
and AND3 (N11038, N11033, N8537, N3744);
nor NOR3 (N11039, N11020, N7040, N4504);
nand NAND3 (N11040, N11031, N6959, N3845);
and AND2 (N11041, N11026, N4200);
not NOT1 (N11042, N11027);
nor NOR3 (N11043, N11039, N1615, N8449);
nand NAND2 (N11044, N11040, N1941);
not NOT1 (N11045, N11036);
buf BUF1 (N11046, N11045);
nor NOR2 (N11047, N11038, N10843);
buf BUF1 (N11048, N11046);
nor NOR2 (N11049, N11041, N453);
or OR4 (N11050, N11047, N2392, N6147, N8436);
buf BUF1 (N11051, N11048);
nand NAND4 (N11052, N11051, N1821, N860, N1353);
or OR2 (N11053, N11034, N283);
or OR3 (N11054, N11053, N1657, N9295);
buf BUF1 (N11055, N11043);
xor XOR2 (N11056, N11042, N5404);
and AND4 (N11057, N11052, N10391, N6283, N3321);
nand NAND2 (N11058, N11049, N1182);
and AND3 (N11059, N11050, N7345, N10624);
and AND2 (N11060, N11054, N8223);
nor NOR4 (N11061, N11055, N8552, N8694, N497);
buf BUF1 (N11062, N11056);
and AND4 (N11063, N11032, N47, N2381, N2988);
nand NAND2 (N11064, N11044, N2835);
and AND3 (N11065, N11057, N103, N10612);
xor XOR2 (N11066, N11060, N3678);
buf BUF1 (N11067, N11063);
nand NAND2 (N11068, N11035, N9417);
xor XOR2 (N11069, N11064, N985);
not NOT1 (N11070, N11065);
xor XOR2 (N11071, N11067, N9448);
and AND2 (N11072, N11069, N4871);
and AND4 (N11073, N11058, N9668, N1928, N10753);
or OR4 (N11074, N11061, N2982, N3963, N1166);
nand NAND3 (N11075, N11073, N755, N4804);
and AND3 (N11076, N11071, N10659, N6787);
xor XOR2 (N11077, N11066, N3572);
buf BUF1 (N11078, N11075);
xor XOR2 (N11079, N11062, N970);
not NOT1 (N11080, N11070);
not NOT1 (N11081, N11078);
not NOT1 (N11082, N11081);
nand NAND4 (N11083, N11074, N9822, N5432, N7754);
buf BUF1 (N11084, N11077);
not NOT1 (N11085, N11076);
and AND4 (N11086, N11083, N8820, N3408, N1825);
not NOT1 (N11087, N11086);
nand NAND2 (N11088, N11059, N5865);
not NOT1 (N11089, N11084);
nor NOR4 (N11090, N11087, N6635, N9334, N1120);
nor NOR4 (N11091, N11072, N3519, N5203, N5712);
or OR3 (N11092, N11082, N1760, N5058);
xor XOR2 (N11093, N11091, N6209);
not NOT1 (N11094, N11080);
and AND2 (N11095, N11088, N217);
nor NOR2 (N11096, N11094, N7523);
nand NAND3 (N11097, N11093, N8768, N3343);
nand NAND4 (N11098, N11090, N7510, N3359, N4585);
nor NOR4 (N11099, N11098, N3469, N2445, N8811);
not NOT1 (N11100, N11089);
nor NOR3 (N11101, N11037, N9113, N8307);
or OR3 (N11102, N11095, N8013, N9410);
buf BUF1 (N11103, N11099);
buf BUF1 (N11104, N11079);
not NOT1 (N11105, N11096);
and AND3 (N11106, N11100, N2500, N4928);
or OR4 (N11107, N11105, N2912, N8275, N6243);
buf BUF1 (N11108, N11107);
and AND3 (N11109, N11104, N3509, N3226);
buf BUF1 (N11110, N11109);
xor XOR2 (N11111, N11085, N7591);
nor NOR2 (N11112, N11092, N2351);
buf BUF1 (N11113, N11097);
or OR2 (N11114, N11103, N6687);
nand NAND4 (N11115, N11102, N1949, N4190, N9767);
and AND3 (N11116, N11114, N908, N1393);
buf BUF1 (N11117, N11108);
buf BUF1 (N11118, N11068);
xor XOR2 (N11119, N11110, N10631);
buf BUF1 (N11120, N11119);
buf BUF1 (N11121, N11116);
not NOT1 (N11122, N11120);
or OR3 (N11123, N11111, N7341, N1186);
xor XOR2 (N11124, N11101, N1395);
not NOT1 (N11125, N11123);
and AND2 (N11126, N11118, N9973);
not NOT1 (N11127, N11113);
nor NOR4 (N11128, N11117, N4320, N8943, N9615);
and AND3 (N11129, N11128, N5331, N7396);
not NOT1 (N11130, N11115);
and AND3 (N11131, N11112, N10739, N417);
not NOT1 (N11132, N11131);
buf BUF1 (N11133, N11129);
not NOT1 (N11134, N11132);
nand NAND4 (N11135, N11125, N7294, N3629, N6902);
nand NAND3 (N11136, N11133, N3588, N8052);
or OR4 (N11137, N11124, N2233, N5186, N10346);
not NOT1 (N11138, N11136);
or OR2 (N11139, N11121, N8268);
nor NOR2 (N11140, N11126, N10871);
or OR4 (N11141, N11138, N452, N9421, N9094);
buf BUF1 (N11142, N11137);
or OR4 (N11143, N11122, N2607, N3043, N3673);
nor NOR3 (N11144, N11130, N8032, N3136);
buf BUF1 (N11145, N11143);
and AND3 (N11146, N11134, N938, N8637);
nor NOR4 (N11147, N11145, N9091, N2321, N1275);
not NOT1 (N11148, N11139);
buf BUF1 (N11149, N11147);
nand NAND2 (N11150, N11142, N10213);
nand NAND4 (N11151, N11146, N1953, N5461, N4418);
xor XOR2 (N11152, N11140, N4619);
and AND3 (N11153, N11148, N8732, N8065);
not NOT1 (N11154, N11151);
xor XOR2 (N11155, N11154, N5868);
and AND2 (N11156, N11144, N367);
or OR3 (N11157, N11135, N2407, N3435);
or OR4 (N11158, N11153, N6316, N8098, N4533);
buf BUF1 (N11159, N11155);
xor XOR2 (N11160, N11158, N3625);
and AND2 (N11161, N11157, N10539);
nor NOR4 (N11162, N11159, N6882, N5602, N2231);
nand NAND2 (N11163, N11160, N9467);
buf BUF1 (N11164, N11156);
buf BUF1 (N11165, N11162);
and AND4 (N11166, N11161, N373, N2202, N811);
buf BUF1 (N11167, N11164);
nand NAND3 (N11168, N11152, N617, N9479);
xor XOR2 (N11169, N11168, N9041);
buf BUF1 (N11170, N11169);
or OR2 (N11171, N11166, N3243);
nand NAND3 (N11172, N11171, N10224, N2390);
or OR4 (N11173, N11172, N10675, N5800, N992);
xor XOR2 (N11174, N11173, N9572);
nand NAND3 (N11175, N11127, N5088, N2055);
xor XOR2 (N11176, N11167, N4891);
not NOT1 (N11177, N11174);
and AND3 (N11178, N11149, N7479, N7551);
buf BUF1 (N11179, N11170);
buf BUF1 (N11180, N11141);
buf BUF1 (N11181, N11150);
not NOT1 (N11182, N11178);
xor XOR2 (N11183, N11175, N5601);
or OR2 (N11184, N11106, N4120);
not NOT1 (N11185, N11180);
nand NAND4 (N11186, N11181, N5985, N3876, N8504);
or OR2 (N11187, N11179, N10845);
and AND3 (N11188, N11163, N7770, N970);
not NOT1 (N11189, N11176);
xor XOR2 (N11190, N11186, N10727);
and AND2 (N11191, N11188, N4028);
and AND3 (N11192, N11183, N1847, N3822);
xor XOR2 (N11193, N11189, N9770);
not NOT1 (N11194, N11177);
xor XOR2 (N11195, N11165, N10438);
and AND3 (N11196, N11193, N5828, N5895);
buf BUF1 (N11197, N11185);
buf BUF1 (N11198, N11195);
or OR3 (N11199, N11191, N6717, N1565);
xor XOR2 (N11200, N11190, N5144);
buf BUF1 (N11201, N11197);
or OR3 (N11202, N11198, N4814, N1761);
not NOT1 (N11203, N11187);
and AND3 (N11204, N11184, N10311, N9758);
not NOT1 (N11205, N11194);
buf BUF1 (N11206, N11204);
and AND2 (N11207, N11182, N5610);
buf BUF1 (N11208, N11192);
nand NAND3 (N11209, N11201, N10412, N10967);
nor NOR3 (N11210, N11196, N8640, N9636);
nand NAND4 (N11211, N11206, N10025, N10687, N7135);
nand NAND2 (N11212, N11200, N4992);
nor NOR3 (N11213, N11209, N9024, N6384);
xor XOR2 (N11214, N11213, N6909);
buf BUF1 (N11215, N11203);
nor NOR3 (N11216, N11212, N7015, N9350);
not NOT1 (N11217, N11215);
nor NOR2 (N11218, N11199, N5605);
not NOT1 (N11219, N11217);
nand NAND3 (N11220, N11216, N9738, N10558);
xor XOR2 (N11221, N11214, N8183);
nand NAND3 (N11222, N11207, N10185, N292);
xor XOR2 (N11223, N11222, N5255);
buf BUF1 (N11224, N11211);
buf BUF1 (N11225, N11210);
xor XOR2 (N11226, N11220, N8682);
or OR4 (N11227, N11221, N1777, N2956, N7569);
xor XOR2 (N11228, N11224, N4895);
xor XOR2 (N11229, N11218, N3100);
nor NOR4 (N11230, N11228, N792, N6004, N5443);
nor NOR2 (N11231, N11227, N4454);
or OR2 (N11232, N11231, N4918);
and AND4 (N11233, N11223, N9948, N10761, N85);
nand NAND4 (N11234, N11219, N825, N2009, N5239);
nand NAND3 (N11235, N11232, N2595, N8880);
not NOT1 (N11236, N11205);
buf BUF1 (N11237, N11208);
nand NAND3 (N11238, N11237, N504, N9931);
buf BUF1 (N11239, N11233);
buf BUF1 (N11240, N11239);
nor NOR3 (N11241, N11202, N7315, N1547);
or OR3 (N11242, N11236, N5070, N905);
and AND4 (N11243, N11225, N8500, N10561, N4147);
not NOT1 (N11244, N11243);
or OR3 (N11245, N11242, N9216, N956);
nor NOR3 (N11246, N11241, N8278, N125);
buf BUF1 (N11247, N11240);
nor NOR4 (N11248, N11229, N5830, N10425, N3400);
nand NAND2 (N11249, N11238, N354);
xor XOR2 (N11250, N11245, N4177);
not NOT1 (N11251, N11247);
or OR4 (N11252, N11251, N8459, N2878, N9625);
nor NOR4 (N11253, N11226, N6334, N9497, N828);
not NOT1 (N11254, N11252);
nor NOR3 (N11255, N11249, N8227, N5573);
not NOT1 (N11256, N11244);
and AND3 (N11257, N11234, N2876, N8342);
or OR4 (N11258, N11235, N5542, N3559, N630);
or OR3 (N11259, N11254, N2679, N9108);
or OR4 (N11260, N11256, N8596, N6012, N1263);
buf BUF1 (N11261, N11255);
and AND2 (N11262, N11261, N6379);
and AND2 (N11263, N11250, N2003);
nor NOR2 (N11264, N11230, N5356);
nand NAND3 (N11265, N11258, N2420, N874);
not NOT1 (N11266, N11248);
and AND2 (N11267, N11257, N9955);
or OR2 (N11268, N11266, N2533);
xor XOR2 (N11269, N11264, N3438);
xor XOR2 (N11270, N11246, N11040);
nand NAND2 (N11271, N11270, N8539);
xor XOR2 (N11272, N11259, N2096);
nor NOR2 (N11273, N11253, N1937);
nor NOR2 (N11274, N11273, N5755);
or OR3 (N11275, N11269, N3140, N3350);
or OR3 (N11276, N11271, N3021, N1575);
nor NOR2 (N11277, N11260, N5543);
and AND3 (N11278, N11276, N6768, N10585);
nand NAND4 (N11279, N11262, N849, N7499, N4285);
xor XOR2 (N11280, N11263, N522);
or OR3 (N11281, N11278, N918, N1822);
nor NOR4 (N11282, N11272, N10576, N130, N4543);
and AND4 (N11283, N11279, N2523, N3670, N4409);
buf BUF1 (N11284, N11265);
or OR2 (N11285, N11282, N5096);
not NOT1 (N11286, N11280);
not NOT1 (N11287, N11267);
not NOT1 (N11288, N11281);
xor XOR2 (N11289, N11288, N8994);
nand NAND2 (N11290, N11277, N4330);
nand NAND2 (N11291, N11289, N11059);
nor NOR2 (N11292, N11283, N9143);
not NOT1 (N11293, N11275);
buf BUF1 (N11294, N11293);
not NOT1 (N11295, N11285);
nand NAND4 (N11296, N11284, N3813, N5665, N1937);
not NOT1 (N11297, N11291);
and AND2 (N11298, N11290, N7712);
nor NOR2 (N11299, N11268, N2134);
or OR4 (N11300, N11296, N8030, N10952, N8149);
not NOT1 (N11301, N11287);
and AND3 (N11302, N11294, N4837, N5093);
and AND2 (N11303, N11298, N6533);
buf BUF1 (N11304, N11297);
nor NOR3 (N11305, N11303, N10015, N8309);
not NOT1 (N11306, N11305);
xor XOR2 (N11307, N11274, N4353);
nand NAND4 (N11308, N11295, N4567, N8971, N7935);
nand NAND4 (N11309, N11306, N6039, N8846, N292);
nand NAND4 (N11310, N11292, N312, N4076, N2118);
not NOT1 (N11311, N11309);
buf BUF1 (N11312, N11301);
or OR2 (N11313, N11286, N6418);
xor XOR2 (N11314, N11304, N7868);
nor NOR3 (N11315, N11308, N4458, N8513);
buf BUF1 (N11316, N11307);
nand NAND3 (N11317, N11312, N843, N7799);
not NOT1 (N11318, N11311);
and AND2 (N11319, N11310, N9533);
nor NOR3 (N11320, N11314, N9388, N3552);
buf BUF1 (N11321, N11316);
or OR3 (N11322, N11315, N788, N5387);
not NOT1 (N11323, N11317);
nand NAND3 (N11324, N11320, N3631, N10862);
nand NAND4 (N11325, N11302, N7660, N11247, N392);
not NOT1 (N11326, N11322);
not NOT1 (N11327, N11326);
buf BUF1 (N11328, N11299);
buf BUF1 (N11329, N11327);
buf BUF1 (N11330, N11329);
nand NAND3 (N11331, N11321, N435, N10392);
or OR3 (N11332, N11319, N7677, N287);
not NOT1 (N11333, N11324);
and AND4 (N11334, N11332, N5186, N2841, N5453);
xor XOR2 (N11335, N11334, N11278);
and AND4 (N11336, N11313, N2197, N7457, N10881);
buf BUF1 (N11337, N11325);
buf BUF1 (N11338, N11328);
buf BUF1 (N11339, N11323);
not NOT1 (N11340, N11318);
buf BUF1 (N11341, N11337);
not NOT1 (N11342, N11333);
or OR3 (N11343, N11339, N4473, N2686);
buf BUF1 (N11344, N11343);
nor NOR3 (N11345, N11331, N8951, N7459);
xor XOR2 (N11346, N11344, N7103);
and AND4 (N11347, N11346, N6412, N4833, N4779);
and AND4 (N11348, N11341, N10103, N730, N8954);
or OR4 (N11349, N11338, N3720, N10862, N4864);
nor NOR4 (N11350, N11345, N9833, N11242, N2911);
xor XOR2 (N11351, N11336, N1269);
nor NOR4 (N11352, N11335, N9883, N2717, N857);
nand NAND3 (N11353, N11340, N5368, N10381);
buf BUF1 (N11354, N11350);
buf BUF1 (N11355, N11351);
nand NAND2 (N11356, N11352, N8492);
buf BUF1 (N11357, N11353);
buf BUF1 (N11358, N11330);
xor XOR2 (N11359, N11357, N10939);
or OR4 (N11360, N11300, N10055, N11324, N9422);
buf BUF1 (N11361, N11355);
xor XOR2 (N11362, N11348, N9369);
or OR2 (N11363, N11361, N6192);
buf BUF1 (N11364, N11358);
buf BUF1 (N11365, N11363);
buf BUF1 (N11366, N11347);
xor XOR2 (N11367, N11354, N4800);
nand NAND3 (N11368, N11356, N6011, N10253);
nand NAND3 (N11369, N11342, N2028, N11006);
or OR2 (N11370, N11364, N4065);
xor XOR2 (N11371, N11365, N1825);
and AND2 (N11372, N11362, N8507);
xor XOR2 (N11373, N11368, N3531);
or OR3 (N11374, N11349, N9990, N1282);
nor NOR3 (N11375, N11373, N5170, N3057);
and AND2 (N11376, N11369, N842);
and AND2 (N11377, N11360, N7706);
nand NAND4 (N11378, N11366, N6129, N5497, N3819);
and AND4 (N11379, N11377, N11358, N4029, N826);
xor XOR2 (N11380, N11367, N10897);
nor NOR3 (N11381, N11379, N8158, N95);
nand NAND2 (N11382, N11375, N1506);
nand NAND4 (N11383, N11370, N9979, N325, N494);
nand NAND3 (N11384, N11378, N10435, N10679);
buf BUF1 (N11385, N11381);
buf BUF1 (N11386, N11380);
nor NOR2 (N11387, N11384, N9100);
not NOT1 (N11388, N11374);
not NOT1 (N11389, N11376);
xor XOR2 (N11390, N11382, N1479);
buf BUF1 (N11391, N11385);
xor XOR2 (N11392, N11390, N1536);
nor NOR2 (N11393, N11371, N6487);
not NOT1 (N11394, N11388);
xor XOR2 (N11395, N11393, N7544);
not NOT1 (N11396, N11392);
nand NAND3 (N11397, N11396, N2100, N10733);
buf BUF1 (N11398, N11389);
not NOT1 (N11399, N11372);
or OR4 (N11400, N11383, N7647, N3958, N1943);
nor NOR4 (N11401, N11395, N848, N6915, N6425);
xor XOR2 (N11402, N11401, N2727);
xor XOR2 (N11403, N11397, N10290);
nor NOR4 (N11404, N11400, N5521, N4301, N9817);
xor XOR2 (N11405, N11386, N7371);
and AND3 (N11406, N11394, N4070, N6903);
and AND2 (N11407, N11359, N7674);
buf BUF1 (N11408, N11406);
and AND2 (N11409, N11407, N6062);
and AND2 (N11410, N11404, N4351);
nor NOR3 (N11411, N11399, N6431, N6794);
nand NAND4 (N11412, N11408, N11227, N9992, N4220);
xor XOR2 (N11413, N11391, N1596);
or OR4 (N11414, N11402, N1428, N8157, N3996);
and AND3 (N11415, N11411, N1475, N10281);
nand NAND4 (N11416, N11409, N903, N4346, N10871);
not NOT1 (N11417, N11387);
buf BUF1 (N11418, N11413);
not NOT1 (N11419, N11417);
xor XOR2 (N11420, N11414, N5648);
xor XOR2 (N11421, N11405, N6778);
xor XOR2 (N11422, N11398, N4101);
not NOT1 (N11423, N11421);
not NOT1 (N11424, N11418);
buf BUF1 (N11425, N11403);
nand NAND2 (N11426, N11423, N2071);
nor NOR4 (N11427, N11425, N7262, N10288, N680);
nand NAND4 (N11428, N11416, N2354, N6543, N3506);
not NOT1 (N11429, N11427);
not NOT1 (N11430, N11419);
xor XOR2 (N11431, N11429, N9286);
buf BUF1 (N11432, N11410);
nor NOR4 (N11433, N11431, N8508, N8925, N7535);
or OR3 (N11434, N11412, N3486, N6425);
or OR3 (N11435, N11424, N134, N7185);
not NOT1 (N11436, N11415);
nor NOR4 (N11437, N11428, N6108, N10905, N8249);
buf BUF1 (N11438, N11433);
buf BUF1 (N11439, N11426);
and AND4 (N11440, N11432, N1484, N683, N183);
not NOT1 (N11441, N11422);
nor NOR4 (N11442, N11420, N10804, N632, N4903);
and AND3 (N11443, N11438, N4184, N4957);
xor XOR2 (N11444, N11439, N2538);
buf BUF1 (N11445, N11434);
and AND2 (N11446, N11442, N3014);
nor NOR2 (N11447, N11445, N3705);
xor XOR2 (N11448, N11446, N10910);
not NOT1 (N11449, N11437);
or OR4 (N11450, N11440, N3160, N3046, N10320);
or OR2 (N11451, N11444, N329);
or OR4 (N11452, N11450, N4490, N10598, N8580);
nand NAND4 (N11453, N11449, N10527, N6561, N10837);
buf BUF1 (N11454, N11430);
nor NOR4 (N11455, N11447, N4281, N4071, N9825);
buf BUF1 (N11456, N11455);
or OR2 (N11457, N11435, N3762);
and AND4 (N11458, N11452, N11160, N8587, N303);
and AND3 (N11459, N11458, N2688, N2825);
nor NOR2 (N11460, N11456, N3529);
and AND3 (N11461, N11448, N11439, N6688);
xor XOR2 (N11462, N11451, N1606);
nand NAND4 (N11463, N11443, N2581, N8676, N1832);
nand NAND2 (N11464, N11453, N9072);
not NOT1 (N11465, N11436);
nor NOR4 (N11466, N11463, N4294, N7636, N11243);
and AND4 (N11467, N11464, N7280, N10113, N7328);
or OR3 (N11468, N11459, N6569, N4650);
not NOT1 (N11469, N11457);
nor NOR3 (N11470, N11467, N11074, N1149);
not NOT1 (N11471, N11470);
nand NAND4 (N11472, N11471, N3139, N8402, N9752);
not NOT1 (N11473, N11460);
xor XOR2 (N11474, N11466, N7438);
or OR2 (N11475, N11441, N2510);
and AND2 (N11476, N11468, N7293);
buf BUF1 (N11477, N11462);
buf BUF1 (N11478, N11474);
nor NOR4 (N11479, N11465, N3624, N4397, N9080);
or OR2 (N11480, N11469, N9586);
not NOT1 (N11481, N11478);
buf BUF1 (N11482, N11472);
xor XOR2 (N11483, N11481, N4273);
xor XOR2 (N11484, N11461, N1765);
and AND4 (N11485, N11475, N1678, N2132, N8663);
and AND4 (N11486, N11484, N1554, N7416, N4595);
xor XOR2 (N11487, N11476, N8283);
xor XOR2 (N11488, N11486, N2326);
nand NAND2 (N11489, N11473, N5462);
nand NAND2 (N11490, N11488, N9942);
or OR3 (N11491, N11477, N1521, N3887);
nor NOR2 (N11492, N11487, N5686);
not NOT1 (N11493, N11454);
buf BUF1 (N11494, N11493);
or OR2 (N11495, N11491, N9664);
or OR2 (N11496, N11495, N7015);
nand NAND4 (N11497, N11479, N946, N4108, N4180);
and AND4 (N11498, N11492, N3692, N9962, N2768);
nor NOR3 (N11499, N11490, N242, N10065);
nand NAND4 (N11500, N11499, N1737, N9704, N7075);
and AND3 (N11501, N11480, N2242, N5195);
nand NAND4 (N11502, N11483, N4440, N7090, N10747);
not NOT1 (N11503, N11489);
nor NOR3 (N11504, N11494, N1409, N735);
xor XOR2 (N11505, N11485, N573);
nand NAND2 (N11506, N11482, N595);
not NOT1 (N11507, N11498);
or OR2 (N11508, N11502, N9100);
not NOT1 (N11509, N11503);
nor NOR2 (N11510, N11496, N1488);
buf BUF1 (N11511, N11501);
nand NAND3 (N11512, N11508, N10651, N11209);
not NOT1 (N11513, N11511);
and AND3 (N11514, N11509, N8539, N8705);
nand NAND3 (N11515, N11497, N315, N3719);
xor XOR2 (N11516, N11510, N4602);
xor XOR2 (N11517, N11516, N10934);
nor NOR4 (N11518, N11512, N9123, N5834, N10920);
nand NAND3 (N11519, N11507, N7124, N4927);
nor NOR3 (N11520, N11515, N9962, N2065);
nor NOR4 (N11521, N11513, N2117, N1882, N2307);
buf BUF1 (N11522, N11519);
buf BUF1 (N11523, N11518);
and AND3 (N11524, N11517, N1851, N9750);
nor NOR3 (N11525, N11504, N4499, N5958);
xor XOR2 (N11526, N11500, N5927);
or OR4 (N11527, N11525, N8236, N1663, N11087);
nor NOR2 (N11528, N11524, N5470);
or OR3 (N11529, N11523, N10501, N4883);
buf BUF1 (N11530, N11522);
not NOT1 (N11531, N11527);
buf BUF1 (N11532, N11528);
nor NOR2 (N11533, N11529, N8814);
or OR4 (N11534, N11520, N971, N2430, N1932);
and AND2 (N11535, N11514, N9705);
buf BUF1 (N11536, N11535);
buf BUF1 (N11537, N11521);
not NOT1 (N11538, N11530);
and AND2 (N11539, N11538, N5900);
nand NAND2 (N11540, N11506, N10399);
not NOT1 (N11541, N11540);
buf BUF1 (N11542, N11536);
nand NAND3 (N11543, N11531, N413, N5213);
or OR2 (N11544, N11542, N11108);
buf BUF1 (N11545, N11543);
or OR3 (N11546, N11532, N3629, N6163);
not NOT1 (N11547, N11546);
nor NOR3 (N11548, N11539, N9837, N8896);
and AND2 (N11549, N11548, N9940);
nor NOR3 (N11550, N11544, N1344, N4133);
buf BUF1 (N11551, N11550);
xor XOR2 (N11552, N11549, N5704);
nor NOR3 (N11553, N11545, N5024, N5927);
nor NOR4 (N11554, N11547, N3740, N3130, N7117);
nand NAND2 (N11555, N11533, N5488);
buf BUF1 (N11556, N11551);
xor XOR2 (N11557, N11526, N3051);
buf BUF1 (N11558, N11534);
nand NAND3 (N11559, N11505, N7200, N970);
nand NAND4 (N11560, N11557, N9276, N9473, N4235);
buf BUF1 (N11561, N11555);
nand NAND4 (N11562, N11554, N2776, N9977, N4945);
or OR2 (N11563, N11560, N5940);
nor NOR3 (N11564, N11541, N2794, N10120);
not NOT1 (N11565, N11553);
or OR2 (N11566, N11561, N3102);
not NOT1 (N11567, N11558);
or OR3 (N11568, N11563, N4761, N855);
not NOT1 (N11569, N11556);
nand NAND2 (N11570, N11568, N7255);
not NOT1 (N11571, N11564);
buf BUF1 (N11572, N11537);
xor XOR2 (N11573, N11552, N10022);
not NOT1 (N11574, N11572);
nand NAND3 (N11575, N11565, N9282, N8761);
not NOT1 (N11576, N11567);
nor NOR3 (N11577, N11569, N1254, N2651);
and AND4 (N11578, N11573, N8341, N7042, N11351);
nand NAND3 (N11579, N11570, N2833, N10632);
not NOT1 (N11580, N11571);
and AND3 (N11581, N11579, N8047, N4175);
nand NAND3 (N11582, N11578, N3960, N2891);
not NOT1 (N11583, N11580);
nor NOR3 (N11584, N11566, N10416, N5581);
nor NOR2 (N11585, N11559, N8735);
nand NAND2 (N11586, N11585, N1776);
buf BUF1 (N11587, N11582);
nor NOR2 (N11588, N11577, N2473);
nor NOR3 (N11589, N11586, N6933, N1572);
or OR2 (N11590, N11562, N10245);
nor NOR2 (N11591, N11581, N26);
buf BUF1 (N11592, N11574);
not NOT1 (N11593, N11591);
not NOT1 (N11594, N11575);
xor XOR2 (N11595, N11576, N1545);
xor XOR2 (N11596, N11587, N6017);
nor NOR3 (N11597, N11596, N1477, N8479);
not NOT1 (N11598, N11595);
nand NAND2 (N11599, N11594, N6348);
buf BUF1 (N11600, N11589);
and AND3 (N11601, N11593, N6418, N11304);
or OR2 (N11602, N11600, N6569);
and AND2 (N11603, N11602, N6076);
and AND2 (N11604, N11597, N5953);
or OR4 (N11605, N11584, N8654, N9269, N6327);
and AND3 (N11606, N11599, N2145, N2525);
xor XOR2 (N11607, N11605, N1347);
buf BUF1 (N11608, N11590);
nand NAND3 (N11609, N11606, N5593, N10071);
or OR3 (N11610, N11592, N7209, N6252);
nor NOR2 (N11611, N11609, N10735);
or OR2 (N11612, N11603, N10726);
xor XOR2 (N11613, N11607, N8777);
or OR2 (N11614, N11613, N2437);
nor NOR4 (N11615, N11588, N3158, N9713, N11405);
nor NOR3 (N11616, N11601, N9073, N7622);
xor XOR2 (N11617, N11598, N4692);
and AND4 (N11618, N11583, N10385, N1095, N1329);
and AND3 (N11619, N11612, N5026, N11433);
not NOT1 (N11620, N11616);
xor XOR2 (N11621, N11610, N11488);
nand NAND2 (N11622, N11618, N89);
and AND4 (N11623, N11622, N537, N6365, N7997);
nand NAND4 (N11624, N11620, N9367, N6412, N3195);
buf BUF1 (N11625, N11621);
nor NOR2 (N11626, N11623, N5661);
not NOT1 (N11627, N11611);
nor NOR2 (N11628, N11624, N1421);
nand NAND3 (N11629, N11628, N5786, N534);
not NOT1 (N11630, N11619);
nand NAND2 (N11631, N11625, N7878);
nor NOR4 (N11632, N11630, N3759, N3102, N4125);
xor XOR2 (N11633, N11627, N4332);
nand NAND2 (N11634, N11614, N7604);
nor NOR3 (N11635, N11632, N7929, N4779);
nor NOR4 (N11636, N11626, N5370, N8065, N8058);
buf BUF1 (N11637, N11635);
xor XOR2 (N11638, N11631, N5458);
or OR2 (N11639, N11638, N7138);
nor NOR4 (N11640, N11617, N10196, N8131, N10799);
and AND2 (N11641, N11640, N421);
buf BUF1 (N11642, N11629);
nand NAND2 (N11643, N11641, N7433);
xor XOR2 (N11644, N11634, N10442);
nand NAND2 (N11645, N11637, N582);
nand NAND2 (N11646, N11639, N11391);
and AND2 (N11647, N11642, N652);
and AND4 (N11648, N11615, N1500, N4297, N10816);
nand NAND3 (N11649, N11636, N3873, N4479);
buf BUF1 (N11650, N11647);
nor NOR3 (N11651, N11646, N3282, N5509);
nor NOR2 (N11652, N11649, N9323);
xor XOR2 (N11653, N11651, N8251);
nor NOR3 (N11654, N11648, N2985, N2720);
not NOT1 (N11655, N11652);
xor XOR2 (N11656, N11654, N658);
xor XOR2 (N11657, N11633, N9345);
or OR3 (N11658, N11645, N3203, N10390);
nor NOR2 (N11659, N11650, N1111);
xor XOR2 (N11660, N11643, N5425);
and AND4 (N11661, N11658, N266, N11505, N1785);
buf BUF1 (N11662, N11644);
buf BUF1 (N11663, N11661);
buf BUF1 (N11664, N11604);
or OR3 (N11665, N11659, N11067, N4635);
nand NAND2 (N11666, N11665, N5982);
not NOT1 (N11667, N11608);
and AND2 (N11668, N11664, N10296);
xor XOR2 (N11669, N11662, N8354);
nor NOR2 (N11670, N11667, N10310);
xor XOR2 (N11671, N11660, N4056);
nand NAND2 (N11672, N11670, N6557);
buf BUF1 (N11673, N11668);
or OR4 (N11674, N11663, N8152, N1756, N9322);
nor NOR3 (N11675, N11673, N1291, N4058);
or OR3 (N11676, N11671, N7175, N6714);
and AND2 (N11677, N11657, N10934);
nand NAND2 (N11678, N11672, N11145);
not NOT1 (N11679, N11653);
buf BUF1 (N11680, N11674);
nand NAND3 (N11681, N11676, N7608, N7038);
nand NAND4 (N11682, N11680, N8145, N8794, N6295);
xor XOR2 (N11683, N11675, N601);
nand NAND3 (N11684, N11683, N9913, N1300);
xor XOR2 (N11685, N11677, N1330);
nand NAND4 (N11686, N11678, N10840, N893, N1575);
nor NOR2 (N11687, N11669, N8364);
buf BUF1 (N11688, N11656);
nor NOR4 (N11689, N11679, N10604, N11343, N9925);
or OR3 (N11690, N11689, N9588, N2165);
buf BUF1 (N11691, N11690);
not NOT1 (N11692, N11688);
and AND2 (N11693, N11691, N9257);
nor NOR4 (N11694, N11687, N1266, N7253, N8288);
not NOT1 (N11695, N11692);
nand NAND2 (N11696, N11655, N352);
buf BUF1 (N11697, N11685);
nand NAND4 (N11698, N11696, N2124, N9396, N9967);
and AND4 (N11699, N11693, N9438, N8933, N7499);
and AND4 (N11700, N11699, N4176, N2179, N1320);
nand NAND2 (N11701, N11700, N11640);
nand NAND4 (N11702, N11666, N10322, N3603, N4686);
and AND2 (N11703, N11698, N5206);
or OR4 (N11704, N11681, N4076, N11606, N244);
nor NOR2 (N11705, N11695, N7906);
not NOT1 (N11706, N11697);
xor XOR2 (N11707, N11706, N8845);
nand NAND4 (N11708, N11705, N9364, N2316, N11288);
nand NAND3 (N11709, N11682, N8606, N7036);
xor XOR2 (N11710, N11704, N2382);
not NOT1 (N11711, N11707);
nor NOR4 (N11712, N11684, N6195, N10580, N3400);
nor NOR3 (N11713, N11708, N5082, N5318);
not NOT1 (N11714, N11711);
nor NOR3 (N11715, N11713, N6023, N10288);
or OR2 (N11716, N11709, N237);
and AND4 (N11717, N11703, N3411, N9014, N7350);
nor NOR2 (N11718, N11702, N8082);
xor XOR2 (N11719, N11717, N7922);
nor NOR3 (N11720, N11716, N11222, N7208);
and AND2 (N11721, N11720, N4146);
buf BUF1 (N11722, N11694);
not NOT1 (N11723, N11718);
and AND2 (N11724, N11715, N3342);
xor XOR2 (N11725, N11686, N5886);
nand NAND4 (N11726, N11714, N7293, N2312, N4057);
or OR4 (N11727, N11712, N3834, N5886, N11190);
xor XOR2 (N11728, N11710, N239);
nand NAND2 (N11729, N11726, N2919);
buf BUF1 (N11730, N11721);
xor XOR2 (N11731, N11730, N2749);
and AND4 (N11732, N11701, N4606, N5482, N4532);
not NOT1 (N11733, N11731);
not NOT1 (N11734, N11719);
nand NAND2 (N11735, N11724, N4439);
nor NOR2 (N11736, N11727, N237);
not NOT1 (N11737, N11732);
xor XOR2 (N11738, N11728, N96);
or OR2 (N11739, N11722, N3922);
nor NOR2 (N11740, N11739, N401);
not NOT1 (N11741, N11723);
xor XOR2 (N11742, N11741, N11453);
or OR2 (N11743, N11725, N7229);
xor XOR2 (N11744, N11734, N2014);
and AND3 (N11745, N11742, N3204, N5339);
buf BUF1 (N11746, N11733);
xor XOR2 (N11747, N11737, N7924);
or OR2 (N11748, N11735, N5106);
or OR4 (N11749, N11748, N10113, N2192, N5381);
buf BUF1 (N11750, N11744);
nand NAND2 (N11751, N11743, N5132);
xor XOR2 (N11752, N11738, N2725);
or OR4 (N11753, N11729, N9121, N4077, N11284);
nor NOR2 (N11754, N11746, N3101);
buf BUF1 (N11755, N11749);
nor NOR2 (N11756, N11755, N5379);
not NOT1 (N11757, N11752);
nand NAND4 (N11758, N11745, N9952, N723, N8237);
nor NOR3 (N11759, N11757, N6271, N6871);
nor NOR4 (N11760, N11753, N2073, N5995, N5152);
not NOT1 (N11761, N11750);
or OR2 (N11762, N11761, N2906);
nor NOR3 (N11763, N11736, N195, N899);
buf BUF1 (N11764, N11756);
not NOT1 (N11765, N11740);
or OR4 (N11766, N11751, N11698, N11186, N6077);
xor XOR2 (N11767, N11754, N3811);
buf BUF1 (N11768, N11759);
not NOT1 (N11769, N11767);
nand NAND2 (N11770, N11762, N11123);
nand NAND4 (N11771, N11769, N10065, N3397, N9812);
nand NAND4 (N11772, N11760, N9606, N3032, N667);
nor NOR3 (N11773, N11758, N10491, N2025);
nor NOR4 (N11774, N11766, N5166, N5779, N6887);
or OR3 (N11775, N11774, N4158, N7078);
xor XOR2 (N11776, N11747, N8252);
not NOT1 (N11777, N11764);
nor NOR2 (N11778, N11775, N4);
xor XOR2 (N11779, N11763, N6917);
nand NAND2 (N11780, N11770, N9356);
or OR3 (N11781, N11776, N5485, N1828);
buf BUF1 (N11782, N11765);
xor XOR2 (N11783, N11777, N6040);
not NOT1 (N11784, N11773);
not NOT1 (N11785, N11783);
not NOT1 (N11786, N11772);
xor XOR2 (N11787, N11785, N2711);
nand NAND4 (N11788, N11784, N8583, N4995, N8699);
not NOT1 (N11789, N11778);
buf BUF1 (N11790, N11768);
buf BUF1 (N11791, N11780);
buf BUF1 (N11792, N11781);
xor XOR2 (N11793, N11771, N10776);
or OR4 (N11794, N11791, N5037, N9886, N7230);
nor NOR4 (N11795, N11788, N9546, N9723, N7864);
xor XOR2 (N11796, N11793, N378);
and AND3 (N11797, N11792, N6465, N10432);
nand NAND3 (N11798, N11790, N330, N6805);
nor NOR2 (N11799, N11782, N8956);
or OR3 (N11800, N11794, N11706, N4877);
nor NOR3 (N11801, N11795, N6269, N11326);
nand NAND3 (N11802, N11779, N10924, N1132);
nand NAND3 (N11803, N11799, N6141, N10818);
nor NOR3 (N11804, N11800, N2550, N665);
buf BUF1 (N11805, N11786);
xor XOR2 (N11806, N11797, N797);
nor NOR3 (N11807, N11787, N3841, N15);
or OR4 (N11808, N11806, N8056, N5739, N7795);
or OR4 (N11809, N11804, N8366, N10496, N2852);
or OR3 (N11810, N11801, N5920, N10503);
and AND2 (N11811, N11807, N5779);
xor XOR2 (N11812, N11809, N181);
not NOT1 (N11813, N11789);
or OR4 (N11814, N11796, N11561, N10492, N5393);
nand NAND4 (N11815, N11803, N6867, N7984, N8431);
nand NAND2 (N11816, N11808, N1106);
nand NAND3 (N11817, N11802, N7515, N4885);
and AND3 (N11818, N11811, N8937, N5861);
not NOT1 (N11819, N11815);
buf BUF1 (N11820, N11816);
or OR4 (N11821, N11818, N4494, N2029, N3037);
or OR3 (N11822, N11819, N1480, N6732);
buf BUF1 (N11823, N11822);
not NOT1 (N11824, N11813);
nand NAND4 (N11825, N11812, N4870, N7122, N6025);
nand NAND2 (N11826, N11825, N11678);
nor NOR2 (N11827, N11814, N890);
buf BUF1 (N11828, N11820);
not NOT1 (N11829, N11827);
nand NAND3 (N11830, N11829, N110, N445);
nor NOR3 (N11831, N11828, N5078, N126);
not NOT1 (N11832, N11805);
or OR4 (N11833, N11830, N760, N1633, N6627);
nor NOR4 (N11834, N11823, N3218, N3271, N1083);
or OR4 (N11835, N11831, N4603, N11016, N3366);
nor NOR3 (N11836, N11798, N2391, N10091);
and AND2 (N11837, N11824, N9642);
buf BUF1 (N11838, N11821);
nand NAND4 (N11839, N11837, N69, N488, N8190);
nand NAND3 (N11840, N11836, N7597, N8051);
and AND3 (N11841, N11833, N3711, N7411);
or OR4 (N11842, N11834, N37, N4847, N779);
nor NOR2 (N11843, N11842, N6689);
buf BUF1 (N11844, N11843);
and AND3 (N11845, N11841, N3763, N2848);
not NOT1 (N11846, N11835);
and AND3 (N11847, N11817, N2600, N5391);
nor NOR3 (N11848, N11838, N371, N8583);
xor XOR2 (N11849, N11832, N10969);
and AND4 (N11850, N11826, N4520, N1917, N6176);
and AND2 (N11851, N11850, N1483);
buf BUF1 (N11852, N11847);
or OR3 (N11853, N11852, N1904, N2996);
and AND4 (N11854, N11844, N8981, N9977, N1003);
nand NAND2 (N11855, N11840, N2569);
nor NOR2 (N11856, N11839, N2670);
nor NOR4 (N11857, N11849, N11252, N6610, N5241);
buf BUF1 (N11858, N11854);
and AND2 (N11859, N11851, N4554);
or OR2 (N11860, N11859, N9171);
not NOT1 (N11861, N11857);
and AND4 (N11862, N11858, N9388, N10063, N10061);
nand NAND2 (N11863, N11846, N2717);
xor XOR2 (N11864, N11855, N4021);
xor XOR2 (N11865, N11864, N5501);
or OR4 (N11866, N11861, N9360, N4103, N6321);
and AND3 (N11867, N11865, N2325, N7788);
xor XOR2 (N11868, N11853, N7443);
or OR3 (N11869, N11845, N2639, N8383);
nor NOR3 (N11870, N11866, N3236, N3710);
nor NOR2 (N11871, N11867, N7201);
buf BUF1 (N11872, N11868);
and AND4 (N11873, N11848, N5666, N10456, N6688);
or OR2 (N11874, N11869, N11701);
nand NAND3 (N11875, N11870, N11495, N6693);
nor NOR2 (N11876, N11874, N8684);
or OR4 (N11877, N11862, N3576, N6603, N8365);
not NOT1 (N11878, N11860);
xor XOR2 (N11879, N11875, N4456);
xor XOR2 (N11880, N11863, N5906);
and AND2 (N11881, N11879, N6177);
nand NAND3 (N11882, N11880, N9018, N2667);
buf BUF1 (N11883, N11882);
or OR4 (N11884, N11810, N11496, N7792, N2513);
nor NOR3 (N11885, N11881, N9112, N1541);
not NOT1 (N11886, N11877);
nand NAND2 (N11887, N11878, N5622);
nor NOR4 (N11888, N11883, N10031, N9406, N9151);
xor XOR2 (N11889, N11885, N2411);
nand NAND2 (N11890, N11872, N11044);
or OR3 (N11891, N11888, N10342, N2097);
xor XOR2 (N11892, N11890, N2903);
not NOT1 (N11893, N11891);
nor NOR3 (N11894, N11893, N559, N11182);
nand NAND4 (N11895, N11856, N11537, N2392, N4118);
not NOT1 (N11896, N11892);
and AND3 (N11897, N11884, N4119, N10279);
xor XOR2 (N11898, N11895, N5521);
or OR3 (N11899, N11894, N10543, N4528);
buf BUF1 (N11900, N11873);
xor XOR2 (N11901, N11889, N9786);
buf BUF1 (N11902, N11901);
or OR2 (N11903, N11900, N10893);
or OR3 (N11904, N11899, N5306, N9305);
buf BUF1 (N11905, N11898);
and AND4 (N11906, N11903, N8907, N9663, N9247);
or OR3 (N11907, N11871, N6232, N3826);
nor NOR3 (N11908, N11902, N1105, N831);
nand NAND3 (N11909, N11907, N10846, N5431);
not NOT1 (N11910, N11905);
xor XOR2 (N11911, N11904, N10816);
not NOT1 (N11912, N11887);
xor XOR2 (N11913, N11911, N5612);
not NOT1 (N11914, N11896);
buf BUF1 (N11915, N11906);
nand NAND3 (N11916, N11915, N10823, N9422);
or OR3 (N11917, N11912, N10654, N11158);
and AND3 (N11918, N11909, N6721, N9253);
nand NAND2 (N11919, N11876, N9867);
nand NAND4 (N11920, N11886, N10536, N8783, N6395);
xor XOR2 (N11921, N11920, N35);
xor XOR2 (N11922, N11921, N469);
not NOT1 (N11923, N11922);
and AND4 (N11924, N11923, N10876, N8639, N10021);
not NOT1 (N11925, N11914);
nor NOR3 (N11926, N11908, N7548, N3065);
nor NOR2 (N11927, N11916, N8479);
nand NAND2 (N11928, N11913, N1234);
and AND4 (N11929, N11917, N9449, N9028, N3627);
nor NOR3 (N11930, N11897, N9508, N8641);
nor NOR4 (N11931, N11927, N4642, N9511, N6793);
not NOT1 (N11932, N11918);
not NOT1 (N11933, N11924);
xor XOR2 (N11934, N11930, N9096);
nor NOR2 (N11935, N11932, N10058);
xor XOR2 (N11936, N11934, N2885);
buf BUF1 (N11937, N11919);
nand NAND4 (N11938, N11929, N1149, N11817, N5129);
nor NOR2 (N11939, N11935, N890);
and AND2 (N11940, N11936, N4233);
buf BUF1 (N11941, N11938);
and AND4 (N11942, N11925, N4130, N3933, N3455);
nor NOR3 (N11943, N11928, N1862, N2352);
or OR2 (N11944, N11940, N2118);
xor XOR2 (N11945, N11910, N2223);
nand NAND2 (N11946, N11937, N10878);
and AND3 (N11947, N11944, N1000, N10396);
and AND4 (N11948, N11926, N5301, N1418, N10702);
or OR2 (N11949, N11946, N5482);
nand NAND3 (N11950, N11933, N8021, N819);
or OR4 (N11951, N11941, N9183, N9392, N1609);
or OR2 (N11952, N11931, N1434);
nor NOR2 (N11953, N11948, N3708);
not NOT1 (N11954, N11953);
and AND2 (N11955, N11954, N11531);
and AND2 (N11956, N11950, N7506);
buf BUF1 (N11957, N11951);
not NOT1 (N11958, N11942);
xor XOR2 (N11959, N11956, N10959);
buf BUF1 (N11960, N11939);
or OR2 (N11961, N11943, N8777);
buf BUF1 (N11962, N11949);
not NOT1 (N11963, N11962);
and AND4 (N11964, N11945, N91, N9690, N5291);
and AND3 (N11965, N11952, N9881, N5284);
nor NOR2 (N11966, N11957, N2431);
not NOT1 (N11967, N11964);
not NOT1 (N11968, N11961);
nand NAND3 (N11969, N11960, N8856, N7087);
not NOT1 (N11970, N11966);
not NOT1 (N11971, N11967);
or OR2 (N11972, N11947, N3497);
xor XOR2 (N11973, N11958, N9960);
buf BUF1 (N11974, N11959);
and AND4 (N11975, N11965, N10976, N5194, N11340);
buf BUF1 (N11976, N11968);
nor NOR2 (N11977, N11963, N10496);
and AND4 (N11978, N11975, N4330, N11169, N11465);
xor XOR2 (N11979, N11969, N3948);
buf BUF1 (N11980, N11979);
not NOT1 (N11981, N11976);
buf BUF1 (N11982, N11974);
buf BUF1 (N11983, N11972);
nor NOR3 (N11984, N11971, N1674, N5963);
or OR4 (N11985, N11978, N8235, N2353, N9028);
nand NAND4 (N11986, N11955, N10404, N9584, N8417);
xor XOR2 (N11987, N11986, N4244);
xor XOR2 (N11988, N11984, N7746);
buf BUF1 (N11989, N11985);
buf BUF1 (N11990, N11987);
xor XOR2 (N11991, N11981, N3729);
or OR2 (N11992, N11970, N7512);
and AND3 (N11993, N11990, N11032, N11239);
xor XOR2 (N11994, N11973, N7007);
and AND3 (N11995, N11994, N8836, N4304);
nand NAND4 (N11996, N11983, N3540, N11466, N10779);
buf BUF1 (N11997, N11982);
nor NOR3 (N11998, N11997, N7494, N961);
and AND3 (N11999, N11989, N2313, N1364);
or OR3 (N12000, N11988, N6626, N10086);
nand NAND3 (N12001, N11991, N4124, N6484);
nand NAND2 (N12002, N11977, N7590);
not NOT1 (N12003, N11995);
nand NAND2 (N12004, N11980, N5773);
not NOT1 (N12005, N12004);
not NOT1 (N12006, N11993);
and AND3 (N12007, N12002, N4451, N1394);
xor XOR2 (N12008, N12000, N9819);
not NOT1 (N12009, N12005);
buf BUF1 (N12010, N12008);
or OR2 (N12011, N11998, N3160);
and AND2 (N12012, N12007, N6175);
nand NAND2 (N12013, N12009, N6749);
and AND2 (N12014, N11999, N6932);
buf BUF1 (N12015, N12003);
not NOT1 (N12016, N12015);
buf BUF1 (N12017, N11992);
nor NOR2 (N12018, N12006, N7745);
and AND3 (N12019, N12001, N2838, N1665);
or OR2 (N12020, N12019, N2348);
xor XOR2 (N12021, N12020, N8554);
nand NAND2 (N12022, N12013, N708);
and AND3 (N12023, N12016, N11370, N4067);
and AND4 (N12024, N12017, N8346, N7973, N665);
nor NOR4 (N12025, N12024, N8126, N4085, N9342);
xor XOR2 (N12026, N12012, N5069);
nand NAND3 (N12027, N12026, N8434, N7618);
not NOT1 (N12028, N12010);
buf BUF1 (N12029, N12011);
or OR2 (N12030, N12014, N8484);
xor XOR2 (N12031, N12027, N579);
buf BUF1 (N12032, N12030);
not NOT1 (N12033, N12021);
buf BUF1 (N12034, N12025);
nand NAND3 (N12035, N12018, N1207, N4257);
or OR2 (N12036, N12029, N3062);
or OR3 (N12037, N12032, N869, N7060);
not NOT1 (N12038, N11996);
not NOT1 (N12039, N12023);
nor NOR2 (N12040, N12031, N10760);
nor NOR2 (N12041, N12033, N2374);
xor XOR2 (N12042, N12028, N390);
nand NAND4 (N12043, N12040, N2940, N4919, N6321);
and AND4 (N12044, N12042, N11403, N210, N6888);
not NOT1 (N12045, N12044);
nor NOR2 (N12046, N12034, N9829);
nand NAND4 (N12047, N12022, N10378, N5765, N7276);
nor NOR2 (N12048, N12046, N1329);
and AND2 (N12049, N12043, N9657);
nand NAND2 (N12050, N12047, N10178);
xor XOR2 (N12051, N12048, N10194);
nand NAND4 (N12052, N12035, N11125, N5995, N10666);
or OR2 (N12053, N12045, N11811);
xor XOR2 (N12054, N12037, N9677);
nor NOR2 (N12055, N12054, N9244);
nand NAND3 (N12056, N12051, N4663, N4587);
xor XOR2 (N12057, N12041, N10121);
or OR3 (N12058, N12057, N6333, N7536);
buf BUF1 (N12059, N12050);
not NOT1 (N12060, N12055);
nor NOR2 (N12061, N12036, N957);
nor NOR2 (N12062, N12053, N11338);
nor NOR4 (N12063, N12052, N7548, N2966, N9738);
nand NAND3 (N12064, N12056, N6149, N2842);
nor NOR3 (N12065, N12049, N7879, N2175);
and AND2 (N12066, N12063, N3395);
nand NAND3 (N12067, N12066, N3931, N2980);
xor XOR2 (N12068, N12065, N3041);
or OR4 (N12069, N12067, N5920, N2622, N2528);
nand NAND3 (N12070, N12062, N5678, N72);
nand NAND4 (N12071, N12038, N5702, N3854, N7407);
or OR2 (N12072, N12068, N11462);
nand NAND4 (N12073, N12070, N10392, N682, N7535);
and AND4 (N12074, N12060, N2153, N10250, N3502);
buf BUF1 (N12075, N12069);
buf BUF1 (N12076, N12071);
nand NAND4 (N12077, N12059, N3953, N8082, N11149);
xor XOR2 (N12078, N12058, N2297);
nand NAND3 (N12079, N12061, N3188, N4029);
nor NOR4 (N12080, N12064, N444, N4271, N4885);
or OR4 (N12081, N12075, N8770, N10919, N10240);
and AND3 (N12082, N12072, N2603, N300);
xor XOR2 (N12083, N12082, N6387);
nor NOR3 (N12084, N12077, N6771, N3475);
not NOT1 (N12085, N12084);
or OR4 (N12086, N12078, N9535, N9103, N4274);
and AND2 (N12087, N12073, N1600);
xor XOR2 (N12088, N12086, N6147);
nor NOR3 (N12089, N12081, N2891, N2705);
or OR3 (N12090, N12079, N6867, N7796);
nand NAND4 (N12091, N12039, N3137, N7730, N9017);
or OR4 (N12092, N12074, N6812, N11745, N4791);
and AND2 (N12093, N12091, N5336);
buf BUF1 (N12094, N12076);
nand NAND2 (N12095, N12080, N8525);
and AND4 (N12096, N12085, N2096, N783, N1614);
buf BUF1 (N12097, N12095);
xor XOR2 (N12098, N12087, N8746);
xor XOR2 (N12099, N12092, N11253);
nand NAND4 (N12100, N12099, N11292, N3334, N99);
or OR3 (N12101, N12097, N10493, N3999);
and AND4 (N12102, N12090, N2318, N12062, N1050);
nand NAND3 (N12103, N12094, N4868, N8562);
not NOT1 (N12104, N12083);
xor XOR2 (N12105, N12103, N10278);
buf BUF1 (N12106, N12089);
nor NOR2 (N12107, N12093, N10750);
xor XOR2 (N12108, N12096, N11903);
not NOT1 (N12109, N12102);
nand NAND2 (N12110, N12108, N10956);
and AND3 (N12111, N12101, N4467, N2772);
and AND4 (N12112, N12106, N7385, N5642, N847);
xor XOR2 (N12113, N12100, N1580);
or OR3 (N12114, N12112, N2982, N8185);
not NOT1 (N12115, N12088);
buf BUF1 (N12116, N12110);
and AND4 (N12117, N12115, N1340, N2640, N9488);
nor NOR4 (N12118, N12098, N8861, N2842, N4929);
or OR4 (N12119, N12109, N9212, N11235, N694);
nand NAND2 (N12120, N12107, N5162);
and AND2 (N12121, N12118, N730);
xor XOR2 (N12122, N12120, N11940);
not NOT1 (N12123, N12114);
not NOT1 (N12124, N12104);
nand NAND2 (N12125, N12119, N4460);
or OR4 (N12126, N12122, N11310, N3088, N5580);
nand NAND2 (N12127, N12111, N324);
nor NOR2 (N12128, N12124, N3990);
and AND3 (N12129, N12105, N903, N11795);
not NOT1 (N12130, N12116);
nor NOR3 (N12131, N12117, N9578, N5178);
and AND4 (N12132, N12130, N4124, N7707, N2463);
not NOT1 (N12133, N12129);
and AND2 (N12134, N12131, N6049);
buf BUF1 (N12135, N12125);
nor NOR3 (N12136, N12135, N89, N9225);
nor NOR4 (N12137, N12123, N9145, N3947, N2821);
not NOT1 (N12138, N12113);
nor NOR3 (N12139, N12126, N7447, N10508);
and AND3 (N12140, N12139, N7337, N1880);
and AND4 (N12141, N12127, N9312, N9741, N1788);
buf BUF1 (N12142, N12133);
buf BUF1 (N12143, N12134);
or OR2 (N12144, N12138, N9084);
and AND2 (N12145, N12121, N8512);
and AND4 (N12146, N12145, N4142, N10158, N870);
and AND3 (N12147, N12137, N2874, N1922);
xor XOR2 (N12148, N12128, N10358);
nand NAND3 (N12149, N12136, N4839, N1150);
xor XOR2 (N12150, N12148, N5643);
buf BUF1 (N12151, N12141);
not NOT1 (N12152, N12149);
xor XOR2 (N12153, N12150, N319);
or OR4 (N12154, N12153, N5652, N3849, N6679);
and AND3 (N12155, N12152, N10567, N5259);
nor NOR3 (N12156, N12146, N486, N749);
and AND2 (N12157, N12132, N1220);
and AND3 (N12158, N12151, N1244, N1104);
nor NOR4 (N12159, N12140, N4790, N10185, N9485);
buf BUF1 (N12160, N12158);
and AND4 (N12161, N12159, N5658, N5224, N10345);
not NOT1 (N12162, N12156);
or OR4 (N12163, N12155, N7811, N7964, N2305);
buf BUF1 (N12164, N12160);
nor NOR3 (N12165, N12163, N9463, N2562);
or OR3 (N12166, N12161, N3508, N2682);
xor XOR2 (N12167, N12144, N6354);
buf BUF1 (N12168, N12162);
buf BUF1 (N12169, N12142);
nand NAND3 (N12170, N12168, N11165, N11892);
nor NOR2 (N12171, N12169, N6145);
and AND2 (N12172, N12164, N8226);
and AND2 (N12173, N12165, N4571);
buf BUF1 (N12174, N12154);
xor XOR2 (N12175, N12166, N4807);
nand NAND3 (N12176, N12171, N3595, N9840);
xor XOR2 (N12177, N12147, N2895);
nor NOR2 (N12178, N12174, N3717);
buf BUF1 (N12179, N12157);
not NOT1 (N12180, N12177);
not NOT1 (N12181, N12143);
buf BUF1 (N12182, N12173);
nor NOR3 (N12183, N12182, N10858, N8558);
not NOT1 (N12184, N12179);
and AND3 (N12185, N12175, N4834, N11462);
nor NOR3 (N12186, N12176, N11003, N2592);
buf BUF1 (N12187, N12180);
buf BUF1 (N12188, N12178);
nand NAND3 (N12189, N12187, N3783, N4403);
not NOT1 (N12190, N12183);
xor XOR2 (N12191, N12181, N1147);
or OR3 (N12192, N12189, N7824, N1071);
xor XOR2 (N12193, N12184, N85);
nand NAND2 (N12194, N12167, N2432);
nor NOR2 (N12195, N12185, N7855);
xor XOR2 (N12196, N12170, N7671);
buf BUF1 (N12197, N12196);
and AND4 (N12198, N12190, N5638, N11510, N9136);
buf BUF1 (N12199, N12191);
not NOT1 (N12200, N12192);
not NOT1 (N12201, N12199);
nor NOR3 (N12202, N12200, N2001, N4466);
nor NOR3 (N12203, N12188, N5995, N2164);
nor NOR2 (N12204, N12198, N5406);
and AND4 (N12205, N12186, N10100, N9247, N6621);
or OR2 (N12206, N12205, N2934);
or OR3 (N12207, N12172, N3332, N11146);
or OR3 (N12208, N12207, N9337, N8162);
or OR3 (N12209, N12197, N10976, N11015);
buf BUF1 (N12210, N12201);
not NOT1 (N12211, N12202);
nand NAND3 (N12212, N12209, N8175, N694);
nor NOR3 (N12213, N12193, N10562, N1856);
not NOT1 (N12214, N12203);
buf BUF1 (N12215, N12208);
not NOT1 (N12216, N12206);
or OR4 (N12217, N12214, N466, N41, N3772);
not NOT1 (N12218, N12213);
and AND2 (N12219, N12217, N8066);
nor NOR3 (N12220, N12210, N9111, N11292);
and AND4 (N12221, N12220, N11310, N592, N10194);
xor XOR2 (N12222, N12195, N7018);
nand NAND4 (N12223, N12212, N7614, N8535, N643);
or OR2 (N12224, N12219, N11874);
nand NAND4 (N12225, N12223, N11416, N7445, N4884);
buf BUF1 (N12226, N12225);
or OR3 (N12227, N12226, N7101, N4556);
or OR4 (N12228, N12215, N1746, N9484, N155);
not NOT1 (N12229, N12224);
buf BUF1 (N12230, N12218);
nand NAND3 (N12231, N12227, N3414, N5266);
buf BUF1 (N12232, N12204);
buf BUF1 (N12233, N12194);
buf BUF1 (N12234, N12233);
nand NAND3 (N12235, N12232, N11626, N7850);
and AND4 (N12236, N12228, N6638, N1993, N6837);
nand NAND2 (N12237, N12235, N7133);
nand NAND2 (N12238, N12231, N9446);
buf BUF1 (N12239, N12237);
nand NAND4 (N12240, N12211, N6133, N11285, N4928);
or OR4 (N12241, N12236, N8187, N6670, N5252);
or OR3 (N12242, N12239, N1756, N10672);
buf BUF1 (N12243, N12221);
xor XOR2 (N12244, N12230, N5145);
not NOT1 (N12245, N12234);
not NOT1 (N12246, N12244);
and AND3 (N12247, N12229, N7034, N4358);
nand NAND3 (N12248, N12216, N3602, N6774);
xor XOR2 (N12249, N12242, N6287);
nand NAND2 (N12250, N12247, N9779);
or OR4 (N12251, N12241, N6063, N1045, N6590);
buf BUF1 (N12252, N12243);
nor NOR4 (N12253, N12252, N4931, N2669, N9801);
nor NOR4 (N12254, N12248, N1479, N1960, N10235);
not NOT1 (N12255, N12238);
xor XOR2 (N12256, N12255, N11477);
nand NAND2 (N12257, N12240, N4288);
or OR4 (N12258, N12250, N723, N2843, N7576);
not NOT1 (N12259, N12253);
xor XOR2 (N12260, N12249, N8844);
nor NOR2 (N12261, N12245, N11787);
and AND4 (N12262, N12261, N11064, N7568, N7251);
xor XOR2 (N12263, N12254, N9253);
nor NOR4 (N12264, N12262, N12169, N3574, N4054);
not NOT1 (N12265, N12222);
or OR3 (N12266, N12251, N7540, N7082);
not NOT1 (N12267, N12256);
nand NAND4 (N12268, N12264, N7323, N7165, N3366);
xor XOR2 (N12269, N12260, N11640);
nand NAND4 (N12270, N12269, N1211, N6184, N10365);
or OR2 (N12271, N12258, N8154);
buf BUF1 (N12272, N12246);
nand NAND4 (N12273, N12272, N1295, N7769, N9864);
not NOT1 (N12274, N12268);
xor XOR2 (N12275, N12270, N499);
and AND4 (N12276, N12259, N1030, N4475, N11924);
and AND4 (N12277, N12265, N5917, N9732, N5537);
or OR3 (N12278, N12267, N7196, N1406);
not NOT1 (N12279, N12257);
xor XOR2 (N12280, N12274, N6063);
or OR4 (N12281, N12278, N3126, N7426, N1982);
or OR4 (N12282, N12280, N7891, N10690, N11609);
not NOT1 (N12283, N12282);
nand NAND4 (N12284, N12281, N4873, N6894, N10719);
or OR3 (N12285, N12266, N4032, N2768);
xor XOR2 (N12286, N12285, N6687);
or OR3 (N12287, N12283, N2047, N9691);
xor XOR2 (N12288, N12275, N356);
nand NAND4 (N12289, N12273, N11533, N5104, N5524);
and AND4 (N12290, N12277, N4446, N10658, N4289);
xor XOR2 (N12291, N12288, N8311);
not NOT1 (N12292, N12287);
xor XOR2 (N12293, N12290, N8167);
nand NAND3 (N12294, N12293, N9920, N4879);
buf BUF1 (N12295, N12292);
not NOT1 (N12296, N12263);
nand NAND2 (N12297, N12271, N3951);
nor NOR3 (N12298, N12297, N11625, N2242);
not NOT1 (N12299, N12294);
or OR2 (N12300, N12276, N3056);
xor XOR2 (N12301, N12286, N3917);
xor XOR2 (N12302, N12289, N9290);
or OR4 (N12303, N12301, N12205, N845, N388);
buf BUF1 (N12304, N12300);
nand NAND4 (N12305, N12295, N1231, N3418, N3317);
nand NAND2 (N12306, N12304, N7595);
buf BUF1 (N12307, N12302);
buf BUF1 (N12308, N12284);
or OR4 (N12309, N12308, N8060, N9735, N12178);
xor XOR2 (N12310, N12303, N12185);
nor NOR3 (N12311, N12291, N330, N11305);
buf BUF1 (N12312, N12310);
not NOT1 (N12313, N12311);
and AND2 (N12314, N12296, N2901);
nand NAND4 (N12315, N12309, N10237, N6579, N4842);
or OR3 (N12316, N12279, N10409, N7308);
nand NAND3 (N12317, N12315, N7368, N11993);
nand NAND3 (N12318, N12316, N6627, N11790);
and AND2 (N12319, N12306, N4021);
xor XOR2 (N12320, N12312, N1229);
not NOT1 (N12321, N12298);
buf BUF1 (N12322, N12299);
buf BUF1 (N12323, N12314);
buf BUF1 (N12324, N12319);
buf BUF1 (N12325, N12324);
not NOT1 (N12326, N12323);
buf BUF1 (N12327, N12305);
or OR4 (N12328, N12325, N10358, N7574, N11247);
xor XOR2 (N12329, N12313, N12162);
and AND2 (N12330, N12318, N3681);
and AND4 (N12331, N12317, N4542, N7638, N2061);
nor NOR2 (N12332, N12322, N1697);
not NOT1 (N12333, N12330);
xor XOR2 (N12334, N12320, N2164);
xor XOR2 (N12335, N12332, N12301);
or OR3 (N12336, N12335, N965, N2401);
xor XOR2 (N12337, N12329, N10602);
not NOT1 (N12338, N12333);
or OR3 (N12339, N12338, N8960, N9296);
or OR2 (N12340, N12337, N7256);
nand NAND2 (N12341, N12326, N4096);
nand NAND3 (N12342, N12341, N4474, N2985);
and AND4 (N12343, N12321, N12342, N11949, N199);
buf BUF1 (N12344, N1596);
buf BUF1 (N12345, N12344);
buf BUF1 (N12346, N12343);
xor XOR2 (N12347, N12334, N4120);
not NOT1 (N12348, N12336);
not NOT1 (N12349, N12339);
or OR2 (N12350, N12328, N10041);
or OR3 (N12351, N12347, N11624, N704);
nand NAND2 (N12352, N12340, N5986);
nand NAND4 (N12353, N12351, N1467, N5713, N2540);
xor XOR2 (N12354, N12346, N2966);
or OR4 (N12355, N12345, N12347, N5882, N286);
nand NAND3 (N12356, N12353, N9107, N8344);
nor NOR4 (N12357, N12307, N12194, N5733, N4180);
nand NAND4 (N12358, N12357, N5691, N6197, N10592);
not NOT1 (N12359, N12349);
and AND4 (N12360, N12354, N10588, N6472, N11470);
or OR2 (N12361, N12352, N4203);
nand NAND2 (N12362, N12356, N12062);
xor XOR2 (N12363, N12359, N9276);
nor NOR3 (N12364, N12362, N5852, N11351);
nor NOR4 (N12365, N12350, N10242, N9477, N8820);
nor NOR3 (N12366, N12331, N4233, N3691);
not NOT1 (N12367, N12360);
nand NAND2 (N12368, N12348, N11106);
or OR2 (N12369, N12365, N2270);
buf BUF1 (N12370, N12368);
xor XOR2 (N12371, N12367, N3756);
xor XOR2 (N12372, N12369, N2006);
or OR2 (N12373, N12364, N2733);
not NOT1 (N12374, N12372);
xor XOR2 (N12375, N12363, N4305);
nor NOR3 (N12376, N12361, N2321, N1234);
not NOT1 (N12377, N12370);
buf BUF1 (N12378, N12376);
not NOT1 (N12379, N12371);
nand NAND3 (N12380, N12379, N12019, N2366);
or OR3 (N12381, N12380, N894, N8496);
or OR4 (N12382, N12377, N9726, N4423, N773);
nand NAND3 (N12383, N12355, N7062, N4760);
or OR2 (N12384, N12375, N11149);
nor NOR2 (N12385, N12381, N11226);
and AND3 (N12386, N12373, N6939, N10423);
nor NOR2 (N12387, N12382, N6685);
buf BUF1 (N12388, N12327);
not NOT1 (N12389, N12387);
buf BUF1 (N12390, N12385);
nor NOR2 (N12391, N12374, N2560);
not NOT1 (N12392, N12378);
buf BUF1 (N12393, N12389);
xor XOR2 (N12394, N12383, N6652);
not NOT1 (N12395, N12384);
xor XOR2 (N12396, N12388, N9203);
nand NAND4 (N12397, N12396, N2496, N8859, N12357);
or OR3 (N12398, N12366, N649, N7032);
nor NOR3 (N12399, N12393, N6107, N1499);
and AND4 (N12400, N12397, N8178, N9883, N8046);
nor NOR2 (N12401, N12395, N8764);
nand NAND2 (N12402, N12401, N6428);
buf BUF1 (N12403, N12399);
not NOT1 (N12404, N12386);
not NOT1 (N12405, N12390);
or OR3 (N12406, N12403, N10873, N10415);
xor XOR2 (N12407, N12392, N1019);
or OR4 (N12408, N12404, N6991, N4542, N11192);
nand NAND2 (N12409, N12407, N4604);
or OR3 (N12410, N12391, N5185, N899);
nor NOR4 (N12411, N12402, N6049, N9002, N10758);
not NOT1 (N12412, N12405);
buf BUF1 (N12413, N12411);
or OR3 (N12414, N12400, N4545, N1990);
not NOT1 (N12415, N12408);
and AND2 (N12416, N12409, N1316);
nor NOR2 (N12417, N12358, N4723);
not NOT1 (N12418, N12410);
and AND4 (N12419, N12398, N5408, N10313, N2692);
and AND4 (N12420, N12416, N5933, N4067, N957);
xor XOR2 (N12421, N12406, N7339);
xor XOR2 (N12422, N12415, N7811);
not NOT1 (N12423, N12421);
nand NAND4 (N12424, N12418, N9640, N12154, N4784);
nand NAND2 (N12425, N12423, N531);
buf BUF1 (N12426, N12414);
or OR4 (N12427, N12422, N1238, N2213, N7285);
or OR2 (N12428, N12425, N10857);
nor NOR4 (N12429, N12394, N12023, N10467, N7255);
nor NOR3 (N12430, N12413, N7551, N11600);
xor XOR2 (N12431, N12428, N1871);
or OR3 (N12432, N12430, N10002, N4606);
or OR2 (N12433, N12424, N6232);
or OR2 (N12434, N12412, N4231);
nor NOR4 (N12435, N12420, N9417, N4645, N9177);
nand NAND2 (N12436, N12435, N5574);
buf BUF1 (N12437, N12436);
buf BUF1 (N12438, N12431);
not NOT1 (N12439, N12427);
nand NAND4 (N12440, N12437, N4228, N5791, N4682);
not NOT1 (N12441, N12417);
nor NOR4 (N12442, N12426, N6370, N11810, N11024);
not NOT1 (N12443, N12419);
or OR2 (N12444, N12433, N1283);
buf BUF1 (N12445, N12442);
xor XOR2 (N12446, N12445, N12110);
and AND2 (N12447, N12438, N7648);
buf BUF1 (N12448, N12429);
xor XOR2 (N12449, N12440, N8424);
or OR3 (N12450, N12434, N1316, N3824);
or OR2 (N12451, N12450, N12411);
buf BUF1 (N12452, N12432);
xor XOR2 (N12453, N12452, N6173);
and AND3 (N12454, N12453, N6839, N8907);
xor XOR2 (N12455, N12451, N394);
and AND3 (N12456, N12454, N3296, N100);
nor NOR3 (N12457, N12443, N11762, N10112);
nor NOR2 (N12458, N12455, N6748);
xor XOR2 (N12459, N12439, N5180);
xor XOR2 (N12460, N12459, N7113);
and AND4 (N12461, N12446, N3735, N12449, N4812);
xor XOR2 (N12462, N3061, N11149);
nor NOR3 (N12463, N12458, N11035, N8686);
or OR2 (N12464, N12463, N3873);
nor NOR4 (N12465, N12448, N4343, N776, N866);
xor XOR2 (N12466, N12456, N7717);
or OR2 (N12467, N12457, N6154);
nor NOR2 (N12468, N12447, N4527);
buf BUF1 (N12469, N12461);
nor NOR2 (N12470, N12464, N11554);
nand NAND3 (N12471, N12465, N3195, N581);
nor NOR4 (N12472, N12441, N1480, N3562, N9628);
or OR2 (N12473, N12467, N147);
buf BUF1 (N12474, N12462);
and AND3 (N12475, N12471, N12140, N5335);
xor XOR2 (N12476, N12469, N5566);
nand NAND3 (N12477, N12476, N2854, N11994);
nand NAND4 (N12478, N12470, N4566, N2668, N121);
buf BUF1 (N12479, N12474);
nor NOR4 (N12480, N12472, N618, N6758, N3005);
buf BUF1 (N12481, N12475);
nand NAND2 (N12482, N12473, N7258);
xor XOR2 (N12483, N12444, N6230);
or OR2 (N12484, N12468, N11774);
xor XOR2 (N12485, N12466, N2839);
nand NAND4 (N12486, N12482, N2917, N8131, N3342);
and AND3 (N12487, N12485, N4049, N11770);
not NOT1 (N12488, N12483);
not NOT1 (N12489, N12484);
or OR2 (N12490, N12460, N7256);
and AND4 (N12491, N12488, N2112, N6018, N444);
xor XOR2 (N12492, N12481, N2117);
or OR3 (N12493, N12479, N10144, N5133);
nand NAND4 (N12494, N12490, N2248, N10835, N6222);
not NOT1 (N12495, N12489);
nor NOR2 (N12496, N12491, N2470);
not NOT1 (N12497, N12496);
nand NAND3 (N12498, N12495, N6539, N2604);
and AND4 (N12499, N12478, N8769, N2726, N11644);
buf BUF1 (N12500, N12493);
not NOT1 (N12501, N12492);
xor XOR2 (N12502, N12486, N1401);
or OR3 (N12503, N12477, N12126, N2185);
nand NAND3 (N12504, N12499, N4571, N2941);
buf BUF1 (N12505, N12503);
nor NOR4 (N12506, N12487, N229, N9918, N12473);
not NOT1 (N12507, N12501);
nand NAND2 (N12508, N12498, N3876);
xor XOR2 (N12509, N12506, N3020);
xor XOR2 (N12510, N12508, N6016);
nor NOR2 (N12511, N12494, N11499);
buf BUF1 (N12512, N12504);
nor NOR4 (N12513, N12512, N11856, N2317, N4269);
not NOT1 (N12514, N12507);
nand NAND3 (N12515, N12500, N11223, N6156);
xor XOR2 (N12516, N12511, N4673);
nand NAND2 (N12517, N12513, N4764);
not NOT1 (N12518, N12480);
not NOT1 (N12519, N12505);
buf BUF1 (N12520, N12516);
nor NOR4 (N12521, N12510, N1296, N10579, N790);
or OR3 (N12522, N12521, N1577, N1829);
xor XOR2 (N12523, N12519, N7804);
or OR3 (N12524, N12518, N1002, N1952);
nand NAND2 (N12525, N12497, N6825);
not NOT1 (N12526, N12522);
and AND3 (N12527, N12524, N7725, N6294);
not NOT1 (N12528, N12509);
nand NAND3 (N12529, N12515, N8444, N9774);
or OR3 (N12530, N12502, N10387, N5374);
and AND3 (N12531, N12525, N6192, N5991);
buf BUF1 (N12532, N12531);
or OR3 (N12533, N12528, N8782, N10591);
nor NOR4 (N12534, N12533, N11801, N2580, N11447);
nor NOR4 (N12535, N12532, N9237, N5788, N10155);
or OR3 (N12536, N12520, N2223, N10312);
xor XOR2 (N12537, N12517, N10307);
or OR3 (N12538, N12535, N2331, N8885);
or OR2 (N12539, N12523, N9983);
not NOT1 (N12540, N12537);
nand NAND2 (N12541, N12530, N5421);
and AND2 (N12542, N12539, N7744);
and AND2 (N12543, N12514, N1234);
xor XOR2 (N12544, N12538, N10945);
nand NAND2 (N12545, N12529, N12186);
or OR4 (N12546, N12545, N3680, N4462, N302);
not NOT1 (N12547, N12541);
not NOT1 (N12548, N12542);
xor XOR2 (N12549, N12527, N2056);
buf BUF1 (N12550, N12549);
not NOT1 (N12551, N12547);
not NOT1 (N12552, N12544);
and AND3 (N12553, N12543, N2539, N7774);
and AND2 (N12554, N12534, N5579);
xor XOR2 (N12555, N12553, N12546);
not NOT1 (N12556, N11604);
or OR4 (N12557, N12550, N15, N9831, N3096);
nand NAND2 (N12558, N12555, N7467);
xor XOR2 (N12559, N12554, N7799);
and AND4 (N12560, N12526, N12109, N2137, N2988);
nor NOR4 (N12561, N12551, N1021, N11825, N9423);
buf BUF1 (N12562, N12558);
nor NOR3 (N12563, N12552, N7719, N5554);
and AND3 (N12564, N12536, N4426, N11044);
or OR2 (N12565, N12557, N8530);
and AND4 (N12566, N12559, N9301, N10019, N6752);
buf BUF1 (N12567, N12556);
nand NAND4 (N12568, N12563, N8682, N1020, N9971);
not NOT1 (N12569, N12562);
or OR4 (N12570, N12560, N660, N8606, N2668);
buf BUF1 (N12571, N12561);
not NOT1 (N12572, N12571);
nand NAND4 (N12573, N12568, N12107, N8286, N9919);
xor XOR2 (N12574, N12573, N5683);
xor XOR2 (N12575, N12567, N11941);
and AND3 (N12576, N12574, N5139, N963);
or OR2 (N12577, N12566, N8543);
nand NAND2 (N12578, N12569, N11164);
xor XOR2 (N12579, N12565, N4162);
and AND3 (N12580, N12575, N7979, N7298);
or OR2 (N12581, N12577, N5980);
xor XOR2 (N12582, N12572, N134);
not NOT1 (N12583, N12564);
buf BUF1 (N12584, N12582);
nand NAND3 (N12585, N12540, N7563, N2884);
nor NOR4 (N12586, N12584, N2158, N6167, N8070);
not NOT1 (N12587, N12581);
not NOT1 (N12588, N12570);
not NOT1 (N12589, N12587);
and AND4 (N12590, N12583, N4405, N4629, N6626);
buf BUF1 (N12591, N12578);
nand NAND2 (N12592, N12591, N11888);
xor XOR2 (N12593, N12585, N3278);
nor NOR4 (N12594, N12580, N12076, N398, N9064);
not NOT1 (N12595, N12590);
not NOT1 (N12596, N12593);
or OR4 (N12597, N12594, N11525, N9145, N8971);
nand NAND3 (N12598, N12588, N9714, N8676);
nor NOR2 (N12599, N12597, N1038);
buf BUF1 (N12600, N12579);
not NOT1 (N12601, N12586);
and AND4 (N12602, N12601, N4404, N12282, N7869);
nand NAND4 (N12603, N12592, N8880, N3280, N2714);
buf BUF1 (N12604, N12602);
and AND3 (N12605, N12598, N1757, N11268);
not NOT1 (N12606, N12576);
or OR3 (N12607, N12596, N6673, N10415);
xor XOR2 (N12608, N12607, N5226);
nand NAND2 (N12609, N12605, N12134);
nor NOR2 (N12610, N12600, N4871);
not NOT1 (N12611, N12606);
nand NAND4 (N12612, N12608, N2113, N9699, N2779);
not NOT1 (N12613, N12548);
or OR4 (N12614, N12611, N660, N2340, N9657);
nor NOR2 (N12615, N12609, N10958);
xor XOR2 (N12616, N12589, N6283);
nor NOR2 (N12617, N12612, N8747);
not NOT1 (N12618, N12610);
or OR2 (N12619, N12599, N521);
xor XOR2 (N12620, N12619, N2795);
or OR4 (N12621, N12613, N10209, N11805, N6063);
xor XOR2 (N12622, N12618, N8526);
nand NAND3 (N12623, N12603, N9953, N4024);
buf BUF1 (N12624, N12615);
xor XOR2 (N12625, N12595, N6063);
buf BUF1 (N12626, N12604);
not NOT1 (N12627, N12624);
and AND2 (N12628, N12627, N9272);
nor NOR3 (N12629, N12626, N9353, N9006);
xor XOR2 (N12630, N12621, N3018);
buf BUF1 (N12631, N12617);
nand NAND2 (N12632, N12631, N8359);
nand NAND3 (N12633, N12614, N979, N5280);
not NOT1 (N12634, N12620);
or OR4 (N12635, N12634, N3604, N3135, N8186);
and AND3 (N12636, N12632, N10283, N8517);
or OR2 (N12637, N12628, N11686);
buf BUF1 (N12638, N12625);
nand NAND4 (N12639, N12623, N2212, N12021, N4421);
nand NAND4 (N12640, N12633, N6160, N4665, N7012);
buf BUF1 (N12641, N12639);
xor XOR2 (N12642, N12629, N9740);
not NOT1 (N12643, N12636);
and AND2 (N12644, N12630, N21);
or OR3 (N12645, N12635, N9522, N2754);
not NOT1 (N12646, N12637);
and AND2 (N12647, N12616, N5440);
buf BUF1 (N12648, N12644);
or OR2 (N12649, N12642, N11391);
or OR3 (N12650, N12640, N4792, N1419);
or OR4 (N12651, N12650, N149, N4414, N8838);
xor XOR2 (N12652, N12647, N12472);
or OR4 (N12653, N12622, N10129, N10678, N4372);
xor XOR2 (N12654, N12651, N7704);
buf BUF1 (N12655, N12652);
or OR3 (N12656, N12655, N4702, N5032);
buf BUF1 (N12657, N12653);
or OR2 (N12658, N12656, N6986);
or OR3 (N12659, N12657, N3704, N61);
not NOT1 (N12660, N12645);
nor NOR2 (N12661, N12646, N2767);
not NOT1 (N12662, N12641);
buf BUF1 (N12663, N12661);
or OR4 (N12664, N12638, N4939, N1284, N7709);
xor XOR2 (N12665, N12648, N7309);
and AND4 (N12666, N12663, N9055, N193, N1081);
and AND3 (N12667, N12665, N1034, N3325);
buf BUF1 (N12668, N12660);
or OR3 (N12669, N12667, N2278, N2689);
or OR3 (N12670, N12662, N4939, N9066);
xor XOR2 (N12671, N12659, N11967);
or OR2 (N12672, N12670, N7154);
nor NOR4 (N12673, N12671, N2177, N11094, N5794);
xor XOR2 (N12674, N12672, N2267);
not NOT1 (N12675, N12669);
and AND4 (N12676, N12666, N10622, N6996, N8081);
nor NOR2 (N12677, N12664, N5113);
or OR3 (N12678, N12654, N1223, N1363);
nor NOR2 (N12679, N12678, N3799);
buf BUF1 (N12680, N12676);
nand NAND2 (N12681, N12674, N1860);
nor NOR4 (N12682, N12675, N1251, N3586, N7205);
nand NAND3 (N12683, N12681, N760, N576);
buf BUF1 (N12684, N12680);
nand NAND3 (N12685, N12684, N4043, N5130);
or OR4 (N12686, N12683, N3557, N2544, N5314);
nand NAND4 (N12687, N12668, N900, N2387, N12469);
nand NAND2 (N12688, N12643, N12260);
or OR2 (N12689, N12687, N5085);
and AND3 (N12690, N12658, N7359, N8930);
or OR3 (N12691, N12679, N11415, N4373);
or OR4 (N12692, N12690, N10116, N9911, N4659);
xor XOR2 (N12693, N12682, N10814);
xor XOR2 (N12694, N12673, N11036);
nor NOR4 (N12695, N12688, N4692, N7133, N5377);
nand NAND4 (N12696, N12689, N9815, N2624, N10112);
not NOT1 (N12697, N12685);
not NOT1 (N12698, N12692);
or OR4 (N12699, N12694, N2130, N7942, N6448);
xor XOR2 (N12700, N12649, N8789);
xor XOR2 (N12701, N12697, N4967);
xor XOR2 (N12702, N12695, N1382);
and AND3 (N12703, N12702, N6596, N12003);
nand NAND4 (N12704, N12703, N941, N12032, N7445);
xor XOR2 (N12705, N12700, N6365);
buf BUF1 (N12706, N12696);
nand NAND2 (N12707, N12705, N9693);
and AND2 (N12708, N12701, N4843);
and AND2 (N12709, N12704, N3484);
buf BUF1 (N12710, N12693);
and AND4 (N12711, N12677, N2590, N9363, N189);
or OR2 (N12712, N12686, N4495);
xor XOR2 (N12713, N12707, N5760);
nor NOR2 (N12714, N12706, N4821);
or OR3 (N12715, N12710, N3488, N4904);
and AND4 (N12716, N12698, N1596, N6473, N6506);
nand NAND4 (N12717, N12708, N2739, N12004, N10633);
xor XOR2 (N12718, N12699, N6674);
nor NOR2 (N12719, N12709, N3310);
or OR3 (N12720, N12713, N6946, N1628);
buf BUF1 (N12721, N12691);
nor NOR4 (N12722, N12714, N12251, N11806, N5078);
and AND3 (N12723, N12716, N9556, N2986);
nor NOR2 (N12724, N12721, N800);
or OR3 (N12725, N12719, N10435, N1009);
xor XOR2 (N12726, N12711, N699);
nand NAND2 (N12727, N12726, N8553);
not NOT1 (N12728, N12725);
nand NAND2 (N12729, N12724, N7923);
nand NAND3 (N12730, N12718, N10997, N8946);
or OR2 (N12731, N12723, N6638);
or OR3 (N12732, N12722, N984, N7636);
nor NOR2 (N12733, N12729, N5983);
not NOT1 (N12734, N12717);
nand NAND2 (N12735, N12712, N6368);
not NOT1 (N12736, N12731);
or OR4 (N12737, N12736, N2504, N7727, N7256);
xor XOR2 (N12738, N12733, N8816);
not NOT1 (N12739, N12715);
xor XOR2 (N12740, N12738, N1205);
nand NAND3 (N12741, N12732, N9389, N11984);
not NOT1 (N12742, N12740);
not NOT1 (N12743, N12734);
xor XOR2 (N12744, N12728, N1848);
nor NOR4 (N12745, N12742, N4972, N7166, N2623);
nor NOR4 (N12746, N12737, N9039, N11932, N5354);
nand NAND2 (N12747, N12739, N8951);
buf BUF1 (N12748, N12747);
buf BUF1 (N12749, N12745);
buf BUF1 (N12750, N12735);
buf BUF1 (N12751, N12746);
or OR2 (N12752, N12720, N9530);
and AND2 (N12753, N12730, N9101);
nand NAND3 (N12754, N12744, N233, N12303);
and AND2 (N12755, N12751, N3455);
nor NOR2 (N12756, N12752, N1294);
nor NOR4 (N12757, N12756, N1682, N9689, N7491);
xor XOR2 (N12758, N12743, N6141);
buf BUF1 (N12759, N12755);
or OR3 (N12760, N12748, N12735, N7054);
and AND3 (N12761, N12760, N7092, N5679);
or OR3 (N12762, N12749, N11, N11984);
xor XOR2 (N12763, N12758, N3652);
nand NAND3 (N12764, N12761, N584, N11339);
not NOT1 (N12765, N12762);
xor XOR2 (N12766, N12741, N8064);
and AND2 (N12767, N12763, N7939);
xor XOR2 (N12768, N12757, N12107);
or OR4 (N12769, N12768, N2416, N2340, N3044);
or OR4 (N12770, N12750, N6981, N11354, N4866);
buf BUF1 (N12771, N12753);
and AND2 (N12772, N12771, N6390);
buf BUF1 (N12773, N12754);
and AND4 (N12774, N12769, N6032, N4921, N2971);
nand NAND2 (N12775, N12764, N12418);
buf BUF1 (N12776, N12770);
or OR4 (N12777, N12727, N5104, N7188, N7834);
nand NAND2 (N12778, N12776, N553);
and AND4 (N12779, N12775, N3788, N12490, N7056);
buf BUF1 (N12780, N12767);
nor NOR2 (N12781, N12765, N864);
nor NOR4 (N12782, N12779, N8414, N8436, N371);
and AND4 (N12783, N12782, N4493, N4015, N10374);
nor NOR2 (N12784, N12780, N10081);
buf BUF1 (N12785, N12778);
nor NOR4 (N12786, N12785, N10514, N8748, N3301);
or OR2 (N12787, N12773, N8716);
buf BUF1 (N12788, N12766);
not NOT1 (N12789, N12788);
and AND4 (N12790, N12789, N11839, N11723, N6208);
or OR4 (N12791, N12772, N6357, N8889, N3970);
or OR3 (N12792, N12784, N9847, N477);
xor XOR2 (N12793, N12777, N323);
or OR2 (N12794, N12774, N5676);
or OR4 (N12795, N12792, N5012, N9996, N6118);
nand NAND4 (N12796, N12781, N10272, N6645, N8954);
xor XOR2 (N12797, N12786, N10233);
not NOT1 (N12798, N12794);
and AND3 (N12799, N12759, N12583, N3634);
buf BUF1 (N12800, N12799);
buf BUF1 (N12801, N12800);
buf BUF1 (N12802, N12797);
nor NOR3 (N12803, N12801, N4007, N80);
and AND2 (N12804, N12793, N4958);
xor XOR2 (N12805, N12798, N2661);
not NOT1 (N12806, N12803);
xor XOR2 (N12807, N12802, N3686);
xor XOR2 (N12808, N12804, N8075);
nor NOR3 (N12809, N12787, N8815, N2252);
or OR3 (N12810, N12809, N6495, N10055);
buf BUF1 (N12811, N12806);
and AND4 (N12812, N12791, N5314, N8519, N3037);
or OR3 (N12813, N12808, N1426, N12208);
nand NAND2 (N12814, N12812, N5174);
not NOT1 (N12815, N12810);
or OR3 (N12816, N12807, N7309, N12549);
not NOT1 (N12817, N12783);
nor NOR4 (N12818, N12790, N1152, N3400, N164);
or OR4 (N12819, N12795, N8843, N11468, N11906);
nand NAND4 (N12820, N12818, N12559, N3270, N11703);
or OR2 (N12821, N12819, N1077);
not NOT1 (N12822, N12816);
xor XOR2 (N12823, N12814, N2202);
not NOT1 (N12824, N12813);
buf BUF1 (N12825, N12823);
or OR4 (N12826, N12817, N6025, N9215, N2038);
xor XOR2 (N12827, N12811, N6345);
and AND3 (N12828, N12815, N542, N1891);
buf BUF1 (N12829, N12805);
or OR3 (N12830, N12820, N1531, N2850);
xor XOR2 (N12831, N12829, N2388);
and AND2 (N12832, N12821, N6369);
xor XOR2 (N12833, N12827, N11780);
or OR2 (N12834, N12796, N11714);
buf BUF1 (N12835, N12831);
xor XOR2 (N12836, N12830, N963);
or OR2 (N12837, N12834, N5225);
buf BUF1 (N12838, N12837);
nand NAND3 (N12839, N12824, N9663, N11788);
xor XOR2 (N12840, N12836, N5504);
or OR4 (N12841, N12832, N6035, N6666, N9424);
xor XOR2 (N12842, N12835, N3969);
nand NAND3 (N12843, N12840, N5088, N11613);
xor XOR2 (N12844, N12838, N12779);
nor NOR2 (N12845, N12844, N7002);
or OR2 (N12846, N12822, N5488);
xor XOR2 (N12847, N12841, N7611);
not NOT1 (N12848, N12839);
xor XOR2 (N12849, N12846, N11359);
xor XOR2 (N12850, N12825, N75);
nand NAND4 (N12851, N12850, N3806, N10243, N10840);
nor NOR4 (N12852, N12845, N9161, N11510, N7605);
not NOT1 (N12853, N12847);
nor NOR2 (N12854, N12849, N5379);
or OR2 (N12855, N12842, N2384);
or OR2 (N12856, N12855, N8354);
xor XOR2 (N12857, N12833, N12552);
nor NOR4 (N12858, N12854, N5696, N7169, N2456);
or OR3 (N12859, N12857, N3305, N12078);
or OR4 (N12860, N12856, N2087, N10316, N9011);
nor NOR2 (N12861, N12828, N10863);
xor XOR2 (N12862, N12851, N9699);
xor XOR2 (N12863, N12853, N6911);
or OR4 (N12864, N12863, N3569, N370, N6193);
xor XOR2 (N12865, N12862, N8077);
xor XOR2 (N12866, N12864, N8505);
xor XOR2 (N12867, N12848, N2703);
buf BUF1 (N12868, N12867);
nor NOR4 (N12869, N12859, N11281, N10644, N9247);
xor XOR2 (N12870, N12861, N1043);
xor XOR2 (N12871, N12870, N11902);
nor NOR4 (N12872, N12826, N3085, N4274, N7552);
and AND2 (N12873, N12860, N2872);
and AND2 (N12874, N12869, N914);
or OR4 (N12875, N12866, N7514, N55, N12870);
nand NAND3 (N12876, N12873, N102, N12469);
nor NOR2 (N12877, N12876, N1612);
not NOT1 (N12878, N12865);
not NOT1 (N12879, N12871);
xor XOR2 (N12880, N12878, N10994);
or OR3 (N12881, N12872, N108, N3688);
or OR3 (N12882, N12877, N745, N418);
or OR3 (N12883, N12868, N4286, N9120);
nand NAND4 (N12884, N12883, N12478, N12471, N9756);
nor NOR4 (N12885, N12875, N12660, N1667, N8187);
nand NAND4 (N12886, N12858, N6984, N7922, N1087);
not NOT1 (N12887, N12881);
xor XOR2 (N12888, N12843, N10773);
and AND3 (N12889, N12888, N5180, N8005);
or OR3 (N12890, N12874, N6041, N3705);
buf BUF1 (N12891, N12885);
buf BUF1 (N12892, N12880);
not NOT1 (N12893, N12882);
nor NOR3 (N12894, N12893, N10450, N1470);
nand NAND4 (N12895, N12884, N4756, N10687, N11644);
nor NOR4 (N12896, N12891, N10323, N10522, N3639);
xor XOR2 (N12897, N12886, N6469);
and AND3 (N12898, N12896, N4520, N6494);
buf BUF1 (N12899, N12852);
xor XOR2 (N12900, N12889, N11138);
buf BUF1 (N12901, N12898);
and AND3 (N12902, N12901, N10200, N12363);
not NOT1 (N12903, N12895);
and AND3 (N12904, N12890, N6277, N5569);
and AND2 (N12905, N12897, N11699);
xor XOR2 (N12906, N12904, N4683);
not NOT1 (N12907, N12905);
or OR3 (N12908, N12894, N3704, N10615);
buf BUF1 (N12909, N12906);
nor NOR3 (N12910, N12900, N3200, N11787);
and AND3 (N12911, N12899, N6683, N4157);
not NOT1 (N12912, N12909);
not NOT1 (N12913, N12892);
and AND3 (N12914, N12910, N7103, N4788);
or OR4 (N12915, N12912, N8385, N3768, N10317);
not NOT1 (N12916, N12915);
or OR3 (N12917, N12911, N4682, N3544);
buf BUF1 (N12918, N12902);
nor NOR4 (N12919, N12913, N1561, N3045, N1448);
xor XOR2 (N12920, N12903, N9454);
not NOT1 (N12921, N12919);
not NOT1 (N12922, N12918);
and AND4 (N12923, N12920, N11445, N9235, N2210);
buf BUF1 (N12924, N12917);
and AND3 (N12925, N12908, N1273, N2021);
not NOT1 (N12926, N12887);
not NOT1 (N12927, N12924);
nor NOR2 (N12928, N12879, N12);
and AND2 (N12929, N12928, N11790);
nand NAND3 (N12930, N12921, N1600, N3591);
buf BUF1 (N12931, N12914);
and AND3 (N12932, N12931, N115, N2572);
nor NOR4 (N12933, N12929, N8434, N3394, N8996);
nor NOR2 (N12934, N12930, N3856);
and AND2 (N12935, N12907, N5908);
or OR4 (N12936, N12925, N11869, N5690, N3054);
not NOT1 (N12937, N12936);
xor XOR2 (N12938, N12934, N5305);
nand NAND3 (N12939, N12922, N9592, N2146);
or OR4 (N12940, N12938, N5623, N6443, N9722);
and AND4 (N12941, N12933, N3852, N10555, N10852);
buf BUF1 (N12942, N12937);
buf BUF1 (N12943, N12923);
nor NOR4 (N12944, N12916, N12126, N2050, N9670);
nor NOR4 (N12945, N12941, N11899, N9712, N8609);
not NOT1 (N12946, N12935);
xor XOR2 (N12947, N12939, N11254);
or OR4 (N12948, N12932, N8202, N7578, N11945);
buf BUF1 (N12949, N12926);
nor NOR3 (N12950, N12948, N6173, N4785);
nor NOR4 (N12951, N12949, N2504, N5210, N10808);
nand NAND2 (N12952, N12944, N8456);
or OR2 (N12953, N12945, N7574);
and AND4 (N12954, N12927, N8103, N788, N11617);
not NOT1 (N12955, N12946);
xor XOR2 (N12956, N12954, N4043);
and AND4 (N12957, N12940, N4107, N2741, N10733);
nor NOR4 (N12958, N12956, N11, N4296, N652);
buf BUF1 (N12959, N12951);
xor XOR2 (N12960, N12950, N1616);
and AND3 (N12961, N12943, N594, N9248);
not NOT1 (N12962, N12942);
buf BUF1 (N12963, N12962);
nor NOR4 (N12964, N12963, N3623, N10559, N8729);
xor XOR2 (N12965, N12960, N7234);
buf BUF1 (N12966, N12964);
or OR2 (N12967, N12959, N11005);
buf BUF1 (N12968, N12955);
or OR4 (N12969, N12967, N4019, N5002, N2277);
nor NOR2 (N12970, N12952, N10593);
nand NAND3 (N12971, N12966, N14, N3401);
or OR4 (N12972, N12957, N5238, N10212, N4679);
not NOT1 (N12973, N12971);
not NOT1 (N12974, N12969);
nor NOR3 (N12975, N12970, N7745, N973);
nor NOR3 (N12976, N12973, N4947, N8832);
or OR3 (N12977, N12968, N9939, N252);
and AND2 (N12978, N12965, N7889);
buf BUF1 (N12979, N12976);
not NOT1 (N12980, N12972);
nand NAND4 (N12981, N12980, N11443, N1489, N2592);
and AND3 (N12982, N12978, N1848, N10307);
and AND4 (N12983, N12953, N3293, N10505, N12162);
nand NAND2 (N12984, N12974, N11914);
xor XOR2 (N12985, N12979, N486);
or OR3 (N12986, N12947, N4504, N7093);
buf BUF1 (N12987, N12983);
not NOT1 (N12988, N12984);
or OR4 (N12989, N12981, N2663, N5562, N8278);
nor NOR2 (N12990, N12975, N5523);
and AND4 (N12991, N12987, N4726, N2467, N12090);
nand NAND4 (N12992, N12977, N10016, N10020, N1567);
not NOT1 (N12993, N12990);
not NOT1 (N12994, N12992);
nor NOR4 (N12995, N12958, N2117, N2504, N11329);
not NOT1 (N12996, N12993);
or OR4 (N12997, N12991, N1242, N7501, N633);
xor XOR2 (N12998, N12997, N3898);
not NOT1 (N12999, N12989);
not NOT1 (N13000, N12994);
buf BUF1 (N13001, N13000);
nand NAND2 (N13002, N12998, N4355);
not NOT1 (N13003, N12985);
not NOT1 (N13004, N12995);
or OR2 (N13005, N13002, N9122);
or OR2 (N13006, N12986, N12012);
or OR2 (N13007, N13001, N11324);
xor XOR2 (N13008, N12988, N4865);
not NOT1 (N13009, N12999);
nand NAND4 (N13010, N12961, N5740, N2206, N10885);
buf BUF1 (N13011, N13004);
xor XOR2 (N13012, N13010, N2565);
or OR2 (N13013, N12982, N12868);
and AND3 (N13014, N13008, N5268, N11577);
nand NAND4 (N13015, N13011, N6721, N1427, N2578);
nor NOR3 (N13016, N13007, N166, N11229);
xor XOR2 (N13017, N13013, N11107);
xor XOR2 (N13018, N13017, N6834);
not NOT1 (N13019, N13016);
nand NAND4 (N13020, N13005, N8626, N3293, N12709);
nor NOR3 (N13021, N13009, N10788, N2234);
nor NOR2 (N13022, N13006, N8385);
not NOT1 (N13023, N13012);
nand NAND2 (N13024, N13015, N11905);
and AND3 (N13025, N13020, N8222, N6619);
or OR4 (N13026, N13018, N7044, N2989, N2210);
or OR2 (N13027, N13025, N7589);
buf BUF1 (N13028, N13003);
nor NOR2 (N13029, N13024, N5659);
nand NAND3 (N13030, N13027, N5196, N6671);
buf BUF1 (N13031, N13014);
nor NOR4 (N13032, N13031, N12145, N687, N7441);
or OR3 (N13033, N13026, N7777, N3647);
buf BUF1 (N13034, N13029);
nor NOR3 (N13035, N13022, N11077, N558);
nand NAND4 (N13036, N13021, N9926, N6751, N3947);
xor XOR2 (N13037, N13030, N11486);
and AND3 (N13038, N13037, N11131, N4248);
and AND4 (N13039, N13038, N7486, N6692, N8773);
and AND4 (N13040, N13036, N11440, N9179, N8097);
nor NOR3 (N13041, N13019, N12285, N6886);
nand NAND2 (N13042, N13032, N11178);
xor XOR2 (N13043, N13041, N11158);
not NOT1 (N13044, N13028);
nor NOR2 (N13045, N13035, N1463);
not NOT1 (N13046, N13045);
and AND3 (N13047, N13046, N12518, N2590);
or OR2 (N13048, N13034, N7099);
nand NAND4 (N13049, N13044, N2261, N12745, N11124);
xor XOR2 (N13050, N13033, N9140);
nor NOR3 (N13051, N12996, N1470, N3813);
or OR4 (N13052, N13023, N1795, N99, N12715);
and AND4 (N13053, N13050, N12073, N4706, N3018);
or OR2 (N13054, N13043, N6365);
or OR4 (N13055, N13039, N9255, N10533, N1516);
xor XOR2 (N13056, N13052, N4387);
and AND4 (N13057, N13051, N12050, N11345, N4318);
and AND4 (N13058, N13040, N249, N7876, N3513);
nand NAND2 (N13059, N13055, N6433);
or OR3 (N13060, N13049, N7472, N2788);
nand NAND3 (N13061, N13048, N11164, N12658);
or OR2 (N13062, N13057, N2394);
or OR4 (N13063, N13059, N12311, N10089, N12230);
and AND3 (N13064, N13047, N12661, N4220);
not NOT1 (N13065, N13061);
nor NOR3 (N13066, N13053, N5294, N1442);
xor XOR2 (N13067, N13066, N5329);
not NOT1 (N13068, N13062);
nor NOR2 (N13069, N13056, N7080);
or OR4 (N13070, N13058, N5275, N6712, N2139);
xor XOR2 (N13071, N13042, N347);
xor XOR2 (N13072, N13064, N6496);
xor XOR2 (N13073, N13069, N10034);
or OR4 (N13074, N13072, N12123, N5530, N5718);
not NOT1 (N13075, N13060);
or OR2 (N13076, N13075, N11141);
and AND2 (N13077, N13074, N3920);
or OR3 (N13078, N13054, N6791, N12251);
not NOT1 (N13079, N13073);
xor XOR2 (N13080, N13068, N11898);
nor NOR2 (N13081, N13063, N12790);
or OR2 (N13082, N13079, N10567);
not NOT1 (N13083, N13080);
nor NOR3 (N13084, N13067, N2992, N8995);
nand NAND3 (N13085, N13082, N5216, N6471);
xor XOR2 (N13086, N13076, N2037);
xor XOR2 (N13087, N13083, N8133);
or OR2 (N13088, N13081, N353);
nand NAND3 (N13089, N13087, N8298, N1232);
or OR4 (N13090, N13089, N7836, N3328, N5972);
nor NOR4 (N13091, N13071, N703, N12869, N3133);
not NOT1 (N13092, N13085);
or OR4 (N13093, N13090, N3666, N8622, N4738);
not NOT1 (N13094, N13077);
or OR4 (N13095, N13092, N3576, N4432, N498);
buf BUF1 (N13096, N13094);
nand NAND3 (N13097, N13095, N6659, N11464);
not NOT1 (N13098, N13088);
xor XOR2 (N13099, N13070, N4047);
xor XOR2 (N13100, N13098, N4951);
not NOT1 (N13101, N13086);
and AND2 (N13102, N13101, N8129);
nand NAND2 (N13103, N13097, N10348);
or OR3 (N13104, N13100, N6439, N11866);
not NOT1 (N13105, N13078);
nand NAND4 (N13106, N13099, N428, N7434, N3044);
not NOT1 (N13107, N13091);
and AND4 (N13108, N13065, N7248, N1060, N4822);
buf BUF1 (N13109, N13106);
xor XOR2 (N13110, N13096, N4867);
nor NOR3 (N13111, N13104, N5065, N5535);
xor XOR2 (N13112, N13107, N10769);
nand NAND3 (N13113, N13110, N11100, N5872);
nand NAND4 (N13114, N13084, N2608, N12105, N3858);
buf BUF1 (N13115, N13108);
or OR2 (N13116, N13105, N4595);
and AND2 (N13117, N13116, N9203);
and AND3 (N13118, N13109, N10849, N10266);
nor NOR2 (N13119, N13114, N1585);
or OR3 (N13120, N13093, N9577, N8206);
or OR4 (N13121, N13111, N6956, N11227, N6408);
nand NAND3 (N13122, N13118, N10641, N2744);
not NOT1 (N13123, N13102);
not NOT1 (N13124, N13123);
xor XOR2 (N13125, N13122, N6775);
nand NAND3 (N13126, N13125, N2214, N6196);
and AND2 (N13127, N13113, N7005);
buf BUF1 (N13128, N13127);
buf BUF1 (N13129, N13126);
and AND3 (N13130, N13121, N6580, N12033);
xor XOR2 (N13131, N13119, N6401);
nand NAND3 (N13132, N13131, N6273, N690);
nor NOR3 (N13133, N13115, N4234, N10788);
or OR4 (N13134, N13117, N10653, N6325, N12696);
not NOT1 (N13135, N13133);
not NOT1 (N13136, N13130);
xor XOR2 (N13137, N13103, N2017);
not NOT1 (N13138, N13128);
nand NAND2 (N13139, N13138, N9450);
buf BUF1 (N13140, N13132);
not NOT1 (N13141, N13120);
not NOT1 (N13142, N13140);
nor NOR3 (N13143, N13112, N8758, N11300);
and AND2 (N13144, N13136, N11884);
not NOT1 (N13145, N13144);
not NOT1 (N13146, N13143);
or OR3 (N13147, N13129, N2943, N4467);
and AND2 (N13148, N13134, N895);
nor NOR2 (N13149, N13142, N60);
or OR2 (N13150, N13141, N12496);
and AND3 (N13151, N13147, N4486, N8005);
not NOT1 (N13152, N13145);
nor NOR4 (N13153, N13148, N4542, N2559, N1836);
not NOT1 (N13154, N13146);
not NOT1 (N13155, N13139);
not NOT1 (N13156, N13154);
xor XOR2 (N13157, N13149, N9371);
or OR4 (N13158, N13135, N6442, N11138, N3520);
nor NOR3 (N13159, N13150, N10996, N9780);
nand NAND2 (N13160, N13159, N12455);
nand NAND4 (N13161, N13152, N10244, N4807, N4651);
xor XOR2 (N13162, N13153, N9189);
buf BUF1 (N13163, N13160);
and AND2 (N13164, N13137, N9973);
and AND2 (N13165, N13124, N10071);
buf BUF1 (N13166, N13162);
nor NOR2 (N13167, N13163, N10426);
nor NOR4 (N13168, N13166, N9618, N9742, N10990);
nand NAND4 (N13169, N13151, N7285, N5362, N12554);
nor NOR3 (N13170, N13165, N10249, N13068);
not NOT1 (N13171, N13155);
and AND2 (N13172, N13168, N10990);
nand NAND4 (N13173, N13157, N4334, N8715, N8571);
nand NAND4 (N13174, N13167, N8021, N1097, N3826);
buf BUF1 (N13175, N13158);
not NOT1 (N13176, N13156);
buf BUF1 (N13177, N13175);
not NOT1 (N13178, N13176);
nand NAND2 (N13179, N13169, N7875);
not NOT1 (N13180, N13173);
nand NAND2 (N13181, N13178, N9305);
and AND4 (N13182, N13177, N11301, N10840, N7465);
or OR3 (N13183, N13170, N13156, N2916);
buf BUF1 (N13184, N13180);
or OR3 (N13185, N13181, N9315, N192);
and AND4 (N13186, N13184, N5569, N2965, N1603);
buf BUF1 (N13187, N13185);
nor NOR4 (N13188, N13183, N4503, N1983, N4955);
buf BUF1 (N13189, N13179);
xor XOR2 (N13190, N13171, N2685);
and AND4 (N13191, N13187, N435, N10923, N288);
not NOT1 (N13192, N13188);
xor XOR2 (N13193, N13174, N10247);
nand NAND3 (N13194, N13190, N10845, N6214);
and AND2 (N13195, N13164, N9423);
buf BUF1 (N13196, N13182);
nor NOR4 (N13197, N13196, N8222, N7371, N11182);
nand NAND4 (N13198, N13194, N11076, N8022, N7229);
nor NOR3 (N13199, N13198, N3520, N12095);
or OR2 (N13200, N13186, N792);
nand NAND2 (N13201, N13191, N12989);
and AND2 (N13202, N13161, N6598);
and AND2 (N13203, N13172, N11532);
and AND4 (N13204, N13192, N11201, N7936, N8586);
and AND3 (N13205, N13199, N12784, N1490);
not NOT1 (N13206, N13195);
and AND4 (N13207, N13201, N11499, N454, N7779);
buf BUF1 (N13208, N13202);
or OR2 (N13209, N13193, N3260);
nor NOR2 (N13210, N13208, N9302);
or OR3 (N13211, N13205, N8658, N11353);
nand NAND4 (N13212, N13206, N1944, N2497, N3246);
not NOT1 (N13213, N13207);
not NOT1 (N13214, N13210);
nor NOR2 (N13215, N13214, N10637);
and AND2 (N13216, N13204, N786);
not NOT1 (N13217, N13200);
nor NOR3 (N13218, N13203, N1708, N9585);
not NOT1 (N13219, N13216);
not NOT1 (N13220, N13215);
xor XOR2 (N13221, N13217, N6162);
nor NOR2 (N13222, N13220, N3012);
or OR4 (N13223, N13213, N11751, N10751, N856);
nand NAND4 (N13224, N13209, N5397, N226, N13180);
not NOT1 (N13225, N13222);
nor NOR2 (N13226, N13211, N235);
and AND2 (N13227, N13224, N8332);
and AND3 (N13228, N13227, N6360, N9645);
and AND4 (N13229, N13226, N6774, N839, N9630);
or OR4 (N13230, N13219, N882, N9397, N12131);
and AND3 (N13231, N13212, N11026, N12925);
and AND2 (N13232, N13230, N2876);
or OR3 (N13233, N13197, N11372, N893);
nor NOR3 (N13234, N13189, N666, N4508);
nor NOR2 (N13235, N13232, N11022);
buf BUF1 (N13236, N13231);
not NOT1 (N13237, N13234);
or OR2 (N13238, N13221, N9125);
xor XOR2 (N13239, N13236, N2634);
buf BUF1 (N13240, N13228);
xor XOR2 (N13241, N13229, N11598);
buf BUF1 (N13242, N13240);
buf BUF1 (N13243, N13241);
xor XOR2 (N13244, N13225, N4692);
or OR3 (N13245, N13239, N307, N586);
nor NOR3 (N13246, N13218, N1191, N4093);
xor XOR2 (N13247, N13237, N10445);
nor NOR2 (N13248, N13233, N11703);
buf BUF1 (N13249, N13247);
xor XOR2 (N13250, N13242, N7520);
xor XOR2 (N13251, N13223, N446);
nand NAND4 (N13252, N13243, N12946, N9233, N13043);
or OR4 (N13253, N13252, N1512, N8154, N7925);
xor XOR2 (N13254, N13235, N6439);
or OR3 (N13255, N13238, N3336, N1961);
buf BUF1 (N13256, N13254);
nor NOR2 (N13257, N13249, N7529);
not NOT1 (N13258, N13255);
nand NAND3 (N13259, N13251, N1209, N9570);
xor XOR2 (N13260, N13244, N6021);
xor XOR2 (N13261, N13260, N7590);
and AND2 (N13262, N13246, N6755);
or OR2 (N13263, N13253, N5215);
buf BUF1 (N13264, N13261);
and AND2 (N13265, N13245, N5073);
xor XOR2 (N13266, N13258, N8328);
and AND4 (N13267, N13248, N10358, N7182, N6160);
and AND4 (N13268, N13264, N180, N4539, N9552);
buf BUF1 (N13269, N13268);
nor NOR2 (N13270, N13256, N10622);
not NOT1 (N13271, N13262);
not NOT1 (N13272, N13271);
not NOT1 (N13273, N13269);
not NOT1 (N13274, N13266);
nor NOR4 (N13275, N13273, N5087, N12966, N6546);
nand NAND2 (N13276, N13263, N2170);
xor XOR2 (N13277, N13265, N12335);
nor NOR3 (N13278, N13267, N6557, N12012);
or OR3 (N13279, N13270, N2706, N3640);
xor XOR2 (N13280, N13279, N11507);
not NOT1 (N13281, N13280);
and AND3 (N13282, N13272, N11340, N3621);
or OR2 (N13283, N13274, N13215);
nand NAND4 (N13284, N13277, N10988, N11818, N1613);
and AND3 (N13285, N13259, N2556, N272);
nand NAND3 (N13286, N13278, N2635, N7095);
nand NAND3 (N13287, N13283, N1440, N10445);
nand NAND4 (N13288, N13287, N12868, N2810, N2310);
not NOT1 (N13289, N13281);
or OR4 (N13290, N13275, N11897, N3178, N10115);
and AND4 (N13291, N13284, N6332, N7201, N1196);
not NOT1 (N13292, N13289);
xor XOR2 (N13293, N13292, N3721);
or OR4 (N13294, N13250, N216, N11743, N973);
buf BUF1 (N13295, N13294);
buf BUF1 (N13296, N13295);
and AND2 (N13297, N13282, N88);
and AND2 (N13298, N13293, N4249);
or OR2 (N13299, N13291, N9878);
nand NAND2 (N13300, N13285, N992);
xor XOR2 (N13301, N13288, N7247);
or OR3 (N13302, N13299, N12490, N10835);
nand NAND3 (N13303, N13300, N3378, N7627);
xor XOR2 (N13304, N13298, N3681);
nand NAND3 (N13305, N13290, N11580, N8825);
xor XOR2 (N13306, N13301, N8050);
and AND3 (N13307, N13296, N4101, N5382);
nor NOR2 (N13308, N13286, N7774);
not NOT1 (N13309, N13305);
nand NAND2 (N13310, N13297, N2920);
nand NAND2 (N13311, N13257, N13092);
or OR2 (N13312, N13306, N324);
not NOT1 (N13313, N13311);
or OR2 (N13314, N13308, N4560);
not NOT1 (N13315, N13276);
xor XOR2 (N13316, N13313, N11634);
nand NAND3 (N13317, N13302, N9099, N2972);
or OR2 (N13318, N13309, N12978);
xor XOR2 (N13319, N13318, N12410);
not NOT1 (N13320, N13316);
buf BUF1 (N13321, N13304);
nand NAND2 (N13322, N13315, N4353);
nor NOR2 (N13323, N13321, N3946);
and AND2 (N13324, N13303, N12128);
or OR3 (N13325, N13312, N1653, N8028);
not NOT1 (N13326, N13307);
not NOT1 (N13327, N13324);
or OR3 (N13328, N13319, N9637, N10044);
or OR3 (N13329, N13327, N9743, N11170);
buf BUF1 (N13330, N13326);
xor XOR2 (N13331, N13325, N12296);
xor XOR2 (N13332, N13328, N11004);
buf BUF1 (N13333, N13331);
xor XOR2 (N13334, N13332, N1094);
xor XOR2 (N13335, N13330, N6754);
nand NAND3 (N13336, N13320, N7553, N3122);
nor NOR3 (N13337, N13336, N13172, N1766);
xor XOR2 (N13338, N13333, N3901);
and AND4 (N13339, N13329, N7178, N4792, N501);
buf BUF1 (N13340, N13314);
nor NOR3 (N13341, N13322, N7613, N9351);
buf BUF1 (N13342, N13335);
or OR2 (N13343, N13334, N9801);
not NOT1 (N13344, N13339);
or OR2 (N13345, N13338, N7118);
buf BUF1 (N13346, N13344);
buf BUF1 (N13347, N13337);
nor NOR3 (N13348, N13347, N12601, N1568);
and AND4 (N13349, N13342, N8811, N4556, N5596);
nor NOR2 (N13350, N13345, N13135);
and AND2 (N13351, N13340, N7270);
xor XOR2 (N13352, N13310, N6574);
xor XOR2 (N13353, N13352, N8942);
and AND2 (N13354, N13346, N11803);
xor XOR2 (N13355, N13341, N1520);
or OR2 (N13356, N13355, N4731);
nand NAND2 (N13357, N13323, N6313);
nand NAND3 (N13358, N13356, N6356, N9704);
xor XOR2 (N13359, N13351, N887);
nand NAND3 (N13360, N13354, N6125, N5416);
or OR3 (N13361, N13358, N8590, N959);
xor XOR2 (N13362, N13343, N2067);
not NOT1 (N13363, N13359);
xor XOR2 (N13364, N13349, N2782);
or OR3 (N13365, N13350, N7883, N3042);
nor NOR2 (N13366, N13348, N8375);
nor NOR2 (N13367, N13357, N2559);
and AND3 (N13368, N13361, N1457, N10009);
or OR3 (N13369, N13317, N3068, N12741);
nor NOR4 (N13370, N13353, N8339, N501, N11140);
xor XOR2 (N13371, N13362, N9135);
not NOT1 (N13372, N13367);
and AND2 (N13373, N13366, N4556);
not NOT1 (N13374, N13370);
or OR3 (N13375, N13368, N7629, N3881);
and AND2 (N13376, N13364, N6914);
xor XOR2 (N13377, N13363, N12312);
nor NOR2 (N13378, N13377, N2873);
or OR4 (N13379, N13374, N1642, N10121, N1175);
buf BUF1 (N13380, N13365);
not NOT1 (N13381, N13372);
nand NAND4 (N13382, N13379, N11336, N4789, N5751);
nand NAND4 (N13383, N13371, N8856, N643, N858);
or OR4 (N13384, N13376, N8898, N10884, N13244);
not NOT1 (N13385, N13378);
buf BUF1 (N13386, N13373);
not NOT1 (N13387, N13360);
and AND3 (N13388, N13381, N3167, N10216);
xor XOR2 (N13389, N13369, N13242);
buf BUF1 (N13390, N13386);
and AND3 (N13391, N13389, N13166, N615);
xor XOR2 (N13392, N13391, N7263);
buf BUF1 (N13393, N13388);
or OR2 (N13394, N13392, N5281);
nor NOR2 (N13395, N13394, N10096);
nor NOR4 (N13396, N13385, N1450, N3412, N11691);
buf BUF1 (N13397, N13375);
nand NAND3 (N13398, N13393, N1840, N5056);
buf BUF1 (N13399, N13396);
nor NOR2 (N13400, N13390, N3165);
buf BUF1 (N13401, N13380);
not NOT1 (N13402, N13384);
not NOT1 (N13403, N13400);
or OR3 (N13404, N13399, N7236, N2321);
and AND4 (N13405, N13398, N7943, N9995, N4123);
or OR4 (N13406, N13402, N3499, N9159, N6978);
nand NAND2 (N13407, N13395, N1789);
xor XOR2 (N13408, N13404, N6565);
nand NAND3 (N13409, N13397, N2258, N5295);
and AND4 (N13410, N13403, N7326, N2499, N7165);
and AND4 (N13411, N13408, N10522, N13203, N9294);
or OR2 (N13412, N13409, N3248);
xor XOR2 (N13413, N13411, N10110);
xor XOR2 (N13414, N13407, N5819);
or OR4 (N13415, N13387, N9435, N2106, N5097);
buf BUF1 (N13416, N13406);
xor XOR2 (N13417, N13410, N11180);
nor NOR2 (N13418, N13412, N541);
nand NAND3 (N13419, N13405, N7232, N11325);
or OR4 (N13420, N13419, N10545, N5731, N1584);
not NOT1 (N13421, N13416);
and AND4 (N13422, N13401, N5817, N7236, N726);
buf BUF1 (N13423, N13383);
xor XOR2 (N13424, N13415, N3118);
nor NOR2 (N13425, N13418, N13150);
not NOT1 (N13426, N13413);
xor XOR2 (N13427, N13422, N7663);
xor XOR2 (N13428, N13382, N1779);
and AND3 (N13429, N13426, N13197, N4714);
xor XOR2 (N13430, N13420, N10967);
or OR3 (N13431, N13429, N4014, N2123);
and AND3 (N13432, N13417, N6904, N10809);
or OR2 (N13433, N13430, N10124);
buf BUF1 (N13434, N13424);
nand NAND3 (N13435, N13427, N8331, N6247);
buf BUF1 (N13436, N13428);
nor NOR3 (N13437, N13435, N12223, N4261);
and AND4 (N13438, N13431, N2687, N2045, N10160);
or OR2 (N13439, N13414, N4703);
buf BUF1 (N13440, N13437);
and AND3 (N13441, N13434, N10851, N393);
nand NAND4 (N13442, N13421, N5470, N116, N4067);
buf BUF1 (N13443, N13438);
or OR3 (N13444, N13425, N680, N3037);
nor NOR2 (N13445, N13432, N12234);
or OR4 (N13446, N13443, N9915, N7302, N4373);
buf BUF1 (N13447, N13444);
nand NAND3 (N13448, N13423, N3271, N7791);
and AND4 (N13449, N13436, N11316, N3026, N10751);
not NOT1 (N13450, N13449);
or OR3 (N13451, N13446, N1477, N10214);
xor XOR2 (N13452, N13433, N8758);
not NOT1 (N13453, N13452);
nor NOR2 (N13454, N13439, N8760);
and AND2 (N13455, N13440, N624);
or OR2 (N13456, N13441, N12845);
buf BUF1 (N13457, N13454);
nand NAND2 (N13458, N13450, N8711);
buf BUF1 (N13459, N13445);
buf BUF1 (N13460, N13448);
or OR2 (N13461, N13456, N5688);
not NOT1 (N13462, N13458);
nor NOR4 (N13463, N13453, N12549, N3328, N9764);
or OR3 (N13464, N13460, N13270, N7912);
or OR4 (N13465, N13447, N7313, N2019, N10097);
or OR3 (N13466, N13464, N3298, N11325);
nor NOR3 (N13467, N13463, N12938, N276);
nand NAND4 (N13468, N13467, N1340, N12431, N12565);
buf BUF1 (N13469, N13451);
and AND4 (N13470, N13466, N1328, N5836, N1990);
nand NAND4 (N13471, N13455, N7063, N12150, N364);
or OR4 (N13472, N13465, N8594, N12381, N11405);
nand NAND3 (N13473, N13442, N9041, N894);
xor XOR2 (N13474, N13468, N5914);
nor NOR3 (N13475, N13473, N7232, N3725);
or OR3 (N13476, N13459, N9391, N4324);
and AND3 (N13477, N13472, N7287, N3452);
not NOT1 (N13478, N13461);
xor XOR2 (N13479, N13478, N6811);
buf BUF1 (N13480, N13457);
nor NOR2 (N13481, N13470, N860);
and AND2 (N13482, N13469, N4225);
nor NOR4 (N13483, N13480, N758, N4503, N5623);
not NOT1 (N13484, N13475);
not NOT1 (N13485, N13474);
xor XOR2 (N13486, N13479, N5550);
not NOT1 (N13487, N13486);
or OR2 (N13488, N13471, N1484);
nand NAND2 (N13489, N13485, N669);
buf BUF1 (N13490, N13481);
nand NAND2 (N13491, N13477, N11394);
nor NOR3 (N13492, N13487, N8455, N8646);
not NOT1 (N13493, N13491);
xor XOR2 (N13494, N13462, N12404);
buf BUF1 (N13495, N13494);
nor NOR2 (N13496, N13483, N3801);
buf BUF1 (N13497, N13476);
buf BUF1 (N13498, N13493);
or OR2 (N13499, N13482, N11181);
xor XOR2 (N13500, N13497, N8017);
or OR2 (N13501, N13498, N11153);
or OR2 (N13502, N13492, N11221);
or OR4 (N13503, N13500, N2159, N5088, N7830);
xor XOR2 (N13504, N13499, N3108);
nor NOR3 (N13505, N13490, N2700, N5858);
buf BUF1 (N13506, N13505);
or OR3 (N13507, N13484, N11712, N3882);
and AND3 (N13508, N13507, N1755, N33);
nand NAND3 (N13509, N13489, N6190, N897);
not NOT1 (N13510, N13506);
nand NAND4 (N13511, N13504, N2749, N5393, N9781);
xor XOR2 (N13512, N13510, N4421);
or OR3 (N13513, N13496, N10040, N10080);
xor XOR2 (N13514, N13511, N915);
buf BUF1 (N13515, N13503);
or OR2 (N13516, N13495, N10603);
nand NAND2 (N13517, N13515, N1263);
not NOT1 (N13518, N13516);
not NOT1 (N13519, N13512);
and AND2 (N13520, N13501, N2946);
nand NAND2 (N13521, N13518, N10868);
or OR3 (N13522, N13508, N7711, N1774);
nand NAND4 (N13523, N13521, N10260, N2560, N9567);
or OR3 (N13524, N13502, N1140, N11400);
nand NAND3 (N13525, N13519, N8317, N404);
nand NAND2 (N13526, N13513, N735);
and AND3 (N13527, N13523, N5520, N9984);
xor XOR2 (N13528, N13488, N523);
not NOT1 (N13529, N13522);
nor NOR3 (N13530, N13520, N8874, N7854);
xor XOR2 (N13531, N13524, N8554);
not NOT1 (N13532, N13528);
buf BUF1 (N13533, N13529);
and AND2 (N13534, N13526, N7950);
xor XOR2 (N13535, N13514, N10333);
and AND2 (N13536, N13534, N6239);
not NOT1 (N13537, N13533);
nor NOR3 (N13538, N13525, N4361, N12536);
buf BUF1 (N13539, N13509);
or OR4 (N13540, N13536, N9200, N13407, N12857);
nand NAND4 (N13541, N13530, N13257, N13535, N920);
or OR4 (N13542, N9477, N3315, N4889, N2707);
buf BUF1 (N13543, N13539);
and AND4 (N13544, N13543, N5608, N6429, N2367);
or OR2 (N13545, N13531, N11308);
nand NAND4 (N13546, N13537, N2115, N6054, N1808);
nand NAND3 (N13547, N13541, N8569, N5098);
nor NOR3 (N13548, N13547, N8297, N13053);
nor NOR4 (N13549, N13527, N2573, N12476, N9340);
xor XOR2 (N13550, N13538, N10691);
xor XOR2 (N13551, N13532, N5561);
and AND3 (N13552, N13545, N7651, N4001);
nor NOR3 (N13553, N13544, N111, N11653);
buf BUF1 (N13554, N13551);
not NOT1 (N13555, N13540);
buf BUF1 (N13556, N13554);
or OR2 (N13557, N13517, N8380);
not NOT1 (N13558, N13549);
nand NAND3 (N13559, N13546, N665, N9662);
nand NAND2 (N13560, N13555, N1413);
nor NOR2 (N13561, N13552, N13107);
buf BUF1 (N13562, N13550);
xor XOR2 (N13563, N13542, N7887);
and AND2 (N13564, N13553, N10335);
nand NAND4 (N13565, N13562, N10582, N4364, N2053);
nor NOR3 (N13566, N13560, N10197, N1923);
and AND4 (N13567, N13564, N2452, N12960, N6967);
nand NAND3 (N13568, N13557, N5817, N6794);
and AND3 (N13569, N13556, N2, N7430);
buf BUF1 (N13570, N13565);
or OR2 (N13571, N13570, N2475);
nor NOR2 (N13572, N13571, N974);
buf BUF1 (N13573, N13572);
and AND3 (N13574, N13573, N2021, N9574);
and AND4 (N13575, N13567, N9821, N7166, N10734);
xor XOR2 (N13576, N13574, N2273);
buf BUF1 (N13577, N13561);
and AND4 (N13578, N13577, N5648, N8630, N10263);
or OR4 (N13579, N13576, N1706, N11919, N8573);
xor XOR2 (N13580, N13558, N3604);
not NOT1 (N13581, N13548);
nand NAND4 (N13582, N13580, N2536, N11438, N1597);
buf BUF1 (N13583, N13568);
nor NOR4 (N13584, N13581, N9034, N10053, N3052);
or OR3 (N13585, N13583, N2802, N12260);
buf BUF1 (N13586, N13575);
not NOT1 (N13587, N13578);
not NOT1 (N13588, N13569);
xor XOR2 (N13589, N13584, N6808);
nor NOR3 (N13590, N13559, N1637, N11853);
buf BUF1 (N13591, N13589);
nor NOR2 (N13592, N13563, N3480);
xor XOR2 (N13593, N13587, N6218);
not NOT1 (N13594, N13579);
buf BUF1 (N13595, N13594);
or OR3 (N13596, N13595, N12284, N11310);
or OR3 (N13597, N13596, N5562, N8890);
buf BUF1 (N13598, N13585);
buf BUF1 (N13599, N13598);
and AND3 (N13600, N13591, N6255, N9560);
and AND4 (N13601, N13582, N1857, N476, N3950);
nand NAND4 (N13602, N13601, N12758, N2542, N9181);
buf BUF1 (N13603, N13586);
nor NOR2 (N13604, N13597, N2477);
xor XOR2 (N13605, N13590, N9517);
nand NAND4 (N13606, N13600, N5214, N4865, N10299);
and AND4 (N13607, N13566, N3386, N6035, N11426);
nand NAND2 (N13608, N13604, N8898);
nor NOR2 (N13609, N13588, N9695);
nand NAND4 (N13610, N13599, N8543, N10637, N2993);
not NOT1 (N13611, N13606);
not NOT1 (N13612, N13605);
nand NAND3 (N13613, N13607, N11466, N9062);
or OR4 (N13614, N13608, N9948, N814, N4146);
not NOT1 (N13615, N13609);
or OR2 (N13616, N13610, N9807);
buf BUF1 (N13617, N13612);
buf BUF1 (N13618, N13617);
and AND2 (N13619, N13613, N12726);
and AND2 (N13620, N13593, N4915);
xor XOR2 (N13621, N13618, N1420);
nor NOR4 (N13622, N13615, N2911, N1864, N11736);
buf BUF1 (N13623, N13621);
buf BUF1 (N13624, N13619);
or OR4 (N13625, N13624, N13200, N3304, N5165);
xor XOR2 (N13626, N13602, N10295);
and AND3 (N13627, N13616, N12927, N12379);
xor XOR2 (N13628, N13611, N8541);
not NOT1 (N13629, N13623);
or OR4 (N13630, N13627, N9724, N9759, N12146);
not NOT1 (N13631, N13630);
and AND2 (N13632, N13622, N2324);
nor NOR3 (N13633, N13603, N6927, N12771);
nor NOR3 (N13634, N13614, N9328, N4595);
not NOT1 (N13635, N13629);
not NOT1 (N13636, N13631);
buf BUF1 (N13637, N13632);
nand NAND2 (N13638, N13634, N11312);
and AND3 (N13639, N13636, N3466, N7465);
nor NOR4 (N13640, N13633, N29, N3548, N7672);
nor NOR3 (N13641, N13635, N3245, N10634);
nand NAND4 (N13642, N13637, N13345, N4407, N5397);
nand NAND3 (N13643, N13628, N11305, N13277);
xor XOR2 (N13644, N13626, N8244);
nor NOR2 (N13645, N13644, N10473);
nand NAND4 (N13646, N13642, N1693, N13604, N7417);
buf BUF1 (N13647, N13640);
or OR3 (N13648, N13638, N8230, N2259);
or OR2 (N13649, N13647, N10833);
nor NOR3 (N13650, N13639, N4026, N5981);
nand NAND2 (N13651, N13646, N72);
nand NAND4 (N13652, N13649, N7689, N7556, N6763);
nand NAND2 (N13653, N13645, N1087);
and AND4 (N13654, N13648, N7783, N2240, N12983);
or OR2 (N13655, N13641, N10048);
nand NAND2 (N13656, N13625, N1520);
buf BUF1 (N13657, N13643);
and AND3 (N13658, N13651, N3057, N8218);
nor NOR3 (N13659, N13653, N13568, N6737);
buf BUF1 (N13660, N13592);
not NOT1 (N13661, N13659);
and AND3 (N13662, N13650, N11842, N7011);
nand NAND4 (N13663, N13655, N3434, N821, N6477);
nor NOR2 (N13664, N13652, N8591);
or OR4 (N13665, N13620, N7734, N12993, N9472);
not NOT1 (N13666, N13660);
or OR4 (N13667, N13662, N8592, N8809, N9603);
nor NOR2 (N13668, N13658, N9756);
not NOT1 (N13669, N13664);
xor XOR2 (N13670, N13665, N12674);
nand NAND4 (N13671, N13654, N9650, N898, N10200);
and AND4 (N13672, N13670, N9076, N10243, N3829);
or OR3 (N13673, N13667, N11130, N9516);
xor XOR2 (N13674, N13672, N7130);
and AND3 (N13675, N13674, N13575, N3717);
not NOT1 (N13676, N13675);
nor NOR2 (N13677, N13668, N2712);
nand NAND3 (N13678, N13657, N12018, N8437);
or OR2 (N13679, N13677, N8261);
or OR2 (N13680, N13671, N13072);
nor NOR3 (N13681, N13656, N10108, N13450);
buf BUF1 (N13682, N13666);
or OR2 (N13683, N13679, N2687);
nor NOR4 (N13684, N13680, N11175, N11989, N414);
buf BUF1 (N13685, N13681);
nor NOR3 (N13686, N13682, N2237, N13110);
or OR2 (N13687, N13663, N7145);
xor XOR2 (N13688, N13686, N879);
or OR3 (N13689, N13685, N644, N707);
or OR4 (N13690, N13689, N9981, N7399, N12546);
nor NOR2 (N13691, N13687, N7167);
not NOT1 (N13692, N13673);
or OR2 (N13693, N13676, N8621);
nor NOR2 (N13694, N13669, N5082);
nor NOR3 (N13695, N13690, N1497, N4717);
not NOT1 (N13696, N13695);
nand NAND2 (N13697, N13661, N12833);
nand NAND3 (N13698, N13692, N10582, N13688);
xor XOR2 (N13699, N3439, N9508);
nand NAND3 (N13700, N13683, N3968, N3412);
not NOT1 (N13701, N13691);
nor NOR2 (N13702, N13698, N9083);
nor NOR3 (N13703, N13697, N8554, N11672);
or OR4 (N13704, N13678, N5279, N13613, N11523);
xor XOR2 (N13705, N13699, N3448);
buf BUF1 (N13706, N13694);
nand NAND4 (N13707, N13706, N992, N11365, N1175);
or OR2 (N13708, N13704, N7213);
and AND2 (N13709, N13696, N4215);
or OR4 (N13710, N13700, N7130, N5578, N4808);
and AND4 (N13711, N13710, N13125, N8002, N5299);
or OR3 (N13712, N13709, N9468, N260);
not NOT1 (N13713, N13711);
nand NAND4 (N13714, N13702, N10241, N1195, N10328);
nor NOR2 (N13715, N13713, N13098);
and AND4 (N13716, N13715, N7193, N6404, N13547);
and AND4 (N13717, N13703, N9435, N8915, N5402);
and AND4 (N13718, N13716, N3980, N859, N1995);
not NOT1 (N13719, N13707);
buf BUF1 (N13720, N13708);
xor XOR2 (N13721, N13712, N3469);
and AND2 (N13722, N13717, N6807);
nor NOR3 (N13723, N13714, N712, N6134);
buf BUF1 (N13724, N13723);
nor NOR3 (N13725, N13722, N1168, N2668);
not NOT1 (N13726, N13693);
nor NOR2 (N13727, N13684, N7872);
buf BUF1 (N13728, N13720);
or OR2 (N13729, N13726, N12024);
and AND3 (N13730, N13701, N6310, N8729);
buf BUF1 (N13731, N13727);
buf BUF1 (N13732, N13721);
buf BUF1 (N13733, N13730);
and AND2 (N13734, N13724, N4072);
and AND3 (N13735, N13705, N8123, N2894);
xor XOR2 (N13736, N13728, N13271);
nand NAND3 (N13737, N13736, N420, N12941);
xor XOR2 (N13738, N13729, N8917);
nor NOR3 (N13739, N13732, N1969, N11514);
buf BUF1 (N13740, N13735);
nor NOR2 (N13741, N13718, N2553);
nand NAND3 (N13742, N13739, N7735, N10638);
buf BUF1 (N13743, N13737);
nand NAND3 (N13744, N13734, N5791, N1038);
nor NOR4 (N13745, N13740, N13385, N189, N5532);
xor XOR2 (N13746, N13745, N3586);
and AND2 (N13747, N13746, N9910);
and AND4 (N13748, N13743, N9236, N6498, N786);
and AND3 (N13749, N13748, N10412, N10348);
nand NAND2 (N13750, N13747, N5642);
and AND4 (N13751, N13744, N2418, N3808, N4431);
nand NAND2 (N13752, N13738, N12353);
buf BUF1 (N13753, N13750);
or OR4 (N13754, N13719, N12269, N5599, N3831);
or OR4 (N13755, N13752, N6049, N6504, N12726);
not NOT1 (N13756, N13753);
nor NOR3 (N13757, N13751, N4378, N4518);
buf BUF1 (N13758, N13757);
not NOT1 (N13759, N13741);
and AND4 (N13760, N13742, N3402, N12926, N1214);
nor NOR3 (N13761, N13758, N13715, N7416);
not NOT1 (N13762, N13760);
and AND2 (N13763, N13749, N283);
xor XOR2 (N13764, N13763, N11655);
nand NAND2 (N13765, N13725, N11552);
or OR2 (N13766, N13761, N12702);
or OR4 (N13767, N13759, N872, N12969, N9888);
nand NAND4 (N13768, N13766, N1612, N11068, N12823);
xor XOR2 (N13769, N13755, N7489);
buf BUF1 (N13770, N13762);
or OR4 (N13771, N13731, N11394, N2685, N10781);
nand NAND2 (N13772, N13765, N4456);
and AND4 (N13773, N13772, N11231, N3195, N10279);
xor XOR2 (N13774, N13771, N6621);
xor XOR2 (N13775, N13767, N742);
and AND3 (N13776, N13773, N4797, N11115);
and AND2 (N13777, N13733, N266);
nor NOR2 (N13778, N13774, N10857);
and AND2 (N13779, N13775, N3071);
nand NAND4 (N13780, N13778, N3406, N5491, N4262);
not NOT1 (N13781, N13764);
nor NOR3 (N13782, N13780, N948, N4384);
buf BUF1 (N13783, N13776);
and AND4 (N13784, N13754, N3381, N3531, N8917);
not NOT1 (N13785, N13779);
and AND3 (N13786, N13785, N938, N3364);
not NOT1 (N13787, N13769);
nand NAND3 (N13788, N13786, N2338, N5977);
nor NOR4 (N13789, N13768, N13581, N8570, N12922);
and AND4 (N13790, N13789, N9083, N2653, N13550);
and AND4 (N13791, N13783, N13689, N3487, N233);
nor NOR2 (N13792, N13788, N1833);
or OR2 (N13793, N13756, N6932);
buf BUF1 (N13794, N13791);
and AND4 (N13795, N13784, N2174, N4716, N13221);
nand NAND3 (N13796, N13795, N12241, N5783);
xor XOR2 (N13797, N13777, N8277);
nand NAND2 (N13798, N13790, N6289);
nand NAND3 (N13799, N13781, N12037, N8993);
nor NOR3 (N13800, N13782, N11431, N11191);
buf BUF1 (N13801, N13794);
xor XOR2 (N13802, N13801, N13209);
buf BUF1 (N13803, N13802);
nor NOR3 (N13804, N13792, N10618, N7794);
nor NOR3 (N13805, N13787, N1642, N12125);
not NOT1 (N13806, N13798);
nand NAND2 (N13807, N13805, N4791);
xor XOR2 (N13808, N13796, N10405);
xor XOR2 (N13809, N13770, N12653);
buf BUF1 (N13810, N13804);
not NOT1 (N13811, N13807);
xor XOR2 (N13812, N13809, N1777);
nand NAND3 (N13813, N13803, N862, N1329);
not NOT1 (N13814, N13810);
buf BUF1 (N13815, N13813);
not NOT1 (N13816, N13811);
nor NOR3 (N13817, N13793, N8931, N1471);
and AND4 (N13818, N13799, N13369, N10553, N1158);
or OR3 (N13819, N13818, N7615, N5657);
buf BUF1 (N13820, N13808);
or OR4 (N13821, N13814, N3159, N5361, N5564);
not NOT1 (N13822, N13797);
nand NAND2 (N13823, N13817, N13813);
xor XOR2 (N13824, N13800, N2354);
or OR4 (N13825, N13824, N402, N3031, N11095);
nand NAND2 (N13826, N13819, N5175);
and AND2 (N13827, N13812, N2457);
or OR3 (N13828, N13826, N4069, N7082);
not NOT1 (N13829, N13816);
nand NAND3 (N13830, N13815, N8579, N8121);
nand NAND2 (N13831, N13828, N1355);
or OR2 (N13832, N13831, N13659);
not NOT1 (N13833, N13822);
nor NOR2 (N13834, N13833, N2368);
and AND3 (N13835, N13834, N4780, N13);
and AND2 (N13836, N13830, N6172);
and AND2 (N13837, N13827, N13159);
not NOT1 (N13838, N13820);
nor NOR3 (N13839, N13832, N13784, N13792);
nor NOR2 (N13840, N13823, N4151);
nand NAND2 (N13841, N13835, N8352);
not NOT1 (N13842, N13839);
not NOT1 (N13843, N13836);
xor XOR2 (N13844, N13829, N11666);
and AND3 (N13845, N13844, N13273, N3804);
not NOT1 (N13846, N13825);
nor NOR2 (N13847, N13837, N9794);
nor NOR3 (N13848, N13846, N9145, N1561);
nor NOR3 (N13849, N13848, N8634, N7844);
and AND4 (N13850, N13838, N6034, N8364, N752);
or OR2 (N13851, N13847, N3573);
or OR4 (N13852, N13849, N1888, N12289, N13482);
and AND2 (N13853, N13840, N4948);
xor XOR2 (N13854, N13851, N8481);
not NOT1 (N13855, N13853);
nor NOR2 (N13856, N13806, N6417);
xor XOR2 (N13857, N13850, N13755);
or OR4 (N13858, N13842, N3397, N1274, N13852);
xor XOR2 (N13859, N7266, N13181);
xor XOR2 (N13860, N13856, N11707);
and AND3 (N13861, N13841, N8612, N13309);
nand NAND3 (N13862, N13855, N5020, N4201);
and AND4 (N13863, N13854, N13391, N12425, N11899);
and AND2 (N13864, N13863, N10401);
not NOT1 (N13865, N13821);
buf BUF1 (N13866, N13860);
xor XOR2 (N13867, N13861, N78);
xor XOR2 (N13868, N13843, N1255);
nand NAND4 (N13869, N13866, N3106, N4757, N4631);
buf BUF1 (N13870, N13862);
buf BUF1 (N13871, N13867);
buf BUF1 (N13872, N13869);
buf BUF1 (N13873, N13871);
and AND2 (N13874, N13870, N5169);
or OR2 (N13875, N13845, N7838);
and AND2 (N13876, N13859, N3981);
xor XOR2 (N13877, N13874, N2842);
or OR4 (N13878, N13873, N10080, N11585, N3780);
nor NOR3 (N13879, N13864, N6760, N8867);
buf BUF1 (N13880, N13872);
and AND4 (N13881, N13857, N1727, N4664, N1030);
xor XOR2 (N13882, N13878, N5160);
not NOT1 (N13883, N13881);
nand NAND3 (N13884, N13880, N7212, N9503);
buf BUF1 (N13885, N13877);
buf BUF1 (N13886, N13875);
nand NAND2 (N13887, N13882, N4681);
or OR2 (N13888, N13883, N7970);
nand NAND3 (N13889, N13884, N5887, N5665);
nand NAND3 (N13890, N13858, N3570, N13580);
xor XOR2 (N13891, N13868, N5127);
buf BUF1 (N13892, N13890);
xor XOR2 (N13893, N13888, N910);
nor NOR4 (N13894, N13879, N6196, N2212, N8740);
nand NAND2 (N13895, N13893, N4340);
nand NAND4 (N13896, N13891, N12513, N2883, N8394);
and AND4 (N13897, N13896, N6853, N3785, N5838);
nor NOR3 (N13898, N13876, N6323, N13598);
nor NOR4 (N13899, N13865, N3914, N2774, N4991);
nand NAND4 (N13900, N13886, N1829, N5413, N4887);
xor XOR2 (N13901, N13897, N13647);
nor NOR4 (N13902, N13889, N6144, N9426, N11646);
buf BUF1 (N13903, N13900);
and AND2 (N13904, N13898, N5701);
nand NAND2 (N13905, N13887, N10446);
or OR3 (N13906, N13901, N12128, N12475);
nor NOR2 (N13907, N13903, N4882);
nand NAND2 (N13908, N13905, N10809);
xor XOR2 (N13909, N13892, N9387);
buf BUF1 (N13910, N13902);
and AND4 (N13911, N13885, N13457, N13504, N10449);
not NOT1 (N13912, N13910);
nand NAND3 (N13913, N13906, N2859, N2580);
and AND2 (N13914, N13909, N9835);
or OR4 (N13915, N13895, N614, N6205, N12528);
buf BUF1 (N13916, N13911);
or OR2 (N13917, N13904, N177);
or OR3 (N13918, N13912, N11521, N11601);
nor NOR3 (N13919, N13908, N10226, N13224);
nand NAND3 (N13920, N13915, N8620, N12960);
nor NOR2 (N13921, N13907, N2355);
or OR3 (N13922, N13914, N10755, N12255);
nor NOR3 (N13923, N13917, N11779, N13249);
not NOT1 (N13924, N13923);
buf BUF1 (N13925, N13922);
nand NAND4 (N13926, N13921, N11979, N6391, N13344);
nand NAND4 (N13927, N13919, N397, N6467, N11231);
buf BUF1 (N13928, N13924);
nand NAND2 (N13929, N13920, N12533);
not NOT1 (N13930, N13913);
not NOT1 (N13931, N13930);
nor NOR3 (N13932, N13927, N10144, N2295);
nor NOR4 (N13933, N13929, N407, N11802, N10741);
and AND4 (N13934, N13928, N236, N11706, N2529);
or OR4 (N13935, N13931, N11970, N4924, N9594);
buf BUF1 (N13936, N13918);
xor XOR2 (N13937, N13935, N12591);
buf BUF1 (N13938, N13933);
nor NOR2 (N13939, N13925, N10087);
or OR4 (N13940, N13899, N13070, N8375, N1604);
or OR4 (N13941, N13926, N4933, N7631, N6770);
not NOT1 (N13942, N13938);
and AND3 (N13943, N13939, N9257, N7969);
nor NOR4 (N13944, N13940, N12977, N2943, N1337);
not NOT1 (N13945, N13944);
nand NAND4 (N13946, N13934, N8390, N1036, N11214);
buf BUF1 (N13947, N13937);
nand NAND4 (N13948, N13894, N8459, N138, N4064);
nand NAND2 (N13949, N13947, N3159);
xor XOR2 (N13950, N13946, N3586);
nand NAND2 (N13951, N13948, N9547);
nand NAND3 (N13952, N13949, N7815, N11515);
xor XOR2 (N13953, N13936, N656);
buf BUF1 (N13954, N13953);
and AND2 (N13955, N13942, N10065);
or OR2 (N13956, N13916, N13695);
nand NAND2 (N13957, N13943, N3719);
or OR4 (N13958, N13932, N12896, N7132, N13489);
or OR3 (N13959, N13952, N1721, N3571);
and AND4 (N13960, N13945, N1191, N3439, N7163);
xor XOR2 (N13961, N13959, N10987);
not NOT1 (N13962, N13954);
nand NAND3 (N13963, N13962, N5152, N8891);
or OR3 (N13964, N13963, N10094, N980);
and AND4 (N13965, N13957, N5948, N5198, N10477);
not NOT1 (N13966, N13964);
nand NAND2 (N13967, N13966, N12913);
or OR2 (N13968, N13961, N4818);
xor XOR2 (N13969, N13956, N6151);
or OR3 (N13970, N13950, N3679, N2572);
not NOT1 (N13971, N13965);
xor XOR2 (N13972, N13968, N12511);
nor NOR3 (N13973, N13971, N12925, N9777);
nor NOR2 (N13974, N13967, N4660);
xor XOR2 (N13975, N13974, N3952);
buf BUF1 (N13976, N13972);
and AND2 (N13977, N13951, N12433);
and AND2 (N13978, N13941, N8956);
nor NOR2 (N13979, N13978, N2996);
buf BUF1 (N13980, N13976);
not NOT1 (N13981, N13970);
buf BUF1 (N13982, N13969);
nand NAND4 (N13983, N13960, N6265, N938, N3681);
buf BUF1 (N13984, N13981);
not NOT1 (N13985, N13980);
nand NAND3 (N13986, N13983, N10010, N6493);
buf BUF1 (N13987, N13975);
xor XOR2 (N13988, N13955, N13759);
or OR2 (N13989, N13977, N13703);
nand NAND2 (N13990, N13988, N13427);
and AND4 (N13991, N13990, N11539, N10783, N506);
not NOT1 (N13992, N13989);
or OR2 (N13993, N13982, N8431);
xor XOR2 (N13994, N13993, N7311);
and AND3 (N13995, N13986, N5092, N1884);
or OR4 (N13996, N13984, N847, N12169, N6750);
and AND4 (N13997, N13995, N8525, N8918, N8776);
nand NAND3 (N13998, N13997, N3370, N2268);
nand NAND3 (N13999, N13958, N1484, N8300);
buf BUF1 (N14000, N13979);
and AND3 (N14001, N13999, N9875, N5167);
buf BUF1 (N14002, N14001);
xor XOR2 (N14003, N13973, N2081);
nand NAND3 (N14004, N13994, N13473, N6852);
buf BUF1 (N14005, N13991);
buf BUF1 (N14006, N13987);
and AND2 (N14007, N14004, N521);
nand NAND3 (N14008, N13985, N5846, N5444);
not NOT1 (N14009, N13992);
and AND3 (N14010, N14008, N8196, N6601);
buf BUF1 (N14011, N14005);
and AND4 (N14012, N14006, N5718, N3746, N2227);
or OR4 (N14013, N14007, N10983, N4275, N13721);
xor XOR2 (N14014, N14012, N783);
xor XOR2 (N14015, N14011, N8195);
buf BUF1 (N14016, N14014);
buf BUF1 (N14017, N14015);
buf BUF1 (N14018, N14016);
or OR2 (N14019, N14003, N5341);
buf BUF1 (N14020, N14017);
and AND4 (N14021, N14002, N13607, N5350, N9792);
and AND4 (N14022, N13998, N13669, N10216, N11681);
not NOT1 (N14023, N14022);
nor NOR4 (N14024, N14023, N13630, N682, N6729);
or OR4 (N14025, N14021, N2403, N3454, N8957);
nor NOR4 (N14026, N14025, N12553, N5121, N12623);
or OR3 (N14027, N14024, N11925, N13516);
nand NAND2 (N14028, N14009, N5041);
nand NAND2 (N14029, N14018, N13176);
xor XOR2 (N14030, N14028, N7002);
nand NAND2 (N14031, N14019, N4404);
nor NOR3 (N14032, N13996, N13296, N7634);
or OR3 (N14033, N14026, N667, N11228);
buf BUF1 (N14034, N14010);
or OR2 (N14035, N14034, N9481);
xor XOR2 (N14036, N14031, N6978);
or OR4 (N14037, N14030, N7087, N4652, N9117);
xor XOR2 (N14038, N14037, N5766);
not NOT1 (N14039, N14000);
nand NAND4 (N14040, N14032, N7275, N14014, N7551);
buf BUF1 (N14041, N14040);
and AND3 (N14042, N14020, N13844, N5690);
or OR4 (N14043, N14036, N3838, N2529, N10639);
nand NAND3 (N14044, N14033, N4183, N7611);
nand NAND4 (N14045, N14035, N8421, N12074, N852);
buf BUF1 (N14046, N14038);
buf BUF1 (N14047, N14029);
nand NAND4 (N14048, N14041, N11877, N6032, N10750);
xor XOR2 (N14049, N14045, N6160);
nor NOR4 (N14050, N14013, N447, N7713, N5459);
xor XOR2 (N14051, N14050, N1512);
not NOT1 (N14052, N14039);
not NOT1 (N14053, N14042);
or OR4 (N14054, N14046, N1815, N2043, N12015);
not NOT1 (N14055, N14053);
nand NAND4 (N14056, N14049, N4114, N7099, N1876);
nor NOR2 (N14057, N14048, N7691);
not NOT1 (N14058, N14056);
xor XOR2 (N14059, N14027, N2652);
nand NAND2 (N14060, N14043, N13200);
and AND4 (N14061, N14047, N6917, N6582, N1039);
or OR2 (N14062, N14059, N2420);
not NOT1 (N14063, N14058);
not NOT1 (N14064, N14061);
xor XOR2 (N14065, N14063, N8914);
or OR3 (N14066, N14064, N1874, N6159);
xor XOR2 (N14067, N14051, N12083);
or OR2 (N14068, N14066, N7003);
and AND4 (N14069, N14054, N7831, N8503, N2465);
and AND3 (N14070, N14060, N11434, N10484);
nand NAND3 (N14071, N14052, N4905, N1377);
or OR3 (N14072, N14055, N2594, N10035);
or OR4 (N14073, N14057, N6677, N9341, N7746);
xor XOR2 (N14074, N14069, N11888);
xor XOR2 (N14075, N14071, N3247);
and AND2 (N14076, N14070, N2622);
or OR3 (N14077, N14073, N6183, N3716);
or OR4 (N14078, N14072, N180, N3236, N7426);
not NOT1 (N14079, N14065);
or OR2 (N14080, N14078, N10473);
and AND4 (N14081, N14062, N5380, N109, N2333);
nand NAND4 (N14082, N14074, N13423, N10407, N4645);
not NOT1 (N14083, N14076);
not NOT1 (N14084, N14083);
and AND3 (N14085, N14080, N6698, N2327);
nand NAND4 (N14086, N14077, N12995, N11489, N9408);
or OR2 (N14087, N14075, N10747);
nand NAND4 (N14088, N14082, N2334, N7269, N12938);
buf BUF1 (N14089, N14067);
xor XOR2 (N14090, N14088, N9263);
or OR3 (N14091, N14044, N8173, N12865);
or OR2 (N14092, N14089, N1816);
not NOT1 (N14093, N14084);
nand NAND2 (N14094, N14081, N9566);
nor NOR3 (N14095, N14085, N4792, N9665);
buf BUF1 (N14096, N14087);
not NOT1 (N14097, N14079);
not NOT1 (N14098, N14068);
nor NOR4 (N14099, N14097, N9511, N10097, N597);
nand NAND2 (N14100, N14099, N12815);
nor NOR2 (N14101, N14094, N10601);
nand NAND3 (N14102, N14096, N4416, N6962);
not NOT1 (N14103, N14102);
nor NOR4 (N14104, N14090, N13502, N69, N2331);
nand NAND4 (N14105, N14098, N9709, N11132, N5350);
buf BUF1 (N14106, N14104);
nor NOR3 (N14107, N14091, N1752, N11654);
xor XOR2 (N14108, N14095, N3833);
nand NAND4 (N14109, N14092, N12049, N11255, N12168);
or OR3 (N14110, N14100, N10838, N6241);
and AND4 (N14111, N14093, N6353, N6225, N9897);
nor NOR4 (N14112, N14106, N134, N8618, N2473);
buf BUF1 (N14113, N14110);
nand NAND3 (N14114, N14111, N12517, N2034);
xor XOR2 (N14115, N14112, N882);
nand NAND3 (N14116, N14113, N4552, N1570);
buf BUF1 (N14117, N14103);
xor XOR2 (N14118, N14116, N7240);
nand NAND2 (N14119, N14105, N502);
nor NOR2 (N14120, N14086, N12347);
not NOT1 (N14121, N14118);
nor NOR2 (N14122, N14101, N4417);
and AND4 (N14123, N14108, N9921, N8578, N12303);
xor XOR2 (N14124, N14122, N12334);
or OR3 (N14125, N14107, N1482, N11656);
xor XOR2 (N14126, N14123, N9561);
or OR3 (N14127, N14120, N11408, N13003);
and AND2 (N14128, N14126, N7817);
or OR3 (N14129, N14127, N10929, N10875);
nand NAND4 (N14130, N14109, N6938, N12132, N2750);
buf BUF1 (N14131, N14114);
nand NAND4 (N14132, N14115, N6939, N12635, N701);
not NOT1 (N14133, N14124);
nor NOR2 (N14134, N14121, N9457);
nor NOR4 (N14135, N14131, N5746, N10194, N8963);
not NOT1 (N14136, N14130);
nand NAND4 (N14137, N14128, N6458, N4791, N1886);
and AND4 (N14138, N14125, N8375, N9701, N6457);
or OR2 (N14139, N14138, N4381);
nand NAND4 (N14140, N14133, N314, N5768, N5682);
not NOT1 (N14141, N14136);
or OR2 (N14142, N14137, N10411);
or OR3 (N14143, N14119, N2041, N1965);
nand NAND4 (N14144, N14134, N13847, N12881, N9040);
buf BUF1 (N14145, N14117);
xor XOR2 (N14146, N14139, N12907);
xor XOR2 (N14147, N14144, N10366);
nor NOR3 (N14148, N14142, N12693, N4581);
nor NOR3 (N14149, N14135, N984, N11524);
nand NAND3 (N14150, N14132, N13745, N5785);
nor NOR4 (N14151, N14140, N537, N6630, N1554);
buf BUF1 (N14152, N14149);
nor NOR2 (N14153, N14152, N9905);
not NOT1 (N14154, N14141);
buf BUF1 (N14155, N14148);
or OR4 (N14156, N14146, N1496, N9198, N10153);
xor XOR2 (N14157, N14151, N11481);
buf BUF1 (N14158, N14145);
nand NAND2 (N14159, N14156, N2019);
not NOT1 (N14160, N14157);
nor NOR2 (N14161, N14160, N1019);
nand NAND4 (N14162, N14150, N7335, N1765, N1284);
buf BUF1 (N14163, N14129);
not NOT1 (N14164, N14143);
not NOT1 (N14165, N14155);
or OR3 (N14166, N14162, N12916, N11139);
or OR3 (N14167, N14147, N4207, N12450);
xor XOR2 (N14168, N14153, N8832);
and AND3 (N14169, N14158, N10280, N7508);
buf BUF1 (N14170, N14159);
and AND3 (N14171, N14154, N2546, N8402);
nand NAND3 (N14172, N14164, N7535, N3227);
nand NAND2 (N14173, N14171, N9013);
nand NAND3 (N14174, N14167, N4188, N3994);
nand NAND3 (N14175, N14169, N4157, N12244);
and AND2 (N14176, N14172, N12927);
xor XOR2 (N14177, N14174, N8593);
xor XOR2 (N14178, N14173, N7807);
xor XOR2 (N14179, N14170, N13741);
not NOT1 (N14180, N14165);
or OR3 (N14181, N14179, N6706, N4915);
not NOT1 (N14182, N14176);
not NOT1 (N14183, N14161);
nor NOR4 (N14184, N14168, N8913, N3364, N10489);
nand NAND4 (N14185, N14178, N1601, N6921, N337);
nor NOR4 (N14186, N14181, N13736, N8271, N4933);
or OR4 (N14187, N14166, N11356, N6222, N13743);
not NOT1 (N14188, N14177);
not NOT1 (N14189, N14188);
and AND4 (N14190, N14180, N9097, N10115, N11971);
xor XOR2 (N14191, N14184, N11588);
or OR3 (N14192, N14191, N6789, N6963);
xor XOR2 (N14193, N14186, N2410);
nor NOR3 (N14194, N14182, N459, N5624);
buf BUF1 (N14195, N14163);
nor NOR3 (N14196, N14175, N847, N11082);
buf BUF1 (N14197, N14183);
xor XOR2 (N14198, N14187, N1078);
xor XOR2 (N14199, N14198, N7356);
or OR3 (N14200, N14193, N1974, N12707);
nor NOR2 (N14201, N14194, N8711);
xor XOR2 (N14202, N14197, N2739);
and AND3 (N14203, N14199, N13430, N752);
nand NAND2 (N14204, N14201, N6262);
not NOT1 (N14205, N14202);
nor NOR4 (N14206, N14190, N8760, N12676, N431);
or OR3 (N14207, N14206, N4740, N2109);
nand NAND2 (N14208, N14185, N5718);
buf BUF1 (N14209, N14205);
or OR2 (N14210, N14196, N64);
buf BUF1 (N14211, N14195);
not NOT1 (N14212, N14209);
buf BUF1 (N14213, N14207);
not NOT1 (N14214, N14192);
or OR2 (N14215, N14208, N9243);
nand NAND2 (N14216, N14214, N10208);
buf BUF1 (N14217, N14210);
or OR3 (N14218, N14217, N5078, N2541);
nand NAND2 (N14219, N14216, N3234);
not NOT1 (N14220, N14213);
nand NAND2 (N14221, N14203, N12743);
or OR4 (N14222, N14220, N2580, N4968, N9784);
or OR3 (N14223, N14212, N7052, N5249);
nand NAND2 (N14224, N14215, N9562);
xor XOR2 (N14225, N14200, N13302);
and AND4 (N14226, N14222, N4175, N10458, N6737);
nor NOR2 (N14227, N14225, N6018);
not NOT1 (N14228, N14204);
or OR2 (N14229, N14227, N3893);
nand NAND4 (N14230, N14211, N8506, N13347, N11238);
buf BUF1 (N14231, N14224);
nor NOR3 (N14232, N14218, N8062, N1849);
nand NAND2 (N14233, N14231, N12779);
buf BUF1 (N14234, N14221);
buf BUF1 (N14235, N14228);
xor XOR2 (N14236, N14234, N7844);
nand NAND2 (N14237, N14233, N5225);
and AND3 (N14238, N14236, N11515, N13892);
buf BUF1 (N14239, N14226);
buf BUF1 (N14240, N14230);
not NOT1 (N14241, N14239);
nand NAND2 (N14242, N14232, N10537);
nor NOR3 (N14243, N14235, N7420, N2793);
buf BUF1 (N14244, N14241);
buf BUF1 (N14245, N14229);
buf BUF1 (N14246, N14237);
xor XOR2 (N14247, N14189, N10763);
or OR3 (N14248, N14243, N5313, N2619);
nand NAND3 (N14249, N14240, N11215, N8888);
or OR4 (N14250, N14245, N7608, N3107, N5553);
nor NOR3 (N14251, N14238, N9417, N3503);
xor XOR2 (N14252, N14248, N6589);
and AND3 (N14253, N14250, N5, N11669);
and AND4 (N14254, N14242, N4890, N6308, N14009);
and AND3 (N14255, N14219, N9857, N514);
not NOT1 (N14256, N14253);
nor NOR2 (N14257, N14246, N12489);
or OR4 (N14258, N14247, N1564, N5796, N11988);
nand NAND3 (N14259, N14249, N11747, N12818);
buf BUF1 (N14260, N14223);
xor XOR2 (N14261, N14254, N9509);
not NOT1 (N14262, N14261);
or OR3 (N14263, N14255, N8601, N8943);
not NOT1 (N14264, N14260);
nor NOR2 (N14265, N14257, N13536);
xor XOR2 (N14266, N14264, N11851);
and AND2 (N14267, N14265, N10260);
buf BUF1 (N14268, N14244);
nor NOR2 (N14269, N14266, N5304);
nor NOR2 (N14270, N14263, N3279);
xor XOR2 (N14271, N14251, N2243);
xor XOR2 (N14272, N14268, N3889);
nor NOR4 (N14273, N14269, N8393, N10452, N12606);
xor XOR2 (N14274, N14256, N2467);
xor XOR2 (N14275, N14272, N6954);
not NOT1 (N14276, N14271);
and AND4 (N14277, N14275, N6736, N5266, N6967);
xor XOR2 (N14278, N14276, N10454);
xor XOR2 (N14279, N14262, N11544);
or OR4 (N14280, N14252, N12622, N5923, N5282);
xor XOR2 (N14281, N14259, N5838);
nand NAND2 (N14282, N14277, N3981);
and AND4 (N14283, N14258, N8493, N12118, N9841);
xor XOR2 (N14284, N14267, N11204);
or OR3 (N14285, N14280, N2664, N5168);
not NOT1 (N14286, N14270);
or OR4 (N14287, N14273, N1176, N6368, N13269);
not NOT1 (N14288, N14287);
xor XOR2 (N14289, N14278, N13376);
nand NAND3 (N14290, N14284, N4284, N8917);
and AND4 (N14291, N14279, N3487, N6573, N1933);
nand NAND4 (N14292, N14291, N3523, N11610, N9403);
not NOT1 (N14293, N14289);
nor NOR3 (N14294, N14288, N11577, N6495);
xor XOR2 (N14295, N14282, N1857);
and AND4 (N14296, N14285, N5327, N10152, N8773);
nor NOR3 (N14297, N14293, N918, N3648);
nand NAND4 (N14298, N14286, N11328, N4459, N12102);
xor XOR2 (N14299, N14281, N7299);
buf BUF1 (N14300, N14283);
xor XOR2 (N14301, N14300, N8114);
nand NAND4 (N14302, N14292, N4190, N3374, N6364);
xor XOR2 (N14303, N14301, N7405);
buf BUF1 (N14304, N14303);
or OR2 (N14305, N14302, N12599);
nor NOR4 (N14306, N14299, N6466, N7604, N14244);
buf BUF1 (N14307, N14274);
not NOT1 (N14308, N14295);
xor XOR2 (N14309, N14296, N13258);
nor NOR3 (N14310, N14305, N2798, N3216);
nand NAND2 (N14311, N14310, N4215);
nor NOR4 (N14312, N14309, N10916, N8123, N8026);
not NOT1 (N14313, N14294);
buf BUF1 (N14314, N14307);
nor NOR4 (N14315, N14304, N504, N3846, N990);
not NOT1 (N14316, N14290);
nand NAND2 (N14317, N14298, N2576);
not NOT1 (N14318, N14311);
buf BUF1 (N14319, N14317);
not NOT1 (N14320, N14318);
buf BUF1 (N14321, N14308);
or OR4 (N14322, N14316, N11621, N5167, N9577);
nand NAND2 (N14323, N14297, N13743);
nor NOR3 (N14324, N14306, N5224, N3349);
or OR3 (N14325, N14315, N10815, N13435);
xor XOR2 (N14326, N14325, N127);
buf BUF1 (N14327, N14314);
and AND4 (N14328, N14321, N2466, N7560, N7105);
nor NOR3 (N14329, N14322, N6698, N13681);
nor NOR4 (N14330, N14327, N10563, N1952, N3508);
nand NAND4 (N14331, N14323, N9791, N9242, N9995);
nand NAND4 (N14332, N14320, N13257, N7060, N8956);
xor XOR2 (N14333, N14331, N10810);
nor NOR3 (N14334, N14312, N1320, N104);
not NOT1 (N14335, N14329);
nor NOR2 (N14336, N14319, N5609);
and AND3 (N14337, N14334, N3654, N4250);
not NOT1 (N14338, N14337);
and AND4 (N14339, N14326, N5894, N13688, N9615);
and AND2 (N14340, N14339, N3887);
nor NOR3 (N14341, N14338, N8970, N10667);
not NOT1 (N14342, N14330);
buf BUF1 (N14343, N14336);
xor XOR2 (N14344, N14333, N8846);
or OR4 (N14345, N14340, N13178, N7005, N8533);
nand NAND3 (N14346, N14344, N14170, N10500);
nor NOR2 (N14347, N14341, N3828);
buf BUF1 (N14348, N14324);
xor XOR2 (N14349, N14345, N4013);
buf BUF1 (N14350, N14346);
and AND3 (N14351, N14335, N8012, N11218);
nor NOR2 (N14352, N14348, N549);
and AND4 (N14353, N14350, N10543, N9315, N9638);
nor NOR3 (N14354, N14347, N2661, N8453);
and AND2 (N14355, N14354, N11530);
not NOT1 (N14356, N14352);
nand NAND2 (N14357, N14351, N8397);
not NOT1 (N14358, N14353);
nor NOR2 (N14359, N14356, N6408);
nor NOR3 (N14360, N14359, N123, N4143);
and AND3 (N14361, N14328, N8843, N2753);
nand NAND3 (N14362, N14358, N6102, N14126);
xor XOR2 (N14363, N14342, N2747);
nor NOR4 (N14364, N14361, N5288, N3754, N10292);
or OR2 (N14365, N14364, N10768);
nor NOR3 (N14366, N14332, N3044, N11173);
xor XOR2 (N14367, N14363, N3770);
and AND2 (N14368, N14349, N13045);
buf BUF1 (N14369, N14360);
xor XOR2 (N14370, N14367, N2308);
nor NOR3 (N14371, N14357, N4081, N1673);
nand NAND3 (N14372, N14365, N12569, N12439);
nor NOR3 (N14373, N14368, N13222, N12693);
or OR2 (N14374, N14343, N5525);
xor XOR2 (N14375, N14313, N2127);
and AND4 (N14376, N14373, N3454, N1850, N13169);
nor NOR3 (N14377, N14372, N11204, N10876);
nand NAND3 (N14378, N14374, N7164, N1633);
nor NOR3 (N14379, N14375, N7220, N902);
not NOT1 (N14380, N14370);
and AND2 (N14381, N14366, N8055);
and AND2 (N14382, N14380, N4249);
buf BUF1 (N14383, N14371);
nor NOR4 (N14384, N14381, N917, N13899, N5417);
nor NOR2 (N14385, N14355, N283);
buf BUF1 (N14386, N14377);
buf BUF1 (N14387, N14379);
or OR4 (N14388, N14382, N10298, N5748, N1321);
buf BUF1 (N14389, N14384);
xor XOR2 (N14390, N14386, N3065);
buf BUF1 (N14391, N14376);
or OR2 (N14392, N14369, N206);
buf BUF1 (N14393, N14387);
and AND3 (N14394, N14392, N8445, N1703);
and AND2 (N14395, N14393, N12059);
nor NOR2 (N14396, N14362, N6091);
not NOT1 (N14397, N14395);
not NOT1 (N14398, N14378);
nor NOR4 (N14399, N14385, N8669, N8852, N10947);
buf BUF1 (N14400, N14389);
nor NOR4 (N14401, N14390, N131, N2415, N4387);
not NOT1 (N14402, N14398);
xor XOR2 (N14403, N14396, N767);
and AND3 (N14404, N14400, N4048, N9567);
nand NAND3 (N14405, N14403, N1760, N12704);
or OR3 (N14406, N14399, N723, N13431);
buf BUF1 (N14407, N14406);
nor NOR3 (N14408, N14404, N6643, N5577);
or OR2 (N14409, N14388, N4395);
not NOT1 (N14410, N14407);
or OR3 (N14411, N14401, N6212, N1351);
xor XOR2 (N14412, N14402, N14058);
xor XOR2 (N14413, N14412, N1737);
xor XOR2 (N14414, N14413, N10946);
buf BUF1 (N14415, N14391);
not NOT1 (N14416, N14397);
buf BUF1 (N14417, N14414);
buf BUF1 (N14418, N14415);
or OR2 (N14419, N14411, N11090);
nand NAND2 (N14420, N14408, N7887);
not NOT1 (N14421, N14409);
nor NOR4 (N14422, N14405, N6944, N3959, N5974);
and AND2 (N14423, N14419, N8028);
not NOT1 (N14424, N14420);
nor NOR3 (N14425, N14421, N2021, N8489);
nand NAND2 (N14426, N14394, N11467);
nand NAND4 (N14427, N14417, N13717, N10924, N1179);
or OR2 (N14428, N14426, N4354);
buf BUF1 (N14429, N14425);
nor NOR4 (N14430, N14418, N527, N10697, N1328);
and AND2 (N14431, N14416, N10797);
xor XOR2 (N14432, N14383, N12989);
or OR4 (N14433, N14427, N5777, N8547, N7514);
xor XOR2 (N14434, N14431, N5807);
buf BUF1 (N14435, N14424);
and AND4 (N14436, N14428, N1884, N8392, N14420);
nand NAND4 (N14437, N14434, N5580, N1317, N6838);
xor XOR2 (N14438, N14432, N479);
nor NOR4 (N14439, N14437, N11195, N4310, N1967);
nand NAND3 (N14440, N14433, N9161, N11695);
nor NOR3 (N14441, N14423, N147, N9149);
not NOT1 (N14442, N14439);
buf BUF1 (N14443, N14440);
or OR4 (N14444, N14429, N915, N2762, N13625);
or OR4 (N14445, N14430, N9377, N13951, N9363);
not NOT1 (N14446, N14422);
or OR2 (N14447, N14438, N13163);
not NOT1 (N14448, N14441);
nand NAND2 (N14449, N14446, N8682);
and AND4 (N14450, N14410, N13537, N12929, N12879);
buf BUF1 (N14451, N14448);
or OR3 (N14452, N14445, N4213, N8123);
nor NOR4 (N14453, N14442, N4686, N9839, N8755);
and AND4 (N14454, N14449, N10171, N7151, N2650);
buf BUF1 (N14455, N14443);
or OR3 (N14456, N14447, N13079, N8870);
xor XOR2 (N14457, N14454, N8886);
nor NOR3 (N14458, N14457, N12008, N4528);
and AND3 (N14459, N14452, N6405, N9546);
not NOT1 (N14460, N14453);
or OR4 (N14461, N14460, N6903, N11651, N2876);
not NOT1 (N14462, N14458);
and AND4 (N14463, N14450, N368, N10026, N282);
and AND3 (N14464, N14451, N12458, N9577);
nand NAND4 (N14465, N14436, N10036, N2738, N4405);
xor XOR2 (N14466, N14444, N5301);
not NOT1 (N14467, N14466);
xor XOR2 (N14468, N14465, N89);
nor NOR2 (N14469, N14455, N9244);
nor NOR3 (N14470, N14464, N10705, N8345);
xor XOR2 (N14471, N14470, N11673);
xor XOR2 (N14472, N14456, N10272);
nand NAND2 (N14473, N14459, N4030);
not NOT1 (N14474, N14463);
not NOT1 (N14475, N14461);
not NOT1 (N14476, N14475);
nand NAND2 (N14477, N14462, N10672);
nand NAND3 (N14478, N14473, N9142, N4953);
nand NAND2 (N14479, N14467, N4078);
nand NAND2 (N14480, N14476, N7755);
nand NAND3 (N14481, N14472, N9653, N13523);
xor XOR2 (N14482, N14471, N13085);
or OR4 (N14483, N14477, N7512, N3393, N13332);
nor NOR4 (N14484, N14478, N6147, N12330, N9484);
nor NOR4 (N14485, N14483, N1949, N9114, N8569);
buf BUF1 (N14486, N14469);
nand NAND3 (N14487, N14435, N423, N4183);
nor NOR2 (N14488, N14474, N939);
or OR2 (N14489, N14486, N5654);
not NOT1 (N14490, N14484);
buf BUF1 (N14491, N14482);
nand NAND4 (N14492, N14485, N5889, N7234, N7598);
xor XOR2 (N14493, N14488, N10241);
or OR4 (N14494, N14493, N4654, N1710, N9438);
nand NAND3 (N14495, N14494, N5678, N6467);
xor XOR2 (N14496, N14490, N8059);
and AND4 (N14497, N14487, N9121, N11248, N11919);
nand NAND4 (N14498, N14480, N5850, N9939, N2447);
buf BUF1 (N14499, N14497);
or OR4 (N14500, N14492, N7761, N5122, N10788);
or OR2 (N14501, N14498, N6529);
nor NOR2 (N14502, N14495, N12785);
buf BUF1 (N14503, N14481);
xor XOR2 (N14504, N14468, N11393);
or OR3 (N14505, N14503, N124, N7046);
buf BUF1 (N14506, N14500);
and AND2 (N14507, N14479, N3147);
nor NOR2 (N14508, N14502, N12838);
or OR2 (N14509, N14496, N12476);
and AND2 (N14510, N14507, N1430);
and AND2 (N14511, N14508, N11345);
nor NOR4 (N14512, N14506, N3315, N12009, N10404);
not NOT1 (N14513, N14511);
nand NAND3 (N14514, N14510, N57, N3214);
buf BUF1 (N14515, N14491);
nor NOR2 (N14516, N14513, N15);
and AND3 (N14517, N14505, N7293, N8088);
or OR4 (N14518, N14501, N10029, N5065, N2658);
buf BUF1 (N14519, N14499);
not NOT1 (N14520, N14515);
buf BUF1 (N14521, N14519);
buf BUF1 (N14522, N14512);
xor XOR2 (N14523, N14509, N2431);
and AND4 (N14524, N14523, N7550, N267, N1654);
buf BUF1 (N14525, N14522);
and AND4 (N14526, N14504, N1360, N13462, N2317);
xor XOR2 (N14527, N14525, N6266);
xor XOR2 (N14528, N14520, N11032);
nand NAND4 (N14529, N14524, N4996, N14099, N12791);
nand NAND4 (N14530, N14521, N141, N8556, N9356);
nor NOR2 (N14531, N14518, N1613);
not NOT1 (N14532, N14516);
buf BUF1 (N14533, N14530);
xor XOR2 (N14534, N14514, N7147);
buf BUF1 (N14535, N14532);
not NOT1 (N14536, N14529);
or OR3 (N14537, N14527, N7644, N5541);
not NOT1 (N14538, N14536);
buf BUF1 (N14539, N14531);
nor NOR4 (N14540, N14517, N6394, N2161, N10340);
buf BUF1 (N14541, N14540);
buf BUF1 (N14542, N14534);
and AND3 (N14543, N14542, N6164, N5282);
nand NAND3 (N14544, N14528, N9848, N5185);
not NOT1 (N14545, N14543);
not NOT1 (N14546, N14533);
and AND3 (N14547, N14535, N1414, N12085);
xor XOR2 (N14548, N14545, N11969);
and AND3 (N14549, N14539, N3011, N10893);
not NOT1 (N14550, N14489);
nand NAND2 (N14551, N14549, N289);
or OR2 (N14552, N14537, N10545);
buf BUF1 (N14553, N14550);
not NOT1 (N14554, N14544);
and AND4 (N14555, N14538, N10659, N6847, N10181);
nor NOR3 (N14556, N14546, N11373, N8642);
xor XOR2 (N14557, N14555, N3025);
or OR3 (N14558, N14547, N13521, N8152);
buf BUF1 (N14559, N14556);
and AND3 (N14560, N14558, N10, N6682);
nand NAND4 (N14561, N14559, N6706, N7623, N4268);
xor XOR2 (N14562, N14557, N4060);
and AND3 (N14563, N14541, N2661, N13639);
buf BUF1 (N14564, N14553);
nand NAND4 (N14565, N14554, N865, N8805, N10850);
nand NAND3 (N14566, N14548, N2098, N5219);
or OR2 (N14567, N14526, N11012);
xor XOR2 (N14568, N14561, N8721);
and AND2 (N14569, N14568, N5113);
xor XOR2 (N14570, N14564, N14016);
and AND2 (N14571, N14570, N3525);
or OR4 (N14572, N14552, N1435, N4578, N13567);
and AND4 (N14573, N14566, N8496, N11677, N4599);
and AND2 (N14574, N14569, N14476);
buf BUF1 (N14575, N14573);
or OR3 (N14576, N14563, N11247, N6015);
buf BUF1 (N14577, N14572);
buf BUF1 (N14578, N14577);
and AND3 (N14579, N14575, N3447, N4550);
xor XOR2 (N14580, N14574, N13641);
nor NOR2 (N14581, N14576, N13147);
or OR2 (N14582, N14571, N6097);
not NOT1 (N14583, N14581);
or OR3 (N14584, N14579, N4179, N6338);
buf BUF1 (N14585, N14584);
buf BUF1 (N14586, N14551);
nor NOR2 (N14587, N14562, N13731);
nor NOR2 (N14588, N14565, N10323);
buf BUF1 (N14589, N14587);
nand NAND2 (N14590, N14589, N188);
and AND2 (N14591, N14567, N9252);
not NOT1 (N14592, N14560);
not NOT1 (N14593, N14588);
not NOT1 (N14594, N14578);
buf BUF1 (N14595, N14580);
nand NAND4 (N14596, N14595, N4491, N13873, N3151);
and AND4 (N14597, N14594, N13040, N8843, N6905);
not NOT1 (N14598, N14590);
buf BUF1 (N14599, N14586);
xor XOR2 (N14600, N14598, N9043);
buf BUF1 (N14601, N14583);
nor NOR3 (N14602, N14601, N4920, N7146);
buf BUF1 (N14603, N14585);
nor NOR3 (N14604, N14599, N1456, N506);
xor XOR2 (N14605, N14593, N6240);
not NOT1 (N14606, N14591);
xor XOR2 (N14607, N14604, N10540);
xor XOR2 (N14608, N14603, N5751);
buf BUF1 (N14609, N14582);
buf BUF1 (N14610, N14607);
nor NOR2 (N14611, N14602, N2668);
and AND3 (N14612, N14605, N4930, N4451);
or OR3 (N14613, N14609, N7652, N11863);
and AND2 (N14614, N14600, N5710);
nand NAND3 (N14615, N14612, N13296, N2851);
xor XOR2 (N14616, N14592, N10316);
xor XOR2 (N14617, N14611, N382);
nor NOR4 (N14618, N14596, N6451, N6731, N7190);
xor XOR2 (N14619, N14615, N14224);
xor XOR2 (N14620, N14618, N3438);
not NOT1 (N14621, N14610);
nor NOR4 (N14622, N14621, N1546, N4067, N12895);
nand NAND4 (N14623, N14622, N3802, N7366, N11897);
buf BUF1 (N14624, N14613);
not NOT1 (N14625, N14606);
and AND4 (N14626, N14619, N5768, N2182, N9326);
or OR3 (N14627, N14623, N423, N5911);
nand NAND2 (N14628, N14614, N8201);
not NOT1 (N14629, N14628);
xor XOR2 (N14630, N14597, N8875);
and AND4 (N14631, N14627, N4148, N3559, N13440);
nor NOR2 (N14632, N14616, N5330);
nand NAND2 (N14633, N14624, N14580);
buf BUF1 (N14634, N14629);
nand NAND3 (N14635, N14631, N10617, N1408);
or OR3 (N14636, N14626, N13841, N5101);
not NOT1 (N14637, N14617);
and AND4 (N14638, N14637, N160, N14081, N9444);
and AND4 (N14639, N14620, N4877, N12336, N6027);
nand NAND2 (N14640, N14636, N14492);
or OR2 (N14641, N14640, N4142);
and AND2 (N14642, N14630, N11153);
nor NOR4 (N14643, N14632, N13779, N1436, N2025);
or OR3 (N14644, N14608, N10004, N4891);
nand NAND2 (N14645, N14633, N1713);
nor NOR2 (N14646, N14638, N5548);
nor NOR4 (N14647, N14644, N592, N1997, N4365);
nor NOR2 (N14648, N14645, N9909);
not NOT1 (N14649, N14648);
xor XOR2 (N14650, N14641, N3829);
nand NAND2 (N14651, N14634, N3338);
and AND2 (N14652, N14642, N12774);
or OR3 (N14653, N14647, N13650, N11808);
nor NOR3 (N14654, N14643, N8108, N3114);
or OR2 (N14655, N14646, N529);
not NOT1 (N14656, N14635);
or OR4 (N14657, N14655, N828, N6238, N22);
nand NAND2 (N14658, N14653, N2481);
xor XOR2 (N14659, N14657, N4730);
nor NOR2 (N14660, N14650, N12927);
nand NAND3 (N14661, N14660, N4757, N10444);
xor XOR2 (N14662, N14654, N13117);
buf BUF1 (N14663, N14639);
buf BUF1 (N14664, N14662);
not NOT1 (N14665, N14658);
or OR3 (N14666, N14663, N14587, N6101);
not NOT1 (N14667, N14652);
nand NAND4 (N14668, N14625, N3413, N7672, N11287);
or OR4 (N14669, N14651, N2252, N9206, N6280);
nand NAND2 (N14670, N14661, N3703);
xor XOR2 (N14671, N14649, N1008);
xor XOR2 (N14672, N14666, N2394);
or OR2 (N14673, N14664, N6481);
nand NAND2 (N14674, N14672, N1310);
and AND4 (N14675, N14670, N3464, N9581, N6795);
nor NOR4 (N14676, N14675, N11689, N4526, N3879);
not NOT1 (N14677, N14671);
and AND3 (N14678, N14673, N1707, N5012);
nand NAND3 (N14679, N14677, N6328, N12669);
or OR4 (N14680, N14659, N5974, N10208, N1302);
or OR3 (N14681, N14667, N6635, N12863);
xor XOR2 (N14682, N14674, N9478);
nand NAND2 (N14683, N14679, N5010);
nand NAND2 (N14684, N14681, N9653);
or OR4 (N14685, N14665, N13972, N12595, N9266);
and AND2 (N14686, N14669, N3995);
buf BUF1 (N14687, N14680);
or OR2 (N14688, N14683, N14025);
buf BUF1 (N14689, N14668);
nand NAND3 (N14690, N14687, N13982, N4870);
nor NOR2 (N14691, N14678, N13183);
or OR4 (N14692, N14688, N13457, N1906, N8228);
and AND4 (N14693, N14656, N5525, N13092, N7072);
and AND2 (N14694, N14686, N4065);
nand NAND4 (N14695, N14692, N6889, N12641, N7402);
nor NOR4 (N14696, N14689, N10497, N7572, N12527);
and AND3 (N14697, N14694, N4128, N3387);
xor XOR2 (N14698, N14691, N11536);
nor NOR2 (N14699, N14693, N1751);
xor XOR2 (N14700, N14699, N10193);
nor NOR3 (N14701, N14698, N9191, N13268);
and AND3 (N14702, N14682, N4341, N12762);
buf BUF1 (N14703, N14685);
xor XOR2 (N14704, N14696, N7028);
xor XOR2 (N14705, N14701, N7204);
nand NAND4 (N14706, N14702, N8113, N13059, N2441);
or OR3 (N14707, N14690, N544, N12682);
nor NOR3 (N14708, N14697, N3386, N1412);
and AND4 (N14709, N14708, N9347, N14438, N13363);
nor NOR2 (N14710, N14705, N4387);
buf BUF1 (N14711, N14707);
nor NOR2 (N14712, N14684, N11208);
and AND2 (N14713, N14704, N9575);
xor XOR2 (N14714, N14700, N10352);
not NOT1 (N14715, N14710);
and AND2 (N14716, N14712, N2506);
and AND2 (N14717, N14711, N7000);
and AND3 (N14718, N14717, N11031, N5807);
not NOT1 (N14719, N14716);
and AND4 (N14720, N14715, N1332, N1282, N9810);
and AND3 (N14721, N14695, N9313, N11274);
nor NOR2 (N14722, N14706, N10768);
not NOT1 (N14723, N14714);
buf BUF1 (N14724, N14713);
nand NAND2 (N14725, N14720, N10908);
xor XOR2 (N14726, N14721, N7750);
nand NAND2 (N14727, N14725, N11558);
nor NOR2 (N14728, N14718, N9983);
nand NAND4 (N14729, N14709, N9153, N3397, N14086);
buf BUF1 (N14730, N14722);
not NOT1 (N14731, N14729);
not NOT1 (N14732, N14730);
or OR4 (N14733, N14724, N4133, N4780, N8623);
not NOT1 (N14734, N14723);
not NOT1 (N14735, N14676);
and AND3 (N14736, N14733, N13815, N4393);
nor NOR4 (N14737, N14726, N3081, N11143, N4376);
xor XOR2 (N14738, N14728, N13021);
or OR3 (N14739, N14737, N226, N14114);
nor NOR4 (N14740, N14738, N5735, N4759, N4795);
xor XOR2 (N14741, N14727, N5002);
not NOT1 (N14742, N14734);
buf BUF1 (N14743, N14719);
xor XOR2 (N14744, N14739, N16);
buf BUF1 (N14745, N14732);
nor NOR4 (N14746, N14736, N11685, N11578, N8345);
buf BUF1 (N14747, N14735);
xor XOR2 (N14748, N14740, N7064);
xor XOR2 (N14749, N14746, N7670);
nor NOR3 (N14750, N14748, N8559, N2662);
nand NAND4 (N14751, N14742, N12593, N7408, N4038);
not NOT1 (N14752, N14731);
nor NOR4 (N14753, N14741, N10847, N12841, N10286);
or OR2 (N14754, N14752, N13843);
buf BUF1 (N14755, N14749);
not NOT1 (N14756, N14755);
and AND3 (N14757, N14754, N8454, N4899);
nor NOR3 (N14758, N14747, N4708, N9064);
not NOT1 (N14759, N14743);
not NOT1 (N14760, N14756);
not NOT1 (N14761, N14760);
or OR3 (N14762, N14757, N3454, N3435);
and AND2 (N14763, N14762, N11364);
and AND4 (N14764, N14745, N3350, N7654, N14115);
or OR4 (N14765, N14750, N2690, N12788, N4190);
xor XOR2 (N14766, N14758, N12127);
and AND4 (N14767, N14751, N5859, N11162, N13779);
not NOT1 (N14768, N14763);
xor XOR2 (N14769, N14766, N9378);
or OR3 (N14770, N14769, N12674, N5126);
or OR2 (N14771, N14744, N8117);
buf BUF1 (N14772, N14767);
xor XOR2 (N14773, N14770, N9500);
xor XOR2 (N14774, N14753, N8596);
xor XOR2 (N14775, N14768, N351);
xor XOR2 (N14776, N14761, N12419);
and AND4 (N14777, N14771, N1601, N10648, N4003);
nor NOR2 (N14778, N14703, N14312);
nor NOR3 (N14779, N14764, N885, N9508);
and AND3 (N14780, N14776, N842, N13750);
not NOT1 (N14781, N14778);
buf BUF1 (N14782, N14765);
and AND4 (N14783, N14781, N14301, N10867, N2891);
nand NAND2 (N14784, N14772, N11817);
not NOT1 (N14785, N14759);
or OR2 (N14786, N14777, N6204);
nor NOR2 (N14787, N14785, N12539);
not NOT1 (N14788, N14773);
not NOT1 (N14789, N14775);
xor XOR2 (N14790, N14786, N1133);
not NOT1 (N14791, N14782);
or OR2 (N14792, N14783, N5619);
not NOT1 (N14793, N14792);
not NOT1 (N14794, N14784);
xor XOR2 (N14795, N14780, N6687);
not NOT1 (N14796, N14794);
xor XOR2 (N14797, N14788, N117);
not NOT1 (N14798, N14791);
nor NOR4 (N14799, N14793, N2801, N6071, N1619);
and AND3 (N14800, N14796, N3771, N2946);
and AND2 (N14801, N14799, N10927);
nor NOR2 (N14802, N14774, N12518);
nand NAND3 (N14803, N14795, N13256, N5418);
nand NAND3 (N14804, N14800, N13869, N4331);
not NOT1 (N14805, N14802);
and AND2 (N14806, N14803, N6967);
xor XOR2 (N14807, N14789, N8917);
nand NAND2 (N14808, N14801, N2283);
nor NOR3 (N14809, N14804, N7107, N13688);
or OR4 (N14810, N14805, N8054, N1464, N9118);
nand NAND2 (N14811, N14808, N6405);
not NOT1 (N14812, N14809);
nand NAND2 (N14813, N14812, N2504);
not NOT1 (N14814, N14807);
nand NAND4 (N14815, N14779, N538, N11612, N1819);
nor NOR3 (N14816, N14790, N14051, N3457);
nand NAND4 (N14817, N14806, N7934, N6603, N7701);
or OR3 (N14818, N14813, N9764, N662);
nand NAND3 (N14819, N14818, N9935, N4581);
or OR3 (N14820, N14787, N10368, N8381);
nor NOR4 (N14821, N14815, N13369, N10310, N10463);
and AND3 (N14822, N14817, N2591, N628);
not NOT1 (N14823, N14822);
not NOT1 (N14824, N14823);
xor XOR2 (N14825, N14814, N8946);
not NOT1 (N14826, N14811);
nand NAND3 (N14827, N14810, N3955, N7364);
and AND2 (N14828, N14819, N9322);
and AND3 (N14829, N14816, N266, N6277);
buf BUF1 (N14830, N14826);
xor XOR2 (N14831, N14830, N10100);
xor XOR2 (N14832, N14831, N14288);
not NOT1 (N14833, N14828);
nor NOR4 (N14834, N14797, N3748, N1655, N5102);
nor NOR4 (N14835, N14834, N1181, N135, N13971);
nand NAND4 (N14836, N14829, N11494, N11818, N988);
not NOT1 (N14837, N14827);
not NOT1 (N14838, N14798);
and AND4 (N14839, N14824, N2547, N7152, N5954);
and AND3 (N14840, N14832, N4860, N12974);
and AND2 (N14841, N14820, N3498);
nor NOR2 (N14842, N14821, N271);
not NOT1 (N14843, N14840);
xor XOR2 (N14844, N14842, N9707);
and AND2 (N14845, N14837, N6007);
nand NAND3 (N14846, N14836, N5918, N3422);
buf BUF1 (N14847, N14825);
nand NAND2 (N14848, N14839, N6725);
or OR3 (N14849, N14844, N8762, N8979);
nand NAND2 (N14850, N14841, N4340);
nor NOR2 (N14851, N14845, N3698);
xor XOR2 (N14852, N14851, N11950);
nor NOR2 (N14853, N14847, N8273);
and AND3 (N14854, N14833, N11492, N12105);
nand NAND3 (N14855, N14849, N10184, N1625);
not NOT1 (N14856, N14854);
and AND3 (N14857, N14853, N13455, N3459);
and AND4 (N14858, N14843, N10372, N13848, N14417);
nand NAND2 (N14859, N14848, N11033);
xor XOR2 (N14860, N14858, N818);
not NOT1 (N14861, N14846);
xor XOR2 (N14862, N14835, N9272);
buf BUF1 (N14863, N14857);
nand NAND3 (N14864, N14862, N5487, N2395);
not NOT1 (N14865, N14850);
nor NOR2 (N14866, N14863, N8095);
and AND3 (N14867, N14865, N1891, N9963);
nand NAND4 (N14868, N14859, N5444, N5162, N11279);
and AND3 (N14869, N14860, N5794, N371);
nand NAND2 (N14870, N14869, N13996);
nor NOR3 (N14871, N14855, N13088, N10686);
or OR4 (N14872, N14861, N10716, N5929, N3430);
xor XOR2 (N14873, N14856, N8928);
nand NAND3 (N14874, N14873, N13120, N5162);
and AND4 (N14875, N14871, N9785, N7144, N14513);
and AND2 (N14876, N14874, N7486);
nand NAND4 (N14877, N14870, N12829, N4955, N12474);
buf BUF1 (N14878, N14877);
not NOT1 (N14879, N14866);
and AND2 (N14880, N14876, N6243);
nor NOR4 (N14881, N14867, N6279, N11284, N6103);
or OR3 (N14882, N14872, N937, N9951);
or OR3 (N14883, N14875, N6914, N12998);
nor NOR2 (N14884, N14868, N1119);
nor NOR4 (N14885, N14882, N1850, N5407, N5370);
and AND2 (N14886, N14852, N8379);
not NOT1 (N14887, N14884);
or OR3 (N14888, N14878, N2608, N402);
xor XOR2 (N14889, N14879, N3935);
buf BUF1 (N14890, N14880);
nor NOR2 (N14891, N14886, N5110);
not NOT1 (N14892, N14891);
nand NAND4 (N14893, N14888, N627, N2490, N8047);
buf BUF1 (N14894, N14892);
buf BUF1 (N14895, N14893);
and AND3 (N14896, N14864, N7093, N9759);
buf BUF1 (N14897, N14890);
nor NOR4 (N14898, N14885, N12139, N11005, N4833);
nor NOR3 (N14899, N14838, N2478, N4281);
nor NOR2 (N14900, N14897, N435);
and AND2 (N14901, N14889, N8679);
and AND4 (N14902, N14894, N2091, N7766, N459);
nand NAND4 (N14903, N14898, N12166, N13017, N2696);
and AND3 (N14904, N14883, N283, N3972);
nand NAND3 (N14905, N14899, N7054, N9686);
buf BUF1 (N14906, N14896);
not NOT1 (N14907, N14901);
nand NAND2 (N14908, N14903, N3323);
not NOT1 (N14909, N14902);
nand NAND3 (N14910, N14909, N11937, N1954);
nand NAND2 (N14911, N14906, N6516);
nand NAND4 (N14912, N14900, N2630, N2824, N3249);
buf BUF1 (N14913, N14908);
and AND2 (N14914, N14904, N13200);
xor XOR2 (N14915, N14911, N5444);
nand NAND2 (N14916, N14912, N3517);
xor XOR2 (N14917, N14887, N3267);
not NOT1 (N14918, N14881);
nor NOR2 (N14919, N14914, N7786);
nand NAND3 (N14920, N14917, N12214, N111);
not NOT1 (N14921, N14905);
buf BUF1 (N14922, N14916);
nand NAND4 (N14923, N14907, N14649, N9669, N8413);
and AND4 (N14924, N14921, N14818, N7349, N13616);
xor XOR2 (N14925, N14919, N14206);
buf BUF1 (N14926, N14910);
and AND4 (N14927, N14918, N5229, N4445, N10816);
buf BUF1 (N14928, N14915);
xor XOR2 (N14929, N14926, N5107);
nand NAND4 (N14930, N14928, N10612, N10854, N10903);
and AND2 (N14931, N14925, N9741);
or OR2 (N14932, N14927, N11210);
nand NAND2 (N14933, N14932, N13331);
not NOT1 (N14934, N14931);
nor NOR3 (N14935, N14895, N185, N6395);
or OR4 (N14936, N14930, N5619, N3435, N4255);
buf BUF1 (N14937, N14922);
not NOT1 (N14938, N14923);
not NOT1 (N14939, N14937);
xor XOR2 (N14940, N14934, N693);
xor XOR2 (N14941, N14939, N13099);
nand NAND4 (N14942, N14940, N8867, N6482, N2294);
xor XOR2 (N14943, N14938, N10603);
or OR3 (N14944, N14929, N7437, N3489);
xor XOR2 (N14945, N14924, N5486);
xor XOR2 (N14946, N14944, N9335);
not NOT1 (N14947, N14933);
xor XOR2 (N14948, N14947, N9379);
xor XOR2 (N14949, N14943, N12442);
not NOT1 (N14950, N14949);
or OR4 (N14951, N14913, N1594, N12961, N11372);
xor XOR2 (N14952, N14920, N7917);
xor XOR2 (N14953, N14935, N12927);
buf BUF1 (N14954, N14948);
and AND3 (N14955, N14941, N13223, N1853);
nand NAND3 (N14956, N14936, N7632, N9729);
and AND4 (N14957, N14950, N13796, N816, N11506);
or OR4 (N14958, N14946, N5644, N8395, N3388);
or OR3 (N14959, N14957, N7797, N936);
and AND3 (N14960, N14955, N9517, N2018);
nor NOR3 (N14961, N14956, N14732, N3352);
and AND3 (N14962, N14960, N2125, N9995);
not NOT1 (N14963, N14953);
nor NOR2 (N14964, N14959, N5911);
not NOT1 (N14965, N14963);
and AND3 (N14966, N14942, N5629, N9316);
or OR2 (N14967, N14951, N13195);
buf BUF1 (N14968, N14967);
nand NAND4 (N14969, N14958, N1054, N10646, N9155);
not NOT1 (N14970, N14969);
xor XOR2 (N14971, N14968, N3998);
nand NAND2 (N14972, N14961, N1591);
buf BUF1 (N14973, N14966);
nand NAND2 (N14974, N14971, N9452);
xor XOR2 (N14975, N14954, N14265);
not NOT1 (N14976, N14975);
nor NOR4 (N14977, N14970, N7563, N12831, N10515);
not NOT1 (N14978, N14952);
xor XOR2 (N14979, N14973, N1281);
nor NOR3 (N14980, N14965, N14128, N12940);
buf BUF1 (N14981, N14962);
and AND2 (N14982, N14979, N4035);
xor XOR2 (N14983, N14981, N12803);
buf BUF1 (N14984, N14980);
not NOT1 (N14985, N14984);
or OR4 (N14986, N14985, N4997, N8664, N14438);
nor NOR2 (N14987, N14974, N6540);
nor NOR4 (N14988, N14964, N11964, N560, N5594);
or OR4 (N14989, N14986, N5097, N13939, N8699);
nor NOR4 (N14990, N14982, N6020, N2109, N1558);
not NOT1 (N14991, N14989);
buf BUF1 (N14992, N14977);
buf BUF1 (N14993, N14988);
and AND2 (N14994, N14993, N8121);
xor XOR2 (N14995, N14976, N12509);
and AND3 (N14996, N14978, N14960, N3403);
or OR2 (N14997, N14945, N6472);
buf BUF1 (N14998, N14994);
xor XOR2 (N14999, N14991, N7580);
not NOT1 (N15000, N14990);
buf BUF1 (N15001, N14987);
buf BUF1 (N15002, N15001);
nand NAND2 (N15003, N14992, N620);
nand NAND3 (N15004, N14996, N14371, N4221);
nand NAND3 (N15005, N14998, N3974, N1074);
or OR4 (N15006, N14995, N11214, N4413, N6828);
buf BUF1 (N15007, N14972);
xor XOR2 (N15008, N15004, N941);
xor XOR2 (N15009, N14997, N10018);
nor NOR3 (N15010, N14983, N2572, N5269);
and AND2 (N15011, N15007, N9485);
nand NAND2 (N15012, N15009, N5642);
and AND4 (N15013, N14999, N330, N13284, N14215);
nor NOR2 (N15014, N15012, N7341);
nand NAND2 (N15015, N15000, N3735);
and AND3 (N15016, N15013, N8147, N11305);
buf BUF1 (N15017, N15005);
xor XOR2 (N15018, N15015, N1188);
not NOT1 (N15019, N15002);
or OR2 (N15020, N15008, N8876);
and AND3 (N15021, N15018, N13576, N9599);
xor XOR2 (N15022, N15010, N9463);
nor NOR2 (N15023, N15011, N10535);
xor XOR2 (N15024, N15003, N10293);
not NOT1 (N15025, N15016);
xor XOR2 (N15026, N15022, N3787);
nand NAND3 (N15027, N15006, N6500, N2497);
and AND3 (N15028, N15014, N11831, N6630);
not NOT1 (N15029, N15019);
buf BUF1 (N15030, N15026);
and AND3 (N15031, N15023, N6472, N6996);
xor XOR2 (N15032, N15017, N12287);
and AND3 (N15033, N15024, N1156, N2444);
nor NOR2 (N15034, N15028, N10331);
xor XOR2 (N15035, N15025, N9850);
xor XOR2 (N15036, N15021, N4843);
nand NAND2 (N15037, N15031, N7158);
and AND2 (N15038, N15030, N6607);
nand NAND3 (N15039, N15033, N11470, N2757);
nand NAND3 (N15040, N15032, N9373, N10979);
buf BUF1 (N15041, N15029);
buf BUF1 (N15042, N15027);
not NOT1 (N15043, N15040);
nand NAND3 (N15044, N15039, N9636, N12662);
buf BUF1 (N15045, N15042);
or OR2 (N15046, N15044, N7625);
not NOT1 (N15047, N15038);
nand NAND3 (N15048, N15047, N12886, N12863);
or OR4 (N15049, N15043, N7506, N7131, N11985);
nand NAND4 (N15050, N15048, N5690, N4396, N305);
nor NOR4 (N15051, N15035, N4685, N10820, N5384);
nor NOR3 (N15052, N15046, N8242, N7841);
buf BUF1 (N15053, N15020);
nor NOR2 (N15054, N15049, N1436);
buf BUF1 (N15055, N15036);
buf BUF1 (N15056, N15051);
or OR4 (N15057, N15055, N5427, N9342, N3764);
buf BUF1 (N15058, N15052);
nand NAND2 (N15059, N15057, N12388);
nand NAND2 (N15060, N15037, N13506);
or OR3 (N15061, N15053, N10113, N12768);
not NOT1 (N15062, N15056);
nand NAND4 (N15063, N15054, N14123, N12008, N1287);
buf BUF1 (N15064, N15041);
or OR2 (N15065, N15034, N12762);
or OR4 (N15066, N15059, N6403, N12554, N7176);
and AND4 (N15067, N15045, N11661, N13512, N14755);
buf BUF1 (N15068, N15064);
xor XOR2 (N15069, N15065, N3670);
nand NAND4 (N15070, N15063, N2891, N7504, N13105);
nand NAND3 (N15071, N15070, N8870, N9161);
xor XOR2 (N15072, N15061, N9662);
or OR3 (N15073, N15067, N4515, N12834);
nor NOR3 (N15074, N15050, N7261, N7988);
nand NAND3 (N15075, N15072, N11583, N9921);
and AND3 (N15076, N15074, N2184, N287);
nor NOR3 (N15077, N15068, N2772, N13939);
or OR4 (N15078, N15069, N964, N13619, N9645);
and AND4 (N15079, N15066, N81, N11498, N2331);
nor NOR3 (N15080, N15077, N1845, N6470);
nand NAND4 (N15081, N15060, N10227, N7956, N11023);
buf BUF1 (N15082, N15079);
nand NAND2 (N15083, N15075, N3411);
xor XOR2 (N15084, N15082, N920);
nor NOR3 (N15085, N15078, N4306, N3884);
xor XOR2 (N15086, N15073, N1710);
buf BUF1 (N15087, N15084);
or OR4 (N15088, N15087, N14346, N366, N3583);
not NOT1 (N15089, N15088);
buf BUF1 (N15090, N15089);
not NOT1 (N15091, N15085);
not NOT1 (N15092, N15086);
xor XOR2 (N15093, N15058, N3114);
and AND2 (N15094, N15076, N14093);
nor NOR3 (N15095, N15094, N5609, N1448);
buf BUF1 (N15096, N15095);
nor NOR4 (N15097, N15090, N463, N9004, N4903);
or OR2 (N15098, N15080, N1077);
xor XOR2 (N15099, N15096, N10987);
nor NOR3 (N15100, N15099, N12221, N7191);
nor NOR3 (N15101, N15100, N6916, N5765);
or OR4 (N15102, N15101, N1002, N12557, N8845);
buf BUF1 (N15103, N15062);
or OR3 (N15104, N15081, N540, N13084);
nand NAND2 (N15105, N15092, N11892);
or OR4 (N15106, N15091, N14572, N11665, N9969);
and AND3 (N15107, N15102, N10799, N5484);
or OR4 (N15108, N15105, N3224, N10943, N4667);
nor NOR4 (N15109, N15107, N2932, N2127, N7617);
buf BUF1 (N15110, N15103);
and AND3 (N15111, N15104, N413, N9254);
nand NAND3 (N15112, N15097, N10081, N2210);
xor XOR2 (N15113, N15108, N7119);
buf BUF1 (N15114, N15093);
buf BUF1 (N15115, N15113);
buf BUF1 (N15116, N15114);
and AND3 (N15117, N15115, N3483, N6273);
nor NOR4 (N15118, N15111, N12147, N14494, N13013);
nor NOR4 (N15119, N15112, N10297, N9705, N5045);
nand NAND2 (N15120, N15118, N11552);
buf BUF1 (N15121, N15120);
nor NOR4 (N15122, N15121, N6931, N6753, N10729);
not NOT1 (N15123, N15119);
and AND4 (N15124, N15123, N2589, N1638, N1439);
buf BUF1 (N15125, N15109);
xor XOR2 (N15126, N15125, N366);
nor NOR2 (N15127, N15116, N2701);
or OR2 (N15128, N15122, N2042);
xor XOR2 (N15129, N15110, N996);
nand NAND2 (N15130, N15106, N9372);
nor NOR4 (N15131, N15098, N13197, N7101, N3754);
xor XOR2 (N15132, N15127, N11293);
or OR4 (N15133, N15128, N406, N6561, N6856);
nand NAND3 (N15134, N15071, N8224, N1597);
and AND4 (N15135, N15133, N11675, N10925, N8381);
nor NOR3 (N15136, N15126, N14696, N2322);
xor XOR2 (N15137, N15132, N4420);
nor NOR2 (N15138, N15135, N12303);
and AND3 (N15139, N15124, N10363, N7388);
not NOT1 (N15140, N15137);
nor NOR3 (N15141, N15131, N13153, N13305);
not NOT1 (N15142, N15139);
not NOT1 (N15143, N15130);
and AND4 (N15144, N15138, N11090, N14427, N10149);
nand NAND2 (N15145, N15083, N9258);
buf BUF1 (N15146, N15142);
and AND4 (N15147, N15144, N316, N6772, N10474);
nor NOR2 (N15148, N15136, N3688);
buf BUF1 (N15149, N15140);
and AND2 (N15150, N15117, N3835);
nand NAND4 (N15151, N15134, N2791, N11654, N3159);
or OR2 (N15152, N15150, N6196);
xor XOR2 (N15153, N15151, N14458);
xor XOR2 (N15154, N15149, N11819);
nor NOR2 (N15155, N15147, N4752);
or OR3 (N15156, N15145, N10196, N8882);
nor NOR4 (N15157, N15129, N3396, N3521, N9607);
nand NAND4 (N15158, N15155, N1837, N8529, N13087);
buf BUF1 (N15159, N15152);
nand NAND4 (N15160, N15141, N6814, N2534, N10050);
not NOT1 (N15161, N15148);
not NOT1 (N15162, N15154);
nand NAND2 (N15163, N15146, N2300);
buf BUF1 (N15164, N15160);
xor XOR2 (N15165, N15143, N14500);
nor NOR2 (N15166, N15153, N6416);
and AND4 (N15167, N15156, N9320, N5173, N13786);
not NOT1 (N15168, N15162);
nor NOR3 (N15169, N15164, N8419, N14532);
nor NOR4 (N15170, N15163, N10063, N1187, N3036);
buf BUF1 (N15171, N15167);
or OR4 (N15172, N15165, N5740, N10875, N10565);
buf BUF1 (N15173, N15161);
or OR3 (N15174, N15171, N8888, N8261);
buf BUF1 (N15175, N15174);
not NOT1 (N15176, N15168);
xor XOR2 (N15177, N15158, N1580);
nor NOR4 (N15178, N15173, N8143, N7424, N14713);
buf BUF1 (N15179, N15175);
nor NOR4 (N15180, N15179, N498, N11102, N887);
xor XOR2 (N15181, N15159, N7996);
nand NAND2 (N15182, N15176, N2574);
not NOT1 (N15183, N15166);
buf BUF1 (N15184, N15170);
or OR4 (N15185, N15178, N14914, N7860, N6334);
nor NOR4 (N15186, N15181, N3829, N15154, N9237);
xor XOR2 (N15187, N15169, N4355);
xor XOR2 (N15188, N15172, N9861);
buf BUF1 (N15189, N15185);
xor XOR2 (N15190, N15187, N11995);
not NOT1 (N15191, N15189);
not NOT1 (N15192, N15183);
xor XOR2 (N15193, N15182, N4465);
xor XOR2 (N15194, N15192, N1036);
buf BUF1 (N15195, N15180);
xor XOR2 (N15196, N15190, N12366);
nand NAND2 (N15197, N15193, N5210);
buf BUF1 (N15198, N15177);
nor NOR4 (N15199, N15157, N3963, N9245, N10437);
buf BUF1 (N15200, N15197);
buf BUF1 (N15201, N15186);
xor XOR2 (N15202, N15201, N4777);
xor XOR2 (N15203, N15184, N7238);
buf BUF1 (N15204, N15202);
buf BUF1 (N15205, N15188);
nand NAND2 (N15206, N15200, N11774);
and AND4 (N15207, N15198, N12012, N2826, N8254);
not NOT1 (N15208, N15205);
not NOT1 (N15209, N15204);
not NOT1 (N15210, N15209);
xor XOR2 (N15211, N15210, N2510);
xor XOR2 (N15212, N15207, N14063);
and AND2 (N15213, N15196, N5336);
nand NAND3 (N15214, N15208, N1636, N4522);
not NOT1 (N15215, N15206);
xor XOR2 (N15216, N15194, N8863);
xor XOR2 (N15217, N15203, N13971);
buf BUF1 (N15218, N15195);
not NOT1 (N15219, N15214);
or OR2 (N15220, N15199, N7933);
nand NAND4 (N15221, N15213, N8811, N1645, N1255);
not NOT1 (N15222, N15215);
not NOT1 (N15223, N15217);
xor XOR2 (N15224, N15191, N9460);
not NOT1 (N15225, N15211);
nand NAND2 (N15226, N15219, N7073);
buf BUF1 (N15227, N15222);
and AND3 (N15228, N15223, N8790, N8229);
buf BUF1 (N15229, N15227);
and AND2 (N15230, N15224, N15073);
nor NOR3 (N15231, N15212, N2139, N10670);
and AND4 (N15232, N15230, N9462, N13408, N5111);
nand NAND4 (N15233, N15229, N11809, N5592, N4898);
and AND3 (N15234, N15218, N615, N4205);
xor XOR2 (N15235, N15220, N10078);
and AND4 (N15236, N15228, N2350, N12451, N812);
or OR3 (N15237, N15226, N6606, N14716);
nand NAND2 (N15238, N15235, N8487);
xor XOR2 (N15239, N15233, N8124);
nand NAND2 (N15240, N15232, N7789);
nand NAND2 (N15241, N15240, N2500);
xor XOR2 (N15242, N15239, N8674);
buf BUF1 (N15243, N15237);
or OR3 (N15244, N15231, N14386, N6900);
and AND4 (N15245, N15243, N15000, N13117, N3672);
and AND2 (N15246, N15244, N1849);
buf BUF1 (N15247, N15246);
and AND3 (N15248, N15245, N1113, N1211);
and AND2 (N15249, N15236, N7420);
nor NOR3 (N15250, N15249, N3785, N11805);
and AND2 (N15251, N15216, N9617);
or OR3 (N15252, N15251, N12661, N11806);
buf BUF1 (N15253, N15238);
buf BUF1 (N15254, N15221);
xor XOR2 (N15255, N15253, N9551);
and AND2 (N15256, N15225, N9456);
xor XOR2 (N15257, N15252, N9204);
nand NAND4 (N15258, N15242, N7242, N8782, N1575);
not NOT1 (N15259, N15254);
and AND3 (N15260, N15255, N14073, N4071);
or OR3 (N15261, N15250, N4589, N264);
xor XOR2 (N15262, N15234, N10936);
buf BUF1 (N15263, N15256);
xor XOR2 (N15264, N15241, N3472);
nor NOR2 (N15265, N15258, N2816);
buf BUF1 (N15266, N15259);
not NOT1 (N15267, N15263);
not NOT1 (N15268, N15262);
or OR4 (N15269, N15257, N10213, N1815, N11162);
not NOT1 (N15270, N15265);
nand NAND4 (N15271, N15260, N5908, N8873, N10239);
xor XOR2 (N15272, N15264, N3323);
and AND2 (N15273, N15269, N4440);
not NOT1 (N15274, N15267);
nor NOR4 (N15275, N15266, N11791, N1710, N8822);
or OR3 (N15276, N15268, N3865, N9897);
xor XOR2 (N15277, N15248, N5875);
nor NOR2 (N15278, N15271, N11701);
and AND2 (N15279, N15247, N9811);
nor NOR2 (N15280, N15270, N11567);
and AND3 (N15281, N15278, N8624, N14235);
xor XOR2 (N15282, N15281, N4997);
buf BUF1 (N15283, N15272);
nand NAND2 (N15284, N15261, N9933);
not NOT1 (N15285, N15283);
buf BUF1 (N15286, N15273);
nand NAND3 (N15287, N15276, N15044, N7207);
nand NAND2 (N15288, N15277, N15150);
and AND4 (N15289, N15280, N14221, N903, N12795);
not NOT1 (N15290, N15284);
nor NOR2 (N15291, N15286, N608);
nor NOR3 (N15292, N15282, N9604, N12398);
not NOT1 (N15293, N15285);
or OR4 (N15294, N15289, N8838, N12362, N13529);
xor XOR2 (N15295, N15291, N14939);
not NOT1 (N15296, N15292);
nor NOR3 (N15297, N15288, N12399, N2045);
and AND3 (N15298, N15287, N8635, N8429);
nor NOR4 (N15299, N15295, N7881, N13898, N12838);
nor NOR3 (N15300, N15299, N10780, N4167);
or OR3 (N15301, N15294, N728, N9581);
xor XOR2 (N15302, N15296, N4459);
nand NAND3 (N15303, N15275, N12761, N10280);
not NOT1 (N15304, N15274);
buf BUF1 (N15305, N15302);
or OR3 (N15306, N15293, N12884, N10314);
nand NAND2 (N15307, N15305, N9437);
nor NOR3 (N15308, N15298, N1787, N6596);
nand NAND2 (N15309, N15297, N8794);
nand NAND3 (N15310, N15290, N3792, N666);
and AND2 (N15311, N15310, N9334);
buf BUF1 (N15312, N15300);
or OR3 (N15313, N15279, N2651, N4922);
xor XOR2 (N15314, N15311, N9213);
nor NOR3 (N15315, N15301, N10753, N5566);
or OR2 (N15316, N15304, N8569);
not NOT1 (N15317, N15306);
nor NOR4 (N15318, N15309, N1272, N14650, N13581);
xor XOR2 (N15319, N15303, N4671);
buf BUF1 (N15320, N15312);
buf BUF1 (N15321, N15307);
buf BUF1 (N15322, N15314);
and AND2 (N15323, N15320, N11770);
nor NOR4 (N15324, N15316, N1747, N2603, N2797);
nor NOR4 (N15325, N15322, N1996, N9806, N4727);
or OR2 (N15326, N15319, N11239);
nand NAND3 (N15327, N15321, N5069, N15290);
not NOT1 (N15328, N15327);
nand NAND4 (N15329, N15326, N6348, N9440, N11576);
nand NAND3 (N15330, N15323, N7811, N10218);
and AND3 (N15331, N15330, N14360, N14467);
and AND4 (N15332, N15313, N13279, N3273, N10167);
buf BUF1 (N15333, N15308);
buf BUF1 (N15334, N15331);
xor XOR2 (N15335, N15325, N14968);
or OR3 (N15336, N15334, N1397, N4665);
and AND3 (N15337, N15336, N10127, N8581);
nand NAND4 (N15338, N15328, N10067, N10198, N10203);
or OR3 (N15339, N15317, N1634, N10474);
nand NAND3 (N15340, N15335, N14296, N8293);
xor XOR2 (N15341, N15337, N4584);
and AND2 (N15342, N15333, N3276);
not NOT1 (N15343, N15341);
nor NOR2 (N15344, N15315, N4367);
not NOT1 (N15345, N15339);
nand NAND2 (N15346, N15343, N9918);
buf BUF1 (N15347, N15329);
nor NOR4 (N15348, N15346, N13571, N14650, N5733);
or OR4 (N15349, N15347, N5476, N10501, N13825);
or OR4 (N15350, N15318, N3992, N13049, N5559);
not NOT1 (N15351, N15345);
or OR2 (N15352, N15342, N11692);
xor XOR2 (N15353, N15332, N10408);
buf BUF1 (N15354, N15353);
not NOT1 (N15355, N15344);
buf BUF1 (N15356, N15352);
nor NOR3 (N15357, N15349, N3046, N8179);
and AND4 (N15358, N15324, N14120, N13484, N15213);
nand NAND4 (N15359, N15350, N13945, N14092, N6961);
nand NAND2 (N15360, N15357, N12246);
xor XOR2 (N15361, N15351, N4959);
and AND4 (N15362, N15360, N4982, N431, N12234);
nor NOR4 (N15363, N15356, N11831, N7791, N10493);
nand NAND4 (N15364, N15358, N7569, N9460, N10561);
or OR2 (N15365, N15359, N8283);
nand NAND3 (N15366, N15363, N5016, N3899);
nand NAND3 (N15367, N15338, N9379, N2134);
buf BUF1 (N15368, N15355);
nor NOR4 (N15369, N15362, N3095, N11411, N5712);
nand NAND3 (N15370, N15367, N12150, N10666);
nand NAND3 (N15371, N15368, N352, N1284);
buf BUF1 (N15372, N15340);
nor NOR2 (N15373, N15348, N4363);
not NOT1 (N15374, N15369);
buf BUF1 (N15375, N15374);
buf BUF1 (N15376, N15371);
nor NOR4 (N15377, N15373, N3597, N3798, N1710);
nor NOR4 (N15378, N15377, N8220, N2574, N15358);
and AND3 (N15379, N15372, N2517, N2882);
or OR4 (N15380, N15378, N1159, N14999, N109);
or OR4 (N15381, N15366, N2235, N2983, N13944);
and AND2 (N15382, N15380, N8736);
buf BUF1 (N15383, N15379);
xor XOR2 (N15384, N15383, N15343);
or OR3 (N15385, N15365, N8173, N1833);
or OR3 (N15386, N15376, N7751, N4140);
or OR4 (N15387, N15364, N10817, N5320, N11952);
not NOT1 (N15388, N15381);
and AND2 (N15389, N15375, N10532);
xor XOR2 (N15390, N15388, N10695);
or OR2 (N15391, N15387, N14342);
and AND4 (N15392, N15389, N13476, N13895, N1609);
nor NOR4 (N15393, N15392, N10173, N8868, N14444);
or OR4 (N15394, N15370, N1970, N5337, N10895);
buf BUF1 (N15395, N15394);
xor XOR2 (N15396, N15385, N8872);
nor NOR4 (N15397, N15396, N258, N14860, N808);
xor XOR2 (N15398, N15390, N7316);
or OR2 (N15399, N15393, N15320);
or OR2 (N15400, N15361, N3307);
nor NOR3 (N15401, N15395, N3695, N11891);
nor NOR2 (N15402, N15397, N8276);
and AND3 (N15403, N15399, N2914, N6117);
xor XOR2 (N15404, N15386, N7860);
and AND2 (N15405, N15403, N1584);
xor XOR2 (N15406, N15354, N2827);
not NOT1 (N15407, N15404);
nor NOR2 (N15408, N15400, N8468);
buf BUF1 (N15409, N15405);
not NOT1 (N15410, N15406);
xor XOR2 (N15411, N15408, N4170);
nand NAND4 (N15412, N15407, N5310, N10482, N88);
or OR2 (N15413, N15411, N8127);
nand NAND3 (N15414, N15410, N10710, N9186);
xor XOR2 (N15415, N15412, N13550);
or OR2 (N15416, N15415, N10127);
nand NAND3 (N15417, N15414, N172, N4786);
xor XOR2 (N15418, N15401, N6401);
nand NAND2 (N15419, N15413, N3039);
buf BUF1 (N15420, N15419);
nor NOR4 (N15421, N15391, N13910, N8682, N4524);
not NOT1 (N15422, N15418);
not NOT1 (N15423, N15398);
and AND4 (N15424, N15417, N10417, N2595, N191);
not NOT1 (N15425, N15382);
nand NAND3 (N15426, N15423, N14877, N10143);
not NOT1 (N15427, N15424);
nand NAND2 (N15428, N15409, N8199);
nor NOR4 (N15429, N15416, N10808, N4824, N3811);
nor NOR2 (N15430, N15420, N14267);
buf BUF1 (N15431, N15428);
and AND3 (N15432, N15427, N14069, N11421);
not NOT1 (N15433, N15429);
xor XOR2 (N15434, N15421, N14354);
xor XOR2 (N15435, N15426, N4988);
xor XOR2 (N15436, N15425, N14400);
buf BUF1 (N15437, N15402);
buf BUF1 (N15438, N15430);
buf BUF1 (N15439, N15432);
nand NAND4 (N15440, N15439, N8098, N5608, N11169);
nand NAND3 (N15441, N15434, N12365, N5588);
nor NOR2 (N15442, N15441, N5341);
nand NAND4 (N15443, N15442, N6460, N2314, N1222);
xor XOR2 (N15444, N15431, N6690);
xor XOR2 (N15445, N15435, N9963);
nor NOR3 (N15446, N15443, N12481, N15204);
buf BUF1 (N15447, N15433);
or OR2 (N15448, N15446, N14429);
nor NOR4 (N15449, N15444, N9345, N2326, N11111);
not NOT1 (N15450, N15384);
nand NAND2 (N15451, N15422, N1090);
buf BUF1 (N15452, N15449);
nor NOR3 (N15453, N15440, N2267, N7748);
xor XOR2 (N15454, N15452, N3604);
nand NAND2 (N15455, N15454, N9219);
not NOT1 (N15456, N15438);
xor XOR2 (N15457, N15448, N8422);
nor NOR2 (N15458, N15457, N15120);
nor NOR2 (N15459, N15453, N5256);
nand NAND2 (N15460, N15447, N14167);
and AND2 (N15461, N15458, N10216);
not NOT1 (N15462, N15445);
nand NAND3 (N15463, N15455, N10272, N9002);
not NOT1 (N15464, N15451);
or OR2 (N15465, N15460, N2767);
xor XOR2 (N15466, N15450, N13835);
nor NOR3 (N15467, N15463, N14393, N1770);
not NOT1 (N15468, N15467);
not NOT1 (N15469, N15436);
xor XOR2 (N15470, N15461, N5676);
and AND2 (N15471, N15464, N4705);
nand NAND4 (N15472, N15462, N10116, N13143, N12262);
not NOT1 (N15473, N15471);
nand NAND4 (N15474, N15466, N8041, N13451, N14198);
nand NAND3 (N15475, N15437, N879, N15055);
nand NAND2 (N15476, N15456, N14299);
nand NAND2 (N15477, N15472, N6046);
nand NAND4 (N15478, N15476, N2587, N1425, N12088);
and AND4 (N15479, N15469, N5861, N13836, N11438);
and AND4 (N15480, N15477, N3086, N11441, N5739);
nor NOR4 (N15481, N15478, N3642, N15474, N7198);
nor NOR3 (N15482, N9436, N2258, N3358);
nand NAND4 (N15483, N15468, N9319, N4680, N1156);
buf BUF1 (N15484, N15482);
xor XOR2 (N15485, N15480, N4394);
nor NOR3 (N15486, N15459, N10369, N14643);
not NOT1 (N15487, N15479);
and AND4 (N15488, N15485, N7629, N13678, N8193);
buf BUF1 (N15489, N15470);
nor NOR2 (N15490, N15486, N3359);
xor XOR2 (N15491, N15481, N7872);
buf BUF1 (N15492, N15491);
nand NAND2 (N15493, N15489, N12797);
nor NOR4 (N15494, N15465, N741, N14312, N9828);
or OR2 (N15495, N15490, N5903);
nor NOR2 (N15496, N15493, N674);
not NOT1 (N15497, N15484);
or OR4 (N15498, N15494, N11334, N9759, N14449);
buf BUF1 (N15499, N15475);
xor XOR2 (N15500, N15498, N14892);
buf BUF1 (N15501, N15488);
not NOT1 (N15502, N15495);
not NOT1 (N15503, N15487);
nor NOR2 (N15504, N15503, N12538);
nand NAND3 (N15505, N15473, N13671, N4570);
nand NAND2 (N15506, N15496, N5072);
xor XOR2 (N15507, N15499, N9107);
and AND3 (N15508, N15504, N908, N679);
not NOT1 (N15509, N15497);
buf BUF1 (N15510, N15505);
not NOT1 (N15511, N15500);
not NOT1 (N15512, N15510);
not NOT1 (N15513, N15501);
nand NAND4 (N15514, N15492, N7313, N9802, N3742);
or OR4 (N15515, N15507, N10253, N2269, N5763);
xor XOR2 (N15516, N15508, N6765);
buf BUF1 (N15517, N15502);
and AND4 (N15518, N15512, N8916, N11801, N7592);
not NOT1 (N15519, N15511);
and AND4 (N15520, N15506, N9205, N9659, N3901);
xor XOR2 (N15521, N15516, N9460);
not NOT1 (N15522, N15515);
and AND4 (N15523, N15514, N5736, N1898, N13947);
or OR3 (N15524, N15523, N8949, N13757);
not NOT1 (N15525, N15522);
buf BUF1 (N15526, N15483);
not NOT1 (N15527, N15524);
buf BUF1 (N15528, N15513);
nor NOR3 (N15529, N15526, N13732, N855);
buf BUF1 (N15530, N15525);
or OR4 (N15531, N15530, N8636, N1880, N15302);
xor XOR2 (N15532, N15531, N7532);
nor NOR2 (N15533, N15528, N9978);
not NOT1 (N15534, N15527);
buf BUF1 (N15535, N15518);
and AND3 (N15536, N15529, N4690, N14788);
and AND2 (N15537, N15509, N7681);
buf BUF1 (N15538, N15520);
or OR4 (N15539, N15521, N13302, N4165, N14584);
and AND2 (N15540, N15534, N6774);
xor XOR2 (N15541, N15535, N8572);
nor NOR4 (N15542, N15540, N2538, N9587, N1755);
nor NOR4 (N15543, N15542, N3965, N4471, N12155);
nand NAND3 (N15544, N15539, N14658, N5533);
nand NAND2 (N15545, N15532, N9182);
and AND3 (N15546, N15519, N12004, N298);
nand NAND3 (N15547, N15544, N5582, N7842);
nand NAND3 (N15548, N15546, N14, N3161);
nor NOR4 (N15549, N15517, N4286, N3690, N13421);
xor XOR2 (N15550, N15537, N7775);
nor NOR4 (N15551, N15543, N9496, N7771, N9560);
nand NAND4 (N15552, N15541, N2967, N522, N9296);
not NOT1 (N15553, N15547);
nor NOR3 (N15554, N15538, N15091, N12420);
nand NAND3 (N15555, N15533, N2283, N9209);
buf BUF1 (N15556, N15553);
not NOT1 (N15557, N15550);
and AND4 (N15558, N15556, N14638, N447, N9193);
nand NAND3 (N15559, N15548, N12297, N14528);
or OR4 (N15560, N15545, N14609, N15206, N10471);
buf BUF1 (N15561, N15536);
buf BUF1 (N15562, N15561);
buf BUF1 (N15563, N15562);
or OR3 (N15564, N15551, N14434, N14249);
buf BUF1 (N15565, N15559);
xor XOR2 (N15566, N15552, N408);
and AND3 (N15567, N15549, N3422, N6390);
or OR3 (N15568, N15566, N14289, N2795);
or OR4 (N15569, N15554, N3549, N4663, N11835);
nand NAND3 (N15570, N15563, N10131, N89);
nor NOR3 (N15571, N15567, N5937, N3264);
not NOT1 (N15572, N15571);
nor NOR2 (N15573, N15570, N5737);
xor XOR2 (N15574, N15564, N2860);
nor NOR3 (N15575, N15574, N4608, N9237);
or OR4 (N15576, N15558, N2276, N4910, N5102);
xor XOR2 (N15577, N15576, N10987);
nor NOR3 (N15578, N15572, N2265, N13593);
or OR3 (N15579, N15573, N6975, N6317);
and AND4 (N15580, N15555, N9904, N8736, N13490);
nor NOR2 (N15581, N15569, N11631);
not NOT1 (N15582, N15565);
and AND3 (N15583, N15568, N2293, N11648);
nand NAND3 (N15584, N15560, N1198, N4266);
xor XOR2 (N15585, N15577, N3280);
and AND4 (N15586, N15584, N4273, N12992, N5909);
not NOT1 (N15587, N15578);
or OR2 (N15588, N15582, N2701);
buf BUF1 (N15589, N15579);
xor XOR2 (N15590, N15588, N11569);
or OR3 (N15591, N15575, N1565, N4588);
and AND3 (N15592, N15581, N13967, N10077);
nand NAND2 (N15593, N15557, N9689);
not NOT1 (N15594, N15591);
and AND2 (N15595, N15594, N6354);
or OR3 (N15596, N15585, N6120, N10103);
and AND3 (N15597, N15590, N1461, N9570);
buf BUF1 (N15598, N15583);
xor XOR2 (N15599, N15593, N14875);
buf BUF1 (N15600, N15586);
buf BUF1 (N15601, N15595);
or OR2 (N15602, N15589, N10211);
buf BUF1 (N15603, N15596);
or OR4 (N15604, N15602, N7554, N3892, N404);
buf BUF1 (N15605, N15580);
nand NAND3 (N15606, N15600, N9989, N3716);
and AND3 (N15607, N15603, N4667, N10544);
not NOT1 (N15608, N15598);
or OR4 (N15609, N15601, N6895, N6485, N9616);
xor XOR2 (N15610, N15592, N2164);
xor XOR2 (N15611, N15597, N1029);
nand NAND2 (N15612, N15609, N9809);
and AND3 (N15613, N15607, N4783, N677);
xor XOR2 (N15614, N15599, N2704);
not NOT1 (N15615, N15610);
and AND4 (N15616, N15612, N3451, N1593, N10448);
or OR3 (N15617, N15614, N5560, N9408);
nand NAND3 (N15618, N15604, N333, N1822);
nor NOR4 (N15619, N15613, N9754, N3673, N9634);
nand NAND4 (N15620, N15606, N11626, N7179, N11468);
nor NOR3 (N15621, N15608, N8284, N14802);
nand NAND2 (N15622, N15621, N2629);
and AND3 (N15623, N15617, N5093, N6304);
xor XOR2 (N15624, N15618, N13392);
not NOT1 (N15625, N15605);
xor XOR2 (N15626, N15620, N2775);
not NOT1 (N15627, N15623);
not NOT1 (N15628, N15615);
and AND3 (N15629, N15626, N12885, N6066);
and AND3 (N15630, N15622, N465, N12903);
not NOT1 (N15631, N15587);
not NOT1 (N15632, N15619);
nand NAND4 (N15633, N15624, N4553, N9856, N11989);
not NOT1 (N15634, N15616);
or OR3 (N15635, N15631, N8043, N5369);
not NOT1 (N15636, N15629);
nor NOR3 (N15637, N15632, N152, N325);
and AND4 (N15638, N15636, N11957, N2889, N11863);
not NOT1 (N15639, N15635);
and AND3 (N15640, N15630, N6634, N393);
buf BUF1 (N15641, N15637);
not NOT1 (N15642, N15625);
and AND2 (N15643, N15641, N10303);
nand NAND4 (N15644, N15611, N10189, N6156, N494);
nand NAND3 (N15645, N15627, N7426, N9943);
buf BUF1 (N15646, N15640);
nand NAND4 (N15647, N15628, N14492, N9734, N11220);
nand NAND2 (N15648, N15633, N3789);
not NOT1 (N15649, N15642);
xor XOR2 (N15650, N15643, N11863);
xor XOR2 (N15651, N15645, N941);
or OR3 (N15652, N15649, N10886, N7443);
and AND3 (N15653, N15646, N4983, N11815);
and AND3 (N15654, N15648, N11026, N15459);
nand NAND4 (N15655, N15638, N14771, N5918, N12885);
not NOT1 (N15656, N15647);
nand NAND2 (N15657, N15651, N14848);
xor XOR2 (N15658, N15634, N8462);
not NOT1 (N15659, N15656);
nor NOR4 (N15660, N15639, N7766, N8621, N3484);
not NOT1 (N15661, N15658);
or OR3 (N15662, N15659, N392, N4133);
and AND4 (N15663, N15644, N12026, N5132, N7498);
xor XOR2 (N15664, N15654, N3404);
xor XOR2 (N15665, N15652, N896);
xor XOR2 (N15666, N15661, N11858);
nand NAND2 (N15667, N15660, N9198);
nor NOR3 (N15668, N15666, N6146, N12698);
xor XOR2 (N15669, N15665, N228);
xor XOR2 (N15670, N15664, N11178);
or OR2 (N15671, N15663, N14726);
nor NOR3 (N15672, N15655, N1480, N4240);
buf BUF1 (N15673, N15657);
or OR4 (N15674, N15662, N1568, N14215, N11063);
and AND2 (N15675, N15672, N2800);
buf BUF1 (N15676, N15650);
xor XOR2 (N15677, N15669, N1588);
nand NAND3 (N15678, N15670, N1566, N15180);
nand NAND3 (N15679, N15675, N6769, N4695);
and AND3 (N15680, N15679, N11494, N7320);
or OR2 (N15681, N15667, N8326);
and AND3 (N15682, N15680, N4139, N13939);
not NOT1 (N15683, N15671);
or OR4 (N15684, N15681, N1370, N6497, N6765);
not NOT1 (N15685, N15673);
and AND2 (N15686, N15682, N7439);
not NOT1 (N15687, N15683);
buf BUF1 (N15688, N15677);
nor NOR4 (N15689, N15684, N14403, N4174, N11362);
and AND4 (N15690, N15668, N5081, N13533, N7188);
buf BUF1 (N15691, N15687);
buf BUF1 (N15692, N15676);
not NOT1 (N15693, N15688);
xor XOR2 (N15694, N15693, N5831);
and AND3 (N15695, N15690, N5066, N14550);
not NOT1 (N15696, N15686);
nor NOR3 (N15697, N15689, N7154, N15054);
not NOT1 (N15698, N15696);
not NOT1 (N15699, N15698);
or OR3 (N15700, N15674, N3510, N14292);
xor XOR2 (N15701, N15691, N14110);
or OR3 (N15702, N15699, N12092, N14984);
or OR3 (N15703, N15694, N14170, N3947);
or OR2 (N15704, N15697, N2572);
xor XOR2 (N15705, N15692, N10494);
or OR4 (N15706, N15700, N3389, N105, N2733);
buf BUF1 (N15707, N15678);
or OR3 (N15708, N15695, N10235, N3999);
or OR4 (N15709, N15702, N12340, N2201, N3946);
nand NAND2 (N15710, N15706, N4517);
and AND4 (N15711, N15701, N4370, N2963, N4212);
not NOT1 (N15712, N15709);
and AND4 (N15713, N15653, N3981, N1537, N11969);
nand NAND3 (N15714, N15705, N8780, N11608);
buf BUF1 (N15715, N15703);
or OR4 (N15716, N15685, N8603, N12541, N2596);
nor NOR3 (N15717, N15713, N6238, N7529);
or OR2 (N15718, N15717, N1535);
not NOT1 (N15719, N15718);
and AND4 (N15720, N15719, N12966, N9140, N4252);
not NOT1 (N15721, N15710);
xor XOR2 (N15722, N15712, N6747);
nand NAND3 (N15723, N15714, N2784, N4147);
nand NAND2 (N15724, N15721, N11451);
or OR4 (N15725, N15704, N6146, N13106, N11256);
or OR2 (N15726, N15720, N9192);
not NOT1 (N15727, N15722);
buf BUF1 (N15728, N15715);
and AND2 (N15729, N15724, N2654);
and AND3 (N15730, N15711, N5791, N5700);
nand NAND4 (N15731, N15725, N14711, N2361, N7275);
not NOT1 (N15732, N15729);
nand NAND2 (N15733, N15708, N4296);
or OR2 (N15734, N15723, N14053);
or OR4 (N15735, N15726, N13442, N1432, N12089);
not NOT1 (N15736, N15732);
xor XOR2 (N15737, N15728, N7178);
or OR3 (N15738, N15716, N15207, N12780);
or OR2 (N15739, N15737, N3533);
or OR2 (N15740, N15733, N1367);
not NOT1 (N15741, N15736);
nor NOR4 (N15742, N15740, N1959, N3039, N11714);
nand NAND4 (N15743, N15730, N7148, N14230, N10004);
buf BUF1 (N15744, N15741);
and AND2 (N15745, N15742, N5130);
and AND4 (N15746, N15727, N586, N45, N11233);
not NOT1 (N15747, N15743);
or OR3 (N15748, N15734, N1188, N10301);
and AND2 (N15749, N15747, N1687);
nand NAND4 (N15750, N15744, N5876, N408, N5598);
xor XOR2 (N15751, N15739, N13853);
nand NAND4 (N15752, N15707, N1592, N1035, N11618);
or OR4 (N15753, N15745, N3539, N2113, N1938);
or OR4 (N15754, N15731, N5195, N6421, N6471);
nand NAND3 (N15755, N15749, N7536, N11088);
nand NAND3 (N15756, N15755, N7061, N761);
nand NAND2 (N15757, N15735, N7668);
nor NOR4 (N15758, N15746, N12381, N15091, N8760);
and AND3 (N15759, N15752, N15388, N104);
xor XOR2 (N15760, N15757, N14253);
nor NOR4 (N15761, N15756, N5684, N9132, N4536);
nor NOR4 (N15762, N15738, N835, N2114, N1203);
or OR4 (N15763, N15760, N8724, N2496, N1378);
nand NAND4 (N15764, N15750, N8913, N11861, N6397);
nor NOR3 (N15765, N15761, N11329, N9776);
or OR4 (N15766, N15751, N12668, N10000, N13957);
nand NAND2 (N15767, N15759, N2293);
or OR2 (N15768, N15762, N9090);
nand NAND3 (N15769, N15758, N7498, N6295);
xor XOR2 (N15770, N15764, N12104);
nand NAND3 (N15771, N15753, N14973, N12069);
nand NAND2 (N15772, N15768, N5016);
buf BUF1 (N15773, N15754);
nor NOR2 (N15774, N15772, N1926);
not NOT1 (N15775, N15767);
xor XOR2 (N15776, N15773, N3695);
buf BUF1 (N15777, N15774);
buf BUF1 (N15778, N15748);
and AND2 (N15779, N15776, N14181);
nand NAND4 (N15780, N15765, N13294, N774, N1883);
or OR4 (N15781, N15763, N5228, N12695, N7657);
not NOT1 (N15782, N15779);
not NOT1 (N15783, N15782);
xor XOR2 (N15784, N15783, N11644);
nor NOR2 (N15785, N15766, N7359);
nand NAND3 (N15786, N15769, N10614, N6012);
xor XOR2 (N15787, N15778, N5250);
xor XOR2 (N15788, N15780, N8391);
buf BUF1 (N15789, N15770);
not NOT1 (N15790, N15786);
nand NAND3 (N15791, N15771, N2192, N11507);
nor NOR2 (N15792, N15784, N8619);
buf BUF1 (N15793, N15791);
or OR3 (N15794, N15777, N14696, N2430);
not NOT1 (N15795, N15788);
or OR2 (N15796, N15787, N5162);
nand NAND3 (N15797, N15785, N14086, N1532);
buf BUF1 (N15798, N15796);
and AND3 (N15799, N15794, N13902, N14030);
nand NAND4 (N15800, N15775, N10357, N6833, N7896);
or OR3 (N15801, N15795, N14347, N14947);
buf BUF1 (N15802, N15798);
and AND2 (N15803, N15797, N1047);
xor XOR2 (N15804, N15792, N4572);
or OR3 (N15805, N15793, N7370, N737);
nand NAND3 (N15806, N15801, N4969, N12441);
buf BUF1 (N15807, N15806);
and AND2 (N15808, N15803, N3925);
or OR4 (N15809, N15790, N9526, N11574, N7910);
xor XOR2 (N15810, N15781, N12822);
or OR4 (N15811, N15809, N6005, N8383, N12531);
xor XOR2 (N15812, N15804, N125);
xor XOR2 (N15813, N15789, N9607);
or OR4 (N15814, N15805, N11365, N348, N5757);
not NOT1 (N15815, N15808);
not NOT1 (N15816, N15810);
nor NOR3 (N15817, N15799, N14940, N3043);
or OR2 (N15818, N15802, N6240);
nor NOR3 (N15819, N15816, N9833, N6840);
nor NOR2 (N15820, N15811, N6310);
buf BUF1 (N15821, N15813);
nor NOR2 (N15822, N15818, N13717);
buf BUF1 (N15823, N15821);
nor NOR3 (N15824, N15812, N14966, N14739);
nor NOR4 (N15825, N15815, N5793, N5523, N8957);
not NOT1 (N15826, N15824);
xor XOR2 (N15827, N15822, N13054);
not NOT1 (N15828, N15826);
not NOT1 (N15829, N15825);
buf BUF1 (N15830, N15823);
nor NOR3 (N15831, N15829, N8487, N5283);
nor NOR4 (N15832, N15827, N3123, N13988, N5757);
and AND3 (N15833, N15832, N7199, N11440);
buf BUF1 (N15834, N15807);
and AND4 (N15835, N15833, N6753, N2886, N871);
and AND4 (N15836, N15819, N11236, N874, N7118);
nand NAND2 (N15837, N15814, N8002);
nor NOR3 (N15838, N15831, N15339, N5053);
and AND3 (N15839, N15830, N3816, N15445);
and AND2 (N15840, N15834, N2019);
nor NOR3 (N15841, N15836, N6590, N13692);
not NOT1 (N15842, N15817);
and AND2 (N15843, N15842, N6817);
nand NAND3 (N15844, N15840, N11099, N438);
and AND2 (N15845, N15844, N6468);
xor XOR2 (N15846, N15800, N4509);
buf BUF1 (N15847, N15837);
buf BUF1 (N15848, N15841);
xor XOR2 (N15849, N15838, N2508);
and AND2 (N15850, N15843, N246);
not NOT1 (N15851, N15849);
buf BUF1 (N15852, N15846);
and AND2 (N15853, N15835, N1938);
and AND4 (N15854, N15828, N13217, N5574, N880);
buf BUF1 (N15855, N15845);
nor NOR3 (N15856, N15853, N112, N7569);
nand NAND4 (N15857, N15855, N157, N2004, N4917);
not NOT1 (N15858, N15839);
not NOT1 (N15859, N15856);
or OR2 (N15860, N15820, N2234);
buf BUF1 (N15861, N15858);
or OR3 (N15862, N15847, N2453, N8519);
buf BUF1 (N15863, N15860);
nor NOR2 (N15864, N15862, N6798);
not NOT1 (N15865, N15848);
not NOT1 (N15866, N15854);
nor NOR4 (N15867, N15865, N2007, N13080, N4594);
and AND3 (N15868, N15852, N4786, N8838);
or OR2 (N15869, N15851, N9087);
buf BUF1 (N15870, N15861);
xor XOR2 (N15871, N15869, N3541);
nor NOR3 (N15872, N15863, N14045, N7103);
and AND3 (N15873, N15871, N9681, N2695);
not NOT1 (N15874, N15867);
not NOT1 (N15875, N15872);
and AND2 (N15876, N15864, N7233);
or OR2 (N15877, N15866, N9003);
not NOT1 (N15878, N15874);
xor XOR2 (N15879, N15857, N6116);
buf BUF1 (N15880, N15878);
xor XOR2 (N15881, N15870, N13796);
xor XOR2 (N15882, N15877, N4800);
nand NAND2 (N15883, N15881, N2119);
xor XOR2 (N15884, N15859, N12926);
not NOT1 (N15885, N15850);
buf BUF1 (N15886, N15879);
nor NOR3 (N15887, N15875, N15830, N12745);
nor NOR4 (N15888, N15884, N15068, N4616, N15859);
or OR2 (N15889, N15882, N622);
and AND3 (N15890, N15873, N12237, N728);
buf BUF1 (N15891, N15868);
not NOT1 (N15892, N15876);
nor NOR4 (N15893, N15889, N8932, N5134, N5948);
not NOT1 (N15894, N15880);
not NOT1 (N15895, N15887);
and AND4 (N15896, N15893, N6317, N7608, N14923);
nor NOR2 (N15897, N15886, N1216);
nor NOR3 (N15898, N15890, N9344, N3120);
and AND3 (N15899, N15891, N5507, N612);
buf BUF1 (N15900, N15899);
xor XOR2 (N15901, N15896, N1766);
buf BUF1 (N15902, N15895);
or OR2 (N15903, N15902, N11192);
not NOT1 (N15904, N15898);
xor XOR2 (N15905, N15900, N14470);
not NOT1 (N15906, N15903);
or OR4 (N15907, N15885, N12220, N14656, N6065);
or OR4 (N15908, N15907, N4757, N4460, N7859);
buf BUF1 (N15909, N15904);
and AND4 (N15910, N15905, N3951, N5038, N12226);
and AND2 (N15911, N15892, N4191);
and AND4 (N15912, N15894, N7439, N4619, N593);
nand NAND3 (N15913, N15911, N3806, N4392);
nor NOR4 (N15914, N15909, N11102, N5791, N2952);
xor XOR2 (N15915, N15888, N13018);
xor XOR2 (N15916, N15912, N12311);
buf BUF1 (N15917, N15908);
buf BUF1 (N15918, N15883);
xor XOR2 (N15919, N15901, N9822);
nor NOR2 (N15920, N15897, N10926);
not NOT1 (N15921, N15917);
not NOT1 (N15922, N15910);
nor NOR3 (N15923, N15913, N7538, N50);
or OR4 (N15924, N15916, N12131, N246, N85);
xor XOR2 (N15925, N15915, N14449);
and AND3 (N15926, N15922, N7286, N660);
nand NAND2 (N15927, N15923, N10847);
or OR4 (N15928, N15914, N8679, N2854, N4146);
xor XOR2 (N15929, N15921, N6718);
nand NAND3 (N15930, N15929, N6456, N9311);
or OR3 (N15931, N15928, N5344, N12037);
not NOT1 (N15932, N15926);
buf BUF1 (N15933, N15925);
and AND2 (N15934, N15906, N7679);
and AND3 (N15935, N15931, N685, N8151);
or OR3 (N15936, N15930, N6484, N2385);
and AND2 (N15937, N15924, N3606);
nor NOR2 (N15938, N15935, N6685);
or OR3 (N15939, N15927, N10588, N1762);
nand NAND2 (N15940, N15918, N14722);
and AND4 (N15941, N15937, N5760, N12371, N6308);
and AND3 (N15942, N15936, N13675, N1438);
or OR3 (N15943, N15942, N1433, N11016);
xor XOR2 (N15944, N15919, N15130);
nand NAND3 (N15945, N15934, N2072, N3817);
not NOT1 (N15946, N15939);
not NOT1 (N15947, N15940);
and AND4 (N15948, N15943, N11146, N6106, N9155);
buf BUF1 (N15949, N15941);
buf BUF1 (N15950, N15920);
and AND4 (N15951, N15947, N535, N1359, N6163);
xor XOR2 (N15952, N15946, N9830);
buf BUF1 (N15953, N15951);
not NOT1 (N15954, N15949);
or OR4 (N15955, N15933, N8675, N11135, N9380);
buf BUF1 (N15956, N15955);
and AND3 (N15957, N15944, N931, N14832);
buf BUF1 (N15958, N15953);
and AND4 (N15959, N15948, N5611, N11520, N3492);
nand NAND4 (N15960, N15957, N152, N6681, N1582);
and AND3 (N15961, N15958, N7426, N1028);
and AND4 (N15962, N15956, N11775, N5280, N8092);
nor NOR4 (N15963, N15959, N15933, N3502, N1228);
or OR4 (N15964, N15938, N2570, N36, N5279);
and AND3 (N15965, N15950, N11567, N13823);
not NOT1 (N15966, N15965);
nand NAND4 (N15967, N15964, N1465, N5882, N15460);
buf BUF1 (N15968, N15967);
or OR2 (N15969, N15968, N7916);
and AND4 (N15970, N15969, N10357, N2171, N12130);
nand NAND2 (N15971, N15962, N14012);
xor XOR2 (N15972, N15954, N11349);
and AND3 (N15973, N15972, N7256, N14203);
xor XOR2 (N15974, N15945, N6702);
nor NOR3 (N15975, N15960, N6979, N1750);
and AND2 (N15976, N15961, N13833);
and AND2 (N15977, N15970, N4785);
not NOT1 (N15978, N15932);
nand NAND4 (N15979, N15973, N532, N4150, N225);
xor XOR2 (N15980, N15975, N9269);
nand NAND4 (N15981, N15974, N7347, N7447, N2319);
nor NOR4 (N15982, N15966, N12493, N8175, N13983);
buf BUF1 (N15983, N15980);
or OR3 (N15984, N15952, N3997, N8762);
buf BUF1 (N15985, N15982);
xor XOR2 (N15986, N15977, N14516);
nor NOR2 (N15987, N15986, N12050);
buf BUF1 (N15988, N15985);
not NOT1 (N15989, N15963);
nor NOR4 (N15990, N15987, N10125, N8413, N11922);
or OR3 (N15991, N15988, N6593, N3408);
not NOT1 (N15992, N15989);
buf BUF1 (N15993, N15984);
buf BUF1 (N15994, N15993);
nand NAND2 (N15995, N15992, N8908);
xor XOR2 (N15996, N15981, N4416);
and AND3 (N15997, N15990, N13860, N5711);
nand NAND2 (N15998, N15997, N15558);
nor NOR4 (N15999, N15976, N5387, N5157, N1372);
xor XOR2 (N16000, N15995, N12723);
buf BUF1 (N16001, N15996);
xor XOR2 (N16002, N15983, N12878);
or OR2 (N16003, N15979, N7159);
nor NOR2 (N16004, N15998, N8228);
buf BUF1 (N16005, N16003);
nor NOR2 (N16006, N15978, N13684);
or OR2 (N16007, N15999, N2967);
and AND2 (N16008, N15971, N10548);
xor XOR2 (N16009, N16004, N4807);
or OR2 (N16010, N16002, N1710);
nor NOR3 (N16011, N15991, N15996, N10983);
not NOT1 (N16012, N16006);
xor XOR2 (N16013, N16009, N7073);
and AND2 (N16014, N16010, N3398);
and AND4 (N16015, N16000, N5441, N91, N11847);
nor NOR3 (N16016, N16005, N10473, N9666);
nand NAND4 (N16017, N16007, N7212, N13041, N6313);
or OR4 (N16018, N15994, N2582, N10271, N3203);
buf BUF1 (N16019, N16013);
and AND4 (N16020, N16018, N98, N6185, N15573);
and AND2 (N16021, N16019, N14715);
nor NOR2 (N16022, N16012, N14278);
buf BUF1 (N16023, N16001);
buf BUF1 (N16024, N16023);
xor XOR2 (N16025, N16021, N223);
buf BUF1 (N16026, N16022);
nand NAND2 (N16027, N16020, N8152);
buf BUF1 (N16028, N16025);
and AND3 (N16029, N16024, N5559, N5757);
buf BUF1 (N16030, N16016);
xor XOR2 (N16031, N16011, N5169);
or OR3 (N16032, N16031, N7129, N9201);
nor NOR2 (N16033, N16026, N5239);
nand NAND3 (N16034, N16033, N1492, N5687);
nor NOR3 (N16035, N16034, N11813, N3717);
and AND2 (N16036, N16035, N15931);
or OR2 (N16037, N16028, N8356);
buf BUF1 (N16038, N16014);
nor NOR4 (N16039, N16038, N9198, N13654, N4847);
nor NOR3 (N16040, N16032, N4555, N8019);
nor NOR2 (N16041, N16030, N707);
nor NOR3 (N16042, N16036, N1574, N12011);
and AND3 (N16043, N16027, N2533, N7584);
not NOT1 (N16044, N16029);
nand NAND4 (N16045, N16008, N4824, N11760, N12023);
not NOT1 (N16046, N16044);
not NOT1 (N16047, N16037);
xor XOR2 (N16048, N16039, N4520);
and AND4 (N16049, N16048, N7479, N2367, N971);
xor XOR2 (N16050, N16046, N6443);
not NOT1 (N16051, N16042);
xor XOR2 (N16052, N16051, N12451);
nand NAND4 (N16053, N16015, N12126, N9299, N12014);
or OR4 (N16054, N16017, N10056, N13452, N3141);
nor NOR3 (N16055, N16047, N11936, N1);
not NOT1 (N16056, N16040);
and AND3 (N16057, N16056, N3155, N4242);
and AND4 (N16058, N16050, N9702, N3884, N11197);
and AND2 (N16059, N16053, N2037);
or OR2 (N16060, N16054, N13524);
not NOT1 (N16061, N16045);
nor NOR4 (N16062, N16061, N3480, N1142, N13625);
not NOT1 (N16063, N16041);
nand NAND4 (N16064, N16055, N1382, N5979, N8015);
xor XOR2 (N16065, N16062, N5620);
nor NOR3 (N16066, N16049, N7337, N9159);
xor XOR2 (N16067, N16064, N5899);
and AND3 (N16068, N16043, N3472, N1210);
not NOT1 (N16069, N16058);
nor NOR2 (N16070, N16059, N5624);
nand NAND4 (N16071, N16060, N14405, N9235, N245);
xor XOR2 (N16072, N16067, N8229);
nor NOR2 (N16073, N16069, N11387);
nor NOR4 (N16074, N16063, N113, N5354, N1654);
buf BUF1 (N16075, N16066);
nor NOR4 (N16076, N16057, N6713, N5868, N14674);
or OR2 (N16077, N16073, N14943);
and AND4 (N16078, N16077, N810, N13035, N4924);
nor NOR4 (N16079, N16052, N7204, N14782, N8654);
and AND4 (N16080, N16068, N1031, N627, N12746);
not NOT1 (N16081, N16075);
nand NAND3 (N16082, N16072, N2364, N650);
and AND3 (N16083, N16074, N788, N4085);
nor NOR4 (N16084, N16071, N3946, N11577, N15833);
nand NAND3 (N16085, N16076, N13389, N6928);
nand NAND4 (N16086, N16082, N6069, N10438, N6372);
or OR4 (N16087, N16070, N1308, N9264, N2606);
and AND3 (N16088, N16083, N14020, N10252);
or OR3 (N16089, N16065, N12139, N8946);
xor XOR2 (N16090, N16084, N12170);
and AND2 (N16091, N16086, N6462);
not NOT1 (N16092, N16088);
nor NOR4 (N16093, N16090, N1984, N3782, N2166);
buf BUF1 (N16094, N16080);
or OR2 (N16095, N16091, N7884);
or OR4 (N16096, N16089, N14782, N2649, N9948);
or OR4 (N16097, N16085, N8880, N11189, N9746);
xor XOR2 (N16098, N16096, N2805);
not NOT1 (N16099, N16097);
and AND4 (N16100, N16087, N5526, N3268, N3957);
or OR4 (N16101, N16079, N8232, N7781, N5709);
or OR3 (N16102, N16093, N15221, N6047);
xor XOR2 (N16103, N16100, N12728);
and AND2 (N16104, N16095, N16051);
nor NOR3 (N16105, N16098, N11287, N5133);
or OR4 (N16106, N16105, N13260, N4281, N7659);
nand NAND4 (N16107, N16102, N9293, N2416, N11829);
xor XOR2 (N16108, N16103, N4147);
nand NAND4 (N16109, N16078, N8683, N14808, N12669);
nand NAND2 (N16110, N16099, N4562);
nor NOR3 (N16111, N16101, N12080, N11546);
buf BUF1 (N16112, N16094);
or OR4 (N16113, N16109, N13463, N1267, N974);
nor NOR4 (N16114, N16107, N991, N893, N6826);
nand NAND4 (N16115, N16110, N380, N6980, N7323);
or OR4 (N16116, N16106, N1777, N9569, N6993);
nor NOR4 (N16117, N16081, N12884, N3372, N3261);
and AND4 (N16118, N16111, N5861, N16062, N5940);
buf BUF1 (N16119, N16113);
buf BUF1 (N16120, N16112);
nor NOR3 (N16121, N16108, N11015, N3426);
nand NAND2 (N16122, N16114, N939);
nor NOR4 (N16123, N16122, N8105, N11183, N6277);
buf BUF1 (N16124, N16123);
xor XOR2 (N16125, N16092, N6500);
xor XOR2 (N16126, N16124, N11877);
nand NAND4 (N16127, N16119, N1260, N15842, N7834);
not NOT1 (N16128, N16116);
nor NOR2 (N16129, N16125, N3883);
nand NAND3 (N16130, N16118, N5394, N1474);
nor NOR4 (N16131, N16128, N3898, N2751, N15654);
nor NOR4 (N16132, N16127, N2526, N6247, N6230);
or OR2 (N16133, N16117, N15501);
xor XOR2 (N16134, N16120, N14174);
not NOT1 (N16135, N16121);
and AND3 (N16136, N16132, N1900, N11294);
nand NAND4 (N16137, N16131, N1761, N13040, N7723);
or OR4 (N16138, N16126, N8770, N1014, N11178);
not NOT1 (N16139, N16135);
and AND2 (N16140, N16138, N12730);
xor XOR2 (N16141, N16129, N9086);
xor XOR2 (N16142, N16134, N10705);
or OR4 (N16143, N16136, N5970, N16132, N11172);
nand NAND4 (N16144, N16130, N14757, N14079, N7216);
buf BUF1 (N16145, N16133);
nor NOR2 (N16146, N16145, N6466);
and AND2 (N16147, N16104, N8063);
not NOT1 (N16148, N16142);
xor XOR2 (N16149, N16137, N6926);
nor NOR4 (N16150, N16144, N3503, N116, N9867);
not NOT1 (N16151, N16147);
not NOT1 (N16152, N16150);
and AND4 (N16153, N16146, N13270, N8845, N7573);
buf BUF1 (N16154, N16115);
or OR4 (N16155, N16154, N3609, N6888, N1876);
and AND2 (N16156, N16140, N13023);
nand NAND3 (N16157, N16156, N4670, N13549);
buf BUF1 (N16158, N16139);
xor XOR2 (N16159, N16157, N1647);
not NOT1 (N16160, N16151);
nor NOR3 (N16161, N16149, N7488, N12081);
nor NOR3 (N16162, N16158, N13873, N3519);
nand NAND3 (N16163, N16153, N12951, N12778);
xor XOR2 (N16164, N16148, N9158);
xor XOR2 (N16165, N16162, N14573);
or OR3 (N16166, N16164, N5647, N1501);
nand NAND3 (N16167, N16163, N4668, N4397);
xor XOR2 (N16168, N16159, N7926);
not NOT1 (N16169, N16161);
nor NOR3 (N16170, N16160, N4790, N15658);
or OR2 (N16171, N16165, N4954);
and AND3 (N16172, N16141, N8268, N6967);
nor NOR3 (N16173, N16155, N10972, N15204);
nor NOR2 (N16174, N16143, N9593);
buf BUF1 (N16175, N16166);
not NOT1 (N16176, N16169);
not NOT1 (N16177, N16175);
xor XOR2 (N16178, N16174, N8935);
and AND3 (N16179, N16176, N1722, N6220);
or OR3 (N16180, N16177, N2024, N12074);
or OR4 (N16181, N16167, N9130, N452, N7300);
nor NOR4 (N16182, N16171, N2739, N7340, N1688);
and AND3 (N16183, N16180, N6115, N12091);
or OR2 (N16184, N16183, N4368);
nand NAND2 (N16185, N16152, N3655);
not NOT1 (N16186, N16185);
nor NOR4 (N16187, N16168, N2006, N12486, N8136);
nor NOR2 (N16188, N16170, N8803);
not NOT1 (N16189, N16173);
buf BUF1 (N16190, N16178);
or OR2 (N16191, N16182, N943);
nor NOR4 (N16192, N16181, N12073, N1660, N15818);
not NOT1 (N16193, N16191);
nor NOR3 (N16194, N16188, N4918, N6563);
and AND2 (N16195, N16184, N7357);
xor XOR2 (N16196, N16172, N628);
nand NAND4 (N16197, N16195, N11786, N12500, N14387);
buf BUF1 (N16198, N16192);
xor XOR2 (N16199, N16197, N4284);
buf BUF1 (N16200, N16187);
xor XOR2 (N16201, N16190, N7526);
nand NAND3 (N16202, N16201, N10729, N14392);
xor XOR2 (N16203, N16186, N1054);
buf BUF1 (N16204, N16189);
and AND3 (N16205, N16193, N2924, N314);
xor XOR2 (N16206, N16199, N13032);
not NOT1 (N16207, N16203);
nor NOR2 (N16208, N16198, N3669);
nor NOR3 (N16209, N16206, N8781, N9995);
not NOT1 (N16210, N16209);
nor NOR3 (N16211, N16204, N864, N3339);
nand NAND4 (N16212, N16200, N4538, N7316, N9087);
and AND3 (N16213, N16212, N12768, N3747);
buf BUF1 (N16214, N16211);
nand NAND3 (N16215, N16202, N4234, N15786);
nor NOR2 (N16216, N16205, N6209);
not NOT1 (N16217, N16207);
not NOT1 (N16218, N16217);
xor XOR2 (N16219, N16213, N6656);
or OR4 (N16220, N16210, N768, N9658, N3730);
not NOT1 (N16221, N16219);
buf BUF1 (N16222, N16194);
and AND4 (N16223, N16222, N10355, N14061, N1789);
nor NOR4 (N16224, N16215, N1936, N11902, N11416);
xor XOR2 (N16225, N16221, N2481);
not NOT1 (N16226, N16216);
not NOT1 (N16227, N16208);
xor XOR2 (N16228, N16214, N807);
buf BUF1 (N16229, N16226);
or OR2 (N16230, N16229, N7476);
and AND4 (N16231, N16223, N7321, N8663, N2479);
not NOT1 (N16232, N16227);
or OR2 (N16233, N16225, N8896);
xor XOR2 (N16234, N16218, N8392);
xor XOR2 (N16235, N16230, N11212);
not NOT1 (N16236, N16233);
nor NOR2 (N16237, N16235, N1917);
and AND3 (N16238, N16179, N13724, N6574);
or OR2 (N16239, N16228, N12705);
nor NOR2 (N16240, N16224, N5206);
or OR3 (N16241, N16236, N13832, N1611);
or OR3 (N16242, N16241, N1102, N11904);
and AND4 (N16243, N16240, N6008, N11096, N2613);
buf BUF1 (N16244, N16232);
xor XOR2 (N16245, N16244, N15734);
not NOT1 (N16246, N16245);
and AND4 (N16247, N16231, N7595, N13832, N139);
or OR2 (N16248, N16237, N12638);
nand NAND4 (N16249, N16242, N13357, N15981, N14323);
nor NOR4 (N16250, N16249, N266, N7961, N2316);
or OR2 (N16251, N16238, N775);
buf BUF1 (N16252, N16220);
or OR3 (N16253, N16246, N2884, N15442);
buf BUF1 (N16254, N16248);
or OR3 (N16255, N16254, N10996, N10798);
or OR3 (N16256, N16247, N13283, N11577);
nand NAND3 (N16257, N16196, N928, N5061);
and AND2 (N16258, N16253, N1602);
not NOT1 (N16259, N16243);
and AND3 (N16260, N16250, N2246, N15711);
or OR3 (N16261, N16251, N12410, N12908);
not NOT1 (N16262, N16261);
or OR3 (N16263, N16257, N5735, N9623);
or OR4 (N16264, N16239, N7183, N6348, N13675);
not NOT1 (N16265, N16234);
nand NAND4 (N16266, N16260, N12400, N8572, N14222);
not NOT1 (N16267, N16263);
nand NAND3 (N16268, N16267, N3111, N8500);
nor NOR2 (N16269, N16262, N12504);
nand NAND4 (N16270, N16268, N13005, N13453, N10013);
or OR3 (N16271, N16270, N13088, N7329);
not NOT1 (N16272, N16266);
or OR2 (N16273, N16258, N4592);
or OR3 (N16274, N16259, N9386, N14438);
and AND2 (N16275, N16273, N5526);
and AND3 (N16276, N16274, N1666, N12989);
nor NOR2 (N16277, N16265, N8406);
nor NOR2 (N16278, N16269, N11687);
nand NAND4 (N16279, N16278, N12217, N8874, N10179);
nand NAND2 (N16280, N16252, N413);
nand NAND2 (N16281, N16277, N10249);
buf BUF1 (N16282, N16276);
nor NOR2 (N16283, N16256, N3341);
nand NAND4 (N16284, N16281, N8174, N11909, N4087);
not NOT1 (N16285, N16255);
and AND2 (N16286, N16284, N13165);
xor XOR2 (N16287, N16271, N597);
xor XOR2 (N16288, N16282, N2380);
nor NOR3 (N16289, N16264, N10969, N9442);
or OR2 (N16290, N16289, N10084);
not NOT1 (N16291, N16275);
nand NAND4 (N16292, N16291, N12258, N1114, N10926);
and AND3 (N16293, N16288, N15762, N11864);
buf BUF1 (N16294, N16290);
and AND4 (N16295, N16285, N12552, N12145, N4570);
and AND3 (N16296, N16287, N4062, N3991);
nor NOR2 (N16297, N16295, N11691);
xor XOR2 (N16298, N16286, N13230);
or OR3 (N16299, N16296, N15589, N7821);
nor NOR3 (N16300, N16280, N12761, N12222);
xor XOR2 (N16301, N16272, N12079);
or OR2 (N16302, N16298, N9573);
xor XOR2 (N16303, N16300, N5136);
and AND3 (N16304, N16302, N12616, N3941);
not NOT1 (N16305, N16294);
nand NAND2 (N16306, N16292, N6612);
xor XOR2 (N16307, N16305, N667);
buf BUF1 (N16308, N16306);
and AND3 (N16309, N16308, N6237, N1702);
not NOT1 (N16310, N16297);
not NOT1 (N16311, N16309);
xor XOR2 (N16312, N16311, N13992);
and AND4 (N16313, N16299, N13864, N10287, N5971);
nand NAND3 (N16314, N16312, N7833, N5929);
or OR2 (N16315, N16307, N7261);
xor XOR2 (N16316, N16313, N6407);
nor NOR3 (N16317, N16304, N14045, N3863);
nand NAND3 (N16318, N16310, N7389, N6001);
nor NOR2 (N16319, N16303, N15711);
buf BUF1 (N16320, N16316);
and AND2 (N16321, N16318, N15629);
not NOT1 (N16322, N16321);
or OR4 (N16323, N16317, N15037, N6087, N7421);
xor XOR2 (N16324, N16319, N940);
nand NAND4 (N16325, N16279, N12185, N2444, N1433);
nand NAND4 (N16326, N16323, N8168, N9212, N4909);
buf BUF1 (N16327, N16325);
or OR4 (N16328, N16315, N4766, N13433, N1554);
not NOT1 (N16329, N16314);
xor XOR2 (N16330, N16293, N14294);
nand NAND4 (N16331, N16326, N7104, N10994, N5991);
nand NAND4 (N16332, N16324, N11073, N1663, N8386);
and AND3 (N16333, N16329, N12991, N4792);
and AND3 (N16334, N16320, N8583, N7306);
or OR3 (N16335, N16283, N10999, N6922);
or OR4 (N16336, N16335, N10571, N2308, N5979);
xor XOR2 (N16337, N16333, N104);
nor NOR2 (N16338, N16332, N949);
nand NAND3 (N16339, N16336, N11151, N12718);
buf BUF1 (N16340, N16330);
nand NAND2 (N16341, N16334, N12582);
xor XOR2 (N16342, N16322, N12469);
nand NAND4 (N16343, N16340, N1854, N16227, N10232);
not NOT1 (N16344, N16337);
xor XOR2 (N16345, N16328, N6545);
and AND4 (N16346, N16345, N15919, N15060, N15308);
and AND3 (N16347, N16341, N14272, N565);
or OR2 (N16348, N16331, N14774);
xor XOR2 (N16349, N16348, N13731);
nor NOR4 (N16350, N16342, N4893, N2730, N780);
buf BUF1 (N16351, N16301);
buf BUF1 (N16352, N16349);
nand NAND2 (N16353, N16352, N16140);
and AND2 (N16354, N16339, N8409);
not NOT1 (N16355, N16350);
xor XOR2 (N16356, N16343, N8924);
and AND2 (N16357, N16338, N11055);
not NOT1 (N16358, N16354);
or OR2 (N16359, N16344, N4583);
and AND2 (N16360, N16353, N2279);
nand NAND3 (N16361, N16357, N6454, N9028);
xor XOR2 (N16362, N16347, N12744);
buf BUF1 (N16363, N16355);
nand NAND3 (N16364, N16362, N9364, N180);
nor NOR4 (N16365, N16361, N12460, N11257, N5047);
or OR4 (N16366, N16346, N11389, N4597, N4576);
buf BUF1 (N16367, N16365);
not NOT1 (N16368, N16360);
or OR2 (N16369, N16358, N6626);
buf BUF1 (N16370, N16351);
or OR4 (N16371, N16327, N16018, N7081, N2538);
and AND2 (N16372, N16366, N16346);
nor NOR3 (N16373, N16364, N14441, N5920);
and AND2 (N16374, N16370, N4015);
or OR2 (N16375, N16372, N10957);
buf BUF1 (N16376, N16356);
or OR4 (N16377, N16373, N3716, N10592, N13272);
buf BUF1 (N16378, N16371);
and AND3 (N16379, N16363, N3048, N9006);
or OR3 (N16380, N16376, N13440, N6557);
not NOT1 (N16381, N16369);
and AND3 (N16382, N16374, N9356, N12889);
buf BUF1 (N16383, N16379);
buf BUF1 (N16384, N16377);
not NOT1 (N16385, N16382);
nand NAND3 (N16386, N16384, N4493, N5230);
nand NAND2 (N16387, N16385, N5132);
or OR2 (N16388, N16387, N11486);
and AND4 (N16389, N16359, N5772, N5775, N2937);
not NOT1 (N16390, N16381);
buf BUF1 (N16391, N16383);
and AND2 (N16392, N16388, N14736);
buf BUF1 (N16393, N16378);
nand NAND3 (N16394, N16386, N14063, N5481);
or OR3 (N16395, N16375, N4367, N2423);
nor NOR2 (N16396, N16389, N2285);
not NOT1 (N16397, N16393);
xor XOR2 (N16398, N16392, N16333);
buf BUF1 (N16399, N16397);
nor NOR2 (N16400, N16395, N8035);
not NOT1 (N16401, N16367);
and AND4 (N16402, N16380, N5756, N15198, N5672);
and AND2 (N16403, N16391, N9217);
or OR2 (N16404, N16390, N2067);
not NOT1 (N16405, N16404);
xor XOR2 (N16406, N16402, N5747);
not NOT1 (N16407, N16398);
and AND2 (N16408, N16400, N8418);
or OR4 (N16409, N16368, N5495, N7151, N5376);
nand NAND4 (N16410, N16409, N3332, N1384, N11389);
not NOT1 (N16411, N16394);
xor XOR2 (N16412, N16405, N3089);
nor NOR4 (N16413, N16403, N948, N6461, N5763);
nand NAND3 (N16414, N16399, N1495, N8267);
not NOT1 (N16415, N16412);
and AND4 (N16416, N16415, N4923, N5461, N15925);
nor NOR4 (N16417, N16407, N2396, N10624, N15037);
nor NOR4 (N16418, N16417, N2113, N5528, N335);
nand NAND2 (N16419, N16401, N566);
xor XOR2 (N16420, N16413, N12925);
xor XOR2 (N16421, N16416, N4659);
xor XOR2 (N16422, N16420, N10761);
nor NOR2 (N16423, N16418, N2889);
nor NOR4 (N16424, N16411, N1148, N9172, N7734);
not NOT1 (N16425, N16424);
nand NAND4 (N16426, N16410, N7027, N5329, N393);
or OR3 (N16427, N16414, N12224, N7543);
or OR3 (N16428, N16396, N8454, N12437);
nand NAND2 (N16429, N16427, N6655);
nor NOR2 (N16430, N16426, N3406);
xor XOR2 (N16431, N16406, N12052);
nor NOR4 (N16432, N16419, N11465, N14672, N4682);
xor XOR2 (N16433, N16429, N11742);
or OR2 (N16434, N16431, N7827);
buf BUF1 (N16435, N16428);
not NOT1 (N16436, N16425);
not NOT1 (N16437, N16435);
nor NOR4 (N16438, N16432, N6478, N11718, N10777);
nor NOR2 (N16439, N16423, N12207);
or OR2 (N16440, N16408, N15925);
not NOT1 (N16441, N16438);
nand NAND2 (N16442, N16437, N12620);
and AND3 (N16443, N16433, N5305, N3613);
not NOT1 (N16444, N16434);
or OR2 (N16445, N16442, N749);
buf BUF1 (N16446, N16421);
or OR4 (N16447, N16445, N6612, N6795, N4832);
buf BUF1 (N16448, N16446);
and AND2 (N16449, N16422, N12037);
buf BUF1 (N16450, N16443);
nor NOR4 (N16451, N16444, N10374, N2109, N737);
or OR3 (N16452, N16449, N13260, N9815);
xor XOR2 (N16453, N16441, N708);
xor XOR2 (N16454, N16439, N8644);
or OR3 (N16455, N16451, N11683, N11081);
nand NAND3 (N16456, N16454, N13691, N6959);
not NOT1 (N16457, N16430);
not NOT1 (N16458, N16436);
xor XOR2 (N16459, N16440, N3367);
not NOT1 (N16460, N16457);
xor XOR2 (N16461, N16453, N8087);
xor XOR2 (N16462, N16450, N296);
not NOT1 (N16463, N16456);
xor XOR2 (N16464, N16447, N11590);
nor NOR2 (N16465, N16459, N11937);
or OR4 (N16466, N16463, N2094, N7679, N3545);
or OR3 (N16467, N16460, N15748, N4580);
xor XOR2 (N16468, N16452, N7867);
and AND3 (N16469, N16462, N9115, N14856);
and AND4 (N16470, N16464, N1020, N231, N2814);
not NOT1 (N16471, N16466);
xor XOR2 (N16472, N16468, N8219);
nand NAND2 (N16473, N16469, N4565);
or OR4 (N16474, N16470, N9453, N12581, N4274);
nor NOR2 (N16475, N16471, N42);
nor NOR4 (N16476, N16474, N5654, N8145, N1337);
not NOT1 (N16477, N16473);
nand NAND3 (N16478, N16461, N12525, N15515);
nor NOR2 (N16479, N16465, N3919);
not NOT1 (N16480, N16478);
nand NAND3 (N16481, N16455, N13809, N9370);
xor XOR2 (N16482, N16479, N11825);
nand NAND4 (N16483, N16467, N14434, N13938, N3592);
and AND3 (N16484, N16458, N10585, N10281);
nor NOR2 (N16485, N16472, N12346);
nor NOR2 (N16486, N16485, N8169);
nand NAND3 (N16487, N16475, N1257, N12758);
nand NAND4 (N16488, N16448, N14501, N10993, N9536);
not NOT1 (N16489, N16486);
buf BUF1 (N16490, N16484);
or OR4 (N16491, N16490, N5510, N11212, N8690);
nand NAND2 (N16492, N16481, N13236);
nor NOR3 (N16493, N16482, N11173, N8289);
nor NOR4 (N16494, N16489, N13182, N13661, N5886);
nor NOR3 (N16495, N16477, N12037, N11189);
nand NAND3 (N16496, N16491, N15025, N15587);
xor XOR2 (N16497, N16493, N1535);
nor NOR3 (N16498, N16483, N10470, N5242);
nand NAND3 (N16499, N16494, N9123, N10190);
nor NOR3 (N16500, N16495, N3630, N6733);
nand NAND4 (N16501, N16500, N3686, N3885, N5468);
nor NOR2 (N16502, N16492, N10323);
and AND2 (N16503, N16498, N5642);
nand NAND3 (N16504, N16488, N7625, N11563);
and AND3 (N16505, N16502, N12129, N7660);
not NOT1 (N16506, N16497);
buf BUF1 (N16507, N16501);
not NOT1 (N16508, N16503);
nand NAND3 (N16509, N16487, N2295, N9591);
buf BUF1 (N16510, N16505);
not NOT1 (N16511, N16510);
nand NAND3 (N16512, N16506, N16200, N13940);
buf BUF1 (N16513, N16476);
buf BUF1 (N16514, N16504);
nor NOR2 (N16515, N16507, N12738);
or OR3 (N16516, N16511, N7729, N2384);
or OR3 (N16517, N16516, N13964, N563);
and AND2 (N16518, N16508, N12497);
or OR2 (N16519, N16509, N7349);
not NOT1 (N16520, N16517);
or OR3 (N16521, N16514, N11013, N5420);
and AND4 (N16522, N16513, N12166, N11336, N1476);
and AND3 (N16523, N16519, N986, N10110);
and AND4 (N16524, N16523, N4644, N9697, N6490);
nand NAND3 (N16525, N16512, N13713, N771);
nand NAND3 (N16526, N16480, N15232, N12294);
or OR3 (N16527, N16522, N439, N3195);
not NOT1 (N16528, N16499);
buf BUF1 (N16529, N16496);
xor XOR2 (N16530, N16528, N8322);
buf BUF1 (N16531, N16524);
buf BUF1 (N16532, N16518);
nand NAND3 (N16533, N16532, N12759, N2671);
or OR4 (N16534, N16529, N9834, N10367, N235);
not NOT1 (N16535, N16521);
not NOT1 (N16536, N16515);
and AND4 (N16537, N16520, N6484, N16090, N4393);
or OR4 (N16538, N16526, N8042, N12250, N9474);
buf BUF1 (N16539, N16533);
and AND2 (N16540, N16531, N5877);
nor NOR3 (N16541, N16530, N971, N7349);
or OR3 (N16542, N16540, N16395, N1581);
buf BUF1 (N16543, N16527);
not NOT1 (N16544, N16542);
nor NOR3 (N16545, N16536, N728, N9099);
nand NAND2 (N16546, N16541, N7473);
or OR4 (N16547, N16545, N10489, N13003, N814);
and AND3 (N16548, N16535, N844, N2171);
not NOT1 (N16549, N16538);
nand NAND4 (N16550, N16537, N8912, N4343, N9645);
or OR3 (N16551, N16543, N13327, N5018);
nor NOR3 (N16552, N16550, N6801, N10428);
nor NOR2 (N16553, N16551, N9005);
xor XOR2 (N16554, N16547, N15985);
nand NAND4 (N16555, N16546, N5095, N2391, N2479);
not NOT1 (N16556, N16554);
xor XOR2 (N16557, N16556, N6396);
not NOT1 (N16558, N16525);
or OR3 (N16559, N16552, N12005, N11572);
and AND3 (N16560, N16534, N5941, N10132);
buf BUF1 (N16561, N16548);
buf BUF1 (N16562, N16553);
nor NOR4 (N16563, N16555, N7422, N10848, N11684);
buf BUF1 (N16564, N16557);
not NOT1 (N16565, N16560);
xor XOR2 (N16566, N16562, N9707);
not NOT1 (N16567, N16539);
nand NAND3 (N16568, N16558, N14672, N11673);
xor XOR2 (N16569, N16544, N10294);
buf BUF1 (N16570, N16564);
xor XOR2 (N16571, N16567, N6448);
and AND3 (N16572, N16571, N713, N9100);
buf BUF1 (N16573, N16572);
nand NAND4 (N16574, N16568, N5083, N1018, N13536);
xor XOR2 (N16575, N16569, N12487);
xor XOR2 (N16576, N16573, N15887);
nand NAND4 (N16577, N16574, N358, N11443, N10682);
and AND2 (N16578, N16559, N6359);
and AND3 (N16579, N16549, N5347, N22);
xor XOR2 (N16580, N16575, N712);
nor NOR2 (N16581, N16579, N15535);
nor NOR3 (N16582, N16570, N6881, N21);
nand NAND2 (N16583, N16563, N5428);
nand NAND2 (N16584, N16581, N15685);
not NOT1 (N16585, N16583);
nand NAND4 (N16586, N16576, N3412, N14395, N5133);
or OR4 (N16587, N16565, N187, N8659, N7838);
buf BUF1 (N16588, N16566);
nand NAND4 (N16589, N16586, N4490, N9479, N8538);
nor NOR3 (N16590, N16561, N13853, N8190);
nand NAND3 (N16591, N16587, N12787, N10073);
nor NOR4 (N16592, N16578, N16341, N2253, N7990);
nand NAND3 (N16593, N16592, N1985, N10151);
or OR2 (N16594, N16577, N8359);
buf BUF1 (N16595, N16582);
nor NOR4 (N16596, N16580, N14843, N1459, N3595);
buf BUF1 (N16597, N16593);
or OR2 (N16598, N16597, N4760);
buf BUF1 (N16599, N16584);
xor XOR2 (N16600, N16594, N718);
nand NAND3 (N16601, N16595, N530, N7909);
nand NAND3 (N16602, N16588, N7407, N11185);
or OR4 (N16603, N16596, N11482, N13088, N7704);
and AND4 (N16604, N16601, N16025, N8702, N491);
buf BUF1 (N16605, N16598);
nand NAND2 (N16606, N16603, N13496);
nor NOR3 (N16607, N16599, N16260, N12089);
nor NOR3 (N16608, N16585, N5133, N16067);
or OR2 (N16609, N16589, N9205);
nand NAND2 (N16610, N16600, N1973);
xor XOR2 (N16611, N16610, N2553);
nand NAND3 (N16612, N16590, N9735, N7334);
or OR2 (N16613, N16606, N8323);
or OR3 (N16614, N16608, N11776, N11759);
buf BUF1 (N16615, N16611);
nor NOR3 (N16616, N16591, N8378, N8275);
nor NOR4 (N16617, N16614, N2663, N9161, N14206);
or OR3 (N16618, N16612, N1251, N11660);
nand NAND2 (N16619, N16617, N2697);
nor NOR4 (N16620, N16609, N12731, N5867, N5730);
xor XOR2 (N16621, N16618, N12236);
or OR2 (N16622, N16613, N15866);
xor XOR2 (N16623, N16605, N3149);
not NOT1 (N16624, N16616);
buf BUF1 (N16625, N16619);
and AND3 (N16626, N16602, N6016, N12529);
nand NAND3 (N16627, N16623, N5263, N10277);
xor XOR2 (N16628, N16624, N16519);
and AND4 (N16629, N16626, N6732, N790, N2796);
nand NAND2 (N16630, N16607, N4221);
xor XOR2 (N16631, N16629, N9279);
and AND3 (N16632, N16625, N3084, N10096);
and AND3 (N16633, N16620, N13519, N8349);
not NOT1 (N16634, N16630);
and AND4 (N16635, N16621, N636, N4262, N10980);
xor XOR2 (N16636, N16635, N7217);
xor XOR2 (N16637, N16627, N14606);
buf BUF1 (N16638, N16631);
or OR4 (N16639, N16637, N2126, N704, N9687);
and AND3 (N16640, N16638, N3620, N9456);
not NOT1 (N16641, N16615);
buf BUF1 (N16642, N16636);
xor XOR2 (N16643, N16604, N3503);
nor NOR2 (N16644, N16628, N789);
buf BUF1 (N16645, N16640);
nand NAND3 (N16646, N16639, N5219, N14652);
not NOT1 (N16647, N16645);
nor NOR3 (N16648, N16622, N4135, N7811);
not NOT1 (N16649, N16641);
and AND4 (N16650, N16649, N11352, N15185, N9533);
nand NAND4 (N16651, N16633, N12046, N13418, N5176);
buf BUF1 (N16652, N16651);
and AND2 (N16653, N16634, N1771);
xor XOR2 (N16654, N16653, N13552);
or OR3 (N16655, N16643, N8128, N546);
nor NOR3 (N16656, N16655, N13654, N12341);
and AND4 (N16657, N16646, N15221, N2013, N12554);
nand NAND2 (N16658, N16642, N7379);
and AND2 (N16659, N16657, N1159);
or OR3 (N16660, N16644, N11694, N15834);
nand NAND3 (N16661, N16648, N10619, N16062);
xor XOR2 (N16662, N16654, N4763);
nand NAND2 (N16663, N16652, N9589);
buf BUF1 (N16664, N16656);
xor XOR2 (N16665, N16663, N5547);
nor NOR2 (N16666, N16660, N2223);
buf BUF1 (N16667, N16650);
and AND2 (N16668, N16667, N2697);
buf BUF1 (N16669, N16664);
nand NAND2 (N16670, N16632, N15236);
nand NAND4 (N16671, N16668, N1760, N8706, N13039);
xor XOR2 (N16672, N16669, N5015);
not NOT1 (N16673, N16665);
nand NAND4 (N16674, N16662, N6872, N16373, N2835);
xor XOR2 (N16675, N16671, N5311);
xor XOR2 (N16676, N16675, N4222);
or OR2 (N16677, N16674, N14320);
not NOT1 (N16678, N16666);
nor NOR3 (N16679, N16672, N7064, N16242);
and AND4 (N16680, N16647, N5988, N1779, N6390);
nor NOR2 (N16681, N16678, N16084);
and AND3 (N16682, N16673, N8396, N15917);
or OR4 (N16683, N16679, N10121, N3235, N3692);
or OR3 (N16684, N16676, N1705, N1468);
nand NAND4 (N16685, N16661, N4732, N5167, N4010);
xor XOR2 (N16686, N16670, N16446);
or OR2 (N16687, N16683, N11160);
xor XOR2 (N16688, N16687, N10130);
buf BUF1 (N16689, N16677);
nand NAND3 (N16690, N16685, N14534, N2552);
buf BUF1 (N16691, N16682);
nand NAND3 (N16692, N16686, N1631, N11860);
not NOT1 (N16693, N16692);
and AND2 (N16694, N16688, N1419);
or OR3 (N16695, N16693, N1736, N5766);
nor NOR2 (N16696, N16691, N12747);
or OR3 (N16697, N16696, N6379, N3599);
buf BUF1 (N16698, N16681);
xor XOR2 (N16699, N16680, N4254);
xor XOR2 (N16700, N16695, N9428);
nand NAND2 (N16701, N16699, N5479);
nand NAND4 (N16702, N16659, N8588, N12740, N13154);
nand NAND2 (N16703, N16698, N4714);
not NOT1 (N16704, N16684);
buf BUF1 (N16705, N16690);
not NOT1 (N16706, N16694);
not NOT1 (N16707, N16689);
xor XOR2 (N16708, N16701, N15274);
and AND3 (N16709, N16697, N15919, N12410);
nor NOR4 (N16710, N16703, N5312, N10293, N14533);
not NOT1 (N16711, N16704);
or OR4 (N16712, N16710, N2043, N12424, N725);
nor NOR3 (N16713, N16658, N2467, N9830);
nor NOR3 (N16714, N16712, N6279, N3149);
and AND2 (N16715, N16711, N3940);
not NOT1 (N16716, N16706);
nor NOR4 (N16717, N16714, N7564, N3168, N16247);
nand NAND3 (N16718, N16700, N12102, N11395);
xor XOR2 (N16719, N16709, N4499);
not NOT1 (N16720, N16716);
nand NAND4 (N16721, N16713, N3645, N14495, N416);
or OR3 (N16722, N16705, N12849, N11954);
nor NOR4 (N16723, N16719, N16584, N5273, N12385);
and AND4 (N16724, N16722, N440, N10137, N10940);
xor XOR2 (N16725, N16707, N8333);
and AND3 (N16726, N16708, N4807, N209);
nand NAND4 (N16727, N16720, N15359, N2678, N11237);
or OR3 (N16728, N16724, N9481, N12836);
not NOT1 (N16729, N16727);
buf BUF1 (N16730, N16715);
nand NAND4 (N16731, N16730, N6609, N10349, N13387);
or OR3 (N16732, N16728, N8658, N7819);
or OR3 (N16733, N16729, N16681, N12792);
nand NAND4 (N16734, N16717, N3954, N11724, N3331);
or OR2 (N16735, N16731, N9965);
nand NAND3 (N16736, N16733, N13275, N11969);
or OR3 (N16737, N16702, N337, N5435);
buf BUF1 (N16738, N16723);
and AND2 (N16739, N16736, N12645);
xor XOR2 (N16740, N16725, N4567);
buf BUF1 (N16741, N16721);
buf BUF1 (N16742, N16734);
buf BUF1 (N16743, N16718);
or OR4 (N16744, N16735, N2856, N5812, N182);
nor NOR3 (N16745, N16741, N15987, N3107);
xor XOR2 (N16746, N16737, N12129);
xor XOR2 (N16747, N16745, N1107);
or OR3 (N16748, N16744, N15403, N15229);
buf BUF1 (N16749, N16732);
nand NAND4 (N16750, N16742, N7707, N5605, N14518);
nand NAND2 (N16751, N16743, N14101);
and AND2 (N16752, N16739, N10552);
buf BUF1 (N16753, N16752);
or OR4 (N16754, N16726, N5395, N547, N15916);
or OR4 (N16755, N16753, N193, N6686, N2680);
or OR3 (N16756, N16754, N10540, N14130);
nor NOR3 (N16757, N16756, N3245, N13645);
nand NAND4 (N16758, N16746, N13963, N10814, N8392);
nand NAND4 (N16759, N16757, N11180, N7598, N1161);
and AND3 (N16760, N16738, N8119, N13431);
and AND4 (N16761, N16750, N4269, N777, N6285);
xor XOR2 (N16762, N16749, N15745);
nand NAND4 (N16763, N16740, N2414, N8328, N8941);
buf BUF1 (N16764, N16748);
not NOT1 (N16765, N16760);
nor NOR3 (N16766, N16751, N11616, N8374);
xor XOR2 (N16767, N16766, N1379);
buf BUF1 (N16768, N16765);
nor NOR3 (N16769, N16758, N10323, N10965);
nor NOR3 (N16770, N16755, N10959, N15698);
buf BUF1 (N16771, N16762);
xor XOR2 (N16772, N16769, N13953);
or OR3 (N16773, N16764, N14193, N12905);
not NOT1 (N16774, N16773);
nand NAND2 (N16775, N16747, N5324);
and AND3 (N16776, N16775, N1830, N9718);
nand NAND2 (N16777, N16771, N10471);
nand NAND2 (N16778, N16761, N3427);
nand NAND3 (N16779, N16770, N11710, N7873);
not NOT1 (N16780, N16776);
buf BUF1 (N16781, N16779);
nand NAND4 (N16782, N16778, N2603, N13534, N7278);
nor NOR4 (N16783, N16759, N12065, N2848, N7453);
nor NOR2 (N16784, N16780, N5107);
and AND2 (N16785, N16763, N10097);
and AND2 (N16786, N16774, N4894);
nor NOR4 (N16787, N16785, N10760, N2607, N15547);
not NOT1 (N16788, N16772);
and AND2 (N16789, N16768, N8756);
not NOT1 (N16790, N16767);
not NOT1 (N16791, N16787);
nand NAND3 (N16792, N16781, N3387, N11258);
nor NOR4 (N16793, N16789, N15701, N3167, N10075);
xor XOR2 (N16794, N16790, N14762);
and AND4 (N16795, N16784, N1847, N14098, N2970);
and AND2 (N16796, N16786, N15555);
nor NOR3 (N16797, N16793, N16121, N4718);
not NOT1 (N16798, N16797);
nor NOR3 (N16799, N16792, N6855, N9894);
and AND2 (N16800, N16783, N5517);
nand NAND2 (N16801, N16800, N2534);
not NOT1 (N16802, N16799);
and AND2 (N16803, N16802, N6365);
or OR3 (N16804, N16795, N9096, N11402);
xor XOR2 (N16805, N16791, N1735);
nor NOR2 (N16806, N16803, N10006);
or OR3 (N16807, N16796, N8721, N16543);
not NOT1 (N16808, N16804);
and AND4 (N16809, N16782, N5767, N5040, N9729);
nand NAND2 (N16810, N16807, N11961);
nor NOR3 (N16811, N16798, N13341, N4943);
nor NOR3 (N16812, N16805, N12091, N2005);
and AND2 (N16813, N16811, N15499);
or OR4 (N16814, N16810, N2351, N15134, N15754);
not NOT1 (N16815, N16801);
xor XOR2 (N16816, N16815, N5891);
nor NOR3 (N16817, N16806, N9717, N7431);
buf BUF1 (N16818, N16809);
not NOT1 (N16819, N16788);
not NOT1 (N16820, N16817);
nand NAND4 (N16821, N16814, N10306, N8234, N16753);
not NOT1 (N16822, N16816);
nor NOR2 (N16823, N16794, N11121);
nor NOR2 (N16824, N16777, N5455);
and AND3 (N16825, N16820, N1803, N5294);
or OR3 (N16826, N16824, N1610, N4232);
xor XOR2 (N16827, N16812, N522);
buf BUF1 (N16828, N16808);
nor NOR3 (N16829, N16818, N14029, N11408);
not NOT1 (N16830, N16827);
or OR3 (N16831, N16819, N266, N15826);
nor NOR4 (N16832, N16828, N14874, N1138, N10646);
and AND4 (N16833, N16830, N12559, N10912, N6688);
nor NOR4 (N16834, N16831, N12452, N15828, N3379);
nand NAND2 (N16835, N16825, N10183);
nor NOR2 (N16836, N16833, N6323);
nor NOR4 (N16837, N16822, N7947, N12702, N642);
buf BUF1 (N16838, N16813);
or OR4 (N16839, N16832, N14466, N15142, N11780);
nand NAND3 (N16840, N16835, N7958, N15778);
nand NAND2 (N16841, N16839, N6757);
xor XOR2 (N16842, N16841, N11301);
and AND3 (N16843, N16836, N2156, N11530);
or OR3 (N16844, N16829, N13672, N2495);
buf BUF1 (N16845, N16821);
and AND3 (N16846, N16843, N3903, N15690);
and AND2 (N16847, N16838, N3409);
not NOT1 (N16848, N16834);
not NOT1 (N16849, N16848);
or OR2 (N16850, N16849, N13668);
buf BUF1 (N16851, N16844);
buf BUF1 (N16852, N16840);
not NOT1 (N16853, N16845);
xor XOR2 (N16854, N16826, N15775);
not NOT1 (N16855, N16853);
xor XOR2 (N16856, N16842, N9187);
buf BUF1 (N16857, N16852);
not NOT1 (N16858, N16850);
xor XOR2 (N16859, N16855, N10019);
not NOT1 (N16860, N16847);
xor XOR2 (N16861, N16837, N3427);
or OR4 (N16862, N16823, N5087, N3741, N10288);
nor NOR3 (N16863, N16862, N5076, N15781);
or OR4 (N16864, N16856, N1274, N5100, N4731);
nand NAND2 (N16865, N16859, N9850);
nand NAND4 (N16866, N16851, N15722, N11376, N638);
or OR4 (N16867, N16858, N9261, N7296, N6055);
nor NOR4 (N16868, N16846, N12507, N293, N13168);
not NOT1 (N16869, N16860);
buf BUF1 (N16870, N16857);
and AND2 (N16871, N16863, N461);
nor NOR4 (N16872, N16866, N8066, N11643, N5768);
xor XOR2 (N16873, N16865, N4055);
and AND4 (N16874, N16868, N551, N11233, N13657);
not NOT1 (N16875, N16874);
xor XOR2 (N16876, N16871, N5544);
or OR4 (N16877, N16861, N15622, N4482, N10962);
or OR4 (N16878, N16867, N13157, N12278, N5556);
nor NOR2 (N16879, N16869, N6471);
or OR4 (N16880, N16873, N6055, N1050, N15319);
or OR2 (N16881, N16875, N7387);
nand NAND2 (N16882, N16879, N8853);
nor NOR4 (N16883, N16880, N5049, N6678, N6677);
or OR4 (N16884, N16870, N3599, N8364, N12607);
not NOT1 (N16885, N16854);
not NOT1 (N16886, N16864);
and AND4 (N16887, N16885, N11303, N6314, N9126);
and AND4 (N16888, N16882, N6784, N15418, N8974);
and AND4 (N16889, N16888, N14272, N10304, N10044);
or OR3 (N16890, N16877, N15197, N684);
buf BUF1 (N16891, N16883);
and AND4 (N16892, N16884, N10527, N14279, N16004);
nor NOR3 (N16893, N16881, N11887, N1726);
nor NOR3 (N16894, N16878, N10525, N2118);
or OR2 (N16895, N16894, N4426);
buf BUF1 (N16896, N16876);
xor XOR2 (N16897, N16891, N6847);
nor NOR4 (N16898, N16895, N255, N15939, N9706);
nor NOR2 (N16899, N16886, N11808);
not NOT1 (N16900, N16892);
xor XOR2 (N16901, N16872, N8768);
buf BUF1 (N16902, N16899);
and AND4 (N16903, N16887, N4501, N15681, N4544);
not NOT1 (N16904, N16889);
or OR3 (N16905, N16901, N10357, N5171);
xor XOR2 (N16906, N16898, N13519);
xor XOR2 (N16907, N16893, N5850);
or OR3 (N16908, N16900, N5741, N6693);
nor NOR2 (N16909, N16896, N3666);
and AND2 (N16910, N16897, N874);
buf BUF1 (N16911, N16904);
xor XOR2 (N16912, N16910, N3965);
buf BUF1 (N16913, N16912);
not NOT1 (N16914, N16906);
and AND4 (N16915, N16911, N11848, N285, N7944);
buf BUF1 (N16916, N16913);
and AND4 (N16917, N16909, N11405, N343, N3528);
and AND4 (N16918, N16903, N8102, N8687, N8120);
nor NOR3 (N16919, N16902, N6941, N1687);
nor NOR2 (N16920, N16905, N1410);
buf BUF1 (N16921, N16907);
nor NOR2 (N16922, N16919, N1656);
xor XOR2 (N16923, N16917, N1884);
xor XOR2 (N16924, N16918, N6038);
xor XOR2 (N16925, N16924, N7203);
xor XOR2 (N16926, N16916, N12704);
buf BUF1 (N16927, N16890);
nand NAND2 (N16928, N16925, N13075);
and AND3 (N16929, N16923, N8428, N9382);
and AND3 (N16930, N16926, N5506, N15765);
buf BUF1 (N16931, N16929);
buf BUF1 (N16932, N16915);
nand NAND2 (N16933, N16922, N2923);
and AND2 (N16934, N16931, N11117);
nand NAND4 (N16935, N16920, N9973, N9061, N2315);
xor XOR2 (N16936, N16928, N13677);
and AND2 (N16937, N16932, N6982);
xor XOR2 (N16938, N16930, N6198);
or OR4 (N16939, N16936, N6460, N2118, N12112);
or OR3 (N16940, N16935, N4190, N8903);
nand NAND4 (N16941, N16937, N7361, N8573, N11629);
or OR4 (N16942, N16938, N9816, N6804, N3882);
or OR3 (N16943, N16908, N14869, N7921);
or OR2 (N16944, N16927, N12133);
not NOT1 (N16945, N16914);
buf BUF1 (N16946, N16943);
nor NOR2 (N16947, N16933, N11828);
nand NAND3 (N16948, N16940, N11109, N653);
and AND4 (N16949, N16947, N13621, N10494, N6499);
buf BUF1 (N16950, N16941);
nor NOR3 (N16951, N16944, N12086, N1209);
buf BUF1 (N16952, N16949);
nor NOR2 (N16953, N16939, N15572);
xor XOR2 (N16954, N16951, N9132);
nor NOR3 (N16955, N16954, N3544, N15525);
xor XOR2 (N16956, N16945, N4769);
xor XOR2 (N16957, N16953, N12682);
and AND4 (N16958, N16957, N16390, N12925, N5029);
and AND2 (N16959, N16958, N4686);
or OR2 (N16960, N16934, N5839);
or OR3 (N16961, N16948, N7606, N6677);
and AND2 (N16962, N16921, N6158);
or OR2 (N16963, N16959, N4694);
xor XOR2 (N16964, N16962, N667);
not NOT1 (N16965, N16961);
and AND3 (N16966, N16955, N106, N16213);
and AND3 (N16967, N16965, N2318, N7180);
and AND2 (N16968, N16952, N12595);
buf BUF1 (N16969, N16942);
buf BUF1 (N16970, N16966);
xor XOR2 (N16971, N16956, N16325);
buf BUF1 (N16972, N16960);
not NOT1 (N16973, N16971);
nand NAND3 (N16974, N16969, N14399, N11918);
or OR3 (N16975, N16950, N594, N4306);
nand NAND2 (N16976, N16972, N1234);
xor XOR2 (N16977, N16970, N13262);
not NOT1 (N16978, N16975);
nand NAND4 (N16979, N16963, N187, N6782, N12591);
xor XOR2 (N16980, N16946, N13906);
nor NOR2 (N16981, N16973, N5522);
nor NOR3 (N16982, N16980, N12982, N11866);
not NOT1 (N16983, N16978);
or OR4 (N16984, N16979, N619, N3394, N3086);
not NOT1 (N16985, N16974);
or OR3 (N16986, N16967, N12106, N7947);
not NOT1 (N16987, N16976);
nor NOR4 (N16988, N16987, N16875, N11785, N16826);
or OR4 (N16989, N16968, N4461, N12949, N6085);
or OR2 (N16990, N16983, N13951);
xor XOR2 (N16991, N16964, N3818);
xor XOR2 (N16992, N16981, N16326);
nor NOR2 (N16993, N16984, N9067);
or OR4 (N16994, N16990, N4994, N636, N14317);
nand NAND4 (N16995, N16986, N13456, N8836, N11665);
not NOT1 (N16996, N16988);
and AND4 (N16997, N16991, N6478, N7550, N3295);
buf BUF1 (N16998, N16989);
xor XOR2 (N16999, N16998, N12309);
buf BUF1 (N17000, N16999);
buf BUF1 (N17001, N16995);
nand NAND4 (N17002, N16993, N4186, N15273, N9000);
or OR3 (N17003, N16992, N13266, N16090);
buf BUF1 (N17004, N17003);
xor XOR2 (N17005, N16982, N14631);
nand NAND2 (N17006, N17000, N15506);
nor NOR3 (N17007, N17006, N24, N1930);
or OR4 (N17008, N17004, N1436, N15360, N16113);
and AND2 (N17009, N17008, N9100);
and AND4 (N17010, N16997, N5664, N15709, N2266);
xor XOR2 (N17011, N16985, N8970);
nand NAND3 (N17012, N17010, N13176, N4357);
or OR4 (N17013, N17007, N7938, N16933, N7755);
nand NAND4 (N17014, N17012, N1349, N14385, N5510);
buf BUF1 (N17015, N16996);
nand NAND4 (N17016, N17013, N12220, N16708, N1335);
not NOT1 (N17017, N16977);
buf BUF1 (N17018, N17002);
or OR3 (N17019, N17014, N3571, N14364);
xor XOR2 (N17020, N17018, N9502);
nor NOR4 (N17021, N17016, N1314, N10496, N9433);
xor XOR2 (N17022, N17019, N13538);
buf BUF1 (N17023, N17021);
buf BUF1 (N17024, N17017);
or OR2 (N17025, N17024, N1228);
buf BUF1 (N17026, N16994);
nand NAND4 (N17027, N17020, N8481, N15538, N2442);
and AND3 (N17028, N17015, N14356, N1642);
not NOT1 (N17029, N17028);
nand NAND4 (N17030, N17027, N11620, N3072, N7964);
not NOT1 (N17031, N17022);
and AND4 (N17032, N17005, N122, N8612, N10586);
nor NOR3 (N17033, N17026, N10962, N3540);
nor NOR3 (N17034, N17033, N8360, N14771);
nor NOR2 (N17035, N17034, N6335);
buf BUF1 (N17036, N17030);
or OR3 (N17037, N17023, N2166, N6496);
not NOT1 (N17038, N17032);
nand NAND3 (N17039, N17025, N8900, N5894);
and AND2 (N17040, N17036, N1700);
not NOT1 (N17041, N17038);
buf BUF1 (N17042, N17040);
not NOT1 (N17043, N17031);
and AND4 (N17044, N17037, N3517, N541, N8742);
nor NOR3 (N17045, N17011, N16031, N14925);
and AND4 (N17046, N17042, N16596, N10954, N12171);
not NOT1 (N17047, N17009);
or OR2 (N17048, N17035, N6435);
buf BUF1 (N17049, N17045);
or OR2 (N17050, N17043, N15442);
xor XOR2 (N17051, N17048, N11097);
xor XOR2 (N17052, N17039, N8558);
nor NOR4 (N17053, N17050, N2149, N12217, N7315);
not NOT1 (N17054, N17029);
or OR2 (N17055, N17053, N705);
nand NAND3 (N17056, N17054, N15879, N10467);
not NOT1 (N17057, N17049);
nor NOR4 (N17058, N17056, N16490, N15291, N707);
nor NOR4 (N17059, N17052, N5121, N8215, N6894);
and AND3 (N17060, N17058, N16307, N4702);
not NOT1 (N17061, N17059);
buf BUF1 (N17062, N17047);
nand NAND3 (N17063, N17041, N1574, N15327);
xor XOR2 (N17064, N17001, N11599);
not NOT1 (N17065, N17062);
buf BUF1 (N17066, N17065);
nor NOR2 (N17067, N17044, N8914);
buf BUF1 (N17068, N17051);
or OR2 (N17069, N17067, N3357);
nor NOR2 (N17070, N17068, N11041);
xor XOR2 (N17071, N17061, N6517);
xor XOR2 (N17072, N17066, N13223);
and AND4 (N17073, N17064, N7024, N188, N2518);
buf BUF1 (N17074, N17060);
or OR2 (N17075, N17069, N4973);
and AND3 (N17076, N17075, N16201, N11414);
or OR2 (N17077, N17070, N9687);
xor XOR2 (N17078, N17057, N7305);
and AND3 (N17079, N17055, N1139, N5436);
buf BUF1 (N17080, N17078);
buf BUF1 (N17081, N17073);
and AND4 (N17082, N17080, N7422, N4707, N4373);
nor NOR4 (N17083, N17046, N6025, N13293, N429);
and AND3 (N17084, N17072, N5221, N1682);
or OR3 (N17085, N17071, N2457, N6612);
not NOT1 (N17086, N17084);
nand NAND3 (N17087, N17077, N14654, N13930);
nor NOR4 (N17088, N17087, N6610, N10146, N11846);
nand NAND3 (N17089, N17074, N366, N411);
or OR3 (N17090, N17088, N1850, N14267);
and AND4 (N17091, N17090, N11027, N11465, N7173);
nand NAND3 (N17092, N17082, N366, N16826);
or OR3 (N17093, N17091, N363, N4032);
nand NAND3 (N17094, N17079, N1766, N8869);
not NOT1 (N17095, N17063);
nor NOR4 (N17096, N17089, N1022, N9240, N14205);
or OR4 (N17097, N17096, N5261, N1786, N15979);
nor NOR4 (N17098, N17085, N4637, N14591, N9003);
or OR2 (N17099, N17083, N5852);
nor NOR3 (N17100, N17092, N16581, N11677);
and AND3 (N17101, N17093, N13096, N14763);
buf BUF1 (N17102, N17086);
nand NAND3 (N17103, N17098, N613, N9100);
nor NOR4 (N17104, N17076, N12478, N11450, N1968);
not NOT1 (N17105, N17097);
buf BUF1 (N17106, N17101);
buf BUF1 (N17107, N17105);
buf BUF1 (N17108, N17081);
nor NOR3 (N17109, N17099, N13002, N10826);
nor NOR4 (N17110, N17094, N2659, N287, N7853);
or OR3 (N17111, N17106, N2294, N2773);
and AND2 (N17112, N17108, N13282);
and AND2 (N17113, N17102, N11415);
nor NOR4 (N17114, N17104, N5828, N14776, N8716);
buf BUF1 (N17115, N17113);
or OR2 (N17116, N17100, N10221);
buf BUF1 (N17117, N17107);
nor NOR3 (N17118, N17111, N11353, N1571);
nor NOR2 (N17119, N17116, N16188);
or OR3 (N17120, N17112, N2688, N11270);
or OR4 (N17121, N17095, N12617, N1586, N7973);
nor NOR3 (N17122, N17109, N7936, N1394);
or OR3 (N17123, N17119, N12402, N11095);
xor XOR2 (N17124, N17117, N12072);
nand NAND3 (N17125, N17120, N2891, N879);
buf BUF1 (N17126, N17110);
and AND4 (N17127, N17126, N921, N15430, N13275);
xor XOR2 (N17128, N17114, N6252);
or OR3 (N17129, N17127, N6321, N12869);
and AND4 (N17130, N17122, N1646, N15337, N14170);
not NOT1 (N17131, N17128);
or OR2 (N17132, N17115, N13117);
xor XOR2 (N17133, N17103, N4903);
nor NOR2 (N17134, N17125, N1909);
xor XOR2 (N17135, N17124, N7835);
xor XOR2 (N17136, N17118, N9012);
and AND3 (N17137, N17132, N16212, N6842);
not NOT1 (N17138, N17131);
nand NAND3 (N17139, N17134, N8538, N823);
xor XOR2 (N17140, N17133, N10681);
nand NAND3 (N17141, N17135, N14128, N11097);
or OR4 (N17142, N17136, N6388, N8598, N5823);
not NOT1 (N17143, N17142);
nor NOR4 (N17144, N17138, N8845, N13384, N10045);
not NOT1 (N17145, N17139);
or OR2 (N17146, N17141, N4426);
xor XOR2 (N17147, N17145, N15941);
and AND2 (N17148, N17147, N12710);
not NOT1 (N17149, N17143);
not NOT1 (N17150, N17148);
or OR2 (N17151, N17149, N13884);
or OR3 (N17152, N17121, N15998, N7258);
or OR3 (N17153, N17140, N10998, N6411);
and AND2 (N17154, N17129, N7921);
buf BUF1 (N17155, N17152);
xor XOR2 (N17156, N17151, N8661);
nor NOR4 (N17157, N17155, N4519, N1247, N16006);
xor XOR2 (N17158, N17130, N760);
or OR3 (N17159, N17144, N8337, N1909);
nor NOR3 (N17160, N17137, N3125, N1417);
not NOT1 (N17161, N17157);
not NOT1 (N17162, N17150);
or OR2 (N17163, N17146, N14328);
nand NAND2 (N17164, N17123, N10362);
nand NAND3 (N17165, N17159, N4228, N14504);
nand NAND4 (N17166, N17160, N15291, N4340, N1953);
nand NAND3 (N17167, N17164, N12093, N7363);
not NOT1 (N17168, N17162);
or OR4 (N17169, N17153, N2235, N13170, N6957);
and AND3 (N17170, N17168, N9060, N12939);
nand NAND2 (N17171, N17154, N431);
or OR2 (N17172, N17163, N1873);
or OR4 (N17173, N17171, N15320, N13105, N13016);
not NOT1 (N17174, N17158);
nand NAND4 (N17175, N17156, N3277, N3114, N5276);
nor NOR4 (N17176, N17174, N10111, N9724, N4961);
buf BUF1 (N17177, N17173);
nand NAND3 (N17178, N17177, N3846, N16670);
buf BUF1 (N17179, N17167);
or OR4 (N17180, N17170, N6639, N5190, N11598);
or OR3 (N17181, N17175, N132, N13351);
nand NAND2 (N17182, N17165, N6801);
xor XOR2 (N17183, N17178, N760);
nand NAND4 (N17184, N17183, N16894, N5887, N9457);
buf BUF1 (N17185, N17172);
nor NOR3 (N17186, N17166, N14268, N15809);
and AND4 (N17187, N17186, N9091, N14264, N2413);
buf BUF1 (N17188, N17182);
xor XOR2 (N17189, N17181, N12566);
and AND3 (N17190, N17184, N4832, N5386);
nand NAND4 (N17191, N17190, N2790, N15803, N16844);
nand NAND4 (N17192, N17169, N13360, N7658, N16428);
buf BUF1 (N17193, N17161);
nand NAND4 (N17194, N17176, N3679, N7679, N13611);
buf BUF1 (N17195, N17180);
nand NAND4 (N17196, N17185, N13867, N2777, N10675);
not NOT1 (N17197, N17194);
not NOT1 (N17198, N17196);
buf BUF1 (N17199, N17197);
or OR3 (N17200, N17187, N13698, N14174);
nor NOR2 (N17201, N17192, N7040);
or OR2 (N17202, N17198, N1310);
not NOT1 (N17203, N17199);
or OR4 (N17204, N17188, N9586, N5436, N1459);
and AND2 (N17205, N17203, N3019);
buf BUF1 (N17206, N17195);
nor NOR4 (N17207, N17205, N13283, N1182, N6153);
nor NOR3 (N17208, N17200, N9448, N5244);
buf BUF1 (N17209, N17204);
not NOT1 (N17210, N17191);
not NOT1 (N17211, N17202);
or OR4 (N17212, N17207, N763, N14465, N11392);
and AND2 (N17213, N17201, N6502);
not NOT1 (N17214, N17211);
xor XOR2 (N17215, N17214, N2011);
xor XOR2 (N17216, N17210, N5529);
nand NAND2 (N17217, N17189, N5689);
xor XOR2 (N17218, N17215, N14950);
nor NOR3 (N17219, N17218, N15158, N8093);
buf BUF1 (N17220, N17208);
and AND3 (N17221, N17179, N14109, N5597);
xor XOR2 (N17222, N17217, N14850);
nand NAND3 (N17223, N17222, N14246, N12252);
xor XOR2 (N17224, N17216, N6387);
or OR2 (N17225, N17221, N12414);
buf BUF1 (N17226, N17212);
xor XOR2 (N17227, N17220, N12350);
nor NOR2 (N17228, N17225, N15242);
nor NOR2 (N17229, N17219, N1477);
nor NOR2 (N17230, N17193, N467);
xor XOR2 (N17231, N17223, N2862);
or OR3 (N17232, N17213, N6116, N5332);
nor NOR2 (N17233, N17229, N14716);
nor NOR2 (N17234, N17231, N5678);
and AND2 (N17235, N17226, N574);
nor NOR4 (N17236, N17209, N6370, N13423, N8876);
nand NAND4 (N17237, N17236, N1227, N13966, N11395);
not NOT1 (N17238, N17227);
buf BUF1 (N17239, N17233);
and AND4 (N17240, N17238, N13987, N13337, N10462);
xor XOR2 (N17241, N17232, N7395);
xor XOR2 (N17242, N17206, N1560);
and AND3 (N17243, N17241, N14065, N246);
nor NOR3 (N17244, N17228, N15990, N6749);
xor XOR2 (N17245, N17224, N10862);
nand NAND4 (N17246, N17237, N10402, N7664, N12762);
and AND4 (N17247, N17242, N6749, N16777, N14910);
xor XOR2 (N17248, N17247, N11906);
not NOT1 (N17249, N17246);
and AND3 (N17250, N17230, N3203, N14261);
xor XOR2 (N17251, N17240, N15083);
not NOT1 (N17252, N17248);
nor NOR4 (N17253, N17235, N14701, N13338, N14216);
not NOT1 (N17254, N17249);
nor NOR4 (N17255, N17239, N10134, N7473, N1648);
and AND3 (N17256, N17243, N2867, N9269);
nand NAND3 (N17257, N17250, N9549, N10654);
buf BUF1 (N17258, N17253);
and AND2 (N17259, N17244, N11312);
xor XOR2 (N17260, N17258, N3823);
nor NOR3 (N17261, N17251, N5335, N13716);
xor XOR2 (N17262, N17245, N15025);
or OR4 (N17263, N17261, N9043, N17249, N9160);
and AND2 (N17264, N17263, N9544);
buf BUF1 (N17265, N17254);
xor XOR2 (N17266, N17234, N16533);
not NOT1 (N17267, N17266);
not NOT1 (N17268, N17259);
or OR3 (N17269, N17256, N4326, N4065);
buf BUF1 (N17270, N17257);
or OR3 (N17271, N17268, N12169, N8860);
or OR4 (N17272, N17267, N915, N17069, N7910);
or OR4 (N17273, N17272, N11285, N15349, N1058);
not NOT1 (N17274, N17265);
buf BUF1 (N17275, N17271);
buf BUF1 (N17276, N17262);
nand NAND2 (N17277, N17252, N738);
not NOT1 (N17278, N17269);
not NOT1 (N17279, N17260);
not NOT1 (N17280, N17264);
nand NAND3 (N17281, N17278, N647, N9515);
nand NAND3 (N17282, N17275, N5852, N16387);
or OR3 (N17283, N17274, N8244, N15729);
nand NAND2 (N17284, N17255, N223);
buf BUF1 (N17285, N17273);
nor NOR2 (N17286, N17282, N1950);
or OR2 (N17287, N17279, N8744);
not NOT1 (N17288, N17283);
not NOT1 (N17289, N17285);
xor XOR2 (N17290, N17288, N2738);
not NOT1 (N17291, N17287);
xor XOR2 (N17292, N17286, N6904);
and AND2 (N17293, N17281, N1080);
not NOT1 (N17294, N17284);
xor XOR2 (N17295, N17290, N635);
buf BUF1 (N17296, N17289);
nand NAND2 (N17297, N17280, N3391);
or OR3 (N17298, N17276, N12380, N3374);
nor NOR4 (N17299, N17298, N8884, N501, N14230);
nand NAND4 (N17300, N17295, N14827, N5080, N11181);
buf BUF1 (N17301, N17297);
or OR4 (N17302, N17300, N14675, N12810, N7506);
or OR4 (N17303, N17291, N8068, N306, N14448);
not NOT1 (N17304, N17294);
nor NOR4 (N17305, N17301, N11249, N5768, N5516);
not NOT1 (N17306, N17299);
xor XOR2 (N17307, N17302, N13862);
or OR3 (N17308, N17292, N2244, N14973);
nand NAND4 (N17309, N17277, N3715, N8132, N7309);
and AND3 (N17310, N17309, N5230, N15107);
and AND4 (N17311, N17304, N522, N11558, N2261);
buf BUF1 (N17312, N17307);
or OR3 (N17313, N17270, N13290, N1461);
not NOT1 (N17314, N17310);
xor XOR2 (N17315, N17305, N12219);
buf BUF1 (N17316, N17314);
nand NAND3 (N17317, N17315, N14926, N5345);
not NOT1 (N17318, N17316);
not NOT1 (N17319, N17311);
not NOT1 (N17320, N17313);
nor NOR3 (N17321, N17317, N13863, N543);
not NOT1 (N17322, N17303);
buf BUF1 (N17323, N17306);
nand NAND3 (N17324, N17312, N15413, N6843);
buf BUF1 (N17325, N17319);
not NOT1 (N17326, N17321);
or OR4 (N17327, N17325, N10120, N4234, N481);
nand NAND3 (N17328, N17324, N3872, N9165);
or OR4 (N17329, N17322, N2565, N10665, N4365);
nand NAND2 (N17330, N17327, N10244);
xor XOR2 (N17331, N17330, N1261);
and AND3 (N17332, N17308, N5464, N2746);
and AND3 (N17333, N17293, N13918, N11779);
and AND3 (N17334, N17326, N1324, N1423);
not NOT1 (N17335, N17296);
buf BUF1 (N17336, N17318);
nand NAND2 (N17337, N17323, N3997);
not NOT1 (N17338, N17329);
or OR3 (N17339, N17337, N16186, N8965);
not NOT1 (N17340, N17339);
not NOT1 (N17341, N17334);
or OR2 (N17342, N17335, N4);
nand NAND2 (N17343, N17332, N14110);
not NOT1 (N17344, N17320);
not NOT1 (N17345, N17336);
and AND4 (N17346, N17328, N13389, N368, N7115);
not NOT1 (N17347, N17343);
not NOT1 (N17348, N17338);
nand NAND2 (N17349, N17347, N10456);
or OR2 (N17350, N17348, N1169);
buf BUF1 (N17351, N17345);
nor NOR3 (N17352, N17342, N13823, N3896);
nor NOR2 (N17353, N17331, N6741);
or OR3 (N17354, N17344, N1340, N12977);
and AND3 (N17355, N17349, N9737, N6897);
and AND4 (N17356, N17346, N3342, N13784, N5260);
xor XOR2 (N17357, N17350, N7422);
or OR3 (N17358, N17355, N14533, N3160);
or OR3 (N17359, N17341, N1482, N10757);
or OR2 (N17360, N17359, N17001);
xor XOR2 (N17361, N17353, N2657);
nand NAND2 (N17362, N17360, N1890);
buf BUF1 (N17363, N17357);
or OR4 (N17364, N17362, N3500, N6160, N6956);
buf BUF1 (N17365, N17354);
xor XOR2 (N17366, N17340, N4806);
nor NOR2 (N17367, N17363, N15036);
buf BUF1 (N17368, N17365);
nor NOR2 (N17369, N17358, N5249);
or OR3 (N17370, N17364, N1716, N2279);
buf BUF1 (N17371, N17351);
buf BUF1 (N17372, N17333);
buf BUF1 (N17373, N17370);
nand NAND4 (N17374, N17352, N14441, N695, N15294);
and AND2 (N17375, N17371, N3025);
and AND4 (N17376, N17368, N17238, N5697, N11992);
and AND4 (N17377, N17372, N8292, N7316, N1969);
nand NAND3 (N17378, N17377, N5309, N13321);
nand NAND4 (N17379, N17361, N16420, N15430, N1061);
not NOT1 (N17380, N17379);
not NOT1 (N17381, N17373);
nor NOR2 (N17382, N17380, N9116);
nand NAND2 (N17383, N17367, N13397);
buf BUF1 (N17384, N17356);
buf BUF1 (N17385, N17375);
buf BUF1 (N17386, N17381);
nand NAND4 (N17387, N17378, N67, N9065, N13974);
and AND2 (N17388, N17384, N8655);
xor XOR2 (N17389, N17374, N14148);
nand NAND3 (N17390, N17385, N10809, N8915);
buf BUF1 (N17391, N17386);
or OR4 (N17392, N17387, N718, N2959, N3468);
xor XOR2 (N17393, N17383, N12253);
nand NAND2 (N17394, N17392, N4481);
nor NOR3 (N17395, N17376, N10153, N15045);
and AND3 (N17396, N17391, N11822, N15830);
and AND2 (N17397, N17390, N14260);
nor NOR4 (N17398, N17388, N7119, N15854, N12361);
nand NAND2 (N17399, N17393, N6434);
xor XOR2 (N17400, N17389, N15510);
xor XOR2 (N17401, N17382, N11269);
nand NAND3 (N17402, N17399, N13433, N6336);
or OR3 (N17403, N17396, N2003, N12335);
buf BUF1 (N17404, N17395);
xor XOR2 (N17405, N17397, N7901);
xor XOR2 (N17406, N17403, N7504);
not NOT1 (N17407, N17398);
xor XOR2 (N17408, N17369, N7362);
xor XOR2 (N17409, N17406, N2653);
buf BUF1 (N17410, N17402);
buf BUF1 (N17411, N17394);
or OR2 (N17412, N17411, N5720);
xor XOR2 (N17413, N17400, N547);
not NOT1 (N17414, N17408);
buf BUF1 (N17415, N17404);
and AND2 (N17416, N17415, N6937);
and AND2 (N17417, N17407, N2692);
xor XOR2 (N17418, N17412, N6597);
nor NOR3 (N17419, N17401, N2723, N15894);
or OR4 (N17420, N17419, N3970, N6100, N15404);
nand NAND2 (N17421, N17410, N9107);
and AND3 (N17422, N17417, N6433, N8854);
nor NOR2 (N17423, N17418, N13473);
nor NOR2 (N17424, N17409, N16810);
nor NOR4 (N17425, N17422, N3824, N4315, N16965);
nand NAND2 (N17426, N17366, N9257);
xor XOR2 (N17427, N17405, N1885);
xor XOR2 (N17428, N17427, N6421);
nand NAND3 (N17429, N17414, N1777, N10707);
and AND3 (N17430, N17416, N17082, N6582);
nor NOR2 (N17431, N17425, N7937);
xor XOR2 (N17432, N17426, N12150);
or OR3 (N17433, N17421, N15574, N6727);
or OR2 (N17434, N17429, N2371);
nor NOR3 (N17435, N17428, N5425, N12016);
buf BUF1 (N17436, N17432);
nand NAND4 (N17437, N17434, N10950, N14475, N7314);
not NOT1 (N17438, N17433);
and AND4 (N17439, N17424, N5668, N16446, N13939);
nand NAND4 (N17440, N17437, N15259, N9487, N6196);
xor XOR2 (N17441, N17439, N16092);
not NOT1 (N17442, N17420);
and AND3 (N17443, N17440, N5212, N3457);
nor NOR2 (N17444, N17442, N2866);
not NOT1 (N17445, N17441);
nand NAND2 (N17446, N17438, N7857);
xor XOR2 (N17447, N17423, N10261);
not NOT1 (N17448, N17447);
not NOT1 (N17449, N17430);
nor NOR4 (N17450, N17446, N1657, N15545, N14686);
xor XOR2 (N17451, N17449, N2530);
xor XOR2 (N17452, N17448, N10782);
or OR2 (N17453, N17452, N2458);
xor XOR2 (N17454, N17436, N7365);
nand NAND3 (N17455, N17431, N3869, N9892);
buf BUF1 (N17456, N17454);
nor NOR4 (N17457, N17453, N1039, N2718, N9146);
not NOT1 (N17458, N17456);
xor XOR2 (N17459, N17435, N629);
xor XOR2 (N17460, N17451, N1515);
buf BUF1 (N17461, N17443);
not NOT1 (N17462, N17461);
nor NOR4 (N17463, N17460, N9413, N3670, N14945);
nand NAND4 (N17464, N17413, N3503, N16168, N9722);
nor NOR4 (N17465, N17462, N2100, N9508, N11139);
nor NOR2 (N17466, N17444, N9442);
and AND4 (N17467, N17455, N11268, N14020, N2529);
not NOT1 (N17468, N17445);
or OR3 (N17469, N17459, N8626, N9615);
xor XOR2 (N17470, N17468, N11178);
and AND2 (N17471, N17469, N14850);
buf BUF1 (N17472, N17465);
buf BUF1 (N17473, N17467);
nand NAND3 (N17474, N17450, N9059, N14857);
not NOT1 (N17475, N17474);
and AND2 (N17476, N17463, N7858);
not NOT1 (N17477, N17471);
buf BUF1 (N17478, N17466);
or OR2 (N17479, N17457, N13650);
and AND2 (N17480, N17464, N15723);
nand NAND4 (N17481, N17480, N9609, N333, N3526);
buf BUF1 (N17482, N17477);
or OR4 (N17483, N17478, N15683, N16605, N8893);
nor NOR2 (N17484, N17470, N3085);
nor NOR3 (N17485, N17476, N1617, N14939);
or OR4 (N17486, N17472, N16318, N558, N14566);
xor XOR2 (N17487, N17473, N13668);
not NOT1 (N17488, N17486);
buf BUF1 (N17489, N17475);
or OR2 (N17490, N17484, N5810);
and AND2 (N17491, N17485, N7718);
not NOT1 (N17492, N17488);
buf BUF1 (N17493, N17492);
not NOT1 (N17494, N17482);
buf BUF1 (N17495, N17481);
nor NOR3 (N17496, N17495, N1358, N6146);
and AND3 (N17497, N17491, N11139, N17401);
buf BUF1 (N17498, N17487);
nand NAND4 (N17499, N17493, N4630, N14250, N6116);
nand NAND2 (N17500, N17479, N13401);
not NOT1 (N17501, N17498);
and AND2 (N17502, N17458, N3165);
xor XOR2 (N17503, N17497, N8807);
nor NOR4 (N17504, N17494, N14843, N8162, N3107);
nor NOR3 (N17505, N17489, N4067, N14695);
buf BUF1 (N17506, N17483);
not NOT1 (N17507, N17502);
buf BUF1 (N17508, N17501);
not NOT1 (N17509, N17505);
buf BUF1 (N17510, N17503);
nor NOR2 (N17511, N17509, N3889);
or OR2 (N17512, N17510, N13748);
or OR2 (N17513, N17499, N9708);
or OR2 (N17514, N17508, N9607);
and AND4 (N17515, N17512, N6534, N8568, N15984);
and AND2 (N17516, N17504, N8952);
nor NOR3 (N17517, N17513, N4373, N8116);
xor XOR2 (N17518, N17490, N3505);
buf BUF1 (N17519, N17516);
buf BUF1 (N17520, N17511);
and AND3 (N17521, N17518, N17504, N8543);
not NOT1 (N17522, N17506);
buf BUF1 (N17523, N17521);
not NOT1 (N17524, N17500);
xor XOR2 (N17525, N17522, N1412);
buf BUF1 (N17526, N17524);
nand NAND2 (N17527, N17519, N14652);
buf BUF1 (N17528, N17527);
buf BUF1 (N17529, N17526);
buf BUF1 (N17530, N17529);
nand NAND2 (N17531, N17517, N2954);
nand NAND3 (N17532, N17523, N14220, N1784);
and AND4 (N17533, N17520, N17130, N8368, N6623);
and AND4 (N17534, N17525, N5837, N15154, N9150);
or OR4 (N17535, N17530, N263, N14677, N3847);
or OR3 (N17536, N17535, N7820, N12204);
buf BUF1 (N17537, N17536);
or OR4 (N17538, N17533, N14038, N5417, N12267);
xor XOR2 (N17539, N17531, N14031);
and AND4 (N17540, N17538, N4434, N9521, N8241);
nor NOR3 (N17541, N17507, N2556, N15243);
nor NOR4 (N17542, N17528, N13867, N2074, N17310);
and AND2 (N17543, N17496, N12654);
xor XOR2 (N17544, N17542, N8029);
nor NOR3 (N17545, N17515, N7744, N4980);
xor XOR2 (N17546, N17514, N7500);
nand NAND3 (N17547, N17545, N10206, N11248);
not NOT1 (N17548, N17544);
xor XOR2 (N17549, N17543, N7033);
and AND3 (N17550, N17539, N12126, N10557);
buf BUF1 (N17551, N17549);
xor XOR2 (N17552, N17547, N1620);
or OR4 (N17553, N17534, N7729, N10731, N1831);
and AND4 (N17554, N17540, N7132, N8367, N13973);
and AND3 (N17555, N17552, N6480, N12007);
and AND2 (N17556, N17537, N15272);
xor XOR2 (N17557, N17546, N10721);
nand NAND4 (N17558, N17557, N17431, N16200, N7656);
or OR2 (N17559, N17532, N4457);
nor NOR4 (N17560, N17550, N8794, N9594, N16274);
and AND4 (N17561, N17559, N9504, N12211, N15331);
or OR2 (N17562, N17556, N626);
and AND4 (N17563, N17560, N2224, N14594, N2200);
not NOT1 (N17564, N17555);
and AND4 (N17565, N17548, N2036, N6635, N94);
not NOT1 (N17566, N17562);
not NOT1 (N17567, N17564);
buf BUF1 (N17568, N17551);
buf BUF1 (N17569, N17558);
or OR3 (N17570, N17561, N1199, N8680);
not NOT1 (N17571, N17541);
not NOT1 (N17572, N17566);
buf BUF1 (N17573, N17567);
not NOT1 (N17574, N17571);
and AND2 (N17575, N17570, N1593);
buf BUF1 (N17576, N17563);
nand NAND3 (N17577, N17569, N10930, N17557);
and AND2 (N17578, N17575, N7740);
nor NOR3 (N17579, N17553, N6301, N10575);
or OR4 (N17580, N17579, N14282, N15823, N3742);
xor XOR2 (N17581, N17577, N14267);
nor NOR2 (N17582, N17572, N632);
not NOT1 (N17583, N17573);
nand NAND3 (N17584, N17580, N15971, N17387);
buf BUF1 (N17585, N17581);
or OR2 (N17586, N17554, N6543);
xor XOR2 (N17587, N17568, N7546);
nor NOR3 (N17588, N17584, N7277, N6072);
not NOT1 (N17589, N17583);
and AND3 (N17590, N17574, N11862, N5049);
or OR2 (N17591, N17578, N17036);
not NOT1 (N17592, N17565);
not NOT1 (N17593, N17576);
and AND4 (N17594, N17589, N14111, N11118, N7069);
or OR3 (N17595, N17591, N11401, N12062);
xor XOR2 (N17596, N17593, N15223);
nand NAND2 (N17597, N17586, N15768);
xor XOR2 (N17598, N17597, N13644);
or OR2 (N17599, N17598, N3618);
not NOT1 (N17600, N17596);
nand NAND2 (N17601, N17588, N10029);
or OR4 (N17602, N17585, N2315, N6442, N4727);
or OR2 (N17603, N17595, N700);
not NOT1 (N17604, N17592);
buf BUF1 (N17605, N17594);
xor XOR2 (N17606, N17601, N6531);
nor NOR3 (N17607, N17599, N10523, N10725);
xor XOR2 (N17608, N17603, N14102);
nor NOR4 (N17609, N17587, N9247, N11199, N7201);
nor NOR2 (N17610, N17607, N10197);
and AND4 (N17611, N17582, N16600, N4038, N10583);
or OR4 (N17612, N17606, N10647, N16252, N2516);
xor XOR2 (N17613, N17600, N9461);
and AND3 (N17614, N17611, N12790, N11007);
or OR2 (N17615, N17604, N7652);
or OR4 (N17616, N17609, N14936, N5243, N13467);
nor NOR2 (N17617, N17613, N15993);
not NOT1 (N17618, N17610);
nor NOR4 (N17619, N17612, N17233, N7932, N6286);
buf BUF1 (N17620, N17616);
not NOT1 (N17621, N17620);
xor XOR2 (N17622, N17590, N174);
and AND4 (N17623, N17608, N3550, N15402, N4319);
and AND4 (N17624, N17602, N5734, N8462, N10386);
xor XOR2 (N17625, N17605, N10369);
buf BUF1 (N17626, N17621);
buf BUF1 (N17627, N17622);
or OR2 (N17628, N17618, N16492);
nand NAND4 (N17629, N17623, N763, N8973, N14168);
xor XOR2 (N17630, N17625, N12288);
or OR3 (N17631, N17624, N4165, N14698);
xor XOR2 (N17632, N17615, N2898);
and AND3 (N17633, N17614, N17367, N16010);
buf BUF1 (N17634, N17626);
not NOT1 (N17635, N17630);
or OR3 (N17636, N17635, N4097, N14608);
xor XOR2 (N17637, N17628, N5343);
not NOT1 (N17638, N17633);
buf BUF1 (N17639, N17638);
xor XOR2 (N17640, N17636, N4073);
nand NAND4 (N17641, N17640, N4283, N17156, N12756);
nand NAND3 (N17642, N17632, N10356, N2873);
nor NOR4 (N17643, N17641, N3383, N1348, N14013);
nand NAND4 (N17644, N17639, N146, N6109, N11916);
or OR2 (N17645, N17644, N516);
xor XOR2 (N17646, N17619, N11943);
or OR3 (N17647, N17646, N3091, N14970);
xor XOR2 (N17648, N17642, N7499);
buf BUF1 (N17649, N17645);
buf BUF1 (N17650, N17637);
buf BUF1 (N17651, N17643);
xor XOR2 (N17652, N17650, N2681);
or OR3 (N17653, N17647, N12590, N5840);
or OR2 (N17654, N17631, N1667);
and AND3 (N17655, N17627, N7712, N9862);
or OR4 (N17656, N17649, N5014, N1652, N9932);
not NOT1 (N17657, N17656);
nor NOR4 (N17658, N17657, N11537, N14512, N7977);
and AND2 (N17659, N17655, N15670);
not NOT1 (N17660, N17652);
not NOT1 (N17661, N17648);
nor NOR3 (N17662, N17659, N228, N2641);
buf BUF1 (N17663, N17634);
not NOT1 (N17664, N17662);
or OR3 (N17665, N17663, N10348, N6943);
or OR3 (N17666, N17664, N6201, N9343);
buf BUF1 (N17667, N17658);
and AND2 (N17668, N17667, N16912);
and AND2 (N17669, N17654, N17297);
nor NOR4 (N17670, N17665, N3657, N16122, N15244);
or OR4 (N17671, N17666, N6163, N17499, N4389);
not NOT1 (N17672, N17669);
buf BUF1 (N17673, N17653);
or OR2 (N17674, N17617, N13288);
and AND4 (N17675, N17651, N8639, N3544, N6655);
xor XOR2 (N17676, N17671, N16739);
nor NOR2 (N17677, N17673, N15512);
buf BUF1 (N17678, N17676);
nand NAND4 (N17679, N17674, N14681, N8921, N1426);
and AND3 (N17680, N17679, N7599, N2758);
nor NOR4 (N17681, N17670, N13565, N15891, N8543);
xor XOR2 (N17682, N17661, N837);
or OR2 (N17683, N17672, N13565);
nor NOR3 (N17684, N17629, N6929, N5544);
and AND2 (N17685, N17668, N16332);
not NOT1 (N17686, N17681);
buf BUF1 (N17687, N17678);
and AND2 (N17688, N17680, N17617);
or OR2 (N17689, N17686, N16503);
xor XOR2 (N17690, N17682, N8537);
or OR2 (N17691, N17689, N2728);
xor XOR2 (N17692, N17685, N2403);
and AND4 (N17693, N17683, N9940, N3861, N10410);
not NOT1 (N17694, N17693);
not NOT1 (N17695, N17660);
nor NOR3 (N17696, N17692, N13724, N2876);
nor NOR3 (N17697, N17675, N8255, N13701);
nand NAND4 (N17698, N17690, N12624, N10143, N69);
or OR4 (N17699, N17695, N12258, N4892, N10591);
and AND2 (N17700, N17688, N2607);
nand NAND2 (N17701, N17691, N2545);
xor XOR2 (N17702, N17684, N16690);
not NOT1 (N17703, N17699);
not NOT1 (N17704, N17698);
and AND2 (N17705, N17696, N13041);
and AND4 (N17706, N17697, N8787, N9515, N7340);
or OR2 (N17707, N17706, N1017);
and AND2 (N17708, N17687, N15561);
and AND2 (N17709, N17694, N12481);
not NOT1 (N17710, N17704);
or OR3 (N17711, N17703, N7787, N13628);
and AND3 (N17712, N17677, N10721, N11642);
nand NAND2 (N17713, N17711, N13262);
or OR3 (N17714, N17701, N10435, N14919);
and AND2 (N17715, N17705, N16097);
not NOT1 (N17716, N17715);
nand NAND4 (N17717, N17716, N11516, N10662, N17226);
and AND3 (N17718, N17707, N16554, N7308);
buf BUF1 (N17719, N17712);
not NOT1 (N17720, N17714);
buf BUF1 (N17721, N17709);
not NOT1 (N17722, N17708);
nor NOR3 (N17723, N17720, N13520, N5449);
nand NAND2 (N17724, N17721, N15231);
not NOT1 (N17725, N17722);
xor XOR2 (N17726, N17702, N4334);
nand NAND2 (N17727, N17724, N10087);
buf BUF1 (N17728, N17719);
buf BUF1 (N17729, N17723);
not NOT1 (N17730, N17729);
not NOT1 (N17731, N17727);
not NOT1 (N17732, N17700);
and AND4 (N17733, N17732, N14320, N5302, N17023);
and AND2 (N17734, N17725, N6547);
not NOT1 (N17735, N17710);
nand NAND2 (N17736, N17731, N9018);
not NOT1 (N17737, N17730);
nor NOR2 (N17738, N17717, N1544);
nor NOR3 (N17739, N17728, N4514, N8181);
buf BUF1 (N17740, N17726);
not NOT1 (N17741, N17735);
xor XOR2 (N17742, N17739, N12736);
nor NOR4 (N17743, N17742, N12210, N5050, N13021);
not NOT1 (N17744, N17737);
and AND3 (N17745, N17740, N16288, N15851);
nand NAND2 (N17746, N17736, N14846);
not NOT1 (N17747, N17744);
nand NAND2 (N17748, N17745, N14714);
buf BUF1 (N17749, N17743);
buf BUF1 (N17750, N17734);
nand NAND4 (N17751, N17738, N10534, N3776, N14715);
or OR3 (N17752, N17748, N9120, N10306);
nand NAND4 (N17753, N17733, N3937, N443, N14560);
not NOT1 (N17754, N17751);
xor XOR2 (N17755, N17753, N15657);
nand NAND3 (N17756, N17754, N4053, N2252);
buf BUF1 (N17757, N17756);
not NOT1 (N17758, N17741);
nand NAND4 (N17759, N17750, N13140, N5843, N8181);
xor XOR2 (N17760, N17747, N1133);
not NOT1 (N17761, N17759);
and AND4 (N17762, N17752, N1798, N2357, N11579);
xor XOR2 (N17763, N17757, N6571);
or OR3 (N17764, N17749, N6930, N12111);
xor XOR2 (N17765, N17755, N8485);
nand NAND3 (N17766, N17763, N16334, N17445);
nor NOR2 (N17767, N17762, N11514);
nor NOR4 (N17768, N17760, N4969, N8501, N5592);
nor NOR2 (N17769, N17718, N757);
or OR4 (N17770, N17761, N9323, N2220, N7858);
nor NOR4 (N17771, N17770, N14561, N12334, N3565);
not NOT1 (N17772, N17746);
nor NOR2 (N17773, N17765, N14135);
xor XOR2 (N17774, N17758, N13175);
xor XOR2 (N17775, N17773, N11032);
and AND3 (N17776, N17713, N2848, N375);
and AND2 (N17777, N17768, N1774);
buf BUF1 (N17778, N17776);
or OR4 (N17779, N17769, N16700, N8201, N17263);
nand NAND4 (N17780, N17775, N7917, N15992, N11635);
and AND3 (N17781, N17767, N1995, N9544);
nor NOR3 (N17782, N17778, N375, N11101);
buf BUF1 (N17783, N17779);
nor NOR4 (N17784, N17777, N4412, N16851, N1228);
and AND3 (N17785, N17780, N16515, N15272);
buf BUF1 (N17786, N17764);
nor NOR2 (N17787, N17766, N16675);
buf BUF1 (N17788, N17785);
or OR4 (N17789, N17786, N5025, N8574, N8832);
xor XOR2 (N17790, N17772, N16982);
nor NOR2 (N17791, N17789, N3381);
or OR2 (N17792, N17787, N3612);
xor XOR2 (N17793, N17771, N16001);
nor NOR4 (N17794, N17782, N11259, N16886, N7141);
and AND3 (N17795, N17794, N3142, N7623);
nor NOR3 (N17796, N17783, N3867, N14246);
and AND4 (N17797, N17784, N6686, N11736, N13595);
nand NAND2 (N17798, N17792, N6304);
nand NAND2 (N17799, N17798, N5560);
and AND2 (N17800, N17788, N12127);
buf BUF1 (N17801, N17797);
buf BUF1 (N17802, N17774);
not NOT1 (N17803, N17790);
buf BUF1 (N17804, N17793);
or OR3 (N17805, N17799, N13929, N1559);
and AND3 (N17806, N17791, N1654, N4555);
xor XOR2 (N17807, N17800, N2402);
buf BUF1 (N17808, N17795);
nand NAND4 (N17809, N17806, N17667, N16512, N4201);
xor XOR2 (N17810, N17781, N11120);
and AND4 (N17811, N17805, N5684, N8658, N5103);
and AND4 (N17812, N17807, N13347, N1107, N5845);
nand NAND2 (N17813, N17804, N57);
nor NOR3 (N17814, N17808, N16991, N11580);
or OR3 (N17815, N17809, N4429, N7169);
xor XOR2 (N17816, N17803, N16280);
or OR2 (N17817, N17802, N14099);
not NOT1 (N17818, N17816);
xor XOR2 (N17819, N17817, N5066);
nand NAND4 (N17820, N17801, N11548, N8944, N10653);
nand NAND3 (N17821, N17810, N13999, N3123);
xor XOR2 (N17822, N17815, N6964);
or OR4 (N17823, N17822, N16357, N14564, N15184);
buf BUF1 (N17824, N17814);
xor XOR2 (N17825, N17820, N7627);
not NOT1 (N17826, N17812);
and AND3 (N17827, N17826, N11338, N1060);
nand NAND4 (N17828, N17823, N13552, N12642, N17415);
buf BUF1 (N17829, N17811);
not NOT1 (N17830, N17821);
nor NOR4 (N17831, N17828, N10540, N13217, N7690);
buf BUF1 (N17832, N17818);
or OR4 (N17833, N17829, N16300, N7593, N9566);
and AND3 (N17834, N17813, N6610, N15926);
or OR4 (N17835, N17796, N301, N4291, N12905);
and AND2 (N17836, N17827, N5273);
xor XOR2 (N17837, N17835, N1331);
xor XOR2 (N17838, N17833, N9933);
nand NAND2 (N17839, N17838, N7423);
and AND3 (N17840, N17832, N14965, N3660);
xor XOR2 (N17841, N17840, N10813);
buf BUF1 (N17842, N17841);
nor NOR4 (N17843, N17824, N324, N2109, N6799);
xor XOR2 (N17844, N17839, N4348);
and AND3 (N17845, N17837, N8952, N8670);
buf BUF1 (N17846, N17825);
and AND3 (N17847, N17831, N8580, N12874);
not NOT1 (N17848, N17834);
or OR2 (N17849, N17836, N5032);
and AND4 (N17850, N17843, N7277, N7809, N9986);
nor NOR2 (N17851, N17846, N16827);
or OR2 (N17852, N17849, N12513);
or OR3 (N17853, N17850, N2942, N5347);
or OR4 (N17854, N17852, N10729, N9226, N17433);
xor XOR2 (N17855, N17845, N14569);
or OR4 (N17856, N17854, N11137, N11039, N844);
xor XOR2 (N17857, N17847, N8735);
or OR2 (N17858, N17857, N7353);
buf BUF1 (N17859, N17819);
nor NOR4 (N17860, N17856, N13709, N8379, N2598);
nand NAND4 (N17861, N17853, N7774, N1328, N13463);
buf BUF1 (N17862, N17844);
nand NAND3 (N17863, N17862, N4150, N8455);
and AND2 (N17864, N17859, N3424);
and AND2 (N17865, N17830, N9625);
xor XOR2 (N17866, N17864, N9090);
nor NOR4 (N17867, N17848, N9676, N5415, N8223);
and AND3 (N17868, N17858, N16290, N14057);
and AND2 (N17869, N17851, N16319);
buf BUF1 (N17870, N17842);
or OR3 (N17871, N17867, N673, N14787);
xor XOR2 (N17872, N17855, N10228);
nor NOR2 (N17873, N17866, N7951);
buf BUF1 (N17874, N17873);
buf BUF1 (N17875, N17860);
nor NOR3 (N17876, N17863, N3400, N13915);
or OR4 (N17877, N17872, N1744, N16164, N10444);
nor NOR2 (N17878, N17861, N9576);
nand NAND2 (N17879, N17870, N10670);
buf BUF1 (N17880, N17868);
xor XOR2 (N17881, N17875, N1970);
not NOT1 (N17882, N17874);
not NOT1 (N17883, N17879);
and AND4 (N17884, N17877, N10226, N3507, N4294);
not NOT1 (N17885, N17881);
and AND3 (N17886, N17884, N10744, N14882);
not NOT1 (N17887, N17869);
not NOT1 (N17888, N17885);
nor NOR4 (N17889, N17883, N4160, N7808, N8073);
and AND2 (N17890, N17882, N16713);
and AND3 (N17891, N17878, N6191, N12780);
not NOT1 (N17892, N17890);
and AND2 (N17893, N17887, N4851);
not NOT1 (N17894, N17893);
not NOT1 (N17895, N17876);
nor NOR4 (N17896, N17894, N10061, N8179, N16533);
xor XOR2 (N17897, N17889, N3953);
not NOT1 (N17898, N17886);
buf BUF1 (N17899, N17888);
buf BUF1 (N17900, N17880);
xor XOR2 (N17901, N17895, N2191);
xor XOR2 (N17902, N17897, N2459);
nand NAND2 (N17903, N17901, N5554);
nor NOR4 (N17904, N17899, N1558, N10552, N11326);
not NOT1 (N17905, N17871);
and AND4 (N17906, N17892, N10897, N6771, N8656);
buf BUF1 (N17907, N17902);
and AND3 (N17908, N17903, N15370, N891);
nand NAND2 (N17909, N17865, N8418);
not NOT1 (N17910, N17904);
buf BUF1 (N17911, N17891);
and AND3 (N17912, N17908, N15648, N8942);
buf BUF1 (N17913, N17905);
not NOT1 (N17914, N17906);
nand NAND2 (N17915, N17909, N2089);
xor XOR2 (N17916, N17896, N15604);
and AND4 (N17917, N17913, N7395, N9309, N15506);
buf BUF1 (N17918, N17898);
and AND4 (N17919, N17912, N4733, N15183, N10055);
nand NAND2 (N17920, N17914, N918);
buf BUF1 (N17921, N17916);
nor NOR2 (N17922, N17911, N14083);
and AND3 (N17923, N17900, N864, N12499);
buf BUF1 (N17924, N17910);
not NOT1 (N17925, N17918);
not NOT1 (N17926, N17917);
or OR3 (N17927, N17922, N12405, N4851);
buf BUF1 (N17928, N17925);
or OR4 (N17929, N17923, N17604, N11065, N13777);
nor NOR3 (N17930, N17926, N17339, N9799);
and AND2 (N17931, N17920, N3410);
not NOT1 (N17932, N17924);
not NOT1 (N17933, N17927);
buf BUF1 (N17934, N17932);
not NOT1 (N17935, N17933);
xor XOR2 (N17936, N17928, N13073);
xor XOR2 (N17937, N17929, N5670);
or OR2 (N17938, N17915, N11291);
nand NAND4 (N17939, N17938, N5240, N10562, N5683);
not NOT1 (N17940, N17937);
buf BUF1 (N17941, N17940);
nand NAND2 (N17942, N17930, N6866);
nand NAND3 (N17943, N17934, N1046, N9568);
nor NOR2 (N17944, N17942, N1334);
nor NOR2 (N17945, N17936, N4431);
nor NOR4 (N17946, N17944, N4678, N2812, N11557);
buf BUF1 (N17947, N17919);
and AND3 (N17948, N17947, N5229, N3351);
not NOT1 (N17949, N17948);
not NOT1 (N17950, N17935);
xor XOR2 (N17951, N17950, N11903);
xor XOR2 (N17952, N17949, N14217);
buf BUF1 (N17953, N17951);
or OR2 (N17954, N17931, N5731);
not NOT1 (N17955, N17946);
not NOT1 (N17956, N17955);
and AND3 (N17957, N17953, N1975, N5787);
xor XOR2 (N17958, N17952, N13796);
not NOT1 (N17959, N17921);
nand NAND3 (N17960, N17907, N14206, N220);
buf BUF1 (N17961, N17958);
xor XOR2 (N17962, N17943, N7927);
nand NAND4 (N17963, N17960, N4642, N10891, N732);
not NOT1 (N17964, N17945);
and AND2 (N17965, N17939, N9337);
buf BUF1 (N17966, N17956);
and AND2 (N17967, N17941, N15974);
not NOT1 (N17968, N17957);
and AND3 (N17969, N17959, N10220, N1526);
xor XOR2 (N17970, N17965, N884);
and AND4 (N17971, N17967, N5182, N12347, N6078);
and AND3 (N17972, N17969, N61, N5192);
buf BUF1 (N17973, N17972);
buf BUF1 (N17974, N17961);
or OR4 (N17975, N17974, N13676, N547, N1860);
nor NOR2 (N17976, N17966, N13456);
not NOT1 (N17977, N17976);
and AND4 (N17978, N17962, N7129, N7645, N3878);
nor NOR4 (N17979, N17977, N11043, N11488, N14688);
not NOT1 (N17980, N17970);
buf BUF1 (N17981, N17978);
not NOT1 (N17982, N17975);
and AND3 (N17983, N17971, N1386, N12351);
xor XOR2 (N17984, N17954, N1520);
not NOT1 (N17985, N17963);
nor NOR4 (N17986, N17981, N13805, N7752, N12376);
nor NOR4 (N17987, N17986, N5947, N10130, N1601);
or OR2 (N17988, N17973, N17210);
xor XOR2 (N17989, N17979, N6035);
nor NOR2 (N17990, N17987, N5986);
not NOT1 (N17991, N17964);
nand NAND3 (N17992, N17985, N1540, N1860);
nand NAND4 (N17993, N17984, N10275, N15216, N2569);
buf BUF1 (N17994, N17990);
and AND2 (N17995, N17980, N13891);
or OR3 (N17996, N17993, N14128, N15265);
and AND4 (N17997, N17968, N4725, N15054, N9640);
nor NOR2 (N17998, N17995, N10852);
or OR2 (N17999, N17982, N10819);
buf BUF1 (N18000, N17997);
nand NAND4 (N18001, N17988, N3705, N6185, N5501);
not NOT1 (N18002, N17991);
or OR4 (N18003, N17994, N6891, N5195, N9118);
not NOT1 (N18004, N18000);
or OR2 (N18005, N17983, N17790);
xor XOR2 (N18006, N17989, N14993);
or OR2 (N18007, N18004, N14714);
xor XOR2 (N18008, N17999, N8171);
not NOT1 (N18009, N18005);
or OR4 (N18010, N17998, N17264, N12059, N8469);
xor XOR2 (N18011, N18008, N12322);
nand NAND2 (N18012, N18010, N13869);
nor NOR4 (N18013, N18002, N13, N9140, N9374);
buf BUF1 (N18014, N18009);
nor NOR4 (N18015, N18001, N17002, N11115, N10598);
buf BUF1 (N18016, N17992);
and AND3 (N18017, N18016, N1775, N5216);
nor NOR3 (N18018, N18014, N8192, N11508);
buf BUF1 (N18019, N18003);
nor NOR2 (N18020, N18007, N5510);
buf BUF1 (N18021, N18006);
not NOT1 (N18022, N17996);
nor NOR3 (N18023, N18019, N1995, N17371);
and AND2 (N18024, N18015, N7105);
nand NAND3 (N18025, N18024, N11797, N2403);
xor XOR2 (N18026, N18012, N14851);
buf BUF1 (N18027, N18025);
or OR4 (N18028, N18021, N10911, N14632, N10387);
or OR4 (N18029, N18022, N6200, N7407, N1936);
buf BUF1 (N18030, N18011);
xor XOR2 (N18031, N18020, N3975);
nor NOR4 (N18032, N18013, N7512, N8652, N10021);
nand NAND4 (N18033, N18032, N17666, N150, N11731);
and AND2 (N18034, N18029, N12526);
and AND2 (N18035, N18031, N8495);
and AND4 (N18036, N18018, N14928, N645, N9523);
and AND4 (N18037, N18027, N15365, N17517, N1793);
and AND4 (N18038, N18028, N6180, N13663, N15292);
and AND2 (N18039, N18030, N863);
buf BUF1 (N18040, N18035);
not NOT1 (N18041, N18017);
nand NAND3 (N18042, N18026, N18038, N4402);
or OR3 (N18043, N10848, N5854, N9218);
xor XOR2 (N18044, N18043, N920);
or OR4 (N18045, N18039, N3803, N10221, N11276);
buf BUF1 (N18046, N18037);
not NOT1 (N18047, N18034);
xor XOR2 (N18048, N18036, N1298);
and AND3 (N18049, N18044, N12612, N17046);
buf BUF1 (N18050, N18046);
nor NOR3 (N18051, N18045, N6694, N3958);
not NOT1 (N18052, N18048);
not NOT1 (N18053, N18052);
buf BUF1 (N18054, N18042);
not NOT1 (N18055, N18033);
nor NOR2 (N18056, N18041, N17320);
and AND2 (N18057, N18055, N3461);
nand NAND4 (N18058, N18051, N5964, N3011, N15688);
and AND2 (N18059, N18053, N7041);
not NOT1 (N18060, N18056);
buf BUF1 (N18061, N18060);
not NOT1 (N18062, N18058);
and AND3 (N18063, N18059, N2841, N3218);
and AND2 (N18064, N18062, N7823);
nand NAND4 (N18065, N18050, N5212, N15525, N331);
xor XOR2 (N18066, N18023, N4380);
buf BUF1 (N18067, N18049);
or OR4 (N18068, N18063, N16997, N16508, N12916);
nand NAND4 (N18069, N18064, N3702, N673, N16473);
xor XOR2 (N18070, N18065, N17051);
and AND2 (N18071, N18068, N4320);
or OR3 (N18072, N18069, N2480, N14131);
xor XOR2 (N18073, N18067, N12839);
nor NOR3 (N18074, N18054, N1932, N11801);
not NOT1 (N18075, N18047);
nor NOR3 (N18076, N18075, N800, N14833);
or OR2 (N18077, N18070, N13712);
nor NOR3 (N18078, N18061, N11217, N524);
or OR3 (N18079, N18057, N17663, N14807);
nor NOR4 (N18080, N18074, N17847, N11388, N17764);
buf BUF1 (N18081, N18080);
and AND4 (N18082, N18081, N17553, N5900, N2644);
nand NAND2 (N18083, N18071, N2504);
nor NOR2 (N18084, N18083, N1677);
or OR2 (N18085, N18082, N17531);
and AND2 (N18086, N18072, N16316);
nor NOR4 (N18087, N18085, N17949, N14995, N17179);
xor XOR2 (N18088, N18078, N6610);
not NOT1 (N18089, N18073);
not NOT1 (N18090, N18079);
not NOT1 (N18091, N18077);
not NOT1 (N18092, N18076);
buf BUF1 (N18093, N18092);
not NOT1 (N18094, N18088);
not NOT1 (N18095, N18094);
or OR3 (N18096, N18089, N12269, N10963);
buf BUF1 (N18097, N18093);
buf BUF1 (N18098, N18086);
and AND2 (N18099, N18095, N13192);
xor XOR2 (N18100, N18090, N12679);
buf BUF1 (N18101, N18097);
or OR3 (N18102, N18040, N4400, N499);
not NOT1 (N18103, N18096);
nand NAND3 (N18104, N18102, N14172, N10050);
and AND2 (N18105, N18104, N4629);
or OR3 (N18106, N18084, N1069, N6660);
nand NAND4 (N18107, N18106, N13126, N4298, N11306);
buf BUF1 (N18108, N18103);
or OR3 (N18109, N18066, N1231, N14240);
nor NOR4 (N18110, N18087, N3737, N5680, N15921);
xor XOR2 (N18111, N18109, N2300);
not NOT1 (N18112, N18091);
xor XOR2 (N18113, N18098, N618);
xor XOR2 (N18114, N18107, N16379);
buf BUF1 (N18115, N18113);
nand NAND4 (N18116, N18101, N8514, N6488, N5226);
xor XOR2 (N18117, N18099, N4422);
nor NOR2 (N18118, N18108, N9633);
or OR2 (N18119, N18114, N10518);
nand NAND4 (N18120, N18111, N3263, N9740, N6649);
buf BUF1 (N18121, N18110);
not NOT1 (N18122, N18119);
xor XOR2 (N18123, N18121, N6195);
or OR3 (N18124, N18115, N14298, N17365);
nor NOR3 (N18125, N18117, N2820, N5546);
nand NAND4 (N18126, N18122, N4850, N9858, N15529);
or OR4 (N18127, N18116, N1014, N10566, N11002);
xor XOR2 (N18128, N18127, N17737);
buf BUF1 (N18129, N18105);
nand NAND2 (N18130, N18100, N14367);
or OR3 (N18131, N18128, N11159, N10280);
not NOT1 (N18132, N18131);
buf BUF1 (N18133, N18129);
nor NOR2 (N18134, N18130, N16758);
not NOT1 (N18135, N18118);
nand NAND4 (N18136, N18123, N8304, N6611, N8676);
and AND4 (N18137, N18132, N15604, N8131, N3848);
or OR2 (N18138, N18137, N1594);
xor XOR2 (N18139, N18136, N15755);
or OR3 (N18140, N18126, N17489, N13760);
nand NAND2 (N18141, N18125, N6890);
or OR3 (N18142, N18112, N4887, N13466);
and AND2 (N18143, N18139, N15661);
buf BUF1 (N18144, N18120);
not NOT1 (N18145, N18133);
buf BUF1 (N18146, N18141);
nor NOR2 (N18147, N18124, N2663);
nor NOR2 (N18148, N18144, N9992);
or OR2 (N18149, N18148, N17979);
nor NOR2 (N18150, N18142, N16846);
xor XOR2 (N18151, N18147, N2141);
xor XOR2 (N18152, N18150, N1998);
not NOT1 (N18153, N18134);
buf BUF1 (N18154, N18140);
buf BUF1 (N18155, N18149);
xor XOR2 (N18156, N18146, N4559);
and AND3 (N18157, N18145, N12085, N11188);
xor XOR2 (N18158, N18152, N10163);
xor XOR2 (N18159, N18157, N8880);
nor NOR2 (N18160, N18154, N12984);
buf BUF1 (N18161, N18151);
or OR2 (N18162, N18138, N16384);
and AND2 (N18163, N18162, N11940);
xor XOR2 (N18164, N18135, N16052);
xor XOR2 (N18165, N18160, N13662);
nor NOR3 (N18166, N18156, N7562, N9909);
and AND2 (N18167, N18153, N16377);
nand NAND3 (N18168, N18165, N555, N10240);
or OR4 (N18169, N18158, N4924, N1682, N9606);
or OR4 (N18170, N18163, N10454, N3308, N9129);
nand NAND4 (N18171, N18159, N4476, N13784, N16842);
xor XOR2 (N18172, N18166, N11757);
xor XOR2 (N18173, N18169, N12911);
nor NOR3 (N18174, N18161, N2319, N13428);
or OR3 (N18175, N18171, N5157, N4521);
buf BUF1 (N18176, N18173);
not NOT1 (N18177, N18168);
xor XOR2 (N18178, N18155, N14353);
and AND3 (N18179, N18176, N6230, N3337);
xor XOR2 (N18180, N18174, N4524);
and AND2 (N18181, N18143, N3328);
not NOT1 (N18182, N18170);
not NOT1 (N18183, N18180);
buf BUF1 (N18184, N18177);
or OR3 (N18185, N18181, N15071, N10149);
buf BUF1 (N18186, N18185);
buf BUF1 (N18187, N18183);
nand NAND2 (N18188, N18178, N17382);
xor XOR2 (N18189, N18188, N3851);
and AND4 (N18190, N18164, N5730, N17637, N6033);
or OR4 (N18191, N18172, N12798, N12511, N6729);
not NOT1 (N18192, N18167);
or OR4 (N18193, N18190, N7851, N13174, N2214);
buf BUF1 (N18194, N18189);
and AND2 (N18195, N18186, N2069);
or OR4 (N18196, N18179, N16190, N227, N9969);
and AND2 (N18197, N18196, N5404);
not NOT1 (N18198, N18191);
nor NOR3 (N18199, N18184, N14200, N5587);
nor NOR2 (N18200, N18194, N3025);
or OR3 (N18201, N18193, N8354, N3278);
nand NAND2 (N18202, N18182, N3115);
or OR4 (N18203, N18198, N1640, N14216, N14894);
nand NAND2 (N18204, N18199, N14457);
not NOT1 (N18205, N18204);
buf BUF1 (N18206, N18175);
buf BUF1 (N18207, N18206);
xor XOR2 (N18208, N18203, N4455);
nor NOR2 (N18209, N18207, N10476);
buf BUF1 (N18210, N18208);
or OR3 (N18211, N18197, N10952, N14824);
not NOT1 (N18212, N18195);
buf BUF1 (N18213, N18201);
and AND4 (N18214, N18200, N18210, N2229, N15386);
not NOT1 (N18215, N269);
nand NAND4 (N18216, N18192, N14298, N6378, N11778);
and AND4 (N18217, N18187, N2286, N1849, N5667);
or OR4 (N18218, N18209, N11675, N10310, N3489);
and AND2 (N18219, N18214, N5590);
and AND3 (N18220, N18217, N1116, N6854);
and AND3 (N18221, N18220, N7038, N10901);
and AND2 (N18222, N18215, N9034);
buf BUF1 (N18223, N18216);
or OR4 (N18224, N18222, N8906, N17016, N6686);
and AND3 (N18225, N18219, N5861, N11000);
buf BUF1 (N18226, N18223);
nand NAND2 (N18227, N18205, N13731);
nor NOR4 (N18228, N18218, N9285, N3888, N5099);
or OR4 (N18229, N18225, N14888, N17479, N9198);
nand NAND3 (N18230, N18227, N14124, N18174);
not NOT1 (N18231, N18211);
and AND3 (N18232, N18221, N10818, N11475);
or OR2 (N18233, N18213, N16839);
buf BUF1 (N18234, N18202);
and AND4 (N18235, N18230, N10564, N8806, N2226);
nand NAND3 (N18236, N18231, N8646, N1780);
nand NAND4 (N18237, N18226, N5164, N15666, N9273);
not NOT1 (N18238, N18229);
nand NAND3 (N18239, N18234, N6213, N11820);
and AND4 (N18240, N18238, N16175, N7712, N16479);
nand NAND4 (N18241, N18232, N7532, N10771, N3593);
or OR4 (N18242, N18241, N2345, N2263, N11192);
not NOT1 (N18243, N18240);
nand NAND4 (N18244, N18237, N9978, N6416, N2206);
xor XOR2 (N18245, N18228, N2365);
xor XOR2 (N18246, N18239, N7675);
buf BUF1 (N18247, N18246);
buf BUF1 (N18248, N18235);
and AND3 (N18249, N18244, N14302, N7230);
or OR3 (N18250, N18236, N10113, N5979);
nor NOR2 (N18251, N18247, N10633);
or OR4 (N18252, N18251, N1874, N14596, N2839);
buf BUF1 (N18253, N18249);
nor NOR3 (N18254, N18250, N4054, N7190);
buf BUF1 (N18255, N18242);
nand NAND3 (N18256, N18254, N16733, N3441);
and AND2 (N18257, N18248, N5880);
buf BUF1 (N18258, N18255);
or OR2 (N18259, N18245, N16542);
nand NAND2 (N18260, N18259, N7266);
nor NOR2 (N18261, N18258, N11417);
xor XOR2 (N18262, N18257, N8870);
buf BUF1 (N18263, N18243);
xor XOR2 (N18264, N18224, N2692);
buf BUF1 (N18265, N18264);
xor XOR2 (N18266, N18212, N17063);
nor NOR3 (N18267, N18265, N7923, N8157);
and AND4 (N18268, N18256, N11212, N3173, N17728);
xor XOR2 (N18269, N18253, N10229);
buf BUF1 (N18270, N18262);
xor XOR2 (N18271, N18261, N13023);
or OR2 (N18272, N18252, N2095);
and AND3 (N18273, N18233, N1927, N12534);
buf BUF1 (N18274, N18269);
and AND4 (N18275, N18270, N15212, N17321, N17392);
buf BUF1 (N18276, N18268);
nand NAND3 (N18277, N18275, N11602, N5314);
nand NAND3 (N18278, N18276, N17304, N13469);
buf BUF1 (N18279, N18260);
not NOT1 (N18280, N18273);
not NOT1 (N18281, N18267);
buf BUF1 (N18282, N18274);
buf BUF1 (N18283, N18271);
nor NOR4 (N18284, N18278, N15719, N4010, N13953);
not NOT1 (N18285, N18282);
buf BUF1 (N18286, N18281);
or OR4 (N18287, N18279, N6749, N8624, N7100);
buf BUF1 (N18288, N18284);
nand NAND2 (N18289, N18277, N13231);
xor XOR2 (N18290, N18287, N16580);
or OR2 (N18291, N18272, N849);
not NOT1 (N18292, N18283);
xor XOR2 (N18293, N18289, N12459);
nand NAND2 (N18294, N18293, N12357);
not NOT1 (N18295, N18266);
nor NOR4 (N18296, N18292, N18228, N5336, N4350);
nor NOR3 (N18297, N18285, N10696, N11908);
buf BUF1 (N18298, N18294);
buf BUF1 (N18299, N18297);
buf BUF1 (N18300, N18296);
or OR4 (N18301, N18291, N11200, N10765, N11824);
xor XOR2 (N18302, N18295, N15401);
buf BUF1 (N18303, N18302);
nor NOR2 (N18304, N18263, N13376);
buf BUF1 (N18305, N18288);
xor XOR2 (N18306, N18280, N7941);
nand NAND3 (N18307, N18299, N8272, N4343);
nand NAND2 (N18308, N18306, N4957);
or OR2 (N18309, N18304, N769);
buf BUF1 (N18310, N18298);
buf BUF1 (N18311, N18309);
xor XOR2 (N18312, N18301, N16909);
or OR4 (N18313, N18303, N16013, N12846, N17857);
not NOT1 (N18314, N18305);
nor NOR3 (N18315, N18307, N13184, N10044);
nand NAND2 (N18316, N18310, N3294);
not NOT1 (N18317, N18315);
not NOT1 (N18318, N18313);
buf BUF1 (N18319, N18290);
nor NOR3 (N18320, N18319, N13108, N12610);
xor XOR2 (N18321, N18286, N6523);
and AND4 (N18322, N18312, N9262, N10104, N17521);
xor XOR2 (N18323, N18321, N17081);
buf BUF1 (N18324, N18316);
nor NOR4 (N18325, N18323, N9117, N11428, N4319);
buf BUF1 (N18326, N18318);
not NOT1 (N18327, N18311);
not NOT1 (N18328, N18317);
nor NOR3 (N18329, N18324, N1112, N7242);
xor XOR2 (N18330, N18322, N17358);
buf BUF1 (N18331, N18308);
buf BUF1 (N18332, N18320);
and AND2 (N18333, N18332, N18130);
xor XOR2 (N18334, N18331, N12872);
buf BUF1 (N18335, N18327);
or OR4 (N18336, N18333, N3997, N11585, N1066);
not NOT1 (N18337, N18336);
buf BUF1 (N18338, N18334);
buf BUF1 (N18339, N18314);
xor XOR2 (N18340, N18337, N15738);
or OR3 (N18341, N18340, N7137, N1531);
buf BUF1 (N18342, N18338);
nor NOR2 (N18343, N18300, N1288);
not NOT1 (N18344, N18343);
not NOT1 (N18345, N18328);
or OR3 (N18346, N18335, N5036, N14149);
and AND4 (N18347, N18346, N14120, N14874, N11099);
and AND2 (N18348, N18344, N13849);
and AND2 (N18349, N18348, N7953);
not NOT1 (N18350, N18347);
nor NOR4 (N18351, N18345, N1279, N17271, N13103);
and AND2 (N18352, N18341, N3368);
and AND3 (N18353, N18326, N13736, N11553);
or OR3 (N18354, N18352, N12414, N12591);
or OR2 (N18355, N18354, N15843);
and AND4 (N18356, N18325, N17202, N6489, N7974);
xor XOR2 (N18357, N18356, N15467);
not NOT1 (N18358, N18349);
nand NAND2 (N18359, N18358, N11862);
not NOT1 (N18360, N18330);
and AND4 (N18361, N18350, N17312, N8280, N829);
nand NAND3 (N18362, N18360, N1983, N4225);
buf BUF1 (N18363, N18329);
or OR3 (N18364, N18353, N18124, N15199);
nand NAND2 (N18365, N18363, N1698);
nand NAND4 (N18366, N18364, N3280, N6665, N10001);
nand NAND2 (N18367, N18366, N6688);
xor XOR2 (N18368, N18339, N8876);
and AND4 (N18369, N18342, N10683, N15123, N3604);
nand NAND2 (N18370, N18367, N11972);
or OR2 (N18371, N18370, N765);
and AND2 (N18372, N18361, N13622);
not NOT1 (N18373, N18357);
nand NAND3 (N18374, N18355, N5415, N11321);
nand NAND4 (N18375, N18365, N17107, N10060, N5054);
not NOT1 (N18376, N18373);
and AND4 (N18377, N18371, N1943, N4339, N6180);
xor XOR2 (N18378, N18375, N7062);
xor XOR2 (N18379, N18377, N6633);
xor XOR2 (N18380, N18372, N13881);
buf BUF1 (N18381, N18362);
xor XOR2 (N18382, N18351, N2138);
nor NOR3 (N18383, N18380, N14777, N15558);
not NOT1 (N18384, N18359);
nor NOR4 (N18385, N18384, N3666, N3883, N10965);
not NOT1 (N18386, N18385);
and AND2 (N18387, N18376, N16496);
xor XOR2 (N18388, N18382, N614);
not NOT1 (N18389, N18369);
and AND2 (N18390, N18379, N11302);
nand NAND4 (N18391, N18390, N4080, N6942, N4637);
and AND4 (N18392, N18387, N7235, N14836, N4795);
xor XOR2 (N18393, N18368, N12200);
xor XOR2 (N18394, N18383, N4096);
buf BUF1 (N18395, N18388);
not NOT1 (N18396, N18389);
not NOT1 (N18397, N18393);
buf BUF1 (N18398, N18392);
buf BUF1 (N18399, N18374);
nand NAND4 (N18400, N18381, N1454, N10281, N11054);
not NOT1 (N18401, N18395);
not NOT1 (N18402, N18400);
nor NOR3 (N18403, N18397, N2287, N5468);
nor NOR4 (N18404, N18386, N6801, N12698, N4321);
buf BUF1 (N18405, N18401);
or OR4 (N18406, N18398, N3763, N17725, N17555);
nand NAND3 (N18407, N18394, N10004, N12923);
xor XOR2 (N18408, N18396, N11021);
nor NOR4 (N18409, N18408, N10323, N14775, N1337);
xor XOR2 (N18410, N18404, N10351);
not NOT1 (N18411, N18402);
not NOT1 (N18412, N18407);
and AND2 (N18413, N18406, N11621);
xor XOR2 (N18414, N18405, N9141);
not NOT1 (N18415, N18391);
and AND4 (N18416, N18410, N15015, N17207, N12930);
nor NOR4 (N18417, N18412, N7161, N14160, N10724);
and AND3 (N18418, N18378, N14540, N4923);
xor XOR2 (N18419, N18409, N7510);
not NOT1 (N18420, N18399);
nor NOR2 (N18421, N18419, N1287);
or OR3 (N18422, N18414, N12944, N6668);
xor XOR2 (N18423, N18403, N14701);
nor NOR4 (N18424, N18421, N2215, N2046, N12715);
not NOT1 (N18425, N18423);
buf BUF1 (N18426, N18416);
not NOT1 (N18427, N18422);
nand NAND2 (N18428, N18415, N4453);
nor NOR4 (N18429, N18417, N5301, N4975, N5018);
and AND3 (N18430, N18425, N4373, N18215);
xor XOR2 (N18431, N18430, N4369);
or OR2 (N18432, N18424, N4199);
xor XOR2 (N18433, N18428, N12117);
and AND3 (N18434, N18433, N16061, N13229);
or OR4 (N18435, N18427, N12552, N18369, N13575);
xor XOR2 (N18436, N18434, N17650);
buf BUF1 (N18437, N18413);
nor NOR4 (N18438, N18420, N17407, N7874, N8868);
xor XOR2 (N18439, N18436, N17511);
and AND4 (N18440, N18426, N2518, N3877, N244);
not NOT1 (N18441, N18429);
nand NAND2 (N18442, N18437, N18218);
or OR3 (N18443, N18431, N3566, N12120);
xor XOR2 (N18444, N18438, N12197);
xor XOR2 (N18445, N18442, N2539);
or OR2 (N18446, N18440, N14275);
nand NAND4 (N18447, N18411, N16120, N14340, N3039);
nand NAND3 (N18448, N18432, N3940, N15428);
and AND3 (N18449, N18435, N16425, N11458);
and AND4 (N18450, N18441, N2133, N10321, N16464);
or OR2 (N18451, N18448, N8293);
and AND4 (N18452, N18449, N13917, N4162, N10344);
nor NOR3 (N18453, N18445, N8401, N15388);
and AND3 (N18454, N18444, N14581, N13885);
and AND4 (N18455, N18447, N8130, N16000, N6555);
or OR4 (N18456, N18451, N3921, N7566, N17015);
not NOT1 (N18457, N18439);
nand NAND4 (N18458, N18452, N2530, N7717, N12078);
and AND3 (N18459, N18456, N12818, N15959);
or OR2 (N18460, N18453, N3641);
not NOT1 (N18461, N18459);
and AND4 (N18462, N18450, N4060, N16126, N14114);
nor NOR3 (N18463, N18446, N10420, N4625);
xor XOR2 (N18464, N18462, N10904);
and AND2 (N18465, N18460, N2704);
xor XOR2 (N18466, N18457, N4678);
or OR4 (N18467, N18464, N211, N5748, N2116);
buf BUF1 (N18468, N18463);
and AND3 (N18469, N18454, N16243, N951);
nand NAND2 (N18470, N18458, N11801);
nand NAND2 (N18471, N18468, N8363);
or OR2 (N18472, N18467, N12952);
not NOT1 (N18473, N18471);
or OR4 (N18474, N18455, N18005, N6676, N18019);
and AND4 (N18475, N18474, N8197, N9434, N1156);
and AND2 (N18476, N18472, N13249);
not NOT1 (N18477, N18418);
or OR4 (N18478, N18473, N9281, N7108, N849);
xor XOR2 (N18479, N18476, N603);
nand NAND4 (N18480, N18469, N6581, N8360, N9471);
nor NOR4 (N18481, N18477, N10950, N16169, N17512);
nor NOR3 (N18482, N18479, N6188, N2880);
buf BUF1 (N18483, N18480);
buf BUF1 (N18484, N18483);
nor NOR4 (N18485, N18466, N7167, N14652, N8681);
nor NOR3 (N18486, N18465, N14950, N13260);
nand NAND3 (N18487, N18478, N16539, N8109);
nand NAND3 (N18488, N18484, N3621, N17971);
or OR3 (N18489, N18488, N4353, N8322);
and AND4 (N18490, N18485, N11068, N15906, N16069);
buf BUF1 (N18491, N18489);
buf BUF1 (N18492, N18470);
and AND4 (N18493, N18481, N5484, N190, N15210);
not NOT1 (N18494, N18443);
nand NAND2 (N18495, N18493, N4045);
nor NOR4 (N18496, N18487, N7140, N738, N578);
or OR4 (N18497, N18495, N8645, N8047, N10148);
nor NOR3 (N18498, N18497, N17107, N332);
xor XOR2 (N18499, N18482, N10321);
not NOT1 (N18500, N18461);
or OR2 (N18501, N18498, N5999);
and AND4 (N18502, N18494, N18500, N17523, N14085);
xor XOR2 (N18503, N14743, N9596);
nor NOR2 (N18504, N18503, N7991);
or OR2 (N18505, N18496, N13241);
or OR3 (N18506, N18501, N6457, N4557);
nand NAND3 (N18507, N18505, N6182, N6553);
nor NOR2 (N18508, N18475, N2398);
xor XOR2 (N18509, N18492, N2643);
buf BUF1 (N18510, N18508);
xor XOR2 (N18511, N18506, N16534);
or OR3 (N18512, N18499, N3545, N15368);
or OR4 (N18513, N18510, N14560, N12634, N2566);
nand NAND2 (N18514, N18512, N18470);
or OR3 (N18515, N18513, N12575, N7469);
buf BUF1 (N18516, N18514);
and AND2 (N18517, N18507, N7814);
nand NAND4 (N18518, N18490, N2701, N10168, N4020);
nor NOR2 (N18519, N18515, N10363);
or OR3 (N18520, N18511, N16092, N9511);
buf BUF1 (N18521, N18509);
or OR2 (N18522, N18486, N13102);
xor XOR2 (N18523, N18520, N10250);
nor NOR2 (N18524, N18521, N15549);
nand NAND4 (N18525, N18517, N8279, N4051, N8699);
nand NAND3 (N18526, N18504, N17515, N8281);
nand NAND3 (N18527, N18526, N661, N8823);
nor NOR2 (N18528, N18502, N1057);
not NOT1 (N18529, N18491);
nand NAND4 (N18530, N18523, N10286, N13773, N14600);
and AND2 (N18531, N18519, N18359);
nor NOR4 (N18532, N18529, N12966, N753, N17696);
or OR2 (N18533, N18522, N9586);
not NOT1 (N18534, N18527);
nand NAND4 (N18535, N18524, N1142, N15555, N7732);
buf BUF1 (N18536, N18535);
nor NOR3 (N18537, N18518, N821, N8059);
nor NOR4 (N18538, N18534, N276, N15517, N5805);
buf BUF1 (N18539, N18516);
and AND4 (N18540, N18539, N12714, N2617, N13584);
and AND3 (N18541, N18532, N8190, N126);
and AND2 (N18542, N18536, N8407);
or OR3 (N18543, N18538, N1631, N732);
or OR4 (N18544, N18542, N1944, N313, N11702);
nor NOR2 (N18545, N18528, N1335);
or OR2 (N18546, N18545, N1210);
and AND2 (N18547, N18546, N7063);
and AND3 (N18548, N18547, N15222, N3070);
xor XOR2 (N18549, N18537, N18074);
xor XOR2 (N18550, N18530, N10862);
nand NAND2 (N18551, N18549, N2370);
buf BUF1 (N18552, N18525);
not NOT1 (N18553, N18541);
not NOT1 (N18554, N18553);
nor NOR3 (N18555, N18550, N6773, N14419);
nand NAND4 (N18556, N18533, N1069, N10296, N6842);
and AND4 (N18557, N18548, N10925, N7077, N5639);
or OR3 (N18558, N18544, N15134, N17288);
nand NAND2 (N18559, N18551, N2804);
buf BUF1 (N18560, N18543);
or OR2 (N18561, N18558, N8574);
not NOT1 (N18562, N18556);
nor NOR4 (N18563, N18540, N12731, N6466, N16063);
nand NAND4 (N18564, N18559, N1934, N15104, N3104);
xor XOR2 (N18565, N18531, N13290);
or OR2 (N18566, N18552, N5600);
and AND4 (N18567, N18555, N18346, N724, N3334);
and AND4 (N18568, N18567, N612, N5907, N12504);
nand NAND2 (N18569, N18563, N16357);
nand NAND3 (N18570, N18554, N2514, N3086);
buf BUF1 (N18571, N18568);
not NOT1 (N18572, N18570);
or OR4 (N18573, N18557, N6204, N8110, N3870);
nor NOR3 (N18574, N18560, N15414, N12423);
nor NOR3 (N18575, N18565, N9108, N7433);
not NOT1 (N18576, N18575);
nor NOR3 (N18577, N18573, N5005, N7846);
not NOT1 (N18578, N18572);
xor XOR2 (N18579, N18576, N18167);
and AND4 (N18580, N18569, N8563, N11809, N5743);
or OR3 (N18581, N18566, N11651, N14259);
or OR4 (N18582, N18580, N11771, N15411, N10055);
not NOT1 (N18583, N18574);
buf BUF1 (N18584, N18582);
nor NOR4 (N18585, N18584, N10484, N8674, N16321);
and AND2 (N18586, N18579, N7566);
nor NOR2 (N18587, N18578, N11763);
nand NAND4 (N18588, N18581, N16451, N6961, N2375);
xor XOR2 (N18589, N18577, N12869);
xor XOR2 (N18590, N18583, N5135);
and AND4 (N18591, N18587, N13723, N13838, N18302);
or OR4 (N18592, N18585, N10310, N16363, N9928);
xor XOR2 (N18593, N18588, N740);
and AND3 (N18594, N18591, N14130, N2394);
buf BUF1 (N18595, N18586);
nor NOR2 (N18596, N18561, N14575);
not NOT1 (N18597, N18562);
nor NOR3 (N18598, N18592, N9820, N8219);
nor NOR3 (N18599, N18598, N9326, N16662);
buf BUF1 (N18600, N18595);
buf BUF1 (N18601, N18599);
not NOT1 (N18602, N18596);
or OR2 (N18603, N18564, N2204);
nand NAND4 (N18604, N18590, N17002, N11479, N11688);
not NOT1 (N18605, N18593);
and AND3 (N18606, N18600, N12228, N5412);
or OR4 (N18607, N18594, N17906, N4437, N14351);
nand NAND3 (N18608, N18602, N9008, N4967);
or OR2 (N18609, N18605, N15876);
and AND2 (N18610, N18603, N759);
nor NOR4 (N18611, N18610, N5248, N17667, N6308);
buf BUF1 (N18612, N18611);
nor NOR4 (N18613, N18601, N8390, N1057, N12170);
nand NAND2 (N18614, N18608, N6553);
nand NAND2 (N18615, N18604, N17722);
or OR2 (N18616, N18615, N2485);
not NOT1 (N18617, N18607);
and AND2 (N18618, N18614, N12645);
and AND3 (N18619, N18609, N9329, N12710);
not NOT1 (N18620, N18616);
nand NAND2 (N18621, N18597, N10577);
xor XOR2 (N18622, N18571, N743);
not NOT1 (N18623, N18622);
nor NOR4 (N18624, N18620, N892, N16590, N3658);
buf BUF1 (N18625, N18619);
nand NAND3 (N18626, N18624, N4561, N493);
and AND3 (N18627, N18626, N5977, N7857);
not NOT1 (N18628, N18618);
not NOT1 (N18629, N18625);
nor NOR2 (N18630, N18627, N16402);
or OR4 (N18631, N18606, N2786, N577, N7760);
or OR4 (N18632, N18628, N14944, N7338, N4008);
or OR3 (N18633, N18631, N2861, N12251);
buf BUF1 (N18634, N18629);
and AND2 (N18635, N18623, N12290);
or OR2 (N18636, N18632, N1875);
not NOT1 (N18637, N18635);
nor NOR2 (N18638, N18634, N17162);
nand NAND2 (N18639, N18636, N17205);
nor NOR3 (N18640, N18617, N872, N16692);
or OR4 (N18641, N18639, N274, N4093, N16000);
not NOT1 (N18642, N18637);
nand NAND2 (N18643, N18641, N6802);
or OR4 (N18644, N18630, N2194, N5892, N13353);
and AND4 (N18645, N18621, N481, N14611, N6398);
not NOT1 (N18646, N18640);
and AND4 (N18647, N18613, N2550, N874, N6171);
nor NOR4 (N18648, N18644, N11542, N3009, N4889);
or OR3 (N18649, N18648, N1352, N4526);
buf BUF1 (N18650, N18633);
and AND3 (N18651, N18642, N1112, N3443);
or OR2 (N18652, N18643, N3943);
or OR3 (N18653, N18650, N1161, N1394);
nand NAND2 (N18654, N18612, N5144);
and AND4 (N18655, N18654, N10880, N5589, N11474);
or OR3 (N18656, N18653, N1821, N15598);
and AND3 (N18657, N18652, N13684, N2941);
xor XOR2 (N18658, N18656, N15433);
buf BUF1 (N18659, N18646);
xor XOR2 (N18660, N18649, N3780);
nor NOR2 (N18661, N18659, N2664);
or OR4 (N18662, N18661, N5932, N7434, N15264);
not NOT1 (N18663, N18655);
nand NAND2 (N18664, N18589, N8954);
buf BUF1 (N18665, N18651);
nor NOR2 (N18666, N18658, N9512);
not NOT1 (N18667, N18666);
nand NAND3 (N18668, N18660, N12953, N9054);
or OR3 (N18669, N18647, N15103, N97);
buf BUF1 (N18670, N18668);
nand NAND3 (N18671, N18665, N2539, N4444);
and AND4 (N18672, N18638, N16740, N5194, N13159);
nor NOR4 (N18673, N18672, N3721, N8116, N3615);
and AND2 (N18674, N18662, N4014);
not NOT1 (N18675, N18657);
and AND4 (N18676, N18673, N2487, N41, N13602);
nor NOR2 (N18677, N18675, N8812);
or OR3 (N18678, N18667, N8945, N8537);
not NOT1 (N18679, N18678);
nor NOR3 (N18680, N18663, N2134, N3406);
or OR4 (N18681, N18671, N18207, N360, N10259);
or OR4 (N18682, N18645, N9479, N16895, N5242);
or OR4 (N18683, N18677, N9369, N9545, N18467);
nor NOR2 (N18684, N18664, N15998);
not NOT1 (N18685, N18679);
and AND4 (N18686, N18685, N17139, N12985, N16898);
nand NAND3 (N18687, N18686, N6850, N1734);
xor XOR2 (N18688, N18669, N11910);
or OR2 (N18689, N18682, N6220);
buf BUF1 (N18690, N18688);
not NOT1 (N18691, N18674);
and AND4 (N18692, N18676, N16902, N15774, N13477);
xor XOR2 (N18693, N18689, N2308);
xor XOR2 (N18694, N18693, N2052);
not NOT1 (N18695, N18687);
not NOT1 (N18696, N18681);
nand NAND3 (N18697, N18692, N12910, N11708);
xor XOR2 (N18698, N18691, N15357);
or OR3 (N18699, N18684, N7270, N8471);
nand NAND3 (N18700, N18670, N6444, N2685);
buf BUF1 (N18701, N18694);
not NOT1 (N18702, N18701);
and AND2 (N18703, N18699, N5583);
and AND3 (N18704, N18697, N11267, N8388);
xor XOR2 (N18705, N18698, N16034);
not NOT1 (N18706, N18704);
xor XOR2 (N18707, N18700, N1451);
nor NOR2 (N18708, N18705, N14967);
or OR3 (N18709, N18702, N4155, N14037);
and AND2 (N18710, N18696, N4151);
xor XOR2 (N18711, N18683, N6276);
and AND2 (N18712, N18711, N13226);
not NOT1 (N18713, N18706);
and AND2 (N18714, N18713, N15337);
xor XOR2 (N18715, N18709, N7083);
buf BUF1 (N18716, N18695);
not NOT1 (N18717, N18712);
not NOT1 (N18718, N18714);
and AND3 (N18719, N18703, N4793, N4485);
nor NOR3 (N18720, N18715, N2547, N958);
or OR3 (N18721, N18680, N13644, N2282);
and AND4 (N18722, N18717, N3566, N11030, N915);
buf BUF1 (N18723, N18719);
or OR4 (N18724, N18720, N10188, N5430, N2459);
or OR3 (N18725, N18707, N8494, N6777);
nor NOR4 (N18726, N18710, N1322, N4593, N11065);
nor NOR2 (N18727, N18718, N4281);
nand NAND2 (N18728, N18725, N1167);
nand NAND4 (N18729, N18726, N10694, N2097, N1972);
or OR4 (N18730, N18716, N7174, N12266, N13735);
or OR3 (N18731, N18724, N1513, N16153);
not NOT1 (N18732, N18722);
nor NOR2 (N18733, N18727, N8890);
nand NAND4 (N18734, N18728, N7619, N13515, N15348);
xor XOR2 (N18735, N18732, N17589);
or OR3 (N18736, N18729, N2079, N16387);
buf BUF1 (N18737, N18734);
or OR3 (N18738, N18735, N2341, N7235);
buf BUF1 (N18739, N18690);
buf BUF1 (N18740, N18721);
not NOT1 (N18741, N18738);
nand NAND3 (N18742, N18730, N1975, N16794);
and AND3 (N18743, N18723, N11556, N16637);
nand NAND2 (N18744, N18743, N17583);
buf BUF1 (N18745, N18741);
not NOT1 (N18746, N18737);
nor NOR2 (N18747, N18740, N4894);
xor XOR2 (N18748, N18747, N11515);
and AND3 (N18749, N18739, N2174, N6615);
xor XOR2 (N18750, N18746, N818);
nand NAND3 (N18751, N18749, N6116, N17330);
nor NOR4 (N18752, N18750, N12453, N1998, N9886);
not NOT1 (N18753, N18742);
not NOT1 (N18754, N18752);
or OR4 (N18755, N18751, N6501, N10187, N10417);
and AND2 (N18756, N18744, N3595);
buf BUF1 (N18757, N18748);
nand NAND2 (N18758, N18756, N9542);
nand NAND3 (N18759, N18736, N1142, N13705);
and AND2 (N18760, N18755, N12515);
and AND3 (N18761, N18733, N13226, N5619);
and AND4 (N18762, N18708, N7238, N14442, N17741);
nand NAND3 (N18763, N18754, N5961, N9462);
buf BUF1 (N18764, N18759);
nor NOR2 (N18765, N18764, N11197);
nand NAND4 (N18766, N18765, N9298, N11802, N1791);
not NOT1 (N18767, N18762);
and AND3 (N18768, N18761, N17218, N1789);
buf BUF1 (N18769, N18758);
nor NOR3 (N18770, N18769, N4177, N16082);
and AND3 (N18771, N18763, N14061, N13866);
not NOT1 (N18772, N18745);
and AND2 (N18773, N18760, N15817);
nand NAND3 (N18774, N18767, N5515, N11040);
not NOT1 (N18775, N18773);
buf BUF1 (N18776, N18766);
not NOT1 (N18777, N18775);
or OR2 (N18778, N18731, N7474);
not NOT1 (N18779, N18768);
or OR4 (N18780, N18778, N12665, N341, N7472);
nor NOR4 (N18781, N18753, N5902, N9899, N5486);
nor NOR2 (N18782, N18777, N14523);
not NOT1 (N18783, N18780);
nand NAND2 (N18784, N18782, N4076);
nand NAND3 (N18785, N18757, N1969, N4971);
nand NAND2 (N18786, N18783, N14110);
xor XOR2 (N18787, N18771, N10835);
not NOT1 (N18788, N18784);
xor XOR2 (N18789, N18788, N14895);
nand NAND4 (N18790, N18785, N13038, N18773, N5656);
nand NAND2 (N18791, N18786, N6023);
and AND4 (N18792, N18791, N13393, N363, N2458);
not NOT1 (N18793, N18774);
nor NOR2 (N18794, N18772, N9728);
nand NAND4 (N18795, N18787, N5861, N7096, N1328);
or OR2 (N18796, N18794, N885);
nor NOR3 (N18797, N18795, N9796, N15414);
not NOT1 (N18798, N18792);
buf BUF1 (N18799, N18797);
nor NOR2 (N18800, N18798, N6478);
nand NAND2 (N18801, N18796, N16537);
or OR4 (N18802, N18790, N673, N8690, N7785);
not NOT1 (N18803, N18779);
not NOT1 (N18804, N18803);
nor NOR4 (N18805, N18776, N5681, N4940, N10388);
nor NOR3 (N18806, N18800, N10065, N6267);
nand NAND4 (N18807, N18802, N17939, N8812, N8189);
nand NAND4 (N18808, N18799, N7217, N12292, N13706);
nand NAND4 (N18809, N18806, N3721, N13929, N16062);
and AND3 (N18810, N18793, N17890, N469);
nand NAND4 (N18811, N18809, N13897, N1124, N4972);
or OR3 (N18812, N18770, N18680, N12006);
nand NAND4 (N18813, N18808, N1776, N3470, N10627);
and AND2 (N18814, N18810, N12222);
not NOT1 (N18815, N18781);
nor NOR3 (N18816, N18814, N18809, N5295);
nor NOR3 (N18817, N18804, N17029, N7492);
nor NOR3 (N18818, N18811, N3433, N1345);
or OR4 (N18819, N18818, N999, N7365, N17455);
and AND4 (N18820, N18807, N16571, N17236, N10931);
and AND4 (N18821, N18789, N14511, N8478, N14425);
nor NOR2 (N18822, N18820, N8549);
buf BUF1 (N18823, N18813);
nand NAND2 (N18824, N18816, N14385);
nor NOR4 (N18825, N18817, N3936, N10251, N16799);
or OR4 (N18826, N18819, N15542, N1015, N3349);
nor NOR3 (N18827, N18826, N7646, N18802);
not NOT1 (N18828, N18823);
and AND4 (N18829, N18812, N8099, N14476, N5711);
and AND2 (N18830, N18822, N11031);
nor NOR3 (N18831, N18821, N5205, N15585);
not NOT1 (N18832, N18825);
not NOT1 (N18833, N18827);
and AND2 (N18834, N18830, N10841);
or OR4 (N18835, N18834, N10773, N18580, N15830);
nand NAND2 (N18836, N18805, N17185);
and AND3 (N18837, N18835, N6734, N9);
nand NAND3 (N18838, N18836, N9318, N1035);
buf BUF1 (N18839, N18829);
nand NAND3 (N18840, N18815, N12768, N5841);
or OR4 (N18841, N18838, N1018, N16220, N2574);
and AND2 (N18842, N18841, N5483);
and AND3 (N18843, N18840, N13344, N9849);
nand NAND4 (N18844, N18824, N17415, N14283, N4334);
nand NAND4 (N18845, N18828, N9838, N8996, N17183);
nand NAND2 (N18846, N18801, N15593);
and AND4 (N18847, N18839, N13428, N8895, N9910);
and AND4 (N18848, N18831, N17487, N16117, N12143);
nor NOR3 (N18849, N18837, N12900, N5171);
buf BUF1 (N18850, N18843);
or OR4 (N18851, N18849, N10432, N17733, N12158);
and AND2 (N18852, N18842, N18632);
nor NOR4 (N18853, N18847, N13967, N2017, N12884);
or OR2 (N18854, N18852, N4059);
buf BUF1 (N18855, N18844);
buf BUF1 (N18856, N18833);
xor XOR2 (N18857, N18853, N7260);
xor XOR2 (N18858, N18856, N7738);
not NOT1 (N18859, N18846);
buf BUF1 (N18860, N18857);
nor NOR2 (N18861, N18855, N2781);
nand NAND3 (N18862, N18858, N16129, N4106);
nand NAND4 (N18863, N18854, N5981, N6062, N18775);
nand NAND4 (N18864, N18845, N3582, N13769, N4361);
xor XOR2 (N18865, N18860, N10621);
buf BUF1 (N18866, N18861);
xor XOR2 (N18867, N18832, N2800);
nand NAND2 (N18868, N18848, N14234);
nor NOR2 (N18869, N18863, N17069);
nor NOR3 (N18870, N18868, N1124, N16992);
buf BUF1 (N18871, N18850);
buf BUF1 (N18872, N18862);
and AND2 (N18873, N18864, N12738);
or OR2 (N18874, N18870, N685);
and AND4 (N18875, N18873, N4866, N210, N15933);
not NOT1 (N18876, N18875);
not NOT1 (N18877, N18871);
nand NAND3 (N18878, N18872, N9602, N15745);
or OR4 (N18879, N18865, N13164, N15103, N17895);
nand NAND4 (N18880, N18877, N11510, N13645, N17691);
not NOT1 (N18881, N18867);
buf BUF1 (N18882, N18859);
nor NOR3 (N18883, N18874, N12000, N18535);
nand NAND3 (N18884, N18869, N11718, N13173);
nor NOR3 (N18885, N18881, N7536, N8219);
xor XOR2 (N18886, N18878, N11450);
or OR3 (N18887, N18885, N1845, N1695);
nor NOR3 (N18888, N18866, N5798, N386);
buf BUF1 (N18889, N18886);
not NOT1 (N18890, N18851);
and AND2 (N18891, N18876, N3918);
xor XOR2 (N18892, N18884, N2399);
xor XOR2 (N18893, N18883, N6018);
nor NOR3 (N18894, N18882, N6900, N11099);
and AND3 (N18895, N18879, N112, N7225);
xor XOR2 (N18896, N18889, N10633);
not NOT1 (N18897, N18891);
or OR2 (N18898, N18888, N3895);
not NOT1 (N18899, N18897);
or OR2 (N18900, N18898, N13409);
buf BUF1 (N18901, N18896);
nand NAND3 (N18902, N18887, N3361, N17863);
nor NOR2 (N18903, N18892, N11001);
and AND4 (N18904, N18893, N1126, N17219, N4812);
not NOT1 (N18905, N18895);
or OR3 (N18906, N18901, N12345, N4148);
nand NAND3 (N18907, N18905, N10866, N2342);
nor NOR2 (N18908, N18880, N115);
nor NOR4 (N18909, N18908, N16738, N18349, N15433);
nand NAND4 (N18910, N18906, N4810, N8285, N6153);
buf BUF1 (N18911, N18894);
nand NAND2 (N18912, N18903, N1652);
nand NAND2 (N18913, N18910, N17765);
nor NOR3 (N18914, N18900, N8058, N505);
nand NAND2 (N18915, N18914, N15175);
and AND2 (N18916, N18890, N1752);
or OR4 (N18917, N18915, N3837, N9368, N17202);
or OR3 (N18918, N18913, N16171, N7778);
or OR2 (N18919, N18907, N3660);
and AND4 (N18920, N18911, N14426, N975, N12448);
xor XOR2 (N18921, N18916, N16584);
and AND4 (N18922, N18909, N13436, N13685, N12813);
buf BUF1 (N18923, N18904);
buf BUF1 (N18924, N18920);
nor NOR4 (N18925, N18912, N2442, N3179, N5548);
buf BUF1 (N18926, N18923);
not NOT1 (N18927, N18917);
buf BUF1 (N18928, N18919);
nor NOR2 (N18929, N18928, N101);
nand NAND3 (N18930, N18918, N8745, N14504);
and AND3 (N18931, N18902, N3539, N8911);
and AND4 (N18932, N18931, N9697, N13356, N18419);
nor NOR2 (N18933, N18932, N9614);
not NOT1 (N18934, N18921);
xor XOR2 (N18935, N18927, N5051);
nor NOR2 (N18936, N18929, N15191);
buf BUF1 (N18937, N18925);
or OR3 (N18938, N18936, N7847, N10684);
and AND3 (N18939, N18899, N8489, N240);
nor NOR3 (N18940, N18934, N13971, N7122);
nor NOR4 (N18941, N18924, N17728, N9890, N3253);
buf BUF1 (N18942, N18939);
nor NOR2 (N18943, N18940, N11577);
nor NOR2 (N18944, N18941, N8670);
buf BUF1 (N18945, N18937);
and AND2 (N18946, N18945, N13789);
nor NOR2 (N18947, N18942, N11593);
buf BUF1 (N18948, N18922);
not NOT1 (N18949, N18933);
or OR4 (N18950, N18948, N15474, N16815, N12105);
and AND2 (N18951, N18935, N18634);
not NOT1 (N18952, N18947);
and AND4 (N18953, N18930, N4323, N1056, N17082);
nand NAND3 (N18954, N18938, N14712, N6764);
buf BUF1 (N18955, N18951);
nor NOR4 (N18956, N18944, N4182, N18287, N6522);
buf BUF1 (N18957, N18956);
or OR3 (N18958, N18954, N5936, N4021);
nand NAND3 (N18959, N18953, N13752, N7343);
nor NOR4 (N18960, N18955, N16960, N3459, N8630);
nor NOR3 (N18961, N18952, N14368, N15852);
not NOT1 (N18962, N18961);
and AND2 (N18963, N18943, N3345);
and AND2 (N18964, N18958, N14833);
nor NOR4 (N18965, N18964, N10882, N5717, N3865);
nor NOR3 (N18966, N18946, N6663, N13653);
or OR4 (N18967, N18949, N7878, N16547, N16800);
not NOT1 (N18968, N18926);
buf BUF1 (N18969, N18967);
and AND3 (N18970, N18963, N4707, N5441);
nor NOR2 (N18971, N18962, N204);
nand NAND4 (N18972, N18957, N5197, N9866, N16955);
buf BUF1 (N18973, N18959);
nand NAND4 (N18974, N18968, N3079, N12110, N4637);
nand NAND2 (N18975, N18972, N9834);
buf BUF1 (N18976, N18974);
and AND3 (N18977, N18969, N1482, N4500);
or OR4 (N18978, N18975, N13931, N15475, N11328);
or OR4 (N18979, N18965, N3334, N15327, N14125);
nor NOR3 (N18980, N18976, N11543, N13085);
buf BUF1 (N18981, N18971);
not NOT1 (N18982, N18980);
nor NOR4 (N18983, N18982, N13758, N8707, N8698);
xor XOR2 (N18984, N18960, N1847);
nor NOR3 (N18985, N18977, N8486, N16995);
xor XOR2 (N18986, N18973, N15973);
xor XOR2 (N18987, N18983, N984);
not NOT1 (N18988, N18985);
buf BUF1 (N18989, N18981);
buf BUF1 (N18990, N18950);
nand NAND3 (N18991, N18966, N10835, N2141);
xor XOR2 (N18992, N18970, N2892);
or OR2 (N18993, N18992, N14065);
or OR3 (N18994, N18986, N15271, N4232);
buf BUF1 (N18995, N18989);
xor XOR2 (N18996, N18984, N1119);
buf BUF1 (N18997, N18991);
or OR2 (N18998, N18997, N15428);
buf BUF1 (N18999, N18993);
or OR2 (N19000, N18979, N1242);
not NOT1 (N19001, N18999);
buf BUF1 (N19002, N18998);
xor XOR2 (N19003, N19000, N1037);
nand NAND3 (N19004, N18987, N6536, N16366);
xor XOR2 (N19005, N19004, N17078);
buf BUF1 (N19006, N18990);
or OR4 (N19007, N19006, N10684, N1972, N4837);
buf BUF1 (N19008, N18988);
and AND2 (N19009, N18996, N12032);
nor NOR3 (N19010, N19008, N1893, N3670);
or OR4 (N19011, N18978, N4548, N5040, N18265);
and AND3 (N19012, N19005, N9980, N15403);
buf BUF1 (N19013, N19001);
xor XOR2 (N19014, N19002, N10846);
not NOT1 (N19015, N18995);
not NOT1 (N19016, N19011);
nand NAND4 (N19017, N19010, N7521, N4750, N10304);
nand NAND4 (N19018, N19009, N7031, N13909, N17829);
or OR3 (N19019, N19018, N9450, N10850);
buf BUF1 (N19020, N19017);
or OR4 (N19021, N18994, N16694, N9505, N17057);
or OR4 (N19022, N19021, N9744, N10734, N14542);
nor NOR2 (N19023, N19020, N14663);
buf BUF1 (N19024, N19014);
not NOT1 (N19025, N19016);
xor XOR2 (N19026, N19013, N7960);
and AND2 (N19027, N19012, N82);
nor NOR3 (N19028, N19024, N15098, N6517);
buf BUF1 (N19029, N19023);
or OR2 (N19030, N19015, N6369);
nor NOR4 (N19031, N19027, N13226, N18357, N17430);
nor NOR4 (N19032, N19026, N17330, N1184, N9931);
buf BUF1 (N19033, N19030);
buf BUF1 (N19034, N19028);
not NOT1 (N19035, N19022);
not NOT1 (N19036, N19034);
not NOT1 (N19037, N19025);
buf BUF1 (N19038, N19003);
or OR4 (N19039, N19031, N11295, N17074, N13697);
and AND2 (N19040, N19036, N5859);
nor NOR3 (N19041, N19029, N13801, N18554);
nand NAND2 (N19042, N19019, N89);
nand NAND3 (N19043, N19040, N17787, N9064);
nand NAND4 (N19044, N19042, N1676, N7741, N122);
or OR2 (N19045, N19044, N15012);
and AND4 (N19046, N19037, N7300, N1967, N16314);
and AND2 (N19047, N19007, N8519);
or OR3 (N19048, N19039, N9959, N5919);
xor XOR2 (N19049, N19041, N9128);
buf BUF1 (N19050, N19038);
and AND2 (N19051, N19045, N1988);
or OR2 (N19052, N19035, N7268);
xor XOR2 (N19053, N19051, N16909);
not NOT1 (N19054, N19046);
nor NOR3 (N19055, N19050, N16711, N7569);
not NOT1 (N19056, N19032);
and AND4 (N19057, N19054, N16681, N3030, N4275);
buf BUF1 (N19058, N19049);
and AND2 (N19059, N19048, N17802);
not NOT1 (N19060, N19053);
xor XOR2 (N19061, N19052, N6903);
and AND4 (N19062, N19060, N11120, N14404, N4751);
xor XOR2 (N19063, N19033, N3437);
nor NOR4 (N19064, N19058, N251, N17179, N7207);
nand NAND3 (N19065, N19064, N4655, N8234);
not NOT1 (N19066, N19047);
and AND2 (N19067, N19063, N13847);
and AND4 (N19068, N19059, N17520, N14835, N9245);
xor XOR2 (N19069, N19068, N16166);
nor NOR4 (N19070, N19056, N2539, N3793, N5533);
nand NAND4 (N19071, N19067, N10668, N2178, N12258);
nor NOR2 (N19072, N19043, N16790);
buf BUF1 (N19073, N19061);
buf BUF1 (N19074, N19065);
xor XOR2 (N19075, N19074, N17137);
or OR4 (N19076, N19070, N18287, N9672, N15045);
buf BUF1 (N19077, N19062);
xor XOR2 (N19078, N19075, N17090);
not NOT1 (N19079, N19069);
xor XOR2 (N19080, N19073, N5789);
or OR3 (N19081, N19077, N4251, N59);
not NOT1 (N19082, N19066);
or OR3 (N19083, N19082, N18794, N6075);
and AND4 (N19084, N19079, N12991, N13507, N17478);
or OR2 (N19085, N19071, N8093);
xor XOR2 (N19086, N19078, N10884);
not NOT1 (N19087, N19072);
xor XOR2 (N19088, N19055, N4919);
and AND2 (N19089, N19057, N8182);
buf BUF1 (N19090, N19084);
xor XOR2 (N19091, N19085, N8191);
or OR3 (N19092, N19076, N8740, N2904);
and AND2 (N19093, N19081, N11808);
and AND3 (N19094, N19091, N17288, N13581);
nor NOR2 (N19095, N19094, N4198);
or OR4 (N19096, N19095, N12303, N6486, N13691);
or OR3 (N19097, N19092, N8220, N6225);
nor NOR4 (N19098, N19083, N1920, N506, N17823);
and AND2 (N19099, N19087, N8589);
nor NOR3 (N19100, N19097, N6538, N11049);
or OR3 (N19101, N19100, N18914, N6914);
not NOT1 (N19102, N19098);
not NOT1 (N19103, N19101);
or OR3 (N19104, N19080, N9536, N6117);
nor NOR4 (N19105, N19099, N9413, N3644, N15611);
nand NAND4 (N19106, N19103, N6348, N2563, N18875);
xor XOR2 (N19107, N19104, N18204);
nand NAND2 (N19108, N19102, N5691);
nor NOR4 (N19109, N19090, N5808, N17140, N11604);
or OR4 (N19110, N19088, N10367, N4022, N6525);
or OR4 (N19111, N19105, N3794, N3213, N11058);
xor XOR2 (N19112, N19110, N7780);
or OR2 (N19113, N19111, N10830);
or OR2 (N19114, N19108, N220);
nand NAND2 (N19115, N19106, N15420);
not NOT1 (N19116, N19107);
xor XOR2 (N19117, N19114, N541);
nor NOR3 (N19118, N19117, N1956, N8891);
nand NAND4 (N19119, N19116, N4117, N8539, N4069);
buf BUF1 (N19120, N19096);
nor NOR4 (N19121, N19118, N8467, N11741, N6502);
nor NOR2 (N19122, N19120, N999);
xor XOR2 (N19123, N19113, N10482);
nor NOR2 (N19124, N19119, N7250);
and AND3 (N19125, N19122, N7223, N5323);
nor NOR4 (N19126, N19112, N5620, N857, N3196);
not NOT1 (N19127, N19125);
nor NOR3 (N19128, N19093, N2056, N9514);
or OR4 (N19129, N19089, N16002, N17654, N19062);
and AND3 (N19130, N19126, N1604, N2975);
and AND3 (N19131, N19124, N14105, N5542);
buf BUF1 (N19132, N19086);
buf BUF1 (N19133, N19131);
buf BUF1 (N19134, N19115);
and AND4 (N19135, N19128, N8952, N16905, N3960);
and AND2 (N19136, N19130, N16989);
buf BUF1 (N19137, N19121);
buf BUF1 (N19138, N19134);
and AND4 (N19139, N19135, N6120, N11783, N8835);
nor NOR3 (N19140, N19139, N15164, N12571);
buf BUF1 (N19141, N19123);
buf BUF1 (N19142, N19132);
and AND2 (N19143, N19138, N14738);
nor NOR4 (N19144, N19136, N1496, N17057, N7107);
and AND3 (N19145, N19140, N170, N16077);
nor NOR4 (N19146, N19142, N5101, N18964, N9792);
buf BUF1 (N19147, N19144);
and AND4 (N19148, N19127, N1391, N8942, N12664);
nand NAND4 (N19149, N19146, N11718, N7397, N6120);
or OR3 (N19150, N19129, N2263, N8473);
nor NOR3 (N19151, N19137, N18285, N16119);
or OR4 (N19152, N19151, N6815, N9746, N8996);
xor XOR2 (N19153, N19150, N10486);
and AND2 (N19154, N19133, N12180);
buf BUF1 (N19155, N19145);
nand NAND3 (N19156, N19141, N12189, N721);
and AND2 (N19157, N19143, N2845);
nor NOR3 (N19158, N19148, N1864, N7904);
and AND3 (N19159, N19155, N12355, N3786);
not NOT1 (N19160, N19152);
buf BUF1 (N19161, N19159);
xor XOR2 (N19162, N19156, N2318);
nand NAND2 (N19163, N19158, N17585);
xor XOR2 (N19164, N19161, N14331);
not NOT1 (N19165, N19154);
nor NOR3 (N19166, N19157, N13977, N14370);
xor XOR2 (N19167, N19166, N14761);
and AND3 (N19168, N19153, N4330, N18116);
buf BUF1 (N19169, N19165);
not NOT1 (N19170, N19163);
buf BUF1 (N19171, N19169);
or OR2 (N19172, N19162, N370);
buf BUF1 (N19173, N19109);
and AND2 (N19174, N19173, N1039);
and AND3 (N19175, N19168, N18680, N11612);
not NOT1 (N19176, N19164);
nand NAND3 (N19177, N19160, N48, N12817);
xor XOR2 (N19178, N19174, N18618);
or OR3 (N19179, N19167, N12303, N6073);
nor NOR4 (N19180, N19149, N4593, N17563, N11149);
not NOT1 (N19181, N19179);
buf BUF1 (N19182, N19147);
xor XOR2 (N19183, N19182, N13264);
and AND4 (N19184, N19176, N12792, N10246, N3062);
and AND2 (N19185, N19180, N3397);
nand NAND3 (N19186, N19184, N10653, N5277);
or OR2 (N19187, N19181, N9080);
nand NAND4 (N19188, N19175, N3291, N11981, N1149);
and AND3 (N19189, N19188, N6838, N19081);
buf BUF1 (N19190, N19170);
and AND3 (N19191, N19172, N14743, N1543);
and AND2 (N19192, N19189, N5555);
nand NAND4 (N19193, N19190, N4575, N12304, N4960);
and AND4 (N19194, N19171, N18339, N17903, N2164);
nand NAND2 (N19195, N19192, N9367);
nor NOR2 (N19196, N19191, N17324);
or OR3 (N19197, N19193, N204, N11896);
xor XOR2 (N19198, N19195, N17821);
xor XOR2 (N19199, N19186, N11062);
xor XOR2 (N19200, N19187, N18355);
not NOT1 (N19201, N19178);
xor XOR2 (N19202, N19185, N13877);
buf BUF1 (N19203, N19177);
xor XOR2 (N19204, N19183, N4342);
or OR3 (N19205, N19199, N18408, N18490);
buf BUF1 (N19206, N19194);
nand NAND3 (N19207, N19203, N16465, N18697);
nand NAND3 (N19208, N19206, N5050, N5219);
and AND3 (N19209, N19197, N17417, N13758);
not NOT1 (N19210, N19200);
not NOT1 (N19211, N19204);
or OR3 (N19212, N19196, N10552, N15483);
buf BUF1 (N19213, N19201);
or OR2 (N19214, N19198, N15757);
or OR3 (N19215, N19211, N15399, N16234);
or OR3 (N19216, N19202, N15380, N15563);
and AND4 (N19217, N19209, N1269, N10712, N11907);
nor NOR4 (N19218, N19214, N9675, N959, N5223);
or OR2 (N19219, N19212, N225);
nor NOR4 (N19220, N19208, N9941, N17327, N13428);
buf BUF1 (N19221, N19219);
xor XOR2 (N19222, N19216, N14511);
not NOT1 (N19223, N19213);
nor NOR3 (N19224, N19223, N10514, N2641);
or OR2 (N19225, N19215, N5619);
nor NOR3 (N19226, N19224, N4039, N17519);
nor NOR4 (N19227, N19226, N12572, N9882, N15505);
xor XOR2 (N19228, N19225, N19211);
or OR4 (N19229, N19205, N17500, N15382, N3070);
buf BUF1 (N19230, N19220);
nor NOR2 (N19231, N19207, N11971);
nor NOR4 (N19232, N19217, N10140, N969, N2774);
buf BUF1 (N19233, N19229);
buf BUF1 (N19234, N19228);
buf BUF1 (N19235, N19218);
not NOT1 (N19236, N19232);
xor XOR2 (N19237, N19236, N2384);
not NOT1 (N19238, N19235);
and AND4 (N19239, N19231, N1883, N12394, N17338);
or OR2 (N19240, N19221, N3503);
xor XOR2 (N19241, N19227, N643);
not NOT1 (N19242, N19230);
or OR4 (N19243, N19222, N11821, N11315, N10955);
xor XOR2 (N19244, N19237, N12843);
nand NAND2 (N19245, N19243, N9785);
xor XOR2 (N19246, N19238, N5365);
buf BUF1 (N19247, N19233);
nor NOR3 (N19248, N19239, N13020, N3416);
and AND4 (N19249, N19242, N8711, N16694, N9467);
nor NOR2 (N19250, N19247, N17392);
xor XOR2 (N19251, N19246, N132);
xor XOR2 (N19252, N19245, N13451);
not NOT1 (N19253, N19210);
xor XOR2 (N19254, N19241, N4029);
and AND3 (N19255, N19251, N18335, N6484);
nand NAND2 (N19256, N19254, N326);
xor XOR2 (N19257, N19248, N2234);
buf BUF1 (N19258, N19240);
xor XOR2 (N19259, N19249, N396);
nor NOR2 (N19260, N19259, N10491);
nand NAND3 (N19261, N19244, N8262, N14572);
and AND2 (N19262, N19260, N12650);
not NOT1 (N19263, N19262);
not NOT1 (N19264, N19263);
xor XOR2 (N19265, N19258, N18913);
and AND3 (N19266, N19257, N1737, N9625);
not NOT1 (N19267, N19252);
and AND2 (N19268, N19267, N1025);
xor XOR2 (N19269, N19265, N1504);
and AND4 (N19270, N19268, N96, N12767, N5815);
xor XOR2 (N19271, N19250, N5881);
xor XOR2 (N19272, N19261, N8798);
and AND4 (N19273, N19266, N17507, N10879, N871);
nor NOR2 (N19274, N19269, N15114);
buf BUF1 (N19275, N19272);
not NOT1 (N19276, N19253);
xor XOR2 (N19277, N19270, N18599);
or OR3 (N19278, N19274, N16928, N3147);
and AND4 (N19279, N19255, N18537, N12693, N12729);
nor NOR4 (N19280, N19277, N6154, N18542, N14976);
not NOT1 (N19281, N19256);
or OR3 (N19282, N19234, N14951, N17046);
nand NAND2 (N19283, N19273, N15590);
and AND2 (N19284, N19279, N1081);
buf BUF1 (N19285, N19271);
not NOT1 (N19286, N19285);
and AND4 (N19287, N19275, N2518, N1980, N855);
nand NAND4 (N19288, N19280, N10074, N14522, N754);
nor NOR4 (N19289, N19278, N12146, N15179, N12957);
buf BUF1 (N19290, N19288);
or OR3 (N19291, N19286, N6049, N3669);
nor NOR3 (N19292, N19289, N12739, N481);
nand NAND3 (N19293, N19264, N16912, N16362);
or OR3 (N19294, N19276, N18597, N18063);
or OR2 (N19295, N19291, N7487);
not NOT1 (N19296, N19287);
xor XOR2 (N19297, N19292, N932);
nor NOR2 (N19298, N19284, N6881);
xor XOR2 (N19299, N19298, N12388);
nand NAND2 (N19300, N19294, N211);
buf BUF1 (N19301, N19293);
and AND4 (N19302, N19301, N1979, N16731, N5871);
nand NAND2 (N19303, N19283, N15274);
or OR2 (N19304, N19290, N15149);
or OR2 (N19305, N19299, N18816);
and AND4 (N19306, N19282, N1239, N11858, N6254);
not NOT1 (N19307, N19306);
nor NOR3 (N19308, N19302, N5698, N13107);
buf BUF1 (N19309, N19297);
not NOT1 (N19310, N19303);
nand NAND4 (N19311, N19296, N8295, N7561, N1427);
not NOT1 (N19312, N19309);
nand NAND4 (N19313, N19281, N11541, N15775, N1536);
nand NAND2 (N19314, N19305, N630);
and AND2 (N19315, N19307, N3043);
and AND3 (N19316, N19308, N5854, N17146);
or OR2 (N19317, N19304, N13009);
nand NAND4 (N19318, N19310, N1044, N12283, N7678);
nor NOR2 (N19319, N19313, N63);
and AND2 (N19320, N19312, N10744);
buf BUF1 (N19321, N19300);
buf BUF1 (N19322, N19317);
buf BUF1 (N19323, N19318);
buf BUF1 (N19324, N19314);
xor XOR2 (N19325, N19321, N4048);
buf BUF1 (N19326, N19311);
nand NAND2 (N19327, N19323, N16288);
xor XOR2 (N19328, N19325, N445);
xor XOR2 (N19329, N19327, N3633);
nor NOR3 (N19330, N19329, N14113, N16102);
or OR3 (N19331, N19315, N6923, N13744);
buf BUF1 (N19332, N19326);
nand NAND3 (N19333, N19319, N3879, N4937);
or OR3 (N19334, N19322, N9756, N15533);
xor XOR2 (N19335, N19330, N4272);
nor NOR3 (N19336, N19332, N8584, N5876);
nand NAND4 (N19337, N19335, N515, N10749, N9007);
xor XOR2 (N19338, N19337, N15987);
and AND2 (N19339, N19334, N3580);
not NOT1 (N19340, N19295);
buf BUF1 (N19341, N19339);
buf BUF1 (N19342, N19336);
nand NAND3 (N19343, N19338, N13930, N7746);
and AND3 (N19344, N19316, N11982, N9104);
buf BUF1 (N19345, N19333);
not NOT1 (N19346, N19324);
nor NOR3 (N19347, N19331, N12006, N10658);
buf BUF1 (N19348, N19347);
not NOT1 (N19349, N19345);
nand NAND3 (N19350, N19341, N15485, N15225);
buf BUF1 (N19351, N19342);
xor XOR2 (N19352, N19320, N15117);
buf BUF1 (N19353, N19346);
and AND4 (N19354, N19352, N13372, N18565, N6335);
buf BUF1 (N19355, N19349);
and AND4 (N19356, N19343, N16389, N15113, N6198);
and AND4 (N19357, N19355, N6936, N14324, N1891);
nand NAND2 (N19358, N19353, N5940);
or OR2 (N19359, N19357, N4349);
or OR2 (N19360, N19356, N13388);
buf BUF1 (N19361, N19344);
nor NOR2 (N19362, N19340, N13944);
nand NAND4 (N19363, N19348, N17654, N18896, N16229);
buf BUF1 (N19364, N19328);
xor XOR2 (N19365, N19363, N13761);
or OR4 (N19366, N19364, N17348, N4204, N4295);
buf BUF1 (N19367, N19366);
nand NAND2 (N19368, N19354, N1780);
or OR3 (N19369, N19358, N16498, N9062);
or OR4 (N19370, N19367, N5104, N2345, N17993);
or OR3 (N19371, N19360, N15851, N16868);
and AND2 (N19372, N19371, N2715);
nor NOR3 (N19373, N19361, N18886, N1312);
buf BUF1 (N19374, N19350);
buf BUF1 (N19375, N19365);
or OR3 (N19376, N19372, N6651, N13750);
nor NOR3 (N19377, N19376, N16463, N15278);
and AND2 (N19378, N19374, N18133);
and AND4 (N19379, N19362, N4522, N4257, N7293);
and AND2 (N19380, N19378, N18979);
xor XOR2 (N19381, N19380, N14921);
and AND3 (N19382, N19381, N15840, N12993);
nand NAND2 (N19383, N19375, N6318);
nor NOR4 (N19384, N19382, N1888, N13314, N6152);
not NOT1 (N19385, N19384);
nand NAND3 (N19386, N19368, N6892, N17195);
nand NAND4 (N19387, N19386, N14665, N6024, N8654);
buf BUF1 (N19388, N19351);
xor XOR2 (N19389, N19369, N14607);
or OR4 (N19390, N19379, N9159, N10578, N10909);
or OR2 (N19391, N19377, N3495);
nor NOR2 (N19392, N19388, N17465);
nand NAND2 (N19393, N19385, N10718);
and AND2 (N19394, N19387, N17433);
xor XOR2 (N19395, N19390, N2157);
and AND4 (N19396, N19383, N11184, N12784, N11382);
not NOT1 (N19397, N19389);
nand NAND4 (N19398, N19373, N845, N5784, N14795);
not NOT1 (N19399, N19397);
nor NOR4 (N19400, N19396, N5605, N16477, N11344);
xor XOR2 (N19401, N19391, N17800);
xor XOR2 (N19402, N19392, N3390);
nand NAND2 (N19403, N19400, N11124);
and AND2 (N19404, N19399, N5822);
xor XOR2 (N19405, N19398, N10950);
and AND3 (N19406, N19402, N10102, N6131);
buf BUF1 (N19407, N19395);
or OR4 (N19408, N19407, N9041, N15589, N13881);
not NOT1 (N19409, N19408);
buf BUF1 (N19410, N19409);
and AND2 (N19411, N19393, N9935);
nor NOR2 (N19412, N19405, N18730);
buf BUF1 (N19413, N19370);
or OR4 (N19414, N19413, N5391, N9566, N8352);
buf BUF1 (N19415, N19414);
or OR4 (N19416, N19412, N8731, N18929, N11363);
and AND2 (N19417, N19411, N7305);
or OR2 (N19418, N19394, N7301);
and AND4 (N19419, N19416, N5111, N17971, N1737);
not NOT1 (N19420, N19410);
nand NAND2 (N19421, N19406, N9991);
nand NAND4 (N19422, N19403, N16490, N15040, N18415);
and AND4 (N19423, N19404, N9290, N656, N12360);
nand NAND2 (N19424, N19359, N11808);
buf BUF1 (N19425, N19415);
or OR2 (N19426, N19418, N16512);
and AND4 (N19427, N19419, N4040, N9100, N8384);
not NOT1 (N19428, N19425);
nand NAND3 (N19429, N19426, N11317, N7856);
nor NOR2 (N19430, N19420, N5421);
nand NAND2 (N19431, N19401, N11746);
not NOT1 (N19432, N19428);
nand NAND2 (N19433, N19417, N8415);
not NOT1 (N19434, N19432);
not NOT1 (N19435, N19422);
and AND2 (N19436, N19435, N6990);
or OR3 (N19437, N19424, N3992, N15124);
xor XOR2 (N19438, N19427, N8578);
xor XOR2 (N19439, N19437, N59);
not NOT1 (N19440, N19436);
nor NOR4 (N19441, N19423, N11362, N9616, N2003);
xor XOR2 (N19442, N19439, N11486);
nand NAND3 (N19443, N19429, N18813, N14062);
or OR2 (N19444, N19438, N18977);
nor NOR3 (N19445, N19441, N4598, N9344);
nor NOR4 (N19446, N19431, N833, N9305, N15527);
buf BUF1 (N19447, N19421);
buf BUF1 (N19448, N19446);
nor NOR2 (N19449, N19443, N11229);
nand NAND4 (N19450, N19440, N11290, N15762, N1241);
not NOT1 (N19451, N19447);
xor XOR2 (N19452, N19451, N17646);
not NOT1 (N19453, N19445);
not NOT1 (N19454, N19444);
nor NOR2 (N19455, N19448, N15594);
xor XOR2 (N19456, N19430, N10944);
and AND2 (N19457, N19454, N12271);
or OR2 (N19458, N19450, N14759);
nor NOR2 (N19459, N19453, N16411);
or OR3 (N19460, N19455, N5370, N6358);
not NOT1 (N19461, N19449);
nor NOR3 (N19462, N19460, N1248, N18424);
nand NAND2 (N19463, N19461, N15605);
not NOT1 (N19464, N19463);
nor NOR4 (N19465, N19458, N8719, N17894, N18527);
and AND2 (N19466, N19465, N5984);
not NOT1 (N19467, N19434);
not NOT1 (N19468, N19467);
xor XOR2 (N19469, N19442, N6725);
nor NOR2 (N19470, N19468, N9163);
and AND3 (N19471, N19462, N16967, N11641);
nand NAND2 (N19472, N19470, N3393);
nor NOR3 (N19473, N19471, N9909, N19428);
not NOT1 (N19474, N19466);
buf BUF1 (N19475, N19452);
or OR4 (N19476, N19459, N2656, N9158, N14121);
or OR2 (N19477, N19474, N7485);
not NOT1 (N19478, N19433);
nand NAND2 (N19479, N19476, N7558);
or OR2 (N19480, N19479, N14507);
nor NOR2 (N19481, N19472, N1214);
not NOT1 (N19482, N19473);
or OR2 (N19483, N19480, N8554);
not NOT1 (N19484, N19482);
xor XOR2 (N19485, N19469, N16495);
xor XOR2 (N19486, N19475, N18738);
not NOT1 (N19487, N19484);
buf BUF1 (N19488, N19477);
nand NAND4 (N19489, N19478, N11121, N3666, N10034);
and AND4 (N19490, N19487, N10776, N16286, N16000);
buf BUF1 (N19491, N19485);
or OR3 (N19492, N19486, N18012, N19103);
nor NOR2 (N19493, N19492, N7589);
xor XOR2 (N19494, N19456, N700);
or OR2 (N19495, N19489, N1480);
not NOT1 (N19496, N19457);
nor NOR3 (N19497, N19491, N4712, N15333);
or OR2 (N19498, N19481, N13181);
buf BUF1 (N19499, N19495);
and AND4 (N19500, N19496, N2736, N10812, N15692);
nand NAND4 (N19501, N19497, N5346, N15772, N10263);
or OR2 (N19502, N19464, N1187);
not NOT1 (N19503, N19490);
not NOT1 (N19504, N19494);
buf BUF1 (N19505, N19500);
and AND4 (N19506, N19503, N6540, N3303, N15076);
nor NOR3 (N19507, N19493, N6723, N10903);
xor XOR2 (N19508, N19506, N6678);
nor NOR3 (N19509, N19504, N7099, N19219);
xor XOR2 (N19510, N19483, N5604);
and AND4 (N19511, N19501, N18103, N9147, N13481);
or OR4 (N19512, N19505, N5031, N12988, N8360);
not NOT1 (N19513, N19512);
and AND4 (N19514, N19511, N15525, N12293, N6213);
nand NAND3 (N19515, N19510, N16355, N12956);
nand NAND2 (N19516, N19508, N17209);
and AND2 (N19517, N19502, N5223);
and AND4 (N19518, N19514, N4442, N4307, N482);
nor NOR2 (N19519, N19518, N17791);
buf BUF1 (N19520, N19513);
and AND2 (N19521, N19509, N15242);
buf BUF1 (N19522, N19507);
nand NAND4 (N19523, N19499, N11130, N14930, N5060);
nor NOR3 (N19524, N19517, N11207, N531);
buf BUF1 (N19525, N19523);
not NOT1 (N19526, N19516);
not NOT1 (N19527, N19498);
or OR3 (N19528, N19527, N19174, N7502);
or OR4 (N19529, N19515, N16998, N17517, N12526);
xor XOR2 (N19530, N19488, N15317);
nand NAND3 (N19531, N19519, N13806, N18416);
nor NOR2 (N19532, N19524, N9584);
xor XOR2 (N19533, N19532, N1189);
not NOT1 (N19534, N19530);
nand NAND3 (N19535, N19531, N7019, N4616);
and AND2 (N19536, N19529, N5703);
not NOT1 (N19537, N19520);
nand NAND2 (N19538, N19535, N18884);
not NOT1 (N19539, N19522);
xor XOR2 (N19540, N19537, N5706);
nor NOR4 (N19541, N19528, N9008, N15252, N3933);
xor XOR2 (N19542, N19536, N4570);
nor NOR3 (N19543, N19542, N9555, N8300);
and AND3 (N19544, N19541, N133, N8762);
nor NOR2 (N19545, N19526, N19457);
or OR2 (N19546, N19543, N16130);
xor XOR2 (N19547, N19540, N5906);
nor NOR4 (N19548, N19521, N14110, N18166, N6738);
nand NAND3 (N19549, N19545, N16311, N13733);
or OR2 (N19550, N19534, N13732);
buf BUF1 (N19551, N19549);
xor XOR2 (N19552, N19544, N18031);
nand NAND4 (N19553, N19548, N7318, N17654, N8161);
nor NOR2 (N19554, N19538, N1535);
xor XOR2 (N19555, N19554, N16556);
not NOT1 (N19556, N19551);
buf BUF1 (N19557, N19533);
not NOT1 (N19558, N19547);
xor XOR2 (N19559, N19555, N7959);
and AND3 (N19560, N19525, N4277, N11024);
nand NAND3 (N19561, N19560, N9057, N1056);
nand NAND3 (N19562, N19557, N18687, N17343);
nor NOR3 (N19563, N19546, N10514, N5426);
not NOT1 (N19564, N19561);
not NOT1 (N19565, N19559);
buf BUF1 (N19566, N19563);
and AND4 (N19567, N19562, N14741, N11017, N9737);
buf BUF1 (N19568, N19558);
nand NAND3 (N19569, N19568, N7881, N17039);
or OR2 (N19570, N19539, N15766);
nor NOR2 (N19571, N19570, N703);
or OR4 (N19572, N19564, N16605, N16047, N4141);
nor NOR4 (N19573, N19567, N18703, N362, N10010);
not NOT1 (N19574, N19573);
not NOT1 (N19575, N19550);
xor XOR2 (N19576, N19552, N8086);
not NOT1 (N19577, N19566);
buf BUF1 (N19578, N19569);
not NOT1 (N19579, N19565);
buf BUF1 (N19580, N19579);
nor NOR2 (N19581, N19571, N9229);
not NOT1 (N19582, N19577);
nand NAND3 (N19583, N19553, N5663, N16603);
xor XOR2 (N19584, N19574, N18466);
or OR2 (N19585, N19578, N2690);
nand NAND3 (N19586, N19556, N18868, N9510);
not NOT1 (N19587, N19576);
not NOT1 (N19588, N19586);
buf BUF1 (N19589, N19572);
buf BUF1 (N19590, N19582);
xor XOR2 (N19591, N19575, N3590);
nor NOR3 (N19592, N19585, N9322, N4298);
or OR2 (N19593, N19592, N9425);
nor NOR4 (N19594, N19593, N1467, N10823, N4273);
or OR4 (N19595, N19584, N3744, N10108, N13587);
and AND2 (N19596, N19595, N1056);
xor XOR2 (N19597, N19590, N2105);
nor NOR2 (N19598, N19588, N9872);
nand NAND4 (N19599, N19589, N10731, N8895, N18588);
xor XOR2 (N19600, N19587, N1849);
buf BUF1 (N19601, N19597);
xor XOR2 (N19602, N19594, N10753);
buf BUF1 (N19603, N19583);
nor NOR4 (N19604, N19598, N5073, N9512, N19351);
buf BUF1 (N19605, N19602);
or OR4 (N19606, N19580, N5744, N10366, N11210);
xor XOR2 (N19607, N19606, N10895);
nand NAND3 (N19608, N19603, N5485, N13158);
or OR2 (N19609, N19607, N12805);
not NOT1 (N19610, N19609);
nand NAND3 (N19611, N19599, N14866, N15203);
or OR3 (N19612, N19610, N828, N7409);
nor NOR2 (N19613, N19591, N1866);
or OR4 (N19614, N19604, N15512, N8736, N280);
not NOT1 (N19615, N19596);
and AND2 (N19616, N19601, N5865);
not NOT1 (N19617, N19614);
nor NOR4 (N19618, N19615, N14055, N5156, N18607);
or OR3 (N19619, N19618, N5820, N15169);
not NOT1 (N19620, N19617);
nor NOR2 (N19621, N19620, N9812);
buf BUF1 (N19622, N19621);
buf BUF1 (N19623, N19605);
xor XOR2 (N19624, N19611, N16076);
nor NOR2 (N19625, N19622, N4502);
not NOT1 (N19626, N19613);
nor NOR2 (N19627, N19619, N50);
xor XOR2 (N19628, N19624, N9625);
nand NAND2 (N19629, N19600, N19438);
or OR3 (N19630, N19616, N2004, N7981);
not NOT1 (N19631, N19581);
nand NAND3 (N19632, N19630, N10368, N12977);
buf BUF1 (N19633, N19631);
xor XOR2 (N19634, N19628, N16596);
nand NAND3 (N19635, N19625, N7918, N6576);
nor NOR2 (N19636, N19635, N16367);
or OR4 (N19637, N19608, N9643, N891, N12675);
buf BUF1 (N19638, N19629);
not NOT1 (N19639, N19627);
nand NAND4 (N19640, N19626, N3669, N14045, N7680);
nand NAND3 (N19641, N19632, N9197, N13141);
or OR4 (N19642, N19639, N13797, N378, N8020);
or OR2 (N19643, N19623, N12335);
nand NAND4 (N19644, N19634, N10444, N10559, N19476);
xor XOR2 (N19645, N19633, N6884);
nand NAND3 (N19646, N19642, N13903, N18455);
buf BUF1 (N19647, N19645);
not NOT1 (N19648, N19640);
or OR4 (N19649, N19648, N11875, N15264, N8524);
buf BUF1 (N19650, N19644);
nor NOR4 (N19651, N19636, N15333, N1203, N19553);
or OR3 (N19652, N19638, N7273, N10836);
nand NAND2 (N19653, N19643, N16554);
nand NAND4 (N19654, N19651, N15007, N11759, N1123);
xor XOR2 (N19655, N19650, N13881);
xor XOR2 (N19656, N19652, N6830);
not NOT1 (N19657, N19654);
nand NAND3 (N19658, N19641, N13753, N11776);
buf BUF1 (N19659, N19656);
nand NAND2 (N19660, N19646, N7461);
nor NOR3 (N19661, N19647, N10893, N9332);
and AND3 (N19662, N19661, N12414, N947);
buf BUF1 (N19663, N19658);
not NOT1 (N19664, N19657);
and AND4 (N19665, N19649, N17348, N11418, N5963);
nor NOR3 (N19666, N19662, N18511, N2024);
buf BUF1 (N19667, N19655);
buf BUF1 (N19668, N19653);
not NOT1 (N19669, N19664);
nand NAND3 (N19670, N19663, N18865, N11698);
buf BUF1 (N19671, N19670);
xor XOR2 (N19672, N19612, N3965);
nor NOR4 (N19673, N19665, N4706, N17957, N6000);
and AND2 (N19674, N19669, N10043);
nand NAND3 (N19675, N19659, N18453, N7854);
buf BUF1 (N19676, N19666);
nor NOR4 (N19677, N19671, N5822, N1806, N8452);
and AND2 (N19678, N19677, N339);
buf BUF1 (N19679, N19668);
or OR3 (N19680, N19637, N4982, N3794);
or OR3 (N19681, N19679, N3677, N4863);
nand NAND3 (N19682, N19681, N14453, N10583);
not NOT1 (N19683, N19675);
or OR2 (N19684, N19682, N1310);
buf BUF1 (N19685, N19667);
nor NOR4 (N19686, N19676, N8883, N17844, N5178);
or OR3 (N19687, N19684, N1618, N5402);
not NOT1 (N19688, N19673);
not NOT1 (N19689, N19672);
and AND4 (N19690, N19674, N15977, N8825, N12562);
and AND3 (N19691, N19685, N14401, N7900);
xor XOR2 (N19692, N19660, N11900);
xor XOR2 (N19693, N19678, N17135);
nor NOR3 (N19694, N19689, N17276, N4021);
xor XOR2 (N19695, N19693, N3723);
buf BUF1 (N19696, N19694);
not NOT1 (N19697, N19680);
buf BUF1 (N19698, N19691);
not NOT1 (N19699, N19695);
nor NOR2 (N19700, N19687, N6829);
or OR4 (N19701, N19692, N16752, N6071, N864);
and AND4 (N19702, N19688, N16897, N19405, N18931);
nor NOR3 (N19703, N19690, N8609, N15388);
not NOT1 (N19704, N19686);
and AND4 (N19705, N19704, N8535, N3004, N15487);
and AND3 (N19706, N19698, N5375, N7044);
buf BUF1 (N19707, N19701);
not NOT1 (N19708, N19700);
and AND4 (N19709, N19697, N4205, N19146, N9536);
and AND4 (N19710, N19708, N3671, N4231, N18682);
and AND2 (N19711, N19706, N19591);
nor NOR3 (N19712, N19703, N2786, N2794);
or OR2 (N19713, N19711, N2192);
nand NAND2 (N19714, N19713, N17879);
xor XOR2 (N19715, N19712, N14230);
or OR4 (N19716, N19705, N19565, N19327, N4936);
nand NAND2 (N19717, N19709, N5346);
nor NOR4 (N19718, N19702, N6381, N12583, N5064);
or OR3 (N19719, N19717, N11786, N543);
xor XOR2 (N19720, N19696, N4725);
buf BUF1 (N19721, N19683);
not NOT1 (N19722, N19715);
and AND4 (N19723, N19719, N16871, N19471, N11120);
nand NAND3 (N19724, N19722, N3129, N5797);
or OR4 (N19725, N19720, N7941, N13642, N16947);
nand NAND3 (N19726, N19716, N1986, N15660);
not NOT1 (N19727, N19710);
xor XOR2 (N19728, N19726, N8722);
not NOT1 (N19729, N19707);
and AND2 (N19730, N19723, N4642);
not NOT1 (N19731, N19729);
nand NAND2 (N19732, N19714, N5357);
and AND4 (N19733, N19721, N14998, N6233, N18286);
nand NAND2 (N19734, N19728, N6393);
buf BUF1 (N19735, N19732);
nand NAND2 (N19736, N19725, N9978);
not NOT1 (N19737, N19718);
buf BUF1 (N19738, N19734);
nor NOR3 (N19739, N19738, N515, N3107);
nand NAND2 (N19740, N19699, N2335);
nand NAND4 (N19741, N19731, N15129, N8656, N17394);
nor NOR3 (N19742, N19739, N4810, N9601);
nand NAND3 (N19743, N19735, N13959, N17534);
or OR2 (N19744, N19727, N836);
nor NOR3 (N19745, N19740, N6804, N3339);
nor NOR4 (N19746, N19744, N17907, N4210, N1419);
nor NOR2 (N19747, N19742, N2728);
or OR4 (N19748, N19747, N18477, N15769, N2648);
nand NAND3 (N19749, N19748, N5964, N3978);
and AND2 (N19750, N19743, N8520);
nor NOR3 (N19751, N19737, N16474, N9571);
or OR4 (N19752, N19724, N11680, N3149, N1834);
and AND2 (N19753, N19749, N15062);
buf BUF1 (N19754, N19745);
not NOT1 (N19755, N19754);
not NOT1 (N19756, N19733);
and AND3 (N19757, N19746, N3660, N12341);
or OR3 (N19758, N19741, N5308, N8874);
nand NAND2 (N19759, N19758, N14811);
not NOT1 (N19760, N19750);
or OR3 (N19761, N19751, N15336, N15396);
and AND2 (N19762, N19761, N14692);
nand NAND3 (N19763, N19736, N9188, N4019);
or OR2 (N19764, N19756, N8269);
xor XOR2 (N19765, N19759, N18952);
and AND4 (N19766, N19752, N10393, N5877, N9214);
nor NOR2 (N19767, N19753, N1811);
buf BUF1 (N19768, N19763);
and AND2 (N19769, N19767, N13751);
nand NAND3 (N19770, N19757, N2579, N15447);
not NOT1 (N19771, N19760);
not NOT1 (N19772, N19770);
nand NAND3 (N19773, N19772, N16506, N19027);
and AND2 (N19774, N19764, N9753);
nor NOR3 (N19775, N19769, N4388, N6898);
nor NOR2 (N19776, N19762, N7986);
buf BUF1 (N19777, N19755);
and AND4 (N19778, N19765, N8558, N6842, N15347);
and AND4 (N19779, N19775, N9348, N11611, N2705);
not NOT1 (N19780, N19777);
nand NAND2 (N19781, N19773, N4678);
and AND3 (N19782, N19771, N6859, N5106);
or OR3 (N19783, N19730, N2052, N1823);
buf BUF1 (N19784, N19782);
or OR2 (N19785, N19779, N17027);
or OR3 (N19786, N19774, N18594, N3599);
nand NAND4 (N19787, N19776, N15224, N11923, N2328);
or OR3 (N19788, N19778, N13303, N17579);
buf BUF1 (N19789, N19766);
not NOT1 (N19790, N19785);
xor XOR2 (N19791, N19790, N10884);
buf BUF1 (N19792, N19768);
not NOT1 (N19793, N19780);
or OR2 (N19794, N19781, N3533);
nor NOR2 (N19795, N19794, N7376);
nand NAND4 (N19796, N19783, N4626, N17671, N4019);
xor XOR2 (N19797, N19789, N8269);
and AND4 (N19798, N19792, N1162, N10924, N799);
xor XOR2 (N19799, N19788, N5659);
and AND2 (N19800, N19797, N1178);
and AND3 (N19801, N19786, N8669, N10234);
nor NOR3 (N19802, N19784, N17751, N6067);
nand NAND4 (N19803, N19793, N10587, N13762, N2482);
not NOT1 (N19804, N19802);
not NOT1 (N19805, N19801);
buf BUF1 (N19806, N19795);
not NOT1 (N19807, N19796);
xor XOR2 (N19808, N19803, N10847);
xor XOR2 (N19809, N19808, N215);
nand NAND3 (N19810, N19805, N13055, N16143);
nor NOR2 (N19811, N19799, N1267);
xor XOR2 (N19812, N19804, N16631);
and AND2 (N19813, N19812, N17774);
not NOT1 (N19814, N19806);
xor XOR2 (N19815, N19810, N10076);
xor XOR2 (N19816, N19798, N13488);
nand NAND3 (N19817, N19791, N767, N15579);
nor NOR3 (N19818, N19787, N35, N19329);
or OR4 (N19819, N19818, N3379, N9060, N7023);
nor NOR2 (N19820, N19819, N18432);
xor XOR2 (N19821, N19800, N18415);
nand NAND4 (N19822, N19821, N12014, N2278, N14409);
xor XOR2 (N19823, N19822, N16257);
or OR3 (N19824, N19815, N10813, N4298);
not NOT1 (N19825, N19824);
or OR4 (N19826, N19816, N12652, N12068, N6012);
nand NAND2 (N19827, N19817, N16845);
and AND4 (N19828, N19826, N11435, N19660, N7400);
or OR4 (N19829, N19820, N12199, N4424, N6148);
or OR2 (N19830, N19823, N11392);
and AND4 (N19831, N19809, N12640, N4004, N11869);
not NOT1 (N19832, N19811);
buf BUF1 (N19833, N19825);
and AND3 (N19834, N19813, N18153, N3370);
not NOT1 (N19835, N19830);
buf BUF1 (N19836, N19835);
and AND4 (N19837, N19807, N5771, N18680, N14090);
buf BUF1 (N19838, N19828);
xor XOR2 (N19839, N19827, N14124);
buf BUF1 (N19840, N19833);
not NOT1 (N19841, N19814);
or OR4 (N19842, N19836, N14160, N3611, N11764);
nand NAND3 (N19843, N19832, N2137, N8480);
buf BUF1 (N19844, N19829);
not NOT1 (N19845, N19841);
and AND4 (N19846, N19840, N2390, N2020, N13532);
and AND2 (N19847, N19844, N14254);
buf BUF1 (N19848, N19843);
xor XOR2 (N19849, N19847, N977);
nor NOR4 (N19850, N19846, N9295, N15590, N590);
nor NOR4 (N19851, N19837, N14819, N7167, N19594);
and AND3 (N19852, N19842, N927, N7713);
xor XOR2 (N19853, N19834, N7327);
or OR3 (N19854, N19839, N10043, N15130);
not NOT1 (N19855, N19848);
not NOT1 (N19856, N19851);
and AND2 (N19857, N19838, N15863);
or OR4 (N19858, N19850, N9826, N16888, N19010);
nand NAND2 (N19859, N19852, N6865);
not NOT1 (N19860, N19849);
nor NOR2 (N19861, N19831, N845);
and AND2 (N19862, N19858, N8566);
nor NOR4 (N19863, N19845, N13164, N3572, N17494);
nor NOR4 (N19864, N19857, N7279, N7470, N386);
nand NAND4 (N19865, N19853, N17589, N19282, N13491);
buf BUF1 (N19866, N19859);
xor XOR2 (N19867, N19856, N12819);
not NOT1 (N19868, N19867);
nor NOR3 (N19869, N19862, N13953, N14519);
nor NOR4 (N19870, N19869, N4949, N9806, N9472);
or OR3 (N19871, N19863, N11279, N5780);
nor NOR2 (N19872, N19855, N1207);
nor NOR4 (N19873, N19868, N3383, N14878, N6354);
nor NOR3 (N19874, N19865, N2578, N865);
not NOT1 (N19875, N19871);
nor NOR2 (N19876, N19870, N19223);
xor XOR2 (N19877, N19873, N14999);
buf BUF1 (N19878, N19877);
not NOT1 (N19879, N19864);
and AND2 (N19880, N19854, N17081);
and AND4 (N19881, N19875, N13150, N73, N16948);
xor XOR2 (N19882, N19878, N15481);
nand NAND2 (N19883, N19874, N8172);
nand NAND4 (N19884, N19861, N10821, N11495, N19307);
and AND4 (N19885, N19880, N9979, N11208, N7162);
nand NAND4 (N19886, N19884, N15958, N14927, N3609);
buf BUF1 (N19887, N19885);
not NOT1 (N19888, N19866);
nand NAND2 (N19889, N19860, N18585);
nand NAND4 (N19890, N19881, N11429, N4247, N7105);
nor NOR4 (N19891, N19876, N4022, N3114, N19808);
nor NOR2 (N19892, N19889, N9249);
buf BUF1 (N19893, N19883);
nor NOR3 (N19894, N19882, N3045, N12621);
xor XOR2 (N19895, N19887, N5006);
and AND2 (N19896, N19872, N2147);
nor NOR4 (N19897, N19893, N828, N4452, N19227);
not NOT1 (N19898, N19891);
nand NAND2 (N19899, N19888, N10219);
buf BUF1 (N19900, N19894);
nand NAND4 (N19901, N19897, N18267, N11885, N11876);
and AND3 (N19902, N19895, N10043, N2683);
nand NAND2 (N19903, N19879, N19400);
and AND2 (N19904, N19886, N3424);
xor XOR2 (N19905, N19902, N19497);
nand NAND3 (N19906, N19904, N8453, N6883);
xor XOR2 (N19907, N19890, N13348);
and AND2 (N19908, N19903, N1719);
xor XOR2 (N19909, N19905, N154);
buf BUF1 (N19910, N19898);
and AND2 (N19911, N19900, N8459);
nor NOR2 (N19912, N19911, N8924);
buf BUF1 (N19913, N19892);
nand NAND3 (N19914, N19913, N13403, N10723);
buf BUF1 (N19915, N19899);
or OR3 (N19916, N19906, N17321, N16060);
and AND3 (N19917, N19912, N13680, N2660);
buf BUF1 (N19918, N19907);
nor NOR3 (N19919, N19901, N14828, N5741);
xor XOR2 (N19920, N19919, N733);
xor XOR2 (N19921, N19920, N8497);
nor NOR2 (N19922, N19916, N18707);
xor XOR2 (N19923, N19915, N4316);
and AND4 (N19924, N19918, N18495, N18286, N19771);
buf BUF1 (N19925, N19910);
and AND3 (N19926, N19896, N4446, N17495);
nand NAND2 (N19927, N19922, N19599);
xor XOR2 (N19928, N19926, N19427);
nand NAND4 (N19929, N19914, N1590, N5840, N8539);
buf BUF1 (N19930, N19909);
nor NOR4 (N19931, N19930, N6385, N5110, N9921);
or OR2 (N19932, N19927, N3193);
xor XOR2 (N19933, N19917, N6077);
buf BUF1 (N19934, N19931);
xor XOR2 (N19935, N19932, N11166);
buf BUF1 (N19936, N19924);
and AND2 (N19937, N19925, N12515);
or OR2 (N19938, N19936, N3344);
xor XOR2 (N19939, N19928, N17976);
not NOT1 (N19940, N19938);
and AND3 (N19941, N19934, N16795, N19395);
buf BUF1 (N19942, N19929);
and AND3 (N19943, N19939, N10425, N14660);
nand NAND4 (N19944, N19937, N3415, N946, N5318);
buf BUF1 (N19945, N19923);
xor XOR2 (N19946, N19940, N17990);
and AND2 (N19947, N19942, N15965);
not NOT1 (N19948, N19933);
and AND2 (N19949, N19908, N9107);
buf BUF1 (N19950, N19949);
nand NAND2 (N19951, N19943, N6997);
or OR4 (N19952, N19944, N243, N539, N15994);
nand NAND3 (N19953, N19945, N14286, N3965);
nor NOR3 (N19954, N19946, N3737, N8642);
or OR2 (N19955, N19941, N12163);
not NOT1 (N19956, N19954);
or OR4 (N19957, N19935, N12007, N9913, N8955);
nor NOR4 (N19958, N19957, N9198, N16603, N13191);
nand NAND2 (N19959, N19950, N18918);
or OR3 (N19960, N19956, N18559, N9323);
nor NOR2 (N19961, N19955, N7439);
nor NOR3 (N19962, N19948, N18520, N10035);
or OR3 (N19963, N19958, N10711, N10346);
buf BUF1 (N19964, N19963);
and AND3 (N19965, N19962, N3115, N4934);
xor XOR2 (N19966, N19947, N1336);
nand NAND2 (N19967, N19953, N8135);
or OR4 (N19968, N19961, N1503, N14678, N19059);
or OR4 (N19969, N19967, N19140, N11547, N13465);
nor NOR4 (N19970, N19965, N15837, N2651, N2765);
nor NOR2 (N19971, N19960, N8972);
xor XOR2 (N19972, N19966, N19836);
and AND2 (N19973, N19972, N2338);
buf BUF1 (N19974, N19968);
and AND2 (N19975, N19951, N19375);
xor XOR2 (N19976, N19973, N13090);
or OR4 (N19977, N19974, N15615, N15677, N6165);
nor NOR3 (N19978, N19969, N16709, N19796);
or OR3 (N19979, N19977, N11423, N17365);
or OR4 (N19980, N19952, N12538, N7182, N16724);
xor XOR2 (N19981, N19959, N3371);
nor NOR3 (N19982, N19964, N14347, N14956);
or OR2 (N19983, N19980, N2196);
buf BUF1 (N19984, N19982);
nor NOR3 (N19985, N19975, N2337, N19186);
xor XOR2 (N19986, N19978, N11533);
nor NOR2 (N19987, N19976, N6328);
xor XOR2 (N19988, N19985, N2629);
and AND4 (N19989, N19979, N17304, N10215, N3804);
or OR3 (N19990, N19987, N53, N4200);
nor NOR4 (N19991, N19981, N18128, N16600, N248);
buf BUF1 (N19992, N19986);
not NOT1 (N19993, N19988);
nand NAND3 (N19994, N19993, N3691, N3628);
or OR4 (N19995, N19990, N18726, N11964, N16674);
or OR4 (N19996, N19994, N4443, N1512, N14022);
buf BUF1 (N19997, N19989);
nand NAND2 (N19998, N19996, N5435);
xor XOR2 (N19999, N19970, N13251);
not NOT1 (N20000, N19971);
not NOT1 (N20001, N19995);
nor NOR2 (N20002, N19997, N10202);
and AND4 (N20003, N19921, N9800, N1993, N17442);
or OR2 (N20004, N20000, N10855);
nor NOR4 (N20005, N19984, N18602, N679, N6499);
not NOT1 (N20006, N20003);
not NOT1 (N20007, N19998);
nand NAND3 (N20008, N20004, N8231, N4090);
nor NOR3 (N20009, N19991, N13099, N15636);
buf BUF1 (N20010, N20006);
not NOT1 (N20011, N20005);
and AND2 (N20012, N20002, N15638);
nor NOR2 (N20013, N20010, N11860);
nand NAND4 (N20014, N20013, N6410, N11590, N13142);
nor NOR2 (N20015, N20009, N11901);
buf BUF1 (N20016, N20001);
not NOT1 (N20017, N20011);
buf BUF1 (N20018, N20016);
and AND3 (N20019, N20012, N1743, N15114);
buf BUF1 (N20020, N20017);
buf BUF1 (N20021, N19999);
not NOT1 (N20022, N20021);
and AND4 (N20023, N20007, N18504, N11077, N5500);
and AND3 (N20024, N20018, N8307, N4772);
nand NAND4 (N20025, N19992, N14111, N14196, N15141);
or OR3 (N20026, N20023, N10935, N17998);
buf BUF1 (N20027, N20008);
nand NAND3 (N20028, N19983, N19978, N14294);
buf BUF1 (N20029, N20024);
or OR4 (N20030, N20029, N7963, N16303, N1927);
and AND2 (N20031, N20014, N4301);
buf BUF1 (N20032, N20019);
xor XOR2 (N20033, N20015, N1749);
nand NAND4 (N20034, N20028, N8227, N1253, N8045);
xor XOR2 (N20035, N20030, N17028);
xor XOR2 (N20036, N20022, N659);
or OR2 (N20037, N20026, N453);
nor NOR3 (N20038, N20035, N9883, N3808);
nor NOR2 (N20039, N20020, N8231);
buf BUF1 (N20040, N20038);
not NOT1 (N20041, N20032);
xor XOR2 (N20042, N20037, N13815);
and AND2 (N20043, N20039, N3670);
buf BUF1 (N20044, N20036);
or OR3 (N20045, N20044, N11311, N19697);
nand NAND4 (N20046, N20045, N13277, N15569, N2938);
nor NOR4 (N20047, N20040, N11053, N2008, N12718);
nand NAND3 (N20048, N20046, N17410, N12434);
xor XOR2 (N20049, N20027, N14163);
buf BUF1 (N20050, N20034);
xor XOR2 (N20051, N20033, N7735);
xor XOR2 (N20052, N20049, N4756);
not NOT1 (N20053, N20052);
xor XOR2 (N20054, N20047, N18849);
buf BUF1 (N20055, N20025);
xor XOR2 (N20056, N20051, N18182);
buf BUF1 (N20057, N20031);
nand NAND4 (N20058, N20053, N6092, N1929, N19316);
xor XOR2 (N20059, N20048, N16173);
buf BUF1 (N20060, N20050);
nor NOR4 (N20061, N20054, N15951, N2452, N10804);
not NOT1 (N20062, N20060);
not NOT1 (N20063, N20061);
nor NOR2 (N20064, N20041, N12074);
and AND4 (N20065, N20063, N6857, N17059, N66);
not NOT1 (N20066, N20065);
xor XOR2 (N20067, N20042, N11461);
buf BUF1 (N20068, N20067);
buf BUF1 (N20069, N20043);
nor NOR3 (N20070, N20068, N15859, N14092);
or OR2 (N20071, N20058, N18164);
xor XOR2 (N20072, N20071, N2838);
or OR2 (N20073, N20072, N4469);
and AND2 (N20074, N20055, N1783);
and AND4 (N20075, N20070, N2576, N250, N17486);
not NOT1 (N20076, N20069);
nor NOR3 (N20077, N20066, N18606, N15337);
or OR2 (N20078, N20077, N3087);
not NOT1 (N20079, N20078);
and AND2 (N20080, N20062, N7762);
buf BUF1 (N20081, N20057);
nand NAND3 (N20082, N20073, N8819, N19015);
nand NAND2 (N20083, N20081, N1961);
or OR4 (N20084, N20074, N1646, N9139, N6543);
and AND3 (N20085, N20076, N13615, N427);
nand NAND3 (N20086, N20059, N19133, N7081);
nor NOR2 (N20087, N20064, N12334);
and AND4 (N20088, N20083, N10534, N8425, N17464);
or OR4 (N20089, N20082, N16253, N5700, N15692);
and AND4 (N20090, N20088, N10371, N4095, N5110);
not NOT1 (N20091, N20080);
nor NOR4 (N20092, N20085, N7872, N13920, N16448);
and AND4 (N20093, N20091, N17810, N10190, N6204);
and AND4 (N20094, N20056, N1309, N19011, N7712);
nor NOR2 (N20095, N20079, N4535);
xor XOR2 (N20096, N20087, N6387);
nor NOR3 (N20097, N20089, N12406, N16680);
nand NAND3 (N20098, N20086, N10531, N9345);
not NOT1 (N20099, N20095);
not NOT1 (N20100, N20084);
nand NAND4 (N20101, N20100, N17125, N19996, N9185);
nand NAND3 (N20102, N20097, N4465, N916);
nand NAND3 (N20103, N20102, N6087, N10206);
not NOT1 (N20104, N20098);
and AND3 (N20105, N20103, N14583, N7869);
nand NAND4 (N20106, N20105, N9984, N9846, N7352);
not NOT1 (N20107, N20099);
and AND3 (N20108, N20107, N3175, N47);
and AND3 (N20109, N20096, N5571, N11931);
or OR3 (N20110, N20075, N104, N3392);
not NOT1 (N20111, N20106);
and AND3 (N20112, N20108, N17426, N731);
nor NOR2 (N20113, N20090, N8273);
xor XOR2 (N20114, N20094, N12974);
nand NAND4 (N20115, N20113, N9560, N1862, N1709);
or OR4 (N20116, N20092, N15123, N3833, N13700);
not NOT1 (N20117, N20101);
and AND4 (N20118, N20116, N5113, N15135, N1197);
buf BUF1 (N20119, N20114);
not NOT1 (N20120, N20112);
buf BUF1 (N20121, N20093);
nor NOR3 (N20122, N20115, N14896, N1923);
xor XOR2 (N20123, N20111, N17083);
nand NAND4 (N20124, N20122, N8049, N1436, N16119);
buf BUF1 (N20125, N20110);
nor NOR2 (N20126, N20117, N17757);
nand NAND4 (N20127, N20126, N10085, N4455, N13116);
and AND2 (N20128, N20124, N12161);
nand NAND4 (N20129, N20125, N13793, N7857, N7744);
xor XOR2 (N20130, N20128, N12659);
nor NOR2 (N20131, N20130, N8792);
or OR4 (N20132, N20121, N16406, N11965, N9304);
not NOT1 (N20133, N20120);
buf BUF1 (N20134, N20119);
buf BUF1 (N20135, N20104);
xor XOR2 (N20136, N20118, N10922);
or OR2 (N20137, N20129, N15227);
buf BUF1 (N20138, N20109);
xor XOR2 (N20139, N20132, N12346);
and AND2 (N20140, N20123, N11889);
nor NOR3 (N20141, N20133, N5317, N7711);
nand NAND2 (N20142, N20139, N5351);
nor NOR3 (N20143, N20142, N6086, N15152);
and AND3 (N20144, N20131, N10174, N4721);
nand NAND4 (N20145, N20135, N17446, N18105, N13265);
nor NOR2 (N20146, N20145, N14218);
buf BUF1 (N20147, N20138);
and AND3 (N20148, N20147, N4563, N14944);
nand NAND4 (N20149, N20141, N6669, N1224, N5072);
nor NOR3 (N20150, N20144, N10953, N8888);
buf BUF1 (N20151, N20140);
nor NOR4 (N20152, N20137, N18502, N13956, N15832);
not NOT1 (N20153, N20149);
xor XOR2 (N20154, N20148, N14341);
or OR3 (N20155, N20127, N227, N18730);
buf BUF1 (N20156, N20146);
xor XOR2 (N20157, N20154, N17563);
nor NOR3 (N20158, N20155, N16061, N14596);
buf BUF1 (N20159, N20134);
or OR3 (N20160, N20153, N18723, N5231);
buf BUF1 (N20161, N20158);
not NOT1 (N20162, N20156);
and AND2 (N20163, N20136, N5623);
nand NAND4 (N20164, N20157, N3402, N16083, N9202);
nor NOR3 (N20165, N20143, N5262, N8134);
and AND4 (N20166, N20159, N16892, N9465, N4651);
or OR4 (N20167, N20163, N60, N8247, N3026);
nor NOR2 (N20168, N20164, N7084);
nor NOR4 (N20169, N20166, N3207, N5094, N15243);
and AND4 (N20170, N20161, N7481, N16220, N16553);
nand NAND2 (N20171, N20152, N12356);
buf BUF1 (N20172, N20160);
or OR4 (N20173, N20150, N3800, N4458, N4230);
not NOT1 (N20174, N20170);
xor XOR2 (N20175, N20172, N12143);
nor NOR4 (N20176, N20173, N11364, N6475, N6716);
not NOT1 (N20177, N20165);
buf BUF1 (N20178, N20175);
nor NOR2 (N20179, N20177, N17779);
not NOT1 (N20180, N20176);
buf BUF1 (N20181, N20171);
buf BUF1 (N20182, N20167);
nor NOR3 (N20183, N20169, N905, N14692);
not NOT1 (N20184, N20182);
xor XOR2 (N20185, N20181, N19094);
buf BUF1 (N20186, N20185);
buf BUF1 (N20187, N20179);
nand NAND2 (N20188, N20162, N17477);
xor XOR2 (N20189, N20178, N13169);
nor NOR4 (N20190, N20186, N17602, N13702, N9347);
xor XOR2 (N20191, N20174, N5374);
xor XOR2 (N20192, N20189, N12307);
and AND2 (N20193, N20191, N10496);
nand NAND4 (N20194, N20183, N10765, N8544, N5919);
or OR2 (N20195, N20180, N14671);
xor XOR2 (N20196, N20151, N16648);
xor XOR2 (N20197, N20193, N15920);
nor NOR2 (N20198, N20184, N19963);
or OR2 (N20199, N20192, N8668);
nor NOR2 (N20200, N20195, N17929);
not NOT1 (N20201, N20199);
or OR4 (N20202, N20196, N5661, N846, N10059);
buf BUF1 (N20203, N20202);
nand NAND2 (N20204, N20198, N9099);
or OR4 (N20205, N20187, N2725, N12143, N7334);
nor NOR3 (N20206, N20205, N966, N17574);
nand NAND3 (N20207, N20203, N3643, N15696);
xor XOR2 (N20208, N20206, N15896);
not NOT1 (N20209, N20207);
not NOT1 (N20210, N20188);
not NOT1 (N20211, N20210);
xor XOR2 (N20212, N20208, N14298);
not NOT1 (N20213, N20209);
nor NOR4 (N20214, N20213, N7195, N3423, N17897);
xor XOR2 (N20215, N20194, N13614);
nand NAND3 (N20216, N20204, N2946, N16252);
nor NOR3 (N20217, N20216, N3484, N19292);
nand NAND2 (N20218, N20212, N9990);
and AND2 (N20219, N20215, N13257);
nor NOR4 (N20220, N20214, N14056, N2360, N8469);
buf BUF1 (N20221, N20217);
and AND4 (N20222, N20221, N13155, N15517, N3795);
nor NOR4 (N20223, N20200, N6334, N1840, N13484);
and AND3 (N20224, N20168, N11265, N10614);
nand NAND3 (N20225, N20201, N1222, N9228);
nor NOR2 (N20226, N20190, N19955);
nor NOR2 (N20227, N20219, N6051);
and AND3 (N20228, N20220, N16155, N16744);
xor XOR2 (N20229, N20224, N10342);
or OR2 (N20230, N20229, N1011);
and AND2 (N20231, N20222, N11024);
nand NAND4 (N20232, N20226, N18530, N9392, N3137);
nand NAND4 (N20233, N20227, N19091, N18773, N3440);
nor NOR2 (N20234, N20233, N15553);
or OR3 (N20235, N20234, N13909, N12597);
buf BUF1 (N20236, N20211);
not NOT1 (N20237, N20232);
nor NOR3 (N20238, N20237, N18143, N2570);
nor NOR2 (N20239, N20223, N10135);
and AND3 (N20240, N20197, N7238, N738);
nand NAND4 (N20241, N20225, N7213, N19460, N18572);
and AND2 (N20242, N20240, N11251);
or OR3 (N20243, N20235, N8976, N3533);
nor NOR2 (N20244, N20238, N3723);
xor XOR2 (N20245, N20231, N1899);
xor XOR2 (N20246, N20236, N2453);
and AND4 (N20247, N20218, N12449, N10439, N12684);
and AND3 (N20248, N20239, N18165, N10267);
xor XOR2 (N20249, N20248, N13430);
not NOT1 (N20250, N20245);
xor XOR2 (N20251, N20241, N12265);
buf BUF1 (N20252, N20250);
nor NOR2 (N20253, N20230, N3318);
and AND2 (N20254, N20249, N2168);
nand NAND4 (N20255, N20254, N18901, N14176, N13997);
not NOT1 (N20256, N20252);
nand NAND3 (N20257, N20228, N3105, N20204);
buf BUF1 (N20258, N20253);
and AND4 (N20259, N20247, N964, N11039, N8291);
nand NAND3 (N20260, N20258, N17405, N12277);
nor NOR4 (N20261, N20256, N17648, N11560, N12740);
buf BUF1 (N20262, N20260);
nor NOR3 (N20263, N20251, N18738, N4206);
buf BUF1 (N20264, N20246);
buf BUF1 (N20265, N20243);
and AND2 (N20266, N20255, N5351);
nor NOR2 (N20267, N20261, N15436);
nand NAND2 (N20268, N20263, N4944);
xor XOR2 (N20269, N20266, N229);
nand NAND4 (N20270, N20268, N12971, N13072, N14002);
and AND3 (N20271, N20265, N10425, N2561);
nand NAND3 (N20272, N20267, N12063, N2526);
not NOT1 (N20273, N20269);
xor XOR2 (N20274, N20259, N1156);
xor XOR2 (N20275, N20264, N1257);
buf BUF1 (N20276, N20242);
nand NAND4 (N20277, N20262, N16735, N2603, N12150);
nand NAND3 (N20278, N20257, N15330, N6865);
nand NAND2 (N20279, N20278, N8599);
not NOT1 (N20280, N20279);
nor NOR3 (N20281, N20272, N18586, N16852);
nor NOR4 (N20282, N20277, N8637, N18463, N17249);
buf BUF1 (N20283, N20275);
not NOT1 (N20284, N20281);
xor XOR2 (N20285, N20280, N2805);
not NOT1 (N20286, N20284);
and AND2 (N20287, N20274, N14241);
or OR3 (N20288, N20282, N6350, N14098);
and AND4 (N20289, N20276, N19053, N11052, N3628);
xor XOR2 (N20290, N20273, N16295);
and AND2 (N20291, N20286, N11781);
nor NOR4 (N20292, N20288, N7402, N4433, N17740);
or OR4 (N20293, N20244, N7805, N17445, N5492);
not NOT1 (N20294, N20283);
nor NOR4 (N20295, N20291, N13210, N19731, N11528);
or OR3 (N20296, N20270, N4192, N11951);
xor XOR2 (N20297, N20294, N12823);
buf BUF1 (N20298, N20287);
not NOT1 (N20299, N20296);
and AND4 (N20300, N20293, N19945, N1668, N19184);
nor NOR3 (N20301, N20289, N5915, N19923);
xor XOR2 (N20302, N20300, N12362);
nand NAND2 (N20303, N20299, N12657);
and AND2 (N20304, N20292, N15884);
not NOT1 (N20305, N20304);
nor NOR4 (N20306, N20285, N5479, N14056, N8454);
xor XOR2 (N20307, N20303, N15965);
nand NAND4 (N20308, N20307, N564, N10136, N5162);
or OR2 (N20309, N20301, N2912);
xor XOR2 (N20310, N20290, N16315);
nand NAND4 (N20311, N20295, N8920, N19989, N16126);
nand NAND2 (N20312, N20305, N3094);
nand NAND3 (N20313, N20309, N10720, N970);
xor XOR2 (N20314, N20306, N8193);
nor NOR4 (N20315, N20312, N420, N706, N11194);
not NOT1 (N20316, N20271);
or OR4 (N20317, N20298, N14421, N13982, N2250);
nor NOR4 (N20318, N20313, N18944, N4179, N13616);
not NOT1 (N20319, N20297);
and AND3 (N20320, N20314, N13758, N187);
not NOT1 (N20321, N20311);
nand NAND4 (N20322, N20310, N5923, N14163, N11566);
nand NAND3 (N20323, N20318, N8037, N10552);
nor NOR3 (N20324, N20308, N8924, N13798);
nand NAND3 (N20325, N20322, N3159, N14527);
buf BUF1 (N20326, N20315);
not NOT1 (N20327, N20323);
or OR2 (N20328, N20324, N20316);
nor NOR2 (N20329, N6765, N3581);
not NOT1 (N20330, N20319);
and AND2 (N20331, N20327, N16145);
not NOT1 (N20332, N20326);
not NOT1 (N20333, N20330);
not NOT1 (N20334, N20333);
xor XOR2 (N20335, N20302, N5867);
and AND3 (N20336, N20320, N20088, N12758);
buf BUF1 (N20337, N20331);
xor XOR2 (N20338, N20325, N2706);
buf BUF1 (N20339, N20337);
nand NAND4 (N20340, N20317, N13006, N2489, N12692);
nor NOR3 (N20341, N20328, N10310, N7176);
xor XOR2 (N20342, N20339, N12458);
xor XOR2 (N20343, N20338, N14387);
or OR2 (N20344, N20329, N6772);
nand NAND2 (N20345, N20343, N19368);
and AND4 (N20346, N20342, N17135, N11739, N565);
xor XOR2 (N20347, N20334, N9510);
not NOT1 (N20348, N20336);
xor XOR2 (N20349, N20340, N15319);
and AND3 (N20350, N20346, N18780, N9809);
xor XOR2 (N20351, N20347, N19761);
nor NOR2 (N20352, N20350, N6497);
buf BUF1 (N20353, N20344);
xor XOR2 (N20354, N20321, N7367);
nand NAND4 (N20355, N20341, N6904, N13106, N10285);
not NOT1 (N20356, N20345);
xor XOR2 (N20357, N20349, N11311);
nand NAND2 (N20358, N20352, N18847);
and AND2 (N20359, N20354, N7792);
xor XOR2 (N20360, N20353, N18507);
not NOT1 (N20361, N20348);
and AND4 (N20362, N20335, N10793, N1854, N10015);
buf BUF1 (N20363, N20361);
nand NAND4 (N20364, N20358, N9217, N2393, N4546);
and AND2 (N20365, N20351, N13418);
not NOT1 (N20366, N20332);
nor NOR4 (N20367, N20363, N3993, N4099, N11672);
nor NOR3 (N20368, N20364, N11365, N5945);
xor XOR2 (N20369, N20357, N16503);
buf BUF1 (N20370, N20368);
nor NOR2 (N20371, N20367, N15447);
xor XOR2 (N20372, N20359, N15580);
or OR3 (N20373, N20372, N11296, N14818);
xor XOR2 (N20374, N20355, N18107);
and AND2 (N20375, N20356, N18883);
and AND2 (N20376, N20360, N18656);
and AND2 (N20377, N20370, N15178);
nand NAND2 (N20378, N20373, N2598);
xor XOR2 (N20379, N20369, N9100);
xor XOR2 (N20380, N20375, N16808);
nor NOR3 (N20381, N20377, N10256, N19881);
buf BUF1 (N20382, N20381);
nor NOR4 (N20383, N20380, N15947, N907, N5356);
buf BUF1 (N20384, N20362);
buf BUF1 (N20385, N20376);
nand NAND4 (N20386, N20365, N10565, N12083, N14428);
xor XOR2 (N20387, N20383, N17455);
nor NOR2 (N20388, N20379, N17873);
buf BUF1 (N20389, N20386);
or OR2 (N20390, N20388, N3504);
xor XOR2 (N20391, N20389, N4871);
or OR3 (N20392, N20385, N6146, N1748);
buf BUF1 (N20393, N20371);
not NOT1 (N20394, N20378);
xor XOR2 (N20395, N20384, N11151);
xor XOR2 (N20396, N20374, N14638);
nor NOR2 (N20397, N20387, N11458);
nor NOR2 (N20398, N20395, N7067);
nor NOR2 (N20399, N20391, N12657);
xor XOR2 (N20400, N20393, N5934);
nor NOR4 (N20401, N20390, N4205, N26, N8627);
and AND4 (N20402, N20366, N20072, N10532, N3262);
xor XOR2 (N20403, N20402, N2413);
buf BUF1 (N20404, N20392);
not NOT1 (N20405, N20401);
not NOT1 (N20406, N20394);
buf BUF1 (N20407, N20397);
or OR2 (N20408, N20407, N2103);
xor XOR2 (N20409, N20406, N3789);
xor XOR2 (N20410, N20405, N8866);
and AND2 (N20411, N20404, N18860);
xor XOR2 (N20412, N20408, N1978);
or OR2 (N20413, N20400, N775);
nor NOR2 (N20414, N20403, N19094);
buf BUF1 (N20415, N20396);
and AND4 (N20416, N20413, N16282, N7184, N15040);
buf BUF1 (N20417, N20414);
and AND4 (N20418, N20398, N665, N14666, N2510);
nand NAND3 (N20419, N20412, N10577, N19405);
not NOT1 (N20420, N20416);
nand NAND4 (N20421, N20415, N2350, N17367, N7541);
nand NAND2 (N20422, N20419, N7253);
nor NOR3 (N20423, N20418, N15531, N10655);
nor NOR2 (N20424, N20422, N10459);
and AND2 (N20425, N20409, N1455);
nor NOR2 (N20426, N20411, N13887);
xor XOR2 (N20427, N20382, N18180);
not NOT1 (N20428, N20427);
nand NAND3 (N20429, N20424, N1354, N13235);
xor XOR2 (N20430, N20429, N14665);
xor XOR2 (N20431, N20399, N7306);
buf BUF1 (N20432, N20426);
buf BUF1 (N20433, N20423);
buf BUF1 (N20434, N20420);
nor NOR2 (N20435, N20431, N4330);
not NOT1 (N20436, N20421);
nand NAND2 (N20437, N20433, N15844);
nor NOR4 (N20438, N20437, N17973, N15723, N14682);
nor NOR4 (N20439, N20436, N18410, N377, N3832);
xor XOR2 (N20440, N20439, N1345);
and AND4 (N20441, N20430, N16740, N14875, N4723);
xor XOR2 (N20442, N20425, N6498);
or OR4 (N20443, N20440, N828, N16198, N19343);
and AND2 (N20444, N20441, N3675);
nor NOR3 (N20445, N20428, N14753, N13396);
buf BUF1 (N20446, N20435);
buf BUF1 (N20447, N20417);
xor XOR2 (N20448, N20443, N64);
nand NAND3 (N20449, N20447, N10015, N2265);
and AND4 (N20450, N20444, N9517, N19509, N8730);
or OR4 (N20451, N20450, N8013, N6947, N9802);
not NOT1 (N20452, N20451);
buf BUF1 (N20453, N20410);
or OR2 (N20454, N20432, N18869);
buf BUF1 (N20455, N20446);
nand NAND3 (N20456, N20455, N7872, N17571);
nor NOR2 (N20457, N20438, N18860);
not NOT1 (N20458, N20453);
or OR3 (N20459, N20448, N5913, N8750);
and AND3 (N20460, N20459, N13221, N8232);
xor XOR2 (N20461, N20458, N6839);
xor XOR2 (N20462, N20445, N4644);
or OR4 (N20463, N20452, N3737, N16700, N16893);
and AND3 (N20464, N20460, N6239, N22);
nor NOR4 (N20465, N20461, N19139, N19122, N6152);
not NOT1 (N20466, N20442);
buf BUF1 (N20467, N20434);
nor NOR2 (N20468, N20467, N7984);
and AND2 (N20469, N20456, N5649);
or OR3 (N20470, N20464, N5412, N18827);
xor XOR2 (N20471, N20469, N2418);
not NOT1 (N20472, N20457);
nor NOR4 (N20473, N20470, N8768, N3828, N2623);
and AND2 (N20474, N20468, N14752);
not NOT1 (N20475, N20471);
or OR3 (N20476, N20462, N5773, N18585);
nand NAND4 (N20477, N20472, N265, N13444, N3976);
and AND3 (N20478, N20477, N17523, N3846);
nor NOR3 (N20479, N20466, N3569, N8364);
and AND4 (N20480, N20463, N20193, N1389, N6569);
buf BUF1 (N20481, N20475);
or OR4 (N20482, N20473, N10670, N3498, N16471);
nand NAND2 (N20483, N20482, N15985);
not NOT1 (N20484, N20480);
not NOT1 (N20485, N20474);
nand NAND3 (N20486, N20465, N11925, N7315);
buf BUF1 (N20487, N20478);
buf BUF1 (N20488, N20454);
nand NAND3 (N20489, N20485, N9919, N8912);
and AND2 (N20490, N20476, N7471);
not NOT1 (N20491, N20479);
or OR2 (N20492, N20481, N7442);
nor NOR3 (N20493, N20483, N7623, N6144);
nand NAND2 (N20494, N20490, N1722);
or OR3 (N20495, N20487, N2358, N9790);
or OR3 (N20496, N20449, N4887, N8639);
nand NAND2 (N20497, N20494, N16712);
and AND2 (N20498, N20496, N7041);
not NOT1 (N20499, N20492);
not NOT1 (N20500, N20488);
buf BUF1 (N20501, N20499);
not NOT1 (N20502, N20491);
xor XOR2 (N20503, N20502, N5205);
nand NAND3 (N20504, N20495, N3787, N15120);
xor XOR2 (N20505, N20504, N1669);
and AND4 (N20506, N20484, N16878, N3323, N13093);
buf BUF1 (N20507, N20486);
not NOT1 (N20508, N20506);
and AND4 (N20509, N20498, N9313, N8505, N16381);
and AND3 (N20510, N20501, N19837, N3287);
nand NAND2 (N20511, N20505, N5236);
buf BUF1 (N20512, N20511);
or OR3 (N20513, N20500, N7389, N12627);
not NOT1 (N20514, N20509);
buf BUF1 (N20515, N20510);
xor XOR2 (N20516, N20512, N11);
nor NOR4 (N20517, N20493, N7298, N3486, N17000);
nor NOR3 (N20518, N20497, N17636, N13659);
buf BUF1 (N20519, N20518);
not NOT1 (N20520, N20519);
or OR2 (N20521, N20507, N18095);
and AND2 (N20522, N20503, N925);
buf BUF1 (N20523, N20508);
and AND2 (N20524, N20520, N4654);
or OR2 (N20525, N20523, N3141);
xor XOR2 (N20526, N20514, N10138);
buf BUF1 (N20527, N20513);
xor XOR2 (N20528, N20517, N6765);
and AND4 (N20529, N20528, N9533, N13740, N3992);
nand NAND3 (N20530, N20525, N12085, N14141);
nor NOR2 (N20531, N20522, N10998);
xor XOR2 (N20532, N20526, N4508);
nand NAND4 (N20533, N20531, N17578, N15763, N9027);
buf BUF1 (N20534, N20529);
and AND4 (N20535, N20532, N18519, N11533, N9069);
nor NOR2 (N20536, N20527, N16564);
nor NOR3 (N20537, N20536, N7874, N9680);
buf BUF1 (N20538, N20489);
nor NOR2 (N20539, N20515, N15815);
nand NAND3 (N20540, N20533, N15804, N15300);
xor XOR2 (N20541, N20534, N14825);
not NOT1 (N20542, N20524);
buf BUF1 (N20543, N20541);
and AND2 (N20544, N20542, N16949);
xor XOR2 (N20545, N20544, N9644);
or OR4 (N20546, N20521, N10022, N5378, N11319);
and AND3 (N20547, N20538, N859, N18196);
nand NAND4 (N20548, N20539, N15656, N124, N19221);
nand NAND2 (N20549, N20516, N20044);
nor NOR4 (N20550, N20549, N19177, N4483, N8224);
nand NAND3 (N20551, N20546, N1625, N5898);
buf BUF1 (N20552, N20537);
or OR4 (N20553, N20547, N20115, N17954, N12907);
and AND2 (N20554, N20543, N17847);
and AND4 (N20555, N20554, N18942, N10117, N6786);
nor NOR3 (N20556, N20550, N17680, N6088);
not NOT1 (N20557, N20540);
xor XOR2 (N20558, N20545, N20126);
and AND3 (N20559, N20552, N10303, N8185);
xor XOR2 (N20560, N20551, N15116);
nor NOR3 (N20561, N20560, N9685, N9761);
nor NOR3 (N20562, N20556, N12940, N3087);
xor XOR2 (N20563, N20555, N19309);
and AND3 (N20564, N20530, N11799, N7756);
nor NOR2 (N20565, N20564, N9072);
and AND4 (N20566, N20562, N7979, N12378, N10582);
and AND3 (N20567, N20559, N5717, N9838);
nand NAND2 (N20568, N20561, N16789);
nor NOR3 (N20569, N20535, N10774, N4647);
nor NOR4 (N20570, N20558, N15991, N12232, N18656);
buf BUF1 (N20571, N20569);
and AND2 (N20572, N20566, N13013);
not NOT1 (N20573, N20567);
xor XOR2 (N20574, N20557, N4035);
and AND4 (N20575, N20568, N12905, N8707, N10690);
and AND2 (N20576, N20575, N6941);
not NOT1 (N20577, N20565);
nor NOR2 (N20578, N20573, N18695);
not NOT1 (N20579, N20572);
not NOT1 (N20580, N20570);
and AND3 (N20581, N20578, N16209, N18014);
and AND3 (N20582, N20553, N4596, N6630);
buf BUF1 (N20583, N20548);
nand NAND2 (N20584, N20576, N419);
or OR3 (N20585, N20581, N12144, N18703);
not NOT1 (N20586, N20579);
buf BUF1 (N20587, N20574);
and AND3 (N20588, N20585, N18090, N12628);
not NOT1 (N20589, N20580);
xor XOR2 (N20590, N20563, N3536);
and AND3 (N20591, N20577, N19917, N8478);
xor XOR2 (N20592, N20590, N2013);
or OR3 (N20593, N20589, N20132, N236);
or OR2 (N20594, N20582, N668);
xor XOR2 (N20595, N20583, N1815);
nor NOR4 (N20596, N20586, N18478, N16591, N18094);
nand NAND3 (N20597, N20596, N1324, N13454);
nand NAND2 (N20598, N20597, N18420);
and AND4 (N20599, N20592, N13448, N3993, N8188);
buf BUF1 (N20600, N20594);
xor XOR2 (N20601, N20598, N12187);
nand NAND3 (N20602, N20593, N3314, N19208);
or OR2 (N20603, N20601, N3159);
nand NAND3 (N20604, N20600, N14840, N3616);
buf BUF1 (N20605, N20588);
buf BUF1 (N20606, N20599);
nor NOR2 (N20607, N20606, N1095);
or OR3 (N20608, N20602, N525, N16520);
not NOT1 (N20609, N20605);
xor XOR2 (N20610, N20609, N11279);
buf BUF1 (N20611, N20587);
and AND4 (N20612, N20611, N1415, N12197, N8522);
or OR3 (N20613, N20610, N14754, N14535);
nor NOR4 (N20614, N20604, N12813, N17328, N14814);
buf BUF1 (N20615, N20591);
xor XOR2 (N20616, N20608, N8604);
nand NAND2 (N20617, N20616, N3045);
xor XOR2 (N20618, N20603, N3366);
nand NAND3 (N20619, N20584, N18771, N18620);
nor NOR3 (N20620, N20613, N11747, N4425);
and AND2 (N20621, N20620, N2993);
nand NAND3 (N20622, N20612, N14355, N13082);
nor NOR4 (N20623, N20571, N2976, N15880, N9491);
not NOT1 (N20624, N20595);
buf BUF1 (N20625, N20624);
not NOT1 (N20626, N20617);
or OR2 (N20627, N20619, N6106);
and AND3 (N20628, N20622, N16861, N6763);
not NOT1 (N20629, N20623);
and AND3 (N20630, N20626, N13863, N3264);
or OR3 (N20631, N20618, N14399, N10820);
not NOT1 (N20632, N20607);
nor NOR3 (N20633, N20631, N5304, N17245);
or OR4 (N20634, N20633, N4047, N11756, N16864);
nor NOR3 (N20635, N20627, N20054, N8991);
and AND2 (N20636, N20615, N1285);
and AND2 (N20637, N20625, N4915);
nor NOR4 (N20638, N20635, N15424, N16091, N5357);
nand NAND2 (N20639, N20628, N20145);
nor NOR2 (N20640, N20629, N1909);
nand NAND2 (N20641, N20632, N5327);
nand NAND2 (N20642, N20634, N4080);
not NOT1 (N20643, N20638);
nor NOR4 (N20644, N20621, N11726, N14202, N7052);
or OR3 (N20645, N20630, N14023, N13854);
not NOT1 (N20646, N20642);
nor NOR3 (N20647, N20640, N8440, N3162);
xor XOR2 (N20648, N20641, N10770);
not NOT1 (N20649, N20646);
or OR3 (N20650, N20639, N5033, N13316);
nor NOR3 (N20651, N20648, N7102, N13275);
or OR4 (N20652, N20644, N7109, N14372, N4385);
nand NAND3 (N20653, N20652, N12459, N2984);
nand NAND3 (N20654, N20647, N15791, N12718);
buf BUF1 (N20655, N20649);
buf BUF1 (N20656, N20653);
and AND3 (N20657, N20651, N19381, N15060);
not NOT1 (N20658, N20614);
buf BUF1 (N20659, N20655);
nor NOR4 (N20660, N20650, N19465, N18293, N4613);
nor NOR3 (N20661, N20658, N18855, N20096);
not NOT1 (N20662, N20654);
nor NOR4 (N20663, N20659, N4851, N12251, N1421);
and AND2 (N20664, N20637, N1322);
xor XOR2 (N20665, N20645, N2644);
and AND4 (N20666, N20662, N7054, N6324, N1658);
nand NAND3 (N20667, N20664, N4555, N9772);
and AND4 (N20668, N20666, N8989, N2902, N8525);
nand NAND3 (N20669, N20663, N3215, N1481);
nor NOR4 (N20670, N20668, N1738, N5442, N18034);
and AND2 (N20671, N20657, N20651);
and AND4 (N20672, N20665, N3578, N3988, N13456);
buf BUF1 (N20673, N20667);
and AND2 (N20674, N20671, N13965);
nand NAND3 (N20675, N20669, N2997, N18221);
buf BUF1 (N20676, N20670);
xor XOR2 (N20677, N20672, N6240);
not NOT1 (N20678, N20676);
nand NAND3 (N20679, N20678, N19344, N12862);
buf BUF1 (N20680, N20673);
and AND3 (N20681, N20636, N7850, N13574);
nor NOR2 (N20682, N20677, N15072);
nand NAND2 (N20683, N20661, N15822);
not NOT1 (N20684, N20681);
nor NOR4 (N20685, N20684, N17055, N12556, N17022);
nand NAND3 (N20686, N20656, N18181, N13708);
or OR4 (N20687, N20643, N9377, N19163, N10336);
nor NOR3 (N20688, N20660, N15315, N5630);
buf BUF1 (N20689, N20686);
buf BUF1 (N20690, N20682);
xor XOR2 (N20691, N20688, N355);
and AND2 (N20692, N20685, N12545);
nand NAND3 (N20693, N20674, N10196, N1781);
nand NAND3 (N20694, N20693, N6740, N8268);
or OR3 (N20695, N20689, N7122, N12303);
buf BUF1 (N20696, N20687);
nor NOR2 (N20697, N20694, N5536);
xor XOR2 (N20698, N20691, N11839);
buf BUF1 (N20699, N20683);
or OR2 (N20700, N20696, N2041);
nand NAND3 (N20701, N20699, N17828, N15308);
buf BUF1 (N20702, N20680);
not NOT1 (N20703, N20702);
or OR3 (N20704, N20697, N982, N10821);
nor NOR4 (N20705, N20690, N20303, N85, N10133);
or OR2 (N20706, N20692, N10026);
not NOT1 (N20707, N20700);
and AND2 (N20708, N20679, N11577);
buf BUF1 (N20709, N20706);
and AND3 (N20710, N20675, N8082, N14398);
buf BUF1 (N20711, N20703);
not NOT1 (N20712, N20695);
or OR4 (N20713, N20701, N13462, N15705, N9725);
buf BUF1 (N20714, N20710);
nor NOR2 (N20715, N20714, N5165);
nand NAND4 (N20716, N20698, N18679, N1192, N19656);
or OR3 (N20717, N20711, N13515, N5539);
not NOT1 (N20718, N20715);
nand NAND4 (N20719, N20708, N2385, N1503, N9800);
nand NAND4 (N20720, N20719, N5534, N8733, N20333);
nand NAND4 (N20721, N20707, N6528, N9013, N13407);
buf BUF1 (N20722, N20705);
or OR2 (N20723, N20716, N3164);
xor XOR2 (N20724, N20717, N13877);
not NOT1 (N20725, N20720);
xor XOR2 (N20726, N20718, N15384);
nor NOR2 (N20727, N20725, N4183);
and AND4 (N20728, N20724, N7300, N3680, N7566);
not NOT1 (N20729, N20728);
not NOT1 (N20730, N20704);
nor NOR2 (N20731, N20729, N650);
nor NOR3 (N20732, N20722, N13240, N13071);
xor XOR2 (N20733, N20713, N6379);
nor NOR4 (N20734, N20731, N1250, N17517, N11707);
nand NAND3 (N20735, N20733, N3040, N3957);
buf BUF1 (N20736, N20734);
nor NOR4 (N20737, N20721, N15159, N6857, N5819);
nor NOR2 (N20738, N20712, N1170);
buf BUF1 (N20739, N20730);
buf BUF1 (N20740, N20709);
nor NOR2 (N20741, N20727, N3806);
nor NOR4 (N20742, N20736, N7006, N6043, N9859);
buf BUF1 (N20743, N20738);
or OR3 (N20744, N20732, N9259, N7157);
or OR4 (N20745, N20735, N2609, N5702, N1817);
or OR4 (N20746, N20739, N14894, N15583, N20607);
nor NOR2 (N20747, N20742, N20347);
nand NAND3 (N20748, N20747, N15833, N16645);
and AND4 (N20749, N20746, N6711, N1652, N20441);
nand NAND3 (N20750, N20743, N5884, N18106);
and AND3 (N20751, N20749, N2226, N3243);
or OR3 (N20752, N20751, N16190, N14514);
xor XOR2 (N20753, N20752, N15814);
xor XOR2 (N20754, N20726, N17000);
or OR4 (N20755, N20744, N15939, N7339, N3815);
nor NOR4 (N20756, N20753, N135, N4323, N239);
or OR2 (N20757, N20745, N9585);
and AND3 (N20758, N20750, N5882, N8347);
nor NOR3 (N20759, N20757, N3665, N1941);
or OR4 (N20760, N20748, N14413, N7921, N17651);
nor NOR3 (N20761, N20754, N17364, N12953);
nor NOR2 (N20762, N20741, N7516);
or OR3 (N20763, N20755, N9227, N12729);
not NOT1 (N20764, N20758);
nand NAND3 (N20765, N20740, N11868, N326);
buf BUF1 (N20766, N20756);
nor NOR4 (N20767, N20764, N15997, N1952, N14105);
or OR4 (N20768, N20765, N10421, N18067, N7158);
nand NAND3 (N20769, N20768, N9196, N2974);
xor XOR2 (N20770, N20760, N18010);
not NOT1 (N20771, N20769);
not NOT1 (N20772, N20771);
or OR3 (N20773, N20766, N1182, N4758);
and AND3 (N20774, N20723, N17031, N8009);
or OR4 (N20775, N20774, N1531, N8004, N11541);
xor XOR2 (N20776, N20773, N18179);
nor NOR2 (N20777, N20775, N6399);
and AND2 (N20778, N20763, N1776);
nor NOR4 (N20779, N20759, N8943, N10082, N3700);
or OR3 (N20780, N20770, N20250, N285);
not NOT1 (N20781, N20778);
not NOT1 (N20782, N20767);
and AND4 (N20783, N20737, N16799, N10826, N451);
buf BUF1 (N20784, N20772);
not NOT1 (N20785, N20780);
nand NAND4 (N20786, N20776, N11425, N16327, N8847);
nand NAND2 (N20787, N20777, N6143);
not NOT1 (N20788, N20785);
or OR3 (N20789, N20781, N14979, N5251);
and AND2 (N20790, N20786, N18726);
nand NAND3 (N20791, N20782, N7513, N5716);
buf BUF1 (N20792, N20791);
or OR4 (N20793, N20792, N15946, N13266, N408);
and AND2 (N20794, N20789, N1886);
and AND3 (N20795, N20779, N7028, N9366);
nor NOR2 (N20796, N20790, N3051);
nor NOR3 (N20797, N20761, N8442, N4868);
not NOT1 (N20798, N20793);
xor XOR2 (N20799, N20798, N15750);
and AND2 (N20800, N20795, N2192);
xor XOR2 (N20801, N20787, N4202);
or OR3 (N20802, N20800, N14758, N11302);
buf BUF1 (N20803, N20788);
buf BUF1 (N20804, N20803);
nor NOR3 (N20805, N20784, N2482, N10642);
and AND3 (N20806, N20796, N11355, N10246);
not NOT1 (N20807, N20762);
not NOT1 (N20808, N20801);
nor NOR4 (N20809, N20808, N2075, N19926, N11373);
nand NAND3 (N20810, N20799, N6888, N9226);
nand NAND3 (N20811, N20804, N19351, N13594);
not NOT1 (N20812, N20794);
not NOT1 (N20813, N20806);
and AND3 (N20814, N20805, N2652, N10761);
nor NOR2 (N20815, N20807, N5538);
xor XOR2 (N20816, N20810, N18274);
buf BUF1 (N20817, N20802);
nand NAND4 (N20818, N20811, N17654, N9639, N5896);
not NOT1 (N20819, N20814);
or OR4 (N20820, N20813, N5845, N19246, N1680);
and AND2 (N20821, N20815, N24);
not NOT1 (N20822, N20809);
xor XOR2 (N20823, N20820, N14612);
and AND2 (N20824, N20797, N4990);
and AND3 (N20825, N20818, N12339, N15949);
and AND4 (N20826, N20822, N10484, N7042, N16566);
or OR2 (N20827, N20825, N10663);
nor NOR3 (N20828, N20824, N8264, N10439);
xor XOR2 (N20829, N20816, N13593);
nand NAND3 (N20830, N20829, N12869, N4912);
not NOT1 (N20831, N20817);
xor XOR2 (N20832, N20783, N221);
or OR2 (N20833, N20826, N12565);
xor XOR2 (N20834, N20827, N15993);
nor NOR4 (N20835, N20819, N17163, N15590, N2776);
not NOT1 (N20836, N20832);
xor XOR2 (N20837, N20812, N11731);
not NOT1 (N20838, N20833);
and AND2 (N20839, N20831, N7969);
xor XOR2 (N20840, N20830, N20141);
buf BUF1 (N20841, N20839);
nor NOR3 (N20842, N20837, N4186, N13624);
buf BUF1 (N20843, N20834);
not NOT1 (N20844, N20821);
xor XOR2 (N20845, N20836, N20363);
and AND2 (N20846, N20843, N10508);
buf BUF1 (N20847, N20845);
not NOT1 (N20848, N20844);
not NOT1 (N20849, N20840);
buf BUF1 (N20850, N20823);
nor NOR4 (N20851, N20842, N14865, N9217, N13046);
xor XOR2 (N20852, N20850, N4662);
buf BUF1 (N20853, N20846);
or OR4 (N20854, N20841, N8815, N11563, N17006);
and AND2 (N20855, N20847, N16032);
nand NAND4 (N20856, N20855, N20496, N13422, N20410);
xor XOR2 (N20857, N20835, N10823);
not NOT1 (N20858, N20848);
nor NOR4 (N20859, N20857, N459, N18435, N4010);
or OR3 (N20860, N20858, N17692, N2513);
nand NAND3 (N20861, N20849, N15589, N1615);
and AND3 (N20862, N20853, N2962, N3755);
buf BUF1 (N20863, N20861);
buf BUF1 (N20864, N20852);
or OR2 (N20865, N20859, N19412);
not NOT1 (N20866, N20856);
and AND4 (N20867, N20863, N1123, N3586, N15546);
nand NAND4 (N20868, N20864, N1152, N11306, N687);
nand NAND3 (N20869, N20860, N20617, N11798);
xor XOR2 (N20870, N20867, N7163);
or OR3 (N20871, N20851, N12620, N9120);
or OR3 (N20872, N20866, N11760, N19620);
or OR3 (N20873, N20838, N6064, N15114);
xor XOR2 (N20874, N20870, N5534);
nor NOR2 (N20875, N20868, N16310);
and AND4 (N20876, N20874, N9354, N6900, N18001);
not NOT1 (N20877, N20871);
and AND3 (N20878, N20876, N17988, N3116);
buf BUF1 (N20879, N20875);
xor XOR2 (N20880, N20869, N15088);
xor XOR2 (N20881, N20880, N9336);
buf BUF1 (N20882, N20873);
buf BUF1 (N20883, N20878);
or OR4 (N20884, N20883, N11633, N11210, N18676);
and AND4 (N20885, N20872, N6819, N12317, N19395);
or OR2 (N20886, N20884, N3818);
buf BUF1 (N20887, N20877);
or OR3 (N20888, N20862, N94, N788);
nand NAND4 (N20889, N20879, N15569, N8696, N1834);
nor NOR2 (N20890, N20865, N11706);
and AND2 (N20891, N20890, N14692);
nor NOR3 (N20892, N20854, N3700, N17642);
nand NAND3 (N20893, N20887, N14335, N9344);
buf BUF1 (N20894, N20828);
or OR2 (N20895, N20891, N476);
xor XOR2 (N20896, N20885, N19256);
nand NAND2 (N20897, N20882, N928);
nand NAND2 (N20898, N20897, N10834);
buf BUF1 (N20899, N20898);
not NOT1 (N20900, N20895);
nor NOR4 (N20901, N20900, N11544, N14853, N14858);
nor NOR2 (N20902, N20896, N15692);
nor NOR4 (N20903, N20899, N6640, N10602, N10327);
and AND4 (N20904, N20892, N3391, N10316, N3284);
not NOT1 (N20905, N20902);
not NOT1 (N20906, N20894);
nor NOR4 (N20907, N20903, N16967, N2296, N18423);
and AND2 (N20908, N20907, N5542);
and AND2 (N20909, N20893, N2694);
or OR4 (N20910, N20886, N20122, N17836, N11094);
not NOT1 (N20911, N20889);
or OR3 (N20912, N20888, N18164, N12828);
nor NOR4 (N20913, N20904, N9360, N12386, N12700);
nor NOR4 (N20914, N20908, N16810, N16964, N9258);
or OR4 (N20915, N20914, N10515, N6964, N5403);
xor XOR2 (N20916, N20906, N7757);
not NOT1 (N20917, N20909);
nand NAND3 (N20918, N20913, N7691, N914);
buf BUF1 (N20919, N20881);
not NOT1 (N20920, N20917);
nand NAND3 (N20921, N20918, N14793, N3855);
and AND2 (N20922, N20915, N20622);
xor XOR2 (N20923, N20911, N11956);
not NOT1 (N20924, N20916);
nand NAND3 (N20925, N20922, N16862, N18430);
and AND3 (N20926, N20924, N20247, N64);
nor NOR4 (N20927, N20912, N4150, N2703, N4892);
buf BUF1 (N20928, N20920);
buf BUF1 (N20929, N20919);
or OR3 (N20930, N20905, N18580, N6313);
and AND4 (N20931, N20925, N9866, N13710, N3089);
and AND3 (N20932, N20910, N14144, N13629);
buf BUF1 (N20933, N20929);
nor NOR4 (N20934, N20931, N3980, N16356, N10878);
not NOT1 (N20935, N20921);
not NOT1 (N20936, N20928);
not NOT1 (N20937, N20901);
not NOT1 (N20938, N20936);
and AND3 (N20939, N20938, N11782, N5382);
or OR2 (N20940, N20933, N8073);
buf BUF1 (N20941, N20937);
buf BUF1 (N20942, N20934);
and AND3 (N20943, N20926, N16779, N2777);
nor NOR3 (N20944, N20930, N12430, N3128);
nand NAND3 (N20945, N20932, N16080, N755);
and AND4 (N20946, N20943, N12128, N9805, N15328);
or OR2 (N20947, N20923, N14291);
or OR4 (N20948, N20941, N1203, N5572, N17545);
xor XOR2 (N20949, N20942, N2991);
xor XOR2 (N20950, N20949, N1927);
not NOT1 (N20951, N20946);
buf BUF1 (N20952, N20948);
not NOT1 (N20953, N20935);
nor NOR2 (N20954, N20944, N3787);
xor XOR2 (N20955, N20950, N5984);
nand NAND3 (N20956, N20951, N7011, N1518);
nand NAND2 (N20957, N20939, N17379);
buf BUF1 (N20958, N20940);
buf BUF1 (N20959, N20945);
xor XOR2 (N20960, N20955, N2768);
or OR4 (N20961, N20959, N5467, N6620, N3427);
nor NOR2 (N20962, N20927, N3928);
buf BUF1 (N20963, N20957);
buf BUF1 (N20964, N20956);
nand NAND3 (N20965, N20947, N6122, N11263);
not NOT1 (N20966, N20960);
xor XOR2 (N20967, N20953, N17199);
xor XOR2 (N20968, N20965, N13864);
not NOT1 (N20969, N20954);
or OR4 (N20970, N20961, N11536, N8140, N11330);
nor NOR4 (N20971, N20969, N285, N19644, N20530);
nor NOR2 (N20972, N20971, N157);
and AND4 (N20973, N20962, N19316, N15184, N20441);
nand NAND3 (N20974, N20964, N20248, N19880);
buf BUF1 (N20975, N20966);
and AND2 (N20976, N20952, N20786);
not NOT1 (N20977, N20973);
nand NAND2 (N20978, N20974, N16014);
nand NAND2 (N20979, N20967, N13231);
nand NAND2 (N20980, N20958, N12580);
or OR2 (N20981, N20972, N6783);
xor XOR2 (N20982, N20978, N1491);
nand NAND3 (N20983, N20981, N9106, N5413);
nor NOR4 (N20984, N20977, N13101, N5727, N9141);
buf BUF1 (N20985, N20970);
nand NAND4 (N20986, N20979, N18448, N4811, N12555);
buf BUF1 (N20987, N20985);
nand NAND2 (N20988, N20983, N15894);
and AND2 (N20989, N20984, N2983);
or OR4 (N20990, N20976, N8883, N3409, N12430);
not NOT1 (N20991, N20968);
not NOT1 (N20992, N20991);
nor NOR2 (N20993, N20975, N12873);
nor NOR2 (N20994, N20980, N9182);
xor XOR2 (N20995, N20988, N12306);
not NOT1 (N20996, N20982);
or OR2 (N20997, N20989, N4526);
nor NOR2 (N20998, N20987, N17708);
buf BUF1 (N20999, N20997);
nand NAND3 (N21000, N20994, N685, N11865);
xor XOR2 (N21001, N20993, N15152);
xor XOR2 (N21002, N20998, N18188);
or OR2 (N21003, N20992, N12166);
nor NOR3 (N21004, N20963, N6078, N1708);
not NOT1 (N21005, N20986);
and AND2 (N21006, N21005, N3440);
not NOT1 (N21007, N21006);
not NOT1 (N21008, N20996);
not NOT1 (N21009, N21008);
nand NAND4 (N21010, N20990, N11993, N20078, N20703);
xor XOR2 (N21011, N21003, N16765);
and AND4 (N21012, N20995, N3275, N11871, N3114);
xor XOR2 (N21013, N21012, N844);
nand NAND4 (N21014, N21007, N2845, N9024, N1353);
xor XOR2 (N21015, N21010, N7063);
buf BUF1 (N21016, N21001);
nand NAND4 (N21017, N21009, N16460, N7995, N18904);
not NOT1 (N21018, N21017);
nor NOR4 (N21019, N21013, N19781, N14655, N10577);
not NOT1 (N21020, N21019);
and AND4 (N21021, N21000, N8463, N1770, N18809);
or OR2 (N21022, N21015, N1923);
and AND2 (N21023, N21011, N20250);
and AND4 (N21024, N21021, N9246, N560, N20621);
nor NOR3 (N21025, N20999, N18282, N762);
and AND3 (N21026, N21014, N11816, N18566);
and AND3 (N21027, N21022, N19358, N13145);
buf BUF1 (N21028, N21023);
buf BUF1 (N21029, N21020);
buf BUF1 (N21030, N21002);
buf BUF1 (N21031, N21028);
and AND4 (N21032, N21024, N17878, N15014, N3379);
not NOT1 (N21033, N21030);
xor XOR2 (N21034, N21004, N15290);
nor NOR4 (N21035, N21034, N20181, N10425, N5130);
and AND2 (N21036, N21016, N20080);
buf BUF1 (N21037, N21033);
or OR2 (N21038, N21035, N17499);
nor NOR2 (N21039, N21029, N20434);
not NOT1 (N21040, N21027);
and AND2 (N21041, N21031, N13179);
xor XOR2 (N21042, N21036, N17367);
nor NOR3 (N21043, N21038, N5736, N3850);
not NOT1 (N21044, N21032);
or OR2 (N21045, N21043, N16908);
nand NAND2 (N21046, N21026, N18112);
not NOT1 (N21047, N21046);
or OR2 (N21048, N21037, N9384);
buf BUF1 (N21049, N21047);
not NOT1 (N21050, N21041);
xor XOR2 (N21051, N21040, N12016);
xor XOR2 (N21052, N21042, N1722);
and AND3 (N21053, N21039, N20039, N19209);
and AND4 (N21054, N21052, N7500, N18717, N12716);
and AND4 (N21055, N21025, N12439, N7318, N4834);
not NOT1 (N21056, N21018);
or OR4 (N21057, N21056, N5338, N18406, N7437);
or OR3 (N21058, N21053, N17487, N5593);
not NOT1 (N21059, N21049);
nor NOR3 (N21060, N21045, N13388, N20880);
or OR3 (N21061, N21044, N4230, N15364);
or OR2 (N21062, N21059, N17030);
not NOT1 (N21063, N21058);
or OR4 (N21064, N21060, N19589, N1565, N10484);
buf BUF1 (N21065, N21062);
xor XOR2 (N21066, N21054, N10331);
xor XOR2 (N21067, N21050, N1634);
and AND3 (N21068, N21055, N1647, N8548);
or OR2 (N21069, N21064, N4580);
or OR4 (N21070, N21048, N5713, N15683, N2539);
nand NAND3 (N21071, N21051, N17251, N16465);
and AND3 (N21072, N21068, N10065, N9596);
and AND2 (N21073, N21063, N8700);
buf BUF1 (N21074, N21067);
nand NAND4 (N21075, N21072, N6650, N18496, N5379);
or OR2 (N21076, N21074, N13538);
nor NOR3 (N21077, N21066, N2399, N11717);
buf BUF1 (N21078, N21061);
buf BUF1 (N21079, N21076);
not NOT1 (N21080, N21075);
and AND2 (N21081, N21057, N9310);
nor NOR3 (N21082, N21077, N104, N820);
buf BUF1 (N21083, N21073);
nor NOR4 (N21084, N21065, N9750, N5803, N14418);
or OR2 (N21085, N21079, N7574);
xor XOR2 (N21086, N21082, N16539);
xor XOR2 (N21087, N21070, N9693);
not NOT1 (N21088, N21080);
buf BUF1 (N21089, N21078);
and AND3 (N21090, N21087, N8324, N13761);
not NOT1 (N21091, N21089);
nor NOR2 (N21092, N21084, N2635);
and AND3 (N21093, N21092, N1871, N13846);
buf BUF1 (N21094, N21091);
not NOT1 (N21095, N21085);
or OR4 (N21096, N21071, N6392, N11816, N8080);
and AND2 (N21097, N21088, N20266);
nand NAND2 (N21098, N21090, N19793);
buf BUF1 (N21099, N21069);
buf BUF1 (N21100, N21086);
xor XOR2 (N21101, N21097, N5958);
or OR3 (N21102, N21093, N13166, N6085);
nand NAND2 (N21103, N21098, N157);
not NOT1 (N21104, N21102);
and AND4 (N21105, N21099, N15758, N19888, N1152);
buf BUF1 (N21106, N21105);
xor XOR2 (N21107, N21096, N17053);
xor XOR2 (N21108, N21104, N19385);
nand NAND2 (N21109, N21095, N2473);
buf BUF1 (N21110, N21083);
not NOT1 (N21111, N21110);
buf BUF1 (N21112, N21107);
not NOT1 (N21113, N21108);
nand NAND3 (N21114, N21081, N17936, N3714);
and AND4 (N21115, N21113, N10071, N9835, N21088);
xor XOR2 (N21116, N21109, N20178);
and AND3 (N21117, N21094, N9127, N14236);
not NOT1 (N21118, N21117);
nor NOR2 (N21119, N21100, N13164);
nand NAND3 (N21120, N21112, N602, N14281);
nand NAND2 (N21121, N21103, N7896);
nand NAND2 (N21122, N21119, N7444);
not NOT1 (N21123, N21111);
nor NOR3 (N21124, N21116, N20964, N11867);
xor XOR2 (N21125, N21114, N18688);
buf BUF1 (N21126, N21124);
buf BUF1 (N21127, N21126);
not NOT1 (N21128, N21120);
buf BUF1 (N21129, N21127);
not NOT1 (N21130, N21118);
nand NAND3 (N21131, N21121, N617, N5438);
buf BUF1 (N21132, N21123);
nand NAND2 (N21133, N21130, N3641);
nand NAND4 (N21134, N21125, N6755, N17548, N7751);
nand NAND2 (N21135, N21132, N3094);
not NOT1 (N21136, N21128);
nor NOR4 (N21137, N21136, N10665, N16101, N12854);
xor XOR2 (N21138, N21131, N20068);
xor XOR2 (N21139, N21122, N1767);
xor XOR2 (N21140, N21115, N12773);
nor NOR3 (N21141, N21138, N6263, N20249);
and AND4 (N21142, N21141, N5456, N7133, N14673);
not NOT1 (N21143, N21134);
or OR3 (N21144, N21137, N14205, N16761);
buf BUF1 (N21145, N21143);
nor NOR3 (N21146, N21145, N16965, N20257);
not NOT1 (N21147, N21106);
not NOT1 (N21148, N21144);
buf BUF1 (N21149, N21142);
or OR2 (N21150, N21148, N18684);
buf BUF1 (N21151, N21133);
nand NAND4 (N21152, N21139, N3057, N4230, N1855);
nand NAND3 (N21153, N21150, N16098, N15155);
xor XOR2 (N21154, N21152, N17852);
xor XOR2 (N21155, N21135, N8637);
buf BUF1 (N21156, N21151);
nor NOR2 (N21157, N21147, N14753);
nand NAND4 (N21158, N21157, N7495, N13791, N12709);
or OR4 (N21159, N21153, N21133, N8463, N10337);
nor NOR4 (N21160, N21159, N11959, N9374, N20165);
buf BUF1 (N21161, N21101);
xor XOR2 (N21162, N21149, N9269);
xor XOR2 (N21163, N21140, N14256);
nor NOR2 (N21164, N21163, N14046);
xor XOR2 (N21165, N21161, N15419);
nor NOR2 (N21166, N21156, N6905);
nand NAND4 (N21167, N21129, N11215, N11949, N7943);
or OR4 (N21168, N21164, N2464, N11039, N12104);
buf BUF1 (N21169, N21168);
xor XOR2 (N21170, N21154, N8141);
buf BUF1 (N21171, N21165);
buf BUF1 (N21172, N21162);
buf BUF1 (N21173, N21172);
nor NOR2 (N21174, N21158, N19377);
buf BUF1 (N21175, N21146);
buf BUF1 (N21176, N21170);
buf BUF1 (N21177, N21169);
buf BUF1 (N21178, N21167);
not NOT1 (N21179, N21174);
nand NAND4 (N21180, N21178, N13045, N13188, N3459);
nor NOR2 (N21181, N21155, N4251);
and AND4 (N21182, N21166, N5700, N9472, N8350);
nand NAND2 (N21183, N21176, N10729);
nand NAND3 (N21184, N21177, N12338, N361);
nor NOR3 (N21185, N21181, N8731, N16401);
nor NOR3 (N21186, N21175, N8275, N16780);
not NOT1 (N21187, N21160);
buf BUF1 (N21188, N21186);
buf BUF1 (N21189, N21179);
or OR4 (N21190, N21182, N8910, N19808, N12812);
not NOT1 (N21191, N21183);
buf BUF1 (N21192, N21185);
and AND4 (N21193, N21189, N6367, N9447, N17551);
buf BUF1 (N21194, N21192);
xor XOR2 (N21195, N21190, N10217);
not NOT1 (N21196, N21191);
not NOT1 (N21197, N21171);
and AND2 (N21198, N21197, N9307);
not NOT1 (N21199, N21173);
not NOT1 (N21200, N21193);
xor XOR2 (N21201, N21188, N18685);
not NOT1 (N21202, N21198);
nand NAND3 (N21203, N21200, N19261, N6620);
not NOT1 (N21204, N21194);
or OR3 (N21205, N21202, N2172, N4105);
and AND2 (N21206, N21195, N12063);
nor NOR2 (N21207, N21205, N15204);
xor XOR2 (N21208, N21206, N5977);
not NOT1 (N21209, N21199);
nor NOR3 (N21210, N21209, N169, N15697);
and AND2 (N21211, N21204, N5097);
or OR2 (N21212, N21201, N14720);
and AND2 (N21213, N21210, N5479);
or OR2 (N21214, N21213, N9534);
nand NAND4 (N21215, N21211, N8237, N1141, N6606);
or OR2 (N21216, N21184, N8464);
or OR4 (N21217, N21214, N7216, N15596, N17716);
xor XOR2 (N21218, N21216, N5353);
or OR2 (N21219, N21217, N7781);
or OR3 (N21220, N21207, N19223, N17672);
xor XOR2 (N21221, N21212, N9818);
not NOT1 (N21222, N21215);
buf BUF1 (N21223, N21203);
nand NAND2 (N21224, N21196, N16041);
and AND4 (N21225, N21187, N12838, N4667, N18905);
nand NAND3 (N21226, N21221, N1989, N14280);
or OR3 (N21227, N21225, N14830, N12435);
xor XOR2 (N21228, N21226, N9362);
not NOT1 (N21229, N21222);
xor XOR2 (N21230, N21208, N6051);
xor XOR2 (N21231, N21223, N14786);
or OR4 (N21232, N21231, N3200, N8024, N7253);
or OR2 (N21233, N21219, N13698);
and AND2 (N21234, N21220, N15970);
nand NAND3 (N21235, N21228, N4185, N20292);
not NOT1 (N21236, N21227);
buf BUF1 (N21237, N21232);
nor NOR4 (N21238, N21218, N10827, N13012, N7094);
buf BUF1 (N21239, N21234);
nand NAND4 (N21240, N21180, N12405, N10620, N3981);
and AND4 (N21241, N21229, N15918, N19812, N10433);
nand NAND2 (N21242, N21239, N9441);
nand NAND3 (N21243, N21241, N9740, N14185);
not NOT1 (N21244, N21235);
xor XOR2 (N21245, N21224, N15388);
or OR2 (N21246, N21230, N9089);
buf BUF1 (N21247, N21243);
not NOT1 (N21248, N21233);
xor XOR2 (N21249, N21246, N12136);
or OR3 (N21250, N21236, N17486, N5660);
xor XOR2 (N21251, N21242, N1698);
nor NOR3 (N21252, N21251, N13800, N7604);
xor XOR2 (N21253, N21250, N9791);
xor XOR2 (N21254, N21253, N12842);
buf BUF1 (N21255, N21240);
or OR3 (N21256, N21255, N3764, N2597);
xor XOR2 (N21257, N21247, N17630);
nand NAND4 (N21258, N21244, N13803, N5936, N8773);
or OR4 (N21259, N21257, N10725, N3360, N8578);
and AND3 (N21260, N21245, N19581, N17301);
xor XOR2 (N21261, N21254, N12992);
or OR3 (N21262, N21258, N66, N12311);
and AND3 (N21263, N21256, N18438, N10762);
xor XOR2 (N21264, N21259, N10822);
buf BUF1 (N21265, N21262);
buf BUF1 (N21266, N21263);
not NOT1 (N21267, N21264);
or OR2 (N21268, N21249, N12521);
xor XOR2 (N21269, N21238, N5534);
xor XOR2 (N21270, N21265, N11557);
not NOT1 (N21271, N21270);
xor XOR2 (N21272, N21252, N8156);
and AND4 (N21273, N21237, N11828, N15213, N20684);
not NOT1 (N21274, N21268);
nand NAND3 (N21275, N21248, N10751, N6941);
not NOT1 (N21276, N21274);
nand NAND4 (N21277, N21266, N16489, N9597, N19314);
nor NOR2 (N21278, N21275, N19706);
xor XOR2 (N21279, N21260, N13721);
buf BUF1 (N21280, N21277);
nand NAND3 (N21281, N21269, N20720, N11620);
not NOT1 (N21282, N21261);
nand NAND4 (N21283, N21279, N3813, N11268, N16685);
nor NOR4 (N21284, N21282, N1189, N13634, N1458);
nor NOR3 (N21285, N21267, N15203, N11345);
or OR3 (N21286, N21276, N20063, N16577);
nor NOR3 (N21287, N21278, N1676, N13069);
nor NOR2 (N21288, N21287, N6618);
not NOT1 (N21289, N21286);
nand NAND3 (N21290, N21271, N11473, N9840);
xor XOR2 (N21291, N21288, N19557);
nand NAND2 (N21292, N21284, N20745);
nor NOR2 (N21293, N21273, N18781);
buf BUF1 (N21294, N21280);
not NOT1 (N21295, N21291);
buf BUF1 (N21296, N21292);
not NOT1 (N21297, N21290);
buf BUF1 (N21298, N21293);
xor XOR2 (N21299, N21296, N4165);
and AND3 (N21300, N21289, N6207, N5189);
xor XOR2 (N21301, N21298, N11948);
nand NAND3 (N21302, N21299, N11628, N19420);
xor XOR2 (N21303, N21294, N11007);
or OR4 (N21304, N21283, N6452, N10407, N12609);
not NOT1 (N21305, N21281);
or OR3 (N21306, N21295, N13338, N4803);
and AND2 (N21307, N21300, N14294);
buf BUF1 (N21308, N21285);
xor XOR2 (N21309, N21307, N12752);
buf BUF1 (N21310, N21304);
xor XOR2 (N21311, N21297, N19263);
buf BUF1 (N21312, N21303);
nand NAND2 (N21313, N21311, N15305);
buf BUF1 (N21314, N21301);
and AND4 (N21315, N21306, N14968, N4, N9698);
nor NOR2 (N21316, N21312, N11454);
buf BUF1 (N21317, N21310);
buf BUF1 (N21318, N21309);
xor XOR2 (N21319, N21305, N6122);
and AND2 (N21320, N21272, N9467);
nor NOR2 (N21321, N21315, N18930);
nor NOR3 (N21322, N21318, N15252, N3818);
xor XOR2 (N21323, N21314, N21062);
buf BUF1 (N21324, N21321);
buf BUF1 (N21325, N21323);
not NOT1 (N21326, N21319);
nor NOR3 (N21327, N21320, N1774, N20276);
xor XOR2 (N21328, N21325, N5329);
buf BUF1 (N21329, N21324);
nor NOR4 (N21330, N21322, N18699, N20466, N2070);
or OR4 (N21331, N21327, N7292, N803, N5682);
or OR3 (N21332, N21308, N7908, N2710);
and AND4 (N21333, N21316, N2429, N18011, N17348);
buf BUF1 (N21334, N21331);
xor XOR2 (N21335, N21329, N244);
or OR2 (N21336, N21313, N9339);
and AND4 (N21337, N21302, N12656, N8585, N14851);
nor NOR3 (N21338, N21326, N14455, N18116);
or OR2 (N21339, N21335, N10008);
nor NOR2 (N21340, N21334, N8798);
nor NOR4 (N21341, N21333, N7299, N225, N13392);
buf BUF1 (N21342, N21328);
nand NAND3 (N21343, N21337, N513, N9644);
not NOT1 (N21344, N21330);
xor XOR2 (N21345, N21338, N1485);
nor NOR3 (N21346, N21344, N10555, N18828);
nor NOR2 (N21347, N21341, N9699);
xor XOR2 (N21348, N21343, N19836);
not NOT1 (N21349, N21348);
not NOT1 (N21350, N21349);
nor NOR3 (N21351, N21347, N2926, N16685);
and AND3 (N21352, N21345, N6366, N17123);
nor NOR3 (N21353, N21340, N9787, N17774);
nand NAND4 (N21354, N21332, N17634, N3873, N5351);
nand NAND3 (N21355, N21353, N18903, N17719);
xor XOR2 (N21356, N21317, N591);
and AND4 (N21357, N21352, N15591, N10025, N14981);
xor XOR2 (N21358, N21354, N720);
buf BUF1 (N21359, N21342);
buf BUF1 (N21360, N21336);
nand NAND2 (N21361, N21357, N2597);
nor NOR4 (N21362, N21350, N10315, N9731, N14831);
nand NAND3 (N21363, N21358, N16228, N15716);
nand NAND3 (N21364, N21339, N20993, N13124);
and AND3 (N21365, N21362, N825, N3261);
nor NOR4 (N21366, N21355, N5829, N18205, N1861);
or OR2 (N21367, N21363, N12605);
nor NOR3 (N21368, N21365, N8952, N20555);
buf BUF1 (N21369, N21367);
and AND4 (N21370, N21361, N6753, N5091, N2760);
not NOT1 (N21371, N21364);
not NOT1 (N21372, N21370);
not NOT1 (N21373, N21371);
xor XOR2 (N21374, N21372, N12485);
or OR4 (N21375, N21374, N17411, N12466, N10995);
nand NAND4 (N21376, N21368, N6265, N17955, N510);
nand NAND2 (N21377, N21351, N18964);
nand NAND4 (N21378, N21359, N2960, N13795, N11006);
and AND3 (N21379, N21360, N4484, N13120);
buf BUF1 (N21380, N21346);
buf BUF1 (N21381, N21376);
nor NOR3 (N21382, N21373, N10551, N9175);
buf BUF1 (N21383, N21379);
xor XOR2 (N21384, N21356, N19359);
and AND2 (N21385, N21381, N18158);
xor XOR2 (N21386, N21385, N15657);
and AND4 (N21387, N21366, N7863, N11961, N4529);
not NOT1 (N21388, N21382);
nand NAND2 (N21389, N21384, N3909);
buf BUF1 (N21390, N21387);
and AND2 (N21391, N21377, N9904);
nand NAND4 (N21392, N21390, N18881, N15084, N10449);
xor XOR2 (N21393, N21378, N1167);
buf BUF1 (N21394, N21375);
and AND2 (N21395, N21380, N16138);
nor NOR2 (N21396, N21391, N10701);
or OR2 (N21397, N21396, N14480);
buf BUF1 (N21398, N21393);
nand NAND3 (N21399, N21397, N18492, N1700);
nor NOR4 (N21400, N21389, N5506, N12548, N18467);
not NOT1 (N21401, N21392);
or OR4 (N21402, N21386, N6938, N19479, N19457);
nor NOR2 (N21403, N21394, N15852);
buf BUF1 (N21404, N21383);
or OR4 (N21405, N21369, N11534, N15911, N10811);
and AND4 (N21406, N21398, N6185, N20333, N18666);
nand NAND4 (N21407, N21402, N6824, N19913, N7620);
buf BUF1 (N21408, N21405);
and AND2 (N21409, N21388, N2718);
xor XOR2 (N21410, N21401, N20184);
xor XOR2 (N21411, N21403, N7814);
buf BUF1 (N21412, N21400);
nor NOR3 (N21413, N21407, N14657, N2847);
nor NOR3 (N21414, N21395, N6244, N3588);
or OR2 (N21415, N21412, N18774);
nand NAND3 (N21416, N21410, N21117, N20017);
or OR2 (N21417, N21408, N4658);
nand NAND2 (N21418, N21404, N18430);
and AND2 (N21419, N21416, N18592);
not NOT1 (N21420, N21419);
not NOT1 (N21421, N21399);
buf BUF1 (N21422, N21417);
or OR4 (N21423, N21411, N15280, N14577, N1774);
buf BUF1 (N21424, N21423);
buf BUF1 (N21425, N21422);
not NOT1 (N21426, N21424);
not NOT1 (N21427, N21409);
buf BUF1 (N21428, N21415);
and AND4 (N21429, N21414, N13834, N148, N9370);
buf BUF1 (N21430, N21429);
not NOT1 (N21431, N21413);
xor XOR2 (N21432, N21427, N20292);
nor NOR3 (N21433, N21406, N13068, N20963);
nand NAND4 (N21434, N21426, N12300, N5616, N8052);
xor XOR2 (N21435, N21433, N17473);
nand NAND3 (N21436, N21430, N342, N9086);
or OR3 (N21437, N21431, N20276, N2673);
or OR3 (N21438, N21421, N14848, N12005);
and AND2 (N21439, N21425, N14709);
and AND2 (N21440, N21437, N9113);
not NOT1 (N21441, N21432);
buf BUF1 (N21442, N21435);
nand NAND4 (N21443, N21420, N8080, N10529, N14318);
xor XOR2 (N21444, N21441, N16619);
or OR4 (N21445, N21442, N15241, N14823, N626);
not NOT1 (N21446, N21445);
nand NAND3 (N21447, N21436, N15240, N1176);
xor XOR2 (N21448, N21447, N4681);
nand NAND4 (N21449, N21448, N6922, N19559, N16258);
xor XOR2 (N21450, N21428, N15795);
nor NOR4 (N21451, N21438, N7051, N19322, N5272);
and AND4 (N21452, N21443, N7891, N17706, N8747);
buf BUF1 (N21453, N21434);
buf BUF1 (N21454, N21452);
nand NAND2 (N21455, N21440, N13025);
buf BUF1 (N21456, N21418);
xor XOR2 (N21457, N21449, N10284);
not NOT1 (N21458, N21444);
not NOT1 (N21459, N21446);
nor NOR4 (N21460, N21457, N6700, N7090, N19496);
buf BUF1 (N21461, N21454);
or OR3 (N21462, N21453, N7565, N20430);
and AND3 (N21463, N21460, N21164, N18427);
and AND3 (N21464, N21458, N20241, N9567);
or OR3 (N21465, N21464, N2450, N19567);
buf BUF1 (N21466, N21461);
or OR4 (N21467, N21439, N12217, N4433, N11195);
not NOT1 (N21468, N21466);
or OR2 (N21469, N21450, N10899);
xor XOR2 (N21470, N21451, N13028);
not NOT1 (N21471, N21468);
buf BUF1 (N21472, N21469);
xor XOR2 (N21473, N21472, N9029);
nor NOR3 (N21474, N21471, N6294, N9747);
not NOT1 (N21475, N21474);
not NOT1 (N21476, N21465);
not NOT1 (N21477, N21455);
xor XOR2 (N21478, N21456, N20948);
not NOT1 (N21479, N21459);
buf BUF1 (N21480, N21477);
and AND2 (N21481, N21478, N9922);
nand NAND4 (N21482, N21475, N1408, N622, N13998);
nor NOR3 (N21483, N21473, N979, N11145);
buf BUF1 (N21484, N21476);
nand NAND4 (N21485, N21481, N1111, N14545, N7055);
not NOT1 (N21486, N21480);
or OR2 (N21487, N21479, N11648);
and AND4 (N21488, N21462, N8471, N18227, N11338);
xor XOR2 (N21489, N21483, N15077);
xor XOR2 (N21490, N21463, N19762);
or OR4 (N21491, N21467, N20586, N1543, N12544);
xor XOR2 (N21492, N21488, N16920);
nand NAND3 (N21493, N21490, N14906, N14005);
buf BUF1 (N21494, N21487);
nand NAND2 (N21495, N21470, N20862);
buf BUF1 (N21496, N21494);
and AND3 (N21497, N21491, N15760, N5584);
xor XOR2 (N21498, N21484, N21414);
or OR4 (N21499, N21486, N17207, N8115, N18711);
or OR3 (N21500, N21496, N4488, N8878);
nor NOR4 (N21501, N21482, N10194, N15625, N16054);
and AND3 (N21502, N21501, N15322, N15500);
and AND2 (N21503, N21500, N11394);
xor XOR2 (N21504, N21499, N2852);
not NOT1 (N21505, N21489);
or OR4 (N21506, N21497, N14723, N11489, N17077);
nor NOR4 (N21507, N21502, N3553, N2876, N11845);
buf BUF1 (N21508, N21498);
and AND3 (N21509, N21503, N15277, N5494);
and AND4 (N21510, N21493, N1392, N18403, N7448);
and AND2 (N21511, N21485, N3504);
xor XOR2 (N21512, N21492, N17326);
nor NOR2 (N21513, N21495, N7670);
nor NOR2 (N21514, N21505, N7680);
not NOT1 (N21515, N21507);
buf BUF1 (N21516, N21510);
nand NAND3 (N21517, N21506, N10444, N726);
not NOT1 (N21518, N21517);
nor NOR3 (N21519, N21511, N8976, N3515);
buf BUF1 (N21520, N21504);
or OR3 (N21521, N21520, N230, N18267);
not NOT1 (N21522, N21519);
and AND4 (N21523, N21514, N7652, N19827, N160);
or OR3 (N21524, N21516, N20316, N6442);
nor NOR2 (N21525, N21508, N15409);
not NOT1 (N21526, N21522);
nor NOR4 (N21527, N21525, N4472, N4893, N6865);
or OR2 (N21528, N21527, N4388);
not NOT1 (N21529, N21513);
or OR2 (N21530, N21529, N20664);
and AND3 (N21531, N21512, N7527, N2160);
not NOT1 (N21532, N21531);
or OR4 (N21533, N21509, N3133, N19066, N13563);
buf BUF1 (N21534, N21533);
not NOT1 (N21535, N21523);
not NOT1 (N21536, N21528);
buf BUF1 (N21537, N21515);
or OR3 (N21538, N21530, N12011, N13961);
or OR4 (N21539, N21538, N6713, N11865, N17231);
xor XOR2 (N21540, N21535, N18904);
nor NOR2 (N21541, N21539, N1737);
and AND3 (N21542, N21537, N16768, N668);
and AND3 (N21543, N21521, N18077, N11169);
not NOT1 (N21544, N21542);
nand NAND4 (N21545, N21536, N7553, N11857, N754);
or OR3 (N21546, N21518, N6267, N2131);
and AND4 (N21547, N21541, N13153, N871, N7890);
or OR4 (N21548, N21540, N10819, N8809, N14616);
nor NOR4 (N21549, N21545, N1497, N3781, N5094);
buf BUF1 (N21550, N21534);
or OR4 (N21551, N21549, N6749, N15983, N3517);
not NOT1 (N21552, N21526);
nand NAND4 (N21553, N21532, N17877, N7175, N16373);
nand NAND4 (N21554, N21553, N149, N9026, N16765);
not NOT1 (N21555, N21547);
xor XOR2 (N21556, N21555, N15605);
nand NAND2 (N21557, N21551, N5772);
not NOT1 (N21558, N21557);
buf BUF1 (N21559, N21543);
buf BUF1 (N21560, N21524);
xor XOR2 (N21561, N21550, N11035);
buf BUF1 (N21562, N21554);
or OR4 (N21563, N21548, N9915, N9027, N20857);
buf BUF1 (N21564, N21546);
nand NAND3 (N21565, N21563, N3064, N14199);
not NOT1 (N21566, N21565);
not NOT1 (N21567, N21558);
not NOT1 (N21568, N21562);
nor NOR2 (N21569, N21544, N8703);
or OR3 (N21570, N21566, N10952, N12607);
or OR2 (N21571, N21567, N1933);
and AND4 (N21572, N21561, N10617, N10245, N9908);
buf BUF1 (N21573, N21560);
buf BUF1 (N21574, N21556);
and AND2 (N21575, N21573, N145);
not NOT1 (N21576, N21572);
or OR4 (N21577, N21574, N6660, N17517, N12959);
nand NAND3 (N21578, N21577, N5117, N8350);
nand NAND2 (N21579, N21552, N4811);
nand NAND4 (N21580, N21568, N14336, N16214, N7614);
nor NOR3 (N21581, N21564, N2709, N4152);
nand NAND4 (N21582, N21579, N20375, N18117, N19084);
nand NAND3 (N21583, N21576, N2214, N16673);
not NOT1 (N21584, N21581);
and AND2 (N21585, N21578, N4653);
nor NOR3 (N21586, N21559, N3760, N10979);
nor NOR3 (N21587, N21583, N19920, N10468);
and AND4 (N21588, N21570, N10399, N10401, N16769);
buf BUF1 (N21589, N21575);
buf BUF1 (N21590, N21588);
or OR3 (N21591, N21582, N8654, N7020);
nor NOR3 (N21592, N21590, N5713, N15550);
and AND3 (N21593, N21580, N13502, N17992);
and AND2 (N21594, N21592, N10130);
nor NOR3 (N21595, N21591, N13932, N18649);
and AND2 (N21596, N21589, N1511);
not NOT1 (N21597, N21571);
nand NAND4 (N21598, N21596, N11476, N18384, N7433);
not NOT1 (N21599, N21598);
and AND2 (N21600, N21595, N5853);
nor NOR3 (N21601, N21569, N13110, N20529);
xor XOR2 (N21602, N21600, N9123);
xor XOR2 (N21603, N21587, N8891);
buf BUF1 (N21604, N21593);
nand NAND3 (N21605, N21585, N19830, N16352);
xor XOR2 (N21606, N21584, N4354);
buf BUF1 (N21607, N21605);
or OR4 (N21608, N21601, N19833, N9995, N1203);
nand NAND3 (N21609, N21607, N8250, N560);
buf BUF1 (N21610, N21609);
nor NOR2 (N21611, N21586, N5839);
and AND4 (N21612, N21608, N16892, N16609, N17250);
or OR3 (N21613, N21606, N14941, N15995);
or OR2 (N21614, N21612, N14847);
xor XOR2 (N21615, N21603, N21054);
and AND2 (N21616, N21594, N7478);
xor XOR2 (N21617, N21611, N15800);
not NOT1 (N21618, N21617);
or OR3 (N21619, N21602, N11933, N17384);
nand NAND4 (N21620, N21610, N5068, N18891, N9002);
or OR4 (N21621, N21615, N10633, N10969, N19530);
not NOT1 (N21622, N21604);
nor NOR3 (N21623, N21618, N12053, N12347);
buf BUF1 (N21624, N21613);
nand NAND2 (N21625, N21620, N1702);
not NOT1 (N21626, N21599);
nand NAND3 (N21627, N21614, N8973, N19562);
nor NOR2 (N21628, N21616, N17603);
buf BUF1 (N21629, N21621);
xor XOR2 (N21630, N21628, N10098);
xor XOR2 (N21631, N21625, N7428);
not NOT1 (N21632, N21627);
xor XOR2 (N21633, N21597, N6936);
buf BUF1 (N21634, N21626);
nor NOR4 (N21635, N21632, N9684, N13445, N19421);
buf BUF1 (N21636, N21633);
or OR3 (N21637, N21619, N11410, N7094);
nand NAND2 (N21638, N21634, N14661);
or OR3 (N21639, N21638, N12513, N9222);
buf BUF1 (N21640, N21622);
nor NOR4 (N21641, N21630, N8607, N11919, N16751);
xor XOR2 (N21642, N21623, N256);
buf BUF1 (N21643, N21642);
and AND4 (N21644, N21637, N19214, N16506, N6504);
nand NAND2 (N21645, N21636, N7668);
nor NOR3 (N21646, N21644, N8867, N8857);
nor NOR4 (N21647, N21631, N10098, N13287, N1456);
not NOT1 (N21648, N21645);
xor XOR2 (N21649, N21635, N21095);
nand NAND3 (N21650, N21648, N11744, N13300);
xor XOR2 (N21651, N21646, N2157);
or OR4 (N21652, N21651, N3582, N19647, N4687);
buf BUF1 (N21653, N21639);
nor NOR3 (N21654, N21624, N14725, N18341);
nand NAND4 (N21655, N21629, N3541, N5543, N20010);
nor NOR3 (N21656, N21655, N875, N14559);
buf BUF1 (N21657, N21649);
not NOT1 (N21658, N21641);
and AND3 (N21659, N21640, N12027, N13883);
nand NAND3 (N21660, N21656, N15895, N14253);
nand NAND2 (N21661, N21659, N17810);
not NOT1 (N21662, N21660);
xor XOR2 (N21663, N21652, N7304);
nand NAND4 (N21664, N21647, N17990, N18015, N17587);
xor XOR2 (N21665, N21663, N10776);
not NOT1 (N21666, N21643);
nand NAND2 (N21667, N21661, N10907);
and AND3 (N21668, N21667, N9610, N12923);
xor XOR2 (N21669, N21658, N2590);
xor XOR2 (N21670, N21669, N16169);
nand NAND3 (N21671, N21670, N7262, N11412);
nand NAND4 (N21672, N21666, N4095, N10345, N1113);
nand NAND4 (N21673, N21668, N8470, N6572, N13726);
nor NOR3 (N21674, N21654, N19517, N5016);
nor NOR3 (N21675, N21671, N6970, N7904);
buf BUF1 (N21676, N21662);
and AND3 (N21677, N21674, N7530, N17581);
and AND3 (N21678, N21664, N1511, N8049);
not NOT1 (N21679, N21676);
nand NAND4 (N21680, N21679, N18605, N14499, N10165);
or OR3 (N21681, N21677, N598, N11647);
not NOT1 (N21682, N21653);
nor NOR3 (N21683, N21682, N7012, N10);
nor NOR2 (N21684, N21683, N4867);
not NOT1 (N21685, N21684);
or OR2 (N21686, N21650, N6623);
buf BUF1 (N21687, N21685);
nand NAND4 (N21688, N21678, N18043, N10833, N16725);
nor NOR3 (N21689, N21657, N6056, N20926);
xor XOR2 (N21690, N21672, N4544);
not NOT1 (N21691, N21689);
not NOT1 (N21692, N21691);
and AND2 (N21693, N21675, N14941);
xor XOR2 (N21694, N21690, N18530);
xor XOR2 (N21695, N21692, N20765);
nor NOR3 (N21696, N21665, N7399, N1911);
nor NOR2 (N21697, N21681, N2551);
or OR4 (N21698, N21693, N6072, N1598, N17629);
xor XOR2 (N21699, N21680, N4304);
buf BUF1 (N21700, N21695);
xor XOR2 (N21701, N21696, N21022);
and AND3 (N21702, N21694, N1320, N12980);
nor NOR4 (N21703, N21697, N16022, N17626, N10669);
buf BUF1 (N21704, N21688);
xor XOR2 (N21705, N21673, N11718);
xor XOR2 (N21706, N21704, N444);
xor XOR2 (N21707, N21705, N6074);
buf BUF1 (N21708, N21701);
not NOT1 (N21709, N21700);
buf BUF1 (N21710, N21687);
buf BUF1 (N21711, N21706);
or OR2 (N21712, N21686, N2641);
not NOT1 (N21713, N21712);
not NOT1 (N21714, N21703);
nor NOR3 (N21715, N21711, N5438, N10525);
and AND4 (N21716, N21699, N7495, N13235, N18577);
xor XOR2 (N21717, N21698, N15782);
buf BUF1 (N21718, N21708);
or OR2 (N21719, N21709, N16090);
nor NOR4 (N21720, N21702, N20756, N15872, N11966);
nand NAND4 (N21721, N21714, N19907, N5907, N18801);
nor NOR4 (N21722, N21715, N2577, N21564, N9102);
xor XOR2 (N21723, N21707, N10946);
nand NAND4 (N21724, N21722, N13616, N53, N18780);
and AND2 (N21725, N21723, N10346);
not NOT1 (N21726, N21721);
not NOT1 (N21727, N21720);
nor NOR4 (N21728, N21727, N15793, N14302, N12427);
not NOT1 (N21729, N21728);
and AND4 (N21730, N21717, N13306, N9376, N4922);
xor XOR2 (N21731, N21713, N11009);
nor NOR4 (N21732, N21724, N14497, N8084, N11124);
and AND4 (N21733, N21718, N8396, N5595, N7073);
nand NAND3 (N21734, N21710, N18186, N5907);
or OR4 (N21735, N21719, N10194, N18845, N2483);
nor NOR3 (N21736, N21735, N6780, N11433);
nand NAND2 (N21737, N21716, N14077);
nor NOR2 (N21738, N21729, N19415);
nand NAND3 (N21739, N21734, N14818, N8635);
nor NOR2 (N21740, N21732, N6921);
nand NAND4 (N21741, N21726, N3247, N8032, N11669);
not NOT1 (N21742, N21725);
nand NAND2 (N21743, N21740, N14885);
or OR4 (N21744, N21743, N8117, N4892, N14270);
buf BUF1 (N21745, N21730);
buf BUF1 (N21746, N21737);
nand NAND2 (N21747, N21736, N17137);
and AND3 (N21748, N21731, N1515, N12828);
nor NOR3 (N21749, N21742, N952, N19586);
nand NAND2 (N21750, N21739, N8641);
buf BUF1 (N21751, N21744);
nor NOR3 (N21752, N21749, N3819, N5058);
buf BUF1 (N21753, N21738);
and AND2 (N21754, N21741, N9571);
and AND3 (N21755, N21748, N13626, N6803);
not NOT1 (N21756, N21755);
and AND2 (N21757, N21746, N6833);
buf BUF1 (N21758, N21753);
not NOT1 (N21759, N21751);
or OR2 (N21760, N21750, N12146);
not NOT1 (N21761, N21759);
and AND2 (N21762, N21733, N21240);
nor NOR2 (N21763, N21760, N6964);
buf BUF1 (N21764, N21762);
nor NOR3 (N21765, N21745, N15701, N18527);
buf BUF1 (N21766, N21752);
or OR3 (N21767, N21765, N15417, N1270);
and AND4 (N21768, N21763, N11278, N1929, N13319);
xor XOR2 (N21769, N21758, N17708);
nor NOR3 (N21770, N21754, N9294, N19763);
nor NOR4 (N21771, N21761, N4891, N13232, N8102);
buf BUF1 (N21772, N21770);
or OR3 (N21773, N21767, N13685, N13398);
xor XOR2 (N21774, N21764, N2798);
nor NOR2 (N21775, N21757, N12841);
or OR4 (N21776, N21766, N12068, N12047, N14573);
and AND4 (N21777, N21768, N5921, N7598, N3995);
nor NOR2 (N21778, N21775, N1114);
nor NOR3 (N21779, N21756, N7551, N10492);
xor XOR2 (N21780, N21779, N17614);
buf BUF1 (N21781, N21772);
or OR2 (N21782, N21778, N11448);
nand NAND2 (N21783, N21774, N13640);
xor XOR2 (N21784, N21782, N4286);
nand NAND3 (N21785, N21771, N18052, N7215);
nand NAND4 (N21786, N21783, N18953, N3479, N18978);
not NOT1 (N21787, N21780);
nand NAND4 (N21788, N21786, N6424, N12916, N6467);
nand NAND3 (N21789, N21747, N15449, N6144);
not NOT1 (N21790, N21773);
buf BUF1 (N21791, N21789);
and AND4 (N21792, N21784, N17747, N14420, N17955);
xor XOR2 (N21793, N21787, N17416);
not NOT1 (N21794, N21781);
xor XOR2 (N21795, N21777, N17275);
nor NOR2 (N21796, N21793, N17084);
nor NOR3 (N21797, N21795, N1028, N3041);
nor NOR2 (N21798, N21794, N14077);
xor XOR2 (N21799, N21785, N21186);
and AND4 (N21800, N21791, N3739, N4891, N1106);
or OR4 (N21801, N21797, N5247, N12877, N6600);
not NOT1 (N21802, N21801);
nand NAND3 (N21803, N21796, N2317, N17475);
buf BUF1 (N21804, N21798);
xor XOR2 (N21805, N21792, N21605);
nand NAND2 (N21806, N21804, N1979);
buf BUF1 (N21807, N21769);
nand NAND2 (N21808, N21776, N10734);
nand NAND2 (N21809, N21803, N9956);
nand NAND2 (N21810, N21788, N19995);
and AND4 (N21811, N21802, N2165, N1228, N16296);
nor NOR2 (N21812, N21805, N11765);
xor XOR2 (N21813, N21790, N7924);
xor XOR2 (N21814, N21807, N15651);
buf BUF1 (N21815, N21808);
xor XOR2 (N21816, N21811, N4600);
xor XOR2 (N21817, N21813, N19424);
and AND3 (N21818, N21814, N13666, N7457);
nor NOR4 (N21819, N21809, N3654, N19254, N15400);
xor XOR2 (N21820, N21817, N10096);
nand NAND3 (N21821, N21818, N7211, N7221);
or OR3 (N21822, N21812, N10743, N7689);
xor XOR2 (N21823, N21815, N10275);
or OR2 (N21824, N21816, N10862);
nor NOR2 (N21825, N21823, N14812);
and AND2 (N21826, N21821, N9709);
and AND4 (N21827, N21810, N7714, N8076, N21181);
and AND3 (N21828, N21824, N18060, N18764);
not NOT1 (N21829, N21825);
or OR3 (N21830, N21827, N4135, N13946);
nor NOR4 (N21831, N21820, N2869, N15014, N13450);
xor XOR2 (N21832, N21830, N18724);
and AND2 (N21833, N21819, N9192);
xor XOR2 (N21834, N21832, N17063);
buf BUF1 (N21835, N21829);
or OR3 (N21836, N21822, N11102, N3027);
not NOT1 (N21837, N21806);
buf BUF1 (N21838, N21837);
or OR4 (N21839, N21835, N10065, N4130, N12048);
buf BUF1 (N21840, N21831);
and AND3 (N21841, N21826, N16083, N10433);
xor XOR2 (N21842, N21838, N11132);
nor NOR2 (N21843, N21828, N9207);
nor NOR2 (N21844, N21839, N12949);
xor XOR2 (N21845, N21800, N7784);
and AND2 (N21846, N21841, N19150);
nor NOR4 (N21847, N21845, N18896, N8341, N3947);
nor NOR2 (N21848, N21833, N3085);
xor XOR2 (N21849, N21834, N14593);
not NOT1 (N21850, N21848);
nor NOR3 (N21851, N21844, N7766, N12364);
and AND2 (N21852, N21846, N4320);
or OR2 (N21853, N21842, N8357);
nor NOR3 (N21854, N21849, N5808, N8731);
xor XOR2 (N21855, N21840, N2878);
not NOT1 (N21856, N21854);
nand NAND3 (N21857, N21851, N11927, N9703);
xor XOR2 (N21858, N21856, N5329);
and AND2 (N21859, N21853, N4882);
or OR2 (N21860, N21843, N8183);
buf BUF1 (N21861, N21852);
nor NOR3 (N21862, N21859, N14796, N8237);
xor XOR2 (N21863, N21862, N10540);
nor NOR3 (N21864, N21860, N13668, N6716);
nand NAND2 (N21865, N21864, N15186);
buf BUF1 (N21866, N21855);
xor XOR2 (N21867, N21863, N19984);
xor XOR2 (N21868, N21799, N12578);
buf BUF1 (N21869, N21858);
not NOT1 (N21870, N21857);
xor XOR2 (N21871, N21869, N17855);
xor XOR2 (N21872, N21865, N14704);
nor NOR4 (N21873, N21861, N9427, N20600, N4846);
buf BUF1 (N21874, N21847);
nor NOR4 (N21875, N21866, N17091, N887, N12356);
nand NAND3 (N21876, N21850, N7377, N614);
not NOT1 (N21877, N21873);
xor XOR2 (N21878, N21872, N19349);
nand NAND2 (N21879, N21867, N17811);
xor XOR2 (N21880, N21878, N9291);
nand NAND2 (N21881, N21879, N7294);
or OR3 (N21882, N21881, N13451, N20745);
and AND2 (N21883, N21882, N7834);
xor XOR2 (N21884, N21876, N2611);
xor XOR2 (N21885, N21874, N18561);
xor XOR2 (N21886, N21883, N17767);
xor XOR2 (N21887, N21868, N11544);
or OR4 (N21888, N21871, N14055, N11492, N5004);
or OR2 (N21889, N21875, N16036);
nand NAND3 (N21890, N21836, N7602, N6566);
not NOT1 (N21891, N21888);
and AND3 (N21892, N21870, N4995, N20480);
or OR4 (N21893, N21886, N14054, N13457, N21788);
buf BUF1 (N21894, N21885);
xor XOR2 (N21895, N21884, N10134);
buf BUF1 (N21896, N21894);
and AND3 (N21897, N21880, N14195, N16432);
buf BUF1 (N21898, N21893);
nand NAND4 (N21899, N21895, N3402, N8520, N18138);
buf BUF1 (N21900, N21890);
not NOT1 (N21901, N21889);
and AND4 (N21902, N21896, N11009, N2299, N13761);
nor NOR2 (N21903, N21892, N6975);
xor XOR2 (N21904, N21898, N4431);
and AND2 (N21905, N21902, N5146);
or OR4 (N21906, N21903, N8993, N16951, N18330);
not NOT1 (N21907, N21887);
xor XOR2 (N21908, N21907, N18853);
or OR4 (N21909, N21905, N8569, N20604, N8989);
not NOT1 (N21910, N21909);
or OR3 (N21911, N21910, N18408, N4749);
not NOT1 (N21912, N21897);
nand NAND2 (N21913, N21901, N16023);
buf BUF1 (N21914, N21912);
xor XOR2 (N21915, N21877, N12421);
buf BUF1 (N21916, N21908);
buf BUF1 (N21917, N21911);
and AND2 (N21918, N21914, N15725);
xor XOR2 (N21919, N21891, N14924);
or OR4 (N21920, N21904, N10966, N12262, N715);
or OR3 (N21921, N21900, N18019, N2157);
and AND2 (N21922, N21913, N13382);
nor NOR3 (N21923, N21899, N4882, N885);
buf BUF1 (N21924, N21922);
or OR4 (N21925, N21906, N20243, N7832, N11438);
nand NAND3 (N21926, N21920, N11436, N6349);
and AND3 (N21927, N21925, N10116, N9868);
and AND4 (N21928, N21921, N6681, N5119, N5908);
nor NOR4 (N21929, N21927, N19761, N9269, N1120);
or OR3 (N21930, N21919, N4941, N20312);
or OR4 (N21931, N21918, N13933, N5972, N15882);
not NOT1 (N21932, N21926);
and AND4 (N21933, N21929, N3762, N11351, N13924);
nand NAND4 (N21934, N21931, N20256, N7088, N14165);
not NOT1 (N21935, N21915);
not NOT1 (N21936, N21930);
xor XOR2 (N21937, N21936, N9227);
nor NOR3 (N21938, N21933, N18630, N20369);
nand NAND3 (N21939, N21932, N5418, N5161);
nand NAND2 (N21940, N21935, N156);
buf BUF1 (N21941, N21938);
and AND3 (N21942, N21940, N6166, N7780);
nor NOR3 (N21943, N21923, N6282, N5397);
or OR2 (N21944, N21916, N17307);
or OR3 (N21945, N21942, N4902, N11751);
nor NOR3 (N21946, N21944, N21405, N11318);
or OR2 (N21947, N21924, N20685);
xor XOR2 (N21948, N21947, N12305);
or OR2 (N21949, N21941, N11830);
buf BUF1 (N21950, N21939);
buf BUF1 (N21951, N21937);
nor NOR2 (N21952, N21950, N9714);
and AND2 (N21953, N21917, N15308);
nand NAND4 (N21954, N21943, N18257, N10396, N7487);
not NOT1 (N21955, N21946);
not NOT1 (N21956, N21954);
buf BUF1 (N21957, N21952);
or OR2 (N21958, N21955, N4381);
nor NOR4 (N21959, N21957, N4705, N13394, N21027);
nor NOR3 (N21960, N21945, N3227, N6701);
and AND2 (N21961, N21951, N66);
not NOT1 (N21962, N21953);
or OR4 (N21963, N21960, N20962, N10423, N13471);
nand NAND2 (N21964, N21928, N13811);
and AND3 (N21965, N21948, N205, N11103);
or OR3 (N21966, N21965, N7350, N10328);
buf BUF1 (N21967, N21961);
or OR3 (N21968, N21959, N2779, N14421);
or OR2 (N21969, N21962, N15983);
buf BUF1 (N21970, N21958);
nor NOR4 (N21971, N21970, N19770, N5513, N16700);
and AND2 (N21972, N21934, N7768);
nor NOR4 (N21973, N21956, N17955, N18408, N16753);
nand NAND4 (N21974, N21971, N11849, N15937, N6676);
nand NAND3 (N21975, N21966, N20039, N11610);
buf BUF1 (N21976, N21963);
buf BUF1 (N21977, N21969);
not NOT1 (N21978, N21974);
nor NOR3 (N21979, N21973, N4221, N17153);
and AND4 (N21980, N21949, N18707, N14315, N7656);
or OR3 (N21981, N21968, N18845, N11311);
or OR2 (N21982, N21981, N12296);
xor XOR2 (N21983, N21975, N3844);
and AND3 (N21984, N21978, N8891, N6220);
nor NOR2 (N21985, N21979, N7556);
not NOT1 (N21986, N21972);
xor XOR2 (N21987, N21964, N5070);
or OR4 (N21988, N21986, N12085, N14862, N10433);
buf BUF1 (N21989, N21980);
xor XOR2 (N21990, N21989, N21804);
not NOT1 (N21991, N21990);
nor NOR3 (N21992, N21984, N10808, N11866);
nand NAND2 (N21993, N21987, N9904);
nand NAND2 (N21994, N21992, N9212);
nand NAND2 (N21995, N21994, N207);
xor XOR2 (N21996, N21988, N4793);
nand NAND3 (N21997, N21993, N17179, N18185);
not NOT1 (N21998, N21967);
or OR3 (N21999, N21991, N15985, N13652);
nand NAND4 (N22000, N21998, N8405, N10843, N8118);
xor XOR2 (N22001, N22000, N15198);
not NOT1 (N22002, N21983);
not NOT1 (N22003, N21995);
not NOT1 (N22004, N21999);
buf BUF1 (N22005, N22002);
nor NOR3 (N22006, N22001, N19195, N2043);
nand NAND3 (N22007, N22003, N270, N11664);
buf BUF1 (N22008, N21976);
and AND4 (N22009, N22006, N14113, N7293, N3628);
nand NAND2 (N22010, N22008, N18308);
nand NAND3 (N22011, N22010, N11347, N3474);
or OR4 (N22012, N22004, N12096, N1487, N1961);
nand NAND4 (N22013, N21977, N10564, N5051, N19834);
xor XOR2 (N22014, N22009, N12849);
buf BUF1 (N22015, N21985);
not NOT1 (N22016, N22013);
and AND2 (N22017, N22015, N4517);
and AND3 (N22018, N21982, N14194, N6100);
buf BUF1 (N22019, N22007);
not NOT1 (N22020, N22017);
nor NOR4 (N22021, N21996, N15134, N8217, N13825);
buf BUF1 (N22022, N22014);
xor XOR2 (N22023, N21997, N4558);
not NOT1 (N22024, N22020);
nand NAND4 (N22025, N22012, N20307, N14897, N17185);
nand NAND4 (N22026, N22019, N18806, N15097, N6419);
nand NAND3 (N22027, N22005, N6004, N16372);
and AND2 (N22028, N22023, N5310);
buf BUF1 (N22029, N22028);
and AND2 (N22030, N22025, N11193);
xor XOR2 (N22031, N22027, N8869);
and AND2 (N22032, N22026, N14725);
not NOT1 (N22033, N22031);
nor NOR3 (N22034, N22029, N22018, N22000);
or OR3 (N22035, N6970, N10774, N20151);
xor XOR2 (N22036, N22033, N3648);
and AND3 (N22037, N22034, N18286, N16865);
not NOT1 (N22038, N22030);
xor XOR2 (N22039, N22032, N1141);
or OR3 (N22040, N22035, N20263, N15460);
not NOT1 (N22041, N22016);
and AND2 (N22042, N22021, N761);
nor NOR2 (N22043, N22022, N8909);
and AND3 (N22044, N22038, N9813, N2026);
nand NAND4 (N22045, N22036, N13388, N18224, N14701);
buf BUF1 (N22046, N22045);
buf BUF1 (N22047, N22044);
nor NOR4 (N22048, N22011, N261, N13932, N5895);
buf BUF1 (N22049, N22042);
and AND3 (N22050, N22039, N11122, N13405);
nand NAND4 (N22051, N22041, N14006, N19903, N2340);
not NOT1 (N22052, N22047);
nor NOR3 (N22053, N22050, N10232, N10572);
xor XOR2 (N22054, N22043, N1570);
not NOT1 (N22055, N22052);
not NOT1 (N22056, N22037);
not NOT1 (N22057, N22053);
buf BUF1 (N22058, N22049);
not NOT1 (N22059, N22040);
nand NAND3 (N22060, N22046, N17372, N13086);
and AND4 (N22061, N22051, N18647, N18420, N7799);
or OR2 (N22062, N22048, N4560);
buf BUF1 (N22063, N22054);
xor XOR2 (N22064, N22057, N14053);
nor NOR2 (N22065, N22064, N21165);
buf BUF1 (N22066, N22024);
or OR3 (N22067, N22063, N243, N9850);
buf BUF1 (N22068, N22065);
and AND2 (N22069, N22062, N16112);
xor XOR2 (N22070, N22066, N6639);
nor NOR2 (N22071, N22067, N20697);
nand NAND3 (N22072, N22069, N20361, N6261);
nand NAND4 (N22073, N22060, N21964, N9289, N1537);
not NOT1 (N22074, N22059);
or OR2 (N22075, N22071, N8505);
nor NOR4 (N22076, N22072, N10542, N8773, N11729);
xor XOR2 (N22077, N22070, N18885);
not NOT1 (N22078, N22076);
nand NAND4 (N22079, N22078, N6894, N16187, N13018);
nor NOR3 (N22080, N22075, N685, N1887);
and AND4 (N22081, N22061, N15345, N12193, N17972);
not NOT1 (N22082, N22073);
nand NAND3 (N22083, N22055, N15185, N13095);
not NOT1 (N22084, N22082);
nand NAND2 (N22085, N22084, N7186);
buf BUF1 (N22086, N22083);
or OR3 (N22087, N22056, N2498, N20951);
nand NAND3 (N22088, N22085, N2485, N18147);
not NOT1 (N22089, N22087);
nor NOR4 (N22090, N22058, N15199, N15964, N3861);
nand NAND4 (N22091, N22080, N19435, N1442, N2153);
nand NAND4 (N22092, N22077, N5236, N1051, N1902);
xor XOR2 (N22093, N22068, N11365);
buf BUF1 (N22094, N22079);
nor NOR4 (N22095, N22086, N9688, N3132, N543);
not NOT1 (N22096, N22091);
xor XOR2 (N22097, N22088, N16883);
not NOT1 (N22098, N22089);
buf BUF1 (N22099, N22095);
or OR4 (N22100, N22093, N21361, N14639, N16594);
nand NAND4 (N22101, N22099, N6717, N17602, N12352);
nand NAND4 (N22102, N22090, N19630, N11905, N3912);
nand NAND2 (N22103, N22096, N20511);
and AND2 (N22104, N22103, N2604);
and AND4 (N22105, N22074, N8835, N3189, N2153);
or OR3 (N22106, N22098, N14481, N12183);
xor XOR2 (N22107, N22105, N5691);
not NOT1 (N22108, N22101);
not NOT1 (N22109, N22107);
nand NAND2 (N22110, N22092, N16987);
nor NOR2 (N22111, N22102, N18857);
nand NAND2 (N22112, N22081, N905);
nand NAND3 (N22113, N22100, N15898, N19179);
buf BUF1 (N22114, N22094);
and AND2 (N22115, N22110, N7663);
or OR3 (N22116, N22111, N18570, N2668);
xor XOR2 (N22117, N22114, N11409);
or OR4 (N22118, N22106, N14868, N11688, N2352);
or OR3 (N22119, N22116, N7739, N8261);
and AND3 (N22120, N22118, N315, N17774);
and AND4 (N22121, N22117, N2802, N11260, N10548);
or OR4 (N22122, N22104, N20385, N19614, N10431);
not NOT1 (N22123, N22097);
and AND3 (N22124, N22109, N3320, N21937);
or OR2 (N22125, N22124, N1020);
or OR4 (N22126, N22108, N17474, N14587, N16639);
or OR4 (N22127, N22125, N706, N7092, N20842);
not NOT1 (N22128, N22112);
nor NOR3 (N22129, N22122, N20750, N4505);
not NOT1 (N22130, N22113);
nor NOR2 (N22131, N22128, N21722);
not NOT1 (N22132, N22119);
not NOT1 (N22133, N22123);
or OR3 (N22134, N22126, N14359, N9666);
nand NAND2 (N22135, N22121, N17918);
and AND2 (N22136, N22127, N14606);
nor NOR3 (N22137, N22115, N8251, N6901);
nand NAND3 (N22138, N22133, N6551, N12822);
or OR4 (N22139, N22129, N18969, N10191, N21205);
or OR3 (N22140, N22131, N9784, N16456);
buf BUF1 (N22141, N22137);
not NOT1 (N22142, N22136);
nor NOR3 (N22143, N22142, N15612, N20898);
and AND3 (N22144, N22138, N12359, N803);
nand NAND3 (N22145, N22139, N4140, N14711);
nor NOR2 (N22146, N22144, N19511);
not NOT1 (N22147, N22134);
buf BUF1 (N22148, N22141);
or OR3 (N22149, N22132, N10390, N6087);
and AND4 (N22150, N22145, N19782, N483, N11664);
and AND2 (N22151, N22120, N12295);
buf BUF1 (N22152, N22148);
and AND4 (N22153, N22149, N8075, N3750, N17401);
nor NOR2 (N22154, N22140, N7001);
or OR4 (N22155, N22130, N16846, N9020, N12600);
not NOT1 (N22156, N22150);
buf BUF1 (N22157, N22151);
not NOT1 (N22158, N22135);
not NOT1 (N22159, N22155);
nor NOR3 (N22160, N22154, N21694, N18262);
nand NAND2 (N22161, N22156, N10616);
not NOT1 (N22162, N22143);
nand NAND3 (N22163, N22152, N21815, N18086);
not NOT1 (N22164, N22146);
xor XOR2 (N22165, N22164, N7307);
nand NAND2 (N22166, N22147, N4505);
nor NOR2 (N22167, N22158, N1517);
and AND3 (N22168, N22166, N3895, N12400);
xor XOR2 (N22169, N22161, N13678);
and AND4 (N22170, N22157, N10372, N13098, N20682);
or OR3 (N22171, N22163, N14451, N1476);
not NOT1 (N22172, N22169);
and AND2 (N22173, N22172, N6213);
or OR3 (N22174, N22159, N2533, N14953);
and AND4 (N22175, N22173, N8031, N5233, N3175);
and AND2 (N22176, N22160, N1208);
buf BUF1 (N22177, N22175);
buf BUF1 (N22178, N22174);
xor XOR2 (N22179, N22165, N22028);
not NOT1 (N22180, N22170);
xor XOR2 (N22181, N22180, N9820);
or OR2 (N22182, N22153, N15723);
xor XOR2 (N22183, N22168, N16990);
xor XOR2 (N22184, N22178, N10982);
nand NAND2 (N22185, N22177, N2723);
nand NAND3 (N22186, N22184, N3382, N20601);
and AND2 (N22187, N22181, N1261);
not NOT1 (N22188, N22182);
nand NAND3 (N22189, N22188, N10204, N11112);
not NOT1 (N22190, N22162);
nor NOR4 (N22191, N22187, N10490, N8589, N18586);
nand NAND4 (N22192, N22186, N15495, N16463, N16323);
nor NOR3 (N22193, N22167, N8186, N7728);
buf BUF1 (N22194, N22189);
nand NAND2 (N22195, N22190, N21906);
buf BUF1 (N22196, N22176);
or OR3 (N22197, N22183, N8578, N9346);
or OR2 (N22198, N22185, N13390);
and AND4 (N22199, N22196, N4089, N6688, N19891);
not NOT1 (N22200, N22199);
buf BUF1 (N22201, N22193);
xor XOR2 (N22202, N22198, N674);
xor XOR2 (N22203, N22179, N11342);
buf BUF1 (N22204, N22203);
nor NOR3 (N22205, N22204, N16087, N5936);
buf BUF1 (N22206, N22195);
buf BUF1 (N22207, N22194);
and AND4 (N22208, N22192, N3258, N14907, N3885);
buf BUF1 (N22209, N22205);
or OR3 (N22210, N22207, N19851, N21881);
nand NAND4 (N22211, N22191, N4786, N17933, N5586);
xor XOR2 (N22212, N22211, N10358);
nand NAND3 (N22213, N22200, N6452, N11372);
nand NAND4 (N22214, N22210, N16683, N2431, N20047);
and AND2 (N22215, N22206, N146);
nand NAND2 (N22216, N22214, N18923);
and AND4 (N22217, N22201, N10936, N20181, N20697);
or OR2 (N22218, N22202, N8593);
buf BUF1 (N22219, N22212);
nand NAND3 (N22220, N22218, N12461, N11615);
xor XOR2 (N22221, N22213, N17251);
or OR2 (N22222, N22217, N7969);
xor XOR2 (N22223, N22219, N747);
and AND4 (N22224, N22197, N15856, N232, N6020);
or OR4 (N22225, N22224, N5473, N7026, N4832);
or OR3 (N22226, N22225, N18193, N17475);
buf BUF1 (N22227, N22223);
and AND4 (N22228, N22209, N10334, N10727, N12328);
not NOT1 (N22229, N22208);
xor XOR2 (N22230, N22220, N15903);
and AND3 (N22231, N22221, N11488, N5492);
xor XOR2 (N22232, N22226, N3350);
nand NAND2 (N22233, N22231, N7212);
or OR4 (N22234, N22233, N3419, N8536, N21674);
and AND2 (N22235, N22222, N6975);
buf BUF1 (N22236, N22235);
nor NOR4 (N22237, N22227, N17261, N2722, N18429);
buf BUF1 (N22238, N22215);
xor XOR2 (N22239, N22216, N12292);
or OR2 (N22240, N22229, N8376);
nor NOR3 (N22241, N22228, N21756, N9599);
not NOT1 (N22242, N22237);
or OR3 (N22243, N22171, N9042, N2798);
or OR4 (N22244, N22240, N21838, N10473, N8363);
buf BUF1 (N22245, N22238);
and AND4 (N22246, N22236, N15099, N14833, N18895);
not NOT1 (N22247, N22245);
not NOT1 (N22248, N22241);
not NOT1 (N22249, N22243);
xor XOR2 (N22250, N22248, N19880);
buf BUF1 (N22251, N22239);
not NOT1 (N22252, N22250);
nor NOR2 (N22253, N22232, N7727);
nor NOR3 (N22254, N22242, N12041, N15268);
not NOT1 (N22255, N22249);
xor XOR2 (N22256, N22253, N8332);
nand NAND4 (N22257, N22256, N7353, N5021, N4404);
not NOT1 (N22258, N22251);
and AND2 (N22259, N22257, N14685);
nor NOR4 (N22260, N22234, N11377, N8764, N8556);
buf BUF1 (N22261, N22247);
and AND4 (N22262, N22255, N6316, N10999, N9317);
or OR2 (N22263, N22230, N21022);
xor XOR2 (N22264, N22252, N12312);
and AND2 (N22265, N22263, N17833);
xor XOR2 (N22266, N22246, N7320);
nor NOR4 (N22267, N22264, N821, N18262, N2528);
not NOT1 (N22268, N22244);
nor NOR3 (N22269, N22260, N8593, N12928);
xor XOR2 (N22270, N22269, N14017);
xor XOR2 (N22271, N22265, N21998);
nand NAND3 (N22272, N22270, N18164, N22057);
xor XOR2 (N22273, N22259, N21759);
or OR4 (N22274, N22262, N18464, N16776, N15060);
not NOT1 (N22275, N22268);
and AND4 (N22276, N22275, N5073, N8650, N13710);
and AND3 (N22277, N22266, N22191, N19569);
nor NOR4 (N22278, N22277, N17760, N894, N10306);
nand NAND2 (N22279, N22271, N7703);
and AND3 (N22280, N22258, N5294, N17781);
or OR2 (N22281, N22278, N3199);
nor NOR2 (N22282, N22261, N18229);
xor XOR2 (N22283, N22282, N10303);
nand NAND2 (N22284, N22279, N19450);
xor XOR2 (N22285, N22267, N4621);
nand NAND2 (N22286, N22272, N13379);
not NOT1 (N22287, N22286);
and AND4 (N22288, N22254, N13330, N14860, N6928);
nor NOR2 (N22289, N22285, N15827);
or OR2 (N22290, N22289, N18418);
and AND3 (N22291, N22283, N14667, N1727);
or OR3 (N22292, N22284, N19277, N15247);
not NOT1 (N22293, N22287);
not NOT1 (N22294, N22281);
nand NAND3 (N22295, N22288, N16819, N3344);
or OR4 (N22296, N22290, N618, N6304, N6217);
xor XOR2 (N22297, N22293, N4295);
or OR4 (N22298, N22280, N897, N4662, N5208);
not NOT1 (N22299, N22294);
not NOT1 (N22300, N22273);
nand NAND2 (N22301, N22298, N18909);
nor NOR2 (N22302, N22276, N15650);
and AND4 (N22303, N22291, N20084, N20049, N19212);
and AND4 (N22304, N22299, N19992, N2993, N16514);
buf BUF1 (N22305, N22295);
nor NOR3 (N22306, N22301, N10934, N14177);
nor NOR4 (N22307, N22305, N7284, N3082, N10065);
and AND3 (N22308, N22292, N447, N17657);
xor XOR2 (N22309, N22307, N18550);
nor NOR2 (N22310, N22300, N5689);
xor XOR2 (N22311, N22304, N847);
and AND4 (N22312, N22297, N8224, N9015, N16762);
or OR2 (N22313, N22310, N5551);
not NOT1 (N22314, N22303);
not NOT1 (N22315, N22312);
buf BUF1 (N22316, N22296);
or OR4 (N22317, N22315, N6370, N3177, N4035);
or OR2 (N22318, N22308, N14088);
not NOT1 (N22319, N22302);
buf BUF1 (N22320, N22306);
and AND2 (N22321, N22309, N17458);
not NOT1 (N22322, N22317);
nor NOR3 (N22323, N22319, N20833, N4825);
xor XOR2 (N22324, N22318, N11225);
nand NAND4 (N22325, N22314, N15553, N14356, N21111);
nor NOR4 (N22326, N22320, N18615, N2431, N15553);
not NOT1 (N22327, N22321);
nand NAND2 (N22328, N22322, N8179);
buf BUF1 (N22329, N22313);
nor NOR2 (N22330, N22328, N12590);
and AND3 (N22331, N22311, N20511, N6621);
or OR4 (N22332, N22329, N3128, N10941, N2888);
not NOT1 (N22333, N22332);
nand NAND3 (N22334, N22274, N5611, N14564);
nand NAND3 (N22335, N22334, N13539, N13254);
not NOT1 (N22336, N22327);
buf BUF1 (N22337, N22335);
not NOT1 (N22338, N22323);
and AND4 (N22339, N22330, N17711, N65, N4807);
and AND4 (N22340, N22316, N3442, N1678, N14893);
buf BUF1 (N22341, N22333);
and AND3 (N22342, N22340, N10378, N4122);
or OR4 (N22343, N22325, N7038, N3405, N10882);
nand NAND3 (N22344, N22326, N21241, N8256);
nand NAND3 (N22345, N22338, N4112, N20496);
nor NOR4 (N22346, N22345, N10130, N5850, N1356);
xor XOR2 (N22347, N22324, N383);
and AND2 (N22348, N22339, N4334);
or OR3 (N22349, N22331, N16765, N15080);
and AND3 (N22350, N22349, N18657, N2149);
not NOT1 (N22351, N22344);
or OR3 (N22352, N22346, N439, N8819);
xor XOR2 (N22353, N22351, N1422);
not NOT1 (N22354, N22350);
nand NAND3 (N22355, N22336, N16842, N19884);
nor NOR4 (N22356, N22352, N18141, N9223, N6414);
xor XOR2 (N22357, N22342, N18104);
or OR2 (N22358, N22341, N8630);
buf BUF1 (N22359, N22348);
nor NOR2 (N22360, N22358, N3352);
nor NOR4 (N22361, N22359, N5720, N6908, N22314);
not NOT1 (N22362, N22353);
buf BUF1 (N22363, N22337);
and AND3 (N22364, N22360, N7455, N18555);
xor XOR2 (N22365, N22347, N13461);
buf BUF1 (N22366, N22362);
or OR3 (N22367, N22363, N11132, N16999);
nand NAND3 (N22368, N22367, N7125, N4052);
nor NOR4 (N22369, N22343, N14153, N208, N7479);
buf BUF1 (N22370, N22364);
xor XOR2 (N22371, N22369, N8239);
buf BUF1 (N22372, N22355);
not NOT1 (N22373, N22365);
nor NOR3 (N22374, N22357, N16370, N7551);
or OR4 (N22375, N22356, N11587, N20310, N13149);
buf BUF1 (N22376, N22354);
or OR4 (N22377, N22375, N8621, N10428, N10672);
not NOT1 (N22378, N22371);
xor XOR2 (N22379, N22368, N7127);
or OR3 (N22380, N22374, N1135, N16752);
or OR4 (N22381, N22373, N7589, N15947, N16458);
nand NAND4 (N22382, N22372, N5418, N338, N4593);
buf BUF1 (N22383, N22377);
nor NOR4 (N22384, N22370, N12161, N14838, N8268);
xor XOR2 (N22385, N22361, N7488);
and AND4 (N22386, N22379, N13545, N933, N979);
xor XOR2 (N22387, N22384, N7149);
xor XOR2 (N22388, N22380, N2367);
not NOT1 (N22389, N22376);
nand NAND4 (N22390, N22388, N14366, N6114, N8916);
not NOT1 (N22391, N22383);
and AND3 (N22392, N22382, N18912, N7396);
nor NOR2 (N22393, N22381, N10036);
nand NAND3 (N22394, N22366, N14328, N4612);
or OR4 (N22395, N22394, N6283, N20538, N18481);
or OR2 (N22396, N22387, N20412);
not NOT1 (N22397, N22392);
buf BUF1 (N22398, N22397);
xor XOR2 (N22399, N22378, N16490);
nand NAND3 (N22400, N22393, N20190, N15087);
xor XOR2 (N22401, N22396, N14431);
or OR4 (N22402, N22385, N21112, N2330, N7906);
nor NOR2 (N22403, N22401, N20843);
nor NOR3 (N22404, N22395, N12828, N4274);
not NOT1 (N22405, N22400);
nand NAND2 (N22406, N22398, N1234);
or OR2 (N22407, N22402, N4860);
and AND3 (N22408, N22386, N4821, N9711);
buf BUF1 (N22409, N22389);
and AND4 (N22410, N22404, N22254, N5272, N14320);
buf BUF1 (N22411, N22408);
nand NAND4 (N22412, N22391, N19119, N15309, N14212);
buf BUF1 (N22413, N22410);
or OR3 (N22414, N22412, N11410, N12272);
buf BUF1 (N22415, N22411);
nand NAND3 (N22416, N22414, N14301, N3177);
buf BUF1 (N22417, N22405);
xor XOR2 (N22418, N22413, N2928);
not NOT1 (N22419, N22416);
and AND4 (N22420, N22409, N6679, N16819, N10293);
not NOT1 (N22421, N22417);
nor NOR4 (N22422, N22406, N7131, N17831, N15884);
nor NOR3 (N22423, N22419, N3227, N9094);
or OR2 (N22424, N22420, N10172);
nor NOR2 (N22425, N22421, N13701);
and AND4 (N22426, N22403, N15506, N12380, N20271);
xor XOR2 (N22427, N22424, N13089);
nand NAND2 (N22428, N22423, N8035);
or OR3 (N22429, N22427, N17860, N3938);
not NOT1 (N22430, N22390);
nor NOR4 (N22431, N22428, N1787, N5849, N18523);
xor XOR2 (N22432, N22418, N8948);
or OR4 (N22433, N22429, N15628, N16119, N9176);
or OR4 (N22434, N22431, N14045, N12720, N6372);
not NOT1 (N22435, N22422);
xor XOR2 (N22436, N22434, N4465);
nand NAND4 (N22437, N22399, N6524, N3857, N15521);
nor NOR2 (N22438, N22436, N6873);
nand NAND4 (N22439, N22435, N20879, N1135, N2077);
or OR4 (N22440, N22439, N9323, N13672, N20900);
buf BUF1 (N22441, N22430);
nand NAND3 (N22442, N22426, N5105, N21256);
nor NOR4 (N22443, N22441, N12564, N4491, N19747);
and AND3 (N22444, N22407, N9695, N16015);
xor XOR2 (N22445, N22432, N14820);
xor XOR2 (N22446, N22425, N21664);
nor NOR3 (N22447, N22440, N19112, N20066);
xor XOR2 (N22448, N22433, N9251);
buf BUF1 (N22449, N22448);
not NOT1 (N22450, N22442);
or OR2 (N22451, N22445, N20473);
buf BUF1 (N22452, N22447);
or OR4 (N22453, N22449, N3553, N6480, N11674);
nand NAND4 (N22454, N22451, N2319, N11503, N14398);
nor NOR4 (N22455, N22438, N13684, N22037, N13666);
nand NAND4 (N22456, N22450, N2499, N20440, N3775);
xor XOR2 (N22457, N22437, N182);
not NOT1 (N22458, N22456);
not NOT1 (N22459, N22458);
and AND3 (N22460, N22457, N14587, N4280);
nor NOR2 (N22461, N22453, N17047);
not NOT1 (N22462, N22446);
buf BUF1 (N22463, N22444);
xor XOR2 (N22464, N22443, N14160);
or OR4 (N22465, N22452, N20156, N19765, N21189);
or OR3 (N22466, N22460, N14738, N4134);
nand NAND2 (N22467, N22455, N7310);
or OR2 (N22468, N22463, N2763);
buf BUF1 (N22469, N22454);
or OR4 (N22470, N22464, N6688, N16339, N7979);
and AND3 (N22471, N22459, N3900, N11262);
or OR4 (N22472, N22468, N81, N14492, N17725);
buf BUF1 (N22473, N22415);
buf BUF1 (N22474, N22462);
xor XOR2 (N22475, N22474, N9000);
xor XOR2 (N22476, N22469, N15178);
xor XOR2 (N22477, N22472, N17015);
nor NOR4 (N22478, N22465, N20631, N10172, N18154);
nand NAND2 (N22479, N22477, N1088);
nor NOR3 (N22480, N22466, N6974, N21237);
nor NOR3 (N22481, N22478, N11534, N19674);
xor XOR2 (N22482, N22470, N19739);
nand NAND2 (N22483, N22482, N12100);
or OR2 (N22484, N22479, N7589);
not NOT1 (N22485, N22476);
buf BUF1 (N22486, N22473);
nand NAND2 (N22487, N22471, N9675);
not NOT1 (N22488, N22484);
not NOT1 (N22489, N22486);
nand NAND2 (N22490, N22487, N12543);
or OR4 (N22491, N22480, N22115, N12458, N10498);
xor XOR2 (N22492, N22491, N15209);
nor NOR2 (N22493, N22467, N4092);
buf BUF1 (N22494, N22461);
buf BUF1 (N22495, N22475);
nor NOR3 (N22496, N22490, N635, N16871);
xor XOR2 (N22497, N22493, N7366);
and AND4 (N22498, N22481, N3984, N6268, N16352);
nand NAND2 (N22499, N22489, N20241);
nand NAND4 (N22500, N22495, N19531, N3331, N20931);
xor XOR2 (N22501, N22488, N1512);
or OR2 (N22502, N22499, N16204);
nor NOR3 (N22503, N22494, N12960, N9075);
buf BUF1 (N22504, N22500);
nand NAND3 (N22505, N22498, N16110, N7801);
xor XOR2 (N22506, N22496, N16214);
and AND3 (N22507, N22504, N6328, N22489);
or OR2 (N22508, N22502, N11142);
or OR4 (N22509, N22503, N5560, N16935, N3096);
nand NAND2 (N22510, N22492, N20832);
not NOT1 (N22511, N22509);
buf BUF1 (N22512, N22485);
and AND3 (N22513, N22505, N3428, N13756);
buf BUF1 (N22514, N22497);
not NOT1 (N22515, N22506);
nand NAND2 (N22516, N22513, N19890);
buf BUF1 (N22517, N22515);
xor XOR2 (N22518, N22483, N15342);
nor NOR4 (N22519, N22516, N11372, N8406, N4922);
buf BUF1 (N22520, N22507);
and AND3 (N22521, N22512, N17219, N13442);
not NOT1 (N22522, N22508);
nand NAND2 (N22523, N22518, N22521);
nand NAND3 (N22524, N21147, N8906, N6359);
not NOT1 (N22525, N22523);
nand NAND4 (N22526, N22524, N21556, N1492, N18321);
xor XOR2 (N22527, N22517, N1985);
nor NOR4 (N22528, N22527, N12993, N4678, N6515);
not NOT1 (N22529, N22519);
buf BUF1 (N22530, N22526);
nand NAND3 (N22531, N22520, N13010, N16416);
and AND4 (N22532, N22529, N6191, N10228, N7370);
nand NAND3 (N22533, N22525, N434, N20126);
buf BUF1 (N22534, N22522);
xor XOR2 (N22535, N22501, N17039);
or OR3 (N22536, N22528, N11704, N21215);
or OR3 (N22537, N22535, N8927, N19260);
xor XOR2 (N22538, N22530, N13105);
not NOT1 (N22539, N22511);
nor NOR3 (N22540, N22539, N22307, N15647);
or OR4 (N22541, N22534, N18330, N9133, N16420);
not NOT1 (N22542, N22510);
and AND3 (N22543, N22540, N5032, N13479);
nand NAND2 (N22544, N22532, N6815);
nor NOR4 (N22545, N22543, N1202, N18941, N21492);
not NOT1 (N22546, N22542);
xor XOR2 (N22547, N22541, N2824);
nor NOR2 (N22548, N22531, N4605);
nand NAND2 (N22549, N22514, N1466);
xor XOR2 (N22550, N22547, N6912);
not NOT1 (N22551, N22548);
nor NOR2 (N22552, N22536, N8574);
nand NAND2 (N22553, N22545, N4474);
nor NOR3 (N22554, N22544, N19197, N5948);
buf BUF1 (N22555, N22553);
not NOT1 (N22556, N22555);
xor XOR2 (N22557, N22537, N9759);
nor NOR4 (N22558, N22549, N19435, N13735, N19408);
and AND3 (N22559, N22546, N4907, N2765);
not NOT1 (N22560, N22552);
nor NOR3 (N22561, N22551, N13854, N12023);
buf BUF1 (N22562, N22557);
nor NOR3 (N22563, N22554, N12681, N20157);
nor NOR3 (N22564, N22562, N14383, N10946);
or OR3 (N22565, N22558, N19769, N17020);
xor XOR2 (N22566, N22538, N18699);
xor XOR2 (N22567, N22566, N3190);
xor XOR2 (N22568, N22563, N13522);
or OR2 (N22569, N22556, N15137);
not NOT1 (N22570, N22565);
not NOT1 (N22571, N22568);
and AND4 (N22572, N22561, N19341, N15342, N7196);
buf BUF1 (N22573, N22572);
nor NOR4 (N22574, N22570, N20416, N18226, N12859);
nand NAND4 (N22575, N22550, N1060, N13370, N13823);
nand NAND4 (N22576, N22533, N12959, N11828, N5532);
not NOT1 (N22577, N22571);
and AND3 (N22578, N22564, N6489, N8648);
and AND3 (N22579, N22569, N10028, N14768);
nor NOR2 (N22580, N22560, N19505);
nor NOR4 (N22581, N22559, N21090, N17544, N4559);
or OR4 (N22582, N22567, N21412, N6572, N6563);
and AND2 (N22583, N22580, N5606);
or OR2 (N22584, N22576, N21594);
not NOT1 (N22585, N22575);
buf BUF1 (N22586, N22573);
and AND2 (N22587, N22585, N21398);
buf BUF1 (N22588, N22578);
xor XOR2 (N22589, N22579, N212);
and AND4 (N22590, N22586, N4896, N4940, N3035);
not NOT1 (N22591, N22584);
not NOT1 (N22592, N22582);
not NOT1 (N22593, N22592);
and AND3 (N22594, N22588, N6585, N4704);
not NOT1 (N22595, N22594);
xor XOR2 (N22596, N22595, N6148);
or OR3 (N22597, N22577, N9366, N14380);
or OR2 (N22598, N22589, N4719);
buf BUF1 (N22599, N22581);
and AND3 (N22600, N22598, N14463, N19821);
nand NAND4 (N22601, N22600, N6066, N6825, N7023);
buf BUF1 (N22602, N22596);
nor NOR3 (N22603, N22587, N8928, N19722);
not NOT1 (N22604, N22597);
not NOT1 (N22605, N22602);
nor NOR2 (N22606, N22599, N2791);
xor XOR2 (N22607, N22603, N778);
buf BUF1 (N22608, N22591);
xor XOR2 (N22609, N22601, N3715);
and AND2 (N22610, N22593, N18735);
and AND2 (N22611, N22606, N14598);
nor NOR3 (N22612, N22607, N20725, N18178);
and AND4 (N22613, N22608, N13935, N6595, N9005);
nor NOR3 (N22614, N22610, N16860, N16844);
buf BUF1 (N22615, N22614);
and AND4 (N22616, N22583, N22011, N5973, N11290);
and AND3 (N22617, N22609, N10816, N2332);
nand NAND4 (N22618, N22613, N11367, N11525, N7491);
and AND3 (N22619, N22616, N4812, N9793);
nand NAND2 (N22620, N22617, N18475);
xor XOR2 (N22621, N22620, N19375);
and AND4 (N22622, N22621, N19731, N18843, N17929);
xor XOR2 (N22623, N22604, N17703);
buf BUF1 (N22624, N22574);
nor NOR2 (N22625, N22590, N285);
or OR3 (N22626, N22624, N11438, N12965);
or OR3 (N22627, N22618, N14426, N19171);
buf BUF1 (N22628, N22619);
nand NAND4 (N22629, N22612, N7023, N3909, N10729);
nand NAND4 (N22630, N22615, N2145, N2524, N7272);
xor XOR2 (N22631, N22625, N18495);
buf BUF1 (N22632, N22628);
nand NAND2 (N22633, N22632, N9607);
buf BUF1 (N22634, N22627);
and AND2 (N22635, N22622, N22596);
not NOT1 (N22636, N22631);
nor NOR4 (N22637, N22634, N14941, N5547, N8693);
buf BUF1 (N22638, N22635);
not NOT1 (N22639, N22623);
nand NAND2 (N22640, N22639, N8384);
xor XOR2 (N22641, N22630, N22351);
buf BUF1 (N22642, N22640);
buf BUF1 (N22643, N22605);
not NOT1 (N22644, N22641);
nor NOR4 (N22645, N22644, N10725, N4452, N2659);
and AND4 (N22646, N22643, N22425, N19704, N7933);
not NOT1 (N22647, N22646);
and AND4 (N22648, N22647, N15119, N9953, N15912);
or OR3 (N22649, N22642, N6596, N18376);
or OR4 (N22650, N22636, N3646, N110, N5777);
or OR2 (N22651, N22611, N20702);
or OR4 (N22652, N22626, N21649, N17445, N22089);
nand NAND3 (N22653, N22637, N16064, N5600);
or OR3 (N22654, N22652, N5841, N20831);
not NOT1 (N22655, N22645);
nand NAND2 (N22656, N22654, N10257);
nand NAND2 (N22657, N22656, N16022);
not NOT1 (N22658, N22633);
or OR2 (N22659, N22638, N16251);
xor XOR2 (N22660, N22651, N20017);
buf BUF1 (N22661, N22657);
nor NOR2 (N22662, N22658, N19125);
or OR3 (N22663, N22660, N1469, N18);
not NOT1 (N22664, N22648);
not NOT1 (N22665, N22653);
nor NOR2 (N22666, N22649, N6368);
or OR2 (N22667, N22665, N3741);
not NOT1 (N22668, N22661);
not NOT1 (N22669, N22659);
and AND2 (N22670, N22629, N6741);
not NOT1 (N22671, N22667);
not NOT1 (N22672, N22650);
or OR2 (N22673, N22668, N6322);
buf BUF1 (N22674, N22663);
and AND3 (N22675, N22671, N18996, N16803);
not NOT1 (N22676, N22673);
nand NAND3 (N22677, N22666, N11043, N7719);
buf BUF1 (N22678, N22677);
or OR4 (N22679, N22664, N15112, N21544, N8738);
nor NOR3 (N22680, N22669, N14050, N20868);
and AND4 (N22681, N22676, N22356, N4386, N20217);
nor NOR3 (N22682, N22674, N6645, N18657);
xor XOR2 (N22683, N22681, N17649);
buf BUF1 (N22684, N22680);
or OR3 (N22685, N22662, N10867, N18521);
not NOT1 (N22686, N22678);
xor XOR2 (N22687, N22655, N2498);
nand NAND3 (N22688, N22685, N4489, N1488);
or OR3 (N22689, N22670, N4941, N19557);
nand NAND2 (N22690, N22682, N8066);
not NOT1 (N22691, N22679);
nand NAND2 (N22692, N22683, N15798);
xor XOR2 (N22693, N22690, N17947);
xor XOR2 (N22694, N22692, N8644);
not NOT1 (N22695, N22693);
buf BUF1 (N22696, N22689);
not NOT1 (N22697, N22696);
nand NAND3 (N22698, N22695, N14955, N21472);
xor XOR2 (N22699, N22684, N11410);
and AND4 (N22700, N22697, N11353, N19140, N17893);
buf BUF1 (N22701, N22672);
not NOT1 (N22702, N22686);
or OR3 (N22703, N22687, N17190, N16702);
and AND4 (N22704, N22694, N9255, N516, N22631);
buf BUF1 (N22705, N22691);
buf BUF1 (N22706, N22705);
nor NOR3 (N22707, N22703, N4101, N14930);
or OR3 (N22708, N22698, N1954, N14723);
not NOT1 (N22709, N22708);
and AND3 (N22710, N22709, N16757, N12604);
and AND2 (N22711, N22702, N5213);
nor NOR4 (N22712, N22710, N14706, N15626, N16480);
and AND3 (N22713, N22712, N14581, N15893);
not NOT1 (N22714, N22706);
xor XOR2 (N22715, N22688, N12261);
nor NOR4 (N22716, N22714, N3101, N14174, N22505);
or OR2 (N22717, N22715, N3718);
nand NAND4 (N22718, N22701, N15313, N20844, N4139);
or OR4 (N22719, N22700, N9647, N18256, N6484);
buf BUF1 (N22720, N22704);
and AND4 (N22721, N22717, N15026, N14965, N139);
not NOT1 (N22722, N22675);
nor NOR4 (N22723, N22721, N2959, N15406, N18039);
not NOT1 (N22724, N22720);
not NOT1 (N22725, N22716);
nand NAND4 (N22726, N22707, N17300, N5078, N14620);
buf BUF1 (N22727, N22726);
or OR2 (N22728, N22725, N3759);
or OR4 (N22729, N22722, N1463, N18061, N11465);
not NOT1 (N22730, N22728);
buf BUF1 (N22731, N22713);
and AND2 (N22732, N22699, N9160);
buf BUF1 (N22733, N22718);
not NOT1 (N22734, N22731);
buf BUF1 (N22735, N22719);
or OR2 (N22736, N22727, N5217);
nand NAND2 (N22737, N22723, N13828);
or OR2 (N22738, N22734, N3364);
and AND4 (N22739, N22737, N11077, N1967, N1274);
xor XOR2 (N22740, N22736, N14847);
and AND2 (N22741, N22732, N2313);
buf BUF1 (N22742, N22738);
and AND2 (N22743, N22742, N22617);
not NOT1 (N22744, N22729);
nor NOR3 (N22745, N22743, N19199, N5401);
or OR4 (N22746, N22740, N18040, N9240, N16306);
or OR2 (N22747, N22711, N17864);
not NOT1 (N22748, N22746);
nand NAND3 (N22749, N22735, N8533, N4266);
nor NOR3 (N22750, N22745, N1497, N1729);
not NOT1 (N22751, N22724);
nand NAND3 (N22752, N22741, N6561, N6961);
buf BUF1 (N22753, N22739);
or OR3 (N22754, N22744, N1182, N1298);
or OR3 (N22755, N22754, N13247, N8125);
or OR2 (N22756, N22747, N16176);
or OR4 (N22757, N22748, N17594, N12955, N19415);
nand NAND4 (N22758, N22751, N16564, N1430, N18780);
nor NOR2 (N22759, N22730, N12514);
not NOT1 (N22760, N22750);
and AND3 (N22761, N22758, N5748, N20288);
not NOT1 (N22762, N22733);
buf BUF1 (N22763, N22762);
nor NOR2 (N22764, N22760, N11805);
nor NOR4 (N22765, N22749, N17463, N484, N15003);
not NOT1 (N22766, N22753);
nand NAND2 (N22767, N22763, N14921);
and AND4 (N22768, N22766, N3435, N2727, N1246);
not NOT1 (N22769, N22759);
not NOT1 (N22770, N22764);
xor XOR2 (N22771, N22765, N2345);
and AND4 (N22772, N22756, N10780, N20199, N12363);
not NOT1 (N22773, N22769);
nor NOR4 (N22774, N22770, N13958, N19473, N10529);
xor XOR2 (N22775, N22771, N16008);
not NOT1 (N22776, N22768);
nor NOR3 (N22777, N22773, N4311, N14936);
not NOT1 (N22778, N22755);
nor NOR3 (N22779, N22777, N3349, N2029);
and AND2 (N22780, N22752, N6641);
not NOT1 (N22781, N22757);
xor XOR2 (N22782, N22776, N10636);
buf BUF1 (N22783, N22780);
xor XOR2 (N22784, N22775, N12993);
buf BUF1 (N22785, N22778);
and AND3 (N22786, N22779, N1506, N870);
nor NOR3 (N22787, N22772, N13619, N5509);
xor XOR2 (N22788, N22781, N22278);
xor XOR2 (N22789, N22783, N18961);
and AND3 (N22790, N22761, N14768, N16089);
nor NOR4 (N22791, N22790, N15295, N17126, N18492);
not NOT1 (N22792, N22789);
not NOT1 (N22793, N22786);
buf BUF1 (N22794, N22793);
and AND4 (N22795, N22792, N15105, N6724, N1193);
and AND2 (N22796, N22788, N14419);
and AND2 (N22797, N22774, N11767);
xor XOR2 (N22798, N22791, N12344);
and AND3 (N22799, N22795, N10434, N2225);
buf BUF1 (N22800, N22787);
nand NAND2 (N22801, N22800, N8701);
buf BUF1 (N22802, N22782);
not NOT1 (N22803, N22798);
buf BUF1 (N22804, N22803);
xor XOR2 (N22805, N22799, N7967);
buf BUF1 (N22806, N22802);
not NOT1 (N22807, N22784);
not NOT1 (N22808, N22805);
and AND4 (N22809, N22785, N17785, N18196, N10078);
xor XOR2 (N22810, N22809, N13127);
buf BUF1 (N22811, N22808);
buf BUF1 (N22812, N22806);
or OR4 (N22813, N22794, N21125, N10767, N22633);
xor XOR2 (N22814, N22807, N3693);
not NOT1 (N22815, N22801);
nor NOR2 (N22816, N22796, N17335);
nand NAND4 (N22817, N22810, N6430, N8293, N7416);
nor NOR3 (N22818, N22813, N10765, N7767);
nor NOR3 (N22819, N22804, N853, N13290);
not NOT1 (N22820, N22815);
nand NAND4 (N22821, N22811, N455, N22762, N10703);
xor XOR2 (N22822, N22812, N3157);
xor XOR2 (N22823, N22767, N17494);
nand NAND3 (N22824, N22819, N19125, N13275);
or OR4 (N22825, N22822, N7679, N10536, N667);
buf BUF1 (N22826, N22816);
nand NAND2 (N22827, N22820, N2957);
nor NOR3 (N22828, N22823, N21487, N13023);
and AND2 (N22829, N22821, N20560);
and AND4 (N22830, N22818, N13605, N14715, N2020);
and AND2 (N22831, N22826, N12738);
xor XOR2 (N22832, N22829, N7806);
nand NAND2 (N22833, N22814, N6985);
nand NAND4 (N22834, N22825, N20408, N19377, N16250);
and AND2 (N22835, N22831, N15771);
buf BUF1 (N22836, N22827);
nor NOR4 (N22837, N22834, N14703, N6954, N12670);
xor XOR2 (N22838, N22824, N13559);
or OR3 (N22839, N22833, N3102, N11106);
xor XOR2 (N22840, N22839, N9586);
nand NAND3 (N22841, N22830, N20030, N11092);
not NOT1 (N22842, N22838);
or OR3 (N22843, N22832, N13902, N13638);
buf BUF1 (N22844, N22797);
or OR4 (N22845, N22843, N4547, N1110, N18429);
not NOT1 (N22846, N22828);
not NOT1 (N22847, N22840);
or OR3 (N22848, N22835, N4530, N13125);
nor NOR3 (N22849, N22845, N2816, N18482);
nor NOR3 (N22850, N22817, N550, N6100);
buf BUF1 (N22851, N22850);
not NOT1 (N22852, N22836);
buf BUF1 (N22853, N22852);
not NOT1 (N22854, N22842);
nor NOR4 (N22855, N22846, N22400, N3080, N1973);
or OR3 (N22856, N22844, N17452, N2460);
not NOT1 (N22857, N22847);
buf BUF1 (N22858, N22856);
not NOT1 (N22859, N22858);
buf BUF1 (N22860, N22857);
xor XOR2 (N22861, N22849, N7108);
nor NOR2 (N22862, N22855, N9844);
and AND2 (N22863, N22854, N21473);
not NOT1 (N22864, N22861);
nor NOR2 (N22865, N22851, N17216);
nor NOR4 (N22866, N22859, N20464, N18835, N7850);
nor NOR4 (N22867, N22866, N4155, N6556, N263);
buf BUF1 (N22868, N22864);
nor NOR2 (N22869, N22848, N7743);
xor XOR2 (N22870, N22865, N2867);
nand NAND4 (N22871, N22870, N4521, N2517, N16967);
nand NAND4 (N22872, N22862, N18719, N2214, N7513);
nand NAND4 (N22873, N22841, N18672, N19429, N122);
not NOT1 (N22874, N22837);
nor NOR4 (N22875, N22874, N18170, N20572, N4776);
xor XOR2 (N22876, N22863, N16366);
nor NOR2 (N22877, N22867, N9798);
xor XOR2 (N22878, N22860, N11246);
buf BUF1 (N22879, N22853);
nor NOR2 (N22880, N22868, N15837);
or OR4 (N22881, N22878, N16505, N14534, N21640);
not NOT1 (N22882, N22880);
nand NAND4 (N22883, N22872, N4233, N22116, N11900);
or OR2 (N22884, N22873, N4568);
nand NAND4 (N22885, N22871, N1594, N13134, N3649);
not NOT1 (N22886, N22875);
xor XOR2 (N22887, N22882, N13261);
nand NAND3 (N22888, N22869, N19842, N15416);
nand NAND3 (N22889, N22879, N12224, N1166);
xor XOR2 (N22890, N22887, N17384);
nor NOR3 (N22891, N22881, N14267, N1446);
nor NOR2 (N22892, N22886, N5764);
not NOT1 (N22893, N22883);
xor XOR2 (N22894, N22884, N16224);
nand NAND2 (N22895, N22885, N14836);
nand NAND3 (N22896, N22892, N5070, N12151);
xor XOR2 (N22897, N22888, N5325);
nor NOR2 (N22898, N22889, N21695);
nand NAND2 (N22899, N22891, N17664);
or OR2 (N22900, N22899, N11484);
nor NOR4 (N22901, N22897, N3330, N16551, N22671);
nand NAND4 (N22902, N22877, N3129, N19101, N19533);
xor XOR2 (N22903, N22898, N11117);
or OR3 (N22904, N22900, N8151, N60);
nor NOR4 (N22905, N22895, N18746, N13169, N10808);
nor NOR3 (N22906, N22890, N10498, N22127);
not NOT1 (N22907, N22903);
nand NAND3 (N22908, N22893, N1229, N7265);
nor NOR3 (N22909, N22902, N17251, N15281);
xor XOR2 (N22910, N22909, N19570);
nor NOR3 (N22911, N22904, N14895, N1762);
buf BUF1 (N22912, N22905);
or OR3 (N22913, N22910, N21615, N15769);
nor NOR4 (N22914, N22876, N666, N16620, N22819);
or OR4 (N22915, N22908, N17126, N6487, N5033);
and AND4 (N22916, N22894, N12988, N4355, N2411);
xor XOR2 (N22917, N22896, N17118);
xor XOR2 (N22918, N22914, N7834);
and AND2 (N22919, N22906, N18770);
and AND3 (N22920, N22915, N19288, N9229);
nand NAND3 (N22921, N22913, N6680, N6976);
nor NOR2 (N22922, N22920, N3714);
or OR3 (N22923, N22917, N20378, N18039);
nand NAND4 (N22924, N22918, N8381, N4099, N16534);
and AND2 (N22925, N22919, N5517);
and AND3 (N22926, N22923, N7845, N12023);
nor NOR2 (N22927, N22911, N6879);
xor XOR2 (N22928, N22927, N16871);
and AND3 (N22929, N22901, N8117, N3954);
and AND4 (N22930, N22925, N15315, N11828, N4247);
xor XOR2 (N22931, N22922, N1491);
xor XOR2 (N22932, N22926, N12898);
or OR4 (N22933, N22912, N2793, N15351, N8792);
nor NOR4 (N22934, N22921, N18354, N15876, N16759);
and AND2 (N22935, N22932, N7445);
xor XOR2 (N22936, N22934, N17810);
or OR2 (N22937, N22928, N21500);
not NOT1 (N22938, N22930);
nand NAND2 (N22939, N22931, N12378);
xor XOR2 (N22940, N22924, N14762);
not NOT1 (N22941, N22937);
buf BUF1 (N22942, N22907);
not NOT1 (N22943, N22929);
xor XOR2 (N22944, N22916, N11621);
and AND4 (N22945, N22933, N8501, N15264, N21208);
or OR3 (N22946, N22942, N12756, N17981);
not NOT1 (N22947, N22940);
nor NOR4 (N22948, N22943, N5685, N15601, N2757);
nand NAND3 (N22949, N22935, N22148, N5081);
buf BUF1 (N22950, N22941);
and AND4 (N22951, N22944, N155, N9203, N22824);
buf BUF1 (N22952, N22945);
nand NAND2 (N22953, N22951, N13187);
buf BUF1 (N22954, N22950);
buf BUF1 (N22955, N22953);
xor XOR2 (N22956, N22954, N6617);
not NOT1 (N22957, N22938);
or OR4 (N22958, N22948, N18913, N7644, N1423);
xor XOR2 (N22959, N22957, N22214);
not NOT1 (N22960, N22936);
buf BUF1 (N22961, N22959);
or OR4 (N22962, N22947, N3945, N17472, N2954);
nand NAND2 (N22963, N22949, N17378);
nand NAND2 (N22964, N22939, N6138);
not NOT1 (N22965, N22960);
xor XOR2 (N22966, N22965, N7910);
buf BUF1 (N22967, N22955);
or OR2 (N22968, N22961, N16822);
buf BUF1 (N22969, N22964);
not NOT1 (N22970, N22967);
and AND3 (N22971, N22968, N14955, N17571);
nor NOR4 (N22972, N22971, N10052, N751, N4729);
and AND4 (N22973, N22956, N2916, N18155, N12566);
and AND2 (N22974, N22952, N6131);
and AND2 (N22975, N22969, N1083);
and AND4 (N22976, N22973, N3032, N22901, N22426);
not NOT1 (N22977, N22976);
or OR2 (N22978, N22946, N18298);
or OR2 (N22979, N22963, N21112);
or OR4 (N22980, N22979, N5852, N7641, N13226);
xor XOR2 (N22981, N22962, N8825);
and AND2 (N22982, N22966, N18788);
or OR3 (N22983, N22975, N18063, N10851);
nor NOR3 (N22984, N22982, N10972, N10939);
buf BUF1 (N22985, N22974);
xor XOR2 (N22986, N22985, N15050);
nand NAND2 (N22987, N22983, N3747);
or OR3 (N22988, N22978, N14345, N14966);
and AND3 (N22989, N22986, N4852, N14305);
or OR4 (N22990, N22988, N6323, N21172, N17206);
and AND3 (N22991, N22981, N13273, N1915);
or OR2 (N22992, N22970, N20163);
not NOT1 (N22993, N22972);
nand NAND2 (N22994, N22977, N5317);
and AND4 (N22995, N22980, N13132, N17827, N21739);
and AND4 (N22996, N22984, N7957, N7865, N6712);
nand NAND4 (N22997, N22996, N17619, N20266, N17250);
not NOT1 (N22998, N22958);
and AND4 (N22999, N22998, N7065, N439, N719);
buf BUF1 (N23000, N22997);
not NOT1 (N23001, N22990);
xor XOR2 (N23002, N22995, N18888);
not NOT1 (N23003, N23002);
nand NAND3 (N23004, N22993, N4402, N21526);
nor NOR3 (N23005, N23003, N15224, N12146);
buf BUF1 (N23006, N22987);
nor NOR4 (N23007, N22992, N5141, N10134, N5891);
nand NAND2 (N23008, N22994, N8860);
or OR2 (N23009, N22989, N17495);
xor XOR2 (N23010, N23000, N6701);
and AND2 (N23011, N23004, N1973);
nand NAND2 (N23012, N22999, N21411);
buf BUF1 (N23013, N23001);
nand NAND3 (N23014, N23010, N8273, N11915);
or OR2 (N23015, N23014, N16471);
nand NAND4 (N23016, N23007, N21239, N2728, N22407);
nand NAND4 (N23017, N23009, N14376, N9926, N19230);
buf BUF1 (N23018, N23017);
xor XOR2 (N23019, N22991, N8451);
or OR3 (N23020, N23011, N16903, N4416);
nor NOR2 (N23021, N23020, N14796);
xor XOR2 (N23022, N23021, N3004);
or OR3 (N23023, N23006, N434, N20281);
nor NOR3 (N23024, N23005, N17130, N20618);
buf BUF1 (N23025, N23022);
xor XOR2 (N23026, N23016, N8110);
nor NOR2 (N23027, N23012, N739);
not NOT1 (N23028, N23024);
buf BUF1 (N23029, N23028);
buf BUF1 (N23030, N23019);
nand NAND4 (N23031, N23026, N13605, N20983, N4840);
buf BUF1 (N23032, N23008);
not NOT1 (N23033, N23030);
or OR4 (N23034, N23033, N4337, N15227, N15785);
xor XOR2 (N23035, N23025, N3560);
nand NAND4 (N23036, N23029, N21282, N17385, N4611);
or OR2 (N23037, N23013, N13482);
nand NAND2 (N23038, N23032, N2148);
nor NOR4 (N23039, N23037, N18146, N22309, N6833);
nor NOR3 (N23040, N23023, N19911, N18689);
and AND2 (N23041, N23035, N14860);
and AND2 (N23042, N23031, N5141);
and AND4 (N23043, N23039, N5783, N686, N13507);
buf BUF1 (N23044, N23040);
and AND3 (N23045, N23018, N19704, N5637);
or OR4 (N23046, N23038, N13029, N15611, N9807);
or OR3 (N23047, N23036, N22106, N13774);
nor NOR4 (N23048, N23043, N8588, N22789, N6202);
nor NOR4 (N23049, N23015, N6987, N7434, N17035);
or OR3 (N23050, N23027, N3710, N15629);
not NOT1 (N23051, N23048);
and AND2 (N23052, N23041, N22618);
not NOT1 (N23053, N23052);
or OR2 (N23054, N23051, N15723);
buf BUF1 (N23055, N23050);
nor NOR3 (N23056, N23053, N6424, N20567);
nand NAND3 (N23057, N23044, N11625, N17587);
or OR2 (N23058, N23054, N7690);
nor NOR2 (N23059, N23055, N16137);
and AND3 (N23060, N23034, N17550, N17461);
nand NAND2 (N23061, N23046, N22642);
nor NOR3 (N23062, N23047, N16542, N16842);
and AND2 (N23063, N23045, N14162);
or OR2 (N23064, N23057, N6528);
and AND4 (N23065, N23062, N3285, N1818, N22622);
nand NAND4 (N23066, N23065, N15560, N4417, N17009);
nor NOR2 (N23067, N23059, N2501);
or OR3 (N23068, N23064, N18248, N8299);
not NOT1 (N23069, N23056);
nand NAND2 (N23070, N23066, N12187);
buf BUF1 (N23071, N23061);
buf BUF1 (N23072, N23060);
nand NAND2 (N23073, N23063, N12738);
xor XOR2 (N23074, N23067, N10321);
not NOT1 (N23075, N23058);
and AND2 (N23076, N23070, N16773);
nand NAND2 (N23077, N23071, N9294);
xor XOR2 (N23078, N23069, N17264);
nand NAND2 (N23079, N23072, N8504);
nand NAND4 (N23080, N23075, N2566, N17471, N22068);
buf BUF1 (N23081, N23068);
buf BUF1 (N23082, N23049);
not NOT1 (N23083, N23079);
buf BUF1 (N23084, N23081);
and AND4 (N23085, N23078, N4418, N18914, N7976);
or OR3 (N23086, N23073, N19356, N11810);
buf BUF1 (N23087, N23084);
nand NAND2 (N23088, N23077, N19294);
not NOT1 (N23089, N23082);
not NOT1 (N23090, N23086);
or OR4 (N23091, N23080, N12692, N14731, N8574);
or OR3 (N23092, N23085, N5690, N5015);
nand NAND3 (N23093, N23042, N15467, N11391);
nor NOR4 (N23094, N23076, N13462, N19789, N10604);
and AND2 (N23095, N23089, N8351);
nor NOR2 (N23096, N23074, N22591);
nor NOR4 (N23097, N23095, N15037, N10263, N19597);
not NOT1 (N23098, N23088);
nor NOR2 (N23099, N23094, N9770);
or OR2 (N23100, N23087, N6373);
xor XOR2 (N23101, N23093, N10139);
xor XOR2 (N23102, N23091, N19084);
buf BUF1 (N23103, N23102);
and AND2 (N23104, N23097, N5117);
nor NOR3 (N23105, N23083, N15781, N12237);
buf BUF1 (N23106, N23104);
nand NAND4 (N23107, N23103, N3509, N10750, N3754);
not NOT1 (N23108, N23092);
and AND3 (N23109, N23101, N5563, N17986);
xor XOR2 (N23110, N23108, N10409);
and AND4 (N23111, N23090, N10434, N19615, N13789);
xor XOR2 (N23112, N23109, N9285);
and AND4 (N23113, N23111, N13713, N5652, N413);
buf BUF1 (N23114, N23106);
and AND2 (N23115, N23105, N14058);
nor NOR3 (N23116, N23113, N22792, N6552);
xor XOR2 (N23117, N23100, N11415);
and AND2 (N23118, N23110, N20847);
buf BUF1 (N23119, N23098);
nor NOR4 (N23120, N23118, N23071, N12679, N18096);
xor XOR2 (N23121, N23112, N11350);
nand NAND2 (N23122, N23119, N3456);
not NOT1 (N23123, N23122);
nand NAND2 (N23124, N23107, N21437);
nand NAND2 (N23125, N23115, N4981);
and AND4 (N23126, N23116, N10769, N5788, N7246);
nor NOR2 (N23127, N23096, N19017);
nor NOR3 (N23128, N23124, N4298, N19565);
nor NOR4 (N23129, N23099, N614, N13204, N12863);
buf BUF1 (N23130, N23128);
or OR3 (N23131, N23121, N16914, N16116);
xor XOR2 (N23132, N23123, N9376);
nand NAND3 (N23133, N23129, N15739, N16313);
xor XOR2 (N23134, N23125, N18937);
buf BUF1 (N23135, N23120);
buf BUF1 (N23136, N23126);
or OR3 (N23137, N23135, N579, N12856);
nor NOR4 (N23138, N23132, N17395, N10881, N488);
buf BUF1 (N23139, N23131);
xor XOR2 (N23140, N23133, N9060);
xor XOR2 (N23141, N23130, N16316);
and AND3 (N23142, N23114, N18685, N1963);
and AND3 (N23143, N23140, N5502, N21109);
buf BUF1 (N23144, N23117);
not NOT1 (N23145, N23144);
not NOT1 (N23146, N23142);
nor NOR3 (N23147, N23137, N18323, N15979);
not NOT1 (N23148, N23127);
nand NAND2 (N23149, N23141, N8399);
not NOT1 (N23150, N23148);
not NOT1 (N23151, N23143);
nand NAND4 (N23152, N23136, N8740, N20015, N18510);
not NOT1 (N23153, N23145);
and AND3 (N23154, N23134, N16862, N21872);
nor NOR3 (N23155, N23153, N16871, N22858);
not NOT1 (N23156, N23147);
and AND3 (N23157, N23151, N8199, N3033);
and AND2 (N23158, N23139, N3909);
and AND4 (N23159, N23157, N16491, N18701, N13206);
nor NOR4 (N23160, N23146, N7400, N8526, N20617);
not NOT1 (N23161, N23154);
nor NOR2 (N23162, N23152, N7791);
not NOT1 (N23163, N23149);
or OR4 (N23164, N23160, N22259, N9296, N16795);
or OR4 (N23165, N23150, N1515, N18834, N9139);
xor XOR2 (N23166, N23162, N130);
xor XOR2 (N23167, N23159, N6873);
xor XOR2 (N23168, N23164, N12471);
and AND4 (N23169, N23165, N9514, N7001, N3599);
nor NOR3 (N23170, N23166, N21989, N3193);
or OR2 (N23171, N23168, N10353);
xor XOR2 (N23172, N23171, N19469);
buf BUF1 (N23173, N23156);
and AND3 (N23174, N23172, N14076, N22605);
not NOT1 (N23175, N23174);
xor XOR2 (N23176, N23170, N11915);
and AND3 (N23177, N23163, N13764, N19132);
buf BUF1 (N23178, N23177);
or OR4 (N23179, N23138, N15308, N11919, N8073);
and AND4 (N23180, N23167, N16513, N13252, N15886);
xor XOR2 (N23181, N23180, N11459);
xor XOR2 (N23182, N23181, N22921);
xor XOR2 (N23183, N23173, N15542);
nand NAND4 (N23184, N23176, N7428, N14326, N21951);
and AND2 (N23185, N23179, N14899);
nor NOR3 (N23186, N23175, N4972, N2034);
and AND3 (N23187, N23183, N11275, N17170);
nor NOR4 (N23188, N23185, N23170, N15971, N3337);
nor NOR3 (N23189, N23158, N10576, N9526);
buf BUF1 (N23190, N23178);
not NOT1 (N23191, N23188);
nor NOR2 (N23192, N23182, N20805);
buf BUF1 (N23193, N23186);
buf BUF1 (N23194, N23193);
not NOT1 (N23195, N23184);
and AND4 (N23196, N23161, N21990, N7704, N22619);
buf BUF1 (N23197, N23191);
not NOT1 (N23198, N23192);
nor NOR2 (N23199, N23189, N22758);
or OR4 (N23200, N23155, N6404, N3226, N7482);
nor NOR3 (N23201, N23195, N17927, N22764);
buf BUF1 (N23202, N23200);
or OR2 (N23203, N23199, N3186);
not NOT1 (N23204, N23202);
nand NAND2 (N23205, N23190, N20340);
nor NOR3 (N23206, N23204, N21898, N21046);
nor NOR2 (N23207, N23203, N705);
nand NAND3 (N23208, N23201, N22153, N2088);
and AND4 (N23209, N23187, N18778, N8915, N8623);
nand NAND4 (N23210, N23207, N3060, N18767, N4780);
and AND3 (N23211, N23196, N4443, N7392);
nand NAND3 (N23212, N23206, N13247, N20942);
nand NAND3 (N23213, N23197, N17319, N14624);
not NOT1 (N23214, N23213);
and AND2 (N23215, N23214, N22317);
not NOT1 (N23216, N23211);
and AND2 (N23217, N23209, N10413);
nor NOR3 (N23218, N23205, N13935, N3164);
buf BUF1 (N23219, N23218);
or OR4 (N23220, N23212, N8887, N20835, N8314);
or OR2 (N23221, N23194, N17476);
nor NOR4 (N23222, N23220, N3590, N18707, N16297);
or OR2 (N23223, N23208, N11797);
not NOT1 (N23224, N23223);
and AND2 (N23225, N23169, N10980);
buf BUF1 (N23226, N23219);
not NOT1 (N23227, N23221);
or OR3 (N23228, N23198, N12529, N10241);
nand NAND4 (N23229, N23225, N6544, N13430, N19397);
not NOT1 (N23230, N23224);
or OR2 (N23231, N23228, N7729);
buf BUF1 (N23232, N23222);
and AND3 (N23233, N23229, N16160, N2286);
nand NAND4 (N23234, N23217, N15481, N746, N18012);
nand NAND4 (N23235, N23231, N5769, N10686, N11507);
not NOT1 (N23236, N23210);
or OR4 (N23237, N23227, N45, N47, N5163);
nor NOR3 (N23238, N23235, N23119, N8887);
or OR3 (N23239, N23234, N4270, N306);
and AND3 (N23240, N23236, N3394, N13882);
or OR4 (N23241, N23226, N12304, N6500, N13197);
and AND3 (N23242, N23240, N12128, N9542);
nor NOR4 (N23243, N23238, N11193, N12522, N7770);
buf BUF1 (N23244, N23237);
nand NAND2 (N23245, N23216, N6059);
nand NAND2 (N23246, N23245, N18459);
and AND4 (N23247, N23215, N19716, N12342, N3478);
buf BUF1 (N23248, N23246);
buf BUF1 (N23249, N23244);
or OR3 (N23250, N23230, N14041, N451);
and AND3 (N23251, N23239, N4060, N7765);
nand NAND4 (N23252, N23243, N1453, N13541, N18967);
buf BUF1 (N23253, N23247);
xor XOR2 (N23254, N23250, N21109);
buf BUF1 (N23255, N23254);
and AND4 (N23256, N23233, N21170, N18309, N5816);
not NOT1 (N23257, N23249);
nand NAND4 (N23258, N23232, N3154, N5198, N9211);
xor XOR2 (N23259, N23248, N1227);
not NOT1 (N23260, N23255);
not NOT1 (N23261, N23251);
nor NOR3 (N23262, N23257, N5995, N17939);
nor NOR2 (N23263, N23256, N209);
and AND3 (N23264, N23258, N6773, N20334);
not NOT1 (N23265, N23253);
and AND2 (N23266, N23265, N7314);
and AND2 (N23267, N23260, N4076);
and AND4 (N23268, N23267, N22349, N2694, N19557);
nor NOR4 (N23269, N23261, N15420, N21312, N12645);
and AND2 (N23270, N23268, N19375);
xor XOR2 (N23271, N23252, N9063);
and AND2 (N23272, N23241, N16742);
nor NOR4 (N23273, N23242, N10428, N10757, N7580);
buf BUF1 (N23274, N23272);
xor XOR2 (N23275, N23269, N1521);
buf BUF1 (N23276, N23262);
nand NAND2 (N23277, N23273, N20370);
xor XOR2 (N23278, N23271, N21405);
buf BUF1 (N23279, N23278);
nor NOR2 (N23280, N23277, N16121);
nand NAND4 (N23281, N23276, N18970, N7915, N8459);
buf BUF1 (N23282, N23266);
not NOT1 (N23283, N23280);
nand NAND3 (N23284, N23279, N19004, N12206);
nand NAND3 (N23285, N23264, N18732, N16310);
not NOT1 (N23286, N23274);
xor XOR2 (N23287, N23263, N13503);
nor NOR3 (N23288, N23275, N12721, N9475);
nand NAND3 (N23289, N23286, N7409, N7529);
or OR3 (N23290, N23282, N10232, N6072);
xor XOR2 (N23291, N23289, N5949);
nor NOR2 (N23292, N23270, N14797);
and AND4 (N23293, N23287, N11142, N2136, N7912);
buf BUF1 (N23294, N23290);
or OR3 (N23295, N23283, N19589, N16739);
nand NAND2 (N23296, N23294, N16055);
nand NAND4 (N23297, N23292, N11832, N19605, N14445);
not NOT1 (N23298, N23288);
not NOT1 (N23299, N23298);
xor XOR2 (N23300, N23259, N3048);
xor XOR2 (N23301, N23285, N6243);
nor NOR3 (N23302, N23293, N12107, N51);
nor NOR3 (N23303, N23284, N13488, N11438);
or OR2 (N23304, N23303, N1429);
nand NAND2 (N23305, N23296, N15425);
buf BUF1 (N23306, N23301);
or OR4 (N23307, N23297, N12763, N13443, N21885);
not NOT1 (N23308, N23306);
nand NAND2 (N23309, N23291, N17644);
nor NOR2 (N23310, N23309, N3122);
nand NAND4 (N23311, N23304, N17020, N12809, N1216);
nand NAND3 (N23312, N23310, N645, N16986);
and AND3 (N23313, N23281, N1961, N5845);
not NOT1 (N23314, N23308);
xor XOR2 (N23315, N23300, N17889);
xor XOR2 (N23316, N23313, N15299);
or OR2 (N23317, N23315, N14923);
nand NAND4 (N23318, N23299, N17548, N8063, N13340);
buf BUF1 (N23319, N23312);
nand NAND2 (N23320, N23307, N10152);
nand NAND4 (N23321, N23316, N6060, N4226, N1680);
nand NAND4 (N23322, N23317, N21280, N6769, N358);
nand NAND3 (N23323, N23322, N9363, N3387);
buf BUF1 (N23324, N23323);
not NOT1 (N23325, N23318);
buf BUF1 (N23326, N23320);
nor NOR3 (N23327, N23325, N8262, N19631);
xor XOR2 (N23328, N23295, N19305);
or OR4 (N23329, N23326, N21184, N13554, N4007);
not NOT1 (N23330, N23328);
not NOT1 (N23331, N23330);
nand NAND3 (N23332, N23327, N20533, N10200);
xor XOR2 (N23333, N23319, N17857);
buf BUF1 (N23334, N23305);
nor NOR2 (N23335, N23302, N4776);
and AND2 (N23336, N23333, N16722);
xor XOR2 (N23337, N23329, N17980);
or OR4 (N23338, N23321, N8626, N11046, N19669);
or OR3 (N23339, N23314, N18888, N10501);
nor NOR4 (N23340, N23337, N10256, N18222, N22123);
nand NAND2 (N23341, N23335, N2886);
or OR2 (N23342, N23334, N20159);
xor XOR2 (N23343, N23342, N13805);
or OR2 (N23344, N23338, N7720);
buf BUF1 (N23345, N23332);
buf BUF1 (N23346, N23339);
nor NOR2 (N23347, N23343, N16797);
nand NAND4 (N23348, N23347, N18081, N16405, N4932);
nor NOR3 (N23349, N23346, N21244, N18908);
nor NOR2 (N23350, N23331, N22097);
not NOT1 (N23351, N23336);
not NOT1 (N23352, N23349);
xor XOR2 (N23353, N23348, N4921);
not NOT1 (N23354, N23340);
xor XOR2 (N23355, N23341, N11343);
or OR2 (N23356, N23354, N14178);
xor XOR2 (N23357, N23352, N4313);
nor NOR2 (N23358, N23324, N20789);
nor NOR3 (N23359, N23356, N5090, N8827);
nor NOR4 (N23360, N23357, N12519, N13922, N16747);
nor NOR4 (N23361, N23311, N2435, N20406, N945);
nor NOR4 (N23362, N23360, N15162, N9414, N364);
nand NAND4 (N23363, N23350, N18322, N2239, N10065);
not NOT1 (N23364, N23353);
xor XOR2 (N23365, N23361, N16830);
or OR4 (N23366, N23358, N9449, N1307, N14204);
and AND4 (N23367, N23355, N5628, N15549, N2085);
buf BUF1 (N23368, N23365);
nor NOR2 (N23369, N23368, N18653);
not NOT1 (N23370, N23362);
nor NOR3 (N23371, N23359, N1115, N20067);
buf BUF1 (N23372, N23344);
buf BUF1 (N23373, N23369);
or OR3 (N23374, N23366, N19457, N21467);
nand NAND3 (N23375, N23373, N4563, N15424);
nand NAND2 (N23376, N23364, N21310);
nand NAND2 (N23377, N23372, N3606);
nor NOR3 (N23378, N23367, N5716, N1988);
nor NOR4 (N23379, N23363, N17908, N11666, N5228);
not NOT1 (N23380, N23371);
buf BUF1 (N23381, N23375);
nand NAND2 (N23382, N23370, N16588);
nand NAND4 (N23383, N23345, N13148, N10638, N5778);
not NOT1 (N23384, N23383);
or OR4 (N23385, N23384, N4594, N13837, N13691);
nand NAND2 (N23386, N23378, N12023);
not NOT1 (N23387, N23377);
not NOT1 (N23388, N23382);
buf BUF1 (N23389, N23379);
and AND4 (N23390, N23381, N13173, N4674, N3830);
nor NOR4 (N23391, N23389, N21652, N6736, N17299);
nand NAND3 (N23392, N23380, N14839, N3316);
nor NOR4 (N23393, N23385, N11782, N23363, N17744);
nand NAND4 (N23394, N23393, N21671, N16131, N17017);
xor XOR2 (N23395, N23376, N20238);
or OR2 (N23396, N23374, N15702);
or OR3 (N23397, N23394, N23295, N2201);
xor XOR2 (N23398, N23387, N21307);
buf BUF1 (N23399, N23388);
buf BUF1 (N23400, N23386);
and AND2 (N23401, N23351, N17894);
nor NOR3 (N23402, N23390, N12073, N14164);
nand NAND2 (N23403, N23401, N19503);
or OR4 (N23404, N23396, N19299, N9884, N1961);
nor NOR2 (N23405, N23391, N18584);
nor NOR2 (N23406, N23402, N13587);
and AND3 (N23407, N23395, N16689, N5584);
nand NAND3 (N23408, N23407, N17708, N14627);
not NOT1 (N23409, N23397);
xor XOR2 (N23410, N23408, N10190);
nand NAND4 (N23411, N23409, N17050, N3450, N13966);
nand NAND2 (N23412, N23399, N15169);
nand NAND2 (N23413, N23410, N2297);
xor XOR2 (N23414, N23411, N13740);
not NOT1 (N23415, N23403);
and AND2 (N23416, N23405, N7743);
or OR3 (N23417, N23414, N7251, N22709);
buf BUF1 (N23418, N23404);
xor XOR2 (N23419, N23406, N7551);
and AND2 (N23420, N23419, N18633);
and AND3 (N23421, N23400, N2742, N13975);
xor XOR2 (N23422, N23417, N9905);
nand NAND2 (N23423, N23420, N2933);
nor NOR3 (N23424, N23418, N17854, N4479);
not NOT1 (N23425, N23424);
and AND2 (N23426, N23421, N9662);
nand NAND4 (N23427, N23413, N16398, N9001, N10566);
and AND3 (N23428, N23425, N11415, N8403);
nor NOR4 (N23429, N23392, N21849, N15725, N17586);
not NOT1 (N23430, N23398);
or OR3 (N23431, N23415, N8140, N13720);
and AND4 (N23432, N23422, N17378, N21122, N10713);
and AND4 (N23433, N23426, N18714, N166, N11950);
or OR4 (N23434, N23429, N849, N11576, N5819);
and AND4 (N23435, N23412, N4419, N18593, N6911);
not NOT1 (N23436, N23432);
buf BUF1 (N23437, N23435);
nor NOR2 (N23438, N23434, N10895);
not NOT1 (N23439, N23438);
buf BUF1 (N23440, N23431);
xor XOR2 (N23441, N23439, N5951);
or OR2 (N23442, N23436, N8123);
nor NOR3 (N23443, N23437, N10900, N9188);
buf BUF1 (N23444, N23433);
and AND2 (N23445, N23444, N21860);
and AND3 (N23446, N23442, N3985, N13808);
buf BUF1 (N23447, N23441);
not NOT1 (N23448, N23443);
xor XOR2 (N23449, N23440, N17709);
nand NAND2 (N23450, N23448, N9602);
buf BUF1 (N23451, N23446);
xor XOR2 (N23452, N23447, N2561);
nor NOR4 (N23453, N23450, N21089, N5448, N17642);
xor XOR2 (N23454, N23445, N787);
buf BUF1 (N23455, N23428);
buf BUF1 (N23456, N23449);
or OR3 (N23457, N23427, N10189, N21914);
or OR2 (N23458, N23454, N8752);
not NOT1 (N23459, N23430);
and AND2 (N23460, N23452, N17736);
nor NOR3 (N23461, N23457, N17193, N1235);
nand NAND4 (N23462, N23453, N10367, N531, N14373);
and AND2 (N23463, N23458, N20303);
nor NOR3 (N23464, N23462, N15798, N7053);
or OR2 (N23465, N23464, N7423);
xor XOR2 (N23466, N23459, N8974);
nand NAND2 (N23467, N23463, N20915);
or OR2 (N23468, N23466, N18161);
not NOT1 (N23469, N23460);
and AND3 (N23470, N23423, N20370, N12098);
nor NOR3 (N23471, N23451, N22772, N18425);
not NOT1 (N23472, N23467);
buf BUF1 (N23473, N23471);
buf BUF1 (N23474, N23416);
nor NOR2 (N23475, N23455, N15686);
or OR2 (N23476, N23470, N6464);
xor XOR2 (N23477, N23476, N12253);
not NOT1 (N23478, N23475);
buf BUF1 (N23479, N23472);
and AND4 (N23480, N23461, N18983, N6504, N17109);
buf BUF1 (N23481, N23473);
xor XOR2 (N23482, N23479, N20293);
not NOT1 (N23483, N23481);
nor NOR2 (N23484, N23477, N22085);
and AND4 (N23485, N23484, N14225, N14875, N9772);
not NOT1 (N23486, N23465);
buf BUF1 (N23487, N23456);
xor XOR2 (N23488, N23468, N14569);
xor XOR2 (N23489, N23486, N21737);
buf BUF1 (N23490, N23478);
or OR2 (N23491, N23485, N19995);
buf BUF1 (N23492, N23469);
nand NAND4 (N23493, N23490, N10080, N3889, N12119);
xor XOR2 (N23494, N23482, N19913);
buf BUF1 (N23495, N23494);
buf BUF1 (N23496, N23491);
xor XOR2 (N23497, N23492, N3157);
not NOT1 (N23498, N23480);
and AND4 (N23499, N23474, N19903, N15146, N1169);
nand NAND3 (N23500, N23483, N19013, N2159);
buf BUF1 (N23501, N23499);
or OR3 (N23502, N23501, N986, N21232);
xor XOR2 (N23503, N23493, N2520);
and AND2 (N23504, N23495, N21692);
buf BUF1 (N23505, N23497);
and AND4 (N23506, N23500, N13981, N12246, N13975);
nor NOR3 (N23507, N23506, N21993, N11556);
or OR2 (N23508, N23503, N22644);
buf BUF1 (N23509, N23489);
and AND3 (N23510, N23508, N7709, N2897);
not NOT1 (N23511, N23498);
buf BUF1 (N23512, N23496);
xor XOR2 (N23513, N23511, N16737);
or OR3 (N23514, N23504, N15905, N20617);
xor XOR2 (N23515, N23512, N8605);
buf BUF1 (N23516, N23507);
and AND2 (N23517, N23515, N11937);
buf BUF1 (N23518, N23516);
xor XOR2 (N23519, N23517, N23431);
nand NAND4 (N23520, N23518, N19753, N21489, N2110);
nor NOR4 (N23521, N23519, N3626, N13321, N23148);
nand NAND3 (N23522, N23505, N9951, N21083);
xor XOR2 (N23523, N23520, N14948);
nor NOR2 (N23524, N23510, N6088);
nor NOR2 (N23525, N23523, N16197);
and AND2 (N23526, N23488, N10877);
or OR4 (N23527, N23522, N7467, N15377, N13320);
xor XOR2 (N23528, N23521, N11504);
nand NAND2 (N23529, N23525, N15142);
buf BUF1 (N23530, N23509);
buf BUF1 (N23531, N23530);
or OR3 (N23532, N23528, N1258, N8829);
buf BUF1 (N23533, N23513);
or OR2 (N23534, N23531, N10763);
nand NAND3 (N23535, N23514, N15750, N22588);
and AND4 (N23536, N23502, N7731, N14363, N5248);
and AND2 (N23537, N23534, N19612);
not NOT1 (N23538, N23527);
and AND2 (N23539, N23536, N22474);
nor NOR4 (N23540, N23487, N3559, N12558, N3976);
buf BUF1 (N23541, N23532);
not NOT1 (N23542, N23529);
buf BUF1 (N23543, N23537);
nor NOR4 (N23544, N23533, N4439, N13074, N6729);
nor NOR3 (N23545, N23543, N1611, N11824);
buf BUF1 (N23546, N23539);
xor XOR2 (N23547, N23538, N18699);
or OR2 (N23548, N23547, N22134);
xor XOR2 (N23549, N23535, N17097);
and AND2 (N23550, N23524, N740);
or OR2 (N23551, N23545, N4779);
xor XOR2 (N23552, N23551, N20121);
not NOT1 (N23553, N23546);
or OR3 (N23554, N23526, N13090, N13195);
xor XOR2 (N23555, N23552, N20629);
xor XOR2 (N23556, N23555, N14272);
buf BUF1 (N23557, N23542);
not NOT1 (N23558, N23556);
and AND3 (N23559, N23557, N7869, N15984);
and AND4 (N23560, N23558, N5926, N8882, N2614);
or OR3 (N23561, N23553, N2342, N2196);
nand NAND2 (N23562, N23549, N1553);
and AND2 (N23563, N23540, N14236);
xor XOR2 (N23564, N23550, N22029);
nand NAND3 (N23565, N23554, N1909, N13274);
nor NOR4 (N23566, N23548, N2096, N13686, N16940);
nand NAND4 (N23567, N23562, N18190, N9540, N9364);
or OR3 (N23568, N23560, N15433, N8714);
xor XOR2 (N23569, N23566, N22305);
not NOT1 (N23570, N23541);
and AND3 (N23571, N23567, N9991, N15614);
not NOT1 (N23572, N23564);
or OR2 (N23573, N23572, N1051);
not NOT1 (N23574, N23561);
xor XOR2 (N23575, N23559, N22064);
xor XOR2 (N23576, N23569, N17858);
nor NOR3 (N23577, N23574, N6442, N7657);
buf BUF1 (N23578, N23571);
buf BUF1 (N23579, N23544);
buf BUF1 (N23580, N23568);
nor NOR2 (N23581, N23563, N10923);
not NOT1 (N23582, N23577);
not NOT1 (N23583, N23580);
xor XOR2 (N23584, N23570, N11342);
nor NOR4 (N23585, N23579, N2028, N21263, N11146);
and AND2 (N23586, N23583, N19321);
and AND4 (N23587, N23573, N22756, N4150, N10766);
not NOT1 (N23588, N23584);
nor NOR4 (N23589, N23585, N16344, N13579, N4199);
xor XOR2 (N23590, N23582, N5420);
xor XOR2 (N23591, N23581, N1012);
xor XOR2 (N23592, N23588, N14257);
or OR2 (N23593, N23592, N11761);
buf BUF1 (N23594, N23590);
buf BUF1 (N23595, N23586);
xor XOR2 (N23596, N23576, N12373);
nand NAND2 (N23597, N23578, N592);
nor NOR3 (N23598, N23587, N5514, N2363);
or OR2 (N23599, N23575, N1930);
buf BUF1 (N23600, N23589);
nand NAND4 (N23601, N23600, N5762, N11501, N9327);
buf BUF1 (N23602, N23594);
xor XOR2 (N23603, N23595, N15008);
or OR2 (N23604, N23593, N21369);
nand NAND3 (N23605, N23565, N19056, N8904);
and AND3 (N23606, N23601, N11419, N14231);
xor XOR2 (N23607, N23596, N15370);
nand NAND4 (N23608, N23606, N8916, N20528, N22578);
buf BUF1 (N23609, N23608);
buf BUF1 (N23610, N23591);
xor XOR2 (N23611, N23605, N11534);
not NOT1 (N23612, N23599);
and AND3 (N23613, N23607, N7498, N3834);
nand NAND2 (N23614, N23598, N16784);
xor XOR2 (N23615, N23609, N8593);
buf BUF1 (N23616, N23613);
or OR3 (N23617, N23602, N9117, N4283);
and AND2 (N23618, N23610, N19402);
nand NAND3 (N23619, N23614, N18972, N22963);
nand NAND3 (N23620, N23604, N10045, N10368);
nor NOR2 (N23621, N23619, N16907);
not NOT1 (N23622, N23616);
or OR3 (N23623, N23621, N12867, N10861);
nand NAND4 (N23624, N23603, N19502, N2946, N15338);
nor NOR3 (N23625, N23611, N18597, N19474);
nand NAND3 (N23626, N23623, N23026, N6286);
or OR3 (N23627, N23618, N14234, N11384);
nand NAND3 (N23628, N23597, N14157, N18639);
not NOT1 (N23629, N23626);
nor NOR3 (N23630, N23629, N15691, N10027);
xor XOR2 (N23631, N23627, N6018);
not NOT1 (N23632, N23624);
xor XOR2 (N23633, N23612, N529);
and AND4 (N23634, N23628, N5989, N17184, N7859);
xor XOR2 (N23635, N23620, N18945);
nor NOR2 (N23636, N23625, N19483);
xor XOR2 (N23637, N23632, N18837);
nor NOR2 (N23638, N23637, N3757);
and AND2 (N23639, N23635, N6189);
xor XOR2 (N23640, N23633, N16747);
buf BUF1 (N23641, N23630);
buf BUF1 (N23642, N23615);
buf BUF1 (N23643, N23631);
xor XOR2 (N23644, N23643, N13621);
nand NAND2 (N23645, N23638, N16400);
and AND2 (N23646, N23641, N16241);
nand NAND3 (N23647, N23642, N9118, N23403);
nor NOR3 (N23648, N23639, N2953, N21858);
not NOT1 (N23649, N23647);
nor NOR3 (N23650, N23649, N10886, N3593);
or OR3 (N23651, N23640, N20027, N7058);
not NOT1 (N23652, N23646);
buf BUF1 (N23653, N23634);
buf BUF1 (N23654, N23636);
not NOT1 (N23655, N23650);
buf BUF1 (N23656, N23654);
nor NOR2 (N23657, N23655, N19210);
xor XOR2 (N23658, N23651, N11949);
buf BUF1 (N23659, N23657);
nor NOR3 (N23660, N23653, N20512, N20724);
buf BUF1 (N23661, N23617);
or OR2 (N23662, N23661, N18789);
nor NOR3 (N23663, N23662, N8232, N1126);
buf BUF1 (N23664, N23622);
or OR3 (N23665, N23658, N20447, N5392);
not NOT1 (N23666, N23656);
nor NOR3 (N23667, N23652, N16248, N1700);
or OR3 (N23668, N23660, N18724, N5321);
not NOT1 (N23669, N23666);
and AND3 (N23670, N23645, N5059, N16556);
or OR3 (N23671, N23667, N1565, N11736);
buf BUF1 (N23672, N23644);
nor NOR2 (N23673, N23663, N12349);
buf BUF1 (N23674, N23648);
nand NAND3 (N23675, N23674, N16945, N13813);
or OR4 (N23676, N23671, N11284, N3347, N8261);
nand NAND4 (N23677, N23675, N10829, N3330, N3161);
and AND4 (N23678, N23673, N19075, N15933, N22823);
nand NAND4 (N23679, N23677, N7399, N8259, N9866);
nand NAND4 (N23680, N23676, N9499, N648, N14580);
or OR2 (N23681, N23678, N13066);
xor XOR2 (N23682, N23664, N16266);
nor NOR2 (N23683, N23670, N20174);
xor XOR2 (N23684, N23680, N4413);
nand NAND4 (N23685, N23668, N13469, N16261, N3543);
nand NAND3 (N23686, N23682, N17502, N8041);
not NOT1 (N23687, N23659);
or OR2 (N23688, N23681, N22822);
xor XOR2 (N23689, N23679, N1361);
or OR2 (N23690, N23685, N14380);
or OR2 (N23691, N23687, N3582);
buf BUF1 (N23692, N23665);
nor NOR3 (N23693, N23669, N2150, N11344);
or OR3 (N23694, N23692, N17892, N23071);
and AND4 (N23695, N23690, N12454, N14494, N21751);
nand NAND2 (N23696, N23688, N7714);
and AND3 (N23697, N23691, N5982, N10010);
nand NAND3 (N23698, N23697, N9897, N8149);
not NOT1 (N23699, N23693);
buf BUF1 (N23700, N23689);
or OR3 (N23701, N23700, N2072, N15945);
and AND3 (N23702, N23684, N17918, N4530);
xor XOR2 (N23703, N23701, N20949);
nand NAND3 (N23704, N23703, N19245, N3747);
nor NOR3 (N23705, N23683, N9816, N21935);
and AND2 (N23706, N23704, N10011);
and AND2 (N23707, N23698, N9861);
not NOT1 (N23708, N23695);
nor NOR2 (N23709, N23686, N21646);
buf BUF1 (N23710, N23699);
and AND3 (N23711, N23702, N17458, N4070);
or OR2 (N23712, N23705, N18166);
and AND3 (N23713, N23707, N1755, N4936);
not NOT1 (N23714, N23696);
and AND4 (N23715, N23706, N7312, N2408, N9803);
and AND2 (N23716, N23715, N2509);
xor XOR2 (N23717, N23716, N13121);
not NOT1 (N23718, N23711);
not NOT1 (N23719, N23717);
not NOT1 (N23720, N23709);
xor XOR2 (N23721, N23672, N6443);
not NOT1 (N23722, N23719);
nand NAND3 (N23723, N23721, N9889, N6375);
not NOT1 (N23724, N23718);
or OR4 (N23725, N23723, N19502, N13984, N7336);
xor XOR2 (N23726, N23708, N10017);
nor NOR3 (N23727, N23720, N22988, N22311);
nor NOR4 (N23728, N23694, N6598, N1943, N15286);
xor XOR2 (N23729, N23726, N15788);
or OR4 (N23730, N23725, N10812, N12002, N13953);
nor NOR4 (N23731, N23712, N207, N21194, N21449);
nor NOR4 (N23732, N23728, N14234, N11185, N3392);
buf BUF1 (N23733, N23713);
buf BUF1 (N23734, N23714);
not NOT1 (N23735, N23731);
not NOT1 (N23736, N23710);
buf BUF1 (N23737, N23736);
xor XOR2 (N23738, N23732, N2669);
nand NAND4 (N23739, N23738, N14740, N14035, N23169);
nor NOR3 (N23740, N23737, N3383, N19506);
xor XOR2 (N23741, N23730, N8445);
not NOT1 (N23742, N23729);
nand NAND2 (N23743, N23724, N19556);
xor XOR2 (N23744, N23739, N755);
nor NOR3 (N23745, N23735, N21544, N21164);
and AND3 (N23746, N23722, N10499, N6480);
nand NAND3 (N23747, N23745, N12244, N2098);
nand NAND2 (N23748, N23740, N19556);
nand NAND2 (N23749, N23734, N4209);
and AND3 (N23750, N23741, N17535, N18620);
not NOT1 (N23751, N23742);
or OR4 (N23752, N23727, N13367, N19260, N1108);
and AND3 (N23753, N23748, N4154, N12969);
or OR4 (N23754, N23746, N19375, N20174, N13908);
nor NOR3 (N23755, N23747, N11684, N18409);
nor NOR3 (N23756, N23750, N8565, N16753);
nor NOR3 (N23757, N23756, N15330, N17596);
buf BUF1 (N23758, N23755);
not NOT1 (N23759, N23754);
buf BUF1 (N23760, N23733);
and AND3 (N23761, N23751, N13177, N18811);
buf BUF1 (N23762, N23760);
buf BUF1 (N23763, N23758);
or OR2 (N23764, N23753, N15670);
nor NOR2 (N23765, N23752, N13798);
xor XOR2 (N23766, N23761, N5529);
or OR4 (N23767, N23749, N1075, N23262, N14334);
or OR4 (N23768, N23765, N23333, N3769, N16967);
nand NAND4 (N23769, N23757, N5386, N226, N3869);
xor XOR2 (N23770, N23743, N19321);
buf BUF1 (N23771, N23764);
nand NAND3 (N23772, N23770, N15612, N592);
nand NAND2 (N23773, N23766, N8428);
not NOT1 (N23774, N23763);
buf BUF1 (N23775, N23774);
nand NAND3 (N23776, N23744, N22722, N14162);
not NOT1 (N23777, N23769);
nor NOR4 (N23778, N23762, N19825, N1364, N5808);
not NOT1 (N23779, N23772);
buf BUF1 (N23780, N23767);
nor NOR4 (N23781, N23771, N10361, N11543, N6179);
nand NAND3 (N23782, N23780, N17831, N3951);
nor NOR3 (N23783, N23768, N2885, N18947);
xor XOR2 (N23784, N23781, N8955);
xor XOR2 (N23785, N23782, N22619);
xor XOR2 (N23786, N23777, N15665);
not NOT1 (N23787, N23759);
and AND3 (N23788, N23779, N19178, N20391);
not NOT1 (N23789, N23775);
or OR3 (N23790, N23788, N23516, N13295);
nor NOR2 (N23791, N23790, N1982);
xor XOR2 (N23792, N23785, N9597);
or OR2 (N23793, N23792, N15476);
nor NOR2 (N23794, N23791, N6294);
nand NAND4 (N23795, N23786, N10543, N9562, N5772);
xor XOR2 (N23796, N23784, N9690);
nand NAND3 (N23797, N23776, N7841, N13082);
or OR4 (N23798, N23797, N19247, N18680, N2415);
nand NAND2 (N23799, N23794, N23097);
xor XOR2 (N23800, N23778, N17569);
nor NOR3 (N23801, N23798, N10611, N10995);
buf BUF1 (N23802, N23789);
xor XOR2 (N23803, N23793, N17268);
and AND2 (N23804, N23796, N11397);
nor NOR3 (N23805, N23799, N2950, N2237);
not NOT1 (N23806, N23773);
xor XOR2 (N23807, N23802, N13811);
or OR3 (N23808, N23795, N3413, N7618);
or OR2 (N23809, N23800, N7689);
xor XOR2 (N23810, N23806, N19272);
buf BUF1 (N23811, N23801);
or OR2 (N23812, N23807, N12215);
not NOT1 (N23813, N23787);
xor XOR2 (N23814, N23813, N16021);
and AND4 (N23815, N23810, N11956, N6455, N16064);
xor XOR2 (N23816, N23804, N7299);
and AND3 (N23817, N23805, N15487, N3824);
and AND4 (N23818, N23816, N12762, N10795, N16117);
nand NAND4 (N23819, N23818, N11167, N8404, N13387);
or OR2 (N23820, N23817, N15145);
not NOT1 (N23821, N23815);
nor NOR4 (N23822, N23808, N10475, N13488, N18230);
not NOT1 (N23823, N23814);
and AND2 (N23824, N23819, N23377);
buf BUF1 (N23825, N23822);
nand NAND3 (N23826, N23803, N10275, N12473);
or OR4 (N23827, N23783, N12335, N19117, N1312);
and AND3 (N23828, N23812, N13250, N822);
xor XOR2 (N23829, N23811, N18264);
or OR4 (N23830, N23829, N21863, N6558, N10454);
and AND4 (N23831, N23827, N19325, N12066, N21174);
nor NOR3 (N23832, N23824, N4710, N8192);
nand NAND3 (N23833, N23831, N11518, N4287);
and AND3 (N23834, N23828, N16117, N3763);
xor XOR2 (N23835, N23821, N14718);
nand NAND2 (N23836, N23825, N8042);
nor NOR2 (N23837, N23826, N1944);
xor XOR2 (N23838, N23832, N3396);
or OR4 (N23839, N23837, N5839, N19059, N20793);
not NOT1 (N23840, N23838);
and AND3 (N23841, N23823, N2168, N525);
or OR2 (N23842, N23840, N19845);
nand NAND4 (N23843, N23830, N7244, N1053, N18650);
xor XOR2 (N23844, N23843, N23383);
nor NOR3 (N23845, N23844, N22211, N14418);
xor XOR2 (N23846, N23839, N3215);
buf BUF1 (N23847, N23809);
nand NAND4 (N23848, N23846, N4195, N2668, N19148);
xor XOR2 (N23849, N23842, N1190);
buf BUF1 (N23850, N23835);
buf BUF1 (N23851, N23849);
not NOT1 (N23852, N23845);
and AND2 (N23853, N23848, N5002);
xor XOR2 (N23854, N23851, N19510);
xor XOR2 (N23855, N23854, N15425);
or OR3 (N23856, N23833, N12649, N15089);
nand NAND2 (N23857, N23856, N13036);
and AND2 (N23858, N23852, N18389);
xor XOR2 (N23859, N23858, N22895);
or OR3 (N23860, N23847, N2517, N7574);
not NOT1 (N23861, N23855);
nand NAND3 (N23862, N23857, N7408, N1904);
nand NAND3 (N23863, N23860, N3763, N16513);
nand NAND2 (N23864, N23850, N22645);
and AND2 (N23865, N23864, N15775);
and AND4 (N23866, N23836, N659, N19229, N13771);
buf BUF1 (N23867, N23841);
nand NAND4 (N23868, N23820, N13844, N7873, N1530);
nor NOR2 (N23869, N23834, N12122);
nand NAND4 (N23870, N23867, N23376, N923, N4652);
not NOT1 (N23871, N23859);
or OR2 (N23872, N23863, N7668);
not NOT1 (N23873, N23868);
nor NOR3 (N23874, N23871, N21679, N13009);
xor XOR2 (N23875, N23866, N8666);
nor NOR4 (N23876, N23869, N3707, N2223, N9139);
and AND4 (N23877, N23876, N13031, N2200, N19158);
nor NOR3 (N23878, N23870, N4823, N291);
and AND4 (N23879, N23862, N14249, N8752, N10082);
nand NAND4 (N23880, N23877, N9994, N155, N6853);
or OR3 (N23881, N23872, N10557, N17350);
xor XOR2 (N23882, N23873, N8816);
or OR4 (N23883, N23875, N16310, N23769, N14540);
buf BUF1 (N23884, N23861);
nand NAND4 (N23885, N23874, N12334, N6706, N18805);
buf BUF1 (N23886, N23880);
nand NAND4 (N23887, N23885, N1744, N5722, N22757);
nor NOR3 (N23888, N23878, N10106, N22783);
xor XOR2 (N23889, N23882, N6624);
and AND2 (N23890, N23879, N2982);
or OR4 (N23891, N23889, N18155, N1108, N18216);
not NOT1 (N23892, N23883);
xor XOR2 (N23893, N23887, N15072);
buf BUF1 (N23894, N23893);
or OR2 (N23895, N23853, N2544);
and AND4 (N23896, N23865, N17120, N210, N9772);
buf BUF1 (N23897, N23888);
xor XOR2 (N23898, N23890, N6094);
nand NAND2 (N23899, N23886, N15469);
buf BUF1 (N23900, N23895);
buf BUF1 (N23901, N23897);
and AND3 (N23902, N23901, N20209, N14091);
nand NAND4 (N23903, N23896, N14490, N9345, N11125);
and AND3 (N23904, N23891, N5709, N58);
nor NOR4 (N23905, N23899, N20757, N5894, N8369);
nor NOR3 (N23906, N23902, N15704, N19790);
and AND2 (N23907, N23884, N15583);
nand NAND2 (N23908, N23905, N10570);
xor XOR2 (N23909, N23906, N10368);
buf BUF1 (N23910, N23892);
buf BUF1 (N23911, N23903);
and AND4 (N23912, N23894, N15658, N23527, N16667);
or OR3 (N23913, N23900, N19471, N1743);
or OR3 (N23914, N23911, N20442, N21991);
buf BUF1 (N23915, N23912);
xor XOR2 (N23916, N23907, N17186);
not NOT1 (N23917, N23916);
not NOT1 (N23918, N23904);
nand NAND2 (N23919, N23913, N7398);
xor XOR2 (N23920, N23918, N23878);
nor NOR3 (N23921, N23919, N1641, N23549);
buf BUF1 (N23922, N23920);
xor XOR2 (N23923, N23908, N9649);
xor XOR2 (N23924, N23921, N354);
not NOT1 (N23925, N23924);
buf BUF1 (N23926, N23917);
nor NOR2 (N23927, N23922, N11049);
xor XOR2 (N23928, N23926, N2751);
xor XOR2 (N23929, N23925, N3597);
nor NOR2 (N23930, N23928, N19387);
nand NAND2 (N23931, N23898, N6053);
buf BUF1 (N23932, N23909);
xor XOR2 (N23933, N23930, N8844);
buf BUF1 (N23934, N23914);
xor XOR2 (N23935, N23910, N979);
nor NOR3 (N23936, N23931, N3920, N8426);
and AND4 (N23937, N23881, N9565, N1152, N3630);
nor NOR2 (N23938, N23932, N6697);
and AND4 (N23939, N23929, N9818, N13394, N6940);
and AND2 (N23940, N23934, N18672);
xor XOR2 (N23941, N23936, N11229);
buf BUF1 (N23942, N23938);
nor NOR3 (N23943, N23915, N11599, N13955);
not NOT1 (N23944, N23923);
not NOT1 (N23945, N23937);
nand NAND4 (N23946, N23940, N1419, N14873, N16006);
and AND3 (N23947, N23939, N21571, N15902);
and AND2 (N23948, N23942, N11582);
or OR4 (N23949, N23946, N12645, N13235, N5466);
or OR2 (N23950, N23944, N12663);
or OR2 (N23951, N23945, N21147);
or OR2 (N23952, N23935, N6386);
and AND3 (N23953, N23943, N3602, N14314);
and AND4 (N23954, N23933, N11704, N17259, N9813);
buf BUF1 (N23955, N23954);
nand NAND2 (N23956, N23953, N10111);
or OR4 (N23957, N23955, N5989, N3352, N9304);
and AND2 (N23958, N23957, N8576);
nor NOR3 (N23959, N23950, N19686, N16709);
nand NAND2 (N23960, N23941, N16393);
not NOT1 (N23961, N23959);
not NOT1 (N23962, N23956);
and AND2 (N23963, N23927, N20304);
buf BUF1 (N23964, N23960);
or OR2 (N23965, N23961, N13588);
buf BUF1 (N23966, N23964);
nor NOR2 (N23967, N23948, N21639);
or OR2 (N23968, N23951, N10773);
nor NOR3 (N23969, N23967, N18178, N14080);
nand NAND2 (N23970, N23947, N4924);
nor NOR3 (N23971, N23963, N17983, N18799);
nand NAND2 (N23972, N23966, N19586);
not NOT1 (N23973, N23962);
or OR4 (N23974, N23949, N11272, N18465, N20318);
or OR3 (N23975, N23958, N10857, N23672);
xor XOR2 (N23976, N23974, N4694);
buf BUF1 (N23977, N23970);
buf BUF1 (N23978, N23971);
and AND4 (N23979, N23952, N10015, N17639, N8554);
nand NAND4 (N23980, N23978, N17412, N18601, N17356);
nand NAND4 (N23981, N23968, N3298, N19287, N15570);
buf BUF1 (N23982, N23979);
not NOT1 (N23983, N23975);
and AND2 (N23984, N23981, N21435);
not NOT1 (N23985, N23982);
and AND3 (N23986, N23984, N15772, N5166);
xor XOR2 (N23987, N23972, N19630);
buf BUF1 (N23988, N23976);
xor XOR2 (N23989, N23988, N21850);
or OR3 (N23990, N23985, N21709, N11039);
nor NOR3 (N23991, N23977, N8145, N13881);
nor NOR4 (N23992, N23969, N5369, N21391, N2899);
not NOT1 (N23993, N23989);
or OR2 (N23994, N23965, N20744);
not NOT1 (N23995, N23983);
nand NAND2 (N23996, N23990, N16302);
and AND4 (N23997, N23991, N20913, N317, N963);
not NOT1 (N23998, N23980);
or OR2 (N23999, N23998, N11130);
buf BUF1 (N24000, N23994);
nor NOR4 (N24001, N23996, N21405, N4895, N18733);
and AND4 (N24002, N23992, N2180, N10451, N7243);
or OR2 (N24003, N23995, N15280);
and AND4 (N24004, N24001, N3714, N20711, N9974);
nor NOR4 (N24005, N23973, N5754, N4815, N7192);
or OR3 (N24006, N24003, N1234, N541);
nor NOR2 (N24007, N23993, N16373);
xor XOR2 (N24008, N24005, N10181);
xor XOR2 (N24009, N24006, N12728);
xor XOR2 (N24010, N24009, N23616);
nor NOR3 (N24011, N24008, N2709, N12465);
nor NOR2 (N24012, N24000, N20311);
nor NOR3 (N24013, N24004, N22251, N6717);
xor XOR2 (N24014, N23986, N10661);
nor NOR4 (N24015, N24014, N1133, N18670, N7900);
nand NAND2 (N24016, N24007, N18048);
buf BUF1 (N24017, N23999);
not NOT1 (N24018, N24010);
nor NOR2 (N24019, N24002, N1625);
buf BUF1 (N24020, N24017);
buf BUF1 (N24021, N23987);
or OR4 (N24022, N24018, N22815, N10894, N5749);
nor NOR3 (N24023, N24019, N23663, N14699);
buf BUF1 (N24024, N24020);
and AND3 (N24025, N24013, N3347, N4677);
nor NOR4 (N24026, N24021, N21451, N17218, N20771);
nand NAND2 (N24027, N23997, N4039);
or OR3 (N24028, N24012, N12089, N3458);
nand NAND3 (N24029, N24024, N3352, N14126);
and AND2 (N24030, N24022, N11148);
xor XOR2 (N24031, N24026, N23022);
not NOT1 (N24032, N24029);
or OR2 (N24033, N24027, N5206);
not NOT1 (N24034, N24023);
buf BUF1 (N24035, N24016);
nor NOR3 (N24036, N24032, N21300, N15119);
nand NAND2 (N24037, N24034, N17073);
nand NAND2 (N24038, N24035, N15922);
xor XOR2 (N24039, N24028, N519);
nor NOR2 (N24040, N24038, N1180);
or OR4 (N24041, N24036, N7428, N7271, N15968);
or OR4 (N24042, N24011, N23073, N16357, N3924);
nand NAND4 (N24043, N24037, N20144, N19328, N7499);
and AND2 (N24044, N24015, N15716);
nand NAND2 (N24045, N24043, N7923);
or OR2 (N24046, N24030, N7528);
nand NAND2 (N24047, N24025, N15489);
nor NOR3 (N24048, N24046, N2592, N8898);
or OR2 (N24049, N24040, N22758);
buf BUF1 (N24050, N24033);
nand NAND2 (N24051, N24048, N12978);
and AND4 (N24052, N24041, N11789, N4522, N7196);
not NOT1 (N24053, N24051);
or OR2 (N24054, N24042, N22459);
buf BUF1 (N24055, N24039);
nand NAND2 (N24056, N24045, N11647);
buf BUF1 (N24057, N24047);
and AND4 (N24058, N24050, N22833, N22062, N8682);
or OR3 (N24059, N24056, N16045, N17579);
nand NAND4 (N24060, N24049, N18169, N17423, N7326);
nor NOR3 (N24061, N24052, N4223, N24003);
buf BUF1 (N24062, N24055);
buf BUF1 (N24063, N24059);
and AND4 (N24064, N24031, N8078, N20909, N20662);
nand NAND2 (N24065, N24060, N2307);
buf BUF1 (N24066, N24064);
and AND3 (N24067, N24066, N19494, N12321);
not NOT1 (N24068, N24067);
xor XOR2 (N24069, N24068, N18219);
nor NOR2 (N24070, N24061, N23324);
nand NAND2 (N24071, N24054, N18042);
and AND4 (N24072, N24063, N21658, N16453, N17390);
and AND2 (N24073, N24053, N22060);
and AND4 (N24074, N24065, N9440, N13197, N6402);
buf BUF1 (N24075, N24069);
not NOT1 (N24076, N24070);
xor XOR2 (N24077, N24073, N20455);
xor XOR2 (N24078, N24044, N2826);
and AND4 (N24079, N24076, N19631, N8189, N4853);
and AND4 (N24080, N24077, N15838, N8458, N3134);
not NOT1 (N24081, N24057);
and AND4 (N24082, N24078, N10956, N11441, N8127);
xor XOR2 (N24083, N24081, N8739);
and AND4 (N24084, N24080, N15902, N1270, N1472);
buf BUF1 (N24085, N24075);
and AND3 (N24086, N24074, N14595, N23224);
xor XOR2 (N24087, N24072, N6572);
or OR2 (N24088, N24079, N2359);
nor NOR4 (N24089, N24058, N11201, N10582, N21684);
or OR4 (N24090, N24071, N5502, N15024, N13841);
or OR3 (N24091, N24084, N13742, N2585);
or OR3 (N24092, N24086, N17466, N1227);
or OR3 (N24093, N24089, N2504, N9383);
xor XOR2 (N24094, N24085, N16556);
nand NAND2 (N24095, N24082, N22648);
or OR3 (N24096, N24094, N11767, N13483);
or OR4 (N24097, N24088, N22611, N14806, N5012);
not NOT1 (N24098, N24096);
nand NAND2 (N24099, N24083, N17405);
xor XOR2 (N24100, N24087, N22679);
and AND2 (N24101, N24090, N8194);
nor NOR3 (N24102, N24095, N23427, N4665);
or OR3 (N24103, N24062, N19306, N12869);
or OR4 (N24104, N24093, N22069, N3334, N1352);
or OR3 (N24105, N24091, N22127, N4656);
buf BUF1 (N24106, N24101);
and AND4 (N24107, N24104, N9833, N7647, N3397);
xor XOR2 (N24108, N24097, N22469);
and AND4 (N24109, N24108, N20185, N20298, N21316);
or OR4 (N24110, N24100, N8925, N14193, N16747);
nand NAND3 (N24111, N24109, N10327, N1651);
not NOT1 (N24112, N24092);
buf BUF1 (N24113, N24110);
nand NAND2 (N24114, N24111, N9068);
or OR2 (N24115, N24113, N21754);
and AND3 (N24116, N24098, N10194, N23441);
not NOT1 (N24117, N24107);
not NOT1 (N24118, N24103);
or OR4 (N24119, N24116, N3415, N5471, N11892);
nor NOR4 (N24120, N24118, N22665, N7650, N22229);
nand NAND2 (N24121, N24120, N13152);
buf BUF1 (N24122, N24121);
nand NAND4 (N24123, N24105, N23889, N21360, N21515);
nand NAND3 (N24124, N24114, N14708, N17797);
xor XOR2 (N24125, N24123, N669);
nor NOR2 (N24126, N24099, N6121);
nand NAND3 (N24127, N24117, N21479, N2692);
not NOT1 (N24128, N24127);
buf BUF1 (N24129, N24119);
xor XOR2 (N24130, N24122, N20447);
nand NAND3 (N24131, N24125, N21993, N5888);
nor NOR4 (N24132, N24124, N14149, N10689, N19039);
buf BUF1 (N24133, N24106);
not NOT1 (N24134, N24126);
nand NAND3 (N24135, N24128, N5548, N14873);
not NOT1 (N24136, N24132);
xor XOR2 (N24137, N24134, N12089);
not NOT1 (N24138, N24129);
not NOT1 (N24139, N24137);
not NOT1 (N24140, N24138);
or OR3 (N24141, N24131, N5956, N2882);
or OR3 (N24142, N24130, N6867, N596);
or OR3 (N24143, N24112, N2024, N14985);
or OR4 (N24144, N24136, N9958, N11164, N6737);
not NOT1 (N24145, N24139);
xor XOR2 (N24146, N24102, N13886);
nor NOR4 (N24147, N24140, N20547, N4617, N2232);
buf BUF1 (N24148, N24141);
nor NOR4 (N24149, N24144, N16028, N19735, N6486);
buf BUF1 (N24150, N24149);
or OR4 (N24151, N24135, N8819, N2656, N10822);
xor XOR2 (N24152, N24143, N23037);
buf BUF1 (N24153, N24115);
nor NOR3 (N24154, N24152, N20223, N9604);
nand NAND2 (N24155, N24142, N22408);
and AND4 (N24156, N24147, N7593, N21270, N14928);
buf BUF1 (N24157, N24151);
and AND2 (N24158, N24153, N10771);
xor XOR2 (N24159, N24146, N4856);
xor XOR2 (N24160, N24157, N21482);
not NOT1 (N24161, N24158);
and AND2 (N24162, N24161, N17598);
or OR2 (N24163, N24162, N10097);
xor XOR2 (N24164, N24156, N6904);
and AND2 (N24165, N24133, N18377);
not NOT1 (N24166, N24159);
and AND3 (N24167, N24148, N15532, N13603);
buf BUF1 (N24168, N24163);
buf BUF1 (N24169, N24154);
xor XOR2 (N24170, N24166, N3948);
buf BUF1 (N24171, N24160);
buf BUF1 (N24172, N24167);
buf BUF1 (N24173, N24172);
nand NAND3 (N24174, N24170, N22076, N7212);
buf BUF1 (N24175, N24174);
nor NOR4 (N24176, N24155, N2575, N19069, N16592);
xor XOR2 (N24177, N24169, N18539);
or OR3 (N24178, N24175, N2949, N17805);
xor XOR2 (N24179, N24173, N238);
nor NOR3 (N24180, N24150, N13, N4059);
nand NAND4 (N24181, N24145, N6406, N6817, N2355);
nand NAND2 (N24182, N24177, N17459);
nand NAND2 (N24183, N24178, N126);
nand NAND3 (N24184, N24164, N18365, N7669);
xor XOR2 (N24185, N24168, N20691);
or OR2 (N24186, N24181, N14475);
nor NOR3 (N24187, N24176, N2117, N22365);
or OR2 (N24188, N24183, N19193);
and AND2 (N24189, N24187, N19549);
and AND3 (N24190, N24182, N20167, N9809);
or OR3 (N24191, N24184, N10146, N9557);
buf BUF1 (N24192, N24191);
buf BUF1 (N24193, N24186);
and AND3 (N24194, N24188, N11001, N1090);
not NOT1 (N24195, N24179);
or OR4 (N24196, N24194, N7405, N20004, N10820);
buf BUF1 (N24197, N24165);
nand NAND3 (N24198, N24192, N12142, N24187);
not NOT1 (N24199, N24171);
and AND2 (N24200, N24193, N20090);
nor NOR4 (N24201, N24199, N14049, N1672, N12950);
or OR2 (N24202, N24201, N16053);
nor NOR4 (N24203, N24202, N9206, N7730, N16699);
or OR3 (N24204, N24198, N2796, N18193);
and AND4 (N24205, N24197, N19906, N8719, N23204);
and AND3 (N24206, N24180, N12168, N3536);
or OR3 (N24207, N24190, N20312, N4127);
and AND3 (N24208, N24204, N11124, N3783);
nor NOR3 (N24209, N24203, N24098, N4815);
and AND3 (N24210, N24208, N3778, N2033);
or OR3 (N24211, N24189, N2343, N7073);
xor XOR2 (N24212, N24195, N6841);
nand NAND4 (N24213, N24196, N22354, N18606, N1872);
or OR4 (N24214, N24185, N12057, N15912, N1023);
xor XOR2 (N24215, N24214, N16423);
nor NOR4 (N24216, N24200, N23249, N15929, N17395);
and AND2 (N24217, N24207, N19769);
and AND2 (N24218, N24217, N21944);
xor XOR2 (N24219, N24213, N23402);
buf BUF1 (N24220, N24216);
nor NOR2 (N24221, N24212, N18638);
buf BUF1 (N24222, N24209);
not NOT1 (N24223, N24219);
or OR3 (N24224, N24223, N12630, N14955);
nand NAND4 (N24225, N24221, N915, N11629, N2685);
not NOT1 (N24226, N24220);
nand NAND2 (N24227, N24211, N785);
not NOT1 (N24228, N24227);
and AND4 (N24229, N24224, N20289, N8702, N10603);
nor NOR2 (N24230, N24206, N20867);
or OR4 (N24231, N24215, N15354, N23689, N5089);
nand NAND4 (N24232, N24210, N19940, N4957, N22991);
xor XOR2 (N24233, N24232, N23704);
not NOT1 (N24234, N24231);
nand NAND2 (N24235, N24222, N23097);
xor XOR2 (N24236, N24235, N22965);
buf BUF1 (N24237, N24225);
and AND2 (N24238, N24237, N12809);
nand NAND4 (N24239, N24228, N12446, N18030, N10814);
xor XOR2 (N24240, N24233, N8971);
nand NAND2 (N24241, N24205, N3128);
xor XOR2 (N24242, N24238, N4232);
xor XOR2 (N24243, N24236, N22385);
nor NOR2 (N24244, N24241, N21520);
nand NAND3 (N24245, N24240, N15498, N21168);
nor NOR4 (N24246, N24239, N9363, N2514, N15710);
not NOT1 (N24247, N24244);
nor NOR2 (N24248, N24226, N3709);
xor XOR2 (N24249, N24242, N22556);
not NOT1 (N24250, N24243);
buf BUF1 (N24251, N24234);
buf BUF1 (N24252, N24250);
not NOT1 (N24253, N24229);
nand NAND3 (N24254, N24218, N1662, N2681);
or OR2 (N24255, N24245, N2398);
not NOT1 (N24256, N24247);
and AND3 (N24257, N24246, N13966, N15664);
nor NOR2 (N24258, N24252, N12203);
and AND3 (N24259, N24256, N14108, N21954);
nor NOR2 (N24260, N24248, N4216);
buf BUF1 (N24261, N24251);
xor XOR2 (N24262, N24249, N6430);
and AND4 (N24263, N24230, N20347, N11835, N7388);
not NOT1 (N24264, N24261);
xor XOR2 (N24265, N24258, N18734);
buf BUF1 (N24266, N24262);
not NOT1 (N24267, N24266);
nand NAND4 (N24268, N24263, N23588, N2367, N11877);
nor NOR3 (N24269, N24264, N14358, N14778);
and AND4 (N24270, N24260, N5655, N8292, N18008);
and AND4 (N24271, N24267, N23979, N7236, N12012);
and AND2 (N24272, N24271, N22540);
xor XOR2 (N24273, N24255, N23436);
nand NAND2 (N24274, N24265, N13704);
and AND3 (N24275, N24269, N4063, N19710);
xor XOR2 (N24276, N24259, N10715);
not NOT1 (N24277, N24254);
buf BUF1 (N24278, N24253);
buf BUF1 (N24279, N24268);
nor NOR4 (N24280, N24275, N13294, N22195, N22453);
or OR4 (N24281, N24280, N4366, N23038, N3774);
xor XOR2 (N24282, N24278, N17325);
buf BUF1 (N24283, N24281);
buf BUF1 (N24284, N24272);
or OR2 (N24285, N24282, N14969);
nand NAND2 (N24286, N24285, N7480);
and AND3 (N24287, N24283, N23036, N4379);
not NOT1 (N24288, N24273);
nand NAND2 (N24289, N24257, N21890);
nand NAND4 (N24290, N24287, N4118, N1677, N19787);
not NOT1 (N24291, N24289);
nand NAND3 (N24292, N24290, N9336, N4208);
buf BUF1 (N24293, N24288);
or OR2 (N24294, N24277, N2952);
xor XOR2 (N24295, N24276, N7488);
and AND2 (N24296, N24270, N16289);
or OR3 (N24297, N24291, N14017, N11713);
xor XOR2 (N24298, N24295, N23300);
buf BUF1 (N24299, N24286);
xor XOR2 (N24300, N24274, N13227);
and AND3 (N24301, N24294, N11207, N13787);
and AND4 (N24302, N24301, N4411, N21981, N7767);
and AND2 (N24303, N24298, N4734);
nor NOR2 (N24304, N24303, N3946);
not NOT1 (N24305, N24292);
nand NAND4 (N24306, N24299, N6920, N19006, N8996);
nand NAND4 (N24307, N24296, N16862, N11379, N13099);
not NOT1 (N24308, N24305);
and AND4 (N24309, N24308, N22475, N8138, N6499);
not NOT1 (N24310, N24300);
and AND3 (N24311, N24310, N12174, N5394);
or OR2 (N24312, N24307, N10696);
and AND4 (N24313, N24311, N8113, N18506, N13170);
nor NOR2 (N24314, N24312, N19713);
not NOT1 (N24315, N24284);
buf BUF1 (N24316, N24306);
nand NAND3 (N24317, N24302, N14005, N8425);
nor NOR2 (N24318, N24316, N22635);
xor XOR2 (N24319, N24293, N4259);
or OR2 (N24320, N24318, N3287);
not NOT1 (N24321, N24297);
xor XOR2 (N24322, N24304, N6278);
and AND3 (N24323, N24322, N225, N7015);
xor XOR2 (N24324, N24320, N17485);
or OR3 (N24325, N24314, N5768, N18174);
and AND2 (N24326, N24317, N7399);
and AND2 (N24327, N24313, N19043);
not NOT1 (N24328, N24319);
nand NAND3 (N24329, N24324, N1158, N9382);
xor XOR2 (N24330, N24328, N21080);
nand NAND2 (N24331, N24327, N6843);
xor XOR2 (N24332, N24325, N14463);
or OR3 (N24333, N24323, N18398, N13628);
nor NOR4 (N24334, N24326, N23285, N22893, N5294);
and AND4 (N24335, N24332, N13184, N1907, N13634);
xor XOR2 (N24336, N24334, N22110);
not NOT1 (N24337, N24279);
xor XOR2 (N24338, N24321, N12436);
not NOT1 (N24339, N24335);
buf BUF1 (N24340, N24330);
nand NAND4 (N24341, N24333, N221, N4284, N5750);
nor NOR3 (N24342, N24315, N22527, N23646);
buf BUF1 (N24343, N24342);
xor XOR2 (N24344, N24338, N22417);
nor NOR4 (N24345, N24343, N10286, N4784, N2081);
not NOT1 (N24346, N24336);
not NOT1 (N24347, N24339);
xor XOR2 (N24348, N24344, N9957);
not NOT1 (N24349, N24309);
xor XOR2 (N24350, N24349, N3200);
not NOT1 (N24351, N24331);
nor NOR3 (N24352, N24329, N10653, N6153);
or OR2 (N24353, N24352, N14230);
or OR2 (N24354, N24337, N20079);
xor XOR2 (N24355, N24351, N15226);
nand NAND2 (N24356, N24341, N18565);
and AND4 (N24357, N24345, N1114, N16879, N19356);
nand NAND3 (N24358, N24348, N9733, N8325);
and AND3 (N24359, N24340, N12548, N4991);
not NOT1 (N24360, N24357);
or OR3 (N24361, N24356, N22174, N4076);
or OR4 (N24362, N24346, N7539, N24305, N14064);
or OR4 (N24363, N24347, N6272, N18766, N4621);
or OR2 (N24364, N24363, N8123);
or OR4 (N24365, N24350, N21511, N6586, N17166);
nand NAND2 (N24366, N24361, N10510);
nand NAND2 (N24367, N24365, N4298);
and AND3 (N24368, N24366, N18035, N13315);
or OR4 (N24369, N24367, N9969, N16733, N21607);
and AND3 (N24370, N24369, N12886, N4726);
nor NOR4 (N24371, N24359, N7520, N6115, N2804);
buf BUF1 (N24372, N24354);
xor XOR2 (N24373, N24353, N10123);
buf BUF1 (N24374, N24371);
nand NAND4 (N24375, N24360, N3694, N5074, N2362);
nand NAND3 (N24376, N24364, N11347, N11219);
nand NAND3 (N24377, N24374, N23201, N14214);
nand NAND2 (N24378, N24372, N3055);
or OR3 (N24379, N24358, N12326, N7439);
xor XOR2 (N24380, N24379, N9702);
or OR3 (N24381, N24377, N18550, N7646);
and AND2 (N24382, N24362, N12939);
or OR3 (N24383, N24376, N16016, N15400);
buf BUF1 (N24384, N24373);
not NOT1 (N24385, N24355);
not NOT1 (N24386, N24383);
nor NOR2 (N24387, N24368, N15709);
or OR2 (N24388, N24370, N4313);
nand NAND4 (N24389, N24382, N9448, N10374, N6033);
xor XOR2 (N24390, N24387, N16029);
nor NOR2 (N24391, N24388, N4196);
not NOT1 (N24392, N24384);
or OR4 (N24393, N24378, N1305, N8537, N8339);
not NOT1 (N24394, N24391);
xor XOR2 (N24395, N24390, N365);
or OR3 (N24396, N24386, N6630, N6662);
nor NOR3 (N24397, N24375, N12385, N449);
nand NAND2 (N24398, N24394, N9107);
nand NAND4 (N24399, N24397, N22987, N13940, N14022);
buf BUF1 (N24400, N24385);
nor NOR4 (N24401, N24395, N14008, N3806, N7994);
buf BUF1 (N24402, N24393);
or OR4 (N24403, N24380, N6062, N18230, N20171);
nand NAND4 (N24404, N24402, N13867, N563, N11649);
nand NAND2 (N24405, N24400, N7051);
nor NOR4 (N24406, N24389, N14492, N11430, N10572);
not NOT1 (N24407, N24399);
not NOT1 (N24408, N24407);
and AND3 (N24409, N24408, N12675, N7336);
and AND4 (N24410, N24381, N24032, N20594, N12294);
nor NOR4 (N24411, N24392, N22895, N14063, N22934);
nor NOR4 (N24412, N24411, N5515, N8559, N16812);
xor XOR2 (N24413, N24396, N16619);
and AND3 (N24414, N24405, N5381, N19178);
xor XOR2 (N24415, N24409, N20530);
buf BUF1 (N24416, N24403);
buf BUF1 (N24417, N24412);
not NOT1 (N24418, N24406);
xor XOR2 (N24419, N24410, N16971);
buf BUF1 (N24420, N24404);
or OR4 (N24421, N24418, N17252, N1885, N9986);
and AND3 (N24422, N24417, N24095, N9114);
nor NOR2 (N24423, N24420, N3636);
nor NOR2 (N24424, N24415, N2360);
and AND3 (N24425, N24413, N13399, N10554);
or OR3 (N24426, N24422, N6478, N15221);
nand NAND4 (N24427, N24424, N17448, N19108, N19894);
not NOT1 (N24428, N24401);
xor XOR2 (N24429, N24423, N18230);
or OR2 (N24430, N24425, N10596);
buf BUF1 (N24431, N24414);
not NOT1 (N24432, N24419);
and AND3 (N24433, N24432, N20581, N15935);
buf BUF1 (N24434, N24430);
buf BUF1 (N24435, N24434);
buf BUF1 (N24436, N24431);
xor XOR2 (N24437, N24428, N3293);
and AND2 (N24438, N24398, N3741);
xor XOR2 (N24439, N24416, N661);
buf BUF1 (N24440, N24437);
nand NAND2 (N24441, N24426, N11381);
not NOT1 (N24442, N24439);
buf BUF1 (N24443, N24433);
and AND2 (N24444, N24427, N22929);
or OR3 (N24445, N24436, N21230, N9451);
or OR3 (N24446, N24429, N19078, N5530);
nand NAND2 (N24447, N24443, N14316);
nor NOR2 (N24448, N24446, N8571);
buf BUF1 (N24449, N24441);
not NOT1 (N24450, N24435);
or OR4 (N24451, N24438, N12638, N15321, N15853);
buf BUF1 (N24452, N24442);
nor NOR2 (N24453, N24444, N23392);
not NOT1 (N24454, N24421);
nor NOR3 (N24455, N24448, N644, N18930);
not NOT1 (N24456, N24449);
or OR4 (N24457, N24447, N2645, N12120, N7676);
or OR3 (N24458, N24440, N9000, N12349);
or OR4 (N24459, N24456, N18396, N13264, N18057);
buf BUF1 (N24460, N24453);
not NOT1 (N24461, N24457);
not NOT1 (N24462, N24461);
buf BUF1 (N24463, N24445);
xor XOR2 (N24464, N24462, N15185);
nor NOR4 (N24465, N24450, N6977, N14419, N7645);
or OR2 (N24466, N24459, N17435);
and AND3 (N24467, N24463, N6604, N12284);
nor NOR2 (N24468, N24455, N20013);
xor XOR2 (N24469, N24466, N21829);
not NOT1 (N24470, N24454);
buf BUF1 (N24471, N24451);
and AND4 (N24472, N24460, N11370, N2195, N10083);
and AND3 (N24473, N24452, N13247, N12635);
xor XOR2 (N24474, N24464, N18531);
nand NAND4 (N24475, N24471, N23706, N2723, N12216);
nor NOR4 (N24476, N24469, N20823, N2345, N22338);
nand NAND3 (N24477, N24470, N3331, N15847);
xor XOR2 (N24478, N24468, N20118);
not NOT1 (N24479, N24465);
xor XOR2 (N24480, N24475, N16386);
xor XOR2 (N24481, N24458, N20057);
nor NOR4 (N24482, N24480, N3100, N20743, N11278);
nand NAND2 (N24483, N24477, N22048);
not NOT1 (N24484, N24482);
xor XOR2 (N24485, N24481, N20480);
or OR4 (N24486, N24474, N16837, N19049, N359);
buf BUF1 (N24487, N24473);
xor XOR2 (N24488, N24484, N8107);
buf BUF1 (N24489, N24472);
not NOT1 (N24490, N24487);
nor NOR2 (N24491, N24467, N20415);
and AND3 (N24492, N24483, N7867, N10405);
xor XOR2 (N24493, N24479, N23847);
or OR4 (N24494, N24492, N14171, N14684, N21159);
or OR3 (N24495, N24489, N6131, N17579);
xor XOR2 (N24496, N24495, N12525);
nor NOR3 (N24497, N24486, N23490, N22226);
not NOT1 (N24498, N24497);
not NOT1 (N24499, N24493);
xor XOR2 (N24500, N24488, N15232);
xor XOR2 (N24501, N24496, N18293);
and AND4 (N24502, N24478, N3418, N6287, N18599);
or OR3 (N24503, N24501, N21843, N16850);
buf BUF1 (N24504, N24498);
not NOT1 (N24505, N24499);
xor XOR2 (N24506, N24505, N21185);
and AND2 (N24507, N24500, N6395);
or OR3 (N24508, N24494, N21221, N7393);
and AND4 (N24509, N24502, N12121, N7661, N23912);
xor XOR2 (N24510, N24504, N22333);
nor NOR3 (N24511, N24491, N8890, N18364);
and AND4 (N24512, N24509, N14652, N538, N12516);
nand NAND3 (N24513, N24503, N19498, N13507);
xor XOR2 (N24514, N24485, N14212);
xor XOR2 (N24515, N24476, N22115);
nor NOR4 (N24516, N24512, N9438, N5990, N8633);
xor XOR2 (N24517, N24515, N14691);
nand NAND3 (N24518, N24517, N8495, N14693);
xor XOR2 (N24519, N24507, N18140);
xor XOR2 (N24520, N24516, N18062);
not NOT1 (N24521, N24519);
and AND2 (N24522, N24506, N690);
or OR2 (N24523, N24518, N19805);
and AND4 (N24524, N24521, N9694, N5394, N12131);
or OR3 (N24525, N24490, N22473, N18345);
xor XOR2 (N24526, N24523, N11261);
xor XOR2 (N24527, N24522, N5124);
and AND2 (N24528, N24511, N23422);
and AND4 (N24529, N24510, N17448, N15294, N17309);
or OR3 (N24530, N24508, N7436, N2534);
nor NOR4 (N24531, N24530, N5868, N9858, N5369);
or OR2 (N24532, N24528, N3159);
buf BUF1 (N24533, N24524);
or OR3 (N24534, N24525, N23562, N452);
or OR4 (N24535, N24532, N13015, N1419, N19783);
nand NAND4 (N24536, N24513, N22643, N7417, N6121);
nor NOR3 (N24537, N24520, N21644, N4815);
or OR4 (N24538, N24514, N8141, N18512, N22248);
or OR4 (N24539, N24534, N7251, N6651, N21901);
nand NAND4 (N24540, N24533, N6066, N15755, N22159);
nand NAND3 (N24541, N24538, N7346, N1099);
not NOT1 (N24542, N24531);
nand NAND4 (N24543, N24536, N19516, N4826, N16140);
or OR2 (N24544, N24535, N10171);
xor XOR2 (N24545, N24527, N3403);
and AND3 (N24546, N24540, N8703, N13980);
not NOT1 (N24547, N24546);
nor NOR4 (N24548, N24529, N9180, N11168, N13991);
not NOT1 (N24549, N24537);
buf BUF1 (N24550, N24544);
nand NAND2 (N24551, N24548, N5049);
buf BUF1 (N24552, N24539);
and AND3 (N24553, N24542, N19656, N7138);
nand NAND4 (N24554, N24552, N10535, N10712, N11019);
nand NAND2 (N24555, N24545, N1895);
and AND2 (N24556, N24550, N1855);
not NOT1 (N24557, N24555);
nor NOR4 (N24558, N24551, N7123, N2741, N17585);
nor NOR2 (N24559, N24557, N15787);
or OR4 (N24560, N24543, N12740, N13030, N2204);
buf BUF1 (N24561, N24556);
xor XOR2 (N24562, N24526, N4307);
not NOT1 (N24563, N24549);
and AND4 (N24564, N24541, N8429, N19842, N12602);
nand NAND2 (N24565, N24547, N178);
xor XOR2 (N24566, N24558, N9705);
and AND3 (N24567, N24562, N20720, N18948);
not NOT1 (N24568, N24561);
not NOT1 (N24569, N24559);
not NOT1 (N24570, N24567);
nor NOR3 (N24571, N24564, N15846, N8866);
nor NOR4 (N24572, N24569, N6589, N12117, N3525);
xor XOR2 (N24573, N24553, N904);
buf BUF1 (N24574, N24560);
or OR2 (N24575, N24571, N2567);
nor NOR2 (N24576, N24565, N1035);
and AND2 (N24577, N24574, N1338);
xor XOR2 (N24578, N24573, N21641);
xor XOR2 (N24579, N24572, N14053);
buf BUF1 (N24580, N24554);
buf BUF1 (N24581, N24577);
not NOT1 (N24582, N24563);
xor XOR2 (N24583, N24579, N22209);
nor NOR3 (N24584, N24566, N15599, N24409);
or OR3 (N24585, N24570, N20301, N19338);
not NOT1 (N24586, N24581);
xor XOR2 (N24587, N24580, N2239);
and AND4 (N24588, N24586, N22599, N11037, N14467);
buf BUF1 (N24589, N24584);
or OR4 (N24590, N24582, N20983, N20109, N7953);
not NOT1 (N24591, N24589);
and AND2 (N24592, N24575, N397);
or OR3 (N24593, N24587, N17854, N23444);
nor NOR4 (N24594, N24585, N24516, N9566, N8393);
or OR2 (N24595, N24593, N13850);
and AND3 (N24596, N24595, N10390, N1355);
nor NOR3 (N24597, N24590, N4704, N9855);
nor NOR3 (N24598, N24588, N22758, N14881);
buf BUF1 (N24599, N24576);
not NOT1 (N24600, N24597);
nand NAND2 (N24601, N24578, N7988);
nor NOR3 (N24602, N24600, N14889, N12341);
buf BUF1 (N24603, N24591);
not NOT1 (N24604, N24568);
and AND2 (N24605, N24602, N1942);
buf BUF1 (N24606, N24604);
or OR2 (N24607, N24601, N21758);
not NOT1 (N24608, N24605);
xor XOR2 (N24609, N24594, N11484);
and AND2 (N24610, N24583, N5710);
not NOT1 (N24611, N24606);
not NOT1 (N24612, N24610);
not NOT1 (N24613, N24608);
nand NAND2 (N24614, N24598, N18837);
xor XOR2 (N24615, N24611, N19041);
buf BUF1 (N24616, N24612);
and AND4 (N24617, N24616, N13533, N21855, N11013);
buf BUF1 (N24618, N24609);
nand NAND2 (N24619, N24617, N24108);
and AND3 (N24620, N24614, N22872, N2335);
xor XOR2 (N24621, N24607, N13666);
or OR4 (N24622, N24596, N12990, N22178, N12039);
xor XOR2 (N24623, N24620, N19214);
not NOT1 (N24624, N24615);
or OR3 (N24625, N24592, N272, N16924);
xor XOR2 (N24626, N24622, N2376);
and AND4 (N24627, N24626, N12943, N18880, N18799);
xor XOR2 (N24628, N24619, N10686);
buf BUF1 (N24629, N24628);
and AND2 (N24630, N24623, N11669);
nor NOR3 (N24631, N24630, N8383, N11193);
and AND4 (N24632, N24621, N17884, N17160, N1266);
xor XOR2 (N24633, N24603, N8365);
buf BUF1 (N24634, N24618);
and AND4 (N24635, N24625, N22582, N9276, N3790);
and AND4 (N24636, N24627, N18177, N13465, N18397);
xor XOR2 (N24637, N24633, N1695);
or OR4 (N24638, N24635, N23182, N7724, N8854);
buf BUF1 (N24639, N24636);
nand NAND4 (N24640, N24639, N20446, N23660, N1533);
buf BUF1 (N24641, N24624);
and AND2 (N24642, N24632, N11352);
and AND2 (N24643, N24638, N24368);
and AND2 (N24644, N24642, N18552);
nor NOR4 (N24645, N24643, N15651, N15522, N184);
not NOT1 (N24646, N24644);
not NOT1 (N24647, N24613);
xor XOR2 (N24648, N24645, N18531);
buf BUF1 (N24649, N24634);
or OR4 (N24650, N24629, N19953, N3018, N16066);
not NOT1 (N24651, N24641);
not NOT1 (N24652, N24637);
or OR2 (N24653, N24652, N13745);
buf BUF1 (N24654, N24599);
xor XOR2 (N24655, N24650, N10735);
and AND2 (N24656, N24651, N4391);
nor NOR3 (N24657, N24649, N15094, N669);
or OR2 (N24658, N24631, N23963);
nor NOR3 (N24659, N24653, N219, N7935);
and AND4 (N24660, N24656, N20565, N22177, N9207);
buf BUF1 (N24661, N24655);
nor NOR3 (N24662, N24654, N16210, N6869);
nor NOR2 (N24663, N24647, N2099);
or OR3 (N24664, N24662, N11651, N21900);
or OR2 (N24665, N24646, N5217);
or OR4 (N24666, N24658, N3080, N23661, N24187);
and AND4 (N24667, N24665, N23268, N878, N22756);
buf BUF1 (N24668, N24657);
xor XOR2 (N24669, N24668, N15514);
nor NOR3 (N24670, N24666, N23712, N208);
or OR2 (N24671, N24640, N14411);
or OR2 (N24672, N24648, N1028);
buf BUF1 (N24673, N24667);
and AND4 (N24674, N24663, N24260, N3479, N13215);
xor XOR2 (N24675, N24661, N22334);
buf BUF1 (N24676, N24674);
nor NOR3 (N24677, N24660, N18885, N13765);
xor XOR2 (N24678, N24675, N8981);
nand NAND3 (N24679, N24659, N3996, N8851);
not NOT1 (N24680, N24678);
buf BUF1 (N24681, N24673);
buf BUF1 (N24682, N24672);
xor XOR2 (N24683, N24679, N13390);
not NOT1 (N24684, N24681);
not NOT1 (N24685, N24676);
not NOT1 (N24686, N24670);
or OR4 (N24687, N24669, N18621, N6605, N13164);
not NOT1 (N24688, N24684);
nand NAND2 (N24689, N24683, N17539);
buf BUF1 (N24690, N24677);
not NOT1 (N24691, N24689);
or OR2 (N24692, N24688, N22436);
and AND4 (N24693, N24664, N12962, N15570, N23739);
buf BUF1 (N24694, N24693);
buf BUF1 (N24695, N24692);
xor XOR2 (N24696, N24695, N15877);
and AND2 (N24697, N24694, N18528);
not NOT1 (N24698, N24680);
buf BUF1 (N24699, N24671);
and AND3 (N24700, N24687, N15930, N8735);
nor NOR4 (N24701, N24686, N12217, N23841, N9778);
and AND4 (N24702, N24697, N6033, N13614, N13839);
and AND4 (N24703, N24701, N4870, N14392, N3168);
nand NAND4 (N24704, N24698, N4174, N11470, N24055);
nand NAND2 (N24705, N24682, N2625);
nor NOR2 (N24706, N24699, N12973);
buf BUF1 (N24707, N24691);
nand NAND2 (N24708, N24707, N12760);
or OR4 (N24709, N24703, N15819, N14732, N21810);
nand NAND3 (N24710, N24702, N18333, N17686);
and AND4 (N24711, N24690, N5064, N5195, N18278);
nand NAND2 (N24712, N24696, N3080);
nand NAND3 (N24713, N24685, N9863, N4336);
buf BUF1 (N24714, N24709);
nand NAND4 (N24715, N24711, N10383, N13624, N17211);
or OR3 (N24716, N24714, N4021, N11102);
nand NAND3 (N24717, N24706, N2236, N619);
and AND3 (N24718, N24712, N11333, N5832);
xor XOR2 (N24719, N24708, N14521);
xor XOR2 (N24720, N24700, N23770);
xor XOR2 (N24721, N24720, N750);
xor XOR2 (N24722, N24718, N19098);
nor NOR4 (N24723, N24719, N14442, N23795, N15443);
and AND2 (N24724, N24710, N9074);
buf BUF1 (N24725, N24713);
xor XOR2 (N24726, N24717, N330);
not NOT1 (N24727, N24715);
not NOT1 (N24728, N24726);
buf BUF1 (N24729, N24722);
nand NAND2 (N24730, N24724, N16076);
and AND2 (N24731, N24727, N22385);
nor NOR3 (N24732, N24731, N3071, N16744);
nand NAND3 (N24733, N24725, N19854, N23289);
nand NAND4 (N24734, N24733, N12769, N10525, N6971);
nand NAND2 (N24735, N24728, N23501);
and AND3 (N24736, N24716, N14586, N8318);
nand NAND2 (N24737, N24723, N16958);
xor XOR2 (N24738, N24729, N20017);
nor NOR2 (N24739, N24705, N18115);
nand NAND2 (N24740, N24732, N3528);
buf BUF1 (N24741, N24734);
or OR4 (N24742, N24735, N23311, N1712, N6473);
buf BUF1 (N24743, N24730);
nand NAND3 (N24744, N24740, N2933, N19077);
xor XOR2 (N24745, N24721, N23646);
not NOT1 (N24746, N24739);
buf BUF1 (N24747, N24741);
nand NAND4 (N24748, N24736, N13963, N20905, N783);
or OR2 (N24749, N24738, N2761);
buf BUF1 (N24750, N24704);
nand NAND2 (N24751, N24750, N21452);
nand NAND4 (N24752, N24747, N8898, N3528, N5767);
nor NOR4 (N24753, N24752, N8820, N19893, N6807);
or OR2 (N24754, N24753, N21408);
nand NAND2 (N24755, N24742, N23293);
and AND3 (N24756, N24755, N5562, N10957);
or OR3 (N24757, N24756, N13779, N7743);
xor XOR2 (N24758, N24749, N18239);
nor NOR3 (N24759, N24743, N17235, N4598);
and AND4 (N24760, N24737, N4567, N10551, N290);
or OR4 (N24761, N24754, N4274, N5271, N13577);
nand NAND4 (N24762, N24759, N1170, N13398, N19153);
xor XOR2 (N24763, N24751, N23268);
and AND4 (N24764, N24758, N3552, N20150, N11432);
buf BUF1 (N24765, N24762);
or OR4 (N24766, N24746, N4470, N3536, N1333);
and AND3 (N24767, N24744, N7253, N8151);
not NOT1 (N24768, N24767);
buf BUF1 (N24769, N24761);
nor NOR2 (N24770, N24766, N8677);
nor NOR3 (N24771, N24748, N24728, N18252);
and AND4 (N24772, N24765, N6421, N9784, N3441);
nand NAND4 (N24773, N24763, N8582, N20841, N22941);
and AND2 (N24774, N24772, N14455);
not NOT1 (N24775, N24769);
buf BUF1 (N24776, N24770);
nand NAND2 (N24777, N24757, N18859);
nand NAND2 (N24778, N24764, N15007);
xor XOR2 (N24779, N24778, N18727);
and AND3 (N24780, N24776, N13777, N20573);
nand NAND2 (N24781, N24775, N5985);
xor XOR2 (N24782, N24745, N2599);
xor XOR2 (N24783, N24777, N3032);
and AND3 (N24784, N24771, N21169, N11655);
buf BUF1 (N24785, N24780);
not NOT1 (N24786, N24773);
nand NAND4 (N24787, N24786, N13957, N6584, N9852);
buf BUF1 (N24788, N24785);
nor NOR4 (N24789, N24788, N13814, N4282, N16205);
and AND3 (N24790, N24774, N21195, N8671);
or OR2 (N24791, N24787, N23945);
or OR2 (N24792, N24782, N9542);
or OR3 (N24793, N24789, N19279, N12738);
xor XOR2 (N24794, N24791, N18828);
nor NOR2 (N24795, N24783, N4570);
nand NAND2 (N24796, N24768, N808);
nor NOR2 (N24797, N24794, N14326);
xor XOR2 (N24798, N24795, N8123);
or OR4 (N24799, N24796, N8712, N12644, N21638);
buf BUF1 (N24800, N24792);
and AND3 (N24801, N24784, N19698, N5596);
buf BUF1 (N24802, N24760);
not NOT1 (N24803, N24802);
or OR2 (N24804, N24779, N3650);
and AND4 (N24805, N24800, N14032, N3358, N5154);
not NOT1 (N24806, N24790);
xor XOR2 (N24807, N24806, N23972);
and AND4 (N24808, N24807, N21180, N23608, N415);
buf BUF1 (N24809, N24797);
xor XOR2 (N24810, N24781, N956);
nand NAND2 (N24811, N24810, N7667);
not NOT1 (N24812, N24804);
nand NAND4 (N24813, N24798, N15708, N19362, N8754);
or OR4 (N24814, N24812, N7773, N10965, N24764);
buf BUF1 (N24815, N24799);
not NOT1 (N24816, N24813);
and AND4 (N24817, N24814, N22208, N3563, N2088);
xor XOR2 (N24818, N24816, N1438);
buf BUF1 (N24819, N24793);
and AND2 (N24820, N24808, N6277);
xor XOR2 (N24821, N24818, N9494);
and AND2 (N24822, N24805, N17668);
not NOT1 (N24823, N24822);
nand NAND4 (N24824, N24819, N22866, N24120, N24369);
xor XOR2 (N24825, N24821, N22214);
nor NOR2 (N24826, N24801, N18483);
and AND3 (N24827, N24820, N5979, N19854);
buf BUF1 (N24828, N24825);
or OR3 (N24829, N24827, N23875, N19645);
buf BUF1 (N24830, N24829);
nand NAND2 (N24831, N24828, N10691);
and AND4 (N24832, N24831, N148, N3822, N780);
buf BUF1 (N24833, N24809);
nor NOR2 (N24834, N24817, N22076);
buf BUF1 (N24835, N24833);
and AND4 (N24836, N24835, N12481, N3243, N3095);
xor XOR2 (N24837, N24811, N7853);
and AND3 (N24838, N24834, N12111, N5461);
xor XOR2 (N24839, N24823, N403);
or OR3 (N24840, N24838, N21055, N7277);
not NOT1 (N24841, N24824);
xor XOR2 (N24842, N24837, N6921);
nand NAND2 (N24843, N24842, N24831);
nor NOR2 (N24844, N24836, N10462);
nand NAND3 (N24845, N24841, N18775, N19106);
nor NOR4 (N24846, N24830, N19926, N16641, N2031);
and AND3 (N24847, N24815, N5144, N23984);
not NOT1 (N24848, N24846);
nand NAND3 (N24849, N24844, N6872, N24801);
not NOT1 (N24850, N24845);
xor XOR2 (N24851, N24847, N10523);
not NOT1 (N24852, N24839);
nand NAND4 (N24853, N24840, N638, N21266, N18430);
nor NOR3 (N24854, N24852, N15730, N17383);
and AND3 (N24855, N24803, N10098, N18805);
or OR3 (N24856, N24848, N21857, N6124);
nor NOR4 (N24857, N24853, N13667, N1957, N14319);
and AND3 (N24858, N24826, N8034, N5422);
xor XOR2 (N24859, N24850, N14319);
xor XOR2 (N24860, N24859, N14175);
nor NOR3 (N24861, N24849, N143, N23764);
not NOT1 (N24862, N24854);
nor NOR4 (N24863, N24857, N2187, N6058, N22652);
xor XOR2 (N24864, N24858, N11579);
or OR4 (N24865, N24855, N18061, N10998, N17151);
not NOT1 (N24866, N24851);
nand NAND2 (N24867, N24865, N397);
xor XOR2 (N24868, N24862, N2038);
or OR4 (N24869, N24868, N2636, N17992, N13760);
and AND4 (N24870, N24861, N3496, N14610, N19300);
or OR2 (N24871, N24843, N18306);
nor NOR3 (N24872, N24864, N21425, N12923);
buf BUF1 (N24873, N24860);
xor XOR2 (N24874, N24856, N12603);
xor XOR2 (N24875, N24832, N6603);
not NOT1 (N24876, N24870);
and AND4 (N24877, N24863, N12662, N3615, N10356);
xor XOR2 (N24878, N24874, N7832);
or OR4 (N24879, N24871, N18050, N1334, N17980);
and AND3 (N24880, N24869, N14099, N1808);
xor XOR2 (N24881, N24867, N15445);
or OR2 (N24882, N24866, N19368);
buf BUF1 (N24883, N24873);
and AND3 (N24884, N24878, N16430, N8534);
not NOT1 (N24885, N24884);
xor XOR2 (N24886, N24879, N24539);
not NOT1 (N24887, N24882);
nand NAND4 (N24888, N24883, N14396, N4758, N11701);
xor XOR2 (N24889, N24886, N641);
nand NAND3 (N24890, N24876, N3725, N17004);
and AND2 (N24891, N24880, N534);
buf BUF1 (N24892, N24890);
buf BUF1 (N24893, N24892);
nand NAND3 (N24894, N24887, N2140, N2874);
xor XOR2 (N24895, N24889, N13914);
buf BUF1 (N24896, N24885);
buf BUF1 (N24897, N24896);
buf BUF1 (N24898, N24891);
nor NOR4 (N24899, N24897, N9974, N9076, N12650);
not NOT1 (N24900, N24875);
xor XOR2 (N24901, N24894, N21262);
and AND4 (N24902, N24901, N24890, N2702, N14199);
xor XOR2 (N24903, N24899, N16193);
nor NOR3 (N24904, N24903, N5390, N2848);
or OR4 (N24905, N24888, N10725, N8189, N9433);
nand NAND2 (N24906, N24872, N3133);
buf BUF1 (N24907, N24895);
not NOT1 (N24908, N24877);
or OR4 (N24909, N24907, N3244, N24255, N1518);
nor NOR3 (N24910, N24908, N3057, N7816);
nor NOR2 (N24911, N24881, N5387);
xor XOR2 (N24912, N24902, N14542);
not NOT1 (N24913, N24910);
nor NOR2 (N24914, N24911, N24891);
and AND3 (N24915, N24905, N3949, N24370);
xor XOR2 (N24916, N24909, N5238);
and AND3 (N24917, N24904, N8417, N23760);
nand NAND2 (N24918, N24900, N21418);
nand NAND2 (N24919, N24918, N11256);
nor NOR3 (N24920, N24919, N21624, N9578);
nand NAND4 (N24921, N24912, N20877, N8052, N907);
nor NOR2 (N24922, N24921, N11910);
not NOT1 (N24923, N24906);
nor NOR2 (N24924, N24922, N20869);
buf BUF1 (N24925, N24916);
buf BUF1 (N24926, N24915);
nand NAND2 (N24927, N24923, N8371);
not NOT1 (N24928, N24926);
not NOT1 (N24929, N24927);
xor XOR2 (N24930, N24898, N21550);
and AND4 (N24931, N24913, N3068, N7228, N15283);
not NOT1 (N24932, N24930);
nand NAND3 (N24933, N24924, N23721, N10224);
xor XOR2 (N24934, N24928, N1292);
or OR3 (N24935, N24925, N24404, N4294);
and AND3 (N24936, N24929, N2405, N11016);
buf BUF1 (N24937, N24931);
buf BUF1 (N24938, N24935);
buf BUF1 (N24939, N24932);
xor XOR2 (N24940, N24893, N1674);
nor NOR2 (N24941, N24917, N623);
xor XOR2 (N24942, N24933, N4637);
xor XOR2 (N24943, N24942, N3430);
or OR2 (N24944, N24920, N121);
and AND3 (N24945, N24941, N4345, N14307);
xor XOR2 (N24946, N24943, N19196);
buf BUF1 (N24947, N24940);
and AND2 (N24948, N24945, N11337);
xor XOR2 (N24949, N24946, N12860);
xor XOR2 (N24950, N24937, N18281);
and AND4 (N24951, N24938, N21774, N22207, N14626);
buf BUF1 (N24952, N24914);
xor XOR2 (N24953, N24947, N2040);
or OR2 (N24954, N24953, N1864);
and AND3 (N24955, N24950, N11342, N14138);
and AND4 (N24956, N24939, N17632, N21165, N17504);
nor NOR3 (N24957, N24951, N13410, N12678);
or OR3 (N24958, N24957, N6447, N23435);
buf BUF1 (N24959, N24948);
xor XOR2 (N24960, N24956, N8553);
and AND4 (N24961, N24955, N818, N13679, N17769);
nand NAND3 (N24962, N24944, N2372, N22328);
buf BUF1 (N24963, N24934);
nand NAND4 (N24964, N24952, N17062, N17618, N8451);
nor NOR2 (N24965, N24959, N6206);
nor NOR4 (N24966, N24964, N126, N24825, N24361);
and AND2 (N24967, N24954, N15080);
nor NOR3 (N24968, N24967, N11936, N2763);
nand NAND4 (N24969, N24966, N18209, N16355, N5907);
nand NAND3 (N24970, N24961, N16436, N18963);
buf BUF1 (N24971, N24968);
xor XOR2 (N24972, N24969, N8027);
nand NAND4 (N24973, N24962, N1957, N2001, N18022);
or OR3 (N24974, N24965, N23940, N18538);
not NOT1 (N24975, N24949);
nor NOR4 (N24976, N24970, N12630, N13153, N12896);
xor XOR2 (N24977, N24936, N12839);
buf BUF1 (N24978, N24972);
buf BUF1 (N24979, N24974);
or OR3 (N24980, N24958, N21223, N5759);
nand NAND3 (N24981, N24977, N9669, N18034);
nor NOR4 (N24982, N24973, N17471, N1990, N12765);
nor NOR4 (N24983, N24980, N9752, N12973, N18535);
or OR3 (N24984, N24981, N23545, N18747);
not NOT1 (N24985, N24960);
buf BUF1 (N24986, N24982);
nand NAND3 (N24987, N24985, N22909, N16815);
nand NAND3 (N24988, N24979, N20950, N4414);
nor NOR3 (N24989, N24963, N1663, N3656);
nand NAND2 (N24990, N24984, N8682);
nor NOR3 (N24991, N24989, N24363, N20344);
nand NAND2 (N24992, N24988, N11263);
buf BUF1 (N24993, N24978);
not NOT1 (N24994, N24992);
buf BUF1 (N24995, N24991);
buf BUF1 (N24996, N24993);
nand NAND2 (N24997, N24987, N24950);
and AND3 (N24998, N24986, N18343, N16321);
and AND4 (N24999, N24990, N9105, N19388, N9950);
or OR2 (N25000, N24983, N23379);
not NOT1 (N25001, N24999);
and AND4 (N25002, N25000, N3963, N23846, N24715);
or OR4 (N25003, N24971, N8900, N19599, N18813);
buf BUF1 (N25004, N24994);
nor NOR4 (N25005, N24976, N9193, N20698, N4427);
nor NOR2 (N25006, N25003, N21463);
or OR4 (N25007, N24998, N9258, N8297, N14231);
xor XOR2 (N25008, N24975, N16670);
nand NAND3 (N25009, N25004, N11399, N13944);
not NOT1 (N25010, N24996);
buf BUF1 (N25011, N25002);
or OR4 (N25012, N25007, N19302, N16784, N15378);
buf BUF1 (N25013, N25012);
nand NAND4 (N25014, N25011, N24454, N24802, N15961);
not NOT1 (N25015, N25001);
or OR2 (N25016, N25013, N12327);
nand NAND2 (N25017, N25009, N19906);
nor NOR3 (N25018, N25010, N18415, N10731);
not NOT1 (N25019, N25008);
not NOT1 (N25020, N24995);
nor NOR2 (N25021, N25017, N14913);
nand NAND4 (N25022, N24997, N7778, N693, N10888);
nand NAND4 (N25023, N25015, N15837, N17258, N11630);
not NOT1 (N25024, N25014);
xor XOR2 (N25025, N25018, N1580);
and AND4 (N25026, N25025, N16734, N4243, N10154);
xor XOR2 (N25027, N25024, N12503);
or OR2 (N25028, N25021, N695);
nand NAND3 (N25029, N25020, N11971, N9830);
not NOT1 (N25030, N25023);
and AND2 (N25031, N25030, N19766);
xor XOR2 (N25032, N25028, N23965);
or OR4 (N25033, N25029, N15148, N15500, N5117);
buf BUF1 (N25034, N25019);
nand NAND3 (N25035, N25032, N5918, N24282);
xor XOR2 (N25036, N25016, N10096);
not NOT1 (N25037, N25035);
nand NAND4 (N25038, N25037, N13711, N20222, N17264);
nor NOR4 (N25039, N25034, N7357, N14868, N8143);
not NOT1 (N25040, N25036);
xor XOR2 (N25041, N25022, N23428);
and AND2 (N25042, N25005, N11008);
or OR3 (N25043, N25041, N20532, N22258);
nor NOR4 (N25044, N25033, N21856, N22747, N18810);
nand NAND3 (N25045, N25044, N5895, N2219);
or OR4 (N25046, N25038, N24874, N18517, N24009);
buf BUF1 (N25047, N25042);
and AND3 (N25048, N25039, N11900, N18918);
not NOT1 (N25049, N25046);
nand NAND2 (N25050, N25043, N896);
xor XOR2 (N25051, N25040, N4167);
nor NOR2 (N25052, N25049, N2977);
xor XOR2 (N25053, N25048, N16909);
and AND2 (N25054, N25031, N6702);
nor NOR2 (N25055, N25006, N17213);
not NOT1 (N25056, N25026);
nand NAND4 (N25057, N25055, N1737, N19, N19690);
and AND2 (N25058, N25054, N24153);
not NOT1 (N25059, N25056);
not NOT1 (N25060, N25053);
nand NAND2 (N25061, N25051, N23130);
not NOT1 (N25062, N25061);
and AND4 (N25063, N25045, N2196, N15032, N23839);
and AND2 (N25064, N25062, N12788);
xor XOR2 (N25065, N25064, N17958);
not NOT1 (N25066, N25065);
and AND3 (N25067, N25050, N18260, N11250);
xor XOR2 (N25068, N25058, N87);
nor NOR4 (N25069, N25059, N17509, N2128, N5538);
nor NOR4 (N25070, N25027, N22244, N1231, N8224);
or OR2 (N25071, N25047, N2445);
buf BUF1 (N25072, N25057);
nand NAND2 (N25073, N25052, N9636);
not NOT1 (N25074, N25073);
xor XOR2 (N25075, N25063, N20280);
not NOT1 (N25076, N25067);
nor NOR3 (N25077, N25069, N13454, N7875);
nor NOR3 (N25078, N25066, N11228, N21820);
nor NOR4 (N25079, N25070, N1893, N11458, N1342);
and AND2 (N25080, N25077, N6029);
nor NOR4 (N25081, N25080, N23180, N6168, N19331);
or OR4 (N25082, N25071, N2559, N2731, N23460);
or OR4 (N25083, N25078, N4314, N6797, N14725);
buf BUF1 (N25084, N25074);
nand NAND2 (N25085, N25081, N3221);
xor XOR2 (N25086, N25060, N23811);
nor NOR2 (N25087, N25083, N5679);
nor NOR4 (N25088, N25087, N7643, N17460, N6281);
nor NOR2 (N25089, N25079, N4172);
buf BUF1 (N25090, N25086);
nor NOR2 (N25091, N25089, N12385);
buf BUF1 (N25092, N25088);
nand NAND4 (N25093, N25084, N6536, N25061, N18544);
nor NOR3 (N25094, N25090, N7230, N527);
buf BUF1 (N25095, N25076);
xor XOR2 (N25096, N25093, N8922);
or OR2 (N25097, N25094, N23657);
not NOT1 (N25098, N25095);
nand NAND3 (N25099, N25075, N8520, N876);
nor NOR3 (N25100, N25092, N1320, N17486);
nand NAND2 (N25101, N25082, N13096);
or OR3 (N25102, N25100, N2449, N12704);
buf BUF1 (N25103, N25102);
buf BUF1 (N25104, N25098);
nor NOR2 (N25105, N25101, N9520);
or OR4 (N25106, N25099, N24710, N18305, N19436);
buf BUF1 (N25107, N25085);
and AND2 (N25108, N25107, N15524);
xor XOR2 (N25109, N25068, N6115);
nand NAND3 (N25110, N25091, N19180, N14932);
buf BUF1 (N25111, N25108);
or OR2 (N25112, N25109, N21869);
nor NOR3 (N25113, N25110, N9898, N5518);
not NOT1 (N25114, N25106);
xor XOR2 (N25115, N25111, N2877);
not NOT1 (N25116, N25096);
buf BUF1 (N25117, N25097);
buf BUF1 (N25118, N25114);
nand NAND3 (N25119, N25118, N12259, N2663);
nor NOR2 (N25120, N25117, N1843);
or OR3 (N25121, N25072, N6416, N23555);
nand NAND2 (N25122, N25104, N12051);
nand NAND2 (N25123, N25115, N1368);
buf BUF1 (N25124, N25121);
nand NAND3 (N25125, N25123, N20980, N2198);
xor XOR2 (N25126, N25112, N4625);
buf BUF1 (N25127, N25125);
or OR2 (N25128, N25113, N18108);
and AND4 (N25129, N25124, N18719, N244, N4419);
and AND4 (N25130, N25103, N3156, N13401, N16653);
xor XOR2 (N25131, N25119, N2443);
not NOT1 (N25132, N25105);
nor NOR2 (N25133, N25129, N9092);
and AND2 (N25134, N25130, N7777);
and AND4 (N25135, N25131, N18728, N22356, N18927);
nor NOR3 (N25136, N25127, N11032, N5910);
buf BUF1 (N25137, N25136);
buf BUF1 (N25138, N25134);
nor NOR3 (N25139, N25132, N25062, N19070);
nor NOR4 (N25140, N25116, N17859, N15815, N5410);
buf BUF1 (N25141, N25122);
nand NAND2 (N25142, N25120, N16402);
not NOT1 (N25143, N25141);
nor NOR4 (N25144, N25142, N12038, N3846, N9227);
and AND3 (N25145, N25126, N309, N15196);
nor NOR4 (N25146, N25140, N8773, N22335, N1795);
xor XOR2 (N25147, N25133, N19745);
or OR4 (N25148, N25145, N7165, N3706, N23269);
buf BUF1 (N25149, N25146);
nor NOR4 (N25150, N25137, N18856, N18402, N9709);
xor XOR2 (N25151, N25144, N5462);
nor NOR3 (N25152, N25139, N9068, N9161);
not NOT1 (N25153, N25128);
nand NAND3 (N25154, N25150, N8802, N3188);
xor XOR2 (N25155, N25148, N3315);
or OR2 (N25156, N25155, N13401);
not NOT1 (N25157, N25154);
nand NAND3 (N25158, N25138, N1960, N10580);
not NOT1 (N25159, N25143);
nand NAND2 (N25160, N25152, N3239);
buf BUF1 (N25161, N25153);
and AND3 (N25162, N25135, N11902, N21502);
not NOT1 (N25163, N25161);
or OR3 (N25164, N25156, N20445, N11419);
xor XOR2 (N25165, N25159, N16364);
not NOT1 (N25166, N25149);
and AND2 (N25167, N25158, N14042);
nand NAND4 (N25168, N25157, N18215, N1970, N25068);
buf BUF1 (N25169, N25164);
nand NAND3 (N25170, N25169, N8000, N19189);
buf BUF1 (N25171, N25165);
xor XOR2 (N25172, N25170, N2289);
and AND4 (N25173, N25151, N13220, N9389, N323);
nand NAND2 (N25174, N25167, N1411);
not NOT1 (N25175, N25172);
buf BUF1 (N25176, N25175);
buf BUF1 (N25177, N25160);
not NOT1 (N25178, N25166);
or OR2 (N25179, N25173, N7083);
nor NOR3 (N25180, N25174, N2527, N8304);
buf BUF1 (N25181, N25162);
nor NOR2 (N25182, N25179, N20961);
buf BUF1 (N25183, N25178);
xor XOR2 (N25184, N25177, N422);
xor XOR2 (N25185, N25168, N4560);
buf BUF1 (N25186, N25183);
nor NOR4 (N25187, N25185, N7954, N2819, N5517);
nand NAND3 (N25188, N25181, N7202, N17380);
buf BUF1 (N25189, N25176);
nand NAND4 (N25190, N25147, N18799, N7709, N24327);
and AND3 (N25191, N25187, N20792, N4097);
nor NOR4 (N25192, N25182, N13788, N11926, N9243);
buf BUF1 (N25193, N25190);
and AND3 (N25194, N25180, N4588, N22595);
not NOT1 (N25195, N25163);
and AND4 (N25196, N25194, N24803, N12672, N6298);
and AND4 (N25197, N25189, N5738, N7836, N3770);
nor NOR2 (N25198, N25184, N2790);
nand NAND4 (N25199, N25196, N4, N17481, N9511);
and AND4 (N25200, N25191, N1585, N10868, N5362);
not NOT1 (N25201, N25186);
and AND3 (N25202, N25197, N18398, N9767);
nand NAND2 (N25203, N25188, N7827);
nand NAND2 (N25204, N25203, N13607);
not NOT1 (N25205, N25171);
nand NAND3 (N25206, N25199, N13552, N24179);
and AND3 (N25207, N25192, N9936, N19284);
not NOT1 (N25208, N25202);
xor XOR2 (N25209, N25206, N20978);
and AND3 (N25210, N25200, N5532, N20930);
not NOT1 (N25211, N25198);
or OR4 (N25212, N25209, N16477, N18783, N19895);
xor XOR2 (N25213, N25195, N6812);
buf BUF1 (N25214, N25208);
and AND2 (N25215, N25214, N24512);
not NOT1 (N25216, N25193);
buf BUF1 (N25217, N25216);
nor NOR2 (N25218, N25213, N8878);
xor XOR2 (N25219, N25218, N13795);
not NOT1 (N25220, N25204);
or OR3 (N25221, N25210, N9571, N17238);
nor NOR2 (N25222, N25201, N15605);
or OR3 (N25223, N25217, N23222, N21829);
or OR4 (N25224, N25222, N5008, N11788, N3544);
and AND2 (N25225, N25215, N24831);
xor XOR2 (N25226, N25223, N13682);
nand NAND2 (N25227, N25220, N16251);
not NOT1 (N25228, N25211);
or OR4 (N25229, N25224, N10413, N21907, N7969);
and AND2 (N25230, N25212, N23210);
buf BUF1 (N25231, N25229);
nand NAND2 (N25232, N25221, N19280);
and AND3 (N25233, N25227, N23899, N6411);
nor NOR4 (N25234, N25230, N23820, N23119, N20484);
xor XOR2 (N25235, N25207, N17838);
buf BUF1 (N25236, N25228);
nor NOR3 (N25237, N25225, N4294, N18383);
or OR4 (N25238, N25219, N24850, N16138, N17552);
and AND2 (N25239, N25234, N2498);
nor NOR2 (N25240, N25236, N5648);
nor NOR4 (N25241, N25231, N23802, N22654, N5010);
nand NAND3 (N25242, N25239, N22095, N8204);
not NOT1 (N25243, N25237);
xor XOR2 (N25244, N25241, N1405);
not NOT1 (N25245, N25244);
xor XOR2 (N25246, N25232, N3243);
buf BUF1 (N25247, N25235);
or OR2 (N25248, N25242, N24224);
buf BUF1 (N25249, N25243);
buf BUF1 (N25250, N25248);
buf BUF1 (N25251, N25233);
not NOT1 (N25252, N25250);
not NOT1 (N25253, N25252);
nor NOR3 (N25254, N25247, N16668, N3872);
nor NOR3 (N25255, N25205, N13963, N25243);
nand NAND3 (N25256, N25255, N4767, N11397);
xor XOR2 (N25257, N25256, N15714);
nor NOR4 (N25258, N25249, N25229, N3839, N23816);
and AND3 (N25259, N25254, N17770, N13622);
and AND4 (N25260, N25240, N20759, N13127, N4951);
nor NOR4 (N25261, N25251, N24505, N6896, N16771);
not NOT1 (N25262, N25257);
nor NOR4 (N25263, N25262, N17479, N20843, N9052);
and AND4 (N25264, N25261, N4704, N21041, N14058);
and AND4 (N25265, N25260, N560, N10575, N8306);
nor NOR2 (N25266, N25238, N11962);
not NOT1 (N25267, N25263);
not NOT1 (N25268, N25253);
nand NAND2 (N25269, N25264, N645);
buf BUF1 (N25270, N25265);
or OR3 (N25271, N25266, N9202, N13500);
nand NAND3 (N25272, N25258, N4875, N24835);
not NOT1 (N25273, N25259);
or OR3 (N25274, N25271, N22887, N14435);
buf BUF1 (N25275, N25273);
not NOT1 (N25276, N25267);
nor NOR4 (N25277, N25272, N291, N1985, N15591);
and AND4 (N25278, N25226, N20432, N10284, N16581);
not NOT1 (N25279, N25278);
nand NAND2 (N25280, N25275, N7623);
nand NAND4 (N25281, N25280, N3398, N22994, N17498);
or OR2 (N25282, N25268, N1508);
buf BUF1 (N25283, N25270);
nand NAND2 (N25284, N25279, N14866);
nor NOR2 (N25285, N25277, N6424);
xor XOR2 (N25286, N25285, N19192);
not NOT1 (N25287, N25286);
nand NAND4 (N25288, N25276, N13053, N7706, N22248);
buf BUF1 (N25289, N25281);
nand NAND4 (N25290, N25282, N18982, N18215, N206);
buf BUF1 (N25291, N25284);
buf BUF1 (N25292, N25289);
or OR4 (N25293, N25291, N5152, N13203, N20235);
nand NAND2 (N25294, N25283, N7666);
and AND2 (N25295, N25274, N12952);
buf BUF1 (N25296, N25245);
xor XOR2 (N25297, N25294, N17947);
not NOT1 (N25298, N25293);
buf BUF1 (N25299, N25295);
nor NOR3 (N25300, N25288, N10540, N22559);
nand NAND4 (N25301, N25299, N24241, N13790, N2935);
nor NOR2 (N25302, N25300, N20322);
and AND4 (N25303, N25290, N12214, N16411, N9872);
xor XOR2 (N25304, N25296, N1309);
and AND3 (N25305, N25304, N21777, N11627);
buf BUF1 (N25306, N25302);
or OR2 (N25307, N25301, N25269);
not NOT1 (N25308, N17898);
nor NOR2 (N25309, N25307, N21974);
or OR4 (N25310, N25246, N18553, N12196, N17424);
buf BUF1 (N25311, N25308);
xor XOR2 (N25312, N25310, N20868);
and AND2 (N25313, N25303, N457);
and AND3 (N25314, N25311, N10033, N19809);
nand NAND4 (N25315, N25287, N14172, N16291, N20877);
or OR3 (N25316, N25297, N21142, N21574);
nand NAND2 (N25317, N25305, N10607);
or OR3 (N25318, N25306, N9986, N7493);
not NOT1 (N25319, N25292);
not NOT1 (N25320, N25319);
xor XOR2 (N25321, N25315, N15578);
and AND2 (N25322, N25314, N4156);
or OR3 (N25323, N25309, N16374, N16680);
not NOT1 (N25324, N25321);
nor NOR3 (N25325, N25317, N142, N20052);
nand NAND4 (N25326, N25323, N23080, N24792, N8510);
and AND2 (N25327, N25320, N9997);
buf BUF1 (N25328, N25324);
or OR2 (N25329, N25325, N22144);
nand NAND3 (N25330, N25318, N570, N10375);
nor NOR4 (N25331, N25312, N1267, N18712, N2581);
nor NOR3 (N25332, N25330, N738, N21982);
and AND3 (N25333, N25322, N10193, N19276);
nor NOR3 (N25334, N25333, N24011, N6681);
not NOT1 (N25335, N25332);
nand NAND2 (N25336, N25327, N7200);
nand NAND4 (N25337, N25334, N20113, N22958, N3292);
not NOT1 (N25338, N25337);
and AND2 (N25339, N25336, N13668);
not NOT1 (N25340, N25316);
not NOT1 (N25341, N25339);
nor NOR4 (N25342, N25340, N18636, N11172, N20786);
buf BUF1 (N25343, N25329);
or OR4 (N25344, N25335, N14657, N8560, N5066);
buf BUF1 (N25345, N25343);
and AND3 (N25346, N25345, N10300, N11372);
nor NOR3 (N25347, N25344, N5047, N11553);
or OR3 (N25348, N25326, N14541, N15734);
not NOT1 (N25349, N25338);
nand NAND2 (N25350, N25313, N14484);
and AND2 (N25351, N25348, N20433);
buf BUF1 (N25352, N25350);
and AND3 (N25353, N25328, N19550, N7722);
not NOT1 (N25354, N25352);
nor NOR3 (N25355, N25346, N21548, N2300);
buf BUF1 (N25356, N25355);
xor XOR2 (N25357, N25354, N2237);
buf BUF1 (N25358, N25331);
nor NOR3 (N25359, N25349, N2262, N18313);
nor NOR3 (N25360, N25359, N23035, N15319);
nand NAND4 (N25361, N25351, N8673, N7712, N4212);
not NOT1 (N25362, N25357);
or OR2 (N25363, N25353, N18478);
not NOT1 (N25364, N25358);
nor NOR3 (N25365, N25361, N15772, N24253);
not NOT1 (N25366, N25360);
buf BUF1 (N25367, N25342);
buf BUF1 (N25368, N25366);
not NOT1 (N25369, N25363);
buf BUF1 (N25370, N25298);
buf BUF1 (N25371, N25364);
nor NOR4 (N25372, N25362, N14828, N4331, N7225);
buf BUF1 (N25373, N25365);
nand NAND3 (N25374, N25371, N4469, N19255);
nor NOR4 (N25375, N25347, N1857, N6687, N18205);
and AND2 (N25376, N25356, N7954);
not NOT1 (N25377, N25376);
or OR2 (N25378, N25341, N9122);
or OR2 (N25379, N25378, N24355);
xor XOR2 (N25380, N25377, N25355);
nand NAND3 (N25381, N25370, N8331, N7145);
nand NAND3 (N25382, N25381, N2385, N7941);
not NOT1 (N25383, N25368);
xor XOR2 (N25384, N25373, N14751);
and AND3 (N25385, N25374, N2289, N4836);
buf BUF1 (N25386, N25369);
not NOT1 (N25387, N25382);
xor XOR2 (N25388, N25386, N6075);
and AND3 (N25389, N25385, N22085, N13308);
or OR3 (N25390, N25389, N21130, N7818);
buf BUF1 (N25391, N25379);
nor NOR3 (N25392, N25391, N21981, N1048);
and AND3 (N25393, N25372, N16062, N823);
and AND2 (N25394, N25388, N1315);
not NOT1 (N25395, N25367);
and AND4 (N25396, N25393, N13154, N13150, N9581);
buf BUF1 (N25397, N25394);
buf BUF1 (N25398, N25387);
and AND4 (N25399, N25397, N18804, N21318, N15952);
not NOT1 (N25400, N25399);
xor XOR2 (N25401, N25400, N23844);
xor XOR2 (N25402, N25390, N21551);
buf BUF1 (N25403, N25402);
xor XOR2 (N25404, N25392, N20347);
and AND2 (N25405, N25395, N12333);
nand NAND3 (N25406, N25401, N14422, N3412);
xor XOR2 (N25407, N25380, N7570);
xor XOR2 (N25408, N25383, N18282);
buf BUF1 (N25409, N25404);
nand NAND3 (N25410, N25384, N14335, N21314);
or OR2 (N25411, N25408, N9340);
not NOT1 (N25412, N25405);
nor NOR4 (N25413, N25411, N21165, N10841, N3048);
nor NOR4 (N25414, N25409, N14925, N5961, N14919);
xor XOR2 (N25415, N25407, N20629);
xor XOR2 (N25416, N25396, N9124);
not NOT1 (N25417, N25410);
nand NAND4 (N25418, N25403, N18335, N19046, N4630);
xor XOR2 (N25419, N25406, N10657);
not NOT1 (N25420, N25414);
buf BUF1 (N25421, N25375);
or OR3 (N25422, N25419, N10066, N19629);
or OR2 (N25423, N25416, N20954);
and AND3 (N25424, N25422, N11110, N833);
and AND4 (N25425, N25415, N9112, N294, N18933);
xor XOR2 (N25426, N25417, N20096);
not NOT1 (N25427, N25413);
or OR4 (N25428, N25420, N12277, N1659, N148);
nor NOR3 (N25429, N25426, N23523, N25275);
nor NOR2 (N25430, N25425, N1356);
nand NAND2 (N25431, N25412, N20711);
nor NOR4 (N25432, N25421, N7374, N19090, N10427);
not NOT1 (N25433, N25432);
buf BUF1 (N25434, N25424);
and AND2 (N25435, N25431, N5867);
xor XOR2 (N25436, N25428, N1564);
or OR2 (N25437, N25436, N18626);
not NOT1 (N25438, N25435);
buf BUF1 (N25439, N25418);
buf BUF1 (N25440, N25427);
not NOT1 (N25441, N25434);
or OR2 (N25442, N25438, N19297);
or OR2 (N25443, N25437, N4998);
not NOT1 (N25444, N25442);
xor XOR2 (N25445, N25439, N21318);
xor XOR2 (N25446, N25429, N18243);
buf BUF1 (N25447, N25430);
or OR2 (N25448, N25398, N24556);
xor XOR2 (N25449, N25433, N13117);
and AND2 (N25450, N25423, N18294);
nor NOR3 (N25451, N25448, N9690, N19050);
nand NAND4 (N25452, N25450, N3000, N15279, N558);
buf BUF1 (N25453, N25444);
and AND4 (N25454, N25440, N21791, N10009, N19817);
buf BUF1 (N25455, N25445);
nand NAND4 (N25456, N25453, N3741, N6563, N15554);
or OR3 (N25457, N25449, N4365, N20711);
and AND4 (N25458, N25447, N1111, N1316, N18318);
nor NOR2 (N25459, N25446, N20819);
buf BUF1 (N25460, N25451);
nand NAND3 (N25461, N25457, N13357, N12787);
and AND2 (N25462, N25460, N1655);
nor NOR2 (N25463, N25455, N18789);
nor NOR2 (N25464, N25443, N21855);
nand NAND4 (N25465, N25462, N20494, N22431, N4218);
nand NAND4 (N25466, N25459, N25092, N12809, N7544);
nor NOR3 (N25467, N25441, N19038, N13862);
nand NAND2 (N25468, N25456, N19306);
nand NAND4 (N25469, N25465, N5183, N8719, N11279);
xor XOR2 (N25470, N25469, N5259);
and AND3 (N25471, N25463, N14395, N1642);
xor XOR2 (N25472, N25468, N11743);
not NOT1 (N25473, N25461);
nand NAND4 (N25474, N25467, N5721, N13208, N24607);
not NOT1 (N25475, N25474);
and AND4 (N25476, N25472, N21187, N9765, N12245);
not NOT1 (N25477, N25470);
buf BUF1 (N25478, N25452);
or OR4 (N25479, N25471, N7838, N15961, N24606);
and AND3 (N25480, N25458, N12805, N23172);
not NOT1 (N25481, N25479);
not NOT1 (N25482, N25481);
buf BUF1 (N25483, N25476);
not NOT1 (N25484, N25477);
buf BUF1 (N25485, N25464);
nor NOR4 (N25486, N25466, N12445, N24789, N22150);
not NOT1 (N25487, N25480);
xor XOR2 (N25488, N25482, N17145);
and AND4 (N25489, N25475, N23618, N21308, N833);
and AND2 (N25490, N25473, N19700);
xor XOR2 (N25491, N25454, N9109);
nand NAND3 (N25492, N25489, N5204, N13105);
buf BUF1 (N25493, N25488);
nor NOR2 (N25494, N25485, N8988);
and AND4 (N25495, N25493, N18477, N15515, N5833);
nand NAND3 (N25496, N25484, N13766, N17364);
nand NAND3 (N25497, N25491, N18659, N4199);
and AND2 (N25498, N25497, N25432);
and AND2 (N25499, N25494, N8194);
xor XOR2 (N25500, N25495, N10576);
nand NAND4 (N25501, N25496, N4779, N7723, N22346);
or OR2 (N25502, N25492, N13976);
buf BUF1 (N25503, N25490);
or OR4 (N25504, N25487, N16821, N15326, N23869);
nor NOR4 (N25505, N25500, N23383, N9408, N1931);
nor NOR4 (N25506, N25502, N15202, N5514, N8326);
not NOT1 (N25507, N25499);
xor XOR2 (N25508, N25498, N9269);
and AND4 (N25509, N25478, N14919, N22062, N14823);
nor NOR4 (N25510, N25483, N2155, N3445, N22888);
nand NAND2 (N25511, N25510, N24021);
and AND4 (N25512, N25505, N4264, N8228, N21480);
buf BUF1 (N25513, N25501);
nand NAND2 (N25514, N25507, N12941);
buf BUF1 (N25515, N25512);
buf BUF1 (N25516, N25509);
nand NAND3 (N25517, N25516, N10447, N12161);
buf BUF1 (N25518, N25511);
nand NAND4 (N25519, N25515, N2897, N9644, N12135);
nor NOR3 (N25520, N25514, N2669, N16133);
xor XOR2 (N25521, N25486, N5709);
xor XOR2 (N25522, N25503, N22);
nand NAND3 (N25523, N25522, N2676, N15243);
nor NOR4 (N25524, N25518, N24623, N19194, N9069);
not NOT1 (N25525, N25513);
and AND3 (N25526, N25519, N2656, N25494);
and AND2 (N25527, N25524, N3990);
nor NOR4 (N25528, N25520, N14124, N2826, N9817);
or OR4 (N25529, N25504, N23967, N4342, N18283);
or OR4 (N25530, N25521, N24241, N22726, N707);
not NOT1 (N25531, N25523);
buf BUF1 (N25532, N25506);
and AND4 (N25533, N25532, N21886, N12611, N5149);
buf BUF1 (N25534, N25529);
or OR3 (N25535, N25534, N25419, N21119);
not NOT1 (N25536, N25533);
xor XOR2 (N25537, N25530, N21177);
nand NAND4 (N25538, N25525, N14823, N19672, N25117);
nor NOR4 (N25539, N25528, N16420, N12747, N4551);
and AND2 (N25540, N25508, N2021);
nor NOR4 (N25541, N25540, N14251, N14001, N6556);
or OR2 (N25542, N25535, N21116);
and AND2 (N25543, N25542, N24126);
or OR2 (N25544, N25527, N23845);
xor XOR2 (N25545, N25541, N2186);
or OR2 (N25546, N25536, N13148);
not NOT1 (N25547, N25539);
nor NOR3 (N25548, N25546, N22142, N24037);
xor XOR2 (N25549, N25537, N8369);
nand NAND3 (N25550, N25517, N13477, N8774);
or OR2 (N25551, N25538, N5618);
not NOT1 (N25552, N25543);
or OR3 (N25553, N25531, N20762, N8766);
not NOT1 (N25554, N25549);
not NOT1 (N25555, N25544);
buf BUF1 (N25556, N25548);
nor NOR2 (N25557, N25545, N17216);
not NOT1 (N25558, N25551);
buf BUF1 (N25559, N25547);
or OR3 (N25560, N25550, N7064, N16403);
and AND4 (N25561, N25526, N19151, N10575, N173);
and AND4 (N25562, N25556, N1470, N6039, N10479);
buf BUF1 (N25563, N25562);
nand NAND2 (N25564, N25560, N23420);
buf BUF1 (N25565, N25564);
or OR2 (N25566, N25559, N83);
nand NAND3 (N25567, N25566, N7520, N738);
xor XOR2 (N25568, N25565, N16918);
not NOT1 (N25569, N25563);
buf BUF1 (N25570, N25568);
buf BUF1 (N25571, N25554);
nand NAND3 (N25572, N25561, N24211, N10257);
nor NOR3 (N25573, N25572, N375, N9041);
nor NOR4 (N25574, N25555, N12760, N5271, N19167);
nand NAND3 (N25575, N25571, N20419, N1017);
buf BUF1 (N25576, N25569);
and AND4 (N25577, N25567, N25152, N19021, N16310);
nand NAND2 (N25578, N25576, N14890);
buf BUF1 (N25579, N25575);
and AND3 (N25580, N25553, N4221, N19503);
and AND2 (N25581, N25558, N10820);
xor XOR2 (N25582, N25580, N23968);
nand NAND3 (N25583, N25552, N14397, N5557);
xor XOR2 (N25584, N25557, N18457);
not NOT1 (N25585, N25577);
and AND3 (N25586, N25584, N884, N19372);
not NOT1 (N25587, N25585);
or OR2 (N25588, N25581, N18055);
xor XOR2 (N25589, N25582, N14536);
or OR2 (N25590, N25586, N7074);
xor XOR2 (N25591, N25579, N21356);
nor NOR3 (N25592, N25588, N15466, N10013);
not NOT1 (N25593, N25570);
not NOT1 (N25594, N25592);
buf BUF1 (N25595, N25583);
and AND2 (N25596, N25574, N7751);
buf BUF1 (N25597, N25573);
and AND2 (N25598, N25596, N19369);
xor XOR2 (N25599, N25597, N8381);
nor NOR3 (N25600, N25590, N5136, N17899);
nor NOR3 (N25601, N25599, N11648, N12209);
buf BUF1 (N25602, N25578);
nor NOR2 (N25603, N25598, N9549);
nand NAND4 (N25604, N25587, N21277, N25368, N22771);
xor XOR2 (N25605, N25603, N1595);
and AND4 (N25606, N25593, N18352, N15584, N7015);
nor NOR4 (N25607, N25604, N3425, N2501, N18761);
or OR4 (N25608, N25595, N24023, N1683, N15485);
nor NOR4 (N25609, N25608, N25062, N16426, N18336);
or OR3 (N25610, N25591, N17808, N5736);
buf BUF1 (N25611, N25601);
nand NAND2 (N25612, N25600, N4394);
not NOT1 (N25613, N25609);
buf BUF1 (N25614, N25594);
and AND2 (N25615, N25605, N21031);
xor XOR2 (N25616, N25606, N7453);
endmodule