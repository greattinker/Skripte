// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23;

output N2006,N2019,N2017,N2012,N1998,N2018,N2021,N2020,N2008,N2023;

nor NOR2 (N24, N22, N8);
buf BUF1 (N25, N13);
buf BUF1 (N26, N4);
nor NOR2 (N27, N22, N26);
buf BUF1 (N28, N22);
nor NOR4 (N29, N11, N28, N9, N3);
xor XOR2 (N30, N17, N20);
not NOT1 (N31, N17);
nand NAND4 (N32, N9, N9, N10, N30);
and AND2 (N33, N3, N2);
not NOT1 (N34, N9);
nor NOR4 (N35, N6, N34, N15, N2);
not NOT1 (N36, N23);
and AND4 (N37, N31, N24, N12, N32);
nand NAND4 (N38, N33, N4, N28, N24);
nand NAND4 (N39, N28, N32, N12, N14);
nand NAND2 (N40, N26, N23);
xor XOR2 (N41, N30, N11);
nor NOR4 (N42, N29, N33, N30, N30);
or OR3 (N43, N27, N32, N22);
and AND4 (N44, N37, N2, N40, N1);
buf BUF1 (N45, N40);
nor NOR2 (N46, N39, N14);
not NOT1 (N47, N25);
nand NAND3 (N48, N46, N37, N31);
nand NAND4 (N49, N41, N37, N19, N44);
or OR4 (N50, N20, N15, N19, N27);
nor NOR4 (N51, N45, N7, N17, N3);
buf BUF1 (N52, N49);
not NOT1 (N53, N35);
buf BUF1 (N54, N50);
nand NAND2 (N55, N51, N1);
nand NAND4 (N56, N55, N51, N2, N40);
xor XOR2 (N57, N54, N45);
not NOT1 (N58, N48);
not NOT1 (N59, N38);
and AND4 (N60, N57, N38, N50, N40);
xor XOR2 (N61, N58, N58);
nand NAND2 (N62, N59, N8);
and AND4 (N63, N47, N24, N56, N43);
nor NOR3 (N64, N54, N56, N37);
buf BUF1 (N65, N8);
or OR4 (N66, N61, N12, N42, N42);
and AND4 (N67, N57, N65, N45, N38);
not NOT1 (N68, N14);
and AND4 (N69, N68, N6, N50, N30);
buf BUF1 (N70, N36);
not NOT1 (N71, N66);
buf BUF1 (N72, N67);
buf BUF1 (N73, N62);
nand NAND3 (N74, N52, N29, N23);
buf BUF1 (N75, N72);
nand NAND2 (N76, N64, N7);
not NOT1 (N77, N63);
nand NAND2 (N78, N53, N12);
buf BUF1 (N79, N76);
or OR3 (N80, N79, N10, N26);
or OR3 (N81, N70, N45, N63);
buf BUF1 (N82, N60);
not NOT1 (N83, N74);
or OR2 (N84, N82, N50);
xor XOR2 (N85, N80, N72);
not NOT1 (N86, N77);
buf BUF1 (N87, N71);
nor NOR4 (N88, N85, N4, N7, N3);
not NOT1 (N89, N88);
buf BUF1 (N90, N87);
or OR3 (N91, N89, N73, N14);
nand NAND2 (N92, N18, N63);
nand NAND3 (N93, N81, N51, N79);
nand NAND2 (N94, N93, N28);
nand NAND2 (N95, N91, N63);
or OR4 (N96, N83, N90, N26, N32);
and AND2 (N97, N28, N33);
not NOT1 (N98, N69);
and AND2 (N99, N95, N37);
or OR3 (N100, N99, N35, N83);
nor NOR4 (N101, N94, N70, N82, N62);
nand NAND2 (N102, N75, N37);
and AND2 (N103, N86, N86);
buf BUF1 (N104, N101);
not NOT1 (N105, N103);
nand NAND4 (N106, N98, N54, N94, N31);
not NOT1 (N107, N100);
xor XOR2 (N108, N106, N73);
and AND2 (N109, N97, N100);
xor XOR2 (N110, N78, N42);
buf BUF1 (N111, N92);
not NOT1 (N112, N105);
nor NOR3 (N113, N109, N24, N82);
nand NAND4 (N114, N107, N98, N87, N105);
nand NAND4 (N115, N113, N75, N81, N2);
buf BUF1 (N116, N108);
buf BUF1 (N117, N102);
not NOT1 (N118, N117);
not NOT1 (N119, N112);
xor XOR2 (N120, N84, N64);
buf BUF1 (N121, N111);
nor NOR3 (N122, N121, N49, N83);
and AND4 (N123, N119, N86, N10, N59);
buf BUF1 (N124, N104);
nor NOR3 (N125, N96, N113, N67);
nor NOR4 (N126, N118, N46, N100, N18);
buf BUF1 (N127, N116);
or OR2 (N128, N123, N71);
or OR2 (N129, N126, N66);
nand NAND3 (N130, N122, N94, N119);
buf BUF1 (N131, N124);
and AND3 (N132, N125, N31, N44);
xor XOR2 (N133, N129, N3);
nor NOR3 (N134, N127, N6, N2);
or OR3 (N135, N130, N67, N35);
xor XOR2 (N136, N131, N56);
buf BUF1 (N137, N115);
or OR3 (N138, N110, N66, N87);
nor NOR2 (N139, N136, N50);
or OR3 (N140, N138, N21, N22);
or OR3 (N141, N140, N99, N12);
or OR3 (N142, N133, N36, N123);
or OR3 (N143, N139, N3, N50);
not NOT1 (N144, N137);
nor NOR2 (N145, N142, N42);
xor XOR2 (N146, N144, N30);
or OR4 (N147, N120, N37, N96, N27);
nand NAND4 (N148, N147, N11, N78, N43);
nand NAND3 (N149, N145, N138, N80);
not NOT1 (N150, N141);
nor NOR2 (N151, N132, N79);
and AND3 (N152, N146, N99, N118);
not NOT1 (N153, N148);
xor XOR2 (N154, N114, N87);
xor XOR2 (N155, N143, N92);
nor NOR3 (N156, N128, N73, N90);
or OR4 (N157, N149, N7, N79, N129);
buf BUF1 (N158, N152);
or OR4 (N159, N155, N136, N107, N118);
nand NAND3 (N160, N151, N19, N37);
xor XOR2 (N161, N159, N121);
xor XOR2 (N162, N135, N56);
nand NAND4 (N163, N162, N36, N16, N95);
buf BUF1 (N164, N161);
not NOT1 (N165, N156);
buf BUF1 (N166, N165);
nor NOR2 (N167, N164, N138);
not NOT1 (N168, N167);
and AND2 (N169, N157, N64);
and AND3 (N170, N134, N72, N154);
nor NOR2 (N171, N25, N138);
and AND3 (N172, N163, N131, N127);
and AND2 (N173, N160, N25);
not NOT1 (N174, N173);
nor NOR2 (N175, N174, N20);
nand NAND2 (N176, N153, N153);
nor NOR2 (N177, N166, N8);
and AND4 (N178, N175, N9, N98, N74);
buf BUF1 (N179, N171);
not NOT1 (N180, N172);
nor NOR2 (N181, N180, N174);
nand NAND3 (N182, N150, N60, N61);
nand NAND2 (N183, N158, N137);
buf BUF1 (N184, N170);
buf BUF1 (N185, N169);
and AND2 (N186, N183, N45);
nor NOR4 (N187, N177, N14, N70, N117);
not NOT1 (N188, N182);
xor XOR2 (N189, N188, N55);
nand NAND2 (N190, N179, N103);
buf BUF1 (N191, N181);
nand NAND2 (N192, N191, N175);
xor XOR2 (N193, N184, N56);
nand NAND3 (N194, N178, N159, N169);
or OR4 (N195, N190, N106, N126, N35);
or OR3 (N196, N187, N109, N116);
nand NAND3 (N197, N168, N121, N160);
nor NOR3 (N198, N192, N20, N28);
xor XOR2 (N199, N185, N145);
or OR3 (N200, N194, N121, N31);
buf BUF1 (N201, N189);
xor XOR2 (N202, N186, N155);
xor XOR2 (N203, N176, N145);
or OR3 (N204, N200, N186, N27);
or OR2 (N205, N203, N31);
nor NOR3 (N206, N195, N3, N76);
not NOT1 (N207, N199);
buf BUF1 (N208, N201);
and AND2 (N209, N207, N169);
nand NAND4 (N210, N209, N48, N25, N161);
buf BUF1 (N211, N197);
xor XOR2 (N212, N206, N59);
or OR3 (N213, N204, N164, N136);
nand NAND3 (N214, N211, N27, N107);
nor NOR3 (N215, N205, N152, N118);
nor NOR3 (N216, N198, N80, N203);
nand NAND2 (N217, N210, N9);
and AND4 (N218, N215, N33, N192, N160);
nor NOR4 (N219, N217, N45, N143, N128);
not NOT1 (N220, N219);
nor NOR3 (N221, N213, N114, N70);
not NOT1 (N222, N202);
or OR2 (N223, N196, N4);
not NOT1 (N224, N222);
nand NAND4 (N225, N218, N224, N197, N30);
not NOT1 (N226, N70);
buf BUF1 (N227, N208);
nand NAND3 (N228, N216, N80, N121);
or OR2 (N229, N220, N114);
buf BUF1 (N230, N228);
nand NAND2 (N231, N226, N153);
or OR2 (N232, N225, N168);
or OR4 (N233, N212, N3, N152, N110);
not NOT1 (N234, N231);
not NOT1 (N235, N214);
or OR2 (N236, N227, N233);
xor XOR2 (N237, N39, N7);
xor XOR2 (N238, N235, N209);
buf BUF1 (N239, N229);
nand NAND3 (N240, N236, N96, N114);
nor NOR3 (N241, N237, N174, N218);
nand NAND2 (N242, N232, N148);
and AND2 (N243, N240, N92);
or OR2 (N244, N238, N192);
nand NAND4 (N245, N244, N23, N128, N100);
and AND4 (N246, N242, N23, N95, N218);
or OR2 (N247, N223, N177);
not NOT1 (N248, N241);
nor NOR3 (N249, N243, N234, N150);
buf BUF1 (N250, N20);
not NOT1 (N251, N250);
and AND3 (N252, N247, N156, N29);
not NOT1 (N253, N251);
not NOT1 (N254, N193);
xor XOR2 (N255, N239, N72);
xor XOR2 (N256, N249, N29);
or OR3 (N257, N256, N134, N227);
xor XOR2 (N258, N246, N171);
nand NAND3 (N259, N258, N58, N193);
xor XOR2 (N260, N248, N225);
buf BUF1 (N261, N253);
or OR3 (N262, N261, N115, N215);
buf BUF1 (N263, N257);
buf BUF1 (N264, N230);
buf BUF1 (N265, N260);
not NOT1 (N266, N265);
buf BUF1 (N267, N221);
xor XOR2 (N268, N245, N72);
nand NAND3 (N269, N259, N65, N81);
buf BUF1 (N270, N268);
xor XOR2 (N271, N262, N168);
not NOT1 (N272, N271);
and AND4 (N273, N269, N57, N209, N5);
buf BUF1 (N274, N272);
xor XOR2 (N275, N270, N53);
buf BUF1 (N276, N263);
or OR2 (N277, N255, N179);
nand NAND3 (N278, N274, N99, N151);
and AND4 (N279, N252, N69, N133, N201);
and AND4 (N280, N277, N63, N82, N26);
nor NOR4 (N281, N264, N234, N236, N195);
buf BUF1 (N282, N280);
nor NOR2 (N283, N267, N85);
buf BUF1 (N284, N282);
and AND2 (N285, N279, N59);
nand NAND3 (N286, N273, N172, N145);
buf BUF1 (N287, N266);
and AND2 (N288, N283, N51);
or OR2 (N289, N288, N193);
nand NAND2 (N290, N276, N187);
xor XOR2 (N291, N254, N290);
buf BUF1 (N292, N42);
buf BUF1 (N293, N284);
nor NOR4 (N294, N281, N88, N264, N132);
not NOT1 (N295, N286);
nor NOR2 (N296, N278, N150);
and AND2 (N297, N285, N267);
xor XOR2 (N298, N275, N56);
nor NOR4 (N299, N297, N225, N245, N150);
xor XOR2 (N300, N295, N88);
and AND4 (N301, N289, N91, N30, N294);
xor XOR2 (N302, N228, N50);
not NOT1 (N303, N293);
or OR3 (N304, N299, N296, N37);
xor XOR2 (N305, N207, N245);
nand NAND3 (N306, N305, N226, N265);
or OR4 (N307, N287, N15, N75, N182);
xor XOR2 (N308, N302, N77);
buf BUF1 (N309, N304);
nand NAND2 (N310, N308, N70);
not NOT1 (N311, N310);
buf BUF1 (N312, N306);
nor NOR4 (N313, N307, N312, N95, N76);
not NOT1 (N314, N280);
or OR3 (N315, N298, N171, N215);
not NOT1 (N316, N291);
buf BUF1 (N317, N300);
and AND4 (N318, N303, N241, N60, N74);
xor XOR2 (N319, N315, N273);
nand NAND3 (N320, N309, N200, N68);
nor NOR4 (N321, N311, N56, N121, N314);
nor NOR4 (N322, N189, N249, N28, N9);
and AND2 (N323, N319, N290);
or OR4 (N324, N322, N231, N169, N10);
not NOT1 (N325, N301);
nand NAND4 (N326, N320, N14, N304, N49);
buf BUF1 (N327, N323);
not NOT1 (N328, N325);
and AND4 (N329, N321, N33, N88, N105);
buf BUF1 (N330, N324);
or OR2 (N331, N326, N36);
not NOT1 (N332, N331);
not NOT1 (N333, N317);
nor NOR4 (N334, N292, N261, N58, N85);
xor XOR2 (N335, N328, N150);
or OR4 (N336, N313, N314, N39, N268);
and AND2 (N337, N318, N254);
and AND3 (N338, N335, N222, N253);
nor NOR2 (N339, N330, N315);
or OR2 (N340, N316, N287);
and AND2 (N341, N340, N335);
or OR2 (N342, N337, N235);
and AND2 (N343, N342, N77);
buf BUF1 (N344, N338);
xor XOR2 (N345, N339, N337);
nand NAND2 (N346, N336, N118);
or OR3 (N347, N329, N30, N193);
nor NOR4 (N348, N344, N21, N226, N331);
nor NOR3 (N349, N333, N163, N48);
or OR3 (N350, N341, N112, N347);
or OR3 (N351, N187, N156, N305);
not NOT1 (N352, N349);
xor XOR2 (N353, N332, N328);
not NOT1 (N354, N348);
buf BUF1 (N355, N346);
nor NOR4 (N356, N351, N149, N259, N335);
and AND3 (N357, N350, N128, N159);
buf BUF1 (N358, N357);
and AND3 (N359, N352, N36, N121);
buf BUF1 (N360, N353);
not NOT1 (N361, N360);
nand NAND3 (N362, N359, N63, N208);
nand NAND2 (N363, N355, N184);
nand NAND4 (N364, N362, N355, N175, N276);
or OR4 (N365, N364, N12, N229, N41);
xor XOR2 (N366, N345, N164);
nand NAND2 (N367, N354, N145);
not NOT1 (N368, N356);
or OR4 (N369, N334, N77, N315, N105);
not NOT1 (N370, N366);
buf BUF1 (N371, N343);
and AND2 (N372, N371, N100);
nor NOR4 (N373, N361, N43, N369, N88);
nor NOR3 (N374, N148, N239, N336);
nand NAND4 (N375, N358, N266, N24, N220);
not NOT1 (N376, N375);
and AND3 (N377, N372, N374, N318);
not NOT1 (N378, N6);
buf BUF1 (N379, N377);
buf BUF1 (N380, N376);
nand NAND3 (N381, N370, N87, N321);
and AND3 (N382, N378, N168, N155);
nor NOR2 (N383, N365, N110);
not NOT1 (N384, N381);
buf BUF1 (N385, N367);
not NOT1 (N386, N385);
xor XOR2 (N387, N379, N164);
not NOT1 (N388, N363);
buf BUF1 (N389, N373);
and AND4 (N390, N383, N346, N327, N142);
nor NOR3 (N391, N249, N16, N88);
and AND4 (N392, N390, N222, N241, N121);
not NOT1 (N393, N386);
nor NOR4 (N394, N384, N50, N326, N364);
nand NAND3 (N395, N388, N114, N392);
buf BUF1 (N396, N23);
not NOT1 (N397, N394);
nor NOR3 (N398, N382, N346, N219);
not NOT1 (N399, N393);
not NOT1 (N400, N391);
not NOT1 (N401, N389);
nor NOR2 (N402, N397, N194);
buf BUF1 (N403, N400);
nand NAND3 (N404, N398, N403, N286);
not NOT1 (N405, N378);
nand NAND3 (N406, N368, N51, N256);
xor XOR2 (N407, N401, N180);
nand NAND4 (N408, N402, N236, N348, N148);
xor XOR2 (N409, N405, N265);
or OR3 (N410, N407, N344, N368);
and AND2 (N411, N408, N201);
nor NOR2 (N412, N409, N338);
or OR3 (N413, N411, N257, N371);
and AND4 (N414, N406, N276, N337, N319);
not NOT1 (N415, N399);
xor XOR2 (N416, N413, N218);
buf BUF1 (N417, N387);
nor NOR2 (N418, N412, N298);
and AND3 (N419, N380, N186, N216);
nand NAND4 (N420, N395, N346, N6, N117);
nor NOR4 (N421, N420, N393, N71, N275);
or OR3 (N422, N421, N16, N331);
nor NOR4 (N423, N416, N2, N32, N129);
or OR3 (N424, N422, N281, N2);
nor NOR3 (N425, N424, N283, N312);
or OR2 (N426, N404, N284);
nand NAND2 (N427, N415, N231);
nor NOR4 (N428, N423, N317, N51, N294);
nand NAND4 (N429, N427, N185, N293, N144);
not NOT1 (N430, N428);
nor NOR2 (N431, N425, N299);
nor NOR3 (N432, N418, N290, N37);
nand NAND4 (N433, N431, N339, N426, N255);
xor XOR2 (N434, N45, N341);
buf BUF1 (N435, N414);
xor XOR2 (N436, N429, N343);
nor NOR2 (N437, N417, N297);
and AND2 (N438, N396, N435);
buf BUF1 (N439, N326);
nor NOR2 (N440, N410, N280);
nand NAND3 (N441, N432, N330, N84);
nor NOR2 (N442, N434, N214);
not NOT1 (N443, N440);
or OR3 (N444, N439, N260, N72);
and AND2 (N445, N430, N172);
nand NAND4 (N446, N419, N374, N188, N261);
not NOT1 (N447, N437);
xor XOR2 (N448, N443, N339);
xor XOR2 (N449, N446, N317);
and AND3 (N450, N448, N417, N230);
buf BUF1 (N451, N445);
nor NOR3 (N452, N451, N380, N345);
nor NOR4 (N453, N436, N297, N65, N338);
buf BUF1 (N454, N442);
and AND2 (N455, N447, N82);
or OR2 (N456, N441, N187);
or OR2 (N457, N453, N186);
xor XOR2 (N458, N444, N331);
nor NOR3 (N459, N450, N128, N273);
nor NOR4 (N460, N457, N311, N55, N456);
xor XOR2 (N461, N249, N359);
and AND4 (N462, N452, N287, N350, N84);
and AND4 (N463, N438, N19, N278, N132);
or OR4 (N464, N463, N419, N255, N113);
and AND4 (N465, N461, N174, N365, N164);
nand NAND4 (N466, N458, N179, N128, N12);
nand NAND4 (N467, N465, N172, N413, N93);
nor NOR3 (N468, N433, N89, N66);
nor NOR3 (N469, N464, N334, N233);
not NOT1 (N470, N469);
nand NAND3 (N471, N460, N457, N467);
nor NOR4 (N472, N171, N98, N125, N418);
or OR3 (N473, N454, N201, N458);
or OR3 (N474, N472, N335, N18);
or OR3 (N475, N459, N156, N474);
nand NAND2 (N476, N280, N284);
or OR2 (N477, N473, N339);
or OR4 (N478, N476, N440, N137, N209);
buf BUF1 (N479, N478);
nor NOR3 (N480, N475, N410, N315);
nor NOR3 (N481, N480, N253, N360);
nand NAND4 (N482, N470, N243, N429, N448);
not NOT1 (N483, N462);
or OR3 (N484, N477, N299, N363);
xor XOR2 (N485, N471, N45);
or OR3 (N486, N468, N234, N315);
nand NAND4 (N487, N485, N324, N300, N75);
or OR4 (N488, N482, N444, N154, N192);
nor NOR4 (N489, N481, N271, N378, N10);
or OR2 (N490, N449, N452);
not NOT1 (N491, N483);
not NOT1 (N492, N487);
or OR3 (N493, N491, N221, N113);
not NOT1 (N494, N489);
buf BUF1 (N495, N494);
or OR2 (N496, N466, N394);
xor XOR2 (N497, N492, N257);
and AND4 (N498, N479, N332, N352, N104);
nor NOR2 (N499, N497, N196);
nor NOR4 (N500, N496, N18, N335, N135);
buf BUF1 (N501, N486);
nand NAND3 (N502, N455, N407, N114);
nand NAND3 (N503, N484, N66, N476);
not NOT1 (N504, N502);
or OR4 (N505, N493, N350, N287, N469);
nor NOR2 (N506, N501, N183);
nand NAND3 (N507, N506, N216, N490);
and AND4 (N508, N290, N55, N117, N461);
nand NAND2 (N509, N500, N342);
nand NAND3 (N510, N504, N83, N462);
buf BUF1 (N511, N498);
buf BUF1 (N512, N505);
nor NOR3 (N513, N499, N434, N413);
xor XOR2 (N514, N509, N497);
and AND4 (N515, N514, N355, N192, N116);
and AND3 (N516, N503, N285, N471);
buf BUF1 (N517, N510);
or OR3 (N518, N516, N269, N230);
or OR4 (N519, N511, N460, N465, N342);
not NOT1 (N520, N507);
or OR2 (N521, N518, N439);
and AND4 (N522, N517, N262, N17, N267);
nor NOR2 (N523, N513, N329);
and AND4 (N524, N523, N336, N229, N40);
and AND2 (N525, N520, N201);
xor XOR2 (N526, N495, N244);
not NOT1 (N527, N512);
xor XOR2 (N528, N508, N384);
or OR4 (N529, N521, N202, N521, N224);
nor NOR3 (N530, N522, N287, N21);
buf BUF1 (N531, N524);
or OR4 (N532, N526, N468, N422, N196);
not NOT1 (N533, N515);
buf BUF1 (N534, N529);
buf BUF1 (N535, N532);
not NOT1 (N536, N530);
xor XOR2 (N537, N488, N455);
not NOT1 (N538, N519);
buf BUF1 (N539, N535);
buf BUF1 (N540, N534);
nand NAND3 (N541, N540, N441, N441);
or OR4 (N542, N537, N27, N126, N326);
xor XOR2 (N543, N542, N160);
buf BUF1 (N544, N543);
buf BUF1 (N545, N536);
nor NOR4 (N546, N531, N56, N145, N388);
nor NOR4 (N547, N533, N48, N12, N114);
and AND3 (N548, N528, N56, N166);
and AND4 (N549, N548, N443, N268, N42);
xor XOR2 (N550, N527, N41);
xor XOR2 (N551, N525, N115);
xor XOR2 (N552, N546, N510);
xor XOR2 (N553, N545, N357);
buf BUF1 (N554, N544);
nand NAND2 (N555, N539, N550);
buf BUF1 (N556, N159);
nor NOR2 (N557, N551, N430);
and AND2 (N558, N553, N265);
buf BUF1 (N559, N541);
buf BUF1 (N560, N554);
buf BUF1 (N561, N557);
nor NOR3 (N562, N559, N337, N400);
buf BUF1 (N563, N555);
not NOT1 (N564, N538);
or OR4 (N565, N547, N553, N542, N269);
buf BUF1 (N566, N565);
nand NAND3 (N567, N558, N250, N459);
nor NOR2 (N568, N552, N193);
xor XOR2 (N569, N561, N229);
not NOT1 (N570, N569);
or OR2 (N571, N564, N366);
not NOT1 (N572, N562);
xor XOR2 (N573, N571, N472);
and AND4 (N574, N567, N271, N346, N548);
nand NAND3 (N575, N568, N265, N235);
nand NAND2 (N576, N570, N13);
nand NAND3 (N577, N576, N200, N305);
not NOT1 (N578, N575);
nor NOR2 (N579, N574, N373);
nand NAND2 (N580, N573, N270);
xor XOR2 (N581, N566, N406);
or OR2 (N582, N549, N363);
buf BUF1 (N583, N580);
xor XOR2 (N584, N577, N353);
buf BUF1 (N585, N584);
nor NOR4 (N586, N582, N254, N406, N154);
xor XOR2 (N587, N556, N427);
or OR4 (N588, N583, N534, N450, N18);
nand NAND2 (N589, N579, N170);
or OR2 (N590, N572, N24);
buf BUF1 (N591, N589);
nand NAND3 (N592, N578, N52, N522);
not NOT1 (N593, N581);
buf BUF1 (N594, N585);
or OR4 (N595, N591, N475, N119, N452);
nor NOR2 (N596, N593, N481);
nor NOR4 (N597, N587, N308, N447, N184);
and AND3 (N598, N586, N544, N550);
or OR3 (N599, N595, N435, N277);
or OR2 (N600, N594, N215);
nor NOR3 (N601, N596, N502, N338);
nor NOR4 (N602, N590, N75, N339, N8);
or OR4 (N603, N600, N503, N188, N139);
xor XOR2 (N604, N599, N221);
nand NAND4 (N605, N601, N236, N433, N469);
or OR3 (N606, N602, N195, N351);
or OR4 (N607, N588, N385, N21, N450);
buf BUF1 (N608, N607);
nand NAND2 (N609, N603, N161);
not NOT1 (N610, N598);
xor XOR2 (N611, N604, N67);
nand NAND2 (N612, N560, N490);
buf BUF1 (N613, N610);
nand NAND2 (N614, N609, N116);
and AND2 (N615, N605, N337);
nor NOR3 (N616, N614, N380, N512);
and AND2 (N617, N563, N326);
or OR2 (N618, N613, N269);
nand NAND3 (N619, N608, N293, N290);
nand NAND4 (N620, N618, N320, N207, N482);
and AND3 (N621, N606, N41, N166);
nand NAND3 (N622, N621, N429, N435);
and AND3 (N623, N616, N307, N8);
nor NOR3 (N624, N622, N443, N51);
and AND3 (N625, N611, N253, N476);
xor XOR2 (N626, N612, N84);
buf BUF1 (N627, N615);
or OR2 (N628, N625, N166);
or OR2 (N629, N626, N498);
nor NOR2 (N630, N617, N580);
not NOT1 (N631, N627);
xor XOR2 (N632, N628, N376);
xor XOR2 (N633, N619, N49);
buf BUF1 (N634, N632);
not NOT1 (N635, N631);
not NOT1 (N636, N635);
buf BUF1 (N637, N636);
not NOT1 (N638, N620);
or OR3 (N639, N638, N493, N30);
xor XOR2 (N640, N623, N220);
not NOT1 (N641, N634);
buf BUF1 (N642, N629);
not NOT1 (N643, N624);
or OR4 (N644, N640, N511, N196, N567);
xor XOR2 (N645, N597, N91);
and AND3 (N646, N645, N250, N621);
not NOT1 (N647, N633);
not NOT1 (N648, N630);
nand NAND4 (N649, N646, N551, N183, N449);
not NOT1 (N650, N637);
nand NAND4 (N651, N592, N491, N203, N53);
and AND3 (N652, N650, N212, N485);
xor XOR2 (N653, N643, N25);
buf BUF1 (N654, N647);
or OR2 (N655, N644, N543);
not NOT1 (N656, N653);
buf BUF1 (N657, N649);
and AND4 (N658, N657, N310, N13, N275);
nor NOR3 (N659, N641, N184, N23);
or OR2 (N660, N648, N275);
and AND4 (N661, N659, N343, N553, N157);
and AND4 (N662, N656, N45, N178, N337);
xor XOR2 (N663, N642, N465);
nand NAND3 (N664, N660, N373, N161);
xor XOR2 (N665, N661, N279);
nand NAND3 (N666, N658, N320, N18);
nand NAND2 (N667, N639, N110);
nand NAND2 (N668, N665, N399);
xor XOR2 (N669, N668, N398);
nor NOR3 (N670, N667, N213, N575);
xor XOR2 (N671, N663, N239);
nand NAND3 (N672, N651, N243, N328);
nand NAND2 (N673, N672, N22);
nor NOR4 (N674, N654, N278, N297, N286);
or OR2 (N675, N662, N282);
xor XOR2 (N676, N675, N271);
nand NAND2 (N677, N664, N218);
nor NOR3 (N678, N652, N386, N454);
not NOT1 (N679, N674);
not NOT1 (N680, N677);
and AND2 (N681, N671, N559);
nand NAND3 (N682, N678, N540, N667);
nor NOR3 (N683, N666, N614, N33);
xor XOR2 (N684, N680, N661);
not NOT1 (N685, N669);
xor XOR2 (N686, N685, N415);
nand NAND2 (N687, N679, N185);
and AND4 (N688, N673, N655, N403, N83);
xor XOR2 (N689, N337, N405);
not NOT1 (N690, N684);
not NOT1 (N691, N676);
or OR4 (N692, N687, N654, N74, N539);
not NOT1 (N693, N681);
or OR4 (N694, N692, N430, N416, N242);
not NOT1 (N695, N693);
or OR4 (N696, N670, N187, N125, N457);
buf BUF1 (N697, N683);
or OR3 (N698, N688, N251, N155);
and AND2 (N699, N695, N310);
not NOT1 (N700, N699);
nor NOR4 (N701, N698, N622, N553, N408);
nor NOR3 (N702, N691, N164, N304);
nor NOR2 (N703, N682, N30);
buf BUF1 (N704, N701);
nand NAND3 (N705, N696, N27, N495);
nand NAND2 (N706, N700, N177);
xor XOR2 (N707, N705, N548);
or OR4 (N708, N707, N492, N183, N15);
buf BUF1 (N709, N686);
buf BUF1 (N710, N690);
not NOT1 (N711, N708);
nor NOR3 (N712, N710, N616, N141);
buf BUF1 (N713, N703);
buf BUF1 (N714, N712);
buf BUF1 (N715, N704);
or OR4 (N716, N706, N510, N668, N631);
buf BUF1 (N717, N702);
and AND3 (N718, N689, N275, N584);
buf BUF1 (N719, N709);
not NOT1 (N720, N718);
or OR4 (N721, N720, N221, N426, N455);
or OR4 (N722, N716, N469, N649, N19);
nand NAND3 (N723, N711, N586, N66);
xor XOR2 (N724, N721, N209);
not NOT1 (N725, N714);
nand NAND4 (N726, N694, N376, N94, N602);
xor XOR2 (N727, N717, N661);
nor NOR2 (N728, N725, N137);
not NOT1 (N729, N715);
buf BUF1 (N730, N713);
or OR4 (N731, N724, N98, N142, N607);
and AND4 (N732, N731, N224, N259, N521);
not NOT1 (N733, N697);
xor XOR2 (N734, N727, N76);
not NOT1 (N735, N734);
and AND4 (N736, N719, N326, N295, N53);
or OR3 (N737, N730, N260, N163);
nor NOR4 (N738, N722, N518, N233, N263);
nand NAND2 (N739, N732, N412);
nor NOR3 (N740, N723, N300, N622);
xor XOR2 (N741, N729, N96);
buf BUF1 (N742, N736);
not NOT1 (N743, N726);
not NOT1 (N744, N738);
buf BUF1 (N745, N735);
xor XOR2 (N746, N745, N207);
buf BUF1 (N747, N740);
or OR3 (N748, N743, N442, N702);
or OR4 (N749, N739, N246, N156, N282);
nand NAND3 (N750, N749, N503, N556);
xor XOR2 (N751, N748, N604);
or OR3 (N752, N728, N612, N748);
buf BUF1 (N753, N741);
nor NOR4 (N754, N751, N37, N621, N149);
buf BUF1 (N755, N752);
nand NAND2 (N756, N747, N645);
not NOT1 (N757, N756);
not NOT1 (N758, N744);
not NOT1 (N759, N755);
buf BUF1 (N760, N759);
buf BUF1 (N761, N754);
nand NAND4 (N762, N737, N163, N279, N38);
and AND2 (N763, N750, N672);
or OR4 (N764, N761, N14, N203, N757);
or OR3 (N765, N224, N627, N222);
not NOT1 (N766, N758);
nor NOR4 (N767, N763, N546, N261, N214);
and AND4 (N768, N753, N310, N211, N473);
and AND2 (N769, N766, N651);
buf BUF1 (N770, N764);
nand NAND2 (N771, N765, N468);
buf BUF1 (N772, N746);
nand NAND4 (N773, N771, N609, N436, N21);
not NOT1 (N774, N760);
or OR3 (N775, N769, N638, N299);
buf BUF1 (N776, N773);
or OR2 (N777, N770, N623);
buf BUF1 (N778, N774);
nor NOR2 (N779, N742, N526);
xor XOR2 (N780, N775, N389);
not NOT1 (N781, N780);
xor XOR2 (N782, N767, N320);
and AND3 (N783, N777, N598, N227);
and AND3 (N784, N781, N346, N298);
nor NOR4 (N785, N733, N168, N170, N635);
or OR2 (N786, N772, N274);
buf BUF1 (N787, N783);
nand NAND3 (N788, N786, N761, N710);
or OR4 (N789, N776, N380, N568, N544);
xor XOR2 (N790, N785, N307);
or OR3 (N791, N787, N470, N64);
or OR2 (N792, N782, N54);
nor NOR4 (N793, N778, N660, N321, N566);
nand NAND2 (N794, N789, N105);
buf BUF1 (N795, N792);
xor XOR2 (N796, N779, N572);
buf BUF1 (N797, N762);
nand NAND2 (N798, N797, N49);
nand NAND4 (N799, N793, N312, N197, N10);
nand NAND2 (N800, N791, N82);
and AND3 (N801, N795, N622, N325);
nor NOR3 (N802, N788, N696, N267);
or OR3 (N803, N800, N661, N494);
and AND2 (N804, N768, N497);
buf BUF1 (N805, N801);
buf BUF1 (N806, N799);
xor XOR2 (N807, N784, N325);
buf BUF1 (N808, N804);
xor XOR2 (N809, N802, N801);
buf BUF1 (N810, N798);
xor XOR2 (N811, N810, N171);
xor XOR2 (N812, N807, N292);
nand NAND4 (N813, N806, N128, N168, N111);
nand NAND2 (N814, N812, N23);
nand NAND2 (N815, N811, N811);
nand NAND3 (N816, N803, N514, N715);
not NOT1 (N817, N813);
and AND2 (N818, N809, N604);
nand NAND2 (N819, N817, N5);
buf BUF1 (N820, N796);
xor XOR2 (N821, N818, N220);
xor XOR2 (N822, N815, N346);
xor XOR2 (N823, N816, N521);
buf BUF1 (N824, N794);
nand NAND2 (N825, N821, N120);
or OR3 (N826, N808, N342, N62);
not NOT1 (N827, N820);
or OR2 (N828, N822, N306);
or OR4 (N829, N827, N622, N743, N566);
nand NAND2 (N830, N824, N675);
or OR2 (N831, N830, N527);
xor XOR2 (N832, N825, N281);
and AND4 (N833, N819, N520, N416, N117);
nor NOR4 (N834, N826, N167, N679, N511);
and AND3 (N835, N834, N808, N90);
buf BUF1 (N836, N832);
xor XOR2 (N837, N805, N135);
not NOT1 (N838, N829);
and AND4 (N839, N833, N832, N297, N215);
or OR2 (N840, N790, N509);
nand NAND3 (N841, N814, N608, N279);
nor NOR4 (N842, N837, N238, N574, N662);
or OR2 (N843, N836, N218);
buf BUF1 (N844, N842);
buf BUF1 (N845, N831);
nand NAND4 (N846, N844, N109, N671, N186);
and AND4 (N847, N843, N490, N19, N246);
nor NOR4 (N848, N839, N150, N646, N406);
buf BUF1 (N849, N838);
nand NAND2 (N850, N848, N236);
not NOT1 (N851, N840);
not NOT1 (N852, N846);
or OR3 (N853, N841, N797, N629);
or OR3 (N854, N835, N206, N161);
nor NOR2 (N855, N852, N50);
nor NOR2 (N856, N855, N402);
or OR3 (N857, N851, N662, N382);
buf BUF1 (N858, N849);
xor XOR2 (N859, N856, N151);
xor XOR2 (N860, N845, N486);
or OR2 (N861, N860, N353);
not NOT1 (N862, N847);
or OR2 (N863, N853, N202);
buf BUF1 (N864, N828);
nand NAND2 (N865, N861, N462);
nand NAND3 (N866, N864, N424, N272);
buf BUF1 (N867, N857);
nor NOR3 (N868, N850, N305, N241);
xor XOR2 (N869, N858, N410);
and AND3 (N870, N868, N253, N788);
xor XOR2 (N871, N863, N276);
nand NAND4 (N872, N871, N127, N409, N762);
xor XOR2 (N873, N872, N719);
not NOT1 (N874, N870);
xor XOR2 (N875, N874, N458);
not NOT1 (N876, N875);
nand NAND3 (N877, N859, N689, N621);
not NOT1 (N878, N823);
nor NOR2 (N879, N854, N200);
not NOT1 (N880, N866);
buf BUF1 (N881, N876);
not NOT1 (N882, N881);
or OR2 (N883, N877, N400);
and AND2 (N884, N867, N257);
nand NAND3 (N885, N884, N524, N255);
or OR4 (N886, N885, N275, N361, N432);
and AND4 (N887, N862, N461, N584, N430);
xor XOR2 (N888, N878, N200);
and AND4 (N889, N869, N205, N225, N633);
xor XOR2 (N890, N886, N113);
buf BUF1 (N891, N890);
nand NAND2 (N892, N889, N603);
nor NOR3 (N893, N891, N368, N495);
nand NAND2 (N894, N887, N497);
nand NAND2 (N895, N893, N351);
xor XOR2 (N896, N865, N770);
nand NAND3 (N897, N882, N315, N290);
xor XOR2 (N898, N892, N155);
not NOT1 (N899, N896);
xor XOR2 (N900, N873, N721);
or OR3 (N901, N888, N491, N186);
and AND2 (N902, N899, N131);
xor XOR2 (N903, N902, N335);
not NOT1 (N904, N897);
or OR4 (N905, N879, N181, N672, N457);
nor NOR2 (N906, N880, N130);
xor XOR2 (N907, N883, N34);
nor NOR3 (N908, N906, N293, N387);
and AND3 (N909, N903, N544, N593);
nand NAND2 (N910, N909, N347);
not NOT1 (N911, N894);
not NOT1 (N912, N910);
and AND2 (N913, N904, N33);
and AND2 (N914, N895, N588);
or OR4 (N915, N908, N574, N475, N442);
buf BUF1 (N916, N912);
nand NAND3 (N917, N900, N726, N529);
not NOT1 (N918, N907);
and AND2 (N919, N915, N374);
buf BUF1 (N920, N913);
nand NAND3 (N921, N914, N726, N811);
or OR2 (N922, N918, N73);
xor XOR2 (N923, N921, N700);
or OR4 (N924, N911, N178, N171, N455);
and AND4 (N925, N923, N504, N156, N499);
nand NAND3 (N926, N901, N827, N327);
nor NOR4 (N927, N924, N223, N741, N203);
and AND2 (N928, N922, N352);
and AND3 (N929, N898, N427, N50);
buf BUF1 (N930, N920);
and AND3 (N931, N905, N878, N355);
or OR2 (N932, N926, N248);
buf BUF1 (N933, N932);
nand NAND4 (N934, N933, N465, N274, N402);
nor NOR3 (N935, N916, N275, N283);
not NOT1 (N936, N930);
not NOT1 (N937, N928);
nand NAND3 (N938, N937, N137, N481);
nor NOR2 (N939, N929, N915);
nand NAND4 (N940, N934, N217, N412, N545);
buf BUF1 (N941, N938);
not NOT1 (N942, N917);
or OR3 (N943, N942, N831, N434);
nor NOR2 (N944, N943, N642);
not NOT1 (N945, N919);
buf BUF1 (N946, N944);
xor XOR2 (N947, N927, N861);
nor NOR3 (N948, N935, N497, N339);
nand NAND4 (N949, N925, N110, N907, N56);
xor XOR2 (N950, N946, N777);
not NOT1 (N951, N948);
and AND2 (N952, N940, N788);
buf BUF1 (N953, N931);
not NOT1 (N954, N939);
and AND4 (N955, N951, N755, N5, N552);
buf BUF1 (N956, N936);
nor NOR4 (N957, N953, N53, N416, N2);
nor NOR4 (N958, N950, N776, N626, N588);
or OR4 (N959, N941, N588, N691, N182);
nor NOR4 (N960, N959, N330, N288, N120);
nand NAND2 (N961, N954, N478);
or OR2 (N962, N945, N734);
buf BUF1 (N963, N949);
nor NOR2 (N964, N958, N907);
nand NAND4 (N965, N963, N34, N503, N776);
nor NOR3 (N966, N957, N416, N426);
and AND4 (N967, N965, N230, N472, N830);
nand NAND2 (N968, N960, N665);
buf BUF1 (N969, N952);
buf BUF1 (N970, N962);
or OR3 (N971, N947, N728, N71);
buf BUF1 (N972, N964);
not NOT1 (N973, N969);
not NOT1 (N974, N966);
not NOT1 (N975, N968);
xor XOR2 (N976, N971, N937);
xor XOR2 (N977, N955, N390);
nor NOR3 (N978, N977, N332, N179);
not NOT1 (N979, N978);
or OR3 (N980, N975, N14, N642);
nor NOR3 (N981, N970, N290, N487);
buf BUF1 (N982, N979);
nor NOR3 (N983, N956, N350, N840);
nand NAND2 (N984, N972, N627);
nor NOR3 (N985, N984, N359, N689);
not NOT1 (N986, N961);
buf BUF1 (N987, N980);
buf BUF1 (N988, N973);
and AND3 (N989, N967, N10, N943);
and AND2 (N990, N983, N282);
nand NAND3 (N991, N985, N662, N990);
nand NAND2 (N992, N615, N43);
and AND2 (N993, N988, N29);
nor NOR4 (N994, N986, N600, N437, N581);
nor NOR2 (N995, N991, N408);
or OR3 (N996, N995, N127, N386);
or OR2 (N997, N992, N717);
nor NOR3 (N998, N989, N814, N387);
xor XOR2 (N999, N993, N320);
nand NAND4 (N1000, N999, N345, N110, N824);
or OR3 (N1001, N982, N258, N190);
and AND2 (N1002, N1000, N85);
not NOT1 (N1003, N1002);
buf BUF1 (N1004, N996);
not NOT1 (N1005, N987);
nand NAND4 (N1006, N1003, N553, N722, N101);
buf BUF1 (N1007, N1006);
nand NAND3 (N1008, N994, N410, N892);
and AND3 (N1009, N997, N404, N840);
buf BUF1 (N1010, N1009);
or OR4 (N1011, N998, N930, N768, N651);
or OR2 (N1012, N1001, N819);
or OR2 (N1013, N981, N591);
nand NAND3 (N1014, N974, N954, N450);
or OR2 (N1015, N1007, N28);
buf BUF1 (N1016, N976);
and AND2 (N1017, N1005, N320);
xor XOR2 (N1018, N1013, N800);
not NOT1 (N1019, N1015);
or OR4 (N1020, N1012, N4, N866, N93);
not NOT1 (N1021, N1016);
and AND3 (N1022, N1010, N526, N215);
xor XOR2 (N1023, N1017, N796);
or OR3 (N1024, N1020, N472, N391);
or OR2 (N1025, N1011, N66);
nor NOR3 (N1026, N1025, N134, N144);
and AND3 (N1027, N1023, N788, N548);
not NOT1 (N1028, N1021);
nor NOR3 (N1029, N1019, N236, N577);
or OR3 (N1030, N1022, N53, N537);
nand NAND3 (N1031, N1030, N222, N362);
not NOT1 (N1032, N1026);
not NOT1 (N1033, N1028);
nand NAND2 (N1034, N1032, N249);
xor XOR2 (N1035, N1008, N802);
buf BUF1 (N1036, N1018);
and AND2 (N1037, N1029, N368);
not NOT1 (N1038, N1035);
nand NAND3 (N1039, N1004, N841, N30);
not NOT1 (N1040, N1027);
xor XOR2 (N1041, N1033, N113);
nor NOR4 (N1042, N1037, N431, N722, N919);
and AND3 (N1043, N1038, N1027, N904);
and AND2 (N1044, N1034, N556);
or OR3 (N1045, N1014, N1021, N740);
not NOT1 (N1046, N1043);
nor NOR3 (N1047, N1024, N92, N976);
not NOT1 (N1048, N1036);
or OR3 (N1049, N1048, N580, N812);
not NOT1 (N1050, N1045);
and AND4 (N1051, N1040, N892, N114, N17);
buf BUF1 (N1052, N1044);
buf BUF1 (N1053, N1050);
buf BUF1 (N1054, N1031);
nand NAND2 (N1055, N1052, N17);
or OR4 (N1056, N1055, N273, N550, N666);
nand NAND2 (N1057, N1041, N512);
nor NOR4 (N1058, N1049, N241, N294, N265);
not NOT1 (N1059, N1039);
and AND4 (N1060, N1047, N860, N29, N272);
nor NOR2 (N1061, N1057, N691);
nand NAND3 (N1062, N1058, N738, N280);
and AND2 (N1063, N1053, N518);
nor NOR3 (N1064, N1062, N493, N1026);
nor NOR3 (N1065, N1056, N724, N778);
xor XOR2 (N1066, N1054, N254);
and AND4 (N1067, N1061, N866, N383, N853);
nand NAND4 (N1068, N1059, N593, N59, N941);
xor XOR2 (N1069, N1065, N635);
buf BUF1 (N1070, N1067);
and AND4 (N1071, N1060, N573, N791, N892);
xor XOR2 (N1072, N1066, N31);
buf BUF1 (N1073, N1070);
nor NOR4 (N1074, N1046, N997, N701, N252);
or OR2 (N1075, N1072, N607);
nand NAND3 (N1076, N1075, N351, N1038);
not NOT1 (N1077, N1042);
and AND2 (N1078, N1063, N413);
not NOT1 (N1079, N1074);
xor XOR2 (N1080, N1076, N330);
and AND3 (N1081, N1078, N48, N614);
nor NOR4 (N1082, N1051, N288, N441, N389);
xor XOR2 (N1083, N1071, N516);
buf BUF1 (N1084, N1073);
xor XOR2 (N1085, N1069, N404);
nand NAND4 (N1086, N1064, N522, N538, N480);
and AND2 (N1087, N1082, N414);
not NOT1 (N1088, N1080);
or OR4 (N1089, N1084, N820, N593, N57);
not NOT1 (N1090, N1085);
nor NOR3 (N1091, N1086, N1081, N959);
xor XOR2 (N1092, N561, N122);
or OR2 (N1093, N1083, N301);
and AND4 (N1094, N1090, N455, N966, N131);
xor XOR2 (N1095, N1091, N7);
not NOT1 (N1096, N1077);
buf BUF1 (N1097, N1094);
buf BUF1 (N1098, N1095);
xor XOR2 (N1099, N1096, N194);
and AND2 (N1100, N1068, N105);
nor NOR4 (N1101, N1093, N908, N777, N522);
not NOT1 (N1102, N1101);
not NOT1 (N1103, N1102);
nand NAND2 (N1104, N1098, N755);
and AND2 (N1105, N1099, N461);
or OR4 (N1106, N1100, N925, N524, N859);
and AND2 (N1107, N1097, N691);
not NOT1 (N1108, N1105);
xor XOR2 (N1109, N1087, N539);
xor XOR2 (N1110, N1089, N399);
or OR3 (N1111, N1106, N872, N314);
and AND4 (N1112, N1092, N719, N346, N40);
buf BUF1 (N1113, N1103);
buf BUF1 (N1114, N1088);
and AND3 (N1115, N1111, N819, N672);
xor XOR2 (N1116, N1112, N100);
and AND3 (N1117, N1107, N848, N68);
and AND2 (N1118, N1113, N930);
and AND2 (N1119, N1110, N675);
nor NOR3 (N1120, N1115, N525, N831);
buf BUF1 (N1121, N1119);
not NOT1 (N1122, N1116);
nor NOR4 (N1123, N1108, N268, N743, N24);
nor NOR4 (N1124, N1114, N156, N741, N691);
and AND2 (N1125, N1122, N925);
xor XOR2 (N1126, N1109, N261);
and AND3 (N1127, N1121, N821, N1106);
and AND2 (N1128, N1127, N171);
buf BUF1 (N1129, N1079);
xor XOR2 (N1130, N1104, N289);
and AND4 (N1131, N1130, N496, N1085, N197);
and AND2 (N1132, N1120, N1013);
xor XOR2 (N1133, N1128, N413);
nor NOR2 (N1134, N1117, N208);
xor XOR2 (N1135, N1126, N54);
nand NAND2 (N1136, N1124, N916);
not NOT1 (N1137, N1131);
xor XOR2 (N1138, N1129, N456);
buf BUF1 (N1139, N1123);
nand NAND4 (N1140, N1136, N856, N777, N1074);
buf BUF1 (N1141, N1125);
nor NOR4 (N1142, N1140, N466, N1014, N197);
buf BUF1 (N1143, N1135);
and AND4 (N1144, N1138, N287, N52, N957);
nand NAND4 (N1145, N1118, N235, N618, N226);
buf BUF1 (N1146, N1137);
xor XOR2 (N1147, N1133, N432);
and AND2 (N1148, N1147, N1089);
or OR3 (N1149, N1148, N905, N1064);
nand NAND2 (N1150, N1141, N411);
xor XOR2 (N1151, N1150, N806);
nor NOR2 (N1152, N1132, N286);
or OR3 (N1153, N1143, N1027, N368);
xor XOR2 (N1154, N1145, N918);
and AND4 (N1155, N1154, N672, N762, N856);
nand NAND3 (N1156, N1155, N1110, N430);
nand NAND2 (N1157, N1134, N628);
not NOT1 (N1158, N1152);
nor NOR4 (N1159, N1153, N237, N648, N692);
nand NAND2 (N1160, N1158, N1098);
not NOT1 (N1161, N1139);
or OR3 (N1162, N1161, N133, N753);
not NOT1 (N1163, N1156);
and AND2 (N1164, N1162, N801);
not NOT1 (N1165, N1144);
not NOT1 (N1166, N1151);
not NOT1 (N1167, N1142);
or OR2 (N1168, N1163, N603);
or OR2 (N1169, N1166, N64);
and AND2 (N1170, N1160, N365);
not NOT1 (N1171, N1157);
not NOT1 (N1172, N1167);
buf BUF1 (N1173, N1172);
not NOT1 (N1174, N1146);
or OR3 (N1175, N1168, N227, N1094);
xor XOR2 (N1176, N1165, N769);
or OR2 (N1177, N1159, N1159);
buf BUF1 (N1178, N1174);
nand NAND2 (N1179, N1149, N859);
not NOT1 (N1180, N1171);
not NOT1 (N1181, N1175);
xor XOR2 (N1182, N1179, N483);
or OR4 (N1183, N1180, N331, N956, N10);
nand NAND2 (N1184, N1182, N732);
buf BUF1 (N1185, N1177);
buf BUF1 (N1186, N1178);
nor NOR4 (N1187, N1184, N240, N883, N604);
not NOT1 (N1188, N1183);
nor NOR2 (N1189, N1186, N47);
not NOT1 (N1190, N1173);
nand NAND2 (N1191, N1187, N323);
nand NAND3 (N1192, N1170, N1171, N505);
nor NOR3 (N1193, N1189, N435, N1021);
buf BUF1 (N1194, N1164);
and AND2 (N1195, N1185, N127);
xor XOR2 (N1196, N1191, N578);
not NOT1 (N1197, N1188);
or OR3 (N1198, N1181, N922, N539);
not NOT1 (N1199, N1176);
and AND3 (N1200, N1199, N239, N294);
xor XOR2 (N1201, N1196, N75);
nor NOR4 (N1202, N1190, N533, N834, N605);
nand NAND2 (N1203, N1200, N754);
not NOT1 (N1204, N1203);
buf BUF1 (N1205, N1193);
not NOT1 (N1206, N1202);
buf BUF1 (N1207, N1205);
xor XOR2 (N1208, N1169, N427);
not NOT1 (N1209, N1201);
or OR4 (N1210, N1207, N212, N74, N30);
xor XOR2 (N1211, N1197, N1093);
not NOT1 (N1212, N1209);
xor XOR2 (N1213, N1211, N889);
and AND2 (N1214, N1206, N328);
and AND3 (N1215, N1214, N1147, N446);
nand NAND4 (N1216, N1215, N352, N919, N1140);
or OR4 (N1217, N1204, N111, N1139, N1161);
and AND2 (N1218, N1212, N282);
xor XOR2 (N1219, N1194, N374);
or OR4 (N1220, N1198, N756, N809, N243);
nor NOR2 (N1221, N1213, N135);
nand NAND4 (N1222, N1220, N1124, N965, N257);
nand NAND3 (N1223, N1195, N1052, N5);
nand NAND4 (N1224, N1216, N155, N698, N49);
nor NOR3 (N1225, N1217, N137, N789);
nand NAND4 (N1226, N1224, N314, N1032, N857);
and AND4 (N1227, N1192, N485, N858, N672);
or OR4 (N1228, N1218, N476, N470, N132);
nand NAND2 (N1229, N1208, N504);
nor NOR2 (N1230, N1229, N275);
nor NOR2 (N1231, N1230, N968);
xor XOR2 (N1232, N1226, N1220);
and AND2 (N1233, N1219, N1086);
xor XOR2 (N1234, N1231, N162);
not NOT1 (N1235, N1227);
xor XOR2 (N1236, N1223, N923);
nor NOR4 (N1237, N1221, N230, N730, N400);
and AND4 (N1238, N1232, N229, N454, N1076);
buf BUF1 (N1239, N1237);
and AND2 (N1240, N1225, N410);
and AND3 (N1241, N1236, N198, N940);
not NOT1 (N1242, N1222);
and AND4 (N1243, N1210, N130, N104, N661);
not NOT1 (N1244, N1242);
or OR4 (N1245, N1241, N409, N845, N673);
and AND2 (N1246, N1228, N1070);
and AND2 (N1247, N1240, N530);
and AND2 (N1248, N1243, N221);
nand NAND2 (N1249, N1238, N91);
nor NOR2 (N1250, N1247, N102);
nor NOR4 (N1251, N1246, N995, N1008, N1129);
or OR4 (N1252, N1234, N423, N907, N1087);
buf BUF1 (N1253, N1250);
not NOT1 (N1254, N1235);
nor NOR4 (N1255, N1239, N811, N662, N502);
or OR2 (N1256, N1233, N466);
xor XOR2 (N1257, N1256, N675);
xor XOR2 (N1258, N1251, N662);
nor NOR3 (N1259, N1255, N580, N375);
buf BUF1 (N1260, N1248);
or OR4 (N1261, N1260, N877, N567, N836);
and AND2 (N1262, N1249, N52);
xor XOR2 (N1263, N1257, N860);
or OR4 (N1264, N1261, N61, N436, N600);
and AND3 (N1265, N1263, N60, N41);
and AND2 (N1266, N1254, N876);
xor XOR2 (N1267, N1264, N97);
xor XOR2 (N1268, N1259, N333);
buf BUF1 (N1269, N1267);
or OR3 (N1270, N1262, N1145, N343);
xor XOR2 (N1271, N1270, N904);
nor NOR3 (N1272, N1253, N1193, N1065);
or OR4 (N1273, N1245, N419, N265, N892);
nor NOR3 (N1274, N1252, N1009, N520);
xor XOR2 (N1275, N1274, N926);
nand NAND3 (N1276, N1265, N1010, N13);
nand NAND2 (N1277, N1258, N1153);
nand NAND2 (N1278, N1273, N578);
buf BUF1 (N1279, N1269);
not NOT1 (N1280, N1272);
nor NOR2 (N1281, N1275, N643);
xor XOR2 (N1282, N1266, N493);
nor NOR3 (N1283, N1268, N1193, N1049);
xor XOR2 (N1284, N1278, N1020);
or OR3 (N1285, N1282, N331, N1140);
nand NAND2 (N1286, N1277, N946);
not NOT1 (N1287, N1244);
not NOT1 (N1288, N1281);
xor XOR2 (N1289, N1286, N1175);
nor NOR4 (N1290, N1276, N749, N428, N1189);
not NOT1 (N1291, N1287);
or OR4 (N1292, N1280, N961, N785, N853);
nand NAND3 (N1293, N1284, N1060, N961);
nor NOR2 (N1294, N1291, N608);
buf BUF1 (N1295, N1292);
or OR4 (N1296, N1295, N1242, N506, N496);
or OR4 (N1297, N1288, N269, N949, N926);
and AND3 (N1298, N1271, N712, N373);
nor NOR4 (N1299, N1293, N658, N257, N374);
or OR4 (N1300, N1289, N928, N1146, N200);
buf BUF1 (N1301, N1290);
nor NOR4 (N1302, N1301, N327, N926, N601);
xor XOR2 (N1303, N1285, N1213);
nand NAND4 (N1304, N1279, N830, N917, N35);
nor NOR2 (N1305, N1300, N644);
not NOT1 (N1306, N1296);
xor XOR2 (N1307, N1303, N670);
or OR4 (N1308, N1302, N624, N124, N786);
nand NAND2 (N1309, N1297, N968);
or OR3 (N1310, N1299, N419, N982);
or OR2 (N1311, N1310, N804);
or OR3 (N1312, N1308, N1291, N1289);
xor XOR2 (N1313, N1305, N1166);
xor XOR2 (N1314, N1307, N311);
buf BUF1 (N1315, N1304);
xor XOR2 (N1316, N1313, N567);
not NOT1 (N1317, N1306);
not NOT1 (N1318, N1315);
or OR2 (N1319, N1298, N489);
nor NOR2 (N1320, N1319, N814);
not NOT1 (N1321, N1316);
xor XOR2 (N1322, N1294, N292);
nand NAND4 (N1323, N1317, N251, N646, N1033);
xor XOR2 (N1324, N1323, N1017);
buf BUF1 (N1325, N1311);
nor NOR4 (N1326, N1318, N497, N425, N131);
xor XOR2 (N1327, N1324, N344);
and AND3 (N1328, N1322, N263, N936);
and AND2 (N1329, N1325, N1288);
nor NOR4 (N1330, N1329, N831, N770, N1151);
not NOT1 (N1331, N1328);
nor NOR4 (N1332, N1309, N794, N1141, N1088);
xor XOR2 (N1333, N1326, N924);
nand NAND4 (N1334, N1330, N849, N872, N46);
buf BUF1 (N1335, N1312);
buf BUF1 (N1336, N1314);
xor XOR2 (N1337, N1327, N14);
or OR2 (N1338, N1321, N1093);
buf BUF1 (N1339, N1334);
nor NOR3 (N1340, N1337, N778, N124);
and AND4 (N1341, N1320, N930, N206, N695);
or OR2 (N1342, N1340, N830);
xor XOR2 (N1343, N1332, N57);
and AND3 (N1344, N1342, N627, N1008);
not NOT1 (N1345, N1335);
nand NAND2 (N1346, N1333, N699);
buf BUF1 (N1347, N1343);
not NOT1 (N1348, N1341);
xor XOR2 (N1349, N1346, N942);
not NOT1 (N1350, N1339);
or OR2 (N1351, N1350, N1157);
buf BUF1 (N1352, N1338);
buf BUF1 (N1353, N1348);
not NOT1 (N1354, N1349);
nor NOR2 (N1355, N1353, N757);
and AND3 (N1356, N1355, N977, N407);
xor XOR2 (N1357, N1352, N1259);
xor XOR2 (N1358, N1336, N325);
not NOT1 (N1359, N1344);
nor NOR4 (N1360, N1354, N918, N188, N1289);
or OR3 (N1361, N1345, N1054, N1313);
not NOT1 (N1362, N1356);
buf BUF1 (N1363, N1362);
not NOT1 (N1364, N1331);
and AND4 (N1365, N1357, N717, N1056, N321);
buf BUF1 (N1366, N1361);
nand NAND4 (N1367, N1364, N1020, N1261, N1327);
not NOT1 (N1368, N1366);
and AND2 (N1369, N1358, N293);
nor NOR3 (N1370, N1363, N1288, N864);
and AND4 (N1371, N1347, N1181, N812, N254);
and AND4 (N1372, N1371, N1190, N882, N1280);
buf BUF1 (N1373, N1369);
buf BUF1 (N1374, N1372);
and AND3 (N1375, N1374, N1369, N1210);
not NOT1 (N1376, N1351);
xor XOR2 (N1377, N1375, N866);
buf BUF1 (N1378, N1365);
not NOT1 (N1379, N1283);
nor NOR2 (N1380, N1378, N894);
buf BUF1 (N1381, N1368);
not NOT1 (N1382, N1373);
nand NAND2 (N1383, N1382, N946);
not NOT1 (N1384, N1380);
nand NAND3 (N1385, N1359, N1055, N667);
nand NAND4 (N1386, N1381, N585, N549, N570);
xor XOR2 (N1387, N1385, N1042);
or OR4 (N1388, N1383, N310, N987, N271);
nand NAND3 (N1389, N1370, N148, N1188);
and AND4 (N1390, N1377, N282, N330, N966);
nand NAND3 (N1391, N1386, N793, N481);
or OR2 (N1392, N1384, N812);
xor XOR2 (N1393, N1392, N4);
nand NAND4 (N1394, N1367, N1307, N1164, N267);
buf BUF1 (N1395, N1391);
not NOT1 (N1396, N1379);
or OR4 (N1397, N1393, N346, N1300, N1124);
xor XOR2 (N1398, N1396, N497);
buf BUF1 (N1399, N1387);
nand NAND3 (N1400, N1399, N984, N545);
not NOT1 (N1401, N1398);
nor NOR4 (N1402, N1400, N640, N420, N1201);
nor NOR3 (N1403, N1390, N501, N923);
or OR4 (N1404, N1360, N999, N2, N993);
nand NAND2 (N1405, N1395, N19);
or OR3 (N1406, N1403, N822, N1302);
nand NAND3 (N1407, N1394, N1120, N55);
buf BUF1 (N1408, N1397);
xor XOR2 (N1409, N1405, N605);
or OR3 (N1410, N1388, N1033, N199);
not NOT1 (N1411, N1410);
or OR2 (N1412, N1409, N898);
xor XOR2 (N1413, N1407, N1003);
xor XOR2 (N1414, N1402, N484);
and AND4 (N1415, N1414, N221, N670, N1270);
nand NAND4 (N1416, N1412, N89, N21, N503);
or OR4 (N1417, N1415, N472, N533, N1298);
buf BUF1 (N1418, N1417);
nand NAND2 (N1419, N1404, N437);
or OR2 (N1420, N1418, N885);
xor XOR2 (N1421, N1389, N254);
nand NAND4 (N1422, N1420, N484, N58, N1135);
or OR2 (N1423, N1411, N1234);
nand NAND3 (N1424, N1408, N711, N1141);
not NOT1 (N1425, N1422);
and AND2 (N1426, N1416, N186);
buf BUF1 (N1427, N1413);
and AND4 (N1428, N1426, N387, N1312, N826);
nor NOR2 (N1429, N1424, N130);
and AND2 (N1430, N1425, N721);
nor NOR2 (N1431, N1428, N1357);
or OR4 (N1432, N1421, N215, N306, N895);
or OR4 (N1433, N1427, N665, N668, N349);
or OR4 (N1434, N1423, N609, N546, N886);
buf BUF1 (N1435, N1429);
xor XOR2 (N1436, N1434, N561);
nor NOR2 (N1437, N1430, N317);
and AND3 (N1438, N1436, N510, N1055);
and AND2 (N1439, N1431, N861);
and AND2 (N1440, N1419, N1367);
and AND2 (N1441, N1437, N1268);
and AND4 (N1442, N1433, N822, N1213, N185);
nor NOR2 (N1443, N1401, N1388);
nor NOR2 (N1444, N1432, N994);
nand NAND2 (N1445, N1438, N783);
nor NOR2 (N1446, N1435, N1192);
not NOT1 (N1447, N1376);
buf BUF1 (N1448, N1406);
or OR2 (N1449, N1445, N795);
or OR4 (N1450, N1444, N37, N571, N316);
or OR4 (N1451, N1446, N554, N100, N120);
xor XOR2 (N1452, N1443, N938);
nand NAND2 (N1453, N1448, N53);
not NOT1 (N1454, N1451);
or OR4 (N1455, N1439, N1042, N1199, N939);
buf BUF1 (N1456, N1452);
nand NAND3 (N1457, N1453, N532, N1440);
buf BUF1 (N1458, N1392);
not NOT1 (N1459, N1450);
xor XOR2 (N1460, N1454, N1130);
xor XOR2 (N1461, N1441, N870);
or OR3 (N1462, N1455, N914, N1171);
or OR3 (N1463, N1447, N75, N451);
xor XOR2 (N1464, N1462, N49);
nor NOR3 (N1465, N1464, N1130, N637);
nand NAND3 (N1466, N1457, N667, N458);
nand NAND3 (N1467, N1461, N1330, N1280);
nand NAND3 (N1468, N1465, N932, N1304);
nand NAND2 (N1469, N1468, N242);
not NOT1 (N1470, N1449);
and AND3 (N1471, N1456, N1442, N1358);
nor NOR3 (N1472, N265, N1168, N372);
nand NAND3 (N1473, N1467, N1205, N30);
not NOT1 (N1474, N1459);
xor XOR2 (N1475, N1466, N761);
and AND2 (N1476, N1469, N16);
xor XOR2 (N1477, N1470, N911);
not NOT1 (N1478, N1475);
and AND2 (N1479, N1477, N156);
not NOT1 (N1480, N1463);
and AND4 (N1481, N1478, N1144, N819, N74);
or OR2 (N1482, N1471, N698);
buf BUF1 (N1483, N1481);
xor XOR2 (N1484, N1479, N62);
not NOT1 (N1485, N1460);
buf BUF1 (N1486, N1474);
not NOT1 (N1487, N1476);
nor NOR3 (N1488, N1473, N346, N1442);
not NOT1 (N1489, N1480);
or OR2 (N1490, N1472, N1219);
nand NAND3 (N1491, N1485, N1332, N1387);
nor NOR4 (N1492, N1486, N1222, N1299, N842);
nand NAND4 (N1493, N1489, N206, N1206, N1262);
or OR4 (N1494, N1488, N1466, N710, N288);
nand NAND2 (N1495, N1487, N644);
not NOT1 (N1496, N1494);
nand NAND4 (N1497, N1491, N1025, N977, N1126);
or OR3 (N1498, N1483, N1121, N757);
xor XOR2 (N1499, N1496, N1069);
or OR3 (N1500, N1492, N1114, N529);
xor XOR2 (N1501, N1499, N1421);
xor XOR2 (N1502, N1500, N1366);
xor XOR2 (N1503, N1501, N221);
or OR3 (N1504, N1502, N30, N725);
or OR4 (N1505, N1504, N627, N78, N1323);
not NOT1 (N1506, N1497);
and AND3 (N1507, N1458, N190, N1306);
or OR3 (N1508, N1482, N306, N112);
not NOT1 (N1509, N1506);
not NOT1 (N1510, N1509);
or OR4 (N1511, N1505, N153, N546, N85);
and AND3 (N1512, N1507, N833, N1434);
xor XOR2 (N1513, N1484, N163);
nand NAND2 (N1514, N1493, N1414);
nand NAND2 (N1515, N1514, N471);
and AND2 (N1516, N1513, N1449);
nor NOR3 (N1517, N1515, N789, N1047);
nor NOR2 (N1518, N1516, N260);
not NOT1 (N1519, N1498);
buf BUF1 (N1520, N1508);
nor NOR4 (N1521, N1517, N285, N560, N1133);
nor NOR3 (N1522, N1490, N858, N970);
nand NAND4 (N1523, N1521, N439, N1420, N1025);
and AND2 (N1524, N1523, N812);
and AND2 (N1525, N1524, N647);
and AND2 (N1526, N1518, N374);
or OR4 (N1527, N1503, N1245, N97, N1351);
not NOT1 (N1528, N1526);
not NOT1 (N1529, N1525);
or OR4 (N1530, N1520, N877, N540, N908);
nand NAND3 (N1531, N1529, N1041, N894);
or OR4 (N1532, N1512, N674, N424, N434);
nand NAND2 (N1533, N1531, N1065);
or OR2 (N1534, N1532, N112);
nand NAND3 (N1535, N1527, N22, N918);
and AND3 (N1536, N1528, N401, N1406);
not NOT1 (N1537, N1519);
buf BUF1 (N1538, N1535);
buf BUF1 (N1539, N1538);
or OR3 (N1540, N1537, N610, N77);
nor NOR3 (N1541, N1540, N952, N336);
and AND3 (N1542, N1541, N40, N1417);
and AND4 (N1543, N1511, N1156, N136, N674);
nor NOR2 (N1544, N1533, N1486);
nor NOR2 (N1545, N1536, N1030);
not NOT1 (N1546, N1530);
nand NAND4 (N1547, N1546, N424, N523, N706);
nand NAND3 (N1548, N1542, N599, N1486);
and AND2 (N1549, N1522, N932);
not NOT1 (N1550, N1545);
or OR4 (N1551, N1550, N413, N818, N7);
not NOT1 (N1552, N1547);
nor NOR2 (N1553, N1551, N1299);
nor NOR2 (N1554, N1548, N529);
buf BUF1 (N1555, N1553);
and AND3 (N1556, N1549, N437, N1297);
nand NAND3 (N1557, N1510, N1484, N820);
not NOT1 (N1558, N1557);
not NOT1 (N1559, N1558);
nor NOR4 (N1560, N1544, N1263, N234, N900);
nand NAND3 (N1561, N1555, N1452, N1147);
or OR2 (N1562, N1559, N154);
buf BUF1 (N1563, N1562);
and AND4 (N1564, N1495, N1527, N61, N473);
buf BUF1 (N1565, N1543);
and AND3 (N1566, N1565, N1561, N417);
buf BUF1 (N1567, N1134);
or OR4 (N1568, N1552, N178, N412, N1426);
and AND4 (N1569, N1560, N752, N443, N521);
nor NOR3 (N1570, N1564, N351, N57);
and AND2 (N1571, N1569, N766);
not NOT1 (N1572, N1554);
and AND2 (N1573, N1556, N1336);
buf BUF1 (N1574, N1568);
buf BUF1 (N1575, N1567);
buf BUF1 (N1576, N1572);
and AND2 (N1577, N1571, N1211);
or OR3 (N1578, N1575, N844, N1047);
nand NAND2 (N1579, N1566, N735);
and AND3 (N1580, N1570, N506, N654);
not NOT1 (N1581, N1576);
buf BUF1 (N1582, N1578);
nor NOR4 (N1583, N1577, N500, N424, N446);
not NOT1 (N1584, N1563);
or OR4 (N1585, N1582, N147, N959, N25);
nand NAND4 (N1586, N1574, N1102, N1177, N703);
buf BUF1 (N1587, N1585);
or OR4 (N1588, N1581, N760, N325, N827);
nor NOR3 (N1589, N1580, N71, N549);
or OR4 (N1590, N1589, N1572, N1425, N440);
and AND4 (N1591, N1583, N815, N1403, N785);
nand NAND4 (N1592, N1539, N724, N924, N1037);
or OR2 (N1593, N1592, N1516);
and AND2 (N1594, N1579, N1397);
nor NOR3 (N1595, N1593, N1287, N812);
nor NOR2 (N1596, N1591, N1228);
xor XOR2 (N1597, N1595, N641);
nor NOR2 (N1598, N1597, N182);
nand NAND2 (N1599, N1586, N1428);
xor XOR2 (N1600, N1596, N151);
xor XOR2 (N1601, N1587, N664);
or OR3 (N1602, N1590, N1373, N1290);
nand NAND3 (N1603, N1600, N762, N411);
nand NAND4 (N1604, N1603, N36, N1596, N266);
xor XOR2 (N1605, N1602, N644);
xor XOR2 (N1606, N1594, N776);
nor NOR4 (N1607, N1588, N885, N1272, N616);
not NOT1 (N1608, N1605);
xor XOR2 (N1609, N1608, N965);
xor XOR2 (N1610, N1604, N641);
and AND3 (N1611, N1599, N892, N704);
or OR4 (N1612, N1534, N654, N477, N687);
not NOT1 (N1613, N1598);
or OR4 (N1614, N1573, N886, N110, N882);
or OR4 (N1615, N1606, N885, N1401, N1446);
and AND3 (N1616, N1615, N257, N1190);
and AND4 (N1617, N1609, N175, N166, N556);
or OR4 (N1618, N1617, N947, N10, N631);
or OR4 (N1619, N1584, N471, N1415, N1311);
or OR3 (N1620, N1607, N467, N234);
not NOT1 (N1621, N1614);
or OR2 (N1622, N1612, N1565);
nand NAND2 (N1623, N1610, N201);
xor XOR2 (N1624, N1623, N1473);
nand NAND4 (N1625, N1619, N1210, N963, N73);
xor XOR2 (N1626, N1618, N241);
and AND3 (N1627, N1625, N439, N893);
buf BUF1 (N1628, N1627);
nor NOR3 (N1629, N1626, N1290, N598);
nor NOR2 (N1630, N1629, N573);
nand NAND3 (N1631, N1628, N803, N878);
nand NAND4 (N1632, N1620, N651, N1367, N1193);
buf BUF1 (N1633, N1613);
nor NOR4 (N1634, N1630, N375, N1071, N390);
or OR4 (N1635, N1616, N1469, N414, N612);
nor NOR3 (N1636, N1611, N48, N986);
or OR2 (N1637, N1636, N1118);
and AND4 (N1638, N1633, N675, N718, N1057);
nor NOR4 (N1639, N1622, N277, N778, N199);
not NOT1 (N1640, N1601);
nand NAND4 (N1641, N1632, N214, N1502, N579);
and AND4 (N1642, N1621, N44, N1096, N77);
nor NOR2 (N1643, N1639, N1503);
buf BUF1 (N1644, N1635);
nand NAND2 (N1645, N1642, N1190);
and AND2 (N1646, N1643, N1313);
xor XOR2 (N1647, N1631, N6);
and AND2 (N1648, N1640, N343);
or OR2 (N1649, N1644, N1206);
nor NOR3 (N1650, N1634, N1316, N170);
xor XOR2 (N1651, N1645, N504);
not NOT1 (N1652, N1649);
nand NAND2 (N1653, N1637, N1024);
nor NOR2 (N1654, N1653, N590);
buf BUF1 (N1655, N1648);
and AND4 (N1656, N1655, N773, N442, N331);
xor XOR2 (N1657, N1651, N68);
nand NAND2 (N1658, N1638, N1262);
or OR3 (N1659, N1647, N333, N2);
and AND4 (N1660, N1652, N1232, N743, N794);
and AND3 (N1661, N1650, N466, N656);
not NOT1 (N1662, N1624);
xor XOR2 (N1663, N1657, N1578);
buf BUF1 (N1664, N1646);
xor XOR2 (N1665, N1660, N721);
nand NAND4 (N1666, N1663, N659, N162, N1308);
xor XOR2 (N1667, N1664, N1133);
nand NAND3 (N1668, N1662, N186, N35);
and AND4 (N1669, N1641, N911, N437, N1541);
nand NAND3 (N1670, N1669, N490, N1640);
not NOT1 (N1671, N1668);
not NOT1 (N1672, N1667);
not NOT1 (N1673, N1665);
xor XOR2 (N1674, N1671, N1293);
not NOT1 (N1675, N1673);
and AND3 (N1676, N1666, N264, N1574);
nor NOR2 (N1677, N1654, N586);
or OR3 (N1678, N1674, N1515, N779);
or OR3 (N1679, N1656, N632, N1602);
buf BUF1 (N1680, N1677);
nor NOR3 (N1681, N1678, N23, N402);
xor XOR2 (N1682, N1672, N1510);
xor XOR2 (N1683, N1681, N790);
xor XOR2 (N1684, N1682, N476);
nand NAND4 (N1685, N1661, N391, N576, N981);
buf BUF1 (N1686, N1675);
xor XOR2 (N1687, N1685, N1279);
xor XOR2 (N1688, N1676, N1553);
not NOT1 (N1689, N1687);
nor NOR3 (N1690, N1670, N1286, N648);
not NOT1 (N1691, N1689);
buf BUF1 (N1692, N1658);
nor NOR4 (N1693, N1686, N964, N591, N1647);
nor NOR3 (N1694, N1691, N845, N756);
nor NOR4 (N1695, N1694, N726, N1494, N196);
nor NOR4 (N1696, N1679, N791, N1378, N445);
buf BUF1 (N1697, N1680);
xor XOR2 (N1698, N1695, N985);
not NOT1 (N1699, N1688);
or OR2 (N1700, N1692, N1382);
nor NOR4 (N1701, N1699, N1362, N1270, N415);
nor NOR2 (N1702, N1701, N203);
and AND3 (N1703, N1700, N933, N1465);
xor XOR2 (N1704, N1693, N1682);
nor NOR4 (N1705, N1690, N83, N67, N1615);
not NOT1 (N1706, N1703);
or OR4 (N1707, N1705, N1472, N311, N1692);
xor XOR2 (N1708, N1696, N125);
xor XOR2 (N1709, N1697, N65);
or OR3 (N1710, N1702, N675, N697);
buf BUF1 (N1711, N1683);
or OR3 (N1712, N1706, N505, N1132);
buf BUF1 (N1713, N1707);
nand NAND3 (N1714, N1710, N1604, N222);
and AND4 (N1715, N1708, N303, N584, N1497);
or OR2 (N1716, N1659, N1679);
not NOT1 (N1717, N1704);
buf BUF1 (N1718, N1715);
and AND2 (N1719, N1711, N1365);
xor XOR2 (N1720, N1716, N1605);
or OR4 (N1721, N1709, N1217, N531, N1271);
nand NAND4 (N1722, N1712, N336, N648, N23);
xor XOR2 (N1723, N1698, N1557);
nand NAND4 (N1724, N1714, N1375, N1496, N222);
buf BUF1 (N1725, N1720);
or OR4 (N1726, N1713, N14, N738, N1063);
not NOT1 (N1727, N1726);
or OR3 (N1728, N1717, N433, N652);
buf BUF1 (N1729, N1724);
or OR4 (N1730, N1728, N1325, N855, N1412);
not NOT1 (N1731, N1719);
nand NAND2 (N1732, N1723, N323);
or OR4 (N1733, N1732, N1059, N1026, N668);
and AND3 (N1734, N1729, N738, N1244);
and AND4 (N1735, N1727, N1020, N757, N729);
xor XOR2 (N1736, N1733, N801);
and AND2 (N1737, N1735, N807);
buf BUF1 (N1738, N1725);
and AND4 (N1739, N1734, N1700, N472, N1655);
or OR2 (N1740, N1722, N1360);
and AND2 (N1741, N1730, N729);
and AND4 (N1742, N1718, N387, N1277, N679);
not NOT1 (N1743, N1721);
nor NOR4 (N1744, N1738, N683, N829, N1642);
and AND2 (N1745, N1742, N1586);
nor NOR4 (N1746, N1731, N1041, N832, N1697);
and AND4 (N1747, N1736, N1255, N1139, N1186);
xor XOR2 (N1748, N1744, N1040);
nor NOR2 (N1749, N1741, N118);
or OR3 (N1750, N1740, N665, N747);
and AND2 (N1751, N1739, N1572);
nor NOR2 (N1752, N1750, N278);
nor NOR2 (N1753, N1737, N1067);
and AND2 (N1754, N1746, N534);
and AND4 (N1755, N1749, N23, N263, N76);
nand NAND2 (N1756, N1755, N36);
and AND3 (N1757, N1748, N1476, N570);
nand NAND4 (N1758, N1743, N201, N1333, N1394);
nand NAND2 (N1759, N1754, N869);
and AND3 (N1760, N1752, N1442, N4);
xor XOR2 (N1761, N1747, N150);
buf BUF1 (N1762, N1758);
not NOT1 (N1763, N1762);
or OR2 (N1764, N1761, N383);
xor XOR2 (N1765, N1753, N945);
not NOT1 (N1766, N1760);
or OR2 (N1767, N1764, N1310);
nand NAND3 (N1768, N1765, N627, N1261);
buf BUF1 (N1769, N1757);
buf BUF1 (N1770, N1751);
not NOT1 (N1771, N1763);
and AND3 (N1772, N1770, N638, N357);
buf BUF1 (N1773, N1766);
xor XOR2 (N1774, N1771, N1389);
xor XOR2 (N1775, N1745, N597);
buf BUF1 (N1776, N1773);
nor NOR4 (N1777, N1776, N561, N330, N570);
nor NOR2 (N1778, N1775, N582);
buf BUF1 (N1779, N1684);
not NOT1 (N1780, N1779);
buf BUF1 (N1781, N1769);
nor NOR2 (N1782, N1759, N40);
xor XOR2 (N1783, N1756, N1613);
nor NOR2 (N1784, N1778, N669);
and AND4 (N1785, N1767, N86, N773, N190);
nand NAND4 (N1786, N1774, N695, N1541, N1210);
not NOT1 (N1787, N1786);
and AND3 (N1788, N1787, N27, N203);
nand NAND4 (N1789, N1782, N268, N100, N1182);
not NOT1 (N1790, N1788);
nor NOR2 (N1791, N1789, N458);
nand NAND4 (N1792, N1777, N146, N1572, N226);
nor NOR4 (N1793, N1790, N1088, N303, N781);
not NOT1 (N1794, N1791);
and AND4 (N1795, N1781, N759, N547, N982);
nand NAND3 (N1796, N1768, N1273, N1456);
xor XOR2 (N1797, N1793, N688);
nand NAND3 (N1798, N1794, N828, N1185);
not NOT1 (N1799, N1783);
not NOT1 (N1800, N1792);
buf BUF1 (N1801, N1795);
nor NOR3 (N1802, N1784, N1590, N399);
buf BUF1 (N1803, N1780);
xor XOR2 (N1804, N1802, N1581);
or OR4 (N1805, N1772, N381, N1484, N1245);
not NOT1 (N1806, N1785);
nor NOR4 (N1807, N1800, N1005, N1032, N1386);
nand NAND2 (N1808, N1798, N218);
xor XOR2 (N1809, N1807, N775);
nor NOR2 (N1810, N1801, N668);
buf BUF1 (N1811, N1796);
not NOT1 (N1812, N1811);
nand NAND3 (N1813, N1804, N283, N522);
and AND4 (N1814, N1805, N415, N55, N524);
xor XOR2 (N1815, N1814, N1340);
nand NAND3 (N1816, N1799, N208, N715);
not NOT1 (N1817, N1810);
or OR4 (N1818, N1813, N1786, N1108, N169);
and AND3 (N1819, N1803, N482, N1176);
nand NAND3 (N1820, N1816, N701, N156);
buf BUF1 (N1821, N1809);
xor XOR2 (N1822, N1815, N1170);
nor NOR3 (N1823, N1806, N326, N328);
or OR3 (N1824, N1808, N1656, N1558);
or OR2 (N1825, N1823, N96);
nand NAND4 (N1826, N1819, N20, N119, N558);
buf BUF1 (N1827, N1821);
and AND4 (N1828, N1825, N1216, N6, N212);
buf BUF1 (N1829, N1826);
xor XOR2 (N1830, N1828, N1372);
nand NAND2 (N1831, N1797, N1519);
and AND4 (N1832, N1829, N1649, N512, N1397);
nand NAND4 (N1833, N1817, N1533, N1451, N1092);
nand NAND3 (N1834, N1822, N1335, N771);
not NOT1 (N1835, N1824);
or OR2 (N1836, N1831, N297);
buf BUF1 (N1837, N1832);
nand NAND2 (N1838, N1837, N1003);
buf BUF1 (N1839, N1836);
not NOT1 (N1840, N1835);
buf BUF1 (N1841, N1838);
not NOT1 (N1842, N1834);
xor XOR2 (N1843, N1839, N538);
or OR2 (N1844, N1842, N1217);
not NOT1 (N1845, N1841);
not NOT1 (N1846, N1843);
nor NOR3 (N1847, N1820, N787, N861);
not NOT1 (N1848, N1840);
buf BUF1 (N1849, N1812);
nand NAND3 (N1850, N1848, N889, N1688);
not NOT1 (N1851, N1846);
or OR3 (N1852, N1827, N683, N586);
and AND3 (N1853, N1830, N253, N1704);
xor XOR2 (N1854, N1850, N279);
xor XOR2 (N1855, N1849, N1598);
nand NAND4 (N1856, N1852, N717, N1594, N937);
or OR4 (N1857, N1853, N699, N1263, N546);
or OR3 (N1858, N1856, N1002, N1053);
nor NOR2 (N1859, N1857, N106);
nand NAND2 (N1860, N1845, N1726);
xor XOR2 (N1861, N1818, N1387);
xor XOR2 (N1862, N1861, N1331);
xor XOR2 (N1863, N1851, N254);
xor XOR2 (N1864, N1863, N1709);
or OR2 (N1865, N1844, N938);
nor NOR2 (N1866, N1864, N453);
not NOT1 (N1867, N1833);
buf BUF1 (N1868, N1865);
nand NAND3 (N1869, N1862, N1158, N559);
nand NAND2 (N1870, N1868, N1866);
and AND3 (N1871, N274, N1031, N434);
or OR4 (N1872, N1858, N674, N549, N1215);
or OR4 (N1873, N1854, N1439, N1833, N822);
not NOT1 (N1874, N1855);
xor XOR2 (N1875, N1867, N818);
buf BUF1 (N1876, N1869);
buf BUF1 (N1877, N1871);
buf BUF1 (N1878, N1875);
xor XOR2 (N1879, N1859, N165);
buf BUF1 (N1880, N1872);
buf BUF1 (N1881, N1878);
and AND3 (N1882, N1873, N456, N1055);
not NOT1 (N1883, N1876);
xor XOR2 (N1884, N1880, N6);
xor XOR2 (N1885, N1874, N1560);
buf BUF1 (N1886, N1883);
xor XOR2 (N1887, N1882, N420);
nand NAND2 (N1888, N1860, N442);
not NOT1 (N1889, N1877);
nand NAND2 (N1890, N1886, N1041);
buf BUF1 (N1891, N1879);
nor NOR3 (N1892, N1847, N1691, N46);
or OR4 (N1893, N1888, N93, N1683, N241);
buf BUF1 (N1894, N1881);
buf BUF1 (N1895, N1893);
xor XOR2 (N1896, N1894, N1139);
not NOT1 (N1897, N1896);
not NOT1 (N1898, N1890);
buf BUF1 (N1899, N1885);
and AND3 (N1900, N1870, N707, N1114);
or OR3 (N1901, N1895, N1743, N1664);
xor XOR2 (N1902, N1897, N1827);
not NOT1 (N1903, N1898);
and AND4 (N1904, N1887, N348, N688, N1242);
buf BUF1 (N1905, N1889);
nor NOR4 (N1906, N1899, N1782, N1074, N914);
buf BUF1 (N1907, N1891);
buf BUF1 (N1908, N1884);
or OR2 (N1909, N1907, N1835);
not NOT1 (N1910, N1901);
nor NOR4 (N1911, N1909, N1729, N1557, N24);
or OR3 (N1912, N1911, N1476, N1272);
and AND3 (N1913, N1903, N1818, N1121);
xor XOR2 (N1914, N1902, N421);
and AND3 (N1915, N1892, N1066, N564);
xor XOR2 (N1916, N1910, N730);
nand NAND4 (N1917, N1908, N422, N1719, N1228);
not NOT1 (N1918, N1915);
nor NOR3 (N1919, N1917, N710, N793);
and AND3 (N1920, N1913, N988, N912);
not NOT1 (N1921, N1912);
not NOT1 (N1922, N1916);
or OR2 (N1923, N1906, N55);
nor NOR3 (N1924, N1923, N412, N793);
xor XOR2 (N1925, N1905, N818);
nand NAND3 (N1926, N1900, N421, N592);
nor NOR4 (N1927, N1925, N1835, N1493, N1897);
or OR2 (N1928, N1918, N38);
buf BUF1 (N1929, N1904);
not NOT1 (N1930, N1929);
xor XOR2 (N1931, N1926, N1633);
or OR3 (N1932, N1930, N1083, N1804);
nor NOR4 (N1933, N1928, N662, N797, N559);
not NOT1 (N1934, N1932);
not NOT1 (N1935, N1920);
buf BUF1 (N1936, N1914);
and AND2 (N1937, N1919, N720);
or OR2 (N1938, N1924, N230);
nand NAND3 (N1939, N1931, N1890, N1485);
not NOT1 (N1940, N1934);
nor NOR2 (N1941, N1938, N512);
or OR4 (N1942, N1921, N949, N600, N712);
buf BUF1 (N1943, N1941);
not NOT1 (N1944, N1942);
or OR3 (N1945, N1927, N1755, N1191);
buf BUF1 (N1946, N1939);
nand NAND2 (N1947, N1945, N531);
xor XOR2 (N1948, N1940, N683);
not NOT1 (N1949, N1946);
nand NAND3 (N1950, N1933, N1846, N865);
and AND3 (N1951, N1947, N43, N1876);
and AND3 (N1952, N1943, N1150, N747);
nor NOR4 (N1953, N1951, N416, N268, N1259);
nor NOR4 (N1954, N1922, N913, N1388, N1839);
and AND3 (N1955, N1950, N1914, N1910);
or OR2 (N1956, N1954, N896);
not NOT1 (N1957, N1935);
and AND3 (N1958, N1949, N935, N91);
buf BUF1 (N1959, N1936);
buf BUF1 (N1960, N1955);
buf BUF1 (N1961, N1952);
buf BUF1 (N1962, N1953);
and AND4 (N1963, N1956, N1167, N1111, N1717);
buf BUF1 (N1964, N1962);
and AND3 (N1965, N1958, N1796, N1308);
or OR4 (N1966, N1957, N140, N495, N288);
nor NOR3 (N1967, N1959, N1722, N1235);
buf BUF1 (N1968, N1944);
not NOT1 (N1969, N1966);
buf BUF1 (N1970, N1967);
buf BUF1 (N1971, N1937);
nand NAND4 (N1972, N1964, N201, N1084, N1588);
or OR4 (N1973, N1963, N1313, N1900, N1600);
or OR3 (N1974, N1948, N1550, N1579);
xor XOR2 (N1975, N1974, N346);
buf BUF1 (N1976, N1965);
not NOT1 (N1977, N1975);
buf BUF1 (N1978, N1961);
nor NOR3 (N1979, N1977, N653, N114);
xor XOR2 (N1980, N1968, N315);
not NOT1 (N1981, N1979);
and AND4 (N1982, N1960, N7, N58, N136);
buf BUF1 (N1983, N1970);
buf BUF1 (N1984, N1981);
xor XOR2 (N1985, N1982, N1920);
nand NAND2 (N1986, N1983, N1171);
and AND4 (N1987, N1969, N681, N119, N1952);
and AND2 (N1988, N1984, N812);
and AND4 (N1989, N1973, N371, N1932, N1605);
buf BUF1 (N1990, N1972);
not NOT1 (N1991, N1989);
nor NOR2 (N1992, N1986, N1802);
buf BUF1 (N1993, N1971);
not NOT1 (N1994, N1980);
xor XOR2 (N1995, N1985, N1713);
not NOT1 (N1996, N1992);
xor XOR2 (N1997, N1994, N1995);
nand NAND2 (N1998, N393, N241);
xor XOR2 (N1999, N1988, N782);
nand NAND3 (N2000, N1993, N209, N1678);
nor NOR2 (N2001, N2000, N1181);
nand NAND3 (N2002, N1987, N787, N610);
not NOT1 (N2003, N1997);
nand NAND2 (N2004, N1996, N267);
nor NOR2 (N2005, N1978, N241);
xor XOR2 (N2006, N1990, N1918);
xor XOR2 (N2007, N1991, N314);
and AND3 (N2008, N1999, N300, N201);
or OR4 (N2009, N2004, N1538, N1866, N253);
buf BUF1 (N2010, N2001);
nor NOR3 (N2011, N1976, N1327, N215);
and AND2 (N2012, N2002, N1617);
or OR2 (N2013, N2009, N1714);
or OR4 (N2014, N2011, N438, N1695, N453);
and AND3 (N2015, N2003, N1693, N1818);
nor NOR4 (N2016, N2005, N1166, N573, N1767);
nand NAND3 (N2017, N2014, N916, N1392);
or OR2 (N2018, N2010, N928);
nand NAND2 (N2019, N2007, N330);
not NOT1 (N2020, N2013);
not NOT1 (N2021, N2015);
or OR3 (N2022, N2016, N1026, N99);
xor XOR2 (N2023, N2022, N1742);
endmodule