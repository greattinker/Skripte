// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20;

output N6418,N6417,N6366,N6397,N6419,N6412,N6408,N6415,N6414,N6420;

nor NOR2 (N21, N6, N13);
nand NAND4 (N22, N1, N6, N4, N3);
not NOT1 (N23, N22);
xor XOR2 (N24, N21, N22);
nand NAND3 (N25, N4, N5, N4);
nand NAND2 (N26, N21, N11);
buf BUF1 (N27, N21);
buf BUF1 (N28, N17);
not NOT1 (N29, N25);
nor NOR3 (N30, N22, N5, N21);
xor XOR2 (N31, N4, N12);
or OR4 (N32, N31, N7, N31, N13);
xor XOR2 (N33, N29, N19);
nor NOR4 (N34, N9, N30, N8, N28);
not NOT1 (N35, N3);
buf BUF1 (N36, N25);
nand NAND4 (N37, N28, N15, N25, N4);
nand NAND2 (N38, N33, N19);
and AND3 (N39, N23, N16, N5);
not NOT1 (N40, N27);
nand NAND3 (N41, N40, N24, N17);
xor XOR2 (N42, N18, N2);
nor NOR2 (N43, N34, N29);
and AND4 (N44, N36, N21, N18, N32);
buf BUF1 (N45, N38);
buf BUF1 (N46, N25);
xor XOR2 (N47, N26, N37);
buf BUF1 (N48, N27);
or OR2 (N49, N35, N41);
not NOT1 (N50, N9);
xor XOR2 (N51, N47, N45);
xor XOR2 (N52, N19, N16);
not NOT1 (N53, N50);
nand NAND3 (N54, N48, N44, N5);
xor XOR2 (N55, N8, N46);
xor XOR2 (N56, N37, N30);
buf BUF1 (N57, N54);
buf BUF1 (N58, N53);
xor XOR2 (N59, N43, N24);
nor NOR4 (N60, N55, N28, N30, N52);
nor NOR3 (N61, N23, N52, N39);
xor XOR2 (N62, N47, N51);
not NOT1 (N63, N6);
not NOT1 (N64, N58);
nor NOR3 (N65, N57, N14, N51);
not NOT1 (N66, N64);
nor NOR3 (N67, N42, N30, N26);
buf BUF1 (N68, N65);
and AND3 (N69, N62, N64, N47);
not NOT1 (N70, N49);
xor XOR2 (N71, N70, N42);
nor NOR3 (N72, N67, N45, N33);
not NOT1 (N73, N59);
or OR4 (N74, N72, N50, N67, N12);
buf BUF1 (N75, N71);
and AND4 (N76, N69, N51, N54, N63);
not NOT1 (N77, N29);
buf BUF1 (N78, N74);
and AND2 (N79, N56, N7);
nand NAND3 (N80, N75, N70, N4);
and AND3 (N81, N66, N63, N49);
and AND2 (N82, N81, N54);
and AND2 (N83, N78, N14);
or OR4 (N84, N79, N39, N15, N73);
nor NOR2 (N85, N81, N61);
nor NOR3 (N86, N84, N20, N62);
nand NAND2 (N87, N16, N45);
and AND2 (N88, N86, N1);
and AND3 (N89, N83, N84, N9);
buf BUF1 (N90, N82);
xor XOR2 (N91, N88, N28);
xor XOR2 (N92, N89, N10);
buf BUF1 (N93, N60);
buf BUF1 (N94, N91);
or OR4 (N95, N92, N37, N92, N37);
buf BUF1 (N96, N94);
not NOT1 (N97, N76);
or OR4 (N98, N96, N89, N60, N91);
nand NAND3 (N99, N98, N64, N37);
not NOT1 (N100, N87);
and AND2 (N101, N77, N35);
or OR2 (N102, N97, N45);
or OR2 (N103, N90, N41);
or OR3 (N104, N95, N7, N90);
not NOT1 (N105, N101);
not NOT1 (N106, N103);
not NOT1 (N107, N105);
xor XOR2 (N108, N68, N107);
or OR3 (N109, N5, N21, N67);
xor XOR2 (N110, N99, N31);
or OR3 (N111, N104, N59, N39);
xor XOR2 (N112, N100, N110);
buf BUF1 (N113, N67);
or OR4 (N114, N106, N91, N84, N74);
or OR3 (N115, N102, N65, N77);
and AND2 (N116, N108, N39);
nor NOR3 (N117, N109, N90, N45);
not NOT1 (N118, N111);
nand NAND4 (N119, N93, N113, N85, N81);
or OR4 (N120, N51, N77, N7, N35);
not NOT1 (N121, N82);
or OR2 (N122, N121, N30);
and AND4 (N123, N112, N10, N92, N120);
xor XOR2 (N124, N84, N53);
not NOT1 (N125, N116);
buf BUF1 (N126, N123);
buf BUF1 (N127, N118);
nand NAND4 (N128, N127, N37, N99, N21);
xor XOR2 (N129, N114, N124);
nand NAND2 (N130, N59, N9);
nand NAND4 (N131, N126, N16, N113, N60);
and AND2 (N132, N115, N5);
xor XOR2 (N133, N129, N80);
and AND3 (N134, N100, N60, N1);
or OR4 (N135, N131, N112, N61, N134);
and AND2 (N136, N83, N101);
and AND4 (N137, N119, N95, N28, N80);
nand NAND2 (N138, N125, N127);
nand NAND3 (N139, N132, N14, N16);
and AND2 (N140, N135, N55);
not NOT1 (N141, N130);
xor XOR2 (N142, N138, N82);
nor NOR3 (N143, N122, N33, N134);
xor XOR2 (N144, N143, N140);
buf BUF1 (N145, N40);
nand NAND3 (N146, N136, N85, N103);
not NOT1 (N147, N137);
or OR2 (N148, N146, N123);
nor NOR4 (N149, N133, N14, N43, N127);
nand NAND4 (N150, N128, N127, N100, N134);
or OR4 (N151, N141, N16, N107, N126);
xor XOR2 (N152, N150, N37);
nand NAND2 (N153, N142, N42);
or OR3 (N154, N149, N107, N48);
nor NOR3 (N155, N152, N14, N78);
or OR3 (N156, N145, N76, N124);
or OR4 (N157, N153, N67, N5, N30);
nor NOR4 (N158, N139, N11, N40, N6);
not NOT1 (N159, N158);
or OR4 (N160, N155, N74, N73, N102);
or OR2 (N161, N157, N81);
or OR2 (N162, N147, N152);
or OR2 (N163, N160, N150);
xor XOR2 (N164, N163, N132);
nand NAND4 (N165, N117, N32, N30, N92);
buf BUF1 (N166, N144);
buf BUF1 (N167, N166);
nand NAND2 (N168, N148, N74);
nor NOR4 (N169, N168, N54, N166, N72);
or OR3 (N170, N164, N25, N134);
xor XOR2 (N171, N165, N117);
nand NAND3 (N172, N161, N65, N98);
buf BUF1 (N173, N159);
and AND3 (N174, N170, N93, N51);
and AND2 (N175, N154, N3);
nand NAND4 (N176, N162, N104, N170, N36);
nor NOR2 (N177, N176, N126);
nand NAND4 (N178, N169, N48, N64, N84);
nor NOR2 (N179, N173, N16);
xor XOR2 (N180, N179, N32);
nor NOR3 (N181, N180, N138, N92);
nand NAND2 (N182, N175, N167);
and AND4 (N183, N179, N10, N68, N135);
xor XOR2 (N184, N178, N181);
buf BUF1 (N185, N17);
buf BUF1 (N186, N171);
nor NOR4 (N187, N172, N49, N136, N31);
buf BUF1 (N188, N177);
buf BUF1 (N189, N151);
xor XOR2 (N190, N189, N12);
not NOT1 (N191, N186);
not NOT1 (N192, N190);
nand NAND2 (N193, N192, N189);
buf BUF1 (N194, N182);
xor XOR2 (N195, N156, N181);
nor NOR4 (N196, N174, N6, N155, N98);
and AND3 (N197, N184, N123, N176);
or OR4 (N198, N188, N173, N159, N8);
or OR2 (N199, N191, N57);
or OR2 (N200, N185, N185);
xor XOR2 (N201, N200, N18);
nor NOR3 (N202, N199, N31, N163);
nor NOR3 (N203, N196, N126, N24);
nor NOR2 (N204, N203, N7);
buf BUF1 (N205, N194);
or OR2 (N206, N195, N2);
or OR2 (N207, N202, N168);
xor XOR2 (N208, N198, N141);
nor NOR2 (N209, N208, N16);
nand NAND4 (N210, N209, N180, N121, N127);
nand NAND2 (N211, N197, N21);
xor XOR2 (N212, N193, N209);
nand NAND4 (N213, N212, N197, N3, N81);
nand NAND3 (N214, N211, N47, N146);
buf BUF1 (N215, N207);
nand NAND4 (N216, N205, N194, N115, N211);
not NOT1 (N217, N187);
or OR3 (N218, N183, N112, N9);
buf BUF1 (N219, N210);
and AND2 (N220, N206, N163);
or OR4 (N221, N213, N119, N71, N1);
nor NOR2 (N222, N219, N27);
nand NAND4 (N223, N222, N136, N148, N53);
xor XOR2 (N224, N223, N209);
or OR3 (N225, N221, N203, N214);
not NOT1 (N226, N199);
or OR3 (N227, N201, N186, N5);
nor NOR4 (N228, N224, N110, N165, N97);
nor NOR2 (N229, N227, N162);
nand NAND3 (N230, N228, N84, N177);
nand NAND3 (N231, N226, N75, N130);
nor NOR3 (N232, N218, N88, N218);
and AND2 (N233, N217, N178);
and AND4 (N234, N220, N60, N8, N74);
nor NOR3 (N235, N232, N42, N19);
and AND3 (N236, N235, N230, N8);
nor NOR4 (N237, N102, N184, N216, N187);
nand NAND2 (N238, N40, N41);
and AND2 (N239, N204, N175);
xor XOR2 (N240, N233, N108);
not NOT1 (N241, N234);
not NOT1 (N242, N231);
not NOT1 (N243, N241);
nor NOR2 (N244, N236, N165);
xor XOR2 (N245, N240, N41);
buf BUF1 (N246, N244);
xor XOR2 (N247, N225, N47);
nand NAND4 (N248, N242, N107, N177, N35);
buf BUF1 (N249, N238);
buf BUF1 (N250, N229);
xor XOR2 (N251, N247, N235);
buf BUF1 (N252, N249);
buf BUF1 (N253, N250);
or OR2 (N254, N237, N170);
xor XOR2 (N255, N243, N150);
and AND3 (N256, N239, N22, N180);
and AND2 (N257, N251, N68);
buf BUF1 (N258, N215);
xor XOR2 (N259, N255, N17);
or OR2 (N260, N252, N247);
not NOT1 (N261, N259);
not NOT1 (N262, N246);
buf BUF1 (N263, N256);
xor XOR2 (N264, N263, N219);
nor NOR2 (N265, N245, N195);
or OR3 (N266, N260, N245, N174);
not NOT1 (N267, N266);
not NOT1 (N268, N248);
or OR4 (N269, N265, N263, N81, N199);
nand NAND4 (N270, N269, N241, N262, N248);
not NOT1 (N271, N213);
xor XOR2 (N272, N267, N177);
nand NAND2 (N273, N271, N104);
xor XOR2 (N274, N257, N167);
xor XOR2 (N275, N274, N85);
buf BUF1 (N276, N261);
and AND2 (N277, N254, N93);
xor XOR2 (N278, N276, N127);
xor XOR2 (N279, N278, N276);
and AND4 (N280, N273, N123, N156, N264);
nor NOR3 (N281, N256, N72, N86);
nor NOR2 (N282, N270, N17);
nand NAND3 (N283, N272, N92, N255);
buf BUF1 (N284, N279);
nand NAND3 (N285, N282, N65, N81);
xor XOR2 (N286, N277, N154);
nand NAND4 (N287, N284, N150, N6, N116);
not NOT1 (N288, N268);
and AND3 (N289, N281, N186, N215);
nor NOR4 (N290, N280, N253, N159, N200);
nor NOR3 (N291, N285, N92, N119);
buf BUF1 (N292, N41);
buf BUF1 (N293, N287);
xor XOR2 (N294, N293, N7);
and AND3 (N295, N289, N127, N126);
and AND3 (N296, N258, N168, N192);
and AND3 (N297, N290, N144, N229);
nor NOR4 (N298, N292, N190, N182, N279);
nand NAND2 (N299, N296, N101);
not NOT1 (N300, N298);
not NOT1 (N301, N275);
xor XOR2 (N302, N300, N227);
nand NAND4 (N303, N299, N250, N138, N241);
xor XOR2 (N304, N297, N176);
nor NOR4 (N305, N283, N243, N99, N88);
or OR3 (N306, N291, N34, N195);
not NOT1 (N307, N305);
nor NOR3 (N308, N286, N35, N42);
and AND2 (N309, N304, N269);
and AND4 (N310, N302, N217, N109, N95);
buf BUF1 (N311, N294);
and AND3 (N312, N307, N274, N103);
nand NAND2 (N313, N306, N206);
buf BUF1 (N314, N312);
xor XOR2 (N315, N313, N42);
not NOT1 (N316, N314);
buf BUF1 (N317, N303);
xor XOR2 (N318, N309, N24);
not NOT1 (N319, N308);
xor XOR2 (N320, N311, N272);
or OR4 (N321, N319, N83, N301, N153);
buf BUF1 (N322, N193);
nor NOR3 (N323, N320, N280, N227);
nand NAND4 (N324, N310, N135, N323, N26);
buf BUF1 (N325, N274);
nor NOR2 (N326, N325, N3);
buf BUF1 (N327, N317);
buf BUF1 (N328, N318);
and AND4 (N329, N324, N125, N129, N109);
not NOT1 (N330, N288);
nor NOR3 (N331, N321, N28, N282);
xor XOR2 (N332, N330, N296);
or OR2 (N333, N329, N317);
or OR4 (N334, N328, N168, N149, N291);
and AND2 (N335, N334, N265);
and AND2 (N336, N335, N320);
buf BUF1 (N337, N327);
and AND3 (N338, N295, N48, N104);
nor NOR3 (N339, N315, N260, N56);
nand NAND3 (N340, N322, N31, N191);
nand NAND4 (N341, N336, N253, N267, N147);
xor XOR2 (N342, N333, N38);
xor XOR2 (N343, N332, N57);
nor NOR3 (N344, N341, N305, N334);
buf BUF1 (N345, N343);
nand NAND4 (N346, N326, N330, N251, N232);
xor XOR2 (N347, N337, N316);
nor NOR2 (N348, N31, N239);
buf BUF1 (N349, N342);
buf BUF1 (N350, N349);
buf BUF1 (N351, N331);
and AND2 (N352, N346, N16);
or OR2 (N353, N350, N340);
or OR2 (N354, N237, N73);
not NOT1 (N355, N353);
xor XOR2 (N356, N348, N103);
buf BUF1 (N357, N352);
or OR4 (N358, N338, N278, N92, N286);
or OR2 (N359, N351, N169);
nand NAND2 (N360, N358, N270);
or OR2 (N361, N359, N154);
or OR4 (N362, N345, N261, N38, N83);
and AND2 (N363, N347, N96);
not NOT1 (N364, N361);
not NOT1 (N365, N355);
or OR3 (N366, N365, N10, N37);
and AND2 (N367, N360, N121);
and AND3 (N368, N362, N154, N21);
not NOT1 (N369, N368);
nor NOR2 (N370, N366, N149);
nand NAND3 (N371, N367, N214, N194);
buf BUF1 (N372, N356);
xor XOR2 (N373, N364, N25);
nand NAND4 (N374, N373, N179, N15, N272);
nand NAND3 (N375, N363, N209, N216);
nand NAND2 (N376, N370, N4);
not NOT1 (N377, N372);
xor XOR2 (N378, N344, N279);
not NOT1 (N379, N339);
or OR4 (N380, N379, N219, N330, N367);
nand NAND3 (N381, N354, N10, N313);
not NOT1 (N382, N375);
buf BUF1 (N383, N378);
nor NOR4 (N384, N382, N209, N268, N73);
xor XOR2 (N385, N380, N1);
buf BUF1 (N386, N371);
nor NOR4 (N387, N384, N41, N7, N334);
and AND4 (N388, N381, N349, N211, N148);
buf BUF1 (N389, N387);
and AND4 (N390, N376, N291, N177, N40);
buf BUF1 (N391, N389);
xor XOR2 (N392, N357, N344);
or OR3 (N393, N369, N171, N155);
nand NAND3 (N394, N383, N192, N87);
buf BUF1 (N395, N391);
not NOT1 (N396, N388);
nor NOR2 (N397, N385, N185);
nor NOR3 (N398, N397, N129, N6);
not NOT1 (N399, N398);
nor NOR2 (N400, N374, N390);
xor XOR2 (N401, N365, N208);
xor XOR2 (N402, N395, N105);
buf BUF1 (N403, N392);
xor XOR2 (N404, N400, N398);
xor XOR2 (N405, N404, N131);
not NOT1 (N406, N402);
and AND4 (N407, N406, N387, N271, N65);
buf BUF1 (N408, N407);
nand NAND4 (N409, N401, N202, N119, N74);
nand NAND4 (N410, N396, N268, N281, N243);
nor NOR3 (N411, N377, N155, N253);
buf BUF1 (N412, N399);
xor XOR2 (N413, N410, N85);
nor NOR4 (N414, N393, N225, N319, N37);
and AND3 (N415, N411, N249, N362);
and AND4 (N416, N405, N229, N176, N70);
not NOT1 (N417, N409);
nor NOR2 (N418, N413, N259);
nor NOR4 (N419, N403, N356, N208, N303);
or OR4 (N420, N414, N326, N63, N230);
or OR3 (N421, N412, N112, N284);
or OR4 (N422, N420, N238, N116, N203);
nand NAND4 (N423, N416, N391, N208, N37);
xor XOR2 (N424, N419, N307);
and AND3 (N425, N424, N184, N28);
and AND2 (N426, N418, N395);
not NOT1 (N427, N422);
xor XOR2 (N428, N427, N119);
or OR3 (N429, N417, N158, N2);
or OR3 (N430, N429, N397, N209);
and AND2 (N431, N415, N122);
nand NAND4 (N432, N408, N274, N241, N175);
buf BUF1 (N433, N426);
or OR2 (N434, N394, N412);
and AND3 (N435, N433, N369, N327);
nand NAND3 (N436, N421, N112, N15);
xor XOR2 (N437, N430, N261);
xor XOR2 (N438, N432, N67);
nand NAND3 (N439, N436, N56, N154);
and AND3 (N440, N437, N53, N373);
and AND4 (N441, N386, N424, N227, N387);
xor XOR2 (N442, N431, N439);
buf BUF1 (N443, N71);
and AND4 (N444, N443, N184, N317, N331);
nor NOR3 (N445, N428, N319, N29);
nor NOR2 (N446, N440, N56);
or OR2 (N447, N425, N124);
buf BUF1 (N448, N423);
not NOT1 (N449, N441);
not NOT1 (N450, N445);
xor XOR2 (N451, N435, N16);
not NOT1 (N452, N450);
not NOT1 (N453, N447);
buf BUF1 (N454, N444);
and AND2 (N455, N442, N200);
nor NOR4 (N456, N448, N246, N364, N68);
not NOT1 (N457, N438);
and AND2 (N458, N457, N457);
xor XOR2 (N459, N451, N119);
and AND4 (N460, N434, N45, N188, N250);
and AND4 (N461, N460, N447, N360, N248);
nor NOR3 (N462, N461, N128, N355);
and AND3 (N463, N446, N441, N92);
buf BUF1 (N464, N455);
xor XOR2 (N465, N456, N195);
xor XOR2 (N466, N464, N354);
xor XOR2 (N467, N459, N37);
nor NOR2 (N468, N463, N441);
xor XOR2 (N469, N449, N342);
xor XOR2 (N470, N469, N230);
not NOT1 (N471, N467);
xor XOR2 (N472, N458, N129);
or OR4 (N473, N472, N467, N252, N173);
nand NAND2 (N474, N465, N218);
buf BUF1 (N475, N454);
nor NOR3 (N476, N466, N252, N439);
buf BUF1 (N477, N468);
xor XOR2 (N478, N477, N119);
nor NOR4 (N479, N474, N313, N337, N328);
xor XOR2 (N480, N475, N72);
nor NOR2 (N481, N453, N362);
not NOT1 (N482, N480);
nor NOR4 (N483, N462, N1, N25, N479);
nand NAND3 (N484, N400, N267, N283);
xor XOR2 (N485, N452, N240);
nor NOR4 (N486, N484, N49, N50, N114);
nand NAND4 (N487, N473, N239, N307, N73);
or OR4 (N488, N478, N364, N414, N310);
or OR4 (N489, N482, N205, N172, N329);
not NOT1 (N490, N483);
nand NAND2 (N491, N470, N74);
xor XOR2 (N492, N490, N19);
buf BUF1 (N493, N491);
or OR3 (N494, N476, N485, N181);
buf BUF1 (N495, N185);
buf BUF1 (N496, N492);
xor XOR2 (N497, N493, N217);
or OR2 (N498, N494, N177);
xor XOR2 (N499, N486, N282);
xor XOR2 (N500, N488, N338);
xor XOR2 (N501, N471, N308);
or OR2 (N502, N499, N307);
nor NOR2 (N503, N481, N448);
or OR2 (N504, N487, N433);
or OR3 (N505, N504, N43, N264);
xor XOR2 (N506, N501, N331);
or OR2 (N507, N505, N427);
xor XOR2 (N508, N506, N383);
not NOT1 (N509, N495);
nor NOR2 (N510, N489, N194);
nand NAND2 (N511, N503, N49);
or OR4 (N512, N500, N425, N481, N269);
nand NAND3 (N513, N498, N330, N110);
xor XOR2 (N514, N497, N156);
nand NAND3 (N515, N509, N319, N274);
or OR3 (N516, N512, N177, N322);
nor NOR3 (N517, N516, N239, N458);
buf BUF1 (N518, N510);
buf BUF1 (N519, N496);
buf BUF1 (N520, N518);
nand NAND2 (N521, N508, N29);
buf BUF1 (N522, N507);
buf BUF1 (N523, N519);
not NOT1 (N524, N511);
nand NAND3 (N525, N523, N92, N148);
and AND2 (N526, N520, N216);
not NOT1 (N527, N526);
nor NOR4 (N528, N517, N147, N386, N207);
xor XOR2 (N529, N515, N289);
buf BUF1 (N530, N513);
and AND3 (N531, N522, N135, N163);
buf BUF1 (N532, N524);
xor XOR2 (N533, N514, N347);
nor NOR4 (N534, N531, N504, N503, N47);
not NOT1 (N535, N525);
or OR2 (N536, N535, N334);
xor XOR2 (N537, N530, N475);
not NOT1 (N538, N533);
or OR3 (N539, N521, N110, N398);
and AND4 (N540, N534, N519, N359, N387);
and AND3 (N541, N532, N332, N538);
nand NAND4 (N542, N254, N93, N352, N186);
buf BUF1 (N543, N540);
nand NAND4 (N544, N502, N185, N483, N167);
and AND4 (N545, N529, N462, N113, N220);
nor NOR2 (N546, N541, N440);
not NOT1 (N547, N527);
buf BUF1 (N548, N539);
buf BUF1 (N549, N543);
and AND2 (N550, N547, N257);
or OR3 (N551, N536, N99, N450);
or OR3 (N552, N537, N428, N469);
or OR4 (N553, N548, N536, N387, N391);
not NOT1 (N554, N544);
nand NAND3 (N555, N553, N5, N366);
buf BUF1 (N556, N545);
not NOT1 (N557, N528);
xor XOR2 (N558, N557, N50);
and AND3 (N559, N552, N68, N175);
nor NOR3 (N560, N551, N226, N386);
not NOT1 (N561, N558);
and AND3 (N562, N546, N157, N51);
and AND4 (N563, N555, N309, N91, N492);
nand NAND2 (N564, N560, N518);
not NOT1 (N565, N549);
buf BUF1 (N566, N564);
or OR3 (N567, N550, N66, N19);
or OR4 (N568, N565, N263, N130, N221);
buf BUF1 (N569, N561);
xor XOR2 (N570, N559, N213);
nand NAND4 (N571, N554, N291, N100, N9);
not NOT1 (N572, N563);
buf BUF1 (N573, N566);
buf BUF1 (N574, N567);
nor NOR3 (N575, N572, N521, N401);
nand NAND4 (N576, N571, N72, N80, N379);
xor XOR2 (N577, N562, N534);
not NOT1 (N578, N569);
not NOT1 (N579, N577);
nand NAND4 (N580, N576, N106, N224, N317);
nand NAND2 (N581, N556, N145);
or OR2 (N582, N578, N477);
or OR2 (N583, N574, N165);
or OR3 (N584, N583, N525, N130);
or OR2 (N585, N579, N288);
buf BUF1 (N586, N585);
nand NAND3 (N587, N573, N250, N20);
nor NOR2 (N588, N575, N489);
nand NAND4 (N589, N580, N551, N323, N21);
nand NAND2 (N590, N570, N85);
buf BUF1 (N591, N590);
and AND2 (N592, N584, N585);
xor XOR2 (N593, N568, N277);
or OR3 (N594, N589, N133, N521);
xor XOR2 (N595, N581, N62);
buf BUF1 (N596, N595);
xor XOR2 (N597, N587, N447);
xor XOR2 (N598, N582, N290);
xor XOR2 (N599, N597, N56);
and AND4 (N600, N594, N118, N295, N452);
nand NAND3 (N601, N598, N328, N299);
xor XOR2 (N602, N593, N59);
buf BUF1 (N603, N592);
not NOT1 (N604, N601);
nand NAND2 (N605, N602, N550);
buf BUF1 (N606, N603);
nand NAND3 (N607, N605, N568, N402);
and AND4 (N608, N586, N258, N237, N95);
not NOT1 (N609, N599);
and AND2 (N610, N606, N253);
and AND3 (N611, N600, N417, N514);
and AND4 (N612, N611, N273, N598, N362);
xor XOR2 (N613, N591, N456);
nor NOR3 (N614, N610, N581, N508);
nand NAND2 (N615, N612, N248);
not NOT1 (N616, N609);
and AND3 (N617, N607, N125, N258);
and AND3 (N618, N604, N65, N191);
and AND4 (N619, N608, N294, N172, N170);
nor NOR3 (N620, N613, N335, N545);
or OR3 (N621, N619, N207, N530);
nor NOR4 (N622, N616, N607, N613, N47);
xor XOR2 (N623, N621, N57);
buf BUF1 (N624, N618);
buf BUF1 (N625, N588);
xor XOR2 (N626, N615, N433);
and AND3 (N627, N625, N532, N511);
buf BUF1 (N628, N626);
and AND2 (N629, N628, N240);
nand NAND3 (N630, N627, N474, N49);
nand NAND3 (N631, N630, N591, N387);
not NOT1 (N632, N614);
xor XOR2 (N633, N629, N305);
or OR2 (N634, N617, N55);
buf BUF1 (N635, N632);
or OR2 (N636, N622, N286);
not NOT1 (N637, N636);
buf BUF1 (N638, N620);
not NOT1 (N639, N637);
and AND3 (N640, N623, N52, N135);
nor NOR2 (N641, N596, N283);
xor XOR2 (N642, N633, N601);
xor XOR2 (N643, N639, N411);
nand NAND2 (N644, N638, N226);
xor XOR2 (N645, N631, N530);
or OR4 (N646, N641, N414, N153, N516);
xor XOR2 (N647, N643, N118);
buf BUF1 (N648, N645);
nand NAND2 (N649, N624, N359);
and AND2 (N650, N647, N323);
nor NOR4 (N651, N650, N193, N359, N323);
nor NOR4 (N652, N644, N275, N439, N513);
not NOT1 (N653, N648);
buf BUF1 (N654, N642);
and AND3 (N655, N640, N433, N252);
xor XOR2 (N656, N655, N647);
nand NAND3 (N657, N653, N304, N69);
or OR4 (N658, N651, N237, N398, N207);
buf BUF1 (N659, N652);
xor XOR2 (N660, N657, N308);
or OR3 (N661, N649, N40, N151);
xor XOR2 (N662, N634, N544);
buf BUF1 (N663, N662);
nor NOR2 (N664, N635, N576);
and AND3 (N665, N663, N165, N203);
xor XOR2 (N666, N664, N518);
and AND2 (N667, N666, N40);
nand NAND4 (N668, N542, N431, N613, N423);
nor NOR2 (N669, N665, N321);
or OR3 (N670, N656, N467, N132);
not NOT1 (N671, N658);
xor XOR2 (N672, N670, N63);
or OR3 (N673, N646, N119, N371);
and AND2 (N674, N671, N17);
nand NAND3 (N675, N654, N534, N110);
or OR4 (N676, N659, N277, N20, N358);
nor NOR3 (N677, N668, N81, N7);
not NOT1 (N678, N673);
and AND4 (N679, N661, N319, N473, N453);
nor NOR3 (N680, N674, N515, N406);
buf BUF1 (N681, N678);
nand NAND2 (N682, N680, N466);
nand NAND2 (N683, N660, N564);
and AND2 (N684, N675, N432);
nor NOR3 (N685, N667, N609, N316);
not NOT1 (N686, N681);
buf BUF1 (N687, N686);
nand NAND4 (N688, N687, N194, N499, N29);
nor NOR2 (N689, N688, N145);
and AND2 (N690, N677, N25);
nand NAND3 (N691, N679, N343, N353);
buf BUF1 (N692, N689);
buf BUF1 (N693, N683);
buf BUF1 (N694, N691);
and AND4 (N695, N682, N358, N444, N27);
nor NOR3 (N696, N693, N421, N653);
nor NOR2 (N697, N694, N56);
xor XOR2 (N698, N697, N50);
or OR4 (N699, N669, N225, N331, N382);
buf BUF1 (N700, N699);
and AND4 (N701, N695, N213, N137, N25);
nor NOR2 (N702, N701, N42);
buf BUF1 (N703, N685);
xor XOR2 (N704, N703, N661);
and AND4 (N705, N690, N254, N84, N638);
not NOT1 (N706, N672);
nor NOR3 (N707, N676, N431, N193);
and AND4 (N708, N706, N462, N513, N671);
buf BUF1 (N709, N707);
nand NAND3 (N710, N684, N151, N678);
buf BUF1 (N711, N700);
not NOT1 (N712, N711);
and AND4 (N713, N708, N524, N278, N200);
or OR3 (N714, N698, N120, N362);
xor XOR2 (N715, N704, N693);
and AND3 (N716, N709, N94, N24);
buf BUF1 (N717, N705);
nand NAND2 (N718, N713, N597);
nor NOR4 (N719, N712, N97, N57, N391);
nor NOR3 (N720, N714, N333, N674);
buf BUF1 (N721, N710);
nand NAND3 (N722, N716, N258, N153);
not NOT1 (N723, N722);
buf BUF1 (N724, N720);
nand NAND3 (N725, N717, N565, N504);
and AND2 (N726, N702, N63);
or OR4 (N727, N723, N64, N491, N508);
or OR2 (N728, N692, N476);
nand NAND3 (N729, N696, N548, N255);
xor XOR2 (N730, N715, N55);
and AND3 (N731, N721, N439, N80);
or OR3 (N732, N730, N578, N345);
nand NAND3 (N733, N727, N564, N632);
not NOT1 (N734, N732);
nor NOR2 (N735, N729, N7);
nor NOR2 (N736, N725, N599);
and AND4 (N737, N726, N648, N475, N57);
nand NAND4 (N738, N718, N637, N712, N443);
nor NOR2 (N739, N734, N646);
or OR2 (N740, N733, N643);
nand NAND4 (N741, N738, N349, N66, N358);
or OR4 (N742, N731, N609, N428, N729);
or OR4 (N743, N739, N428, N365, N310);
not NOT1 (N744, N728);
not NOT1 (N745, N743);
not NOT1 (N746, N745);
or OR2 (N747, N741, N362);
and AND2 (N748, N746, N590);
not NOT1 (N749, N744);
not NOT1 (N750, N742);
nand NAND3 (N751, N750, N633, N317);
or OR3 (N752, N748, N135, N471);
nand NAND2 (N753, N749, N699);
not NOT1 (N754, N752);
nand NAND2 (N755, N737, N180);
buf BUF1 (N756, N747);
xor XOR2 (N757, N719, N645);
nand NAND4 (N758, N724, N21, N464, N39);
nand NAND3 (N759, N751, N44, N19);
nor NOR2 (N760, N759, N753);
nor NOR4 (N761, N509, N571, N299, N207);
nand NAND3 (N762, N736, N572, N720);
nor NOR3 (N763, N740, N180, N691);
or OR2 (N764, N760, N578);
not NOT1 (N765, N761);
and AND3 (N766, N756, N682, N578);
not NOT1 (N767, N735);
or OR3 (N768, N765, N508, N264);
buf BUF1 (N769, N762);
or OR2 (N770, N764, N560);
or OR3 (N771, N768, N474, N528);
xor XOR2 (N772, N758, N366);
xor XOR2 (N773, N757, N328);
buf BUF1 (N774, N767);
buf BUF1 (N775, N754);
xor XOR2 (N776, N755, N183);
nor NOR4 (N777, N770, N722, N503, N220);
xor XOR2 (N778, N763, N74);
nor NOR4 (N779, N777, N345, N388, N55);
and AND4 (N780, N775, N368, N433, N201);
buf BUF1 (N781, N780);
nor NOR4 (N782, N776, N510, N261, N64);
buf BUF1 (N783, N772);
and AND2 (N784, N782, N761);
buf BUF1 (N785, N784);
and AND4 (N786, N769, N173, N83, N782);
or OR2 (N787, N766, N256);
xor XOR2 (N788, N783, N463);
not NOT1 (N789, N781);
not NOT1 (N790, N789);
or OR4 (N791, N785, N358, N164, N766);
buf BUF1 (N792, N791);
or OR4 (N793, N773, N93, N315, N580);
nor NOR2 (N794, N788, N599);
nand NAND4 (N795, N779, N653, N651, N663);
nand NAND2 (N796, N794, N449);
nand NAND2 (N797, N796, N113);
not NOT1 (N798, N787);
and AND3 (N799, N798, N730, N755);
buf BUF1 (N800, N786);
or OR3 (N801, N799, N564, N623);
buf BUF1 (N802, N771);
buf BUF1 (N803, N801);
or OR3 (N804, N778, N562, N536);
nand NAND4 (N805, N790, N375, N516, N493);
xor XOR2 (N806, N805, N751);
xor XOR2 (N807, N806, N101);
nor NOR4 (N808, N807, N178, N86, N14);
and AND3 (N809, N808, N706, N663);
not NOT1 (N810, N792);
not NOT1 (N811, N793);
nor NOR2 (N812, N800, N666);
nor NOR2 (N813, N810, N196);
not NOT1 (N814, N803);
nor NOR4 (N815, N813, N459, N364, N475);
buf BUF1 (N816, N774);
or OR2 (N817, N814, N807);
nor NOR4 (N818, N809, N77, N285, N738);
or OR4 (N819, N811, N456, N94, N363);
nor NOR2 (N820, N797, N286);
not NOT1 (N821, N815);
nand NAND3 (N822, N816, N437, N668);
xor XOR2 (N823, N819, N183);
buf BUF1 (N824, N823);
xor XOR2 (N825, N804, N647);
nand NAND3 (N826, N802, N379, N77);
nor NOR3 (N827, N825, N298, N826);
not NOT1 (N828, N233);
and AND2 (N829, N795, N407);
or OR4 (N830, N822, N241, N60, N292);
buf BUF1 (N831, N818);
or OR3 (N832, N831, N206, N321);
buf BUF1 (N833, N824);
buf BUF1 (N834, N829);
xor XOR2 (N835, N833, N533);
and AND4 (N836, N830, N44, N484, N427);
not NOT1 (N837, N820);
and AND2 (N838, N836, N367);
buf BUF1 (N839, N817);
not NOT1 (N840, N821);
not NOT1 (N841, N838);
buf BUF1 (N842, N827);
and AND2 (N843, N834, N385);
not NOT1 (N844, N837);
nand NAND2 (N845, N843, N459);
not NOT1 (N846, N842);
nand NAND4 (N847, N812, N563, N127, N822);
nor NOR4 (N848, N846, N694, N9, N493);
nor NOR3 (N849, N840, N171, N300);
nand NAND4 (N850, N849, N570, N669, N667);
nand NAND3 (N851, N844, N429, N807);
or OR4 (N852, N845, N707, N352, N7);
xor XOR2 (N853, N848, N409);
nand NAND2 (N854, N839, N514);
not NOT1 (N855, N847);
nor NOR2 (N856, N853, N397);
or OR2 (N857, N850, N54);
or OR3 (N858, N852, N326, N269);
xor XOR2 (N859, N857, N265);
buf BUF1 (N860, N835);
nand NAND3 (N861, N854, N544, N438);
and AND3 (N862, N828, N47, N559);
xor XOR2 (N863, N856, N648);
xor XOR2 (N864, N860, N87);
xor XOR2 (N865, N864, N138);
and AND2 (N866, N859, N225);
or OR2 (N867, N855, N51);
xor XOR2 (N868, N866, N207);
not NOT1 (N869, N868);
xor XOR2 (N870, N865, N476);
nor NOR2 (N871, N867, N424);
or OR4 (N872, N869, N741, N233, N84);
xor XOR2 (N873, N862, N593);
and AND2 (N874, N861, N364);
xor XOR2 (N875, N832, N299);
and AND3 (N876, N863, N667, N81);
nand NAND2 (N877, N858, N320);
not NOT1 (N878, N873);
nand NAND4 (N879, N841, N121, N818, N96);
buf BUF1 (N880, N871);
nor NOR3 (N881, N876, N467, N612);
xor XOR2 (N882, N872, N189);
not NOT1 (N883, N875);
nor NOR2 (N884, N851, N74);
xor XOR2 (N885, N878, N410);
xor XOR2 (N886, N870, N153);
or OR4 (N887, N885, N378, N210, N626);
nand NAND2 (N888, N886, N684);
or OR4 (N889, N883, N22, N435, N144);
and AND3 (N890, N888, N217, N539);
not NOT1 (N891, N879);
nand NAND4 (N892, N884, N666, N523, N62);
and AND3 (N893, N889, N416, N585);
nor NOR2 (N894, N891, N107);
nor NOR4 (N895, N882, N671, N791, N59);
not NOT1 (N896, N880);
buf BUF1 (N897, N893);
and AND4 (N898, N881, N757, N702, N72);
xor XOR2 (N899, N877, N577);
nor NOR3 (N900, N894, N552, N850);
buf BUF1 (N901, N890);
or OR4 (N902, N897, N134, N811, N316);
nand NAND3 (N903, N899, N319, N569);
xor XOR2 (N904, N903, N327);
nor NOR2 (N905, N887, N362);
buf BUF1 (N906, N898);
xor XOR2 (N907, N905, N395);
or OR3 (N908, N895, N710, N819);
nand NAND3 (N909, N902, N451, N236);
xor XOR2 (N910, N909, N41);
not NOT1 (N911, N892);
nor NOR3 (N912, N906, N166, N858);
nor NOR2 (N913, N901, N868);
or OR2 (N914, N911, N569);
nor NOR4 (N915, N907, N209, N182, N426);
or OR2 (N916, N912, N327);
nand NAND4 (N917, N916, N3, N87, N732);
or OR3 (N918, N908, N516, N201);
buf BUF1 (N919, N915);
not NOT1 (N920, N917);
or OR2 (N921, N900, N647);
xor XOR2 (N922, N874, N713);
nand NAND3 (N923, N914, N89, N713);
nand NAND4 (N924, N913, N402, N196, N42);
xor XOR2 (N925, N918, N924);
buf BUF1 (N926, N652);
or OR2 (N927, N910, N652);
nor NOR4 (N928, N926, N158, N2, N428);
nor NOR3 (N929, N927, N924, N797);
xor XOR2 (N930, N920, N283);
or OR3 (N931, N919, N114, N613);
nor NOR3 (N932, N925, N744, N548);
not NOT1 (N933, N922);
nand NAND3 (N934, N928, N298, N683);
nor NOR2 (N935, N934, N685);
buf BUF1 (N936, N929);
and AND4 (N937, N933, N737, N737, N290);
or OR2 (N938, N936, N387);
not NOT1 (N939, N935);
nor NOR3 (N940, N930, N247, N505);
or OR2 (N941, N932, N629);
and AND4 (N942, N937, N912, N308, N801);
xor XOR2 (N943, N940, N110);
or OR3 (N944, N939, N878, N488);
xor XOR2 (N945, N943, N942);
buf BUF1 (N946, N371);
nand NAND2 (N947, N904, N694);
nand NAND4 (N948, N923, N806, N32, N84);
and AND4 (N949, N896, N112, N854, N288);
nand NAND4 (N950, N931, N285, N406, N163);
nand NAND3 (N951, N941, N730, N90);
buf BUF1 (N952, N949);
or OR4 (N953, N950, N778, N88, N304);
nand NAND2 (N954, N946, N156);
nand NAND4 (N955, N948, N450, N626, N472);
and AND4 (N956, N945, N442, N777, N550);
nand NAND4 (N957, N944, N253, N260, N133);
xor XOR2 (N958, N955, N763);
and AND4 (N959, N957, N946, N35, N273);
and AND2 (N960, N947, N333);
nor NOR3 (N961, N958, N627, N214);
nand NAND3 (N962, N959, N229, N272);
nor NOR2 (N963, N951, N409);
xor XOR2 (N964, N963, N449);
not NOT1 (N965, N921);
and AND3 (N966, N953, N346, N410);
or OR3 (N967, N962, N509, N147);
or OR4 (N968, N967, N151, N651, N729);
xor XOR2 (N969, N965, N270);
buf BUF1 (N970, N968);
or OR2 (N971, N960, N575);
nor NOR4 (N972, N961, N326, N561, N888);
and AND3 (N973, N956, N7, N311);
xor XOR2 (N974, N938, N865);
not NOT1 (N975, N970);
xor XOR2 (N976, N964, N786);
xor XOR2 (N977, N973, N522);
not NOT1 (N978, N966);
not NOT1 (N979, N974);
buf BUF1 (N980, N972);
nand NAND4 (N981, N971, N947, N707, N282);
xor XOR2 (N982, N979, N931);
nor NOR4 (N983, N982, N34, N907, N873);
not NOT1 (N984, N952);
and AND2 (N985, N954, N767);
buf BUF1 (N986, N977);
nor NOR3 (N987, N976, N433, N825);
or OR4 (N988, N983, N843, N930, N15);
xor XOR2 (N989, N986, N196);
not NOT1 (N990, N988);
nand NAND4 (N991, N989, N192, N661, N46);
or OR4 (N992, N991, N399, N931, N955);
nand NAND2 (N993, N975, N730);
nor NOR4 (N994, N987, N476, N963, N167);
not NOT1 (N995, N981);
xor XOR2 (N996, N984, N37);
xor XOR2 (N997, N969, N511);
buf BUF1 (N998, N985);
buf BUF1 (N999, N997);
buf BUF1 (N1000, N996);
xor XOR2 (N1001, N993, N994);
and AND4 (N1002, N42, N955, N750, N888);
xor XOR2 (N1003, N1002, N628);
or OR4 (N1004, N1001, N407, N70, N238);
nor NOR3 (N1005, N999, N401, N52);
xor XOR2 (N1006, N980, N273);
and AND4 (N1007, N1006, N737, N833, N591);
not NOT1 (N1008, N1005);
xor XOR2 (N1009, N1003, N662);
or OR2 (N1010, N992, N1003);
xor XOR2 (N1011, N1007, N347);
buf BUF1 (N1012, N990);
or OR2 (N1013, N1008, N349);
and AND2 (N1014, N1009, N520);
nand NAND2 (N1015, N1014, N540);
and AND3 (N1016, N1012, N111, N516);
nand NAND4 (N1017, N998, N454, N1006, N966);
and AND2 (N1018, N1004, N165);
nand NAND4 (N1019, N1016, N665, N632, N488);
nand NAND3 (N1020, N1013, N205, N686);
or OR2 (N1021, N1018, N749);
buf BUF1 (N1022, N1019);
xor XOR2 (N1023, N1017, N805);
and AND3 (N1024, N1022, N145, N520);
nand NAND4 (N1025, N978, N786, N377, N985);
or OR4 (N1026, N1024, N286, N423, N267);
and AND2 (N1027, N1000, N540);
or OR2 (N1028, N995, N917);
buf BUF1 (N1029, N1023);
and AND2 (N1030, N1025, N165);
not NOT1 (N1031, N1010);
buf BUF1 (N1032, N1030);
nand NAND3 (N1033, N1026, N968, N897);
not NOT1 (N1034, N1015);
buf BUF1 (N1035, N1032);
and AND2 (N1036, N1034, N208);
nand NAND3 (N1037, N1021, N87, N248);
buf BUF1 (N1038, N1036);
xor XOR2 (N1039, N1037, N1017);
not NOT1 (N1040, N1027);
and AND3 (N1041, N1031, N45, N239);
and AND3 (N1042, N1020, N914, N722);
or OR3 (N1043, N1041, N205, N874);
nor NOR4 (N1044, N1039, N362, N628, N473);
nor NOR2 (N1045, N1044, N965);
not NOT1 (N1046, N1043);
xor XOR2 (N1047, N1011, N236);
nor NOR3 (N1048, N1028, N400, N203);
or OR4 (N1049, N1046, N560, N19, N178);
xor XOR2 (N1050, N1047, N424);
nor NOR4 (N1051, N1045, N673, N1028, N529);
nand NAND3 (N1052, N1042, N550, N1);
buf BUF1 (N1053, N1029);
and AND4 (N1054, N1035, N391, N487, N791);
or OR4 (N1055, N1053, N788, N883, N545);
buf BUF1 (N1056, N1054);
buf BUF1 (N1057, N1052);
nand NAND2 (N1058, N1049, N647);
buf BUF1 (N1059, N1056);
nor NOR4 (N1060, N1040, N688, N9, N400);
nor NOR4 (N1061, N1048, N599, N599, N1051);
nor NOR2 (N1062, N533, N608);
not NOT1 (N1063, N1055);
nand NAND2 (N1064, N1062, N984);
not NOT1 (N1065, N1038);
buf BUF1 (N1066, N1061);
nor NOR4 (N1067, N1065, N423, N184, N324);
nand NAND2 (N1068, N1059, N1047);
nor NOR2 (N1069, N1058, N727);
nand NAND3 (N1070, N1064, N392, N510);
nand NAND3 (N1071, N1070, N336, N835);
or OR4 (N1072, N1033, N154, N782, N234);
buf BUF1 (N1073, N1069);
or OR3 (N1074, N1073, N97, N274);
xor XOR2 (N1075, N1057, N844);
nand NAND3 (N1076, N1067, N863, N1041);
or OR3 (N1077, N1071, N359, N571);
xor XOR2 (N1078, N1060, N1022);
not NOT1 (N1079, N1078);
xor XOR2 (N1080, N1077, N173);
or OR2 (N1081, N1050, N882);
xor XOR2 (N1082, N1080, N951);
nor NOR3 (N1083, N1079, N347, N107);
and AND3 (N1084, N1063, N693, N389);
buf BUF1 (N1085, N1074);
or OR3 (N1086, N1066, N489, N236);
nor NOR2 (N1087, N1068, N606);
or OR2 (N1088, N1084, N6);
nor NOR4 (N1089, N1087, N715, N513, N403);
and AND4 (N1090, N1085, N343, N300, N156);
not NOT1 (N1091, N1083);
nor NOR3 (N1092, N1076, N819, N1055);
not NOT1 (N1093, N1075);
or OR2 (N1094, N1082, N185);
nor NOR3 (N1095, N1090, N27, N735);
nand NAND2 (N1096, N1081, N1042);
buf BUF1 (N1097, N1072);
and AND2 (N1098, N1095, N140);
not NOT1 (N1099, N1096);
not NOT1 (N1100, N1086);
xor XOR2 (N1101, N1098, N258);
buf BUF1 (N1102, N1088);
nand NAND3 (N1103, N1092, N21, N935);
and AND3 (N1104, N1094, N645, N1102);
buf BUF1 (N1105, N454);
buf BUF1 (N1106, N1104);
buf BUF1 (N1107, N1091);
xor XOR2 (N1108, N1101, N551);
or OR2 (N1109, N1108, N351);
xor XOR2 (N1110, N1089, N935);
or OR4 (N1111, N1100, N671, N347, N576);
nand NAND3 (N1112, N1110, N985, N151);
and AND2 (N1113, N1097, N170);
nor NOR3 (N1114, N1107, N811, N660);
nand NAND2 (N1115, N1093, N51);
buf BUF1 (N1116, N1105);
xor XOR2 (N1117, N1113, N811);
xor XOR2 (N1118, N1109, N450);
buf BUF1 (N1119, N1118);
nor NOR4 (N1120, N1099, N39, N842, N1109);
xor XOR2 (N1121, N1106, N380);
and AND2 (N1122, N1120, N441);
buf BUF1 (N1123, N1117);
nand NAND4 (N1124, N1111, N794, N62, N675);
or OR2 (N1125, N1123, N17);
nand NAND2 (N1126, N1116, N499);
or OR3 (N1127, N1122, N802, N808);
buf BUF1 (N1128, N1103);
or OR3 (N1129, N1119, N25, N233);
xor XOR2 (N1130, N1129, N234);
or OR4 (N1131, N1130, N507, N185, N94);
nand NAND4 (N1132, N1114, N506, N245, N1107);
nor NOR3 (N1133, N1115, N140, N795);
nor NOR3 (N1134, N1112, N289, N53);
nor NOR3 (N1135, N1125, N717, N723);
nand NAND4 (N1136, N1132, N161, N967, N489);
buf BUF1 (N1137, N1135);
or OR3 (N1138, N1134, N1074, N600);
xor XOR2 (N1139, N1133, N369);
or OR2 (N1140, N1127, N755);
or OR3 (N1141, N1136, N744, N472);
nor NOR2 (N1142, N1140, N1028);
nand NAND3 (N1143, N1139, N107, N1070);
nand NAND4 (N1144, N1124, N364, N1008, N738);
nor NOR4 (N1145, N1144, N371, N1014, N694);
and AND4 (N1146, N1142, N381, N12, N528);
not NOT1 (N1147, N1146);
and AND3 (N1148, N1145, N811, N311);
buf BUF1 (N1149, N1148);
buf BUF1 (N1150, N1137);
nor NOR4 (N1151, N1143, N393, N888, N456);
xor XOR2 (N1152, N1150, N147);
and AND4 (N1153, N1138, N835, N566, N738);
nor NOR3 (N1154, N1152, N72, N905);
nand NAND3 (N1155, N1151, N1055, N706);
nand NAND3 (N1156, N1141, N275, N685);
nor NOR3 (N1157, N1128, N794, N304);
xor XOR2 (N1158, N1149, N797);
nor NOR3 (N1159, N1126, N1153, N1086);
nor NOR2 (N1160, N569, N709);
buf BUF1 (N1161, N1147);
nand NAND2 (N1162, N1156, N1153);
xor XOR2 (N1163, N1162, N583);
xor XOR2 (N1164, N1154, N742);
not NOT1 (N1165, N1163);
or OR3 (N1166, N1131, N933, N239);
not NOT1 (N1167, N1164);
or OR2 (N1168, N1159, N156);
nor NOR4 (N1169, N1160, N228, N1060, N212);
buf BUF1 (N1170, N1167);
and AND3 (N1171, N1170, N741, N864);
buf BUF1 (N1172, N1168);
or OR3 (N1173, N1157, N153, N710);
and AND3 (N1174, N1161, N521, N129);
not NOT1 (N1175, N1169);
or OR2 (N1176, N1174, N155);
nor NOR2 (N1177, N1166, N851);
buf BUF1 (N1178, N1176);
xor XOR2 (N1179, N1173, N95);
not NOT1 (N1180, N1172);
nor NOR3 (N1181, N1165, N772, N706);
xor XOR2 (N1182, N1178, N1);
buf BUF1 (N1183, N1180);
xor XOR2 (N1184, N1181, N878);
or OR2 (N1185, N1158, N281);
and AND4 (N1186, N1177, N20, N722, N161);
nor NOR4 (N1187, N1183, N1153, N841, N454);
and AND2 (N1188, N1121, N447);
and AND3 (N1189, N1155, N929, N151);
nor NOR2 (N1190, N1189, N510);
or OR2 (N1191, N1184, N1038);
or OR3 (N1192, N1186, N664, N988);
or OR3 (N1193, N1188, N826, N1003);
xor XOR2 (N1194, N1175, N522);
nor NOR3 (N1195, N1185, N437, N670);
buf BUF1 (N1196, N1195);
or OR4 (N1197, N1193, N635, N577, N857);
nand NAND4 (N1198, N1190, N722, N211, N938);
buf BUF1 (N1199, N1196);
and AND2 (N1200, N1198, N514);
nand NAND2 (N1201, N1199, N268);
nor NOR3 (N1202, N1194, N1067, N124);
or OR4 (N1203, N1197, N1070, N208, N586);
buf BUF1 (N1204, N1192);
xor XOR2 (N1205, N1171, N383);
nor NOR2 (N1206, N1205, N620);
nor NOR3 (N1207, N1201, N588, N213);
buf BUF1 (N1208, N1179);
xor XOR2 (N1209, N1207, N175);
xor XOR2 (N1210, N1200, N1134);
buf BUF1 (N1211, N1203);
buf BUF1 (N1212, N1208);
and AND4 (N1213, N1202, N178, N918, N1091);
or OR2 (N1214, N1209, N955);
xor XOR2 (N1215, N1214, N448);
nor NOR4 (N1216, N1210, N1110, N750, N224);
and AND4 (N1217, N1182, N1083, N681, N1020);
nand NAND3 (N1218, N1213, N657, N830);
xor XOR2 (N1219, N1206, N759);
nand NAND4 (N1220, N1191, N113, N1158, N971);
buf BUF1 (N1221, N1220);
xor XOR2 (N1222, N1219, N227);
xor XOR2 (N1223, N1204, N614);
and AND2 (N1224, N1221, N1084);
or OR4 (N1225, N1223, N162, N427, N90);
nand NAND2 (N1226, N1211, N965);
or OR4 (N1227, N1222, N502, N659, N778);
and AND3 (N1228, N1217, N160, N1084);
not NOT1 (N1229, N1215);
or OR3 (N1230, N1227, N202, N117);
and AND2 (N1231, N1225, N10);
xor XOR2 (N1232, N1218, N1061);
buf BUF1 (N1233, N1228);
not NOT1 (N1234, N1233);
xor XOR2 (N1235, N1226, N917);
buf BUF1 (N1236, N1232);
and AND4 (N1237, N1230, N565, N1020, N943);
nor NOR2 (N1238, N1234, N228);
and AND3 (N1239, N1224, N325, N1078);
not NOT1 (N1240, N1235);
nor NOR3 (N1241, N1231, N567, N392);
or OR2 (N1242, N1236, N493);
not NOT1 (N1243, N1240);
buf BUF1 (N1244, N1212);
buf BUF1 (N1245, N1238);
xor XOR2 (N1246, N1244, N1063);
nand NAND2 (N1247, N1242, N1039);
buf BUF1 (N1248, N1229);
or OR4 (N1249, N1237, N402, N770, N520);
nor NOR3 (N1250, N1243, N214, N668);
and AND2 (N1251, N1247, N180);
nor NOR4 (N1252, N1187, N897, N567, N569);
buf BUF1 (N1253, N1241);
or OR3 (N1254, N1239, N1085, N964);
and AND3 (N1255, N1253, N709, N818);
and AND3 (N1256, N1254, N249, N639);
not NOT1 (N1257, N1251);
not NOT1 (N1258, N1245);
nor NOR4 (N1259, N1250, N356, N515, N441);
or OR4 (N1260, N1216, N379, N369, N201);
buf BUF1 (N1261, N1258);
or OR4 (N1262, N1248, N264, N173, N210);
nor NOR2 (N1263, N1255, N145);
and AND2 (N1264, N1263, N729);
nor NOR4 (N1265, N1260, N750, N1001, N588);
xor XOR2 (N1266, N1252, N13);
xor XOR2 (N1267, N1246, N304);
or OR4 (N1268, N1267, N338, N1258, N565);
not NOT1 (N1269, N1266);
nand NAND3 (N1270, N1265, N846, N1037);
nand NAND2 (N1271, N1261, N148);
nor NOR4 (N1272, N1268, N1133, N597, N1152);
and AND4 (N1273, N1259, N1006, N608, N152);
or OR2 (N1274, N1257, N305);
nor NOR2 (N1275, N1273, N324);
buf BUF1 (N1276, N1256);
not NOT1 (N1277, N1270);
buf BUF1 (N1278, N1271);
buf BUF1 (N1279, N1262);
xor XOR2 (N1280, N1249, N192);
nor NOR3 (N1281, N1279, N21, N709);
nor NOR4 (N1282, N1280, N738, N532, N356);
and AND3 (N1283, N1264, N601, N809);
or OR2 (N1284, N1281, N632);
xor XOR2 (N1285, N1272, N843);
nand NAND3 (N1286, N1284, N258, N129);
or OR2 (N1287, N1285, N1064);
and AND2 (N1288, N1277, N1103);
and AND4 (N1289, N1278, N904, N533, N219);
nor NOR4 (N1290, N1282, N219, N637, N897);
nand NAND4 (N1291, N1288, N749, N7, N150);
xor XOR2 (N1292, N1286, N695);
or OR2 (N1293, N1289, N206);
nand NAND3 (N1294, N1293, N1128, N1008);
xor XOR2 (N1295, N1294, N468);
xor XOR2 (N1296, N1276, N1117);
or OR4 (N1297, N1296, N932, N25, N252);
and AND3 (N1298, N1269, N244, N1110);
nand NAND2 (N1299, N1274, N1016);
buf BUF1 (N1300, N1290);
xor XOR2 (N1301, N1295, N810);
xor XOR2 (N1302, N1275, N49);
nor NOR3 (N1303, N1301, N346, N1232);
or OR2 (N1304, N1302, N812);
buf BUF1 (N1305, N1298);
nor NOR3 (N1306, N1303, N1012, N429);
buf BUF1 (N1307, N1283);
or OR3 (N1308, N1307, N1102, N380);
nor NOR4 (N1309, N1305, N1123, N1273, N1061);
xor XOR2 (N1310, N1309, N864);
xor XOR2 (N1311, N1291, N1007);
nand NAND3 (N1312, N1310, N587, N132);
xor XOR2 (N1313, N1300, N529);
nor NOR3 (N1314, N1297, N638, N460);
not NOT1 (N1315, N1313);
nand NAND2 (N1316, N1304, N713);
buf BUF1 (N1317, N1314);
nor NOR2 (N1318, N1299, N952);
not NOT1 (N1319, N1316);
nand NAND4 (N1320, N1287, N881, N878, N454);
nand NAND3 (N1321, N1306, N114, N1220);
nor NOR3 (N1322, N1311, N1047, N541);
nor NOR2 (N1323, N1312, N740);
or OR2 (N1324, N1308, N858);
and AND2 (N1325, N1323, N89);
or OR4 (N1326, N1319, N1117, N134, N981);
and AND2 (N1327, N1324, N116);
nor NOR4 (N1328, N1318, N1087, N623, N376);
not NOT1 (N1329, N1327);
buf BUF1 (N1330, N1325);
and AND3 (N1331, N1330, N380, N120);
nor NOR4 (N1332, N1317, N1295, N791, N780);
not NOT1 (N1333, N1328);
or OR3 (N1334, N1315, N399, N573);
or OR2 (N1335, N1321, N1326);
not NOT1 (N1336, N849);
and AND4 (N1337, N1335, N541, N1064, N832);
not NOT1 (N1338, N1332);
nand NAND2 (N1339, N1337, N612);
nand NAND4 (N1340, N1338, N811, N1337, N439);
nand NAND3 (N1341, N1340, N385, N479);
not NOT1 (N1342, N1322);
xor XOR2 (N1343, N1333, N109);
not NOT1 (N1344, N1292);
and AND3 (N1345, N1343, N1307, N1211);
xor XOR2 (N1346, N1336, N17);
buf BUF1 (N1347, N1345);
nand NAND4 (N1348, N1347, N754, N904, N162);
xor XOR2 (N1349, N1344, N756);
nand NAND2 (N1350, N1329, N1319);
or OR2 (N1351, N1350, N779);
nor NOR3 (N1352, N1339, N165, N521);
not NOT1 (N1353, N1346);
nand NAND3 (N1354, N1341, N992, N1035);
xor XOR2 (N1355, N1331, N1347);
or OR3 (N1356, N1349, N592, N1159);
nor NOR2 (N1357, N1352, N273);
xor XOR2 (N1358, N1348, N1048);
buf BUF1 (N1359, N1354);
or OR4 (N1360, N1320, N108, N29, N391);
buf BUF1 (N1361, N1357);
xor XOR2 (N1362, N1342, N109);
xor XOR2 (N1363, N1356, N508);
not NOT1 (N1364, N1334);
buf BUF1 (N1365, N1362);
not NOT1 (N1366, N1361);
nand NAND2 (N1367, N1358, N235);
or OR3 (N1368, N1366, N229, N1351);
and AND4 (N1369, N1030, N250, N766, N920);
not NOT1 (N1370, N1368);
xor XOR2 (N1371, N1359, N54);
and AND3 (N1372, N1364, N1132, N1124);
nor NOR2 (N1373, N1360, N39);
nor NOR3 (N1374, N1355, N524, N1265);
xor XOR2 (N1375, N1370, N136);
not NOT1 (N1376, N1363);
nor NOR3 (N1377, N1372, N981, N829);
not NOT1 (N1378, N1371);
buf BUF1 (N1379, N1369);
buf BUF1 (N1380, N1367);
xor XOR2 (N1381, N1380, N337);
nor NOR4 (N1382, N1375, N1150, N247, N220);
not NOT1 (N1383, N1379);
nor NOR3 (N1384, N1382, N1026, N272);
and AND4 (N1385, N1378, N736, N929, N1103);
buf BUF1 (N1386, N1377);
nor NOR4 (N1387, N1383, N799, N864, N798);
nor NOR3 (N1388, N1385, N227, N1220);
or OR3 (N1389, N1381, N188, N293);
xor XOR2 (N1390, N1376, N804);
or OR2 (N1391, N1389, N909);
or OR2 (N1392, N1388, N694);
not NOT1 (N1393, N1392);
xor XOR2 (N1394, N1391, N695);
xor XOR2 (N1395, N1393, N69);
and AND4 (N1396, N1387, N1246, N644, N197);
nand NAND2 (N1397, N1365, N852);
xor XOR2 (N1398, N1395, N1268);
xor XOR2 (N1399, N1373, N95);
or OR2 (N1400, N1394, N303);
and AND3 (N1401, N1400, N1253, N34);
and AND3 (N1402, N1386, N686, N130);
nor NOR4 (N1403, N1353, N472, N1139, N82);
xor XOR2 (N1404, N1403, N240);
or OR4 (N1405, N1384, N1370, N202, N347);
nor NOR3 (N1406, N1405, N811, N361);
buf BUF1 (N1407, N1397);
nor NOR2 (N1408, N1402, N1126);
nor NOR3 (N1409, N1408, N77, N1377);
xor XOR2 (N1410, N1401, N797);
xor XOR2 (N1411, N1398, N705);
buf BUF1 (N1412, N1411);
nand NAND2 (N1413, N1407, N332);
nand NAND4 (N1414, N1412, N655, N952, N406);
not NOT1 (N1415, N1410);
nand NAND4 (N1416, N1374, N89, N706, N47);
buf BUF1 (N1417, N1413);
nor NOR2 (N1418, N1415, N771);
and AND4 (N1419, N1406, N12, N971, N559);
not NOT1 (N1420, N1390);
buf BUF1 (N1421, N1396);
buf BUF1 (N1422, N1414);
buf BUF1 (N1423, N1409);
or OR2 (N1424, N1423, N1317);
not NOT1 (N1425, N1417);
buf BUF1 (N1426, N1425);
and AND4 (N1427, N1421, N371, N1339, N801);
nand NAND3 (N1428, N1426, N92, N1201);
not NOT1 (N1429, N1418);
nor NOR2 (N1430, N1428, N902);
nor NOR4 (N1431, N1424, N1092, N226, N230);
nor NOR3 (N1432, N1427, N202, N452);
or OR4 (N1433, N1429, N537, N994, N874);
nand NAND2 (N1434, N1420, N601);
or OR4 (N1435, N1433, N1117, N1330, N588);
buf BUF1 (N1436, N1404);
xor XOR2 (N1437, N1399, N145);
xor XOR2 (N1438, N1437, N376);
nor NOR4 (N1439, N1422, N766, N534, N1109);
nand NAND3 (N1440, N1435, N927, N146);
not NOT1 (N1441, N1440);
nor NOR2 (N1442, N1439, N1400);
and AND2 (N1443, N1436, N1354);
and AND2 (N1444, N1419, N1012);
or OR2 (N1445, N1416, N1433);
xor XOR2 (N1446, N1444, N915);
not NOT1 (N1447, N1434);
xor XOR2 (N1448, N1445, N481);
nand NAND2 (N1449, N1448, N195);
nor NOR3 (N1450, N1432, N361, N30);
nand NAND4 (N1451, N1442, N403, N1317, N1362);
nand NAND4 (N1452, N1441, N1201, N997, N671);
or OR3 (N1453, N1431, N676, N304);
buf BUF1 (N1454, N1443);
not NOT1 (N1455, N1450);
xor XOR2 (N1456, N1455, N1366);
and AND3 (N1457, N1438, N990, N375);
nand NAND3 (N1458, N1447, N8, N1002);
nor NOR2 (N1459, N1456, N133);
not NOT1 (N1460, N1452);
xor XOR2 (N1461, N1458, N930);
and AND4 (N1462, N1453, N852, N172, N1079);
buf BUF1 (N1463, N1449);
nor NOR4 (N1464, N1430, N1117, N868, N227);
nand NAND4 (N1465, N1457, N904, N179, N250);
nand NAND4 (N1466, N1465, N396, N79, N828);
not NOT1 (N1467, N1466);
or OR3 (N1468, N1463, N900, N1385);
or OR2 (N1469, N1467, N650);
xor XOR2 (N1470, N1460, N198);
or OR2 (N1471, N1468, N1065);
nand NAND4 (N1472, N1461, N1415, N49, N342);
nand NAND3 (N1473, N1470, N252, N913);
nor NOR3 (N1474, N1462, N849, N318);
nor NOR3 (N1475, N1446, N1373, N546);
nand NAND2 (N1476, N1464, N437);
buf BUF1 (N1477, N1475);
and AND3 (N1478, N1473, N204, N1182);
and AND3 (N1479, N1469, N859, N975);
nor NOR4 (N1480, N1479, N293, N361, N375);
buf BUF1 (N1481, N1451);
nor NOR4 (N1482, N1476, N1261, N1165, N671);
and AND3 (N1483, N1482, N633, N662);
nand NAND2 (N1484, N1459, N390);
nand NAND3 (N1485, N1484, N64, N1195);
not NOT1 (N1486, N1480);
and AND3 (N1487, N1485, N459, N139);
xor XOR2 (N1488, N1472, N663);
or OR4 (N1489, N1471, N1451, N655, N832);
not NOT1 (N1490, N1486);
nand NAND2 (N1491, N1487, N240);
or OR4 (N1492, N1478, N253, N461, N111);
nand NAND3 (N1493, N1492, N841, N1161);
buf BUF1 (N1494, N1481);
or OR4 (N1495, N1490, N1099, N830, N195);
and AND2 (N1496, N1477, N608);
nand NAND3 (N1497, N1488, N248, N1026);
buf BUF1 (N1498, N1494);
nand NAND3 (N1499, N1493, N1239, N217);
nor NOR2 (N1500, N1454, N1212);
nand NAND3 (N1501, N1483, N937, N692);
nand NAND3 (N1502, N1474, N1043, N1105);
buf BUF1 (N1503, N1491);
and AND3 (N1504, N1499, N1501, N1486);
nand NAND3 (N1505, N662, N535, N1274);
or OR2 (N1506, N1503, N771);
xor XOR2 (N1507, N1498, N1407);
not NOT1 (N1508, N1489);
buf BUF1 (N1509, N1504);
and AND4 (N1510, N1502, N597, N261, N857);
or OR3 (N1511, N1496, N594, N212);
xor XOR2 (N1512, N1505, N25);
nand NAND4 (N1513, N1511, N438, N1452, N718);
nor NOR4 (N1514, N1495, N1129, N808, N1068);
nand NAND2 (N1515, N1512, N414);
buf BUF1 (N1516, N1514);
not NOT1 (N1517, N1513);
or OR3 (N1518, N1516, N385, N97);
or OR3 (N1519, N1515, N10, N706);
nand NAND4 (N1520, N1500, N629, N1503, N707);
not NOT1 (N1521, N1517);
not NOT1 (N1522, N1506);
nor NOR3 (N1523, N1497, N556, N759);
nand NAND4 (N1524, N1521, N158, N445, N607);
or OR2 (N1525, N1524, N532);
buf BUF1 (N1526, N1507);
nand NAND2 (N1527, N1522, N275);
nand NAND4 (N1528, N1526, N992, N781, N10);
nand NAND2 (N1529, N1525, N1161);
and AND4 (N1530, N1508, N930, N1518, N741);
buf BUF1 (N1531, N184);
or OR2 (N1532, N1527, N233);
xor XOR2 (N1533, N1509, N67);
or OR2 (N1534, N1533, N1434);
not NOT1 (N1535, N1531);
and AND3 (N1536, N1535, N645, N1376);
not NOT1 (N1537, N1523);
buf BUF1 (N1538, N1537);
nand NAND3 (N1539, N1538, N427, N819);
xor XOR2 (N1540, N1510, N1487);
nor NOR4 (N1541, N1530, N942, N1093, N359);
nor NOR3 (N1542, N1534, N1287, N797);
buf BUF1 (N1543, N1532);
and AND4 (N1544, N1543, N279, N350, N440);
and AND3 (N1545, N1520, N882, N407);
nor NOR4 (N1546, N1528, N1071, N548, N452);
and AND3 (N1547, N1540, N1375, N991);
nor NOR4 (N1548, N1546, N1362, N1094, N997);
nand NAND4 (N1549, N1548, N299, N1387, N663);
xor XOR2 (N1550, N1539, N79);
nor NOR3 (N1551, N1529, N1153, N281);
xor XOR2 (N1552, N1541, N1258);
not NOT1 (N1553, N1547);
nand NAND2 (N1554, N1549, N1189);
nor NOR4 (N1555, N1553, N594, N1455, N1377);
and AND2 (N1556, N1542, N690);
buf BUF1 (N1557, N1544);
nor NOR2 (N1558, N1555, N1350);
buf BUF1 (N1559, N1551);
or OR3 (N1560, N1545, N1348, N1431);
nor NOR3 (N1561, N1556, N1383, N1083);
not NOT1 (N1562, N1554);
xor XOR2 (N1563, N1550, N817);
and AND4 (N1564, N1552, N940, N775, N1210);
or OR2 (N1565, N1564, N1304);
nand NAND3 (N1566, N1519, N583, N332);
or OR4 (N1567, N1558, N1452, N40, N1353);
xor XOR2 (N1568, N1562, N1515);
not NOT1 (N1569, N1561);
and AND4 (N1570, N1557, N1318, N1203, N359);
nand NAND3 (N1571, N1559, N1143, N1164);
buf BUF1 (N1572, N1568);
and AND4 (N1573, N1570, N886, N426, N49);
nand NAND2 (N1574, N1572, N79);
buf BUF1 (N1575, N1574);
nand NAND2 (N1576, N1563, N1489);
not NOT1 (N1577, N1571);
not NOT1 (N1578, N1575);
and AND4 (N1579, N1569, N1131, N1220, N914);
xor XOR2 (N1580, N1536, N1291);
nor NOR3 (N1581, N1560, N493, N1294);
not NOT1 (N1582, N1576);
buf BUF1 (N1583, N1582);
nor NOR2 (N1584, N1566, N850);
buf BUF1 (N1585, N1580);
or OR4 (N1586, N1581, N623, N641, N1261);
nor NOR4 (N1587, N1578, N1020, N1549, N1523);
not NOT1 (N1588, N1585);
nor NOR4 (N1589, N1565, N636, N349, N1164);
and AND3 (N1590, N1583, N1107, N906);
nor NOR4 (N1591, N1587, N6, N1224, N87);
or OR4 (N1592, N1589, N14, N563, N336);
not NOT1 (N1593, N1577);
buf BUF1 (N1594, N1584);
not NOT1 (N1595, N1588);
and AND4 (N1596, N1586, N1003, N843, N1108);
nand NAND2 (N1597, N1593, N41);
buf BUF1 (N1598, N1594);
not NOT1 (N1599, N1591);
not NOT1 (N1600, N1597);
not NOT1 (N1601, N1579);
and AND2 (N1602, N1598, N49);
and AND4 (N1603, N1596, N497, N688, N588);
and AND2 (N1604, N1603, N268);
not NOT1 (N1605, N1604);
or OR2 (N1606, N1573, N904);
and AND4 (N1607, N1567, N1505, N468, N980);
nand NAND2 (N1608, N1590, N872);
buf BUF1 (N1609, N1599);
xor XOR2 (N1610, N1605, N609);
and AND3 (N1611, N1592, N1136, N1285);
buf BUF1 (N1612, N1606);
nand NAND4 (N1613, N1608, N1591, N1241, N830);
nand NAND4 (N1614, N1595, N1153, N1123, N1454);
xor XOR2 (N1615, N1611, N21);
nand NAND2 (N1616, N1615, N532);
nor NOR3 (N1617, N1616, N101, N964);
xor XOR2 (N1618, N1609, N464);
not NOT1 (N1619, N1613);
xor XOR2 (N1620, N1610, N1112);
xor XOR2 (N1621, N1601, N1528);
or OR4 (N1622, N1612, N1099, N855, N381);
and AND3 (N1623, N1619, N999, N1219);
buf BUF1 (N1624, N1622);
nor NOR2 (N1625, N1620, N873);
xor XOR2 (N1626, N1621, N652);
nand NAND4 (N1627, N1614, N762, N658, N1475);
xor XOR2 (N1628, N1602, N23);
not NOT1 (N1629, N1618);
nor NOR4 (N1630, N1624, N1305, N957, N1514);
not NOT1 (N1631, N1626);
and AND4 (N1632, N1631, N1291, N499, N1485);
nand NAND4 (N1633, N1623, N788, N576, N411);
or OR4 (N1634, N1630, N133, N1337, N25);
nor NOR2 (N1635, N1627, N1597);
not NOT1 (N1636, N1600);
or OR3 (N1637, N1636, N1505, N362);
or OR2 (N1638, N1637, N1326);
not NOT1 (N1639, N1633);
nor NOR2 (N1640, N1628, N1407);
nor NOR4 (N1641, N1639, N347, N1457, N554);
xor XOR2 (N1642, N1638, N502);
and AND4 (N1643, N1642, N5, N470, N918);
nor NOR3 (N1644, N1640, N682, N962);
buf BUF1 (N1645, N1634);
nor NOR2 (N1646, N1607, N235);
or OR2 (N1647, N1635, N1265);
nand NAND2 (N1648, N1641, N1570);
nor NOR4 (N1649, N1643, N1113, N952, N1215);
or OR2 (N1650, N1617, N1044);
buf BUF1 (N1651, N1646);
buf BUF1 (N1652, N1650);
nor NOR2 (N1653, N1632, N885);
buf BUF1 (N1654, N1644);
nand NAND4 (N1655, N1649, N799, N670, N819);
xor XOR2 (N1656, N1652, N241);
nor NOR3 (N1657, N1651, N18, N656);
buf BUF1 (N1658, N1648);
nand NAND4 (N1659, N1657, N686, N35, N833);
xor XOR2 (N1660, N1653, N1241);
buf BUF1 (N1661, N1660);
or OR3 (N1662, N1625, N532, N324);
not NOT1 (N1663, N1662);
nor NOR2 (N1664, N1661, N602);
buf BUF1 (N1665, N1629);
nor NOR3 (N1666, N1664, N240, N995);
buf BUF1 (N1667, N1666);
xor XOR2 (N1668, N1667, N171);
or OR2 (N1669, N1665, N452);
and AND4 (N1670, N1658, N444, N1545, N1249);
or OR2 (N1671, N1659, N530);
nand NAND4 (N1672, N1645, N1247, N1648, N1141);
nor NOR3 (N1673, N1670, N263, N892);
nand NAND3 (N1674, N1672, N1553, N745);
nor NOR4 (N1675, N1674, N930, N669, N581);
xor XOR2 (N1676, N1675, N683);
xor XOR2 (N1677, N1669, N1202);
not NOT1 (N1678, N1676);
buf BUF1 (N1679, N1678);
buf BUF1 (N1680, N1655);
xor XOR2 (N1681, N1673, N1169);
or OR4 (N1682, N1654, N1561, N346, N785);
or OR2 (N1683, N1663, N874);
nor NOR3 (N1684, N1668, N1380, N525);
nand NAND3 (N1685, N1684, N644, N321);
xor XOR2 (N1686, N1677, N560);
buf BUF1 (N1687, N1686);
nor NOR4 (N1688, N1680, N740, N1039, N16);
xor XOR2 (N1689, N1681, N1056);
not NOT1 (N1690, N1679);
buf BUF1 (N1691, N1682);
or OR3 (N1692, N1685, N441, N1003);
not NOT1 (N1693, N1683);
nand NAND2 (N1694, N1688, N918);
nor NOR3 (N1695, N1656, N1257, N1593);
xor XOR2 (N1696, N1694, N1097);
or OR2 (N1697, N1693, N877);
or OR3 (N1698, N1647, N148, N391);
xor XOR2 (N1699, N1696, N890);
and AND4 (N1700, N1698, N1485, N376, N114);
nor NOR3 (N1701, N1687, N1442, N1514);
not NOT1 (N1702, N1697);
nand NAND2 (N1703, N1699, N582);
nand NAND4 (N1704, N1703, N271, N1592, N989);
xor XOR2 (N1705, N1702, N881);
buf BUF1 (N1706, N1692);
or OR4 (N1707, N1706, N491, N849, N894);
nor NOR2 (N1708, N1700, N1162);
nand NAND4 (N1709, N1704, N1405, N1689, N43);
nor NOR2 (N1710, N1682, N483);
or OR4 (N1711, N1709, N372, N905, N580);
xor XOR2 (N1712, N1705, N427);
and AND2 (N1713, N1708, N426);
and AND3 (N1714, N1710, N428, N228);
and AND3 (N1715, N1712, N1150, N141);
not NOT1 (N1716, N1714);
xor XOR2 (N1717, N1691, N1086);
xor XOR2 (N1718, N1671, N719);
xor XOR2 (N1719, N1717, N281);
nand NAND2 (N1720, N1719, N1380);
nand NAND4 (N1721, N1690, N794, N944, N1293);
not NOT1 (N1722, N1711);
nor NOR4 (N1723, N1720, N424, N1465, N82);
nand NAND2 (N1724, N1695, N610);
nor NOR3 (N1725, N1701, N1183, N79);
or OR3 (N1726, N1713, N660, N259);
nand NAND4 (N1727, N1725, N1198, N1446, N1358);
not NOT1 (N1728, N1723);
nor NOR3 (N1729, N1727, N765, N950);
nor NOR2 (N1730, N1715, N602);
nor NOR2 (N1731, N1707, N242);
and AND2 (N1732, N1721, N282);
buf BUF1 (N1733, N1722);
xor XOR2 (N1734, N1718, N828);
buf BUF1 (N1735, N1728);
nor NOR4 (N1736, N1735, N1725, N1387, N748);
and AND2 (N1737, N1730, N1412);
not NOT1 (N1738, N1734);
buf BUF1 (N1739, N1732);
nor NOR2 (N1740, N1736, N1567);
or OR2 (N1741, N1716, N1506);
xor XOR2 (N1742, N1737, N985);
nor NOR3 (N1743, N1739, N290, N588);
or OR3 (N1744, N1741, N706, N1152);
and AND4 (N1745, N1731, N820, N285, N100);
nor NOR3 (N1746, N1724, N745, N1450);
xor XOR2 (N1747, N1746, N241);
nand NAND3 (N1748, N1744, N1385, N612);
not NOT1 (N1749, N1738);
not NOT1 (N1750, N1745);
not NOT1 (N1751, N1749);
nand NAND4 (N1752, N1747, N865, N170, N441);
nand NAND2 (N1753, N1752, N17);
and AND3 (N1754, N1740, N1447, N926);
and AND3 (N1755, N1733, N1079, N1262);
and AND3 (N1756, N1755, N956, N1583);
buf BUF1 (N1757, N1748);
nor NOR2 (N1758, N1742, N588);
not NOT1 (N1759, N1754);
or OR3 (N1760, N1757, N221, N1544);
buf BUF1 (N1761, N1729);
nor NOR4 (N1762, N1760, N1493, N920, N1353);
not NOT1 (N1763, N1751);
nand NAND2 (N1764, N1743, N1301);
nor NOR2 (N1765, N1756, N1165);
nor NOR2 (N1766, N1753, N812);
and AND2 (N1767, N1750, N962);
or OR2 (N1768, N1759, N470);
xor XOR2 (N1769, N1767, N933);
not NOT1 (N1770, N1726);
nor NOR4 (N1771, N1761, N1544, N268, N829);
xor XOR2 (N1772, N1770, N1166);
buf BUF1 (N1773, N1763);
nand NAND4 (N1774, N1762, N696, N1002, N1243);
or OR4 (N1775, N1773, N1188, N1158, N1581);
not NOT1 (N1776, N1775);
not NOT1 (N1777, N1768);
nand NAND3 (N1778, N1777, N136, N679);
nand NAND3 (N1779, N1765, N1724, N1433);
or OR2 (N1780, N1776, N553);
buf BUF1 (N1781, N1758);
nor NOR3 (N1782, N1764, N972, N1382);
xor XOR2 (N1783, N1772, N234);
buf BUF1 (N1784, N1779);
nor NOR2 (N1785, N1781, N1712);
xor XOR2 (N1786, N1769, N194);
nor NOR4 (N1787, N1786, N639, N177, N1230);
xor XOR2 (N1788, N1780, N1454);
and AND3 (N1789, N1782, N892, N497);
not NOT1 (N1790, N1787);
xor XOR2 (N1791, N1789, N866);
nor NOR3 (N1792, N1783, N1679, N622);
nor NOR3 (N1793, N1792, N716, N1213);
not NOT1 (N1794, N1791);
not NOT1 (N1795, N1788);
not NOT1 (N1796, N1795);
not NOT1 (N1797, N1794);
buf BUF1 (N1798, N1797);
nor NOR3 (N1799, N1798, N1580, N990);
nor NOR3 (N1800, N1784, N1556, N1491);
and AND4 (N1801, N1800, N146, N448, N1165);
nand NAND3 (N1802, N1796, N320, N335);
and AND2 (N1803, N1793, N1403);
xor XOR2 (N1804, N1766, N1743);
xor XOR2 (N1805, N1778, N842);
not NOT1 (N1806, N1771);
or OR4 (N1807, N1804, N583, N746, N890);
nor NOR2 (N1808, N1805, N1211);
xor XOR2 (N1809, N1802, N710);
nor NOR2 (N1810, N1799, N677);
and AND2 (N1811, N1803, N160);
nand NAND3 (N1812, N1809, N1033, N1706);
and AND2 (N1813, N1801, N436);
and AND2 (N1814, N1806, N260);
xor XOR2 (N1815, N1790, N969);
xor XOR2 (N1816, N1814, N28);
or OR3 (N1817, N1810, N1464, N707);
buf BUF1 (N1818, N1811);
not NOT1 (N1819, N1817);
not NOT1 (N1820, N1819);
nand NAND2 (N1821, N1785, N276);
nor NOR2 (N1822, N1815, N1037);
buf BUF1 (N1823, N1807);
not NOT1 (N1824, N1816);
xor XOR2 (N1825, N1820, N561);
buf BUF1 (N1826, N1823);
xor XOR2 (N1827, N1821, N1711);
nand NAND3 (N1828, N1827, N1222, N1690);
nand NAND2 (N1829, N1808, N1442);
xor XOR2 (N1830, N1828, N596);
nor NOR3 (N1831, N1825, N71, N1560);
nand NAND3 (N1832, N1818, N1473, N148);
or OR4 (N1833, N1812, N1745, N1720, N1542);
or OR4 (N1834, N1826, N198, N1542, N621);
buf BUF1 (N1835, N1822);
or OR4 (N1836, N1834, N581, N1072, N65);
buf BUF1 (N1837, N1813);
buf BUF1 (N1838, N1836);
not NOT1 (N1839, N1824);
xor XOR2 (N1840, N1829, N729);
xor XOR2 (N1841, N1774, N1650);
not NOT1 (N1842, N1831);
and AND4 (N1843, N1840, N252, N14, N1811);
xor XOR2 (N1844, N1833, N130);
xor XOR2 (N1845, N1832, N1213);
buf BUF1 (N1846, N1841);
buf BUF1 (N1847, N1844);
not NOT1 (N1848, N1830);
buf BUF1 (N1849, N1847);
nor NOR2 (N1850, N1842, N815);
xor XOR2 (N1851, N1838, N702);
nand NAND3 (N1852, N1848, N525, N1780);
nor NOR2 (N1853, N1846, N42);
or OR2 (N1854, N1850, N202);
nand NAND4 (N1855, N1837, N1807, N1320, N515);
nand NAND2 (N1856, N1851, N1414);
or OR3 (N1857, N1855, N1246, N546);
or OR2 (N1858, N1839, N935);
buf BUF1 (N1859, N1835);
or OR4 (N1860, N1854, N1475, N865, N1585);
nor NOR3 (N1861, N1849, N247, N987);
xor XOR2 (N1862, N1853, N20);
nor NOR4 (N1863, N1858, N1152, N1657, N109);
or OR2 (N1864, N1843, N1406);
nor NOR2 (N1865, N1863, N1430);
nor NOR2 (N1866, N1862, N708);
buf BUF1 (N1867, N1859);
and AND2 (N1868, N1861, N819);
buf BUF1 (N1869, N1860);
nand NAND3 (N1870, N1867, N1752, N968);
and AND4 (N1871, N1856, N218, N274, N1568);
and AND2 (N1872, N1869, N1678);
and AND2 (N1873, N1864, N436);
nand NAND4 (N1874, N1872, N1622, N1372, N1477);
not NOT1 (N1875, N1873);
nand NAND2 (N1876, N1871, N1738);
and AND3 (N1877, N1865, N1755, N858);
and AND2 (N1878, N1876, N992);
or OR4 (N1879, N1857, N436, N1846, N833);
and AND4 (N1880, N1878, N1577, N1096, N1144);
xor XOR2 (N1881, N1875, N949);
nand NAND2 (N1882, N1881, N533);
or OR2 (N1883, N1877, N1224);
nand NAND4 (N1884, N1870, N190, N669, N650);
xor XOR2 (N1885, N1879, N1446);
not NOT1 (N1886, N1882);
or OR4 (N1887, N1884, N296, N485, N506);
nor NOR3 (N1888, N1866, N843, N1448);
or OR3 (N1889, N1868, N483, N947);
nand NAND4 (N1890, N1845, N888, N50, N79);
buf BUF1 (N1891, N1885);
or OR3 (N1892, N1891, N1440, N1547);
not NOT1 (N1893, N1852);
and AND2 (N1894, N1888, N1460);
not NOT1 (N1895, N1894);
nand NAND2 (N1896, N1874, N811);
or OR4 (N1897, N1890, N980, N501, N316);
nor NOR2 (N1898, N1892, N1668);
not NOT1 (N1899, N1896);
not NOT1 (N1900, N1886);
not NOT1 (N1901, N1898);
nor NOR4 (N1902, N1895, N929, N512, N647);
nor NOR3 (N1903, N1901, N263, N883);
buf BUF1 (N1904, N1899);
nor NOR3 (N1905, N1902, N1510, N1492);
nand NAND4 (N1906, N1880, N885, N1106, N776);
and AND3 (N1907, N1883, N559, N1799);
not NOT1 (N1908, N1893);
xor XOR2 (N1909, N1907, N1863);
not NOT1 (N1910, N1909);
nand NAND4 (N1911, N1906, N795, N789, N1243);
buf BUF1 (N1912, N1900);
nor NOR4 (N1913, N1905, N1203, N1623, N552);
xor XOR2 (N1914, N1897, N859);
and AND3 (N1915, N1913, N1732, N1015);
or OR2 (N1916, N1912, N1736);
nor NOR2 (N1917, N1916, N525);
nand NAND4 (N1918, N1889, N763, N1249, N1471);
not NOT1 (N1919, N1917);
buf BUF1 (N1920, N1904);
nor NOR4 (N1921, N1919, N521, N1888, N1721);
or OR4 (N1922, N1887, N155, N1734, N773);
nor NOR3 (N1923, N1922, N1101, N1175);
buf BUF1 (N1924, N1920);
and AND3 (N1925, N1918, N1849, N784);
nand NAND2 (N1926, N1925, N937);
buf BUF1 (N1927, N1908);
and AND4 (N1928, N1921, N1189, N1849, N1370);
buf BUF1 (N1929, N1927);
nand NAND3 (N1930, N1926, N1434, N754);
nor NOR4 (N1931, N1928, N497, N215, N1007);
buf BUF1 (N1932, N1930);
nand NAND3 (N1933, N1929, N1621, N362);
nand NAND3 (N1934, N1914, N1771, N194);
xor XOR2 (N1935, N1923, N1042);
or OR3 (N1936, N1915, N953, N512);
xor XOR2 (N1937, N1911, N293);
nor NOR3 (N1938, N1931, N1847, N1745);
buf BUF1 (N1939, N1937);
or OR3 (N1940, N1934, N75, N1835);
or OR4 (N1941, N1903, N633, N291, N1122);
and AND3 (N1942, N1924, N601, N1225);
and AND4 (N1943, N1939, N565, N492, N1288);
or OR3 (N1944, N1933, N1061, N1818);
and AND4 (N1945, N1942, N799, N1759, N1910);
and AND2 (N1946, N1501, N1036);
not NOT1 (N1947, N1938);
xor XOR2 (N1948, N1943, N1021);
and AND3 (N1949, N1936, N1257, N1326);
nor NOR4 (N1950, N1949, N1527, N1263, N1567);
xor XOR2 (N1951, N1935, N1474);
not NOT1 (N1952, N1941);
nor NOR3 (N1953, N1932, N1375, N595);
buf BUF1 (N1954, N1946);
or OR2 (N1955, N1951, N548);
nand NAND2 (N1956, N1953, N854);
or OR3 (N1957, N1948, N621, N1575);
xor XOR2 (N1958, N1954, N347);
buf BUF1 (N1959, N1940);
buf BUF1 (N1960, N1944);
and AND4 (N1961, N1945, N539, N1634, N1762);
buf BUF1 (N1962, N1955);
nor NOR2 (N1963, N1947, N334);
nand NAND4 (N1964, N1962, N1464, N483, N1127);
buf BUF1 (N1965, N1958);
or OR4 (N1966, N1952, N1944, N1917, N1799);
buf BUF1 (N1967, N1957);
buf BUF1 (N1968, N1950);
xor XOR2 (N1969, N1963, N19);
or OR4 (N1970, N1965, N191, N92, N392);
not NOT1 (N1971, N1959);
buf BUF1 (N1972, N1966);
xor XOR2 (N1973, N1956, N1797);
buf BUF1 (N1974, N1972);
nor NOR2 (N1975, N1969, N972);
or OR2 (N1976, N1971, N282);
xor XOR2 (N1977, N1973, N1363);
not NOT1 (N1978, N1975);
nand NAND2 (N1979, N1960, N873);
nand NAND3 (N1980, N1977, N1598, N350);
or OR4 (N1981, N1964, N588, N350, N141);
nand NAND2 (N1982, N1980, N1327);
buf BUF1 (N1983, N1961);
xor XOR2 (N1984, N1983, N1976);
or OR2 (N1985, N937, N1720);
and AND4 (N1986, N1967, N58, N1573, N787);
xor XOR2 (N1987, N1985, N1569);
nor NOR2 (N1988, N1986, N1281);
not NOT1 (N1989, N1978);
nor NOR2 (N1990, N1988, N1663);
xor XOR2 (N1991, N1984, N95);
nor NOR4 (N1992, N1987, N858, N1350, N174);
nor NOR2 (N1993, N1979, N1499);
xor XOR2 (N1994, N1981, N1168);
nand NAND4 (N1995, N1989, N1191, N82, N1694);
nor NOR3 (N1996, N1982, N771, N50);
xor XOR2 (N1997, N1970, N707);
or OR3 (N1998, N1995, N1361, N1703);
and AND2 (N1999, N1992, N1769);
xor XOR2 (N2000, N1974, N39);
nor NOR4 (N2001, N1991, N1585, N1424, N1219);
buf BUF1 (N2002, N1999);
nor NOR3 (N2003, N2001, N1737, N1697);
nor NOR4 (N2004, N1990, N657, N1135, N88);
and AND4 (N2005, N1997, N43, N1908, N870);
not NOT1 (N2006, N1998);
or OR4 (N2007, N1968, N1658, N1530, N708);
nor NOR4 (N2008, N1996, N333, N253, N937);
and AND3 (N2009, N1994, N418, N1604);
nand NAND2 (N2010, N2005, N1921);
or OR3 (N2011, N2000, N386, N1002);
buf BUF1 (N2012, N1993);
buf BUF1 (N2013, N2004);
nand NAND4 (N2014, N2007, N1075, N889, N426);
nand NAND2 (N2015, N2011, N1811);
buf BUF1 (N2016, N2003);
nand NAND3 (N2017, N2008, N1539, N16);
not NOT1 (N2018, N2009);
nor NOR2 (N2019, N2002, N1886);
not NOT1 (N2020, N2019);
not NOT1 (N2021, N2017);
and AND2 (N2022, N2020, N267);
not NOT1 (N2023, N2012);
xor XOR2 (N2024, N2015, N1850);
xor XOR2 (N2025, N2016, N998);
buf BUF1 (N2026, N2022);
and AND4 (N2027, N2018, N1509, N458, N1653);
or OR2 (N2028, N2027, N1346);
nor NOR4 (N2029, N2010, N1602, N1376, N335);
not NOT1 (N2030, N2028);
not NOT1 (N2031, N2025);
buf BUF1 (N2032, N2030);
nor NOR4 (N2033, N2032, N1955, N62, N1603);
nand NAND3 (N2034, N2033, N753, N373);
not NOT1 (N2035, N2006);
xor XOR2 (N2036, N2024, N49);
and AND2 (N2037, N2021, N1745);
xor XOR2 (N2038, N2036, N615);
and AND2 (N2039, N2029, N412);
xor XOR2 (N2040, N2026, N579);
nand NAND4 (N2041, N2034, N712, N646, N1343);
nand NAND3 (N2042, N2014, N1453, N609);
xor XOR2 (N2043, N2023, N1403);
or OR2 (N2044, N2035, N697);
not NOT1 (N2045, N2037);
nand NAND3 (N2046, N2043, N1709, N220);
buf BUF1 (N2047, N2044);
and AND3 (N2048, N2013, N721, N1936);
buf BUF1 (N2049, N2046);
xor XOR2 (N2050, N2038, N1632);
buf BUF1 (N2051, N2047);
xor XOR2 (N2052, N2049, N1268);
and AND4 (N2053, N2040, N1066, N680, N1386);
and AND4 (N2054, N2053, N1682, N391, N1888);
not NOT1 (N2055, N2041);
buf BUF1 (N2056, N2031);
buf BUF1 (N2057, N2045);
or OR3 (N2058, N2039, N1308, N10);
buf BUF1 (N2059, N2054);
buf BUF1 (N2060, N2057);
and AND3 (N2061, N2059, N1085, N1053);
xor XOR2 (N2062, N2055, N1664);
xor XOR2 (N2063, N2050, N1590);
xor XOR2 (N2064, N2048, N1330);
or OR2 (N2065, N2056, N1002);
nand NAND2 (N2066, N2062, N272);
or OR4 (N2067, N2042, N643, N814, N1071);
nand NAND2 (N2068, N2052, N1073);
buf BUF1 (N2069, N2064);
or OR4 (N2070, N2069, N461, N1690, N1950);
nor NOR3 (N2071, N2051, N487, N885);
xor XOR2 (N2072, N2058, N506);
xor XOR2 (N2073, N2066, N518);
xor XOR2 (N2074, N2073, N371);
not NOT1 (N2075, N2060);
and AND3 (N2076, N2072, N1865, N1652);
nor NOR3 (N2077, N2068, N315, N2061);
buf BUF1 (N2078, N1410);
xor XOR2 (N2079, N2078, N1470);
buf BUF1 (N2080, N2075);
nor NOR3 (N2081, N2074, N71, N538);
or OR3 (N2082, N2076, N893, N765);
nand NAND3 (N2083, N2070, N543, N1414);
or OR4 (N2084, N2079, N544, N830, N2018);
nor NOR2 (N2085, N2063, N1740);
nand NAND2 (N2086, N2083, N821);
or OR2 (N2087, N2084, N1756);
or OR2 (N2088, N2082, N628);
not NOT1 (N2089, N2085);
nand NAND2 (N2090, N2080, N718);
and AND3 (N2091, N2071, N367, N1074);
and AND3 (N2092, N2089, N952, N272);
nor NOR4 (N2093, N2067, N53, N285, N2043);
and AND2 (N2094, N2092, N1918);
or OR2 (N2095, N2077, N681);
and AND3 (N2096, N2091, N1884, N1770);
xor XOR2 (N2097, N2096, N1591);
xor XOR2 (N2098, N2097, N667);
not NOT1 (N2099, N2098);
nor NOR4 (N2100, N2090, N1554, N608, N2034);
xor XOR2 (N2101, N2081, N1675);
nand NAND2 (N2102, N2088, N148);
xor XOR2 (N2103, N2102, N1528);
nor NOR2 (N2104, N2099, N1909);
nand NAND4 (N2105, N2093, N605, N603, N1306);
and AND4 (N2106, N2095, N624, N1810, N1147);
xor XOR2 (N2107, N2103, N1027);
or OR4 (N2108, N2106, N1219, N1798, N852);
xor XOR2 (N2109, N2100, N725);
and AND4 (N2110, N2101, N999, N209, N388);
and AND3 (N2111, N2087, N1963, N891);
nor NOR2 (N2112, N2110, N33);
nor NOR2 (N2113, N2107, N84);
or OR4 (N2114, N2094, N283, N1775, N1363);
nor NOR2 (N2115, N2114, N971);
nand NAND4 (N2116, N2086, N1956, N489, N1984);
and AND2 (N2117, N2112, N913);
or OR3 (N2118, N2116, N146, N1413);
and AND4 (N2119, N2065, N55, N910, N1852);
nor NOR3 (N2120, N2119, N1796, N1692);
xor XOR2 (N2121, N2117, N967);
xor XOR2 (N2122, N2109, N260);
nor NOR4 (N2123, N2105, N361, N458, N1713);
or OR2 (N2124, N2108, N625);
xor XOR2 (N2125, N2104, N529);
nand NAND2 (N2126, N2124, N1086);
nor NOR3 (N2127, N2120, N1957, N1461);
not NOT1 (N2128, N2118);
nor NOR3 (N2129, N2113, N1031, N658);
xor XOR2 (N2130, N2122, N2042);
and AND2 (N2131, N2123, N550);
buf BUF1 (N2132, N2128);
or OR4 (N2133, N2115, N675, N661, N427);
and AND2 (N2134, N2111, N957);
or OR2 (N2135, N2129, N2003);
nand NAND2 (N2136, N2126, N797);
nor NOR4 (N2137, N2133, N882, N699, N1408);
nand NAND4 (N2138, N2135, N1509, N1942, N173);
nand NAND4 (N2139, N2134, N652, N1386, N913);
and AND4 (N2140, N2136, N921, N1096, N1758);
or OR2 (N2141, N2121, N1135);
xor XOR2 (N2142, N2131, N1220);
xor XOR2 (N2143, N2141, N916);
and AND4 (N2144, N2127, N1206, N944, N149);
and AND3 (N2145, N2140, N476, N1466);
buf BUF1 (N2146, N2125);
xor XOR2 (N2147, N2144, N1207);
not NOT1 (N2148, N2137);
nand NAND2 (N2149, N2143, N793);
nand NAND4 (N2150, N2146, N646, N1306, N982);
nand NAND3 (N2151, N2139, N712, N1734);
xor XOR2 (N2152, N2149, N650);
nand NAND2 (N2153, N2150, N528);
not NOT1 (N2154, N2148);
xor XOR2 (N2155, N2142, N299);
not NOT1 (N2156, N2154);
not NOT1 (N2157, N2138);
xor XOR2 (N2158, N2132, N847);
nor NOR3 (N2159, N2158, N2048, N363);
or OR3 (N2160, N2130, N998, N1901);
not NOT1 (N2161, N2147);
nand NAND3 (N2162, N2145, N2092, N283);
and AND2 (N2163, N2151, N1531);
not NOT1 (N2164, N2161);
and AND4 (N2165, N2160, N1211, N832, N189);
or OR4 (N2166, N2162, N189, N1461, N325);
not NOT1 (N2167, N2166);
buf BUF1 (N2168, N2156);
nand NAND4 (N2169, N2159, N1074, N1198, N307);
or OR2 (N2170, N2167, N121);
or OR4 (N2171, N2155, N149, N1095, N1544);
xor XOR2 (N2172, N2165, N1149);
nand NAND4 (N2173, N2170, N1263, N1901, N804);
not NOT1 (N2174, N2172);
and AND3 (N2175, N2152, N1205, N1418);
or OR2 (N2176, N2163, N583);
not NOT1 (N2177, N2157);
xor XOR2 (N2178, N2153, N778);
buf BUF1 (N2179, N2175);
and AND3 (N2180, N2179, N636, N1126);
not NOT1 (N2181, N2177);
or OR3 (N2182, N2174, N112, N271);
buf BUF1 (N2183, N2164);
buf BUF1 (N2184, N2182);
xor XOR2 (N2185, N2176, N1039);
buf BUF1 (N2186, N2171);
not NOT1 (N2187, N2168);
buf BUF1 (N2188, N2173);
or OR2 (N2189, N2183, N1931);
nand NAND4 (N2190, N2181, N2102, N683, N1170);
xor XOR2 (N2191, N2184, N1452);
nand NAND4 (N2192, N2187, N226, N1538, N2177);
buf BUF1 (N2193, N2188);
nor NOR3 (N2194, N2189, N2157, N1499);
or OR4 (N2195, N2192, N554, N760, N1210);
nor NOR4 (N2196, N2185, N206, N854, N569);
not NOT1 (N2197, N2191);
not NOT1 (N2198, N2194);
not NOT1 (N2199, N2186);
xor XOR2 (N2200, N2169, N1161);
nand NAND3 (N2201, N2197, N1878, N1093);
nor NOR4 (N2202, N2195, N1516, N926, N602);
xor XOR2 (N2203, N2202, N67);
buf BUF1 (N2204, N2198);
buf BUF1 (N2205, N2204);
and AND3 (N2206, N2180, N1120, N1333);
and AND2 (N2207, N2193, N423);
nand NAND3 (N2208, N2178, N2160, N1814);
xor XOR2 (N2209, N2200, N830);
nand NAND2 (N2210, N2207, N1004);
or OR2 (N2211, N2196, N1393);
xor XOR2 (N2212, N2208, N1217);
not NOT1 (N2213, N2201);
xor XOR2 (N2214, N2190, N2003);
nor NOR4 (N2215, N2203, N683, N941, N2202);
not NOT1 (N2216, N2212);
nand NAND4 (N2217, N2205, N1668, N399, N774);
xor XOR2 (N2218, N2216, N1280);
or OR3 (N2219, N2210, N38, N523);
buf BUF1 (N2220, N2199);
or OR2 (N2221, N2209, N1881);
or OR2 (N2222, N2219, N49);
or OR2 (N2223, N2214, N2020);
not NOT1 (N2224, N2220);
and AND3 (N2225, N2211, N344, N2136);
and AND3 (N2226, N2223, N409, N702);
or OR2 (N2227, N2226, N639);
nand NAND3 (N2228, N2215, N327, N1050);
and AND4 (N2229, N2206, N372, N1236, N2083);
buf BUF1 (N2230, N2224);
nor NOR4 (N2231, N2217, N1151, N1360, N1687);
xor XOR2 (N2232, N2222, N1160);
nand NAND2 (N2233, N2228, N1462);
xor XOR2 (N2234, N2232, N2063);
not NOT1 (N2235, N2225);
nor NOR3 (N2236, N2213, N547, N894);
buf BUF1 (N2237, N2231);
and AND4 (N2238, N2229, N915, N1490, N1418);
buf BUF1 (N2239, N2233);
and AND2 (N2240, N2235, N929);
xor XOR2 (N2241, N2237, N1618);
or OR2 (N2242, N2236, N250);
or OR2 (N2243, N2227, N686);
or OR4 (N2244, N2230, N1723, N701, N631);
or OR2 (N2245, N2238, N1846);
buf BUF1 (N2246, N2239);
not NOT1 (N2247, N2246);
and AND4 (N2248, N2245, N1624, N141, N985);
not NOT1 (N2249, N2247);
nor NOR4 (N2250, N2242, N1960, N1283, N735);
xor XOR2 (N2251, N2250, N661);
or OR4 (N2252, N2221, N594, N711, N2173);
or OR2 (N2253, N2234, N1510);
nand NAND4 (N2254, N2252, N1662, N153, N784);
nor NOR4 (N2255, N2244, N314, N2101, N1509);
buf BUF1 (N2256, N2218);
not NOT1 (N2257, N2251);
or OR3 (N2258, N2254, N1515, N463);
nor NOR3 (N2259, N2243, N1581, N1797);
and AND4 (N2260, N2249, N88, N2038, N971);
nand NAND3 (N2261, N2259, N399, N326);
or OR4 (N2262, N2258, N1697, N742, N118);
buf BUF1 (N2263, N2262);
or OR4 (N2264, N2260, N1812, N141, N1587);
and AND3 (N2265, N2253, N415, N2155);
or OR3 (N2266, N2265, N1415, N1364);
and AND2 (N2267, N2263, N802);
and AND4 (N2268, N2267, N428, N1855, N1634);
not NOT1 (N2269, N2256);
nor NOR4 (N2270, N2261, N2142, N1857, N1414);
xor XOR2 (N2271, N2241, N1823);
or OR2 (N2272, N2270, N1351);
xor XOR2 (N2273, N2269, N1742);
and AND3 (N2274, N2264, N1174, N339);
buf BUF1 (N2275, N2268);
nor NOR4 (N2276, N2240, N953, N139, N1832);
xor XOR2 (N2277, N2274, N1853);
not NOT1 (N2278, N2273);
nor NOR4 (N2279, N2257, N922, N1379, N1504);
buf BUF1 (N2280, N2276);
buf BUF1 (N2281, N2278);
xor XOR2 (N2282, N2275, N1460);
not NOT1 (N2283, N2271);
nand NAND3 (N2284, N2280, N2206, N1913);
or OR2 (N2285, N2281, N2137);
or OR2 (N2286, N2277, N876);
nand NAND3 (N2287, N2286, N1969, N2231);
not NOT1 (N2288, N2282);
not NOT1 (N2289, N2287);
and AND2 (N2290, N2285, N1477);
xor XOR2 (N2291, N2266, N758);
nand NAND3 (N2292, N2279, N2186, N2089);
and AND2 (N2293, N2283, N395);
nand NAND3 (N2294, N2289, N2224, N711);
nand NAND4 (N2295, N2284, N680, N716, N551);
or OR4 (N2296, N2294, N1935, N1170, N20);
buf BUF1 (N2297, N2272);
xor XOR2 (N2298, N2290, N1928);
buf BUF1 (N2299, N2295);
nor NOR3 (N2300, N2298, N1098, N1304);
or OR2 (N2301, N2255, N101);
and AND4 (N2302, N2248, N1829, N1017, N842);
nand NAND2 (N2303, N2301, N2021);
nand NAND2 (N2304, N2299, N63);
nand NAND2 (N2305, N2296, N665);
nand NAND4 (N2306, N2293, N315, N992, N203);
nor NOR3 (N2307, N2291, N1855, N239);
or OR2 (N2308, N2297, N1061);
buf BUF1 (N2309, N2305);
nor NOR3 (N2310, N2306, N1903, N554);
and AND2 (N2311, N2300, N1152);
and AND3 (N2312, N2311, N1779, N1982);
xor XOR2 (N2313, N2302, N1101);
and AND2 (N2314, N2307, N2022);
buf BUF1 (N2315, N2303);
not NOT1 (N2316, N2314);
buf BUF1 (N2317, N2288);
or OR3 (N2318, N2308, N1791, N1800);
xor XOR2 (N2319, N2310, N314);
and AND3 (N2320, N2315, N1813, N661);
nand NAND4 (N2321, N2316, N969, N487, N693);
or OR2 (N2322, N2309, N1373);
not NOT1 (N2323, N2318);
not NOT1 (N2324, N2292);
xor XOR2 (N2325, N2312, N392);
nor NOR3 (N2326, N2321, N1943, N821);
or OR3 (N2327, N2323, N988, N1076);
and AND2 (N2328, N2304, N2258);
buf BUF1 (N2329, N2325);
buf BUF1 (N2330, N2319);
or OR3 (N2331, N2329, N1452, N786);
and AND3 (N2332, N2324, N367, N401);
and AND2 (N2333, N2332, N1820);
nand NAND4 (N2334, N2320, N1887, N1838, N2058);
or OR4 (N2335, N2330, N866, N681, N493);
not NOT1 (N2336, N2317);
and AND2 (N2337, N2335, N2152);
buf BUF1 (N2338, N2313);
not NOT1 (N2339, N2327);
xor XOR2 (N2340, N2337, N1418);
nand NAND4 (N2341, N2328, N1703, N953, N1073);
nand NAND2 (N2342, N2334, N675);
or OR3 (N2343, N2341, N1175, N2022);
or OR3 (N2344, N2326, N1419, N1466);
xor XOR2 (N2345, N2331, N2308);
xor XOR2 (N2346, N2342, N25);
buf BUF1 (N2347, N2346);
or OR4 (N2348, N2333, N88, N44, N1886);
and AND3 (N2349, N2347, N2111, N1840);
nor NOR2 (N2350, N2343, N587);
buf BUF1 (N2351, N2348);
not NOT1 (N2352, N2338);
and AND2 (N2353, N2340, N646);
or OR2 (N2354, N2322, N1378);
buf BUF1 (N2355, N2354);
not NOT1 (N2356, N2352);
not NOT1 (N2357, N2349);
and AND2 (N2358, N2336, N859);
nand NAND4 (N2359, N2351, N414, N2160, N1639);
nand NAND3 (N2360, N2356, N2307, N1383);
or OR3 (N2361, N2353, N1369, N746);
nor NOR3 (N2362, N2344, N855, N76);
nor NOR2 (N2363, N2345, N1700);
and AND2 (N2364, N2360, N1383);
nor NOR4 (N2365, N2355, N481, N422, N1381);
buf BUF1 (N2366, N2359);
xor XOR2 (N2367, N2364, N428);
xor XOR2 (N2368, N2365, N2238);
not NOT1 (N2369, N2362);
or OR4 (N2370, N2366, N817, N1232, N1517);
not NOT1 (N2371, N2370);
xor XOR2 (N2372, N2368, N1093);
or OR2 (N2373, N2350, N1043);
nor NOR2 (N2374, N2372, N1412);
or OR2 (N2375, N2369, N1884);
or OR4 (N2376, N2371, N1077, N2084, N1579);
nand NAND4 (N2377, N2363, N735, N2268, N788);
or OR3 (N2378, N2339, N579, N1451);
nor NOR2 (N2379, N2358, N1676);
buf BUF1 (N2380, N2374);
nor NOR3 (N2381, N2378, N762, N2268);
not NOT1 (N2382, N2367);
nand NAND3 (N2383, N2382, N1497, N1612);
or OR2 (N2384, N2383, N1773);
or OR3 (N2385, N2375, N158, N1555);
xor XOR2 (N2386, N2384, N1242);
or OR2 (N2387, N2380, N1756);
not NOT1 (N2388, N2373);
and AND2 (N2389, N2376, N2363);
xor XOR2 (N2390, N2385, N2328);
xor XOR2 (N2391, N2377, N1953);
nor NOR2 (N2392, N2390, N260);
or OR3 (N2393, N2357, N860, N2187);
or OR4 (N2394, N2392, N817, N264, N613);
or OR3 (N2395, N2393, N245, N759);
and AND4 (N2396, N2386, N177, N1395, N347);
nor NOR4 (N2397, N2387, N2307, N1034, N639);
not NOT1 (N2398, N2394);
buf BUF1 (N2399, N2361);
or OR2 (N2400, N2381, N321);
or OR4 (N2401, N2389, N900, N621, N2237);
xor XOR2 (N2402, N2400, N1814);
nand NAND3 (N2403, N2396, N296, N2388);
and AND4 (N2404, N2092, N2307, N56, N770);
buf BUF1 (N2405, N2398);
buf BUF1 (N2406, N2404);
not NOT1 (N2407, N2401);
and AND2 (N2408, N2399, N1035);
xor XOR2 (N2409, N2406, N2395);
or OR4 (N2410, N916, N22, N1772, N89);
nand NAND2 (N2411, N2397, N1425);
or OR4 (N2412, N2408, N433, N241, N2197);
not NOT1 (N2413, N2405);
nor NOR4 (N2414, N2409, N1218, N967, N954);
or OR3 (N2415, N2379, N2196, N2374);
and AND2 (N2416, N2410, N1980);
not NOT1 (N2417, N2411);
or OR2 (N2418, N2417, N1987);
xor XOR2 (N2419, N2391, N879);
not NOT1 (N2420, N2419);
nor NOR2 (N2421, N2415, N2361);
nor NOR4 (N2422, N2402, N1611, N413, N1059);
xor XOR2 (N2423, N2420, N1367);
buf BUF1 (N2424, N2421);
not NOT1 (N2425, N2423);
or OR3 (N2426, N2414, N310, N685);
not NOT1 (N2427, N2425);
buf BUF1 (N2428, N2427);
buf BUF1 (N2429, N2412);
or OR2 (N2430, N2429, N2367);
or OR4 (N2431, N2430, N121, N2080, N1899);
xor XOR2 (N2432, N2403, N1699);
not NOT1 (N2433, N2428);
buf BUF1 (N2434, N2433);
buf BUF1 (N2435, N2432);
or OR4 (N2436, N2407, N587, N1167, N1873);
nor NOR2 (N2437, N2424, N1560);
and AND3 (N2438, N2435, N1055, N2031);
nor NOR3 (N2439, N2426, N1380, N363);
or OR3 (N2440, N2437, N1898, N1878);
nor NOR2 (N2441, N2438, N1863);
and AND3 (N2442, N2436, N752, N1261);
and AND2 (N2443, N2441, N337);
xor XOR2 (N2444, N2413, N1178);
not NOT1 (N2445, N2416);
not NOT1 (N2446, N2442);
not NOT1 (N2447, N2439);
nor NOR4 (N2448, N2443, N2069, N497, N96);
not NOT1 (N2449, N2448);
buf BUF1 (N2450, N2445);
nor NOR4 (N2451, N2450, N1096, N1749, N2068);
nand NAND4 (N2452, N2444, N2341, N588, N864);
or OR4 (N2453, N2434, N502, N160, N2144);
or OR2 (N2454, N2431, N2350);
nand NAND3 (N2455, N2449, N17, N1390);
nor NOR3 (N2456, N2455, N858, N219);
buf BUF1 (N2457, N2454);
not NOT1 (N2458, N2451);
or OR3 (N2459, N2422, N86, N678);
not NOT1 (N2460, N2457);
xor XOR2 (N2461, N2446, N1415);
xor XOR2 (N2462, N2447, N152);
nand NAND3 (N2463, N2452, N1026, N1376);
xor XOR2 (N2464, N2459, N413);
and AND2 (N2465, N2440, N1362);
or OR2 (N2466, N2418, N36);
not NOT1 (N2467, N2462);
xor XOR2 (N2468, N2461, N1027);
xor XOR2 (N2469, N2458, N149);
nand NAND3 (N2470, N2463, N2467, N1676);
buf BUF1 (N2471, N1045);
buf BUF1 (N2472, N2466);
nor NOR4 (N2473, N2456, N1787, N2414, N1810);
xor XOR2 (N2474, N2473, N1562);
or OR3 (N2475, N2474, N2409, N2124);
buf BUF1 (N2476, N2460);
nor NOR2 (N2477, N2476, N1914);
or OR2 (N2478, N2472, N987);
or OR2 (N2479, N2475, N161);
not NOT1 (N2480, N2471);
buf BUF1 (N2481, N2477);
not NOT1 (N2482, N2453);
or OR2 (N2483, N2469, N722);
or OR4 (N2484, N2468, N1609, N1821, N995);
nor NOR3 (N2485, N2483, N2368, N932);
not NOT1 (N2486, N2484);
buf BUF1 (N2487, N2480);
buf BUF1 (N2488, N2479);
xor XOR2 (N2489, N2478, N1100);
buf BUF1 (N2490, N2487);
or OR3 (N2491, N2464, N1133, N527);
or OR4 (N2492, N2482, N22, N650, N525);
nand NAND3 (N2493, N2491, N297, N1461);
not NOT1 (N2494, N2490);
and AND4 (N2495, N2492, N212, N92, N2097);
and AND3 (N2496, N2489, N883, N1170);
xor XOR2 (N2497, N2485, N1540);
or OR3 (N2498, N2497, N395, N521);
nor NOR4 (N2499, N2465, N2318, N2449, N728);
nor NOR3 (N2500, N2498, N2048, N449);
not NOT1 (N2501, N2470);
and AND2 (N2502, N2500, N594);
not NOT1 (N2503, N2496);
buf BUF1 (N2504, N2495);
or OR3 (N2505, N2481, N1458, N1684);
nor NOR3 (N2506, N2501, N447, N2336);
nand NAND4 (N2507, N2503, N728, N480, N1313);
xor XOR2 (N2508, N2488, N506);
and AND4 (N2509, N2502, N81, N671, N543);
buf BUF1 (N2510, N2507);
nand NAND2 (N2511, N2499, N2424);
not NOT1 (N2512, N2506);
and AND4 (N2513, N2508, N720, N1170, N1612);
nor NOR4 (N2514, N2494, N1795, N344, N1583);
and AND3 (N2515, N2510, N597, N1833);
nand NAND4 (N2516, N2486, N1290, N1482, N2170);
buf BUF1 (N2517, N2512);
nand NAND3 (N2518, N2514, N1451, N1846);
and AND4 (N2519, N2517, N200, N2448, N1369);
xor XOR2 (N2520, N2516, N2239);
nand NAND3 (N2521, N2520, N1728, N364);
and AND3 (N2522, N2504, N639, N2391);
or OR4 (N2523, N2519, N1521, N183, N827);
xor XOR2 (N2524, N2493, N37);
and AND2 (N2525, N2523, N1028);
not NOT1 (N2526, N2509);
nand NAND2 (N2527, N2511, N369);
xor XOR2 (N2528, N2505, N2223);
buf BUF1 (N2529, N2524);
and AND2 (N2530, N2525, N1488);
not NOT1 (N2531, N2518);
nor NOR4 (N2532, N2531, N671, N313, N1006);
nor NOR4 (N2533, N2521, N1360, N2185, N441);
buf BUF1 (N2534, N2513);
nor NOR2 (N2535, N2522, N386);
nor NOR3 (N2536, N2535, N155, N1506);
or OR2 (N2537, N2536, N672);
and AND2 (N2538, N2534, N443);
not NOT1 (N2539, N2532);
not NOT1 (N2540, N2526);
and AND2 (N2541, N2537, N1022);
nand NAND3 (N2542, N2530, N2215, N2200);
nor NOR4 (N2543, N2529, N1901, N1078, N2236);
and AND3 (N2544, N2527, N841, N1062);
or OR4 (N2545, N2533, N655, N2063, N447);
nor NOR3 (N2546, N2540, N2517, N964);
or OR4 (N2547, N2528, N898, N328, N6);
buf BUF1 (N2548, N2542);
xor XOR2 (N2549, N2538, N2454);
and AND2 (N2550, N2515, N574);
and AND2 (N2551, N2539, N1453);
or OR2 (N2552, N2544, N1107);
xor XOR2 (N2553, N2550, N1312);
nor NOR2 (N2554, N2551, N1959);
and AND4 (N2555, N2541, N1537, N1902, N1662);
and AND3 (N2556, N2547, N1940, N1488);
nand NAND3 (N2557, N2553, N1412, N66);
and AND2 (N2558, N2554, N567);
or OR2 (N2559, N2552, N2143);
not NOT1 (N2560, N2558);
nor NOR3 (N2561, N2559, N542, N261);
nor NOR4 (N2562, N2543, N1253, N2528, N1185);
and AND2 (N2563, N2556, N2071);
or OR3 (N2564, N2555, N968, N337);
buf BUF1 (N2565, N2562);
xor XOR2 (N2566, N2548, N1202);
and AND2 (N2567, N2564, N337);
buf BUF1 (N2568, N2557);
nand NAND4 (N2569, N2566, N481, N2330, N322);
buf BUF1 (N2570, N2567);
and AND2 (N2571, N2561, N1889);
buf BUF1 (N2572, N2545);
nor NOR4 (N2573, N2568, N1848, N2102, N2250);
nand NAND4 (N2574, N2565, N770, N2000, N1582);
xor XOR2 (N2575, N2574, N1469);
buf BUF1 (N2576, N2549);
xor XOR2 (N2577, N2575, N119);
buf BUF1 (N2578, N2576);
not NOT1 (N2579, N2560);
not NOT1 (N2580, N2571);
or OR3 (N2581, N2579, N2076, N69);
buf BUF1 (N2582, N2572);
or OR2 (N2583, N2573, N140);
xor XOR2 (N2584, N2583, N900);
not NOT1 (N2585, N2570);
nand NAND3 (N2586, N2546, N1009, N2270);
nand NAND4 (N2587, N2585, N1889, N2036, N869);
nor NOR2 (N2588, N2580, N2487);
or OR3 (N2589, N2578, N2104, N1770);
nor NOR3 (N2590, N2586, N2368, N1779);
xor XOR2 (N2591, N2582, N260);
buf BUF1 (N2592, N2569);
not NOT1 (N2593, N2590);
nand NAND4 (N2594, N2584, N1989, N1402, N649);
not NOT1 (N2595, N2593);
buf BUF1 (N2596, N2588);
nor NOR3 (N2597, N2581, N1017, N2416);
not NOT1 (N2598, N2589);
nand NAND3 (N2599, N2597, N1212, N1361);
xor XOR2 (N2600, N2577, N1783);
nand NAND3 (N2601, N2596, N2048, N1997);
buf BUF1 (N2602, N2601);
buf BUF1 (N2603, N2595);
nor NOR3 (N2604, N2594, N2429, N780);
nor NOR3 (N2605, N2587, N2245, N2465);
xor XOR2 (N2606, N2598, N1620);
xor XOR2 (N2607, N2591, N2276);
nor NOR3 (N2608, N2604, N1354, N218);
nor NOR3 (N2609, N2563, N1570, N1943);
nor NOR2 (N2610, N2603, N1878);
and AND3 (N2611, N2606, N52, N2420);
xor XOR2 (N2612, N2610, N1909);
not NOT1 (N2613, N2608);
xor XOR2 (N2614, N2613, N252);
nor NOR3 (N2615, N2599, N118, N1242);
buf BUF1 (N2616, N2600);
nor NOR3 (N2617, N2602, N406, N2303);
nand NAND3 (N2618, N2615, N2086, N2541);
or OR2 (N2619, N2592, N2578);
nor NOR2 (N2620, N2616, N307);
not NOT1 (N2621, N2612);
not NOT1 (N2622, N2605);
buf BUF1 (N2623, N2621);
or OR4 (N2624, N2607, N1085, N1603, N474);
xor XOR2 (N2625, N2622, N1328);
and AND4 (N2626, N2617, N1099, N2337, N1635);
buf BUF1 (N2627, N2623);
not NOT1 (N2628, N2626);
xor XOR2 (N2629, N2628, N2091);
nor NOR4 (N2630, N2614, N1469, N1692, N918);
xor XOR2 (N2631, N2620, N681);
nor NOR4 (N2632, N2624, N95, N2093, N2222);
or OR3 (N2633, N2611, N407, N2259);
nor NOR2 (N2634, N2630, N2416);
nor NOR4 (N2635, N2633, N2476, N1873, N973);
or OR3 (N2636, N2618, N643, N104);
nor NOR2 (N2637, N2625, N83);
buf BUF1 (N2638, N2609);
not NOT1 (N2639, N2627);
or OR3 (N2640, N2635, N535, N1421);
not NOT1 (N2641, N2631);
xor XOR2 (N2642, N2641, N802);
nor NOR4 (N2643, N2636, N2286, N2580, N1410);
buf BUF1 (N2644, N2638);
xor XOR2 (N2645, N2619, N2487);
nand NAND3 (N2646, N2629, N1495, N537);
buf BUF1 (N2647, N2645);
nand NAND2 (N2648, N2637, N157);
xor XOR2 (N2649, N2646, N1927);
buf BUF1 (N2650, N2634);
xor XOR2 (N2651, N2632, N2467);
not NOT1 (N2652, N2651);
nor NOR4 (N2653, N2640, N2168, N363, N436);
nand NAND2 (N2654, N2642, N1008);
and AND3 (N2655, N2647, N2449, N439);
or OR4 (N2656, N2649, N1370, N2109, N2591);
nor NOR2 (N2657, N2639, N2537);
not NOT1 (N2658, N2650);
and AND4 (N2659, N2653, N2586, N1999, N703);
not NOT1 (N2660, N2644);
or OR4 (N2661, N2657, N2351, N1377, N90);
or OR2 (N2662, N2648, N961);
or OR2 (N2663, N2658, N757);
not NOT1 (N2664, N2659);
buf BUF1 (N2665, N2654);
and AND2 (N2666, N2660, N1343);
and AND2 (N2667, N2665, N467);
and AND4 (N2668, N2664, N415, N1778, N795);
nor NOR2 (N2669, N2652, N1020);
nor NOR2 (N2670, N2656, N1560);
nor NOR4 (N2671, N2661, N1191, N1697, N2607);
nor NOR4 (N2672, N2662, N2650, N1995, N218);
or OR4 (N2673, N2655, N1376, N1667, N1028);
or OR4 (N2674, N2672, N2647, N2561, N761);
buf BUF1 (N2675, N2673);
and AND2 (N2676, N2671, N643);
not NOT1 (N2677, N2675);
xor XOR2 (N2678, N2676, N478);
not NOT1 (N2679, N2677);
or OR3 (N2680, N2643, N1261, N525);
or OR3 (N2681, N2678, N2083, N2018);
xor XOR2 (N2682, N2680, N1994);
buf BUF1 (N2683, N2679);
nor NOR3 (N2684, N2682, N608, N543);
xor XOR2 (N2685, N2681, N1991);
and AND4 (N2686, N2683, N290, N660, N97);
nand NAND3 (N2687, N2684, N989, N1693);
nand NAND2 (N2688, N2669, N2380);
nand NAND3 (N2689, N2674, N896, N2595);
buf BUF1 (N2690, N2663);
and AND2 (N2691, N2690, N448);
and AND3 (N2692, N2667, N324, N2056);
buf BUF1 (N2693, N2670);
or OR2 (N2694, N2693, N738);
and AND4 (N2695, N2688, N2196, N2379, N1791);
xor XOR2 (N2696, N2685, N2486);
not NOT1 (N2697, N2668);
or OR4 (N2698, N2691, N295, N731, N35);
or OR3 (N2699, N2687, N383, N768);
nor NOR2 (N2700, N2694, N612);
buf BUF1 (N2701, N2698);
and AND4 (N2702, N2686, N2026, N1447, N1333);
buf BUF1 (N2703, N2702);
not NOT1 (N2704, N2703);
xor XOR2 (N2705, N2700, N2423);
nand NAND4 (N2706, N2704, N1130, N844, N462);
or OR3 (N2707, N2666, N706, N1618);
buf BUF1 (N2708, N2697);
xor XOR2 (N2709, N2708, N1355);
nor NOR3 (N2710, N2699, N440, N799);
not NOT1 (N2711, N2707);
nor NOR3 (N2712, N2696, N432, N478);
nor NOR3 (N2713, N2706, N368, N1255);
not NOT1 (N2714, N2701);
and AND3 (N2715, N2689, N2473, N2216);
not NOT1 (N2716, N2712);
xor XOR2 (N2717, N2715, N1459);
buf BUF1 (N2718, N2717);
buf BUF1 (N2719, N2711);
nor NOR2 (N2720, N2705, N2157);
nand NAND4 (N2721, N2719, N2048, N1402, N1801);
nor NOR3 (N2722, N2692, N1026, N2663);
buf BUF1 (N2723, N2720);
and AND3 (N2724, N2722, N892, N1709);
nor NOR3 (N2725, N2710, N803, N205);
and AND3 (N2726, N2716, N2304, N1890);
buf BUF1 (N2727, N2725);
not NOT1 (N2728, N2713);
and AND2 (N2729, N2718, N2345);
nor NOR2 (N2730, N2721, N2441);
nor NOR2 (N2731, N2695, N1257);
not NOT1 (N2732, N2730);
or OR3 (N2733, N2724, N791, N2170);
and AND3 (N2734, N2733, N1380, N757);
and AND2 (N2735, N2727, N1268);
nand NAND2 (N2736, N2732, N107);
nand NAND3 (N2737, N2709, N918, N452);
buf BUF1 (N2738, N2728);
or OR3 (N2739, N2723, N975, N1171);
and AND4 (N2740, N2731, N1108, N476, N2368);
buf BUF1 (N2741, N2726);
or OR3 (N2742, N2737, N300, N1153);
or OR4 (N2743, N2741, N439, N1212, N940);
buf BUF1 (N2744, N2743);
not NOT1 (N2745, N2714);
and AND3 (N2746, N2739, N399, N2743);
not NOT1 (N2747, N2746);
not NOT1 (N2748, N2735);
nand NAND4 (N2749, N2745, N885, N95, N2528);
nor NOR3 (N2750, N2729, N1831, N1272);
nand NAND4 (N2751, N2738, N730, N1227, N2243);
and AND2 (N2752, N2736, N2509);
not NOT1 (N2753, N2749);
nand NAND4 (N2754, N2748, N576, N2283, N2137);
not NOT1 (N2755, N2734);
not NOT1 (N2756, N2740);
xor XOR2 (N2757, N2753, N1449);
nor NOR2 (N2758, N2752, N1791);
or OR4 (N2759, N2744, N1543, N1939, N166);
nand NAND2 (N2760, N2751, N2019);
nor NOR3 (N2761, N2754, N807, N592);
nand NAND2 (N2762, N2756, N299);
nor NOR4 (N2763, N2761, N1564, N1081, N1726);
xor XOR2 (N2764, N2763, N2479);
nor NOR4 (N2765, N2758, N2005, N838, N2503);
not NOT1 (N2766, N2750);
nor NOR4 (N2767, N2766, N1205, N667, N2263);
nand NAND3 (N2768, N2764, N2465, N2464);
nand NAND2 (N2769, N2759, N1855);
buf BUF1 (N2770, N2757);
buf BUF1 (N2771, N2767);
xor XOR2 (N2772, N2765, N42);
not NOT1 (N2773, N2768);
or OR4 (N2774, N2772, N2705, N893, N2274);
nand NAND4 (N2775, N2742, N1571, N555, N1917);
nor NOR2 (N2776, N2771, N107);
buf BUF1 (N2777, N2770);
or OR3 (N2778, N2777, N1334, N1614);
buf BUF1 (N2779, N2775);
and AND3 (N2780, N2776, N854, N2035);
xor XOR2 (N2781, N2779, N2331);
nor NOR2 (N2782, N2760, N2674);
nand NAND3 (N2783, N2782, N627, N1572);
nor NOR2 (N2784, N2783, N2509);
buf BUF1 (N2785, N2747);
nor NOR2 (N2786, N2781, N2300);
or OR3 (N2787, N2784, N11, N1206);
or OR2 (N2788, N2755, N2627);
or OR2 (N2789, N2774, N149);
or OR2 (N2790, N2778, N723);
not NOT1 (N2791, N2780);
buf BUF1 (N2792, N2787);
buf BUF1 (N2793, N2792);
buf BUF1 (N2794, N2788);
nand NAND4 (N2795, N2793, N1539, N1750, N692);
or OR4 (N2796, N2791, N610, N1785, N773);
or OR3 (N2797, N2769, N2708, N2250);
nor NOR2 (N2798, N2796, N1776);
not NOT1 (N2799, N2797);
xor XOR2 (N2800, N2762, N1474);
and AND2 (N2801, N2790, N2640);
nor NOR2 (N2802, N2800, N2033);
not NOT1 (N2803, N2785);
buf BUF1 (N2804, N2786);
nand NAND4 (N2805, N2801, N965, N1723, N1202);
and AND4 (N2806, N2803, N1379, N654, N1701);
buf BUF1 (N2807, N2773);
not NOT1 (N2808, N2806);
and AND3 (N2809, N2794, N553, N2692);
nand NAND3 (N2810, N2805, N2274, N2766);
xor XOR2 (N2811, N2798, N960);
or OR3 (N2812, N2802, N1087, N484);
nor NOR4 (N2813, N2795, N992, N614, N1941);
xor XOR2 (N2814, N2811, N2272);
buf BUF1 (N2815, N2813);
xor XOR2 (N2816, N2807, N450);
and AND4 (N2817, N2808, N164, N362, N2736);
nor NOR3 (N2818, N2809, N207, N2556);
not NOT1 (N2819, N2815);
not NOT1 (N2820, N2789);
nor NOR2 (N2821, N2818, N563);
not NOT1 (N2822, N2816);
nor NOR4 (N2823, N2814, N2759, N2770, N2644);
xor XOR2 (N2824, N2819, N378);
xor XOR2 (N2825, N2812, N2626);
nor NOR4 (N2826, N2823, N2093, N591, N1081);
nor NOR3 (N2827, N2810, N2651, N1187);
not NOT1 (N2828, N2826);
and AND4 (N2829, N2821, N1829, N2617, N858);
nor NOR2 (N2830, N2822, N1977);
and AND2 (N2831, N2799, N312);
or OR4 (N2832, N2829, N300, N1450, N1059);
nor NOR2 (N2833, N2817, N357);
or OR4 (N2834, N2830, N2169, N425, N397);
xor XOR2 (N2835, N2827, N1496);
xor XOR2 (N2836, N2834, N1498);
buf BUF1 (N2837, N2825);
nand NAND3 (N2838, N2835, N550, N463);
not NOT1 (N2839, N2828);
xor XOR2 (N2840, N2820, N2791);
nand NAND2 (N2841, N2804, N2599);
not NOT1 (N2842, N2839);
nand NAND3 (N2843, N2840, N1117, N850);
nand NAND3 (N2844, N2841, N1685, N2063);
buf BUF1 (N2845, N2843);
buf BUF1 (N2846, N2824);
xor XOR2 (N2847, N2832, N1220);
or OR3 (N2848, N2847, N932, N184);
nor NOR2 (N2849, N2848, N2327);
xor XOR2 (N2850, N2837, N2085);
nand NAND3 (N2851, N2836, N267, N628);
not NOT1 (N2852, N2833);
nand NAND2 (N2853, N2844, N1446);
or OR2 (N2854, N2851, N221);
or OR3 (N2855, N2852, N2478, N1284);
buf BUF1 (N2856, N2849);
xor XOR2 (N2857, N2856, N727);
or OR2 (N2858, N2855, N1092);
and AND4 (N2859, N2846, N174, N1656, N2114);
buf BUF1 (N2860, N2838);
buf BUF1 (N2861, N2857);
or OR2 (N2862, N2845, N2518);
buf BUF1 (N2863, N2860);
nand NAND4 (N2864, N2863, N2353, N933, N2179);
nor NOR3 (N2865, N2858, N1810, N2542);
buf BUF1 (N2866, N2865);
nor NOR4 (N2867, N2866, N1630, N2038, N2342);
or OR3 (N2868, N2867, N2417, N1504);
and AND3 (N2869, N2853, N763, N2751);
or OR4 (N2870, N2864, N957, N1039, N1831);
and AND3 (N2871, N2870, N1817, N1972);
nand NAND4 (N2872, N2850, N454, N2513, N920);
buf BUF1 (N2873, N2842);
and AND3 (N2874, N2831, N1000, N1989);
nor NOR2 (N2875, N2862, N681);
xor XOR2 (N2876, N2872, N203);
not NOT1 (N2877, N2859);
xor XOR2 (N2878, N2871, N2766);
or OR4 (N2879, N2854, N2488, N2662, N1875);
not NOT1 (N2880, N2869);
and AND2 (N2881, N2876, N2382);
and AND3 (N2882, N2880, N1595, N2087);
and AND4 (N2883, N2861, N768, N674, N1169);
and AND2 (N2884, N2873, N1514);
or OR2 (N2885, N2877, N2507);
and AND3 (N2886, N2884, N1355, N1901);
buf BUF1 (N2887, N2879);
xor XOR2 (N2888, N2881, N2089);
or OR3 (N2889, N2882, N2032, N137);
xor XOR2 (N2890, N2886, N2820);
not NOT1 (N2891, N2890);
nor NOR3 (N2892, N2878, N833, N23);
not NOT1 (N2893, N2889);
or OR4 (N2894, N2883, N457, N1360, N655);
not NOT1 (N2895, N2887);
not NOT1 (N2896, N2892);
buf BUF1 (N2897, N2868);
not NOT1 (N2898, N2891);
or OR2 (N2899, N2893, N200);
or OR3 (N2900, N2874, N905, N952);
nor NOR2 (N2901, N2888, N1401);
and AND2 (N2902, N2896, N18);
nor NOR4 (N2903, N2897, N2475, N1675, N1679);
buf BUF1 (N2904, N2898);
nor NOR4 (N2905, N2902, N643, N73, N1561);
or OR4 (N2906, N2894, N2292, N2586, N2624);
or OR3 (N2907, N2906, N2210, N2807);
and AND4 (N2908, N2903, N827, N2314, N2906);
nor NOR2 (N2909, N2907, N2898);
and AND2 (N2910, N2904, N2485);
nor NOR4 (N2911, N2909, N1531, N1953, N1189);
buf BUF1 (N2912, N2901);
and AND4 (N2913, N2905, N2018, N657, N1565);
xor XOR2 (N2914, N2908, N2894);
xor XOR2 (N2915, N2914, N2331);
nor NOR3 (N2916, N2900, N2678, N1661);
or OR3 (N2917, N2915, N486, N695);
nand NAND2 (N2918, N2913, N2139);
not NOT1 (N2919, N2916);
xor XOR2 (N2920, N2918, N2605);
not NOT1 (N2921, N2885);
buf BUF1 (N2922, N2919);
or OR3 (N2923, N2910, N748, N2155);
nor NOR3 (N2924, N2895, N1003, N1031);
or OR4 (N2925, N2875, N2093, N1962, N2119);
or OR3 (N2926, N2925, N733, N1250);
buf BUF1 (N2927, N2911);
nor NOR2 (N2928, N2922, N183);
nor NOR3 (N2929, N2926, N653, N1522);
xor XOR2 (N2930, N2912, N1622);
not NOT1 (N2931, N2921);
nor NOR2 (N2932, N2929, N443);
not NOT1 (N2933, N2917);
nor NOR3 (N2934, N2924, N590, N1197);
xor XOR2 (N2935, N2932, N285);
xor XOR2 (N2936, N2927, N1636);
and AND2 (N2937, N2933, N1327);
xor XOR2 (N2938, N2923, N2781);
nand NAND3 (N2939, N2934, N2702, N1029);
or OR3 (N2940, N2931, N2283, N1773);
xor XOR2 (N2941, N2928, N2089);
and AND2 (N2942, N2899, N629);
xor XOR2 (N2943, N2941, N556);
nand NAND3 (N2944, N2942, N2463, N1389);
and AND3 (N2945, N2938, N1838, N1922);
or OR2 (N2946, N2939, N344);
xor XOR2 (N2947, N2920, N742);
or OR3 (N2948, N2944, N1722, N1361);
and AND2 (N2949, N2943, N844);
nor NOR4 (N2950, N2946, N2240, N2454, N2776);
not NOT1 (N2951, N2936);
or OR2 (N2952, N2930, N1344);
xor XOR2 (N2953, N2949, N2872);
and AND4 (N2954, N2940, N2170, N46, N2947);
nand NAND2 (N2955, N561, N2639);
not NOT1 (N2956, N2945);
or OR4 (N2957, N2951, N1096, N2109, N1819);
not NOT1 (N2958, N2948);
or OR2 (N2959, N2952, N1109);
nand NAND4 (N2960, N2955, N1857, N1480, N2377);
buf BUF1 (N2961, N2960);
or OR2 (N2962, N2957, N2085);
and AND4 (N2963, N2953, N1874, N2385, N348);
or OR4 (N2964, N2954, N2505, N1065, N678);
nand NAND4 (N2965, N2937, N887, N2525, N1273);
nor NOR3 (N2966, N2950, N267, N2002);
not NOT1 (N2967, N2964);
or OR3 (N2968, N2962, N157, N2475);
not NOT1 (N2969, N2961);
nand NAND3 (N2970, N2935, N895, N217);
not NOT1 (N2971, N2965);
or OR4 (N2972, N2958, N1351, N1117, N2671);
not NOT1 (N2973, N2972);
buf BUF1 (N2974, N2970);
xor XOR2 (N2975, N2967, N1090);
or OR2 (N2976, N2973, N289);
or OR2 (N2977, N2966, N1803);
xor XOR2 (N2978, N2974, N1322);
not NOT1 (N2979, N2975);
or OR4 (N2980, N2968, N727, N2539, N640);
or OR2 (N2981, N2980, N211);
nor NOR2 (N2982, N2971, N1535);
and AND3 (N2983, N2969, N2152, N1128);
and AND3 (N2984, N2978, N847, N2033);
nor NOR2 (N2985, N2979, N2509);
nand NAND2 (N2986, N2981, N591);
xor XOR2 (N2987, N2956, N1998);
not NOT1 (N2988, N2977);
and AND2 (N2989, N2988, N2596);
xor XOR2 (N2990, N2976, N1827);
nor NOR4 (N2991, N2987, N2429, N929, N1075);
nand NAND4 (N2992, N2983, N1003, N383, N799);
and AND3 (N2993, N2986, N1470, N2785);
or OR3 (N2994, N2982, N1940, N2852);
not NOT1 (N2995, N2993);
nor NOR4 (N2996, N2992, N512, N2817, N2894);
buf BUF1 (N2997, N2959);
nor NOR3 (N2998, N2997, N1290, N2396);
or OR3 (N2999, N2990, N2640, N2698);
nor NOR3 (N3000, N2999, N2598, N1881);
nor NOR4 (N3001, N2991, N464, N304, N2794);
xor XOR2 (N3002, N2985, N2612);
nor NOR4 (N3003, N2998, N780, N1047, N2447);
nand NAND4 (N3004, N3001, N1621, N2172, N32);
nand NAND2 (N3005, N2963, N1502);
xor XOR2 (N3006, N3002, N2330);
or OR4 (N3007, N2994, N555, N991, N2383);
xor XOR2 (N3008, N3003, N214);
nor NOR4 (N3009, N3007, N1464, N1053, N814);
and AND3 (N3010, N3008, N2021, N2491);
xor XOR2 (N3011, N3005, N266);
and AND2 (N3012, N2989, N665);
buf BUF1 (N3013, N3011);
nand NAND3 (N3014, N3004, N401, N2342);
or OR4 (N3015, N2984, N1346, N1713, N1857);
buf BUF1 (N3016, N3015);
not NOT1 (N3017, N3000);
and AND3 (N3018, N2995, N1182, N802);
nand NAND4 (N3019, N2996, N1175, N805, N2965);
nor NOR2 (N3020, N3019, N857);
or OR4 (N3021, N3020, N1169, N994, N839);
or OR2 (N3022, N3021, N1981);
nor NOR4 (N3023, N3016, N2597, N882, N2915);
nor NOR4 (N3024, N3013, N1061, N1272, N377);
buf BUF1 (N3025, N3017);
xor XOR2 (N3026, N3025, N1073);
nor NOR3 (N3027, N3010, N2453, N1256);
or OR4 (N3028, N3018, N771, N211, N1800);
xor XOR2 (N3029, N3012, N2602);
nor NOR4 (N3030, N3022, N2044, N2386, N1992);
and AND2 (N3031, N3009, N1465);
nor NOR4 (N3032, N3031, N825, N1885, N1469);
not NOT1 (N3033, N3027);
and AND2 (N3034, N3032, N357);
not NOT1 (N3035, N3033);
nor NOR3 (N3036, N3023, N2094, N167);
nor NOR2 (N3037, N3034, N757);
and AND3 (N3038, N3037, N1547, N2963);
nor NOR2 (N3039, N3006, N2533);
xor XOR2 (N3040, N3038, N2295);
nor NOR4 (N3041, N3040, N2538, N3024, N1034);
not NOT1 (N3042, N1330);
nand NAND2 (N3043, N3028, N2117);
not NOT1 (N3044, N3041);
buf BUF1 (N3045, N3014);
not NOT1 (N3046, N3029);
and AND2 (N3047, N3046, N2102);
or OR3 (N3048, N3047, N683, N2725);
and AND4 (N3049, N3030, N884, N2403, N836);
or OR3 (N3050, N3036, N2574, N318);
nand NAND2 (N3051, N3044, N2858);
buf BUF1 (N3052, N3051);
and AND4 (N3053, N3043, N2515, N2186, N1874);
not NOT1 (N3054, N3035);
or OR4 (N3055, N3052, N73, N2950, N266);
nor NOR2 (N3056, N3049, N944);
buf BUF1 (N3057, N3050);
or OR2 (N3058, N3045, N1804);
buf BUF1 (N3059, N3039);
buf BUF1 (N3060, N3054);
xor XOR2 (N3061, N3042, N2901);
xor XOR2 (N3062, N3026, N859);
nor NOR2 (N3063, N3055, N1128);
nor NOR2 (N3064, N3048, N123);
not NOT1 (N3065, N3060);
nor NOR3 (N3066, N3065, N2289, N1204);
or OR3 (N3067, N3064, N1264, N704);
buf BUF1 (N3068, N3066);
nor NOR4 (N3069, N3056, N2477, N1712, N985);
nand NAND4 (N3070, N3062, N2347, N2796, N1989);
and AND4 (N3071, N3069, N1212, N178, N880);
or OR3 (N3072, N3058, N404, N1794);
and AND4 (N3073, N3067, N1017, N2093, N902);
or OR3 (N3074, N3072, N2387, N1488);
and AND3 (N3075, N3063, N2515, N2630);
buf BUF1 (N3076, N3073);
buf BUF1 (N3077, N3070);
nor NOR3 (N3078, N3059, N1351, N1595);
nor NOR3 (N3079, N3061, N1071, N792);
xor XOR2 (N3080, N3079, N1721);
or OR4 (N3081, N3053, N2807, N1581, N317);
and AND2 (N3082, N3074, N497);
xor XOR2 (N3083, N3068, N2946);
not NOT1 (N3084, N3078);
xor XOR2 (N3085, N3071, N144);
and AND3 (N3086, N3081, N2820, N2111);
and AND2 (N3087, N3084, N1414);
buf BUF1 (N3088, N3080);
xor XOR2 (N3089, N3077, N36);
nand NAND4 (N3090, N3082, N2122, N1386, N331);
xor XOR2 (N3091, N3090, N99);
nor NOR2 (N3092, N3086, N2500);
or OR2 (N3093, N3076, N435);
xor XOR2 (N3094, N3057, N953);
buf BUF1 (N3095, N3092);
xor XOR2 (N3096, N3088, N1863);
or OR4 (N3097, N3089, N2182, N718, N917);
nor NOR4 (N3098, N3091, N1492, N878, N999);
or OR2 (N3099, N3096, N764);
not NOT1 (N3100, N3099);
and AND2 (N3101, N3085, N3011);
nand NAND4 (N3102, N3075, N2055, N2603, N12);
buf BUF1 (N3103, N3100);
xor XOR2 (N3104, N3098, N2034);
nand NAND4 (N3105, N3102, N2640, N2996, N2719);
or OR4 (N3106, N3103, N808, N1102, N1040);
and AND4 (N3107, N3093, N710, N1467, N1690);
or OR2 (N3108, N3106, N943);
not NOT1 (N3109, N3101);
buf BUF1 (N3110, N3083);
not NOT1 (N3111, N3107);
nand NAND2 (N3112, N3104, N34);
nor NOR2 (N3113, N3109, N577);
or OR3 (N3114, N3110, N2205, N3059);
or OR2 (N3115, N3114, N1989);
or OR2 (N3116, N3111, N645);
xor XOR2 (N3117, N3116, N1494);
and AND3 (N3118, N3117, N2801, N341);
and AND3 (N3119, N3094, N3117, N229);
or OR3 (N3120, N3105, N2671, N867);
buf BUF1 (N3121, N3119);
nor NOR2 (N3122, N3095, N2049);
xor XOR2 (N3123, N3113, N449);
xor XOR2 (N3124, N3122, N760);
buf BUF1 (N3125, N3087);
or OR4 (N3126, N3125, N473, N524, N131);
not NOT1 (N3127, N3112);
nand NAND3 (N3128, N3124, N794, N1949);
xor XOR2 (N3129, N3108, N1635);
not NOT1 (N3130, N3126);
xor XOR2 (N3131, N3129, N680);
buf BUF1 (N3132, N3127);
xor XOR2 (N3133, N3130, N440);
nor NOR3 (N3134, N3118, N843, N1059);
nor NOR4 (N3135, N3115, N2636, N2835, N2786);
buf BUF1 (N3136, N3123);
nor NOR2 (N3137, N3097, N224);
nand NAND4 (N3138, N3121, N2390, N1227, N2261);
buf BUF1 (N3139, N3132);
nand NAND4 (N3140, N3133, N1173, N1679, N2492);
not NOT1 (N3141, N3136);
nor NOR4 (N3142, N3137, N2607, N729, N2581);
nand NAND4 (N3143, N3138, N2656, N60, N142);
not NOT1 (N3144, N3135);
nor NOR2 (N3145, N3128, N286);
nand NAND2 (N3146, N3134, N2670);
not NOT1 (N3147, N3120);
nand NAND3 (N3148, N3146, N2710, N2678);
buf BUF1 (N3149, N3131);
nand NAND4 (N3150, N3142, N1966, N2534, N2201);
not NOT1 (N3151, N3148);
and AND2 (N3152, N3141, N2906);
not NOT1 (N3153, N3143);
nand NAND4 (N3154, N3153, N1587, N2660, N2552);
xor XOR2 (N3155, N3149, N223);
buf BUF1 (N3156, N3140);
nand NAND4 (N3157, N3147, N2333, N1329, N1986);
nor NOR4 (N3158, N3139, N1612, N2986, N1496);
or OR2 (N3159, N3145, N2850);
xor XOR2 (N3160, N3158, N2338);
nand NAND2 (N3161, N3160, N1804);
and AND3 (N3162, N3161, N631, N2543);
or OR4 (N3163, N3155, N2917, N1197, N2501);
xor XOR2 (N3164, N3154, N89);
nand NAND3 (N3165, N3156, N875, N2425);
or OR3 (N3166, N3163, N936, N2200);
nor NOR3 (N3167, N3165, N2818, N887);
and AND3 (N3168, N3151, N3155, N1327);
nor NOR4 (N3169, N3159, N779, N2125, N463);
and AND3 (N3170, N3144, N2137, N1706);
buf BUF1 (N3171, N3150);
or OR3 (N3172, N3170, N2076, N913);
and AND3 (N3173, N3164, N1261, N224);
nor NOR4 (N3174, N3173, N414, N2253, N16);
xor XOR2 (N3175, N3172, N515);
nor NOR2 (N3176, N3166, N2454);
or OR2 (N3177, N3157, N885);
nand NAND4 (N3178, N3176, N3083, N2713, N675);
buf BUF1 (N3179, N3167);
and AND4 (N3180, N3171, N1221, N478, N868);
or OR2 (N3181, N3177, N2489);
nand NAND4 (N3182, N3174, N1833, N2835, N747);
nor NOR3 (N3183, N3162, N477, N2362);
buf BUF1 (N3184, N3181);
and AND2 (N3185, N3179, N851);
nand NAND2 (N3186, N3183, N2270);
buf BUF1 (N3187, N3186);
and AND2 (N3188, N3187, N127);
and AND3 (N3189, N3188, N2827, N2784);
not NOT1 (N3190, N3180);
or OR3 (N3191, N3152, N1497, N2570);
buf BUF1 (N3192, N3182);
nor NOR2 (N3193, N3168, N1527);
nand NAND2 (N3194, N3169, N2899);
buf BUF1 (N3195, N3178);
and AND3 (N3196, N3190, N2562, N2645);
or OR2 (N3197, N3196, N2846);
nand NAND2 (N3198, N3194, N734);
xor XOR2 (N3199, N3191, N224);
or OR4 (N3200, N3199, N2650, N2092, N1041);
xor XOR2 (N3201, N3184, N1105);
nor NOR4 (N3202, N3195, N451, N68, N2586);
buf BUF1 (N3203, N3192);
and AND3 (N3204, N3202, N166, N2058);
nor NOR4 (N3205, N3200, N3195, N1, N1091);
and AND3 (N3206, N3197, N1131, N1795);
nand NAND3 (N3207, N3204, N3184, N1078);
or OR4 (N3208, N3198, N1132, N861, N2489);
nor NOR2 (N3209, N3193, N2677);
or OR4 (N3210, N3209, N1198, N1283, N3066);
and AND3 (N3211, N3207, N2174, N185);
xor XOR2 (N3212, N3210, N2262);
nand NAND2 (N3213, N3175, N1170);
and AND4 (N3214, N3189, N2588, N1293, N1130);
xor XOR2 (N3215, N3213, N2529);
buf BUF1 (N3216, N3208);
and AND2 (N3217, N3205, N681);
xor XOR2 (N3218, N3201, N566);
xor XOR2 (N3219, N3217, N900);
or OR3 (N3220, N3212, N1534, N2080);
nand NAND2 (N3221, N3214, N1668);
or OR2 (N3222, N3216, N2318);
nor NOR4 (N3223, N3203, N1308, N342, N470);
not NOT1 (N3224, N3220);
xor XOR2 (N3225, N3211, N2799);
nand NAND4 (N3226, N3185, N487, N1490, N1945);
nor NOR4 (N3227, N3222, N2428, N2325, N179);
xor XOR2 (N3228, N3221, N2483);
nand NAND4 (N3229, N3227, N1367, N937, N1348);
nand NAND4 (N3230, N3226, N1354, N2139, N2458);
not NOT1 (N3231, N3219);
not NOT1 (N3232, N3229);
not NOT1 (N3233, N3224);
buf BUF1 (N3234, N3218);
or OR3 (N3235, N3232, N2234, N86);
xor XOR2 (N3236, N3225, N1332);
nand NAND3 (N3237, N3206, N3118, N637);
xor XOR2 (N3238, N3234, N2721);
not NOT1 (N3239, N3223);
or OR2 (N3240, N3237, N2821);
or OR2 (N3241, N3238, N282);
and AND2 (N3242, N3239, N3148);
buf BUF1 (N3243, N3235);
or OR3 (N3244, N3236, N1525, N3237);
or OR2 (N3245, N3241, N1195);
not NOT1 (N3246, N3231);
xor XOR2 (N3247, N3243, N1321);
xor XOR2 (N3248, N3246, N487);
xor XOR2 (N3249, N3240, N2978);
or OR2 (N3250, N3249, N107);
not NOT1 (N3251, N3244);
xor XOR2 (N3252, N3247, N1413);
nand NAND4 (N3253, N3233, N1967, N2829, N448);
and AND3 (N3254, N3252, N1853, N1056);
or OR3 (N3255, N3230, N1724, N2887);
or OR2 (N3256, N3253, N1479);
nand NAND4 (N3257, N3248, N1542, N655, N1307);
nor NOR3 (N3258, N3215, N859, N2055);
nor NOR3 (N3259, N3255, N3205, N1696);
not NOT1 (N3260, N3242);
nand NAND2 (N3261, N3254, N2566);
or OR4 (N3262, N3245, N219, N1096, N991);
or OR3 (N3263, N3251, N2177, N3214);
or OR3 (N3264, N3262, N1363, N2508);
not NOT1 (N3265, N3250);
buf BUF1 (N3266, N3263);
buf BUF1 (N3267, N3261);
or OR3 (N3268, N3264, N927, N1192);
not NOT1 (N3269, N3258);
and AND2 (N3270, N3269, N2474);
xor XOR2 (N3271, N3270, N2360);
and AND3 (N3272, N3266, N1090, N2619);
buf BUF1 (N3273, N3228);
nand NAND2 (N3274, N3267, N3012);
buf BUF1 (N3275, N3265);
buf BUF1 (N3276, N3275);
and AND3 (N3277, N3274, N434, N352);
nand NAND4 (N3278, N3271, N107, N1522, N1108);
not NOT1 (N3279, N3277);
nand NAND4 (N3280, N3276, N1108, N2911, N2359);
nor NOR4 (N3281, N3273, N818, N2351, N713);
nand NAND4 (N3282, N3257, N954, N2431, N2427);
nor NOR2 (N3283, N3280, N840);
and AND3 (N3284, N3259, N1871, N1800);
not NOT1 (N3285, N3279);
xor XOR2 (N3286, N3256, N2835);
buf BUF1 (N3287, N3268);
or OR3 (N3288, N3278, N2247, N3159);
and AND3 (N3289, N3287, N1421, N1718);
nor NOR4 (N3290, N3282, N1296, N596, N1781);
buf BUF1 (N3291, N3289);
nor NOR3 (N3292, N3288, N2704, N2898);
or OR3 (N3293, N3281, N1005, N2275);
and AND4 (N3294, N3272, N1899, N32, N553);
nor NOR2 (N3295, N3283, N274);
and AND3 (N3296, N3292, N177, N2711);
xor XOR2 (N3297, N3290, N452);
not NOT1 (N3298, N3294);
nand NAND4 (N3299, N3286, N836, N2398, N439);
or OR3 (N3300, N3291, N2095, N53);
nor NOR3 (N3301, N3295, N1985, N463);
xor XOR2 (N3302, N3285, N1885);
buf BUF1 (N3303, N3296);
nand NAND2 (N3304, N3301, N2922);
buf BUF1 (N3305, N3284);
xor XOR2 (N3306, N3299, N1789);
or OR4 (N3307, N3304, N989, N436, N2044);
and AND3 (N3308, N3305, N855, N208);
xor XOR2 (N3309, N3260, N450);
nand NAND2 (N3310, N3293, N2752);
not NOT1 (N3311, N3297);
nand NAND4 (N3312, N3311, N968, N2315, N3201);
xor XOR2 (N3313, N3312, N474);
not NOT1 (N3314, N3313);
not NOT1 (N3315, N3306);
xor XOR2 (N3316, N3300, N2481);
xor XOR2 (N3317, N3316, N3179);
nand NAND3 (N3318, N3307, N270, N764);
xor XOR2 (N3319, N3318, N2874);
and AND3 (N3320, N3302, N2589, N1835);
and AND2 (N3321, N3320, N2851);
nor NOR3 (N3322, N3308, N1228, N638);
xor XOR2 (N3323, N3309, N1077);
or OR3 (N3324, N3298, N1232, N2326);
xor XOR2 (N3325, N3314, N1638);
and AND4 (N3326, N3322, N2901, N384, N1157);
xor XOR2 (N3327, N3321, N1321);
nor NOR4 (N3328, N3303, N2535, N506, N1856);
not NOT1 (N3329, N3315);
or OR2 (N3330, N3328, N128);
buf BUF1 (N3331, N3327);
xor XOR2 (N3332, N3329, N2454);
xor XOR2 (N3333, N3325, N2934);
and AND3 (N3334, N3331, N1593, N1101);
nand NAND3 (N3335, N3326, N2048, N1603);
xor XOR2 (N3336, N3310, N2665);
or OR3 (N3337, N3319, N2268, N2646);
not NOT1 (N3338, N3323);
xor XOR2 (N3339, N3335, N1363);
not NOT1 (N3340, N3334);
nor NOR3 (N3341, N3340, N2725, N1999);
and AND4 (N3342, N3332, N2385, N2547, N1502);
nand NAND2 (N3343, N3333, N2628);
nor NOR2 (N3344, N3342, N792);
or OR2 (N3345, N3344, N3334);
and AND4 (N3346, N3330, N2333, N2687, N608);
xor XOR2 (N3347, N3338, N3165);
buf BUF1 (N3348, N3347);
nor NOR4 (N3349, N3339, N959, N1201, N2347);
buf BUF1 (N3350, N3336);
nor NOR4 (N3351, N3345, N565, N3128, N1635);
and AND4 (N3352, N3324, N3029, N3155, N1159);
buf BUF1 (N3353, N3350);
or OR4 (N3354, N3352, N3023, N768, N2220);
or OR3 (N3355, N3346, N1126, N376);
xor XOR2 (N3356, N3348, N2268);
or OR4 (N3357, N3356, N1023, N2566, N3155);
buf BUF1 (N3358, N3341);
and AND4 (N3359, N3357, N869, N3018, N2530);
nor NOR4 (N3360, N3337, N3190, N3087, N2098);
nor NOR3 (N3361, N3360, N2561, N1620);
xor XOR2 (N3362, N3354, N1411);
buf BUF1 (N3363, N3355);
buf BUF1 (N3364, N3353);
buf BUF1 (N3365, N3358);
buf BUF1 (N3366, N3349);
and AND4 (N3367, N3365, N86, N1713, N3040);
not NOT1 (N3368, N3351);
not NOT1 (N3369, N3343);
or OR2 (N3370, N3367, N921);
and AND4 (N3371, N3363, N488, N571, N1745);
xor XOR2 (N3372, N3366, N2565);
not NOT1 (N3373, N3359);
or OR3 (N3374, N3317, N3063, N1547);
not NOT1 (N3375, N3374);
nor NOR3 (N3376, N3364, N2643, N3353);
nand NAND4 (N3377, N3372, N2210, N894, N1953);
nand NAND2 (N3378, N3368, N3245);
buf BUF1 (N3379, N3369);
nor NOR3 (N3380, N3370, N761, N1003);
xor XOR2 (N3381, N3380, N1767);
not NOT1 (N3382, N3379);
xor XOR2 (N3383, N3373, N1774);
buf BUF1 (N3384, N3378);
not NOT1 (N3385, N3382);
nand NAND2 (N3386, N3377, N1406);
not NOT1 (N3387, N3362);
and AND3 (N3388, N3371, N2446, N1763);
xor XOR2 (N3389, N3376, N2346);
not NOT1 (N3390, N3387);
nand NAND4 (N3391, N3389, N2293, N2546, N1586);
buf BUF1 (N3392, N3385);
nand NAND3 (N3393, N3388, N1488, N2491);
nor NOR3 (N3394, N3386, N2912, N2219);
nand NAND3 (N3395, N3394, N2895, N3013);
buf BUF1 (N3396, N3395);
xor XOR2 (N3397, N3390, N2951);
not NOT1 (N3398, N3381);
nor NOR3 (N3399, N3398, N621, N1630);
xor XOR2 (N3400, N3399, N2660);
xor XOR2 (N3401, N3397, N463);
or OR4 (N3402, N3384, N214, N1937, N1297);
and AND2 (N3403, N3361, N3381);
nor NOR2 (N3404, N3392, N2253);
not NOT1 (N3405, N3396);
and AND4 (N3406, N3404, N283, N58, N432);
or OR2 (N3407, N3403, N3001);
nor NOR3 (N3408, N3407, N746, N767);
buf BUF1 (N3409, N3400);
nor NOR3 (N3410, N3401, N851, N2474);
nor NOR3 (N3411, N3391, N2015, N1032);
and AND3 (N3412, N3383, N2505, N2882);
nor NOR2 (N3413, N3375, N1463);
not NOT1 (N3414, N3393);
not NOT1 (N3415, N3406);
and AND4 (N3416, N3405, N1103, N1381, N3350);
nor NOR3 (N3417, N3411, N1645, N667);
buf BUF1 (N3418, N3402);
and AND4 (N3419, N3409, N3026, N1426, N2512);
not NOT1 (N3420, N3412);
nand NAND3 (N3421, N3415, N1009, N1360);
not NOT1 (N3422, N3421);
and AND3 (N3423, N3413, N2440, N1194);
and AND3 (N3424, N3410, N1897, N2201);
or OR2 (N3425, N3423, N439);
nand NAND4 (N3426, N3419, N1148, N3258, N2398);
buf BUF1 (N3427, N3426);
buf BUF1 (N3428, N3414);
xor XOR2 (N3429, N3424, N3246);
nand NAND3 (N3430, N3416, N2574, N2431);
not NOT1 (N3431, N3418);
nand NAND3 (N3432, N3430, N1288, N1280);
nand NAND3 (N3433, N3432, N2160, N1274);
buf BUF1 (N3434, N3429);
xor XOR2 (N3435, N3434, N2873);
nand NAND3 (N3436, N3427, N1258, N625);
not NOT1 (N3437, N3425);
buf BUF1 (N3438, N3428);
not NOT1 (N3439, N3438);
nor NOR4 (N3440, N3439, N2677, N575, N2946);
nor NOR2 (N3441, N3431, N3118);
or OR2 (N3442, N3440, N1691);
nand NAND2 (N3443, N3417, N2488);
and AND2 (N3444, N3443, N779);
xor XOR2 (N3445, N3420, N1223);
xor XOR2 (N3446, N3445, N1454);
buf BUF1 (N3447, N3435);
and AND3 (N3448, N3436, N535, N2650);
and AND3 (N3449, N3444, N822, N411);
xor XOR2 (N3450, N3433, N1719);
nor NOR4 (N3451, N3408, N1597, N1542, N1549);
or OR3 (N3452, N3451, N3049, N353);
not NOT1 (N3453, N3437);
nor NOR3 (N3454, N3452, N1590, N889);
or OR4 (N3455, N3442, N2927, N3248, N1239);
and AND4 (N3456, N3448, N2299, N1229, N461);
buf BUF1 (N3457, N3454);
xor XOR2 (N3458, N3457, N2756);
not NOT1 (N3459, N3441);
buf BUF1 (N3460, N3446);
or OR3 (N3461, N3460, N1545, N735);
not NOT1 (N3462, N3459);
or OR4 (N3463, N3456, N3164, N256, N3022);
buf BUF1 (N3464, N3449);
and AND2 (N3465, N3461, N279);
not NOT1 (N3466, N3455);
nor NOR2 (N3467, N3462, N1851);
not NOT1 (N3468, N3463);
buf BUF1 (N3469, N3450);
not NOT1 (N3470, N3453);
and AND4 (N3471, N3464, N1566, N3167, N450);
not NOT1 (N3472, N3471);
xor XOR2 (N3473, N3466, N1258);
or OR2 (N3474, N3470, N2569);
xor XOR2 (N3475, N3468, N3057);
not NOT1 (N3476, N3469);
nor NOR2 (N3477, N3473, N1555);
nand NAND2 (N3478, N3465, N2140);
nor NOR2 (N3479, N3422, N667);
nor NOR4 (N3480, N3476, N3464, N2234, N2616);
nor NOR4 (N3481, N3467, N3392, N3334, N786);
nand NAND3 (N3482, N3477, N2985, N846);
and AND4 (N3483, N3481, N1382, N37, N297);
or OR3 (N3484, N3472, N3430, N860);
nor NOR3 (N3485, N3480, N193, N3220);
or OR3 (N3486, N3475, N1867, N3384);
buf BUF1 (N3487, N3447);
nand NAND4 (N3488, N3474, N2945, N2898, N2964);
xor XOR2 (N3489, N3485, N2587);
xor XOR2 (N3490, N3484, N1018);
xor XOR2 (N3491, N3487, N401);
buf BUF1 (N3492, N3479);
nor NOR3 (N3493, N3490, N1496, N3349);
not NOT1 (N3494, N3482);
nand NAND4 (N3495, N3458, N1246, N2681, N1712);
nor NOR2 (N3496, N3478, N3124);
nand NAND3 (N3497, N3495, N2911, N2003);
and AND2 (N3498, N3493, N2667);
or OR4 (N3499, N3483, N1629, N1964, N925);
and AND2 (N3500, N3489, N1463);
not NOT1 (N3501, N3494);
not NOT1 (N3502, N3501);
buf BUF1 (N3503, N3497);
buf BUF1 (N3504, N3503);
and AND3 (N3505, N3500, N3090, N642);
and AND3 (N3506, N3486, N3460, N2358);
not NOT1 (N3507, N3505);
xor XOR2 (N3508, N3488, N1109);
nand NAND2 (N3509, N3491, N1755);
buf BUF1 (N3510, N3492);
not NOT1 (N3511, N3496);
nor NOR4 (N3512, N3507, N162, N1361, N354);
nand NAND3 (N3513, N3512, N1356, N115);
and AND3 (N3514, N3509, N285, N595);
or OR2 (N3515, N3499, N1115);
or OR2 (N3516, N3508, N2813);
nand NAND4 (N3517, N3515, N3481, N1485, N1755);
or OR2 (N3518, N3516, N1398);
nand NAND2 (N3519, N3498, N3263);
nor NOR2 (N3520, N3502, N1062);
xor XOR2 (N3521, N3506, N1201);
or OR2 (N3522, N3518, N3078);
xor XOR2 (N3523, N3519, N2296);
nor NOR4 (N3524, N3510, N962, N1512, N1757);
or OR3 (N3525, N3522, N854, N2163);
or OR4 (N3526, N3525, N706, N2400, N244);
and AND3 (N3527, N3517, N2650, N1340);
and AND3 (N3528, N3526, N1288, N2310);
nor NOR4 (N3529, N3511, N1447, N2720, N3304);
nand NAND4 (N3530, N3514, N3219, N368, N2243);
nor NOR2 (N3531, N3529, N1836);
or OR2 (N3532, N3520, N2358);
and AND4 (N3533, N3531, N163, N1574, N517);
buf BUF1 (N3534, N3527);
or OR4 (N3535, N3528, N2663, N2083, N308);
nand NAND4 (N3536, N3521, N509, N1997, N335);
not NOT1 (N3537, N3504);
buf BUF1 (N3538, N3537);
and AND4 (N3539, N3523, N2708, N3037, N2136);
or OR3 (N3540, N3539, N3417, N3008);
buf BUF1 (N3541, N3530);
buf BUF1 (N3542, N3538);
nand NAND3 (N3543, N3524, N959, N1340);
nand NAND4 (N3544, N3513, N1195, N2536, N643);
nand NAND4 (N3545, N3534, N1514, N1868, N3136);
nand NAND3 (N3546, N3542, N288, N1728);
not NOT1 (N3547, N3536);
and AND3 (N3548, N3532, N165, N1727);
not NOT1 (N3549, N3541);
xor XOR2 (N3550, N3548, N1766);
or OR2 (N3551, N3549, N2227);
and AND4 (N3552, N3540, N884, N2450, N390);
nor NOR2 (N3553, N3535, N651);
xor XOR2 (N3554, N3550, N1350);
or OR3 (N3555, N3546, N3109, N678);
buf BUF1 (N3556, N3551);
and AND4 (N3557, N3544, N1409, N666, N3435);
buf BUF1 (N3558, N3547);
not NOT1 (N3559, N3543);
buf BUF1 (N3560, N3533);
and AND2 (N3561, N3555, N3122);
or OR2 (N3562, N3559, N861);
or OR2 (N3563, N3553, N1464);
not NOT1 (N3564, N3561);
nand NAND2 (N3565, N3563, N1260);
nor NOR3 (N3566, N3562, N805, N1746);
nor NOR4 (N3567, N3560, N2830, N2484, N1316);
xor XOR2 (N3568, N3567, N3123);
and AND4 (N3569, N3557, N770, N161, N2010);
nor NOR2 (N3570, N3566, N2647);
xor XOR2 (N3571, N3554, N1711);
nand NAND2 (N3572, N3545, N2074);
buf BUF1 (N3573, N3570);
not NOT1 (N3574, N3558);
nor NOR3 (N3575, N3565, N3431, N2631);
and AND3 (N3576, N3556, N3573, N2923);
or OR4 (N3577, N2863, N2056, N2708, N1651);
buf BUF1 (N3578, N3569);
xor XOR2 (N3579, N3578, N2363);
buf BUF1 (N3580, N3576);
nor NOR4 (N3581, N3572, N2518, N197, N1385);
xor XOR2 (N3582, N3568, N1585);
or OR3 (N3583, N3574, N302, N70);
or OR2 (N3584, N3579, N1027);
and AND3 (N3585, N3584, N1596, N2384);
or OR2 (N3586, N3582, N3138);
nand NAND2 (N3587, N3585, N2299);
not NOT1 (N3588, N3586);
nor NOR4 (N3589, N3580, N1277, N3216, N3421);
buf BUF1 (N3590, N3564);
or OR2 (N3591, N3590, N1142);
nor NOR4 (N3592, N3581, N1782, N714, N3422);
buf BUF1 (N3593, N3592);
buf BUF1 (N3594, N3552);
buf BUF1 (N3595, N3575);
buf BUF1 (N3596, N3587);
xor XOR2 (N3597, N3593, N655);
not NOT1 (N3598, N3588);
nor NOR4 (N3599, N3596, N551, N2019, N3113);
xor XOR2 (N3600, N3583, N194);
buf BUF1 (N3601, N3597);
and AND3 (N3602, N3600, N3442, N964);
not NOT1 (N3603, N3591);
nor NOR3 (N3604, N3598, N20, N382);
not NOT1 (N3605, N3603);
or OR3 (N3606, N3589, N1145, N1031);
nand NAND3 (N3607, N3602, N1175, N3296);
or OR4 (N3608, N3606, N622, N975, N1822);
not NOT1 (N3609, N3577);
buf BUF1 (N3610, N3595);
or OR3 (N3611, N3594, N170, N2610);
buf BUF1 (N3612, N3610);
not NOT1 (N3613, N3607);
xor XOR2 (N3614, N3601, N3277);
buf BUF1 (N3615, N3599);
nand NAND4 (N3616, N3611, N1865, N1497, N1852);
nand NAND3 (N3617, N3612, N1562, N1393);
nand NAND3 (N3618, N3617, N1066, N2358);
xor XOR2 (N3619, N3616, N946);
or OR2 (N3620, N3609, N3045);
or OR4 (N3621, N3618, N3126, N2011, N2595);
xor XOR2 (N3622, N3608, N17);
buf BUF1 (N3623, N3620);
buf BUF1 (N3624, N3614);
buf BUF1 (N3625, N3621);
not NOT1 (N3626, N3623);
nor NOR3 (N3627, N3613, N2325, N136);
or OR2 (N3628, N3627, N290);
buf BUF1 (N3629, N3622);
buf BUF1 (N3630, N3605);
buf BUF1 (N3631, N3628);
and AND4 (N3632, N3619, N1821, N3471, N3325);
not NOT1 (N3633, N3626);
not NOT1 (N3634, N3630);
nor NOR4 (N3635, N3631, N64, N1578, N711);
xor XOR2 (N3636, N3633, N3507);
not NOT1 (N3637, N3634);
nor NOR4 (N3638, N3604, N3241, N739, N2579);
xor XOR2 (N3639, N3638, N549);
nor NOR4 (N3640, N3629, N3334, N273, N1869);
nand NAND4 (N3641, N3637, N3218, N772, N573);
xor XOR2 (N3642, N3632, N2379);
nor NOR4 (N3643, N3615, N45, N967, N2658);
not NOT1 (N3644, N3636);
nor NOR4 (N3645, N3635, N858, N3122, N2484);
or OR4 (N3646, N3642, N143, N46, N171);
xor XOR2 (N3647, N3571, N765);
xor XOR2 (N3648, N3640, N2240);
nand NAND3 (N3649, N3645, N3259, N665);
nor NOR4 (N3650, N3644, N550, N3302, N3327);
nor NOR4 (N3651, N3649, N1319, N74, N3518);
not NOT1 (N3652, N3650);
not NOT1 (N3653, N3652);
nand NAND4 (N3654, N3639, N499, N1681, N3381);
not NOT1 (N3655, N3643);
not NOT1 (N3656, N3651);
xor XOR2 (N3657, N3656, N3379);
xor XOR2 (N3658, N3641, N560);
xor XOR2 (N3659, N3658, N1532);
nand NAND3 (N3660, N3655, N1188, N281);
not NOT1 (N3661, N3646);
nand NAND4 (N3662, N3624, N3106, N3126, N2034);
and AND4 (N3663, N3653, N3254, N784, N2775);
nor NOR4 (N3664, N3648, N3163, N1641, N1150);
xor XOR2 (N3665, N3654, N2453);
buf BUF1 (N3666, N3625);
xor XOR2 (N3667, N3662, N252);
nor NOR2 (N3668, N3660, N3483);
xor XOR2 (N3669, N3657, N2115);
xor XOR2 (N3670, N3667, N573);
nor NOR2 (N3671, N3664, N2094);
and AND2 (N3672, N3668, N1189);
nand NAND3 (N3673, N3672, N1371, N1783);
or OR4 (N3674, N3669, N2683, N1501, N3288);
nand NAND4 (N3675, N3659, N984, N1903, N3285);
nor NOR3 (N3676, N3673, N407, N302);
not NOT1 (N3677, N3663);
nand NAND2 (N3678, N3671, N2632);
or OR4 (N3679, N3647, N3001, N3433, N1470);
not NOT1 (N3680, N3666);
and AND3 (N3681, N3680, N2256, N687);
and AND4 (N3682, N3661, N1928, N2912, N434);
buf BUF1 (N3683, N3665);
or OR4 (N3684, N3678, N897, N3375, N1758);
not NOT1 (N3685, N3683);
or OR4 (N3686, N3677, N79, N1746, N279);
buf BUF1 (N3687, N3685);
and AND3 (N3688, N3686, N3029, N2649);
xor XOR2 (N3689, N3688, N3298);
and AND3 (N3690, N3675, N647, N1568);
xor XOR2 (N3691, N3679, N205);
xor XOR2 (N3692, N3674, N3497);
and AND2 (N3693, N3684, N2296);
nand NAND3 (N3694, N3676, N1931, N1738);
nand NAND4 (N3695, N3693, N942, N2669, N392);
buf BUF1 (N3696, N3689);
and AND3 (N3697, N3694, N3072, N52);
nor NOR4 (N3698, N3670, N2494, N1074, N3628);
buf BUF1 (N3699, N3690);
or OR3 (N3700, N3695, N460, N2641);
nand NAND2 (N3701, N3682, N2392);
buf BUF1 (N3702, N3692);
buf BUF1 (N3703, N3701);
xor XOR2 (N3704, N3698, N2212);
or OR4 (N3705, N3696, N2998, N3173, N1076);
not NOT1 (N3706, N3705);
nor NOR3 (N3707, N3687, N220, N566);
not NOT1 (N3708, N3703);
xor XOR2 (N3709, N3691, N3377);
nand NAND3 (N3710, N3704, N996, N1982);
nand NAND2 (N3711, N3708, N214);
nor NOR2 (N3712, N3707, N1124);
nand NAND3 (N3713, N3697, N996, N3033);
xor XOR2 (N3714, N3702, N3684);
buf BUF1 (N3715, N3709);
xor XOR2 (N3716, N3710, N681);
nand NAND4 (N3717, N3706, N1129, N2586, N1451);
xor XOR2 (N3718, N3714, N1682);
xor XOR2 (N3719, N3717, N1856);
nand NAND2 (N3720, N3711, N562);
nor NOR4 (N3721, N3715, N3385, N2377, N2644);
and AND4 (N3722, N3718, N1917, N2117, N2148);
and AND4 (N3723, N3699, N2544, N1816, N329);
or OR4 (N3724, N3721, N3582, N3496, N3578);
nand NAND3 (N3725, N3719, N3254, N1948);
and AND2 (N3726, N3713, N334);
xor XOR2 (N3727, N3716, N2374);
xor XOR2 (N3728, N3725, N3610);
not NOT1 (N3729, N3681);
buf BUF1 (N3730, N3722);
xor XOR2 (N3731, N3700, N1036);
xor XOR2 (N3732, N3726, N3171);
or OR2 (N3733, N3712, N2839);
buf BUF1 (N3734, N3720);
nand NAND3 (N3735, N3730, N169, N27);
buf BUF1 (N3736, N3732);
xor XOR2 (N3737, N3736, N540);
buf BUF1 (N3738, N3735);
buf BUF1 (N3739, N3727);
nand NAND4 (N3740, N3737, N2984, N3305, N3553);
and AND3 (N3741, N3723, N444, N2528);
or OR4 (N3742, N3724, N2569, N2965, N254);
not NOT1 (N3743, N3731);
nor NOR3 (N3744, N3740, N1531, N1002);
xor XOR2 (N3745, N3741, N1068);
xor XOR2 (N3746, N3745, N2615);
xor XOR2 (N3747, N3733, N2750);
nor NOR2 (N3748, N3747, N3246);
and AND2 (N3749, N3739, N69);
not NOT1 (N3750, N3734);
xor XOR2 (N3751, N3728, N2713);
nand NAND3 (N3752, N3749, N3133, N2119);
buf BUF1 (N3753, N3743);
or OR4 (N3754, N3750, N2942, N118, N3279);
buf BUF1 (N3755, N3742);
nor NOR3 (N3756, N3752, N4, N3276);
nor NOR3 (N3757, N3755, N2038, N1621);
or OR3 (N3758, N3729, N220, N2478);
buf BUF1 (N3759, N3751);
nor NOR3 (N3760, N3738, N2782, N1756);
buf BUF1 (N3761, N3756);
not NOT1 (N3762, N3757);
nand NAND3 (N3763, N3753, N1630, N3166);
not NOT1 (N3764, N3761);
or OR3 (N3765, N3759, N2995, N2032);
xor XOR2 (N3766, N3746, N1750);
nor NOR2 (N3767, N3765, N315);
or OR4 (N3768, N3748, N1587, N3415, N1367);
nor NOR4 (N3769, N3744, N466, N1558, N2358);
nor NOR4 (N3770, N3767, N213, N2561, N914);
or OR4 (N3771, N3768, N3006, N1905, N2212);
xor XOR2 (N3772, N3771, N2132);
nor NOR2 (N3773, N3763, N499);
or OR4 (N3774, N3758, N1099, N952, N1200);
and AND4 (N3775, N3766, N2147, N3039, N769);
nand NAND2 (N3776, N3773, N3585);
nor NOR4 (N3777, N3776, N3666, N976, N1363);
buf BUF1 (N3778, N3760);
and AND4 (N3779, N3777, N727, N2250, N2165);
nor NOR3 (N3780, N3775, N3490, N1398);
not NOT1 (N3781, N3770);
not NOT1 (N3782, N3772);
xor XOR2 (N3783, N3779, N3321);
or OR4 (N3784, N3781, N1456, N2028, N2174);
not NOT1 (N3785, N3784);
nand NAND2 (N3786, N3762, N2745);
and AND2 (N3787, N3769, N1034);
nor NOR3 (N3788, N3778, N1913, N555);
and AND4 (N3789, N3783, N3588, N2980, N3289);
nor NOR2 (N3790, N3788, N1709);
buf BUF1 (N3791, N3786);
nor NOR4 (N3792, N3791, N2684, N47, N3027);
buf BUF1 (N3793, N3785);
nand NAND3 (N3794, N3789, N1713, N3397);
buf BUF1 (N3795, N3794);
nor NOR3 (N3796, N3787, N2727, N1709);
nand NAND3 (N3797, N3782, N253, N3655);
or OR2 (N3798, N3793, N1473);
buf BUF1 (N3799, N3796);
nor NOR2 (N3800, N3774, N1620);
buf BUF1 (N3801, N3754);
xor XOR2 (N3802, N3792, N1484);
nor NOR3 (N3803, N3780, N1274, N2158);
not NOT1 (N3804, N3797);
nand NAND2 (N3805, N3799, N306);
nor NOR3 (N3806, N3800, N3632, N2576);
and AND2 (N3807, N3802, N2932);
nand NAND3 (N3808, N3806, N3178, N1104);
nor NOR2 (N3809, N3808, N2226);
nand NAND4 (N3810, N3805, N2631, N2623, N2130);
nand NAND3 (N3811, N3803, N3664, N2475);
nor NOR2 (N3812, N3790, N3615);
not NOT1 (N3813, N3764);
buf BUF1 (N3814, N3801);
xor XOR2 (N3815, N3814, N1940);
xor XOR2 (N3816, N3809, N2565);
xor XOR2 (N3817, N3812, N1990);
or OR3 (N3818, N3798, N302, N1795);
xor XOR2 (N3819, N3804, N1516);
nand NAND3 (N3820, N3810, N375, N1476);
buf BUF1 (N3821, N3813);
nand NAND3 (N3822, N3811, N1538, N980);
and AND2 (N3823, N3820, N1193);
nand NAND3 (N3824, N3819, N2966, N106);
and AND4 (N3825, N3823, N2896, N320, N3137);
xor XOR2 (N3826, N3815, N2126);
nor NOR2 (N3827, N3825, N2919);
or OR4 (N3828, N3795, N1736, N218, N1005);
buf BUF1 (N3829, N3817);
nor NOR3 (N3830, N3818, N148, N501);
not NOT1 (N3831, N3807);
or OR4 (N3832, N3829, N1423, N3658, N3693);
xor XOR2 (N3833, N3827, N3476);
nor NOR2 (N3834, N3830, N497);
buf BUF1 (N3835, N3828);
or OR4 (N3836, N3824, N2587, N784, N1859);
xor XOR2 (N3837, N3816, N849);
and AND4 (N3838, N3822, N446, N3023, N2736);
nand NAND2 (N3839, N3826, N2556);
nand NAND3 (N3840, N3821, N3023, N3438);
or OR4 (N3841, N3839, N437, N2717, N2530);
xor XOR2 (N3842, N3832, N437);
not NOT1 (N3843, N3837);
or OR4 (N3844, N3835, N672, N3115, N2653);
not NOT1 (N3845, N3836);
not NOT1 (N3846, N3831);
buf BUF1 (N3847, N3843);
and AND4 (N3848, N3845, N1660, N3319, N2009);
nand NAND3 (N3849, N3842, N223, N2689);
nand NAND3 (N3850, N3838, N160, N1660);
xor XOR2 (N3851, N3847, N3507);
nor NOR4 (N3852, N3850, N12, N1164, N2238);
xor XOR2 (N3853, N3841, N2641);
buf BUF1 (N3854, N3833);
and AND2 (N3855, N3852, N545);
nand NAND3 (N3856, N3840, N2986, N3636);
and AND4 (N3857, N3844, N664, N3247, N1059);
and AND2 (N3858, N3856, N1035);
buf BUF1 (N3859, N3846);
nand NAND4 (N3860, N3857, N576, N1821, N782);
nor NOR3 (N3861, N3858, N2173, N2327);
nand NAND4 (N3862, N3834, N3286, N2568, N2935);
buf BUF1 (N3863, N3851);
not NOT1 (N3864, N3848);
nor NOR3 (N3865, N3859, N1444, N2098);
or OR3 (N3866, N3853, N2625, N865);
or OR4 (N3867, N3866, N3733, N756, N22);
and AND2 (N3868, N3849, N1303);
nor NOR2 (N3869, N3865, N3709);
nand NAND3 (N3870, N3861, N3075, N304);
not NOT1 (N3871, N3862);
nand NAND4 (N3872, N3864, N529, N1009, N2023);
nor NOR4 (N3873, N3860, N3374, N2756, N2493);
buf BUF1 (N3874, N3863);
not NOT1 (N3875, N3872);
nand NAND4 (N3876, N3873, N420, N515, N481);
or OR3 (N3877, N3869, N1680, N755);
xor XOR2 (N3878, N3867, N64);
or OR4 (N3879, N3855, N285, N3660, N3203);
nor NOR3 (N3880, N3877, N462, N1280);
nand NAND2 (N3881, N3880, N3342);
buf BUF1 (N3882, N3854);
xor XOR2 (N3883, N3882, N2060);
xor XOR2 (N3884, N3875, N311);
not NOT1 (N3885, N3879);
nand NAND3 (N3886, N3870, N3517, N3221);
xor XOR2 (N3887, N3881, N3158);
or OR3 (N3888, N3886, N1278, N411);
nand NAND4 (N3889, N3887, N515, N725, N1061);
or OR3 (N3890, N3871, N3343, N3663);
or OR2 (N3891, N3883, N1499);
buf BUF1 (N3892, N3876);
xor XOR2 (N3893, N3888, N2113);
nor NOR4 (N3894, N3885, N3451, N1952, N1960);
nand NAND4 (N3895, N3894, N2556, N3185, N2643);
nand NAND2 (N3896, N3884, N3212);
or OR4 (N3897, N3895, N2842, N1021, N3197);
xor XOR2 (N3898, N3891, N1780);
not NOT1 (N3899, N3897);
nor NOR3 (N3900, N3868, N1011, N626);
not NOT1 (N3901, N3893);
buf BUF1 (N3902, N3874);
or OR2 (N3903, N3902, N844);
not NOT1 (N3904, N3899);
nor NOR4 (N3905, N3904, N2844, N64, N1025);
nor NOR3 (N3906, N3890, N2648, N1993);
nor NOR2 (N3907, N3896, N780);
or OR3 (N3908, N3889, N916, N3296);
nand NAND2 (N3909, N3898, N1606);
or OR2 (N3910, N3908, N3881);
and AND2 (N3911, N3909, N1397);
and AND2 (N3912, N3878, N1000);
and AND2 (N3913, N3911, N263);
nor NOR4 (N3914, N3912, N2501, N3237, N3460);
or OR3 (N3915, N3907, N3192, N3256);
and AND4 (N3916, N3914, N3376, N676, N728);
and AND2 (N3917, N3901, N315);
nand NAND4 (N3918, N3905, N2979, N1011, N42);
nor NOR2 (N3919, N3918, N1010);
nor NOR2 (N3920, N3900, N1567);
buf BUF1 (N3921, N3916);
buf BUF1 (N3922, N3906);
nor NOR3 (N3923, N3892, N3659, N3486);
nor NOR4 (N3924, N3923, N561, N2219, N2506);
nand NAND3 (N3925, N3917, N2642, N3285);
buf BUF1 (N3926, N3919);
nand NAND2 (N3927, N3913, N2019);
or OR3 (N3928, N3910, N3646, N116);
nor NOR4 (N3929, N3921, N859, N3418, N2578);
not NOT1 (N3930, N3927);
not NOT1 (N3931, N3925);
nor NOR2 (N3932, N3930, N502);
xor XOR2 (N3933, N3931, N1311);
not NOT1 (N3934, N3932);
xor XOR2 (N3935, N3903, N1340);
buf BUF1 (N3936, N3915);
not NOT1 (N3937, N3920);
nor NOR3 (N3938, N3926, N655, N2287);
and AND3 (N3939, N3922, N3413, N3457);
or OR3 (N3940, N3937, N505, N3194);
nor NOR4 (N3941, N3938, N1466, N3418, N199);
xor XOR2 (N3942, N3929, N3156);
and AND2 (N3943, N3940, N2874);
buf BUF1 (N3944, N3935);
nand NAND3 (N3945, N3934, N1226, N239);
nor NOR3 (N3946, N3933, N2973, N711);
not NOT1 (N3947, N3943);
not NOT1 (N3948, N3946);
not NOT1 (N3949, N3928);
and AND3 (N3950, N3924, N2974, N1967);
and AND4 (N3951, N3942, N2380, N2223, N2899);
xor XOR2 (N3952, N3949, N2225);
nand NAND4 (N3953, N3936, N3680, N2500, N1712);
buf BUF1 (N3954, N3948);
nand NAND2 (N3955, N3941, N54);
nor NOR4 (N3956, N3952, N1804, N3315, N711);
or OR4 (N3957, N3944, N862, N1008, N2420);
or OR3 (N3958, N3950, N2192, N2584);
nor NOR4 (N3959, N3954, N2682, N1380, N1743);
nor NOR4 (N3960, N3956, N381, N1189, N335);
nor NOR3 (N3961, N3959, N2760, N1895);
buf BUF1 (N3962, N3958);
and AND4 (N3963, N3961, N3383, N2169, N2052);
buf BUF1 (N3964, N3957);
or OR2 (N3965, N3945, N3123);
nor NOR2 (N3966, N3964, N2255);
buf BUF1 (N3967, N3962);
or OR2 (N3968, N3960, N1916);
nor NOR3 (N3969, N3967, N3830, N47);
nor NOR4 (N3970, N3966, N1329, N2567, N2223);
not NOT1 (N3971, N3970);
not NOT1 (N3972, N3939);
xor XOR2 (N3973, N3953, N1621);
and AND2 (N3974, N3965, N87);
nor NOR4 (N3975, N3973, N813, N782, N3522);
buf BUF1 (N3976, N3972);
nand NAND4 (N3977, N3968, N1947, N3236, N1530);
not NOT1 (N3978, N3951);
buf BUF1 (N3979, N3963);
or OR4 (N3980, N3955, N3197, N464, N2228);
nand NAND3 (N3981, N3975, N3660, N3612);
or OR3 (N3982, N3979, N3621, N1529);
nand NAND4 (N3983, N3971, N1339, N137, N758);
not NOT1 (N3984, N3947);
nand NAND2 (N3985, N3984, N862);
buf BUF1 (N3986, N3977);
and AND2 (N3987, N3982, N862);
and AND4 (N3988, N3981, N1102, N1670, N2927);
buf BUF1 (N3989, N3978);
nand NAND4 (N3990, N3976, N1505, N22, N3151);
nor NOR4 (N3991, N3989, N2365, N1005, N3052);
nor NOR2 (N3992, N3980, N1958);
nor NOR3 (N3993, N3992, N1444, N2497);
or OR3 (N3994, N3983, N592, N1046);
buf BUF1 (N3995, N3974);
nand NAND3 (N3996, N3994, N1807, N3611);
xor XOR2 (N3997, N3995, N2189);
or OR3 (N3998, N3988, N1711, N708);
and AND2 (N3999, N3985, N2501);
xor XOR2 (N4000, N3997, N2684);
not NOT1 (N4001, N3986);
not NOT1 (N4002, N3993);
nand NAND3 (N4003, N3999, N487, N2291);
xor XOR2 (N4004, N3990, N1239);
not NOT1 (N4005, N4002);
or OR2 (N4006, N3987, N2952);
or OR2 (N4007, N4003, N454);
not NOT1 (N4008, N3969);
or OR3 (N4009, N4007, N1690, N2561);
nand NAND2 (N4010, N3998, N1206);
nor NOR2 (N4011, N3996, N2623);
nand NAND4 (N4012, N4005, N1410, N210, N1575);
nand NAND2 (N4013, N4004, N2762);
and AND3 (N4014, N4010, N2117, N1270);
xor XOR2 (N4015, N4006, N451);
not NOT1 (N4016, N4001);
and AND4 (N4017, N4012, N729, N3264, N1752);
nand NAND4 (N4018, N4013, N2363, N3652, N2835);
and AND3 (N4019, N4000, N1611, N1618);
or OR4 (N4020, N4018, N1438, N3454, N3455);
nor NOR4 (N4021, N4009, N3990, N1137, N3089);
nor NOR4 (N4022, N4019, N3641, N3764, N595);
and AND4 (N4023, N4017, N517, N1554, N3643);
nor NOR3 (N4024, N4011, N1690, N860);
nand NAND3 (N4025, N4022, N803, N1028);
and AND4 (N4026, N4024, N2135, N1320, N2151);
xor XOR2 (N4027, N4016, N3707);
or OR4 (N4028, N4020, N100, N1858, N2203);
not NOT1 (N4029, N4027);
buf BUF1 (N4030, N4021);
xor XOR2 (N4031, N4008, N3097);
buf BUF1 (N4032, N4015);
nor NOR4 (N4033, N4029, N3342, N2795, N1427);
xor XOR2 (N4034, N4031, N1496);
nor NOR2 (N4035, N4028, N1117);
nand NAND3 (N4036, N4035, N387, N1708);
and AND3 (N4037, N4023, N2502, N3956);
xor XOR2 (N4038, N4014, N3928);
or OR4 (N4039, N4025, N1005, N905, N2266);
nand NAND4 (N4040, N4039, N3928, N1699, N240);
nand NAND2 (N4041, N4026, N2490);
xor XOR2 (N4042, N4030, N1452);
or OR3 (N4043, N4037, N262, N2015);
not NOT1 (N4044, N4032);
xor XOR2 (N4045, N3991, N2443);
nor NOR3 (N4046, N4045, N3764, N2674);
nand NAND4 (N4047, N4046, N2006, N693, N2004);
nand NAND3 (N4048, N4033, N813, N3508);
nand NAND4 (N4049, N4043, N836, N1468, N19);
xor XOR2 (N4050, N4049, N4020);
xor XOR2 (N4051, N4050, N1950);
xor XOR2 (N4052, N4051, N1156);
nand NAND4 (N4053, N4044, N3879, N3379, N234);
nor NOR3 (N4054, N4038, N653, N754);
not NOT1 (N4055, N4048);
nand NAND3 (N4056, N4052, N2154, N1036);
or OR2 (N4057, N4055, N1823);
buf BUF1 (N4058, N4041);
not NOT1 (N4059, N4042);
xor XOR2 (N4060, N4034, N1456);
xor XOR2 (N4061, N4058, N2520);
and AND2 (N4062, N4054, N145);
buf BUF1 (N4063, N4062);
nor NOR2 (N4064, N4047, N1654);
buf BUF1 (N4065, N4053);
buf BUF1 (N4066, N4056);
buf BUF1 (N4067, N4066);
and AND4 (N4068, N4040, N2294, N2474, N3887);
xor XOR2 (N4069, N4061, N1943);
not NOT1 (N4070, N4059);
xor XOR2 (N4071, N4069, N2746);
xor XOR2 (N4072, N4063, N1971);
or OR4 (N4073, N4060, N1049, N1681, N1331);
nor NOR4 (N4074, N4036, N3490, N708, N3629);
xor XOR2 (N4075, N4057, N2199);
and AND4 (N4076, N4075, N945, N2794, N3573);
not NOT1 (N4077, N4065);
buf BUF1 (N4078, N4064);
and AND4 (N4079, N4068, N1999, N2297, N681);
buf BUF1 (N4080, N4072);
or OR2 (N4081, N4071, N1646);
nand NAND3 (N4082, N4081, N431, N1960);
nor NOR4 (N4083, N4074, N825, N1976, N903);
and AND3 (N4084, N4082, N3600, N1203);
or OR3 (N4085, N4080, N3074, N1886);
xor XOR2 (N4086, N4070, N1624);
and AND3 (N4087, N4079, N829, N3832);
and AND2 (N4088, N4085, N158);
nor NOR3 (N4089, N4084, N1941, N180);
and AND3 (N4090, N4088, N326, N910);
nor NOR4 (N4091, N4089, N1418, N3394, N2130);
not NOT1 (N4092, N4083);
nand NAND3 (N4093, N4086, N253, N3450);
nand NAND3 (N4094, N4078, N1882, N3551);
xor XOR2 (N4095, N4077, N3559);
buf BUF1 (N4096, N4076);
or OR2 (N4097, N4073, N1087);
buf BUF1 (N4098, N4094);
buf BUF1 (N4099, N4097);
not NOT1 (N4100, N4096);
xor XOR2 (N4101, N4092, N3904);
and AND4 (N4102, N4095, N848, N3641, N3515);
buf BUF1 (N4103, N4101);
and AND4 (N4104, N4102, N1858, N1680, N2458);
xor XOR2 (N4105, N4091, N75);
and AND3 (N4106, N4104, N1170, N1274);
buf BUF1 (N4107, N4087);
nor NOR3 (N4108, N4098, N2943, N2517);
not NOT1 (N4109, N4105);
nor NOR4 (N4110, N4067, N865, N3771, N1644);
nand NAND3 (N4111, N4106, N1307, N1199);
or OR4 (N4112, N4100, N3577, N800, N1876);
and AND4 (N4113, N4107, N853, N2119, N3344);
nand NAND4 (N4114, N4112, N2678, N1635, N3291);
and AND3 (N4115, N4114, N1061, N1961);
xor XOR2 (N4116, N4113, N722);
not NOT1 (N4117, N4115);
nor NOR4 (N4118, N4108, N3641, N2242, N3135);
or OR4 (N4119, N4090, N1775, N2729, N2995);
not NOT1 (N4120, N4118);
not NOT1 (N4121, N4103);
or OR2 (N4122, N4119, N830);
and AND4 (N4123, N4111, N1610, N596, N1361);
not NOT1 (N4124, N4116);
buf BUF1 (N4125, N4120);
not NOT1 (N4126, N4117);
buf BUF1 (N4127, N4123);
or OR2 (N4128, N4110, N2161);
buf BUF1 (N4129, N4125);
nor NOR3 (N4130, N4124, N659, N154);
not NOT1 (N4131, N4093);
and AND4 (N4132, N4122, N3886, N2633, N2309);
nand NAND3 (N4133, N4121, N1862, N1646);
buf BUF1 (N4134, N4129);
not NOT1 (N4135, N4099);
nor NOR4 (N4136, N4133, N2214, N2469, N2474);
not NOT1 (N4137, N4135);
nand NAND3 (N4138, N4137, N3654, N3458);
xor XOR2 (N4139, N4109, N224);
and AND2 (N4140, N4138, N1006);
xor XOR2 (N4141, N4130, N2498);
and AND2 (N4142, N4134, N3283);
buf BUF1 (N4143, N4141);
buf BUF1 (N4144, N4136);
and AND4 (N4145, N4131, N2410, N4114, N3581);
and AND4 (N4146, N4142, N2757, N2915, N914);
or OR4 (N4147, N4132, N2025, N2576, N3001);
nand NAND3 (N4148, N4128, N1328, N2429);
buf BUF1 (N4149, N4144);
and AND3 (N4150, N4127, N293, N2177);
and AND4 (N4151, N4150, N724, N1180, N1211);
nor NOR3 (N4152, N4149, N913, N2228);
or OR3 (N4153, N4152, N3490, N245);
not NOT1 (N4154, N4139);
nor NOR3 (N4155, N4145, N1653, N1792);
xor XOR2 (N4156, N4155, N2058);
nand NAND4 (N4157, N4148, N1571, N1714, N4111);
xor XOR2 (N4158, N4143, N1060);
xor XOR2 (N4159, N4151, N2914);
nand NAND2 (N4160, N4159, N3923);
nor NOR2 (N4161, N4158, N166);
and AND3 (N4162, N4157, N1103, N3413);
and AND3 (N4163, N4146, N2261, N2337);
and AND3 (N4164, N4161, N283, N108);
and AND4 (N4165, N4156, N2162, N91, N1283);
and AND4 (N4166, N4163, N1713, N1856, N2710);
nor NOR3 (N4167, N4162, N517, N2413);
not NOT1 (N4168, N4160);
nand NAND4 (N4169, N4126, N3207, N3670, N1170);
and AND3 (N4170, N4168, N2020, N2184);
nand NAND2 (N4171, N4165, N536);
not NOT1 (N4172, N4167);
nor NOR3 (N4173, N4166, N2676, N3238);
nor NOR4 (N4174, N4147, N1246, N1527, N2552);
and AND2 (N4175, N4164, N738);
not NOT1 (N4176, N4170);
and AND2 (N4177, N4171, N501);
and AND4 (N4178, N4154, N4101, N3272, N786);
xor XOR2 (N4179, N4174, N330);
nor NOR4 (N4180, N4175, N4071, N3218, N1563);
nand NAND2 (N4181, N4177, N1587);
nand NAND3 (N4182, N4153, N291, N1676);
xor XOR2 (N4183, N4169, N1757);
nor NOR4 (N4184, N4179, N686, N2478, N1418);
and AND3 (N4185, N4140, N1356, N3942);
nand NAND2 (N4186, N4173, N1380);
not NOT1 (N4187, N4172);
buf BUF1 (N4188, N4187);
buf BUF1 (N4189, N4176);
not NOT1 (N4190, N4182);
and AND2 (N4191, N4184, N691);
xor XOR2 (N4192, N4186, N3215);
buf BUF1 (N4193, N4189);
xor XOR2 (N4194, N4183, N234);
buf BUF1 (N4195, N4192);
xor XOR2 (N4196, N4181, N546);
and AND3 (N4197, N4185, N72, N2733);
buf BUF1 (N4198, N4188);
xor XOR2 (N4199, N4197, N3230);
nor NOR3 (N4200, N4193, N305, N3188);
buf BUF1 (N4201, N4199);
nand NAND2 (N4202, N4196, N3595);
xor XOR2 (N4203, N4190, N1935);
nand NAND4 (N4204, N4202, N3600, N4152, N3155);
xor XOR2 (N4205, N4194, N1704);
and AND3 (N4206, N4195, N1268, N4181);
or OR3 (N4207, N4178, N227, N2041);
not NOT1 (N4208, N4200);
or OR4 (N4209, N4191, N1748, N490, N3883);
nand NAND2 (N4210, N4198, N1397);
not NOT1 (N4211, N4210);
nor NOR3 (N4212, N4201, N130, N3143);
buf BUF1 (N4213, N4211);
buf BUF1 (N4214, N4206);
buf BUF1 (N4215, N4213);
nor NOR3 (N4216, N4209, N4163, N705);
xor XOR2 (N4217, N4212, N2364);
nor NOR2 (N4218, N4180, N1716);
and AND4 (N4219, N4205, N1806, N1958, N4204);
buf BUF1 (N4220, N3273);
buf BUF1 (N4221, N4220);
not NOT1 (N4222, N4219);
or OR3 (N4223, N4216, N3646, N3072);
buf BUF1 (N4224, N4215);
buf BUF1 (N4225, N4207);
buf BUF1 (N4226, N4203);
nor NOR2 (N4227, N4208, N2585);
buf BUF1 (N4228, N4227);
nor NOR4 (N4229, N4221, N1757, N559, N2605);
nand NAND2 (N4230, N4226, N1900);
or OR3 (N4231, N4223, N3610, N1525);
nand NAND4 (N4232, N4228, N3722, N722, N472);
nand NAND3 (N4233, N4230, N235, N3597);
not NOT1 (N4234, N4233);
nor NOR2 (N4235, N4229, N3640);
nand NAND2 (N4236, N4222, N2431);
nor NOR3 (N4237, N4231, N821, N3670);
or OR3 (N4238, N4225, N661, N963);
nor NOR2 (N4239, N4234, N1708);
nand NAND4 (N4240, N4235, N2557, N366, N661);
xor XOR2 (N4241, N4237, N3950);
or OR4 (N4242, N4239, N657, N1615, N246);
and AND4 (N4243, N4238, N2975, N599, N2881);
xor XOR2 (N4244, N4224, N4154);
nand NAND2 (N4245, N4243, N3058);
nand NAND3 (N4246, N4236, N1825, N1434);
and AND4 (N4247, N4214, N3178, N3173, N3649);
nand NAND4 (N4248, N4246, N1044, N1106, N1028);
not NOT1 (N4249, N4248);
xor XOR2 (N4250, N4244, N3870);
xor XOR2 (N4251, N4241, N4178);
xor XOR2 (N4252, N4245, N162);
nand NAND2 (N4253, N4247, N4233);
not NOT1 (N4254, N4253);
or OR2 (N4255, N4254, N4224);
or OR2 (N4256, N4255, N3721);
nand NAND4 (N4257, N4218, N4155, N3065, N3441);
nand NAND4 (N4258, N4232, N1566, N3348, N1263);
or OR3 (N4259, N4242, N1957, N3442);
nand NAND3 (N4260, N4249, N3746, N1535);
buf BUF1 (N4261, N4240);
or OR3 (N4262, N4261, N1682, N1585);
and AND4 (N4263, N4262, N3359, N2050, N3398);
buf BUF1 (N4264, N4250);
xor XOR2 (N4265, N4264, N2810);
not NOT1 (N4266, N4258);
and AND2 (N4267, N4260, N752);
nor NOR2 (N4268, N4256, N2824);
nand NAND3 (N4269, N4259, N397, N2605);
and AND2 (N4270, N4257, N28);
xor XOR2 (N4271, N4267, N252);
nor NOR3 (N4272, N4268, N2838, N3486);
nor NOR4 (N4273, N4251, N173, N3110, N344);
and AND2 (N4274, N4263, N359);
xor XOR2 (N4275, N4271, N2347);
xor XOR2 (N4276, N4270, N4044);
or OR3 (N4277, N4252, N4169, N350);
or OR3 (N4278, N4269, N3709, N1068);
xor XOR2 (N4279, N4272, N349);
buf BUF1 (N4280, N4278);
not NOT1 (N4281, N4273);
not NOT1 (N4282, N4276);
xor XOR2 (N4283, N4280, N3918);
not NOT1 (N4284, N4265);
and AND2 (N4285, N4275, N508);
nand NAND2 (N4286, N4284, N3462);
xor XOR2 (N4287, N4286, N490);
and AND3 (N4288, N4266, N596, N2230);
buf BUF1 (N4289, N4282);
and AND4 (N4290, N4287, N808, N3943, N583);
nand NAND2 (N4291, N4289, N3487);
buf BUF1 (N4292, N4277);
not NOT1 (N4293, N4291);
buf BUF1 (N4294, N4279);
buf BUF1 (N4295, N4294);
buf BUF1 (N4296, N4217);
not NOT1 (N4297, N4290);
not NOT1 (N4298, N4281);
nand NAND4 (N4299, N4285, N2157, N1682, N3301);
and AND3 (N4300, N4283, N177, N1345);
xor XOR2 (N4301, N4299, N186);
nor NOR2 (N4302, N4292, N2516);
xor XOR2 (N4303, N4298, N3614);
nor NOR2 (N4304, N4296, N1361);
nor NOR4 (N4305, N4274, N1118, N2188, N3431);
xor XOR2 (N4306, N4297, N4103);
nor NOR2 (N4307, N4306, N2428);
and AND2 (N4308, N4300, N1301);
and AND4 (N4309, N4293, N4044, N901, N164);
not NOT1 (N4310, N4301);
or OR3 (N4311, N4304, N1769, N634);
nor NOR4 (N4312, N4303, N110, N3545, N1199);
nor NOR3 (N4313, N4307, N3721, N3578);
nor NOR2 (N4314, N4310, N154);
buf BUF1 (N4315, N4295);
not NOT1 (N4316, N4314);
xor XOR2 (N4317, N4309, N2853);
buf BUF1 (N4318, N4317);
not NOT1 (N4319, N4302);
nor NOR4 (N4320, N4305, N2010, N1921, N460);
xor XOR2 (N4321, N4318, N3507);
not NOT1 (N4322, N4320);
not NOT1 (N4323, N4321);
and AND4 (N4324, N4313, N2084, N3907, N1994);
nand NAND2 (N4325, N4319, N1286);
nand NAND2 (N4326, N4324, N223);
xor XOR2 (N4327, N4323, N2115);
nor NOR2 (N4328, N4312, N2744);
and AND2 (N4329, N4311, N410);
and AND3 (N4330, N4308, N4038, N3749);
buf BUF1 (N4331, N4329);
xor XOR2 (N4332, N4322, N3880);
buf BUF1 (N4333, N4332);
not NOT1 (N4334, N4315);
or OR3 (N4335, N4328, N3812, N4026);
and AND3 (N4336, N4335, N1667, N682);
or OR2 (N4337, N4330, N12);
and AND2 (N4338, N4327, N2763);
not NOT1 (N4339, N4336);
xor XOR2 (N4340, N4339, N2587);
and AND4 (N4341, N4340, N1039, N892, N3393);
not NOT1 (N4342, N4326);
nand NAND4 (N4343, N4331, N2428, N1836, N4036);
or OR3 (N4344, N4343, N3711, N1707);
xor XOR2 (N4345, N4333, N2018);
xor XOR2 (N4346, N4325, N2805);
not NOT1 (N4347, N4337);
nand NAND2 (N4348, N4341, N296);
nand NAND4 (N4349, N4338, N2356, N2971, N2654);
not NOT1 (N4350, N4316);
and AND3 (N4351, N4344, N4210, N2442);
buf BUF1 (N4352, N4350);
nand NAND3 (N4353, N4342, N2503, N2114);
xor XOR2 (N4354, N4352, N601);
xor XOR2 (N4355, N4349, N3232);
or OR4 (N4356, N4348, N3237, N1199, N3531);
xor XOR2 (N4357, N4347, N3076);
nand NAND2 (N4358, N4351, N4257);
nor NOR3 (N4359, N4353, N4070, N3008);
and AND2 (N4360, N4356, N1856);
not NOT1 (N4361, N4345);
not NOT1 (N4362, N4288);
and AND4 (N4363, N4346, N116, N3711, N248);
or OR4 (N4364, N4362, N1892, N4118, N548);
not NOT1 (N4365, N4358);
or OR4 (N4366, N4359, N415, N3217, N874);
and AND4 (N4367, N4366, N4077, N3394, N3292);
nor NOR4 (N4368, N4361, N1530, N2206, N3128);
buf BUF1 (N4369, N4360);
and AND3 (N4370, N4357, N3606, N2280);
buf BUF1 (N4371, N4365);
xor XOR2 (N4372, N4364, N406);
xor XOR2 (N4373, N4334, N3167);
xor XOR2 (N4374, N4372, N1705);
nand NAND3 (N4375, N4370, N2213, N3909);
xor XOR2 (N4376, N4368, N1279);
or OR3 (N4377, N4355, N2959, N2656);
buf BUF1 (N4378, N4377);
nor NOR3 (N4379, N4354, N3530, N3468);
nor NOR2 (N4380, N4371, N3865);
nor NOR2 (N4381, N4369, N2521);
nand NAND4 (N4382, N4376, N4074, N4253, N1551);
nor NOR3 (N4383, N4380, N550, N3968);
xor XOR2 (N4384, N4382, N2851);
nor NOR2 (N4385, N4383, N1667);
nand NAND2 (N4386, N4367, N2740);
or OR3 (N4387, N4378, N904, N2479);
and AND2 (N4388, N4387, N115);
or OR4 (N4389, N4375, N3809, N96, N2056);
nand NAND4 (N4390, N4374, N3547, N4359, N1167);
nor NOR2 (N4391, N4385, N4106);
and AND4 (N4392, N4390, N4193, N8, N321);
nand NAND3 (N4393, N4389, N4332, N3746);
nand NAND2 (N4394, N4363, N772);
nor NOR3 (N4395, N4393, N3875, N1029);
nor NOR2 (N4396, N4392, N335);
nor NOR3 (N4397, N4386, N1379, N2344);
nor NOR3 (N4398, N4391, N3810, N2379);
nor NOR3 (N4399, N4381, N2599, N4209);
nor NOR4 (N4400, N4395, N4131, N708, N4208);
nor NOR2 (N4401, N4384, N2752);
nor NOR3 (N4402, N4394, N970, N3259);
not NOT1 (N4403, N4396);
and AND4 (N4404, N4403, N1761, N4030, N4358);
and AND3 (N4405, N4398, N1976, N3426);
not NOT1 (N4406, N4402);
nand NAND4 (N4407, N4397, N3419, N1637, N4016);
and AND3 (N4408, N4404, N3344, N3810);
or OR2 (N4409, N4400, N4309);
nand NAND3 (N4410, N4408, N2062, N1507);
nand NAND3 (N4411, N4409, N1840, N3841);
or OR3 (N4412, N4373, N4028, N2432);
buf BUF1 (N4413, N4407);
xor XOR2 (N4414, N4410, N314);
buf BUF1 (N4415, N4405);
nand NAND4 (N4416, N4412, N4274, N1203, N3182);
buf BUF1 (N4417, N4413);
or OR4 (N4418, N4379, N1564, N1810, N3148);
xor XOR2 (N4419, N4415, N3619);
or OR4 (N4420, N4401, N4261, N2411, N2535);
buf BUF1 (N4421, N4388);
nor NOR4 (N4422, N4414, N2975, N520, N4017);
nand NAND3 (N4423, N4411, N1419, N3237);
xor XOR2 (N4424, N4419, N3123);
nor NOR3 (N4425, N4423, N2915, N2091);
not NOT1 (N4426, N4421);
nor NOR3 (N4427, N4422, N607, N2982);
and AND2 (N4428, N4418, N3791);
not NOT1 (N4429, N4399);
nor NOR3 (N4430, N4420, N1004, N2392);
nor NOR2 (N4431, N4425, N4168);
or OR2 (N4432, N4429, N2161);
buf BUF1 (N4433, N4430);
buf BUF1 (N4434, N4427);
xor XOR2 (N4435, N4434, N1497);
and AND2 (N4436, N4428, N1022);
nor NOR4 (N4437, N4435, N258, N3572, N1048);
nor NOR3 (N4438, N4406, N2460, N3864);
not NOT1 (N4439, N4437);
nor NOR2 (N4440, N4424, N2993);
and AND2 (N4441, N4417, N1512);
not NOT1 (N4442, N4436);
buf BUF1 (N4443, N4426);
not NOT1 (N4444, N4440);
and AND2 (N4445, N4442, N3349);
or OR4 (N4446, N4439, N1234, N1219, N2182);
xor XOR2 (N4447, N4446, N519);
nor NOR2 (N4448, N4441, N250);
and AND3 (N4449, N4445, N393, N3261);
and AND4 (N4450, N4433, N3253, N242, N3754);
buf BUF1 (N4451, N4450);
xor XOR2 (N4452, N4416, N693);
not NOT1 (N4453, N4444);
xor XOR2 (N4454, N4448, N4181);
not NOT1 (N4455, N4431);
nor NOR4 (N4456, N4447, N2475, N1472, N2940);
not NOT1 (N4457, N4449);
xor XOR2 (N4458, N4432, N478);
nand NAND4 (N4459, N4455, N2672, N2555, N3069);
not NOT1 (N4460, N4443);
nor NOR2 (N4461, N4459, N900);
xor XOR2 (N4462, N4438, N817);
not NOT1 (N4463, N4451);
and AND2 (N4464, N4453, N3758);
not NOT1 (N4465, N4457);
nand NAND2 (N4466, N4461, N1388);
xor XOR2 (N4467, N4460, N766);
nand NAND3 (N4468, N4454, N83, N1569);
nor NOR4 (N4469, N4456, N3378, N800, N2764);
xor XOR2 (N4470, N4462, N1951);
not NOT1 (N4471, N4467);
buf BUF1 (N4472, N4470);
nand NAND4 (N4473, N4466, N2757, N395, N2740);
buf BUF1 (N4474, N4471);
nor NOR3 (N4475, N4464, N818, N4469);
not NOT1 (N4476, N2568);
xor XOR2 (N4477, N4468, N1854);
not NOT1 (N4478, N4475);
nor NOR3 (N4479, N4476, N3148, N231);
not NOT1 (N4480, N4458);
not NOT1 (N4481, N4480);
not NOT1 (N4482, N4481);
and AND4 (N4483, N4482, N3769, N1031, N2318);
and AND3 (N4484, N4479, N3980, N2385);
buf BUF1 (N4485, N4473);
not NOT1 (N4486, N4477);
or OR3 (N4487, N4463, N4294, N3765);
buf BUF1 (N4488, N4486);
or OR4 (N4489, N4484, N3289, N7, N33);
buf BUF1 (N4490, N4474);
or OR3 (N4491, N4488, N3841, N3189);
or OR4 (N4492, N4487, N891, N1462, N193);
or OR4 (N4493, N4452, N2342, N2842, N1499);
or OR2 (N4494, N4485, N3523);
xor XOR2 (N4495, N4490, N3407);
xor XOR2 (N4496, N4493, N771);
nand NAND3 (N4497, N4495, N4361, N3058);
and AND4 (N4498, N4494, N2685, N753, N906);
and AND4 (N4499, N4492, N4106, N1603, N4330);
nand NAND2 (N4500, N4496, N3634);
not NOT1 (N4501, N4491);
xor XOR2 (N4502, N4489, N1331);
not NOT1 (N4503, N4478);
nand NAND4 (N4504, N4498, N1141, N2397, N2927);
not NOT1 (N4505, N4502);
or OR3 (N4506, N4504, N1026, N1174);
nand NAND2 (N4507, N4503, N1703);
or OR4 (N4508, N4472, N110, N5, N1299);
xor XOR2 (N4509, N4506, N1846);
nor NOR2 (N4510, N4505, N3951);
nand NAND2 (N4511, N4509, N128);
and AND4 (N4512, N4507, N2807, N405, N2312);
not NOT1 (N4513, N4500);
nand NAND2 (N4514, N4497, N245);
nand NAND3 (N4515, N4511, N2679, N2385);
or OR4 (N4516, N4499, N1544, N791, N4373);
nand NAND2 (N4517, N4465, N4478);
not NOT1 (N4518, N4483);
and AND3 (N4519, N4517, N3952, N80);
xor XOR2 (N4520, N4514, N2475);
not NOT1 (N4521, N4515);
nor NOR3 (N4522, N4510, N723, N269);
buf BUF1 (N4523, N4508);
or OR3 (N4524, N4521, N104, N718);
buf BUF1 (N4525, N4501);
or OR2 (N4526, N4524, N2911);
and AND4 (N4527, N4518, N1178, N2273, N1145);
xor XOR2 (N4528, N4520, N3828);
nand NAND4 (N4529, N4512, N2491, N3565, N803);
nand NAND3 (N4530, N4526, N1689, N3991);
nor NOR2 (N4531, N4528, N923);
nand NAND2 (N4532, N4530, N288);
or OR3 (N4533, N4525, N2963, N515);
or OR2 (N4534, N4516, N1182);
not NOT1 (N4535, N4522);
xor XOR2 (N4536, N4533, N2025);
and AND2 (N4537, N4519, N3872);
xor XOR2 (N4538, N4531, N3961);
xor XOR2 (N4539, N4534, N1127);
and AND3 (N4540, N4537, N1453, N3014);
nand NAND2 (N4541, N4527, N2458);
buf BUF1 (N4542, N4536);
not NOT1 (N4543, N4541);
not NOT1 (N4544, N4532);
buf BUF1 (N4545, N4535);
and AND3 (N4546, N4540, N3463, N4297);
and AND3 (N4547, N4542, N622, N1478);
and AND2 (N4548, N4513, N3361);
nand NAND4 (N4549, N4548, N317, N2113, N2272);
and AND3 (N4550, N4546, N790, N2069);
nor NOR4 (N4551, N4539, N3765, N3806, N628);
nor NOR4 (N4552, N4551, N2815, N3989, N2291);
buf BUF1 (N4553, N4529);
and AND3 (N4554, N4544, N3130, N2072);
or OR3 (N4555, N4554, N3148, N2398);
and AND2 (N4556, N4538, N3435);
buf BUF1 (N4557, N4549);
not NOT1 (N4558, N4557);
nor NOR4 (N4559, N4552, N78, N2097, N219);
nand NAND3 (N4560, N4558, N4169, N4212);
not NOT1 (N4561, N4556);
buf BUF1 (N4562, N4547);
not NOT1 (N4563, N4555);
buf BUF1 (N4564, N4563);
nor NOR3 (N4565, N4543, N1300, N545);
nor NOR3 (N4566, N4550, N4073, N4489);
not NOT1 (N4567, N4559);
and AND3 (N4568, N4562, N3116, N3434);
nand NAND3 (N4569, N4553, N826, N91);
xor XOR2 (N4570, N4564, N145);
and AND4 (N4571, N4560, N140, N3014, N2147);
nand NAND2 (N4572, N4565, N4089);
not NOT1 (N4573, N4571);
xor XOR2 (N4574, N4570, N1796);
xor XOR2 (N4575, N4561, N1415);
buf BUF1 (N4576, N4573);
xor XOR2 (N4577, N4576, N2894);
buf BUF1 (N4578, N4572);
not NOT1 (N4579, N4578);
not NOT1 (N4580, N4567);
or OR2 (N4581, N4566, N4226);
not NOT1 (N4582, N4545);
or OR2 (N4583, N4581, N2965);
buf BUF1 (N4584, N4579);
buf BUF1 (N4585, N4582);
or OR4 (N4586, N4585, N809, N1689, N1212);
nand NAND2 (N4587, N4586, N3839);
and AND2 (N4588, N4569, N4552);
nand NAND4 (N4589, N4588, N2336, N4401, N2854);
and AND2 (N4590, N4574, N1828);
nand NAND2 (N4591, N4587, N2286);
not NOT1 (N4592, N4523);
nor NOR4 (N4593, N4590, N890, N3602, N2648);
nor NOR3 (N4594, N4568, N1889, N2302);
buf BUF1 (N4595, N4591);
or OR3 (N4596, N4593, N2454, N822);
buf BUF1 (N4597, N4592);
not NOT1 (N4598, N4580);
buf BUF1 (N4599, N4583);
nand NAND3 (N4600, N4594, N1235, N1892);
and AND2 (N4601, N4597, N3703);
nor NOR4 (N4602, N4584, N2343, N323, N2147);
xor XOR2 (N4603, N4595, N841);
not NOT1 (N4604, N4603);
buf BUF1 (N4605, N4575);
nor NOR4 (N4606, N4604, N1600, N3099, N1138);
and AND4 (N4607, N4600, N2179, N3137, N2484);
buf BUF1 (N4608, N4577);
nand NAND2 (N4609, N4601, N1664);
buf BUF1 (N4610, N4605);
and AND4 (N4611, N4607, N813, N4589, N504);
nor NOR4 (N4612, N1296, N992, N4126, N1691);
nor NOR4 (N4613, N4612, N716, N2800, N2760);
nand NAND2 (N4614, N4610, N3280);
xor XOR2 (N4615, N4614, N3624);
nor NOR2 (N4616, N4611, N1568);
nand NAND4 (N4617, N4596, N2498, N2303, N1965);
and AND2 (N4618, N4598, N4183);
nor NOR2 (N4619, N4613, N180);
nor NOR3 (N4620, N4617, N382, N97);
or OR2 (N4621, N4619, N3158);
or OR4 (N4622, N4618, N3566, N4226, N2990);
nor NOR4 (N4623, N4620, N3977, N266, N2916);
or OR2 (N4624, N4616, N4287);
or OR2 (N4625, N4624, N182);
xor XOR2 (N4626, N4621, N2051);
not NOT1 (N4627, N4622);
buf BUF1 (N4628, N4608);
nand NAND3 (N4629, N4609, N4434, N2324);
xor XOR2 (N4630, N4602, N4438);
or OR2 (N4631, N4625, N2061);
not NOT1 (N4632, N4630);
nand NAND2 (N4633, N4599, N4333);
or OR4 (N4634, N4633, N312, N2764, N1592);
and AND3 (N4635, N4631, N309, N4498);
nand NAND3 (N4636, N4615, N360, N4125);
and AND4 (N4637, N4632, N2132, N4351, N2047);
or OR4 (N4638, N4635, N1000, N3756, N832);
and AND4 (N4639, N4629, N3087, N3614, N256);
nor NOR4 (N4640, N4637, N3774, N2187, N1240);
buf BUF1 (N4641, N4640);
xor XOR2 (N4642, N4628, N4085);
or OR3 (N4643, N4606, N2871, N96);
nand NAND3 (N4644, N4638, N2158, N325);
buf BUF1 (N4645, N4644);
not NOT1 (N4646, N4626);
not NOT1 (N4647, N4623);
not NOT1 (N4648, N4634);
buf BUF1 (N4649, N4639);
nand NAND4 (N4650, N4648, N1586, N3196, N3445);
or OR4 (N4651, N4646, N175, N3013, N1304);
buf BUF1 (N4652, N4636);
and AND4 (N4653, N4641, N3659, N1590, N851);
or OR3 (N4654, N4627, N843, N1551);
or OR2 (N4655, N4643, N3006);
or OR2 (N4656, N4650, N1660);
nor NOR3 (N4657, N4653, N663, N2403);
not NOT1 (N4658, N4647);
and AND4 (N4659, N4657, N2851, N4001, N1585);
and AND4 (N4660, N4651, N2675, N37, N3195);
not NOT1 (N4661, N4655);
xor XOR2 (N4662, N4660, N1141);
xor XOR2 (N4663, N4654, N1733);
nand NAND2 (N4664, N4663, N1054);
nand NAND4 (N4665, N4659, N3193, N2965, N3683);
nand NAND3 (N4666, N4658, N3772, N3658);
and AND3 (N4667, N4649, N1334, N4124);
not NOT1 (N4668, N4656);
nand NAND3 (N4669, N4645, N3177, N1171);
not NOT1 (N4670, N4664);
buf BUF1 (N4671, N4669);
xor XOR2 (N4672, N4668, N2826);
nand NAND4 (N4673, N4665, N3089, N3315, N3569);
nand NAND2 (N4674, N4642, N1034);
or OR2 (N4675, N4652, N855);
not NOT1 (N4676, N4666);
or OR4 (N4677, N4662, N3767, N1058, N999);
not NOT1 (N4678, N4675);
not NOT1 (N4679, N4673);
or OR3 (N4680, N4676, N1572, N4596);
nor NOR4 (N4681, N4672, N1868, N3316, N4680);
buf BUF1 (N4682, N979);
and AND4 (N4683, N4661, N2538, N4303, N1340);
not NOT1 (N4684, N4667);
buf BUF1 (N4685, N4670);
xor XOR2 (N4686, N4671, N2547);
buf BUF1 (N4687, N4685);
or OR3 (N4688, N4679, N2193, N3292);
and AND2 (N4689, N4687, N768);
buf BUF1 (N4690, N4689);
nand NAND2 (N4691, N4686, N1499);
nand NAND4 (N4692, N4683, N887, N192, N4252);
and AND2 (N4693, N4681, N1061);
not NOT1 (N4694, N4674);
nand NAND3 (N4695, N4688, N3462, N2994);
nand NAND3 (N4696, N4691, N3038, N3109);
buf BUF1 (N4697, N4695);
not NOT1 (N4698, N4682);
buf BUF1 (N4699, N4692);
not NOT1 (N4700, N4684);
or OR2 (N4701, N4699, N4631);
xor XOR2 (N4702, N4701, N3880);
nor NOR3 (N4703, N4693, N4347, N306);
and AND3 (N4704, N4677, N3789, N449);
nand NAND3 (N4705, N4697, N3684, N3833);
buf BUF1 (N4706, N4698);
not NOT1 (N4707, N4703);
not NOT1 (N4708, N4706);
buf BUF1 (N4709, N4696);
or OR4 (N4710, N4702, N4514, N3821, N4088);
buf BUF1 (N4711, N4705);
nor NOR3 (N4712, N4694, N4322, N1847);
not NOT1 (N4713, N4709);
xor XOR2 (N4714, N4712, N4190);
and AND3 (N4715, N4711, N1877, N1742);
and AND2 (N4716, N4690, N274);
nor NOR4 (N4717, N4714, N2090, N3009, N1164);
not NOT1 (N4718, N4715);
or OR4 (N4719, N4713, N562, N4141, N1002);
xor XOR2 (N4720, N4710, N4490);
nor NOR2 (N4721, N4700, N3791);
xor XOR2 (N4722, N4707, N1322);
nor NOR2 (N4723, N4720, N1736);
nor NOR4 (N4724, N4678, N1203, N2107, N3358);
or OR4 (N4725, N4722, N2168, N4649, N853);
or OR2 (N4726, N4716, N1977);
xor XOR2 (N4727, N4723, N1189);
not NOT1 (N4728, N4721);
or OR2 (N4729, N4717, N437);
and AND3 (N4730, N4724, N3169, N3784);
not NOT1 (N4731, N4718);
not NOT1 (N4732, N4719);
nand NAND4 (N4733, N4726, N709, N4119, N1173);
xor XOR2 (N4734, N4704, N1454);
xor XOR2 (N4735, N4734, N2747);
xor XOR2 (N4736, N4733, N4699);
and AND4 (N4737, N4727, N1133, N4069, N1973);
and AND4 (N4738, N4730, N1153, N3015, N1681);
xor XOR2 (N4739, N4728, N1026);
nand NAND3 (N4740, N4708, N3962, N3223);
or OR2 (N4741, N4739, N50);
and AND2 (N4742, N4731, N744);
xor XOR2 (N4743, N4741, N3769);
not NOT1 (N4744, N4729);
and AND4 (N4745, N4743, N3896, N4031, N4318);
nor NOR3 (N4746, N4745, N694, N1915);
nor NOR4 (N4747, N4742, N4259, N3863, N3151);
nand NAND2 (N4748, N4747, N2255);
not NOT1 (N4749, N4748);
not NOT1 (N4750, N4740);
xor XOR2 (N4751, N4750, N624);
or OR4 (N4752, N4744, N4557, N2390, N3817);
not NOT1 (N4753, N4738);
xor XOR2 (N4754, N4735, N69);
and AND3 (N4755, N4753, N2523, N4683);
and AND4 (N4756, N4754, N843, N2153, N3460);
xor XOR2 (N4757, N4755, N1569);
nor NOR3 (N4758, N4749, N228, N965);
buf BUF1 (N4759, N4736);
buf BUF1 (N4760, N4758);
buf BUF1 (N4761, N4751);
xor XOR2 (N4762, N4761, N270);
nor NOR3 (N4763, N4737, N2680, N1561);
nor NOR3 (N4764, N4762, N3056, N3518);
buf BUF1 (N4765, N4760);
xor XOR2 (N4766, N4764, N971);
not NOT1 (N4767, N4759);
nor NOR4 (N4768, N4765, N2676, N3108, N3466);
xor XOR2 (N4769, N4767, N2842);
or OR3 (N4770, N4746, N3818, N2002);
buf BUF1 (N4771, N4766);
nor NOR3 (N4772, N4770, N653, N1749);
nor NOR4 (N4773, N4772, N563, N3359, N4617);
or OR2 (N4774, N4757, N2979);
nand NAND2 (N4775, N4752, N4181);
nor NOR4 (N4776, N4725, N1462, N1647, N720);
nor NOR4 (N4777, N4775, N147, N2670, N293);
or OR4 (N4778, N4771, N17, N3726, N2999);
and AND4 (N4779, N4763, N1611, N2399, N3375);
buf BUF1 (N4780, N4769);
nor NOR3 (N4781, N4776, N2733, N4548);
and AND3 (N4782, N4778, N3515, N4773);
and AND2 (N4783, N1973, N3764);
buf BUF1 (N4784, N4777);
nor NOR4 (N4785, N4781, N2219, N2298, N2745);
nand NAND4 (N4786, N4783, N2719, N4152, N787);
or OR4 (N4787, N4780, N174, N3191, N4332);
buf BUF1 (N4788, N4782);
and AND4 (N4789, N4756, N3343, N3760, N4299);
buf BUF1 (N4790, N4785);
nand NAND3 (N4791, N4784, N650, N2539);
xor XOR2 (N4792, N4774, N4137);
or OR2 (N4793, N4779, N500);
and AND3 (N4794, N4768, N3744, N1782);
or OR3 (N4795, N4732, N2394, N1484);
not NOT1 (N4796, N4789);
nand NAND4 (N4797, N4793, N1403, N1767, N3592);
nor NOR2 (N4798, N4791, N663);
not NOT1 (N4799, N4788);
not NOT1 (N4800, N4794);
not NOT1 (N4801, N4797);
nor NOR4 (N4802, N4787, N3763, N1537, N2234);
xor XOR2 (N4803, N4792, N1779);
nand NAND3 (N4804, N4800, N3118, N1514);
or OR3 (N4805, N4795, N573, N2726);
xor XOR2 (N4806, N4805, N4285);
and AND4 (N4807, N4801, N682, N3896, N957);
buf BUF1 (N4808, N4804);
nor NOR4 (N4809, N4796, N2697, N4253, N4421);
not NOT1 (N4810, N4790);
buf BUF1 (N4811, N4806);
nor NOR2 (N4812, N4786, N4380);
buf BUF1 (N4813, N4810);
or OR4 (N4814, N4813, N3161, N4687, N1746);
or OR2 (N4815, N4798, N2577);
xor XOR2 (N4816, N4815, N3526);
xor XOR2 (N4817, N4814, N1128);
nand NAND3 (N4818, N4811, N495, N3435);
and AND4 (N4819, N4818, N1978, N1487, N4208);
not NOT1 (N4820, N4816);
not NOT1 (N4821, N4808);
buf BUF1 (N4822, N4809);
not NOT1 (N4823, N4812);
not NOT1 (N4824, N4821);
xor XOR2 (N4825, N4820, N1784);
or OR2 (N4826, N4807, N854);
or OR4 (N4827, N4826, N2999, N386, N4274);
nor NOR3 (N4828, N4824, N3504, N3783);
buf BUF1 (N4829, N4828);
and AND2 (N4830, N4817, N3945);
and AND2 (N4831, N4819, N3916);
nor NOR3 (N4832, N4822, N4001, N775);
and AND2 (N4833, N4823, N1709);
nor NOR3 (N4834, N4799, N773, N3016);
not NOT1 (N4835, N4831);
nor NOR3 (N4836, N4825, N1905, N1239);
buf BUF1 (N4837, N4803);
not NOT1 (N4838, N4830);
nor NOR4 (N4839, N4833, N1042, N4726, N4602);
not NOT1 (N4840, N4839);
xor XOR2 (N4841, N4829, N289);
nor NOR4 (N4842, N4827, N3628, N2465, N1279);
nand NAND2 (N4843, N4836, N4394);
xor XOR2 (N4844, N4841, N1667);
or OR4 (N4845, N4844, N3595, N2420, N2501);
xor XOR2 (N4846, N4832, N4263);
nor NOR4 (N4847, N4840, N1592, N4772, N3660);
xor XOR2 (N4848, N4847, N4433);
not NOT1 (N4849, N4835);
xor XOR2 (N4850, N4843, N606);
not NOT1 (N4851, N4842);
buf BUF1 (N4852, N4851);
nand NAND4 (N4853, N4849, N1107, N1669, N4257);
and AND3 (N4854, N4850, N4089, N3822);
buf BUF1 (N4855, N4802);
nor NOR2 (N4856, N4838, N1552);
xor XOR2 (N4857, N4852, N2071);
and AND4 (N4858, N4848, N2170, N45, N159);
nand NAND4 (N4859, N4853, N417, N2999, N1250);
xor XOR2 (N4860, N4837, N4855);
nand NAND4 (N4861, N4754, N2058, N3271, N555);
or OR2 (N4862, N4858, N1439);
buf BUF1 (N4863, N4857);
and AND4 (N4864, N4860, N3578, N4376, N652);
nor NOR2 (N4865, N4859, N909);
or OR4 (N4866, N4862, N397, N2238, N3321);
nand NAND3 (N4867, N4863, N142, N4862);
buf BUF1 (N4868, N4864);
or OR2 (N4869, N4867, N1165);
and AND3 (N4870, N4866, N272, N1043);
buf BUF1 (N4871, N4856);
and AND2 (N4872, N4846, N4580);
not NOT1 (N4873, N4871);
nor NOR2 (N4874, N4870, N1286);
not NOT1 (N4875, N4873);
or OR2 (N4876, N4872, N1821);
xor XOR2 (N4877, N4845, N3009);
xor XOR2 (N4878, N4875, N3126);
nor NOR2 (N4879, N4854, N1108);
buf BUF1 (N4880, N4869);
nor NOR2 (N4881, N4880, N2284);
xor XOR2 (N4882, N4879, N229);
and AND4 (N4883, N4878, N1128, N2969, N1289);
not NOT1 (N4884, N4882);
nor NOR2 (N4885, N4834, N2521);
or OR4 (N4886, N4876, N3577, N3687, N552);
nand NAND3 (N4887, N4877, N4379, N629);
not NOT1 (N4888, N4886);
not NOT1 (N4889, N4888);
nand NAND3 (N4890, N4874, N1217, N1983);
xor XOR2 (N4891, N4883, N749);
xor XOR2 (N4892, N4861, N2599);
xor XOR2 (N4893, N4865, N857);
nor NOR3 (N4894, N4891, N1698, N3799);
xor XOR2 (N4895, N4893, N1443);
xor XOR2 (N4896, N4885, N719);
not NOT1 (N4897, N4889);
not NOT1 (N4898, N4890);
and AND3 (N4899, N4896, N2709, N1338);
and AND3 (N4900, N4894, N3224, N3886);
not NOT1 (N4901, N4900);
or OR3 (N4902, N4901, N4662, N3263);
and AND2 (N4903, N4895, N1398);
buf BUF1 (N4904, N4892);
nand NAND4 (N4905, N4884, N276, N1616, N2232);
xor XOR2 (N4906, N4868, N1657);
nor NOR4 (N4907, N4899, N984, N1339, N2995);
nor NOR3 (N4908, N4897, N354, N2138);
nor NOR2 (N4909, N4902, N3852);
nand NAND2 (N4910, N4906, N2289);
nor NOR4 (N4911, N4887, N1221, N2943, N4152);
not NOT1 (N4912, N4907);
xor XOR2 (N4913, N4909, N1616);
xor XOR2 (N4914, N4908, N3174);
buf BUF1 (N4915, N4905);
nand NAND3 (N4916, N4912, N1493, N3877);
xor XOR2 (N4917, N4915, N2018);
nand NAND3 (N4918, N4914, N4428, N795);
nor NOR4 (N4919, N4881, N55, N2875, N2575);
not NOT1 (N4920, N4918);
and AND4 (N4921, N4910, N2850, N4316, N2511);
nor NOR2 (N4922, N4903, N4277);
not NOT1 (N4923, N4913);
and AND2 (N4924, N4920, N1236);
nand NAND2 (N4925, N4922, N3429);
not NOT1 (N4926, N4921);
buf BUF1 (N4927, N4926);
or OR3 (N4928, N4898, N4085, N4837);
nor NOR3 (N4929, N4911, N1328, N2616);
xor XOR2 (N4930, N4929, N2703);
and AND2 (N4931, N4917, N1818);
and AND2 (N4932, N4924, N3381);
nand NAND3 (N4933, N4930, N450, N4791);
nand NAND3 (N4934, N4925, N2293, N2518);
or OR4 (N4935, N4904, N430, N3692, N3419);
buf BUF1 (N4936, N4923);
and AND2 (N4937, N4927, N3315);
xor XOR2 (N4938, N4919, N4574);
nor NOR2 (N4939, N4933, N3780);
or OR4 (N4940, N4934, N107, N1879, N1325);
and AND3 (N4941, N4916, N4026, N3839);
xor XOR2 (N4942, N4937, N4221);
nand NAND3 (N4943, N4932, N959, N4222);
and AND3 (N4944, N4939, N3983, N4226);
xor XOR2 (N4945, N4928, N1345);
and AND4 (N4946, N4943, N2062, N3082, N3541);
buf BUF1 (N4947, N4935);
nand NAND3 (N4948, N4945, N4846, N1416);
nor NOR4 (N4949, N4940, N2761, N3473, N4606);
nand NAND2 (N4950, N4949, N3424);
nand NAND4 (N4951, N4948, N164, N3039, N1112);
buf BUF1 (N4952, N4936);
nor NOR3 (N4953, N4946, N2126, N1057);
or OR2 (N4954, N4938, N3552);
or OR3 (N4955, N4941, N2855, N984);
not NOT1 (N4956, N4952);
or OR2 (N4957, N4955, N394);
nor NOR2 (N4958, N4956, N3580);
and AND4 (N4959, N4953, N3459, N3439, N2804);
nand NAND4 (N4960, N4959, N1843, N3959, N1212);
not NOT1 (N4961, N4957);
buf BUF1 (N4962, N4947);
not NOT1 (N4963, N4961);
xor XOR2 (N4964, N4960, N923);
nand NAND4 (N4965, N4942, N3881, N4057, N3140);
nand NAND2 (N4966, N4931, N1734);
nand NAND4 (N4967, N4964, N2408, N3479, N431);
buf BUF1 (N4968, N4967);
buf BUF1 (N4969, N4962);
xor XOR2 (N4970, N4944, N3607);
buf BUF1 (N4971, N4969);
buf BUF1 (N4972, N4951);
and AND3 (N4973, N4971, N1941, N690);
not NOT1 (N4974, N4970);
or OR4 (N4975, N4968, N4136, N3849, N3572);
nor NOR2 (N4976, N4973, N4455);
nor NOR3 (N4977, N4958, N38, N1329);
nor NOR4 (N4978, N4976, N4921, N1411, N664);
or OR3 (N4979, N4966, N2859, N1422);
xor XOR2 (N4980, N4975, N1485);
and AND3 (N4981, N4974, N1467, N1741);
nor NOR2 (N4982, N4950, N2853);
nor NOR3 (N4983, N4979, N4084, N4474);
xor XOR2 (N4984, N4977, N4348);
or OR3 (N4985, N4982, N3627, N1148);
or OR3 (N4986, N4980, N2605, N4088);
nand NAND3 (N4987, N4972, N1679, N3748);
and AND3 (N4988, N4985, N2413, N2784);
xor XOR2 (N4989, N4965, N397);
not NOT1 (N4990, N4963);
and AND3 (N4991, N4983, N2981, N551);
not NOT1 (N4992, N4978);
xor XOR2 (N4993, N4986, N953);
xor XOR2 (N4994, N4992, N2906);
xor XOR2 (N4995, N4984, N755);
nand NAND3 (N4996, N4994, N1931, N3205);
not NOT1 (N4997, N4981);
nand NAND3 (N4998, N4988, N1432, N308);
and AND3 (N4999, N4987, N3783, N3175);
xor XOR2 (N5000, N4995, N4673);
nor NOR3 (N5001, N4998, N678, N1824);
not NOT1 (N5002, N4993);
not NOT1 (N5003, N5001);
xor XOR2 (N5004, N4996, N2523);
or OR3 (N5005, N5003, N3026, N1165);
or OR2 (N5006, N5004, N267);
or OR3 (N5007, N4999, N3946, N1578);
buf BUF1 (N5008, N4997);
not NOT1 (N5009, N5008);
not NOT1 (N5010, N5000);
and AND4 (N5011, N5009, N1375, N4493, N4975);
or OR3 (N5012, N5005, N425, N3179);
nand NAND3 (N5013, N5006, N2526, N3349);
buf BUF1 (N5014, N5002);
or OR4 (N5015, N5012, N743, N3363, N3773);
or OR3 (N5016, N5010, N2318, N638);
buf BUF1 (N5017, N5015);
xor XOR2 (N5018, N5017, N3698);
nor NOR3 (N5019, N5018, N1636, N4547);
or OR3 (N5020, N4954, N370, N4824);
and AND2 (N5021, N4989, N4726);
or OR4 (N5022, N5011, N4711, N4165, N4903);
and AND2 (N5023, N5016, N3271);
and AND3 (N5024, N5020, N947, N3988);
xor XOR2 (N5025, N5021, N1664);
not NOT1 (N5026, N4990);
nor NOR4 (N5027, N5023, N2038, N482, N2892);
xor XOR2 (N5028, N5013, N3278);
xor XOR2 (N5029, N5026, N1282);
nand NAND2 (N5030, N5029, N4100);
not NOT1 (N5031, N5024);
nand NAND2 (N5032, N5027, N4823);
nand NAND2 (N5033, N5032, N512);
nand NAND3 (N5034, N5025, N4040, N1624);
nor NOR3 (N5035, N4991, N1288, N4983);
not NOT1 (N5036, N5014);
or OR3 (N5037, N5019, N4394, N2632);
not NOT1 (N5038, N5028);
buf BUF1 (N5039, N5022);
or OR4 (N5040, N5033, N2972, N701, N3560);
xor XOR2 (N5041, N5007, N4700);
not NOT1 (N5042, N5034);
buf BUF1 (N5043, N5042);
xor XOR2 (N5044, N5039, N4475);
and AND2 (N5045, N5038, N3594);
xor XOR2 (N5046, N5041, N2590);
buf BUF1 (N5047, N5046);
nor NOR3 (N5048, N5045, N3214, N3046);
not NOT1 (N5049, N5031);
buf BUF1 (N5050, N5049);
or OR4 (N5051, N5047, N2314, N2602, N1128);
and AND3 (N5052, N5044, N2934, N2595);
nand NAND2 (N5053, N5048, N867);
buf BUF1 (N5054, N5050);
and AND2 (N5055, N5035, N3951);
xor XOR2 (N5056, N5036, N1860);
nor NOR4 (N5057, N5043, N1218, N4347, N605);
nor NOR3 (N5058, N5057, N2467, N2874);
nand NAND2 (N5059, N5037, N2249);
not NOT1 (N5060, N5059);
buf BUF1 (N5061, N5060);
or OR2 (N5062, N5056, N3354);
buf BUF1 (N5063, N5062);
and AND4 (N5064, N5055, N375, N2133, N1229);
buf BUF1 (N5065, N5051);
and AND2 (N5066, N5065, N135);
buf BUF1 (N5067, N5063);
nor NOR3 (N5068, N5052, N3971, N4427);
xor XOR2 (N5069, N5061, N1460);
nand NAND2 (N5070, N5054, N2127);
or OR2 (N5071, N5058, N4246);
buf BUF1 (N5072, N5064);
nor NOR2 (N5073, N5030, N330);
or OR3 (N5074, N5066, N3116, N4406);
not NOT1 (N5075, N5071);
nor NOR2 (N5076, N5067, N4270);
xor XOR2 (N5077, N5074, N19);
xor XOR2 (N5078, N5077, N1076);
and AND4 (N5079, N5040, N484, N1197, N3029);
not NOT1 (N5080, N5070);
and AND3 (N5081, N5076, N1045, N4758);
not NOT1 (N5082, N5072);
buf BUF1 (N5083, N5053);
nor NOR4 (N5084, N5081, N4362, N1004, N1453);
or OR4 (N5085, N5078, N4298, N3926, N2226);
buf BUF1 (N5086, N5068);
nor NOR2 (N5087, N5075, N2899);
buf BUF1 (N5088, N5086);
nor NOR2 (N5089, N5082, N4618);
xor XOR2 (N5090, N5069, N859);
xor XOR2 (N5091, N5090, N1786);
buf BUF1 (N5092, N5089);
buf BUF1 (N5093, N5084);
xor XOR2 (N5094, N5083, N754);
buf BUF1 (N5095, N5087);
not NOT1 (N5096, N5094);
nand NAND2 (N5097, N5093, N4717);
nand NAND4 (N5098, N5085, N3579, N672, N4319);
not NOT1 (N5099, N5091);
not NOT1 (N5100, N5096);
not NOT1 (N5101, N5088);
not NOT1 (N5102, N5097);
xor XOR2 (N5103, N5079, N1148);
nand NAND4 (N5104, N5073, N3782, N330, N2545);
and AND3 (N5105, N5099, N2011, N3832);
xor XOR2 (N5106, N5101, N1327);
buf BUF1 (N5107, N5102);
buf BUF1 (N5108, N5105);
or OR4 (N5109, N5100, N5013, N3965, N2889);
nor NOR4 (N5110, N5104, N3340, N5034, N2891);
buf BUF1 (N5111, N5110);
or OR4 (N5112, N5111, N2051, N3765, N2170);
nand NAND2 (N5113, N5103, N4442);
and AND3 (N5114, N5092, N10, N2566);
xor XOR2 (N5115, N5114, N1688);
nand NAND3 (N5116, N5106, N3986, N4391);
nand NAND4 (N5117, N5109, N4733, N5096, N2869);
nor NOR3 (N5118, N5112, N994, N1103);
or OR2 (N5119, N5107, N1957);
nor NOR4 (N5120, N5118, N3110, N881, N3086);
and AND2 (N5121, N5095, N1841);
and AND4 (N5122, N5120, N3439, N1017, N2615);
or OR3 (N5123, N5108, N2332, N3547);
and AND4 (N5124, N5119, N2095, N2521, N2997);
xor XOR2 (N5125, N5116, N4314);
nand NAND2 (N5126, N5124, N3728);
xor XOR2 (N5127, N5125, N4336);
nor NOR4 (N5128, N5126, N959, N4167, N165);
and AND4 (N5129, N5123, N1433, N1009, N4239);
not NOT1 (N5130, N5115);
buf BUF1 (N5131, N5122);
or OR4 (N5132, N5129, N3328, N3484, N210);
nor NOR4 (N5133, N5130, N3318, N4956, N1074);
nor NOR2 (N5134, N5080, N288);
nand NAND4 (N5135, N5127, N2791, N1599, N1860);
nor NOR4 (N5136, N5131, N1337, N4035, N2898);
and AND3 (N5137, N5121, N1204, N5128);
not NOT1 (N5138, N2690);
xor XOR2 (N5139, N5134, N4418);
not NOT1 (N5140, N5098);
and AND2 (N5141, N5133, N719);
or OR2 (N5142, N5132, N2304);
buf BUF1 (N5143, N5138);
not NOT1 (N5144, N5139);
nand NAND2 (N5145, N5140, N989);
and AND2 (N5146, N5142, N3821);
not NOT1 (N5147, N5141);
nor NOR3 (N5148, N5145, N2661, N3104);
or OR2 (N5149, N5137, N3971);
not NOT1 (N5150, N5149);
or OR3 (N5151, N5146, N3841, N2844);
not NOT1 (N5152, N5117);
and AND3 (N5153, N5143, N967, N2244);
not NOT1 (N5154, N5153);
not NOT1 (N5155, N5144);
not NOT1 (N5156, N5136);
xor XOR2 (N5157, N5113, N3904);
nor NOR3 (N5158, N5157, N3607, N432);
or OR2 (N5159, N5158, N4844);
and AND2 (N5160, N5135, N4873);
nor NOR4 (N5161, N5150, N3755, N3050, N1923);
or OR2 (N5162, N5147, N13);
or OR2 (N5163, N5159, N227);
and AND3 (N5164, N5152, N1605, N4694);
not NOT1 (N5165, N5160);
nand NAND4 (N5166, N5156, N2194, N1609, N987);
buf BUF1 (N5167, N5162);
buf BUF1 (N5168, N5166);
or OR3 (N5169, N5148, N4515, N1613);
nor NOR3 (N5170, N5161, N2317, N3323);
or OR4 (N5171, N5163, N1196, N575, N654);
and AND2 (N5172, N5155, N2096);
and AND4 (N5173, N5167, N3021, N3636, N802);
buf BUF1 (N5174, N5154);
nor NOR4 (N5175, N5174, N2442, N2708, N3944);
not NOT1 (N5176, N5171);
nand NAND4 (N5177, N5164, N4512, N2881, N1150);
nor NOR4 (N5178, N5176, N3492, N496, N733);
not NOT1 (N5179, N5151);
buf BUF1 (N5180, N5165);
and AND4 (N5181, N5173, N760, N5072, N1006);
xor XOR2 (N5182, N5175, N2394);
nor NOR3 (N5183, N5182, N2720, N493);
nand NAND2 (N5184, N5168, N478);
nand NAND2 (N5185, N5183, N1866);
xor XOR2 (N5186, N5179, N489);
xor XOR2 (N5187, N5177, N4166);
and AND2 (N5188, N5169, N715);
nor NOR3 (N5189, N5170, N4470, N4954);
nor NOR4 (N5190, N5187, N3263, N2723, N3245);
buf BUF1 (N5191, N5189);
buf BUF1 (N5192, N5181);
not NOT1 (N5193, N5192);
not NOT1 (N5194, N5185);
or OR3 (N5195, N5190, N3479, N4286);
buf BUF1 (N5196, N5188);
nor NOR3 (N5197, N5191, N4713, N2792);
or OR3 (N5198, N5172, N4564, N4434);
xor XOR2 (N5199, N5196, N5176);
nor NOR2 (N5200, N5197, N3240);
buf BUF1 (N5201, N5193);
nor NOR3 (N5202, N5194, N2705, N1072);
not NOT1 (N5203, N5184);
buf BUF1 (N5204, N5178);
not NOT1 (N5205, N5199);
nor NOR2 (N5206, N5198, N345);
buf BUF1 (N5207, N5186);
or OR3 (N5208, N5202, N3969, N3383);
buf BUF1 (N5209, N5205);
not NOT1 (N5210, N5208);
xor XOR2 (N5211, N5201, N49);
buf BUF1 (N5212, N5180);
xor XOR2 (N5213, N5209, N4163);
or OR4 (N5214, N5195, N364, N4646, N413);
nand NAND2 (N5215, N5212, N3846);
buf BUF1 (N5216, N5207);
nand NAND3 (N5217, N5214, N4374, N4305);
and AND4 (N5218, N5203, N1828, N843, N3019);
nand NAND3 (N5219, N5211, N609, N2588);
and AND2 (N5220, N5213, N2685);
nand NAND2 (N5221, N5200, N3139);
and AND4 (N5222, N5215, N1975, N3496, N2239);
xor XOR2 (N5223, N5217, N160);
and AND4 (N5224, N5221, N1258, N3569, N4024);
or OR2 (N5225, N5218, N1742);
buf BUF1 (N5226, N5224);
nor NOR2 (N5227, N5210, N2811);
xor XOR2 (N5228, N5226, N5171);
nor NOR2 (N5229, N5228, N3057);
nor NOR2 (N5230, N5204, N3685);
xor XOR2 (N5231, N5216, N4596);
buf BUF1 (N5232, N5223);
and AND2 (N5233, N5230, N4006);
and AND4 (N5234, N5206, N2792, N4661, N2387);
and AND2 (N5235, N5231, N1420);
and AND2 (N5236, N5219, N4622);
not NOT1 (N5237, N5222);
not NOT1 (N5238, N5225);
and AND2 (N5239, N5235, N3793);
and AND2 (N5240, N5229, N3310);
not NOT1 (N5241, N5237);
not NOT1 (N5242, N5234);
and AND4 (N5243, N5233, N5209, N764, N3718);
xor XOR2 (N5244, N5242, N40);
or OR2 (N5245, N5232, N1015);
nor NOR4 (N5246, N5245, N5184, N3278, N1844);
and AND4 (N5247, N5243, N462, N2418, N5246);
xor XOR2 (N5248, N3392, N2685);
or OR3 (N5249, N5236, N2173, N41);
buf BUF1 (N5250, N5249);
nand NAND2 (N5251, N5238, N4646);
nor NOR2 (N5252, N5241, N1576);
buf BUF1 (N5253, N5220);
xor XOR2 (N5254, N5240, N1307);
nand NAND4 (N5255, N5248, N3511, N3201, N3933);
xor XOR2 (N5256, N5250, N4217);
and AND4 (N5257, N5239, N3061, N2176, N2528);
nand NAND4 (N5258, N5251, N3574, N3532, N4518);
nand NAND3 (N5259, N5256, N354, N4085);
xor XOR2 (N5260, N5247, N3709);
xor XOR2 (N5261, N5255, N665);
or OR3 (N5262, N5259, N4151, N4200);
not NOT1 (N5263, N5252);
nand NAND3 (N5264, N5261, N4890, N5137);
nand NAND4 (N5265, N5260, N2550, N398, N3544);
buf BUF1 (N5266, N5257);
nor NOR3 (N5267, N5254, N3522, N1838);
nand NAND4 (N5268, N5262, N30, N4307, N3028);
not NOT1 (N5269, N5266);
nand NAND4 (N5270, N5244, N2445, N3097, N3509);
buf BUF1 (N5271, N5269);
nand NAND4 (N5272, N5267, N3767, N1274, N1524);
and AND2 (N5273, N5263, N679);
and AND2 (N5274, N5227, N4375);
buf BUF1 (N5275, N5270);
nand NAND4 (N5276, N5253, N3027, N1204, N70);
nor NOR3 (N5277, N5264, N5152, N457);
nand NAND3 (N5278, N5274, N3266, N2037);
buf BUF1 (N5279, N5265);
buf BUF1 (N5280, N5275);
and AND2 (N5281, N5258, N1132);
buf BUF1 (N5282, N5272);
and AND3 (N5283, N5280, N4015, N2556);
or OR3 (N5284, N5277, N643, N473);
buf BUF1 (N5285, N5284);
nor NOR2 (N5286, N5279, N3427);
buf BUF1 (N5287, N5273);
xor XOR2 (N5288, N5283, N3570);
nand NAND2 (N5289, N5268, N1385);
and AND2 (N5290, N5289, N5);
not NOT1 (N5291, N5276);
nand NAND2 (N5292, N5281, N1490);
buf BUF1 (N5293, N5271);
nor NOR3 (N5294, N5288, N568, N3211);
buf BUF1 (N5295, N5293);
or OR3 (N5296, N5282, N428, N1037);
nor NOR2 (N5297, N5294, N3523);
nand NAND4 (N5298, N5287, N4826, N4262, N2659);
or OR3 (N5299, N5292, N2202, N5104);
and AND2 (N5300, N5290, N5253);
buf BUF1 (N5301, N5295);
nand NAND4 (N5302, N5299, N2325, N4871, N2516);
nand NAND4 (N5303, N5300, N4623, N3404, N4843);
nor NOR3 (N5304, N5302, N287, N2674);
or OR3 (N5305, N5301, N3603, N31);
xor XOR2 (N5306, N5278, N4927);
not NOT1 (N5307, N5285);
not NOT1 (N5308, N5297);
or OR3 (N5309, N5291, N1839, N5137);
or OR3 (N5310, N5286, N144, N2639);
nor NOR2 (N5311, N5304, N918);
or OR4 (N5312, N5311, N481, N1954, N969);
nor NOR4 (N5313, N5309, N4671, N409, N2401);
buf BUF1 (N5314, N5308);
buf BUF1 (N5315, N5307);
nor NOR4 (N5316, N5298, N1954, N3610, N2572);
or OR4 (N5317, N5315, N4883, N4311, N4045);
or OR3 (N5318, N5314, N2620, N174);
and AND3 (N5319, N5303, N1603, N2925);
nor NOR3 (N5320, N5319, N2819, N2537);
or OR2 (N5321, N5296, N4494);
or OR4 (N5322, N5310, N2080, N2944, N2421);
and AND4 (N5323, N5305, N4347, N2939, N5283);
nand NAND3 (N5324, N5321, N1564, N3141);
xor XOR2 (N5325, N5313, N2424);
nand NAND2 (N5326, N5322, N3996);
or OR3 (N5327, N5320, N3394, N4353);
buf BUF1 (N5328, N5324);
buf BUF1 (N5329, N5327);
nor NOR4 (N5330, N5312, N2035, N4812, N381);
nor NOR4 (N5331, N5329, N2960, N2134, N2441);
and AND3 (N5332, N5330, N4298, N4824);
and AND4 (N5333, N5326, N3647, N1139, N2660);
nor NOR4 (N5334, N5306, N4246, N4118, N4318);
and AND2 (N5335, N5331, N5262);
not NOT1 (N5336, N5333);
not NOT1 (N5337, N5328);
or OR2 (N5338, N5318, N4319);
nand NAND3 (N5339, N5334, N5047, N2924);
and AND4 (N5340, N5337, N3327, N1018, N510);
not NOT1 (N5341, N5323);
nor NOR2 (N5342, N5335, N2611);
xor XOR2 (N5343, N5339, N14);
nand NAND4 (N5344, N5338, N4602, N2685, N3640);
xor XOR2 (N5345, N5316, N3601);
nor NOR2 (N5346, N5317, N5174);
xor XOR2 (N5347, N5343, N2267);
and AND3 (N5348, N5336, N5113, N5063);
xor XOR2 (N5349, N5325, N2490);
or OR3 (N5350, N5340, N4693, N2311);
or OR3 (N5351, N5346, N1498, N2405);
xor XOR2 (N5352, N5344, N879);
or OR3 (N5353, N5351, N1425, N5295);
not NOT1 (N5354, N5349);
not NOT1 (N5355, N5342);
buf BUF1 (N5356, N5348);
or OR3 (N5357, N5355, N151, N3);
xor XOR2 (N5358, N5350, N1595);
not NOT1 (N5359, N5358);
xor XOR2 (N5360, N5332, N1507);
nor NOR3 (N5361, N5359, N280, N2502);
and AND2 (N5362, N5347, N4742);
and AND3 (N5363, N5356, N1503, N2460);
and AND2 (N5364, N5341, N3606);
nand NAND2 (N5365, N5364, N3772);
xor XOR2 (N5366, N5345, N4044);
or OR2 (N5367, N5362, N1038);
nor NOR3 (N5368, N5352, N670, N230);
xor XOR2 (N5369, N5365, N5080);
xor XOR2 (N5370, N5357, N2912);
nand NAND2 (N5371, N5369, N2091);
or OR3 (N5372, N5354, N405, N3174);
xor XOR2 (N5373, N5372, N3022);
xor XOR2 (N5374, N5368, N1095);
or OR4 (N5375, N5361, N4917, N1553, N122);
xor XOR2 (N5376, N5366, N2102);
buf BUF1 (N5377, N5360);
xor XOR2 (N5378, N5353, N1314);
nand NAND3 (N5379, N5374, N4232, N729);
nand NAND2 (N5380, N5377, N2867);
buf BUF1 (N5381, N5367);
and AND3 (N5382, N5381, N1384, N2335);
buf BUF1 (N5383, N5379);
not NOT1 (N5384, N5373);
nand NAND2 (N5385, N5363, N2850);
buf BUF1 (N5386, N5376);
or OR4 (N5387, N5375, N864, N4497, N3532);
not NOT1 (N5388, N5378);
nor NOR3 (N5389, N5383, N4990, N3106);
or OR2 (N5390, N5389, N332);
or OR4 (N5391, N5382, N1222, N2439, N2731);
nand NAND4 (N5392, N5384, N1493, N1330, N4577);
and AND3 (N5393, N5371, N4262, N2764);
not NOT1 (N5394, N5370);
not NOT1 (N5395, N5391);
buf BUF1 (N5396, N5380);
buf BUF1 (N5397, N5385);
nor NOR4 (N5398, N5386, N803, N420, N730);
nor NOR4 (N5399, N5390, N1905, N498, N1233);
nand NAND4 (N5400, N5399, N4286, N5136, N3606);
not NOT1 (N5401, N5395);
nand NAND2 (N5402, N5400, N4267);
xor XOR2 (N5403, N5401, N4056);
buf BUF1 (N5404, N5398);
not NOT1 (N5405, N5403);
nor NOR2 (N5406, N5396, N1380);
xor XOR2 (N5407, N5402, N4274);
buf BUF1 (N5408, N5397);
and AND4 (N5409, N5394, N4389, N5113, N4699);
xor XOR2 (N5410, N5405, N260);
and AND2 (N5411, N5406, N4176);
or OR2 (N5412, N5387, N277);
not NOT1 (N5413, N5393);
buf BUF1 (N5414, N5409);
nand NAND4 (N5415, N5413, N1845, N4620, N4283);
nand NAND4 (N5416, N5407, N1810, N5097, N807);
nand NAND4 (N5417, N5416, N920, N1376, N974);
nand NAND3 (N5418, N5410, N4572, N5057);
not NOT1 (N5419, N5417);
nor NOR4 (N5420, N5392, N1301, N4964, N12);
nor NOR2 (N5421, N5419, N1866);
nand NAND3 (N5422, N5388, N4717, N1059);
nor NOR4 (N5423, N5408, N4510, N2467, N237);
and AND4 (N5424, N5418, N4721, N4385, N5167);
and AND4 (N5425, N5420, N170, N4934, N2090);
not NOT1 (N5426, N5424);
nand NAND3 (N5427, N5411, N642, N5051);
or OR3 (N5428, N5423, N2542, N2225);
nand NAND2 (N5429, N5428, N2764);
or OR4 (N5430, N5422, N5104, N2442, N4655);
nor NOR3 (N5431, N5404, N3202, N2809);
nand NAND2 (N5432, N5415, N4898);
not NOT1 (N5433, N5432);
buf BUF1 (N5434, N5433);
nor NOR3 (N5435, N5431, N4399, N4760);
not NOT1 (N5436, N5435);
buf BUF1 (N5437, N5436);
nor NOR2 (N5438, N5427, N4924);
xor XOR2 (N5439, N5438, N4214);
nand NAND3 (N5440, N5434, N2026, N3978);
and AND3 (N5441, N5412, N4420, N3842);
buf BUF1 (N5442, N5430);
or OR4 (N5443, N5425, N35, N131, N4557);
and AND4 (N5444, N5440, N4507, N4211, N3590);
buf BUF1 (N5445, N5437);
buf BUF1 (N5446, N5442);
nand NAND3 (N5447, N5443, N4560, N4006);
and AND2 (N5448, N5447, N3288);
and AND4 (N5449, N5429, N3236, N22, N2479);
nor NOR2 (N5450, N5446, N2187);
and AND2 (N5451, N5439, N2601);
xor XOR2 (N5452, N5445, N2762);
xor XOR2 (N5453, N5421, N416);
nor NOR4 (N5454, N5448, N2051, N3384, N4820);
buf BUF1 (N5455, N5452);
nor NOR2 (N5456, N5426, N3752);
or OR4 (N5457, N5455, N3721, N320, N595);
not NOT1 (N5458, N5450);
buf BUF1 (N5459, N5451);
not NOT1 (N5460, N5454);
and AND4 (N5461, N5457, N5228, N1620, N4391);
or OR4 (N5462, N5456, N4291, N734, N4290);
nand NAND2 (N5463, N5460, N5265);
not NOT1 (N5464, N5463);
xor XOR2 (N5465, N5464, N5090);
not NOT1 (N5466, N5458);
nand NAND3 (N5467, N5414, N46, N5155);
buf BUF1 (N5468, N5465);
not NOT1 (N5469, N5461);
or OR4 (N5470, N5462, N3646, N3176, N3289);
or OR4 (N5471, N5449, N3835, N509, N1015);
or OR2 (N5472, N5453, N732);
buf BUF1 (N5473, N5469);
xor XOR2 (N5474, N5459, N263);
nor NOR4 (N5475, N5468, N3750, N4617, N1143);
or OR2 (N5476, N5470, N4700);
nand NAND3 (N5477, N5475, N3972, N3228);
or OR2 (N5478, N5471, N4088);
xor XOR2 (N5479, N5472, N4619);
not NOT1 (N5480, N5444);
nor NOR2 (N5481, N5479, N441);
not NOT1 (N5482, N5467);
not NOT1 (N5483, N5476);
xor XOR2 (N5484, N5478, N2199);
and AND2 (N5485, N5481, N1457);
buf BUF1 (N5486, N5466);
not NOT1 (N5487, N5484);
buf BUF1 (N5488, N5474);
buf BUF1 (N5489, N5485);
or OR4 (N5490, N5441, N3472, N4194, N1696);
xor XOR2 (N5491, N5480, N3185);
nand NAND4 (N5492, N5486, N3638, N5248, N1515);
nand NAND3 (N5493, N5492, N4183, N4777);
buf BUF1 (N5494, N5488);
buf BUF1 (N5495, N5473);
and AND2 (N5496, N5482, N1157);
or OR4 (N5497, N5490, N5352, N2267, N4206);
xor XOR2 (N5498, N5497, N2227);
nor NOR4 (N5499, N5495, N3394, N216, N1133);
xor XOR2 (N5500, N5477, N4624);
xor XOR2 (N5501, N5498, N4745);
nor NOR2 (N5502, N5487, N243);
nor NOR4 (N5503, N5489, N4687, N1797, N981);
xor XOR2 (N5504, N5500, N3642);
xor XOR2 (N5505, N5501, N5027);
nand NAND2 (N5506, N5499, N5464);
xor XOR2 (N5507, N5483, N335);
not NOT1 (N5508, N5504);
nand NAND4 (N5509, N5496, N78, N198, N3407);
xor XOR2 (N5510, N5502, N992);
nand NAND4 (N5511, N5491, N4684, N816, N1375);
and AND2 (N5512, N5509, N2065);
nor NOR4 (N5513, N5493, N761, N2777, N3099);
nor NOR3 (N5514, N5511, N4405, N1952);
or OR2 (N5515, N5508, N4270);
and AND4 (N5516, N5513, N2067, N1217, N4263);
and AND4 (N5517, N5494, N3889, N5238, N1385);
nand NAND2 (N5518, N5516, N2028);
xor XOR2 (N5519, N5507, N360);
not NOT1 (N5520, N5514);
buf BUF1 (N5521, N5503);
nand NAND3 (N5522, N5515, N4426, N4033);
nor NOR3 (N5523, N5506, N5175, N1186);
not NOT1 (N5524, N5510);
nand NAND3 (N5525, N5519, N3540, N2399);
and AND4 (N5526, N5525, N4670, N1228, N2461);
buf BUF1 (N5527, N5517);
or OR4 (N5528, N5520, N2666, N5484, N2824);
and AND3 (N5529, N5526, N1428, N4376);
not NOT1 (N5530, N5512);
nor NOR3 (N5531, N5518, N1070, N3711);
nand NAND4 (N5532, N5524, N510, N349, N2649);
nand NAND4 (N5533, N5531, N794, N843, N3525);
not NOT1 (N5534, N5529);
buf BUF1 (N5535, N5530);
not NOT1 (N5536, N5521);
buf BUF1 (N5537, N5534);
or OR4 (N5538, N5537, N1456, N2720, N4305);
buf BUF1 (N5539, N5527);
buf BUF1 (N5540, N5538);
and AND4 (N5541, N5540, N4521, N974, N3991);
nand NAND2 (N5542, N5539, N1446);
not NOT1 (N5543, N5532);
nor NOR3 (N5544, N5505, N360, N66);
and AND3 (N5545, N5541, N600, N2385);
and AND2 (N5546, N5543, N4776);
buf BUF1 (N5547, N5522);
nand NAND4 (N5548, N5545, N3835, N1962, N897);
buf BUF1 (N5549, N5542);
buf BUF1 (N5550, N5548);
or OR3 (N5551, N5535, N3891, N4219);
or OR2 (N5552, N5547, N5251);
nor NOR2 (N5553, N5550, N1505);
nor NOR2 (N5554, N5523, N5313);
nand NAND4 (N5555, N5544, N3631, N417, N1914);
nor NOR3 (N5556, N5555, N304, N4558);
buf BUF1 (N5557, N5536);
xor XOR2 (N5558, N5533, N1001);
buf BUF1 (N5559, N5528);
buf BUF1 (N5560, N5556);
xor XOR2 (N5561, N5546, N1216);
nand NAND4 (N5562, N5554, N5211, N3625, N1034);
xor XOR2 (N5563, N5561, N1182);
or OR4 (N5564, N5551, N3285, N2446, N4643);
nand NAND4 (N5565, N5563, N1291, N1357, N448);
or OR4 (N5566, N5558, N3732, N1168, N110);
or OR4 (N5567, N5552, N2754, N1255, N4346);
xor XOR2 (N5568, N5553, N1947);
buf BUF1 (N5569, N5549);
or OR3 (N5570, N5566, N267, N640);
nor NOR3 (N5571, N5564, N5336, N3122);
buf BUF1 (N5572, N5567);
buf BUF1 (N5573, N5557);
or OR2 (N5574, N5568, N4179);
nand NAND2 (N5575, N5562, N4042);
xor XOR2 (N5576, N5565, N2770);
not NOT1 (N5577, N5569);
xor XOR2 (N5578, N5571, N1968);
or OR2 (N5579, N5572, N2447);
and AND3 (N5580, N5570, N2484, N1953);
buf BUF1 (N5581, N5576);
xor XOR2 (N5582, N5575, N2908);
xor XOR2 (N5583, N5560, N2054);
xor XOR2 (N5584, N5578, N2659);
xor XOR2 (N5585, N5581, N2453);
xor XOR2 (N5586, N5583, N1656);
or OR2 (N5587, N5559, N5409);
nor NOR3 (N5588, N5577, N2440, N5179);
or OR2 (N5589, N5585, N1787);
and AND2 (N5590, N5582, N1437);
buf BUF1 (N5591, N5574);
not NOT1 (N5592, N5587);
not NOT1 (N5593, N5591);
or OR2 (N5594, N5579, N630);
or OR2 (N5595, N5573, N4142);
xor XOR2 (N5596, N5595, N958);
not NOT1 (N5597, N5586);
not NOT1 (N5598, N5596);
nor NOR4 (N5599, N5589, N3301, N1786, N1938);
not NOT1 (N5600, N5588);
and AND3 (N5601, N5580, N1036, N1299);
and AND2 (N5602, N5601, N4078);
buf BUF1 (N5603, N5597);
not NOT1 (N5604, N5584);
buf BUF1 (N5605, N5592);
and AND3 (N5606, N5600, N271, N2021);
nor NOR3 (N5607, N5598, N1081, N5266);
not NOT1 (N5608, N5603);
not NOT1 (N5609, N5606);
xor XOR2 (N5610, N5599, N5484);
nand NAND2 (N5611, N5605, N851);
xor XOR2 (N5612, N5602, N5267);
nand NAND2 (N5613, N5607, N2140);
and AND3 (N5614, N5593, N5393, N5185);
nand NAND3 (N5615, N5594, N3536, N2383);
not NOT1 (N5616, N5604);
and AND4 (N5617, N5590, N1820, N5148, N812);
nand NAND3 (N5618, N5609, N5318, N1556);
and AND4 (N5619, N5616, N2212, N846, N3981);
or OR3 (N5620, N5610, N4119, N1655);
or OR4 (N5621, N5608, N3774, N3881, N745);
and AND2 (N5622, N5619, N1286);
nand NAND4 (N5623, N5613, N4838, N3384, N284);
buf BUF1 (N5624, N5618);
not NOT1 (N5625, N5623);
and AND2 (N5626, N5624, N2751);
or OR4 (N5627, N5617, N4033, N457, N1730);
buf BUF1 (N5628, N5611);
or OR4 (N5629, N5614, N5192, N3184, N5030);
xor XOR2 (N5630, N5612, N4092);
nor NOR3 (N5631, N5627, N5043, N4410);
xor XOR2 (N5632, N5620, N1838);
nor NOR2 (N5633, N5625, N159);
and AND2 (N5634, N5632, N4971);
not NOT1 (N5635, N5626);
buf BUF1 (N5636, N5622);
nand NAND2 (N5637, N5630, N4544);
nor NOR2 (N5638, N5628, N3081);
xor XOR2 (N5639, N5621, N2663);
or OR3 (N5640, N5629, N4556, N2483);
xor XOR2 (N5641, N5640, N3875);
nor NOR4 (N5642, N5615, N1237, N4276, N3974);
not NOT1 (N5643, N5633);
not NOT1 (N5644, N5641);
not NOT1 (N5645, N5637);
and AND4 (N5646, N5644, N3424, N1936, N3949);
not NOT1 (N5647, N5635);
nor NOR4 (N5648, N5647, N5326, N263, N5619);
nand NAND4 (N5649, N5634, N4382, N1576, N2369);
nand NAND2 (N5650, N5642, N4708);
and AND4 (N5651, N5636, N83, N2279, N1333);
not NOT1 (N5652, N5650);
xor XOR2 (N5653, N5631, N876);
nand NAND2 (N5654, N5648, N4637);
xor XOR2 (N5655, N5643, N3929);
not NOT1 (N5656, N5652);
buf BUF1 (N5657, N5646);
nand NAND4 (N5658, N5649, N5444, N2538, N5657);
and AND2 (N5659, N662, N3610);
and AND3 (N5660, N5639, N800, N2857);
nor NOR4 (N5661, N5656, N945, N1737, N1899);
xor XOR2 (N5662, N5654, N2695);
not NOT1 (N5663, N5662);
buf BUF1 (N5664, N5659);
xor XOR2 (N5665, N5658, N1277);
or OR4 (N5666, N5660, N2735, N3338, N3718);
xor XOR2 (N5667, N5645, N1900);
and AND4 (N5668, N5663, N505, N1006, N74);
and AND2 (N5669, N5655, N4384);
and AND2 (N5670, N5664, N3286);
or OR3 (N5671, N5668, N785, N2377);
and AND4 (N5672, N5661, N145, N2150, N3583);
xor XOR2 (N5673, N5667, N2194);
and AND2 (N5674, N5672, N990);
nor NOR3 (N5675, N5666, N2931, N295);
xor XOR2 (N5676, N5665, N5018);
xor XOR2 (N5677, N5676, N601);
and AND2 (N5678, N5638, N5366);
not NOT1 (N5679, N5673);
nand NAND3 (N5680, N5674, N3423, N710);
nor NOR2 (N5681, N5680, N2355);
xor XOR2 (N5682, N5681, N3164);
nor NOR2 (N5683, N5678, N2586);
nand NAND4 (N5684, N5670, N3220, N3579, N909);
or OR3 (N5685, N5675, N2097, N1021);
buf BUF1 (N5686, N5671);
nand NAND3 (N5687, N5679, N2132, N4128);
xor XOR2 (N5688, N5683, N4261);
nor NOR4 (N5689, N5653, N4613, N1713, N1090);
xor XOR2 (N5690, N5689, N1391);
and AND4 (N5691, N5687, N2894, N1537, N2074);
nor NOR4 (N5692, N5690, N4963, N713, N4586);
and AND2 (N5693, N5651, N3937);
and AND4 (N5694, N5684, N4580, N5066, N1143);
nand NAND4 (N5695, N5688, N3708, N2968, N3625);
or OR2 (N5696, N5694, N3615);
nor NOR3 (N5697, N5692, N2871, N4706);
not NOT1 (N5698, N5696);
buf BUF1 (N5699, N5677);
xor XOR2 (N5700, N5695, N5100);
nand NAND3 (N5701, N5691, N1181, N2618);
buf BUF1 (N5702, N5698);
and AND2 (N5703, N5700, N3458);
or OR2 (N5704, N5699, N2360);
nor NOR2 (N5705, N5704, N121);
buf BUF1 (N5706, N5686);
nor NOR3 (N5707, N5682, N3374, N1006);
and AND4 (N5708, N5697, N4106, N4853, N2958);
not NOT1 (N5709, N5685);
nor NOR3 (N5710, N5701, N3964, N5214);
or OR2 (N5711, N5669, N5031);
nand NAND4 (N5712, N5705, N989, N4073, N1085);
or OR2 (N5713, N5710, N2542);
xor XOR2 (N5714, N5702, N3381);
xor XOR2 (N5715, N5714, N5086);
or OR4 (N5716, N5707, N1215, N1254, N3338);
xor XOR2 (N5717, N5712, N4186);
xor XOR2 (N5718, N5716, N503);
buf BUF1 (N5719, N5715);
xor XOR2 (N5720, N5713, N3235);
nor NOR3 (N5721, N5719, N4764, N987);
buf BUF1 (N5722, N5721);
nand NAND4 (N5723, N5711, N1977, N3225, N2249);
and AND2 (N5724, N5722, N2201);
or OR3 (N5725, N5720, N402, N4170);
xor XOR2 (N5726, N5717, N4926);
buf BUF1 (N5727, N5725);
nor NOR2 (N5728, N5706, N3612);
buf BUF1 (N5729, N5709);
or OR2 (N5730, N5693, N1429);
xor XOR2 (N5731, N5729, N1557);
buf BUF1 (N5732, N5730);
or OR4 (N5733, N5723, N1867, N3119, N1716);
xor XOR2 (N5734, N5728, N5214);
or OR3 (N5735, N5708, N5012, N3503);
buf BUF1 (N5736, N5735);
xor XOR2 (N5737, N5731, N4567);
buf BUF1 (N5738, N5737);
nor NOR2 (N5739, N5727, N4912);
nand NAND4 (N5740, N5724, N224, N225, N4126);
nand NAND4 (N5741, N5736, N5211, N5109, N4587);
and AND3 (N5742, N5718, N5499, N3266);
xor XOR2 (N5743, N5740, N2130);
nand NAND4 (N5744, N5742, N2401, N117, N3207);
buf BUF1 (N5745, N5744);
and AND3 (N5746, N5734, N3302, N1560);
xor XOR2 (N5747, N5745, N3241);
nor NOR4 (N5748, N5747, N2910, N802, N3771);
buf BUF1 (N5749, N5743);
xor XOR2 (N5750, N5739, N1854);
buf BUF1 (N5751, N5726);
xor XOR2 (N5752, N5750, N5241);
not NOT1 (N5753, N5748);
buf BUF1 (N5754, N5738);
and AND2 (N5755, N5732, N3751);
not NOT1 (N5756, N5752);
buf BUF1 (N5757, N5756);
nor NOR2 (N5758, N5753, N751);
xor XOR2 (N5759, N5746, N5687);
xor XOR2 (N5760, N5755, N3406);
or OR2 (N5761, N5751, N3356);
xor XOR2 (N5762, N5758, N2271);
not NOT1 (N5763, N5754);
or OR3 (N5764, N5749, N4855, N2461);
nor NOR3 (N5765, N5733, N3728, N4895);
buf BUF1 (N5766, N5757);
and AND2 (N5767, N5764, N2373);
and AND4 (N5768, N5762, N5286, N3806, N5349);
xor XOR2 (N5769, N5760, N4574);
nor NOR2 (N5770, N5767, N3300);
not NOT1 (N5771, N5741);
or OR2 (N5772, N5769, N2676);
not NOT1 (N5773, N5768);
nor NOR2 (N5774, N5759, N3941);
and AND4 (N5775, N5772, N2611, N5324, N4632);
buf BUF1 (N5776, N5773);
buf BUF1 (N5777, N5761);
not NOT1 (N5778, N5776);
xor XOR2 (N5779, N5775, N672);
nor NOR3 (N5780, N5778, N1992, N2362);
buf BUF1 (N5781, N5703);
or OR3 (N5782, N5765, N534, N349);
nor NOR3 (N5783, N5781, N2611, N5590);
nand NAND4 (N5784, N5779, N214, N4653, N4664);
not NOT1 (N5785, N5784);
or OR4 (N5786, N5780, N5208, N2494, N4296);
not NOT1 (N5787, N5783);
xor XOR2 (N5788, N5766, N4599);
buf BUF1 (N5789, N5785);
or OR3 (N5790, N5786, N3753, N4007);
nor NOR2 (N5791, N5770, N4091);
and AND2 (N5792, N5777, N1086);
nor NOR2 (N5793, N5763, N2310);
or OR4 (N5794, N5791, N4043, N4375, N3860);
nand NAND2 (N5795, N5788, N979);
or OR4 (N5796, N5792, N4340, N447, N3561);
or OR2 (N5797, N5789, N5175);
xor XOR2 (N5798, N5774, N5559);
and AND4 (N5799, N5790, N3692, N5511, N1613);
and AND4 (N5800, N5771, N3896, N2859, N3264);
nand NAND3 (N5801, N5798, N1201, N2097);
nand NAND4 (N5802, N5796, N1225, N58, N1098);
not NOT1 (N5803, N5795);
not NOT1 (N5804, N5793);
buf BUF1 (N5805, N5803);
nand NAND2 (N5806, N5800, N3419);
nand NAND3 (N5807, N5794, N4545, N2208);
xor XOR2 (N5808, N5804, N3738);
nor NOR3 (N5809, N5787, N2272, N1024);
not NOT1 (N5810, N5807);
not NOT1 (N5811, N5797);
or OR3 (N5812, N5801, N3855, N5804);
buf BUF1 (N5813, N5806);
not NOT1 (N5814, N5810);
nand NAND2 (N5815, N5811, N5540);
not NOT1 (N5816, N5808);
or OR2 (N5817, N5799, N4648);
nor NOR4 (N5818, N5805, N4159, N1944, N5224);
or OR2 (N5819, N5813, N1721);
nand NAND4 (N5820, N5817, N2774, N2347, N1353);
or OR4 (N5821, N5814, N2500, N2558, N4180);
or OR3 (N5822, N5821, N912, N2655);
and AND3 (N5823, N5782, N1525, N763);
and AND2 (N5824, N5812, N5078);
or OR4 (N5825, N5824, N2921, N3725, N5392);
nand NAND3 (N5826, N5809, N1548, N422);
not NOT1 (N5827, N5823);
nor NOR3 (N5828, N5827, N1348, N1488);
not NOT1 (N5829, N5818);
and AND2 (N5830, N5826, N3063);
nor NOR4 (N5831, N5829, N4381, N2183, N4118);
nor NOR4 (N5832, N5820, N4414, N1075, N2900);
or OR3 (N5833, N5819, N2126, N4845);
and AND4 (N5834, N5830, N1162, N2160, N2582);
xor XOR2 (N5835, N5831, N3999);
not NOT1 (N5836, N5832);
nor NOR3 (N5837, N5815, N1526, N3088);
not NOT1 (N5838, N5816);
xor XOR2 (N5839, N5838, N5692);
not NOT1 (N5840, N5839);
not NOT1 (N5841, N5822);
and AND3 (N5842, N5837, N5815, N4220);
buf BUF1 (N5843, N5840);
not NOT1 (N5844, N5842);
or OR4 (N5845, N5802, N2288, N1778, N1880);
nor NOR2 (N5846, N5834, N5657);
xor XOR2 (N5847, N5825, N3904);
not NOT1 (N5848, N5841);
not NOT1 (N5849, N5843);
or OR2 (N5850, N5836, N1361);
or OR4 (N5851, N5844, N3975, N5399, N3481);
xor XOR2 (N5852, N5846, N1479);
xor XOR2 (N5853, N5852, N3603);
nand NAND4 (N5854, N5850, N4351, N989, N2007);
nand NAND3 (N5855, N5849, N5116, N3492);
or OR4 (N5856, N5851, N2269, N5147, N723);
not NOT1 (N5857, N5856);
nand NAND3 (N5858, N5857, N4865, N2408);
nand NAND3 (N5859, N5853, N3783, N879);
and AND4 (N5860, N5835, N4192, N5035, N5573);
nand NAND2 (N5861, N5848, N3536);
not NOT1 (N5862, N5828);
buf BUF1 (N5863, N5860);
and AND2 (N5864, N5855, N3071);
and AND4 (N5865, N5854, N5102, N4466, N980);
nor NOR2 (N5866, N5847, N1535);
nor NOR3 (N5867, N5861, N135, N334);
and AND2 (N5868, N5864, N1987);
or OR3 (N5869, N5866, N4092, N1907);
not NOT1 (N5870, N5865);
and AND2 (N5871, N5858, N2469);
nor NOR2 (N5872, N5868, N5468);
nand NAND3 (N5873, N5863, N1972, N605);
buf BUF1 (N5874, N5862);
nand NAND3 (N5875, N5869, N1544, N665);
xor XOR2 (N5876, N5871, N4136);
nand NAND4 (N5877, N5833, N1574, N2102, N4890);
or OR2 (N5878, N5877, N3513);
xor XOR2 (N5879, N5859, N1360);
nand NAND2 (N5880, N5872, N5238);
nor NOR4 (N5881, N5875, N3431, N4086, N1518);
nor NOR2 (N5882, N5881, N4595);
nand NAND3 (N5883, N5882, N4630, N5156);
not NOT1 (N5884, N5880);
nor NOR2 (N5885, N5867, N4827);
nand NAND2 (N5886, N5845, N3909);
xor XOR2 (N5887, N5874, N3329);
or OR3 (N5888, N5883, N1090, N3285);
and AND3 (N5889, N5878, N2225, N1302);
not NOT1 (N5890, N5884);
nand NAND4 (N5891, N5873, N5663, N5650, N3230);
xor XOR2 (N5892, N5890, N3809);
nor NOR2 (N5893, N5876, N435);
buf BUF1 (N5894, N5888);
and AND4 (N5895, N5886, N3201, N1100, N84);
nor NOR4 (N5896, N5891, N4015, N2219, N346);
or OR3 (N5897, N5896, N5825, N1151);
or OR4 (N5898, N5885, N3820, N3374, N1411);
not NOT1 (N5899, N5894);
not NOT1 (N5900, N5889);
nor NOR4 (N5901, N5887, N5466, N4375, N4838);
nor NOR4 (N5902, N5879, N4482, N2364, N4487);
nor NOR4 (N5903, N5901, N2103, N1134, N2252);
xor XOR2 (N5904, N5899, N794);
nor NOR3 (N5905, N5900, N1058, N2092);
xor XOR2 (N5906, N5893, N3358);
xor XOR2 (N5907, N5870, N1653);
nor NOR2 (N5908, N5898, N415);
nand NAND2 (N5909, N5905, N3634);
nor NOR2 (N5910, N5892, N1082);
or OR3 (N5911, N5902, N2084, N267);
buf BUF1 (N5912, N5906);
nor NOR2 (N5913, N5907, N2661);
nor NOR4 (N5914, N5913, N4162, N1066, N5279);
buf BUF1 (N5915, N5911);
buf BUF1 (N5916, N5904);
and AND2 (N5917, N5912, N437);
buf BUF1 (N5918, N5909);
nor NOR4 (N5919, N5903, N1065, N5246, N79);
nor NOR2 (N5920, N5915, N199);
and AND3 (N5921, N5920, N3006, N1642);
not NOT1 (N5922, N5918);
and AND3 (N5923, N5895, N3340, N770);
nand NAND2 (N5924, N5908, N192);
xor XOR2 (N5925, N5916, N5280);
nor NOR4 (N5926, N5922, N4889, N3185, N4467);
and AND4 (N5927, N5925, N4893, N5468, N5581);
nand NAND3 (N5928, N5923, N4066, N5333);
xor XOR2 (N5929, N5928, N5218);
xor XOR2 (N5930, N5921, N5780);
or OR2 (N5931, N5926, N3257);
xor XOR2 (N5932, N5924, N883);
xor XOR2 (N5933, N5927, N4889);
buf BUF1 (N5934, N5932);
nand NAND3 (N5935, N5917, N4712, N1783);
nor NOR2 (N5936, N5910, N174);
nand NAND4 (N5937, N5914, N5437, N1229, N1598);
and AND2 (N5938, N5930, N2739);
nand NAND2 (N5939, N5936, N4254);
buf BUF1 (N5940, N5919);
buf BUF1 (N5941, N5934);
nor NOR3 (N5942, N5931, N1910, N1769);
or OR3 (N5943, N5937, N2957, N2758);
or OR3 (N5944, N5938, N1687, N1394);
nor NOR2 (N5945, N5944, N1643);
nor NOR3 (N5946, N5897, N4002, N3597);
not NOT1 (N5947, N5945);
buf BUF1 (N5948, N5943);
and AND2 (N5949, N5948, N2621);
xor XOR2 (N5950, N5929, N4881);
or OR3 (N5951, N5941, N4873, N2515);
xor XOR2 (N5952, N5942, N4041);
nor NOR4 (N5953, N5949, N1928, N2902, N3755);
and AND2 (N5954, N5952, N4596);
and AND2 (N5955, N5933, N3291);
and AND2 (N5956, N5935, N159);
and AND4 (N5957, N5953, N5516, N2739, N2565);
nand NAND2 (N5958, N5956, N2814);
not NOT1 (N5959, N5957);
nor NOR4 (N5960, N5946, N5723, N364, N1297);
or OR3 (N5961, N5940, N1781, N364);
buf BUF1 (N5962, N5954);
or OR4 (N5963, N5961, N966, N2494, N5312);
and AND2 (N5964, N5958, N554);
nand NAND3 (N5965, N5950, N30, N4870);
xor XOR2 (N5966, N5963, N3467);
xor XOR2 (N5967, N5959, N3669);
or OR4 (N5968, N5947, N3814, N8, N5532);
nand NAND4 (N5969, N5964, N1759, N399, N2563);
or OR3 (N5970, N5965, N5323, N3871);
nand NAND3 (N5971, N5951, N3749, N4366);
and AND4 (N5972, N5955, N4456, N1947, N968);
nor NOR2 (N5973, N5970, N1639);
or OR2 (N5974, N5939, N272);
nor NOR3 (N5975, N5967, N27, N2939);
nand NAND2 (N5976, N5966, N4120);
and AND4 (N5977, N5960, N5154, N3884, N5802);
buf BUF1 (N5978, N5969);
nand NAND4 (N5979, N5971, N3526, N2541, N626);
xor XOR2 (N5980, N5968, N3415);
nand NAND4 (N5981, N5976, N1094, N2943, N989);
nor NOR3 (N5982, N5975, N5368, N1035);
nand NAND2 (N5983, N5962, N2389);
buf BUF1 (N5984, N5973);
and AND3 (N5985, N5974, N4267, N3252);
xor XOR2 (N5986, N5984, N5965);
nand NAND3 (N5987, N5981, N4570, N4836);
xor XOR2 (N5988, N5979, N5206);
or OR3 (N5989, N5986, N5213, N4147);
not NOT1 (N5990, N5977);
buf BUF1 (N5991, N5989);
nand NAND3 (N5992, N5972, N3528, N2525);
or OR2 (N5993, N5987, N4830);
buf BUF1 (N5994, N5980);
not NOT1 (N5995, N5982);
buf BUF1 (N5996, N5995);
nand NAND4 (N5997, N5990, N2689, N5268, N3575);
and AND3 (N5998, N5992, N5556, N3310);
buf BUF1 (N5999, N5996);
not NOT1 (N6000, N5993);
xor XOR2 (N6001, N5997, N373);
and AND4 (N6002, N6000, N4715, N5011, N127);
or OR4 (N6003, N5998, N412, N5732, N2332);
nand NAND2 (N6004, N5991, N1720);
buf BUF1 (N6005, N6002);
nor NOR3 (N6006, N5994, N394, N4057);
not NOT1 (N6007, N5988);
not NOT1 (N6008, N6007);
nand NAND2 (N6009, N6006, N2286);
not NOT1 (N6010, N6005);
not NOT1 (N6011, N5999);
nand NAND4 (N6012, N6001, N2165, N3498, N2649);
nand NAND2 (N6013, N6009, N1464);
nor NOR4 (N6014, N6004, N5224, N2356, N2516);
or OR3 (N6015, N6013, N4073, N5780);
xor XOR2 (N6016, N5978, N981);
buf BUF1 (N6017, N6008);
or OR4 (N6018, N6010, N4533, N3106, N2744);
nor NOR2 (N6019, N6003, N5821);
xor XOR2 (N6020, N6018, N1882);
nand NAND2 (N6021, N6017, N980);
xor XOR2 (N6022, N6020, N3089);
or OR2 (N6023, N6022, N1249);
nor NOR3 (N6024, N6012, N4879, N1151);
or OR2 (N6025, N5985, N3799);
nor NOR3 (N6026, N6019, N2340, N96);
nand NAND4 (N6027, N6026, N942, N901, N3523);
not NOT1 (N6028, N6027);
not NOT1 (N6029, N6016);
nor NOR3 (N6030, N6025, N1845, N1780);
nand NAND4 (N6031, N6023, N2728, N315, N4911);
not NOT1 (N6032, N6015);
nor NOR2 (N6033, N6030, N3410);
xor XOR2 (N6034, N5983, N4615);
buf BUF1 (N6035, N6034);
buf BUF1 (N6036, N6014);
xor XOR2 (N6037, N6021, N5300);
not NOT1 (N6038, N6032);
nand NAND3 (N6039, N6031, N1083, N474);
and AND4 (N6040, N6033, N619, N4677, N613);
nor NOR2 (N6041, N6011, N2443);
not NOT1 (N6042, N6040);
nor NOR4 (N6043, N6029, N704, N267, N2034);
and AND3 (N6044, N6039, N2862, N1562);
and AND4 (N6045, N6037, N5538, N3495, N3003);
buf BUF1 (N6046, N6043);
xor XOR2 (N6047, N6036, N1096);
nor NOR4 (N6048, N6046, N5328, N556, N4545);
and AND3 (N6049, N6028, N5691, N295);
buf BUF1 (N6050, N6048);
and AND3 (N6051, N6024, N4699, N2747);
or OR4 (N6052, N6045, N4791, N1494, N4486);
and AND3 (N6053, N6047, N1398, N2546);
xor XOR2 (N6054, N6042, N934);
or OR4 (N6055, N6044, N4633, N1993, N5235);
not NOT1 (N6056, N6051);
xor XOR2 (N6057, N6041, N2020);
or OR2 (N6058, N6057, N1042);
buf BUF1 (N6059, N6035);
or OR4 (N6060, N6058, N1515, N5948, N2479);
xor XOR2 (N6061, N6049, N1016);
not NOT1 (N6062, N6053);
and AND2 (N6063, N6055, N614);
or OR4 (N6064, N6061, N1401, N4394, N3150);
nor NOR2 (N6065, N6038, N2167);
nand NAND2 (N6066, N6064, N3301);
xor XOR2 (N6067, N6062, N3828);
nand NAND3 (N6068, N6054, N3144, N4243);
nor NOR3 (N6069, N6060, N3559, N3288);
buf BUF1 (N6070, N6056);
or OR4 (N6071, N6065, N5814, N1344, N6059);
and AND4 (N6072, N3119, N3745, N3598, N5944);
not NOT1 (N6073, N6050);
nor NOR2 (N6074, N6069, N1636);
and AND2 (N6075, N6063, N337);
and AND4 (N6076, N6072, N158, N1982, N4467);
and AND2 (N6077, N6066, N217);
not NOT1 (N6078, N6067);
and AND2 (N6079, N6052, N1465);
or OR2 (N6080, N6075, N1205);
or OR2 (N6081, N6076, N77);
xor XOR2 (N6082, N6078, N1342);
nand NAND2 (N6083, N6073, N4975);
buf BUF1 (N6084, N6079);
buf BUF1 (N6085, N6080);
not NOT1 (N6086, N6083);
nor NOR3 (N6087, N6070, N807, N5406);
not NOT1 (N6088, N6068);
and AND2 (N6089, N6088, N443);
or OR4 (N6090, N6077, N2798, N3430, N862);
or OR2 (N6091, N6074, N2238);
or OR4 (N6092, N6085, N4271, N65, N1296);
xor XOR2 (N6093, N6089, N4415);
xor XOR2 (N6094, N6081, N432);
not NOT1 (N6095, N6071);
or OR3 (N6096, N6093, N424, N5093);
or OR4 (N6097, N6094, N1077, N745, N5017);
not NOT1 (N6098, N6087);
not NOT1 (N6099, N6091);
nand NAND3 (N6100, N6090, N3709, N5967);
and AND3 (N6101, N6092, N2485, N1656);
and AND3 (N6102, N6097, N1521, N2705);
buf BUF1 (N6103, N6084);
buf BUF1 (N6104, N6103);
and AND4 (N6105, N6096, N5936, N930, N2567);
buf BUF1 (N6106, N6105);
nand NAND3 (N6107, N6095, N270, N726);
not NOT1 (N6108, N6098);
nand NAND3 (N6109, N6108, N3635, N1568);
nor NOR4 (N6110, N6106, N2330, N1109, N5159);
and AND3 (N6111, N6109, N3360, N3643);
and AND3 (N6112, N6082, N2534, N1699);
or OR2 (N6113, N6111, N5302);
nor NOR4 (N6114, N6113, N775, N413, N5094);
xor XOR2 (N6115, N6107, N4906);
nor NOR3 (N6116, N6086, N1634, N2605);
and AND2 (N6117, N6115, N4222);
and AND3 (N6118, N6110, N4531, N186);
nor NOR2 (N6119, N6112, N980);
or OR3 (N6120, N6116, N4819, N3717);
buf BUF1 (N6121, N6099);
nand NAND3 (N6122, N6101, N2626, N4204);
not NOT1 (N6123, N6119);
nor NOR2 (N6124, N6122, N3884);
nor NOR4 (N6125, N6104, N5924, N3053, N1763);
nand NAND3 (N6126, N6123, N4241, N2200);
not NOT1 (N6127, N6100);
xor XOR2 (N6128, N6124, N615);
buf BUF1 (N6129, N6120);
buf BUF1 (N6130, N6117);
and AND3 (N6131, N6114, N5216, N402);
nor NOR2 (N6132, N6128, N2325);
or OR2 (N6133, N6121, N4280);
and AND2 (N6134, N6129, N1152);
or OR4 (N6135, N6133, N5965, N4529, N4613);
not NOT1 (N6136, N6132);
and AND4 (N6137, N6125, N4572, N5342, N5336);
not NOT1 (N6138, N6102);
buf BUF1 (N6139, N6134);
nor NOR4 (N6140, N6138, N1792, N1105, N4238);
not NOT1 (N6141, N6130);
not NOT1 (N6142, N6141);
or OR3 (N6143, N6137, N861, N4379);
buf BUF1 (N6144, N6136);
and AND3 (N6145, N6118, N3384, N329);
and AND4 (N6146, N6139, N3949, N4688, N3044);
or OR4 (N6147, N6144, N245, N4739, N2022);
and AND3 (N6148, N6127, N5638, N3306);
not NOT1 (N6149, N6147);
nor NOR4 (N6150, N6131, N3754, N4859, N1783);
xor XOR2 (N6151, N6126, N2932);
xor XOR2 (N6152, N6142, N6117);
nor NOR3 (N6153, N6146, N2176, N2095);
buf BUF1 (N6154, N6149);
or OR3 (N6155, N6154, N3309, N1971);
buf BUF1 (N6156, N6153);
xor XOR2 (N6157, N6155, N1404);
and AND3 (N6158, N6151, N4826, N4832);
nand NAND3 (N6159, N6148, N4656, N4119);
buf BUF1 (N6160, N6140);
xor XOR2 (N6161, N6160, N5628);
xor XOR2 (N6162, N6161, N3912);
or OR3 (N6163, N6158, N2503, N4899);
or OR2 (N6164, N6159, N4890);
not NOT1 (N6165, N6143);
xor XOR2 (N6166, N6164, N1341);
not NOT1 (N6167, N6152);
not NOT1 (N6168, N6145);
buf BUF1 (N6169, N6157);
xor XOR2 (N6170, N6165, N1334);
xor XOR2 (N6171, N6169, N4050);
nand NAND2 (N6172, N6166, N2951);
not NOT1 (N6173, N6168);
xor XOR2 (N6174, N6173, N2204);
nand NAND4 (N6175, N6163, N3559, N4549, N5171);
or OR4 (N6176, N6171, N498, N807, N4604);
buf BUF1 (N6177, N6167);
and AND4 (N6178, N6156, N618, N628, N5998);
buf BUF1 (N6179, N6176);
or OR4 (N6180, N6162, N3555, N2687, N4513);
or OR4 (N6181, N6178, N1025, N4006, N5519);
xor XOR2 (N6182, N6150, N5129);
buf BUF1 (N6183, N6174);
nand NAND4 (N6184, N6170, N5578, N5482, N4194);
nand NAND2 (N6185, N6180, N4585);
nor NOR3 (N6186, N6182, N1077, N2943);
buf BUF1 (N6187, N6172);
and AND3 (N6188, N6185, N2661, N2972);
and AND4 (N6189, N6187, N233, N304, N4825);
not NOT1 (N6190, N6183);
buf BUF1 (N6191, N6135);
and AND4 (N6192, N6181, N2049, N4849, N4179);
not NOT1 (N6193, N6184);
nor NOR2 (N6194, N6191, N917);
nor NOR2 (N6195, N6194, N2689);
nor NOR4 (N6196, N6192, N1935, N2061, N32);
xor XOR2 (N6197, N6190, N2746);
or OR4 (N6198, N6196, N2399, N1204, N2174);
or OR2 (N6199, N6189, N4275);
buf BUF1 (N6200, N6186);
xor XOR2 (N6201, N6193, N2890);
nor NOR3 (N6202, N6195, N1176, N4156);
and AND2 (N6203, N6200, N1097);
not NOT1 (N6204, N6188);
buf BUF1 (N6205, N6203);
not NOT1 (N6206, N6197);
nand NAND3 (N6207, N6206, N1390, N1982);
and AND2 (N6208, N6204, N4842);
not NOT1 (N6209, N6205);
nand NAND3 (N6210, N6199, N2808, N2037);
nor NOR2 (N6211, N6202, N5668);
buf BUF1 (N6212, N6201);
or OR2 (N6213, N6211, N4374);
nor NOR4 (N6214, N6177, N1974, N1899, N4134);
xor XOR2 (N6215, N6210, N203);
buf BUF1 (N6216, N6198);
and AND2 (N6217, N6175, N4933);
nor NOR2 (N6218, N6217, N530);
or OR3 (N6219, N6215, N6094, N520);
or OR3 (N6220, N6212, N3413, N2575);
and AND3 (N6221, N6207, N2337, N2629);
and AND2 (N6222, N6214, N3244);
nor NOR2 (N6223, N6218, N2150);
buf BUF1 (N6224, N6221);
buf BUF1 (N6225, N6220);
nand NAND2 (N6226, N6223, N4840);
not NOT1 (N6227, N6219);
or OR2 (N6228, N6216, N2144);
xor XOR2 (N6229, N6228, N3826);
not NOT1 (N6230, N6213);
not NOT1 (N6231, N6209);
not NOT1 (N6232, N6222);
nand NAND4 (N6233, N6208, N6025, N2266, N878);
nor NOR4 (N6234, N6226, N2091, N2336, N4013);
nand NAND3 (N6235, N6232, N1990, N784);
buf BUF1 (N6236, N6224);
buf BUF1 (N6237, N6229);
nor NOR3 (N6238, N6237, N4936, N3144);
buf BUF1 (N6239, N6238);
or OR2 (N6240, N6239, N2369);
nand NAND2 (N6241, N6240, N2293);
nand NAND3 (N6242, N6227, N2328, N6049);
nand NAND2 (N6243, N6233, N1888);
not NOT1 (N6244, N6242);
xor XOR2 (N6245, N6234, N4555);
not NOT1 (N6246, N6179);
nor NOR4 (N6247, N6243, N2072, N3191, N1510);
and AND4 (N6248, N6230, N5975, N2509, N5492);
buf BUF1 (N6249, N6241);
and AND2 (N6250, N6231, N598);
nor NOR3 (N6251, N6249, N4456, N2334);
or OR4 (N6252, N6235, N491, N5695, N4680);
or OR2 (N6253, N6252, N130);
nand NAND4 (N6254, N6236, N3669, N5966, N1759);
buf BUF1 (N6255, N6225);
nand NAND4 (N6256, N6247, N1658, N5747, N4110);
not NOT1 (N6257, N6253);
xor XOR2 (N6258, N6251, N2023);
nand NAND3 (N6259, N6258, N5424, N6016);
nand NAND2 (N6260, N6245, N3154);
nor NOR4 (N6261, N6260, N31, N3325, N3955);
not NOT1 (N6262, N6255);
or OR4 (N6263, N6250, N4388, N1751, N2180);
nand NAND3 (N6264, N6261, N3114, N4018);
not NOT1 (N6265, N6259);
nor NOR2 (N6266, N6248, N6128);
and AND2 (N6267, N6262, N4580);
nand NAND2 (N6268, N6263, N4132);
and AND2 (N6269, N6265, N378);
nand NAND4 (N6270, N6264, N291, N6223, N1778);
xor XOR2 (N6271, N6244, N4653);
buf BUF1 (N6272, N6270);
or OR4 (N6273, N6268, N3813, N2906, N1899);
nand NAND3 (N6274, N6267, N886, N3005);
not NOT1 (N6275, N6246);
nor NOR2 (N6276, N6256, N6263);
not NOT1 (N6277, N6274);
nand NAND3 (N6278, N6272, N1372, N3974);
and AND2 (N6279, N6276, N1540);
not NOT1 (N6280, N6266);
or OR4 (N6281, N6273, N2947, N5207, N2867);
nor NOR3 (N6282, N6277, N2815, N2285);
buf BUF1 (N6283, N6278);
xor XOR2 (N6284, N6281, N5792);
buf BUF1 (N6285, N6275);
not NOT1 (N6286, N6284);
buf BUF1 (N6287, N6282);
xor XOR2 (N6288, N6283, N5566);
buf BUF1 (N6289, N6288);
nand NAND2 (N6290, N6269, N2486);
or OR2 (N6291, N6280, N5906);
not NOT1 (N6292, N6257);
nor NOR2 (N6293, N6292, N3895);
not NOT1 (N6294, N6287);
buf BUF1 (N6295, N6294);
nand NAND3 (N6296, N6289, N55, N981);
xor XOR2 (N6297, N6290, N5914);
buf BUF1 (N6298, N6296);
and AND4 (N6299, N6254, N20, N6156, N3466);
not NOT1 (N6300, N6279);
and AND2 (N6301, N6298, N5334);
or OR4 (N6302, N6295, N2899, N1364, N5476);
nand NAND3 (N6303, N6299, N3307, N4775);
nor NOR2 (N6304, N6297, N4490);
and AND3 (N6305, N6302, N1279, N4885);
not NOT1 (N6306, N6286);
and AND4 (N6307, N6303, N1551, N60, N2616);
nand NAND2 (N6308, N6300, N1391);
not NOT1 (N6309, N6271);
buf BUF1 (N6310, N6305);
and AND3 (N6311, N6307, N3031, N2860);
xor XOR2 (N6312, N6309, N364);
xor XOR2 (N6313, N6310, N4344);
and AND2 (N6314, N6304, N4191);
buf BUF1 (N6315, N6312);
nand NAND4 (N6316, N6313, N5126, N3406, N5365);
not NOT1 (N6317, N6291);
not NOT1 (N6318, N6315);
buf BUF1 (N6319, N6316);
nand NAND4 (N6320, N6285, N6039, N3502, N4344);
buf BUF1 (N6321, N6314);
xor XOR2 (N6322, N6321, N5393);
nand NAND2 (N6323, N6301, N1012);
not NOT1 (N6324, N6319);
xor XOR2 (N6325, N6293, N933);
or OR2 (N6326, N6311, N2124);
and AND4 (N6327, N6318, N1056, N4121, N5886);
not NOT1 (N6328, N6320);
nand NAND3 (N6329, N6326, N3221, N1170);
not NOT1 (N6330, N6322);
nor NOR3 (N6331, N6330, N6135, N4544);
or OR2 (N6332, N6306, N3346);
nor NOR2 (N6333, N6331, N834);
and AND2 (N6334, N6324, N2258);
and AND4 (N6335, N6333, N907, N2561, N4085);
nand NAND4 (N6336, N6327, N4693, N1285, N1957);
xor XOR2 (N6337, N6335, N5688);
not NOT1 (N6338, N6334);
nor NOR4 (N6339, N6332, N3460, N6306, N487);
buf BUF1 (N6340, N6325);
or OR2 (N6341, N6323, N518);
nand NAND4 (N6342, N6336, N3333, N1980, N2189);
xor XOR2 (N6343, N6338, N5426);
not NOT1 (N6344, N6329);
nor NOR3 (N6345, N6317, N2014, N2693);
nor NOR4 (N6346, N6341, N5324, N870, N4115);
nor NOR4 (N6347, N6308, N2099, N1449, N4712);
nand NAND3 (N6348, N6346, N3959, N3397);
not NOT1 (N6349, N6340);
buf BUF1 (N6350, N6345);
and AND4 (N6351, N6328, N4338, N807, N5457);
buf BUF1 (N6352, N6350);
not NOT1 (N6353, N6343);
or OR4 (N6354, N6347, N4045, N862, N6033);
buf BUF1 (N6355, N6349);
not NOT1 (N6356, N6342);
nor NOR3 (N6357, N6356, N2495, N1300);
and AND4 (N6358, N6353, N1318, N5743, N4440);
not NOT1 (N6359, N6337);
nor NOR4 (N6360, N6352, N344, N1150, N5541);
not NOT1 (N6361, N6351);
nor NOR3 (N6362, N6359, N124, N2898);
not NOT1 (N6363, N6360);
and AND3 (N6364, N6357, N1094, N4444);
or OR3 (N6365, N6364, N5759, N5525);
nand NAND3 (N6366, N6365, N2201, N2166);
nand NAND2 (N6367, N6358, N2985);
xor XOR2 (N6368, N6363, N5509);
nor NOR2 (N6369, N6354, N3952);
or OR2 (N6370, N6362, N3958);
nand NAND2 (N6371, N6355, N5313);
nor NOR3 (N6372, N6344, N5544, N2769);
buf BUF1 (N6373, N6367);
buf BUF1 (N6374, N6373);
buf BUF1 (N6375, N6371);
buf BUF1 (N6376, N6374);
not NOT1 (N6377, N6339);
or OR3 (N6378, N6368, N5001, N5336);
not NOT1 (N6379, N6376);
and AND4 (N6380, N6378, N4421, N3563, N4493);
nand NAND3 (N6381, N6348, N3486, N5708);
or OR3 (N6382, N6369, N5481, N4176);
and AND3 (N6383, N6380, N4672, N2156);
nand NAND2 (N6384, N6381, N3845);
nor NOR2 (N6385, N6379, N1304);
and AND4 (N6386, N6384, N1907, N5426, N2108);
nor NOR4 (N6387, N6386, N569, N2790, N4361);
nor NOR2 (N6388, N6383, N1598);
nand NAND4 (N6389, N6372, N5760, N3705, N3602);
and AND4 (N6390, N6387, N971, N5953, N1101);
or OR4 (N6391, N6390, N3103, N4630, N1916);
and AND4 (N6392, N6382, N411, N3498, N2096);
not NOT1 (N6393, N6389);
nand NAND2 (N6394, N6377, N4658);
nand NAND2 (N6395, N6391, N6225);
or OR4 (N6396, N6370, N3688, N5808, N4030);
or OR2 (N6397, N6393, N2443);
not NOT1 (N6398, N6392);
not NOT1 (N6399, N6388);
and AND4 (N6400, N6385, N2553, N5616, N880);
nand NAND3 (N6401, N6396, N1447, N4461);
or OR3 (N6402, N6400, N5745, N4880);
buf BUF1 (N6403, N6398);
buf BUF1 (N6404, N6401);
or OR2 (N6405, N6399, N619);
xor XOR2 (N6406, N6395, N271);
or OR2 (N6407, N6405, N1225);
nand NAND3 (N6408, N6375, N4087, N6119);
and AND2 (N6409, N6402, N3408);
xor XOR2 (N6410, N6409, N980);
nand NAND3 (N6411, N6403, N4511, N1112);
and AND4 (N6412, N6411, N4742, N4886, N4316);
nor NOR2 (N6413, N6407, N924);
and AND4 (N6414, N6410, N163, N2254, N5239);
not NOT1 (N6415, N6404);
or OR2 (N6416, N6361, N3393);
nand NAND4 (N6417, N6413, N2918, N911, N2510);
or OR3 (N6418, N6394, N1673, N3780);
or OR3 (N6419, N6416, N4965, N2454);
and AND4 (N6420, N6406, N4690, N3571, N715);
endmodule