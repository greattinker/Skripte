// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15;

output N297,N303,N314,N307,N313,N306,N312,N298,N311,N315;

or OR2 (N16, N15, N8);
and AND3 (N17, N12, N11, N8);
buf BUF1 (N18, N4);
not NOT1 (N19, N4);
buf BUF1 (N20, N5);
buf BUF1 (N21, N11);
buf BUF1 (N22, N13);
nand NAND2 (N23, N18, N17);
xor XOR2 (N24, N15, N7);
not NOT1 (N25, N23);
nand NAND4 (N26, N14, N9, N17, N4);
nand NAND3 (N27, N22, N22, N6);
buf BUF1 (N28, N12);
or OR3 (N29, N1, N24, N19);
xor XOR2 (N30, N20, N4);
or OR3 (N31, N7, N14, N18);
buf BUF1 (N32, N1);
or OR4 (N33, N31, N28, N31, N14);
not NOT1 (N34, N28);
xor XOR2 (N35, N21, N22);
nor NOR4 (N36, N35, N23, N7, N35);
xor XOR2 (N37, N26, N17);
xor XOR2 (N38, N33, N17);
or OR4 (N39, N36, N31, N37, N38);
xor XOR2 (N40, N2, N1);
xor XOR2 (N41, N13, N27);
buf BUF1 (N42, N5);
nor NOR2 (N43, N34, N13);
or OR2 (N44, N39, N37);
not NOT1 (N45, N44);
buf BUF1 (N46, N41);
buf BUF1 (N47, N25);
not NOT1 (N48, N32);
nor NOR3 (N49, N43, N41, N47);
xor XOR2 (N50, N1, N16);
xor XOR2 (N51, N17, N4);
nand NAND4 (N52, N30, N39, N18, N11);
buf BUF1 (N53, N46);
and AND4 (N54, N40, N25, N21, N53);
not NOT1 (N55, N48);
or OR4 (N56, N20, N34, N39, N12);
or OR3 (N57, N52, N22, N56);
xor XOR2 (N58, N57, N1);
and AND3 (N59, N41, N44, N53);
xor XOR2 (N60, N58, N56);
and AND4 (N61, N60, N29, N32, N54);
or OR3 (N62, N52, N13, N5);
or OR4 (N63, N22, N29, N8, N8);
buf BUF1 (N64, N45);
buf BUF1 (N65, N59);
or OR4 (N66, N62, N29, N36, N10);
and AND2 (N67, N55, N6);
or OR3 (N68, N65, N57, N15);
buf BUF1 (N69, N61);
or OR4 (N70, N66, N35, N29, N58);
and AND3 (N71, N68, N37, N66);
buf BUF1 (N72, N63);
xor XOR2 (N73, N70, N10);
buf BUF1 (N74, N69);
and AND3 (N75, N67, N32, N26);
xor XOR2 (N76, N51, N52);
or OR4 (N77, N72, N43, N5, N22);
not NOT1 (N78, N77);
nor NOR4 (N79, N75, N53, N74, N45);
nand NAND4 (N80, N37, N31, N8, N8);
and AND2 (N81, N42, N26);
or OR2 (N82, N71, N21);
xor XOR2 (N83, N80, N23);
xor XOR2 (N84, N78, N34);
buf BUF1 (N85, N82);
buf BUF1 (N86, N64);
and AND4 (N87, N49, N74, N15, N59);
or OR4 (N88, N79, N21, N30, N63);
nor NOR3 (N89, N85, N1, N41);
xor XOR2 (N90, N81, N41);
and AND3 (N91, N87, N80, N40);
buf BUF1 (N92, N84);
or OR4 (N93, N88, N29, N24, N69);
and AND4 (N94, N92, N66, N60, N26);
xor XOR2 (N95, N86, N92);
nand NAND4 (N96, N91, N84, N46, N73);
nor NOR2 (N97, N46, N20);
xor XOR2 (N98, N89, N91);
nor NOR2 (N99, N90, N74);
nor NOR2 (N100, N96, N31);
nand NAND4 (N101, N95, N31, N45, N95);
nand NAND2 (N102, N100, N66);
xor XOR2 (N103, N98, N28);
and AND2 (N104, N83, N83);
buf BUF1 (N105, N101);
not NOT1 (N106, N104);
or OR4 (N107, N103, N93, N101, N54);
or OR3 (N108, N66, N19, N80);
or OR4 (N109, N108, N14, N46, N87);
nor NOR2 (N110, N50, N44);
nand NAND3 (N111, N110, N94, N54);
and AND3 (N112, N21, N104, N10);
nor NOR4 (N113, N97, N18, N78, N87);
nor NOR3 (N114, N113, N45, N84);
or OR2 (N115, N102, N87);
and AND4 (N116, N106, N111, N20, N75);
nand NAND3 (N117, N86, N91, N109);
not NOT1 (N118, N48);
nand NAND4 (N119, N114, N18, N59, N108);
and AND2 (N120, N117, N101);
nand NAND4 (N121, N107, N23, N51, N71);
and AND4 (N122, N121, N80, N13, N101);
nand NAND4 (N123, N120, N51, N82, N44);
buf BUF1 (N124, N118);
buf BUF1 (N125, N112);
or OR4 (N126, N122, N9, N120, N96);
xor XOR2 (N127, N76, N105);
xor XOR2 (N128, N8, N74);
buf BUF1 (N129, N125);
or OR2 (N130, N126, N115);
buf BUF1 (N131, N106);
or OR2 (N132, N129, N72);
nand NAND2 (N133, N130, N117);
not NOT1 (N134, N99);
and AND3 (N135, N132, N58, N68);
and AND3 (N136, N123, N54, N37);
xor XOR2 (N137, N134, N84);
buf BUF1 (N138, N131);
or OR3 (N139, N116, N105, N12);
xor XOR2 (N140, N133, N117);
not NOT1 (N141, N140);
or OR4 (N142, N141, N15, N94, N129);
and AND4 (N143, N128, N99, N25, N106);
buf BUF1 (N144, N136);
and AND2 (N145, N119, N59);
buf BUF1 (N146, N144);
xor XOR2 (N147, N124, N73);
nand NAND4 (N148, N147, N135, N52, N6);
xor XOR2 (N149, N14, N64);
nor NOR3 (N150, N148, N41, N16);
not NOT1 (N151, N143);
nand NAND4 (N152, N146, N89, N145, N63);
or OR4 (N153, N91, N99, N9, N111);
buf BUF1 (N154, N150);
nor NOR3 (N155, N151, N145, N108);
or OR4 (N156, N139, N61, N138, N90);
nor NOR4 (N157, N148, N69, N44, N51);
xor XOR2 (N158, N137, N54);
buf BUF1 (N159, N153);
buf BUF1 (N160, N156);
xor XOR2 (N161, N160, N18);
and AND4 (N162, N154, N77, N34, N92);
and AND3 (N163, N158, N108, N25);
and AND2 (N164, N162, N122);
nand NAND4 (N165, N157, N12, N163, N70);
xor XOR2 (N166, N14, N145);
buf BUF1 (N167, N149);
nand NAND2 (N168, N165, N34);
or OR4 (N169, N167, N48, N106, N50);
xor XOR2 (N170, N168, N101);
nand NAND4 (N171, N166, N22, N43, N88);
or OR3 (N172, N170, N58, N28);
and AND2 (N173, N152, N125);
and AND3 (N174, N161, N123, N11);
and AND2 (N175, N169, N72);
not NOT1 (N176, N174);
not NOT1 (N177, N173);
nor NOR2 (N178, N142, N72);
xor XOR2 (N179, N127, N167);
xor XOR2 (N180, N164, N85);
buf BUF1 (N181, N179);
not NOT1 (N182, N172);
nor NOR4 (N183, N178, N94, N132, N10);
or OR3 (N184, N155, N171, N84);
or OR3 (N185, N157, N34, N33);
and AND4 (N186, N181, N173, N148, N74);
buf BUF1 (N187, N177);
or OR3 (N188, N184, N93, N30);
or OR4 (N189, N176, N184, N104, N38);
not NOT1 (N190, N186);
buf BUF1 (N191, N187);
buf BUF1 (N192, N188);
xor XOR2 (N193, N180, N91);
and AND2 (N194, N183, N68);
not NOT1 (N195, N182);
and AND4 (N196, N159, N174, N171, N30);
buf BUF1 (N197, N195);
buf BUF1 (N198, N197);
buf BUF1 (N199, N175);
and AND2 (N200, N196, N175);
xor XOR2 (N201, N192, N39);
not NOT1 (N202, N199);
xor XOR2 (N203, N185, N164);
or OR3 (N204, N194, N37, N78);
not NOT1 (N205, N201);
nand NAND2 (N206, N205, N109);
buf BUF1 (N207, N204);
or OR2 (N208, N203, N64);
not NOT1 (N209, N206);
not NOT1 (N210, N193);
nand NAND2 (N211, N190, N204);
not NOT1 (N212, N202);
buf BUF1 (N213, N189);
xor XOR2 (N214, N208, N40);
xor XOR2 (N215, N200, N161);
not NOT1 (N216, N210);
not NOT1 (N217, N191);
nor NOR3 (N218, N215, N1, N89);
xor XOR2 (N219, N217, N105);
and AND3 (N220, N211, N168, N78);
buf BUF1 (N221, N209);
nor NOR4 (N222, N213, N99, N101, N17);
nor NOR3 (N223, N218, N28, N171);
xor XOR2 (N224, N222, N1);
xor XOR2 (N225, N223, N27);
xor XOR2 (N226, N216, N93);
nand NAND3 (N227, N225, N144, N25);
not NOT1 (N228, N220);
not NOT1 (N229, N224);
buf BUF1 (N230, N226);
xor XOR2 (N231, N227, N165);
and AND4 (N232, N212, N187, N177, N24);
nor NOR3 (N233, N198, N154, N148);
nor NOR2 (N234, N232, N89);
not NOT1 (N235, N230);
not NOT1 (N236, N207);
xor XOR2 (N237, N236, N171);
nor NOR2 (N238, N233, N20);
and AND3 (N239, N214, N47, N40);
and AND2 (N240, N229, N117);
or OR4 (N241, N238, N191, N158, N107);
nor NOR3 (N242, N231, N148, N89);
xor XOR2 (N243, N240, N237);
nand NAND3 (N244, N35, N220, N216);
nand NAND2 (N245, N243, N61);
xor XOR2 (N246, N245, N132);
nor NOR4 (N247, N244, N7, N32, N150);
nor NOR3 (N248, N234, N61, N6);
or OR4 (N249, N228, N206, N58, N179);
xor XOR2 (N250, N219, N61);
xor XOR2 (N251, N242, N211);
and AND3 (N252, N235, N175, N153);
nor NOR4 (N253, N247, N86, N9, N86);
nor NOR4 (N254, N250, N40, N159, N94);
xor XOR2 (N255, N249, N210);
or OR3 (N256, N239, N61, N107);
and AND3 (N257, N221, N45, N171);
not NOT1 (N258, N254);
buf BUF1 (N259, N241);
nor NOR2 (N260, N256, N206);
not NOT1 (N261, N259);
xor XOR2 (N262, N258, N181);
and AND3 (N263, N260, N5, N128);
buf BUF1 (N264, N251);
buf BUF1 (N265, N262);
buf BUF1 (N266, N248);
not NOT1 (N267, N252);
buf BUF1 (N268, N265);
and AND2 (N269, N264, N164);
or OR2 (N270, N255, N115);
xor XOR2 (N271, N257, N75);
and AND2 (N272, N246, N23);
or OR3 (N273, N270, N42, N56);
nor NOR4 (N274, N266, N189, N235, N37);
buf BUF1 (N275, N263);
xor XOR2 (N276, N261, N40);
xor XOR2 (N277, N268, N34);
not NOT1 (N278, N274);
or OR2 (N279, N276, N191);
buf BUF1 (N280, N271);
xor XOR2 (N281, N280, N10);
not NOT1 (N282, N281);
or OR2 (N283, N279, N209);
not NOT1 (N284, N283);
not NOT1 (N285, N267);
nor NOR2 (N286, N285, N138);
not NOT1 (N287, N253);
nor NOR2 (N288, N269, N252);
or OR2 (N289, N286, N65);
nor NOR3 (N290, N275, N58, N120);
not NOT1 (N291, N289);
xor XOR2 (N292, N282, N112);
buf BUF1 (N293, N290);
buf BUF1 (N294, N292);
buf BUF1 (N295, N273);
nand NAND2 (N296, N293, N227);
not NOT1 (N297, N284);
xor XOR2 (N298, N272, N272);
or OR3 (N299, N294, N47, N100);
nand NAND2 (N300, N278, N274);
or OR2 (N301, N295, N152);
buf BUF1 (N302, N301);
nand NAND3 (N303, N302, N209, N184);
nor NOR4 (N304, N291, N41, N137, N217);
nor NOR3 (N305, N299, N20, N58);
not NOT1 (N306, N305);
buf BUF1 (N307, N288);
not NOT1 (N308, N287);
and AND2 (N309, N296, N116);
xor XOR2 (N310, N309, N205);
nand NAND2 (N311, N304, N7);
not NOT1 (N312, N300);
xor XOR2 (N313, N277, N93);
nor NOR4 (N314, N310, N161, N31, N267);
not NOT1 (N315, N308);
endmodule