// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24;

output N117,N95,N110,N121,N113,N105,N123,N114,N119,N124;

nand NAND2 (N25, N24, N16);
and AND2 (N26, N9, N15);
xor XOR2 (N27, N5, N17);
nand NAND2 (N28, N16, N9);
nand NAND3 (N29, N3, N22, N3);
buf BUF1 (N30, N17);
not NOT1 (N31, N6);
not NOT1 (N32, N8);
and AND4 (N33, N31, N17, N3, N15);
xor XOR2 (N34, N19, N28);
nand NAND2 (N35, N24, N31);
or OR3 (N36, N22, N31, N27);
or OR2 (N37, N18, N27);
nand NAND2 (N38, N34, N2);
and AND2 (N39, N37, N21);
and AND2 (N40, N35, N1);
or OR4 (N41, N33, N24, N15, N31);
or OR4 (N42, N32, N20, N17, N36);
not NOT1 (N43, N14);
not NOT1 (N44, N30);
nor NOR2 (N45, N38, N6);
nor NOR3 (N46, N43, N33, N45);
nand NAND3 (N47, N24, N38, N23);
not NOT1 (N48, N29);
nand NAND4 (N49, N41, N34, N5, N18);
not NOT1 (N50, N39);
or OR2 (N51, N50, N45);
or OR3 (N52, N25, N7, N15);
not NOT1 (N53, N52);
nor NOR3 (N54, N48, N17, N35);
xor XOR2 (N55, N51, N23);
nor NOR4 (N56, N47, N54, N41, N29);
or OR2 (N57, N9, N23);
or OR3 (N58, N55, N39, N24);
and AND3 (N59, N57, N23, N37);
nor NOR3 (N60, N26, N23, N51);
or OR3 (N61, N46, N19, N19);
not NOT1 (N62, N59);
nor NOR3 (N63, N60, N22, N21);
and AND2 (N64, N42, N16);
nand NAND4 (N65, N61, N44, N5, N18);
nor NOR4 (N66, N43, N31, N9, N48);
not NOT1 (N67, N56);
or OR2 (N68, N67, N39);
and AND2 (N69, N68, N23);
nor NOR2 (N70, N40, N21);
not NOT1 (N71, N49);
nor NOR2 (N72, N64, N70);
buf BUF1 (N73, N36);
nor NOR3 (N74, N62, N70, N6);
not NOT1 (N75, N63);
and AND2 (N76, N75, N75);
nand NAND4 (N77, N69, N4, N45, N40);
not NOT1 (N78, N65);
or OR4 (N79, N76, N43, N22, N15);
and AND2 (N80, N66, N6);
nand NAND4 (N81, N80, N79, N34, N19);
or OR3 (N82, N58, N39, N2);
and AND3 (N83, N63, N9, N62);
nand NAND3 (N84, N74, N75, N56);
buf BUF1 (N85, N73);
not NOT1 (N86, N71);
and AND4 (N87, N84, N41, N34, N19);
xor XOR2 (N88, N72, N83);
buf BUF1 (N89, N10);
nand NAND4 (N90, N86, N11, N60, N78);
xor XOR2 (N91, N9, N35);
xor XOR2 (N92, N82, N85);
nor NOR2 (N93, N46, N82);
nor NOR3 (N94, N93, N89, N67);
and AND2 (N95, N62, N83);
and AND2 (N96, N91, N35);
not NOT1 (N97, N88);
nand NAND3 (N98, N97, N46, N79);
buf BUF1 (N99, N92);
and AND2 (N100, N81, N15);
or OR2 (N101, N53, N19);
nor NOR2 (N102, N96, N78);
xor XOR2 (N103, N101, N99);
xor XOR2 (N104, N58, N93);
not NOT1 (N105, N98);
xor XOR2 (N106, N104, N78);
not NOT1 (N107, N106);
and AND2 (N108, N100, N11);
and AND2 (N109, N107, N77);
nor NOR3 (N110, N30, N92, N17);
nor NOR4 (N111, N90, N47, N70, N77);
buf BUF1 (N112, N102);
not NOT1 (N113, N87);
buf BUF1 (N114, N108);
or OR3 (N115, N109, N67, N11);
or OR4 (N116, N112, N111, N42, N53);
nor NOR4 (N117, N46, N97, N116, N63);
nor NOR2 (N118, N99, N54);
not NOT1 (N119, N94);
or OR2 (N120, N103, N61);
or OR3 (N121, N115, N43, N97);
nand NAND2 (N122, N120, N64);
xor XOR2 (N123, N118, N51);
and AND3 (N124, N122, N29, N47);
endmodule