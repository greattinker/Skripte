// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12;

output N501,N511,N503,N490,N509,N510,N496,N508,N495,N512;

nor NOR3 (N13, N8, N7, N11);
xor XOR2 (N14, N12, N9);
xor XOR2 (N15, N6, N5);
xor XOR2 (N16, N14, N6);
nor NOR4 (N17, N15, N2, N14, N4);
or OR2 (N18, N11, N7);
buf BUF1 (N19, N7);
xor XOR2 (N20, N11, N6);
not NOT1 (N21, N8);
nand NAND4 (N22, N9, N6, N4, N16);
not NOT1 (N23, N5);
nand NAND3 (N24, N22, N6, N18);
not NOT1 (N25, N24);
buf BUF1 (N26, N1);
xor XOR2 (N27, N3, N26);
or OR4 (N28, N2, N4, N3, N15);
or OR3 (N29, N1, N28, N19);
and AND2 (N30, N12, N11);
nand NAND2 (N31, N3, N18);
xor XOR2 (N32, N31, N1);
and AND3 (N33, N30, N24, N27);
buf BUF1 (N34, N7);
nor NOR2 (N35, N23, N9);
not NOT1 (N36, N35);
not NOT1 (N37, N32);
not NOT1 (N38, N21);
and AND3 (N39, N29, N12, N31);
not NOT1 (N40, N25);
or OR3 (N41, N34, N26, N4);
not NOT1 (N42, N41);
nor NOR2 (N43, N37, N36);
buf BUF1 (N44, N26);
and AND3 (N45, N43, N6, N10);
nor NOR4 (N46, N13, N19, N12, N43);
or OR3 (N47, N20, N19, N19);
or OR4 (N48, N46, N8, N18, N23);
buf BUF1 (N49, N44);
or OR2 (N50, N40, N41);
and AND3 (N51, N48, N15, N41);
and AND2 (N52, N17, N39);
buf BUF1 (N53, N9);
buf BUF1 (N54, N47);
and AND3 (N55, N42, N38, N50);
or OR3 (N56, N24, N54, N4);
not NOT1 (N57, N33);
or OR3 (N58, N1, N42, N43);
not NOT1 (N59, N40);
buf BUF1 (N60, N53);
buf BUF1 (N61, N51);
and AND3 (N62, N56, N23, N3);
xor XOR2 (N63, N60, N40);
and AND4 (N64, N57, N27, N6, N60);
xor XOR2 (N65, N52, N16);
buf BUF1 (N66, N45);
buf BUF1 (N67, N61);
nand NAND4 (N68, N55, N59, N56, N65);
or OR3 (N69, N27, N25, N2);
or OR2 (N70, N27, N64);
and AND4 (N71, N10, N32, N50, N60);
and AND3 (N72, N71, N27, N63);
nor NOR4 (N73, N46, N15, N56, N31);
buf BUF1 (N74, N69);
not NOT1 (N75, N68);
buf BUF1 (N76, N62);
nand NAND2 (N77, N49, N34);
not NOT1 (N78, N75);
nand NAND3 (N79, N78, N55, N26);
buf BUF1 (N80, N67);
or OR2 (N81, N70, N38);
or OR4 (N82, N74, N59, N52, N45);
buf BUF1 (N83, N73);
nand NAND3 (N84, N77, N59, N46);
xor XOR2 (N85, N76, N63);
buf BUF1 (N86, N80);
or OR3 (N87, N58, N21, N6);
and AND3 (N88, N79, N79, N43);
nor NOR4 (N89, N82, N44, N54, N49);
buf BUF1 (N90, N85);
or OR3 (N91, N87, N60, N5);
or OR2 (N92, N88, N41);
and AND2 (N93, N92, N79);
xor XOR2 (N94, N72, N5);
or OR2 (N95, N90, N39);
xor XOR2 (N96, N89, N91);
not NOT1 (N97, N66);
buf BUF1 (N98, N69);
xor XOR2 (N99, N96, N11);
nor NOR2 (N100, N94, N15);
not NOT1 (N101, N100);
not NOT1 (N102, N98);
nor NOR4 (N103, N83, N67, N20, N42);
xor XOR2 (N104, N84, N90);
and AND3 (N105, N97, N72, N39);
buf BUF1 (N106, N99);
nand NAND3 (N107, N103, N99, N54);
buf BUF1 (N108, N86);
not NOT1 (N109, N106);
and AND3 (N110, N108, N59, N108);
nor NOR3 (N111, N101, N22, N53);
or OR2 (N112, N102, N12);
buf BUF1 (N113, N95);
buf BUF1 (N114, N113);
nand NAND2 (N115, N93, N25);
not NOT1 (N116, N105);
not NOT1 (N117, N111);
nand NAND3 (N118, N116, N46, N43);
buf BUF1 (N119, N104);
xor XOR2 (N120, N109, N34);
not NOT1 (N121, N81);
and AND3 (N122, N118, N114, N120);
or OR3 (N123, N58, N30, N108);
buf BUF1 (N124, N120);
nand NAND2 (N125, N122, N79);
nand NAND3 (N126, N121, N77, N69);
xor XOR2 (N127, N107, N29);
not NOT1 (N128, N115);
nor NOR2 (N129, N125, N13);
nor NOR4 (N130, N129, N122, N2, N16);
or OR2 (N131, N112, N86);
buf BUF1 (N132, N128);
nand NAND4 (N133, N132, N9, N23, N102);
xor XOR2 (N134, N123, N107);
xor XOR2 (N135, N130, N105);
xor XOR2 (N136, N134, N21);
xor XOR2 (N137, N136, N73);
not NOT1 (N138, N135);
and AND4 (N139, N117, N16, N122, N89);
not NOT1 (N140, N131);
not NOT1 (N141, N140);
buf BUF1 (N142, N110);
buf BUF1 (N143, N133);
nand NAND2 (N144, N119, N112);
buf BUF1 (N145, N127);
xor XOR2 (N146, N139, N35);
xor XOR2 (N147, N142, N101);
xor XOR2 (N148, N137, N35);
xor XOR2 (N149, N138, N114);
not NOT1 (N150, N147);
buf BUF1 (N151, N144);
nand NAND4 (N152, N145, N78, N125, N73);
not NOT1 (N153, N152);
nor NOR4 (N154, N151, N113, N45, N30);
not NOT1 (N155, N143);
and AND4 (N156, N153, N70, N61, N137);
xor XOR2 (N157, N149, N55);
xor XOR2 (N158, N150, N125);
nor NOR2 (N159, N156, N54);
xor XOR2 (N160, N148, N114);
nor NOR4 (N161, N155, N159, N64, N81);
buf BUF1 (N162, N155);
nor NOR2 (N163, N162, N60);
buf BUF1 (N164, N141);
nor NOR2 (N165, N146, N18);
nand NAND2 (N166, N124, N20);
and AND2 (N167, N160, N124);
nor NOR4 (N168, N166, N113, N27, N66);
or OR3 (N169, N163, N168, N131);
or OR3 (N170, N110, N74, N11);
xor XOR2 (N171, N126, N29);
or OR2 (N172, N158, N61);
nand NAND3 (N173, N167, N30, N21);
and AND4 (N174, N154, N113, N135, N151);
not NOT1 (N175, N164);
buf BUF1 (N176, N171);
not NOT1 (N177, N176);
not NOT1 (N178, N165);
buf BUF1 (N179, N172);
nor NOR4 (N180, N170, N80, N14, N77);
buf BUF1 (N181, N157);
nor NOR2 (N182, N173, N66);
nand NAND4 (N183, N179, N90, N53, N76);
xor XOR2 (N184, N181, N28);
or OR4 (N185, N184, N74, N8, N54);
not NOT1 (N186, N177);
not NOT1 (N187, N182);
buf BUF1 (N188, N174);
xor XOR2 (N189, N161, N40);
not NOT1 (N190, N186);
not NOT1 (N191, N189);
nand NAND3 (N192, N169, N146, N14);
buf BUF1 (N193, N180);
xor XOR2 (N194, N193, N163);
buf BUF1 (N195, N187);
and AND3 (N196, N178, N33, N167);
xor XOR2 (N197, N195, N107);
nor NOR2 (N198, N190, N147);
or OR4 (N199, N192, N168, N103, N91);
xor XOR2 (N200, N194, N123);
nand NAND3 (N201, N191, N171, N154);
buf BUF1 (N202, N199);
and AND3 (N203, N200, N100, N47);
not NOT1 (N204, N201);
and AND2 (N205, N203, N90);
and AND2 (N206, N198, N34);
nor NOR3 (N207, N205, N176, N83);
nand NAND4 (N208, N188, N134, N66, N42);
not NOT1 (N209, N183);
buf BUF1 (N210, N206);
xor XOR2 (N211, N197, N121);
nor NOR2 (N212, N196, N133);
nor NOR4 (N213, N204, N43, N139, N177);
nor NOR4 (N214, N202, N151, N92, N191);
buf BUF1 (N215, N211);
nor NOR2 (N216, N213, N72);
nor NOR2 (N217, N208, N166);
nand NAND4 (N218, N209, N89, N32, N167);
nand NAND4 (N219, N218, N161, N179, N179);
nand NAND3 (N220, N219, N129, N217);
xor XOR2 (N221, N94, N22);
nor NOR4 (N222, N215, N167, N74, N166);
nand NAND2 (N223, N207, N68);
xor XOR2 (N224, N220, N147);
nor NOR4 (N225, N185, N221, N100, N174);
nor NOR4 (N226, N165, N26, N140, N200);
buf BUF1 (N227, N216);
buf BUF1 (N228, N212);
nor NOR2 (N229, N228, N127);
buf BUF1 (N230, N226);
nand NAND4 (N231, N227, N62, N87, N118);
not NOT1 (N232, N230);
and AND4 (N233, N214, N52, N197, N116);
nand NAND2 (N234, N224, N111);
or OR2 (N235, N234, N46);
buf BUF1 (N236, N229);
not NOT1 (N237, N210);
and AND3 (N238, N222, N152, N30);
nor NOR4 (N239, N232, N235, N126, N67);
buf BUF1 (N240, N198);
and AND4 (N241, N236, N39, N59, N237);
and AND3 (N242, N73, N194, N44);
nor NOR2 (N243, N239, N51);
and AND2 (N244, N231, N140);
buf BUF1 (N245, N223);
and AND2 (N246, N245, N119);
xor XOR2 (N247, N225, N103);
not NOT1 (N248, N241);
buf BUF1 (N249, N244);
or OR3 (N250, N233, N138, N37);
not NOT1 (N251, N248);
xor XOR2 (N252, N251, N135);
or OR3 (N253, N175, N96, N120);
nor NOR4 (N254, N250, N247, N62, N2);
not NOT1 (N255, N141);
nor NOR3 (N256, N246, N254, N79);
nor NOR3 (N257, N175, N218, N72);
nand NAND3 (N258, N255, N158, N190);
and AND4 (N259, N252, N182, N167, N116);
and AND4 (N260, N242, N161, N56, N117);
nand NAND3 (N261, N259, N186, N117);
not NOT1 (N262, N253);
nor NOR2 (N263, N262, N196);
not NOT1 (N264, N243);
xor XOR2 (N265, N260, N46);
buf BUF1 (N266, N258);
and AND4 (N267, N263, N18, N207, N53);
and AND4 (N268, N256, N111, N252, N61);
xor XOR2 (N269, N240, N239);
not NOT1 (N270, N261);
and AND2 (N271, N269, N207);
buf BUF1 (N272, N268);
not NOT1 (N273, N257);
buf BUF1 (N274, N249);
and AND2 (N275, N264, N2);
buf BUF1 (N276, N266);
nor NOR2 (N277, N273, N150);
nand NAND2 (N278, N277, N36);
nor NOR4 (N279, N238, N189, N74, N227);
or OR4 (N280, N278, N147, N242, N150);
nand NAND3 (N281, N274, N84, N172);
nor NOR3 (N282, N275, N39, N223);
buf BUF1 (N283, N271);
xor XOR2 (N284, N282, N23);
nor NOR2 (N285, N279, N137);
xor XOR2 (N286, N267, N142);
xor XOR2 (N287, N285, N39);
not NOT1 (N288, N284);
not NOT1 (N289, N288);
nor NOR3 (N290, N281, N73, N252);
buf BUF1 (N291, N289);
xor XOR2 (N292, N290, N274);
nand NAND2 (N293, N283, N257);
or OR2 (N294, N286, N237);
buf BUF1 (N295, N280);
and AND2 (N296, N295, N280);
buf BUF1 (N297, N265);
and AND4 (N298, N287, N212, N78, N247);
or OR4 (N299, N294, N169, N219, N154);
and AND4 (N300, N293, N229, N298, N15);
and AND4 (N301, N10, N290, N230, N117);
xor XOR2 (N302, N291, N1);
not NOT1 (N303, N301);
or OR2 (N304, N296, N26);
or OR4 (N305, N270, N208, N288, N151);
or OR3 (N306, N299, N9, N198);
nor NOR2 (N307, N302, N211);
nor NOR4 (N308, N297, N155, N257, N242);
not NOT1 (N309, N292);
and AND4 (N310, N305, N241, N177, N222);
buf BUF1 (N311, N306);
and AND4 (N312, N276, N139, N28, N209);
xor XOR2 (N313, N308, N219);
or OR3 (N314, N311, N227, N294);
and AND2 (N315, N313, N104);
xor XOR2 (N316, N314, N202);
xor XOR2 (N317, N303, N109);
nor NOR3 (N318, N309, N10, N282);
buf BUF1 (N319, N312);
or OR3 (N320, N316, N239, N46);
or OR4 (N321, N307, N82, N76, N37);
not NOT1 (N322, N320);
and AND4 (N323, N322, N290, N139, N298);
and AND3 (N324, N310, N185, N30);
buf BUF1 (N325, N318);
not NOT1 (N326, N321);
nand NAND4 (N327, N300, N14, N117, N53);
not NOT1 (N328, N326);
nor NOR2 (N329, N323, N252);
buf BUF1 (N330, N315);
nand NAND3 (N331, N324, N308, N117);
not NOT1 (N332, N317);
buf BUF1 (N333, N319);
buf BUF1 (N334, N330);
nor NOR3 (N335, N334, N225, N17);
nor NOR4 (N336, N272, N232, N215, N263);
not NOT1 (N337, N327);
nor NOR3 (N338, N329, N118, N199);
nor NOR4 (N339, N338, N313, N76, N232);
buf BUF1 (N340, N331);
xor XOR2 (N341, N339, N321);
and AND4 (N342, N332, N166, N185, N301);
buf BUF1 (N343, N328);
nand NAND3 (N344, N335, N332, N155);
nand NAND3 (N345, N325, N107, N106);
xor XOR2 (N346, N340, N139);
nor NOR3 (N347, N336, N86, N288);
and AND2 (N348, N342, N256);
not NOT1 (N349, N333);
not NOT1 (N350, N341);
xor XOR2 (N351, N304, N236);
nor NOR3 (N352, N343, N229, N328);
buf BUF1 (N353, N347);
not NOT1 (N354, N350);
not NOT1 (N355, N352);
not NOT1 (N356, N337);
not NOT1 (N357, N348);
or OR3 (N358, N346, N9, N236);
nand NAND2 (N359, N354, N79);
nand NAND2 (N360, N351, N170);
or OR3 (N361, N349, N241, N301);
not NOT1 (N362, N355);
and AND3 (N363, N359, N29, N190);
or OR3 (N364, N353, N225, N62);
or OR3 (N365, N358, N185, N217);
buf BUF1 (N366, N356);
nor NOR3 (N367, N363, N129, N320);
or OR3 (N368, N361, N130, N278);
buf BUF1 (N369, N357);
nor NOR3 (N370, N369, N298, N207);
and AND2 (N371, N366, N305);
nand NAND2 (N372, N365, N41);
or OR3 (N373, N367, N294, N42);
and AND3 (N374, N360, N238, N273);
and AND4 (N375, N370, N136, N130, N107);
nand NAND3 (N376, N374, N46, N223);
or OR4 (N377, N376, N233, N333, N90);
nor NOR2 (N378, N364, N139);
xor XOR2 (N379, N377, N193);
nor NOR4 (N380, N373, N19, N127, N88);
xor XOR2 (N381, N362, N337);
nor NOR2 (N382, N372, N80);
or OR2 (N383, N381, N244);
or OR4 (N384, N383, N140, N140, N36);
and AND4 (N385, N379, N35, N307, N51);
nor NOR2 (N386, N384, N159);
or OR3 (N387, N368, N1, N210);
xor XOR2 (N388, N375, N221);
and AND3 (N389, N345, N284, N93);
or OR3 (N390, N371, N97, N34);
not NOT1 (N391, N387);
or OR4 (N392, N390, N226, N265, N37);
and AND4 (N393, N382, N269, N237, N17);
buf BUF1 (N394, N380);
and AND2 (N395, N378, N203);
and AND2 (N396, N389, N240);
nand NAND2 (N397, N386, N33);
not NOT1 (N398, N395);
nand NAND4 (N399, N388, N1, N131, N79);
nand NAND3 (N400, N344, N321, N357);
buf BUF1 (N401, N396);
buf BUF1 (N402, N401);
xor XOR2 (N403, N392, N293);
buf BUF1 (N404, N400);
not NOT1 (N405, N385);
xor XOR2 (N406, N394, N312);
nand NAND3 (N407, N405, N112, N167);
and AND4 (N408, N406, N218, N179, N304);
nand NAND4 (N409, N407, N146, N321, N83);
or OR2 (N410, N391, N221);
xor XOR2 (N411, N393, N293);
buf BUF1 (N412, N411);
nor NOR4 (N413, N402, N36, N69, N118);
nand NAND4 (N414, N412, N39, N356, N360);
and AND3 (N415, N399, N379, N141);
not NOT1 (N416, N403);
nor NOR3 (N417, N413, N78, N221);
xor XOR2 (N418, N416, N214);
xor XOR2 (N419, N398, N206);
nor NOR2 (N420, N415, N231);
xor XOR2 (N421, N417, N244);
nand NAND3 (N422, N414, N37, N25);
and AND3 (N423, N421, N248, N44);
nand NAND2 (N424, N420, N18);
nand NAND4 (N425, N419, N338, N213, N128);
not NOT1 (N426, N425);
buf BUF1 (N427, N418);
xor XOR2 (N428, N404, N94);
nor NOR2 (N429, N408, N300);
xor XOR2 (N430, N426, N353);
xor XOR2 (N431, N427, N61);
or OR2 (N432, N397, N408);
xor XOR2 (N433, N423, N186);
or OR2 (N434, N410, N333);
buf BUF1 (N435, N428);
and AND2 (N436, N435, N360);
nor NOR4 (N437, N432, N63, N38, N344);
buf BUF1 (N438, N430);
xor XOR2 (N439, N437, N270);
nor NOR3 (N440, N422, N378, N129);
or OR4 (N441, N433, N400, N53, N152);
nand NAND3 (N442, N431, N44, N189);
nand NAND3 (N443, N441, N110, N41);
not NOT1 (N444, N439);
nor NOR3 (N445, N429, N281, N388);
buf BUF1 (N446, N443);
nand NAND4 (N447, N409, N434, N141, N79);
not NOT1 (N448, N87);
buf BUF1 (N449, N446);
nand NAND4 (N450, N447, N13, N360, N246);
or OR3 (N451, N438, N304, N117);
nor NOR4 (N452, N449, N56, N27, N327);
nor NOR3 (N453, N440, N286, N309);
nand NAND2 (N454, N450, N65);
and AND4 (N455, N448, N329, N7, N106);
or OR3 (N456, N455, N360, N17);
xor XOR2 (N457, N452, N169);
nor NOR2 (N458, N456, N371);
and AND3 (N459, N454, N112, N284);
buf BUF1 (N460, N457);
xor XOR2 (N461, N444, N85);
xor XOR2 (N462, N424, N119);
or OR4 (N463, N453, N341, N63, N327);
nand NAND2 (N464, N436, N261);
and AND3 (N465, N464, N201, N161);
nor NOR4 (N466, N459, N72, N241, N376);
buf BUF1 (N467, N461);
xor XOR2 (N468, N445, N309);
nor NOR3 (N469, N468, N414, N121);
buf BUF1 (N470, N467);
or OR3 (N471, N463, N340, N346);
nor NOR3 (N472, N469, N178, N332);
and AND3 (N473, N462, N227, N318);
nor NOR4 (N474, N470, N386, N281, N236);
buf BUF1 (N475, N442);
nand NAND4 (N476, N475, N301, N410, N180);
buf BUF1 (N477, N476);
not NOT1 (N478, N472);
and AND2 (N479, N458, N230);
not NOT1 (N480, N466);
xor XOR2 (N481, N465, N26);
xor XOR2 (N482, N479, N395);
nor NOR4 (N483, N480, N319, N68, N66);
nand NAND3 (N484, N478, N29, N398);
nand NAND2 (N485, N482, N412);
buf BUF1 (N486, N471);
or OR3 (N487, N486, N232, N471);
xor XOR2 (N488, N487, N133);
nor NOR2 (N489, N473, N52);
not NOT1 (N490, N451);
or OR4 (N491, N483, N264, N354, N172);
and AND2 (N492, N474, N86);
and AND2 (N493, N484, N251);
nand NAND4 (N494, N492, N402, N428, N241);
and AND2 (N495, N488, N69);
nor NOR3 (N496, N485, N446, N122);
nor NOR2 (N497, N460, N382);
nor NOR2 (N498, N477, N394);
or OR4 (N499, N494, N325, N398, N42);
buf BUF1 (N500, N499);
xor XOR2 (N501, N497, N134);
nor NOR4 (N502, N498, N284, N477, N356);
and AND4 (N503, N481, N15, N440, N358);
nor NOR3 (N504, N489, N187, N428);
or OR3 (N505, N500, N54, N157);
or OR2 (N506, N502, N309);
or OR2 (N507, N504, N287);
or OR4 (N508, N493, N420, N468, N358);
not NOT1 (N509, N506);
xor XOR2 (N510, N491, N294);
nor NOR2 (N511, N505, N24);
xor XOR2 (N512, N507, N376);
endmodule