// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19;

output N6418,N6416,N6414,N6410,N6411,N6412,N6403,N6415,N6413,N6419;

nor NOR2 (N20, N17, N11);
not NOT1 (N21, N17);
nor NOR4 (N22, N2, N3, N13, N9);
nor NOR3 (N23, N12, N17, N14);
xor XOR2 (N24, N3, N9);
not NOT1 (N25, N19);
xor XOR2 (N26, N6, N25);
buf BUF1 (N27, N1);
buf BUF1 (N28, N14);
nand NAND3 (N29, N3, N24, N26);
nand NAND3 (N30, N18, N13, N7);
or OR4 (N31, N9, N13, N13, N7);
buf BUF1 (N32, N29);
nor NOR2 (N33, N32, N3);
and AND2 (N34, N32, N30);
buf BUF1 (N35, N9);
or OR3 (N36, N22, N2, N10);
and AND2 (N37, N21, N3);
nor NOR4 (N38, N35, N12, N16, N25);
xor XOR2 (N39, N33, N18);
not NOT1 (N40, N37);
not NOT1 (N41, N23);
buf BUF1 (N42, N36);
nand NAND2 (N43, N20, N11);
xor XOR2 (N44, N31, N14);
nand NAND4 (N45, N27, N6, N7, N34);
or OR3 (N46, N6, N25, N1);
nor NOR3 (N47, N41, N32, N45);
nand NAND4 (N48, N16, N44, N9, N13);
nor NOR3 (N49, N36, N25, N44);
buf BUF1 (N50, N49);
and AND3 (N51, N47, N27, N8);
nand NAND3 (N52, N28, N42, N10);
nand NAND4 (N53, N29, N7, N40, N15);
or OR3 (N54, N46, N30, N13);
xor XOR2 (N55, N24, N27);
and AND2 (N56, N39, N10);
buf BUF1 (N57, N56);
nor NOR2 (N58, N50, N35);
buf BUF1 (N59, N57);
buf BUF1 (N60, N59);
xor XOR2 (N61, N54, N57);
and AND3 (N62, N48, N51, N61);
xor XOR2 (N63, N34, N58);
nor NOR4 (N64, N17, N18, N63, N39);
nand NAND3 (N65, N22, N62, N56);
not NOT1 (N66, N14);
not NOT1 (N67, N39);
buf BUF1 (N68, N38);
not NOT1 (N69, N64);
nand NAND4 (N70, N52, N31, N8, N43);
xor XOR2 (N71, N27, N70);
or OR4 (N72, N35, N14, N43, N63);
xor XOR2 (N73, N55, N20);
nand NAND3 (N74, N68, N19, N47);
xor XOR2 (N75, N71, N50);
nand NAND2 (N76, N67, N36);
nand NAND3 (N77, N66, N59, N61);
and AND2 (N78, N72, N16);
or OR3 (N79, N77, N42, N14);
buf BUF1 (N80, N74);
buf BUF1 (N81, N79);
nor NOR2 (N82, N81, N21);
or OR4 (N83, N60, N82, N46, N5);
not NOT1 (N84, N4);
and AND3 (N85, N73, N65, N57);
or OR2 (N86, N72, N60);
nor NOR2 (N87, N85, N13);
xor XOR2 (N88, N86, N19);
nand NAND3 (N89, N80, N59, N63);
or OR3 (N90, N78, N6, N64);
buf BUF1 (N91, N83);
nor NOR3 (N92, N88, N27, N65);
and AND2 (N93, N75, N31);
nor NOR4 (N94, N53, N66, N58, N80);
or OR3 (N95, N91, N93, N50);
or OR3 (N96, N11, N88, N73);
buf BUF1 (N97, N84);
or OR2 (N98, N94, N51);
nand NAND4 (N99, N89, N72, N35, N37);
not NOT1 (N100, N69);
nand NAND4 (N101, N96, N2, N70, N100);
and AND3 (N102, N50, N57, N43);
and AND4 (N103, N98, N10, N18, N51);
xor XOR2 (N104, N87, N74);
nor NOR2 (N105, N103, N84);
or OR2 (N106, N102, N10);
not NOT1 (N107, N95);
xor XOR2 (N108, N106, N39);
nor NOR3 (N109, N101, N17, N33);
and AND4 (N110, N109, N52, N26, N94);
buf BUF1 (N111, N99);
and AND2 (N112, N92, N37);
nand NAND2 (N113, N104, N13);
or OR3 (N114, N76, N95, N32);
or OR4 (N115, N110, N49, N85, N32);
buf BUF1 (N116, N111);
xor XOR2 (N117, N116, N111);
nor NOR2 (N118, N114, N90);
nand NAND4 (N119, N36, N2, N9, N55);
buf BUF1 (N120, N108);
nor NOR3 (N121, N97, N87, N25);
or OR2 (N122, N117, N21);
xor XOR2 (N123, N118, N97);
and AND2 (N124, N107, N120);
buf BUF1 (N125, N91);
nor NOR2 (N126, N115, N78);
and AND2 (N127, N124, N1);
xor XOR2 (N128, N127, N113);
xor XOR2 (N129, N74, N30);
and AND2 (N130, N105, N116);
xor XOR2 (N131, N122, N38);
xor XOR2 (N132, N131, N28);
or OR4 (N133, N128, N58, N44, N23);
nand NAND4 (N134, N132, N80, N79, N49);
and AND2 (N135, N125, N62);
nand NAND2 (N136, N133, N4);
or OR2 (N137, N130, N46);
nor NOR4 (N138, N126, N27, N56, N125);
not NOT1 (N139, N135);
nand NAND3 (N140, N138, N108, N10);
or OR2 (N141, N134, N37);
xor XOR2 (N142, N129, N42);
buf BUF1 (N143, N141);
xor XOR2 (N144, N142, N87);
xor XOR2 (N145, N119, N141);
or OR3 (N146, N121, N39, N58);
xor XOR2 (N147, N140, N92);
buf BUF1 (N148, N112);
nor NOR2 (N149, N139, N35);
xor XOR2 (N150, N145, N86);
or OR2 (N151, N149, N134);
xor XOR2 (N152, N147, N54);
nor NOR4 (N153, N151, N142, N89, N29);
not NOT1 (N154, N148);
not NOT1 (N155, N152);
or OR4 (N156, N146, N27, N110, N154);
and AND3 (N157, N12, N102, N101);
and AND2 (N158, N136, N142);
buf BUF1 (N159, N150);
not NOT1 (N160, N158);
nand NAND2 (N161, N143, N131);
nand NAND4 (N162, N160, N71, N158, N113);
or OR3 (N163, N159, N8, N13);
or OR3 (N164, N157, N99, N8);
and AND3 (N165, N161, N25, N97);
nand NAND4 (N166, N155, N46, N148, N7);
nand NAND3 (N167, N164, N141, N10);
or OR4 (N168, N144, N159, N5, N98);
nor NOR3 (N169, N167, N20, N118);
not NOT1 (N170, N137);
or OR3 (N171, N163, N50, N168);
xor XOR2 (N172, N129, N91);
not NOT1 (N173, N166);
and AND2 (N174, N153, N150);
nor NOR4 (N175, N170, N35, N90, N59);
or OR2 (N176, N173, N1);
not NOT1 (N177, N174);
buf BUF1 (N178, N156);
xor XOR2 (N179, N162, N161);
or OR2 (N180, N171, N141);
not NOT1 (N181, N176);
not NOT1 (N182, N181);
nand NAND4 (N183, N165, N59, N43, N23);
not NOT1 (N184, N179);
xor XOR2 (N185, N177, N66);
and AND3 (N186, N184, N17, N49);
nor NOR4 (N187, N185, N178, N22, N186);
buf BUF1 (N188, N37);
and AND2 (N189, N58, N71);
xor XOR2 (N190, N183, N122);
buf BUF1 (N191, N188);
xor XOR2 (N192, N180, N121);
nor NOR4 (N193, N175, N89, N25, N92);
not NOT1 (N194, N169);
nor NOR2 (N195, N192, N42);
and AND3 (N196, N190, N102, N21);
not NOT1 (N197, N187);
not NOT1 (N198, N197);
or OR3 (N199, N193, N119, N27);
nand NAND2 (N200, N182, N185);
and AND4 (N201, N198, N160, N64, N53);
buf BUF1 (N202, N199);
or OR4 (N203, N202, N167, N114, N126);
nor NOR3 (N204, N172, N59, N6);
buf BUF1 (N205, N195);
nor NOR4 (N206, N189, N3, N62, N97);
and AND2 (N207, N203, N31);
not NOT1 (N208, N123);
nor NOR3 (N209, N206, N6, N153);
not NOT1 (N210, N200);
nand NAND2 (N211, N205, N123);
xor XOR2 (N212, N201, N172);
xor XOR2 (N213, N196, N145);
or OR3 (N214, N207, N174, N107);
buf BUF1 (N215, N204);
and AND4 (N216, N215, N61, N57, N167);
and AND4 (N217, N212, N128, N193, N81);
and AND4 (N218, N194, N32, N35, N100);
nand NAND2 (N219, N209, N210);
xor XOR2 (N220, N87, N113);
not NOT1 (N221, N191);
nor NOR3 (N222, N217, N114, N221);
not NOT1 (N223, N101);
and AND3 (N224, N213, N188, N85);
nand NAND3 (N225, N214, N111, N45);
xor XOR2 (N226, N216, N136);
buf BUF1 (N227, N218);
xor XOR2 (N228, N208, N29);
xor XOR2 (N229, N222, N69);
nor NOR2 (N230, N229, N28);
buf BUF1 (N231, N226);
buf BUF1 (N232, N219);
or OR3 (N233, N232, N104, N227);
nor NOR4 (N234, N66, N138, N199, N152);
nor NOR2 (N235, N223, N226);
buf BUF1 (N236, N224);
nor NOR4 (N237, N211, N218, N222, N115);
nor NOR4 (N238, N233, N147, N10, N222);
xor XOR2 (N239, N231, N120);
buf BUF1 (N240, N236);
or OR4 (N241, N234, N198, N93, N121);
buf BUF1 (N242, N225);
and AND3 (N243, N241, N100, N74);
nor NOR2 (N244, N228, N51);
buf BUF1 (N245, N220);
nand NAND4 (N246, N244, N16, N55, N243);
not NOT1 (N247, N40);
nand NAND2 (N248, N242, N89);
and AND4 (N249, N247, N81, N95, N1);
and AND4 (N250, N230, N239, N244, N10);
or OR4 (N251, N208, N160, N72, N140);
nor NOR2 (N252, N235, N160);
xor XOR2 (N253, N251, N250);
or OR4 (N254, N249, N68, N217, N16);
not NOT1 (N255, N221);
or OR4 (N256, N253, N80, N28, N82);
buf BUF1 (N257, N246);
xor XOR2 (N258, N248, N46);
or OR4 (N259, N237, N188, N132, N9);
not NOT1 (N260, N259);
nor NOR2 (N261, N254, N71);
nand NAND3 (N262, N257, N181, N250);
xor XOR2 (N263, N260, N113);
buf BUF1 (N264, N263);
nand NAND4 (N265, N238, N63, N111, N64);
nand NAND3 (N266, N264, N20, N211);
nand NAND4 (N267, N261, N99, N95, N157);
and AND3 (N268, N256, N202, N132);
and AND3 (N269, N245, N36, N120);
not NOT1 (N270, N269);
nand NAND3 (N271, N252, N233, N263);
not NOT1 (N272, N265);
or OR2 (N273, N255, N25);
and AND2 (N274, N266, N177);
and AND3 (N275, N262, N101, N264);
nor NOR2 (N276, N268, N205);
and AND2 (N277, N272, N273);
xor XOR2 (N278, N156, N161);
not NOT1 (N279, N275);
not NOT1 (N280, N274);
buf BUF1 (N281, N270);
xor XOR2 (N282, N278, N269);
nand NAND3 (N283, N277, N90, N282);
xor XOR2 (N284, N249, N174);
or OR2 (N285, N283, N214);
buf BUF1 (N286, N285);
xor XOR2 (N287, N279, N220);
xor XOR2 (N288, N284, N269);
nor NOR4 (N289, N286, N287, N100, N112);
nor NOR2 (N290, N289, N249);
nand NAND2 (N291, N48, N163);
nor NOR2 (N292, N281, N28);
buf BUF1 (N293, N276);
xor XOR2 (N294, N240, N206);
or OR2 (N295, N258, N34);
nor NOR4 (N296, N292, N149, N73, N140);
buf BUF1 (N297, N296);
buf BUF1 (N298, N271);
buf BUF1 (N299, N294);
xor XOR2 (N300, N293, N16);
buf BUF1 (N301, N299);
not NOT1 (N302, N295);
xor XOR2 (N303, N298, N158);
and AND4 (N304, N297, N229, N174, N204);
nor NOR3 (N305, N301, N144, N272);
nand NAND2 (N306, N305, N293);
buf BUF1 (N307, N280);
nand NAND2 (N308, N291, N165);
nor NOR3 (N309, N302, N124, N53);
nor NOR4 (N310, N288, N250, N281, N81);
and AND2 (N311, N308, N295);
buf BUF1 (N312, N303);
buf BUF1 (N313, N300);
not NOT1 (N314, N307);
or OR2 (N315, N267, N254);
and AND4 (N316, N315, N103, N53, N6);
nand NAND4 (N317, N313, N266, N217, N305);
and AND3 (N318, N311, N113, N66);
nor NOR3 (N319, N304, N60, N68);
or OR4 (N320, N314, N214, N269, N276);
and AND4 (N321, N320, N294, N162, N301);
and AND4 (N322, N310, N143, N11, N89);
nor NOR2 (N323, N309, N244);
xor XOR2 (N324, N323, N87);
nand NAND3 (N325, N324, N20, N257);
nor NOR4 (N326, N317, N237, N321, N207);
nand NAND2 (N327, N49, N220);
nand NAND3 (N328, N322, N68, N83);
nor NOR3 (N329, N326, N23, N12);
xor XOR2 (N330, N328, N253);
xor XOR2 (N331, N290, N219);
not NOT1 (N332, N327);
nand NAND2 (N333, N325, N134);
buf BUF1 (N334, N333);
xor XOR2 (N335, N331, N22);
and AND4 (N336, N318, N198, N167, N161);
nor NOR4 (N337, N329, N3, N182, N186);
buf BUF1 (N338, N332);
not NOT1 (N339, N336);
buf BUF1 (N340, N338);
and AND4 (N341, N316, N86, N236, N162);
nor NOR4 (N342, N339, N309, N161, N338);
nor NOR4 (N343, N312, N213, N15, N341);
nand NAND3 (N344, N147, N67, N287);
xor XOR2 (N345, N330, N255);
nand NAND3 (N346, N343, N321, N198);
or OR3 (N347, N344, N4, N327);
buf BUF1 (N348, N340);
nor NOR3 (N349, N346, N167, N216);
nand NAND3 (N350, N348, N262, N39);
nor NOR2 (N351, N349, N23);
xor XOR2 (N352, N350, N230);
nor NOR4 (N353, N352, N170, N78, N106);
nand NAND4 (N354, N342, N148, N221, N23);
xor XOR2 (N355, N345, N73);
nor NOR2 (N356, N353, N186);
not NOT1 (N357, N351);
not NOT1 (N358, N334);
and AND4 (N359, N357, N17, N140, N312);
and AND4 (N360, N358, N188, N198, N141);
or OR2 (N361, N306, N240);
or OR2 (N362, N356, N260);
buf BUF1 (N363, N337);
or OR3 (N364, N362, N219, N194);
buf BUF1 (N365, N347);
not NOT1 (N366, N363);
not NOT1 (N367, N360);
xor XOR2 (N368, N355, N108);
and AND2 (N369, N361, N56);
or OR3 (N370, N369, N352, N72);
and AND2 (N371, N335, N301);
or OR3 (N372, N319, N289, N262);
nand NAND3 (N373, N371, N357, N97);
or OR4 (N374, N364, N99, N173, N162);
xor XOR2 (N375, N359, N38);
nand NAND2 (N376, N366, N9);
not NOT1 (N377, N374);
xor XOR2 (N378, N368, N58);
not NOT1 (N379, N378);
nor NOR2 (N380, N375, N41);
nand NAND4 (N381, N370, N31, N250, N191);
or OR4 (N382, N377, N106, N218, N100);
and AND3 (N383, N373, N192, N250);
nand NAND4 (N384, N367, N77, N377, N70);
xor XOR2 (N385, N365, N330);
nor NOR3 (N386, N372, N168, N169);
or OR2 (N387, N385, N125);
nor NOR2 (N388, N384, N244);
or OR3 (N389, N381, N9, N24);
nor NOR3 (N390, N388, N385, N99);
nand NAND3 (N391, N354, N65, N341);
not NOT1 (N392, N380);
buf BUF1 (N393, N387);
nand NAND4 (N394, N379, N311, N189, N216);
nor NOR2 (N395, N383, N297);
and AND3 (N396, N382, N67, N376);
nor NOR4 (N397, N258, N87, N161, N389);
not NOT1 (N398, N94);
xor XOR2 (N399, N391, N33);
buf BUF1 (N400, N386);
and AND4 (N401, N390, N379, N77, N292);
nand NAND2 (N402, N396, N255);
and AND4 (N403, N393, N49, N23, N307);
or OR2 (N404, N392, N154);
and AND4 (N405, N402, N295, N351, N77);
and AND4 (N406, N397, N299, N206, N209);
nor NOR2 (N407, N394, N52);
nor NOR2 (N408, N395, N220);
nor NOR4 (N409, N404, N386, N68, N283);
and AND3 (N410, N399, N26, N103);
nor NOR4 (N411, N408, N251, N362, N358);
xor XOR2 (N412, N411, N89);
nand NAND4 (N413, N403, N80, N43, N382);
xor XOR2 (N414, N410, N390);
nand NAND2 (N415, N413, N216);
not NOT1 (N416, N398);
and AND4 (N417, N416, N10, N112, N36);
nand NAND4 (N418, N409, N403, N102, N268);
not NOT1 (N419, N407);
nor NOR2 (N420, N406, N75);
nor NOR2 (N421, N415, N281);
and AND3 (N422, N418, N53, N122);
nand NAND3 (N423, N412, N177, N217);
and AND4 (N424, N400, N383, N237, N262);
or OR3 (N425, N417, N53, N246);
and AND2 (N426, N421, N5);
nand NAND4 (N427, N422, N299, N198, N262);
xor XOR2 (N428, N427, N409);
and AND4 (N429, N426, N426, N350, N36);
and AND3 (N430, N429, N148, N262);
nor NOR2 (N431, N423, N224);
xor XOR2 (N432, N430, N407);
and AND3 (N433, N419, N431, N350);
nand NAND4 (N434, N6, N106, N249, N122);
buf BUF1 (N435, N425);
and AND3 (N436, N424, N313, N402);
nand NAND2 (N437, N436, N5);
nand NAND2 (N438, N405, N167);
xor XOR2 (N439, N435, N149);
buf BUF1 (N440, N438);
xor XOR2 (N441, N428, N199);
and AND2 (N442, N437, N396);
or OR2 (N443, N440, N4);
not NOT1 (N444, N442);
buf BUF1 (N445, N444);
nand NAND3 (N446, N432, N90, N353);
xor XOR2 (N447, N441, N419);
buf BUF1 (N448, N420);
not NOT1 (N449, N434);
nor NOR2 (N450, N439, N428);
nand NAND2 (N451, N447, N449);
xor XOR2 (N452, N281, N232);
nor NOR2 (N453, N450, N315);
buf BUF1 (N454, N401);
nor NOR3 (N455, N414, N84, N326);
nand NAND2 (N456, N455, N194);
or OR4 (N457, N443, N448, N347, N100);
not NOT1 (N458, N73);
and AND2 (N459, N458, N321);
or OR3 (N460, N456, N29, N189);
nor NOR2 (N461, N445, N8);
buf BUF1 (N462, N452);
and AND2 (N463, N433, N133);
xor XOR2 (N464, N454, N154);
and AND3 (N465, N464, N102, N242);
not NOT1 (N466, N461);
nor NOR3 (N467, N460, N113, N404);
not NOT1 (N468, N467);
not NOT1 (N469, N462);
and AND3 (N470, N453, N3, N297);
or OR2 (N471, N470, N340);
or OR3 (N472, N457, N196, N231);
not NOT1 (N473, N469);
xor XOR2 (N474, N468, N471);
xor XOR2 (N475, N340, N87);
nor NOR4 (N476, N472, N234, N429, N323);
not NOT1 (N477, N459);
xor XOR2 (N478, N475, N384);
xor XOR2 (N479, N474, N206);
and AND4 (N480, N479, N339, N236, N463);
and AND3 (N481, N211, N254, N278);
nor NOR2 (N482, N446, N57);
buf BUF1 (N483, N478);
and AND3 (N484, N465, N223, N148);
and AND4 (N485, N484, N277, N195, N289);
nand NAND4 (N486, N483, N478, N405, N480);
nor NOR2 (N487, N449, N446);
xor XOR2 (N488, N473, N154);
nor NOR4 (N489, N481, N190, N375, N329);
nor NOR2 (N490, N451, N278);
not NOT1 (N491, N466);
or OR3 (N492, N487, N54, N292);
buf BUF1 (N493, N492);
or OR3 (N494, N491, N481, N315);
not NOT1 (N495, N477);
nand NAND3 (N496, N489, N421, N97);
nor NOR4 (N497, N490, N249, N121, N171);
not NOT1 (N498, N482);
nand NAND2 (N499, N493, N277);
xor XOR2 (N500, N488, N138);
not NOT1 (N501, N499);
nor NOR4 (N502, N501, N452, N205, N194);
and AND3 (N503, N497, N257, N73);
buf BUF1 (N504, N498);
not NOT1 (N505, N495);
or OR3 (N506, N504, N191, N193);
nor NOR3 (N507, N485, N327, N19);
not NOT1 (N508, N494);
and AND3 (N509, N486, N356, N216);
nor NOR4 (N510, N506, N129, N267, N390);
or OR4 (N511, N505, N309, N87, N484);
nor NOR4 (N512, N511, N271, N268, N354);
not NOT1 (N513, N510);
nor NOR4 (N514, N509, N169, N455, N318);
nand NAND2 (N515, N507, N245);
nor NOR4 (N516, N514, N29, N4, N497);
buf BUF1 (N517, N513);
and AND2 (N518, N515, N355);
and AND4 (N519, N516, N484, N85, N163);
nor NOR4 (N520, N476, N63, N28, N410);
or OR3 (N521, N500, N439, N334);
nor NOR4 (N522, N521, N185, N510, N262);
buf BUF1 (N523, N522);
and AND4 (N524, N520, N273, N42, N482);
buf BUF1 (N525, N508);
or OR3 (N526, N518, N433, N339);
nor NOR4 (N527, N512, N27, N411, N332);
xor XOR2 (N528, N503, N250);
buf BUF1 (N529, N502);
and AND3 (N530, N524, N126, N204);
nand NAND4 (N531, N526, N432, N199, N350);
nand NAND3 (N532, N529, N497, N96);
buf BUF1 (N533, N527);
buf BUF1 (N534, N530);
nand NAND4 (N535, N525, N364, N231, N102);
and AND3 (N536, N531, N50, N254);
not NOT1 (N537, N496);
xor XOR2 (N538, N533, N486);
and AND2 (N539, N523, N477);
and AND2 (N540, N517, N153);
nor NOR2 (N541, N535, N28);
nand NAND2 (N542, N537, N86);
and AND2 (N543, N538, N2);
xor XOR2 (N544, N528, N75);
not NOT1 (N545, N519);
buf BUF1 (N546, N534);
not NOT1 (N547, N536);
xor XOR2 (N548, N539, N277);
nor NOR2 (N549, N542, N516);
and AND2 (N550, N545, N171);
nor NOR4 (N551, N541, N248, N259, N103);
buf BUF1 (N552, N540);
and AND3 (N553, N550, N162, N487);
not NOT1 (N554, N552);
nand NAND4 (N555, N543, N474, N46, N179);
buf BUF1 (N556, N544);
xor XOR2 (N557, N556, N437);
nand NAND4 (N558, N548, N318, N182, N34);
nor NOR2 (N559, N553, N333);
nor NOR3 (N560, N547, N388, N406);
or OR4 (N561, N546, N28, N414, N511);
nand NAND4 (N562, N551, N118, N369, N138);
nand NAND2 (N563, N554, N479);
xor XOR2 (N564, N555, N337);
and AND2 (N565, N564, N512);
nor NOR4 (N566, N549, N39, N504, N78);
xor XOR2 (N567, N566, N140);
nand NAND3 (N568, N561, N15, N546);
not NOT1 (N569, N568);
or OR3 (N570, N532, N220, N321);
and AND2 (N571, N563, N317);
xor XOR2 (N572, N571, N532);
not NOT1 (N573, N572);
nor NOR4 (N574, N558, N215, N464, N243);
xor XOR2 (N575, N574, N562);
nand NAND2 (N576, N411, N407);
nor NOR4 (N577, N569, N282, N46, N341);
not NOT1 (N578, N557);
nand NAND3 (N579, N567, N563, N5);
not NOT1 (N580, N565);
nand NAND3 (N581, N570, N419, N508);
or OR4 (N582, N576, N304, N382, N17);
xor XOR2 (N583, N579, N364);
nand NAND2 (N584, N573, N329);
nor NOR3 (N585, N577, N147, N244);
buf BUF1 (N586, N560);
or OR3 (N587, N575, N418, N61);
and AND4 (N588, N585, N587, N97, N56);
nor NOR4 (N589, N129, N137, N122, N56);
xor XOR2 (N590, N578, N51);
and AND2 (N591, N586, N269);
and AND3 (N592, N588, N204, N156);
xor XOR2 (N593, N592, N71);
nand NAND2 (N594, N583, N87);
and AND2 (N595, N581, N285);
nor NOR4 (N596, N591, N218, N227, N589);
nand NAND4 (N597, N502, N375, N596, N37);
nor NOR4 (N598, N72, N86, N168, N86);
and AND2 (N599, N590, N430);
nand NAND2 (N600, N597, N472);
nor NOR2 (N601, N584, N180);
nand NAND4 (N602, N559, N182, N429, N457);
nand NAND3 (N603, N602, N303, N338);
not NOT1 (N604, N599);
not NOT1 (N605, N600);
xor XOR2 (N606, N582, N372);
xor XOR2 (N607, N580, N333);
nor NOR4 (N608, N605, N260, N195, N455);
xor XOR2 (N609, N598, N29);
nor NOR2 (N610, N609, N357);
buf BUF1 (N611, N608);
and AND3 (N612, N611, N136, N44);
xor XOR2 (N613, N594, N607);
nor NOR4 (N614, N106, N431, N154, N284);
and AND3 (N615, N606, N490, N55);
and AND2 (N616, N601, N467);
nand NAND3 (N617, N613, N401, N278);
buf BUF1 (N618, N617);
buf BUF1 (N619, N618);
and AND2 (N620, N615, N616);
and AND3 (N621, N282, N547, N86);
not NOT1 (N622, N620);
nor NOR2 (N623, N621, N333);
buf BUF1 (N624, N610);
nor NOR4 (N625, N624, N436, N12, N377);
xor XOR2 (N626, N593, N598);
not NOT1 (N627, N614);
and AND4 (N628, N623, N621, N462, N460);
xor XOR2 (N629, N612, N45);
not NOT1 (N630, N603);
not NOT1 (N631, N630);
not NOT1 (N632, N622);
or OR3 (N633, N628, N143, N3);
xor XOR2 (N634, N631, N113);
or OR2 (N635, N633, N275);
nand NAND3 (N636, N635, N492, N24);
not NOT1 (N637, N625);
nor NOR3 (N638, N629, N424, N549);
not NOT1 (N639, N637);
nand NAND4 (N640, N638, N452, N117, N301);
nand NAND2 (N641, N626, N329);
not NOT1 (N642, N634);
buf BUF1 (N643, N595);
buf BUF1 (N644, N642);
not NOT1 (N645, N641);
not NOT1 (N646, N636);
or OR3 (N647, N645, N209, N288);
xor XOR2 (N648, N639, N518);
and AND3 (N649, N646, N476, N440);
or OR2 (N650, N604, N597);
and AND3 (N651, N650, N468, N242);
nor NOR4 (N652, N632, N543, N516, N418);
xor XOR2 (N653, N652, N359);
nand NAND3 (N654, N619, N71, N540);
nand NAND2 (N655, N651, N320);
nor NOR4 (N656, N655, N472, N494, N18);
nand NAND2 (N657, N648, N630);
nand NAND2 (N658, N644, N396);
not NOT1 (N659, N656);
and AND2 (N660, N627, N333);
not NOT1 (N661, N640);
xor XOR2 (N662, N660, N467);
nor NOR2 (N663, N653, N144);
and AND4 (N664, N658, N178, N596, N388);
nand NAND2 (N665, N649, N63);
and AND2 (N666, N661, N401);
or OR4 (N667, N662, N193, N335, N257);
nor NOR4 (N668, N667, N369, N256, N151);
and AND2 (N669, N664, N531);
not NOT1 (N670, N643);
nor NOR4 (N671, N668, N59, N85, N570);
nand NAND2 (N672, N671, N368);
xor XOR2 (N673, N663, N85);
or OR3 (N674, N669, N50, N4);
buf BUF1 (N675, N659);
not NOT1 (N676, N672);
not NOT1 (N677, N676);
not NOT1 (N678, N647);
buf BUF1 (N679, N677);
not NOT1 (N680, N673);
nor NOR3 (N681, N678, N146, N163);
nor NOR4 (N682, N654, N204, N231, N91);
not NOT1 (N683, N674);
or OR2 (N684, N670, N14);
buf BUF1 (N685, N675);
or OR3 (N686, N683, N613, N463);
nand NAND3 (N687, N665, N598, N169);
nor NOR2 (N688, N666, N225);
nand NAND4 (N689, N688, N100, N338, N462);
nor NOR4 (N690, N679, N189, N362, N612);
nor NOR4 (N691, N685, N488, N297, N276);
and AND4 (N692, N684, N145, N557, N91);
not NOT1 (N693, N690);
buf BUF1 (N694, N657);
nand NAND4 (N695, N680, N639, N365, N48);
xor XOR2 (N696, N686, N267);
not NOT1 (N697, N693);
xor XOR2 (N698, N687, N319);
buf BUF1 (N699, N697);
nand NAND3 (N700, N689, N617, N446);
nor NOR3 (N701, N694, N68, N40);
nor NOR2 (N702, N700, N263);
not NOT1 (N703, N681);
and AND3 (N704, N702, N304, N88);
and AND2 (N705, N698, N391);
nand NAND2 (N706, N705, N25);
or OR2 (N707, N682, N660);
buf BUF1 (N708, N691);
nor NOR3 (N709, N701, N88, N288);
or OR4 (N710, N703, N284, N100, N340);
buf BUF1 (N711, N707);
buf BUF1 (N712, N695);
and AND4 (N713, N704, N623, N225, N73);
and AND2 (N714, N712, N692);
or OR3 (N715, N207, N325, N104);
or OR2 (N716, N699, N639);
not NOT1 (N717, N708);
not NOT1 (N718, N710);
and AND4 (N719, N716, N368, N145, N224);
and AND4 (N720, N696, N672, N97, N636);
nor NOR4 (N721, N711, N477, N84, N111);
not NOT1 (N722, N720);
not NOT1 (N723, N717);
and AND4 (N724, N722, N191, N36, N128);
buf BUF1 (N725, N706);
nor NOR4 (N726, N719, N31, N149, N433);
and AND2 (N727, N713, N203);
nand NAND4 (N728, N715, N233, N419, N489);
and AND2 (N729, N714, N287);
nand NAND3 (N730, N725, N77, N184);
nor NOR4 (N731, N728, N155, N277, N350);
or OR4 (N732, N724, N421, N108, N1);
xor XOR2 (N733, N709, N176);
nand NAND4 (N734, N733, N298, N516, N306);
xor XOR2 (N735, N732, N188);
xor XOR2 (N736, N730, N336);
or OR3 (N737, N726, N420, N434);
and AND3 (N738, N718, N581, N114);
or OR2 (N739, N731, N612);
or OR2 (N740, N738, N285);
buf BUF1 (N741, N729);
nor NOR4 (N742, N739, N684, N550, N724);
nor NOR4 (N743, N741, N337, N65, N559);
buf BUF1 (N744, N734);
and AND4 (N745, N737, N594, N360, N637);
nand NAND4 (N746, N736, N560, N639, N645);
nand NAND3 (N747, N743, N253, N287);
xor XOR2 (N748, N744, N574);
xor XOR2 (N749, N747, N227);
and AND4 (N750, N745, N188, N186, N15);
nor NOR2 (N751, N748, N276);
or OR2 (N752, N721, N576);
nand NAND2 (N753, N751, N213);
buf BUF1 (N754, N752);
nand NAND2 (N755, N735, N461);
not NOT1 (N756, N754);
not NOT1 (N757, N753);
buf BUF1 (N758, N723);
buf BUF1 (N759, N749);
buf BUF1 (N760, N746);
xor XOR2 (N761, N759, N701);
and AND4 (N762, N755, N661, N503, N761);
nor NOR3 (N763, N672, N737, N482);
buf BUF1 (N764, N742);
nor NOR3 (N765, N757, N433, N745);
and AND4 (N766, N750, N344, N245, N668);
or OR3 (N767, N740, N633, N676);
nand NAND2 (N768, N765, N259);
or OR4 (N769, N727, N383, N627, N521);
nor NOR3 (N770, N769, N686, N702);
or OR3 (N771, N768, N635, N242);
and AND4 (N772, N762, N298, N735, N713);
xor XOR2 (N773, N771, N680);
nor NOR4 (N774, N773, N540, N608, N538);
nand NAND2 (N775, N764, N535);
buf BUF1 (N776, N775);
nor NOR3 (N777, N776, N3, N161);
nand NAND2 (N778, N777, N755);
or OR2 (N779, N778, N571);
or OR2 (N780, N774, N156);
or OR2 (N781, N772, N192);
nor NOR4 (N782, N758, N454, N151, N733);
nand NAND2 (N783, N781, N229);
and AND4 (N784, N782, N301, N52, N81);
buf BUF1 (N785, N760);
buf BUF1 (N786, N785);
and AND3 (N787, N756, N321, N520);
xor XOR2 (N788, N767, N674);
nor NOR2 (N789, N784, N219);
and AND2 (N790, N766, N190);
not NOT1 (N791, N763);
or OR4 (N792, N788, N123, N145, N54);
or OR2 (N793, N789, N77);
xor XOR2 (N794, N780, N197);
not NOT1 (N795, N791);
and AND2 (N796, N795, N335);
buf BUF1 (N797, N779);
nor NOR2 (N798, N787, N448);
xor XOR2 (N799, N793, N337);
nor NOR2 (N800, N796, N743);
nor NOR3 (N801, N792, N785, N134);
nand NAND3 (N802, N799, N593, N660);
or OR3 (N803, N800, N205, N9);
not NOT1 (N804, N797);
or OR4 (N805, N798, N73, N543, N447);
xor XOR2 (N806, N802, N162);
and AND3 (N807, N805, N426, N265);
buf BUF1 (N808, N807);
not NOT1 (N809, N783);
xor XOR2 (N810, N803, N791);
not NOT1 (N811, N794);
buf BUF1 (N812, N806);
and AND3 (N813, N790, N744, N373);
nand NAND2 (N814, N770, N213);
and AND2 (N815, N812, N764);
not NOT1 (N816, N814);
xor XOR2 (N817, N804, N449);
or OR4 (N818, N815, N423, N588, N639);
xor XOR2 (N819, N801, N738);
or OR4 (N820, N786, N338, N454, N643);
and AND3 (N821, N820, N106, N364);
nor NOR4 (N822, N811, N674, N192, N780);
and AND2 (N823, N821, N29);
nand NAND4 (N824, N822, N499, N675, N415);
buf BUF1 (N825, N818);
nand NAND3 (N826, N816, N347, N447);
not NOT1 (N827, N819);
and AND3 (N828, N827, N166, N616);
not NOT1 (N829, N817);
or OR2 (N830, N824, N580);
or OR4 (N831, N810, N290, N406, N472);
nand NAND2 (N832, N829, N539);
nand NAND3 (N833, N828, N108, N316);
nand NAND4 (N834, N808, N409, N665, N691);
xor XOR2 (N835, N830, N479);
buf BUF1 (N836, N831);
and AND3 (N837, N826, N123, N685);
or OR2 (N838, N832, N546);
nor NOR3 (N839, N825, N606, N630);
nand NAND2 (N840, N839, N310);
or OR4 (N841, N836, N463, N166, N167);
xor XOR2 (N842, N833, N574);
nand NAND2 (N843, N823, N773);
nand NAND4 (N844, N837, N796, N54, N315);
nor NOR3 (N845, N809, N600, N574);
buf BUF1 (N846, N835);
nand NAND4 (N847, N844, N257, N496, N165);
buf BUF1 (N848, N840);
nor NOR2 (N849, N847, N201);
or OR2 (N850, N846, N698);
nor NOR3 (N851, N845, N145, N163);
and AND3 (N852, N851, N473, N224);
nor NOR3 (N853, N842, N767, N825);
nor NOR2 (N854, N849, N236);
or OR4 (N855, N813, N125, N353, N88);
nor NOR4 (N856, N834, N495, N415, N818);
and AND2 (N857, N838, N503);
xor XOR2 (N858, N852, N57);
nor NOR4 (N859, N850, N174, N392, N538);
or OR4 (N860, N853, N189, N528, N388);
xor XOR2 (N861, N857, N527);
nor NOR3 (N862, N861, N771, N354);
or OR3 (N863, N841, N170, N360);
or OR4 (N864, N858, N663, N478, N708);
xor XOR2 (N865, N854, N327);
nand NAND4 (N866, N856, N608, N475, N552);
xor XOR2 (N867, N860, N630);
or OR3 (N868, N863, N90, N619);
nand NAND4 (N869, N848, N94, N714, N361);
buf BUF1 (N870, N866);
nand NAND4 (N871, N870, N103, N804, N491);
nor NOR3 (N872, N855, N91, N106);
and AND3 (N873, N869, N852, N228);
and AND4 (N874, N871, N475, N601, N320);
xor XOR2 (N875, N843, N77);
buf BUF1 (N876, N862);
buf BUF1 (N877, N872);
not NOT1 (N878, N877);
nor NOR2 (N879, N875, N629);
or OR3 (N880, N864, N504, N505);
and AND3 (N881, N874, N66, N218);
nand NAND4 (N882, N881, N129, N422, N139);
nand NAND4 (N883, N859, N803, N188, N565);
buf BUF1 (N884, N865);
not NOT1 (N885, N873);
xor XOR2 (N886, N884, N421);
nor NOR3 (N887, N879, N309, N413);
or OR4 (N888, N887, N332, N56, N810);
nor NOR2 (N889, N886, N283);
buf BUF1 (N890, N868);
xor XOR2 (N891, N880, N29);
not NOT1 (N892, N890);
or OR3 (N893, N892, N730, N78);
and AND3 (N894, N883, N731, N286);
buf BUF1 (N895, N891);
or OR2 (N896, N882, N226);
buf BUF1 (N897, N896);
nor NOR4 (N898, N876, N554, N547, N172);
nor NOR4 (N899, N867, N454, N736, N709);
xor XOR2 (N900, N885, N503);
nand NAND2 (N901, N894, N541);
and AND4 (N902, N893, N746, N423, N323);
or OR4 (N903, N900, N631, N134, N550);
buf BUF1 (N904, N903);
buf BUF1 (N905, N878);
nand NAND3 (N906, N902, N598, N874);
nor NOR3 (N907, N901, N153, N627);
xor XOR2 (N908, N906, N26);
or OR3 (N909, N899, N310, N174);
buf BUF1 (N910, N895);
nand NAND2 (N911, N898, N83);
not NOT1 (N912, N905);
nand NAND4 (N913, N912, N233, N213, N236);
nor NOR3 (N914, N907, N505, N824);
or OR3 (N915, N911, N298, N557);
not NOT1 (N916, N914);
and AND3 (N917, N916, N734, N325);
or OR4 (N918, N915, N322, N453, N88);
not NOT1 (N919, N908);
or OR2 (N920, N917, N321);
buf BUF1 (N921, N909);
nand NAND2 (N922, N889, N146);
xor XOR2 (N923, N919, N326);
xor XOR2 (N924, N888, N833);
not NOT1 (N925, N910);
or OR3 (N926, N925, N184, N79);
nand NAND2 (N927, N921, N633);
and AND4 (N928, N904, N871, N834, N119);
xor XOR2 (N929, N918, N645);
buf BUF1 (N930, N897);
nor NOR2 (N931, N923, N623);
or OR2 (N932, N927, N400);
nor NOR4 (N933, N926, N724, N391, N276);
or OR4 (N934, N933, N1, N399, N237);
xor XOR2 (N935, N913, N904);
nor NOR4 (N936, N929, N98, N278, N868);
xor XOR2 (N937, N924, N790);
xor XOR2 (N938, N934, N596);
or OR3 (N939, N931, N626, N116);
and AND4 (N940, N920, N369, N174, N20);
buf BUF1 (N941, N940);
nand NAND4 (N942, N937, N155, N421, N33);
or OR4 (N943, N935, N559, N397, N659);
not NOT1 (N944, N941);
nor NOR2 (N945, N942, N393);
or OR3 (N946, N938, N571, N830);
not NOT1 (N947, N945);
xor XOR2 (N948, N946, N71);
and AND4 (N949, N948, N893, N604, N545);
nor NOR2 (N950, N928, N190);
not NOT1 (N951, N936);
nand NAND4 (N952, N939, N428, N821, N696);
nor NOR3 (N953, N947, N350, N360);
not NOT1 (N954, N951);
and AND3 (N955, N953, N584, N388);
nor NOR3 (N956, N950, N497, N93);
nand NAND4 (N957, N930, N620, N152, N277);
xor XOR2 (N958, N932, N222);
nor NOR4 (N959, N922, N175, N672, N633);
buf BUF1 (N960, N954);
nor NOR3 (N961, N949, N100, N728);
and AND2 (N962, N944, N171);
xor XOR2 (N963, N957, N461);
and AND3 (N964, N961, N658, N460);
and AND3 (N965, N958, N712, N196);
and AND3 (N966, N959, N517, N959);
or OR2 (N967, N956, N672);
nand NAND2 (N968, N965, N174);
buf BUF1 (N969, N962);
not NOT1 (N970, N964);
buf BUF1 (N971, N968);
nand NAND3 (N972, N952, N805, N366);
xor XOR2 (N973, N960, N494);
buf BUF1 (N974, N971);
buf BUF1 (N975, N969);
nor NOR4 (N976, N970, N593, N565, N705);
buf BUF1 (N977, N963);
nand NAND2 (N978, N973, N106);
nand NAND2 (N979, N976, N83);
and AND4 (N980, N977, N465, N278, N216);
buf BUF1 (N981, N943);
and AND3 (N982, N974, N513, N261);
xor XOR2 (N983, N979, N208);
or OR2 (N984, N982, N943);
xor XOR2 (N985, N984, N541);
buf BUF1 (N986, N983);
nor NOR4 (N987, N955, N841, N385, N986);
xor XOR2 (N988, N341, N284);
buf BUF1 (N989, N981);
nand NAND3 (N990, N972, N840, N681);
buf BUF1 (N991, N975);
or OR4 (N992, N967, N748, N9, N450);
and AND3 (N993, N966, N451, N337);
nor NOR2 (N994, N987, N618);
buf BUF1 (N995, N985);
xor XOR2 (N996, N994, N209);
nor NOR4 (N997, N988, N149, N474, N48);
buf BUF1 (N998, N978);
or OR3 (N999, N996, N641, N270);
and AND3 (N1000, N991, N911, N795);
nor NOR3 (N1001, N990, N160, N504);
xor XOR2 (N1002, N999, N618);
and AND3 (N1003, N989, N85, N850);
or OR2 (N1004, N1002, N947);
and AND2 (N1005, N980, N614);
not NOT1 (N1006, N1000);
nor NOR3 (N1007, N998, N481, N770);
and AND3 (N1008, N993, N518, N266);
nand NAND4 (N1009, N1006, N831, N195, N73);
xor XOR2 (N1010, N995, N875);
xor XOR2 (N1011, N1008, N513);
xor XOR2 (N1012, N1001, N724);
and AND2 (N1013, N1012, N952);
nor NOR2 (N1014, N1011, N135);
or OR3 (N1015, N1013, N902, N382);
nand NAND3 (N1016, N1005, N923, N1006);
buf BUF1 (N1017, N1007);
not NOT1 (N1018, N1017);
xor XOR2 (N1019, N997, N86);
buf BUF1 (N1020, N1003);
xor XOR2 (N1021, N1020, N332);
and AND3 (N1022, N1018, N444, N933);
and AND3 (N1023, N1016, N423, N286);
nand NAND3 (N1024, N1004, N309, N907);
not NOT1 (N1025, N1019);
nand NAND2 (N1026, N1010, N532);
or OR3 (N1027, N1009, N852, N79);
and AND3 (N1028, N992, N584, N827);
nand NAND2 (N1029, N1028, N474);
buf BUF1 (N1030, N1027);
not NOT1 (N1031, N1014);
not NOT1 (N1032, N1025);
not NOT1 (N1033, N1023);
buf BUF1 (N1034, N1031);
buf BUF1 (N1035, N1026);
xor XOR2 (N1036, N1022, N199);
nand NAND3 (N1037, N1021, N621, N869);
not NOT1 (N1038, N1030);
not NOT1 (N1039, N1032);
and AND4 (N1040, N1038, N206, N744, N744);
nand NAND3 (N1041, N1035, N920, N896);
not NOT1 (N1042, N1024);
not NOT1 (N1043, N1033);
and AND4 (N1044, N1034, N512, N219, N615);
nor NOR3 (N1045, N1015, N982, N755);
not NOT1 (N1046, N1036);
xor XOR2 (N1047, N1044, N314);
or OR4 (N1048, N1043, N324, N635, N96);
not NOT1 (N1049, N1037);
xor XOR2 (N1050, N1040, N1047);
or OR4 (N1051, N295, N545, N461, N743);
nand NAND3 (N1052, N1039, N643, N964);
xor XOR2 (N1053, N1049, N104);
and AND2 (N1054, N1041, N815);
nand NAND2 (N1055, N1052, N932);
not NOT1 (N1056, N1029);
buf BUF1 (N1057, N1046);
nor NOR2 (N1058, N1055, N889);
xor XOR2 (N1059, N1053, N738);
nand NAND4 (N1060, N1057, N444, N778, N467);
or OR4 (N1061, N1059, N147, N831, N386);
nor NOR4 (N1062, N1042, N238, N919, N515);
not NOT1 (N1063, N1050);
and AND4 (N1064, N1054, N877, N215, N22);
buf BUF1 (N1065, N1056);
or OR3 (N1066, N1060, N930, N245);
xor XOR2 (N1067, N1062, N284);
or OR2 (N1068, N1058, N346);
and AND2 (N1069, N1051, N686);
nor NOR2 (N1070, N1064, N375);
or OR3 (N1071, N1067, N140, N22);
nor NOR3 (N1072, N1070, N560, N858);
buf BUF1 (N1073, N1065);
nand NAND2 (N1074, N1045, N696);
nand NAND2 (N1075, N1066, N205);
not NOT1 (N1076, N1072);
buf BUF1 (N1077, N1063);
or OR2 (N1078, N1075, N167);
not NOT1 (N1079, N1074);
not NOT1 (N1080, N1077);
nand NAND3 (N1081, N1073, N200, N242);
and AND4 (N1082, N1080, N269, N858, N425);
nor NOR3 (N1083, N1048, N501, N355);
nand NAND3 (N1084, N1076, N594, N710);
and AND4 (N1085, N1071, N76, N22, N96);
not NOT1 (N1086, N1078);
buf BUF1 (N1087, N1085);
not NOT1 (N1088, N1087);
xor XOR2 (N1089, N1082, N1032);
not NOT1 (N1090, N1081);
nand NAND2 (N1091, N1061, N759);
nand NAND3 (N1092, N1088, N430, N1043);
and AND4 (N1093, N1091, N348, N195, N375);
or OR4 (N1094, N1090, N559, N675, N842);
not NOT1 (N1095, N1079);
buf BUF1 (N1096, N1086);
and AND2 (N1097, N1095, N149);
xor XOR2 (N1098, N1093, N186);
xor XOR2 (N1099, N1092, N785);
nor NOR4 (N1100, N1098, N207, N384, N687);
or OR3 (N1101, N1089, N121, N1045);
and AND3 (N1102, N1097, N888, N517);
or OR2 (N1103, N1100, N284);
nor NOR2 (N1104, N1096, N158);
not NOT1 (N1105, N1084);
nor NOR3 (N1106, N1102, N620, N801);
nor NOR4 (N1107, N1068, N239, N172, N484);
or OR3 (N1108, N1107, N739, N406);
or OR3 (N1109, N1103, N549, N928);
and AND2 (N1110, N1083, N481);
not NOT1 (N1111, N1109);
and AND2 (N1112, N1108, N632);
xor XOR2 (N1113, N1104, N324);
and AND3 (N1114, N1113, N1086, N957);
xor XOR2 (N1115, N1069, N145);
or OR4 (N1116, N1099, N5, N125, N90);
or OR2 (N1117, N1110, N388);
or OR4 (N1118, N1106, N210, N558, N11);
nand NAND4 (N1119, N1118, N511, N736, N490);
or OR3 (N1120, N1115, N159, N557);
nor NOR3 (N1121, N1101, N492, N649);
or OR3 (N1122, N1120, N511, N1035);
and AND2 (N1123, N1111, N72);
or OR2 (N1124, N1116, N216);
nor NOR2 (N1125, N1124, N778);
and AND3 (N1126, N1121, N130, N1051);
and AND4 (N1127, N1119, N333, N131, N1048);
not NOT1 (N1128, N1094);
nor NOR4 (N1129, N1125, N90, N1015, N586);
nor NOR2 (N1130, N1117, N940);
not NOT1 (N1131, N1105);
not NOT1 (N1132, N1127);
buf BUF1 (N1133, N1128);
nor NOR4 (N1134, N1123, N961, N45, N221);
nand NAND2 (N1135, N1114, N364);
or OR4 (N1136, N1130, N1090, N842, N500);
not NOT1 (N1137, N1134);
nand NAND2 (N1138, N1126, N503);
buf BUF1 (N1139, N1133);
not NOT1 (N1140, N1137);
buf BUF1 (N1141, N1112);
buf BUF1 (N1142, N1129);
and AND2 (N1143, N1131, N688);
and AND2 (N1144, N1141, N927);
or OR2 (N1145, N1144, N697);
nor NOR3 (N1146, N1140, N21, N394);
and AND2 (N1147, N1132, N900);
and AND2 (N1148, N1122, N189);
nand NAND2 (N1149, N1136, N225);
and AND4 (N1150, N1138, N165, N912, N791);
xor XOR2 (N1151, N1142, N524);
buf BUF1 (N1152, N1145);
and AND4 (N1153, N1151, N386, N831, N988);
xor XOR2 (N1154, N1149, N102);
or OR2 (N1155, N1152, N1054);
or OR3 (N1156, N1155, N537, N1039);
nand NAND4 (N1157, N1153, N817, N260, N603);
buf BUF1 (N1158, N1148);
and AND4 (N1159, N1146, N230, N629, N1047);
or OR2 (N1160, N1135, N1036);
buf BUF1 (N1161, N1150);
buf BUF1 (N1162, N1154);
buf BUF1 (N1163, N1162);
and AND3 (N1164, N1158, N1155, N321);
not NOT1 (N1165, N1147);
not NOT1 (N1166, N1160);
xor XOR2 (N1167, N1139, N748);
or OR2 (N1168, N1166, N939);
xor XOR2 (N1169, N1157, N1028);
buf BUF1 (N1170, N1168);
not NOT1 (N1171, N1156);
nor NOR3 (N1172, N1159, N539, N863);
or OR4 (N1173, N1165, N807, N1033, N455);
and AND2 (N1174, N1169, N1063);
nand NAND3 (N1175, N1167, N390, N242);
not NOT1 (N1176, N1143);
buf BUF1 (N1177, N1172);
nand NAND3 (N1178, N1170, N764, N916);
xor XOR2 (N1179, N1171, N629);
buf BUF1 (N1180, N1173);
or OR4 (N1181, N1176, N656, N609, N949);
and AND2 (N1182, N1181, N752);
and AND4 (N1183, N1163, N412, N877, N728);
or OR2 (N1184, N1175, N899);
xor XOR2 (N1185, N1164, N622);
and AND3 (N1186, N1184, N17, N1114);
buf BUF1 (N1187, N1161);
xor XOR2 (N1188, N1185, N471);
buf BUF1 (N1189, N1186);
nor NOR4 (N1190, N1189, N1019, N692, N1074);
xor XOR2 (N1191, N1174, N156);
and AND2 (N1192, N1178, N445);
or OR3 (N1193, N1182, N370, N515);
and AND4 (N1194, N1193, N852, N620, N681);
and AND2 (N1195, N1179, N707);
or OR2 (N1196, N1177, N77);
not NOT1 (N1197, N1190);
xor XOR2 (N1198, N1196, N1114);
nand NAND3 (N1199, N1188, N929, N634);
nand NAND4 (N1200, N1192, N568, N694, N884);
or OR4 (N1201, N1198, N361, N835, N1158);
not NOT1 (N1202, N1195);
and AND3 (N1203, N1200, N1037, N1182);
buf BUF1 (N1204, N1187);
nand NAND2 (N1205, N1199, N1138);
nand NAND2 (N1206, N1191, N20);
nand NAND4 (N1207, N1194, N359, N29, N225);
not NOT1 (N1208, N1201);
buf BUF1 (N1209, N1202);
not NOT1 (N1210, N1183);
not NOT1 (N1211, N1204);
not NOT1 (N1212, N1211);
not NOT1 (N1213, N1203);
not NOT1 (N1214, N1213);
xor XOR2 (N1215, N1208, N995);
or OR4 (N1216, N1180, N83, N726, N948);
buf BUF1 (N1217, N1206);
nand NAND4 (N1218, N1216, N456, N89, N34);
buf BUF1 (N1219, N1210);
not NOT1 (N1220, N1218);
nand NAND3 (N1221, N1214, N463, N1192);
not NOT1 (N1222, N1209);
buf BUF1 (N1223, N1219);
xor XOR2 (N1224, N1197, N1197);
and AND2 (N1225, N1222, N1068);
not NOT1 (N1226, N1217);
not NOT1 (N1227, N1226);
or OR4 (N1228, N1215, N973, N458, N426);
not NOT1 (N1229, N1205);
and AND4 (N1230, N1228, N75, N162, N226);
nor NOR3 (N1231, N1207, N927, N307);
not NOT1 (N1232, N1230);
buf BUF1 (N1233, N1212);
buf BUF1 (N1234, N1232);
not NOT1 (N1235, N1234);
nand NAND3 (N1236, N1220, N142, N728);
buf BUF1 (N1237, N1231);
or OR4 (N1238, N1229, N883, N881, N738);
buf BUF1 (N1239, N1224);
nand NAND4 (N1240, N1237, N473, N119, N611);
or OR4 (N1241, N1235, N452, N1060, N1116);
not NOT1 (N1242, N1240);
not NOT1 (N1243, N1242);
buf BUF1 (N1244, N1239);
xor XOR2 (N1245, N1244, N524);
not NOT1 (N1246, N1223);
nor NOR4 (N1247, N1241, N927, N578, N1064);
nor NOR4 (N1248, N1246, N1016, N303, N61);
not NOT1 (N1249, N1243);
nor NOR4 (N1250, N1247, N7, N639, N593);
nand NAND3 (N1251, N1227, N936, N1156);
nor NOR4 (N1252, N1248, N547, N38, N532);
and AND4 (N1253, N1238, N479, N751, N342);
and AND2 (N1254, N1252, N716);
xor XOR2 (N1255, N1245, N671);
or OR2 (N1256, N1251, N515);
buf BUF1 (N1257, N1225);
nand NAND2 (N1258, N1257, N58);
not NOT1 (N1259, N1254);
and AND3 (N1260, N1259, N496, N280);
nor NOR4 (N1261, N1255, N1144, N719, N1256);
nand NAND3 (N1262, N1107, N1127, N677);
xor XOR2 (N1263, N1221, N699);
nand NAND4 (N1264, N1253, N101, N202, N939);
nor NOR4 (N1265, N1258, N94, N862, N689);
xor XOR2 (N1266, N1261, N456);
and AND4 (N1267, N1260, N625, N998, N1110);
not NOT1 (N1268, N1236);
buf BUF1 (N1269, N1250);
and AND3 (N1270, N1266, N514, N847);
nand NAND3 (N1271, N1264, N613, N996);
xor XOR2 (N1272, N1270, N349);
nand NAND4 (N1273, N1265, N580, N577, N1227);
xor XOR2 (N1274, N1269, N425);
not NOT1 (N1275, N1262);
nand NAND2 (N1276, N1275, N834);
nand NAND2 (N1277, N1249, N1042);
not NOT1 (N1278, N1263);
nand NAND2 (N1279, N1273, N1087);
buf BUF1 (N1280, N1272);
buf BUF1 (N1281, N1274);
nand NAND3 (N1282, N1277, N554, N584);
xor XOR2 (N1283, N1282, N1046);
nor NOR3 (N1284, N1278, N1184, N1043);
nand NAND3 (N1285, N1283, N1067, N56);
and AND3 (N1286, N1267, N490, N38);
nor NOR4 (N1287, N1276, N268, N398, N488);
and AND4 (N1288, N1271, N161, N846, N478);
xor XOR2 (N1289, N1285, N108);
or OR4 (N1290, N1281, N596, N603, N1251);
nand NAND4 (N1291, N1279, N627, N486, N1229);
and AND2 (N1292, N1268, N1265);
and AND3 (N1293, N1286, N226, N1191);
xor XOR2 (N1294, N1280, N907);
nor NOR2 (N1295, N1292, N282);
and AND3 (N1296, N1233, N518, N1229);
and AND3 (N1297, N1293, N899, N567);
or OR3 (N1298, N1287, N1049, N1);
nor NOR4 (N1299, N1289, N774, N511, N583);
not NOT1 (N1300, N1296);
or OR2 (N1301, N1284, N313);
not NOT1 (N1302, N1291);
buf BUF1 (N1303, N1302);
or OR4 (N1304, N1297, N742, N649, N935);
not NOT1 (N1305, N1295);
or OR2 (N1306, N1298, N729);
nor NOR3 (N1307, N1301, N279, N886);
buf BUF1 (N1308, N1290);
and AND2 (N1309, N1307, N1139);
nand NAND2 (N1310, N1308, N69);
not NOT1 (N1311, N1310);
xor XOR2 (N1312, N1304, N1277);
or OR2 (N1313, N1300, N631);
or OR4 (N1314, N1311, N271, N963, N288);
xor XOR2 (N1315, N1313, N766);
and AND3 (N1316, N1299, N1086, N1207);
buf BUF1 (N1317, N1312);
buf BUF1 (N1318, N1294);
not NOT1 (N1319, N1314);
not NOT1 (N1320, N1315);
nand NAND4 (N1321, N1319, N541, N874, N1205);
not NOT1 (N1322, N1321);
nand NAND2 (N1323, N1309, N303);
and AND3 (N1324, N1316, N451, N332);
or OR4 (N1325, N1303, N868, N174, N596);
and AND4 (N1326, N1322, N72, N988, N40);
nand NAND4 (N1327, N1326, N365, N154, N1012);
buf BUF1 (N1328, N1324);
buf BUF1 (N1329, N1288);
xor XOR2 (N1330, N1327, N506);
nand NAND3 (N1331, N1305, N817, N912);
buf BUF1 (N1332, N1329);
and AND3 (N1333, N1331, N1226, N41);
buf BUF1 (N1334, N1332);
not NOT1 (N1335, N1318);
not NOT1 (N1336, N1317);
not NOT1 (N1337, N1330);
nand NAND4 (N1338, N1334, N594, N717, N753);
or OR4 (N1339, N1337, N1013, N228, N999);
or OR3 (N1340, N1339, N1217, N823);
xor XOR2 (N1341, N1325, N270);
or OR2 (N1342, N1306, N945);
not NOT1 (N1343, N1336);
nand NAND4 (N1344, N1338, N751, N387, N195);
not NOT1 (N1345, N1323);
nand NAND2 (N1346, N1320, N1124);
or OR2 (N1347, N1341, N857);
xor XOR2 (N1348, N1344, N945);
nor NOR4 (N1349, N1335, N49, N1341, N411);
buf BUF1 (N1350, N1345);
and AND4 (N1351, N1340, N284, N184, N1125);
or OR2 (N1352, N1349, N891);
and AND4 (N1353, N1347, N320, N1248, N259);
not NOT1 (N1354, N1351);
buf BUF1 (N1355, N1352);
nor NOR4 (N1356, N1354, N415, N1201, N350);
buf BUF1 (N1357, N1333);
or OR2 (N1358, N1357, N839);
nand NAND3 (N1359, N1358, N615, N788);
nand NAND3 (N1360, N1359, N76, N380);
not NOT1 (N1361, N1356);
nor NOR3 (N1362, N1350, N376, N114);
buf BUF1 (N1363, N1328);
nor NOR3 (N1364, N1362, N1319, N819);
buf BUF1 (N1365, N1355);
and AND4 (N1366, N1342, N32, N532, N173);
not NOT1 (N1367, N1366);
not NOT1 (N1368, N1360);
buf BUF1 (N1369, N1353);
and AND4 (N1370, N1369, N305, N58, N885);
buf BUF1 (N1371, N1367);
not NOT1 (N1372, N1364);
nand NAND4 (N1373, N1370, N647, N829, N1187);
and AND2 (N1374, N1346, N867);
and AND4 (N1375, N1372, N362, N165, N732);
nand NAND4 (N1376, N1375, N305, N1236, N570);
not NOT1 (N1377, N1343);
or OR2 (N1378, N1376, N696);
nand NAND4 (N1379, N1377, N614, N602, N982);
buf BUF1 (N1380, N1348);
nand NAND3 (N1381, N1371, N155, N481);
buf BUF1 (N1382, N1361);
xor XOR2 (N1383, N1378, N404);
buf BUF1 (N1384, N1383);
or OR3 (N1385, N1380, N903, N803);
and AND4 (N1386, N1385, N670, N472, N634);
and AND3 (N1387, N1379, N1368, N1134);
not NOT1 (N1388, N1323);
nand NAND2 (N1389, N1381, N1207);
nor NOR2 (N1390, N1384, N25);
buf BUF1 (N1391, N1373);
buf BUF1 (N1392, N1386);
nor NOR2 (N1393, N1363, N846);
nand NAND4 (N1394, N1387, N1340, N901, N830);
or OR3 (N1395, N1382, N999, N246);
not NOT1 (N1396, N1365);
and AND2 (N1397, N1374, N1086);
nand NAND3 (N1398, N1389, N1068, N371);
and AND4 (N1399, N1388, N723, N965, N24);
or OR4 (N1400, N1390, N249, N489, N1296);
and AND4 (N1401, N1391, N574, N1205, N986);
and AND3 (N1402, N1392, N982, N542);
nor NOR4 (N1403, N1395, N955, N744, N401);
buf BUF1 (N1404, N1403);
nand NAND3 (N1405, N1401, N27, N1135);
not NOT1 (N1406, N1400);
and AND3 (N1407, N1405, N1382, N1307);
nand NAND3 (N1408, N1406, N171, N523);
nor NOR4 (N1409, N1398, N1155, N1386, N586);
and AND2 (N1410, N1394, N1037);
not NOT1 (N1411, N1402);
nor NOR3 (N1412, N1410, N260, N518);
nand NAND2 (N1413, N1407, N660);
buf BUF1 (N1414, N1399);
buf BUF1 (N1415, N1393);
and AND4 (N1416, N1396, N8, N85, N154);
and AND3 (N1417, N1411, N1096, N846);
buf BUF1 (N1418, N1416);
nand NAND3 (N1419, N1404, N961, N488);
buf BUF1 (N1420, N1419);
or OR3 (N1421, N1408, N700, N302);
nor NOR2 (N1422, N1397, N864);
or OR3 (N1423, N1422, N1231, N137);
not NOT1 (N1424, N1423);
not NOT1 (N1425, N1414);
nand NAND2 (N1426, N1425, N1144);
buf BUF1 (N1427, N1426);
buf BUF1 (N1428, N1417);
xor XOR2 (N1429, N1427, N760);
or OR3 (N1430, N1424, N1032, N793);
and AND4 (N1431, N1428, N885, N1064, N540);
or OR4 (N1432, N1409, N246, N1375, N1370);
or OR4 (N1433, N1430, N590, N1396, N168);
or OR4 (N1434, N1412, N588, N302, N1095);
buf BUF1 (N1435, N1420);
or OR2 (N1436, N1429, N142);
nand NAND2 (N1437, N1418, N908);
or OR3 (N1438, N1435, N1415, N364);
nand NAND4 (N1439, N175, N1251, N982, N1396);
and AND2 (N1440, N1431, N165);
buf BUF1 (N1441, N1438);
or OR3 (N1442, N1421, N369, N838);
nand NAND2 (N1443, N1440, N1053);
and AND4 (N1444, N1443, N141, N647, N1216);
nand NAND4 (N1445, N1442, N1163, N1295, N693);
nor NOR2 (N1446, N1445, N1275);
and AND2 (N1447, N1436, N278);
nor NOR3 (N1448, N1413, N27, N210);
or OR2 (N1449, N1448, N439);
buf BUF1 (N1450, N1444);
or OR4 (N1451, N1446, N242, N857, N1354);
or OR4 (N1452, N1449, N246, N253, N12);
buf BUF1 (N1453, N1432);
or OR4 (N1454, N1447, N24, N22, N886);
and AND4 (N1455, N1454, N342, N689, N465);
or OR2 (N1456, N1451, N412);
buf BUF1 (N1457, N1434);
not NOT1 (N1458, N1441);
xor XOR2 (N1459, N1453, N170);
not NOT1 (N1460, N1452);
or OR4 (N1461, N1450, N1007, N768, N1438);
or OR2 (N1462, N1456, N910);
buf BUF1 (N1463, N1439);
xor XOR2 (N1464, N1455, N695);
or OR3 (N1465, N1461, N1374, N221);
or OR4 (N1466, N1465, N445, N148, N1169);
xor XOR2 (N1467, N1466, N819);
and AND2 (N1468, N1437, N35);
and AND2 (N1469, N1458, N584);
not NOT1 (N1470, N1462);
not NOT1 (N1471, N1468);
or OR4 (N1472, N1470, N1334, N1044, N1239);
nor NOR2 (N1473, N1457, N1332);
and AND4 (N1474, N1433, N357, N377, N441);
nand NAND4 (N1475, N1472, N845, N682, N147);
buf BUF1 (N1476, N1467);
and AND3 (N1477, N1469, N69, N909);
and AND4 (N1478, N1464, N937, N1334, N358);
nand NAND4 (N1479, N1474, N189, N1019, N384);
nand NAND2 (N1480, N1476, N800);
or OR4 (N1481, N1459, N1425, N665, N342);
nor NOR4 (N1482, N1475, N537, N436, N529);
or OR4 (N1483, N1463, N298, N888, N733);
and AND2 (N1484, N1481, N535);
nor NOR3 (N1485, N1477, N457, N1087);
and AND4 (N1486, N1460, N979, N450, N901);
and AND4 (N1487, N1471, N727, N1236, N490);
xor XOR2 (N1488, N1484, N226);
nor NOR4 (N1489, N1483, N1374, N1195, N1030);
nand NAND4 (N1490, N1478, N569, N71, N606);
xor XOR2 (N1491, N1487, N1155);
and AND3 (N1492, N1480, N276, N562);
and AND2 (N1493, N1489, N1340);
nor NOR3 (N1494, N1479, N786, N1413);
nor NOR3 (N1495, N1482, N993, N1079);
not NOT1 (N1496, N1485);
nand NAND3 (N1497, N1490, N20, N203);
nor NOR2 (N1498, N1494, N1069);
nor NOR3 (N1499, N1493, N1248, N56);
and AND2 (N1500, N1486, N601);
or OR4 (N1501, N1492, N467, N1008, N636);
not NOT1 (N1502, N1498);
nand NAND4 (N1503, N1501, N93, N6, N823);
and AND2 (N1504, N1500, N451);
nand NAND4 (N1505, N1499, N112, N1013, N526);
nor NOR3 (N1506, N1502, N328, N224);
and AND4 (N1507, N1488, N353, N1372, N1107);
or OR3 (N1508, N1505, N420, N193);
nor NOR2 (N1509, N1507, N489);
nor NOR4 (N1510, N1509, N1206, N518, N247);
or OR2 (N1511, N1491, N422);
not NOT1 (N1512, N1497);
nor NOR4 (N1513, N1512, N97, N857, N961);
xor XOR2 (N1514, N1495, N1143);
and AND4 (N1515, N1511, N790, N1332, N262);
not NOT1 (N1516, N1510);
not NOT1 (N1517, N1504);
not NOT1 (N1518, N1473);
nor NOR2 (N1519, N1506, N298);
xor XOR2 (N1520, N1516, N906);
and AND4 (N1521, N1508, N814, N1080, N587);
nand NAND2 (N1522, N1520, N1379);
and AND4 (N1523, N1522, N1363, N370, N1190);
buf BUF1 (N1524, N1518);
nor NOR2 (N1525, N1519, N1468);
not NOT1 (N1526, N1521);
nor NOR2 (N1527, N1496, N429);
not NOT1 (N1528, N1515);
or OR2 (N1529, N1528, N1212);
or OR4 (N1530, N1525, N703, N1419, N620);
xor XOR2 (N1531, N1503, N851);
buf BUF1 (N1532, N1526);
buf BUF1 (N1533, N1513);
nand NAND4 (N1534, N1531, N1127, N529, N1291);
and AND2 (N1535, N1534, N37);
or OR4 (N1536, N1535, N1276, N542, N318);
or OR4 (N1537, N1529, N421, N695, N1258);
nor NOR3 (N1538, N1532, N1411, N1381);
buf BUF1 (N1539, N1530);
or OR2 (N1540, N1538, N1010);
or OR4 (N1541, N1533, N1007, N1190, N684);
not NOT1 (N1542, N1540);
and AND2 (N1543, N1524, N284);
nor NOR4 (N1544, N1523, N912, N487, N963);
xor XOR2 (N1545, N1537, N379);
or OR2 (N1546, N1541, N325);
nor NOR3 (N1547, N1514, N1345, N261);
not NOT1 (N1548, N1547);
nand NAND2 (N1549, N1548, N1305);
buf BUF1 (N1550, N1545);
nor NOR3 (N1551, N1542, N581, N1530);
and AND4 (N1552, N1527, N921, N1213, N389);
nand NAND2 (N1553, N1549, N1339);
or OR4 (N1554, N1544, N77, N731, N1394);
or OR4 (N1555, N1539, N439, N727, N1355);
buf BUF1 (N1556, N1536);
nand NAND3 (N1557, N1556, N1521, N44);
and AND3 (N1558, N1552, N128, N499);
and AND2 (N1559, N1557, N379);
xor XOR2 (N1560, N1555, N1164);
and AND3 (N1561, N1554, N894, N1458);
buf BUF1 (N1562, N1560);
nand NAND3 (N1563, N1558, N556, N829);
xor XOR2 (N1564, N1563, N1460);
buf BUF1 (N1565, N1562);
buf BUF1 (N1566, N1559);
not NOT1 (N1567, N1546);
nand NAND2 (N1568, N1561, N142);
buf BUF1 (N1569, N1517);
or OR2 (N1570, N1566, N232);
and AND4 (N1571, N1570, N63, N121, N251);
or OR2 (N1572, N1553, N53);
xor XOR2 (N1573, N1550, N1207);
xor XOR2 (N1574, N1551, N9);
xor XOR2 (N1575, N1567, N1434);
and AND2 (N1576, N1571, N476);
nand NAND2 (N1577, N1575, N1521);
and AND4 (N1578, N1543, N1154, N125, N996);
nand NAND4 (N1579, N1577, N24, N1210, N1190);
xor XOR2 (N1580, N1578, N1316);
xor XOR2 (N1581, N1580, N445);
buf BUF1 (N1582, N1573);
buf BUF1 (N1583, N1582);
or OR2 (N1584, N1565, N1126);
nor NOR4 (N1585, N1569, N155, N551, N820);
nor NOR2 (N1586, N1581, N1477);
xor XOR2 (N1587, N1568, N145);
buf BUF1 (N1588, N1574);
not NOT1 (N1589, N1586);
not NOT1 (N1590, N1584);
not NOT1 (N1591, N1585);
and AND3 (N1592, N1590, N370, N694);
or OR4 (N1593, N1564, N21, N1502, N1037);
xor XOR2 (N1594, N1591, N985);
xor XOR2 (N1595, N1583, N40);
buf BUF1 (N1596, N1595);
or OR2 (N1597, N1587, N1439);
nor NOR3 (N1598, N1596, N642, N23);
nand NAND4 (N1599, N1593, N897, N728, N817);
xor XOR2 (N1600, N1576, N222);
buf BUF1 (N1601, N1572);
buf BUF1 (N1602, N1601);
buf BUF1 (N1603, N1602);
nor NOR3 (N1604, N1579, N711, N726);
nand NAND2 (N1605, N1592, N201);
not NOT1 (N1606, N1605);
nand NAND2 (N1607, N1603, N1552);
nor NOR2 (N1608, N1597, N1527);
not NOT1 (N1609, N1607);
nand NAND4 (N1610, N1589, N906, N716, N1166);
or OR2 (N1611, N1598, N365);
or OR4 (N1612, N1610, N908, N695, N1102);
xor XOR2 (N1613, N1604, N810);
buf BUF1 (N1614, N1612);
not NOT1 (N1615, N1614);
and AND4 (N1616, N1599, N509, N544, N348);
not NOT1 (N1617, N1600);
buf BUF1 (N1618, N1616);
xor XOR2 (N1619, N1608, N907);
not NOT1 (N1620, N1613);
xor XOR2 (N1621, N1609, N1491);
xor XOR2 (N1622, N1615, N71);
and AND4 (N1623, N1617, N956, N334, N372);
not NOT1 (N1624, N1622);
and AND3 (N1625, N1623, N1160, N513);
nor NOR3 (N1626, N1625, N28, N56);
and AND3 (N1627, N1618, N86, N218);
xor XOR2 (N1628, N1627, N938);
nand NAND3 (N1629, N1621, N1540, N418);
xor XOR2 (N1630, N1606, N1180);
and AND3 (N1631, N1628, N803, N116);
buf BUF1 (N1632, N1629);
buf BUF1 (N1633, N1588);
nand NAND3 (N1634, N1631, N479, N986);
nand NAND2 (N1635, N1594, N517);
nand NAND4 (N1636, N1619, N653, N1319, N837);
and AND3 (N1637, N1626, N485, N1048);
or OR2 (N1638, N1637, N444);
or OR4 (N1639, N1632, N1346, N1626, N1025);
not NOT1 (N1640, N1636);
nand NAND3 (N1641, N1611, N470, N276);
nand NAND4 (N1642, N1633, N1357, N738, N872);
nor NOR3 (N1643, N1638, N318, N556);
nor NOR4 (N1644, N1620, N966, N213, N1303);
buf BUF1 (N1645, N1643);
buf BUF1 (N1646, N1639);
nand NAND2 (N1647, N1645, N680);
not NOT1 (N1648, N1635);
xor XOR2 (N1649, N1624, N1584);
nand NAND4 (N1650, N1634, N1122, N767, N551);
buf BUF1 (N1651, N1646);
and AND4 (N1652, N1649, N443, N676, N80);
not NOT1 (N1653, N1647);
or OR4 (N1654, N1641, N428, N1630, N1159);
not NOT1 (N1655, N1189);
buf BUF1 (N1656, N1640);
nand NAND2 (N1657, N1654, N66);
nor NOR2 (N1658, N1644, N1108);
xor XOR2 (N1659, N1652, N191);
xor XOR2 (N1660, N1656, N378);
or OR4 (N1661, N1655, N633, N337, N481);
nor NOR4 (N1662, N1660, N1128, N1025, N1152);
nand NAND2 (N1663, N1651, N656);
buf BUF1 (N1664, N1661);
buf BUF1 (N1665, N1650);
nand NAND2 (N1666, N1658, N125);
and AND2 (N1667, N1653, N1638);
xor XOR2 (N1668, N1665, N1641);
not NOT1 (N1669, N1667);
not NOT1 (N1670, N1664);
not NOT1 (N1671, N1662);
buf BUF1 (N1672, N1659);
nor NOR2 (N1673, N1666, N1004);
or OR3 (N1674, N1642, N78, N1442);
not NOT1 (N1675, N1648);
or OR3 (N1676, N1668, N159, N274);
buf BUF1 (N1677, N1670);
or OR4 (N1678, N1663, N1604, N358, N11);
and AND2 (N1679, N1678, N307);
or OR4 (N1680, N1673, N565, N1375, N545);
or OR2 (N1681, N1669, N381);
nor NOR3 (N1682, N1675, N284, N1157);
and AND3 (N1683, N1674, N1203, N657);
buf BUF1 (N1684, N1677);
nand NAND2 (N1685, N1671, N1532);
and AND3 (N1686, N1657, N835, N237);
buf BUF1 (N1687, N1683);
nand NAND2 (N1688, N1679, N149);
not NOT1 (N1689, N1688);
xor XOR2 (N1690, N1682, N694);
and AND4 (N1691, N1684, N1255, N171, N1461);
not NOT1 (N1692, N1690);
and AND3 (N1693, N1672, N1686, N84);
buf BUF1 (N1694, N1153);
buf BUF1 (N1695, N1687);
and AND2 (N1696, N1691, N489);
or OR3 (N1697, N1696, N646, N658);
nor NOR2 (N1698, N1681, N679);
buf BUF1 (N1699, N1676);
buf BUF1 (N1700, N1698);
nand NAND4 (N1701, N1700, N460, N519, N523);
xor XOR2 (N1702, N1697, N95);
buf BUF1 (N1703, N1702);
nor NOR2 (N1704, N1692, N1484);
nor NOR4 (N1705, N1685, N1338, N1567, N1325);
not NOT1 (N1706, N1705);
xor XOR2 (N1707, N1703, N1237);
nand NAND4 (N1708, N1699, N544, N120, N694);
not NOT1 (N1709, N1701);
nand NAND2 (N1710, N1704, N1440);
xor XOR2 (N1711, N1693, N821);
not NOT1 (N1712, N1707);
xor XOR2 (N1713, N1706, N1364);
nand NAND2 (N1714, N1709, N198);
nor NOR2 (N1715, N1711, N1201);
and AND4 (N1716, N1694, N1059, N1426, N1587);
xor XOR2 (N1717, N1710, N1483);
xor XOR2 (N1718, N1714, N999);
buf BUF1 (N1719, N1680);
and AND3 (N1720, N1715, N395, N622);
xor XOR2 (N1721, N1719, N466);
or OR3 (N1722, N1708, N368, N577);
nor NOR4 (N1723, N1720, N860, N1001, N210);
or OR2 (N1724, N1695, N1025);
or OR4 (N1725, N1689, N1122, N1012, N1062);
buf BUF1 (N1726, N1712);
xor XOR2 (N1727, N1721, N379);
not NOT1 (N1728, N1717);
or OR2 (N1729, N1723, N436);
nor NOR4 (N1730, N1718, N1104, N417, N747);
buf BUF1 (N1731, N1730);
nor NOR4 (N1732, N1726, N560, N516, N1405);
xor XOR2 (N1733, N1724, N1263);
or OR2 (N1734, N1733, N1228);
and AND3 (N1735, N1731, N1019, N768);
xor XOR2 (N1736, N1729, N1179);
xor XOR2 (N1737, N1716, N1427);
nor NOR4 (N1738, N1737, N1643, N1381, N1045);
not NOT1 (N1739, N1722);
and AND2 (N1740, N1732, N1620);
or OR3 (N1741, N1727, N920, N309);
nor NOR2 (N1742, N1736, N1492);
xor XOR2 (N1743, N1735, N225);
and AND4 (N1744, N1734, N1448, N313, N794);
xor XOR2 (N1745, N1742, N734);
xor XOR2 (N1746, N1725, N1319);
xor XOR2 (N1747, N1713, N65);
nand NAND4 (N1748, N1740, N623, N138, N84);
buf BUF1 (N1749, N1747);
or OR2 (N1750, N1748, N516);
or OR4 (N1751, N1728, N803, N875, N747);
and AND2 (N1752, N1743, N574);
not NOT1 (N1753, N1746);
buf BUF1 (N1754, N1752);
buf BUF1 (N1755, N1754);
xor XOR2 (N1756, N1745, N498);
and AND4 (N1757, N1755, N1713, N710, N1136);
and AND2 (N1758, N1741, N849);
xor XOR2 (N1759, N1758, N1386);
nand NAND2 (N1760, N1756, N726);
buf BUF1 (N1761, N1749);
or OR2 (N1762, N1738, N1219);
buf BUF1 (N1763, N1760);
and AND2 (N1764, N1739, N325);
or OR4 (N1765, N1750, N1155, N639, N468);
xor XOR2 (N1766, N1762, N1280);
and AND4 (N1767, N1764, N1335, N865, N829);
or OR2 (N1768, N1767, N1307);
buf BUF1 (N1769, N1766);
nand NAND2 (N1770, N1757, N1675);
nor NOR2 (N1771, N1751, N983);
and AND2 (N1772, N1765, N1110);
or OR3 (N1773, N1769, N1569, N1381);
xor XOR2 (N1774, N1768, N158);
nand NAND3 (N1775, N1761, N1161, N1271);
nor NOR4 (N1776, N1771, N1510, N1609, N1563);
or OR3 (N1777, N1774, N1237, N1703);
or OR3 (N1778, N1775, N757, N1638);
xor XOR2 (N1779, N1772, N1588);
and AND2 (N1780, N1759, N683);
xor XOR2 (N1781, N1777, N1343);
buf BUF1 (N1782, N1753);
or OR4 (N1783, N1779, N1432, N763, N964);
nor NOR2 (N1784, N1773, N1481);
nor NOR2 (N1785, N1783, N965);
not NOT1 (N1786, N1781);
not NOT1 (N1787, N1780);
and AND3 (N1788, N1770, N834, N424);
nand NAND4 (N1789, N1778, N471, N1550, N831);
or OR3 (N1790, N1789, N1659, N945);
not NOT1 (N1791, N1763);
or OR3 (N1792, N1744, N870, N216);
nand NAND2 (N1793, N1776, N542);
xor XOR2 (N1794, N1787, N1530);
xor XOR2 (N1795, N1788, N902);
or OR4 (N1796, N1792, N1044, N857, N1356);
xor XOR2 (N1797, N1782, N378);
nor NOR3 (N1798, N1793, N823, N654);
and AND2 (N1799, N1796, N644);
xor XOR2 (N1800, N1794, N1151);
and AND2 (N1801, N1795, N1117);
nand NAND3 (N1802, N1786, N11, N263);
nor NOR3 (N1803, N1798, N1785, N1782);
or OR3 (N1804, N1598, N570, N1527);
or OR4 (N1805, N1801, N1443, N1009, N39);
xor XOR2 (N1806, N1804, N869);
nand NAND3 (N1807, N1800, N502, N155);
or OR3 (N1808, N1803, N283, N481);
buf BUF1 (N1809, N1805);
and AND2 (N1810, N1807, N1518);
buf BUF1 (N1811, N1808);
nand NAND4 (N1812, N1806, N992, N829, N1270);
not NOT1 (N1813, N1810);
nor NOR3 (N1814, N1784, N1227, N1181);
nor NOR3 (N1815, N1802, N803, N731);
or OR4 (N1816, N1809, N722, N655, N575);
not NOT1 (N1817, N1813);
nor NOR3 (N1818, N1815, N63, N631);
not NOT1 (N1819, N1790);
or OR2 (N1820, N1814, N412);
buf BUF1 (N1821, N1797);
buf BUF1 (N1822, N1816);
nand NAND2 (N1823, N1818, N832);
xor XOR2 (N1824, N1811, N70);
not NOT1 (N1825, N1820);
nor NOR3 (N1826, N1822, N1554, N712);
xor XOR2 (N1827, N1819, N1388);
nand NAND4 (N1828, N1826, N727, N1032, N861);
and AND2 (N1829, N1799, N14);
or OR3 (N1830, N1791, N1003, N835);
and AND4 (N1831, N1823, N1167, N1652, N1614);
xor XOR2 (N1832, N1825, N1474);
or OR3 (N1833, N1812, N9, N598);
nand NAND4 (N1834, N1833, N1419, N85, N723);
not NOT1 (N1835, N1831);
buf BUF1 (N1836, N1821);
buf BUF1 (N1837, N1835);
and AND3 (N1838, N1832, N322, N886);
not NOT1 (N1839, N1827);
nand NAND2 (N1840, N1828, N1797);
xor XOR2 (N1841, N1834, N1651);
or OR4 (N1842, N1830, N590, N177, N371);
nand NAND2 (N1843, N1824, N1146);
buf BUF1 (N1844, N1836);
nor NOR3 (N1845, N1841, N1192, N1479);
xor XOR2 (N1846, N1838, N381);
not NOT1 (N1847, N1840);
buf BUF1 (N1848, N1846);
nand NAND4 (N1849, N1837, N340, N1376, N705);
xor XOR2 (N1850, N1844, N360);
or OR2 (N1851, N1829, N966);
and AND3 (N1852, N1843, N1386, N1136);
and AND3 (N1853, N1848, N96, N1091);
or OR4 (N1854, N1845, N1343, N1798, N1439);
and AND4 (N1855, N1817, N743, N982, N809);
not NOT1 (N1856, N1851);
xor XOR2 (N1857, N1842, N988);
xor XOR2 (N1858, N1847, N1408);
not NOT1 (N1859, N1849);
nand NAND3 (N1860, N1857, N1122, N125);
buf BUF1 (N1861, N1855);
or OR3 (N1862, N1853, N410, N1228);
xor XOR2 (N1863, N1862, N356);
buf BUF1 (N1864, N1863);
xor XOR2 (N1865, N1859, N393);
xor XOR2 (N1866, N1854, N329);
not NOT1 (N1867, N1852);
not NOT1 (N1868, N1866);
xor XOR2 (N1869, N1864, N1204);
not NOT1 (N1870, N1860);
not NOT1 (N1871, N1867);
not NOT1 (N1872, N1858);
xor XOR2 (N1873, N1839, N1362);
not NOT1 (N1874, N1873);
not NOT1 (N1875, N1850);
not NOT1 (N1876, N1875);
nand NAND2 (N1877, N1856, N657);
or OR3 (N1878, N1861, N639, N515);
not NOT1 (N1879, N1878);
not NOT1 (N1880, N1879);
nand NAND3 (N1881, N1871, N627, N1715);
not NOT1 (N1882, N1872);
not NOT1 (N1883, N1869);
nand NAND4 (N1884, N1868, N1028, N687, N1583);
buf BUF1 (N1885, N1884);
and AND4 (N1886, N1880, N1046, N925, N99);
nand NAND4 (N1887, N1883, N166, N860, N14);
nor NOR3 (N1888, N1865, N360, N183);
not NOT1 (N1889, N1881);
nand NAND3 (N1890, N1876, N1197, N1271);
and AND3 (N1891, N1874, N1352, N641);
xor XOR2 (N1892, N1870, N356);
not NOT1 (N1893, N1890);
nor NOR2 (N1894, N1886, N608);
not NOT1 (N1895, N1891);
nor NOR2 (N1896, N1892, N1377);
not NOT1 (N1897, N1887);
or OR4 (N1898, N1893, N1690, N1576, N670);
or OR2 (N1899, N1895, N66);
buf BUF1 (N1900, N1885);
or OR3 (N1901, N1897, N925, N1210);
and AND4 (N1902, N1882, N13, N190, N1144);
or OR2 (N1903, N1899, N1490);
nor NOR3 (N1904, N1877, N1053, N1535);
nand NAND3 (N1905, N1904, N244, N1015);
nor NOR4 (N1906, N1903, N935, N928, N633);
and AND3 (N1907, N1889, N80, N120);
and AND4 (N1908, N1888, N1327, N90, N176);
not NOT1 (N1909, N1906);
or OR2 (N1910, N1908, N1278);
not NOT1 (N1911, N1896);
and AND4 (N1912, N1909, N1308, N1831, N663);
xor XOR2 (N1913, N1902, N1345);
or OR3 (N1914, N1898, N1195, N49);
not NOT1 (N1915, N1910);
buf BUF1 (N1916, N1901);
not NOT1 (N1917, N1912);
nand NAND2 (N1918, N1914, N870);
not NOT1 (N1919, N1894);
nor NOR3 (N1920, N1915, N1479, N957);
nor NOR3 (N1921, N1905, N1713, N1582);
or OR2 (N1922, N1920, N1273);
nor NOR2 (N1923, N1913, N1794);
or OR2 (N1924, N1919, N1719);
nand NAND2 (N1925, N1918, N67);
not NOT1 (N1926, N1924);
not NOT1 (N1927, N1917);
xor XOR2 (N1928, N1907, N148);
buf BUF1 (N1929, N1923);
nor NOR4 (N1930, N1921, N340, N1811, N741);
or OR2 (N1931, N1928, N257);
nand NAND2 (N1932, N1922, N3);
xor XOR2 (N1933, N1931, N113);
nor NOR4 (N1934, N1927, N1279, N1736, N777);
buf BUF1 (N1935, N1911);
or OR3 (N1936, N1935, N95, N230);
buf BUF1 (N1937, N1916);
nand NAND2 (N1938, N1934, N278);
xor XOR2 (N1939, N1938, N496);
xor XOR2 (N1940, N1925, N1916);
buf BUF1 (N1941, N1926);
not NOT1 (N1942, N1936);
not NOT1 (N1943, N1900);
and AND4 (N1944, N1932, N527, N552, N938);
nor NOR2 (N1945, N1940, N1450);
nand NAND4 (N1946, N1933, N1900, N1017, N1940);
nand NAND3 (N1947, N1929, N1554, N1345);
and AND3 (N1948, N1947, N1174, N1360);
buf BUF1 (N1949, N1939);
nor NOR4 (N1950, N1937, N124, N555, N56);
nand NAND4 (N1951, N1941, N252, N1183, N1315);
buf BUF1 (N1952, N1949);
xor XOR2 (N1953, N1944, N613);
or OR2 (N1954, N1950, N1758);
nand NAND4 (N1955, N1943, N1713, N612, N582);
buf BUF1 (N1956, N1955);
buf BUF1 (N1957, N1946);
not NOT1 (N1958, N1953);
or OR2 (N1959, N1954, N1607);
nor NOR3 (N1960, N1945, N979, N186);
or OR3 (N1961, N1930, N707, N294);
and AND4 (N1962, N1952, N1052, N118, N1135);
buf BUF1 (N1963, N1962);
buf BUF1 (N1964, N1956);
nor NOR3 (N1965, N1948, N184, N1889);
nor NOR4 (N1966, N1964, N1620, N94, N1064);
or OR2 (N1967, N1957, N310);
xor XOR2 (N1968, N1942, N565);
not NOT1 (N1969, N1961);
or OR2 (N1970, N1958, N624);
or OR2 (N1971, N1970, N1749);
or OR3 (N1972, N1951, N385, N1721);
buf BUF1 (N1973, N1971);
or OR2 (N1974, N1968, N573);
buf BUF1 (N1975, N1965);
not NOT1 (N1976, N1959);
nand NAND2 (N1977, N1966, N572);
not NOT1 (N1978, N1976);
and AND3 (N1979, N1969, N1165, N1812);
not NOT1 (N1980, N1977);
and AND4 (N1981, N1980, N400, N1828, N1397);
xor XOR2 (N1982, N1978, N1214);
nor NOR4 (N1983, N1967, N1671, N1175, N395);
buf BUF1 (N1984, N1960);
nor NOR4 (N1985, N1979, N830, N1117, N1779);
nand NAND3 (N1986, N1963, N193, N281);
nor NOR2 (N1987, N1983, N1642);
not NOT1 (N1988, N1972);
or OR3 (N1989, N1987, N1963, N1097);
nor NOR2 (N1990, N1985, N769);
not NOT1 (N1991, N1988);
and AND3 (N1992, N1981, N1113, N1477);
nand NAND3 (N1993, N1986, N1614, N449);
nand NAND4 (N1994, N1989, N1230, N1087, N1488);
nor NOR4 (N1995, N1984, N937, N1167, N755);
nor NOR3 (N1996, N1982, N217, N175);
or OR3 (N1997, N1974, N1434, N131);
buf BUF1 (N1998, N1990);
not NOT1 (N1999, N1973);
nor NOR4 (N2000, N1975, N843, N1963, N1647);
buf BUF1 (N2001, N1991);
xor XOR2 (N2002, N1993, N123);
buf BUF1 (N2003, N1995);
xor XOR2 (N2004, N1998, N493);
and AND2 (N2005, N2003, N986);
not NOT1 (N2006, N1999);
xor XOR2 (N2007, N2001, N1590);
or OR2 (N2008, N2006, N861);
and AND2 (N2009, N1992, N483);
xor XOR2 (N2010, N2000, N1460);
nand NAND4 (N2011, N2008, N51, N1237, N1553);
and AND3 (N2012, N2009, N1277, N43);
nor NOR2 (N2013, N2005, N1756);
not NOT1 (N2014, N1996);
buf BUF1 (N2015, N2010);
nor NOR2 (N2016, N2015, N1218);
not NOT1 (N2017, N2004);
nor NOR2 (N2018, N2014, N910);
nor NOR2 (N2019, N2007, N536);
and AND3 (N2020, N2002, N424, N1244);
nor NOR4 (N2021, N2016, N1252, N1097, N1007);
xor XOR2 (N2022, N2013, N1257);
nor NOR4 (N2023, N2011, N1173, N1249, N1629);
or OR2 (N2024, N2021, N910);
nand NAND3 (N2025, N2020, N1568, N933);
xor XOR2 (N2026, N2018, N748);
xor XOR2 (N2027, N2017, N1351);
buf BUF1 (N2028, N2019);
not NOT1 (N2029, N2027);
buf BUF1 (N2030, N1994);
or OR3 (N2031, N2024, N312, N1387);
not NOT1 (N2032, N2029);
not NOT1 (N2033, N2031);
xor XOR2 (N2034, N2025, N189);
buf BUF1 (N2035, N2034);
buf BUF1 (N2036, N1997);
or OR2 (N2037, N2036, N77);
buf BUF1 (N2038, N2026);
and AND2 (N2039, N2012, N903);
nor NOR2 (N2040, N2022, N1121);
and AND2 (N2041, N2023, N1429);
xor XOR2 (N2042, N2040, N728);
or OR3 (N2043, N2038, N253, N464);
or OR2 (N2044, N2033, N277);
and AND4 (N2045, N2041, N631, N685, N1739);
or OR4 (N2046, N2028, N1881, N1452, N107);
not NOT1 (N2047, N2039);
xor XOR2 (N2048, N2030, N901);
buf BUF1 (N2049, N2037);
buf BUF1 (N2050, N2047);
and AND2 (N2051, N2045, N398);
and AND2 (N2052, N2048, N1824);
or OR2 (N2053, N2050, N794);
xor XOR2 (N2054, N2052, N940);
and AND2 (N2055, N2054, N1490);
not NOT1 (N2056, N2044);
nand NAND4 (N2057, N2055, N36, N774, N157);
nand NAND4 (N2058, N2051, N1971, N496, N1172);
buf BUF1 (N2059, N2043);
and AND2 (N2060, N2049, N1009);
nor NOR4 (N2061, N2057, N498, N580, N1945);
xor XOR2 (N2062, N2053, N959);
not NOT1 (N2063, N2042);
not NOT1 (N2064, N2062);
nor NOR3 (N2065, N2058, N1795, N1024);
nor NOR3 (N2066, N2032, N1233, N355);
nand NAND4 (N2067, N2066, N1791, N1803, N604);
nor NOR2 (N2068, N2056, N56);
nor NOR2 (N2069, N2035, N1130);
xor XOR2 (N2070, N2065, N996);
xor XOR2 (N2071, N2063, N1238);
or OR3 (N2072, N2071, N1620, N515);
buf BUF1 (N2073, N2064);
and AND3 (N2074, N2072, N803, N833);
not NOT1 (N2075, N2046);
xor XOR2 (N2076, N2067, N252);
and AND2 (N2077, N2060, N1095);
or OR4 (N2078, N2061, N1648, N1804, N1366);
buf BUF1 (N2079, N2069);
nor NOR4 (N2080, N2068, N1730, N294, N1366);
nor NOR4 (N2081, N2080, N1979, N1291, N738);
buf BUF1 (N2082, N2074);
xor XOR2 (N2083, N2079, N855);
and AND3 (N2084, N2076, N1513, N1687);
not NOT1 (N2085, N2070);
xor XOR2 (N2086, N2078, N1477);
not NOT1 (N2087, N2082);
buf BUF1 (N2088, N2075);
nand NAND3 (N2089, N2088, N248, N663);
and AND2 (N2090, N2059, N1729);
and AND2 (N2091, N2083, N1619);
nand NAND2 (N2092, N2090, N1283);
xor XOR2 (N2093, N2086, N77);
not NOT1 (N2094, N2091);
buf BUF1 (N2095, N2084);
nor NOR3 (N2096, N2093, N1395, N1770);
nand NAND2 (N2097, N2077, N1195);
buf BUF1 (N2098, N2087);
nand NAND3 (N2099, N2073, N469, N479);
nor NOR3 (N2100, N2085, N2043, N1192);
or OR2 (N2101, N2097, N749);
xor XOR2 (N2102, N2089, N656);
xor XOR2 (N2103, N2081, N1676);
nand NAND4 (N2104, N2100, N2077, N768, N485);
nor NOR4 (N2105, N2092, N503, N487, N1893);
nand NAND3 (N2106, N2095, N1547, N1738);
buf BUF1 (N2107, N2096);
and AND3 (N2108, N2099, N47, N1729);
or OR4 (N2109, N2106, N428, N887, N2106);
nor NOR2 (N2110, N2102, N1598);
xor XOR2 (N2111, N2109, N1376);
buf BUF1 (N2112, N2105);
not NOT1 (N2113, N2103);
and AND3 (N2114, N2112, N606, N1947);
nor NOR2 (N2115, N2101, N229);
or OR3 (N2116, N2113, N233, N1088);
nor NOR3 (N2117, N2114, N615, N526);
or OR3 (N2118, N2104, N1522, N31);
buf BUF1 (N2119, N2117);
not NOT1 (N2120, N2107);
nand NAND2 (N2121, N2111, N1436);
not NOT1 (N2122, N2098);
and AND2 (N2123, N2108, N181);
or OR3 (N2124, N2115, N551, N1928);
xor XOR2 (N2125, N2124, N2070);
xor XOR2 (N2126, N2116, N1103);
not NOT1 (N2127, N2121);
xor XOR2 (N2128, N2094, N919);
not NOT1 (N2129, N2126);
buf BUF1 (N2130, N2122);
buf BUF1 (N2131, N2130);
or OR4 (N2132, N2125, N753, N952, N1774);
nor NOR4 (N2133, N2110, N844, N1777, N1298);
not NOT1 (N2134, N2128);
or OR3 (N2135, N2127, N1548, N929);
xor XOR2 (N2136, N2134, N540);
buf BUF1 (N2137, N2133);
nand NAND2 (N2138, N2123, N1688);
nand NAND4 (N2139, N2137, N1828, N1989, N1754);
xor XOR2 (N2140, N2132, N187);
nor NOR2 (N2141, N2136, N54);
or OR4 (N2142, N2135, N1839, N1597, N2140);
nand NAND3 (N2143, N1330, N1508, N1633);
or OR3 (N2144, N2129, N546, N1674);
buf BUF1 (N2145, N2144);
or OR2 (N2146, N2131, N2025);
not NOT1 (N2147, N2139);
not NOT1 (N2148, N2119);
xor XOR2 (N2149, N2147, N1732);
buf BUF1 (N2150, N2141);
not NOT1 (N2151, N2120);
nor NOR4 (N2152, N2145, N1161, N178, N590);
buf BUF1 (N2153, N2151);
not NOT1 (N2154, N2149);
buf BUF1 (N2155, N2148);
nand NAND4 (N2156, N2118, N640, N1406, N2137);
buf BUF1 (N2157, N2154);
nor NOR3 (N2158, N2143, N324, N429);
buf BUF1 (N2159, N2156);
nor NOR3 (N2160, N2159, N273, N504);
or OR3 (N2161, N2155, N1666, N579);
buf BUF1 (N2162, N2160);
or OR3 (N2163, N2161, N563, N1648);
or OR3 (N2164, N2153, N812, N717);
buf BUF1 (N2165, N2146);
and AND2 (N2166, N2158, N1105);
nor NOR4 (N2167, N2138, N406, N1569, N2084);
not NOT1 (N2168, N2157);
nand NAND4 (N2169, N2152, N1479, N944, N1483);
or OR4 (N2170, N2167, N117, N1190, N640);
buf BUF1 (N2171, N2162);
buf BUF1 (N2172, N2171);
nor NOR3 (N2173, N2172, N1312, N441);
and AND4 (N2174, N2163, N1139, N494, N454);
nor NOR2 (N2175, N2173, N374);
xor XOR2 (N2176, N2168, N55);
xor XOR2 (N2177, N2176, N691);
nor NOR4 (N2178, N2166, N1349, N255, N381);
and AND2 (N2179, N2164, N1710);
or OR4 (N2180, N2170, N810, N1736, N695);
not NOT1 (N2181, N2180);
xor XOR2 (N2182, N2174, N779);
nor NOR2 (N2183, N2181, N888);
or OR2 (N2184, N2178, N1597);
and AND3 (N2185, N2177, N1772, N1844);
nand NAND2 (N2186, N2150, N2094);
and AND2 (N2187, N2185, N1032);
and AND2 (N2188, N2187, N1685);
not NOT1 (N2189, N2182);
not NOT1 (N2190, N2184);
xor XOR2 (N2191, N2142, N345);
nand NAND3 (N2192, N2183, N367, N2158);
xor XOR2 (N2193, N2179, N1317);
buf BUF1 (N2194, N2169);
and AND2 (N2195, N2165, N1245);
and AND2 (N2196, N2186, N1098);
nor NOR2 (N2197, N2191, N1084);
nor NOR3 (N2198, N2190, N221, N1010);
buf BUF1 (N2199, N2196);
not NOT1 (N2200, N2197);
or OR2 (N2201, N2175, N1164);
nand NAND2 (N2202, N2189, N1667);
buf BUF1 (N2203, N2195);
xor XOR2 (N2204, N2188, N751);
and AND4 (N2205, N2199, N1732, N1123, N2059);
buf BUF1 (N2206, N2198);
buf BUF1 (N2207, N2202);
and AND3 (N2208, N2192, N1912, N41);
xor XOR2 (N2209, N2193, N1950);
not NOT1 (N2210, N2208);
nand NAND4 (N2211, N2210, N297, N693, N963);
nor NOR4 (N2212, N2206, N1133, N807, N2014);
nand NAND2 (N2213, N2207, N2212);
nor NOR3 (N2214, N1158, N391, N835);
or OR2 (N2215, N2213, N2070);
xor XOR2 (N2216, N2209, N1238);
buf BUF1 (N2217, N2200);
not NOT1 (N2218, N2211);
and AND2 (N2219, N2214, N1474);
not NOT1 (N2220, N2194);
and AND3 (N2221, N2218, N1974, N1215);
buf BUF1 (N2222, N2219);
nor NOR2 (N2223, N2220, N954);
buf BUF1 (N2224, N2217);
nand NAND4 (N2225, N2204, N250, N1035, N216);
and AND4 (N2226, N2224, N1906, N911, N687);
and AND3 (N2227, N2215, N1004, N1418);
xor XOR2 (N2228, N2226, N626);
buf BUF1 (N2229, N2223);
or OR2 (N2230, N2221, N1140);
and AND2 (N2231, N2201, N103);
nor NOR2 (N2232, N2203, N1960);
not NOT1 (N2233, N2229);
buf BUF1 (N2234, N2233);
or OR2 (N2235, N2234, N6);
buf BUF1 (N2236, N2227);
buf BUF1 (N2237, N2228);
and AND2 (N2238, N2222, N2072);
buf BUF1 (N2239, N2238);
buf BUF1 (N2240, N2236);
or OR2 (N2241, N2205, N2175);
not NOT1 (N2242, N2237);
nand NAND2 (N2243, N2239, N2175);
nor NOR4 (N2244, N2231, N1945, N915, N2040);
or OR3 (N2245, N2240, N1972, N1422);
buf BUF1 (N2246, N2244);
xor XOR2 (N2247, N2230, N1477);
or OR3 (N2248, N2243, N1358, N1048);
and AND3 (N2249, N2242, N632, N1490);
nand NAND3 (N2250, N2216, N948, N493);
and AND2 (N2251, N2245, N522);
nor NOR4 (N2252, N2232, N1883, N1570, N239);
and AND2 (N2253, N2247, N1899);
nand NAND4 (N2254, N2249, N483, N1606, N810);
not NOT1 (N2255, N2235);
not NOT1 (N2256, N2250);
xor XOR2 (N2257, N2241, N2031);
and AND3 (N2258, N2255, N1327, N675);
and AND4 (N2259, N2253, N1352, N1200, N1739);
or OR2 (N2260, N2258, N1807);
not NOT1 (N2261, N2260);
buf BUF1 (N2262, N2246);
not NOT1 (N2263, N2225);
not NOT1 (N2264, N2251);
and AND4 (N2265, N2254, N125, N712, N876);
nand NAND2 (N2266, N2263, N1718);
nand NAND4 (N2267, N2257, N2067, N1634, N1145);
nand NAND2 (N2268, N2252, N531);
buf BUF1 (N2269, N2256);
and AND4 (N2270, N2268, N94, N766, N170);
buf BUF1 (N2271, N2266);
and AND2 (N2272, N2261, N1481);
buf BUF1 (N2273, N2265);
not NOT1 (N2274, N2264);
nand NAND2 (N2275, N2269, N471);
and AND2 (N2276, N2267, N923);
or OR3 (N2277, N2276, N290, N1679);
or OR3 (N2278, N2277, N632, N897);
nor NOR2 (N2279, N2248, N1365);
or OR2 (N2280, N2272, N1915);
or OR2 (N2281, N2270, N46);
or OR4 (N2282, N2278, N134, N1686, N1732);
nand NAND4 (N2283, N2279, N413, N1488, N482);
nor NOR3 (N2284, N2275, N1192, N642);
or OR4 (N2285, N2283, N219, N2149, N831);
nor NOR2 (N2286, N2271, N352);
buf BUF1 (N2287, N2281);
buf BUF1 (N2288, N2285);
xor XOR2 (N2289, N2284, N843);
or OR3 (N2290, N2282, N646, N607);
and AND3 (N2291, N2287, N1387, N458);
xor XOR2 (N2292, N2259, N1261);
buf BUF1 (N2293, N2291);
or OR2 (N2294, N2262, N874);
nor NOR4 (N2295, N2273, N1973, N624, N905);
nor NOR3 (N2296, N2274, N1866, N1781);
nor NOR4 (N2297, N2288, N1307, N1132, N581);
nor NOR4 (N2298, N2292, N653, N1385, N531);
or OR2 (N2299, N2298, N127);
nor NOR2 (N2300, N2289, N332);
xor XOR2 (N2301, N2295, N1837);
not NOT1 (N2302, N2290);
not NOT1 (N2303, N2301);
and AND3 (N2304, N2297, N1331, N834);
and AND2 (N2305, N2294, N1890);
buf BUF1 (N2306, N2296);
and AND2 (N2307, N2299, N366);
or OR4 (N2308, N2307, N1257, N2057, N98);
xor XOR2 (N2309, N2303, N2305);
xor XOR2 (N2310, N2094, N1169);
not NOT1 (N2311, N2286);
xor XOR2 (N2312, N2311, N1379);
nor NOR2 (N2313, N2302, N889);
or OR3 (N2314, N2300, N630, N240);
or OR2 (N2315, N2280, N1632);
nand NAND4 (N2316, N2315, N1901, N1501, N1971);
or OR2 (N2317, N2313, N2069);
nand NAND4 (N2318, N2316, N1048, N1955, N2232);
nand NAND4 (N2319, N2309, N973, N847, N55);
nor NOR3 (N2320, N2314, N1871, N815);
buf BUF1 (N2321, N2319);
nand NAND4 (N2322, N2293, N2071, N1651, N1715);
and AND2 (N2323, N2318, N1597);
nor NOR2 (N2324, N2312, N1764);
not NOT1 (N2325, N2322);
nand NAND3 (N2326, N2304, N1505, N1835);
nand NAND2 (N2327, N2320, N2159);
and AND4 (N2328, N2321, N1957, N1591, N694);
nor NOR3 (N2329, N2328, N623, N563);
or OR4 (N2330, N2323, N312, N1635, N27);
buf BUF1 (N2331, N2330);
xor XOR2 (N2332, N2306, N536);
and AND4 (N2333, N2332, N294, N653, N904);
buf BUF1 (N2334, N2329);
buf BUF1 (N2335, N2331);
or OR4 (N2336, N2334, N597, N2331, N598);
or OR3 (N2337, N2317, N138, N2182);
and AND2 (N2338, N2336, N1445);
nand NAND4 (N2339, N2335, N1254, N1772, N1727);
not NOT1 (N2340, N2327);
xor XOR2 (N2341, N2339, N1154);
nor NOR2 (N2342, N2340, N1185);
not NOT1 (N2343, N2310);
or OR4 (N2344, N2338, N271, N444, N151);
and AND3 (N2345, N2343, N1331, N1154);
not NOT1 (N2346, N2308);
not NOT1 (N2347, N2324);
nor NOR4 (N2348, N2325, N429, N344, N498);
nor NOR2 (N2349, N2341, N1769);
or OR2 (N2350, N2333, N450);
nor NOR2 (N2351, N2345, N2240);
xor XOR2 (N2352, N2342, N305);
xor XOR2 (N2353, N2349, N1793);
nand NAND3 (N2354, N2348, N1196, N859);
not NOT1 (N2355, N2354);
nor NOR2 (N2356, N2353, N148);
xor XOR2 (N2357, N2356, N575);
or OR3 (N2358, N2344, N1774, N216);
nor NOR4 (N2359, N2358, N2148, N953, N1449);
nor NOR4 (N2360, N2351, N1795, N1445, N1212);
or OR3 (N2361, N2326, N95, N1139);
and AND4 (N2362, N2346, N2277, N2090, N2074);
or OR3 (N2363, N2355, N1451, N544);
not NOT1 (N2364, N2359);
and AND2 (N2365, N2352, N1172);
nor NOR3 (N2366, N2361, N1925, N750);
not NOT1 (N2367, N2357);
or OR4 (N2368, N2362, N1398, N1940, N1771);
xor XOR2 (N2369, N2363, N693);
or OR3 (N2370, N2337, N926, N136);
nand NAND2 (N2371, N2370, N1864);
buf BUF1 (N2372, N2347);
xor XOR2 (N2373, N2365, N2362);
xor XOR2 (N2374, N2364, N1305);
xor XOR2 (N2375, N2371, N990);
xor XOR2 (N2376, N2373, N459);
or OR3 (N2377, N2367, N937, N1495);
and AND4 (N2378, N2375, N285, N1631, N1240);
not NOT1 (N2379, N2377);
not NOT1 (N2380, N2378);
and AND2 (N2381, N2379, N1137);
xor XOR2 (N2382, N2374, N924);
nand NAND3 (N2383, N2369, N559, N357);
or OR4 (N2384, N2381, N1275, N720, N1052);
xor XOR2 (N2385, N2382, N1591);
not NOT1 (N2386, N2360);
nand NAND3 (N2387, N2376, N173, N874);
and AND2 (N2388, N2368, N1356);
and AND3 (N2389, N2388, N48, N264);
xor XOR2 (N2390, N2366, N744);
buf BUF1 (N2391, N2350);
xor XOR2 (N2392, N2390, N1669);
xor XOR2 (N2393, N2389, N440);
not NOT1 (N2394, N2391);
not NOT1 (N2395, N2393);
nand NAND4 (N2396, N2383, N1016, N735, N1372);
or OR4 (N2397, N2392, N1838, N71, N771);
nand NAND2 (N2398, N2397, N2243);
or OR2 (N2399, N2398, N873);
or OR3 (N2400, N2395, N220, N20);
or OR3 (N2401, N2385, N196, N1318);
not NOT1 (N2402, N2394);
buf BUF1 (N2403, N2372);
or OR3 (N2404, N2384, N2042, N1322);
or OR4 (N2405, N2386, N533, N518, N963);
nor NOR3 (N2406, N2380, N284, N1311);
nand NAND2 (N2407, N2402, N629);
or OR2 (N2408, N2400, N2214);
or OR4 (N2409, N2404, N622, N1337, N931);
nand NAND2 (N2410, N2409, N490);
nor NOR4 (N2411, N2405, N1755, N2228, N1868);
buf BUF1 (N2412, N2403);
or OR4 (N2413, N2401, N906, N889, N8);
nor NOR4 (N2414, N2411, N585, N1254, N1472);
buf BUF1 (N2415, N2408);
xor XOR2 (N2416, N2399, N1630);
xor XOR2 (N2417, N2414, N78);
buf BUF1 (N2418, N2416);
buf BUF1 (N2419, N2413);
or OR2 (N2420, N2396, N234);
and AND4 (N2421, N2412, N1188, N1269, N1890);
nand NAND3 (N2422, N2421, N1563, N304);
and AND2 (N2423, N2406, N950);
or OR3 (N2424, N2387, N1838, N326);
not NOT1 (N2425, N2418);
or OR3 (N2426, N2422, N1697, N2328);
not NOT1 (N2427, N2424);
and AND3 (N2428, N2425, N1589, N1517);
nor NOR2 (N2429, N2428, N494);
or OR2 (N2430, N2427, N269);
buf BUF1 (N2431, N2415);
nand NAND4 (N2432, N2423, N517, N862, N1900);
nor NOR2 (N2433, N2407, N1689);
xor XOR2 (N2434, N2420, N1164);
nor NOR4 (N2435, N2429, N2273, N1206, N1073);
nand NAND4 (N2436, N2417, N846, N1593, N217);
or OR3 (N2437, N2419, N627, N447);
or OR3 (N2438, N2431, N368, N2211);
nor NOR2 (N2439, N2426, N569);
not NOT1 (N2440, N2437);
nand NAND2 (N2441, N2430, N746);
nand NAND3 (N2442, N2436, N1099, N863);
not NOT1 (N2443, N2441);
buf BUF1 (N2444, N2443);
buf BUF1 (N2445, N2438);
and AND4 (N2446, N2442, N2415, N511, N1222);
buf BUF1 (N2447, N2410);
nand NAND3 (N2448, N2432, N1431, N1061);
xor XOR2 (N2449, N2439, N1323);
or OR4 (N2450, N2433, N1031, N2349, N1048);
xor XOR2 (N2451, N2448, N496);
or OR4 (N2452, N2445, N728, N413, N705);
or OR3 (N2453, N2434, N898, N1155);
nand NAND4 (N2454, N2440, N791, N1087, N1092);
not NOT1 (N2455, N2454);
xor XOR2 (N2456, N2449, N1381);
buf BUF1 (N2457, N2444);
xor XOR2 (N2458, N2435, N1596);
nand NAND4 (N2459, N2457, N2403, N1972, N1606);
or OR2 (N2460, N2447, N2195);
not NOT1 (N2461, N2459);
xor XOR2 (N2462, N2461, N158);
or OR4 (N2463, N2462, N2208, N507, N198);
buf BUF1 (N2464, N2456);
xor XOR2 (N2465, N2460, N31);
xor XOR2 (N2466, N2450, N457);
xor XOR2 (N2467, N2455, N2293);
nand NAND4 (N2468, N2463, N1273, N676, N1958);
nor NOR4 (N2469, N2465, N712, N2017, N1482);
and AND3 (N2470, N2446, N201, N193);
and AND2 (N2471, N2468, N1896);
nor NOR3 (N2472, N2470, N2427, N2455);
or OR4 (N2473, N2458, N1445, N748, N1920);
or OR2 (N2474, N2469, N611);
or OR4 (N2475, N2474, N275, N1168, N2439);
nand NAND3 (N2476, N2472, N850, N583);
or OR3 (N2477, N2452, N435, N499);
or OR4 (N2478, N2467, N573, N946, N2378);
xor XOR2 (N2479, N2464, N2072);
xor XOR2 (N2480, N2479, N1080);
buf BUF1 (N2481, N2478);
buf BUF1 (N2482, N2475);
or OR4 (N2483, N2451, N1235, N2046, N672);
xor XOR2 (N2484, N2476, N1256);
not NOT1 (N2485, N2473);
buf BUF1 (N2486, N2483);
and AND4 (N2487, N2471, N1124, N1794, N2021);
not NOT1 (N2488, N2484);
or OR4 (N2489, N2486, N268, N244, N102);
nor NOR3 (N2490, N2466, N1967, N1935);
nor NOR4 (N2491, N2488, N455, N25, N1091);
xor XOR2 (N2492, N2489, N502);
buf BUF1 (N2493, N2487);
or OR2 (N2494, N2493, N1574);
nor NOR4 (N2495, N2490, N2453, N421, N1166);
not NOT1 (N2496, N2254);
xor XOR2 (N2497, N2480, N27);
nand NAND4 (N2498, N2482, N344, N432, N2464);
or OR4 (N2499, N2491, N1050, N755, N815);
and AND2 (N2500, N2497, N200);
or OR3 (N2501, N2499, N2006, N493);
nand NAND3 (N2502, N2485, N1438, N599);
or OR2 (N2503, N2477, N1717);
nand NAND2 (N2504, N2494, N1716);
nor NOR4 (N2505, N2496, N717, N1145, N2210);
nor NOR2 (N2506, N2501, N1908);
nor NOR2 (N2507, N2500, N293);
not NOT1 (N2508, N2502);
nor NOR4 (N2509, N2498, N701, N2166, N1248);
nand NAND2 (N2510, N2495, N1764);
nand NAND2 (N2511, N2509, N2125);
buf BUF1 (N2512, N2503);
nand NAND4 (N2513, N2506, N90, N1442, N23);
and AND2 (N2514, N2481, N2353);
nand NAND4 (N2515, N2508, N2497, N1939, N1984);
and AND2 (N2516, N2512, N830);
and AND3 (N2517, N2515, N2313, N938);
not NOT1 (N2518, N2516);
buf BUF1 (N2519, N2517);
xor XOR2 (N2520, N2518, N177);
nor NOR2 (N2521, N2510, N2044);
buf BUF1 (N2522, N2513);
nor NOR3 (N2523, N2507, N155, N1754);
and AND4 (N2524, N2511, N335, N845, N623);
not NOT1 (N2525, N2521);
or OR2 (N2526, N2514, N812);
nand NAND4 (N2527, N2504, N1355, N841, N926);
nand NAND2 (N2528, N2519, N2132);
nor NOR4 (N2529, N2523, N1692, N1179, N75);
nor NOR2 (N2530, N2505, N167);
and AND4 (N2531, N2530, N1253, N769, N69);
or OR2 (N2532, N2526, N735);
buf BUF1 (N2533, N2492);
nor NOR2 (N2534, N2532, N1846);
buf BUF1 (N2535, N2524);
nor NOR4 (N2536, N2525, N1192, N1650, N1089);
and AND3 (N2537, N2529, N1771, N138);
xor XOR2 (N2538, N2531, N2282);
and AND2 (N2539, N2537, N2529);
and AND2 (N2540, N2534, N2534);
nor NOR2 (N2541, N2540, N1437);
buf BUF1 (N2542, N2535);
or OR2 (N2543, N2522, N1745);
or OR3 (N2544, N2527, N1875, N582);
not NOT1 (N2545, N2543);
nor NOR4 (N2546, N2533, N1528, N873, N1511);
buf BUF1 (N2547, N2528);
and AND4 (N2548, N2542, N1307, N939, N1493);
buf BUF1 (N2549, N2548);
not NOT1 (N2550, N2546);
xor XOR2 (N2551, N2544, N2053);
not NOT1 (N2552, N2538);
xor XOR2 (N2553, N2547, N2240);
buf BUF1 (N2554, N2551);
xor XOR2 (N2555, N2554, N888);
and AND3 (N2556, N2549, N438, N190);
xor XOR2 (N2557, N2536, N799);
and AND2 (N2558, N2550, N12);
and AND4 (N2559, N2545, N335, N1263, N654);
and AND3 (N2560, N2553, N1419, N1601);
nor NOR2 (N2561, N2559, N1888);
buf BUF1 (N2562, N2561);
and AND2 (N2563, N2558, N556);
nor NOR3 (N2564, N2563, N1627, N788);
xor XOR2 (N2565, N2541, N1489);
nor NOR2 (N2566, N2520, N868);
buf BUF1 (N2567, N2562);
nor NOR2 (N2568, N2566, N480);
xor XOR2 (N2569, N2560, N89);
and AND3 (N2570, N2568, N1230, N1972);
xor XOR2 (N2571, N2556, N1468);
nor NOR3 (N2572, N2555, N1930, N1409);
not NOT1 (N2573, N2571);
nor NOR4 (N2574, N2557, N1019, N1839, N1609);
xor XOR2 (N2575, N2564, N2499);
nand NAND4 (N2576, N2567, N1667, N649, N2527);
nand NAND3 (N2577, N2576, N1178, N1556);
not NOT1 (N2578, N2572);
and AND2 (N2579, N2569, N562);
not NOT1 (N2580, N2579);
buf BUF1 (N2581, N2580);
nor NOR2 (N2582, N2581, N2246);
nand NAND4 (N2583, N2573, N1812, N937, N1144);
nor NOR4 (N2584, N2565, N2359, N995, N971);
nand NAND2 (N2585, N2574, N2357);
nand NAND2 (N2586, N2539, N1988);
nor NOR3 (N2587, N2577, N2157, N7);
not NOT1 (N2588, N2585);
and AND2 (N2589, N2584, N2356);
nand NAND4 (N2590, N2589, N587, N2445, N1960);
nand NAND4 (N2591, N2590, N86, N1744, N1010);
buf BUF1 (N2592, N2570);
nor NOR2 (N2593, N2552, N1649);
and AND3 (N2594, N2578, N1062, N840);
not NOT1 (N2595, N2594);
not NOT1 (N2596, N2592);
not NOT1 (N2597, N2583);
nor NOR2 (N2598, N2591, N178);
nand NAND4 (N2599, N2582, N234, N935, N1647);
or OR3 (N2600, N2596, N1980, N167);
or OR2 (N2601, N2586, N930);
not NOT1 (N2602, N2588);
nor NOR4 (N2603, N2602, N1965, N712, N2158);
buf BUF1 (N2604, N2598);
or OR2 (N2605, N2587, N2325);
and AND3 (N2606, N2597, N1493, N208);
nor NOR2 (N2607, N2599, N166);
and AND3 (N2608, N2605, N1739, N1531);
and AND4 (N2609, N2600, N169, N451, N1766);
xor XOR2 (N2610, N2607, N100);
buf BUF1 (N2611, N2603);
xor XOR2 (N2612, N2606, N258);
or OR3 (N2613, N2595, N2187, N2537);
xor XOR2 (N2614, N2593, N2516);
and AND4 (N2615, N2612, N453, N1954, N1248);
buf BUF1 (N2616, N2610);
xor XOR2 (N2617, N2601, N607);
buf BUF1 (N2618, N2609);
and AND3 (N2619, N2575, N1392, N131);
xor XOR2 (N2620, N2614, N1617);
xor XOR2 (N2621, N2615, N480);
not NOT1 (N2622, N2619);
nand NAND2 (N2623, N2617, N2167);
nand NAND2 (N2624, N2613, N2567);
xor XOR2 (N2625, N2623, N1591);
or OR4 (N2626, N2624, N1830, N633, N723);
xor XOR2 (N2627, N2621, N618);
not NOT1 (N2628, N2611);
and AND4 (N2629, N2604, N1379, N1533, N503);
or OR4 (N2630, N2608, N858, N1909, N2378);
xor XOR2 (N2631, N2628, N1003);
not NOT1 (N2632, N2626);
xor XOR2 (N2633, N2629, N1298);
or OR3 (N2634, N2620, N1509, N2629);
xor XOR2 (N2635, N2618, N1937);
not NOT1 (N2636, N2616);
nand NAND4 (N2637, N2635, N837, N1016, N2528);
xor XOR2 (N2638, N2637, N1008);
nor NOR3 (N2639, N2630, N51, N1947);
and AND2 (N2640, N2627, N1878);
buf BUF1 (N2641, N2622);
or OR4 (N2642, N2625, N734, N892, N817);
xor XOR2 (N2643, N2632, N847);
nor NOR3 (N2644, N2640, N938, N1039);
nor NOR3 (N2645, N2636, N2235, N2545);
nand NAND3 (N2646, N2634, N609, N1016);
nor NOR3 (N2647, N2642, N752, N1156);
xor XOR2 (N2648, N2647, N649);
and AND2 (N2649, N2639, N1792);
or OR4 (N2650, N2644, N1379, N183, N1852);
and AND4 (N2651, N2641, N394, N1062, N805);
and AND3 (N2652, N2648, N491, N745);
nor NOR2 (N2653, N2651, N816);
buf BUF1 (N2654, N2643);
nand NAND2 (N2655, N2633, N1216);
buf BUF1 (N2656, N2652);
or OR3 (N2657, N2655, N1097, N294);
nor NOR2 (N2658, N2649, N1613);
nor NOR4 (N2659, N2645, N962, N995, N2403);
or OR2 (N2660, N2654, N2087);
buf BUF1 (N2661, N2659);
and AND3 (N2662, N2661, N2100, N1321);
buf BUF1 (N2663, N2631);
buf BUF1 (N2664, N2663);
xor XOR2 (N2665, N2658, N290);
or OR4 (N2666, N2662, N994, N290, N1619);
not NOT1 (N2667, N2665);
nor NOR4 (N2668, N2667, N1368, N280, N1806);
nor NOR2 (N2669, N2646, N2605);
not NOT1 (N2670, N2638);
nand NAND4 (N2671, N2668, N643, N1137, N697);
xor XOR2 (N2672, N2653, N2200);
buf BUF1 (N2673, N2670);
xor XOR2 (N2674, N2657, N797);
not NOT1 (N2675, N2666);
and AND2 (N2676, N2660, N277);
or OR4 (N2677, N2656, N1546, N1978, N2522);
nand NAND4 (N2678, N2674, N1683, N1684, N1573);
nand NAND3 (N2679, N2650, N1621, N714);
buf BUF1 (N2680, N2675);
nor NOR4 (N2681, N2676, N647, N2555, N2212);
xor XOR2 (N2682, N2679, N1025);
nand NAND3 (N2683, N2673, N2640, N1110);
nor NOR2 (N2684, N2681, N2294);
not NOT1 (N2685, N2672);
nor NOR3 (N2686, N2664, N583, N317);
nor NOR4 (N2687, N2680, N2384, N721, N543);
nand NAND2 (N2688, N2677, N393);
and AND3 (N2689, N2678, N2285, N2073);
not NOT1 (N2690, N2671);
or OR2 (N2691, N2685, N918);
nor NOR2 (N2692, N2690, N856);
buf BUF1 (N2693, N2684);
buf BUF1 (N2694, N2669);
buf BUF1 (N2695, N2692);
not NOT1 (N2696, N2689);
nand NAND3 (N2697, N2695, N1026, N2676);
nor NOR3 (N2698, N2696, N412, N72);
not NOT1 (N2699, N2683);
or OR2 (N2700, N2688, N1895);
and AND2 (N2701, N2700, N474);
and AND4 (N2702, N2686, N1801, N463, N547);
and AND2 (N2703, N2691, N2569);
nor NOR2 (N2704, N2702, N1077);
not NOT1 (N2705, N2694);
nand NAND3 (N2706, N2697, N481, N1605);
nor NOR4 (N2707, N2703, N1938, N2583, N2215);
xor XOR2 (N2708, N2701, N2052);
buf BUF1 (N2709, N2707);
buf BUF1 (N2710, N2698);
xor XOR2 (N2711, N2687, N341);
buf BUF1 (N2712, N2710);
and AND4 (N2713, N2708, N1735, N1946, N1328);
xor XOR2 (N2714, N2711, N2065);
nand NAND2 (N2715, N2699, N1089);
nand NAND4 (N2716, N2693, N1721, N452, N960);
xor XOR2 (N2717, N2709, N2112);
nor NOR3 (N2718, N2706, N1875, N1034);
not NOT1 (N2719, N2718);
nor NOR4 (N2720, N2682, N1119, N1756, N2257);
and AND4 (N2721, N2714, N1142, N897, N1718);
xor XOR2 (N2722, N2704, N710);
buf BUF1 (N2723, N2722);
not NOT1 (N2724, N2716);
buf BUF1 (N2725, N2721);
not NOT1 (N2726, N2719);
and AND3 (N2727, N2705, N1221, N123);
nor NOR3 (N2728, N2724, N1158, N1443);
not NOT1 (N2729, N2728);
buf BUF1 (N2730, N2713);
or OR4 (N2731, N2729, N2588, N69, N2682);
xor XOR2 (N2732, N2726, N1270);
and AND3 (N2733, N2727, N2165, N395);
nor NOR4 (N2734, N2712, N793, N2133, N1661);
xor XOR2 (N2735, N2715, N2525);
not NOT1 (N2736, N2735);
and AND2 (N2737, N2731, N1448);
or OR3 (N2738, N2720, N1413, N1700);
not NOT1 (N2739, N2737);
xor XOR2 (N2740, N2725, N502);
buf BUF1 (N2741, N2734);
and AND2 (N2742, N2733, N2176);
and AND3 (N2743, N2730, N323, N957);
xor XOR2 (N2744, N2740, N1541);
or OR4 (N2745, N2723, N1420, N2168, N1770);
not NOT1 (N2746, N2732);
not NOT1 (N2747, N2739);
or OR2 (N2748, N2738, N312);
xor XOR2 (N2749, N2748, N2365);
xor XOR2 (N2750, N2747, N1379);
nand NAND3 (N2751, N2742, N2722, N1956);
nand NAND4 (N2752, N2745, N1730, N1236, N634);
and AND2 (N2753, N2752, N1355);
nand NAND4 (N2754, N2744, N603, N511, N1160);
not NOT1 (N2755, N2746);
or OR2 (N2756, N2753, N194);
xor XOR2 (N2757, N2741, N134);
or OR3 (N2758, N2757, N1749, N1271);
and AND3 (N2759, N2717, N246, N2559);
and AND4 (N2760, N2754, N1265, N115, N2359);
nor NOR4 (N2761, N2756, N1452, N1934, N1556);
and AND4 (N2762, N2759, N963, N2636, N1918);
xor XOR2 (N2763, N2755, N2417);
and AND3 (N2764, N2763, N80, N1818);
and AND2 (N2765, N2764, N1994);
nor NOR4 (N2766, N2760, N468, N1430, N1675);
buf BUF1 (N2767, N2743);
and AND2 (N2768, N2750, N2044);
nand NAND4 (N2769, N2751, N847, N1909, N1132);
and AND2 (N2770, N2767, N753);
or OR2 (N2771, N2736, N1616);
xor XOR2 (N2772, N2769, N1052);
or OR2 (N2773, N2761, N63);
or OR4 (N2774, N2766, N859, N464, N1589);
nand NAND2 (N2775, N2768, N2625);
buf BUF1 (N2776, N2758);
not NOT1 (N2777, N2765);
not NOT1 (N2778, N2771);
or OR4 (N2779, N2772, N1081, N434, N2390);
buf BUF1 (N2780, N2773);
xor XOR2 (N2781, N2774, N2681);
nor NOR4 (N2782, N2776, N1972, N405, N42);
or OR3 (N2783, N2778, N884, N379);
nor NOR3 (N2784, N2781, N2476, N725);
nand NAND4 (N2785, N2783, N1777, N348, N2101);
nor NOR2 (N2786, N2775, N1581);
not NOT1 (N2787, N2782);
nand NAND3 (N2788, N2762, N498, N174);
xor XOR2 (N2789, N2770, N68);
or OR2 (N2790, N2749, N698);
nor NOR2 (N2791, N2780, N1270);
nor NOR4 (N2792, N2787, N600, N335, N1370);
buf BUF1 (N2793, N2791);
nand NAND3 (N2794, N2789, N2545, N2391);
and AND4 (N2795, N2792, N2621, N1813, N1032);
nor NOR2 (N2796, N2790, N887);
nand NAND3 (N2797, N2794, N2672, N1739);
nand NAND2 (N2798, N2784, N22);
not NOT1 (N2799, N2788);
not NOT1 (N2800, N2777);
nand NAND3 (N2801, N2785, N2567, N1532);
nor NOR2 (N2802, N2799, N1230);
nor NOR3 (N2803, N2793, N780, N1797);
not NOT1 (N2804, N2798);
nand NAND3 (N2805, N2800, N2611, N716);
nor NOR2 (N2806, N2804, N472);
nand NAND2 (N2807, N2803, N1956);
xor XOR2 (N2808, N2805, N556);
buf BUF1 (N2809, N2801);
and AND4 (N2810, N2797, N1198, N2144, N1828);
and AND4 (N2811, N2779, N2585, N1588, N995);
and AND3 (N2812, N2811, N393, N853);
nand NAND2 (N2813, N2807, N384);
xor XOR2 (N2814, N2808, N112);
xor XOR2 (N2815, N2812, N1059);
nand NAND4 (N2816, N2796, N1039, N236, N2492);
not NOT1 (N2817, N2816);
buf BUF1 (N2818, N2813);
nor NOR2 (N2819, N2810, N2211);
and AND2 (N2820, N2786, N1113);
buf BUF1 (N2821, N2802);
nand NAND3 (N2822, N2809, N1171, N390);
and AND4 (N2823, N2815, N492, N1833, N2217);
or OR4 (N2824, N2822, N117, N1912, N2656);
buf BUF1 (N2825, N2820);
not NOT1 (N2826, N2814);
or OR3 (N2827, N2825, N908, N1141);
buf BUF1 (N2828, N2827);
buf BUF1 (N2829, N2819);
not NOT1 (N2830, N2828);
nand NAND4 (N2831, N2823, N2564, N1118, N122);
and AND3 (N2832, N2795, N300, N145);
nor NOR3 (N2833, N2832, N2729, N1434);
nor NOR3 (N2834, N2830, N2535, N746);
not NOT1 (N2835, N2826);
nand NAND2 (N2836, N2817, N2471);
nand NAND4 (N2837, N2821, N2148, N552, N2340);
nand NAND3 (N2838, N2806, N1690, N891);
buf BUF1 (N2839, N2836);
buf BUF1 (N2840, N2838);
not NOT1 (N2841, N2834);
nand NAND4 (N2842, N2833, N1661, N1466, N2038);
nor NOR4 (N2843, N2835, N1859, N2805, N2801);
nand NAND4 (N2844, N2837, N2007, N2302, N389);
not NOT1 (N2845, N2844);
buf BUF1 (N2846, N2843);
not NOT1 (N2847, N2831);
or OR2 (N2848, N2842, N1750);
nor NOR3 (N2849, N2845, N1707, N1598);
nor NOR4 (N2850, N2839, N2688, N1065, N2475);
xor XOR2 (N2851, N2850, N2112);
not NOT1 (N2852, N2847);
nor NOR4 (N2853, N2840, N683, N2799, N86);
not NOT1 (N2854, N2849);
not NOT1 (N2855, N2848);
buf BUF1 (N2856, N2852);
xor XOR2 (N2857, N2851, N2551);
or OR4 (N2858, N2853, N1660, N2791, N722);
not NOT1 (N2859, N2858);
or OR3 (N2860, N2829, N166, N2157);
and AND4 (N2861, N2841, N261, N2746, N462);
nor NOR3 (N2862, N2855, N148, N1327);
not NOT1 (N2863, N2824);
buf BUF1 (N2864, N2862);
buf BUF1 (N2865, N2854);
or OR2 (N2866, N2860, N876);
not NOT1 (N2867, N2846);
nand NAND4 (N2868, N2867, N904, N1120, N2019);
nand NAND2 (N2869, N2864, N1224);
and AND4 (N2870, N2866, N2357, N1281, N1479);
not NOT1 (N2871, N2857);
or OR3 (N2872, N2856, N2344, N1549);
nor NOR3 (N2873, N2863, N2683, N276);
nand NAND4 (N2874, N2872, N1983, N1096, N279);
nor NOR4 (N2875, N2861, N2198, N454, N564);
not NOT1 (N2876, N2868);
and AND2 (N2877, N2873, N575);
xor XOR2 (N2878, N2871, N2271);
nor NOR4 (N2879, N2859, N798, N1776, N2552);
nand NAND4 (N2880, N2879, N1671, N191, N403);
nor NOR3 (N2881, N2865, N315, N2120);
xor XOR2 (N2882, N2881, N1149);
buf BUF1 (N2883, N2877);
xor XOR2 (N2884, N2876, N145);
nor NOR3 (N2885, N2869, N2718, N210);
not NOT1 (N2886, N2874);
nor NOR3 (N2887, N2880, N1788, N187);
nand NAND3 (N2888, N2818, N1607, N2855);
nor NOR2 (N2889, N2888, N218);
nand NAND4 (N2890, N2875, N1571, N2563, N2673);
not NOT1 (N2891, N2884);
xor XOR2 (N2892, N2885, N829);
xor XOR2 (N2893, N2870, N2145);
not NOT1 (N2894, N2889);
and AND4 (N2895, N2892, N277, N2499, N2167);
nor NOR4 (N2896, N2893, N2442, N132, N591);
and AND3 (N2897, N2896, N1861, N2409);
nand NAND3 (N2898, N2890, N1199, N2132);
not NOT1 (N2899, N2894);
xor XOR2 (N2900, N2878, N732);
not NOT1 (N2901, N2895);
nor NOR2 (N2902, N2899, N352);
and AND3 (N2903, N2901, N2187, N1807);
or OR4 (N2904, N2886, N2577, N2743, N875);
nor NOR3 (N2905, N2900, N2820, N1144);
nor NOR2 (N2906, N2905, N1393);
nor NOR3 (N2907, N2891, N2316, N1912);
nor NOR3 (N2908, N2903, N1448, N1978);
or OR4 (N2909, N2902, N1430, N518, N2248);
xor XOR2 (N2910, N2898, N1523);
not NOT1 (N2911, N2906);
or OR4 (N2912, N2907, N542, N2117, N752);
buf BUF1 (N2913, N2908);
buf BUF1 (N2914, N2883);
and AND2 (N2915, N2911, N2822);
not NOT1 (N2916, N2882);
nand NAND3 (N2917, N2909, N1224, N210);
nand NAND2 (N2918, N2914, N2278);
or OR3 (N2919, N2897, N1157, N1778);
nand NAND3 (N2920, N2904, N1777, N193);
xor XOR2 (N2921, N2910, N396);
nor NOR4 (N2922, N2916, N1798, N2649, N2439);
or OR3 (N2923, N2917, N261, N623);
nor NOR3 (N2924, N2887, N208, N592);
buf BUF1 (N2925, N2919);
nor NOR3 (N2926, N2915, N1783, N1833);
nor NOR3 (N2927, N2918, N2116, N1062);
xor XOR2 (N2928, N2921, N1213);
nor NOR2 (N2929, N2920, N1278);
nand NAND3 (N2930, N2913, N1848, N1783);
not NOT1 (N2931, N2925);
buf BUF1 (N2932, N2926);
xor XOR2 (N2933, N2932, N2749);
xor XOR2 (N2934, N2931, N2339);
not NOT1 (N2935, N2930);
xor XOR2 (N2936, N2924, N2415);
or OR2 (N2937, N2929, N657);
nand NAND4 (N2938, N2933, N2145, N837, N128);
and AND3 (N2939, N2927, N1578, N48);
nand NAND3 (N2940, N2935, N9, N1273);
and AND3 (N2941, N2928, N2126, N2432);
xor XOR2 (N2942, N2940, N2904);
and AND2 (N2943, N2934, N574);
nor NOR2 (N2944, N2943, N1137);
not NOT1 (N2945, N2938);
xor XOR2 (N2946, N2912, N365);
buf BUF1 (N2947, N2945);
and AND2 (N2948, N2922, N2233);
and AND4 (N2949, N2948, N45, N1876, N2309);
or OR3 (N2950, N2936, N2222, N1069);
xor XOR2 (N2951, N2939, N215);
nand NAND3 (N2952, N2947, N2928, N786);
and AND2 (N2953, N2949, N1454);
or OR4 (N2954, N2946, N276, N681, N641);
or OR3 (N2955, N2951, N1862, N1346);
or OR4 (N2956, N2955, N2789, N2441, N1507);
not NOT1 (N2957, N2952);
and AND3 (N2958, N2953, N440, N2143);
xor XOR2 (N2959, N2954, N67);
not NOT1 (N2960, N2950);
xor XOR2 (N2961, N2941, N899);
nor NOR2 (N2962, N2956, N2473);
xor XOR2 (N2963, N2960, N659);
buf BUF1 (N2964, N2923);
xor XOR2 (N2965, N2962, N835);
or OR2 (N2966, N2963, N1565);
not NOT1 (N2967, N2957);
not NOT1 (N2968, N2961);
nand NAND3 (N2969, N2959, N934, N2638);
buf BUF1 (N2970, N2965);
nand NAND4 (N2971, N2966, N2317, N2948, N117);
buf BUF1 (N2972, N2937);
xor XOR2 (N2973, N2944, N1092);
nand NAND4 (N2974, N2967, N974, N1912, N2026);
and AND3 (N2975, N2970, N2711, N2523);
not NOT1 (N2976, N2968);
and AND3 (N2977, N2972, N2078, N613);
nor NOR3 (N2978, N2942, N2912, N1302);
not NOT1 (N2979, N2971);
nor NOR3 (N2980, N2975, N861, N2887);
nand NAND4 (N2981, N2976, N602, N990, N811);
nand NAND4 (N2982, N2978, N152, N1566, N2410);
nand NAND3 (N2983, N2958, N103, N2511);
buf BUF1 (N2984, N2981);
nor NOR4 (N2985, N2983, N563, N819, N126);
and AND3 (N2986, N2979, N2456, N1224);
nor NOR4 (N2987, N2974, N12, N564, N2068);
nor NOR2 (N2988, N2964, N2318);
not NOT1 (N2989, N2985);
xor XOR2 (N2990, N2984, N2385);
and AND3 (N2991, N2973, N1820, N1573);
not NOT1 (N2992, N2969);
not NOT1 (N2993, N2988);
buf BUF1 (N2994, N2982);
or OR3 (N2995, N2993, N1402, N297);
buf BUF1 (N2996, N2995);
nor NOR2 (N2997, N2991, N2625);
xor XOR2 (N2998, N2989, N2637);
and AND3 (N2999, N2987, N2182, N180);
or OR4 (N3000, N2980, N1956, N1029, N451);
xor XOR2 (N3001, N2999, N227);
or OR3 (N3002, N2994, N144, N895);
buf BUF1 (N3003, N2992);
nor NOR2 (N3004, N2986, N989);
buf BUF1 (N3005, N3001);
nor NOR2 (N3006, N2998, N195);
and AND4 (N3007, N2977, N2109, N248, N1782);
xor XOR2 (N3008, N3002, N1894);
and AND3 (N3009, N3006, N2550, N1852);
or OR3 (N3010, N2990, N1530, N2566);
nor NOR3 (N3011, N2996, N2424, N2920);
nor NOR4 (N3012, N3009, N2598, N1571, N1976);
not NOT1 (N3013, N3003);
not NOT1 (N3014, N3011);
and AND2 (N3015, N3013, N1000);
buf BUF1 (N3016, N3000);
buf BUF1 (N3017, N3005);
not NOT1 (N3018, N3007);
nor NOR3 (N3019, N3014, N91, N1352);
and AND4 (N3020, N3019, N2095, N1547, N1853);
xor XOR2 (N3021, N3012, N270);
buf BUF1 (N3022, N3010);
not NOT1 (N3023, N3022);
nor NOR3 (N3024, N3021, N2135, N2104);
nor NOR3 (N3025, N3016, N2071, N2668);
and AND4 (N3026, N3004, N913, N2013, N1652);
and AND4 (N3027, N3017, N2469, N1117, N2904);
and AND2 (N3028, N3018, N495);
nand NAND2 (N3029, N3020, N1632);
or OR4 (N3030, N3029, N1666, N2410, N540);
nor NOR2 (N3031, N2997, N2425);
and AND3 (N3032, N3026, N814, N1618);
not NOT1 (N3033, N3032);
nand NAND2 (N3034, N3008, N913);
and AND2 (N3035, N3025, N456);
and AND3 (N3036, N3024, N3035, N2639);
xor XOR2 (N3037, N953, N2413);
or OR4 (N3038, N3027, N1374, N428, N2387);
xor XOR2 (N3039, N3037, N1081);
buf BUF1 (N3040, N3039);
nand NAND4 (N3041, N3033, N1491, N254, N2765);
nor NOR2 (N3042, N3030, N2757);
nand NAND4 (N3043, N3034, N1266, N2672, N786);
nor NOR4 (N3044, N3038, N656, N1337, N2219);
not NOT1 (N3045, N3043);
nor NOR2 (N3046, N3042, N446);
nor NOR4 (N3047, N3015, N2079, N2085, N737);
and AND3 (N3048, N3041, N2799, N2733);
xor XOR2 (N3049, N3040, N2455);
and AND2 (N3050, N3047, N764);
nor NOR2 (N3051, N3028, N2900);
and AND3 (N3052, N3044, N299, N526);
nor NOR4 (N3053, N3050, N3050, N1396, N1790);
xor XOR2 (N3054, N3031, N375);
nor NOR2 (N3055, N3051, N1208);
or OR3 (N3056, N3036, N2654, N2545);
or OR4 (N3057, N3045, N605, N565, N830);
or OR2 (N3058, N3052, N1052);
nor NOR3 (N3059, N3055, N2007, N2909);
xor XOR2 (N3060, N3049, N1869);
xor XOR2 (N3061, N3056, N967);
or OR3 (N3062, N3048, N1779, N374);
and AND4 (N3063, N3060, N2919, N2814, N601);
buf BUF1 (N3064, N3061);
and AND2 (N3065, N3057, N2432);
nor NOR3 (N3066, N3023, N2233, N1556);
not NOT1 (N3067, N3053);
and AND4 (N3068, N3046, N772, N591, N2581);
xor XOR2 (N3069, N3063, N2852);
xor XOR2 (N3070, N3054, N787);
buf BUF1 (N3071, N3064);
nand NAND4 (N3072, N3071, N158, N43, N2168);
nor NOR3 (N3073, N3067, N388, N1172);
or OR4 (N3074, N3062, N512, N540, N309);
or OR3 (N3075, N3072, N500, N2980);
buf BUF1 (N3076, N3075);
xor XOR2 (N3077, N3074, N2552);
nor NOR2 (N3078, N3073, N2276);
not NOT1 (N3079, N3070);
nor NOR4 (N3080, N3068, N634, N226, N2013);
nor NOR3 (N3081, N3065, N1445, N278);
not NOT1 (N3082, N3059);
and AND4 (N3083, N3081, N1137, N2474, N985);
or OR3 (N3084, N3082, N219, N2540);
nor NOR4 (N3085, N3076, N1957, N1742, N1405);
nand NAND3 (N3086, N3083, N13, N2226);
nor NOR4 (N3087, N3077, N745, N2322, N1530);
xor XOR2 (N3088, N3086, N2521);
not NOT1 (N3089, N3087);
not NOT1 (N3090, N3069);
or OR4 (N3091, N3090, N1431, N3037, N2027);
nor NOR2 (N3092, N3079, N2804);
buf BUF1 (N3093, N3089);
or OR2 (N3094, N3088, N482);
or OR4 (N3095, N3078, N1939, N2524, N930);
buf BUF1 (N3096, N3080);
buf BUF1 (N3097, N3095);
xor XOR2 (N3098, N3092, N852);
and AND3 (N3099, N3085, N2863, N820);
buf BUF1 (N3100, N3096);
nor NOR4 (N3101, N3100, N411, N1712, N700);
xor XOR2 (N3102, N3094, N1037);
nor NOR4 (N3103, N3093, N2951, N1865, N1517);
not NOT1 (N3104, N3084);
xor XOR2 (N3105, N3098, N2495);
nor NOR4 (N3106, N3066, N1425, N310, N534);
buf BUF1 (N3107, N3105);
not NOT1 (N3108, N3103);
or OR4 (N3109, N3108, N2823, N1169, N1065);
not NOT1 (N3110, N3091);
nor NOR3 (N3111, N3109, N452, N1300);
nand NAND2 (N3112, N3111, N2460);
not NOT1 (N3113, N3106);
buf BUF1 (N3114, N3113);
and AND3 (N3115, N3107, N1736, N1381);
xor XOR2 (N3116, N3114, N1689);
nand NAND2 (N3117, N3099, N270);
nand NAND2 (N3118, N3101, N2808);
nor NOR4 (N3119, N3117, N1547, N2003, N963);
buf BUF1 (N3120, N3116);
or OR3 (N3121, N3058, N778, N1082);
buf BUF1 (N3122, N3110);
xor XOR2 (N3123, N3118, N2683);
and AND3 (N3124, N3122, N649, N1943);
not NOT1 (N3125, N3124);
nand NAND2 (N3126, N3102, N2707);
or OR4 (N3127, N3115, N2116, N2440, N777);
not NOT1 (N3128, N3120);
or OR2 (N3129, N3128, N2259);
or OR2 (N3130, N3126, N4);
not NOT1 (N3131, N3097);
xor XOR2 (N3132, N3112, N1209);
and AND2 (N3133, N3121, N3045);
nand NAND2 (N3134, N3130, N1800);
xor XOR2 (N3135, N3127, N2166);
buf BUF1 (N3136, N3131);
nor NOR3 (N3137, N3125, N154, N200);
not NOT1 (N3138, N3135);
xor XOR2 (N3139, N3119, N1012);
nor NOR2 (N3140, N3138, N1185);
and AND2 (N3141, N3133, N508);
nor NOR4 (N3142, N3136, N456, N1473, N440);
nand NAND2 (N3143, N3137, N2018);
and AND4 (N3144, N3140, N1541, N566, N2376);
nand NAND2 (N3145, N3129, N756);
nand NAND4 (N3146, N3144, N3008, N2161, N1910);
or OR2 (N3147, N3123, N1017);
nor NOR3 (N3148, N3145, N2023, N1343);
buf BUF1 (N3149, N3139);
not NOT1 (N3150, N3149);
not NOT1 (N3151, N3147);
and AND4 (N3152, N3143, N53, N1498, N305);
xor XOR2 (N3153, N3152, N246);
nor NOR3 (N3154, N3153, N3140, N748);
buf BUF1 (N3155, N3154);
or OR4 (N3156, N3155, N788, N1893, N115);
xor XOR2 (N3157, N3104, N1542);
or OR4 (N3158, N3151, N2858, N319, N1953);
buf BUF1 (N3159, N3146);
or OR3 (N3160, N3158, N412, N320);
or OR3 (N3161, N3142, N2081, N1368);
and AND3 (N3162, N3156, N986, N1330);
and AND3 (N3163, N3134, N1588, N1620);
and AND4 (N3164, N3159, N956, N972, N3048);
not NOT1 (N3165, N3141);
xor XOR2 (N3166, N3164, N933);
not NOT1 (N3167, N3150);
xor XOR2 (N3168, N3161, N2104);
buf BUF1 (N3169, N3160);
nand NAND2 (N3170, N3169, N1375);
buf BUF1 (N3171, N3132);
buf BUF1 (N3172, N3148);
or OR3 (N3173, N3172, N1815, N542);
not NOT1 (N3174, N3157);
nand NAND2 (N3175, N3174, N1861);
nor NOR2 (N3176, N3162, N717);
and AND3 (N3177, N3175, N1895, N2444);
not NOT1 (N3178, N3167);
nand NAND4 (N3179, N3173, N2496, N1103, N2002);
xor XOR2 (N3180, N3168, N612);
buf BUF1 (N3181, N3170);
not NOT1 (N3182, N3171);
buf BUF1 (N3183, N3166);
and AND4 (N3184, N3182, N1090, N752, N2798);
not NOT1 (N3185, N3165);
and AND3 (N3186, N3176, N2233, N204);
and AND3 (N3187, N3186, N373, N451);
or OR4 (N3188, N3184, N1374, N391, N1549);
nor NOR3 (N3189, N3179, N1887, N1304);
or OR4 (N3190, N3188, N987, N1834, N1212);
nor NOR4 (N3191, N3180, N2514, N2372, N2193);
buf BUF1 (N3192, N3187);
and AND4 (N3193, N3192, N464, N166, N2605);
buf BUF1 (N3194, N3190);
or OR3 (N3195, N3185, N2884, N885);
nand NAND2 (N3196, N3193, N2479);
buf BUF1 (N3197, N3178);
not NOT1 (N3198, N3194);
nor NOR4 (N3199, N3177, N708, N1128, N1621);
buf BUF1 (N3200, N3181);
and AND3 (N3201, N3198, N2530, N2822);
nor NOR4 (N3202, N3163, N1176, N751, N2669);
not NOT1 (N3203, N3197);
nand NAND3 (N3204, N3189, N1677, N789);
buf BUF1 (N3205, N3200);
xor XOR2 (N3206, N3202, N348);
nand NAND2 (N3207, N3206, N2195);
and AND2 (N3208, N3196, N305);
xor XOR2 (N3209, N3205, N462);
or OR3 (N3210, N3204, N578, N109);
and AND3 (N3211, N3207, N517, N3039);
or OR2 (N3212, N3199, N2694);
nor NOR2 (N3213, N3201, N29);
nand NAND4 (N3214, N3183, N2057, N1193, N1381);
not NOT1 (N3215, N3203);
nor NOR2 (N3216, N3195, N2499);
or OR3 (N3217, N3213, N1034, N2772);
and AND2 (N3218, N3215, N207);
or OR3 (N3219, N3214, N1000, N1592);
not NOT1 (N3220, N3219);
xor XOR2 (N3221, N3210, N1597);
xor XOR2 (N3222, N3216, N2402);
xor XOR2 (N3223, N3212, N3140);
nor NOR3 (N3224, N3223, N1574, N1270);
not NOT1 (N3225, N3209);
buf BUF1 (N3226, N3191);
nand NAND2 (N3227, N3225, N429);
xor XOR2 (N3228, N3211, N2192);
buf BUF1 (N3229, N3217);
xor XOR2 (N3230, N3226, N1939);
buf BUF1 (N3231, N3208);
not NOT1 (N3232, N3220);
not NOT1 (N3233, N3231);
buf BUF1 (N3234, N3222);
xor XOR2 (N3235, N3234, N2713);
not NOT1 (N3236, N3221);
xor XOR2 (N3237, N3230, N2927);
nor NOR3 (N3238, N3237, N2532, N787);
or OR3 (N3239, N3224, N3190, N1515);
xor XOR2 (N3240, N3236, N1684);
nand NAND3 (N3241, N3240, N1856, N1155);
nand NAND2 (N3242, N3229, N213);
xor XOR2 (N3243, N3242, N1084);
buf BUF1 (N3244, N3241);
not NOT1 (N3245, N3227);
and AND2 (N3246, N3232, N548);
buf BUF1 (N3247, N3238);
xor XOR2 (N3248, N3247, N2782);
and AND2 (N3249, N3218, N59);
xor XOR2 (N3250, N3235, N1378);
nand NAND2 (N3251, N3244, N59);
nand NAND3 (N3252, N3249, N633, N1975);
not NOT1 (N3253, N3250);
nand NAND4 (N3254, N3253, N1048, N3125, N3040);
xor XOR2 (N3255, N3245, N3185);
nand NAND3 (N3256, N3252, N3090, N1253);
xor XOR2 (N3257, N3233, N1723);
not NOT1 (N3258, N3246);
buf BUF1 (N3259, N3255);
nor NOR4 (N3260, N3248, N1234, N298, N3223);
and AND3 (N3261, N3260, N1362, N277);
buf BUF1 (N3262, N3228);
nor NOR4 (N3263, N3254, N2871, N2669, N1683);
and AND4 (N3264, N3262, N3190, N1055, N2061);
not NOT1 (N3265, N3264);
nand NAND2 (N3266, N3257, N186);
or OR4 (N3267, N3243, N2984, N3171, N1690);
nand NAND3 (N3268, N3259, N1575, N3141);
nand NAND2 (N3269, N3251, N1451);
not NOT1 (N3270, N3263);
nor NOR2 (N3271, N3267, N1705);
not NOT1 (N3272, N3256);
nand NAND4 (N3273, N3265, N1814, N1799, N439);
xor XOR2 (N3274, N3269, N1317);
not NOT1 (N3275, N3258);
nand NAND3 (N3276, N3275, N1922, N2408);
nand NAND2 (N3277, N3271, N396);
not NOT1 (N3278, N3268);
not NOT1 (N3279, N3261);
or OR2 (N3280, N3278, N345);
buf BUF1 (N3281, N3277);
and AND3 (N3282, N3266, N3168, N625);
not NOT1 (N3283, N3276);
and AND4 (N3284, N3279, N733, N470, N2041);
buf BUF1 (N3285, N3281);
nand NAND2 (N3286, N3272, N1230);
or OR3 (N3287, N3270, N3245, N1241);
buf BUF1 (N3288, N3239);
buf BUF1 (N3289, N3274);
nor NOR4 (N3290, N3289, N119, N1667, N1357);
or OR3 (N3291, N3283, N2005, N1598);
nor NOR3 (N3292, N3286, N1094, N1840);
not NOT1 (N3293, N3292);
not NOT1 (N3294, N3290);
nor NOR2 (N3295, N3280, N554);
or OR2 (N3296, N3295, N133);
buf BUF1 (N3297, N3285);
not NOT1 (N3298, N3288);
and AND4 (N3299, N3273, N177, N2509, N1778);
nor NOR3 (N3300, N3298, N1394, N1193);
and AND4 (N3301, N3297, N1619, N2112, N1724);
xor XOR2 (N3302, N3296, N470);
or OR2 (N3303, N3301, N605);
nor NOR4 (N3304, N3302, N1117, N710, N102);
xor XOR2 (N3305, N3294, N439);
and AND2 (N3306, N3291, N2639);
nor NOR2 (N3307, N3304, N184);
not NOT1 (N3308, N3284);
or OR3 (N3309, N3306, N3284, N311);
not NOT1 (N3310, N3300);
and AND4 (N3311, N3309, N1137, N627, N3013);
or OR3 (N3312, N3303, N1050, N647);
xor XOR2 (N3313, N3308, N2342);
not NOT1 (N3314, N3299);
and AND2 (N3315, N3305, N2689);
nor NOR4 (N3316, N3282, N2383, N2350, N2423);
buf BUF1 (N3317, N3314);
not NOT1 (N3318, N3316);
not NOT1 (N3319, N3313);
nand NAND4 (N3320, N3293, N366, N598, N3053);
xor XOR2 (N3321, N3315, N1476);
nor NOR4 (N3322, N3307, N1292, N611, N1905);
not NOT1 (N3323, N3321);
or OR2 (N3324, N3311, N1091);
nor NOR2 (N3325, N3317, N649);
nor NOR4 (N3326, N3287, N1264, N14, N515);
and AND4 (N3327, N3322, N3289, N1700, N1293);
xor XOR2 (N3328, N3327, N1283);
not NOT1 (N3329, N3324);
nor NOR2 (N3330, N3319, N2563);
nor NOR3 (N3331, N3320, N806, N494);
and AND3 (N3332, N3326, N1841, N1389);
nand NAND4 (N3333, N3332, N1526, N1181, N1385);
buf BUF1 (N3334, N3312);
or OR2 (N3335, N3325, N3003);
and AND4 (N3336, N3328, N2835, N1034, N1667);
xor XOR2 (N3337, N3323, N163);
nand NAND2 (N3338, N3333, N2463);
not NOT1 (N3339, N3330);
xor XOR2 (N3340, N3331, N1773);
and AND4 (N3341, N3318, N2527, N3194, N3240);
xor XOR2 (N3342, N3341, N1534);
nor NOR3 (N3343, N3335, N2345, N2042);
nand NAND2 (N3344, N3343, N2043);
nand NAND2 (N3345, N3310, N1195);
not NOT1 (N3346, N3345);
nor NOR4 (N3347, N3336, N1160, N318, N389);
or OR2 (N3348, N3338, N784);
and AND3 (N3349, N3340, N2358, N2816);
xor XOR2 (N3350, N3342, N2320);
and AND2 (N3351, N3346, N1802);
or OR4 (N3352, N3349, N2130, N1309, N2607);
nand NAND3 (N3353, N3339, N3018, N3176);
xor XOR2 (N3354, N3347, N2643);
nand NAND2 (N3355, N3344, N1287);
xor XOR2 (N3356, N3348, N2317);
xor XOR2 (N3357, N3337, N40);
buf BUF1 (N3358, N3356);
and AND3 (N3359, N3353, N2203, N306);
and AND3 (N3360, N3350, N2473, N2645);
nor NOR4 (N3361, N3358, N489, N395, N1082);
or OR2 (N3362, N3355, N2622);
or OR2 (N3363, N3329, N298);
xor XOR2 (N3364, N3354, N1247);
or OR3 (N3365, N3363, N2534, N2469);
buf BUF1 (N3366, N3362);
and AND3 (N3367, N3361, N1274, N1654);
not NOT1 (N3368, N3357);
not NOT1 (N3369, N3364);
nor NOR4 (N3370, N3352, N42, N590, N1577);
buf BUF1 (N3371, N3365);
buf BUF1 (N3372, N3370);
xor XOR2 (N3373, N3360, N3141);
nand NAND2 (N3374, N3373, N478);
nand NAND3 (N3375, N3359, N1258, N2119);
and AND3 (N3376, N3351, N599, N870);
nand NAND2 (N3377, N3374, N2545);
nor NOR4 (N3378, N3377, N276, N1067, N1321);
or OR4 (N3379, N3334, N2236, N2362, N139);
and AND2 (N3380, N3371, N381);
not NOT1 (N3381, N3366);
nand NAND2 (N3382, N3367, N59);
nand NAND4 (N3383, N3382, N2413, N2642, N857);
or OR3 (N3384, N3379, N2071, N1266);
and AND3 (N3385, N3376, N2453, N1801);
and AND3 (N3386, N3384, N1043, N1915);
or OR2 (N3387, N3369, N2505);
or OR2 (N3388, N3387, N2919);
nand NAND4 (N3389, N3388, N3050, N158, N1337);
and AND4 (N3390, N3389, N3087, N2979, N322);
or OR3 (N3391, N3380, N3247, N372);
and AND3 (N3392, N3383, N340, N2001);
not NOT1 (N3393, N3375);
not NOT1 (N3394, N3386);
and AND2 (N3395, N3368, N467);
xor XOR2 (N3396, N3391, N1944);
nand NAND3 (N3397, N3372, N2614, N3327);
buf BUF1 (N3398, N3381);
and AND3 (N3399, N3378, N697, N1812);
buf BUF1 (N3400, N3392);
buf BUF1 (N3401, N3390);
nor NOR4 (N3402, N3395, N104, N2470, N152);
buf BUF1 (N3403, N3400);
nor NOR2 (N3404, N3403, N1186);
and AND2 (N3405, N3385, N2957);
buf BUF1 (N3406, N3404);
and AND3 (N3407, N3398, N1724, N2078);
buf BUF1 (N3408, N3401);
nor NOR2 (N3409, N3397, N2456);
and AND4 (N3410, N3408, N1369, N512, N1965);
not NOT1 (N3411, N3394);
nor NOR3 (N3412, N3411, N202, N342);
buf BUF1 (N3413, N3407);
nand NAND2 (N3414, N3413, N1539);
nor NOR4 (N3415, N3399, N3304, N2355, N1000);
xor XOR2 (N3416, N3410, N1842);
not NOT1 (N3417, N3415);
or OR2 (N3418, N3406, N1274);
not NOT1 (N3419, N3416);
and AND2 (N3420, N3402, N2525);
or OR3 (N3421, N3418, N730, N2631);
and AND2 (N3422, N3396, N1154);
or OR4 (N3423, N3405, N240, N2677, N1405);
nand NAND4 (N3424, N3422, N3392, N297, N2692);
buf BUF1 (N3425, N3409);
xor XOR2 (N3426, N3424, N3104);
nand NAND3 (N3427, N3414, N3150, N345);
nand NAND3 (N3428, N3426, N2067, N3052);
buf BUF1 (N3429, N3421);
and AND4 (N3430, N3419, N1368, N399, N700);
nand NAND4 (N3431, N3425, N2683, N1357, N2210);
not NOT1 (N3432, N3428);
not NOT1 (N3433, N3412);
not NOT1 (N3434, N3433);
nand NAND3 (N3435, N3434, N2739, N1603);
and AND3 (N3436, N3393, N1384, N1922);
not NOT1 (N3437, N3423);
xor XOR2 (N3438, N3420, N2356);
not NOT1 (N3439, N3427);
not NOT1 (N3440, N3436);
xor XOR2 (N3441, N3439, N1129);
nor NOR4 (N3442, N3430, N211, N80, N821);
and AND2 (N3443, N3432, N2117);
nand NAND2 (N3444, N3429, N145);
or OR3 (N3445, N3435, N232, N519);
not NOT1 (N3446, N3431);
nor NOR3 (N3447, N3442, N1583, N1097);
buf BUF1 (N3448, N3440);
xor XOR2 (N3449, N3444, N549);
xor XOR2 (N3450, N3448, N371);
and AND3 (N3451, N3445, N841, N3132);
nor NOR2 (N3452, N3447, N466);
nand NAND4 (N3453, N3446, N2299, N3118, N2816);
not NOT1 (N3454, N3417);
xor XOR2 (N3455, N3451, N2767);
buf BUF1 (N3456, N3455);
buf BUF1 (N3457, N3443);
buf BUF1 (N3458, N3449);
nand NAND3 (N3459, N3457, N950, N2990);
nor NOR4 (N3460, N3452, N533, N2790, N1836);
or OR4 (N3461, N3454, N502, N1027, N1157);
nor NOR4 (N3462, N3459, N1445, N2051, N2790);
or OR3 (N3463, N3441, N2215, N3131);
nand NAND3 (N3464, N3463, N523, N249);
buf BUF1 (N3465, N3453);
nor NOR4 (N3466, N3437, N2357, N2541, N1636);
nor NOR3 (N3467, N3450, N2846, N45);
and AND4 (N3468, N3466, N3127, N2605, N2692);
or OR2 (N3469, N3460, N559);
nand NAND4 (N3470, N3462, N2745, N224, N1947);
not NOT1 (N3471, N3464);
and AND3 (N3472, N3465, N3262, N2212);
buf BUF1 (N3473, N3471);
and AND4 (N3474, N3468, N729, N965, N495);
buf BUF1 (N3475, N3438);
not NOT1 (N3476, N3458);
or OR2 (N3477, N3472, N264);
not NOT1 (N3478, N3461);
nand NAND3 (N3479, N3476, N2269, N3053);
nand NAND3 (N3480, N3479, N216, N262);
or OR4 (N3481, N3477, N540, N910, N2853);
buf BUF1 (N3482, N3475);
and AND3 (N3483, N3473, N536, N1647);
and AND2 (N3484, N3481, N914);
nand NAND4 (N3485, N3469, N929, N2040, N2770);
buf BUF1 (N3486, N3474);
nand NAND4 (N3487, N3470, N921, N512, N550);
buf BUF1 (N3488, N3478);
or OR2 (N3489, N3487, N3161);
buf BUF1 (N3490, N3482);
and AND3 (N3491, N3467, N22, N2455);
nor NOR3 (N3492, N3483, N624, N2518);
not NOT1 (N3493, N3490);
nor NOR2 (N3494, N3488, N1240);
or OR3 (N3495, N3492, N933, N2544);
and AND2 (N3496, N3456, N488);
nand NAND4 (N3497, N3489, N2234, N648, N857);
or OR3 (N3498, N3494, N3193, N2806);
buf BUF1 (N3499, N3485);
and AND3 (N3500, N3486, N1053, N1966);
xor XOR2 (N3501, N3497, N3159);
xor XOR2 (N3502, N3495, N1466);
nand NAND2 (N3503, N3500, N2283);
buf BUF1 (N3504, N3491);
buf BUF1 (N3505, N3498);
xor XOR2 (N3506, N3504, N362);
not NOT1 (N3507, N3496);
nor NOR3 (N3508, N3480, N1726, N1506);
or OR2 (N3509, N3501, N3234);
nor NOR3 (N3510, N3509, N1854, N2210);
buf BUF1 (N3511, N3484);
not NOT1 (N3512, N3507);
or OR3 (N3513, N3508, N2650, N2023);
or OR2 (N3514, N3493, N23);
or OR3 (N3515, N3511, N1226, N1791);
nand NAND2 (N3516, N3515, N174);
nand NAND3 (N3517, N3502, N2403, N2732);
buf BUF1 (N3518, N3510);
or OR2 (N3519, N3514, N2386);
buf BUF1 (N3520, N3516);
and AND3 (N3521, N3519, N1440, N2215);
nor NOR2 (N3522, N3517, N2510);
nor NOR4 (N3523, N3522, N1891, N3320, N1717);
and AND4 (N3524, N3503, N2753, N3036, N1383);
nand NAND4 (N3525, N3512, N260, N469, N2882);
nand NAND2 (N3526, N3506, N2714);
nor NOR3 (N3527, N3499, N69, N79);
xor XOR2 (N3528, N3521, N2606);
not NOT1 (N3529, N3526);
or OR4 (N3530, N3524, N1243, N3364, N1810);
not NOT1 (N3531, N3520);
not NOT1 (N3532, N3531);
or OR4 (N3533, N3529, N17, N941, N45);
or OR3 (N3534, N3532, N3294, N3285);
nor NOR3 (N3535, N3523, N419, N2548);
or OR2 (N3536, N3528, N1620);
nand NAND2 (N3537, N3535, N1370);
not NOT1 (N3538, N3537);
or OR3 (N3539, N3505, N3048, N1586);
nor NOR4 (N3540, N3539, N923, N2220, N1155);
not NOT1 (N3541, N3536);
not NOT1 (N3542, N3534);
or OR2 (N3543, N3518, N2488);
and AND4 (N3544, N3540, N3288, N1737, N2487);
and AND4 (N3545, N3542, N3396, N869, N245);
nor NOR3 (N3546, N3533, N222, N925);
buf BUF1 (N3547, N3543);
nor NOR2 (N3548, N3525, N407);
and AND4 (N3549, N3538, N2422, N1817, N1032);
not NOT1 (N3550, N3548);
nor NOR2 (N3551, N3544, N1030);
buf BUF1 (N3552, N3549);
nand NAND4 (N3553, N3530, N2105, N3276, N2248);
nand NAND4 (N3554, N3513, N2355, N2355, N2294);
not NOT1 (N3555, N3547);
buf BUF1 (N3556, N3550);
xor XOR2 (N3557, N3553, N1600);
or OR4 (N3558, N3554, N884, N1122, N761);
and AND3 (N3559, N3545, N1057, N58);
and AND4 (N3560, N3555, N1914, N1189, N2333);
nand NAND4 (N3561, N3558, N1925, N2446, N2338);
xor XOR2 (N3562, N3552, N1330);
nand NAND2 (N3563, N3556, N2588);
and AND4 (N3564, N3560, N1323, N3050, N595);
buf BUF1 (N3565, N3551);
buf BUF1 (N3566, N3565);
or OR4 (N3567, N3566, N3118, N1941, N110);
nand NAND4 (N3568, N3563, N3114, N1015, N2165);
buf BUF1 (N3569, N3559);
xor XOR2 (N3570, N3546, N3285);
buf BUF1 (N3571, N3570);
buf BUF1 (N3572, N3527);
nor NOR3 (N3573, N3541, N2224, N3309);
nand NAND4 (N3574, N3562, N785, N2050, N873);
nand NAND2 (N3575, N3572, N73);
xor XOR2 (N3576, N3575, N3410);
nor NOR2 (N3577, N3569, N355);
nand NAND2 (N3578, N3573, N1515);
xor XOR2 (N3579, N3571, N1624);
and AND4 (N3580, N3564, N1845, N1522, N2300);
xor XOR2 (N3581, N3574, N2214);
or OR2 (N3582, N3579, N332);
not NOT1 (N3583, N3567);
or OR4 (N3584, N3561, N175, N1839, N1473);
not NOT1 (N3585, N3580);
not NOT1 (N3586, N3585);
nor NOR4 (N3587, N3583, N1422, N1733, N1862);
nor NOR4 (N3588, N3586, N2039, N1340, N3457);
nor NOR4 (N3589, N3577, N3196, N1981, N2267);
buf BUF1 (N3590, N3576);
or OR3 (N3591, N3587, N1768, N219);
and AND3 (N3592, N3568, N2142, N3471);
xor XOR2 (N3593, N3581, N735);
and AND4 (N3594, N3590, N37, N2523, N407);
not NOT1 (N3595, N3593);
nor NOR3 (N3596, N3584, N1984, N2549);
xor XOR2 (N3597, N3596, N1188);
and AND3 (N3598, N3589, N187, N1500);
or OR3 (N3599, N3588, N3171, N1080);
buf BUF1 (N3600, N3582);
xor XOR2 (N3601, N3600, N2423);
and AND2 (N3602, N3599, N2331);
not NOT1 (N3603, N3592);
not NOT1 (N3604, N3591);
or OR3 (N3605, N3594, N1100, N561);
not NOT1 (N3606, N3605);
nand NAND3 (N3607, N3598, N962, N1833);
and AND2 (N3608, N3604, N1053);
buf BUF1 (N3609, N3602);
and AND2 (N3610, N3603, N3269);
not NOT1 (N3611, N3609);
nor NOR4 (N3612, N3597, N3024, N3485, N667);
nor NOR4 (N3613, N3578, N500, N2147, N1824);
not NOT1 (N3614, N3607);
xor XOR2 (N3615, N3557, N650);
nand NAND2 (N3616, N3608, N2596);
and AND3 (N3617, N3616, N2426, N769);
buf BUF1 (N3618, N3606);
xor XOR2 (N3619, N3601, N2620);
buf BUF1 (N3620, N3612);
nand NAND2 (N3621, N3619, N380);
nor NOR3 (N3622, N3621, N950, N3592);
nand NAND2 (N3623, N3613, N2527);
not NOT1 (N3624, N3595);
or OR2 (N3625, N3620, N2718);
xor XOR2 (N3626, N3624, N2464);
nand NAND2 (N3627, N3626, N2156);
buf BUF1 (N3628, N3617);
and AND2 (N3629, N3611, N2484);
nor NOR4 (N3630, N3629, N2295, N2619, N1422);
nand NAND3 (N3631, N3630, N3366, N3465);
and AND4 (N3632, N3615, N699, N817, N2259);
and AND4 (N3633, N3622, N3059, N2550, N448);
buf BUF1 (N3634, N3623);
xor XOR2 (N3635, N3625, N2486);
not NOT1 (N3636, N3632);
or OR2 (N3637, N3628, N2847);
nor NOR4 (N3638, N3610, N842, N318, N674);
nor NOR3 (N3639, N3618, N1249, N51);
or OR3 (N3640, N3636, N939, N781);
nand NAND3 (N3641, N3635, N1510, N1216);
not NOT1 (N3642, N3614);
or OR3 (N3643, N3638, N2965, N2299);
and AND4 (N3644, N3641, N715, N3215, N3177);
not NOT1 (N3645, N3639);
or OR3 (N3646, N3640, N2866, N396);
not NOT1 (N3647, N3631);
xor XOR2 (N3648, N3646, N2046);
buf BUF1 (N3649, N3647);
buf BUF1 (N3650, N3648);
nand NAND3 (N3651, N3644, N531, N3301);
and AND4 (N3652, N3634, N1346, N2784, N645);
or OR2 (N3653, N3650, N2876);
xor XOR2 (N3654, N3643, N3340);
not NOT1 (N3655, N3637);
not NOT1 (N3656, N3645);
not NOT1 (N3657, N3652);
xor XOR2 (N3658, N3627, N2664);
nand NAND2 (N3659, N3651, N1668);
and AND2 (N3660, N3658, N1150);
xor XOR2 (N3661, N3656, N269);
nor NOR2 (N3662, N3661, N3613);
and AND4 (N3663, N3633, N2903, N3025, N312);
and AND2 (N3664, N3642, N2456);
or OR2 (N3665, N3653, N1486);
not NOT1 (N3666, N3660);
buf BUF1 (N3667, N3664);
nand NAND3 (N3668, N3662, N2954, N3021);
not NOT1 (N3669, N3657);
nand NAND4 (N3670, N3666, N3039, N2205, N1608);
not NOT1 (N3671, N3649);
and AND4 (N3672, N3665, N2653, N1906, N241);
nand NAND4 (N3673, N3668, N2959, N2165, N1650);
and AND2 (N3674, N3671, N858);
xor XOR2 (N3675, N3674, N1303);
buf BUF1 (N3676, N3675);
xor XOR2 (N3677, N3663, N597);
nor NOR3 (N3678, N3676, N3023, N1690);
buf BUF1 (N3679, N3672);
and AND3 (N3680, N3678, N2330, N3622);
buf BUF1 (N3681, N3669);
buf BUF1 (N3682, N3667);
nor NOR2 (N3683, N3673, N90);
and AND3 (N3684, N3683, N782, N1287);
not NOT1 (N3685, N3655);
not NOT1 (N3686, N3685);
nand NAND3 (N3687, N3679, N1109, N1405);
xor XOR2 (N3688, N3677, N895);
nand NAND3 (N3689, N3670, N750, N3604);
nor NOR3 (N3690, N3680, N3418, N2914);
xor XOR2 (N3691, N3687, N2738);
xor XOR2 (N3692, N3684, N1812);
not NOT1 (N3693, N3682);
buf BUF1 (N3694, N3654);
or OR3 (N3695, N3689, N459, N3105);
xor XOR2 (N3696, N3659, N60);
buf BUF1 (N3697, N3688);
nand NAND3 (N3698, N3686, N2520, N2445);
or OR2 (N3699, N3681, N1373);
xor XOR2 (N3700, N3691, N429);
or OR2 (N3701, N3699, N1276);
not NOT1 (N3702, N3698);
nand NAND2 (N3703, N3697, N371);
and AND3 (N3704, N3692, N2083, N154);
xor XOR2 (N3705, N3693, N83);
or OR3 (N3706, N3694, N1321, N2164);
nor NOR3 (N3707, N3702, N1995, N814);
xor XOR2 (N3708, N3701, N2375);
buf BUF1 (N3709, N3696);
not NOT1 (N3710, N3706);
or OR2 (N3711, N3704, N2356);
and AND2 (N3712, N3711, N485);
nor NOR3 (N3713, N3703, N1942, N2214);
not NOT1 (N3714, N3712);
nand NAND4 (N3715, N3700, N2274, N3072, N1085);
and AND4 (N3716, N3705, N2252, N2125, N3235);
and AND3 (N3717, N3708, N1979, N1916);
nor NOR4 (N3718, N3714, N44, N602, N2401);
buf BUF1 (N3719, N3715);
nand NAND2 (N3720, N3717, N1338);
nand NAND4 (N3721, N3690, N2610, N595, N1497);
xor XOR2 (N3722, N3721, N2113);
and AND4 (N3723, N3707, N3128, N2781, N2591);
buf BUF1 (N3724, N3723);
not NOT1 (N3725, N3695);
or OR2 (N3726, N3713, N3335);
buf BUF1 (N3727, N3710);
not NOT1 (N3728, N3709);
not NOT1 (N3729, N3722);
xor XOR2 (N3730, N3718, N438);
and AND2 (N3731, N3726, N177);
nor NOR2 (N3732, N3724, N3512);
buf BUF1 (N3733, N3731);
xor XOR2 (N3734, N3729, N2975);
and AND3 (N3735, N3733, N292, N607);
or OR3 (N3736, N3727, N3616, N3325);
xor XOR2 (N3737, N3725, N786);
nor NOR3 (N3738, N3736, N3165, N3736);
nand NAND3 (N3739, N3719, N2161, N1938);
or OR2 (N3740, N3737, N1130);
nor NOR4 (N3741, N3740, N2190, N2721, N3346);
nand NAND3 (N3742, N3732, N186, N1983);
and AND4 (N3743, N3738, N1656, N2782, N426);
buf BUF1 (N3744, N3730);
and AND4 (N3745, N3728, N1899, N3268, N3437);
not NOT1 (N3746, N3742);
nor NOR2 (N3747, N3743, N1172);
nand NAND3 (N3748, N3744, N449, N1939);
or OR2 (N3749, N3747, N1452);
and AND2 (N3750, N3741, N2891);
not NOT1 (N3751, N3720);
nor NOR4 (N3752, N3751, N1321, N2188, N1551);
nand NAND3 (N3753, N3752, N2086, N802);
and AND2 (N3754, N3734, N3399);
nor NOR4 (N3755, N3745, N1684, N2962, N3275);
nor NOR3 (N3756, N3739, N530, N715);
or OR4 (N3757, N3735, N681, N975, N1238);
nor NOR2 (N3758, N3748, N3284);
or OR4 (N3759, N3746, N315, N2230, N1751);
xor XOR2 (N3760, N3758, N620);
and AND3 (N3761, N3754, N3540, N3585);
not NOT1 (N3762, N3755);
xor XOR2 (N3763, N3756, N2643);
not NOT1 (N3764, N3760);
and AND3 (N3765, N3716, N862, N1863);
and AND3 (N3766, N3762, N3494, N3028);
not NOT1 (N3767, N3766);
and AND4 (N3768, N3765, N3, N22, N360);
or OR2 (N3769, N3763, N3673);
nor NOR4 (N3770, N3749, N1403, N1947, N2207);
nand NAND4 (N3771, N3759, N102, N2858, N3306);
nor NOR4 (N3772, N3764, N3412, N317, N606);
xor XOR2 (N3773, N3771, N3158);
nor NOR4 (N3774, N3753, N3273, N3412, N1870);
or OR4 (N3775, N3773, N1514, N3286, N2091);
buf BUF1 (N3776, N3757);
buf BUF1 (N3777, N3772);
buf BUF1 (N3778, N3750);
and AND3 (N3779, N3777, N1690, N450);
or OR3 (N3780, N3770, N3450, N1610);
nor NOR2 (N3781, N3780, N803);
not NOT1 (N3782, N3774);
and AND3 (N3783, N3775, N998, N3478);
buf BUF1 (N3784, N3778);
nand NAND3 (N3785, N3781, N2672, N3594);
or OR4 (N3786, N3785, N463, N3279, N2686);
or OR2 (N3787, N3776, N441);
not NOT1 (N3788, N3786);
nand NAND3 (N3789, N3784, N2229, N72);
xor XOR2 (N3790, N3761, N2031);
xor XOR2 (N3791, N3787, N3619);
nor NOR3 (N3792, N3790, N1805, N2565);
buf BUF1 (N3793, N3782);
and AND4 (N3794, N3767, N96, N1044, N2597);
nand NAND3 (N3795, N3789, N3350, N1829);
xor XOR2 (N3796, N3795, N2393);
buf BUF1 (N3797, N3794);
nand NAND3 (N3798, N3768, N3054, N3697);
not NOT1 (N3799, N3791);
or OR4 (N3800, N3788, N712, N1781, N841);
buf BUF1 (N3801, N3783);
nor NOR2 (N3802, N3798, N2048);
nor NOR2 (N3803, N3802, N959);
and AND3 (N3804, N3797, N1370, N3257);
nor NOR2 (N3805, N3804, N3372);
nor NOR4 (N3806, N3769, N1784, N2829, N3782);
xor XOR2 (N3807, N3800, N675);
xor XOR2 (N3808, N3805, N2470);
and AND2 (N3809, N3803, N316);
nand NAND3 (N3810, N3792, N890, N102);
nor NOR3 (N3811, N3809, N1239, N1434);
nand NAND3 (N3812, N3793, N3392, N1372);
or OR2 (N3813, N3806, N3114);
or OR4 (N3814, N3801, N1936, N3731, N308);
nand NAND2 (N3815, N3779, N3607);
and AND2 (N3816, N3799, N1818);
and AND4 (N3817, N3807, N2075, N2865, N2292);
nor NOR4 (N3818, N3817, N455, N2550, N1058);
or OR3 (N3819, N3816, N3275, N1124);
nor NOR3 (N3820, N3815, N2027, N2101);
or OR3 (N3821, N3813, N3634, N2388);
or OR4 (N3822, N3796, N3778, N1200, N3814);
xor XOR2 (N3823, N1922, N852);
and AND4 (N3824, N3821, N3681, N1793, N3798);
not NOT1 (N3825, N3824);
buf BUF1 (N3826, N3820);
xor XOR2 (N3827, N3808, N4);
not NOT1 (N3828, N3810);
not NOT1 (N3829, N3823);
nor NOR2 (N3830, N3811, N3556);
or OR4 (N3831, N3812, N3047, N1227, N1044);
nor NOR2 (N3832, N3822, N660);
not NOT1 (N3833, N3818);
or OR2 (N3834, N3825, N1844);
or OR3 (N3835, N3827, N3555, N3678);
nand NAND2 (N3836, N3819, N2097);
buf BUF1 (N3837, N3832);
nand NAND4 (N3838, N3826, N86, N1475, N3454);
not NOT1 (N3839, N3835);
buf BUF1 (N3840, N3834);
nand NAND3 (N3841, N3839, N3727, N3705);
not NOT1 (N3842, N3841);
nor NOR2 (N3843, N3836, N1321);
buf BUF1 (N3844, N3831);
or OR4 (N3845, N3830, N1134, N2520, N3375);
nor NOR4 (N3846, N3833, N2586, N1591, N3471);
nor NOR3 (N3847, N3843, N2139, N3238);
nor NOR4 (N3848, N3846, N2683, N753, N429);
not NOT1 (N3849, N3844);
xor XOR2 (N3850, N3849, N2623);
buf BUF1 (N3851, N3828);
nand NAND4 (N3852, N3840, N849, N1732, N1292);
nand NAND2 (N3853, N3838, N3271);
xor XOR2 (N3854, N3837, N3238);
nor NOR4 (N3855, N3852, N970, N684, N2051);
nor NOR2 (N3856, N3850, N388);
or OR3 (N3857, N3854, N589, N2129);
nor NOR3 (N3858, N3851, N90, N2290);
or OR3 (N3859, N3858, N1234, N3224);
or OR4 (N3860, N3857, N2844, N2801, N3687);
nand NAND2 (N3861, N3853, N247);
xor XOR2 (N3862, N3848, N1524);
xor XOR2 (N3863, N3860, N3403);
not NOT1 (N3864, N3861);
or OR3 (N3865, N3845, N857, N2579);
not NOT1 (N3866, N3862);
and AND2 (N3867, N3866, N3269);
and AND3 (N3868, N3863, N677, N1420);
not NOT1 (N3869, N3856);
buf BUF1 (N3870, N3869);
xor XOR2 (N3871, N3829, N3804);
nand NAND3 (N3872, N3870, N2338, N3132);
nor NOR2 (N3873, N3867, N1624);
nor NOR2 (N3874, N3859, N2500);
not NOT1 (N3875, N3868);
not NOT1 (N3876, N3865);
not NOT1 (N3877, N3872);
buf BUF1 (N3878, N3871);
nor NOR3 (N3879, N3855, N1703, N2694);
not NOT1 (N3880, N3864);
buf BUF1 (N3881, N3877);
and AND2 (N3882, N3879, N3057);
buf BUF1 (N3883, N3873);
and AND2 (N3884, N3881, N2631);
xor XOR2 (N3885, N3880, N196);
or OR2 (N3886, N3885, N1692);
nand NAND3 (N3887, N3874, N3357, N1333);
not NOT1 (N3888, N3886);
nor NOR2 (N3889, N3888, N1080);
nor NOR4 (N3890, N3887, N1777, N2230, N3424);
not NOT1 (N3891, N3890);
buf BUF1 (N3892, N3889);
or OR3 (N3893, N3875, N3003, N3470);
or OR3 (N3894, N3892, N3301, N3350);
nor NOR4 (N3895, N3894, N78, N3146, N1133);
buf BUF1 (N3896, N3893);
nor NOR2 (N3897, N3895, N989);
not NOT1 (N3898, N3878);
buf BUF1 (N3899, N3897);
not NOT1 (N3900, N3882);
buf BUF1 (N3901, N3898);
or OR2 (N3902, N3900, N2228);
nand NAND2 (N3903, N3842, N119);
nand NAND2 (N3904, N3899, N599);
or OR3 (N3905, N3883, N450, N1806);
not NOT1 (N3906, N3847);
buf BUF1 (N3907, N3904);
not NOT1 (N3908, N3876);
or OR3 (N3909, N3896, N3864, N3421);
nor NOR4 (N3910, N3902, N2790, N1980, N1445);
not NOT1 (N3911, N3891);
and AND3 (N3912, N3907, N168, N2090);
buf BUF1 (N3913, N3884);
and AND2 (N3914, N3909, N3302);
xor XOR2 (N3915, N3905, N3753);
or OR3 (N3916, N3910, N982, N1999);
and AND2 (N3917, N3906, N1478);
nand NAND3 (N3918, N3908, N399, N1270);
and AND4 (N3919, N3912, N1286, N1986, N687);
not NOT1 (N3920, N3915);
or OR3 (N3921, N3901, N3754, N3903);
nand NAND4 (N3922, N1999, N740, N3493, N2876);
xor XOR2 (N3923, N3918, N3292);
or OR2 (N3924, N3916, N172);
not NOT1 (N3925, N3917);
xor XOR2 (N3926, N3925, N3888);
nor NOR3 (N3927, N3914, N2580, N3670);
buf BUF1 (N3928, N3927);
not NOT1 (N3929, N3920);
nor NOR4 (N3930, N3921, N2950, N103, N1336);
nand NAND2 (N3931, N3924, N660);
nand NAND2 (N3932, N3922, N2929);
nand NAND3 (N3933, N3928, N3116, N1704);
and AND2 (N3934, N3913, N2816);
nand NAND4 (N3935, N3931, N144, N287, N2760);
and AND2 (N3936, N3935, N2225);
and AND4 (N3937, N3911, N1877, N3660, N2558);
xor XOR2 (N3938, N3919, N3789);
buf BUF1 (N3939, N3936);
nand NAND2 (N3940, N3934, N399);
and AND4 (N3941, N3940, N1684, N1505, N51);
nand NAND3 (N3942, N3929, N3106, N3420);
or OR3 (N3943, N3939, N1235, N926);
and AND3 (N3944, N3938, N3744, N277);
and AND2 (N3945, N3930, N1823);
not NOT1 (N3946, N3926);
xor XOR2 (N3947, N3946, N3749);
not NOT1 (N3948, N3942);
nand NAND2 (N3949, N3923, N2296);
not NOT1 (N3950, N3943);
nor NOR3 (N3951, N3947, N2655, N2653);
nor NOR3 (N3952, N3950, N2046, N2592);
nand NAND2 (N3953, N3932, N886);
xor XOR2 (N3954, N3941, N193);
nor NOR4 (N3955, N3952, N1977, N154, N1939);
buf BUF1 (N3956, N3937);
or OR4 (N3957, N3951, N303, N208, N1532);
nor NOR4 (N3958, N3945, N3062, N3500, N3574);
not NOT1 (N3959, N3956);
nor NOR4 (N3960, N3959, N2452, N587, N1829);
nand NAND4 (N3961, N3960, N586, N32, N238);
nand NAND3 (N3962, N3948, N901, N1595);
buf BUF1 (N3963, N3961);
or OR4 (N3964, N3955, N80, N2367, N1785);
nand NAND3 (N3965, N3957, N1435, N1262);
buf BUF1 (N3966, N3965);
buf BUF1 (N3967, N3953);
nand NAND2 (N3968, N3958, N2117);
or OR2 (N3969, N3963, N69);
and AND2 (N3970, N3969, N1761);
buf BUF1 (N3971, N3964);
buf BUF1 (N3972, N3966);
nand NAND3 (N3973, N3944, N2139, N1659);
buf BUF1 (N3974, N3933);
or OR2 (N3975, N3954, N1373);
or OR4 (N3976, N3949, N2027, N3638, N2968);
and AND2 (N3977, N3975, N825);
xor XOR2 (N3978, N3974, N2630);
not NOT1 (N3979, N3973);
or OR3 (N3980, N3967, N2462, N853);
buf BUF1 (N3981, N3976);
and AND4 (N3982, N3962, N502, N3867, N1686);
nor NOR3 (N3983, N3977, N2580, N2113);
or OR3 (N3984, N3980, N2153, N337);
or OR4 (N3985, N3971, N2908, N1148, N726);
or OR2 (N3986, N3981, N1693);
and AND4 (N3987, N3968, N213, N2491, N98);
nand NAND4 (N3988, N3986, N2269, N255, N428);
and AND4 (N3989, N3987, N2461, N2241, N2340);
or OR4 (N3990, N3979, N3774, N1004, N1349);
or OR3 (N3991, N3982, N1434, N2888);
not NOT1 (N3992, N3988);
nor NOR3 (N3993, N3983, N2975, N1239);
not NOT1 (N3994, N3985);
and AND4 (N3995, N3972, N3609, N3713, N118);
xor XOR2 (N3996, N3990, N2908);
and AND3 (N3997, N3989, N2684, N3319);
xor XOR2 (N3998, N3995, N2648);
and AND2 (N3999, N3978, N825);
nor NOR3 (N4000, N3993, N743, N1532);
buf BUF1 (N4001, N3970);
not NOT1 (N4002, N3997);
nor NOR4 (N4003, N3984, N1075, N2424, N3180);
and AND2 (N4004, N3991, N1113);
or OR4 (N4005, N4001, N844, N3778, N708);
buf BUF1 (N4006, N4000);
nor NOR2 (N4007, N3996, N3665);
nor NOR2 (N4008, N4007, N3133);
not NOT1 (N4009, N4005);
nor NOR4 (N4010, N3999, N2279, N2109, N1324);
nand NAND3 (N4011, N4009, N1080, N655);
nand NAND2 (N4012, N4011, N75);
nand NAND2 (N4013, N3994, N1336);
nand NAND3 (N4014, N4003, N2727, N279);
xor XOR2 (N4015, N4010, N805);
and AND4 (N4016, N3998, N2633, N2630, N3630);
not NOT1 (N4017, N4006);
xor XOR2 (N4018, N4004, N963);
buf BUF1 (N4019, N4002);
nand NAND2 (N4020, N3992, N2484);
buf BUF1 (N4021, N4008);
xor XOR2 (N4022, N4017, N494);
not NOT1 (N4023, N4018);
and AND2 (N4024, N4014, N342);
and AND3 (N4025, N4024, N622, N1589);
not NOT1 (N4026, N4025);
nor NOR3 (N4027, N4013, N645, N1547);
not NOT1 (N4028, N4012);
xor XOR2 (N4029, N4022, N283);
buf BUF1 (N4030, N4029);
nand NAND2 (N4031, N4026, N328);
nand NAND2 (N4032, N4030, N346);
xor XOR2 (N4033, N4021, N1389);
nor NOR3 (N4034, N4023, N2734, N2970);
nor NOR4 (N4035, N4031, N2282, N2960, N439);
buf BUF1 (N4036, N4019);
xor XOR2 (N4037, N4015, N3019);
nor NOR3 (N4038, N4016, N528, N1414);
xor XOR2 (N4039, N4033, N2789);
nand NAND3 (N4040, N4037, N3865, N3649);
not NOT1 (N4041, N4020);
nor NOR2 (N4042, N4039, N612);
nand NAND4 (N4043, N4040, N84, N1088, N271);
nor NOR3 (N4044, N4038, N3705, N1014);
nand NAND2 (N4045, N4035, N3882);
xor XOR2 (N4046, N4027, N2734);
nand NAND2 (N4047, N4036, N2868);
not NOT1 (N4048, N4028);
nand NAND2 (N4049, N4043, N3946);
nand NAND2 (N4050, N4032, N4035);
nor NOR2 (N4051, N4049, N3149);
not NOT1 (N4052, N4045);
nand NAND4 (N4053, N4034, N1583, N2988, N113);
or OR4 (N4054, N4044, N612, N392, N3324);
nor NOR2 (N4055, N4046, N2890);
nand NAND2 (N4056, N4051, N1037);
or OR3 (N4057, N4055, N2291, N2950);
not NOT1 (N4058, N4056);
and AND2 (N4059, N4042, N3777);
and AND3 (N4060, N4053, N1937, N896);
buf BUF1 (N4061, N4050);
xor XOR2 (N4062, N4052, N1150);
buf BUF1 (N4063, N4060);
nor NOR2 (N4064, N4059, N3686);
nor NOR3 (N4065, N4058, N3273, N2243);
buf BUF1 (N4066, N4041);
buf BUF1 (N4067, N4061);
xor XOR2 (N4068, N4047, N3172);
buf BUF1 (N4069, N4054);
buf BUF1 (N4070, N4062);
xor XOR2 (N4071, N4068, N2735);
not NOT1 (N4072, N4064);
buf BUF1 (N4073, N4066);
or OR2 (N4074, N4073, N1836);
and AND3 (N4075, N4069, N2934, N2024);
buf BUF1 (N4076, N4048);
and AND3 (N4077, N4057, N950, N3895);
nor NOR4 (N4078, N4067, N260, N1387, N3320);
nor NOR4 (N4079, N4065, N773, N2902, N3326);
nand NAND2 (N4080, N4076, N2265);
buf BUF1 (N4081, N4070);
xor XOR2 (N4082, N4074, N796);
nand NAND2 (N4083, N4078, N1966);
xor XOR2 (N4084, N4082, N1546);
xor XOR2 (N4085, N4063, N3913);
or OR3 (N4086, N4085, N1678, N2233);
nor NOR2 (N4087, N4075, N2728);
or OR2 (N4088, N4083, N649);
nor NOR3 (N4089, N4080, N976, N801);
or OR2 (N4090, N4081, N3755);
not NOT1 (N4091, N4086);
or OR2 (N4092, N4090, N1149);
and AND3 (N4093, N4089, N25, N3787);
xor XOR2 (N4094, N4084, N429);
nor NOR3 (N4095, N4093, N1404, N2911);
nand NAND2 (N4096, N4088, N2060);
not NOT1 (N4097, N4072);
xor XOR2 (N4098, N4095, N411);
nand NAND3 (N4099, N4079, N3987, N3091);
xor XOR2 (N4100, N4097, N773);
or OR3 (N4101, N4091, N1800, N493);
xor XOR2 (N4102, N4087, N87);
nand NAND4 (N4103, N4099, N1270, N2390, N2915);
not NOT1 (N4104, N4101);
buf BUF1 (N4105, N4096);
buf BUF1 (N4106, N4104);
and AND3 (N4107, N4103, N3312, N2092);
and AND2 (N4108, N4106, N2259);
buf BUF1 (N4109, N4108);
or OR2 (N4110, N4098, N1793);
nor NOR2 (N4111, N4107, N4098);
nor NOR2 (N4112, N4111, N788);
or OR3 (N4113, N4092, N474, N3339);
or OR4 (N4114, N4077, N2386, N1539, N2019);
not NOT1 (N4115, N4071);
not NOT1 (N4116, N4113);
nand NAND2 (N4117, N4110, N2962);
or OR4 (N4118, N4094, N1814, N2953, N2906);
nand NAND4 (N4119, N4118, N2854, N276, N830);
nand NAND2 (N4120, N4112, N1808);
or OR3 (N4121, N4120, N2029, N306);
or OR3 (N4122, N4100, N1614, N1700);
or OR2 (N4123, N4102, N3996);
buf BUF1 (N4124, N4105);
nor NOR4 (N4125, N4116, N3631, N3608, N645);
nand NAND2 (N4126, N4125, N2662);
not NOT1 (N4127, N4126);
not NOT1 (N4128, N4109);
buf BUF1 (N4129, N4114);
xor XOR2 (N4130, N4128, N266);
xor XOR2 (N4131, N4115, N3645);
not NOT1 (N4132, N4130);
buf BUF1 (N4133, N4129);
nand NAND4 (N4134, N4122, N1847, N2420, N1027);
or OR4 (N4135, N4132, N193, N2779, N3267);
xor XOR2 (N4136, N4127, N1626);
and AND3 (N4137, N4124, N2036, N1134);
xor XOR2 (N4138, N4121, N3540);
and AND4 (N4139, N4137, N1661, N3637, N463);
xor XOR2 (N4140, N4138, N40);
nand NAND4 (N4141, N4117, N356, N3940, N2822);
xor XOR2 (N4142, N4139, N213);
nor NOR2 (N4143, N4119, N1318);
xor XOR2 (N4144, N4141, N1171);
or OR4 (N4145, N4133, N3024, N1238, N975);
buf BUF1 (N4146, N4135);
and AND4 (N4147, N4144, N3836, N1957, N2894);
not NOT1 (N4148, N4136);
buf BUF1 (N4149, N4148);
nand NAND3 (N4150, N4134, N154, N2870);
buf BUF1 (N4151, N4140);
or OR3 (N4152, N4131, N483, N1695);
nand NAND3 (N4153, N4145, N1977, N1762);
nand NAND3 (N4154, N4150, N767, N62);
not NOT1 (N4155, N4152);
nand NAND4 (N4156, N4151, N2636, N1159, N1022);
nand NAND3 (N4157, N4147, N1185, N1282);
xor XOR2 (N4158, N4142, N3157);
nand NAND4 (N4159, N4155, N3362, N1386, N840);
and AND4 (N4160, N4154, N3347, N1852, N1398);
not NOT1 (N4161, N4157);
nand NAND2 (N4162, N4160, N1286);
and AND3 (N4163, N4149, N2856, N3094);
nor NOR3 (N4164, N4163, N839, N1727);
buf BUF1 (N4165, N4146);
nor NOR4 (N4166, N4159, N1207, N3712, N2415);
xor XOR2 (N4167, N4166, N2596);
nor NOR3 (N4168, N4164, N3408, N2531);
xor XOR2 (N4169, N4161, N1191);
not NOT1 (N4170, N4153);
nand NAND4 (N4171, N4158, N2111, N3943, N1347);
and AND3 (N4172, N4162, N1422, N3008);
or OR2 (N4173, N4143, N3554);
xor XOR2 (N4174, N4167, N2534);
nand NAND3 (N4175, N4165, N3641, N1087);
buf BUF1 (N4176, N4175);
or OR3 (N4177, N4172, N699, N3633);
buf BUF1 (N4178, N4171);
buf BUF1 (N4179, N4123);
xor XOR2 (N4180, N4176, N1021);
nand NAND3 (N4181, N4169, N2408, N603);
nand NAND2 (N4182, N4180, N406);
buf BUF1 (N4183, N4170);
and AND2 (N4184, N4173, N232);
buf BUF1 (N4185, N4177);
and AND3 (N4186, N4182, N1576, N2020);
not NOT1 (N4187, N4185);
buf BUF1 (N4188, N4174);
not NOT1 (N4189, N4181);
xor XOR2 (N4190, N4189, N1899);
nor NOR3 (N4191, N4187, N2389, N1935);
nand NAND2 (N4192, N4190, N519);
and AND3 (N4193, N4184, N101, N2444);
and AND2 (N4194, N4168, N4120);
nor NOR2 (N4195, N4191, N3000);
or OR3 (N4196, N4179, N1883, N3502);
nand NAND3 (N4197, N4156, N1897, N2487);
or OR4 (N4198, N4183, N3400, N1097, N2404);
or OR3 (N4199, N4195, N1264, N1956);
nor NOR4 (N4200, N4188, N2736, N2865, N1397);
buf BUF1 (N4201, N4197);
xor XOR2 (N4202, N4194, N836);
nand NAND4 (N4203, N4201, N1891, N985, N2089);
not NOT1 (N4204, N4202);
not NOT1 (N4205, N4193);
not NOT1 (N4206, N4198);
xor XOR2 (N4207, N4178, N1629);
or OR4 (N4208, N4204, N1380, N3763, N2681);
nor NOR3 (N4209, N4192, N91, N2557);
xor XOR2 (N4210, N4199, N1678);
nand NAND3 (N4211, N4203, N1709, N421);
or OR3 (N4212, N4205, N1430, N671);
xor XOR2 (N4213, N4211, N2481);
nor NOR2 (N4214, N4207, N2660);
not NOT1 (N4215, N4213);
nand NAND4 (N4216, N4208, N2661, N3713, N2067);
xor XOR2 (N4217, N4186, N1665);
xor XOR2 (N4218, N4209, N1953);
not NOT1 (N4219, N4218);
or OR2 (N4220, N4216, N3339);
xor XOR2 (N4221, N4212, N4009);
xor XOR2 (N4222, N4217, N2709);
buf BUF1 (N4223, N4215);
nor NOR3 (N4224, N4222, N991, N219);
and AND2 (N4225, N4224, N1504);
and AND4 (N4226, N4225, N2886, N2323, N76);
not NOT1 (N4227, N4214);
nand NAND3 (N4228, N4200, N185, N3191);
xor XOR2 (N4229, N4228, N3665);
or OR4 (N4230, N4221, N3009, N3667, N5);
and AND2 (N4231, N4210, N31);
buf BUF1 (N4232, N4227);
and AND3 (N4233, N4232, N4028, N318);
nand NAND2 (N4234, N4231, N2995);
xor XOR2 (N4235, N4196, N2065);
xor XOR2 (N4236, N4219, N4077);
and AND4 (N4237, N4220, N784, N2776, N55);
nor NOR4 (N4238, N4234, N3907, N3155, N1627);
not NOT1 (N4239, N4236);
nand NAND4 (N4240, N4237, N2249, N3015, N2499);
nor NOR3 (N4241, N4240, N282, N3351);
nor NOR3 (N4242, N4241, N1648, N678);
not NOT1 (N4243, N4230);
or OR3 (N4244, N4226, N3015, N1207);
and AND3 (N4245, N4239, N3281, N2793);
nand NAND3 (N4246, N4245, N1130, N1035);
not NOT1 (N4247, N4246);
not NOT1 (N4248, N4247);
buf BUF1 (N4249, N4235);
buf BUF1 (N4250, N4229);
not NOT1 (N4251, N4250);
nor NOR2 (N4252, N4248, N3127);
nand NAND3 (N4253, N4206, N2647, N3226);
or OR2 (N4254, N4244, N2880);
and AND3 (N4255, N4249, N1665, N4015);
nand NAND2 (N4256, N4253, N3711);
nor NOR4 (N4257, N4238, N1660, N826, N7);
or OR3 (N4258, N4255, N4092, N1250);
not NOT1 (N4259, N4254);
or OR3 (N4260, N4258, N1557, N450);
or OR2 (N4261, N4252, N1790);
and AND2 (N4262, N4261, N2880);
nor NOR3 (N4263, N4260, N3191, N1175);
xor XOR2 (N4264, N4233, N2895);
xor XOR2 (N4265, N4256, N3740);
not NOT1 (N4266, N4257);
nand NAND2 (N4267, N4251, N3947);
not NOT1 (N4268, N4266);
or OR2 (N4269, N4263, N453);
buf BUF1 (N4270, N4264);
not NOT1 (N4271, N4265);
xor XOR2 (N4272, N4262, N4143);
nor NOR2 (N4273, N4259, N1991);
xor XOR2 (N4274, N4269, N2343);
nor NOR3 (N4275, N4243, N286, N1202);
xor XOR2 (N4276, N4275, N3867);
or OR4 (N4277, N4270, N304, N55, N1031);
buf BUF1 (N4278, N4277);
and AND4 (N4279, N4274, N3396, N1230, N1118);
nand NAND4 (N4280, N4242, N4228, N2313, N1787);
nand NAND3 (N4281, N4280, N190, N4197);
or OR3 (N4282, N4278, N3110, N2025);
buf BUF1 (N4283, N4272);
and AND2 (N4284, N4276, N970);
nor NOR4 (N4285, N4271, N1316, N2256, N2265);
or OR4 (N4286, N4283, N1061, N949, N1357);
buf BUF1 (N4287, N4273);
buf BUF1 (N4288, N4279);
buf BUF1 (N4289, N4281);
or OR4 (N4290, N4289, N3008, N3571, N266);
nor NOR4 (N4291, N4288, N789, N3133, N2544);
xor XOR2 (N4292, N4284, N1087);
nand NAND4 (N4293, N4287, N1488, N3827, N2186);
buf BUF1 (N4294, N4282);
xor XOR2 (N4295, N4267, N3942);
nor NOR4 (N4296, N4286, N1079, N1042, N1185);
xor XOR2 (N4297, N4223, N1868);
nor NOR3 (N4298, N4294, N2464, N379);
and AND4 (N4299, N4298, N1926, N2762, N3511);
nor NOR2 (N4300, N4296, N1048);
nand NAND4 (N4301, N4285, N2300, N3473, N777);
not NOT1 (N4302, N4297);
or OR4 (N4303, N4302, N2466, N1420, N575);
xor XOR2 (N4304, N4292, N2054);
buf BUF1 (N4305, N4291);
nor NOR4 (N4306, N4305, N2954, N3936, N1479);
and AND4 (N4307, N4301, N2676, N2620, N891);
not NOT1 (N4308, N4307);
or OR3 (N4309, N4306, N3309, N1795);
buf BUF1 (N4310, N4293);
or OR3 (N4311, N4268, N1202, N4196);
or OR2 (N4312, N4310, N3105);
and AND3 (N4313, N4311, N3377, N3581);
nor NOR3 (N4314, N4308, N1324, N2631);
nand NAND4 (N4315, N4300, N1632, N3882, N837);
and AND2 (N4316, N4299, N1214);
or OR2 (N4317, N4312, N2835);
or OR3 (N4318, N4317, N3326, N1935);
nand NAND3 (N4319, N4313, N685, N588);
nand NAND2 (N4320, N4318, N3516);
or OR4 (N4321, N4295, N961, N2869, N2400);
or OR4 (N4322, N4316, N2862, N1463, N1257);
and AND3 (N4323, N4304, N1706, N2038);
not NOT1 (N4324, N4314);
nor NOR2 (N4325, N4290, N3752);
not NOT1 (N4326, N4321);
buf BUF1 (N4327, N4326);
nor NOR3 (N4328, N4315, N1117, N1239);
and AND3 (N4329, N4309, N2418, N1590);
not NOT1 (N4330, N4319);
nand NAND2 (N4331, N4329, N516);
and AND4 (N4332, N4320, N4169, N3886, N2575);
xor XOR2 (N4333, N4332, N3659);
nand NAND3 (N4334, N4323, N954, N3175);
not NOT1 (N4335, N4325);
nor NOR2 (N4336, N4324, N431);
nor NOR4 (N4337, N4327, N1270, N1668, N1950);
not NOT1 (N4338, N4334);
buf BUF1 (N4339, N4337);
buf BUF1 (N4340, N4333);
nand NAND3 (N4341, N4335, N3313, N3207);
xor XOR2 (N4342, N4340, N3811);
nand NAND4 (N4343, N4303, N452, N2576, N2481);
buf BUF1 (N4344, N4338);
nand NAND2 (N4345, N4344, N469);
and AND4 (N4346, N4342, N2436, N1169, N2435);
buf BUF1 (N4347, N4343);
buf BUF1 (N4348, N4322);
xor XOR2 (N4349, N4348, N3791);
buf BUF1 (N4350, N4328);
nand NAND2 (N4351, N4331, N1719);
or OR3 (N4352, N4336, N775, N2566);
buf BUF1 (N4353, N4347);
and AND3 (N4354, N4339, N1935, N3314);
nand NAND4 (N4355, N4346, N2439, N803, N346);
buf BUF1 (N4356, N4352);
and AND2 (N4357, N4349, N3128);
nand NAND4 (N4358, N4357, N2202, N3856, N1895);
or OR4 (N4359, N4355, N4346, N96, N4172);
or OR3 (N4360, N4353, N723, N2769);
not NOT1 (N4361, N4358);
and AND4 (N4362, N4330, N1689, N1818, N229);
or OR3 (N4363, N4345, N37, N4118);
nor NOR3 (N4364, N4351, N3654, N1469);
nor NOR3 (N4365, N4354, N526, N1478);
not NOT1 (N4366, N4362);
xor XOR2 (N4367, N4364, N2309);
xor XOR2 (N4368, N4365, N2429);
or OR3 (N4369, N4360, N174, N862);
buf BUF1 (N4370, N4350);
nor NOR3 (N4371, N4361, N1012, N644);
not NOT1 (N4372, N4359);
or OR4 (N4373, N4356, N1990, N1342, N1544);
xor XOR2 (N4374, N4366, N3817);
nand NAND3 (N4375, N4363, N78, N3898);
and AND2 (N4376, N4369, N1048);
buf BUF1 (N4377, N4373);
or OR2 (N4378, N4341, N3713);
nor NOR2 (N4379, N4378, N4117);
nor NOR2 (N4380, N4367, N4311);
xor XOR2 (N4381, N4380, N3170);
or OR3 (N4382, N4371, N1325, N4028);
not NOT1 (N4383, N4376);
buf BUF1 (N4384, N4370);
buf BUF1 (N4385, N4382);
not NOT1 (N4386, N4385);
nand NAND2 (N4387, N4383, N43);
buf BUF1 (N4388, N4375);
nor NOR2 (N4389, N4384, N3151);
not NOT1 (N4390, N4368);
or OR3 (N4391, N4379, N561, N807);
or OR3 (N4392, N4374, N436, N4155);
nor NOR3 (N4393, N4386, N2450, N2129);
nand NAND3 (N4394, N4377, N3898, N1795);
and AND4 (N4395, N4392, N1281, N1228, N3411);
buf BUF1 (N4396, N4395);
xor XOR2 (N4397, N4390, N1539);
buf BUF1 (N4398, N4391);
not NOT1 (N4399, N4398);
and AND3 (N4400, N4372, N4267, N4040);
and AND3 (N4401, N4399, N1779, N1129);
xor XOR2 (N4402, N4389, N3712);
nand NAND3 (N4403, N4397, N47, N3882);
or OR4 (N4404, N4388, N2021, N41, N3327);
not NOT1 (N4405, N4402);
and AND3 (N4406, N4396, N3337, N3460);
nor NOR3 (N4407, N4406, N1283, N2718);
buf BUF1 (N4408, N4381);
nor NOR4 (N4409, N4405, N1723, N160, N2776);
nand NAND3 (N4410, N4387, N1585, N2549);
nor NOR4 (N4411, N4394, N1102, N2209, N2818);
xor XOR2 (N4412, N4410, N4006);
or OR4 (N4413, N4409, N2331, N1149, N890);
not NOT1 (N4414, N4400);
and AND2 (N4415, N4412, N3135);
or OR3 (N4416, N4393, N2777, N3409);
and AND4 (N4417, N4401, N362, N2231, N1635);
and AND3 (N4418, N4411, N2552, N1325);
or OR4 (N4419, N4404, N1906, N2844, N1753);
not NOT1 (N4420, N4417);
xor XOR2 (N4421, N4413, N3251);
nand NAND4 (N4422, N4415, N3114, N1842, N211);
nand NAND4 (N4423, N4408, N3739, N2315, N1554);
and AND2 (N4424, N4403, N2672);
or OR2 (N4425, N4419, N2767);
or OR4 (N4426, N4418, N1409, N777, N3518);
xor XOR2 (N4427, N4426, N348);
nand NAND2 (N4428, N4425, N644);
nor NOR3 (N4429, N4407, N2379, N1948);
nand NAND2 (N4430, N4422, N2065);
and AND2 (N4431, N4414, N3402);
nand NAND2 (N4432, N4420, N504);
or OR2 (N4433, N4428, N4123);
and AND3 (N4434, N4433, N2591, N4187);
nand NAND2 (N4435, N4431, N635);
buf BUF1 (N4436, N4432);
or OR3 (N4437, N4424, N432, N2640);
nand NAND2 (N4438, N4430, N4235);
or OR4 (N4439, N4436, N724, N2342, N229);
buf BUF1 (N4440, N4434);
nand NAND2 (N4441, N4440, N4095);
nand NAND3 (N4442, N4421, N3245, N4087);
nor NOR3 (N4443, N4438, N43, N4417);
buf BUF1 (N4444, N4429);
nand NAND2 (N4445, N4423, N750);
and AND4 (N4446, N4427, N1084, N2085, N4305);
nor NOR4 (N4447, N4442, N1574, N1839, N320);
buf BUF1 (N4448, N4445);
buf BUF1 (N4449, N4444);
buf BUF1 (N4450, N4446);
nor NOR4 (N4451, N4448, N3666, N401, N2195);
buf BUF1 (N4452, N4447);
not NOT1 (N4453, N4416);
buf BUF1 (N4454, N4452);
buf BUF1 (N4455, N4437);
and AND2 (N4456, N4451, N45);
nor NOR4 (N4457, N4454, N77, N906, N1857);
buf BUF1 (N4458, N4439);
and AND2 (N4459, N4435, N2263);
not NOT1 (N4460, N4453);
xor XOR2 (N4461, N4450, N2835);
nor NOR4 (N4462, N4458, N704, N3785, N1708);
and AND3 (N4463, N4443, N1705, N4111);
not NOT1 (N4464, N4462);
xor XOR2 (N4465, N4455, N2725);
nand NAND4 (N4466, N4456, N2659, N2085, N18);
xor XOR2 (N4467, N4459, N3368);
nor NOR3 (N4468, N4464, N2528, N2200);
and AND3 (N4469, N4457, N1519, N601);
xor XOR2 (N4470, N4463, N4026);
buf BUF1 (N4471, N4466);
or OR2 (N4472, N4460, N2002);
xor XOR2 (N4473, N4470, N2024);
buf BUF1 (N4474, N4469);
buf BUF1 (N4475, N4467);
and AND2 (N4476, N4468, N3254);
buf BUF1 (N4477, N4475);
or OR3 (N4478, N4476, N4026, N3320);
buf BUF1 (N4479, N4477);
and AND4 (N4480, N4478, N112, N295, N4293);
nor NOR3 (N4481, N4461, N2988, N1803);
xor XOR2 (N4482, N4465, N10);
buf BUF1 (N4483, N4479);
nand NAND3 (N4484, N4480, N2861, N3943);
or OR4 (N4485, N4484, N1493, N3888, N1494);
and AND3 (N4486, N4481, N1639, N4002);
and AND2 (N4487, N4482, N917);
not NOT1 (N4488, N4474);
or OR4 (N4489, N4485, N2413, N3316, N605);
nor NOR3 (N4490, N4489, N974, N4040);
nand NAND4 (N4491, N4486, N2733, N4319, N1559);
xor XOR2 (N4492, N4487, N2977);
or OR2 (N4493, N4490, N1808);
nor NOR4 (N4494, N4472, N562, N2442, N1578);
xor XOR2 (N4495, N4471, N3268);
nand NAND4 (N4496, N4473, N2939, N2367, N1889);
nor NOR2 (N4497, N4494, N2503);
or OR4 (N4498, N4483, N545, N1029, N847);
not NOT1 (N4499, N4441);
buf BUF1 (N4500, N4497);
buf BUF1 (N4501, N4493);
buf BUF1 (N4502, N4488);
buf BUF1 (N4503, N4491);
or OR2 (N4504, N4502, N2003);
buf BUF1 (N4505, N4449);
nand NAND4 (N4506, N4492, N2752, N791, N2203);
and AND2 (N4507, N4500, N3501);
and AND3 (N4508, N4496, N3537, N3241);
or OR2 (N4509, N4503, N3742);
not NOT1 (N4510, N4495);
not NOT1 (N4511, N4507);
nor NOR3 (N4512, N4499, N1998, N1591);
nor NOR3 (N4513, N4501, N4112, N2280);
not NOT1 (N4514, N4509);
and AND3 (N4515, N4514, N1863, N4470);
xor XOR2 (N4516, N4510, N1616);
or OR3 (N4517, N4505, N2979, N3318);
or OR2 (N4518, N4517, N1556);
and AND2 (N4519, N4504, N2825);
buf BUF1 (N4520, N4513);
nor NOR2 (N4521, N4511, N2210);
buf BUF1 (N4522, N4515);
xor XOR2 (N4523, N4521, N3485);
or OR2 (N4524, N4506, N3792);
nand NAND3 (N4525, N4524, N3091, N4462);
xor XOR2 (N4526, N4519, N2150);
not NOT1 (N4527, N4508);
nand NAND4 (N4528, N4522, N3719, N1787, N3676);
buf BUF1 (N4529, N4523);
xor XOR2 (N4530, N4512, N2863);
not NOT1 (N4531, N4498);
buf BUF1 (N4532, N4529);
nor NOR3 (N4533, N4532, N346, N3598);
not NOT1 (N4534, N4533);
nand NAND4 (N4535, N4528, N621, N575, N782);
buf BUF1 (N4536, N4527);
and AND3 (N4537, N4530, N3572, N1554);
and AND3 (N4538, N4531, N1211, N1487);
nor NOR3 (N4539, N4536, N2712, N3840);
and AND2 (N4540, N4526, N3746);
nor NOR3 (N4541, N4525, N3620, N566);
not NOT1 (N4542, N4534);
or OR2 (N4543, N4520, N4056);
nor NOR2 (N4544, N4518, N858);
and AND3 (N4545, N4543, N2478, N4362);
nor NOR4 (N4546, N4542, N3727, N590, N4423);
not NOT1 (N4547, N4541);
xor XOR2 (N4548, N4537, N3691);
nand NAND4 (N4549, N4516, N995, N1975, N3299);
nor NOR4 (N4550, N4539, N2425, N2038, N3551);
and AND3 (N4551, N4544, N1852, N1426);
not NOT1 (N4552, N4545);
buf BUF1 (N4553, N4549);
or OR2 (N4554, N4550, N2699);
buf BUF1 (N4555, N4547);
xor XOR2 (N4556, N4540, N1207);
buf BUF1 (N4557, N4556);
xor XOR2 (N4558, N4548, N1283);
nor NOR4 (N4559, N4554, N3224, N3260, N3274);
nand NAND4 (N4560, N4559, N880, N2507, N2129);
xor XOR2 (N4561, N4555, N907);
and AND2 (N4562, N4535, N3616);
nor NOR4 (N4563, N4551, N3371, N2219, N497);
or OR4 (N4564, N4538, N2122, N3530, N1675);
and AND2 (N4565, N4564, N4274);
nand NAND3 (N4566, N4562, N4503, N1057);
nand NAND2 (N4567, N4561, N2361);
xor XOR2 (N4568, N4553, N1248);
or OR3 (N4569, N4567, N995, N1112);
nor NOR3 (N4570, N4558, N1660, N2670);
nor NOR4 (N4571, N4570, N4543, N2447, N3031);
buf BUF1 (N4572, N4546);
nor NOR3 (N4573, N4569, N1110, N4256);
nand NAND2 (N4574, N4572, N124);
and AND4 (N4575, N4573, N645, N977, N1054);
and AND3 (N4576, N4566, N4071, N3232);
buf BUF1 (N4577, N4565);
or OR4 (N4578, N4552, N2257, N2853, N3367);
nor NOR3 (N4579, N4557, N416, N4081);
xor XOR2 (N4580, N4578, N308);
buf BUF1 (N4581, N4577);
xor XOR2 (N4582, N4575, N3696);
nand NAND2 (N4583, N4568, N60);
and AND2 (N4584, N4583, N104);
and AND3 (N4585, N4560, N2013, N702);
or OR4 (N4586, N4582, N446, N2156, N1585);
buf BUF1 (N4587, N4574);
nor NOR4 (N4588, N4571, N2432, N4453, N1725);
nor NOR3 (N4589, N4580, N3626, N3406);
or OR2 (N4590, N4585, N264);
buf BUF1 (N4591, N4586);
xor XOR2 (N4592, N4591, N2009);
nor NOR3 (N4593, N4584, N469, N2338);
nor NOR4 (N4594, N4563, N3125, N2849, N4504);
and AND3 (N4595, N4589, N3762, N1073);
xor XOR2 (N4596, N4592, N1289);
buf BUF1 (N4597, N4595);
nand NAND2 (N4598, N4576, N2781);
not NOT1 (N4599, N4594);
buf BUF1 (N4600, N4598);
not NOT1 (N4601, N4581);
nor NOR2 (N4602, N4588, N3995);
buf BUF1 (N4603, N4593);
buf BUF1 (N4604, N4597);
nor NOR2 (N4605, N4601, N1567);
buf BUF1 (N4606, N4602);
nand NAND3 (N4607, N4579, N3469, N2721);
or OR2 (N4608, N4603, N103);
nand NAND3 (N4609, N4607, N3365, N4312);
not NOT1 (N4610, N4604);
nor NOR2 (N4611, N4608, N3315);
and AND4 (N4612, N4605, N4075, N3396, N997);
and AND4 (N4613, N4609, N2533, N4482, N4094);
buf BUF1 (N4614, N4606);
buf BUF1 (N4615, N4612);
not NOT1 (N4616, N4611);
xor XOR2 (N4617, N4599, N2638);
or OR2 (N4618, N4587, N2722);
nand NAND3 (N4619, N4590, N2855, N2914);
nand NAND4 (N4620, N4596, N3039, N780, N1973);
not NOT1 (N4621, N4620);
and AND2 (N4622, N4616, N2085);
xor XOR2 (N4623, N4615, N352);
or OR3 (N4624, N4621, N1533, N1726);
nor NOR2 (N4625, N4623, N574);
nor NOR4 (N4626, N4624, N1791, N32, N4466);
or OR2 (N4627, N4600, N2366);
nand NAND2 (N4628, N4619, N1406);
nand NAND2 (N4629, N4626, N1567);
and AND2 (N4630, N4622, N2041);
nand NAND2 (N4631, N4613, N1414);
not NOT1 (N4632, N4625);
and AND2 (N4633, N4630, N184);
xor XOR2 (N4634, N4631, N3387);
or OR2 (N4635, N4629, N2416);
and AND3 (N4636, N4610, N2382, N3864);
not NOT1 (N4637, N4614);
buf BUF1 (N4638, N4636);
nand NAND3 (N4639, N4627, N3571, N3037);
xor XOR2 (N4640, N4638, N55);
xor XOR2 (N4641, N4618, N4563);
or OR3 (N4642, N4640, N3707, N3303);
buf BUF1 (N4643, N4632);
nor NOR2 (N4644, N4639, N3009);
or OR2 (N4645, N4635, N1437);
not NOT1 (N4646, N4643);
buf BUF1 (N4647, N4642);
and AND2 (N4648, N4617, N2873);
and AND2 (N4649, N4644, N1809);
buf BUF1 (N4650, N4637);
nor NOR4 (N4651, N4628, N2824, N4558, N4337);
nor NOR2 (N4652, N4634, N4159);
xor XOR2 (N4653, N4647, N1768);
or OR2 (N4654, N4646, N4381);
not NOT1 (N4655, N4651);
buf BUF1 (N4656, N4654);
nand NAND2 (N4657, N4645, N2225);
nor NOR3 (N4658, N4652, N3132, N3954);
and AND3 (N4659, N4655, N437, N4128);
and AND2 (N4660, N4648, N661);
xor XOR2 (N4661, N4650, N4261);
nand NAND3 (N4662, N4660, N2431, N3558);
not NOT1 (N4663, N4656);
and AND4 (N4664, N4658, N2784, N323, N615);
not NOT1 (N4665, N4649);
and AND3 (N4666, N4661, N3686, N1178);
nand NAND3 (N4667, N4657, N2094, N666);
nor NOR3 (N4668, N4662, N2714, N3033);
or OR4 (N4669, N4665, N534, N390, N2569);
and AND2 (N4670, N4669, N2205);
and AND4 (N4671, N4653, N2802, N3022, N3958);
buf BUF1 (N4672, N4641);
not NOT1 (N4673, N4668);
xor XOR2 (N4674, N4672, N3469);
xor XOR2 (N4675, N4633, N2926);
buf BUF1 (N4676, N4674);
nand NAND4 (N4677, N4667, N3126, N3074, N700);
nand NAND4 (N4678, N4671, N644, N1164, N2001);
or OR2 (N4679, N4676, N1718);
buf BUF1 (N4680, N4679);
nor NOR4 (N4681, N4659, N1557, N1605, N3764);
nand NAND3 (N4682, N4680, N2000, N1464);
nand NAND2 (N4683, N4664, N3028);
buf BUF1 (N4684, N4670);
and AND4 (N4685, N4675, N928, N1381, N1685);
buf BUF1 (N4686, N4673);
not NOT1 (N4687, N4663);
xor XOR2 (N4688, N4678, N2544);
nand NAND4 (N4689, N4666, N2311, N3069, N3159);
or OR2 (N4690, N4689, N4625);
not NOT1 (N4691, N4682);
buf BUF1 (N4692, N4683);
not NOT1 (N4693, N4681);
and AND3 (N4694, N4691, N1041, N950);
not NOT1 (N4695, N4690);
xor XOR2 (N4696, N4687, N1464);
buf BUF1 (N4697, N4684);
or OR4 (N4698, N4685, N2161, N3329, N2869);
buf BUF1 (N4699, N4694);
and AND3 (N4700, N4696, N4026, N3806);
and AND3 (N4701, N4688, N2095, N700);
nor NOR2 (N4702, N4693, N3365);
xor XOR2 (N4703, N4699, N3745);
xor XOR2 (N4704, N4677, N2771);
nand NAND2 (N4705, N4700, N612);
xor XOR2 (N4706, N4695, N806);
and AND3 (N4707, N4686, N3213, N4432);
nand NAND2 (N4708, N4702, N3662);
nand NAND2 (N4709, N4704, N584);
and AND2 (N4710, N4692, N4126);
buf BUF1 (N4711, N4705);
buf BUF1 (N4712, N4703);
nor NOR4 (N4713, N4698, N1815, N2771, N3568);
and AND4 (N4714, N4709, N556, N4073, N4358);
nor NOR3 (N4715, N4708, N1883, N4444);
or OR3 (N4716, N4706, N1973, N1901);
nand NAND4 (N4717, N4713, N1177, N2762, N4124);
buf BUF1 (N4718, N4717);
nor NOR3 (N4719, N4718, N3666, N2283);
and AND4 (N4720, N4714, N4505, N78, N2573);
xor XOR2 (N4721, N4710, N3613);
buf BUF1 (N4722, N4721);
nand NAND3 (N4723, N4707, N4703, N1102);
not NOT1 (N4724, N4723);
buf BUF1 (N4725, N4715);
nand NAND4 (N4726, N4701, N998, N1883, N1946);
buf BUF1 (N4727, N4712);
not NOT1 (N4728, N4726);
nand NAND2 (N4729, N4727, N3491);
not NOT1 (N4730, N4697);
nand NAND4 (N4731, N4729, N460, N549, N1255);
xor XOR2 (N4732, N4731, N4525);
nor NOR2 (N4733, N4725, N3159);
or OR4 (N4734, N4728, N379, N3003, N128);
nand NAND4 (N4735, N4732, N3912, N710, N4224);
nand NAND2 (N4736, N4734, N4260);
buf BUF1 (N4737, N4711);
buf BUF1 (N4738, N4722);
and AND4 (N4739, N4738, N2051, N4576, N2528);
buf BUF1 (N4740, N4737);
nand NAND3 (N4741, N4720, N3931, N3592);
buf BUF1 (N4742, N4739);
or OR2 (N4743, N4736, N4533);
or OR3 (N4744, N4741, N4043, N1302);
or OR2 (N4745, N4735, N49);
buf BUF1 (N4746, N4730);
nor NOR4 (N4747, N4719, N3695, N3686, N2356);
and AND2 (N4748, N4743, N1310);
nor NOR4 (N4749, N4746, N582, N1765, N28);
and AND3 (N4750, N4749, N1146, N41);
and AND2 (N4751, N4740, N3127);
buf BUF1 (N4752, N4742);
buf BUF1 (N4753, N4724);
nor NOR2 (N4754, N4748, N4583);
buf BUF1 (N4755, N4750);
and AND2 (N4756, N4755, N4518);
and AND4 (N4757, N4752, N3482, N2046, N100);
or OR4 (N4758, N4744, N1751, N1317, N746);
not NOT1 (N4759, N4733);
and AND2 (N4760, N4745, N3998);
nand NAND3 (N4761, N4716, N2308, N3171);
nor NOR3 (N4762, N4747, N238, N791);
buf BUF1 (N4763, N4757);
nor NOR3 (N4764, N4753, N3652, N4763);
nor NOR3 (N4765, N2714, N3952, N642);
xor XOR2 (N4766, N4756, N1081);
or OR2 (N4767, N4760, N1673);
nor NOR4 (N4768, N4767, N4595, N4566, N2532);
and AND3 (N4769, N4751, N3065, N2777);
nor NOR2 (N4770, N4765, N2849);
or OR4 (N4771, N4768, N3756, N650, N3078);
not NOT1 (N4772, N4770);
xor XOR2 (N4773, N4769, N3516);
or OR4 (N4774, N4758, N1357, N4745, N2574);
or OR3 (N4775, N4761, N2608, N3694);
or OR2 (N4776, N4773, N807);
xor XOR2 (N4777, N4764, N1847);
not NOT1 (N4778, N4772);
not NOT1 (N4779, N4775);
and AND3 (N4780, N4774, N319, N105);
buf BUF1 (N4781, N4771);
nor NOR2 (N4782, N4777, N2993);
nor NOR3 (N4783, N4780, N399, N2141);
or OR2 (N4784, N4779, N4232);
nor NOR2 (N4785, N4759, N2130);
and AND4 (N4786, N4785, N2294, N4474, N2827);
xor XOR2 (N4787, N4784, N2952);
or OR2 (N4788, N4783, N658);
buf BUF1 (N4789, N4776);
and AND3 (N4790, N4781, N4590, N2734);
or OR2 (N4791, N4778, N3416);
nor NOR4 (N4792, N4789, N2633, N3884, N1481);
not NOT1 (N4793, N4762);
not NOT1 (N4794, N4788);
and AND2 (N4795, N4790, N2926);
or OR3 (N4796, N4792, N119, N1357);
and AND4 (N4797, N4766, N2132, N880, N4239);
not NOT1 (N4798, N4795);
or OR2 (N4799, N4794, N2666);
or OR3 (N4800, N4754, N1196, N3438);
nand NAND4 (N4801, N4796, N4287, N4646, N3779);
buf BUF1 (N4802, N4782);
nand NAND2 (N4803, N4802, N2040);
nor NOR3 (N4804, N4787, N1372, N1980);
not NOT1 (N4805, N4791);
not NOT1 (N4806, N4805);
or OR3 (N4807, N4806, N2849, N3308);
nor NOR4 (N4808, N4797, N2354, N1096, N2180);
not NOT1 (N4809, N4799);
nand NAND2 (N4810, N4793, N2401);
not NOT1 (N4811, N4786);
buf BUF1 (N4812, N4803);
nor NOR3 (N4813, N4801, N2017, N74);
xor XOR2 (N4814, N4811, N3445);
and AND4 (N4815, N4813, N4526, N4617, N1716);
nor NOR3 (N4816, N4804, N3465, N139);
or OR2 (N4817, N4800, N1375);
buf BUF1 (N4818, N4810);
xor XOR2 (N4819, N4817, N4729);
nand NAND3 (N4820, N4815, N3213, N1573);
xor XOR2 (N4821, N4798, N1348);
xor XOR2 (N4822, N4820, N3337);
xor XOR2 (N4823, N4808, N4020);
xor XOR2 (N4824, N4816, N2799);
buf BUF1 (N4825, N4821);
not NOT1 (N4826, N4812);
and AND3 (N4827, N4823, N4526, N3870);
not NOT1 (N4828, N4825);
not NOT1 (N4829, N4819);
buf BUF1 (N4830, N4814);
buf BUF1 (N4831, N4827);
not NOT1 (N4832, N4828);
nand NAND2 (N4833, N4829, N4665);
buf BUF1 (N4834, N4832);
or OR2 (N4835, N4809, N3980);
buf BUF1 (N4836, N4826);
buf BUF1 (N4837, N4831);
nor NOR4 (N4838, N4807, N1953, N3180, N3914);
nand NAND3 (N4839, N4830, N4163, N1065);
or OR2 (N4840, N4822, N3447);
or OR3 (N4841, N4818, N3432, N4770);
not NOT1 (N4842, N4838);
nor NOR4 (N4843, N4836, N293, N1708, N4284);
or OR4 (N4844, N4834, N3834, N4755, N348);
or OR3 (N4845, N4840, N2342, N343);
or OR3 (N4846, N4835, N2427, N3455);
nand NAND3 (N4847, N4846, N342, N474);
and AND3 (N4848, N4837, N52, N790);
buf BUF1 (N4849, N4824);
nor NOR4 (N4850, N4849, N4204, N1676, N3510);
or OR2 (N4851, N4848, N105);
xor XOR2 (N4852, N4843, N4149);
not NOT1 (N4853, N4833);
buf BUF1 (N4854, N4841);
buf BUF1 (N4855, N4851);
not NOT1 (N4856, N4844);
and AND2 (N4857, N4847, N3036);
xor XOR2 (N4858, N4839, N4556);
buf BUF1 (N4859, N4856);
or OR4 (N4860, N4858, N4698, N1945, N2845);
or OR3 (N4861, N4857, N1558, N4318);
buf BUF1 (N4862, N4853);
xor XOR2 (N4863, N4862, N4142);
or OR4 (N4864, N4842, N4075, N4450, N1311);
nor NOR2 (N4865, N4850, N2632);
and AND2 (N4866, N4855, N3405);
and AND3 (N4867, N4854, N1761, N3616);
nor NOR3 (N4868, N4860, N1615, N2828);
xor XOR2 (N4869, N4859, N3895);
or OR3 (N4870, N4866, N430, N2318);
not NOT1 (N4871, N4868);
and AND4 (N4872, N4845, N1916, N2225, N3028);
and AND4 (N4873, N4867, N4853, N1571, N3416);
nor NOR4 (N4874, N4861, N1837, N1562, N3995);
nand NAND4 (N4875, N4852, N3010, N895, N2007);
xor XOR2 (N4876, N4871, N4321);
buf BUF1 (N4877, N4873);
or OR3 (N4878, N4875, N1080, N448);
nor NOR4 (N4879, N4864, N96, N3620, N4708);
nor NOR4 (N4880, N4869, N4678, N1017, N79);
or OR4 (N4881, N4863, N212, N2891, N3000);
not NOT1 (N4882, N4872);
buf BUF1 (N4883, N4865);
nor NOR3 (N4884, N4876, N727, N1235);
not NOT1 (N4885, N4881);
buf BUF1 (N4886, N4882);
xor XOR2 (N4887, N4870, N210);
or OR4 (N4888, N4883, N2846, N3836, N2839);
xor XOR2 (N4889, N4880, N436);
nor NOR3 (N4890, N4887, N4845, N2355);
not NOT1 (N4891, N4884);
and AND2 (N4892, N4878, N416);
xor XOR2 (N4893, N4885, N1008);
buf BUF1 (N4894, N4886);
nand NAND3 (N4895, N4889, N4202, N1054);
and AND2 (N4896, N4893, N4309);
xor XOR2 (N4897, N4890, N4581);
nor NOR4 (N4898, N4891, N2938, N335, N1175);
nand NAND3 (N4899, N4879, N1815, N2938);
and AND2 (N4900, N4897, N725);
xor XOR2 (N4901, N4892, N1387);
nand NAND3 (N4902, N4895, N1555, N4692);
nor NOR3 (N4903, N4899, N3521, N2398);
buf BUF1 (N4904, N4898);
not NOT1 (N4905, N4904);
or OR2 (N4906, N4902, N1499);
not NOT1 (N4907, N4874);
or OR4 (N4908, N4905, N3706, N2188, N4489);
not NOT1 (N4909, N4901);
nand NAND3 (N4910, N4894, N1104, N4752);
xor XOR2 (N4911, N4896, N2547);
nand NAND4 (N4912, N4910, N2581, N3829, N2654);
and AND2 (N4913, N4907, N2163);
nor NOR2 (N4914, N4913, N2785);
xor XOR2 (N4915, N4914, N1726);
nand NAND4 (N4916, N4909, N1988, N1252, N6);
nor NOR3 (N4917, N4888, N2283, N966);
xor XOR2 (N4918, N4903, N2890);
or OR3 (N4919, N4877, N1566, N641);
not NOT1 (N4920, N4911);
buf BUF1 (N4921, N4900);
buf BUF1 (N4922, N4919);
or OR2 (N4923, N4916, N2205);
or OR3 (N4924, N4922, N915, N3389);
nand NAND3 (N4925, N4908, N3925, N1761);
not NOT1 (N4926, N4925);
buf BUF1 (N4927, N4917);
and AND2 (N4928, N4923, N533);
not NOT1 (N4929, N4924);
and AND2 (N4930, N4927, N4386);
nor NOR2 (N4931, N4926, N1138);
buf BUF1 (N4932, N4921);
nand NAND4 (N4933, N4930, N1006, N3088, N457);
nor NOR4 (N4934, N4929, N638, N677, N4835);
or OR2 (N4935, N4932, N1606);
xor XOR2 (N4936, N4934, N4155);
or OR3 (N4937, N4936, N4329, N475);
nand NAND3 (N4938, N4928, N4588, N3336);
not NOT1 (N4939, N4931);
nor NOR4 (N4940, N4920, N3709, N1826, N212);
not NOT1 (N4941, N4906);
buf BUF1 (N4942, N4912);
nor NOR3 (N4943, N4942, N1601, N309);
buf BUF1 (N4944, N4915);
xor XOR2 (N4945, N4935, N4801);
not NOT1 (N4946, N4940);
not NOT1 (N4947, N4941);
nand NAND3 (N4948, N4945, N839, N851);
nor NOR3 (N4949, N4947, N566, N387);
and AND2 (N4950, N4944, N2742);
and AND4 (N4951, N4943, N3677, N2099, N610);
nand NAND2 (N4952, N4933, N4287);
not NOT1 (N4953, N4946);
and AND4 (N4954, N4953, N1065, N6, N2712);
and AND3 (N4955, N4938, N929, N2731);
or OR4 (N4956, N4949, N1287, N4880, N4107);
nor NOR4 (N4957, N4939, N400, N3443, N3646);
and AND4 (N4958, N4950, N971, N2657, N435);
or OR3 (N4959, N4918, N3979, N199);
xor XOR2 (N4960, N4937, N3046);
buf BUF1 (N4961, N4959);
xor XOR2 (N4962, N4957, N2530);
xor XOR2 (N4963, N4956, N1377);
buf BUF1 (N4964, N4948);
not NOT1 (N4965, N4962);
nand NAND2 (N4966, N4955, N3928);
not NOT1 (N4967, N4963);
or OR2 (N4968, N4964, N1685);
nand NAND4 (N4969, N4952, N1968, N3551, N4882);
not NOT1 (N4970, N4954);
xor XOR2 (N4971, N4970, N678);
buf BUF1 (N4972, N4968);
nor NOR3 (N4973, N4971, N3683, N1940);
not NOT1 (N4974, N4973);
nor NOR2 (N4975, N4966, N3380);
or OR4 (N4976, N4961, N4046, N2304, N880);
or OR4 (N4977, N4974, N2583, N2192, N2683);
or OR3 (N4978, N4975, N4086, N341);
nand NAND4 (N4979, N4969, N4188, N1782, N1041);
and AND2 (N4980, N4979, N2656);
buf BUF1 (N4981, N4978);
nand NAND4 (N4982, N4967, N4591, N2656, N144);
and AND3 (N4983, N4981, N3453, N1095);
buf BUF1 (N4984, N4983);
buf BUF1 (N4985, N4951);
and AND2 (N4986, N4985, N3937);
or OR2 (N4987, N4977, N661);
nand NAND3 (N4988, N4982, N4446, N3530);
or OR3 (N4989, N4987, N3833, N4408);
or OR3 (N4990, N4989, N4665, N1679);
xor XOR2 (N4991, N4965, N2810);
and AND3 (N4992, N4972, N4928, N4206);
nor NOR3 (N4993, N4958, N3531, N3337);
nor NOR3 (N4994, N4986, N4929, N714);
and AND2 (N4995, N4984, N4806);
nor NOR4 (N4996, N4992, N2479, N1424, N2897);
or OR2 (N4997, N4995, N3813);
and AND4 (N4998, N4980, N1087, N643, N1562);
xor XOR2 (N4999, N4991, N2107);
not NOT1 (N5000, N4976);
nor NOR4 (N5001, N4990, N2562, N1576, N4555);
xor XOR2 (N5002, N5000, N1446);
buf BUF1 (N5003, N4988);
nand NAND2 (N5004, N4960, N4913);
and AND4 (N5005, N4993, N1751, N49, N2466);
nor NOR3 (N5006, N5005, N549, N2991);
nor NOR4 (N5007, N4996, N3198, N4521, N4515);
or OR4 (N5008, N5007, N4587, N2755, N3000);
buf BUF1 (N5009, N5006);
nor NOR4 (N5010, N4998, N749, N711, N4806);
or OR3 (N5011, N5010, N3861, N1967);
or OR3 (N5012, N5002, N630, N1719);
nor NOR4 (N5013, N5001, N2284, N727, N910);
buf BUF1 (N5014, N5004);
xor XOR2 (N5015, N5009, N3879);
nand NAND3 (N5016, N5012, N3043, N2611);
not NOT1 (N5017, N5003);
not NOT1 (N5018, N5013);
nand NAND2 (N5019, N4999, N280);
nand NAND4 (N5020, N5019, N3448, N1242, N4802);
nor NOR2 (N5021, N5016, N2343);
not NOT1 (N5022, N5020);
nand NAND2 (N5023, N5021, N1292);
and AND4 (N5024, N5008, N2241, N2326, N1308);
and AND4 (N5025, N5024, N21, N1911, N606);
not NOT1 (N5026, N5017);
nand NAND3 (N5027, N5022, N3192, N808);
not NOT1 (N5028, N5025);
and AND4 (N5029, N5015, N1116, N4475, N445);
buf BUF1 (N5030, N5027);
xor XOR2 (N5031, N5014, N3012);
or OR4 (N5032, N5026, N851, N3010, N3582);
and AND3 (N5033, N5018, N98, N4165);
not NOT1 (N5034, N5023);
nor NOR2 (N5035, N4994, N3212);
not NOT1 (N5036, N5011);
nand NAND3 (N5037, N5033, N514, N1217);
or OR4 (N5038, N5036, N4421, N476, N2029);
nor NOR4 (N5039, N5037, N485, N4160, N844);
not NOT1 (N5040, N5034);
or OR4 (N5041, N5030, N3014, N2367, N2621);
nand NAND2 (N5042, N5035, N4266);
nor NOR2 (N5043, N5031, N2197);
buf BUF1 (N5044, N5042);
buf BUF1 (N5045, N5041);
nor NOR3 (N5046, N5043, N4365, N2699);
and AND4 (N5047, N5039, N2671, N2764, N4505);
not NOT1 (N5048, N5046);
nand NAND4 (N5049, N5044, N4435, N2272, N3065);
buf BUF1 (N5050, N5048);
and AND4 (N5051, N5038, N1210, N264, N1357);
and AND3 (N5052, N5047, N132, N4547);
nand NAND2 (N5053, N4997, N1530);
nor NOR4 (N5054, N5051, N1163, N3614, N3065);
nand NAND3 (N5055, N5053, N3680, N4629);
xor XOR2 (N5056, N5054, N3925);
or OR2 (N5057, N5050, N3968);
nand NAND4 (N5058, N5055, N899, N3278, N1000);
and AND3 (N5059, N5058, N4205, N2972);
xor XOR2 (N5060, N5032, N4172);
not NOT1 (N5061, N5060);
nand NAND2 (N5062, N5040, N4660);
nand NAND4 (N5063, N5029, N662, N4081, N4838);
xor XOR2 (N5064, N5045, N985);
or OR4 (N5065, N5049, N167, N3453, N166);
xor XOR2 (N5066, N5063, N2082);
nand NAND3 (N5067, N5061, N1179, N918);
nand NAND2 (N5068, N5066, N2081);
buf BUF1 (N5069, N5059);
nand NAND4 (N5070, N5065, N161, N2970, N1910);
and AND3 (N5071, N5062, N2480, N3607);
nor NOR2 (N5072, N5064, N1873);
and AND4 (N5073, N5070, N838, N853, N1083);
not NOT1 (N5074, N5069);
nand NAND3 (N5075, N5073, N3993, N3579);
xor XOR2 (N5076, N5072, N2240);
buf BUF1 (N5077, N5056);
not NOT1 (N5078, N5077);
nand NAND4 (N5079, N5057, N459, N3123, N351);
or OR4 (N5080, N5067, N2891, N3966, N698);
buf BUF1 (N5081, N5068);
and AND3 (N5082, N5052, N642, N3168);
nand NAND3 (N5083, N5078, N1635, N400);
nand NAND3 (N5084, N5082, N2023, N1301);
and AND4 (N5085, N5028, N3137, N1821, N10);
or OR4 (N5086, N5080, N1292, N549, N4845);
or OR3 (N5087, N5071, N3344, N855);
nand NAND4 (N5088, N5087, N3769, N1118, N2753);
xor XOR2 (N5089, N5085, N230);
buf BUF1 (N5090, N5081);
or OR3 (N5091, N5083, N3556, N4401);
and AND3 (N5092, N5074, N3782, N2657);
xor XOR2 (N5093, N5089, N1774);
or OR4 (N5094, N5092, N1327, N2394, N2812);
buf BUF1 (N5095, N5086);
or OR2 (N5096, N5079, N4628);
nor NOR2 (N5097, N5091, N2106);
not NOT1 (N5098, N5095);
xor XOR2 (N5099, N5093, N870);
nor NOR4 (N5100, N5075, N260, N2116, N4608);
buf BUF1 (N5101, N5094);
xor XOR2 (N5102, N5088, N4447);
xor XOR2 (N5103, N5099, N1364);
not NOT1 (N5104, N5103);
nor NOR2 (N5105, N5090, N1348);
xor XOR2 (N5106, N5100, N4203);
nor NOR4 (N5107, N5084, N1807, N4092, N1251);
xor XOR2 (N5108, N5107, N2119);
xor XOR2 (N5109, N5102, N1802);
buf BUF1 (N5110, N5104);
or OR3 (N5111, N5105, N4882, N80);
nand NAND4 (N5112, N5109, N2003, N1498, N1660);
nand NAND3 (N5113, N5111, N5109, N3488);
xor XOR2 (N5114, N5076, N4103);
nor NOR2 (N5115, N5106, N4527);
buf BUF1 (N5116, N5101);
or OR4 (N5117, N5108, N1035, N3949, N3423);
nor NOR2 (N5118, N5116, N2277);
nor NOR3 (N5119, N5096, N4376, N865);
nand NAND4 (N5120, N5113, N4349, N1058, N1543);
xor XOR2 (N5121, N5118, N1476);
not NOT1 (N5122, N5115);
or OR4 (N5123, N5110, N336, N150, N3695);
nand NAND4 (N5124, N5122, N2665, N2734, N1510);
or OR2 (N5125, N5117, N1279);
not NOT1 (N5126, N5119);
or OR2 (N5127, N5097, N4111);
nor NOR3 (N5128, N5120, N2062, N2621);
or OR4 (N5129, N5114, N501, N1350, N873);
and AND4 (N5130, N5098, N3755, N3809, N4677);
xor XOR2 (N5131, N5127, N164);
nand NAND4 (N5132, N5131, N2104, N3727, N968);
nand NAND4 (N5133, N5128, N5129, N2932, N3365);
and AND2 (N5134, N4111, N13);
buf BUF1 (N5135, N5121);
not NOT1 (N5136, N5125);
nand NAND4 (N5137, N5132, N3782, N4259, N699);
or OR3 (N5138, N5130, N45, N4557);
not NOT1 (N5139, N5137);
or OR2 (N5140, N5138, N686);
not NOT1 (N5141, N5139);
not NOT1 (N5142, N5136);
buf BUF1 (N5143, N5141);
xor XOR2 (N5144, N5140, N2428);
not NOT1 (N5145, N5134);
buf BUF1 (N5146, N5123);
or OR2 (N5147, N5126, N2137);
nand NAND3 (N5148, N5124, N3347, N2313);
or OR4 (N5149, N5133, N2382, N2573, N863);
xor XOR2 (N5150, N5147, N1182);
xor XOR2 (N5151, N5148, N4652);
buf BUF1 (N5152, N5149);
and AND3 (N5153, N5135, N4127, N2541);
buf BUF1 (N5154, N5150);
not NOT1 (N5155, N5144);
not NOT1 (N5156, N5112);
and AND2 (N5157, N5143, N4909);
nand NAND2 (N5158, N5155, N2877);
nand NAND3 (N5159, N5145, N3855, N2679);
or OR3 (N5160, N5142, N4351, N1241);
nand NAND2 (N5161, N5157, N3599);
nand NAND3 (N5162, N5151, N3413, N4571);
buf BUF1 (N5163, N5159);
nand NAND2 (N5164, N5153, N892);
not NOT1 (N5165, N5160);
or OR2 (N5166, N5152, N1806);
nand NAND3 (N5167, N5165, N3768, N1018);
xor XOR2 (N5168, N5162, N5036);
xor XOR2 (N5169, N5168, N2839);
nand NAND2 (N5170, N5164, N2108);
and AND3 (N5171, N5146, N2852, N2863);
not NOT1 (N5172, N5169);
xor XOR2 (N5173, N5163, N5120);
nor NOR3 (N5174, N5161, N4697, N1639);
or OR2 (N5175, N5170, N1963);
buf BUF1 (N5176, N5158);
not NOT1 (N5177, N5156);
nor NOR3 (N5178, N5167, N1203, N2397);
nand NAND2 (N5179, N5171, N3009);
buf BUF1 (N5180, N5174);
and AND3 (N5181, N5179, N1454, N302);
nor NOR2 (N5182, N5175, N3887);
xor XOR2 (N5183, N5177, N4830);
buf BUF1 (N5184, N5181);
nand NAND2 (N5185, N5172, N5088);
and AND3 (N5186, N5185, N626, N1335);
buf BUF1 (N5187, N5154);
nor NOR4 (N5188, N5186, N4615, N1468, N3005);
nor NOR4 (N5189, N5184, N1113, N205, N3090);
xor XOR2 (N5190, N5166, N3638);
or OR4 (N5191, N5182, N3688, N1868, N329);
or OR4 (N5192, N5191, N5043, N1215, N1906);
xor XOR2 (N5193, N5173, N2980);
not NOT1 (N5194, N5187);
xor XOR2 (N5195, N5188, N3578);
nand NAND2 (N5196, N5183, N3790);
and AND3 (N5197, N5180, N2547, N2422);
and AND3 (N5198, N5197, N4711, N141);
buf BUF1 (N5199, N5195);
or OR3 (N5200, N5192, N3107, N2974);
and AND4 (N5201, N5194, N3890, N3860, N3470);
or OR3 (N5202, N5176, N4629, N2693);
or OR4 (N5203, N5199, N1264, N2390, N4741);
nand NAND2 (N5204, N5189, N2896);
or OR4 (N5205, N5196, N2137, N3791, N4818);
not NOT1 (N5206, N5204);
nor NOR4 (N5207, N5201, N4636, N2136, N2606);
xor XOR2 (N5208, N5207, N1837);
xor XOR2 (N5209, N5205, N1758);
xor XOR2 (N5210, N5203, N758);
or OR2 (N5211, N5202, N1546);
or OR2 (N5212, N5178, N1848);
nor NOR4 (N5213, N5212, N4290, N4500, N4057);
xor XOR2 (N5214, N5208, N4878);
or OR2 (N5215, N5190, N1683);
xor XOR2 (N5216, N5210, N474);
xor XOR2 (N5217, N5213, N966);
nor NOR2 (N5218, N5206, N766);
xor XOR2 (N5219, N5198, N4767);
not NOT1 (N5220, N5214);
xor XOR2 (N5221, N5193, N4582);
nor NOR2 (N5222, N5211, N4125);
nand NAND3 (N5223, N5215, N4206, N2739);
buf BUF1 (N5224, N5220);
and AND2 (N5225, N5221, N4715);
nor NOR4 (N5226, N5209, N3637, N1663, N4513);
xor XOR2 (N5227, N5218, N3439);
nand NAND4 (N5228, N5222, N3550, N1215, N2226);
xor XOR2 (N5229, N5224, N3195);
nand NAND4 (N5230, N5227, N5015, N2628, N4430);
or OR3 (N5231, N5229, N4644, N3049);
xor XOR2 (N5232, N5223, N1572);
and AND2 (N5233, N5217, N1717);
xor XOR2 (N5234, N5219, N1533);
buf BUF1 (N5235, N5231);
xor XOR2 (N5236, N5233, N4483);
xor XOR2 (N5237, N5236, N1101);
nand NAND2 (N5238, N5226, N1079);
and AND3 (N5239, N5228, N2948, N3236);
buf BUF1 (N5240, N5230);
not NOT1 (N5241, N5200);
buf BUF1 (N5242, N5216);
buf BUF1 (N5243, N5232);
xor XOR2 (N5244, N5239, N4898);
nor NOR4 (N5245, N5238, N4220, N3586, N466);
not NOT1 (N5246, N5237);
xor XOR2 (N5247, N5234, N3014);
not NOT1 (N5248, N5245);
or OR2 (N5249, N5246, N1700);
not NOT1 (N5250, N5242);
and AND4 (N5251, N5247, N1243, N2957, N410);
xor XOR2 (N5252, N5248, N4780);
nor NOR4 (N5253, N5240, N933, N4276, N1541);
nor NOR2 (N5254, N5241, N4289);
and AND4 (N5255, N5235, N3574, N2972, N3708);
and AND3 (N5256, N5253, N4934, N3453);
or OR4 (N5257, N5249, N1492, N3848, N1798);
not NOT1 (N5258, N5243);
not NOT1 (N5259, N5254);
xor XOR2 (N5260, N5258, N273);
buf BUF1 (N5261, N5260);
nand NAND3 (N5262, N5257, N567, N1120);
not NOT1 (N5263, N5225);
and AND2 (N5264, N5255, N1117);
and AND3 (N5265, N5264, N157, N3380);
buf BUF1 (N5266, N5259);
not NOT1 (N5267, N5261);
xor XOR2 (N5268, N5263, N1813);
not NOT1 (N5269, N5268);
not NOT1 (N5270, N5251);
not NOT1 (N5271, N5244);
or OR2 (N5272, N5269, N2295);
and AND4 (N5273, N5266, N1896, N2575, N4924);
not NOT1 (N5274, N5271);
buf BUF1 (N5275, N5252);
and AND2 (N5276, N5265, N315);
nand NAND3 (N5277, N5272, N445, N3999);
and AND4 (N5278, N5273, N4948, N763, N717);
not NOT1 (N5279, N5274);
xor XOR2 (N5280, N5270, N4758);
xor XOR2 (N5281, N5262, N1224);
nand NAND4 (N5282, N5276, N377, N2469, N1286);
nand NAND4 (N5283, N5279, N4057, N1307, N5068);
not NOT1 (N5284, N5256);
and AND4 (N5285, N5280, N2361, N1699, N785);
not NOT1 (N5286, N5283);
or OR2 (N5287, N5275, N3521);
nand NAND3 (N5288, N5267, N1506, N5149);
or OR2 (N5289, N5250, N885);
buf BUF1 (N5290, N5285);
nor NOR3 (N5291, N5277, N490, N626);
xor XOR2 (N5292, N5288, N4045);
not NOT1 (N5293, N5281);
nor NOR2 (N5294, N5286, N3662);
nor NOR4 (N5295, N5293, N472, N1622, N3600);
nor NOR4 (N5296, N5292, N3201, N277, N599);
nor NOR4 (N5297, N5278, N4576, N3169, N3922);
and AND3 (N5298, N5289, N1080, N2571);
nand NAND3 (N5299, N5291, N818, N2575);
and AND4 (N5300, N5299, N2192, N3943, N4157);
buf BUF1 (N5301, N5282);
and AND3 (N5302, N5287, N2255, N4735);
or OR2 (N5303, N5284, N3130);
or OR4 (N5304, N5302, N733, N2853, N1996);
nor NOR3 (N5305, N5297, N4052, N4071);
nor NOR4 (N5306, N5290, N2167, N5010, N2761);
buf BUF1 (N5307, N5296);
not NOT1 (N5308, N5304);
buf BUF1 (N5309, N5303);
or OR2 (N5310, N5306, N4148);
and AND3 (N5311, N5295, N559, N3034);
nor NOR2 (N5312, N5310, N1478);
and AND4 (N5313, N5298, N2940, N2933, N2444);
and AND2 (N5314, N5307, N614);
and AND3 (N5315, N5294, N4010, N1087);
not NOT1 (N5316, N5308);
nor NOR2 (N5317, N5309, N4803);
xor XOR2 (N5318, N5316, N2320);
xor XOR2 (N5319, N5317, N4635);
or OR2 (N5320, N5313, N4480);
nand NAND2 (N5321, N5300, N4330);
not NOT1 (N5322, N5315);
xor XOR2 (N5323, N5311, N1316);
not NOT1 (N5324, N5314);
and AND3 (N5325, N5323, N4211, N402);
and AND4 (N5326, N5301, N2719, N4572, N233);
not NOT1 (N5327, N5324);
buf BUF1 (N5328, N5305);
or OR3 (N5329, N5326, N1413, N5017);
nand NAND4 (N5330, N5329, N996, N2871, N4625);
nand NAND4 (N5331, N5312, N940, N5152, N3718);
nor NOR4 (N5332, N5322, N4999, N2921, N3133);
or OR3 (N5333, N5321, N1474, N5098);
xor XOR2 (N5334, N5327, N3885);
nand NAND3 (N5335, N5331, N1448, N2013);
xor XOR2 (N5336, N5320, N4088);
nand NAND2 (N5337, N5325, N2756);
not NOT1 (N5338, N5337);
xor XOR2 (N5339, N5334, N3714);
not NOT1 (N5340, N5339);
xor XOR2 (N5341, N5318, N4413);
buf BUF1 (N5342, N5332);
and AND3 (N5343, N5338, N1021, N4947);
nor NOR4 (N5344, N5335, N5341, N2881, N2990);
or OR3 (N5345, N960, N1400, N2045);
nand NAND2 (N5346, N5344, N3663);
or OR4 (N5347, N5340, N5325, N4381, N2459);
nor NOR4 (N5348, N5328, N31, N2196, N2198);
xor XOR2 (N5349, N5319, N266);
xor XOR2 (N5350, N5333, N2570);
and AND2 (N5351, N5343, N675);
and AND3 (N5352, N5342, N4545, N3301);
and AND2 (N5353, N5336, N2450);
nand NAND4 (N5354, N5347, N5132, N499, N4215);
nand NAND4 (N5355, N5330, N3519, N5243, N3546);
or OR2 (N5356, N5354, N256);
and AND4 (N5357, N5346, N1942, N1939, N1955);
and AND2 (N5358, N5353, N2323);
and AND4 (N5359, N5357, N804, N1566, N517);
xor XOR2 (N5360, N5345, N3785);
and AND2 (N5361, N5351, N2532);
buf BUF1 (N5362, N5349);
nand NAND3 (N5363, N5356, N1590, N1160);
buf BUF1 (N5364, N5352);
nor NOR2 (N5365, N5362, N1215);
and AND2 (N5366, N5360, N2146);
xor XOR2 (N5367, N5364, N410);
buf BUF1 (N5368, N5366);
nor NOR3 (N5369, N5367, N1967, N5309);
or OR3 (N5370, N5365, N2018, N1606);
xor XOR2 (N5371, N5355, N2106);
and AND2 (N5372, N5370, N3887);
nor NOR2 (N5373, N5348, N1214);
xor XOR2 (N5374, N5350, N4617);
xor XOR2 (N5375, N5361, N1396);
nor NOR3 (N5376, N5372, N3791, N4676);
xor XOR2 (N5377, N5374, N1709);
not NOT1 (N5378, N5358);
or OR3 (N5379, N5363, N2306, N3970);
buf BUF1 (N5380, N5371);
and AND3 (N5381, N5373, N3203, N3049);
buf BUF1 (N5382, N5378);
not NOT1 (N5383, N5377);
and AND2 (N5384, N5381, N2684);
and AND2 (N5385, N5383, N830);
nand NAND4 (N5386, N5369, N3173, N2280, N3934);
buf BUF1 (N5387, N5385);
xor XOR2 (N5388, N5384, N4633);
nand NAND4 (N5389, N5375, N5287, N2155, N5073);
and AND4 (N5390, N5387, N4623, N1061, N621);
buf BUF1 (N5391, N5382);
nor NOR3 (N5392, N5380, N893, N2989);
xor XOR2 (N5393, N5376, N5330);
buf BUF1 (N5394, N5379);
not NOT1 (N5395, N5393);
or OR4 (N5396, N5394, N1129, N4888, N3478);
xor XOR2 (N5397, N5388, N3690);
not NOT1 (N5398, N5390);
buf BUF1 (N5399, N5386);
buf BUF1 (N5400, N5397);
not NOT1 (N5401, N5399);
xor XOR2 (N5402, N5401, N1308);
nand NAND2 (N5403, N5398, N5024);
nand NAND4 (N5404, N5402, N4368, N1239, N3399);
and AND4 (N5405, N5396, N1640, N3626, N4435);
not NOT1 (N5406, N5405);
and AND2 (N5407, N5406, N3448);
buf BUF1 (N5408, N5392);
not NOT1 (N5409, N5368);
xor XOR2 (N5410, N5404, N1081);
nor NOR2 (N5411, N5410, N1693);
not NOT1 (N5412, N5389);
nor NOR2 (N5413, N5412, N3472);
buf BUF1 (N5414, N5395);
and AND3 (N5415, N5400, N3686, N152);
xor XOR2 (N5416, N5407, N2424);
nand NAND2 (N5417, N5359, N4589);
nor NOR3 (N5418, N5415, N1830, N3094);
and AND3 (N5419, N5418, N1923, N1627);
nor NOR3 (N5420, N5413, N2298, N560);
nor NOR3 (N5421, N5416, N1478, N5029);
nand NAND3 (N5422, N5421, N3608, N887);
nor NOR3 (N5423, N5411, N4142, N800);
buf BUF1 (N5424, N5419);
buf BUF1 (N5425, N5403);
buf BUF1 (N5426, N5420);
nand NAND2 (N5427, N5414, N974);
not NOT1 (N5428, N5391);
not NOT1 (N5429, N5417);
buf BUF1 (N5430, N5425);
buf BUF1 (N5431, N5426);
xor XOR2 (N5432, N5424, N3393);
nor NOR2 (N5433, N5409, N3166);
nor NOR2 (N5434, N5427, N1523);
buf BUF1 (N5435, N5433);
not NOT1 (N5436, N5435);
or OR3 (N5437, N5436, N1059, N1807);
and AND3 (N5438, N5422, N5407, N2761);
nor NOR4 (N5439, N5432, N2753, N2208, N237);
xor XOR2 (N5440, N5431, N3066);
or OR2 (N5441, N5440, N4977);
xor XOR2 (N5442, N5423, N3249);
nand NAND3 (N5443, N5441, N3860, N998);
xor XOR2 (N5444, N5408, N3345);
xor XOR2 (N5445, N5439, N3197);
nand NAND4 (N5446, N5445, N2363, N5154, N4707);
or OR3 (N5447, N5429, N3836, N5215);
nor NOR4 (N5448, N5434, N575, N2850, N523);
buf BUF1 (N5449, N5446);
nand NAND3 (N5450, N5447, N1271, N4225);
xor XOR2 (N5451, N5438, N1441);
xor XOR2 (N5452, N5448, N2716);
and AND2 (N5453, N5452, N532);
not NOT1 (N5454, N5442);
buf BUF1 (N5455, N5444);
and AND2 (N5456, N5453, N2626);
xor XOR2 (N5457, N5428, N3627);
and AND4 (N5458, N5449, N5053, N3895, N482);
nor NOR4 (N5459, N5455, N4886, N2969, N4558);
nand NAND2 (N5460, N5450, N1999);
xor XOR2 (N5461, N5459, N484);
and AND3 (N5462, N5461, N1358, N2929);
xor XOR2 (N5463, N5437, N1436);
and AND3 (N5464, N5443, N3783, N2487);
not NOT1 (N5465, N5451);
or OR4 (N5466, N5460, N2079, N2490, N3209);
xor XOR2 (N5467, N5466, N507);
nor NOR4 (N5468, N5467, N4522, N1236, N743);
buf BUF1 (N5469, N5430);
and AND2 (N5470, N5468, N4035);
and AND4 (N5471, N5464, N4967, N4813, N2053);
xor XOR2 (N5472, N5465, N5200);
xor XOR2 (N5473, N5470, N4353);
not NOT1 (N5474, N5472);
nand NAND4 (N5475, N5473, N1464, N1149, N660);
nor NOR2 (N5476, N5463, N4631);
and AND4 (N5477, N5458, N4248, N155, N5213);
and AND2 (N5478, N5475, N2208);
xor XOR2 (N5479, N5457, N4235);
nor NOR2 (N5480, N5477, N2601);
xor XOR2 (N5481, N5462, N4285);
not NOT1 (N5482, N5476);
nor NOR3 (N5483, N5479, N2388, N1038);
nor NOR2 (N5484, N5480, N1254);
nor NOR2 (N5485, N5478, N5333);
buf BUF1 (N5486, N5454);
or OR3 (N5487, N5485, N445, N1364);
not NOT1 (N5488, N5469);
buf BUF1 (N5489, N5481);
or OR3 (N5490, N5487, N1208, N2236);
nor NOR3 (N5491, N5489, N3033, N4603);
nor NOR3 (N5492, N5488, N1053, N3318);
or OR2 (N5493, N5483, N5285);
and AND4 (N5494, N5492, N4824, N3905, N418);
nand NAND4 (N5495, N5474, N3853, N1776, N1385);
or OR2 (N5496, N5494, N1730);
nand NAND2 (N5497, N5495, N1088);
nand NAND3 (N5498, N5484, N3196, N3206);
buf BUF1 (N5499, N5490);
nand NAND2 (N5500, N5486, N3980);
or OR4 (N5501, N5496, N2365, N3688, N2457);
and AND4 (N5502, N5493, N1686, N4116, N1129);
not NOT1 (N5503, N5482);
xor XOR2 (N5504, N5502, N1154);
or OR3 (N5505, N5497, N859, N2823);
xor XOR2 (N5506, N5501, N2754);
not NOT1 (N5507, N5498);
not NOT1 (N5508, N5499);
nand NAND4 (N5509, N5491, N4487, N4114, N2188);
not NOT1 (N5510, N5507);
nand NAND4 (N5511, N5506, N2854, N117, N5043);
buf BUF1 (N5512, N5511);
and AND3 (N5513, N5500, N1479, N4456);
buf BUF1 (N5514, N5504);
xor XOR2 (N5515, N5514, N1391);
nor NOR4 (N5516, N5456, N4834, N2458, N1650);
not NOT1 (N5517, N5471);
buf BUF1 (N5518, N5503);
xor XOR2 (N5519, N5513, N3404);
not NOT1 (N5520, N5509);
nor NOR3 (N5521, N5512, N2083, N490);
xor XOR2 (N5522, N5516, N524);
buf BUF1 (N5523, N5515);
buf BUF1 (N5524, N5517);
nor NOR2 (N5525, N5522, N4993);
nor NOR4 (N5526, N5524, N5169, N4019, N2697);
and AND3 (N5527, N5505, N2796, N5221);
nor NOR4 (N5528, N5525, N2476, N5296, N4975);
not NOT1 (N5529, N5523);
nor NOR3 (N5530, N5529, N2360, N629);
not NOT1 (N5531, N5527);
and AND3 (N5532, N5518, N628, N1952);
and AND4 (N5533, N5508, N4577, N4352, N644);
not NOT1 (N5534, N5531);
nand NAND2 (N5535, N5528, N2563);
buf BUF1 (N5536, N5526);
not NOT1 (N5537, N5532);
nand NAND4 (N5538, N5530, N3972, N4631, N4432);
xor XOR2 (N5539, N5537, N1339);
nand NAND2 (N5540, N5539, N600);
or OR3 (N5541, N5519, N664, N3690);
nor NOR3 (N5542, N5510, N4693, N2007);
or OR4 (N5543, N5533, N2298, N4998, N5221);
or OR2 (N5544, N5534, N4311);
or OR4 (N5545, N5542, N4055, N3024, N4453);
nand NAND4 (N5546, N5538, N4187, N1456, N1796);
nand NAND4 (N5547, N5544, N4305, N4659, N2505);
xor XOR2 (N5548, N5545, N2217);
buf BUF1 (N5549, N5546);
nand NAND3 (N5550, N5547, N2174, N908);
buf BUF1 (N5551, N5541);
or OR4 (N5552, N5543, N1007, N270, N1581);
buf BUF1 (N5553, N5550);
buf BUF1 (N5554, N5521);
not NOT1 (N5555, N5535);
xor XOR2 (N5556, N5553, N5157);
xor XOR2 (N5557, N5536, N5109);
xor XOR2 (N5558, N5554, N17);
buf BUF1 (N5559, N5520);
and AND3 (N5560, N5540, N2272, N593);
and AND3 (N5561, N5555, N664, N3397);
nor NOR3 (N5562, N5558, N335, N4947);
nand NAND4 (N5563, N5549, N3243, N2338, N214);
nor NOR2 (N5564, N5557, N4845);
or OR3 (N5565, N5548, N1094, N2032);
not NOT1 (N5566, N5551);
xor XOR2 (N5567, N5563, N3996);
or OR4 (N5568, N5567, N4578, N4221, N2203);
buf BUF1 (N5569, N5559);
not NOT1 (N5570, N5566);
buf BUF1 (N5571, N5560);
or OR3 (N5572, N5565, N2344, N838);
not NOT1 (N5573, N5552);
and AND4 (N5574, N5569, N996, N2549, N3128);
or OR4 (N5575, N5571, N1709, N965, N3633);
and AND2 (N5576, N5561, N602);
nand NAND4 (N5577, N5573, N3113, N4117, N3625);
not NOT1 (N5578, N5572);
buf BUF1 (N5579, N5576);
nand NAND3 (N5580, N5568, N320, N1861);
and AND3 (N5581, N5562, N3680, N3848);
and AND3 (N5582, N5575, N2092, N1930);
nor NOR2 (N5583, N5564, N4658);
not NOT1 (N5584, N5583);
xor XOR2 (N5585, N5570, N3136);
buf BUF1 (N5586, N5577);
xor XOR2 (N5587, N5584, N816);
xor XOR2 (N5588, N5581, N4435);
not NOT1 (N5589, N5578);
not NOT1 (N5590, N5579);
xor XOR2 (N5591, N5590, N4397);
nand NAND4 (N5592, N5587, N4746, N2981, N1071);
and AND4 (N5593, N5592, N2518, N5282, N5185);
not NOT1 (N5594, N5574);
or OR2 (N5595, N5582, N2385);
buf BUF1 (N5596, N5586);
buf BUF1 (N5597, N5588);
or OR3 (N5598, N5594, N2256, N4747);
nand NAND3 (N5599, N5596, N1058, N4124);
or OR2 (N5600, N5598, N4373);
xor XOR2 (N5601, N5593, N5440);
or OR2 (N5602, N5580, N4182);
buf BUF1 (N5603, N5556);
xor XOR2 (N5604, N5599, N1935);
nand NAND2 (N5605, N5601, N4442);
buf BUF1 (N5606, N5595);
nand NAND3 (N5607, N5600, N3574, N62);
xor XOR2 (N5608, N5589, N3779);
xor XOR2 (N5609, N5603, N105);
nand NAND2 (N5610, N5597, N2885);
not NOT1 (N5611, N5591);
xor XOR2 (N5612, N5611, N2176);
xor XOR2 (N5613, N5585, N2212);
xor XOR2 (N5614, N5604, N2690);
buf BUF1 (N5615, N5613);
or OR4 (N5616, N5615, N3875, N955, N4112);
buf BUF1 (N5617, N5602);
not NOT1 (N5618, N5609);
nand NAND3 (N5619, N5616, N254, N3225);
or OR2 (N5620, N5612, N3588);
and AND3 (N5621, N5617, N3459, N594);
or OR3 (N5622, N5621, N1622, N4187);
and AND2 (N5623, N5607, N4241);
not NOT1 (N5624, N5614);
nand NAND3 (N5625, N5620, N4188, N3527);
and AND2 (N5626, N5619, N5470);
xor XOR2 (N5627, N5626, N5545);
and AND4 (N5628, N5618, N1553, N5487, N1021);
and AND4 (N5629, N5608, N1026, N719, N926);
not NOT1 (N5630, N5610);
nand NAND4 (N5631, N5605, N3604, N5270, N2112);
and AND4 (N5632, N5624, N839, N1845, N1723);
buf BUF1 (N5633, N5623);
xor XOR2 (N5634, N5628, N4050);
xor XOR2 (N5635, N5633, N4393);
and AND4 (N5636, N5627, N1976, N4111, N4007);
not NOT1 (N5637, N5631);
not NOT1 (N5638, N5634);
or OR4 (N5639, N5630, N1563, N1790, N2552);
or OR3 (N5640, N5622, N5487, N2405);
not NOT1 (N5641, N5632);
or OR3 (N5642, N5638, N2285, N4728);
xor XOR2 (N5643, N5639, N2155);
or OR4 (N5644, N5637, N4652, N1940, N3318);
buf BUF1 (N5645, N5636);
or OR3 (N5646, N5645, N868, N4081);
or OR2 (N5647, N5635, N5464);
not NOT1 (N5648, N5647);
nor NOR4 (N5649, N5625, N1610, N1800, N457);
nand NAND2 (N5650, N5644, N2761);
xor XOR2 (N5651, N5648, N2663);
buf BUF1 (N5652, N5629);
not NOT1 (N5653, N5651);
xor XOR2 (N5654, N5650, N730);
or OR2 (N5655, N5649, N2079);
and AND4 (N5656, N5654, N1159, N4174, N179);
buf BUF1 (N5657, N5642);
nand NAND4 (N5658, N5643, N2357, N3584, N2157);
or OR4 (N5659, N5640, N3446, N1325, N4220);
nor NOR2 (N5660, N5655, N2457);
nand NAND2 (N5661, N5646, N4599);
xor XOR2 (N5662, N5657, N1741);
buf BUF1 (N5663, N5606);
or OR2 (N5664, N5652, N3876);
not NOT1 (N5665, N5660);
xor XOR2 (N5666, N5665, N3670);
xor XOR2 (N5667, N5656, N4242);
or OR2 (N5668, N5661, N864);
nor NOR4 (N5669, N5663, N2698, N4010, N2475);
and AND2 (N5670, N5668, N1219);
nand NAND2 (N5671, N5658, N2358);
or OR2 (N5672, N5659, N3249);
and AND3 (N5673, N5666, N1660, N5325);
xor XOR2 (N5674, N5672, N5371);
and AND2 (N5675, N5674, N3477);
and AND2 (N5676, N5662, N4050);
or OR4 (N5677, N5669, N602, N3761, N2635);
xor XOR2 (N5678, N5641, N364);
buf BUF1 (N5679, N5664);
and AND2 (N5680, N5667, N4955);
and AND3 (N5681, N5670, N4932, N4234);
buf BUF1 (N5682, N5671);
or OR2 (N5683, N5673, N1716);
xor XOR2 (N5684, N5653, N3645);
or OR2 (N5685, N5677, N814);
buf BUF1 (N5686, N5679);
and AND3 (N5687, N5680, N877, N1494);
not NOT1 (N5688, N5676);
nand NAND3 (N5689, N5682, N3120, N3834);
xor XOR2 (N5690, N5678, N380);
or OR4 (N5691, N5689, N1784, N2341, N3020);
nor NOR2 (N5692, N5688, N1951);
buf BUF1 (N5693, N5690);
and AND3 (N5694, N5687, N5263, N13);
nand NAND3 (N5695, N5693, N223, N5224);
not NOT1 (N5696, N5695);
not NOT1 (N5697, N5681);
xor XOR2 (N5698, N5675, N3300);
nor NOR4 (N5699, N5698, N1727, N721, N3434);
or OR2 (N5700, N5694, N1487);
xor XOR2 (N5701, N5691, N5059);
nor NOR3 (N5702, N5685, N2612, N2525);
not NOT1 (N5703, N5701);
nor NOR4 (N5704, N5686, N5303, N2236, N3154);
and AND2 (N5705, N5703, N3408);
and AND4 (N5706, N5684, N2944, N5638, N1402);
and AND3 (N5707, N5683, N4933, N984);
nor NOR4 (N5708, N5704, N2034, N3959, N951);
or OR4 (N5709, N5699, N2898, N2260, N2130);
and AND3 (N5710, N5708, N3437, N1728);
xor XOR2 (N5711, N5697, N1463);
nand NAND4 (N5712, N5711, N2193, N3872, N3477);
nand NAND3 (N5713, N5710, N1407, N2788);
xor XOR2 (N5714, N5712, N618);
buf BUF1 (N5715, N5705);
nand NAND4 (N5716, N5702, N2634, N174, N3007);
xor XOR2 (N5717, N5692, N2603);
nor NOR2 (N5718, N5709, N4444);
xor XOR2 (N5719, N5718, N5511);
nor NOR2 (N5720, N5715, N1071);
nand NAND3 (N5721, N5696, N2986, N207);
nand NAND4 (N5722, N5716, N3327, N533, N259);
buf BUF1 (N5723, N5713);
nor NOR2 (N5724, N5714, N2806);
nand NAND3 (N5725, N5717, N2779, N2242);
xor XOR2 (N5726, N5722, N2871);
buf BUF1 (N5727, N5724);
nand NAND4 (N5728, N5707, N792, N732, N2474);
not NOT1 (N5729, N5700);
nor NOR2 (N5730, N5720, N3634);
nand NAND4 (N5731, N5723, N2576, N3372, N5274);
or OR4 (N5732, N5706, N4607, N5246, N4972);
not NOT1 (N5733, N5731);
nor NOR4 (N5734, N5733, N2811, N2526, N3342);
or OR3 (N5735, N5727, N4145, N2754);
xor XOR2 (N5736, N5729, N869);
or OR3 (N5737, N5732, N4672, N514);
or OR2 (N5738, N5728, N2745);
nor NOR2 (N5739, N5730, N160);
nand NAND3 (N5740, N5721, N4440, N1945);
buf BUF1 (N5741, N5719);
buf BUF1 (N5742, N5741);
xor XOR2 (N5743, N5740, N4599);
xor XOR2 (N5744, N5743, N5660);
or OR2 (N5745, N5738, N2523);
nand NAND4 (N5746, N5736, N5528, N83, N3070);
buf BUF1 (N5747, N5739);
and AND4 (N5748, N5745, N5434, N1349, N4701);
nand NAND4 (N5749, N5734, N3693, N42, N4039);
and AND4 (N5750, N5742, N5077, N2337, N4654);
and AND2 (N5751, N5744, N2862);
xor XOR2 (N5752, N5725, N3947);
buf BUF1 (N5753, N5750);
and AND2 (N5754, N5737, N4235);
nand NAND2 (N5755, N5726, N362);
and AND2 (N5756, N5755, N5448);
and AND3 (N5757, N5752, N2552, N1676);
nor NOR3 (N5758, N5749, N3578, N2828);
nor NOR3 (N5759, N5758, N3048, N3853);
not NOT1 (N5760, N5751);
xor XOR2 (N5761, N5753, N401);
not NOT1 (N5762, N5757);
nand NAND3 (N5763, N5747, N1665, N2510);
buf BUF1 (N5764, N5763);
not NOT1 (N5765, N5735);
not NOT1 (N5766, N5754);
or OR3 (N5767, N5761, N1857, N4380);
and AND4 (N5768, N5762, N5327, N2101, N3224);
xor XOR2 (N5769, N5767, N4596);
and AND3 (N5770, N5764, N314, N5545);
nand NAND2 (N5771, N5768, N633);
and AND2 (N5772, N5748, N3712);
buf BUF1 (N5773, N5771);
not NOT1 (N5774, N5772);
nor NOR3 (N5775, N5774, N1958, N335);
not NOT1 (N5776, N5759);
nand NAND2 (N5777, N5756, N1580);
xor XOR2 (N5778, N5776, N3721);
xor XOR2 (N5779, N5775, N3826);
nor NOR4 (N5780, N5766, N1832, N3736, N2641);
not NOT1 (N5781, N5769);
or OR4 (N5782, N5781, N2564, N2552, N1708);
not NOT1 (N5783, N5770);
xor XOR2 (N5784, N5783, N3151);
xor XOR2 (N5785, N5760, N5090);
xor XOR2 (N5786, N5746, N562);
or OR3 (N5787, N5779, N1956, N4630);
nor NOR4 (N5788, N5773, N1443, N3902, N5650);
nand NAND4 (N5789, N5784, N16, N3391, N2851);
xor XOR2 (N5790, N5780, N5302);
nand NAND2 (N5791, N5778, N923);
and AND3 (N5792, N5782, N4885, N5754);
buf BUF1 (N5793, N5791);
nand NAND3 (N5794, N5788, N5264, N1402);
or OR3 (N5795, N5793, N5123, N49);
buf BUF1 (N5796, N5787);
nor NOR2 (N5797, N5777, N528);
nor NOR4 (N5798, N5795, N692, N1849, N3844);
nand NAND4 (N5799, N5765, N4175, N5782, N4501);
buf BUF1 (N5800, N5794);
buf BUF1 (N5801, N5798);
xor XOR2 (N5802, N5786, N1172);
and AND4 (N5803, N5790, N4251, N5212, N578);
nor NOR2 (N5804, N5802, N1411);
nor NOR3 (N5805, N5789, N4454, N2562);
xor XOR2 (N5806, N5801, N3172);
nand NAND4 (N5807, N5806, N4193, N1817, N195);
buf BUF1 (N5808, N5799);
buf BUF1 (N5809, N5808);
buf BUF1 (N5810, N5797);
or OR2 (N5811, N5809, N1062);
buf BUF1 (N5812, N5804);
or OR4 (N5813, N5805, N5562, N2617, N760);
xor XOR2 (N5814, N5812, N5523);
nand NAND4 (N5815, N5800, N1567, N4403, N5324);
and AND3 (N5816, N5813, N5660, N4693);
nor NOR3 (N5817, N5811, N4196, N2041);
not NOT1 (N5818, N5816);
or OR2 (N5819, N5803, N1237);
nand NAND3 (N5820, N5818, N3243, N5603);
nor NOR2 (N5821, N5815, N1192);
nand NAND2 (N5822, N5807, N3475);
nor NOR2 (N5823, N5785, N3550);
nor NOR2 (N5824, N5823, N4532);
and AND4 (N5825, N5817, N5232, N3858, N4746);
nand NAND4 (N5826, N5824, N1207, N3649, N1583);
nor NOR3 (N5827, N5792, N3360, N1682);
nand NAND2 (N5828, N5822, N4145);
or OR2 (N5829, N5814, N4546);
nand NAND3 (N5830, N5826, N4871, N4368);
nand NAND2 (N5831, N5810, N2712);
nand NAND4 (N5832, N5821, N2289, N5230, N1466);
not NOT1 (N5833, N5831);
and AND2 (N5834, N5825, N1271);
nor NOR3 (N5835, N5796, N3692, N4179);
nand NAND4 (N5836, N5820, N2053, N4601, N3356);
nor NOR4 (N5837, N5828, N4439, N5538, N4189);
xor XOR2 (N5838, N5832, N5540);
xor XOR2 (N5839, N5836, N1854);
or OR2 (N5840, N5835, N1026);
or OR3 (N5841, N5837, N2960, N2930);
nand NAND4 (N5842, N5827, N3707, N4900, N5735);
and AND2 (N5843, N5841, N4205);
or OR3 (N5844, N5838, N3540, N557);
nor NOR2 (N5845, N5844, N547);
or OR4 (N5846, N5842, N1121, N4687, N2590);
nand NAND3 (N5847, N5829, N4828, N5805);
buf BUF1 (N5848, N5845);
not NOT1 (N5849, N5843);
or OR3 (N5850, N5839, N4100, N1134);
nand NAND3 (N5851, N5847, N1864, N5211);
or OR3 (N5852, N5833, N373, N1842);
not NOT1 (N5853, N5846);
and AND2 (N5854, N5849, N3455);
xor XOR2 (N5855, N5851, N651);
nand NAND4 (N5856, N5834, N2781, N2464, N4472);
buf BUF1 (N5857, N5856);
nor NOR4 (N5858, N5855, N2075, N2379, N2920);
xor XOR2 (N5859, N5848, N2858);
nor NOR4 (N5860, N5853, N5107, N5529, N5403);
and AND4 (N5861, N5850, N1566, N875, N4420);
nor NOR2 (N5862, N5830, N3442);
xor XOR2 (N5863, N5840, N4507);
and AND2 (N5864, N5858, N4258);
nor NOR4 (N5865, N5819, N3764, N1965, N557);
not NOT1 (N5866, N5861);
xor XOR2 (N5867, N5866, N3337);
nand NAND3 (N5868, N5857, N2900, N4085);
not NOT1 (N5869, N5865);
and AND3 (N5870, N5862, N1367, N3165);
xor XOR2 (N5871, N5864, N1787);
nor NOR4 (N5872, N5869, N2420, N275, N1993);
and AND4 (N5873, N5868, N1024, N804, N4453);
and AND3 (N5874, N5870, N657, N2239);
not NOT1 (N5875, N5872);
and AND3 (N5876, N5860, N2537, N2011);
nand NAND3 (N5877, N5863, N826, N4883);
nand NAND2 (N5878, N5859, N5458);
or OR3 (N5879, N5877, N3685, N465);
xor XOR2 (N5880, N5852, N2615);
buf BUF1 (N5881, N5871);
or OR4 (N5882, N5873, N3096, N5248, N3673);
and AND3 (N5883, N5876, N5301, N4093);
nor NOR2 (N5884, N5854, N3916);
xor XOR2 (N5885, N5879, N3248);
buf BUF1 (N5886, N5882);
buf BUF1 (N5887, N5878);
buf BUF1 (N5888, N5880);
or OR4 (N5889, N5875, N3989, N4256, N3307);
xor XOR2 (N5890, N5889, N3993);
buf BUF1 (N5891, N5885);
and AND4 (N5892, N5881, N1196, N283, N3006);
and AND3 (N5893, N5874, N1512, N2726);
and AND4 (N5894, N5890, N4140, N356, N4102);
buf BUF1 (N5895, N5883);
not NOT1 (N5896, N5891);
buf BUF1 (N5897, N5892);
not NOT1 (N5898, N5897);
buf BUF1 (N5899, N5887);
or OR3 (N5900, N5893, N2567, N553);
xor XOR2 (N5901, N5867, N4702);
xor XOR2 (N5902, N5884, N2658);
buf BUF1 (N5903, N5899);
xor XOR2 (N5904, N5898, N4740);
nand NAND4 (N5905, N5888, N139, N2449, N5756);
nand NAND2 (N5906, N5886, N2376);
nand NAND3 (N5907, N5906, N2880, N1245);
or OR4 (N5908, N5905, N2620, N4785, N3059);
nor NOR4 (N5909, N5900, N3570, N473, N2759);
or OR2 (N5910, N5895, N4907);
xor XOR2 (N5911, N5908, N1504);
not NOT1 (N5912, N5902);
nand NAND4 (N5913, N5903, N5156, N246, N818);
nor NOR2 (N5914, N5910, N4333);
not NOT1 (N5915, N5907);
nor NOR3 (N5916, N5911, N2461, N4843);
buf BUF1 (N5917, N5913);
nand NAND2 (N5918, N5916, N4172);
and AND2 (N5919, N5901, N507);
or OR2 (N5920, N5894, N4926);
or OR3 (N5921, N5904, N1386, N935);
and AND4 (N5922, N5918, N3182, N3118, N5392);
xor XOR2 (N5923, N5914, N4730);
nor NOR2 (N5924, N5920, N4403);
and AND2 (N5925, N5922, N1341);
xor XOR2 (N5926, N5912, N692);
xor XOR2 (N5927, N5896, N1866);
nand NAND3 (N5928, N5926, N436, N968);
xor XOR2 (N5929, N5915, N293);
nor NOR2 (N5930, N5928, N937);
not NOT1 (N5931, N5923);
or OR3 (N5932, N5927, N4969, N2352);
or OR3 (N5933, N5931, N107, N4550);
not NOT1 (N5934, N5930);
nand NAND4 (N5935, N5924, N4498, N58, N461);
xor XOR2 (N5936, N5934, N872);
not NOT1 (N5937, N5933);
and AND2 (N5938, N5936, N5058);
not NOT1 (N5939, N5932);
nor NOR4 (N5940, N5909, N1999, N4416, N3717);
or OR2 (N5941, N5937, N1319);
xor XOR2 (N5942, N5919, N5224);
nand NAND3 (N5943, N5929, N454, N2341);
nor NOR2 (N5944, N5941, N4015);
and AND4 (N5945, N5944, N4733, N5050, N2766);
nand NAND3 (N5946, N5939, N1984, N80);
not NOT1 (N5947, N5945);
nand NAND4 (N5948, N5946, N3170, N5331, N2848);
not NOT1 (N5949, N5948);
xor XOR2 (N5950, N5925, N4095);
nand NAND3 (N5951, N5935, N1450, N833);
nor NOR2 (N5952, N5950, N2779);
nor NOR4 (N5953, N5951, N3373, N5644, N5633);
or OR4 (N5954, N5949, N1880, N4185, N5231);
buf BUF1 (N5955, N5952);
and AND4 (N5956, N5943, N4666, N607, N4472);
xor XOR2 (N5957, N5917, N2182);
buf BUF1 (N5958, N5921);
xor XOR2 (N5959, N5956, N756);
and AND2 (N5960, N5958, N2060);
or OR4 (N5961, N5954, N5253, N2693, N491);
xor XOR2 (N5962, N5957, N3778);
and AND2 (N5963, N5962, N5342);
and AND2 (N5964, N5938, N779);
xor XOR2 (N5965, N5960, N1332);
not NOT1 (N5966, N5964);
and AND3 (N5967, N5947, N3218, N5765);
buf BUF1 (N5968, N5965);
nor NOR2 (N5969, N5961, N1353);
or OR2 (N5970, N5968, N2757);
and AND3 (N5971, N5953, N5255, N3109);
buf BUF1 (N5972, N5966);
not NOT1 (N5973, N5942);
not NOT1 (N5974, N5970);
and AND3 (N5975, N5963, N1593, N4911);
buf BUF1 (N5976, N5959);
not NOT1 (N5977, N5975);
buf BUF1 (N5978, N5955);
not NOT1 (N5979, N5971);
not NOT1 (N5980, N5972);
not NOT1 (N5981, N5969);
nor NOR2 (N5982, N5977, N2037);
nand NAND3 (N5983, N5940, N3063, N3686);
nand NAND4 (N5984, N5980, N5127, N1433, N172);
buf BUF1 (N5985, N5981);
or OR4 (N5986, N5974, N1128, N2007, N4600);
not NOT1 (N5987, N5978);
or OR2 (N5988, N5986, N2265);
buf BUF1 (N5989, N5984);
and AND3 (N5990, N5983, N3523, N3265);
xor XOR2 (N5991, N5988, N1291);
and AND3 (N5992, N5990, N5019, N5723);
xor XOR2 (N5993, N5976, N5344);
not NOT1 (N5994, N5989);
not NOT1 (N5995, N5967);
and AND3 (N5996, N5994, N3332, N5956);
nand NAND4 (N5997, N5995, N4014, N3354, N5634);
or OR4 (N5998, N5973, N646, N3910, N3819);
nand NAND3 (N5999, N5998, N2730, N5293);
not NOT1 (N6000, N5982);
not NOT1 (N6001, N5985);
nor NOR2 (N6002, N5979, N5221);
nor NOR4 (N6003, N6001, N1674, N5820, N426);
xor XOR2 (N6004, N6000, N3179);
nand NAND2 (N6005, N5993, N1302);
xor XOR2 (N6006, N5997, N3691);
and AND3 (N6007, N5992, N1345, N4747);
xor XOR2 (N6008, N6002, N2218);
nor NOR3 (N6009, N5987, N2483, N3104);
buf BUF1 (N6010, N5999);
or OR2 (N6011, N6004, N1131);
nand NAND4 (N6012, N6006, N1752, N3901, N2927);
nand NAND2 (N6013, N6011, N3415);
not NOT1 (N6014, N6009);
nand NAND2 (N6015, N6013, N3396);
not NOT1 (N6016, N6003);
and AND3 (N6017, N5991, N3683, N3233);
not NOT1 (N6018, N6016);
and AND2 (N6019, N6010, N1002);
nor NOR2 (N6020, N6015, N2240);
and AND2 (N6021, N6018, N3147);
nand NAND4 (N6022, N6012, N4732, N4532, N1317);
or OR3 (N6023, N6005, N3838, N3185);
and AND3 (N6024, N5996, N5729, N3093);
buf BUF1 (N6025, N6007);
or OR2 (N6026, N6022, N968);
xor XOR2 (N6027, N6020, N2215);
nor NOR2 (N6028, N6019, N2445);
nor NOR2 (N6029, N6014, N874);
nor NOR3 (N6030, N6026, N4197, N4262);
nand NAND2 (N6031, N6025, N5310);
or OR3 (N6032, N6023, N2011, N5373);
xor XOR2 (N6033, N6031, N2800);
nand NAND2 (N6034, N6029, N1849);
not NOT1 (N6035, N6017);
xor XOR2 (N6036, N6033, N2899);
xor XOR2 (N6037, N6030, N2848);
not NOT1 (N6038, N6036);
or OR2 (N6039, N6028, N4078);
nor NOR3 (N6040, N6035, N4265, N4906);
or OR2 (N6041, N6032, N337);
nor NOR3 (N6042, N6008, N4313, N235);
or OR3 (N6043, N6038, N266, N5857);
xor XOR2 (N6044, N6037, N4739);
not NOT1 (N6045, N6040);
nand NAND3 (N6046, N6041, N4513, N3463);
xor XOR2 (N6047, N6046, N1254);
buf BUF1 (N6048, N6034);
xor XOR2 (N6049, N6027, N757);
nand NAND3 (N6050, N6043, N5469, N3424);
nor NOR2 (N6051, N6021, N3007);
xor XOR2 (N6052, N6047, N5754);
or OR3 (N6053, N6050, N5523, N4993);
not NOT1 (N6054, N6042);
nand NAND4 (N6055, N6052, N3844, N208, N4593);
and AND4 (N6056, N6045, N2563, N5508, N3555);
or OR4 (N6057, N6049, N4634, N745, N4199);
nand NAND2 (N6058, N6056, N5685);
or OR4 (N6059, N6048, N1339, N6008, N1337);
buf BUF1 (N6060, N6024);
or OR4 (N6061, N6058, N5356, N779, N3790);
nor NOR3 (N6062, N6039, N2107, N4232);
and AND2 (N6063, N6055, N495);
not NOT1 (N6064, N6059);
or OR3 (N6065, N6053, N2430, N3293);
nand NAND3 (N6066, N6060, N5821, N3345);
nor NOR4 (N6067, N6063, N5975, N4455, N4660);
nor NOR3 (N6068, N6061, N5729, N4508);
buf BUF1 (N6069, N6051);
nand NAND2 (N6070, N6057, N1866);
nand NAND3 (N6071, N6064, N4712, N2000);
nor NOR2 (N6072, N6068, N430);
xor XOR2 (N6073, N6062, N5055);
xor XOR2 (N6074, N6070, N3807);
nand NAND3 (N6075, N6073, N353, N2622);
and AND4 (N6076, N6075, N1356, N4881, N5732);
xor XOR2 (N6077, N6069, N4621);
not NOT1 (N6078, N6066);
and AND3 (N6079, N6067, N2912, N3448);
buf BUF1 (N6080, N6079);
xor XOR2 (N6081, N6074, N4871);
and AND3 (N6082, N6078, N4484, N5567);
or OR2 (N6083, N6082, N3692);
not NOT1 (N6084, N6044);
not NOT1 (N6085, N6084);
nand NAND2 (N6086, N6072, N24);
xor XOR2 (N6087, N6080, N4732);
xor XOR2 (N6088, N6076, N3568);
and AND4 (N6089, N6085, N5170, N5150, N1672);
or OR4 (N6090, N6071, N2877, N3126, N5903);
buf BUF1 (N6091, N6089);
nand NAND4 (N6092, N6081, N2968, N3550, N1453);
buf BUF1 (N6093, N6054);
and AND4 (N6094, N6065, N3408, N5498, N4200);
buf BUF1 (N6095, N6093);
nand NAND2 (N6096, N6087, N3405);
buf BUF1 (N6097, N6077);
not NOT1 (N6098, N6088);
or OR4 (N6099, N6091, N247, N1109, N2531);
or OR3 (N6100, N6094, N3848, N2165);
xor XOR2 (N6101, N6098, N3154);
nand NAND4 (N6102, N6100, N2455, N5522, N3927);
nor NOR2 (N6103, N6096, N2339);
and AND3 (N6104, N6099, N4010, N4289);
xor XOR2 (N6105, N6104, N2315);
nand NAND3 (N6106, N6090, N2095, N176);
not NOT1 (N6107, N6083);
and AND4 (N6108, N6103, N3171, N838, N3750);
nand NAND2 (N6109, N6107, N1306);
not NOT1 (N6110, N6095);
nor NOR2 (N6111, N6110, N883);
nand NAND2 (N6112, N6101, N5548);
nor NOR3 (N6113, N6102, N894, N5660);
nand NAND2 (N6114, N6086, N1199);
xor XOR2 (N6115, N6105, N3649);
buf BUF1 (N6116, N6106);
not NOT1 (N6117, N6092);
nand NAND2 (N6118, N6115, N1677);
nor NOR4 (N6119, N6118, N1614, N3482, N4124);
buf BUF1 (N6120, N6111);
not NOT1 (N6121, N6119);
nand NAND4 (N6122, N6120, N3787, N1669, N5319);
and AND2 (N6123, N6113, N2220);
xor XOR2 (N6124, N6117, N3077);
nor NOR2 (N6125, N6097, N4664);
and AND4 (N6126, N6109, N5290, N308, N5630);
buf BUF1 (N6127, N6125);
or OR2 (N6128, N6121, N4829);
not NOT1 (N6129, N6127);
nand NAND2 (N6130, N6124, N2443);
xor XOR2 (N6131, N6114, N3610);
or OR2 (N6132, N6122, N4074);
nand NAND4 (N6133, N6112, N5506, N560, N205);
buf BUF1 (N6134, N6129);
nor NOR2 (N6135, N6126, N1282);
nand NAND4 (N6136, N6131, N5257, N2738, N1570);
nand NAND2 (N6137, N6133, N6082);
buf BUF1 (N6138, N6128);
nand NAND4 (N6139, N6134, N3107, N1269, N324);
nand NAND3 (N6140, N6137, N5466, N3055);
and AND3 (N6141, N6140, N343, N3498);
nand NAND2 (N6142, N6132, N5391);
nor NOR4 (N6143, N6130, N2161, N4576, N2597);
xor XOR2 (N6144, N6138, N1355);
buf BUF1 (N6145, N6141);
not NOT1 (N6146, N6108);
nor NOR4 (N6147, N6139, N1728, N2359, N1794);
and AND2 (N6148, N6145, N2552);
not NOT1 (N6149, N6146);
and AND3 (N6150, N6135, N1238, N252);
not NOT1 (N6151, N6116);
not NOT1 (N6152, N6150);
nand NAND2 (N6153, N6147, N3150);
nand NAND4 (N6154, N6153, N5964, N4670, N1940);
xor XOR2 (N6155, N6143, N2308);
and AND2 (N6156, N6151, N1566);
nor NOR2 (N6157, N6142, N4334);
not NOT1 (N6158, N6144);
buf BUF1 (N6159, N6148);
and AND4 (N6160, N6136, N984, N1249, N1441);
buf BUF1 (N6161, N6155);
buf BUF1 (N6162, N6160);
xor XOR2 (N6163, N6158, N3061);
xor XOR2 (N6164, N6163, N1314);
and AND3 (N6165, N6164, N286, N5234);
buf BUF1 (N6166, N6162);
and AND2 (N6167, N6165, N791);
buf BUF1 (N6168, N6157);
not NOT1 (N6169, N6167);
xor XOR2 (N6170, N6154, N3329);
nand NAND3 (N6171, N6169, N142, N4480);
nor NOR3 (N6172, N6156, N1604, N926);
xor XOR2 (N6173, N6172, N2797);
not NOT1 (N6174, N6161);
xor XOR2 (N6175, N6171, N5951);
and AND4 (N6176, N6175, N2199, N3102, N3763);
buf BUF1 (N6177, N6173);
or OR3 (N6178, N6123, N1156, N5688);
nand NAND2 (N6179, N6166, N317);
buf BUF1 (N6180, N6152);
nor NOR4 (N6181, N6174, N3228, N4582, N1574);
or OR4 (N6182, N6179, N2974, N349, N4710);
buf BUF1 (N6183, N6159);
and AND4 (N6184, N6176, N5522, N660, N6107);
nor NOR2 (N6185, N6180, N2924);
nor NOR2 (N6186, N6185, N2861);
xor XOR2 (N6187, N6183, N3906);
xor XOR2 (N6188, N6182, N3470);
buf BUF1 (N6189, N6187);
buf BUF1 (N6190, N6178);
nand NAND4 (N6191, N6177, N2711, N3404, N3658);
or OR2 (N6192, N6186, N4131);
nand NAND2 (N6193, N6170, N2346);
not NOT1 (N6194, N6149);
buf BUF1 (N6195, N6188);
and AND3 (N6196, N6181, N3817, N1458);
or OR4 (N6197, N6184, N5278, N3973, N4780);
not NOT1 (N6198, N6197);
nor NOR2 (N6199, N6196, N1920);
nand NAND3 (N6200, N6191, N2244, N5325);
not NOT1 (N6201, N6192);
and AND3 (N6202, N6189, N3843, N6044);
nor NOR4 (N6203, N6200, N1430, N6086, N3034);
or OR2 (N6204, N6202, N6089);
nor NOR2 (N6205, N6201, N622);
xor XOR2 (N6206, N6198, N4399);
nand NAND3 (N6207, N6193, N1425, N386);
and AND2 (N6208, N6204, N105);
buf BUF1 (N6209, N6206);
buf BUF1 (N6210, N6205);
not NOT1 (N6211, N6208);
nor NOR4 (N6212, N6194, N3932, N5886, N858);
nand NAND2 (N6213, N6207, N215);
nand NAND3 (N6214, N6213, N1529, N4974);
or OR3 (N6215, N6212, N4308, N551);
nand NAND4 (N6216, N6168, N4728, N2145, N6198);
nand NAND4 (N6217, N6214, N3649, N1266, N2995);
not NOT1 (N6218, N6217);
buf BUF1 (N6219, N6190);
nor NOR2 (N6220, N6219, N242);
nand NAND3 (N6221, N6195, N607, N2290);
nor NOR4 (N6222, N6220, N314, N2405, N114);
not NOT1 (N6223, N6222);
and AND3 (N6224, N6215, N5009, N3501);
nand NAND3 (N6225, N6211, N5100, N3451);
nand NAND2 (N6226, N6225, N4004);
and AND3 (N6227, N6224, N3544, N4838);
or OR3 (N6228, N6218, N913, N1755);
not NOT1 (N6229, N6223);
or OR3 (N6230, N6227, N3565, N5009);
nor NOR3 (N6231, N6216, N2875, N244);
nor NOR4 (N6232, N6226, N5817, N266, N3745);
nand NAND3 (N6233, N6210, N1590, N5646);
nand NAND2 (N6234, N6229, N3082);
and AND2 (N6235, N6209, N5963);
nand NAND3 (N6236, N6232, N2757, N4444);
xor XOR2 (N6237, N6235, N4266);
nor NOR4 (N6238, N6233, N5049, N5383, N4614);
nor NOR3 (N6239, N6234, N2214, N2225);
nor NOR2 (N6240, N6221, N3296);
not NOT1 (N6241, N6231);
xor XOR2 (N6242, N6239, N3760);
buf BUF1 (N6243, N6241);
xor XOR2 (N6244, N6243, N4147);
xor XOR2 (N6245, N6236, N2877);
or OR4 (N6246, N6242, N3894, N2019, N2044);
nor NOR2 (N6247, N6244, N440);
not NOT1 (N6248, N6240);
nor NOR4 (N6249, N6246, N4596, N1591, N2794);
buf BUF1 (N6250, N6248);
nor NOR3 (N6251, N6250, N3814, N137);
not NOT1 (N6252, N6199);
buf BUF1 (N6253, N6247);
not NOT1 (N6254, N6252);
nand NAND3 (N6255, N6253, N4539, N416);
nand NAND3 (N6256, N6245, N6102, N498);
or OR4 (N6257, N6255, N836, N2315, N196);
or OR2 (N6258, N6203, N2431);
buf BUF1 (N6259, N6257);
not NOT1 (N6260, N6230);
xor XOR2 (N6261, N6258, N4742);
or OR2 (N6262, N6249, N188);
not NOT1 (N6263, N6261);
and AND3 (N6264, N6259, N5996, N3286);
not NOT1 (N6265, N6263);
nand NAND2 (N6266, N6260, N392);
xor XOR2 (N6267, N6237, N3740);
buf BUF1 (N6268, N6238);
or OR4 (N6269, N6265, N5940, N5993, N5631);
nor NOR2 (N6270, N6228, N1726);
or OR3 (N6271, N6264, N5294, N5530);
not NOT1 (N6272, N6262);
nor NOR2 (N6273, N6269, N2078);
nand NAND2 (N6274, N6256, N2739);
or OR4 (N6275, N6270, N3728, N6252, N5584);
nor NOR3 (N6276, N6266, N4231, N5328);
buf BUF1 (N6277, N6276);
nand NAND3 (N6278, N6272, N3738, N256);
and AND4 (N6279, N6268, N690, N5833, N1490);
nand NAND4 (N6280, N6251, N2832, N3663, N1276);
and AND2 (N6281, N6254, N3772);
xor XOR2 (N6282, N6278, N3151);
and AND2 (N6283, N6279, N842);
xor XOR2 (N6284, N6275, N556);
or OR3 (N6285, N6277, N44, N2961);
nand NAND2 (N6286, N6273, N2373);
nor NOR3 (N6287, N6274, N4538, N1686);
buf BUF1 (N6288, N6284);
not NOT1 (N6289, N6287);
or OR2 (N6290, N6267, N2413);
nor NOR3 (N6291, N6282, N3791, N4009);
nor NOR3 (N6292, N6289, N462, N6119);
xor XOR2 (N6293, N6290, N702);
not NOT1 (N6294, N6286);
nor NOR3 (N6295, N6292, N4302, N5416);
buf BUF1 (N6296, N6281);
nand NAND3 (N6297, N6293, N4500, N654);
nand NAND4 (N6298, N6297, N5434, N4725, N1711);
xor XOR2 (N6299, N6271, N1154);
nand NAND2 (N6300, N6288, N4729);
and AND4 (N6301, N6283, N1004, N3964, N1781);
and AND4 (N6302, N6294, N2972, N4017, N1940);
nand NAND2 (N6303, N6300, N1989);
and AND4 (N6304, N6298, N4745, N5984, N5830);
and AND3 (N6305, N6285, N2679, N1470);
or OR4 (N6306, N6304, N2406, N6043, N1643);
nand NAND2 (N6307, N6305, N2573);
and AND3 (N6308, N6301, N3065, N4511);
nor NOR4 (N6309, N6307, N2707, N2465, N1672);
xor XOR2 (N6310, N6302, N135);
nor NOR3 (N6311, N6295, N2453, N423);
nor NOR4 (N6312, N6291, N5355, N60, N5247);
and AND3 (N6313, N6309, N4025, N1744);
and AND2 (N6314, N6306, N5776);
nor NOR3 (N6315, N6312, N4910, N5483);
nor NOR4 (N6316, N6296, N2382, N3040, N1787);
buf BUF1 (N6317, N6316);
or OR3 (N6318, N6303, N209, N4770);
not NOT1 (N6319, N6317);
xor XOR2 (N6320, N6315, N4410);
and AND4 (N6321, N6308, N5164, N3482, N1750);
or OR4 (N6322, N6320, N4991, N462, N3928);
not NOT1 (N6323, N6319);
or OR2 (N6324, N6318, N3255);
or OR3 (N6325, N6314, N2756, N2901);
xor XOR2 (N6326, N6324, N3868);
buf BUF1 (N6327, N6280);
or OR4 (N6328, N6313, N6145, N5465, N3846);
nor NOR4 (N6329, N6321, N4536, N1803, N597);
and AND4 (N6330, N6327, N851, N3441, N5868);
not NOT1 (N6331, N6322);
nand NAND2 (N6332, N6311, N1472);
buf BUF1 (N6333, N6326);
or OR4 (N6334, N6332, N3076, N4440, N514);
xor XOR2 (N6335, N6325, N2551);
xor XOR2 (N6336, N6335, N1225);
buf BUF1 (N6337, N6323);
nand NAND3 (N6338, N6310, N4892, N41);
and AND3 (N6339, N6330, N3926, N3481);
not NOT1 (N6340, N6339);
xor XOR2 (N6341, N6331, N6123);
nand NAND4 (N6342, N6328, N1714, N4029, N3883);
not NOT1 (N6343, N6341);
xor XOR2 (N6344, N6333, N1666);
xor XOR2 (N6345, N6340, N3155);
and AND2 (N6346, N6345, N4513);
nand NAND4 (N6347, N6343, N1946, N4264, N150);
or OR3 (N6348, N6344, N913, N1314);
and AND4 (N6349, N6336, N2135, N1077, N812);
or OR4 (N6350, N6329, N4096, N109, N2997);
xor XOR2 (N6351, N6334, N6105);
not NOT1 (N6352, N6351);
buf BUF1 (N6353, N6337);
buf BUF1 (N6354, N6338);
and AND4 (N6355, N6350, N697, N6273, N3101);
not NOT1 (N6356, N6346);
nor NOR2 (N6357, N6348, N6097);
buf BUF1 (N6358, N6355);
not NOT1 (N6359, N6299);
nor NOR3 (N6360, N6358, N1669, N3285);
nor NOR3 (N6361, N6359, N4743, N4878);
xor XOR2 (N6362, N6342, N2590);
nand NAND3 (N6363, N6362, N4890, N1606);
or OR2 (N6364, N6360, N163);
buf BUF1 (N6365, N6349);
nand NAND4 (N6366, N6347, N4914, N4460, N5811);
nor NOR4 (N6367, N6353, N4042, N5182, N2060);
xor XOR2 (N6368, N6366, N525);
and AND3 (N6369, N6361, N4933, N3326);
and AND4 (N6370, N6368, N6264, N6238, N1571);
nor NOR3 (N6371, N6370, N2938, N5588);
nand NAND2 (N6372, N6369, N2153);
not NOT1 (N6373, N6352);
not NOT1 (N6374, N6372);
xor XOR2 (N6375, N6371, N5841);
xor XOR2 (N6376, N6356, N6114);
and AND3 (N6377, N6357, N464, N3857);
not NOT1 (N6378, N6364);
xor XOR2 (N6379, N6375, N288);
not NOT1 (N6380, N6378);
and AND4 (N6381, N6377, N3998, N3190, N3103);
buf BUF1 (N6382, N6376);
and AND2 (N6383, N6354, N1536);
buf BUF1 (N6384, N6373);
xor XOR2 (N6385, N6379, N3285);
not NOT1 (N6386, N6380);
or OR3 (N6387, N6384, N1568, N2619);
not NOT1 (N6388, N6374);
nor NOR4 (N6389, N6367, N2400, N5578, N1531);
nor NOR4 (N6390, N6365, N1614, N1929, N1210);
buf BUF1 (N6391, N6363);
nor NOR2 (N6392, N6387, N2644);
xor XOR2 (N6393, N6391, N1330);
nand NAND3 (N6394, N6388, N2800, N2894);
not NOT1 (N6395, N6382);
not NOT1 (N6396, N6390);
xor XOR2 (N6397, N6396, N4416);
nand NAND2 (N6398, N6395, N5706);
and AND3 (N6399, N6386, N5697, N3938);
and AND3 (N6400, N6399, N4722, N99);
nand NAND4 (N6401, N6398, N4972, N4682, N3261);
buf BUF1 (N6402, N6393);
and AND3 (N6403, N6397, N6343, N4040);
buf BUF1 (N6404, N6401);
xor XOR2 (N6405, N6402, N4598);
xor XOR2 (N6406, N6383, N2677);
or OR3 (N6407, N6385, N4000, N3820);
or OR2 (N6408, N6404, N5171);
not NOT1 (N6409, N6406);
and AND2 (N6410, N6381, N2986);
nand NAND2 (N6411, N6407, N1977);
and AND2 (N6412, N6408, N3604);
nand NAND3 (N6413, N6389, N1256, N114);
nand NAND2 (N6414, N6394, N85);
nor NOR2 (N6415, N6400, N5127);
xor XOR2 (N6416, N6392, N2327);
nand NAND4 (N6417, N6409, N5418, N2879, N526);
buf BUF1 (N6418, N6417);
buf BUF1 (N6419, N6405);
endmodule