// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12;

output N707,N689,N706,N710,N705,N690,N708,N691,N711,N712;

or OR3 (N13, N10, N10, N3);
nor NOR2 (N14, N10, N3);
or OR3 (N15, N4, N8, N8);
and AND4 (N16, N8, N9, N12, N13);
or OR4 (N17, N4, N2, N15, N13);
nand NAND3 (N18, N2, N11, N5);
xor XOR2 (N19, N2, N18);
nand NAND4 (N20, N19, N15, N4, N12);
nor NOR2 (N21, N4, N20);
or OR4 (N22, N3, N13, N20, N4);
not NOT1 (N23, N12);
not NOT1 (N24, N16);
not NOT1 (N25, N9);
nand NAND3 (N26, N11, N6, N15);
or OR2 (N27, N4, N3);
and AND3 (N28, N19, N24, N13);
and AND3 (N29, N28, N5, N25);
nor NOR3 (N30, N23, N23, N11);
buf BUF1 (N31, N20);
and AND2 (N32, N14, N6);
or OR2 (N33, N12, N22);
nand NAND3 (N34, N7, N30, N16);
and AND4 (N35, N22, N10, N6, N34);
and AND3 (N36, N11, N13, N14);
nor NOR2 (N37, N27, N29);
and AND2 (N38, N28, N29);
nand NAND4 (N39, N36, N19, N24, N18);
xor XOR2 (N40, N33, N11);
or OR2 (N41, N38, N10);
nand NAND3 (N42, N37, N21, N10);
nor NOR3 (N43, N1, N3, N19);
xor XOR2 (N44, N41, N27);
xor XOR2 (N45, N39, N8);
nor NOR4 (N46, N17, N7, N11, N30);
xor XOR2 (N47, N31, N14);
and AND4 (N48, N44, N39, N19, N2);
xor XOR2 (N49, N46, N20);
nor NOR4 (N50, N47, N46, N24, N39);
or OR3 (N51, N42, N8, N16);
and AND2 (N52, N49, N24);
nand NAND4 (N53, N26, N21, N36, N3);
and AND2 (N54, N50, N7);
buf BUF1 (N55, N54);
and AND2 (N56, N52, N33);
buf BUF1 (N57, N32);
and AND4 (N58, N43, N9, N11, N50);
nor NOR3 (N59, N51, N18, N8);
and AND2 (N60, N40, N18);
or OR4 (N61, N45, N39, N1, N37);
or OR2 (N62, N57, N10);
xor XOR2 (N63, N62, N48);
and AND4 (N64, N11, N39, N27, N26);
or OR2 (N65, N35, N18);
and AND3 (N66, N64, N10, N44);
and AND2 (N67, N58, N39);
nand NAND4 (N68, N65, N27, N14, N20);
nor NOR4 (N69, N59, N42, N20, N41);
and AND2 (N70, N53, N49);
nor NOR2 (N71, N63, N64);
and AND4 (N72, N71, N6, N64, N36);
nand NAND2 (N73, N72, N19);
nor NOR2 (N74, N69, N57);
nand NAND4 (N75, N68, N72, N22, N74);
or OR4 (N76, N22, N71, N13, N35);
xor XOR2 (N77, N60, N22);
and AND2 (N78, N66, N56);
or OR3 (N79, N29, N28, N66);
and AND3 (N80, N55, N66, N21);
nand NAND3 (N81, N67, N73, N78);
xor XOR2 (N82, N81, N9);
nand NAND2 (N83, N43, N44);
or OR2 (N84, N3, N25);
nand NAND3 (N85, N61, N11, N83);
xor XOR2 (N86, N45, N34);
xor XOR2 (N87, N84, N33);
and AND4 (N88, N86, N77, N34, N34);
and AND4 (N89, N26, N11, N46, N58);
and AND4 (N90, N89, N34, N84, N31);
and AND2 (N91, N70, N66);
xor XOR2 (N92, N88, N76);
nor NOR2 (N93, N6, N7);
and AND4 (N94, N87, N26, N87, N4);
nand NAND4 (N95, N91, N37, N66, N82);
and AND4 (N96, N36, N25, N15, N42);
nand NAND2 (N97, N95, N16);
and AND2 (N98, N90, N49);
xor XOR2 (N99, N75, N1);
buf BUF1 (N100, N94);
and AND3 (N101, N79, N85, N53);
xor XOR2 (N102, N36, N83);
buf BUF1 (N103, N102);
or OR4 (N104, N80, N35, N46, N79);
buf BUF1 (N105, N97);
or OR3 (N106, N99, N34, N1);
not NOT1 (N107, N93);
xor XOR2 (N108, N105, N11);
not NOT1 (N109, N106);
buf BUF1 (N110, N108);
buf BUF1 (N111, N101);
buf BUF1 (N112, N98);
and AND4 (N113, N103, N52, N26, N55);
not NOT1 (N114, N112);
buf BUF1 (N115, N107);
nand NAND4 (N116, N104, N101, N103, N63);
xor XOR2 (N117, N92, N39);
xor XOR2 (N118, N114, N79);
nor NOR3 (N119, N115, N36, N81);
buf BUF1 (N120, N110);
or OR3 (N121, N117, N96, N15);
buf BUF1 (N122, N20);
nand NAND3 (N123, N116, N14, N26);
buf BUF1 (N124, N118);
and AND4 (N125, N121, N117, N113, N120);
nand NAND2 (N126, N120, N14);
buf BUF1 (N127, N83);
nand NAND2 (N128, N122, N113);
nand NAND4 (N129, N125, N85, N60, N76);
buf BUF1 (N130, N128);
buf BUF1 (N131, N119);
buf BUF1 (N132, N131);
or OR2 (N133, N132, N93);
buf BUF1 (N134, N123);
nand NAND4 (N135, N124, N13, N99, N119);
and AND3 (N136, N133, N116, N59);
and AND3 (N137, N130, N2, N39);
nor NOR3 (N138, N100, N122, N97);
and AND2 (N139, N126, N124);
not NOT1 (N140, N109);
nor NOR4 (N141, N127, N55, N46, N133);
and AND2 (N142, N137, N45);
or OR2 (N143, N138, N139);
not NOT1 (N144, N105);
buf BUF1 (N145, N136);
nand NAND4 (N146, N134, N137, N27, N120);
nor NOR2 (N147, N135, N141);
xor XOR2 (N148, N12, N57);
nand NAND4 (N149, N147, N109, N64, N39);
xor XOR2 (N150, N148, N132);
xor XOR2 (N151, N144, N150);
or OR4 (N152, N62, N125, N30, N107);
buf BUF1 (N153, N143);
not NOT1 (N154, N149);
buf BUF1 (N155, N145);
not NOT1 (N156, N152);
nand NAND2 (N157, N140, N136);
not NOT1 (N158, N142);
xor XOR2 (N159, N157, N71);
or OR2 (N160, N155, N89);
and AND2 (N161, N111, N8);
buf BUF1 (N162, N151);
not NOT1 (N163, N160);
or OR4 (N164, N159, N62, N148, N85);
or OR3 (N165, N161, N5, N83);
xor XOR2 (N166, N154, N119);
or OR3 (N167, N153, N31, N65);
buf BUF1 (N168, N164);
not NOT1 (N169, N162);
buf BUF1 (N170, N168);
nor NOR2 (N171, N165, N20);
nor NOR4 (N172, N158, N51, N85, N60);
not NOT1 (N173, N163);
and AND3 (N174, N173, N62, N36);
nor NOR4 (N175, N129, N141, N117, N108);
nor NOR2 (N176, N156, N2);
nor NOR2 (N177, N167, N64);
or OR4 (N178, N171, N110, N159, N47);
xor XOR2 (N179, N178, N49);
xor XOR2 (N180, N170, N170);
or OR2 (N181, N172, N136);
nand NAND3 (N182, N181, N30, N176);
or OR2 (N183, N113, N66);
or OR4 (N184, N179, N47, N168, N7);
not NOT1 (N185, N174);
nand NAND2 (N186, N183, N148);
buf BUF1 (N187, N185);
buf BUF1 (N188, N182);
or OR3 (N189, N186, N27, N61);
not NOT1 (N190, N146);
xor XOR2 (N191, N175, N114);
not NOT1 (N192, N169);
and AND2 (N193, N189, N121);
and AND4 (N194, N188, N154, N161, N157);
buf BUF1 (N195, N193);
xor XOR2 (N196, N177, N43);
and AND4 (N197, N196, N44, N4, N170);
and AND3 (N198, N197, N66, N89);
or OR3 (N199, N190, N143, N35);
and AND3 (N200, N195, N72, N182);
or OR2 (N201, N184, N167);
or OR2 (N202, N201, N27);
or OR4 (N203, N166, N177, N83, N67);
nor NOR2 (N204, N202, N72);
buf BUF1 (N205, N199);
buf BUF1 (N206, N204);
not NOT1 (N207, N194);
nand NAND4 (N208, N198, N166, N106, N73);
not NOT1 (N209, N205);
xor XOR2 (N210, N187, N12);
nand NAND4 (N211, N206, N16, N54, N60);
nand NAND3 (N212, N192, N4, N210);
buf BUF1 (N213, N182);
not NOT1 (N214, N212);
and AND2 (N215, N214, N8);
nor NOR2 (N216, N200, N148);
nor NOR2 (N217, N208, N30);
xor XOR2 (N218, N213, N31);
buf BUF1 (N219, N209);
not NOT1 (N220, N207);
or OR4 (N221, N180, N168, N156, N74);
nor NOR2 (N222, N203, N200);
xor XOR2 (N223, N215, N188);
not NOT1 (N224, N220);
or OR3 (N225, N223, N86, N214);
not NOT1 (N226, N224);
or OR3 (N227, N219, N169, N146);
xor XOR2 (N228, N191, N161);
nand NAND3 (N229, N211, N35, N4);
or OR2 (N230, N222, N200);
or OR4 (N231, N225, N143, N11, N156);
buf BUF1 (N232, N228);
xor XOR2 (N233, N232, N142);
not NOT1 (N234, N229);
xor XOR2 (N235, N231, N173);
and AND4 (N236, N218, N13, N201, N200);
not NOT1 (N237, N236);
buf BUF1 (N238, N216);
xor XOR2 (N239, N221, N164);
nand NAND2 (N240, N234, N202);
nand NAND3 (N241, N233, N108, N178);
nand NAND3 (N242, N238, N93, N163);
or OR2 (N243, N239, N165);
nand NAND2 (N244, N230, N148);
nor NOR4 (N245, N226, N116, N79, N217);
buf BUF1 (N246, N133);
nand NAND3 (N247, N246, N87, N10);
buf BUF1 (N248, N244);
nand NAND3 (N249, N235, N177, N81);
buf BUF1 (N250, N227);
not NOT1 (N251, N245);
nand NAND3 (N252, N248, N107, N129);
or OR4 (N253, N242, N88, N181, N148);
nor NOR2 (N254, N241, N231);
xor XOR2 (N255, N237, N162);
xor XOR2 (N256, N254, N189);
not NOT1 (N257, N249);
buf BUF1 (N258, N251);
not NOT1 (N259, N252);
not NOT1 (N260, N243);
nor NOR2 (N261, N250, N177);
xor XOR2 (N262, N258, N90);
buf BUF1 (N263, N240);
buf BUF1 (N264, N261);
nor NOR2 (N265, N257, N156);
nand NAND2 (N266, N260, N116);
nor NOR3 (N267, N253, N187, N188);
nor NOR2 (N268, N255, N146);
and AND4 (N269, N262, N233, N162, N262);
or OR2 (N270, N266, N228);
buf BUF1 (N271, N256);
or OR2 (N272, N267, N60);
buf BUF1 (N273, N265);
and AND4 (N274, N269, N70, N31, N100);
and AND4 (N275, N274, N35, N245, N140);
or OR4 (N276, N247, N60, N254, N170);
not NOT1 (N277, N270);
nor NOR3 (N278, N277, N227, N114);
not NOT1 (N279, N259);
or OR4 (N280, N275, N221, N124, N151);
and AND4 (N281, N271, N243, N147, N46);
nand NAND2 (N282, N268, N238);
and AND3 (N283, N279, N270, N176);
nand NAND2 (N284, N281, N27);
and AND3 (N285, N280, N173, N255);
nand NAND4 (N286, N272, N38, N37, N5);
buf BUF1 (N287, N284);
and AND2 (N288, N276, N241);
nand NAND2 (N289, N283, N178);
xor XOR2 (N290, N288, N289);
nand NAND4 (N291, N280, N277, N47, N284);
or OR3 (N292, N263, N233, N213);
buf BUF1 (N293, N282);
not NOT1 (N294, N273);
nor NOR3 (N295, N293, N44, N126);
and AND4 (N296, N264, N191, N8, N205);
buf BUF1 (N297, N295);
buf BUF1 (N298, N294);
nand NAND4 (N299, N278, N230, N82, N234);
and AND2 (N300, N286, N157);
nor NOR3 (N301, N291, N143, N207);
or OR2 (N302, N287, N287);
nor NOR3 (N303, N301, N124, N55);
or OR2 (N304, N303, N13);
buf BUF1 (N305, N298);
xor XOR2 (N306, N285, N236);
nor NOR3 (N307, N302, N252, N83);
and AND3 (N308, N290, N128, N55);
buf BUF1 (N309, N292);
buf BUF1 (N310, N305);
xor XOR2 (N311, N308, N56);
nand NAND3 (N312, N307, N310, N144);
buf BUF1 (N313, N207);
buf BUF1 (N314, N313);
not NOT1 (N315, N300);
and AND4 (N316, N306, N180, N275, N12);
nor NOR3 (N317, N304, N64, N311);
nand NAND3 (N318, N47, N278, N11);
or OR3 (N319, N314, N267, N204);
buf BUF1 (N320, N315);
and AND4 (N321, N318, N317, N116, N210);
not NOT1 (N322, N242);
nor NOR3 (N323, N322, N257, N133);
buf BUF1 (N324, N319);
xor XOR2 (N325, N297, N114);
xor XOR2 (N326, N323, N7);
nor NOR4 (N327, N299, N134, N287, N133);
and AND2 (N328, N320, N325);
buf BUF1 (N329, N302);
not NOT1 (N330, N312);
or OR2 (N331, N316, N228);
nand NAND2 (N332, N328, N51);
nand NAND3 (N333, N330, N152, N148);
xor XOR2 (N334, N333, N61);
not NOT1 (N335, N309);
buf BUF1 (N336, N335);
and AND4 (N337, N334, N332, N209, N100);
xor XOR2 (N338, N133, N92);
and AND4 (N339, N336, N134, N181, N309);
or OR2 (N340, N324, N267);
or OR2 (N341, N321, N88);
and AND2 (N342, N340, N339);
not NOT1 (N343, N241);
buf BUF1 (N344, N343);
buf BUF1 (N345, N344);
nand NAND3 (N346, N341, N294, N91);
nor NOR2 (N347, N338, N159);
buf BUF1 (N348, N345);
xor XOR2 (N349, N326, N208);
not NOT1 (N350, N337);
buf BUF1 (N351, N329);
xor XOR2 (N352, N350, N258);
nor NOR4 (N353, N349, N214, N149, N90);
nor NOR4 (N354, N346, N154, N308, N164);
buf BUF1 (N355, N354);
buf BUF1 (N356, N296);
and AND4 (N357, N327, N237, N332, N333);
buf BUF1 (N358, N342);
not NOT1 (N359, N358);
and AND2 (N360, N356, N299);
not NOT1 (N361, N331);
xor XOR2 (N362, N357, N289);
or OR3 (N363, N360, N192, N212);
not NOT1 (N364, N361);
nor NOR2 (N365, N364, N65);
or OR2 (N366, N355, N62);
and AND2 (N367, N366, N19);
or OR3 (N368, N365, N67, N286);
not NOT1 (N369, N348);
or OR4 (N370, N353, N98, N53, N155);
not NOT1 (N371, N351);
or OR2 (N372, N371, N278);
or OR3 (N373, N363, N131, N107);
not NOT1 (N374, N347);
and AND4 (N375, N372, N321, N181, N194);
not NOT1 (N376, N373);
nor NOR3 (N377, N359, N108, N208);
not NOT1 (N378, N352);
not NOT1 (N379, N375);
or OR3 (N380, N378, N294, N201);
nand NAND2 (N381, N377, N234);
not NOT1 (N382, N367);
or OR2 (N383, N362, N204);
nand NAND4 (N384, N383, N209, N306, N169);
buf BUF1 (N385, N384);
nand NAND2 (N386, N376, N178);
or OR3 (N387, N386, N154, N124);
not NOT1 (N388, N374);
nand NAND2 (N389, N381, N93);
not NOT1 (N390, N389);
nor NOR3 (N391, N388, N70, N359);
not NOT1 (N392, N391);
or OR3 (N393, N379, N276, N54);
and AND3 (N394, N368, N6, N255);
and AND4 (N395, N385, N61, N153, N123);
nor NOR3 (N396, N382, N370, N219);
nor NOR3 (N397, N11, N150, N87);
xor XOR2 (N398, N394, N343);
or OR3 (N399, N393, N374, N330);
buf BUF1 (N400, N380);
xor XOR2 (N401, N392, N205);
not NOT1 (N402, N390);
or OR2 (N403, N387, N54);
xor XOR2 (N404, N399, N54);
and AND4 (N405, N401, N82, N269, N101);
and AND4 (N406, N398, N233, N174, N62);
and AND3 (N407, N404, N122, N387);
nand NAND2 (N408, N395, N356);
buf BUF1 (N409, N406);
not NOT1 (N410, N409);
buf BUF1 (N411, N402);
nor NOR3 (N412, N405, N41, N56);
and AND2 (N413, N403, N160);
buf BUF1 (N414, N396);
xor XOR2 (N415, N412, N373);
and AND4 (N416, N414, N28, N287, N345);
nand NAND2 (N417, N415, N183);
xor XOR2 (N418, N408, N268);
or OR3 (N419, N418, N383, N291);
or OR3 (N420, N397, N291, N337);
or OR4 (N421, N400, N147, N231, N255);
buf BUF1 (N422, N413);
buf BUF1 (N423, N411);
and AND3 (N424, N419, N112, N125);
and AND4 (N425, N410, N46, N85, N53);
and AND4 (N426, N417, N258, N182, N120);
or OR2 (N427, N420, N271);
and AND2 (N428, N427, N310);
nand NAND2 (N429, N407, N6);
nor NOR4 (N430, N424, N137, N365, N290);
or OR4 (N431, N429, N206, N106, N297);
buf BUF1 (N432, N425);
and AND3 (N433, N422, N236, N199);
xor XOR2 (N434, N416, N17);
xor XOR2 (N435, N426, N19);
not NOT1 (N436, N428);
nor NOR4 (N437, N432, N419, N206, N259);
xor XOR2 (N438, N433, N194);
xor XOR2 (N439, N436, N87);
and AND3 (N440, N421, N214, N255);
not NOT1 (N441, N439);
xor XOR2 (N442, N437, N293);
not NOT1 (N443, N441);
not NOT1 (N444, N435);
and AND2 (N445, N434, N190);
nand NAND2 (N446, N430, N179);
xor XOR2 (N447, N431, N302);
or OR4 (N448, N446, N188, N72, N195);
xor XOR2 (N449, N448, N440);
nand NAND2 (N450, N178, N70);
nor NOR3 (N451, N423, N328, N154);
nor NOR2 (N452, N438, N334);
and AND2 (N453, N450, N440);
and AND2 (N454, N452, N214);
nor NOR3 (N455, N447, N191, N317);
not NOT1 (N456, N455);
or OR4 (N457, N445, N308, N429, N369);
xor XOR2 (N458, N333, N262);
not NOT1 (N459, N458);
nand NAND4 (N460, N454, N404, N420, N418);
or OR3 (N461, N460, N432, N140);
or OR3 (N462, N449, N218, N173);
buf BUF1 (N463, N451);
or OR2 (N464, N463, N371);
and AND3 (N465, N461, N327, N54);
nand NAND2 (N466, N443, N236);
buf BUF1 (N467, N465);
buf BUF1 (N468, N466);
or OR4 (N469, N468, N129, N430, N350);
buf BUF1 (N470, N456);
not NOT1 (N471, N459);
or OR3 (N472, N467, N45, N325);
not NOT1 (N473, N470);
or OR2 (N474, N442, N264);
or OR2 (N475, N469, N89);
or OR3 (N476, N471, N34, N333);
buf BUF1 (N477, N472);
buf BUF1 (N478, N462);
xor XOR2 (N479, N475, N146);
and AND2 (N480, N476, N262);
xor XOR2 (N481, N477, N394);
or OR4 (N482, N473, N136, N175, N158);
xor XOR2 (N483, N453, N222);
xor XOR2 (N484, N457, N451);
not NOT1 (N485, N464);
and AND2 (N486, N482, N1);
nor NOR3 (N487, N478, N70, N126);
nor NOR4 (N488, N480, N432, N459, N136);
or OR4 (N489, N487, N299, N208, N407);
and AND3 (N490, N481, N421, N157);
not NOT1 (N491, N489);
nand NAND2 (N492, N479, N233);
buf BUF1 (N493, N486);
xor XOR2 (N494, N491, N117);
nand NAND4 (N495, N492, N455, N79, N107);
or OR4 (N496, N485, N289, N44, N430);
nand NAND4 (N497, N474, N250, N221, N43);
nand NAND4 (N498, N490, N55, N436, N332);
and AND2 (N499, N444, N137);
nand NAND4 (N500, N494, N63, N397, N448);
xor XOR2 (N501, N497, N257);
or OR3 (N502, N500, N61, N120);
buf BUF1 (N503, N488);
and AND2 (N504, N496, N209);
nand NAND4 (N505, N495, N183, N96, N134);
and AND2 (N506, N503, N76);
xor XOR2 (N507, N498, N25);
xor XOR2 (N508, N483, N308);
and AND3 (N509, N508, N392, N484);
or OR2 (N510, N19, N48);
or OR4 (N511, N502, N231, N426, N143);
xor XOR2 (N512, N501, N224);
and AND4 (N513, N506, N6, N349, N23);
buf BUF1 (N514, N512);
or OR2 (N515, N510, N114);
and AND2 (N516, N493, N473);
nand NAND3 (N517, N511, N465, N516);
nand NAND3 (N518, N35, N142, N496);
not NOT1 (N519, N505);
buf BUF1 (N520, N504);
not NOT1 (N521, N520);
not NOT1 (N522, N499);
buf BUF1 (N523, N521);
not NOT1 (N524, N518);
or OR4 (N525, N517, N327, N343, N11);
or OR4 (N526, N522, N372, N465, N364);
or OR2 (N527, N525, N282);
nor NOR3 (N528, N524, N200, N134);
and AND4 (N529, N526, N48, N99, N47);
or OR3 (N530, N513, N364, N486);
nand NAND3 (N531, N528, N3, N161);
not NOT1 (N532, N514);
nor NOR3 (N533, N519, N39, N379);
and AND2 (N534, N515, N373);
nor NOR2 (N535, N509, N531);
nor NOR3 (N536, N525, N286, N149);
or OR2 (N537, N535, N455);
buf BUF1 (N538, N527);
not NOT1 (N539, N533);
and AND4 (N540, N530, N11, N60, N174);
xor XOR2 (N541, N536, N160);
buf BUF1 (N542, N523);
not NOT1 (N543, N532);
and AND3 (N544, N542, N484, N157);
not NOT1 (N545, N537);
nor NOR2 (N546, N529, N379);
xor XOR2 (N547, N541, N91);
not NOT1 (N548, N539);
or OR4 (N549, N544, N39, N235, N409);
or OR2 (N550, N546, N271);
nand NAND3 (N551, N549, N289, N120);
not NOT1 (N552, N534);
xor XOR2 (N553, N547, N26);
and AND3 (N554, N550, N426, N449);
and AND3 (N555, N554, N228, N463);
nand NAND2 (N556, N555, N178);
nor NOR4 (N557, N553, N404, N445, N133);
nor NOR2 (N558, N552, N360);
or OR4 (N559, N545, N85, N256, N8);
buf BUF1 (N560, N559);
xor XOR2 (N561, N507, N298);
buf BUF1 (N562, N538);
and AND4 (N563, N548, N225, N247, N201);
and AND2 (N564, N557, N196);
or OR4 (N565, N540, N247, N245, N336);
buf BUF1 (N566, N562);
xor XOR2 (N567, N565, N292);
and AND2 (N568, N560, N424);
or OR3 (N569, N568, N45, N276);
xor XOR2 (N570, N543, N128);
or OR4 (N571, N569, N46, N77, N174);
nor NOR2 (N572, N566, N495);
not NOT1 (N573, N567);
nand NAND3 (N574, N564, N218, N382);
buf BUF1 (N575, N563);
and AND2 (N576, N575, N109);
nor NOR3 (N577, N561, N195, N244);
xor XOR2 (N578, N576, N536);
buf BUF1 (N579, N577);
xor XOR2 (N580, N570, N552);
not NOT1 (N581, N573);
not NOT1 (N582, N580);
nor NOR2 (N583, N574, N386);
nor NOR4 (N584, N581, N135, N408, N101);
nor NOR2 (N585, N584, N442);
xor XOR2 (N586, N585, N367);
nor NOR3 (N587, N583, N445, N284);
and AND4 (N588, N578, N133, N535, N372);
not NOT1 (N589, N571);
nand NAND2 (N590, N586, N125);
or OR4 (N591, N589, N422, N543, N111);
not NOT1 (N592, N556);
nor NOR2 (N593, N558, N527);
xor XOR2 (N594, N590, N478);
buf BUF1 (N595, N588);
not NOT1 (N596, N579);
nor NOR2 (N597, N572, N137);
xor XOR2 (N598, N592, N523);
xor XOR2 (N599, N582, N168);
nor NOR3 (N600, N599, N467, N293);
and AND4 (N601, N596, N361, N18, N424);
nand NAND4 (N602, N600, N66, N343, N327);
or OR2 (N603, N551, N265);
or OR4 (N604, N601, N52, N413, N305);
buf BUF1 (N605, N604);
nor NOR3 (N606, N602, N242, N67);
xor XOR2 (N607, N605, N280);
buf BUF1 (N608, N591);
and AND2 (N609, N608, N420);
not NOT1 (N610, N607);
buf BUF1 (N611, N603);
not NOT1 (N612, N609);
buf BUF1 (N613, N594);
nor NOR3 (N614, N598, N561, N170);
xor XOR2 (N615, N614, N110);
nand NAND3 (N616, N613, N512, N145);
nand NAND4 (N617, N615, N571, N48, N513);
nor NOR2 (N618, N617, N7);
and AND4 (N619, N595, N325, N94, N452);
nand NAND3 (N620, N612, N124, N295);
and AND2 (N621, N611, N432);
xor XOR2 (N622, N619, N73);
or OR4 (N623, N622, N433, N86, N185);
xor XOR2 (N624, N620, N326);
xor XOR2 (N625, N624, N332);
or OR4 (N626, N618, N413, N48, N322);
and AND3 (N627, N610, N535, N357);
xor XOR2 (N628, N616, N467);
not NOT1 (N629, N628);
or OR2 (N630, N597, N33);
nand NAND2 (N631, N623, N288);
nand NAND3 (N632, N606, N239, N213);
not NOT1 (N633, N632);
or OR2 (N634, N631, N166);
nand NAND4 (N635, N625, N305, N367, N46);
xor XOR2 (N636, N621, N354);
or OR4 (N637, N587, N58, N447, N185);
and AND2 (N638, N593, N281);
buf BUF1 (N639, N637);
or OR4 (N640, N639, N198, N197, N106);
buf BUF1 (N641, N635);
not NOT1 (N642, N641);
and AND2 (N643, N634, N429);
not NOT1 (N644, N627);
and AND4 (N645, N626, N613, N453, N213);
xor XOR2 (N646, N636, N579);
xor XOR2 (N647, N638, N454);
buf BUF1 (N648, N630);
nor NOR2 (N649, N644, N49);
or OR3 (N650, N643, N506, N592);
and AND4 (N651, N642, N555, N574, N616);
nand NAND3 (N652, N646, N222, N309);
and AND2 (N653, N650, N573);
nand NAND3 (N654, N649, N14, N591);
not NOT1 (N655, N653);
nor NOR2 (N656, N652, N32);
nand NAND2 (N657, N629, N262);
nand NAND3 (N658, N647, N284, N291);
buf BUF1 (N659, N633);
and AND3 (N660, N655, N420, N344);
buf BUF1 (N661, N660);
nor NOR4 (N662, N657, N71, N222, N497);
buf BUF1 (N663, N661);
and AND2 (N664, N658, N288);
and AND2 (N665, N640, N373);
xor XOR2 (N666, N659, N50);
and AND2 (N667, N648, N517);
nand NAND4 (N668, N651, N402, N216, N597);
not NOT1 (N669, N654);
buf BUF1 (N670, N645);
nor NOR4 (N671, N669, N502, N472, N66);
nand NAND2 (N672, N667, N517);
not NOT1 (N673, N662);
not NOT1 (N674, N670);
and AND4 (N675, N663, N531, N173, N592);
nand NAND2 (N676, N664, N546);
buf BUF1 (N677, N676);
nand NAND4 (N678, N671, N585, N397, N652);
xor XOR2 (N679, N672, N39);
nor NOR3 (N680, N675, N75, N608);
xor XOR2 (N681, N668, N468);
buf BUF1 (N682, N673);
nand NAND2 (N683, N666, N676);
buf BUF1 (N684, N681);
and AND4 (N685, N665, N565, N550, N473);
xor XOR2 (N686, N679, N358);
or OR4 (N687, N680, N131, N233, N26);
and AND4 (N688, N656, N460, N480, N11);
not NOT1 (N689, N687);
buf BUF1 (N690, N684);
buf BUF1 (N691, N677);
and AND4 (N692, N686, N211, N275, N232);
xor XOR2 (N693, N682, N528);
not NOT1 (N694, N692);
buf BUF1 (N695, N693);
nand NAND4 (N696, N688, N287, N354, N62);
not NOT1 (N697, N685);
xor XOR2 (N698, N696, N134);
and AND4 (N699, N697, N137, N649, N412);
not NOT1 (N700, N674);
nand NAND2 (N701, N678, N17);
not NOT1 (N702, N694);
xor XOR2 (N703, N698, N643);
xor XOR2 (N704, N695, N265);
buf BUF1 (N705, N700);
and AND4 (N706, N701, N380, N37, N234);
nor NOR2 (N707, N699, N8);
nor NOR2 (N708, N704, N402);
nand NAND3 (N709, N702, N387, N44);
and AND3 (N710, N709, N605, N241);
not NOT1 (N711, N703);
and AND4 (N712, N683, N392, N513, N223);
endmodule