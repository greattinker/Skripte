// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23;

output N699,N720,N709,N716,N719,N707,N712,N722,N708,N723;

nor NOR2 (N24, N15, N22);
and AND4 (N25, N11, N19, N15, N20);
nand NAND4 (N26, N17, N12, N7, N8);
xor XOR2 (N27, N3, N3);
and AND3 (N28, N4, N12, N1);
buf BUF1 (N29, N24);
not NOT1 (N30, N19);
and AND4 (N31, N26, N20, N2, N15);
not NOT1 (N32, N18);
not NOT1 (N33, N5);
or OR3 (N34, N7, N6, N20);
buf BUF1 (N35, N11);
and AND2 (N36, N27, N12);
or OR3 (N37, N34, N22, N4);
not NOT1 (N38, N32);
not NOT1 (N39, N29);
not NOT1 (N40, N31);
nor NOR4 (N41, N37, N1, N18, N20);
nand NAND3 (N42, N25, N1, N1);
not NOT1 (N43, N41);
xor XOR2 (N44, N39, N40);
or OR4 (N45, N35, N10, N35, N44);
not NOT1 (N46, N9);
nor NOR3 (N47, N2, N11, N46);
not NOT1 (N48, N26);
xor XOR2 (N49, N38, N24);
or OR2 (N50, N30, N34);
nand NAND3 (N51, N47, N35, N43);
buf BUF1 (N52, N39);
xor XOR2 (N53, N36, N36);
nor NOR3 (N54, N51, N49, N22);
xor XOR2 (N55, N46, N51);
or OR4 (N56, N42, N16, N44, N34);
or OR2 (N57, N53, N6);
not NOT1 (N58, N28);
and AND2 (N59, N54, N45);
or OR4 (N60, N34, N21, N17, N21);
not NOT1 (N61, N48);
not NOT1 (N62, N60);
xor XOR2 (N63, N52, N39);
not NOT1 (N64, N33);
and AND2 (N65, N59, N6);
nor NOR4 (N66, N50, N61, N60, N3);
not NOT1 (N67, N42);
and AND4 (N68, N67, N65, N42, N64);
xor XOR2 (N69, N21, N3);
and AND4 (N70, N56, N35, N32, N43);
xor XOR2 (N71, N36, N58);
xor XOR2 (N72, N46, N69);
xor XOR2 (N73, N36, N25);
or OR2 (N74, N68, N61);
nor NOR3 (N75, N70, N8, N33);
xor XOR2 (N76, N63, N56);
buf BUF1 (N77, N71);
not NOT1 (N78, N76);
and AND4 (N79, N62, N77, N55, N45);
buf BUF1 (N80, N4);
and AND4 (N81, N39, N72, N31, N79);
nor NOR2 (N82, N63, N39);
buf BUF1 (N83, N27);
or OR4 (N84, N57, N83, N80, N70);
nor NOR2 (N85, N82, N63);
nand NAND3 (N86, N14, N31, N13);
nor NOR3 (N87, N62, N53, N28);
or OR3 (N88, N85, N18, N37);
xor XOR2 (N89, N73, N74);
xor XOR2 (N90, N64, N40);
and AND3 (N91, N89, N71, N45);
buf BUF1 (N92, N84);
not NOT1 (N93, N78);
or OR2 (N94, N93, N83);
xor XOR2 (N95, N81, N50);
and AND4 (N96, N92, N86, N2, N44);
xor XOR2 (N97, N63, N36);
or OR3 (N98, N97, N97, N71);
or OR4 (N99, N66, N96, N56, N74);
xor XOR2 (N100, N18, N76);
not NOT1 (N101, N100);
or OR3 (N102, N94, N75, N53);
xor XOR2 (N103, N86, N75);
not NOT1 (N104, N91);
nor NOR4 (N105, N88, N83, N12, N51);
buf BUF1 (N106, N98);
buf BUF1 (N107, N102);
nor NOR3 (N108, N90, N107, N91);
buf BUF1 (N109, N58);
nand NAND4 (N110, N103, N99, N45, N100);
xor XOR2 (N111, N101, N32);
not NOT1 (N112, N8);
or OR2 (N113, N87, N88);
nor NOR2 (N114, N105, N108);
not NOT1 (N115, N74);
xor XOR2 (N116, N113, N54);
not NOT1 (N117, N104);
or OR3 (N118, N106, N3, N26);
xor XOR2 (N119, N110, N64);
buf BUF1 (N120, N115);
nand NAND4 (N121, N95, N43, N98, N63);
xor XOR2 (N122, N114, N14);
buf BUF1 (N123, N121);
not NOT1 (N124, N118);
xor XOR2 (N125, N119, N104);
buf BUF1 (N126, N124);
nor NOR4 (N127, N111, N92, N44, N25);
nor NOR4 (N128, N109, N95, N92, N9);
or OR2 (N129, N117, N37);
and AND4 (N130, N127, N94, N71, N129);
not NOT1 (N131, N93);
xor XOR2 (N132, N130, N17);
or OR3 (N133, N126, N36, N74);
nor NOR3 (N134, N132, N96, N51);
not NOT1 (N135, N123);
not NOT1 (N136, N131);
not NOT1 (N137, N128);
or OR3 (N138, N122, N109, N73);
nand NAND3 (N139, N135, N127, N59);
not NOT1 (N140, N138);
nor NOR2 (N141, N133, N75);
xor XOR2 (N142, N112, N60);
and AND2 (N143, N125, N134);
xor XOR2 (N144, N122, N75);
or OR3 (N145, N116, N114, N65);
buf BUF1 (N146, N140);
and AND3 (N147, N141, N43, N78);
not NOT1 (N148, N144);
and AND2 (N149, N148, N142);
nand NAND2 (N150, N13, N36);
nand NAND2 (N151, N147, N110);
xor XOR2 (N152, N150, N89);
nor NOR2 (N153, N143, N147);
buf BUF1 (N154, N120);
nor NOR3 (N155, N137, N62, N13);
and AND4 (N156, N155, N64, N106, N19);
nor NOR2 (N157, N146, N88);
and AND3 (N158, N149, N19, N89);
xor XOR2 (N159, N153, N67);
not NOT1 (N160, N139);
or OR4 (N161, N152, N78, N137, N15);
buf BUF1 (N162, N156);
nand NAND4 (N163, N160, N102, N3, N38);
or OR2 (N164, N151, N40);
nand NAND4 (N165, N154, N87, N58, N48);
nor NOR2 (N166, N165, N141);
xor XOR2 (N167, N166, N82);
or OR4 (N168, N159, N58, N142, N57);
or OR4 (N169, N167, N151, N12, N136);
xor XOR2 (N170, N150, N11);
and AND4 (N171, N169, N143, N113, N159);
and AND2 (N172, N164, N121);
not NOT1 (N173, N170);
nor NOR3 (N174, N163, N44, N67);
buf BUF1 (N175, N168);
nor NOR2 (N176, N173, N59);
nand NAND3 (N177, N145, N70, N37);
not NOT1 (N178, N177);
and AND4 (N179, N162, N24, N148, N28);
nor NOR3 (N180, N178, N76, N122);
and AND4 (N181, N172, N46, N91, N59);
or OR3 (N182, N158, N87, N18);
buf BUF1 (N183, N161);
and AND4 (N184, N183, N86, N81, N136);
buf BUF1 (N185, N180);
nor NOR4 (N186, N184, N33, N23, N88);
not NOT1 (N187, N174);
buf BUF1 (N188, N187);
and AND2 (N189, N182, N91);
nor NOR4 (N190, N175, N149, N88, N156);
and AND4 (N191, N188, N47, N68, N66);
buf BUF1 (N192, N191);
nand NAND3 (N193, N185, N104, N38);
and AND4 (N194, N189, N166, N96, N174);
xor XOR2 (N195, N193, N68);
or OR2 (N196, N171, N32);
nand NAND3 (N197, N186, N132, N103);
nand NAND4 (N198, N179, N35, N180, N121);
xor XOR2 (N199, N181, N100);
or OR4 (N200, N157, N80, N66, N182);
not NOT1 (N201, N200);
and AND3 (N202, N197, N122, N30);
or OR2 (N203, N194, N199);
or OR2 (N204, N152, N56);
buf BUF1 (N205, N198);
xor XOR2 (N206, N192, N65);
or OR2 (N207, N205, N204);
not NOT1 (N208, N115);
nand NAND4 (N209, N208, N182, N156, N6);
and AND3 (N210, N201, N145, N156);
nor NOR3 (N211, N209, N148, N93);
xor XOR2 (N212, N190, N44);
not NOT1 (N213, N210);
not NOT1 (N214, N195);
xor XOR2 (N215, N211, N196);
nor NOR2 (N216, N10, N18);
not NOT1 (N217, N206);
not NOT1 (N218, N203);
not NOT1 (N219, N216);
or OR2 (N220, N218, N45);
buf BUF1 (N221, N213);
buf BUF1 (N222, N215);
or OR3 (N223, N207, N36, N190);
or OR2 (N224, N219, N18);
nor NOR4 (N225, N217, N32, N65, N164);
xor XOR2 (N226, N214, N68);
and AND2 (N227, N221, N211);
xor XOR2 (N228, N176, N114);
or OR4 (N229, N225, N165, N81, N156);
or OR2 (N230, N223, N33);
not NOT1 (N231, N229);
xor XOR2 (N232, N202, N230);
and AND3 (N233, N136, N152, N156);
nor NOR2 (N234, N222, N184);
nand NAND3 (N235, N228, N152, N154);
nor NOR4 (N236, N220, N195, N65, N2);
xor XOR2 (N237, N233, N75);
and AND2 (N238, N237, N202);
or OR2 (N239, N236, N80);
nor NOR4 (N240, N235, N228, N152, N35);
xor XOR2 (N241, N224, N168);
not NOT1 (N242, N239);
nand NAND3 (N243, N234, N76, N4);
and AND4 (N244, N212, N216, N193, N110);
buf BUF1 (N245, N238);
xor XOR2 (N246, N243, N183);
nor NOR2 (N247, N227, N28);
or OR2 (N248, N247, N45);
nand NAND4 (N249, N245, N109, N55, N94);
nor NOR3 (N250, N241, N212, N42);
xor XOR2 (N251, N242, N25);
xor XOR2 (N252, N250, N148);
and AND3 (N253, N240, N14, N156);
and AND4 (N254, N226, N167, N62, N21);
nor NOR4 (N255, N252, N210, N98, N10);
nand NAND2 (N256, N255, N175);
buf BUF1 (N257, N253);
nor NOR3 (N258, N249, N23, N8);
buf BUF1 (N259, N257);
and AND3 (N260, N258, N192, N105);
or OR3 (N261, N232, N105, N215);
not NOT1 (N262, N244);
xor XOR2 (N263, N261, N17);
or OR3 (N264, N260, N141, N64);
nor NOR4 (N265, N262, N166, N72, N95);
and AND2 (N266, N246, N247);
or OR3 (N267, N264, N210, N18);
xor XOR2 (N268, N259, N32);
buf BUF1 (N269, N263);
xor XOR2 (N270, N254, N73);
and AND4 (N271, N269, N23, N231, N63);
buf BUF1 (N272, N73);
xor XOR2 (N273, N272, N212);
or OR2 (N274, N270, N181);
not NOT1 (N275, N268);
xor XOR2 (N276, N274, N210);
xor XOR2 (N277, N256, N243);
nor NOR3 (N278, N267, N78, N109);
not NOT1 (N279, N251);
buf BUF1 (N280, N276);
nand NAND4 (N281, N266, N115, N151, N198);
xor XOR2 (N282, N265, N207);
xor XOR2 (N283, N248, N16);
xor XOR2 (N284, N281, N16);
or OR4 (N285, N284, N95, N270, N198);
and AND2 (N286, N275, N172);
buf BUF1 (N287, N283);
or OR4 (N288, N286, N58, N208, N57);
nor NOR4 (N289, N278, N219, N194, N61);
and AND3 (N290, N273, N134, N131);
nand NAND4 (N291, N289, N28, N68, N165);
xor XOR2 (N292, N271, N241);
and AND4 (N293, N290, N291, N53, N141);
or OR3 (N294, N156, N229, N253);
and AND2 (N295, N279, N81);
and AND4 (N296, N292, N143, N216, N129);
buf BUF1 (N297, N287);
and AND2 (N298, N285, N225);
nand NAND2 (N299, N280, N114);
buf BUF1 (N300, N282);
not NOT1 (N301, N298);
or OR2 (N302, N300, N206);
not NOT1 (N303, N296);
not NOT1 (N304, N277);
nand NAND4 (N305, N288, N273, N144, N291);
or OR3 (N306, N297, N24, N172);
buf BUF1 (N307, N299);
and AND3 (N308, N295, N223, N155);
xor XOR2 (N309, N308, N92);
buf BUF1 (N310, N309);
not NOT1 (N311, N310);
xor XOR2 (N312, N304, N307);
or OR4 (N313, N271, N270, N86, N219);
nor NOR3 (N314, N313, N73, N290);
nand NAND3 (N315, N311, N61, N238);
nand NAND3 (N316, N314, N279, N108);
nor NOR3 (N317, N301, N65, N99);
nand NAND2 (N318, N306, N109);
and AND3 (N319, N316, N259, N110);
xor XOR2 (N320, N303, N251);
nor NOR2 (N321, N319, N134);
buf BUF1 (N322, N302);
buf BUF1 (N323, N318);
nor NOR2 (N324, N305, N71);
not NOT1 (N325, N322);
buf BUF1 (N326, N323);
or OR2 (N327, N320, N77);
or OR2 (N328, N321, N9);
xor XOR2 (N329, N326, N226);
not NOT1 (N330, N317);
nand NAND3 (N331, N312, N205, N242);
and AND3 (N332, N315, N256, N51);
nand NAND4 (N333, N329, N75, N72, N306);
xor XOR2 (N334, N331, N44);
nand NAND2 (N335, N325, N69);
buf BUF1 (N336, N333);
and AND2 (N337, N332, N250);
and AND2 (N338, N328, N101);
nor NOR3 (N339, N335, N122, N316);
and AND2 (N340, N338, N32);
buf BUF1 (N341, N330);
not NOT1 (N342, N336);
xor XOR2 (N343, N341, N141);
buf BUF1 (N344, N343);
nand NAND2 (N345, N334, N209);
nand NAND3 (N346, N293, N302, N96);
buf BUF1 (N347, N337);
buf BUF1 (N348, N327);
or OR2 (N349, N347, N81);
nor NOR2 (N350, N340, N36);
or OR3 (N351, N344, N329, N227);
nor NOR2 (N352, N324, N111);
buf BUF1 (N353, N348);
not NOT1 (N354, N351);
not NOT1 (N355, N354);
or OR4 (N356, N342, N140, N197, N123);
xor XOR2 (N357, N345, N22);
and AND2 (N358, N339, N4);
nor NOR4 (N359, N352, N278, N127, N109);
not NOT1 (N360, N358);
xor XOR2 (N361, N349, N3);
nor NOR4 (N362, N353, N46, N188, N291);
nor NOR2 (N363, N346, N276);
not NOT1 (N364, N362);
nand NAND4 (N365, N364, N352, N117, N172);
and AND3 (N366, N356, N220, N351);
buf BUF1 (N367, N361);
not NOT1 (N368, N355);
buf BUF1 (N369, N367);
not NOT1 (N370, N357);
nor NOR4 (N371, N365, N283, N171, N153);
and AND3 (N372, N366, N265, N111);
buf BUF1 (N373, N370);
xor XOR2 (N374, N369, N306);
nor NOR4 (N375, N374, N27, N83, N115);
not NOT1 (N376, N350);
nand NAND3 (N377, N372, N278, N183);
nand NAND2 (N378, N373, N267);
buf BUF1 (N379, N375);
nor NOR4 (N380, N368, N305, N79, N196);
or OR2 (N381, N360, N376);
nor NOR3 (N382, N289, N110, N59);
xor XOR2 (N383, N294, N148);
not NOT1 (N384, N359);
xor XOR2 (N385, N371, N260);
buf BUF1 (N386, N363);
nor NOR2 (N387, N383, N65);
and AND2 (N388, N378, N92);
nor NOR4 (N389, N386, N38, N345, N183);
and AND2 (N390, N387, N250);
and AND3 (N391, N385, N343, N98);
or OR4 (N392, N382, N77, N377, N104);
nand NAND2 (N393, N215, N337);
buf BUF1 (N394, N393);
nor NOR3 (N395, N379, N179, N300);
or OR2 (N396, N389, N343);
nand NAND4 (N397, N394, N51, N168, N33);
and AND3 (N398, N397, N174, N24);
nand NAND4 (N399, N392, N150, N285, N365);
xor XOR2 (N400, N388, N333);
or OR4 (N401, N380, N369, N163, N69);
xor XOR2 (N402, N400, N127);
buf BUF1 (N403, N402);
and AND2 (N404, N395, N129);
not NOT1 (N405, N403);
and AND2 (N406, N384, N189);
not NOT1 (N407, N390);
and AND3 (N408, N391, N288, N320);
xor XOR2 (N409, N407, N179);
or OR4 (N410, N404, N159, N60, N337);
not NOT1 (N411, N408);
and AND4 (N412, N406, N318, N290, N74);
nand NAND2 (N413, N399, N181);
nor NOR3 (N414, N412, N226, N295);
buf BUF1 (N415, N409);
not NOT1 (N416, N381);
not NOT1 (N417, N398);
buf BUF1 (N418, N414);
and AND3 (N419, N418, N177, N48);
buf BUF1 (N420, N415);
not NOT1 (N421, N405);
nor NOR3 (N422, N396, N173, N23);
nor NOR4 (N423, N420, N309, N143, N117);
xor XOR2 (N424, N423, N154);
xor XOR2 (N425, N411, N398);
nand NAND2 (N426, N416, N98);
or OR3 (N427, N425, N2, N244);
nor NOR2 (N428, N401, N240);
nor NOR2 (N429, N413, N238);
xor XOR2 (N430, N424, N35);
xor XOR2 (N431, N428, N278);
nor NOR4 (N432, N421, N256, N171, N230);
not NOT1 (N433, N432);
not NOT1 (N434, N410);
and AND2 (N435, N427, N72);
nand NAND2 (N436, N435, N231);
not NOT1 (N437, N436);
and AND2 (N438, N419, N299);
buf BUF1 (N439, N433);
nor NOR2 (N440, N439, N115);
buf BUF1 (N441, N440);
xor XOR2 (N442, N437, N245);
not NOT1 (N443, N431);
nor NOR4 (N444, N443, N332, N140, N279);
buf BUF1 (N445, N430);
and AND3 (N446, N442, N329, N276);
buf BUF1 (N447, N446);
xor XOR2 (N448, N444, N169);
buf BUF1 (N449, N441);
and AND3 (N450, N447, N313, N340);
nor NOR4 (N451, N450, N58, N293, N430);
buf BUF1 (N452, N438);
xor XOR2 (N453, N452, N207);
or OR4 (N454, N422, N139, N409, N60);
and AND4 (N455, N417, N16, N446, N294);
buf BUF1 (N456, N448);
or OR4 (N457, N445, N180, N394, N180);
xor XOR2 (N458, N455, N64);
and AND3 (N459, N434, N141, N151);
and AND3 (N460, N429, N67, N384);
or OR4 (N461, N459, N51, N328, N20);
buf BUF1 (N462, N451);
not NOT1 (N463, N454);
buf BUF1 (N464, N462);
and AND2 (N465, N460, N43);
or OR3 (N466, N456, N175, N359);
and AND3 (N467, N426, N106, N307);
xor XOR2 (N468, N467, N10);
nor NOR4 (N469, N461, N14, N218, N37);
and AND3 (N470, N464, N211, N359);
or OR2 (N471, N470, N250);
or OR3 (N472, N466, N188, N362);
buf BUF1 (N473, N472);
nand NAND2 (N474, N453, N20);
nor NOR4 (N475, N471, N299, N229, N285);
or OR3 (N476, N475, N139, N289);
nor NOR2 (N477, N449, N88);
xor XOR2 (N478, N463, N380);
not NOT1 (N479, N457);
or OR4 (N480, N474, N399, N247, N58);
not NOT1 (N481, N480);
xor XOR2 (N482, N479, N146);
nor NOR3 (N483, N469, N94, N386);
nand NAND2 (N484, N483, N410);
xor XOR2 (N485, N458, N81);
nand NAND2 (N486, N485, N430);
xor XOR2 (N487, N481, N125);
or OR4 (N488, N473, N111, N374, N213);
nand NAND4 (N489, N484, N323, N269, N34);
or OR2 (N490, N488, N270);
nor NOR2 (N491, N487, N246);
and AND2 (N492, N468, N451);
not NOT1 (N493, N465);
nand NAND3 (N494, N476, N216, N354);
or OR4 (N495, N493, N383, N35, N490);
xor XOR2 (N496, N203, N193);
not NOT1 (N497, N494);
nor NOR2 (N498, N478, N483);
buf BUF1 (N499, N486);
and AND3 (N500, N477, N315, N78);
xor XOR2 (N501, N492, N445);
xor XOR2 (N502, N498, N418);
nor NOR4 (N503, N501, N495, N128, N367);
buf BUF1 (N504, N382);
and AND2 (N505, N482, N159);
buf BUF1 (N506, N500);
xor XOR2 (N507, N506, N244);
not NOT1 (N508, N504);
or OR4 (N509, N497, N301, N202, N505);
or OR3 (N510, N333, N92, N2);
xor XOR2 (N511, N491, N187);
not NOT1 (N512, N499);
nand NAND4 (N513, N507, N132, N407, N195);
and AND4 (N514, N508, N364, N512, N218);
and AND4 (N515, N416, N287, N180, N509);
not NOT1 (N516, N347);
xor XOR2 (N517, N513, N304);
nand NAND4 (N518, N503, N234, N31, N219);
not NOT1 (N519, N517);
or OR4 (N520, N511, N70, N68, N242);
and AND4 (N521, N496, N353, N65, N17);
not NOT1 (N522, N489);
xor XOR2 (N523, N514, N467);
xor XOR2 (N524, N521, N511);
buf BUF1 (N525, N520);
xor XOR2 (N526, N510, N81);
buf BUF1 (N527, N502);
buf BUF1 (N528, N522);
nor NOR4 (N529, N526, N288, N99, N411);
and AND2 (N530, N523, N256);
not NOT1 (N531, N515);
buf BUF1 (N532, N525);
buf BUF1 (N533, N529);
xor XOR2 (N534, N524, N180);
xor XOR2 (N535, N527, N151);
nand NAND4 (N536, N518, N522, N345, N392);
or OR4 (N537, N535, N440, N131, N166);
and AND2 (N538, N533, N468);
xor XOR2 (N539, N534, N12);
and AND2 (N540, N537, N25);
xor XOR2 (N541, N528, N251);
or OR2 (N542, N541, N175);
not NOT1 (N543, N536);
or OR2 (N544, N539, N254);
nor NOR3 (N545, N538, N183, N265);
and AND4 (N546, N540, N207, N5, N424);
buf BUF1 (N547, N519);
nand NAND3 (N548, N544, N534, N135);
xor XOR2 (N549, N543, N49);
not NOT1 (N550, N546);
and AND2 (N551, N547, N236);
xor XOR2 (N552, N542, N489);
and AND4 (N553, N549, N374, N45, N322);
and AND3 (N554, N516, N107, N56);
and AND4 (N555, N548, N197, N539, N259);
and AND3 (N556, N532, N360, N510);
xor XOR2 (N557, N530, N107);
or OR2 (N558, N550, N284);
not NOT1 (N559, N558);
buf BUF1 (N560, N551);
buf BUF1 (N561, N559);
not NOT1 (N562, N561);
buf BUF1 (N563, N531);
nor NOR2 (N564, N552, N48);
and AND4 (N565, N564, N492, N85, N541);
buf BUF1 (N566, N545);
xor XOR2 (N567, N555, N105);
buf BUF1 (N568, N562);
buf BUF1 (N569, N563);
xor XOR2 (N570, N554, N193);
not NOT1 (N571, N569);
nand NAND3 (N572, N560, N484, N398);
xor XOR2 (N573, N553, N151);
nand NAND2 (N574, N557, N152);
or OR4 (N575, N568, N106, N224, N340);
nor NOR2 (N576, N566, N21);
buf BUF1 (N577, N576);
not NOT1 (N578, N575);
nor NOR4 (N579, N565, N33, N394, N252);
nor NOR2 (N580, N572, N391);
and AND3 (N581, N578, N329, N393);
nor NOR3 (N582, N567, N429, N266);
or OR2 (N583, N579, N504);
xor XOR2 (N584, N580, N406);
xor XOR2 (N585, N584, N447);
xor XOR2 (N586, N556, N127);
nor NOR3 (N587, N585, N465, N572);
nor NOR4 (N588, N583, N311, N19, N227);
xor XOR2 (N589, N587, N423);
buf BUF1 (N590, N589);
or OR2 (N591, N570, N396);
not NOT1 (N592, N577);
buf BUF1 (N593, N581);
or OR2 (N594, N571, N277);
and AND4 (N595, N592, N39, N119, N510);
nand NAND4 (N596, N594, N316, N210, N467);
not NOT1 (N597, N595);
or OR4 (N598, N573, N439, N421, N134);
nor NOR4 (N599, N588, N225, N446, N150);
buf BUF1 (N600, N582);
nand NAND3 (N601, N597, N124, N323);
xor XOR2 (N602, N590, N228);
and AND4 (N603, N586, N59, N36, N522);
xor XOR2 (N604, N601, N410);
xor XOR2 (N605, N596, N360);
buf BUF1 (N606, N598);
or OR4 (N607, N605, N363, N206, N425);
nand NAND2 (N608, N593, N217);
not NOT1 (N609, N591);
not NOT1 (N610, N608);
not NOT1 (N611, N609);
not NOT1 (N612, N611);
nand NAND2 (N613, N612, N348);
nor NOR4 (N614, N606, N320, N590, N244);
or OR4 (N615, N599, N348, N286, N176);
not NOT1 (N616, N607);
and AND2 (N617, N610, N47);
nand NAND4 (N618, N617, N200, N299, N105);
and AND3 (N619, N613, N9, N568);
nand NAND4 (N620, N618, N114, N331, N490);
buf BUF1 (N621, N600);
buf BUF1 (N622, N615);
nand NAND4 (N623, N621, N347, N40, N351);
and AND4 (N624, N623, N455, N26, N521);
nor NOR3 (N625, N602, N464, N395);
buf BUF1 (N626, N616);
nor NOR4 (N627, N625, N125, N65, N312);
or OR3 (N628, N620, N567, N322);
and AND3 (N629, N622, N49, N181);
buf BUF1 (N630, N626);
or OR3 (N631, N603, N6, N423);
and AND3 (N632, N624, N9, N124);
and AND4 (N633, N619, N137, N247, N109);
nor NOR4 (N634, N629, N521, N177, N115);
and AND4 (N635, N614, N504, N607, N83);
nand NAND3 (N636, N635, N234, N223);
or OR4 (N637, N634, N213, N555, N260);
not NOT1 (N638, N637);
nand NAND2 (N639, N638, N145);
and AND2 (N640, N627, N4);
not NOT1 (N641, N632);
or OR2 (N642, N574, N158);
and AND2 (N643, N642, N514);
and AND3 (N644, N641, N70, N297);
or OR4 (N645, N643, N551, N366, N546);
xor XOR2 (N646, N628, N639);
not NOT1 (N647, N628);
nand NAND2 (N648, N636, N351);
or OR3 (N649, N604, N232, N349);
xor XOR2 (N650, N645, N368);
xor XOR2 (N651, N633, N447);
nand NAND4 (N652, N651, N573, N424, N206);
not NOT1 (N653, N646);
xor XOR2 (N654, N631, N8);
nor NOR4 (N655, N653, N361, N226, N379);
not NOT1 (N656, N654);
and AND3 (N657, N656, N502, N124);
buf BUF1 (N658, N644);
not NOT1 (N659, N650);
nand NAND4 (N660, N655, N646, N238, N27);
not NOT1 (N661, N657);
nand NAND2 (N662, N659, N251);
or OR3 (N663, N662, N576, N280);
not NOT1 (N664, N630);
nor NOR3 (N665, N663, N366, N587);
or OR4 (N666, N661, N83, N455, N355);
nor NOR4 (N667, N648, N432, N21, N6);
xor XOR2 (N668, N649, N49);
and AND3 (N669, N665, N157, N209);
nor NOR2 (N670, N668, N71);
and AND3 (N671, N670, N395, N363);
not NOT1 (N672, N666);
and AND4 (N673, N669, N389, N436, N193);
nand NAND3 (N674, N673, N429, N330);
or OR2 (N675, N674, N115);
not NOT1 (N676, N671);
nand NAND2 (N677, N640, N581);
or OR4 (N678, N660, N259, N676, N41);
not NOT1 (N679, N48);
nor NOR4 (N680, N647, N350, N614, N407);
and AND3 (N681, N658, N559, N395);
xor XOR2 (N682, N667, N639);
not NOT1 (N683, N672);
buf BUF1 (N684, N675);
buf BUF1 (N685, N684);
not NOT1 (N686, N679);
not NOT1 (N687, N681);
nand NAND3 (N688, N680, N637, N48);
buf BUF1 (N689, N652);
or OR2 (N690, N689, N663);
xor XOR2 (N691, N678, N283);
nor NOR2 (N692, N682, N584);
buf BUF1 (N693, N690);
xor XOR2 (N694, N664, N588);
and AND2 (N695, N686, N668);
or OR2 (N696, N683, N32);
or OR3 (N697, N685, N577, N393);
and AND4 (N698, N687, N608, N486, N143);
not NOT1 (N699, N696);
nand NAND4 (N700, N695, N134, N278, N691);
xor XOR2 (N701, N486, N627);
nand NAND2 (N702, N688, N446);
xor XOR2 (N703, N701, N529);
buf BUF1 (N704, N697);
not NOT1 (N705, N694);
buf BUF1 (N706, N705);
and AND2 (N707, N704, N483);
not NOT1 (N708, N677);
nor NOR2 (N709, N693, N235);
not NOT1 (N710, N698);
buf BUF1 (N711, N710);
buf BUF1 (N712, N706);
buf BUF1 (N713, N692);
or OR3 (N714, N702, N488, N109);
not NOT1 (N715, N711);
or OR4 (N716, N715, N600, N221, N532);
nand NAND4 (N717, N714, N53, N351, N329);
not NOT1 (N718, N717);
and AND3 (N719, N700, N502, N685);
nand NAND4 (N720, N718, N111, N6, N213);
and AND2 (N721, N713, N715);
xor XOR2 (N722, N721, N530);
and AND4 (N723, N703, N333, N525, N584);
endmodule