// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15;

output N2510,N2499,N2511,N2496,N2512,N2506,N2495,N2513,N2514,N2515;

and AND4 (N16, N13, N3, N2, N8);
or OR2 (N17, N11, N1);
nor NOR4 (N18, N5, N14, N4, N13);
and AND4 (N19, N11, N10, N10, N14);
buf BUF1 (N20, N3);
nor NOR4 (N21, N9, N17, N11, N14);
or OR2 (N22, N15, N21);
nor NOR3 (N23, N3, N13, N12);
or OR2 (N24, N5, N10);
or OR2 (N25, N14, N18);
and AND4 (N26, N3, N1, N13, N11);
buf BUF1 (N27, N18);
or OR2 (N28, N19, N1);
buf BUF1 (N29, N22);
not NOT1 (N30, N22);
nand NAND2 (N31, N25, N18);
nand NAND2 (N32, N23, N16);
and AND3 (N33, N18, N1, N30);
buf BUF1 (N34, N13);
nand NAND2 (N35, N31, N18);
buf BUF1 (N36, N20);
nor NOR3 (N37, N28, N4, N9);
buf BUF1 (N38, N29);
or OR3 (N39, N35, N5, N25);
buf BUF1 (N40, N33);
xor XOR2 (N41, N40, N32);
xor XOR2 (N42, N40, N31);
and AND2 (N43, N27, N21);
or OR2 (N44, N42, N36);
xor XOR2 (N45, N27, N18);
nand NAND3 (N46, N37, N27, N11);
or OR4 (N47, N45, N33, N9, N23);
not NOT1 (N48, N26);
or OR2 (N49, N44, N4);
or OR4 (N50, N41, N2, N37, N42);
buf BUF1 (N51, N24);
or OR4 (N52, N48, N46, N51, N31);
not NOT1 (N53, N13);
or OR4 (N54, N41, N45, N39, N43);
nor NOR2 (N55, N27, N28);
not NOT1 (N56, N29);
and AND4 (N57, N53, N53, N38, N30);
not NOT1 (N58, N3);
not NOT1 (N59, N49);
nand NAND2 (N60, N55, N31);
xor XOR2 (N61, N56, N58);
nor NOR4 (N62, N34, N3, N51, N33);
not NOT1 (N63, N6);
and AND4 (N64, N52, N2, N46, N17);
or OR4 (N65, N50, N35, N56, N2);
and AND3 (N66, N59, N32, N60);
and AND2 (N67, N44, N22);
or OR3 (N68, N54, N8, N45);
nor NOR4 (N69, N65, N16, N3, N13);
xor XOR2 (N70, N63, N61);
or OR3 (N71, N13, N39, N54);
buf BUF1 (N72, N67);
not NOT1 (N73, N69);
buf BUF1 (N74, N72);
buf BUF1 (N75, N66);
or OR3 (N76, N70, N36, N37);
not NOT1 (N77, N47);
xor XOR2 (N78, N62, N26);
nor NOR2 (N79, N73, N24);
nand NAND4 (N80, N68, N43, N17, N68);
not NOT1 (N81, N71);
not NOT1 (N82, N80);
xor XOR2 (N83, N81, N39);
buf BUF1 (N84, N78);
buf BUF1 (N85, N77);
not NOT1 (N86, N57);
or OR3 (N87, N79, N22, N69);
buf BUF1 (N88, N84);
xor XOR2 (N89, N86, N41);
not NOT1 (N90, N82);
not NOT1 (N91, N85);
or OR3 (N92, N88, N12, N6);
buf BUF1 (N93, N89);
xor XOR2 (N94, N87, N69);
buf BUF1 (N95, N74);
nor NOR4 (N96, N90, N25, N9, N16);
buf BUF1 (N97, N75);
and AND3 (N98, N97, N48, N73);
buf BUF1 (N99, N98);
not NOT1 (N100, N91);
buf BUF1 (N101, N96);
nand NAND3 (N102, N95, N10, N28);
buf BUF1 (N103, N99);
not NOT1 (N104, N83);
and AND2 (N105, N64, N55);
nor NOR3 (N106, N76, N98, N19);
or OR4 (N107, N94, N53, N34, N57);
and AND3 (N108, N102, N91, N48);
buf BUF1 (N109, N100);
nor NOR4 (N110, N106, N50, N3, N41);
nor NOR3 (N111, N105, N99, N55);
nor NOR4 (N112, N111, N25, N91, N68);
xor XOR2 (N113, N93, N56);
and AND3 (N114, N108, N86, N109);
or OR4 (N115, N60, N11, N36, N17);
and AND3 (N116, N103, N107, N73);
xor XOR2 (N117, N68, N51);
not NOT1 (N118, N101);
and AND4 (N119, N117, N36, N117, N88);
xor XOR2 (N120, N92, N69);
not NOT1 (N121, N118);
not NOT1 (N122, N113);
xor XOR2 (N123, N120, N51);
not NOT1 (N124, N121);
buf BUF1 (N125, N104);
not NOT1 (N126, N122);
and AND2 (N127, N126, N51);
buf BUF1 (N128, N127);
and AND3 (N129, N115, N36, N98);
nor NOR2 (N130, N125, N53);
not NOT1 (N131, N116);
or OR3 (N132, N112, N73, N38);
nand NAND3 (N133, N131, N113, N130);
and AND2 (N134, N50, N95);
or OR3 (N135, N133, N11, N107);
buf BUF1 (N136, N114);
or OR4 (N137, N124, N50, N114, N129);
not NOT1 (N138, N13);
xor XOR2 (N139, N137, N35);
not NOT1 (N140, N139);
buf BUF1 (N141, N110);
or OR4 (N142, N119, N54, N97, N141);
and AND2 (N143, N77, N99);
nand NAND4 (N144, N135, N83, N18, N66);
not NOT1 (N145, N144);
and AND2 (N146, N132, N52);
or OR3 (N147, N134, N137, N99);
and AND3 (N148, N147, N104, N34);
nand NAND4 (N149, N143, N16, N132, N63);
nor NOR3 (N150, N149, N128, N6);
xor XOR2 (N151, N50, N44);
or OR2 (N152, N140, N132);
and AND4 (N153, N146, N32, N41, N65);
xor XOR2 (N154, N136, N131);
nand NAND3 (N155, N148, N76, N140);
or OR3 (N156, N145, N117, N63);
nand NAND3 (N157, N155, N132, N138);
not NOT1 (N158, N37);
nor NOR2 (N159, N156, N116);
not NOT1 (N160, N158);
buf BUF1 (N161, N160);
buf BUF1 (N162, N150);
and AND2 (N163, N142, N67);
xor XOR2 (N164, N123, N75);
nand NAND4 (N165, N159, N104, N155, N137);
nand NAND2 (N166, N164, N95);
nor NOR2 (N167, N152, N50);
nor NOR2 (N168, N157, N23);
nand NAND3 (N169, N166, N146, N37);
buf BUF1 (N170, N163);
buf BUF1 (N171, N169);
and AND3 (N172, N151, N10, N159);
not NOT1 (N173, N171);
nand NAND3 (N174, N162, N27, N66);
nor NOR4 (N175, N174, N35, N75, N152);
not NOT1 (N176, N172);
nor NOR2 (N177, N175, N44);
or OR2 (N178, N167, N15);
or OR2 (N179, N170, N10);
buf BUF1 (N180, N178);
nand NAND4 (N181, N161, N111, N102, N175);
nor NOR3 (N182, N168, N137, N33);
or OR4 (N183, N177, N5, N75, N83);
or OR2 (N184, N165, N80);
nor NOR2 (N185, N176, N71);
not NOT1 (N186, N183);
not NOT1 (N187, N184);
nand NAND2 (N188, N185, N124);
or OR4 (N189, N179, N74, N155, N104);
or OR2 (N190, N181, N121);
nand NAND2 (N191, N190, N96);
and AND4 (N192, N191, N155, N66, N150);
nor NOR4 (N193, N186, N109, N11, N21);
buf BUF1 (N194, N192);
nor NOR4 (N195, N189, N100, N17, N15);
nor NOR3 (N196, N193, N55, N122);
xor XOR2 (N197, N188, N39);
nor NOR2 (N198, N182, N5);
nor NOR3 (N199, N153, N67, N185);
and AND2 (N200, N154, N102);
buf BUF1 (N201, N200);
and AND3 (N202, N196, N122, N155);
or OR4 (N203, N194, N34, N49, N138);
buf BUF1 (N204, N198);
buf BUF1 (N205, N195);
and AND2 (N206, N173, N86);
xor XOR2 (N207, N206, N67);
nand NAND4 (N208, N199, N21, N2, N85);
and AND2 (N209, N205, N113);
nand NAND4 (N210, N187, N129, N166, N68);
nand NAND3 (N211, N208, N50, N199);
nand NAND2 (N212, N210, N180);
xor XOR2 (N213, N210, N103);
not NOT1 (N214, N203);
buf BUF1 (N215, N202);
nand NAND2 (N216, N207, N143);
not NOT1 (N217, N212);
nand NAND4 (N218, N201, N106, N184, N87);
buf BUF1 (N219, N197);
not NOT1 (N220, N209);
buf BUF1 (N221, N220);
nand NAND4 (N222, N217, N181, N122, N2);
not NOT1 (N223, N222);
buf BUF1 (N224, N214);
nor NOR3 (N225, N204, N83, N12);
nand NAND4 (N226, N223, N122, N182, N39);
xor XOR2 (N227, N216, N89);
or OR3 (N228, N215, N129, N62);
buf BUF1 (N229, N227);
nor NOR2 (N230, N228, N115);
or OR2 (N231, N221, N4);
buf BUF1 (N232, N229);
not NOT1 (N233, N224);
not NOT1 (N234, N211);
not NOT1 (N235, N226);
buf BUF1 (N236, N232);
buf BUF1 (N237, N219);
or OR3 (N238, N218, N96, N4);
xor XOR2 (N239, N233, N176);
buf BUF1 (N240, N230);
nand NAND4 (N241, N238, N71, N99, N188);
and AND4 (N242, N239, N73, N60, N171);
buf BUF1 (N243, N234);
nand NAND3 (N244, N225, N21, N218);
xor XOR2 (N245, N244, N74);
and AND2 (N246, N243, N49);
buf BUF1 (N247, N237);
xor XOR2 (N248, N235, N247);
xor XOR2 (N249, N41, N25);
xor XOR2 (N250, N242, N190);
nor NOR2 (N251, N246, N230);
not NOT1 (N252, N240);
nand NAND3 (N253, N251, N113, N206);
and AND2 (N254, N248, N122);
and AND2 (N255, N245, N101);
buf BUF1 (N256, N249);
not NOT1 (N257, N250);
and AND3 (N258, N253, N91, N143);
buf BUF1 (N259, N258);
nor NOR3 (N260, N236, N224, N72);
xor XOR2 (N261, N256, N127);
buf BUF1 (N262, N261);
nor NOR3 (N263, N231, N53, N189);
or OR4 (N264, N260, N19, N52, N203);
not NOT1 (N265, N262);
buf BUF1 (N266, N257);
nor NOR4 (N267, N254, N201, N112, N10);
nand NAND4 (N268, N259, N234, N236, N121);
nand NAND4 (N269, N241, N187, N93, N148);
and AND2 (N270, N266, N245);
nor NOR3 (N271, N255, N262, N143);
and AND4 (N272, N213, N112, N168, N141);
or OR2 (N273, N272, N83);
nand NAND3 (N274, N273, N72, N250);
nand NAND4 (N275, N263, N261, N85, N245);
buf BUF1 (N276, N268);
not NOT1 (N277, N270);
not NOT1 (N278, N269);
or OR2 (N279, N276, N19);
or OR3 (N280, N271, N196, N89);
xor XOR2 (N281, N275, N212);
nor NOR4 (N282, N281, N89, N26, N146);
not NOT1 (N283, N277);
nand NAND2 (N284, N283, N205);
or OR2 (N285, N280, N179);
not NOT1 (N286, N285);
nor NOR4 (N287, N267, N242, N45, N48);
nor NOR2 (N288, N274, N83);
buf BUF1 (N289, N287);
buf BUF1 (N290, N278);
or OR2 (N291, N290, N219);
not NOT1 (N292, N279);
xor XOR2 (N293, N289, N104);
not NOT1 (N294, N293);
nor NOR3 (N295, N265, N18, N87);
nand NAND2 (N296, N288, N294);
xor XOR2 (N297, N233, N222);
not NOT1 (N298, N282);
nor NOR3 (N299, N286, N195, N7);
or OR3 (N300, N295, N247, N56);
xor XOR2 (N301, N252, N242);
xor XOR2 (N302, N291, N73);
buf BUF1 (N303, N264);
xor XOR2 (N304, N302, N232);
or OR4 (N305, N296, N144, N99, N42);
buf BUF1 (N306, N303);
nand NAND3 (N307, N298, N47, N202);
nor NOR2 (N308, N307, N257);
or OR4 (N309, N284, N109, N178, N126);
nor NOR2 (N310, N297, N121);
xor XOR2 (N311, N309, N241);
and AND4 (N312, N301, N263, N107, N204);
nor NOR4 (N313, N312, N95, N305, N300);
and AND4 (N314, N135, N115, N297, N54);
buf BUF1 (N315, N289);
nand NAND4 (N316, N306, N102, N212, N42);
and AND2 (N317, N316, N169);
and AND4 (N318, N314, N80, N250, N305);
buf BUF1 (N319, N308);
or OR2 (N320, N319, N311);
nand NAND4 (N321, N234, N31, N173, N29);
not NOT1 (N322, N317);
nor NOR4 (N323, N310, N230, N140, N216);
or OR2 (N324, N320, N234);
buf BUF1 (N325, N318);
buf BUF1 (N326, N315);
and AND4 (N327, N324, N273, N137, N309);
or OR4 (N328, N325, N310, N253, N315);
not NOT1 (N329, N299);
xor XOR2 (N330, N326, N178);
or OR3 (N331, N328, N181, N263);
and AND3 (N332, N321, N319, N146);
nor NOR4 (N333, N330, N119, N302, N71);
nor NOR4 (N334, N322, N291, N252, N228);
not NOT1 (N335, N292);
buf BUF1 (N336, N335);
nand NAND4 (N337, N332, N225, N150, N73);
or OR4 (N338, N333, N310, N310, N327);
and AND3 (N339, N318, N275, N209);
not NOT1 (N340, N329);
nor NOR2 (N341, N336, N32);
nand NAND3 (N342, N304, N33, N244);
not NOT1 (N343, N339);
xor XOR2 (N344, N323, N302);
buf BUF1 (N345, N334);
xor XOR2 (N346, N340, N70);
and AND3 (N347, N337, N301, N203);
and AND2 (N348, N346, N281);
or OR4 (N349, N341, N135, N229, N249);
xor XOR2 (N350, N343, N21);
or OR4 (N351, N338, N251, N7, N310);
buf BUF1 (N352, N344);
not NOT1 (N353, N352);
xor XOR2 (N354, N350, N98);
nand NAND3 (N355, N353, N334, N144);
and AND2 (N356, N354, N227);
nor NOR3 (N357, N345, N4, N57);
xor XOR2 (N358, N355, N37);
buf BUF1 (N359, N356);
not NOT1 (N360, N349);
xor XOR2 (N361, N331, N315);
xor XOR2 (N362, N342, N37);
buf BUF1 (N363, N351);
xor XOR2 (N364, N361, N281);
nand NAND3 (N365, N360, N308, N188);
or OR2 (N366, N347, N325);
nor NOR3 (N367, N359, N328, N98);
or OR2 (N368, N364, N267);
nand NAND4 (N369, N367, N21, N288, N148);
not NOT1 (N370, N368);
buf BUF1 (N371, N366);
or OR2 (N372, N365, N78);
and AND3 (N373, N358, N14, N369);
nand NAND4 (N374, N179, N348, N144, N177);
buf BUF1 (N375, N355);
nand NAND4 (N376, N374, N319, N365, N346);
not NOT1 (N377, N376);
xor XOR2 (N378, N362, N8);
and AND4 (N379, N371, N376, N14, N297);
and AND2 (N380, N377, N122);
xor XOR2 (N381, N378, N171);
xor XOR2 (N382, N372, N326);
not NOT1 (N383, N357);
xor XOR2 (N384, N382, N187);
xor XOR2 (N385, N380, N98);
nor NOR2 (N386, N381, N160);
buf BUF1 (N387, N379);
not NOT1 (N388, N386);
nor NOR3 (N389, N375, N304, N333);
buf BUF1 (N390, N383);
nand NAND4 (N391, N385, N68, N176, N163);
nor NOR4 (N392, N390, N197, N336, N354);
nor NOR4 (N393, N363, N291, N202, N35);
xor XOR2 (N394, N387, N182);
xor XOR2 (N395, N389, N236);
nor NOR4 (N396, N395, N109, N57, N178);
or OR4 (N397, N392, N271, N116, N87);
nand NAND3 (N398, N393, N277, N331);
xor XOR2 (N399, N394, N328);
or OR2 (N400, N388, N346);
nor NOR2 (N401, N384, N9);
and AND4 (N402, N373, N340, N149, N297);
and AND4 (N403, N391, N291, N358, N272);
nand NAND4 (N404, N399, N270, N29, N107);
or OR3 (N405, N313, N49, N371);
nand NAND4 (N406, N400, N165, N364, N29);
buf BUF1 (N407, N403);
nand NAND4 (N408, N370, N102, N378, N169);
nand NAND2 (N409, N398, N294);
nand NAND4 (N410, N407, N119, N115, N196);
nor NOR2 (N411, N410, N43);
xor XOR2 (N412, N404, N377);
nand NAND3 (N413, N405, N212, N397);
not NOT1 (N414, N8);
buf BUF1 (N415, N396);
or OR2 (N416, N412, N57);
nor NOR2 (N417, N411, N273);
or OR3 (N418, N401, N324, N384);
xor XOR2 (N419, N406, N290);
not NOT1 (N420, N418);
buf BUF1 (N421, N417);
or OR3 (N422, N409, N284, N10);
or OR3 (N423, N420, N206, N220);
and AND4 (N424, N419, N284, N117, N328);
or OR4 (N425, N423, N333, N10, N205);
nor NOR2 (N426, N414, N159);
xor XOR2 (N427, N413, N145);
and AND2 (N428, N415, N87);
and AND2 (N429, N424, N374);
nor NOR3 (N430, N425, N50, N98);
buf BUF1 (N431, N422);
or OR4 (N432, N408, N293, N208, N345);
and AND2 (N433, N427, N320);
nor NOR3 (N434, N432, N329, N338);
xor XOR2 (N435, N428, N157);
nor NOR4 (N436, N433, N433, N24, N125);
and AND2 (N437, N426, N175);
or OR2 (N438, N437, N136);
nand NAND4 (N439, N431, N206, N7, N26);
nor NOR2 (N440, N416, N350);
nand NAND3 (N441, N429, N244, N373);
buf BUF1 (N442, N438);
or OR3 (N443, N439, N294, N116);
nand NAND4 (N444, N430, N440, N346, N364);
buf BUF1 (N445, N221);
not NOT1 (N446, N436);
and AND4 (N447, N444, N136, N352, N409);
not NOT1 (N448, N402);
not NOT1 (N449, N446);
not NOT1 (N450, N421);
buf BUF1 (N451, N434);
and AND4 (N452, N441, N416, N332, N246);
buf BUF1 (N453, N450);
or OR2 (N454, N443, N78);
nor NOR4 (N455, N454, N333, N117, N445);
nand NAND3 (N456, N4, N367, N32);
xor XOR2 (N457, N449, N436);
or OR4 (N458, N447, N385, N390, N22);
not NOT1 (N459, N457);
buf BUF1 (N460, N452);
not NOT1 (N461, N458);
or OR4 (N462, N459, N402, N133, N120);
nand NAND4 (N463, N456, N402, N406, N50);
or OR4 (N464, N435, N406, N56, N37);
or OR2 (N465, N462, N259);
nand NAND4 (N466, N465, N73, N8, N19);
and AND2 (N467, N442, N102);
buf BUF1 (N468, N451);
buf BUF1 (N469, N463);
or OR2 (N470, N448, N203);
buf BUF1 (N471, N455);
nand NAND4 (N472, N471, N397, N192, N330);
and AND4 (N473, N472, N203, N258, N43);
and AND2 (N474, N460, N149);
or OR3 (N475, N468, N462, N119);
nand NAND3 (N476, N467, N47, N168);
nor NOR3 (N477, N476, N237, N69);
xor XOR2 (N478, N466, N301);
or OR2 (N479, N474, N81);
and AND2 (N480, N453, N215);
xor XOR2 (N481, N464, N143);
not NOT1 (N482, N461);
not NOT1 (N483, N479);
buf BUF1 (N484, N470);
nand NAND3 (N485, N475, N244, N110);
not NOT1 (N486, N469);
buf BUF1 (N487, N478);
and AND3 (N488, N483, N294, N89);
and AND3 (N489, N481, N117, N458);
buf BUF1 (N490, N480);
not NOT1 (N491, N487);
or OR2 (N492, N485, N414);
not NOT1 (N493, N492);
xor XOR2 (N494, N488, N464);
nand NAND4 (N495, N473, N245, N415, N322);
and AND4 (N496, N486, N201, N347, N391);
or OR3 (N497, N477, N258, N274);
nand NAND4 (N498, N496, N455, N241, N257);
buf BUF1 (N499, N491);
or OR3 (N500, N497, N367, N433);
nor NOR4 (N501, N500, N460, N242, N11);
or OR4 (N502, N489, N154, N473, N139);
or OR4 (N503, N502, N379, N399, N474);
or OR3 (N504, N493, N54, N59);
and AND3 (N505, N503, N504, N382);
nand NAND3 (N506, N50, N326, N203);
nor NOR3 (N507, N490, N471, N501);
buf BUF1 (N508, N409);
xor XOR2 (N509, N498, N15);
and AND3 (N510, N494, N369, N123);
xor XOR2 (N511, N510, N377);
xor XOR2 (N512, N506, N73);
nor NOR2 (N513, N505, N238);
nor NOR3 (N514, N512, N436, N481);
nor NOR2 (N515, N495, N139);
not NOT1 (N516, N511);
not NOT1 (N517, N514);
not NOT1 (N518, N482);
buf BUF1 (N519, N507);
and AND4 (N520, N509, N289, N236, N449);
xor XOR2 (N521, N508, N118);
or OR4 (N522, N484, N158, N97, N488);
nor NOR4 (N523, N516, N240, N520, N498);
buf BUF1 (N524, N270);
buf BUF1 (N525, N515);
buf BUF1 (N526, N523);
and AND2 (N527, N518, N432);
xor XOR2 (N528, N519, N210);
buf BUF1 (N529, N517);
buf BUF1 (N530, N499);
xor XOR2 (N531, N525, N516);
or OR2 (N532, N524, N179);
and AND2 (N533, N531, N352);
or OR3 (N534, N533, N119, N9);
and AND4 (N535, N513, N245, N269, N446);
or OR4 (N536, N528, N150, N321, N109);
and AND2 (N537, N527, N515);
xor XOR2 (N538, N522, N28);
nor NOR3 (N539, N534, N33, N112);
xor XOR2 (N540, N521, N298);
buf BUF1 (N541, N538);
xor XOR2 (N542, N530, N96);
xor XOR2 (N543, N536, N393);
and AND2 (N544, N535, N348);
nor NOR4 (N545, N539, N78, N241, N449);
not NOT1 (N546, N544);
nand NAND4 (N547, N532, N50, N301, N393);
buf BUF1 (N548, N546);
and AND4 (N549, N547, N172, N66, N163);
not NOT1 (N550, N537);
nor NOR3 (N551, N545, N460, N314);
not NOT1 (N552, N550);
nor NOR4 (N553, N540, N314, N516, N438);
xor XOR2 (N554, N551, N347);
nor NOR4 (N555, N552, N63, N418, N319);
not NOT1 (N556, N548);
not NOT1 (N557, N549);
not NOT1 (N558, N554);
buf BUF1 (N559, N553);
nand NAND3 (N560, N559, N126, N159);
xor XOR2 (N561, N555, N24);
or OR2 (N562, N529, N452);
and AND2 (N563, N541, N189);
nand NAND2 (N564, N562, N179);
not NOT1 (N565, N563);
nand NAND3 (N566, N556, N97, N214);
nor NOR2 (N567, N561, N5);
nor NOR4 (N568, N543, N51, N111, N86);
buf BUF1 (N569, N557);
not NOT1 (N570, N564);
not NOT1 (N571, N566);
or OR3 (N572, N568, N153, N518);
or OR2 (N573, N571, N329);
and AND4 (N574, N560, N69, N255, N237);
xor XOR2 (N575, N542, N484);
and AND3 (N576, N567, N73, N234);
nor NOR3 (N577, N526, N31, N470);
and AND3 (N578, N570, N286, N154);
nand NAND3 (N579, N558, N254, N191);
nand NAND2 (N580, N573, N513);
buf BUF1 (N581, N574);
and AND2 (N582, N575, N204);
nand NAND4 (N583, N582, N383, N37, N109);
xor XOR2 (N584, N579, N140);
and AND4 (N585, N569, N309, N414, N245);
buf BUF1 (N586, N581);
buf BUF1 (N587, N580);
and AND3 (N588, N576, N290, N19);
nor NOR2 (N589, N577, N253);
not NOT1 (N590, N585);
buf BUF1 (N591, N590);
and AND2 (N592, N588, N373);
buf BUF1 (N593, N591);
not NOT1 (N594, N578);
or OR4 (N595, N594, N120, N563, N256);
not NOT1 (N596, N586);
or OR2 (N597, N587, N121);
nor NOR4 (N598, N583, N108, N564, N303);
and AND2 (N599, N593, N322);
buf BUF1 (N600, N596);
xor XOR2 (N601, N599, N342);
nor NOR3 (N602, N595, N291, N270);
nand NAND3 (N603, N600, N21, N216);
not NOT1 (N604, N589);
or OR3 (N605, N584, N371, N380);
or OR4 (N606, N604, N411, N302, N129);
xor XOR2 (N607, N572, N419);
buf BUF1 (N608, N603);
nor NOR3 (N609, N565, N72, N301);
buf BUF1 (N610, N592);
buf BUF1 (N611, N609);
nand NAND2 (N612, N597, N298);
buf BUF1 (N613, N608);
buf BUF1 (N614, N602);
and AND2 (N615, N613, N520);
not NOT1 (N616, N614);
not NOT1 (N617, N601);
xor XOR2 (N618, N615, N119);
or OR3 (N619, N617, N552, N504);
or OR2 (N620, N607, N59);
nand NAND2 (N621, N619, N467);
or OR3 (N622, N621, N46, N208);
or OR2 (N623, N616, N520);
buf BUF1 (N624, N598);
nor NOR4 (N625, N618, N59, N190, N193);
buf BUF1 (N626, N623);
buf BUF1 (N627, N624);
not NOT1 (N628, N612);
nor NOR4 (N629, N610, N345, N8, N298);
buf BUF1 (N630, N628);
not NOT1 (N631, N611);
xor XOR2 (N632, N626, N338);
nor NOR3 (N633, N630, N233, N521);
xor XOR2 (N634, N629, N220);
not NOT1 (N635, N620);
and AND3 (N636, N635, N77, N17);
or OR4 (N637, N631, N302, N243, N506);
and AND2 (N638, N633, N409);
and AND3 (N639, N622, N544, N252);
and AND2 (N640, N625, N197);
nor NOR2 (N641, N638, N54);
or OR2 (N642, N639, N402);
nand NAND3 (N643, N627, N593, N54);
xor XOR2 (N644, N637, N460);
or OR4 (N645, N642, N508, N417, N273);
nand NAND3 (N646, N605, N135, N602);
and AND3 (N647, N644, N305, N480);
buf BUF1 (N648, N640);
or OR2 (N649, N647, N4);
xor XOR2 (N650, N634, N620);
buf BUF1 (N651, N643);
nor NOR2 (N652, N650, N211);
or OR4 (N653, N636, N233, N400, N524);
and AND3 (N654, N649, N530, N10);
buf BUF1 (N655, N654);
not NOT1 (N656, N652);
not NOT1 (N657, N632);
or OR2 (N658, N651, N150);
or OR2 (N659, N648, N355);
nor NOR2 (N660, N653, N581);
not NOT1 (N661, N646);
xor XOR2 (N662, N656, N117);
nand NAND4 (N663, N662, N242, N101, N635);
nor NOR2 (N664, N606, N493);
nand NAND3 (N665, N641, N118, N33);
and AND3 (N666, N665, N319, N227);
or OR4 (N667, N660, N588, N550, N589);
not NOT1 (N668, N666);
buf BUF1 (N669, N658);
buf BUF1 (N670, N661);
not NOT1 (N671, N668);
nor NOR4 (N672, N671, N477, N374, N131);
not NOT1 (N673, N657);
nand NAND3 (N674, N670, N434, N361);
and AND2 (N675, N659, N539);
nor NOR3 (N676, N655, N343, N473);
not NOT1 (N677, N675);
or OR4 (N678, N669, N600, N623, N77);
or OR3 (N679, N672, N534, N187);
and AND3 (N680, N663, N169, N44);
not NOT1 (N681, N674);
not NOT1 (N682, N676);
not NOT1 (N683, N645);
nor NOR3 (N684, N677, N255, N53);
buf BUF1 (N685, N681);
not NOT1 (N686, N678);
and AND3 (N687, N664, N624, N448);
nor NOR4 (N688, N683, N539, N459, N522);
not NOT1 (N689, N682);
and AND3 (N690, N667, N371, N32);
nand NAND2 (N691, N679, N351);
nand NAND2 (N692, N690, N480);
nand NAND3 (N693, N673, N287, N569);
nand NAND4 (N694, N684, N227, N518, N407);
nand NAND3 (N695, N692, N394, N206);
or OR4 (N696, N695, N465, N5, N474);
not NOT1 (N697, N686);
xor XOR2 (N698, N696, N74);
nor NOR4 (N699, N687, N290, N141, N627);
nand NAND3 (N700, N685, N187, N197);
not NOT1 (N701, N691);
and AND2 (N702, N688, N362);
xor XOR2 (N703, N698, N246);
nand NAND2 (N704, N701, N498);
xor XOR2 (N705, N680, N93);
and AND2 (N706, N697, N620);
buf BUF1 (N707, N702);
or OR3 (N708, N700, N494, N238);
xor XOR2 (N709, N705, N495);
xor XOR2 (N710, N693, N349);
buf BUF1 (N711, N689);
buf BUF1 (N712, N708);
not NOT1 (N713, N694);
nor NOR4 (N714, N699, N356, N557, N492);
nor NOR3 (N715, N713, N168, N501);
nor NOR2 (N716, N710, N321);
not NOT1 (N717, N704);
xor XOR2 (N718, N706, N136);
or OR4 (N719, N712, N292, N414, N109);
and AND3 (N720, N719, N432, N381);
or OR4 (N721, N703, N582, N717, N22);
xor XOR2 (N722, N408, N478);
not NOT1 (N723, N709);
and AND2 (N724, N716, N154);
buf BUF1 (N725, N707);
and AND4 (N726, N715, N569, N685, N39);
not NOT1 (N727, N711);
or OR3 (N728, N726, N426, N197);
or OR3 (N729, N718, N468, N127);
or OR4 (N730, N727, N528, N300, N209);
nand NAND3 (N731, N728, N559, N329);
or OR2 (N732, N731, N187);
xor XOR2 (N733, N730, N436);
buf BUF1 (N734, N721);
not NOT1 (N735, N725);
xor XOR2 (N736, N720, N387);
xor XOR2 (N737, N729, N65);
not NOT1 (N738, N737);
or OR4 (N739, N714, N528, N8, N86);
xor XOR2 (N740, N736, N516);
buf BUF1 (N741, N734);
xor XOR2 (N742, N735, N223);
xor XOR2 (N743, N739, N538);
nand NAND4 (N744, N740, N303, N427, N496);
nor NOR2 (N745, N723, N78);
or OR3 (N746, N722, N671, N144);
xor XOR2 (N747, N738, N96);
nand NAND4 (N748, N744, N460, N232, N708);
buf BUF1 (N749, N742);
or OR4 (N750, N749, N559, N175, N403);
buf BUF1 (N751, N750);
and AND3 (N752, N733, N494, N225);
nor NOR4 (N753, N747, N295, N28, N299);
nor NOR2 (N754, N753, N238);
buf BUF1 (N755, N745);
or OR2 (N756, N732, N29);
xor XOR2 (N757, N743, N33);
and AND4 (N758, N746, N238, N514, N92);
buf BUF1 (N759, N741);
nor NOR3 (N760, N755, N286, N620);
not NOT1 (N761, N752);
or OR2 (N762, N754, N247);
or OR2 (N763, N756, N479);
nand NAND3 (N764, N757, N382, N719);
nor NOR2 (N765, N760, N612);
not NOT1 (N766, N759);
buf BUF1 (N767, N763);
and AND3 (N768, N761, N742, N102);
xor XOR2 (N769, N724, N39);
or OR3 (N770, N748, N603, N255);
or OR2 (N771, N768, N331);
buf BUF1 (N772, N764);
nand NAND3 (N773, N751, N118, N388);
nand NAND3 (N774, N766, N64, N27);
or OR2 (N775, N772, N1);
buf BUF1 (N776, N770);
or OR4 (N777, N765, N197, N50, N5);
xor XOR2 (N778, N762, N301);
not NOT1 (N779, N776);
and AND4 (N780, N775, N770, N601, N388);
or OR2 (N781, N779, N621);
xor XOR2 (N782, N769, N734);
and AND4 (N783, N767, N158, N119, N14);
and AND3 (N784, N758, N218, N86);
buf BUF1 (N785, N771);
xor XOR2 (N786, N783, N339);
or OR4 (N787, N781, N233, N640, N245);
and AND4 (N788, N785, N126, N609, N32);
xor XOR2 (N789, N788, N192);
nor NOR4 (N790, N786, N182, N600, N585);
xor XOR2 (N791, N780, N687);
and AND4 (N792, N791, N417, N190, N743);
not NOT1 (N793, N790);
or OR2 (N794, N774, N200);
nand NAND2 (N795, N784, N28);
nand NAND2 (N796, N794, N155);
xor XOR2 (N797, N796, N387);
not NOT1 (N798, N795);
buf BUF1 (N799, N777);
not NOT1 (N800, N798);
not NOT1 (N801, N799);
nor NOR3 (N802, N782, N393, N537);
nor NOR2 (N803, N801, N664);
xor XOR2 (N804, N773, N492);
or OR4 (N805, N789, N424, N790, N440);
nand NAND3 (N806, N797, N755, N658);
and AND4 (N807, N804, N1, N596, N129);
nor NOR4 (N808, N800, N129, N507, N751);
buf BUF1 (N809, N803);
or OR4 (N810, N793, N517, N581, N182);
or OR4 (N811, N805, N324, N626, N626);
or OR3 (N812, N808, N484, N564);
and AND2 (N813, N811, N61);
nand NAND2 (N814, N812, N677);
nand NAND3 (N815, N806, N439, N430);
or OR4 (N816, N787, N312, N631, N207);
not NOT1 (N817, N807);
nand NAND2 (N818, N809, N81);
not NOT1 (N819, N778);
buf BUF1 (N820, N810);
not NOT1 (N821, N815);
buf BUF1 (N822, N816);
or OR4 (N823, N792, N641, N738, N101);
and AND3 (N824, N821, N800, N253);
xor XOR2 (N825, N817, N269);
and AND3 (N826, N813, N186, N279);
xor XOR2 (N827, N814, N174);
nor NOR3 (N828, N822, N771, N328);
not NOT1 (N829, N825);
nor NOR4 (N830, N819, N727, N277, N734);
buf BUF1 (N831, N823);
not NOT1 (N832, N829);
and AND2 (N833, N830, N399);
or OR3 (N834, N824, N54, N639);
and AND3 (N835, N826, N337, N472);
xor XOR2 (N836, N833, N628);
nand NAND3 (N837, N827, N453, N706);
xor XOR2 (N838, N832, N452);
and AND3 (N839, N820, N498, N245);
not NOT1 (N840, N818);
not NOT1 (N841, N831);
nand NAND2 (N842, N802, N385);
xor XOR2 (N843, N841, N330);
or OR4 (N844, N839, N119, N555, N828);
buf BUF1 (N845, N265);
nand NAND4 (N846, N834, N32, N684, N314);
and AND4 (N847, N842, N485, N422, N52);
buf BUF1 (N848, N843);
nor NOR4 (N849, N844, N54, N614, N517);
or OR4 (N850, N845, N296, N703, N654);
or OR2 (N851, N838, N770);
or OR2 (N852, N850, N618);
and AND2 (N853, N848, N41);
not NOT1 (N854, N852);
or OR3 (N855, N854, N751, N729);
or OR2 (N856, N840, N557);
or OR3 (N857, N849, N187, N609);
nor NOR2 (N858, N847, N558);
nor NOR4 (N859, N851, N853, N62, N646);
buf BUF1 (N860, N434);
and AND2 (N861, N836, N615);
not NOT1 (N862, N857);
nand NAND4 (N863, N861, N844, N631, N73);
and AND3 (N864, N859, N110, N131);
not NOT1 (N865, N863);
and AND3 (N866, N865, N145, N434);
nand NAND3 (N867, N866, N178, N333);
and AND3 (N868, N846, N636, N511);
nor NOR2 (N869, N860, N223);
buf BUF1 (N870, N868);
and AND2 (N871, N867, N390);
or OR3 (N872, N864, N766, N645);
or OR2 (N873, N856, N171);
not NOT1 (N874, N858);
nand NAND2 (N875, N871, N183);
nand NAND2 (N876, N869, N410);
buf BUF1 (N877, N855);
and AND3 (N878, N877, N228, N69);
and AND3 (N879, N878, N53, N586);
and AND4 (N880, N875, N795, N180, N256);
nor NOR2 (N881, N835, N340);
or OR4 (N882, N874, N786, N878, N127);
not NOT1 (N883, N880);
nor NOR3 (N884, N872, N70, N322);
and AND4 (N885, N881, N231, N184, N181);
buf BUF1 (N886, N876);
and AND4 (N887, N879, N794, N34, N33);
and AND4 (N888, N886, N765, N825, N513);
xor XOR2 (N889, N873, N481);
or OR3 (N890, N882, N372, N348);
or OR3 (N891, N883, N14, N584);
buf BUF1 (N892, N884);
xor XOR2 (N893, N889, N190);
buf BUF1 (N894, N892);
and AND4 (N895, N837, N474, N863, N60);
and AND2 (N896, N888, N718);
and AND3 (N897, N862, N257, N425);
xor XOR2 (N898, N896, N224);
buf BUF1 (N899, N893);
nor NOR4 (N900, N898, N66, N10, N166);
xor XOR2 (N901, N885, N668);
or OR4 (N902, N870, N623, N475, N594);
not NOT1 (N903, N895);
and AND3 (N904, N894, N169, N481);
nor NOR4 (N905, N902, N41, N143, N446);
buf BUF1 (N906, N887);
nor NOR2 (N907, N904, N196);
nor NOR3 (N908, N901, N726, N19);
xor XOR2 (N909, N897, N80);
buf BUF1 (N910, N906);
and AND3 (N911, N899, N85, N889);
and AND3 (N912, N900, N584, N457);
not NOT1 (N913, N910);
not NOT1 (N914, N905);
xor XOR2 (N915, N914, N419);
nor NOR3 (N916, N912, N225, N568);
xor XOR2 (N917, N916, N72);
and AND2 (N918, N907, N722);
not NOT1 (N919, N911);
nor NOR3 (N920, N903, N430, N657);
xor XOR2 (N921, N919, N167);
nand NAND3 (N922, N921, N858, N468);
xor XOR2 (N923, N909, N797);
xor XOR2 (N924, N908, N66);
buf BUF1 (N925, N891);
and AND3 (N926, N917, N726, N99);
nor NOR4 (N927, N913, N149, N748, N825);
not NOT1 (N928, N923);
and AND4 (N929, N918, N511, N803, N688);
or OR4 (N930, N927, N798, N771, N621);
nor NOR3 (N931, N930, N908, N684);
buf BUF1 (N932, N890);
xor XOR2 (N933, N925, N874);
nand NAND2 (N934, N931, N384);
or OR4 (N935, N922, N230, N934, N413);
nand NAND2 (N936, N526, N232);
or OR4 (N937, N936, N385, N115, N882);
and AND2 (N938, N929, N240);
and AND4 (N939, N915, N113, N839, N518);
nand NAND2 (N940, N926, N313);
not NOT1 (N941, N933);
nor NOR2 (N942, N941, N595);
xor XOR2 (N943, N940, N97);
nand NAND3 (N944, N924, N320, N446);
xor XOR2 (N945, N920, N870);
nor NOR4 (N946, N935, N483, N583, N791);
not NOT1 (N947, N937);
buf BUF1 (N948, N944);
nor NOR4 (N949, N938, N577, N236, N305);
or OR4 (N950, N928, N364, N682, N879);
and AND3 (N951, N948, N519, N299);
not NOT1 (N952, N945);
not NOT1 (N953, N946);
or OR3 (N954, N949, N132, N537);
or OR3 (N955, N951, N79, N855);
and AND2 (N956, N953, N820);
or OR3 (N957, N955, N668, N72);
nor NOR4 (N958, N954, N922, N689, N567);
buf BUF1 (N959, N950);
and AND2 (N960, N943, N874);
or OR3 (N961, N932, N377, N78);
and AND4 (N962, N939, N568, N715, N697);
or OR2 (N963, N962, N132);
or OR4 (N964, N957, N656, N510, N524);
buf BUF1 (N965, N952);
nor NOR4 (N966, N960, N321, N20, N763);
nor NOR2 (N967, N956, N878);
nand NAND3 (N968, N963, N648, N643);
nor NOR4 (N969, N961, N22, N304, N71);
and AND4 (N970, N968, N122, N284, N185);
or OR3 (N971, N959, N968, N783);
nand NAND4 (N972, N967, N175, N447, N464);
not NOT1 (N973, N971);
not NOT1 (N974, N965);
and AND2 (N975, N958, N409);
xor XOR2 (N976, N966, N696);
buf BUF1 (N977, N969);
not NOT1 (N978, N976);
or OR4 (N979, N947, N685, N218, N122);
and AND4 (N980, N973, N411, N770, N809);
xor XOR2 (N981, N978, N97);
buf BUF1 (N982, N979);
nand NAND3 (N983, N981, N378, N900);
nor NOR3 (N984, N977, N597, N757);
nand NAND3 (N985, N974, N794, N842);
nor NOR2 (N986, N975, N158);
or OR2 (N987, N984, N175);
nor NOR3 (N988, N987, N885, N116);
xor XOR2 (N989, N985, N795);
not NOT1 (N990, N983);
or OR2 (N991, N989, N839);
not NOT1 (N992, N982);
xor XOR2 (N993, N942, N510);
nor NOR4 (N994, N991, N836, N514, N355);
and AND2 (N995, N994, N138);
xor XOR2 (N996, N990, N591);
nand NAND2 (N997, N988, N509);
not NOT1 (N998, N970);
buf BUF1 (N999, N993);
nand NAND2 (N1000, N998, N201);
or OR2 (N1001, N995, N429);
not NOT1 (N1002, N964);
xor XOR2 (N1003, N1001, N968);
buf BUF1 (N1004, N986);
not NOT1 (N1005, N1000);
xor XOR2 (N1006, N1004, N672);
or OR2 (N1007, N1003, N909);
nand NAND4 (N1008, N1007, N191, N364, N65);
nand NAND2 (N1009, N972, N837);
nand NAND3 (N1010, N992, N300, N366);
nor NOR3 (N1011, N999, N631, N931);
xor XOR2 (N1012, N996, N827);
not NOT1 (N1013, N997);
not NOT1 (N1014, N1002);
nor NOR3 (N1015, N1008, N567, N22);
or OR4 (N1016, N1011, N318, N524, N723);
nand NAND3 (N1017, N1005, N147, N972);
nand NAND4 (N1018, N1016, N330, N485, N124);
nor NOR4 (N1019, N1012, N82, N309, N248);
and AND4 (N1020, N1014, N906, N320, N515);
nand NAND2 (N1021, N1013, N317);
and AND2 (N1022, N1015, N873);
nor NOR3 (N1023, N1010, N1004, N40);
and AND4 (N1024, N1009, N170, N97, N134);
not NOT1 (N1025, N1022);
nor NOR2 (N1026, N1019, N873);
and AND2 (N1027, N1024, N537);
nand NAND3 (N1028, N1018, N932, N62);
buf BUF1 (N1029, N1021);
or OR2 (N1030, N1017, N482);
or OR2 (N1031, N1027, N913);
not NOT1 (N1032, N1028);
and AND3 (N1033, N1006, N728, N294);
and AND3 (N1034, N1032, N29, N236);
buf BUF1 (N1035, N1026);
xor XOR2 (N1036, N1029, N587);
not NOT1 (N1037, N1030);
buf BUF1 (N1038, N1025);
not NOT1 (N1039, N980);
xor XOR2 (N1040, N1033, N200);
xor XOR2 (N1041, N1036, N260);
and AND2 (N1042, N1023, N674);
not NOT1 (N1043, N1038);
nand NAND3 (N1044, N1039, N490, N541);
not NOT1 (N1045, N1044);
xor XOR2 (N1046, N1045, N106);
nand NAND3 (N1047, N1042, N921, N440);
or OR2 (N1048, N1043, N914);
buf BUF1 (N1049, N1037);
or OR2 (N1050, N1041, N605);
nor NOR4 (N1051, N1035, N177, N761, N697);
nor NOR2 (N1052, N1046, N400);
or OR4 (N1053, N1052, N525, N131, N670);
nand NAND2 (N1054, N1049, N21);
xor XOR2 (N1055, N1034, N88);
buf BUF1 (N1056, N1053);
xor XOR2 (N1057, N1050, N710);
and AND4 (N1058, N1047, N656, N957, N214);
or OR3 (N1059, N1048, N213, N35);
buf BUF1 (N1060, N1020);
nand NAND4 (N1061, N1060, N164, N554, N586);
or OR2 (N1062, N1061, N812);
nor NOR2 (N1063, N1062, N804);
and AND4 (N1064, N1054, N286, N426, N417);
and AND2 (N1065, N1056, N82);
xor XOR2 (N1066, N1051, N30);
or OR4 (N1067, N1064, N43, N289, N1047);
not NOT1 (N1068, N1063);
nand NAND2 (N1069, N1031, N642);
nand NAND3 (N1070, N1059, N723, N548);
and AND3 (N1071, N1069, N416, N1048);
buf BUF1 (N1072, N1070);
nor NOR4 (N1073, N1067, N397, N852, N512);
nand NAND3 (N1074, N1058, N588, N147);
or OR4 (N1075, N1071, N608, N976, N1040);
nand NAND4 (N1076, N120, N695, N334, N377);
not NOT1 (N1077, N1066);
not NOT1 (N1078, N1076);
or OR4 (N1079, N1055, N902, N957, N863);
not NOT1 (N1080, N1078);
not NOT1 (N1081, N1080);
buf BUF1 (N1082, N1073);
and AND4 (N1083, N1072, N301, N273, N708);
nand NAND3 (N1084, N1081, N860, N719);
buf BUF1 (N1085, N1065);
buf BUF1 (N1086, N1083);
xor XOR2 (N1087, N1086, N408);
and AND2 (N1088, N1082, N161);
or OR4 (N1089, N1057, N923, N168, N162);
not NOT1 (N1090, N1085);
nand NAND3 (N1091, N1089, N187, N390);
xor XOR2 (N1092, N1088, N661);
not NOT1 (N1093, N1074);
xor XOR2 (N1094, N1092, N290);
and AND2 (N1095, N1084, N221);
or OR2 (N1096, N1093, N436);
buf BUF1 (N1097, N1075);
buf BUF1 (N1098, N1087);
nand NAND4 (N1099, N1079, N408, N958, N816);
nor NOR4 (N1100, N1098, N10, N324, N950);
xor XOR2 (N1101, N1090, N823);
buf BUF1 (N1102, N1096);
xor XOR2 (N1103, N1091, N488);
or OR2 (N1104, N1101, N268);
xor XOR2 (N1105, N1094, N343);
buf BUF1 (N1106, N1099);
nand NAND4 (N1107, N1068, N646, N72, N720);
or OR3 (N1108, N1107, N532, N1038);
nand NAND2 (N1109, N1103, N705);
nand NAND4 (N1110, N1106, N791, N509, N194);
nor NOR4 (N1111, N1108, N38, N597, N40);
or OR4 (N1112, N1104, N276, N1060, N588);
nor NOR2 (N1113, N1097, N838);
and AND4 (N1114, N1100, N1076, N784, N500);
or OR3 (N1115, N1111, N658, N516);
xor XOR2 (N1116, N1077, N264);
or OR4 (N1117, N1114, N811, N211, N570);
nor NOR3 (N1118, N1110, N184, N373);
nor NOR3 (N1119, N1112, N42, N646);
buf BUF1 (N1120, N1109);
buf BUF1 (N1121, N1120);
buf BUF1 (N1122, N1119);
nand NAND4 (N1123, N1102, N48, N151, N45);
not NOT1 (N1124, N1121);
buf BUF1 (N1125, N1124);
nand NAND2 (N1126, N1105, N281);
nand NAND4 (N1127, N1126, N644, N86, N935);
not NOT1 (N1128, N1125);
and AND2 (N1129, N1127, N764);
xor XOR2 (N1130, N1116, N244);
or OR3 (N1131, N1118, N690, N175);
or OR4 (N1132, N1128, N148, N273, N902);
nor NOR4 (N1133, N1117, N784, N133, N1123);
buf BUF1 (N1134, N673);
buf BUF1 (N1135, N1115);
not NOT1 (N1136, N1122);
xor XOR2 (N1137, N1130, N859);
and AND3 (N1138, N1095, N602, N1102);
nand NAND2 (N1139, N1129, N107);
not NOT1 (N1140, N1136);
not NOT1 (N1141, N1137);
or OR2 (N1142, N1141, N1109);
nand NAND4 (N1143, N1142, N29, N839, N735);
nand NAND3 (N1144, N1138, N583, N714);
not NOT1 (N1145, N1139);
not NOT1 (N1146, N1135);
or OR2 (N1147, N1140, N561);
not NOT1 (N1148, N1144);
nand NAND2 (N1149, N1146, N904);
nand NAND4 (N1150, N1133, N130, N15, N469);
and AND3 (N1151, N1132, N282, N634);
and AND3 (N1152, N1150, N411, N186);
and AND3 (N1153, N1148, N380, N428);
nand NAND4 (N1154, N1113, N166, N917, N964);
not NOT1 (N1155, N1143);
nand NAND2 (N1156, N1131, N542);
xor XOR2 (N1157, N1156, N744);
buf BUF1 (N1158, N1157);
and AND2 (N1159, N1145, N650);
or OR2 (N1160, N1153, N190);
not NOT1 (N1161, N1155);
and AND2 (N1162, N1147, N875);
buf BUF1 (N1163, N1160);
nand NAND4 (N1164, N1134, N529, N177, N723);
or OR4 (N1165, N1154, N847, N791, N165);
nor NOR2 (N1166, N1149, N333);
nor NOR4 (N1167, N1162, N920, N618, N82);
buf BUF1 (N1168, N1151);
buf BUF1 (N1169, N1165);
not NOT1 (N1170, N1167);
and AND4 (N1171, N1166, N257, N902, N338);
not NOT1 (N1172, N1152);
and AND4 (N1173, N1159, N964, N541, N375);
and AND3 (N1174, N1161, N438, N382);
buf BUF1 (N1175, N1168);
nand NAND4 (N1176, N1173, N982, N837, N622);
buf BUF1 (N1177, N1163);
nor NOR2 (N1178, N1170, N1083);
nand NAND4 (N1179, N1177, N32, N433, N334);
not NOT1 (N1180, N1179);
nand NAND2 (N1181, N1169, N132);
not NOT1 (N1182, N1164);
and AND4 (N1183, N1158, N204, N109, N558);
xor XOR2 (N1184, N1180, N470);
or OR4 (N1185, N1174, N798, N643, N679);
buf BUF1 (N1186, N1175);
buf BUF1 (N1187, N1171);
xor XOR2 (N1188, N1176, N422);
buf BUF1 (N1189, N1178);
nand NAND4 (N1190, N1181, N503, N496, N1083);
nor NOR3 (N1191, N1185, N1006, N1025);
buf BUF1 (N1192, N1190);
or OR4 (N1193, N1187, N184, N333, N761);
buf BUF1 (N1194, N1189);
or OR3 (N1195, N1184, N1096, N1139);
or OR4 (N1196, N1182, N938, N925, N886);
xor XOR2 (N1197, N1172, N988);
not NOT1 (N1198, N1183);
xor XOR2 (N1199, N1198, N5);
xor XOR2 (N1200, N1197, N681);
or OR3 (N1201, N1192, N202, N1169);
and AND3 (N1202, N1199, N62, N175);
xor XOR2 (N1203, N1200, N80);
or OR4 (N1204, N1201, N433, N838, N26);
buf BUF1 (N1205, N1195);
xor XOR2 (N1206, N1193, N220);
not NOT1 (N1207, N1205);
xor XOR2 (N1208, N1207, N1018);
or OR2 (N1209, N1208, N619);
nor NOR2 (N1210, N1209, N68);
nand NAND4 (N1211, N1186, N664, N1169, N808);
buf BUF1 (N1212, N1191);
xor XOR2 (N1213, N1203, N645);
buf BUF1 (N1214, N1210);
or OR3 (N1215, N1212, N454, N779);
and AND2 (N1216, N1213, N836);
xor XOR2 (N1217, N1204, N551);
nor NOR2 (N1218, N1217, N485);
buf BUF1 (N1219, N1214);
or OR4 (N1220, N1188, N576, N49, N558);
xor XOR2 (N1221, N1211, N1094);
not NOT1 (N1222, N1194);
and AND2 (N1223, N1220, N83);
or OR3 (N1224, N1196, N955, N801);
or OR4 (N1225, N1216, N990, N55, N735);
nor NOR3 (N1226, N1225, N985, N288);
or OR3 (N1227, N1218, N1208, N1073);
and AND2 (N1228, N1224, N425);
nand NAND3 (N1229, N1202, N1106, N902);
and AND3 (N1230, N1215, N635, N187);
and AND4 (N1231, N1229, N438, N867, N927);
not NOT1 (N1232, N1231);
nand NAND2 (N1233, N1221, N30);
buf BUF1 (N1234, N1227);
and AND3 (N1235, N1234, N610, N189);
xor XOR2 (N1236, N1235, N322);
nand NAND2 (N1237, N1230, N84);
nand NAND4 (N1238, N1226, N1107, N678, N399);
nand NAND3 (N1239, N1238, N1096, N867);
and AND3 (N1240, N1237, N772, N973);
buf BUF1 (N1241, N1232);
or OR3 (N1242, N1206, N583, N740);
nor NOR4 (N1243, N1233, N557, N730, N654);
or OR4 (N1244, N1239, N963, N354, N1121);
nand NAND2 (N1245, N1240, N628);
nand NAND2 (N1246, N1243, N374);
and AND3 (N1247, N1236, N195, N1120);
nand NAND4 (N1248, N1245, N733, N622, N1067);
and AND3 (N1249, N1242, N68, N84);
buf BUF1 (N1250, N1248);
not NOT1 (N1251, N1250);
xor XOR2 (N1252, N1222, N860);
or OR4 (N1253, N1251, N1238, N679, N1059);
not NOT1 (N1254, N1246);
nor NOR2 (N1255, N1249, N284);
nand NAND4 (N1256, N1244, N891, N374, N1149);
nand NAND3 (N1257, N1219, N159, N338);
nor NOR3 (N1258, N1228, N575, N866);
nand NAND3 (N1259, N1254, N199, N436);
not NOT1 (N1260, N1256);
nor NOR4 (N1261, N1241, N453, N1178, N1028);
buf BUF1 (N1262, N1258);
buf BUF1 (N1263, N1259);
or OR4 (N1264, N1262, N936, N994, N159);
nor NOR4 (N1265, N1257, N729, N996, N198);
buf BUF1 (N1266, N1261);
nand NAND4 (N1267, N1247, N709, N1003, N1095);
or OR2 (N1268, N1263, N1008);
xor XOR2 (N1269, N1265, N1019);
or OR4 (N1270, N1268, N500, N1247, N121);
or OR2 (N1271, N1269, N322);
nor NOR3 (N1272, N1255, N67, N176);
buf BUF1 (N1273, N1270);
xor XOR2 (N1274, N1266, N760);
xor XOR2 (N1275, N1252, N232);
or OR4 (N1276, N1264, N1096, N1103, N544);
or OR4 (N1277, N1267, N1244, N304, N1077);
buf BUF1 (N1278, N1271);
nor NOR3 (N1279, N1273, N935, N498);
nand NAND3 (N1280, N1277, N1236, N984);
or OR3 (N1281, N1272, N501, N482);
buf BUF1 (N1282, N1274);
not NOT1 (N1283, N1223);
and AND2 (N1284, N1260, N879);
xor XOR2 (N1285, N1281, N1089);
xor XOR2 (N1286, N1279, N430);
nand NAND3 (N1287, N1282, N770, N651);
and AND4 (N1288, N1276, N543, N897, N143);
nor NOR2 (N1289, N1288, N542);
or OR3 (N1290, N1286, N129, N1051);
not NOT1 (N1291, N1290);
nand NAND3 (N1292, N1285, N326, N46);
not NOT1 (N1293, N1284);
nor NOR3 (N1294, N1280, N1198, N756);
nand NAND3 (N1295, N1278, N426, N278);
nor NOR2 (N1296, N1289, N42);
nor NOR3 (N1297, N1287, N186, N344);
or OR4 (N1298, N1291, N837, N312, N1059);
xor XOR2 (N1299, N1298, N173);
or OR4 (N1300, N1293, N150, N619, N180);
nand NAND4 (N1301, N1292, N795, N330, N767);
nand NAND3 (N1302, N1299, N987, N710);
or OR2 (N1303, N1253, N548);
xor XOR2 (N1304, N1283, N422);
not NOT1 (N1305, N1303);
not NOT1 (N1306, N1295);
nand NAND2 (N1307, N1304, N293);
or OR3 (N1308, N1296, N71, N1199);
buf BUF1 (N1309, N1275);
xor XOR2 (N1310, N1294, N1024);
nand NAND4 (N1311, N1300, N287, N1010, N364);
buf BUF1 (N1312, N1301);
buf BUF1 (N1313, N1307);
nand NAND4 (N1314, N1308, N75, N905, N346);
or OR2 (N1315, N1302, N436);
or OR2 (N1316, N1314, N377);
not NOT1 (N1317, N1297);
and AND3 (N1318, N1305, N540, N509);
xor XOR2 (N1319, N1317, N315);
nor NOR4 (N1320, N1316, N196, N650, N543);
nand NAND2 (N1321, N1315, N43);
not NOT1 (N1322, N1319);
xor XOR2 (N1323, N1322, N1293);
nor NOR2 (N1324, N1310, N657);
not NOT1 (N1325, N1321);
buf BUF1 (N1326, N1313);
or OR4 (N1327, N1306, N860, N632, N1303);
not NOT1 (N1328, N1312);
and AND2 (N1329, N1325, N309);
xor XOR2 (N1330, N1318, N333);
and AND2 (N1331, N1326, N916);
nor NOR3 (N1332, N1309, N203, N212);
and AND3 (N1333, N1324, N946, N797);
nor NOR4 (N1334, N1328, N904, N549, N1010);
or OR2 (N1335, N1320, N612);
xor XOR2 (N1336, N1323, N38);
not NOT1 (N1337, N1331);
and AND3 (N1338, N1335, N776, N1064);
not NOT1 (N1339, N1311);
nand NAND4 (N1340, N1327, N1250, N253, N1037);
or OR4 (N1341, N1336, N456, N203, N73);
and AND4 (N1342, N1338, N315, N559, N1149);
nor NOR2 (N1343, N1339, N516);
not NOT1 (N1344, N1341);
not NOT1 (N1345, N1332);
not NOT1 (N1346, N1330);
buf BUF1 (N1347, N1334);
nand NAND3 (N1348, N1329, N870, N1116);
xor XOR2 (N1349, N1340, N752);
or OR2 (N1350, N1345, N1020);
not NOT1 (N1351, N1350);
buf BUF1 (N1352, N1337);
xor XOR2 (N1353, N1333, N547);
xor XOR2 (N1354, N1348, N229);
buf BUF1 (N1355, N1354);
nor NOR3 (N1356, N1342, N13, N396);
nor NOR3 (N1357, N1352, N1190, N1288);
nand NAND4 (N1358, N1357, N1141, N1056, N1289);
nand NAND3 (N1359, N1353, N115, N407);
nand NAND2 (N1360, N1356, N543);
not NOT1 (N1361, N1351);
and AND3 (N1362, N1358, N1002, N559);
or OR2 (N1363, N1347, N1081);
nand NAND4 (N1364, N1346, N70, N1, N696);
not NOT1 (N1365, N1361);
nor NOR2 (N1366, N1362, N1289);
nand NAND4 (N1367, N1349, N1277, N1257, N615);
or OR3 (N1368, N1360, N783, N544);
and AND4 (N1369, N1344, N513, N897, N695);
nand NAND4 (N1370, N1367, N1093, N100, N273);
or OR4 (N1371, N1370, N1357, N1370, N1090);
or OR4 (N1372, N1368, N781, N656, N962);
or OR4 (N1373, N1359, N1019, N447, N935);
nor NOR2 (N1374, N1364, N177);
not NOT1 (N1375, N1366);
nand NAND3 (N1376, N1363, N929, N575);
buf BUF1 (N1377, N1374);
not NOT1 (N1378, N1376);
buf BUF1 (N1379, N1355);
not NOT1 (N1380, N1377);
nor NOR2 (N1381, N1343, N1280);
nor NOR2 (N1382, N1378, N387);
or OR4 (N1383, N1365, N1310, N8, N1363);
or OR4 (N1384, N1371, N1126, N629, N847);
or OR4 (N1385, N1382, N639, N509, N279);
not NOT1 (N1386, N1381);
nor NOR4 (N1387, N1383, N22, N1230, N807);
or OR4 (N1388, N1379, N533, N729, N1203);
nand NAND3 (N1389, N1384, N606, N519);
buf BUF1 (N1390, N1373);
nand NAND3 (N1391, N1372, N822, N1048);
not NOT1 (N1392, N1385);
or OR2 (N1393, N1392, N539);
or OR3 (N1394, N1389, N1131, N9);
xor XOR2 (N1395, N1386, N1218);
nor NOR2 (N1396, N1395, N1036);
and AND3 (N1397, N1369, N1141, N42);
not NOT1 (N1398, N1394);
buf BUF1 (N1399, N1390);
and AND3 (N1400, N1387, N210, N614);
nor NOR3 (N1401, N1393, N446, N882);
not NOT1 (N1402, N1396);
nor NOR3 (N1403, N1402, N520, N674);
or OR2 (N1404, N1380, N372);
nor NOR3 (N1405, N1391, N479, N1157);
and AND3 (N1406, N1375, N232, N181);
xor XOR2 (N1407, N1403, N1111);
xor XOR2 (N1408, N1406, N246);
not NOT1 (N1409, N1401);
not NOT1 (N1410, N1408);
or OR2 (N1411, N1399, N640);
nor NOR4 (N1412, N1410, N1281, N481, N474);
and AND2 (N1413, N1411, N863);
xor XOR2 (N1414, N1412, N69);
or OR2 (N1415, N1400, N219);
nand NAND2 (N1416, N1407, N253);
nand NAND3 (N1417, N1405, N1215, N617);
not NOT1 (N1418, N1416);
nor NOR2 (N1419, N1417, N704);
and AND3 (N1420, N1409, N885, N1270);
xor XOR2 (N1421, N1418, N546);
xor XOR2 (N1422, N1397, N1002);
or OR4 (N1423, N1404, N652, N1359, N285);
nor NOR4 (N1424, N1423, N124, N607, N864);
not NOT1 (N1425, N1398);
and AND4 (N1426, N1421, N80, N225, N1003);
buf BUF1 (N1427, N1420);
not NOT1 (N1428, N1422);
and AND4 (N1429, N1413, N1335, N1065, N899);
xor XOR2 (N1430, N1419, N1336);
or OR2 (N1431, N1428, N995);
nor NOR3 (N1432, N1388, N935, N9);
buf BUF1 (N1433, N1425);
nor NOR2 (N1434, N1433, N443);
not NOT1 (N1435, N1424);
nor NOR4 (N1436, N1429, N1037, N644, N634);
nor NOR3 (N1437, N1426, N323, N433);
not NOT1 (N1438, N1432);
buf BUF1 (N1439, N1430);
xor XOR2 (N1440, N1427, N309);
xor XOR2 (N1441, N1436, N339);
nand NAND4 (N1442, N1441, N871, N499, N765);
not NOT1 (N1443, N1437);
nor NOR3 (N1444, N1414, N948, N443);
nor NOR3 (N1445, N1444, N1080, N1309);
nor NOR4 (N1446, N1415, N840, N159, N411);
not NOT1 (N1447, N1445);
nand NAND2 (N1448, N1434, N1284);
or OR2 (N1449, N1431, N905);
not NOT1 (N1450, N1449);
nor NOR4 (N1451, N1439, N465, N782, N945);
or OR3 (N1452, N1446, N677, N425);
or OR3 (N1453, N1443, N221, N45);
nor NOR3 (N1454, N1451, N775, N196);
and AND2 (N1455, N1454, N1327);
buf BUF1 (N1456, N1442);
nor NOR3 (N1457, N1453, N545, N496);
nand NAND3 (N1458, N1438, N1206, N1158);
xor XOR2 (N1459, N1440, N464);
and AND4 (N1460, N1455, N1162, N844, N1457);
not NOT1 (N1461, N656);
not NOT1 (N1462, N1435);
buf BUF1 (N1463, N1456);
nor NOR3 (N1464, N1462, N1039, N536);
xor XOR2 (N1465, N1463, N223);
xor XOR2 (N1466, N1450, N1111);
nor NOR4 (N1467, N1459, N933, N1346, N349);
buf BUF1 (N1468, N1466);
xor XOR2 (N1469, N1447, N380);
nand NAND4 (N1470, N1469, N212, N665, N382);
buf BUF1 (N1471, N1464);
nand NAND4 (N1472, N1452, N1118, N404, N244);
not NOT1 (N1473, N1461);
not NOT1 (N1474, N1467);
or OR2 (N1475, N1468, N786);
nor NOR2 (N1476, N1470, N1176);
buf BUF1 (N1477, N1476);
nand NAND2 (N1478, N1471, N1449);
buf BUF1 (N1479, N1473);
not NOT1 (N1480, N1472);
or OR4 (N1481, N1480, N448, N135, N405);
buf BUF1 (N1482, N1478);
nor NOR3 (N1483, N1474, N1188, N918);
buf BUF1 (N1484, N1479);
nand NAND2 (N1485, N1482, N371);
nor NOR4 (N1486, N1485, N559, N1410, N1125);
buf BUF1 (N1487, N1477);
and AND4 (N1488, N1448, N366, N986, N1480);
nand NAND2 (N1489, N1458, N366);
nor NOR2 (N1490, N1465, N1287);
buf BUF1 (N1491, N1487);
nor NOR3 (N1492, N1460, N1049, N963);
or OR2 (N1493, N1490, N828);
nor NOR2 (N1494, N1489, N654);
and AND3 (N1495, N1484, N46, N233);
nor NOR4 (N1496, N1494, N109, N1258, N1104);
not NOT1 (N1497, N1491);
nor NOR2 (N1498, N1486, N1462);
not NOT1 (N1499, N1495);
not NOT1 (N1500, N1498);
nand NAND4 (N1501, N1492, N630, N1259, N115);
buf BUF1 (N1502, N1488);
or OR2 (N1503, N1481, N459);
buf BUF1 (N1504, N1500);
and AND3 (N1505, N1475, N601, N877);
buf BUF1 (N1506, N1504);
or OR3 (N1507, N1503, N1154, N328);
nand NAND4 (N1508, N1502, N944, N1468, N213);
and AND4 (N1509, N1496, N947, N1328, N1484);
and AND2 (N1510, N1501, N282);
nor NOR4 (N1511, N1505, N598, N76, N169);
buf BUF1 (N1512, N1508);
xor XOR2 (N1513, N1483, N529);
or OR3 (N1514, N1497, N1121, N130);
not NOT1 (N1515, N1510);
nand NAND3 (N1516, N1507, N299, N397);
or OR3 (N1517, N1493, N1037, N979);
buf BUF1 (N1518, N1516);
nor NOR3 (N1519, N1513, N817, N981);
xor XOR2 (N1520, N1499, N768);
nor NOR4 (N1521, N1519, N818, N891, N584);
not NOT1 (N1522, N1512);
nor NOR4 (N1523, N1506, N1477, N1170, N999);
buf BUF1 (N1524, N1518);
nor NOR3 (N1525, N1524, N808, N1499);
or OR2 (N1526, N1521, N300);
not NOT1 (N1527, N1523);
not NOT1 (N1528, N1511);
nand NAND2 (N1529, N1520, N236);
and AND3 (N1530, N1514, N572, N1043);
nand NAND4 (N1531, N1525, N1051, N1093, N609);
or OR2 (N1532, N1526, N918);
xor XOR2 (N1533, N1527, N266);
buf BUF1 (N1534, N1515);
xor XOR2 (N1535, N1532, N129);
nor NOR2 (N1536, N1533, N302);
and AND3 (N1537, N1529, N540, N595);
xor XOR2 (N1538, N1522, N1388);
or OR2 (N1539, N1530, N602);
not NOT1 (N1540, N1509);
nand NAND2 (N1541, N1536, N1391);
and AND3 (N1542, N1534, N425, N967);
not NOT1 (N1543, N1517);
not NOT1 (N1544, N1540);
and AND3 (N1545, N1541, N1354, N579);
and AND4 (N1546, N1535, N820, N609, N854);
and AND4 (N1547, N1531, N108, N432, N335);
nand NAND4 (N1548, N1538, N277, N785, N1420);
not NOT1 (N1549, N1545);
buf BUF1 (N1550, N1547);
xor XOR2 (N1551, N1544, N1349);
not NOT1 (N1552, N1549);
buf BUF1 (N1553, N1546);
nand NAND4 (N1554, N1543, N1455, N1172, N658);
nand NAND3 (N1555, N1552, N595, N628);
buf BUF1 (N1556, N1542);
buf BUF1 (N1557, N1556);
buf BUF1 (N1558, N1555);
or OR3 (N1559, N1554, N636, N179);
nor NOR4 (N1560, N1553, N554, N1260, N418);
and AND4 (N1561, N1548, N1554, N1424, N741);
and AND4 (N1562, N1528, N63, N334, N1019);
and AND2 (N1563, N1557, N294);
xor XOR2 (N1564, N1562, N58);
not NOT1 (N1565, N1550);
not NOT1 (N1566, N1558);
nor NOR4 (N1567, N1564, N515, N379, N1432);
buf BUF1 (N1568, N1566);
buf BUF1 (N1569, N1537);
nand NAND2 (N1570, N1569, N1211);
or OR4 (N1571, N1551, N580, N702, N183);
and AND3 (N1572, N1565, N1564, N1116);
nand NAND2 (N1573, N1560, N1563);
buf BUF1 (N1574, N194);
and AND2 (N1575, N1561, N645);
not NOT1 (N1576, N1573);
nand NAND2 (N1577, N1567, N1556);
nand NAND2 (N1578, N1577, N882);
not NOT1 (N1579, N1578);
not NOT1 (N1580, N1568);
buf BUF1 (N1581, N1576);
nor NOR2 (N1582, N1580, N745);
nand NAND2 (N1583, N1571, N184);
and AND2 (N1584, N1572, N1439);
or OR4 (N1585, N1583, N666, N554, N82);
and AND3 (N1586, N1539, N49, N1160);
xor XOR2 (N1587, N1579, N39);
buf BUF1 (N1588, N1581);
xor XOR2 (N1589, N1570, N288);
or OR4 (N1590, N1588, N262, N1292, N1527);
and AND4 (N1591, N1585, N505, N545, N69);
nor NOR2 (N1592, N1587, N1228);
nor NOR2 (N1593, N1584, N313);
and AND4 (N1594, N1590, N511, N372, N977);
buf BUF1 (N1595, N1592);
nand NAND2 (N1596, N1575, N135);
buf BUF1 (N1597, N1589);
xor XOR2 (N1598, N1596, N99);
not NOT1 (N1599, N1559);
xor XOR2 (N1600, N1591, N260);
or OR3 (N1601, N1593, N450, N1401);
buf BUF1 (N1602, N1601);
xor XOR2 (N1603, N1595, N812);
xor XOR2 (N1604, N1574, N1177);
nor NOR3 (N1605, N1582, N693, N709);
or OR2 (N1606, N1594, N1553);
nand NAND2 (N1607, N1599, N834);
not NOT1 (N1608, N1604);
nor NOR3 (N1609, N1606, N472, N1547);
nor NOR3 (N1610, N1609, N810, N510);
nor NOR4 (N1611, N1605, N262, N1365, N1436);
or OR2 (N1612, N1600, N953);
or OR4 (N1613, N1612, N570, N253, N97);
or OR2 (N1614, N1603, N1248);
or OR4 (N1615, N1607, N189, N55, N496);
nor NOR4 (N1616, N1608, N872, N34, N1599);
nand NAND2 (N1617, N1602, N1211);
xor XOR2 (N1618, N1613, N1243);
nand NAND3 (N1619, N1611, N351, N1226);
nand NAND2 (N1620, N1618, N1320);
xor XOR2 (N1621, N1620, N952);
and AND3 (N1622, N1598, N1256, N188);
xor XOR2 (N1623, N1619, N637);
nand NAND3 (N1624, N1615, N798, N680);
nand NAND3 (N1625, N1614, N1365, N1497);
or OR3 (N1626, N1624, N1366, N499);
or OR4 (N1627, N1621, N834, N190, N212);
not NOT1 (N1628, N1617);
and AND3 (N1629, N1628, N725, N1382);
nand NAND2 (N1630, N1626, N803);
and AND3 (N1631, N1630, N357, N70);
or OR3 (N1632, N1627, N1413, N371);
not NOT1 (N1633, N1629);
not NOT1 (N1634, N1610);
nor NOR3 (N1635, N1633, N1555, N1612);
not NOT1 (N1636, N1634);
or OR4 (N1637, N1623, N1062, N302, N128);
or OR2 (N1638, N1631, N60);
buf BUF1 (N1639, N1597);
nor NOR3 (N1640, N1586, N1155, N1167);
nor NOR4 (N1641, N1636, N579, N783, N406);
and AND4 (N1642, N1639, N1084, N1569, N1453);
buf BUF1 (N1643, N1635);
and AND4 (N1644, N1622, N1425, N287, N432);
xor XOR2 (N1645, N1644, N825);
nand NAND3 (N1646, N1645, N1487, N524);
nor NOR3 (N1647, N1640, N644, N635);
nor NOR2 (N1648, N1642, N895);
nor NOR4 (N1649, N1632, N24, N310, N95);
nand NAND3 (N1650, N1638, N695, N812);
or OR2 (N1651, N1648, N112);
not NOT1 (N1652, N1650);
nand NAND2 (N1653, N1625, N883);
nand NAND3 (N1654, N1651, N159, N1635);
nand NAND4 (N1655, N1637, N1376, N1307, N1050);
and AND3 (N1656, N1653, N68, N164);
not NOT1 (N1657, N1656);
and AND4 (N1658, N1646, N193, N821, N913);
nand NAND2 (N1659, N1641, N307);
nand NAND2 (N1660, N1643, N1635);
or OR4 (N1661, N1616, N308, N1559, N597);
and AND4 (N1662, N1655, N1054, N1378, N1421);
and AND2 (N1663, N1658, N753);
buf BUF1 (N1664, N1663);
nor NOR4 (N1665, N1657, N732, N1438, N66);
nand NAND3 (N1666, N1652, N1490, N1600);
xor XOR2 (N1667, N1647, N572);
xor XOR2 (N1668, N1649, N648);
nand NAND3 (N1669, N1654, N1378, N330);
and AND3 (N1670, N1664, N480, N524);
and AND3 (N1671, N1665, N1416, N1116);
buf BUF1 (N1672, N1670);
xor XOR2 (N1673, N1668, N497);
nand NAND2 (N1674, N1661, N1249);
and AND4 (N1675, N1659, N506, N573, N813);
nand NAND4 (N1676, N1667, N829, N1446, N354);
or OR2 (N1677, N1672, N593);
nand NAND3 (N1678, N1674, N919, N338);
or OR4 (N1679, N1662, N672, N584, N307);
xor XOR2 (N1680, N1673, N1401);
not NOT1 (N1681, N1660);
nor NOR3 (N1682, N1666, N351, N728);
buf BUF1 (N1683, N1682);
buf BUF1 (N1684, N1681);
or OR3 (N1685, N1680, N1127, N1613);
not NOT1 (N1686, N1683);
or OR3 (N1687, N1671, N1158, N400);
xor XOR2 (N1688, N1677, N571);
buf BUF1 (N1689, N1675);
nor NOR2 (N1690, N1684, N1496);
nand NAND2 (N1691, N1687, N99);
or OR3 (N1692, N1690, N698, N1091);
buf BUF1 (N1693, N1679);
buf BUF1 (N1694, N1676);
not NOT1 (N1695, N1678);
nand NAND3 (N1696, N1669, N694, N1142);
not NOT1 (N1697, N1686);
not NOT1 (N1698, N1694);
not NOT1 (N1699, N1697);
not NOT1 (N1700, N1698);
nor NOR4 (N1701, N1699, N1478, N1214, N928);
nor NOR2 (N1702, N1701, N232);
not NOT1 (N1703, N1692);
and AND4 (N1704, N1688, N679, N691, N508);
nor NOR4 (N1705, N1702, N427, N788, N1002);
buf BUF1 (N1706, N1693);
not NOT1 (N1707, N1685);
buf BUF1 (N1708, N1689);
and AND2 (N1709, N1696, N767);
not NOT1 (N1710, N1700);
nand NAND3 (N1711, N1705, N1179, N483);
and AND4 (N1712, N1708, N966, N1064, N1290);
nor NOR4 (N1713, N1695, N440, N1238, N1176);
nor NOR3 (N1714, N1691, N149, N165);
nor NOR2 (N1715, N1712, N972);
not NOT1 (N1716, N1709);
and AND4 (N1717, N1711, N748, N475, N792);
nor NOR2 (N1718, N1706, N1479);
nor NOR3 (N1719, N1714, N959, N340);
nor NOR4 (N1720, N1703, N550, N579, N1292);
xor XOR2 (N1721, N1719, N1023);
not NOT1 (N1722, N1704);
xor XOR2 (N1723, N1718, N1180);
or OR2 (N1724, N1710, N741);
xor XOR2 (N1725, N1720, N1350);
not NOT1 (N1726, N1717);
xor XOR2 (N1727, N1726, N1203);
buf BUF1 (N1728, N1725);
buf BUF1 (N1729, N1713);
buf BUF1 (N1730, N1727);
and AND2 (N1731, N1730, N334);
nand NAND2 (N1732, N1724, N497);
nand NAND3 (N1733, N1728, N1326, N130);
not NOT1 (N1734, N1731);
not NOT1 (N1735, N1733);
nand NAND4 (N1736, N1707, N713, N339, N1373);
buf BUF1 (N1737, N1721);
nor NOR2 (N1738, N1722, N1571);
and AND4 (N1739, N1729, N600, N997, N84);
buf BUF1 (N1740, N1736);
and AND3 (N1741, N1734, N369, N1188);
and AND3 (N1742, N1740, N1551, N114);
nor NOR4 (N1743, N1737, N1295, N656, N459);
nor NOR2 (N1744, N1715, N412);
xor XOR2 (N1745, N1735, N583);
and AND2 (N1746, N1745, N865);
xor XOR2 (N1747, N1716, N1003);
and AND4 (N1748, N1732, N380, N1557, N1348);
nand NAND2 (N1749, N1748, N1084);
nor NOR3 (N1750, N1749, N80, N576);
buf BUF1 (N1751, N1743);
nand NAND3 (N1752, N1738, N1121, N910);
and AND2 (N1753, N1739, N740);
nor NOR2 (N1754, N1753, N876);
and AND4 (N1755, N1754, N993, N1521, N1103);
not NOT1 (N1756, N1747);
and AND4 (N1757, N1744, N430, N325, N853);
or OR2 (N1758, N1723, N603);
nor NOR2 (N1759, N1741, N1502);
nand NAND2 (N1760, N1742, N1122);
or OR3 (N1761, N1759, N1086, N1720);
buf BUF1 (N1762, N1751);
and AND2 (N1763, N1750, N495);
xor XOR2 (N1764, N1762, N1647);
and AND2 (N1765, N1760, N407);
not NOT1 (N1766, N1757);
and AND2 (N1767, N1758, N1150);
xor XOR2 (N1768, N1746, N1577);
xor XOR2 (N1769, N1766, N481);
nand NAND4 (N1770, N1755, N278, N1632, N349);
not NOT1 (N1771, N1763);
nor NOR4 (N1772, N1752, N704, N1140, N318);
xor XOR2 (N1773, N1761, N996);
or OR2 (N1774, N1773, N781);
nor NOR2 (N1775, N1772, N359);
xor XOR2 (N1776, N1771, N1632);
nand NAND3 (N1777, N1774, N1222, N931);
nand NAND4 (N1778, N1769, N1097, N746, N1295);
not NOT1 (N1779, N1764);
nor NOR4 (N1780, N1767, N626, N146, N455);
or OR4 (N1781, N1770, N1103, N1738, N211);
not NOT1 (N1782, N1768);
and AND2 (N1783, N1781, N1105);
buf BUF1 (N1784, N1776);
or OR4 (N1785, N1780, N448, N19, N1538);
buf BUF1 (N1786, N1765);
or OR2 (N1787, N1756, N1277);
xor XOR2 (N1788, N1779, N1046);
nand NAND4 (N1789, N1786, N444, N741, N1010);
not NOT1 (N1790, N1788);
nor NOR4 (N1791, N1784, N1556, N611, N1240);
not NOT1 (N1792, N1789);
or OR2 (N1793, N1783, N158);
xor XOR2 (N1794, N1775, N1306);
or OR2 (N1795, N1777, N667);
nand NAND4 (N1796, N1792, N1332, N1372, N276);
nand NAND2 (N1797, N1782, N1112);
not NOT1 (N1798, N1797);
or OR4 (N1799, N1798, N225, N607, N578);
nor NOR3 (N1800, N1787, N875, N309);
nor NOR2 (N1801, N1790, N326);
xor XOR2 (N1802, N1801, N1052);
nor NOR3 (N1803, N1802, N1209, N1460);
nand NAND2 (N1804, N1791, N232);
xor XOR2 (N1805, N1794, N881);
xor XOR2 (N1806, N1799, N644);
xor XOR2 (N1807, N1795, N1613);
xor XOR2 (N1808, N1793, N241);
or OR2 (N1809, N1796, N370);
or OR4 (N1810, N1806, N1352, N179, N81);
nand NAND4 (N1811, N1810, N872, N522, N1377);
nand NAND2 (N1812, N1811, N627);
and AND4 (N1813, N1808, N1027, N1698, N431);
and AND4 (N1814, N1778, N263, N363, N406);
not NOT1 (N1815, N1804);
nand NAND3 (N1816, N1809, N1245, N856);
or OR3 (N1817, N1813, N673, N356);
nor NOR3 (N1818, N1807, N1055, N626);
or OR4 (N1819, N1814, N315, N164, N1704);
not NOT1 (N1820, N1812);
xor XOR2 (N1821, N1805, N573);
buf BUF1 (N1822, N1815);
buf BUF1 (N1823, N1821);
nor NOR3 (N1824, N1785, N318, N979);
buf BUF1 (N1825, N1803);
xor XOR2 (N1826, N1823, N1501);
nand NAND4 (N1827, N1816, N1505, N674, N167);
buf BUF1 (N1828, N1820);
buf BUF1 (N1829, N1824);
buf BUF1 (N1830, N1817);
or OR4 (N1831, N1827, N1074, N928, N1263);
buf BUF1 (N1832, N1819);
buf BUF1 (N1833, N1828);
and AND2 (N1834, N1830, N1186);
xor XOR2 (N1835, N1833, N580);
xor XOR2 (N1836, N1829, N1077);
not NOT1 (N1837, N1832);
nor NOR4 (N1838, N1836, N1168, N1700, N484);
nor NOR2 (N1839, N1834, N470);
nand NAND3 (N1840, N1837, N1699, N1804);
nor NOR3 (N1841, N1839, N1265, N898);
nand NAND4 (N1842, N1840, N268, N397, N149);
buf BUF1 (N1843, N1825);
buf BUF1 (N1844, N1838);
and AND4 (N1845, N1818, N55, N657, N1230);
not NOT1 (N1846, N1831);
buf BUF1 (N1847, N1845);
not NOT1 (N1848, N1826);
nor NOR3 (N1849, N1822, N191, N66);
nand NAND2 (N1850, N1842, N371);
buf BUF1 (N1851, N1841);
not NOT1 (N1852, N1851);
and AND4 (N1853, N1850, N1310, N575, N1562);
or OR4 (N1854, N1844, N390, N788, N1238);
xor XOR2 (N1855, N1853, N1496);
nor NOR4 (N1856, N1855, N253, N1848, N1190);
or OR4 (N1857, N213, N983, N1458, N1289);
not NOT1 (N1858, N1846);
nand NAND4 (N1859, N1800, N870, N145, N318);
nand NAND3 (N1860, N1843, N857, N300);
xor XOR2 (N1861, N1856, N558);
xor XOR2 (N1862, N1861, N797);
nand NAND4 (N1863, N1849, N1430, N1260, N1664);
nor NOR4 (N1864, N1854, N1358, N945, N1537);
nand NAND4 (N1865, N1852, N1497, N503, N1398);
xor XOR2 (N1866, N1858, N269);
not NOT1 (N1867, N1865);
or OR2 (N1868, N1867, N71);
and AND2 (N1869, N1864, N730);
nor NOR3 (N1870, N1862, N1508, N1144);
not NOT1 (N1871, N1868);
xor XOR2 (N1872, N1860, N1111);
nor NOR4 (N1873, N1857, N165, N708, N1499);
or OR4 (N1874, N1859, N92, N1820, N771);
nand NAND2 (N1875, N1863, N1440);
xor XOR2 (N1876, N1873, N494);
nor NOR2 (N1877, N1871, N751);
or OR2 (N1878, N1870, N475);
and AND4 (N1879, N1835, N1450, N1632, N1627);
buf BUF1 (N1880, N1866);
and AND3 (N1881, N1875, N611, N148);
buf BUF1 (N1882, N1876);
nor NOR3 (N1883, N1882, N1421, N402);
and AND4 (N1884, N1879, N1167, N121, N775);
xor XOR2 (N1885, N1877, N565);
not NOT1 (N1886, N1869);
xor XOR2 (N1887, N1874, N1724);
and AND4 (N1888, N1884, N536, N110, N479);
xor XOR2 (N1889, N1880, N920);
xor XOR2 (N1890, N1888, N982);
or OR4 (N1891, N1885, N345, N715, N123);
nor NOR3 (N1892, N1872, N1084, N1101);
buf BUF1 (N1893, N1891);
not NOT1 (N1894, N1881);
nor NOR4 (N1895, N1890, N80, N308, N1217);
not NOT1 (N1896, N1895);
nor NOR4 (N1897, N1878, N1543, N753, N969);
nor NOR2 (N1898, N1847, N1450);
nor NOR3 (N1899, N1892, N1280, N1582);
buf BUF1 (N1900, N1897);
not NOT1 (N1901, N1886);
nor NOR3 (N1902, N1899, N1076, N397);
nor NOR2 (N1903, N1889, N1646);
not NOT1 (N1904, N1887);
and AND2 (N1905, N1898, N334);
xor XOR2 (N1906, N1904, N664);
nand NAND2 (N1907, N1901, N1638);
nor NOR2 (N1908, N1900, N1694);
nand NAND4 (N1909, N1906, N404, N57, N142);
nand NAND2 (N1910, N1909, N349);
and AND3 (N1911, N1902, N1155, N1645);
not NOT1 (N1912, N1908);
not NOT1 (N1913, N1903);
nor NOR3 (N1914, N1894, N835, N1195);
nor NOR4 (N1915, N1914, N1130, N1104, N1909);
not NOT1 (N1916, N1905);
xor XOR2 (N1917, N1910, N1551);
nor NOR2 (N1918, N1907, N1563);
or OR4 (N1919, N1912, N1628, N583, N1782);
not NOT1 (N1920, N1913);
buf BUF1 (N1921, N1919);
nor NOR3 (N1922, N1883, N1752, N1062);
or OR3 (N1923, N1918, N804, N154);
xor XOR2 (N1924, N1921, N63);
nand NAND3 (N1925, N1911, N800, N1705);
and AND4 (N1926, N1923, N1001, N273, N568);
not NOT1 (N1927, N1920);
buf BUF1 (N1928, N1917);
and AND3 (N1929, N1924, N1200, N1223);
or OR4 (N1930, N1896, N1625, N590, N574);
nor NOR4 (N1931, N1916, N402, N851, N1065);
not NOT1 (N1932, N1922);
nand NAND4 (N1933, N1928, N1784, N1158, N678);
not NOT1 (N1934, N1926);
buf BUF1 (N1935, N1893);
nand NAND2 (N1936, N1930, N836);
not NOT1 (N1937, N1915);
buf BUF1 (N1938, N1927);
nand NAND2 (N1939, N1935, N1462);
nor NOR3 (N1940, N1925, N1158, N17);
xor XOR2 (N1941, N1929, N1429);
and AND2 (N1942, N1936, N150);
nor NOR2 (N1943, N1938, N1266);
not NOT1 (N1944, N1937);
and AND4 (N1945, N1934, N1309, N119, N614);
and AND4 (N1946, N1940, N893, N137, N1272);
buf BUF1 (N1947, N1931);
not NOT1 (N1948, N1932);
nor NOR3 (N1949, N1933, N696, N1699);
xor XOR2 (N1950, N1942, N1000);
not NOT1 (N1951, N1945);
xor XOR2 (N1952, N1941, N620);
nor NOR2 (N1953, N1944, N1811);
and AND4 (N1954, N1953, N1750, N1412, N1189);
not NOT1 (N1955, N1949);
nand NAND2 (N1956, N1947, N1553);
not NOT1 (N1957, N1956);
or OR4 (N1958, N1957, N491, N1683, N1475);
xor XOR2 (N1959, N1939, N1090);
and AND2 (N1960, N1954, N1079);
and AND3 (N1961, N1958, N478, N1377);
xor XOR2 (N1962, N1961, N561);
and AND2 (N1963, N1950, N1698);
nor NOR3 (N1964, N1948, N1749, N786);
nor NOR2 (N1965, N1951, N410);
nand NAND2 (N1966, N1955, N1854);
or OR4 (N1967, N1960, N1122, N1418, N64);
nor NOR3 (N1968, N1965, N278, N1523);
or OR2 (N1969, N1967, N954);
nand NAND3 (N1970, N1946, N47, N545);
or OR4 (N1971, N1962, N1038, N1183, N205);
nand NAND3 (N1972, N1971, N243, N224);
xor XOR2 (N1973, N1972, N942);
buf BUF1 (N1974, N1964);
nor NOR3 (N1975, N1966, N939, N419);
or OR4 (N1976, N1970, N827, N1869, N1733);
buf BUF1 (N1977, N1969);
buf BUF1 (N1978, N1943);
nand NAND4 (N1979, N1977, N530, N1138, N338);
nor NOR4 (N1980, N1959, N1086, N140, N1099);
not NOT1 (N1981, N1980);
buf BUF1 (N1982, N1968);
and AND3 (N1983, N1978, N1929, N137);
nand NAND3 (N1984, N1976, N112, N455);
buf BUF1 (N1985, N1983);
buf BUF1 (N1986, N1982);
buf BUF1 (N1987, N1985);
xor XOR2 (N1988, N1952, N1829);
xor XOR2 (N1989, N1987, N674);
not NOT1 (N1990, N1979);
buf BUF1 (N1991, N1975);
not NOT1 (N1992, N1990);
xor XOR2 (N1993, N1963, N1828);
not NOT1 (N1994, N1989);
and AND3 (N1995, N1992, N1298, N138);
and AND2 (N1996, N1974, N450);
nand NAND3 (N1997, N1988, N111, N235);
nor NOR4 (N1998, N1997, N690, N1267, N1562);
and AND4 (N1999, N1994, N1440, N1569, N1170);
nor NOR3 (N2000, N1996, N609, N1438);
nor NOR4 (N2001, N2000, N1409, N313, N451);
not NOT1 (N2002, N1984);
xor XOR2 (N2003, N1998, N276);
nor NOR4 (N2004, N1993, N1186, N1276, N939);
or OR3 (N2005, N2003, N406, N1211);
xor XOR2 (N2006, N1991, N463);
buf BUF1 (N2007, N1981);
nand NAND3 (N2008, N2002, N242, N603);
nor NOR3 (N2009, N2004, N722, N889);
nand NAND3 (N2010, N1973, N970, N1832);
or OR4 (N2011, N2005, N92, N1378, N680);
buf BUF1 (N2012, N2006);
xor XOR2 (N2013, N2012, N70);
nand NAND2 (N2014, N2011, N457);
buf BUF1 (N2015, N2001);
and AND3 (N2016, N2013, N744, N1165);
nand NAND2 (N2017, N2007, N1253);
and AND2 (N2018, N2010, N1630);
nand NAND3 (N2019, N2017, N1697, N1249);
not NOT1 (N2020, N1999);
not NOT1 (N2021, N2020);
buf BUF1 (N2022, N2019);
nand NAND4 (N2023, N2009, N549, N710, N602);
nor NOR2 (N2024, N2016, N1531);
and AND3 (N2025, N2023, N1624, N851);
xor XOR2 (N2026, N2008, N41);
xor XOR2 (N2027, N1986, N1722);
xor XOR2 (N2028, N2021, N1389);
nor NOR4 (N2029, N2018, N2002, N864, N1475);
nor NOR2 (N2030, N2024, N616);
nand NAND4 (N2031, N2027, N276, N608, N1369);
nand NAND3 (N2032, N2026, N1857, N1252);
buf BUF1 (N2033, N2015);
nand NAND4 (N2034, N1995, N1384, N810, N389);
or OR2 (N2035, N2022, N1280);
or OR2 (N2036, N2025, N361);
buf BUF1 (N2037, N2028);
nand NAND2 (N2038, N2014, N2011);
or OR4 (N2039, N2030, N1864, N45, N1669);
nand NAND3 (N2040, N2031, N1314, N1220);
or OR3 (N2041, N2038, N854, N350);
or OR2 (N2042, N2037, N578);
nor NOR3 (N2043, N2039, N1963, N1648);
or OR2 (N2044, N2035, N1666);
and AND3 (N2045, N2033, N1142, N1494);
xor XOR2 (N2046, N2029, N451);
not NOT1 (N2047, N2032);
buf BUF1 (N2048, N2036);
nor NOR2 (N2049, N2044, N737);
nor NOR4 (N2050, N2049, N1180, N1100, N1196);
or OR3 (N2051, N2040, N963, N806);
xor XOR2 (N2052, N2034, N1570);
nor NOR3 (N2053, N2046, N342, N1655);
nor NOR3 (N2054, N2052, N1160, N973);
buf BUF1 (N2055, N2053);
nor NOR4 (N2056, N2051, N1956, N878, N772);
nor NOR3 (N2057, N2055, N794, N787);
xor XOR2 (N2058, N2057, N1140);
not NOT1 (N2059, N2058);
nand NAND4 (N2060, N2050, N929, N137, N532);
nor NOR2 (N2061, N2047, N1668);
nand NAND3 (N2062, N2060, N572, N964);
and AND2 (N2063, N2054, N597);
xor XOR2 (N2064, N2042, N1306);
nand NAND4 (N2065, N2041, N700, N2033, N292);
buf BUF1 (N2066, N2045);
buf BUF1 (N2067, N2062);
buf BUF1 (N2068, N2059);
buf BUF1 (N2069, N2056);
buf BUF1 (N2070, N2066);
not NOT1 (N2071, N2064);
xor XOR2 (N2072, N2043, N1165);
xor XOR2 (N2073, N2061, N1437);
nor NOR4 (N2074, N2065, N760, N1499, N244);
not NOT1 (N2075, N2072);
or OR4 (N2076, N2074, N645, N1716, N1623);
nand NAND2 (N2077, N2073, N887);
xor XOR2 (N2078, N2069, N1585);
nand NAND2 (N2079, N2063, N480);
nor NOR3 (N2080, N2067, N659, N738);
or OR3 (N2081, N2077, N628, N2068);
and AND3 (N2082, N921, N955, N19);
and AND4 (N2083, N2081, N301, N1635, N1734);
nand NAND2 (N2084, N2078, N1103);
not NOT1 (N2085, N2080);
nand NAND4 (N2086, N2048, N562, N1197, N1829);
not NOT1 (N2087, N2084);
xor XOR2 (N2088, N2071, N1294);
nand NAND2 (N2089, N2087, N960);
or OR2 (N2090, N2083, N1494);
not NOT1 (N2091, N2085);
or OR2 (N2092, N2076, N1371);
buf BUF1 (N2093, N2082);
and AND4 (N2094, N2088, N194, N1082, N1842);
nor NOR2 (N2095, N2075, N1389);
not NOT1 (N2096, N2095);
and AND3 (N2097, N2092, N242, N60);
or OR3 (N2098, N2096, N1046, N1712);
buf BUF1 (N2099, N2093);
nand NAND2 (N2100, N2086, N1768);
xor XOR2 (N2101, N2091, N1041);
not NOT1 (N2102, N2090);
xor XOR2 (N2103, N2079, N1849);
nand NAND3 (N2104, N2089, N1629, N601);
not NOT1 (N2105, N2102);
and AND2 (N2106, N2070, N1124);
or OR4 (N2107, N2099, N1997, N1067, N963);
and AND3 (N2108, N2094, N676, N1127);
not NOT1 (N2109, N2107);
nor NOR2 (N2110, N2103, N1809);
nor NOR4 (N2111, N2109, N2068, N1126, N923);
or OR4 (N2112, N2097, N1430, N659, N203);
or OR4 (N2113, N2112, N1175, N776, N1918);
or OR2 (N2114, N2106, N1250);
nand NAND4 (N2115, N2108, N1392, N860, N829);
or OR4 (N2116, N2111, N1750, N828, N906);
nor NOR2 (N2117, N2100, N1278);
or OR2 (N2118, N2114, N1574);
xor XOR2 (N2119, N2118, N1258);
and AND2 (N2120, N2117, N1111);
nor NOR3 (N2121, N2113, N1142, N953);
or OR4 (N2122, N2098, N1957, N252, N1721);
not NOT1 (N2123, N2105);
and AND4 (N2124, N2104, N998, N1548, N1993);
and AND2 (N2125, N2115, N1166);
xor XOR2 (N2126, N2123, N1515);
xor XOR2 (N2127, N2121, N131);
or OR2 (N2128, N2110, N941);
not NOT1 (N2129, N2126);
xor XOR2 (N2130, N2116, N1211);
buf BUF1 (N2131, N2120);
nor NOR2 (N2132, N2129, N764);
nor NOR3 (N2133, N2132, N1814, N1837);
nor NOR4 (N2134, N2124, N966, N1250, N1569);
nand NAND3 (N2135, N2119, N1591, N1937);
nor NOR3 (N2136, N2101, N650, N1206);
nand NAND3 (N2137, N2135, N1026, N578);
not NOT1 (N2138, N2128);
nand NAND4 (N2139, N2134, N1815, N1893, N1223);
nor NOR3 (N2140, N2127, N629, N39);
nor NOR3 (N2141, N2130, N907, N2030);
or OR2 (N2142, N2122, N1203);
and AND3 (N2143, N2137, N341, N973);
or OR3 (N2144, N2139, N1976, N529);
or OR2 (N2145, N2131, N1218);
and AND4 (N2146, N2143, N1920, N865, N976);
nand NAND2 (N2147, N2138, N1764);
not NOT1 (N2148, N2136);
nand NAND3 (N2149, N2125, N1958, N309);
or OR2 (N2150, N2141, N1179);
and AND3 (N2151, N2148, N125, N347);
and AND4 (N2152, N2150, N1533, N2140, N689);
or OR4 (N2153, N1167, N835, N1208, N1355);
not NOT1 (N2154, N2151);
buf BUF1 (N2155, N2153);
nand NAND4 (N2156, N2155, N898, N1997, N1759);
xor XOR2 (N2157, N2154, N1838);
buf BUF1 (N2158, N2144);
not NOT1 (N2159, N2145);
and AND2 (N2160, N2133, N1643);
and AND2 (N2161, N2146, N1899);
and AND4 (N2162, N2161, N881, N865, N172);
xor XOR2 (N2163, N2157, N671);
nor NOR3 (N2164, N2156, N501, N1713);
and AND3 (N2165, N2158, N2134, N1247);
xor XOR2 (N2166, N2152, N1701);
or OR4 (N2167, N2142, N703, N1988, N700);
buf BUF1 (N2168, N2147);
not NOT1 (N2169, N2167);
nand NAND4 (N2170, N2168, N1874, N1617, N1862);
not NOT1 (N2171, N2164);
nand NAND3 (N2172, N2171, N1276, N656);
and AND3 (N2173, N2159, N695, N1536);
nor NOR3 (N2174, N2160, N2044, N1656);
xor XOR2 (N2175, N2172, N739);
not NOT1 (N2176, N2162);
nand NAND4 (N2177, N2173, N1121, N1009, N1057);
and AND2 (N2178, N2174, N1757);
xor XOR2 (N2179, N2165, N1559);
nor NOR4 (N2180, N2177, N53, N1269, N533);
buf BUF1 (N2181, N2163);
buf BUF1 (N2182, N2180);
xor XOR2 (N2183, N2175, N1408);
buf BUF1 (N2184, N2179);
xor XOR2 (N2185, N2183, N421);
buf BUF1 (N2186, N2169);
buf BUF1 (N2187, N2178);
buf BUF1 (N2188, N2170);
not NOT1 (N2189, N2185);
buf BUF1 (N2190, N2182);
not NOT1 (N2191, N2149);
xor XOR2 (N2192, N2176, N1448);
not NOT1 (N2193, N2184);
xor XOR2 (N2194, N2188, N1494);
nand NAND3 (N2195, N2187, N2153, N542);
xor XOR2 (N2196, N2189, N1719);
xor XOR2 (N2197, N2195, N696);
nor NOR2 (N2198, N2166, N324);
or OR2 (N2199, N2198, N1833);
nor NOR3 (N2200, N2192, N1653, N924);
nand NAND3 (N2201, N2199, N1642, N1503);
not NOT1 (N2202, N2193);
buf BUF1 (N2203, N2200);
nand NAND2 (N2204, N2201, N1863);
or OR2 (N2205, N2181, N1298);
not NOT1 (N2206, N2204);
or OR3 (N2207, N2191, N675, N1669);
nand NAND2 (N2208, N2207, N1433);
nor NOR2 (N2209, N2186, N1525);
not NOT1 (N2210, N2205);
nand NAND4 (N2211, N2210, N293, N1141, N1517);
nand NAND4 (N2212, N2211, N2120, N735, N411);
not NOT1 (N2213, N2209);
or OR4 (N2214, N2213, N1693, N157, N589);
and AND4 (N2215, N2197, N1828, N495, N569);
not NOT1 (N2216, N2214);
and AND4 (N2217, N2194, N470, N1612, N1484);
not NOT1 (N2218, N2212);
nor NOR4 (N2219, N2202, N1278, N239, N302);
not NOT1 (N2220, N2217);
not NOT1 (N2221, N2216);
nand NAND4 (N2222, N2208, N1019, N1216, N493);
and AND2 (N2223, N2206, N1454);
or OR4 (N2224, N2190, N1385, N955, N2161);
or OR2 (N2225, N2221, N1797);
nor NOR3 (N2226, N2196, N360, N664);
xor XOR2 (N2227, N2219, N1548);
nand NAND2 (N2228, N2222, N2164);
or OR4 (N2229, N2227, N1885, N1067, N1680);
not NOT1 (N2230, N2215);
and AND4 (N2231, N2203, N2216, N1094, N2007);
nand NAND4 (N2232, N2220, N64, N1286, N482);
xor XOR2 (N2233, N2228, N183);
not NOT1 (N2234, N2224);
and AND3 (N2235, N2233, N906, N1038);
xor XOR2 (N2236, N2223, N1496);
not NOT1 (N2237, N2218);
nor NOR4 (N2238, N2235, N1125, N1822, N914);
nand NAND4 (N2239, N2229, N1519, N1137, N1893);
nand NAND2 (N2240, N2234, N422);
and AND4 (N2241, N2237, N279, N1251, N1208);
and AND2 (N2242, N2241, N381);
buf BUF1 (N2243, N2242);
nand NAND4 (N2244, N2236, N350, N201, N177);
nand NAND2 (N2245, N2244, N43);
nand NAND3 (N2246, N2226, N1124, N176);
nand NAND3 (N2247, N2230, N1941, N379);
buf BUF1 (N2248, N2246);
and AND4 (N2249, N2240, N1849, N2111, N507);
not NOT1 (N2250, N2247);
not NOT1 (N2251, N2245);
nor NOR3 (N2252, N2239, N1841, N1649);
buf BUF1 (N2253, N2248);
not NOT1 (N2254, N2249);
nor NOR4 (N2255, N2254, N202, N990, N1754);
not NOT1 (N2256, N2232);
not NOT1 (N2257, N2256);
not NOT1 (N2258, N2243);
not NOT1 (N2259, N2225);
nand NAND2 (N2260, N2253, N729);
and AND2 (N2261, N2260, N717);
buf BUF1 (N2262, N2231);
and AND3 (N2263, N2259, N146, N116);
or OR4 (N2264, N2258, N1787, N1377, N1220);
xor XOR2 (N2265, N2263, N715);
or OR2 (N2266, N2265, N1235);
or OR3 (N2267, N2250, N404, N957);
and AND3 (N2268, N2252, N2010, N249);
xor XOR2 (N2269, N2268, N940);
or OR3 (N2270, N2257, N382, N830);
xor XOR2 (N2271, N2264, N2266);
and AND3 (N2272, N1016, N1353, N314);
buf BUF1 (N2273, N2271);
and AND3 (N2274, N2262, N1281, N475);
nand NAND3 (N2275, N2272, N1816, N427);
xor XOR2 (N2276, N2275, N154);
or OR4 (N2277, N2261, N2175, N371, N613);
xor XOR2 (N2278, N2238, N1698);
or OR2 (N2279, N2270, N308);
nor NOR4 (N2280, N2267, N2005, N900, N1630);
buf BUF1 (N2281, N2280);
xor XOR2 (N2282, N2278, N1447);
not NOT1 (N2283, N2255);
xor XOR2 (N2284, N2251, N421);
nor NOR4 (N2285, N2274, N1695, N880, N359);
or OR3 (N2286, N2284, N710, N573);
buf BUF1 (N2287, N2283);
nor NOR4 (N2288, N2273, N1611, N381, N958);
xor XOR2 (N2289, N2279, N1590);
or OR3 (N2290, N2276, N1060, N1094);
buf BUF1 (N2291, N2281);
nor NOR2 (N2292, N2282, N526);
or OR3 (N2293, N2288, N1793, N1778);
buf BUF1 (N2294, N2289);
nor NOR3 (N2295, N2277, N2182, N1802);
xor XOR2 (N2296, N2269, N1295);
nand NAND3 (N2297, N2287, N443, N2189);
xor XOR2 (N2298, N2294, N275);
nand NAND3 (N2299, N2290, N1747, N1374);
not NOT1 (N2300, N2286);
not NOT1 (N2301, N2297);
and AND2 (N2302, N2298, N561);
buf BUF1 (N2303, N2291);
not NOT1 (N2304, N2296);
and AND4 (N2305, N2304, N1520, N552, N1299);
nand NAND2 (N2306, N2299, N1452);
not NOT1 (N2307, N2300);
or OR3 (N2308, N2303, N2266, N978);
xor XOR2 (N2309, N2306, N2085);
nand NAND2 (N2310, N2307, N390);
nor NOR4 (N2311, N2305, N319, N2142, N1560);
not NOT1 (N2312, N2301);
buf BUF1 (N2313, N2308);
not NOT1 (N2314, N2311);
and AND2 (N2315, N2309, N650);
not NOT1 (N2316, N2302);
not NOT1 (N2317, N2310);
and AND4 (N2318, N2315, N1534, N750, N437);
nor NOR2 (N2319, N2292, N1185);
buf BUF1 (N2320, N2317);
nand NAND4 (N2321, N2320, N1392, N198, N671);
not NOT1 (N2322, N2285);
or OR4 (N2323, N2295, N1745, N864, N1454);
nor NOR2 (N2324, N2319, N356);
nand NAND3 (N2325, N2313, N818, N579);
and AND3 (N2326, N2324, N498, N2163);
buf BUF1 (N2327, N2322);
or OR4 (N2328, N2323, N160, N196, N600);
and AND3 (N2329, N2327, N2090, N199);
nand NAND2 (N2330, N2293, N627);
nor NOR2 (N2331, N2326, N1656);
buf BUF1 (N2332, N2321);
nand NAND4 (N2333, N2316, N1860, N411, N1338);
and AND3 (N2334, N2325, N116, N941);
xor XOR2 (N2335, N2314, N1179);
xor XOR2 (N2336, N2329, N1408);
xor XOR2 (N2337, N2332, N1085);
buf BUF1 (N2338, N2331);
and AND2 (N2339, N2330, N1798);
buf BUF1 (N2340, N2334);
or OR3 (N2341, N2339, N745, N1502);
xor XOR2 (N2342, N2335, N350);
nand NAND4 (N2343, N2333, N706, N1809, N2088);
xor XOR2 (N2344, N2328, N185);
nand NAND2 (N2345, N2336, N1232);
xor XOR2 (N2346, N2343, N97);
buf BUF1 (N2347, N2345);
buf BUF1 (N2348, N2341);
or OR2 (N2349, N2342, N2106);
buf BUF1 (N2350, N2318);
or OR2 (N2351, N2338, N1025);
nor NOR2 (N2352, N2346, N1861);
nor NOR3 (N2353, N2351, N772, N774);
nand NAND4 (N2354, N2348, N117, N1125, N1963);
or OR2 (N2355, N2337, N374);
nand NAND3 (N2356, N2349, N218, N1613);
and AND4 (N2357, N2347, N376, N1289, N646);
nand NAND2 (N2358, N2344, N663);
xor XOR2 (N2359, N2355, N340);
nor NOR4 (N2360, N2353, N2113, N1535, N757);
xor XOR2 (N2361, N2352, N1932);
buf BUF1 (N2362, N2356);
nand NAND2 (N2363, N2360, N313);
buf BUF1 (N2364, N2312);
buf BUF1 (N2365, N2364);
buf BUF1 (N2366, N2354);
and AND2 (N2367, N2359, N2176);
xor XOR2 (N2368, N2367, N368);
buf BUF1 (N2369, N2363);
nor NOR2 (N2370, N2340, N1979);
nand NAND2 (N2371, N2358, N319);
not NOT1 (N2372, N2368);
and AND3 (N2373, N2362, N1702, N631);
nor NOR4 (N2374, N2369, N1825, N2146, N161);
nor NOR3 (N2375, N2373, N864, N548);
nor NOR2 (N2376, N2350, N2120);
xor XOR2 (N2377, N2357, N1671);
and AND4 (N2378, N2366, N1142, N1021, N1279);
and AND2 (N2379, N2370, N975);
buf BUF1 (N2380, N2365);
nand NAND4 (N2381, N2377, N1305, N1214, N971);
and AND3 (N2382, N2371, N1099, N525);
and AND2 (N2383, N2380, N1660);
not NOT1 (N2384, N2383);
and AND2 (N2385, N2372, N2342);
or OR2 (N2386, N2382, N1497);
nor NOR4 (N2387, N2379, N100, N55, N1273);
xor XOR2 (N2388, N2375, N1659);
and AND4 (N2389, N2388, N1264, N1334, N820);
buf BUF1 (N2390, N2384);
nand NAND2 (N2391, N2386, N1864);
and AND2 (N2392, N2376, N2220);
not NOT1 (N2393, N2389);
and AND2 (N2394, N2391, N1501);
and AND4 (N2395, N2374, N946, N1842, N2044);
and AND3 (N2396, N2393, N2230, N54);
buf BUF1 (N2397, N2394);
nor NOR4 (N2398, N2396, N1413, N1125, N2058);
xor XOR2 (N2399, N2397, N140);
xor XOR2 (N2400, N2385, N628);
nor NOR3 (N2401, N2390, N1407, N686);
not NOT1 (N2402, N2361);
or OR4 (N2403, N2387, N167, N782, N1899);
not NOT1 (N2404, N2395);
not NOT1 (N2405, N2400);
and AND4 (N2406, N2401, N764, N52, N1375);
or OR3 (N2407, N2392, N876, N692);
xor XOR2 (N2408, N2403, N110);
and AND4 (N2409, N2381, N1398, N2143, N401);
and AND4 (N2410, N2409, N1514, N609, N682);
nand NAND3 (N2411, N2404, N225, N329);
or OR2 (N2412, N2398, N253);
xor XOR2 (N2413, N2412, N997);
nor NOR4 (N2414, N2378, N923, N845, N1891);
and AND2 (N2415, N2399, N2032);
buf BUF1 (N2416, N2407);
buf BUF1 (N2417, N2406);
nor NOR2 (N2418, N2413, N1663);
or OR2 (N2419, N2410, N2402);
nand NAND4 (N2420, N2398, N1251, N952, N1293);
and AND4 (N2421, N2416, N556, N205, N2236);
not NOT1 (N2422, N2405);
buf BUF1 (N2423, N2421);
nor NOR3 (N2424, N2418, N2333, N1135);
buf BUF1 (N2425, N2414);
nor NOR3 (N2426, N2424, N2337, N2397);
not NOT1 (N2427, N2422);
nor NOR4 (N2428, N2423, N1237, N593, N1511);
nor NOR2 (N2429, N2427, N91);
xor XOR2 (N2430, N2419, N2183);
nor NOR2 (N2431, N2430, N1536);
nand NAND2 (N2432, N2431, N653);
and AND2 (N2433, N2415, N405);
not NOT1 (N2434, N2417);
or OR4 (N2435, N2426, N2057, N2149, N794);
and AND2 (N2436, N2420, N2108);
and AND2 (N2437, N2411, N804);
or OR3 (N2438, N2435, N1198, N1584);
xor XOR2 (N2439, N2437, N2105);
nor NOR3 (N2440, N2429, N686, N1806);
nand NAND3 (N2441, N2436, N2422, N817);
nand NAND2 (N2442, N2408, N1969);
or OR3 (N2443, N2441, N995, N1831);
nor NOR3 (N2444, N2439, N1083, N1346);
xor XOR2 (N2445, N2434, N575);
not NOT1 (N2446, N2428);
nand NAND2 (N2447, N2445, N2099);
buf BUF1 (N2448, N2425);
nand NAND3 (N2449, N2447, N2281, N856);
xor XOR2 (N2450, N2432, N809);
or OR3 (N2451, N2433, N197, N225);
nor NOR3 (N2452, N2440, N2003, N1581);
nand NAND2 (N2453, N2448, N1793);
not NOT1 (N2454, N2452);
buf BUF1 (N2455, N2453);
nor NOR2 (N2456, N2443, N780);
and AND3 (N2457, N2446, N1377, N1086);
nor NOR4 (N2458, N2456, N617, N780, N1534);
or OR2 (N2459, N2451, N1532);
not NOT1 (N2460, N2458);
nor NOR4 (N2461, N2450, N2455, N1453, N2150);
nand NAND2 (N2462, N1708, N503);
or OR2 (N2463, N2459, N199);
buf BUF1 (N2464, N2461);
and AND3 (N2465, N2463, N2403, N2407);
or OR2 (N2466, N2454, N1762);
and AND3 (N2467, N2438, N1914, N695);
buf BUF1 (N2468, N2466);
and AND4 (N2469, N2465, N1305, N268, N2468);
nand NAND2 (N2470, N1582, N2442);
or OR4 (N2471, N2080, N2002, N352, N557);
and AND4 (N2472, N2444, N1385, N1994, N1986);
xor XOR2 (N2473, N2464, N207);
nand NAND2 (N2474, N2457, N2432);
and AND4 (N2475, N2462, N1751, N1972, N2177);
buf BUF1 (N2476, N2475);
xor XOR2 (N2477, N2476, N7);
nor NOR4 (N2478, N2472, N845, N741, N1226);
or OR3 (N2479, N2471, N1286, N571);
and AND3 (N2480, N2477, N1121, N971);
nor NOR2 (N2481, N2473, N1820);
and AND3 (N2482, N2479, N459, N1489);
and AND2 (N2483, N2481, N498);
nand NAND3 (N2484, N2460, N1732, N625);
buf BUF1 (N2485, N2484);
nor NOR4 (N2486, N2449, N611, N1618, N720);
and AND3 (N2487, N2486, N2430, N1405);
xor XOR2 (N2488, N2480, N1043);
nand NAND3 (N2489, N2487, N2131, N2394);
not NOT1 (N2490, N2478);
nand NAND4 (N2491, N2467, N696, N58, N62);
or OR3 (N2492, N2485, N944, N168);
and AND4 (N2493, N2470, N1729, N862, N100);
xor XOR2 (N2494, N2491, N1949);
nand NAND2 (N2495, N2490, N1275);
buf BUF1 (N2496, N2482);
nor NOR2 (N2497, N2483, N1513);
xor XOR2 (N2498, N2489, N2131);
and AND3 (N2499, N2469, N729, N1773);
nor NOR4 (N2500, N2493, N920, N2450, N713);
xor XOR2 (N2501, N2497, N961);
nor NOR4 (N2502, N2498, N1161, N45, N1468);
nor NOR2 (N2503, N2500, N989);
not NOT1 (N2504, N2503);
and AND2 (N2505, N2494, N1460);
xor XOR2 (N2506, N2474, N1233);
and AND2 (N2507, N2501, N107);
nand NAND4 (N2508, N2502, N426, N2103, N802);
nor NOR3 (N2509, N2488, N2225, N447);
and AND2 (N2510, N2505, N2357);
and AND2 (N2511, N2509, N1599);
nor NOR3 (N2512, N2504, N369, N1161);
xor XOR2 (N2513, N2507, N1307);
and AND3 (N2514, N2508, N583, N2268);
and AND2 (N2515, N2492, N1079);
endmodule