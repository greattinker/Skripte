// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20;

output N3203,N3218,N3209,N3215,N3211,N3210,N3219,N3201,N3216,N3220;

xor XOR2 (N21, N9, N6);
or OR3 (N22, N12, N12, N19);
nor NOR4 (N23, N10, N17, N9, N10);
nor NOR2 (N24, N7, N15);
nor NOR2 (N25, N15, N7);
nor NOR4 (N26, N24, N6, N20, N22);
xor XOR2 (N27, N3, N17);
or OR2 (N28, N16, N6);
xor XOR2 (N29, N28, N26);
not NOT1 (N30, N8);
nand NAND2 (N31, N18, N5);
buf BUF1 (N32, N26);
not NOT1 (N33, N13);
nand NAND2 (N34, N33, N5);
nand NAND4 (N35, N33, N2, N18, N22);
nor NOR4 (N36, N34, N26, N8, N32);
buf BUF1 (N37, N5);
xor XOR2 (N38, N37, N10);
xor XOR2 (N39, N27, N5);
xor XOR2 (N40, N38, N1);
or OR4 (N41, N25, N17, N34, N17);
and AND3 (N42, N35, N12, N28);
buf BUF1 (N43, N39);
xor XOR2 (N44, N41, N32);
xor XOR2 (N45, N21, N16);
and AND3 (N46, N44, N25, N7);
not NOT1 (N47, N42);
nand NAND2 (N48, N29, N15);
or OR3 (N49, N43, N20, N35);
buf BUF1 (N50, N46);
not NOT1 (N51, N45);
not NOT1 (N52, N23);
buf BUF1 (N53, N47);
buf BUF1 (N54, N51);
buf BUF1 (N55, N50);
xor XOR2 (N56, N48, N48);
nand NAND2 (N57, N55, N24);
or OR4 (N58, N56, N47, N19, N41);
nand NAND3 (N59, N58, N46, N24);
or OR4 (N60, N52, N32, N56, N39);
or OR3 (N61, N59, N15, N5);
nand NAND3 (N62, N40, N13, N21);
not NOT1 (N63, N54);
and AND4 (N64, N57, N29, N2, N42);
nand NAND2 (N65, N49, N43);
nor NOR4 (N66, N60, N37, N13, N32);
and AND2 (N67, N63, N22);
buf BUF1 (N68, N66);
or OR4 (N69, N31, N32, N33, N19);
and AND3 (N70, N61, N13, N44);
or OR3 (N71, N68, N12, N36);
xor XOR2 (N72, N3, N19);
not NOT1 (N73, N64);
nor NOR4 (N74, N71, N72, N46, N27);
not NOT1 (N75, N55);
xor XOR2 (N76, N74, N6);
and AND4 (N77, N62, N4, N71, N30);
nand NAND2 (N78, N35, N61);
buf BUF1 (N79, N53);
and AND4 (N80, N67, N35, N26, N61);
nor NOR4 (N81, N65, N44, N39, N12);
nand NAND2 (N82, N79, N72);
nor NOR3 (N83, N78, N22, N36);
buf BUF1 (N84, N83);
xor XOR2 (N85, N76, N10);
not NOT1 (N86, N69);
xor XOR2 (N87, N81, N36);
nand NAND4 (N88, N84, N1, N65, N16);
nand NAND4 (N89, N73, N72, N63, N4);
buf BUF1 (N90, N75);
not NOT1 (N91, N85);
or OR3 (N92, N86, N47, N18);
not NOT1 (N93, N87);
nand NAND3 (N94, N82, N88, N8);
xor XOR2 (N95, N26, N26);
buf BUF1 (N96, N95);
buf BUF1 (N97, N96);
buf BUF1 (N98, N80);
and AND4 (N99, N92, N50, N80, N72);
nor NOR3 (N100, N90, N59, N62);
xor XOR2 (N101, N93, N71);
not NOT1 (N102, N89);
nand NAND4 (N103, N77, N100, N11, N71);
xor XOR2 (N104, N85, N25);
not NOT1 (N105, N104);
and AND3 (N106, N91, N9, N14);
or OR3 (N107, N101, N49, N70);
nand NAND2 (N108, N7, N63);
and AND3 (N109, N107, N8, N50);
and AND3 (N110, N97, N40, N90);
nand NAND4 (N111, N98, N67, N67, N99);
not NOT1 (N112, N62);
xor XOR2 (N113, N94, N27);
and AND3 (N114, N110, N4, N19);
or OR2 (N115, N108, N76);
buf BUF1 (N116, N103);
nand NAND3 (N117, N114, N76, N8);
nor NOR3 (N118, N117, N49, N34);
buf BUF1 (N119, N118);
and AND3 (N120, N116, N49, N13);
nor NOR4 (N121, N112, N88, N35, N15);
and AND4 (N122, N113, N48, N72, N83);
or OR4 (N123, N109, N40, N109, N77);
xor XOR2 (N124, N111, N84);
not NOT1 (N125, N120);
not NOT1 (N126, N119);
nand NAND4 (N127, N115, N15, N12, N126);
nand NAND4 (N128, N53, N127, N50, N17);
and AND4 (N129, N5, N108, N54, N40);
nor NOR2 (N130, N124, N24);
nor NOR3 (N131, N123, N42, N32);
nor NOR4 (N132, N129, N33, N26, N84);
nor NOR4 (N133, N128, N56, N51, N28);
buf BUF1 (N134, N102);
not NOT1 (N135, N132);
buf BUF1 (N136, N106);
and AND2 (N137, N136, N24);
and AND4 (N138, N130, N1, N37, N101);
nand NAND3 (N139, N121, N74, N79);
nor NOR2 (N140, N138, N31);
or OR2 (N141, N122, N67);
and AND4 (N142, N134, N14, N11, N98);
nor NOR2 (N143, N142, N136);
buf BUF1 (N144, N105);
not NOT1 (N145, N131);
not NOT1 (N146, N140);
xor XOR2 (N147, N146, N44);
nor NOR2 (N148, N145, N66);
or OR4 (N149, N133, N134, N24, N12);
buf BUF1 (N150, N143);
nor NOR3 (N151, N150, N59, N65);
nand NAND2 (N152, N137, N146);
xor XOR2 (N153, N144, N44);
nand NAND2 (N154, N135, N99);
and AND3 (N155, N139, N91, N24);
nor NOR2 (N156, N155, N95);
and AND3 (N157, N152, N58, N13);
buf BUF1 (N158, N157);
nor NOR4 (N159, N149, N3, N86, N48);
or OR3 (N160, N159, N112, N153);
nor NOR4 (N161, N98, N154, N83, N89);
nand NAND2 (N162, N80, N49);
nor NOR4 (N163, N156, N81, N135, N76);
nand NAND4 (N164, N158, N132, N129, N29);
buf BUF1 (N165, N160);
nand NAND4 (N166, N163, N53, N141, N64);
xor XOR2 (N167, N15, N33);
nor NOR3 (N168, N147, N28, N93);
buf BUF1 (N169, N161);
nor NOR4 (N170, N125, N155, N134, N140);
nor NOR3 (N171, N164, N88, N94);
nor NOR2 (N172, N148, N94);
nor NOR2 (N173, N166, N171);
xor XOR2 (N174, N114, N160);
and AND3 (N175, N169, N70, N18);
nand NAND2 (N176, N165, N78);
or OR3 (N177, N174, N49, N54);
or OR2 (N178, N175, N119);
xor XOR2 (N179, N168, N178);
xor XOR2 (N180, N155, N144);
nor NOR2 (N181, N179, N82);
buf BUF1 (N182, N167);
buf BUF1 (N183, N173);
xor XOR2 (N184, N176, N60);
nand NAND2 (N185, N182, N42);
not NOT1 (N186, N184);
buf BUF1 (N187, N186);
buf BUF1 (N188, N181);
not NOT1 (N189, N180);
or OR3 (N190, N170, N31, N186);
and AND3 (N191, N190, N157, N152);
buf BUF1 (N192, N189);
or OR3 (N193, N177, N142, N19);
xor XOR2 (N194, N162, N182);
xor XOR2 (N195, N193, N54);
or OR2 (N196, N191, N115);
not NOT1 (N197, N183);
not NOT1 (N198, N151);
buf BUF1 (N199, N194);
not NOT1 (N200, N187);
nor NOR2 (N201, N196, N4);
xor XOR2 (N202, N195, N30);
and AND3 (N203, N200, N201, N190);
or OR4 (N204, N32, N170, N199, N127);
or OR2 (N205, N97, N140);
buf BUF1 (N206, N202);
not NOT1 (N207, N192);
nand NAND3 (N208, N206, N91, N77);
buf BUF1 (N209, N188);
not NOT1 (N210, N204);
buf BUF1 (N211, N172);
or OR4 (N212, N205, N92, N139, N143);
and AND2 (N213, N210, N150);
nor NOR4 (N214, N211, N88, N197, N136);
or OR3 (N215, N95, N128, N189);
buf BUF1 (N216, N209);
and AND4 (N217, N216, N33, N72, N164);
or OR2 (N218, N203, N157);
buf BUF1 (N219, N208);
xor XOR2 (N220, N185, N85);
xor XOR2 (N221, N213, N154);
or OR3 (N222, N220, N105, N179);
nor NOR2 (N223, N218, N145);
nor NOR3 (N224, N214, N66, N38);
not NOT1 (N225, N198);
buf BUF1 (N226, N222);
nor NOR4 (N227, N224, N46, N197, N87);
or OR4 (N228, N219, N217, N171, N43);
nor NOR4 (N229, N20, N36, N37, N205);
nand NAND2 (N230, N215, N107);
or OR3 (N231, N207, N167, N124);
nand NAND4 (N232, N231, N72, N126, N199);
buf BUF1 (N233, N230);
xor XOR2 (N234, N221, N195);
xor XOR2 (N235, N227, N221);
and AND4 (N236, N229, N227, N224, N16);
nor NOR4 (N237, N235, N83, N167, N109);
not NOT1 (N238, N212);
and AND3 (N239, N234, N94, N32);
or OR3 (N240, N225, N24, N15);
and AND3 (N241, N233, N74, N182);
not NOT1 (N242, N241);
and AND2 (N243, N236, N1);
buf BUF1 (N244, N238);
not NOT1 (N245, N242);
xor XOR2 (N246, N232, N238);
and AND3 (N247, N246, N128, N87);
or OR3 (N248, N244, N212, N175);
and AND4 (N249, N228, N152, N127, N7);
xor XOR2 (N250, N249, N169);
nor NOR2 (N251, N245, N180);
xor XOR2 (N252, N250, N78);
xor XOR2 (N253, N252, N63);
not NOT1 (N254, N237);
nor NOR3 (N255, N239, N104, N18);
or OR2 (N256, N255, N215);
or OR4 (N257, N251, N222, N131, N37);
buf BUF1 (N258, N256);
nor NOR2 (N259, N258, N177);
xor XOR2 (N260, N257, N137);
nor NOR4 (N261, N260, N162, N239, N12);
buf BUF1 (N262, N254);
or OR4 (N263, N253, N117, N40, N34);
nand NAND2 (N264, N248, N52);
not NOT1 (N265, N240);
and AND2 (N266, N261, N35);
and AND3 (N267, N266, N78, N73);
xor XOR2 (N268, N226, N126);
nand NAND2 (N269, N265, N233);
nand NAND2 (N270, N267, N183);
and AND2 (N271, N269, N96);
or OR2 (N272, N271, N196);
or OR2 (N273, N272, N32);
and AND4 (N274, N268, N254, N149, N16);
not NOT1 (N275, N262);
nand NAND2 (N276, N275, N38);
nor NOR3 (N277, N259, N271, N31);
nand NAND3 (N278, N273, N59, N51);
not NOT1 (N279, N276);
nand NAND2 (N280, N279, N184);
not NOT1 (N281, N278);
and AND2 (N282, N277, N167);
nor NOR4 (N283, N264, N44, N159, N251);
or OR2 (N284, N270, N67);
and AND3 (N285, N281, N41, N220);
xor XOR2 (N286, N247, N275);
xor XOR2 (N287, N223, N79);
and AND3 (N288, N263, N28, N184);
nor NOR2 (N289, N286, N279);
buf BUF1 (N290, N243);
nor NOR3 (N291, N280, N119, N165);
nor NOR3 (N292, N284, N223, N101);
buf BUF1 (N293, N288);
xor XOR2 (N294, N274, N201);
buf BUF1 (N295, N294);
not NOT1 (N296, N293);
or OR2 (N297, N291, N82);
or OR3 (N298, N285, N205, N13);
buf BUF1 (N299, N295);
nor NOR2 (N300, N283, N107);
and AND3 (N301, N289, N129, N147);
or OR3 (N302, N298, N93, N60);
buf BUF1 (N303, N301);
xor XOR2 (N304, N290, N60);
nor NOR2 (N305, N300, N164);
not NOT1 (N306, N302);
nor NOR2 (N307, N282, N80);
nor NOR3 (N308, N307, N258, N92);
buf BUF1 (N309, N308);
nand NAND4 (N310, N309, N127, N75, N6);
nor NOR3 (N311, N296, N228, N79);
and AND3 (N312, N292, N87, N119);
xor XOR2 (N313, N311, N235);
nor NOR3 (N314, N305, N216, N35);
buf BUF1 (N315, N287);
and AND2 (N316, N312, N127);
nor NOR4 (N317, N310, N233, N70, N114);
not NOT1 (N318, N314);
nor NOR2 (N319, N316, N125);
xor XOR2 (N320, N304, N79);
xor XOR2 (N321, N320, N250);
buf BUF1 (N322, N306);
nand NAND4 (N323, N319, N182, N272, N122);
or OR4 (N324, N318, N174, N81, N123);
or OR2 (N325, N317, N91);
xor XOR2 (N326, N324, N142);
nand NAND4 (N327, N321, N192, N218, N71);
buf BUF1 (N328, N297);
xor XOR2 (N329, N326, N207);
buf BUF1 (N330, N323);
buf BUF1 (N331, N329);
xor XOR2 (N332, N330, N262);
xor XOR2 (N333, N332, N88);
nor NOR4 (N334, N303, N142, N45, N92);
and AND4 (N335, N331, N72, N133, N142);
or OR3 (N336, N335, N107, N174);
buf BUF1 (N337, N322);
nor NOR4 (N338, N333, N309, N166, N160);
nand NAND2 (N339, N334, N128);
not NOT1 (N340, N337);
and AND4 (N341, N327, N152, N77, N306);
not NOT1 (N342, N315);
or OR2 (N343, N338, N68);
buf BUF1 (N344, N313);
or OR2 (N345, N343, N138);
not NOT1 (N346, N344);
or OR2 (N347, N328, N126);
and AND3 (N348, N346, N279, N315);
buf BUF1 (N349, N348);
and AND2 (N350, N347, N100);
or OR2 (N351, N345, N24);
not NOT1 (N352, N350);
not NOT1 (N353, N342);
nand NAND4 (N354, N341, N264, N131, N279);
buf BUF1 (N355, N336);
xor XOR2 (N356, N351, N305);
buf BUF1 (N357, N354);
or OR2 (N358, N299, N203);
or OR4 (N359, N339, N185, N22, N241);
or OR3 (N360, N349, N347, N335);
nor NOR4 (N361, N357, N66, N260, N333);
nor NOR2 (N362, N353, N87);
not NOT1 (N363, N361);
xor XOR2 (N364, N362, N189);
buf BUF1 (N365, N356);
xor XOR2 (N366, N340, N175);
or OR2 (N367, N365, N232);
nor NOR3 (N368, N364, N183, N152);
not NOT1 (N369, N352);
buf BUF1 (N370, N363);
or OR2 (N371, N368, N284);
and AND4 (N372, N360, N21, N360, N281);
and AND2 (N373, N366, N111);
xor XOR2 (N374, N372, N347);
and AND4 (N375, N355, N84, N339, N150);
and AND2 (N376, N371, N256);
not NOT1 (N377, N359);
and AND3 (N378, N369, N23, N17);
or OR2 (N379, N375, N355);
buf BUF1 (N380, N370);
and AND4 (N381, N358, N357, N190, N138);
or OR2 (N382, N377, N215);
nand NAND3 (N383, N325, N282, N56);
and AND3 (N384, N374, N74, N45);
or OR2 (N385, N383, N299);
xor XOR2 (N386, N367, N218);
xor XOR2 (N387, N379, N321);
xor XOR2 (N388, N376, N67);
nor NOR4 (N389, N384, N8, N52, N109);
nor NOR3 (N390, N387, N313, N215);
buf BUF1 (N391, N381);
not NOT1 (N392, N388);
nor NOR3 (N393, N390, N9, N7);
not NOT1 (N394, N385);
or OR3 (N395, N380, N94, N374);
not NOT1 (N396, N391);
nand NAND2 (N397, N378, N140);
or OR2 (N398, N394, N76);
nor NOR2 (N399, N373, N128);
nor NOR2 (N400, N386, N182);
nor NOR4 (N401, N389, N105, N378, N383);
and AND4 (N402, N397, N90, N227, N34);
nand NAND4 (N403, N393, N184, N356, N331);
nor NOR3 (N404, N400, N115, N155);
nand NAND2 (N405, N395, N349);
buf BUF1 (N406, N396);
or OR3 (N407, N402, N386, N246);
and AND3 (N408, N405, N30, N11);
nor NOR4 (N409, N398, N205, N360, N352);
not NOT1 (N410, N406);
xor XOR2 (N411, N408, N266);
or OR2 (N412, N382, N92);
xor XOR2 (N413, N392, N124);
nor NOR3 (N414, N411, N93, N236);
and AND4 (N415, N409, N315, N140, N330);
not NOT1 (N416, N415);
or OR2 (N417, N401, N316);
or OR2 (N418, N403, N403);
not NOT1 (N419, N417);
and AND4 (N420, N414, N159, N268, N257);
not NOT1 (N421, N416);
or OR3 (N422, N418, N90, N368);
xor XOR2 (N423, N420, N188);
nor NOR3 (N424, N410, N128, N330);
buf BUF1 (N425, N412);
buf BUF1 (N426, N421);
nor NOR3 (N427, N407, N421, N101);
or OR2 (N428, N425, N13);
nand NAND4 (N429, N422, N409, N92, N383);
not NOT1 (N430, N419);
not NOT1 (N431, N404);
or OR3 (N432, N424, N56, N32);
and AND2 (N433, N426, N143);
xor XOR2 (N434, N428, N164);
nand NAND4 (N435, N423, N408, N390, N371);
and AND2 (N436, N431, N16);
or OR2 (N437, N429, N226);
or OR2 (N438, N435, N162);
not NOT1 (N439, N399);
nand NAND3 (N440, N427, N260, N35);
buf BUF1 (N441, N430);
or OR4 (N442, N440, N307, N432, N311);
nand NAND3 (N443, N395, N421, N108);
and AND3 (N444, N413, N270, N159);
nand NAND3 (N445, N438, N102, N199);
xor XOR2 (N446, N441, N404);
not NOT1 (N447, N437);
not NOT1 (N448, N444);
or OR4 (N449, N433, N437, N278, N349);
and AND4 (N450, N445, N243, N153, N39);
nor NOR2 (N451, N446, N33);
nor NOR3 (N452, N449, N216, N138);
not NOT1 (N453, N439);
xor XOR2 (N454, N452, N43);
xor XOR2 (N455, N451, N43);
nand NAND2 (N456, N447, N453);
nand NAND2 (N457, N448, N302);
xor XOR2 (N458, N337, N97);
buf BUF1 (N459, N456);
nand NAND4 (N460, N443, N437, N331, N183);
or OR3 (N461, N450, N180, N85);
and AND4 (N462, N455, N164, N11, N29);
xor XOR2 (N463, N460, N94);
nand NAND4 (N464, N463, N130, N85, N152);
and AND3 (N465, N434, N37, N311);
and AND3 (N466, N465, N153, N271);
nor NOR4 (N467, N466, N308, N438, N290);
not NOT1 (N468, N467);
buf BUF1 (N469, N468);
nand NAND2 (N470, N464, N271);
and AND4 (N471, N470, N42, N233, N409);
not NOT1 (N472, N457);
nand NAND2 (N473, N436, N268);
not NOT1 (N474, N454);
nor NOR2 (N475, N458, N2);
and AND3 (N476, N472, N387, N305);
or OR2 (N477, N474, N83);
and AND2 (N478, N442, N415);
xor XOR2 (N479, N461, N411);
and AND4 (N480, N478, N139, N107, N189);
xor XOR2 (N481, N469, N292);
and AND4 (N482, N476, N95, N134, N431);
nand NAND4 (N483, N473, N359, N472, N466);
buf BUF1 (N484, N475);
or OR2 (N485, N480, N266);
and AND4 (N486, N471, N363, N84, N150);
xor XOR2 (N487, N486, N61);
nand NAND2 (N488, N482, N225);
buf BUF1 (N489, N477);
and AND4 (N490, N487, N255, N327, N69);
nand NAND3 (N491, N459, N462, N34);
not NOT1 (N492, N333);
and AND2 (N493, N479, N13);
xor XOR2 (N494, N488, N321);
xor XOR2 (N495, N485, N228);
nand NAND4 (N496, N490, N273, N381, N474);
buf BUF1 (N497, N492);
nand NAND2 (N498, N481, N417);
xor XOR2 (N499, N496, N60);
not NOT1 (N500, N497);
buf BUF1 (N501, N499);
and AND2 (N502, N491, N72);
or OR2 (N503, N498, N479);
not NOT1 (N504, N495);
or OR4 (N505, N502, N338, N334, N409);
or OR2 (N506, N493, N96);
nor NOR4 (N507, N483, N339, N199, N101);
and AND4 (N508, N494, N449, N99, N83);
xor XOR2 (N509, N484, N185);
and AND3 (N510, N503, N140, N432);
or OR4 (N511, N504, N424, N119, N345);
nand NAND4 (N512, N511, N283, N381, N51);
and AND4 (N513, N510, N84, N72, N352);
and AND4 (N514, N501, N315, N119, N415);
and AND4 (N515, N500, N155, N447, N266);
and AND4 (N516, N508, N183, N133, N508);
and AND3 (N517, N506, N249, N477);
xor XOR2 (N518, N516, N167);
and AND4 (N519, N515, N418, N109, N246);
and AND4 (N520, N513, N366, N50, N342);
xor XOR2 (N521, N518, N377);
or OR3 (N522, N512, N503, N15);
not NOT1 (N523, N507);
not NOT1 (N524, N519);
nand NAND3 (N525, N509, N204, N337);
not NOT1 (N526, N517);
not NOT1 (N527, N522);
nand NAND3 (N528, N520, N349, N107);
nor NOR4 (N529, N521, N318, N498, N308);
xor XOR2 (N530, N525, N82);
not NOT1 (N531, N523);
or OR2 (N532, N528, N296);
and AND3 (N533, N489, N141, N188);
or OR4 (N534, N530, N432, N403, N423);
and AND4 (N535, N524, N447, N312, N90);
not NOT1 (N536, N529);
not NOT1 (N537, N532);
and AND4 (N538, N534, N508, N212, N475);
nand NAND3 (N539, N531, N434, N520);
buf BUF1 (N540, N514);
buf BUF1 (N541, N533);
not NOT1 (N542, N541);
and AND3 (N543, N526, N21, N347);
or OR2 (N544, N505, N89);
xor XOR2 (N545, N543, N48);
nor NOR3 (N546, N544, N40, N283);
nor NOR4 (N547, N537, N408, N132, N79);
xor XOR2 (N548, N536, N339);
nor NOR3 (N549, N545, N465, N435);
buf BUF1 (N550, N539);
nor NOR2 (N551, N550, N161);
and AND2 (N552, N540, N234);
buf BUF1 (N553, N551);
nor NOR4 (N554, N548, N303, N259, N194);
or OR3 (N555, N546, N357, N534);
xor XOR2 (N556, N535, N432);
nand NAND3 (N557, N552, N301, N217);
not NOT1 (N558, N527);
buf BUF1 (N559, N555);
nand NAND4 (N560, N553, N63, N71, N60);
nand NAND2 (N561, N559, N336);
buf BUF1 (N562, N560);
or OR2 (N563, N549, N10);
not NOT1 (N564, N538);
nand NAND2 (N565, N562, N256);
or OR3 (N566, N556, N83, N291);
nand NAND3 (N567, N564, N285, N396);
or OR4 (N568, N567, N393, N220, N331);
nand NAND4 (N569, N547, N437, N272, N213);
buf BUF1 (N570, N565);
xor XOR2 (N571, N566, N72);
not NOT1 (N572, N557);
nor NOR4 (N573, N558, N269, N485, N363);
or OR3 (N574, N570, N264, N337);
nand NAND2 (N575, N563, N335);
nor NOR2 (N576, N575, N39);
not NOT1 (N577, N569);
nor NOR3 (N578, N574, N351, N221);
and AND4 (N579, N578, N218, N97, N530);
not NOT1 (N580, N579);
not NOT1 (N581, N571);
not NOT1 (N582, N580);
xor XOR2 (N583, N577, N203);
buf BUF1 (N584, N582);
nand NAND2 (N585, N572, N331);
nand NAND2 (N586, N568, N525);
not NOT1 (N587, N586);
not NOT1 (N588, N581);
buf BUF1 (N589, N561);
nor NOR2 (N590, N576, N385);
xor XOR2 (N591, N542, N458);
xor XOR2 (N592, N588, N262);
not NOT1 (N593, N585);
not NOT1 (N594, N593);
not NOT1 (N595, N590);
xor XOR2 (N596, N587, N298);
not NOT1 (N597, N584);
nor NOR4 (N598, N596, N186, N549, N511);
nand NAND2 (N599, N591, N3);
or OR4 (N600, N592, N148, N326, N122);
buf BUF1 (N601, N573);
nor NOR4 (N602, N601, N396, N193, N119);
xor XOR2 (N603, N595, N217);
xor XOR2 (N604, N554, N1);
nor NOR2 (N605, N604, N365);
nor NOR4 (N606, N602, N549, N219, N72);
nand NAND2 (N607, N583, N602);
not NOT1 (N608, N606);
nor NOR2 (N609, N600, N414);
not NOT1 (N610, N607);
or OR3 (N611, N594, N493, N480);
and AND2 (N612, N605, N102);
and AND3 (N613, N599, N54, N438);
or OR4 (N614, N589, N216, N600, N547);
nor NOR4 (N615, N609, N556, N598, N398);
and AND2 (N616, N589, N183);
buf BUF1 (N617, N616);
and AND2 (N618, N615, N439);
or OR4 (N619, N611, N200, N108, N25);
and AND3 (N620, N613, N432, N169);
or OR4 (N621, N612, N292, N131, N201);
buf BUF1 (N622, N614);
not NOT1 (N623, N608);
or OR4 (N624, N621, N202, N233, N447);
nor NOR2 (N625, N622, N426);
buf BUF1 (N626, N625);
and AND4 (N627, N624, N112, N612, N167);
and AND3 (N628, N617, N402, N451);
buf BUF1 (N629, N627);
nand NAND4 (N630, N597, N323, N309, N264);
buf BUF1 (N631, N620);
or OR3 (N632, N618, N401, N575);
xor XOR2 (N633, N631, N243);
nor NOR3 (N634, N630, N223, N368);
xor XOR2 (N635, N633, N413);
nand NAND4 (N636, N634, N568, N307, N84);
or OR3 (N637, N626, N116, N424);
xor XOR2 (N638, N623, N134);
buf BUF1 (N639, N635);
not NOT1 (N640, N638);
xor XOR2 (N641, N610, N610);
nor NOR3 (N642, N639, N505, N343);
nor NOR3 (N643, N641, N68, N168);
and AND3 (N644, N636, N448, N353);
nor NOR4 (N645, N642, N118, N568, N559);
nor NOR2 (N646, N629, N430);
nand NAND4 (N647, N603, N68, N429, N484);
not NOT1 (N648, N619);
buf BUF1 (N649, N644);
and AND2 (N650, N628, N157);
nand NAND2 (N651, N643, N269);
nor NOR2 (N652, N640, N221);
nor NOR3 (N653, N652, N236, N191);
nand NAND3 (N654, N646, N387, N113);
or OR4 (N655, N645, N304, N640, N614);
buf BUF1 (N656, N655);
xor XOR2 (N657, N653, N520);
not NOT1 (N658, N657);
nor NOR4 (N659, N650, N268, N396, N487);
and AND4 (N660, N648, N138, N254, N653);
xor XOR2 (N661, N659, N207);
and AND3 (N662, N661, N262, N645);
not NOT1 (N663, N651);
xor XOR2 (N664, N663, N451);
nand NAND4 (N665, N637, N283, N664, N113);
and AND3 (N666, N185, N247, N516);
nor NOR2 (N667, N654, N57);
buf BUF1 (N668, N667);
and AND3 (N669, N660, N237, N612);
nor NOR4 (N670, N662, N380, N298, N299);
nand NAND2 (N671, N656, N535);
and AND3 (N672, N665, N95, N358);
nor NOR3 (N673, N668, N567, N201);
nor NOR3 (N674, N666, N29, N429);
buf BUF1 (N675, N632);
buf BUF1 (N676, N647);
not NOT1 (N677, N676);
nor NOR3 (N678, N671, N199, N579);
not NOT1 (N679, N675);
nand NAND4 (N680, N672, N287, N439, N26);
or OR4 (N681, N674, N318, N330, N363);
or OR3 (N682, N677, N31, N422);
buf BUF1 (N683, N682);
not NOT1 (N684, N681);
nor NOR3 (N685, N678, N511, N70);
or OR3 (N686, N649, N575, N17);
nand NAND2 (N687, N683, N651);
nand NAND2 (N688, N658, N182);
buf BUF1 (N689, N687);
xor XOR2 (N690, N689, N535);
buf BUF1 (N691, N690);
buf BUF1 (N692, N684);
or OR2 (N693, N679, N259);
and AND2 (N694, N670, N39);
nand NAND3 (N695, N693, N364, N665);
not NOT1 (N696, N669);
buf BUF1 (N697, N696);
xor XOR2 (N698, N688, N523);
buf BUF1 (N699, N698);
not NOT1 (N700, N699);
not NOT1 (N701, N680);
not NOT1 (N702, N701);
not NOT1 (N703, N700);
nand NAND3 (N704, N692, N158, N502);
nand NAND2 (N705, N673, N161);
and AND2 (N706, N691, N126);
or OR2 (N707, N704, N410);
or OR2 (N708, N703, N494);
buf BUF1 (N709, N697);
nor NOR2 (N710, N709, N358);
not NOT1 (N711, N708);
and AND3 (N712, N694, N84, N632);
nand NAND2 (N713, N707, N379);
nor NOR3 (N714, N695, N184, N138);
nand NAND2 (N715, N713, N380);
and AND2 (N716, N685, N446);
nand NAND2 (N717, N715, N632);
and AND4 (N718, N711, N26, N468, N495);
nor NOR2 (N719, N702, N54);
or OR3 (N720, N706, N712, N638);
or OR2 (N721, N154, N586);
not NOT1 (N722, N721);
or OR2 (N723, N705, N194);
nor NOR2 (N724, N723, N367);
and AND4 (N725, N724, N248, N245, N478);
buf BUF1 (N726, N714);
buf BUF1 (N727, N725);
nand NAND4 (N728, N726, N721, N605, N655);
nand NAND3 (N729, N727, N187, N508);
and AND3 (N730, N729, N679, N466);
nand NAND3 (N731, N686, N661, N609);
not NOT1 (N732, N719);
nor NOR3 (N733, N718, N500, N99);
xor XOR2 (N734, N710, N376);
nor NOR4 (N735, N728, N465, N323, N513);
buf BUF1 (N736, N720);
buf BUF1 (N737, N716);
xor XOR2 (N738, N735, N732);
not NOT1 (N739, N272);
nor NOR2 (N740, N736, N393);
nand NAND2 (N741, N722, N94);
buf BUF1 (N742, N730);
and AND4 (N743, N742, N658, N149, N670);
nand NAND2 (N744, N741, N164);
or OR4 (N745, N738, N59, N139, N727);
buf BUF1 (N746, N744);
or OR3 (N747, N737, N428, N189);
nand NAND3 (N748, N731, N690, N149);
and AND3 (N749, N733, N649, N714);
buf BUF1 (N750, N748);
and AND2 (N751, N717, N285);
xor XOR2 (N752, N745, N347);
not NOT1 (N753, N743);
nand NAND4 (N754, N749, N12, N357, N590);
not NOT1 (N755, N746);
nor NOR4 (N756, N754, N447, N591, N303);
nand NAND2 (N757, N755, N212);
and AND4 (N758, N757, N14, N670, N352);
nand NAND2 (N759, N758, N406);
and AND4 (N760, N734, N552, N722, N144);
nor NOR4 (N761, N752, N542, N452, N442);
buf BUF1 (N762, N740);
or OR4 (N763, N739, N528, N243, N621);
or OR4 (N764, N750, N557, N124, N112);
and AND3 (N765, N751, N269, N7);
and AND4 (N766, N761, N247, N447, N549);
and AND3 (N767, N762, N66, N157);
nand NAND2 (N768, N763, N433);
not NOT1 (N769, N747);
or OR2 (N770, N766, N627);
or OR2 (N771, N753, N458);
nand NAND4 (N772, N760, N376, N283, N336);
xor XOR2 (N773, N759, N623);
xor XOR2 (N774, N764, N627);
and AND2 (N775, N770, N227);
or OR3 (N776, N769, N605, N358);
nand NAND3 (N777, N776, N154, N626);
buf BUF1 (N778, N774);
and AND3 (N779, N775, N537, N307);
and AND2 (N780, N756, N319);
xor XOR2 (N781, N772, N542);
or OR4 (N782, N768, N513, N499, N201);
xor XOR2 (N783, N781, N549);
nand NAND4 (N784, N771, N703, N626, N405);
xor XOR2 (N785, N765, N619);
not NOT1 (N786, N785);
buf BUF1 (N787, N784);
and AND2 (N788, N780, N86);
buf BUF1 (N789, N788);
or OR3 (N790, N779, N21, N671);
buf BUF1 (N791, N786);
nand NAND4 (N792, N767, N427, N351, N122);
not NOT1 (N793, N773);
or OR2 (N794, N790, N711);
or OR4 (N795, N792, N442, N290, N136);
or OR2 (N796, N791, N726);
buf BUF1 (N797, N787);
nand NAND4 (N798, N777, N28, N33, N64);
nand NAND2 (N799, N796, N36);
nor NOR4 (N800, N789, N414, N271, N343);
buf BUF1 (N801, N783);
and AND2 (N802, N798, N567);
xor XOR2 (N803, N799, N490);
and AND3 (N804, N801, N548, N450);
not NOT1 (N805, N778);
nor NOR4 (N806, N803, N240, N426, N494);
nor NOR3 (N807, N795, N499, N200);
or OR2 (N808, N802, N191);
buf BUF1 (N809, N782);
or OR2 (N810, N794, N495);
or OR4 (N811, N804, N228, N662, N55);
and AND2 (N812, N808, N572);
buf BUF1 (N813, N806);
or OR2 (N814, N797, N33);
not NOT1 (N815, N800);
and AND3 (N816, N809, N320, N329);
nand NAND4 (N817, N816, N210, N461, N545);
nor NOR3 (N818, N817, N381, N390);
nand NAND4 (N819, N807, N780, N401, N246);
not NOT1 (N820, N805);
xor XOR2 (N821, N819, N403);
buf BUF1 (N822, N821);
nand NAND3 (N823, N793, N636, N77);
nor NOR4 (N824, N814, N13, N515, N442);
xor XOR2 (N825, N820, N499);
nor NOR2 (N826, N815, N16);
xor XOR2 (N827, N812, N670);
nor NOR3 (N828, N813, N152, N22);
buf BUF1 (N829, N818);
nor NOR2 (N830, N811, N70);
and AND3 (N831, N810, N635, N585);
nor NOR3 (N832, N831, N735, N758);
xor XOR2 (N833, N828, N536);
not NOT1 (N834, N825);
nand NAND4 (N835, N832, N547, N523, N46);
or OR4 (N836, N823, N254, N802, N774);
nand NAND4 (N837, N835, N508, N507, N377);
buf BUF1 (N838, N833);
nor NOR3 (N839, N826, N24, N472);
not NOT1 (N840, N837);
and AND2 (N841, N834, N687);
nand NAND2 (N842, N822, N623);
nand NAND3 (N843, N839, N540, N214);
buf BUF1 (N844, N827);
or OR3 (N845, N844, N815, N647);
xor XOR2 (N846, N843, N828);
not NOT1 (N847, N830);
nand NAND4 (N848, N840, N81, N697, N348);
and AND4 (N849, N829, N839, N412, N298);
xor XOR2 (N850, N824, N5);
or OR3 (N851, N845, N772, N401);
and AND3 (N852, N846, N484, N318);
nor NOR3 (N853, N852, N710, N194);
and AND3 (N854, N836, N619, N480);
nand NAND3 (N855, N850, N339, N675);
xor XOR2 (N856, N855, N571);
xor XOR2 (N857, N842, N164);
and AND4 (N858, N849, N645, N832, N698);
xor XOR2 (N859, N854, N108);
nor NOR4 (N860, N851, N577, N22, N484);
or OR4 (N861, N856, N701, N158, N503);
xor XOR2 (N862, N858, N451);
not NOT1 (N863, N847);
nor NOR2 (N864, N857, N760);
nand NAND3 (N865, N838, N61, N433);
buf BUF1 (N866, N860);
xor XOR2 (N867, N848, N710);
and AND3 (N868, N867, N639, N728);
nor NOR2 (N869, N863, N701);
buf BUF1 (N870, N865);
nor NOR4 (N871, N870, N177, N440, N690);
buf BUF1 (N872, N841);
xor XOR2 (N873, N871, N522);
nand NAND3 (N874, N861, N333, N838);
and AND4 (N875, N869, N189, N827, N635);
or OR2 (N876, N853, N335);
nor NOR3 (N877, N866, N758, N868);
not NOT1 (N878, N680);
or OR2 (N879, N859, N222);
buf BUF1 (N880, N872);
and AND2 (N881, N879, N346);
nor NOR3 (N882, N880, N181, N597);
xor XOR2 (N883, N878, N96);
or OR2 (N884, N873, N261);
buf BUF1 (N885, N876);
nor NOR2 (N886, N883, N393);
not NOT1 (N887, N886);
nand NAND4 (N888, N875, N285, N661, N662);
nand NAND4 (N889, N877, N316, N762, N162);
and AND3 (N890, N874, N399, N402);
not NOT1 (N891, N889);
buf BUF1 (N892, N890);
buf BUF1 (N893, N891);
nor NOR3 (N894, N881, N279, N628);
and AND4 (N895, N884, N612, N490, N20);
buf BUF1 (N896, N894);
not NOT1 (N897, N893);
nand NAND2 (N898, N887, N228);
nor NOR3 (N899, N895, N245, N861);
and AND4 (N900, N896, N680, N573, N359);
nor NOR2 (N901, N898, N102);
nand NAND2 (N902, N897, N693);
or OR2 (N903, N862, N592);
nor NOR2 (N904, N864, N440);
not NOT1 (N905, N899);
nand NAND3 (N906, N902, N253, N331);
xor XOR2 (N907, N901, N797);
nand NAND2 (N908, N907, N170);
xor XOR2 (N909, N903, N2);
nand NAND2 (N910, N882, N49);
not NOT1 (N911, N910);
nand NAND3 (N912, N908, N261, N25);
or OR3 (N913, N885, N386, N509);
xor XOR2 (N914, N913, N852);
and AND3 (N915, N904, N295, N731);
xor XOR2 (N916, N914, N82);
xor XOR2 (N917, N912, N114);
buf BUF1 (N918, N892);
nand NAND2 (N919, N900, N78);
nand NAND2 (N920, N918, N609);
xor XOR2 (N921, N888, N836);
xor XOR2 (N922, N915, N429);
xor XOR2 (N923, N917, N543);
or OR2 (N924, N922, N53);
and AND2 (N925, N916, N65);
nor NOR2 (N926, N925, N173);
or OR4 (N927, N926, N1, N347, N339);
nor NOR4 (N928, N920, N71, N413, N411);
buf BUF1 (N929, N906);
buf BUF1 (N930, N911);
xor XOR2 (N931, N919, N622);
buf BUF1 (N932, N931);
nand NAND3 (N933, N909, N177, N522);
nor NOR4 (N934, N923, N725, N211, N538);
buf BUF1 (N935, N928);
not NOT1 (N936, N932);
xor XOR2 (N937, N921, N4);
buf BUF1 (N938, N935);
and AND3 (N939, N937, N104, N309);
and AND2 (N940, N927, N598);
nor NOR3 (N941, N929, N872, N279);
not NOT1 (N942, N905);
or OR3 (N943, N939, N908, N438);
and AND4 (N944, N934, N713, N832, N380);
nor NOR2 (N945, N936, N382);
or OR2 (N946, N943, N132);
nor NOR4 (N947, N946, N237, N31, N597);
not NOT1 (N948, N924);
nand NAND4 (N949, N941, N358, N587, N777);
nor NOR2 (N950, N930, N430);
and AND4 (N951, N942, N178, N416, N815);
nand NAND2 (N952, N945, N460);
nor NOR3 (N953, N951, N82, N879);
not NOT1 (N954, N938);
buf BUF1 (N955, N953);
nor NOR2 (N956, N933, N117);
and AND2 (N957, N940, N736);
or OR2 (N958, N950, N267);
not NOT1 (N959, N955);
and AND3 (N960, N959, N148, N298);
buf BUF1 (N961, N944);
nand NAND2 (N962, N952, N74);
nand NAND2 (N963, N957, N780);
xor XOR2 (N964, N963, N262);
or OR3 (N965, N948, N270, N806);
buf BUF1 (N966, N965);
or OR4 (N967, N947, N834, N466, N395);
buf BUF1 (N968, N958);
not NOT1 (N969, N968);
nor NOR2 (N970, N962, N237);
nand NAND4 (N971, N961, N258, N566, N3);
nand NAND3 (N972, N964, N437, N191);
or OR3 (N973, N967, N4, N594);
or OR4 (N974, N954, N925, N774, N297);
buf BUF1 (N975, N956);
nand NAND4 (N976, N969, N545, N743, N963);
nor NOR4 (N977, N975, N300, N533, N363);
and AND4 (N978, N949, N931, N486, N852);
buf BUF1 (N979, N976);
nand NAND2 (N980, N979, N69);
xor XOR2 (N981, N970, N596);
and AND3 (N982, N977, N967, N770);
nand NAND2 (N983, N974, N692);
nand NAND3 (N984, N978, N474, N931);
or OR4 (N985, N960, N810, N47, N201);
buf BUF1 (N986, N971);
nor NOR2 (N987, N983, N616);
buf BUF1 (N988, N981);
xor XOR2 (N989, N980, N674);
not NOT1 (N990, N987);
nor NOR3 (N991, N972, N270, N531);
nor NOR2 (N992, N991, N332);
nor NOR2 (N993, N982, N864);
buf BUF1 (N994, N986);
or OR4 (N995, N992, N424, N282, N195);
and AND3 (N996, N973, N471, N142);
nand NAND4 (N997, N995, N175, N916, N331);
nor NOR2 (N998, N996, N750);
buf BUF1 (N999, N990);
nand NAND2 (N1000, N998, N184);
nand NAND2 (N1001, N966, N870);
buf BUF1 (N1002, N993);
not NOT1 (N1003, N997);
xor XOR2 (N1004, N989, N883);
nand NAND4 (N1005, N1002, N86, N993, N210);
buf BUF1 (N1006, N984);
buf BUF1 (N1007, N1005);
not NOT1 (N1008, N1000);
not NOT1 (N1009, N985);
buf BUF1 (N1010, N1001);
and AND3 (N1011, N988, N226, N922);
not NOT1 (N1012, N1007);
and AND3 (N1013, N1012, N608, N359);
buf BUF1 (N1014, N1009);
nand NAND4 (N1015, N999, N702, N45, N558);
nand NAND3 (N1016, N1010, N71, N725);
and AND3 (N1017, N1011, N292, N745);
or OR4 (N1018, N1016, N753, N907, N170);
and AND2 (N1019, N1015, N105);
not NOT1 (N1020, N1004);
or OR3 (N1021, N1014, N648, N881);
xor XOR2 (N1022, N1006, N944);
not NOT1 (N1023, N1003);
not NOT1 (N1024, N1013);
nand NAND3 (N1025, N1022, N152, N558);
nor NOR3 (N1026, N1008, N604, N571);
nand NAND2 (N1027, N1025, N750);
nor NOR2 (N1028, N1024, N833);
or OR3 (N1029, N1020, N259, N324);
nand NAND2 (N1030, N1026, N1022);
nor NOR3 (N1031, N1029, N302, N810);
or OR4 (N1032, N1019, N926, N707, N749);
not NOT1 (N1033, N1021);
xor XOR2 (N1034, N1031, N545);
and AND4 (N1035, N1027, N561, N262, N38);
buf BUF1 (N1036, N1017);
buf BUF1 (N1037, N1030);
buf BUF1 (N1038, N1018);
or OR3 (N1039, N1032, N594, N68);
and AND4 (N1040, N1033, N510, N402, N737);
nor NOR2 (N1041, N1028, N535);
or OR2 (N1042, N1034, N949);
nor NOR4 (N1043, N1038, N422, N816, N1024);
nand NAND2 (N1044, N1037, N164);
and AND2 (N1045, N1039, N955);
buf BUF1 (N1046, N1023);
not NOT1 (N1047, N1046);
nand NAND4 (N1048, N1047, N750, N1010, N926);
nand NAND3 (N1049, N1048, N493, N971);
buf BUF1 (N1050, N1042);
nand NAND2 (N1051, N1036, N595);
xor XOR2 (N1052, N1045, N812);
nor NOR2 (N1053, N1049, N329);
buf BUF1 (N1054, N1050);
xor XOR2 (N1055, N1044, N356);
xor XOR2 (N1056, N1040, N365);
nor NOR3 (N1057, N1054, N804, N905);
xor XOR2 (N1058, N1055, N696);
and AND3 (N1059, N994, N952, N688);
xor XOR2 (N1060, N1057, N86);
nor NOR3 (N1061, N1053, N278, N187);
nand NAND4 (N1062, N1043, N162, N1027, N307);
nand NAND2 (N1063, N1056, N633);
nand NAND3 (N1064, N1035, N30, N614);
buf BUF1 (N1065, N1063);
buf BUF1 (N1066, N1064);
buf BUF1 (N1067, N1052);
buf BUF1 (N1068, N1060);
xor XOR2 (N1069, N1067, N1044);
and AND2 (N1070, N1058, N591);
nor NOR3 (N1071, N1068, N575, N589);
or OR2 (N1072, N1069, N598);
nor NOR2 (N1073, N1041, N937);
and AND4 (N1074, N1051, N3, N292, N503);
nor NOR3 (N1075, N1070, N659, N359);
xor XOR2 (N1076, N1065, N163);
buf BUF1 (N1077, N1066);
and AND4 (N1078, N1072, N26, N466, N544);
xor XOR2 (N1079, N1059, N969);
nor NOR4 (N1080, N1077, N989, N997, N481);
nor NOR2 (N1081, N1071, N584);
nor NOR2 (N1082, N1076, N887);
not NOT1 (N1083, N1061);
nor NOR2 (N1084, N1080, N1050);
and AND2 (N1085, N1082, N769);
buf BUF1 (N1086, N1079);
and AND3 (N1087, N1081, N305, N98);
not NOT1 (N1088, N1062);
nor NOR4 (N1089, N1075, N464, N423, N831);
nor NOR3 (N1090, N1088, N949, N212);
not NOT1 (N1091, N1074);
xor XOR2 (N1092, N1078, N671);
nand NAND3 (N1093, N1084, N596, N54);
nand NAND3 (N1094, N1086, N937, N42);
nor NOR4 (N1095, N1085, N810, N109, N764);
nor NOR4 (N1096, N1087, N763, N502, N355);
xor XOR2 (N1097, N1096, N757);
xor XOR2 (N1098, N1095, N789);
buf BUF1 (N1099, N1092);
nor NOR2 (N1100, N1073, N979);
buf BUF1 (N1101, N1094);
or OR2 (N1102, N1091, N63);
not NOT1 (N1103, N1083);
and AND3 (N1104, N1102, N475, N724);
nand NAND3 (N1105, N1099, N100, N188);
xor XOR2 (N1106, N1089, N233);
nand NAND4 (N1107, N1103, N754, N991, N867);
nor NOR2 (N1108, N1105, N529);
or OR2 (N1109, N1097, N372);
buf BUF1 (N1110, N1106);
nor NOR2 (N1111, N1101, N344);
or OR2 (N1112, N1090, N639);
nand NAND2 (N1113, N1112, N2);
nor NOR4 (N1114, N1100, N406, N680, N374);
nor NOR3 (N1115, N1110, N454, N24);
not NOT1 (N1116, N1104);
xor XOR2 (N1117, N1098, N745);
buf BUF1 (N1118, N1109);
or OR2 (N1119, N1111, N791);
xor XOR2 (N1120, N1114, N529);
not NOT1 (N1121, N1113);
buf BUF1 (N1122, N1093);
nand NAND3 (N1123, N1116, N1006, N1098);
xor XOR2 (N1124, N1118, N318);
or OR4 (N1125, N1117, N500, N354, N241);
not NOT1 (N1126, N1125);
and AND4 (N1127, N1123, N1002, N111, N227);
xor XOR2 (N1128, N1124, N346);
xor XOR2 (N1129, N1108, N144);
xor XOR2 (N1130, N1127, N546);
xor XOR2 (N1131, N1122, N403);
xor XOR2 (N1132, N1131, N599);
and AND2 (N1133, N1115, N204);
and AND2 (N1134, N1119, N903);
or OR4 (N1135, N1134, N587, N230, N492);
nor NOR2 (N1136, N1126, N985);
not NOT1 (N1137, N1121);
and AND2 (N1138, N1130, N160);
buf BUF1 (N1139, N1132);
nand NAND4 (N1140, N1137, N54, N117, N380);
and AND3 (N1141, N1139, N10, N246);
nand NAND3 (N1142, N1141, N317, N222);
buf BUF1 (N1143, N1133);
nor NOR3 (N1144, N1143, N1053, N396);
not NOT1 (N1145, N1140);
or OR4 (N1146, N1145, N553, N982, N268);
nand NAND4 (N1147, N1136, N857, N981, N54);
nand NAND3 (N1148, N1135, N1120, N1145);
nor NOR4 (N1149, N587, N265, N1057, N666);
or OR3 (N1150, N1146, N94, N642);
nor NOR2 (N1151, N1150, N546);
and AND3 (N1152, N1128, N608, N55);
or OR4 (N1153, N1147, N1067, N7, N598);
nor NOR3 (N1154, N1107, N477, N664);
not NOT1 (N1155, N1138);
and AND2 (N1156, N1129, N989);
or OR2 (N1157, N1144, N107);
or OR2 (N1158, N1156, N260);
nor NOR3 (N1159, N1155, N164, N907);
and AND4 (N1160, N1158, N609, N781, N501);
and AND2 (N1161, N1159, N539);
not NOT1 (N1162, N1152);
or OR4 (N1163, N1142, N678, N289, N162);
xor XOR2 (N1164, N1153, N1069);
buf BUF1 (N1165, N1154);
xor XOR2 (N1166, N1149, N406);
or OR2 (N1167, N1166, N899);
not NOT1 (N1168, N1161);
nor NOR3 (N1169, N1148, N206, N984);
and AND3 (N1170, N1151, N577, N350);
not NOT1 (N1171, N1157);
and AND3 (N1172, N1170, N269, N386);
or OR4 (N1173, N1164, N666, N946, N32);
xor XOR2 (N1174, N1168, N476);
not NOT1 (N1175, N1172);
or OR4 (N1176, N1163, N1175, N240, N1116);
nor NOR2 (N1177, N772, N740);
and AND4 (N1178, N1174, N829, N540, N300);
not NOT1 (N1179, N1178);
nor NOR4 (N1180, N1179, N868, N258, N147);
buf BUF1 (N1181, N1165);
or OR4 (N1182, N1167, N565, N622, N96);
xor XOR2 (N1183, N1180, N84);
or OR4 (N1184, N1171, N985, N1130, N643);
nand NAND3 (N1185, N1160, N553, N246);
xor XOR2 (N1186, N1162, N844);
or OR3 (N1187, N1177, N682, N129);
or OR4 (N1188, N1182, N387, N132, N357);
nand NAND4 (N1189, N1181, N734, N1027, N858);
or OR3 (N1190, N1176, N300, N776);
nand NAND4 (N1191, N1184, N813, N677, N588);
buf BUF1 (N1192, N1191);
nor NOR4 (N1193, N1189, N685, N634, N669);
or OR4 (N1194, N1193, N996, N996, N31);
and AND4 (N1195, N1194, N27, N565, N144);
buf BUF1 (N1196, N1190);
buf BUF1 (N1197, N1196);
nand NAND3 (N1198, N1192, N596, N1149);
and AND3 (N1199, N1195, N969, N615);
or OR4 (N1200, N1198, N559, N1068, N487);
not NOT1 (N1201, N1200);
or OR3 (N1202, N1187, N668, N1107);
xor XOR2 (N1203, N1197, N461);
xor XOR2 (N1204, N1203, N794);
or OR4 (N1205, N1201, N1089, N1117, N23);
nor NOR4 (N1206, N1205, N264, N164, N505);
not NOT1 (N1207, N1188);
and AND4 (N1208, N1169, N741, N159, N937);
nand NAND2 (N1209, N1199, N318);
nor NOR2 (N1210, N1209, N250);
xor XOR2 (N1211, N1186, N482);
not NOT1 (N1212, N1206);
nand NAND3 (N1213, N1211, N1056, N644);
not NOT1 (N1214, N1173);
xor XOR2 (N1215, N1212, N658);
or OR3 (N1216, N1202, N118, N897);
nor NOR2 (N1217, N1214, N23);
xor XOR2 (N1218, N1215, N618);
xor XOR2 (N1219, N1207, N560);
nand NAND2 (N1220, N1217, N1059);
and AND4 (N1221, N1183, N812, N56, N869);
or OR4 (N1222, N1220, N74, N554, N84);
or OR4 (N1223, N1218, N66, N697, N158);
not NOT1 (N1224, N1208);
nand NAND3 (N1225, N1216, N274, N793);
nor NOR4 (N1226, N1219, N584, N336, N380);
buf BUF1 (N1227, N1221);
buf BUF1 (N1228, N1222);
nor NOR3 (N1229, N1210, N1125, N982);
nand NAND3 (N1230, N1226, N354, N816);
nand NAND2 (N1231, N1227, N891);
not NOT1 (N1232, N1213);
and AND4 (N1233, N1229, N417, N972, N1207);
not NOT1 (N1234, N1228);
nand NAND2 (N1235, N1231, N865);
nor NOR2 (N1236, N1233, N1189);
buf BUF1 (N1237, N1225);
and AND4 (N1238, N1236, N1188, N800, N450);
or OR2 (N1239, N1234, N494);
nand NAND3 (N1240, N1224, N622, N468);
not NOT1 (N1241, N1239);
and AND4 (N1242, N1185, N375, N35, N74);
and AND3 (N1243, N1241, N503, N413);
and AND4 (N1244, N1243, N455, N80, N1227);
not NOT1 (N1245, N1244);
and AND4 (N1246, N1238, N212, N426, N320);
not NOT1 (N1247, N1240);
xor XOR2 (N1248, N1246, N650);
buf BUF1 (N1249, N1204);
and AND4 (N1250, N1235, N973, N1180, N261);
not NOT1 (N1251, N1245);
and AND4 (N1252, N1247, N451, N748, N498);
xor XOR2 (N1253, N1230, N759);
or OR4 (N1254, N1252, N1125, N1203, N456);
nand NAND3 (N1255, N1223, N249, N323);
buf BUF1 (N1256, N1253);
or OR3 (N1257, N1254, N473, N62);
or OR4 (N1258, N1248, N1253, N907, N261);
xor XOR2 (N1259, N1258, N852);
xor XOR2 (N1260, N1255, N487);
nor NOR2 (N1261, N1256, N1007);
nand NAND4 (N1262, N1251, N1244, N489, N102);
or OR3 (N1263, N1242, N532, N1132);
and AND2 (N1264, N1250, N210);
and AND4 (N1265, N1263, N951, N1076, N992);
buf BUF1 (N1266, N1265);
xor XOR2 (N1267, N1262, N886);
and AND4 (N1268, N1232, N731, N1094, N191);
nor NOR2 (N1269, N1259, N561);
nand NAND2 (N1270, N1268, N543);
nor NOR3 (N1271, N1266, N1101, N603);
nand NAND4 (N1272, N1267, N866, N758, N225);
or OR4 (N1273, N1261, N299, N245, N336);
nand NAND2 (N1274, N1249, N1258);
or OR3 (N1275, N1272, N444, N189);
not NOT1 (N1276, N1271);
not NOT1 (N1277, N1269);
xor XOR2 (N1278, N1270, N731);
buf BUF1 (N1279, N1278);
xor XOR2 (N1280, N1273, N503);
nand NAND2 (N1281, N1275, N49);
or OR4 (N1282, N1280, N402, N1122, N318);
xor XOR2 (N1283, N1282, N805);
or OR4 (N1284, N1264, N872, N277, N1132);
not NOT1 (N1285, N1260);
and AND3 (N1286, N1279, N1252, N726);
nor NOR3 (N1287, N1257, N422, N1103);
xor XOR2 (N1288, N1284, N1183);
buf BUF1 (N1289, N1276);
not NOT1 (N1290, N1237);
and AND4 (N1291, N1285, N792, N735, N218);
not NOT1 (N1292, N1289);
nand NAND3 (N1293, N1286, N1020, N181);
not NOT1 (N1294, N1290);
or OR4 (N1295, N1283, N1081, N395, N1019);
and AND2 (N1296, N1277, N594);
nor NOR2 (N1297, N1281, N1043);
or OR4 (N1298, N1294, N330, N1281, N212);
nand NAND4 (N1299, N1288, N4, N798, N539);
xor XOR2 (N1300, N1287, N339);
and AND3 (N1301, N1292, N965, N1109);
buf BUF1 (N1302, N1274);
not NOT1 (N1303, N1293);
not NOT1 (N1304, N1291);
nor NOR2 (N1305, N1299, N1256);
xor XOR2 (N1306, N1295, N1234);
buf BUF1 (N1307, N1300);
nor NOR3 (N1308, N1298, N70, N1191);
xor XOR2 (N1309, N1307, N790);
or OR4 (N1310, N1301, N542, N446, N628);
or OR2 (N1311, N1310, N832);
nand NAND3 (N1312, N1297, N607, N346);
not NOT1 (N1313, N1304);
and AND4 (N1314, N1313, N1300, N658, N483);
not NOT1 (N1315, N1312);
buf BUF1 (N1316, N1303);
xor XOR2 (N1317, N1315, N1054);
nor NOR3 (N1318, N1309, N971, N451);
nor NOR4 (N1319, N1316, N677, N1181, N1218);
buf BUF1 (N1320, N1305);
nor NOR2 (N1321, N1296, N1185);
buf BUF1 (N1322, N1321);
nor NOR4 (N1323, N1311, N263, N109, N874);
nor NOR2 (N1324, N1320, N204);
not NOT1 (N1325, N1318);
and AND2 (N1326, N1308, N691);
and AND3 (N1327, N1302, N1267, N462);
nor NOR4 (N1328, N1323, N944, N238, N312);
xor XOR2 (N1329, N1306, N1141);
buf BUF1 (N1330, N1317);
not NOT1 (N1331, N1324);
and AND4 (N1332, N1319, N1246, N476, N21);
not NOT1 (N1333, N1327);
nor NOR2 (N1334, N1328, N127);
not NOT1 (N1335, N1332);
xor XOR2 (N1336, N1314, N758);
nand NAND3 (N1337, N1336, N230, N469);
buf BUF1 (N1338, N1335);
nand NAND4 (N1339, N1331, N648, N526, N822);
or OR3 (N1340, N1337, N779, N309);
nor NOR3 (N1341, N1333, N1153, N538);
nor NOR2 (N1342, N1339, N705);
not NOT1 (N1343, N1340);
not NOT1 (N1344, N1325);
nand NAND4 (N1345, N1322, N647, N1075, N131);
nor NOR2 (N1346, N1341, N708);
and AND3 (N1347, N1345, N920, N368);
nand NAND2 (N1348, N1346, N607);
nand NAND4 (N1349, N1330, N653, N244, N991);
and AND4 (N1350, N1349, N475, N502, N555);
xor XOR2 (N1351, N1326, N881);
not NOT1 (N1352, N1351);
or OR4 (N1353, N1350, N95, N1164, N79);
xor XOR2 (N1354, N1342, N928);
and AND2 (N1355, N1329, N996);
buf BUF1 (N1356, N1355);
and AND4 (N1357, N1352, N549, N450, N536);
xor XOR2 (N1358, N1334, N1328);
buf BUF1 (N1359, N1347);
not NOT1 (N1360, N1359);
nor NOR3 (N1361, N1356, N967, N587);
buf BUF1 (N1362, N1357);
nor NOR3 (N1363, N1353, N39, N1312);
xor XOR2 (N1364, N1362, N297);
not NOT1 (N1365, N1363);
buf BUF1 (N1366, N1343);
nor NOR3 (N1367, N1338, N1249, N757);
and AND2 (N1368, N1354, N991);
nor NOR3 (N1369, N1367, N1274, N720);
and AND4 (N1370, N1365, N673, N736, N1090);
or OR3 (N1371, N1344, N333, N95);
not NOT1 (N1372, N1371);
not NOT1 (N1373, N1368);
or OR4 (N1374, N1358, N511, N983, N822);
xor XOR2 (N1375, N1348, N602);
xor XOR2 (N1376, N1372, N1067);
nand NAND4 (N1377, N1360, N26, N1369, N285);
buf BUF1 (N1378, N805);
nand NAND3 (N1379, N1376, N1338, N1166);
and AND4 (N1380, N1377, N1007, N752, N268);
nand NAND2 (N1381, N1378, N12);
and AND4 (N1382, N1374, N1044, N346, N946);
not NOT1 (N1383, N1375);
buf BUF1 (N1384, N1380);
buf BUF1 (N1385, N1383);
xor XOR2 (N1386, N1385, N1337);
buf BUF1 (N1387, N1373);
and AND3 (N1388, N1384, N539, N485);
buf BUF1 (N1389, N1387);
nand NAND2 (N1390, N1370, N1065);
nand NAND4 (N1391, N1382, N657, N652, N1193);
not NOT1 (N1392, N1386);
or OR2 (N1393, N1388, N84);
not NOT1 (N1394, N1393);
and AND3 (N1395, N1379, N471, N462);
buf BUF1 (N1396, N1361);
nor NOR4 (N1397, N1396, N960, N911, N875);
not NOT1 (N1398, N1364);
buf BUF1 (N1399, N1392);
and AND4 (N1400, N1395, N535, N322, N693);
not NOT1 (N1401, N1398);
and AND4 (N1402, N1394, N1122, N721, N1013);
or OR3 (N1403, N1397, N778, N295);
xor XOR2 (N1404, N1366, N1052);
nor NOR2 (N1405, N1404, N109);
or OR3 (N1406, N1389, N381, N676);
xor XOR2 (N1407, N1401, N1344);
or OR3 (N1408, N1406, N1111, N1282);
nor NOR3 (N1409, N1408, N364, N1180);
nor NOR2 (N1410, N1402, N1130);
xor XOR2 (N1411, N1405, N32);
and AND3 (N1412, N1399, N1399, N552);
and AND3 (N1413, N1412, N537, N1165);
xor XOR2 (N1414, N1410, N548);
or OR4 (N1415, N1409, N643, N774, N621);
buf BUF1 (N1416, N1411);
and AND3 (N1417, N1400, N44, N650);
nor NOR4 (N1418, N1390, N277, N1148, N765);
and AND3 (N1419, N1415, N1144, N822);
not NOT1 (N1420, N1413);
nand NAND2 (N1421, N1420, N1352);
not NOT1 (N1422, N1416);
xor XOR2 (N1423, N1381, N410);
nand NAND3 (N1424, N1423, N283, N1199);
or OR3 (N1425, N1417, N853, N789);
or OR2 (N1426, N1407, N769);
xor XOR2 (N1427, N1421, N1375);
and AND4 (N1428, N1424, N594, N180, N1178);
xor XOR2 (N1429, N1427, N260);
buf BUF1 (N1430, N1425);
or OR2 (N1431, N1426, N534);
and AND3 (N1432, N1431, N181, N1411);
buf BUF1 (N1433, N1432);
and AND2 (N1434, N1429, N292);
nor NOR4 (N1435, N1403, N1295, N1156, N588);
nor NOR4 (N1436, N1428, N1308, N90, N866);
nand NAND2 (N1437, N1422, N1039);
xor XOR2 (N1438, N1437, N511);
not NOT1 (N1439, N1436);
and AND4 (N1440, N1418, N1416, N929, N400);
xor XOR2 (N1441, N1419, N56);
nand NAND2 (N1442, N1438, N790);
and AND2 (N1443, N1439, N191);
xor XOR2 (N1444, N1441, N653);
and AND2 (N1445, N1440, N347);
not NOT1 (N1446, N1430);
not NOT1 (N1447, N1442);
not NOT1 (N1448, N1443);
not NOT1 (N1449, N1414);
not NOT1 (N1450, N1444);
not NOT1 (N1451, N1450);
nand NAND3 (N1452, N1446, N118, N675);
or OR4 (N1453, N1452, N1333, N133, N57);
nand NAND2 (N1454, N1451, N95);
nand NAND4 (N1455, N1433, N395, N1330, N647);
nor NOR3 (N1456, N1445, N486, N1374);
nand NAND3 (N1457, N1449, N1407, N1375);
and AND4 (N1458, N1447, N504, N1000, N23);
and AND4 (N1459, N1457, N1073, N427, N9);
or OR3 (N1460, N1458, N1355, N1148);
xor XOR2 (N1461, N1448, N81);
xor XOR2 (N1462, N1391, N125);
and AND4 (N1463, N1453, N380, N376, N1031);
not NOT1 (N1464, N1463);
not NOT1 (N1465, N1434);
nor NOR3 (N1466, N1464, N1253, N933);
nand NAND2 (N1467, N1461, N631);
xor XOR2 (N1468, N1462, N156);
xor XOR2 (N1469, N1466, N302);
nand NAND4 (N1470, N1468, N1175, N1347, N1040);
and AND2 (N1471, N1435, N783);
nor NOR4 (N1472, N1470, N347, N661, N929);
not NOT1 (N1473, N1471);
buf BUF1 (N1474, N1467);
not NOT1 (N1475, N1465);
not NOT1 (N1476, N1456);
buf BUF1 (N1477, N1469);
and AND2 (N1478, N1474, N630);
nor NOR3 (N1479, N1459, N605, N1006);
buf BUF1 (N1480, N1476);
not NOT1 (N1481, N1480);
not NOT1 (N1482, N1473);
not NOT1 (N1483, N1482);
not NOT1 (N1484, N1454);
and AND2 (N1485, N1483, N102);
nor NOR2 (N1486, N1478, N541);
nand NAND4 (N1487, N1455, N419, N318, N1463);
nand NAND4 (N1488, N1477, N1160, N1356, N486);
buf BUF1 (N1489, N1487);
or OR3 (N1490, N1489, N1259, N407);
xor XOR2 (N1491, N1488, N227);
not NOT1 (N1492, N1486);
and AND3 (N1493, N1460, N614, N385);
xor XOR2 (N1494, N1490, N1045);
xor XOR2 (N1495, N1485, N100);
or OR2 (N1496, N1481, N854);
nor NOR3 (N1497, N1491, N1099, N1475);
not NOT1 (N1498, N1481);
nand NAND4 (N1499, N1496, N1293, N135, N1084);
or OR3 (N1500, N1493, N736, N1045);
not NOT1 (N1501, N1484);
xor XOR2 (N1502, N1494, N325);
and AND2 (N1503, N1501, N125);
xor XOR2 (N1504, N1500, N782);
nand NAND2 (N1505, N1499, N312);
or OR2 (N1506, N1502, N645);
not NOT1 (N1507, N1492);
not NOT1 (N1508, N1504);
nand NAND3 (N1509, N1505, N187, N621);
and AND2 (N1510, N1506, N1008);
or OR4 (N1511, N1479, N349, N1418, N147);
xor XOR2 (N1512, N1511, N1301);
xor XOR2 (N1513, N1512, N979);
buf BUF1 (N1514, N1497);
xor XOR2 (N1515, N1509, N1321);
or OR4 (N1516, N1514, N1466, N1151, N1443);
nor NOR4 (N1517, N1503, N1453, N1316, N365);
or OR4 (N1518, N1517, N1081, N536, N564);
nor NOR3 (N1519, N1498, N130, N197);
nand NAND3 (N1520, N1507, N1304, N627);
and AND4 (N1521, N1520, N606, N22, N566);
and AND2 (N1522, N1510, N1266);
not NOT1 (N1523, N1508);
xor XOR2 (N1524, N1513, N76);
buf BUF1 (N1525, N1472);
nand NAND2 (N1526, N1515, N541);
nor NOR3 (N1527, N1526, N1090, N273);
or OR4 (N1528, N1516, N831, N89, N1389);
nand NAND2 (N1529, N1523, N643);
buf BUF1 (N1530, N1521);
xor XOR2 (N1531, N1530, N1195);
and AND4 (N1532, N1518, N403, N1397, N29);
nand NAND4 (N1533, N1495, N1459, N1006, N2);
nand NAND4 (N1534, N1519, N93, N666, N54);
or OR3 (N1535, N1522, N1104, N807);
and AND2 (N1536, N1528, N1493);
or OR3 (N1537, N1535, N457, N499);
buf BUF1 (N1538, N1524);
nor NOR3 (N1539, N1527, N404, N396);
not NOT1 (N1540, N1525);
xor XOR2 (N1541, N1533, N1008);
and AND4 (N1542, N1541, N1453, N134, N278);
buf BUF1 (N1543, N1539);
not NOT1 (N1544, N1529);
and AND3 (N1545, N1542, N676, N382);
or OR3 (N1546, N1531, N1236, N771);
nand NAND4 (N1547, N1546, N558, N109, N1320);
buf BUF1 (N1548, N1537);
or OR2 (N1549, N1548, N857);
xor XOR2 (N1550, N1532, N1223);
and AND2 (N1551, N1550, N1414);
and AND2 (N1552, N1549, N1227);
and AND3 (N1553, N1543, N195, N503);
xor XOR2 (N1554, N1534, N1283);
xor XOR2 (N1555, N1536, N1265);
nor NOR4 (N1556, N1554, N183, N944, N412);
nor NOR2 (N1557, N1547, N1177);
not NOT1 (N1558, N1538);
not NOT1 (N1559, N1552);
buf BUF1 (N1560, N1557);
and AND2 (N1561, N1540, N809);
and AND4 (N1562, N1553, N928, N1129, N1392);
nor NOR4 (N1563, N1559, N542, N35, N856);
buf BUF1 (N1564, N1562);
xor XOR2 (N1565, N1561, N426);
and AND3 (N1566, N1544, N343, N240);
xor XOR2 (N1567, N1560, N1508);
or OR3 (N1568, N1551, N678, N75);
not NOT1 (N1569, N1555);
nor NOR4 (N1570, N1568, N1202, N1299, N102);
not NOT1 (N1571, N1566);
not NOT1 (N1572, N1556);
or OR2 (N1573, N1572, N993);
or OR2 (N1574, N1573, N931);
not NOT1 (N1575, N1569);
nand NAND2 (N1576, N1575, N479);
not NOT1 (N1577, N1558);
or OR2 (N1578, N1570, N1224);
nor NOR4 (N1579, N1545, N1276, N1236, N20);
not NOT1 (N1580, N1564);
or OR4 (N1581, N1580, N437, N206, N1443);
xor XOR2 (N1582, N1578, N1049);
or OR2 (N1583, N1563, N352);
nand NAND2 (N1584, N1577, N278);
xor XOR2 (N1585, N1571, N1542);
buf BUF1 (N1586, N1583);
nand NAND2 (N1587, N1565, N1241);
buf BUF1 (N1588, N1586);
xor XOR2 (N1589, N1567, N469);
xor XOR2 (N1590, N1585, N736);
buf BUF1 (N1591, N1579);
buf BUF1 (N1592, N1588);
buf BUF1 (N1593, N1582);
xor XOR2 (N1594, N1590, N874);
buf BUF1 (N1595, N1576);
nor NOR4 (N1596, N1584, N635, N1180, N131);
xor XOR2 (N1597, N1594, N563);
nand NAND3 (N1598, N1587, N1018, N577);
and AND2 (N1599, N1597, N183);
nand NAND3 (N1600, N1599, N827, N864);
not NOT1 (N1601, N1600);
nor NOR2 (N1602, N1596, N530);
and AND3 (N1603, N1598, N519, N202);
xor XOR2 (N1604, N1589, N1286);
not NOT1 (N1605, N1593);
xor XOR2 (N1606, N1602, N1165);
or OR2 (N1607, N1605, N273);
buf BUF1 (N1608, N1601);
nand NAND2 (N1609, N1574, N1445);
and AND3 (N1610, N1606, N481, N552);
and AND3 (N1611, N1609, N1268, N687);
not NOT1 (N1612, N1591);
buf BUF1 (N1613, N1604);
and AND2 (N1614, N1608, N1121);
buf BUF1 (N1615, N1611);
xor XOR2 (N1616, N1592, N1585);
xor XOR2 (N1617, N1616, N566);
nor NOR3 (N1618, N1607, N468, N368);
nand NAND3 (N1619, N1617, N626, N1228);
nand NAND4 (N1620, N1610, N1311, N955, N1499);
nor NOR4 (N1621, N1613, N345, N189, N192);
nand NAND2 (N1622, N1621, N464);
xor XOR2 (N1623, N1581, N1129);
buf BUF1 (N1624, N1618);
buf BUF1 (N1625, N1620);
not NOT1 (N1626, N1623);
nand NAND4 (N1627, N1595, N1571, N1589, N1255);
or OR2 (N1628, N1622, N673);
nand NAND2 (N1629, N1614, N541);
or OR2 (N1630, N1619, N1076);
xor XOR2 (N1631, N1627, N1474);
buf BUF1 (N1632, N1630);
nand NAND2 (N1633, N1603, N116);
nand NAND4 (N1634, N1626, N1357, N72, N58);
nor NOR2 (N1635, N1612, N984);
xor XOR2 (N1636, N1615, N1565);
buf BUF1 (N1637, N1629);
not NOT1 (N1638, N1625);
and AND4 (N1639, N1634, N1219, N1405, N811);
nand NAND3 (N1640, N1638, N1081, N203);
and AND2 (N1641, N1635, N1012);
nand NAND3 (N1642, N1636, N642, N185);
not NOT1 (N1643, N1640);
nand NAND4 (N1644, N1642, N374, N943, N943);
nand NAND4 (N1645, N1639, N274, N477, N1036);
and AND2 (N1646, N1624, N1105);
buf BUF1 (N1647, N1631);
buf BUF1 (N1648, N1641);
or OR3 (N1649, N1646, N1523, N312);
xor XOR2 (N1650, N1633, N178);
not NOT1 (N1651, N1648);
and AND2 (N1652, N1645, N273);
nand NAND3 (N1653, N1643, N1429, N908);
xor XOR2 (N1654, N1637, N320);
nor NOR4 (N1655, N1653, N381, N842, N1606);
xor XOR2 (N1656, N1650, N810);
not NOT1 (N1657, N1651);
buf BUF1 (N1658, N1647);
or OR3 (N1659, N1655, N1489, N105);
or OR4 (N1660, N1657, N909, N1365, N792);
not NOT1 (N1661, N1628);
buf BUF1 (N1662, N1644);
and AND2 (N1663, N1661, N326);
or OR3 (N1664, N1660, N1112, N1058);
or OR2 (N1665, N1649, N1237);
nor NOR4 (N1666, N1662, N35, N493, N1135);
buf BUF1 (N1667, N1659);
or OR2 (N1668, N1666, N501);
not NOT1 (N1669, N1632);
and AND2 (N1670, N1669, N1165);
buf BUF1 (N1671, N1664);
or OR2 (N1672, N1658, N700);
and AND2 (N1673, N1654, N1273);
and AND2 (N1674, N1652, N279);
nor NOR4 (N1675, N1663, N55, N1542, N85);
not NOT1 (N1676, N1665);
buf BUF1 (N1677, N1673);
not NOT1 (N1678, N1656);
nand NAND2 (N1679, N1677, N229);
and AND3 (N1680, N1674, N508, N335);
and AND2 (N1681, N1668, N693);
nand NAND3 (N1682, N1667, N206, N660);
nand NAND4 (N1683, N1676, N342, N1162, N1038);
nand NAND2 (N1684, N1680, N1062);
xor XOR2 (N1685, N1675, N437);
or OR4 (N1686, N1679, N1032, N978, N44);
xor XOR2 (N1687, N1678, N867);
or OR4 (N1688, N1670, N1158, N1161, N1679);
buf BUF1 (N1689, N1684);
not NOT1 (N1690, N1683);
or OR4 (N1691, N1682, N259, N1109, N1274);
nor NOR4 (N1692, N1691, N1183, N769, N1021);
buf BUF1 (N1693, N1687);
xor XOR2 (N1694, N1686, N283);
buf BUF1 (N1695, N1681);
and AND3 (N1696, N1671, N1689, N279);
nand NAND2 (N1697, N1501, N125);
nor NOR2 (N1698, N1685, N1300);
xor XOR2 (N1699, N1696, N464);
and AND4 (N1700, N1688, N779, N559, N852);
not NOT1 (N1701, N1690);
nand NAND3 (N1702, N1694, N35, N1158);
or OR2 (N1703, N1672, N191);
xor XOR2 (N1704, N1701, N386);
buf BUF1 (N1705, N1698);
nor NOR2 (N1706, N1702, N1066);
and AND2 (N1707, N1703, N1498);
xor XOR2 (N1708, N1693, N1474);
not NOT1 (N1709, N1708);
nand NAND3 (N1710, N1692, N1455, N443);
nor NOR2 (N1711, N1699, N694);
or OR2 (N1712, N1695, N168);
not NOT1 (N1713, N1711);
or OR3 (N1714, N1710, N962, N1207);
or OR4 (N1715, N1704, N166, N159, N46);
xor XOR2 (N1716, N1707, N480);
xor XOR2 (N1717, N1716, N781);
not NOT1 (N1718, N1697);
not NOT1 (N1719, N1714);
nor NOR2 (N1720, N1709, N591);
xor XOR2 (N1721, N1720, N297);
not NOT1 (N1722, N1700);
buf BUF1 (N1723, N1719);
buf BUF1 (N1724, N1717);
and AND3 (N1725, N1713, N885, N57);
and AND4 (N1726, N1706, N1612, N425, N1708);
buf BUF1 (N1727, N1723);
nand NAND4 (N1728, N1721, N533, N1386, N526);
nor NOR3 (N1729, N1726, N1390, N956);
xor XOR2 (N1730, N1729, N42);
and AND2 (N1731, N1727, N1562);
buf BUF1 (N1732, N1712);
not NOT1 (N1733, N1722);
and AND3 (N1734, N1730, N1426, N1533);
nor NOR4 (N1735, N1731, N81, N719, N936);
or OR2 (N1736, N1734, N1313);
nor NOR4 (N1737, N1732, N36, N641, N1349);
or OR2 (N1738, N1733, N718);
buf BUF1 (N1739, N1718);
not NOT1 (N1740, N1739);
nor NOR4 (N1741, N1736, N1241, N1556, N633);
and AND4 (N1742, N1715, N219, N419, N986);
nor NOR2 (N1743, N1740, N598);
nor NOR3 (N1744, N1735, N1655, N396);
nor NOR4 (N1745, N1742, N928, N1250, N589);
xor XOR2 (N1746, N1744, N410);
nor NOR2 (N1747, N1724, N1185);
nand NAND3 (N1748, N1746, N1722, N806);
and AND4 (N1749, N1705, N1434, N702, N680);
or OR3 (N1750, N1728, N1107, N634);
nand NAND4 (N1751, N1743, N458, N1139, N465);
not NOT1 (N1752, N1725);
nand NAND3 (N1753, N1741, N80, N1700);
xor XOR2 (N1754, N1751, N295);
buf BUF1 (N1755, N1752);
xor XOR2 (N1756, N1747, N1390);
nor NOR3 (N1757, N1749, N921, N342);
not NOT1 (N1758, N1737);
or OR4 (N1759, N1745, N143, N1422, N1429);
nor NOR3 (N1760, N1738, N1570, N617);
xor XOR2 (N1761, N1753, N929);
or OR2 (N1762, N1750, N476);
or OR2 (N1763, N1758, N751);
nand NAND4 (N1764, N1760, N1077, N1478, N1288);
not NOT1 (N1765, N1761);
not NOT1 (N1766, N1764);
not NOT1 (N1767, N1757);
nor NOR2 (N1768, N1766, N932);
not NOT1 (N1769, N1767);
xor XOR2 (N1770, N1769, N870);
nor NOR3 (N1771, N1755, N779, N759);
nand NAND3 (N1772, N1771, N1067, N1588);
nor NOR4 (N1773, N1772, N611, N913, N45);
buf BUF1 (N1774, N1770);
not NOT1 (N1775, N1765);
nand NAND3 (N1776, N1756, N1664, N1314);
buf BUF1 (N1777, N1776);
or OR4 (N1778, N1775, N1203, N298, N1297);
nor NOR3 (N1779, N1777, N1628, N858);
nand NAND2 (N1780, N1748, N1568);
not NOT1 (N1781, N1774);
xor XOR2 (N1782, N1754, N603);
nor NOR3 (N1783, N1781, N1715, N298);
xor XOR2 (N1784, N1779, N1753);
not NOT1 (N1785, N1768);
not NOT1 (N1786, N1778);
or OR3 (N1787, N1762, N1016, N726);
and AND4 (N1788, N1785, N1002, N938, N866);
not NOT1 (N1789, N1759);
and AND4 (N1790, N1787, N947, N914, N1215);
or OR3 (N1791, N1780, N485, N150);
nor NOR4 (N1792, N1773, N1447, N383, N277);
and AND3 (N1793, N1782, N926, N1546);
nand NAND2 (N1794, N1788, N137);
buf BUF1 (N1795, N1790);
xor XOR2 (N1796, N1784, N1742);
buf BUF1 (N1797, N1793);
not NOT1 (N1798, N1794);
not NOT1 (N1799, N1795);
or OR2 (N1800, N1763, N682);
or OR4 (N1801, N1797, N670, N480, N406);
nor NOR3 (N1802, N1791, N1067, N1089);
nand NAND3 (N1803, N1786, N1375, N935);
or OR2 (N1804, N1799, N1489);
or OR3 (N1805, N1804, N251, N1272);
and AND4 (N1806, N1789, N970, N483, N587);
and AND3 (N1807, N1798, N1639, N618);
not NOT1 (N1808, N1800);
not NOT1 (N1809, N1796);
nor NOR3 (N1810, N1807, N1268, N1277);
nor NOR2 (N1811, N1805, N937);
buf BUF1 (N1812, N1802);
not NOT1 (N1813, N1801);
and AND3 (N1814, N1792, N1722, N483);
and AND3 (N1815, N1811, N1260, N1558);
or OR4 (N1816, N1783, N1749, N860, N1539);
xor XOR2 (N1817, N1808, N534);
or OR2 (N1818, N1806, N170);
not NOT1 (N1819, N1812);
nor NOR4 (N1820, N1810, N1637, N218, N798);
nand NAND3 (N1821, N1809, N537, N298);
nand NAND4 (N1822, N1817, N184, N1728, N1424);
nor NOR2 (N1823, N1814, N1569);
not NOT1 (N1824, N1813);
xor XOR2 (N1825, N1823, N785);
buf BUF1 (N1826, N1815);
and AND4 (N1827, N1825, N1441, N400, N214);
xor XOR2 (N1828, N1803, N105);
xor XOR2 (N1829, N1816, N8);
and AND2 (N1830, N1818, N678);
not NOT1 (N1831, N1819);
and AND2 (N1832, N1820, N703);
or OR3 (N1833, N1828, N615, N56);
not NOT1 (N1834, N1826);
buf BUF1 (N1835, N1821);
nand NAND4 (N1836, N1833, N897, N1543, N1272);
and AND2 (N1837, N1827, N294);
nand NAND2 (N1838, N1830, N922);
nor NOR2 (N1839, N1838, N86);
not NOT1 (N1840, N1831);
or OR4 (N1841, N1835, N1332, N1047, N1830);
not NOT1 (N1842, N1837);
xor XOR2 (N1843, N1832, N950);
buf BUF1 (N1844, N1829);
and AND2 (N1845, N1836, N940);
buf BUF1 (N1846, N1840);
and AND4 (N1847, N1846, N1016, N44, N1771);
not NOT1 (N1848, N1845);
and AND4 (N1849, N1848, N237, N1461, N574);
not NOT1 (N1850, N1843);
xor XOR2 (N1851, N1850, N834);
xor XOR2 (N1852, N1839, N213);
not NOT1 (N1853, N1822);
buf BUF1 (N1854, N1842);
and AND4 (N1855, N1849, N692, N316, N1692);
or OR2 (N1856, N1853, N1555);
nor NOR3 (N1857, N1841, N510, N1769);
buf BUF1 (N1858, N1824);
and AND4 (N1859, N1844, N284, N837, N803);
or OR4 (N1860, N1857, N1124, N910, N165);
or OR4 (N1861, N1851, N1479, N536, N425);
nand NAND2 (N1862, N1860, N1543);
nand NAND4 (N1863, N1856, N1384, N739, N88);
nor NOR2 (N1864, N1852, N457);
buf BUF1 (N1865, N1864);
and AND2 (N1866, N1854, N246);
not NOT1 (N1867, N1834);
not NOT1 (N1868, N1847);
buf BUF1 (N1869, N1865);
xor XOR2 (N1870, N1863, N1693);
buf BUF1 (N1871, N1868);
and AND3 (N1872, N1870, N1497, N837);
and AND2 (N1873, N1872, N149);
nor NOR2 (N1874, N1871, N828);
or OR4 (N1875, N1866, N768, N1054, N938);
not NOT1 (N1876, N1859);
buf BUF1 (N1877, N1873);
nor NOR4 (N1878, N1874, N1452, N656, N948);
nor NOR4 (N1879, N1878, N43, N1070, N1525);
not NOT1 (N1880, N1858);
or OR4 (N1881, N1879, N448, N1253, N171);
nand NAND4 (N1882, N1867, N865, N1492, N1093);
and AND4 (N1883, N1869, N1692, N1735, N1156);
xor XOR2 (N1884, N1882, N945);
or OR3 (N1885, N1881, N252, N1799);
buf BUF1 (N1886, N1875);
nand NAND4 (N1887, N1883, N812, N1770, N1135);
xor XOR2 (N1888, N1877, N1321);
or OR3 (N1889, N1861, N990, N794);
buf BUF1 (N1890, N1885);
buf BUF1 (N1891, N1888);
buf BUF1 (N1892, N1876);
nand NAND3 (N1893, N1862, N1277, N758);
xor XOR2 (N1894, N1890, N550);
buf BUF1 (N1895, N1889);
not NOT1 (N1896, N1887);
nor NOR4 (N1897, N1896, N1467, N443, N146);
nand NAND4 (N1898, N1897, N19, N721, N1719);
not NOT1 (N1899, N1894);
xor XOR2 (N1900, N1891, N318);
and AND4 (N1901, N1880, N198, N1091, N960);
and AND4 (N1902, N1884, N185, N1838, N1348);
nand NAND2 (N1903, N1900, N425);
xor XOR2 (N1904, N1855, N297);
nor NOR2 (N1905, N1892, N279);
not NOT1 (N1906, N1886);
nand NAND4 (N1907, N1906, N846, N1439, N1539);
nand NAND3 (N1908, N1899, N1774, N497);
not NOT1 (N1909, N1901);
or OR4 (N1910, N1908, N532, N215, N546);
not NOT1 (N1911, N1893);
buf BUF1 (N1912, N1903);
xor XOR2 (N1913, N1912, N1738);
buf BUF1 (N1914, N1909);
and AND3 (N1915, N1907, N53, N1209);
nand NAND3 (N1916, N1913, N1315, N945);
nand NAND2 (N1917, N1898, N1730);
buf BUF1 (N1918, N1915);
not NOT1 (N1919, N1918);
nand NAND2 (N1920, N1895, N592);
nand NAND2 (N1921, N1916, N696);
or OR2 (N1922, N1902, N599);
nand NAND4 (N1923, N1917, N1743, N623, N72);
and AND2 (N1924, N1911, N1048);
and AND3 (N1925, N1919, N1170, N1616);
or OR3 (N1926, N1923, N442, N1781);
nand NAND4 (N1927, N1905, N904, N1156, N1673);
nor NOR4 (N1928, N1920, N60, N601, N1622);
not NOT1 (N1929, N1921);
not NOT1 (N1930, N1925);
not NOT1 (N1931, N1926);
buf BUF1 (N1932, N1927);
nand NAND3 (N1933, N1924, N686, N1042);
xor XOR2 (N1934, N1929, N1245);
buf BUF1 (N1935, N1910);
xor XOR2 (N1936, N1930, N1228);
and AND3 (N1937, N1936, N937, N616);
nor NOR4 (N1938, N1914, N123, N1596, N476);
not NOT1 (N1939, N1938);
xor XOR2 (N1940, N1931, N1735);
or OR2 (N1941, N1935, N1139);
and AND4 (N1942, N1939, N1468, N250, N441);
buf BUF1 (N1943, N1922);
nand NAND2 (N1944, N1941, N1776);
and AND2 (N1945, N1934, N1649);
buf BUF1 (N1946, N1942);
xor XOR2 (N1947, N1945, N763);
and AND4 (N1948, N1928, N130, N344, N759);
not NOT1 (N1949, N1943);
not NOT1 (N1950, N1904);
buf BUF1 (N1951, N1947);
or OR2 (N1952, N1950, N1702);
nor NOR2 (N1953, N1940, N1579);
not NOT1 (N1954, N1932);
nand NAND4 (N1955, N1954, N1152, N1025, N368);
buf BUF1 (N1956, N1937);
nor NOR3 (N1957, N1948, N965, N1777);
buf BUF1 (N1958, N1933);
and AND4 (N1959, N1951, N1087, N221, N1839);
nor NOR3 (N1960, N1946, N1644, N1232);
xor XOR2 (N1961, N1944, N235);
xor XOR2 (N1962, N1955, N49);
xor XOR2 (N1963, N1958, N450);
and AND3 (N1964, N1957, N107, N672);
nand NAND3 (N1965, N1961, N1477, N73);
not NOT1 (N1966, N1962);
not NOT1 (N1967, N1966);
buf BUF1 (N1968, N1952);
and AND3 (N1969, N1949, N1529, N1178);
or OR3 (N1970, N1960, N1758, N220);
xor XOR2 (N1971, N1959, N1106);
not NOT1 (N1972, N1963);
nor NOR2 (N1973, N1956, N1724);
nor NOR4 (N1974, N1968, N1720, N1401, N720);
xor XOR2 (N1975, N1964, N394);
nand NAND3 (N1976, N1970, N502, N1341);
buf BUF1 (N1977, N1971);
nand NAND3 (N1978, N1977, N998, N1900);
nor NOR2 (N1979, N1953, N711);
nand NAND3 (N1980, N1973, N275, N1633);
or OR2 (N1981, N1965, N148);
nor NOR4 (N1982, N1976, N1566, N1823, N1377);
xor XOR2 (N1983, N1981, N827);
buf BUF1 (N1984, N1967);
buf BUF1 (N1985, N1983);
buf BUF1 (N1986, N1985);
xor XOR2 (N1987, N1979, N402);
xor XOR2 (N1988, N1969, N1918);
and AND3 (N1989, N1975, N18, N500);
nor NOR3 (N1990, N1984, N1624, N781);
nor NOR4 (N1991, N1989, N1848, N766, N922);
nor NOR2 (N1992, N1986, N1951);
and AND4 (N1993, N1988, N856, N780, N1374);
or OR3 (N1994, N1980, N988, N1203);
nor NOR3 (N1995, N1972, N1898, N366);
nand NAND2 (N1996, N1990, N238);
nor NOR4 (N1997, N1996, N233, N1608, N1994);
nand NAND2 (N1998, N930, N1694);
nand NAND4 (N1999, N1995, N44, N1702, N155);
buf BUF1 (N2000, N1999);
and AND4 (N2001, N1991, N786, N1451, N62);
xor XOR2 (N2002, N1987, N1505);
and AND4 (N2003, N1982, N542, N22, N1315);
nand NAND3 (N2004, N1998, N29, N288);
nor NOR2 (N2005, N1978, N1512);
xor XOR2 (N2006, N2003, N132);
buf BUF1 (N2007, N2000);
nand NAND3 (N2008, N2004, N78, N763);
buf BUF1 (N2009, N1974);
and AND3 (N2010, N2005, N1126, N826);
or OR4 (N2011, N2009, N1340, N443, N1739);
or OR2 (N2012, N2007, N880);
buf BUF1 (N2013, N2012);
not NOT1 (N2014, N1992);
and AND2 (N2015, N2013, N404);
and AND3 (N2016, N1993, N1743, N497);
not NOT1 (N2017, N2010);
xor XOR2 (N2018, N2015, N376);
nand NAND3 (N2019, N2016, N1714, N1818);
and AND3 (N2020, N2011, N628, N89);
or OR2 (N2021, N2018, N139);
or OR2 (N2022, N2006, N341);
xor XOR2 (N2023, N2019, N1916);
buf BUF1 (N2024, N2017);
nand NAND4 (N2025, N2021, N1598, N1930, N1911);
buf BUF1 (N2026, N2001);
xor XOR2 (N2027, N2025, N1977);
not NOT1 (N2028, N2027);
not NOT1 (N2029, N2008);
nor NOR3 (N2030, N2026, N730, N1929);
nor NOR4 (N2031, N1997, N1854, N494, N561);
nor NOR3 (N2032, N2028, N1587, N853);
nor NOR2 (N2033, N2020, N1132);
or OR4 (N2034, N2032, N1416, N1517, N1);
buf BUF1 (N2035, N2022);
nand NAND2 (N2036, N2024, N1692);
not NOT1 (N2037, N2029);
nand NAND2 (N2038, N2002, N832);
nand NAND4 (N2039, N2030, N218, N1259, N1658);
nor NOR3 (N2040, N2037, N1342, N1613);
not NOT1 (N2041, N2039);
and AND2 (N2042, N2023, N1766);
and AND4 (N2043, N2033, N650, N275, N1407);
buf BUF1 (N2044, N2043);
and AND3 (N2045, N2041, N1011, N1144);
buf BUF1 (N2046, N2034);
nand NAND3 (N2047, N2046, N1100, N1430);
xor XOR2 (N2048, N2044, N1614);
buf BUF1 (N2049, N2047);
and AND3 (N2050, N2045, N1905, N493);
or OR2 (N2051, N2035, N1126);
nor NOR3 (N2052, N2038, N244, N759);
and AND4 (N2053, N2051, N1518, N1721, N1727);
nand NAND4 (N2054, N2036, N1438, N1486, N1844);
and AND4 (N2055, N2040, N1411, N402, N1764);
nor NOR3 (N2056, N2014, N1581, N1109);
not NOT1 (N2057, N2050);
and AND2 (N2058, N2042, N1690);
xor XOR2 (N2059, N2049, N1666);
or OR4 (N2060, N2031, N313, N777, N1897);
or OR3 (N2061, N2052, N1043, N1449);
and AND2 (N2062, N2055, N679);
or OR3 (N2063, N2062, N1139, N284);
xor XOR2 (N2064, N2054, N87);
nor NOR2 (N2065, N2048, N596);
buf BUF1 (N2066, N2053);
nor NOR4 (N2067, N2066, N1231, N1205, N1675);
nand NAND4 (N2068, N2065, N553, N589, N1499);
not NOT1 (N2069, N2064);
buf BUF1 (N2070, N2059);
xor XOR2 (N2071, N2068, N1352);
buf BUF1 (N2072, N2057);
nand NAND3 (N2073, N2070, N1510, N87);
and AND2 (N2074, N2058, N652);
buf BUF1 (N2075, N2061);
or OR4 (N2076, N2074, N105, N450, N1573);
and AND3 (N2077, N2063, N1995, N1502);
and AND2 (N2078, N2060, N360);
nand NAND3 (N2079, N2069, N547, N322);
nand NAND2 (N2080, N2077, N1730);
nor NOR4 (N2081, N2080, N742, N758, N549);
xor XOR2 (N2082, N2081, N1898);
buf BUF1 (N2083, N2067);
and AND4 (N2084, N2056, N1605, N906, N1825);
xor XOR2 (N2085, N2082, N812);
xor XOR2 (N2086, N2078, N635);
nand NAND2 (N2087, N2071, N110);
not NOT1 (N2088, N2075);
buf BUF1 (N2089, N2073);
nand NAND3 (N2090, N2086, N716, N310);
or OR2 (N2091, N2087, N327);
xor XOR2 (N2092, N2076, N501);
xor XOR2 (N2093, N2092, N863);
or OR4 (N2094, N2093, N1802, N51, N891);
or OR4 (N2095, N2084, N1911, N44, N1196);
nand NAND4 (N2096, N2091, N1510, N1341, N1640);
and AND3 (N2097, N2085, N1807, N1166);
not NOT1 (N2098, N2079);
nand NAND4 (N2099, N2088, N841, N1300, N1389);
nand NAND4 (N2100, N2096, N414, N552, N88);
nand NAND4 (N2101, N2090, N1767, N1924, N1031);
and AND4 (N2102, N2083, N1403, N1608, N374);
not NOT1 (N2103, N2094);
not NOT1 (N2104, N2103);
buf BUF1 (N2105, N2100);
xor XOR2 (N2106, N2098, N856);
or OR2 (N2107, N2101, N1834);
and AND3 (N2108, N2106, N768, N583);
xor XOR2 (N2109, N2095, N199);
or OR3 (N2110, N2109, N943, N1339);
buf BUF1 (N2111, N2097);
and AND4 (N2112, N2099, N357, N45, N1214);
nand NAND4 (N2113, N2108, N1531, N1770, N1278);
nor NOR2 (N2114, N2107, N201);
xor XOR2 (N2115, N2113, N1433);
buf BUF1 (N2116, N2114);
nor NOR2 (N2117, N2115, N1276);
and AND4 (N2118, N2072, N493, N665, N840);
not NOT1 (N2119, N2105);
buf BUF1 (N2120, N2117);
not NOT1 (N2121, N2116);
nand NAND4 (N2122, N2119, N963, N1575, N1150);
nand NAND3 (N2123, N2122, N669, N1733);
or OR3 (N2124, N2111, N383, N602);
buf BUF1 (N2125, N2104);
nand NAND4 (N2126, N2120, N1663, N1046, N1752);
and AND3 (N2127, N2112, N324, N1406);
not NOT1 (N2128, N2121);
buf BUF1 (N2129, N2128);
buf BUF1 (N2130, N2125);
xor XOR2 (N2131, N2110, N1658);
buf BUF1 (N2132, N2102);
not NOT1 (N2133, N2127);
not NOT1 (N2134, N2131);
not NOT1 (N2135, N2124);
buf BUF1 (N2136, N2126);
not NOT1 (N2137, N2132);
buf BUF1 (N2138, N2118);
buf BUF1 (N2139, N2135);
xor XOR2 (N2140, N2089, N94);
nor NOR3 (N2141, N2133, N1187, N90);
nor NOR4 (N2142, N2123, N656, N1889, N188);
nand NAND2 (N2143, N2139, N2062);
and AND4 (N2144, N2136, N778, N1564, N758);
nand NAND3 (N2145, N2142, N559, N1876);
not NOT1 (N2146, N2129);
buf BUF1 (N2147, N2143);
or OR3 (N2148, N2134, N1002, N238);
nand NAND3 (N2149, N2145, N707, N724);
nor NOR3 (N2150, N2137, N1013, N498);
xor XOR2 (N2151, N2149, N465);
or OR2 (N2152, N2148, N1545);
and AND3 (N2153, N2150, N1878, N1216);
xor XOR2 (N2154, N2141, N1909);
and AND2 (N2155, N2151, N2036);
and AND3 (N2156, N2146, N703, N647);
or OR4 (N2157, N2154, N24, N473, N2130);
xor XOR2 (N2158, N1804, N1031);
xor XOR2 (N2159, N2155, N2134);
nand NAND4 (N2160, N2138, N1143, N351, N865);
and AND4 (N2161, N2157, N198, N899, N869);
buf BUF1 (N2162, N2147);
buf BUF1 (N2163, N2162);
or OR3 (N2164, N2156, N1186, N1029);
nand NAND3 (N2165, N2152, N1535, N359);
not NOT1 (N2166, N2165);
nand NAND4 (N2167, N2164, N1642, N228, N2156);
nand NAND4 (N2168, N2140, N433, N1030, N297);
and AND3 (N2169, N2159, N550, N1820);
not NOT1 (N2170, N2169);
buf BUF1 (N2171, N2160);
nor NOR2 (N2172, N2158, N1063);
not NOT1 (N2173, N2172);
xor XOR2 (N2174, N2173, N316);
or OR2 (N2175, N2144, N207);
xor XOR2 (N2176, N2171, N922);
nand NAND3 (N2177, N2176, N1499, N132);
not NOT1 (N2178, N2177);
not NOT1 (N2179, N2166);
buf BUF1 (N2180, N2163);
not NOT1 (N2181, N2161);
xor XOR2 (N2182, N2181, N978);
xor XOR2 (N2183, N2153, N20);
and AND2 (N2184, N2178, N1533);
buf BUF1 (N2185, N2175);
or OR2 (N2186, N2167, N1304);
buf BUF1 (N2187, N2168);
nor NOR3 (N2188, N2183, N1441, N323);
buf BUF1 (N2189, N2184);
buf BUF1 (N2190, N2187);
nor NOR2 (N2191, N2170, N1990);
nand NAND3 (N2192, N2179, N386, N603);
xor XOR2 (N2193, N2188, N1835);
buf BUF1 (N2194, N2191);
xor XOR2 (N2195, N2189, N1265);
nand NAND3 (N2196, N2195, N1963, N308);
nand NAND3 (N2197, N2186, N1668, N221);
nor NOR3 (N2198, N2197, N778, N853);
buf BUF1 (N2199, N2182);
or OR3 (N2200, N2193, N1427, N1170);
xor XOR2 (N2201, N2196, N1919);
nor NOR4 (N2202, N2194, N1918, N185, N910);
and AND4 (N2203, N2202, N1753, N1524, N1611);
buf BUF1 (N2204, N2180);
and AND2 (N2205, N2200, N1384);
nor NOR3 (N2206, N2190, N1875, N852);
nor NOR2 (N2207, N2205, N792);
buf BUF1 (N2208, N2203);
nand NAND2 (N2209, N2207, N1919);
not NOT1 (N2210, N2204);
nand NAND3 (N2211, N2208, N1598, N2151);
or OR3 (N2212, N2209, N1075, N679);
xor XOR2 (N2213, N2206, N1314);
and AND4 (N2214, N2199, N1959, N835, N1585);
not NOT1 (N2215, N2174);
buf BUF1 (N2216, N2215);
xor XOR2 (N2217, N2212, N717);
nand NAND3 (N2218, N2201, N1266, N218);
not NOT1 (N2219, N2216);
and AND4 (N2220, N2210, N989, N903, N1295);
xor XOR2 (N2221, N2185, N106);
xor XOR2 (N2222, N2218, N1243);
nand NAND3 (N2223, N2198, N327, N414);
xor XOR2 (N2224, N2217, N1161);
nor NOR3 (N2225, N2220, N2106, N58);
and AND3 (N2226, N2211, N214, N559);
nand NAND2 (N2227, N2221, N1145);
and AND3 (N2228, N2225, N1843, N1148);
not NOT1 (N2229, N2228);
nand NAND2 (N2230, N2229, N193);
or OR4 (N2231, N2222, N1622, N1412, N2001);
nand NAND4 (N2232, N2226, N2212, N1701, N295);
buf BUF1 (N2233, N2230);
nand NAND3 (N2234, N2214, N507, N1436);
and AND2 (N2235, N2213, N223);
nor NOR3 (N2236, N2235, N203, N1384);
buf BUF1 (N2237, N2233);
nand NAND3 (N2238, N2219, N1402, N1267);
xor XOR2 (N2239, N2234, N785);
xor XOR2 (N2240, N2239, N1772);
nand NAND2 (N2241, N2238, N1595);
not NOT1 (N2242, N2240);
or OR3 (N2243, N2241, N1662, N1258);
or OR3 (N2244, N2236, N2128, N2113);
xor XOR2 (N2245, N2232, N668);
xor XOR2 (N2246, N2192, N1804);
or OR3 (N2247, N2224, N627, N2187);
xor XOR2 (N2248, N2237, N1424);
nand NAND3 (N2249, N2245, N1910, N1606);
buf BUF1 (N2250, N2247);
not NOT1 (N2251, N2223);
not NOT1 (N2252, N2249);
nor NOR3 (N2253, N2250, N592, N580);
or OR2 (N2254, N2246, N796);
buf BUF1 (N2255, N2248);
or OR2 (N2256, N2253, N1276);
buf BUF1 (N2257, N2231);
not NOT1 (N2258, N2255);
or OR4 (N2259, N2258, N1501, N2189, N2099);
xor XOR2 (N2260, N2259, N1288);
buf BUF1 (N2261, N2257);
and AND3 (N2262, N2227, N712, N1999);
nand NAND3 (N2263, N2261, N1941, N299);
xor XOR2 (N2264, N2263, N677);
and AND4 (N2265, N2252, N1757, N278, N1868);
not NOT1 (N2266, N2260);
nand NAND3 (N2267, N2243, N249, N381);
buf BUF1 (N2268, N2244);
xor XOR2 (N2269, N2268, N1791);
and AND3 (N2270, N2242, N295, N811);
xor XOR2 (N2271, N2262, N1841);
nand NAND3 (N2272, N2265, N648, N528);
or OR3 (N2273, N2256, N383, N818);
nand NAND2 (N2274, N2272, N195);
xor XOR2 (N2275, N2271, N1569);
and AND3 (N2276, N2269, N1314, N536);
nand NAND2 (N2277, N2275, N1417);
buf BUF1 (N2278, N2274);
nand NAND2 (N2279, N2254, N1837);
xor XOR2 (N2280, N2273, N401);
and AND3 (N2281, N2277, N89, N716);
nand NAND4 (N2282, N2276, N1377, N881, N1364);
and AND3 (N2283, N2251, N1564, N1033);
not NOT1 (N2284, N2267);
not NOT1 (N2285, N2266);
not NOT1 (N2286, N2282);
nor NOR3 (N2287, N2286, N716, N3);
or OR2 (N2288, N2279, N1140);
buf BUF1 (N2289, N2285);
buf BUF1 (N2290, N2287);
nor NOR4 (N2291, N2290, N957, N392, N1987);
not NOT1 (N2292, N2270);
not NOT1 (N2293, N2281);
nor NOR3 (N2294, N2288, N1746, N1785);
nor NOR2 (N2295, N2264, N817);
not NOT1 (N2296, N2278);
or OR3 (N2297, N2284, N1711, N909);
xor XOR2 (N2298, N2291, N892);
not NOT1 (N2299, N2297);
nand NAND2 (N2300, N2298, N2108);
nand NAND4 (N2301, N2283, N1249, N1811, N582);
not NOT1 (N2302, N2295);
not NOT1 (N2303, N2296);
not NOT1 (N2304, N2299);
xor XOR2 (N2305, N2292, N1930);
and AND2 (N2306, N2304, N1623);
not NOT1 (N2307, N2306);
buf BUF1 (N2308, N2302);
buf BUF1 (N2309, N2301);
and AND2 (N2310, N2308, N582);
or OR4 (N2311, N2280, N981, N182, N1074);
or OR3 (N2312, N2294, N477, N1307);
not NOT1 (N2313, N2312);
nor NOR2 (N2314, N2307, N1791);
nor NOR3 (N2315, N2293, N1150, N137);
nand NAND3 (N2316, N2289, N646, N987);
not NOT1 (N2317, N2311);
xor XOR2 (N2318, N2309, N1187);
and AND3 (N2319, N2303, N1936, N477);
and AND3 (N2320, N2310, N1046, N665);
nor NOR4 (N2321, N2318, N1101, N964, N1655);
or OR3 (N2322, N2300, N2160, N1546);
nand NAND4 (N2323, N2315, N792, N124, N382);
nand NAND2 (N2324, N2314, N558);
nor NOR2 (N2325, N2320, N1995);
or OR4 (N2326, N2313, N922, N115, N1612);
or OR4 (N2327, N2317, N691, N314, N1442);
and AND3 (N2328, N2322, N1884, N926);
or OR4 (N2329, N2327, N1971, N1581, N1608);
buf BUF1 (N2330, N2316);
nor NOR3 (N2331, N2329, N947, N1904);
or OR4 (N2332, N2326, N335, N83, N1990);
xor XOR2 (N2333, N2323, N1327);
xor XOR2 (N2334, N2324, N1822);
buf BUF1 (N2335, N2321);
or OR2 (N2336, N2325, N65);
or OR3 (N2337, N2336, N1945, N1808);
buf BUF1 (N2338, N2337);
not NOT1 (N2339, N2305);
and AND2 (N2340, N2335, N137);
buf BUF1 (N2341, N2330);
nor NOR3 (N2342, N2319, N1520, N1995);
buf BUF1 (N2343, N2328);
not NOT1 (N2344, N2331);
and AND3 (N2345, N2343, N2053, N2192);
or OR3 (N2346, N2340, N1434, N411);
buf BUF1 (N2347, N2342);
nand NAND4 (N2348, N2345, N1656, N2064, N311);
or OR4 (N2349, N2332, N772, N548, N367);
buf BUF1 (N2350, N2334);
xor XOR2 (N2351, N2349, N1544);
and AND2 (N2352, N2351, N2189);
xor XOR2 (N2353, N2348, N2156);
buf BUF1 (N2354, N2344);
buf BUF1 (N2355, N2346);
not NOT1 (N2356, N2339);
not NOT1 (N2357, N2341);
or OR4 (N2358, N2353, N729, N129, N950);
nor NOR4 (N2359, N2352, N624, N386, N138);
xor XOR2 (N2360, N2358, N730);
xor XOR2 (N2361, N2350, N1472);
nor NOR2 (N2362, N2338, N690);
and AND3 (N2363, N2359, N321, N191);
nand NAND3 (N2364, N2362, N1840, N712);
xor XOR2 (N2365, N2356, N65);
or OR4 (N2366, N2363, N1979, N1780, N94);
buf BUF1 (N2367, N2357);
xor XOR2 (N2368, N2364, N1627);
not NOT1 (N2369, N2360);
not NOT1 (N2370, N2368);
or OR3 (N2371, N2366, N1152, N1632);
or OR3 (N2372, N2354, N1800, N2178);
nand NAND3 (N2373, N2369, N563, N1698);
and AND4 (N2374, N2367, N1280, N1120, N216);
nor NOR3 (N2375, N2372, N203, N1046);
xor XOR2 (N2376, N2355, N1696);
nand NAND3 (N2377, N2370, N1100, N1440);
or OR4 (N2378, N2377, N1172, N1010, N1346);
buf BUF1 (N2379, N2371);
and AND4 (N2380, N2373, N2058, N208, N2169);
nand NAND4 (N2381, N2378, N927, N1426, N936);
and AND2 (N2382, N2361, N140);
nand NAND2 (N2383, N2347, N1367);
buf BUF1 (N2384, N2375);
not NOT1 (N2385, N2384);
buf BUF1 (N2386, N2379);
nand NAND3 (N2387, N2380, N279, N891);
xor XOR2 (N2388, N2381, N1193);
and AND4 (N2389, N2365, N1003, N1950, N1460);
nand NAND3 (N2390, N2389, N1823, N339);
and AND2 (N2391, N2333, N133);
and AND3 (N2392, N2387, N217, N497);
and AND2 (N2393, N2374, N786);
and AND3 (N2394, N2391, N1960, N2172);
not NOT1 (N2395, N2390);
not NOT1 (N2396, N2383);
nand NAND4 (N2397, N2395, N2246, N1680, N1855);
xor XOR2 (N2398, N2388, N742);
xor XOR2 (N2399, N2396, N915);
xor XOR2 (N2400, N2392, N1193);
or OR3 (N2401, N2393, N369, N1109);
nand NAND4 (N2402, N2385, N240, N1189, N787);
nand NAND3 (N2403, N2394, N1989, N476);
or OR3 (N2404, N2401, N1638, N1843);
xor XOR2 (N2405, N2399, N1527);
not NOT1 (N2406, N2404);
not NOT1 (N2407, N2402);
and AND4 (N2408, N2386, N2254, N1105, N1018);
xor XOR2 (N2409, N2398, N2275);
and AND3 (N2410, N2400, N785, N1817);
nor NOR2 (N2411, N2403, N2052);
not NOT1 (N2412, N2376);
xor XOR2 (N2413, N2409, N998);
and AND3 (N2414, N2410, N798, N1337);
xor XOR2 (N2415, N2412, N2170);
nor NOR4 (N2416, N2382, N1655, N114, N1447);
and AND4 (N2417, N2407, N1792, N1775, N1204);
nand NAND3 (N2418, N2405, N795, N46);
nor NOR4 (N2419, N2411, N970, N328, N2080);
buf BUF1 (N2420, N2419);
nand NAND3 (N2421, N2415, N1867, N1895);
buf BUF1 (N2422, N2414);
nand NAND2 (N2423, N2397, N651);
nand NAND3 (N2424, N2418, N942, N2022);
buf BUF1 (N2425, N2416);
nor NOR3 (N2426, N2417, N1451, N1284);
nor NOR2 (N2427, N2424, N1139);
buf BUF1 (N2428, N2425);
and AND3 (N2429, N2422, N339, N170);
or OR2 (N2430, N2421, N1197);
buf BUF1 (N2431, N2427);
nand NAND4 (N2432, N2428, N899, N733, N1441);
or OR2 (N2433, N2406, N1506);
nor NOR2 (N2434, N2423, N51);
and AND3 (N2435, N2426, N815, N2343);
buf BUF1 (N2436, N2434);
not NOT1 (N2437, N2435);
nand NAND4 (N2438, N2413, N256, N533, N1147);
or OR2 (N2439, N2420, N1850);
nand NAND4 (N2440, N2432, N305, N832, N2226);
or OR2 (N2441, N2433, N1050);
xor XOR2 (N2442, N2429, N1455);
xor XOR2 (N2443, N2439, N54);
or OR2 (N2444, N2431, N836);
not NOT1 (N2445, N2438);
nor NOR4 (N2446, N2441, N2236, N2210, N22);
not NOT1 (N2447, N2408);
and AND4 (N2448, N2440, N292, N347, N716);
or OR3 (N2449, N2446, N2050, N1811);
and AND2 (N2450, N2449, N612);
and AND4 (N2451, N2436, N920, N778, N83);
nor NOR4 (N2452, N2450, N2073, N1451, N2223);
nand NAND4 (N2453, N2452, N1186, N503, N546);
buf BUF1 (N2454, N2453);
buf BUF1 (N2455, N2454);
or OR3 (N2456, N2444, N440, N1506);
nand NAND4 (N2457, N2451, N1743, N623, N1001);
and AND2 (N2458, N2447, N1243);
and AND2 (N2459, N2448, N357);
buf BUF1 (N2460, N2430);
buf BUF1 (N2461, N2455);
not NOT1 (N2462, N2456);
nand NAND2 (N2463, N2445, N1702);
buf BUF1 (N2464, N2442);
and AND4 (N2465, N2460, N964, N2180, N306);
and AND3 (N2466, N2465, N230, N1821);
or OR4 (N2467, N2466, N1359, N531, N2350);
nand NAND3 (N2468, N2458, N2076, N1659);
nor NOR4 (N2469, N2468, N924, N2331, N415);
not NOT1 (N2470, N2463);
xor XOR2 (N2471, N2470, N123);
nand NAND3 (N2472, N2461, N1983, N202);
not NOT1 (N2473, N2437);
xor XOR2 (N2474, N2457, N1984);
nand NAND2 (N2475, N2467, N2313);
or OR4 (N2476, N2474, N1593, N1288, N1529);
and AND4 (N2477, N2476, N652, N2364, N2105);
or OR3 (N2478, N2471, N2, N328);
buf BUF1 (N2479, N2464);
or OR4 (N2480, N2478, N1691, N579, N1743);
and AND4 (N2481, N2479, N141, N1576, N1128);
buf BUF1 (N2482, N2477);
buf BUF1 (N2483, N2459);
xor XOR2 (N2484, N2481, N1396);
and AND3 (N2485, N2472, N522, N1245);
nor NOR3 (N2486, N2485, N1778, N2082);
xor XOR2 (N2487, N2483, N1209);
xor XOR2 (N2488, N2469, N1784);
and AND2 (N2489, N2462, N2244);
xor XOR2 (N2490, N2484, N1051);
not NOT1 (N2491, N2487);
nor NOR2 (N2492, N2490, N887);
nor NOR3 (N2493, N2473, N1111, N1610);
not NOT1 (N2494, N2488);
nor NOR4 (N2495, N2492, N590, N750, N2386);
xor XOR2 (N2496, N2443, N1269);
or OR3 (N2497, N2495, N1733, N624);
and AND2 (N2498, N2494, N2020);
buf BUF1 (N2499, N2496);
nand NAND2 (N2500, N2493, N116);
buf BUF1 (N2501, N2497);
nor NOR3 (N2502, N2500, N2210, N1246);
nor NOR3 (N2503, N2501, N669, N905);
nor NOR4 (N2504, N2498, N848, N1993, N1845);
buf BUF1 (N2505, N2502);
nor NOR3 (N2506, N2475, N1747, N1419);
buf BUF1 (N2507, N2480);
or OR3 (N2508, N2489, N883, N2438);
buf BUF1 (N2509, N2503);
and AND2 (N2510, N2499, N783);
nor NOR3 (N2511, N2491, N1962, N5);
and AND2 (N2512, N2504, N1593);
and AND4 (N2513, N2510, N1892, N2120, N1318);
xor XOR2 (N2514, N2505, N1621);
buf BUF1 (N2515, N2509);
nand NAND3 (N2516, N2513, N555, N2165);
and AND4 (N2517, N2516, N306, N2438, N72);
and AND3 (N2518, N2515, N119, N547);
buf BUF1 (N2519, N2518);
or OR4 (N2520, N2512, N2259, N1525, N2154);
and AND4 (N2521, N2519, N501, N2154, N482);
buf BUF1 (N2522, N2482);
nand NAND2 (N2523, N2514, N644);
buf BUF1 (N2524, N2507);
and AND3 (N2525, N2524, N2483, N1669);
nand NAND2 (N2526, N2520, N1480);
not NOT1 (N2527, N2508);
not NOT1 (N2528, N2522);
xor XOR2 (N2529, N2521, N2091);
xor XOR2 (N2530, N2486, N2028);
xor XOR2 (N2531, N2529, N1748);
xor XOR2 (N2532, N2523, N1393);
not NOT1 (N2533, N2525);
and AND2 (N2534, N2527, N1676);
not NOT1 (N2535, N2528);
buf BUF1 (N2536, N2530);
xor XOR2 (N2537, N2506, N2157);
nor NOR2 (N2538, N2531, N356);
and AND3 (N2539, N2535, N506, N1597);
nand NAND3 (N2540, N2517, N1030, N1477);
nand NAND3 (N2541, N2534, N564, N518);
not NOT1 (N2542, N2536);
nand NAND4 (N2543, N2526, N2162, N704, N1711);
xor XOR2 (N2544, N2532, N176);
buf BUF1 (N2545, N2542);
buf BUF1 (N2546, N2539);
or OR3 (N2547, N2540, N1888, N1954);
nor NOR4 (N2548, N2546, N783, N1726, N1814);
and AND2 (N2549, N2541, N1229);
not NOT1 (N2550, N2538);
nand NAND3 (N2551, N2533, N712, N823);
buf BUF1 (N2552, N2543);
or OR3 (N2553, N2545, N1361, N2005);
not NOT1 (N2554, N2549);
buf BUF1 (N2555, N2552);
buf BUF1 (N2556, N2537);
xor XOR2 (N2557, N2550, N326);
nand NAND4 (N2558, N2551, N1309, N1345, N639);
and AND4 (N2559, N2544, N1063, N2401, N1090);
and AND2 (N2560, N2558, N366);
buf BUF1 (N2561, N2547);
xor XOR2 (N2562, N2557, N116);
nor NOR3 (N2563, N2554, N2338, N797);
nand NAND3 (N2564, N2560, N944, N806);
nand NAND4 (N2565, N2561, N35, N1918, N2027);
or OR4 (N2566, N2565, N550, N76, N1794);
and AND2 (N2567, N2511, N1381);
xor XOR2 (N2568, N2559, N1761);
not NOT1 (N2569, N2548);
buf BUF1 (N2570, N2564);
or OR3 (N2571, N2563, N236, N2356);
buf BUF1 (N2572, N2569);
nand NAND3 (N2573, N2568, N2354, N1421);
and AND4 (N2574, N2571, N2207, N275, N2259);
not NOT1 (N2575, N2567);
xor XOR2 (N2576, N2575, N2275);
nor NOR4 (N2577, N2556, N138, N498, N1087);
buf BUF1 (N2578, N2573);
buf BUF1 (N2579, N2574);
or OR4 (N2580, N2579, N1601, N1101, N2300);
nor NOR3 (N2581, N2578, N1791, N2325);
nand NAND4 (N2582, N2580, N1662, N905, N1856);
xor XOR2 (N2583, N2562, N219);
or OR3 (N2584, N2577, N1467, N2441);
or OR2 (N2585, N2581, N2050);
buf BUF1 (N2586, N2553);
or OR4 (N2587, N2572, N2348, N1573, N1104);
and AND4 (N2588, N2555, N1240, N1066, N400);
or OR3 (N2589, N2587, N1093, N62);
not NOT1 (N2590, N2566);
or OR4 (N2591, N2590, N1761, N478, N2445);
xor XOR2 (N2592, N2584, N534);
nand NAND3 (N2593, N2576, N465, N463);
nor NOR2 (N2594, N2592, N415);
or OR2 (N2595, N2582, N1617);
nor NOR2 (N2596, N2570, N2389);
nand NAND2 (N2597, N2583, N180);
xor XOR2 (N2598, N2596, N1757);
or OR4 (N2599, N2585, N2060, N1831, N1097);
nor NOR4 (N2600, N2595, N1967, N732, N2060);
or OR4 (N2601, N2591, N2311, N182, N1223);
not NOT1 (N2602, N2588);
and AND3 (N2603, N2598, N1501, N2403);
not NOT1 (N2604, N2594);
nand NAND2 (N2605, N2603, N1478);
nor NOR4 (N2606, N2604, N2019, N1624, N1623);
nand NAND4 (N2607, N2589, N1368, N145, N2279);
buf BUF1 (N2608, N2607);
nand NAND2 (N2609, N2597, N1134);
and AND4 (N2610, N2586, N1169, N499, N905);
nor NOR3 (N2611, N2609, N339, N284);
or OR4 (N2612, N2605, N397, N2392, N833);
nor NOR3 (N2613, N2600, N628, N1850);
not NOT1 (N2614, N2610);
nand NAND4 (N2615, N2614, N30, N2426, N326);
nor NOR4 (N2616, N2593, N1768, N998, N2383);
nand NAND4 (N2617, N2608, N766, N1706, N2534);
not NOT1 (N2618, N2602);
xor XOR2 (N2619, N2617, N374);
nor NOR4 (N2620, N2601, N411, N1963, N2033);
nor NOR2 (N2621, N2615, N972);
not NOT1 (N2622, N2606);
buf BUF1 (N2623, N2619);
buf BUF1 (N2624, N2621);
nand NAND4 (N2625, N2599, N1320, N39, N2594);
nor NOR3 (N2626, N2612, N156, N2545);
buf BUF1 (N2627, N2618);
xor XOR2 (N2628, N2622, N1092);
not NOT1 (N2629, N2623);
or OR4 (N2630, N2611, N2399, N1345, N1717);
and AND3 (N2631, N2627, N217, N1676);
xor XOR2 (N2632, N2630, N1287);
nor NOR3 (N2633, N2624, N2319, N494);
and AND3 (N2634, N2620, N572, N2244);
nor NOR3 (N2635, N2632, N2026, N2120);
nand NAND4 (N2636, N2631, N968, N1200, N1654);
nand NAND4 (N2637, N2634, N1057, N990, N1303);
buf BUF1 (N2638, N2626);
or OR4 (N2639, N2625, N2343, N1969, N2380);
or OR3 (N2640, N2638, N1604, N1935);
nand NAND2 (N2641, N2629, N1776);
nand NAND2 (N2642, N2635, N2261);
or OR2 (N2643, N2640, N423);
nor NOR2 (N2644, N2641, N1694);
and AND2 (N2645, N2639, N2499);
nand NAND4 (N2646, N2637, N865, N363, N627);
or OR3 (N2647, N2628, N2503, N688);
and AND4 (N2648, N2645, N1153, N479, N1613);
or OR4 (N2649, N2636, N1351, N1512, N193);
or OR4 (N2650, N2646, N1250, N1943, N315);
nor NOR3 (N2651, N2648, N1941, N2566);
buf BUF1 (N2652, N2644);
buf BUF1 (N2653, N2647);
and AND3 (N2654, N2650, N678, N107);
and AND3 (N2655, N2649, N1, N186);
not NOT1 (N2656, N2613);
not NOT1 (N2657, N2633);
and AND2 (N2658, N2643, N111);
and AND2 (N2659, N2616, N2142);
and AND3 (N2660, N2642, N1746, N1163);
or OR4 (N2661, N2657, N2376, N2425, N2395);
not NOT1 (N2662, N2659);
buf BUF1 (N2663, N2662);
and AND2 (N2664, N2660, N1713);
nor NOR4 (N2665, N2651, N1798, N617, N490);
buf BUF1 (N2666, N2654);
and AND3 (N2667, N2661, N843, N1402);
nand NAND3 (N2668, N2652, N771, N680);
nand NAND4 (N2669, N2668, N592, N595, N1923);
not NOT1 (N2670, N2666);
and AND4 (N2671, N2663, N1480, N1207, N824);
and AND3 (N2672, N2658, N1068, N1564);
and AND2 (N2673, N2656, N1405);
and AND4 (N2674, N2655, N2319, N2404, N1303);
nand NAND3 (N2675, N2671, N1381, N596);
nand NAND4 (N2676, N2675, N1049, N1830, N331);
and AND4 (N2677, N2673, N1095, N45, N1765);
buf BUF1 (N2678, N2669);
buf BUF1 (N2679, N2653);
or OR4 (N2680, N2678, N86, N2498, N1110);
xor XOR2 (N2681, N2676, N1125);
xor XOR2 (N2682, N2677, N2460);
buf BUF1 (N2683, N2667);
nor NOR4 (N2684, N2683, N2412, N1710, N2498);
buf BUF1 (N2685, N2684);
buf BUF1 (N2686, N2670);
nor NOR2 (N2687, N2672, N343);
or OR4 (N2688, N2664, N1604, N2168, N1702);
nand NAND3 (N2689, N2679, N425, N97);
or OR4 (N2690, N2682, N2616, N2274, N1023);
not NOT1 (N2691, N2680);
and AND2 (N2692, N2681, N2184);
or OR3 (N2693, N2687, N1390, N1553);
nor NOR2 (N2694, N2688, N999);
nor NOR4 (N2695, N2665, N2174, N2637, N747);
nand NAND4 (N2696, N2674, N2609, N200, N880);
and AND4 (N2697, N2689, N1694, N997, N2332);
xor XOR2 (N2698, N2685, N1754);
nor NOR2 (N2699, N2695, N1654);
or OR4 (N2700, N2699, N1515, N1813, N1562);
xor XOR2 (N2701, N2698, N58);
nand NAND3 (N2702, N2694, N1318, N643);
and AND4 (N2703, N2696, N2043, N2623, N2030);
not NOT1 (N2704, N2700);
not NOT1 (N2705, N2703);
or OR3 (N2706, N2693, N845, N1606);
and AND4 (N2707, N2697, N1755, N1674, N1927);
or OR3 (N2708, N2690, N999, N1727);
or OR4 (N2709, N2701, N2611, N2124, N2463);
or OR3 (N2710, N2692, N167, N56);
xor XOR2 (N2711, N2709, N2552);
and AND2 (N2712, N2711, N2468);
xor XOR2 (N2713, N2705, N920);
nor NOR2 (N2714, N2706, N280);
nor NOR2 (N2715, N2710, N2150);
xor XOR2 (N2716, N2708, N220);
and AND2 (N2717, N2714, N1609);
not NOT1 (N2718, N2691);
nand NAND3 (N2719, N2704, N2198, N1146);
buf BUF1 (N2720, N2718);
xor XOR2 (N2721, N2713, N617);
not NOT1 (N2722, N2716);
not NOT1 (N2723, N2720);
nand NAND3 (N2724, N2702, N1573, N34);
buf BUF1 (N2725, N2722);
nand NAND2 (N2726, N2712, N277);
or OR4 (N2727, N2719, N1875, N1949, N415);
not NOT1 (N2728, N2725);
or OR4 (N2729, N2717, N1352, N371, N2318);
and AND2 (N2730, N2729, N2340);
xor XOR2 (N2731, N2726, N2240);
xor XOR2 (N2732, N2730, N579);
buf BUF1 (N2733, N2724);
xor XOR2 (N2734, N2707, N1558);
buf BUF1 (N2735, N2686);
nor NOR2 (N2736, N2723, N2179);
not NOT1 (N2737, N2728);
xor XOR2 (N2738, N2727, N290);
buf BUF1 (N2739, N2733);
nor NOR3 (N2740, N2721, N1391, N1176);
xor XOR2 (N2741, N2731, N2495);
nand NAND4 (N2742, N2737, N1749, N106, N903);
xor XOR2 (N2743, N2739, N2643);
nand NAND3 (N2744, N2740, N2011, N2723);
buf BUF1 (N2745, N2736);
or OR3 (N2746, N2734, N1484, N548);
buf BUF1 (N2747, N2741);
nand NAND4 (N2748, N2735, N1512, N1352, N2483);
or OR4 (N2749, N2748, N1476, N1542, N524);
or OR3 (N2750, N2749, N2602, N814);
or OR4 (N2751, N2744, N38, N572, N1612);
or OR3 (N2752, N2746, N1611, N855);
and AND3 (N2753, N2738, N335, N1708);
not NOT1 (N2754, N2732);
and AND3 (N2755, N2750, N2487, N1538);
nand NAND2 (N2756, N2745, N1659);
nand NAND4 (N2757, N2751, N2587, N242, N1066);
not NOT1 (N2758, N2747);
and AND3 (N2759, N2742, N591, N2331);
nand NAND3 (N2760, N2759, N1408, N178);
xor XOR2 (N2761, N2753, N2553);
buf BUF1 (N2762, N2754);
not NOT1 (N2763, N2762);
nor NOR4 (N2764, N2755, N1283, N2618, N1734);
not NOT1 (N2765, N2763);
buf BUF1 (N2766, N2757);
xor XOR2 (N2767, N2758, N385);
and AND4 (N2768, N2767, N453, N2549, N1880);
nand NAND2 (N2769, N2761, N1381);
nor NOR3 (N2770, N2765, N372, N1300);
buf BUF1 (N2771, N2760);
xor XOR2 (N2772, N2756, N1679);
and AND2 (N2773, N2768, N1554);
nand NAND4 (N2774, N2752, N1459, N1617, N944);
not NOT1 (N2775, N2766);
nand NAND4 (N2776, N2764, N326, N76, N2150);
and AND2 (N2777, N2772, N342);
or OR3 (N2778, N2774, N1602, N1958);
xor XOR2 (N2779, N2776, N2368);
nor NOR3 (N2780, N2775, N1503, N1238);
or OR3 (N2781, N2770, N1190, N1631);
buf BUF1 (N2782, N2715);
xor XOR2 (N2783, N2743, N104);
buf BUF1 (N2784, N2783);
not NOT1 (N2785, N2782);
nand NAND4 (N2786, N2780, N709, N1396, N568);
nor NOR4 (N2787, N2785, N629, N1976, N244);
and AND4 (N2788, N2779, N1337, N1968, N955);
and AND4 (N2789, N2786, N1276, N1238, N1622);
and AND3 (N2790, N2771, N701, N589);
xor XOR2 (N2791, N2784, N2264);
nand NAND4 (N2792, N2781, N2020, N2297, N693);
buf BUF1 (N2793, N2787);
nor NOR3 (N2794, N2773, N1328, N1295);
or OR4 (N2795, N2778, N1300, N1774, N1296);
not NOT1 (N2796, N2794);
nand NAND4 (N2797, N2789, N1924, N2358, N121);
nand NAND3 (N2798, N2795, N1446, N1681);
not NOT1 (N2799, N2788);
xor XOR2 (N2800, N2797, N1187);
xor XOR2 (N2801, N2791, N1892);
xor XOR2 (N2802, N2799, N1763);
not NOT1 (N2803, N2790);
xor XOR2 (N2804, N2800, N2508);
xor XOR2 (N2805, N2804, N1905);
buf BUF1 (N2806, N2802);
not NOT1 (N2807, N2803);
not NOT1 (N2808, N2807);
xor XOR2 (N2809, N2777, N2585);
and AND2 (N2810, N2796, N601);
nor NOR2 (N2811, N2801, N40);
not NOT1 (N2812, N2809);
not NOT1 (N2813, N2805);
or OR4 (N2814, N2806, N2490, N1631, N1150);
nand NAND4 (N2815, N2808, N1106, N732, N2393);
or OR2 (N2816, N2792, N2108);
nor NOR4 (N2817, N2810, N99, N839, N955);
nor NOR3 (N2818, N2798, N148, N238);
or OR2 (N2819, N2818, N1866);
and AND3 (N2820, N2812, N1882, N2254);
not NOT1 (N2821, N2817);
nor NOR3 (N2822, N2819, N2285, N261);
nor NOR2 (N2823, N2811, N1472);
not NOT1 (N2824, N2822);
buf BUF1 (N2825, N2815);
not NOT1 (N2826, N2825);
nand NAND2 (N2827, N2826, N1753);
buf BUF1 (N2828, N2793);
or OR3 (N2829, N2820, N362, N2214);
buf BUF1 (N2830, N2813);
and AND3 (N2831, N2816, N1951, N1867);
buf BUF1 (N2832, N2828);
xor XOR2 (N2833, N2831, N1268);
not NOT1 (N2834, N2832);
or OR3 (N2835, N2834, N1847, N463);
nor NOR3 (N2836, N2833, N2727, N1098);
or OR2 (N2837, N2814, N795);
xor XOR2 (N2838, N2821, N99);
or OR3 (N2839, N2829, N657, N1758);
nand NAND3 (N2840, N2823, N32, N2703);
not NOT1 (N2841, N2836);
nand NAND3 (N2842, N2839, N2317, N982);
not NOT1 (N2843, N2837);
xor XOR2 (N2844, N2842, N1436);
and AND4 (N2845, N2840, N1243, N138, N1677);
nor NOR2 (N2846, N2841, N1946);
xor XOR2 (N2847, N2824, N2758);
xor XOR2 (N2848, N2830, N366);
buf BUF1 (N2849, N2848);
not NOT1 (N2850, N2846);
nand NAND4 (N2851, N2843, N866, N912, N1799);
xor XOR2 (N2852, N2850, N1145);
and AND3 (N2853, N2838, N2669, N2473);
xor XOR2 (N2854, N2847, N2774);
nor NOR4 (N2855, N2851, N2791, N812, N1154);
nand NAND4 (N2856, N2844, N1339, N897, N416);
buf BUF1 (N2857, N2856);
nor NOR3 (N2858, N2849, N249, N185);
buf BUF1 (N2859, N2835);
and AND2 (N2860, N2858, N65);
nand NAND4 (N2861, N2855, N2792, N1802, N1800);
or OR2 (N2862, N2859, N1203);
nor NOR2 (N2863, N2852, N1450);
not NOT1 (N2864, N2862);
buf BUF1 (N2865, N2860);
not NOT1 (N2866, N2864);
xor XOR2 (N2867, N2853, N904);
and AND4 (N2868, N2865, N2127, N2341, N419);
nor NOR2 (N2869, N2866, N665);
and AND3 (N2870, N2868, N604, N2671);
or OR2 (N2871, N2861, N676);
not NOT1 (N2872, N2867);
xor XOR2 (N2873, N2863, N1925);
nor NOR2 (N2874, N2857, N119);
buf BUF1 (N2875, N2869);
nor NOR4 (N2876, N2769, N2739, N750, N633);
and AND4 (N2877, N2875, N610, N1463, N1544);
buf BUF1 (N2878, N2871);
nor NOR3 (N2879, N2827, N813, N1088);
not NOT1 (N2880, N2845);
nor NOR4 (N2881, N2873, N391, N1679, N2838);
nand NAND3 (N2882, N2878, N2272, N1509);
or OR4 (N2883, N2874, N1, N1981, N1311);
not NOT1 (N2884, N2882);
not NOT1 (N2885, N2877);
nor NOR3 (N2886, N2870, N2355, N2018);
not NOT1 (N2887, N2881);
buf BUF1 (N2888, N2872);
xor XOR2 (N2889, N2876, N1615);
or OR2 (N2890, N2889, N899);
not NOT1 (N2891, N2887);
nand NAND3 (N2892, N2854, N1641, N2113);
or OR4 (N2893, N2883, N2655, N692, N848);
nand NAND4 (N2894, N2888, N2545, N1623, N1323);
buf BUF1 (N2895, N2885);
and AND2 (N2896, N2880, N103);
not NOT1 (N2897, N2890);
nand NAND2 (N2898, N2879, N1031);
and AND4 (N2899, N2893, N596, N1598, N2234);
xor XOR2 (N2900, N2895, N2829);
nor NOR3 (N2901, N2897, N1034, N1340);
not NOT1 (N2902, N2901);
nor NOR2 (N2903, N2899, N2547);
xor XOR2 (N2904, N2892, N1068);
not NOT1 (N2905, N2900);
not NOT1 (N2906, N2884);
nand NAND2 (N2907, N2903, N2760);
or OR4 (N2908, N2886, N841, N636, N628);
not NOT1 (N2909, N2908);
not NOT1 (N2910, N2896);
and AND3 (N2911, N2905, N1219, N1110);
not NOT1 (N2912, N2902);
buf BUF1 (N2913, N2910);
xor XOR2 (N2914, N2891, N623);
and AND3 (N2915, N2904, N176, N2902);
not NOT1 (N2916, N2906);
not NOT1 (N2917, N2913);
xor XOR2 (N2918, N2898, N872);
xor XOR2 (N2919, N2911, N877);
or OR4 (N2920, N2907, N2569, N1095, N2549);
not NOT1 (N2921, N2912);
nand NAND2 (N2922, N2916, N264);
nor NOR4 (N2923, N2894, N226, N2531, N2158);
buf BUF1 (N2924, N2922);
or OR3 (N2925, N2919, N71, N2451);
not NOT1 (N2926, N2909);
xor XOR2 (N2927, N2923, N2847);
xor XOR2 (N2928, N2926, N798);
or OR4 (N2929, N2920, N2506, N2130, N2668);
xor XOR2 (N2930, N2924, N2148);
and AND3 (N2931, N2929, N2082, N1589);
xor XOR2 (N2932, N2917, N1205);
nand NAND4 (N2933, N2928, N1548, N74, N1765);
xor XOR2 (N2934, N2914, N2493);
or OR3 (N2935, N2918, N126, N855);
nor NOR4 (N2936, N2915, N446, N2597, N1465);
not NOT1 (N2937, N2936);
not NOT1 (N2938, N2927);
buf BUF1 (N2939, N2932);
nand NAND3 (N2940, N2939, N1246, N2849);
buf BUF1 (N2941, N2921);
nor NOR4 (N2942, N2933, N235, N417, N329);
xor XOR2 (N2943, N2935, N2131);
or OR2 (N2944, N2940, N669);
nand NAND2 (N2945, N2930, N111);
buf BUF1 (N2946, N2943);
and AND3 (N2947, N2942, N2339, N1489);
xor XOR2 (N2948, N2941, N579);
xor XOR2 (N2949, N2947, N102);
buf BUF1 (N2950, N2934);
nand NAND3 (N2951, N2944, N1577, N2424);
not NOT1 (N2952, N2945);
or OR3 (N2953, N2948, N2806, N984);
and AND3 (N2954, N2946, N668, N2882);
nand NAND3 (N2955, N2949, N1541, N2626);
not NOT1 (N2956, N2953);
or OR4 (N2957, N2955, N1881, N908, N110);
nand NAND4 (N2958, N2925, N1115, N1149, N2077);
nor NOR2 (N2959, N2938, N1745);
xor XOR2 (N2960, N2931, N791);
or OR3 (N2961, N2952, N2957, N1846);
xor XOR2 (N2962, N934, N2009);
buf BUF1 (N2963, N2951);
nor NOR3 (N2964, N2963, N1582, N294);
and AND3 (N2965, N2937, N1428, N1683);
nor NOR4 (N2966, N2964, N2806, N608, N2208);
buf BUF1 (N2967, N2966);
nor NOR4 (N2968, N2956, N191, N2706, N1957);
xor XOR2 (N2969, N2950, N2592);
nand NAND4 (N2970, N2961, N1588, N1445, N383);
nand NAND2 (N2971, N2954, N1147);
not NOT1 (N2972, N2960);
and AND2 (N2973, N2965, N469);
buf BUF1 (N2974, N2972);
not NOT1 (N2975, N2971);
buf BUF1 (N2976, N2974);
and AND4 (N2977, N2959, N174, N867, N979);
not NOT1 (N2978, N2967);
or OR2 (N2979, N2973, N168);
nand NAND4 (N2980, N2977, N1494, N232, N2444);
nor NOR2 (N2981, N2976, N2635);
xor XOR2 (N2982, N2979, N536);
xor XOR2 (N2983, N2962, N524);
and AND4 (N2984, N2968, N2558, N2457, N2612);
buf BUF1 (N2985, N2969);
and AND3 (N2986, N2982, N567, N2104);
nor NOR2 (N2987, N2980, N2029);
xor XOR2 (N2988, N2970, N2021);
nand NAND3 (N2989, N2984, N862, N831);
not NOT1 (N2990, N2958);
nand NAND2 (N2991, N2985, N2261);
or OR2 (N2992, N2975, N841);
nor NOR2 (N2993, N2992, N1863);
buf BUF1 (N2994, N2983);
nand NAND2 (N2995, N2987, N201);
nor NOR2 (N2996, N2990, N2423);
nand NAND2 (N2997, N2989, N309);
or OR4 (N2998, N2996, N2711, N809, N263);
xor XOR2 (N2999, N2986, N301);
and AND2 (N3000, N2999, N1104);
buf BUF1 (N3001, N2981);
nand NAND2 (N3002, N2991, N2433);
not NOT1 (N3003, N2998);
nor NOR3 (N3004, N2995, N2203, N1668);
buf BUF1 (N3005, N3000);
xor XOR2 (N3006, N3004, N1261);
not NOT1 (N3007, N2997);
nand NAND4 (N3008, N2994, N2039, N1426, N1782);
nor NOR2 (N3009, N3001, N2430);
nor NOR2 (N3010, N3007, N1643);
nor NOR3 (N3011, N3003, N418, N2546);
nand NAND2 (N3012, N3005, N552);
and AND3 (N3013, N2978, N142, N840);
nor NOR2 (N3014, N3013, N2252);
xor XOR2 (N3015, N2988, N968);
or OR3 (N3016, N3014, N2035, N417);
nor NOR4 (N3017, N2993, N2941, N531, N1674);
nor NOR2 (N3018, N3011, N2720);
xor XOR2 (N3019, N3018, N1619);
nor NOR3 (N3020, N3012, N1972, N2814);
nand NAND2 (N3021, N3002, N1540);
xor XOR2 (N3022, N3009, N2000);
buf BUF1 (N3023, N3022);
nand NAND4 (N3024, N3021, N1375, N2311, N432);
nor NOR3 (N3025, N3015, N3001, N350);
or OR3 (N3026, N3023, N2157, N415);
nor NOR4 (N3027, N3024, N1649, N461, N2027);
not NOT1 (N3028, N3027);
buf BUF1 (N3029, N3016);
nand NAND3 (N3030, N3017, N1200, N2283);
not NOT1 (N3031, N3025);
or OR4 (N3032, N3019, N341, N2974, N2715);
nand NAND4 (N3033, N3008, N1920, N2570, N2132);
not NOT1 (N3034, N3033);
xor XOR2 (N3035, N3034, N2125);
or OR4 (N3036, N3020, N1204, N446, N988);
not NOT1 (N3037, N3006);
xor XOR2 (N3038, N3036, N2384);
buf BUF1 (N3039, N3032);
buf BUF1 (N3040, N3030);
or OR3 (N3041, N3039, N955, N1360);
and AND4 (N3042, N3035, N2291, N2645, N579);
or OR3 (N3043, N3029, N703, N2944);
and AND3 (N3044, N3028, N2488, N2685);
not NOT1 (N3045, N3041);
xor XOR2 (N3046, N3045, N543);
buf BUF1 (N3047, N3043);
nand NAND4 (N3048, N3038, N1772, N1969, N525);
buf BUF1 (N3049, N3010);
or OR3 (N3050, N3047, N2111, N506);
and AND2 (N3051, N3040, N2689);
or OR3 (N3052, N3031, N248, N931);
and AND3 (N3053, N3042, N1179, N1757);
xor XOR2 (N3054, N3026, N602);
not NOT1 (N3055, N3049);
not NOT1 (N3056, N3046);
not NOT1 (N3057, N3051);
not NOT1 (N3058, N3050);
not NOT1 (N3059, N3048);
and AND4 (N3060, N3053, N920, N25, N2157);
not NOT1 (N3061, N3058);
buf BUF1 (N3062, N3056);
nor NOR4 (N3063, N3052, N1884, N1268, N2515);
nor NOR2 (N3064, N3054, N2281);
or OR2 (N3065, N3057, N2932);
xor XOR2 (N3066, N3061, N59);
nand NAND4 (N3067, N3044, N1585, N1528, N2494);
nor NOR3 (N3068, N3063, N995, N100);
buf BUF1 (N3069, N3068);
buf BUF1 (N3070, N3055);
buf BUF1 (N3071, N3060);
nor NOR2 (N3072, N3066, N274);
and AND2 (N3073, N3059, N646);
and AND4 (N3074, N3070, N2820, N1192, N594);
xor XOR2 (N3075, N3069, N2693);
and AND3 (N3076, N3075, N1014, N573);
xor XOR2 (N3077, N3073, N2452);
buf BUF1 (N3078, N3067);
and AND2 (N3079, N3065, N22);
and AND3 (N3080, N3076, N705, N1753);
nand NAND4 (N3081, N3071, N1353, N1343, N1700);
nor NOR3 (N3082, N3079, N651, N2473);
not NOT1 (N3083, N3062);
or OR3 (N3084, N3074, N736, N299);
xor XOR2 (N3085, N3082, N537);
nand NAND3 (N3086, N3064, N2654, N1400);
nand NAND3 (N3087, N3085, N1750, N2272);
not NOT1 (N3088, N3080);
buf BUF1 (N3089, N3072);
not NOT1 (N3090, N3081);
not NOT1 (N3091, N3037);
or OR3 (N3092, N3088, N1757, N1070);
not NOT1 (N3093, N3087);
xor XOR2 (N3094, N3092, N1946);
xor XOR2 (N3095, N3078, N1579);
nor NOR4 (N3096, N3094, N2367, N1564, N353);
xor XOR2 (N3097, N3096, N2059);
nand NAND2 (N3098, N3089, N2074);
or OR3 (N3099, N3090, N2822, N2150);
not NOT1 (N3100, N3086);
buf BUF1 (N3101, N3083);
nor NOR2 (N3102, N3077, N2781);
buf BUF1 (N3103, N3091);
nand NAND2 (N3104, N3098, N1316);
xor XOR2 (N3105, N3103, N695);
xor XOR2 (N3106, N3104, N2853);
and AND3 (N3107, N3106, N263, N2402);
nand NAND2 (N3108, N3107, N1812);
nand NAND3 (N3109, N3108, N2786, N2221);
xor XOR2 (N3110, N3097, N2865);
not NOT1 (N3111, N3109);
nor NOR2 (N3112, N3102, N328);
buf BUF1 (N3113, N3093);
nand NAND3 (N3114, N3100, N1853, N3064);
xor XOR2 (N3115, N3105, N2519);
xor XOR2 (N3116, N3101, N1668);
buf BUF1 (N3117, N3095);
or OR3 (N3118, N3084, N186, N1906);
not NOT1 (N3119, N3111);
nor NOR2 (N3120, N3114, N2983);
buf BUF1 (N3121, N3120);
nor NOR4 (N3122, N3099, N2788, N2918, N400);
buf BUF1 (N3123, N3122);
buf BUF1 (N3124, N3110);
not NOT1 (N3125, N3118);
nor NOR4 (N3126, N3113, N1454, N1190, N2893);
nor NOR4 (N3127, N3126, N2617, N3024, N2000);
nor NOR3 (N3128, N3115, N2160, N1456);
and AND3 (N3129, N3119, N1626, N638);
buf BUF1 (N3130, N3123);
not NOT1 (N3131, N3121);
nand NAND3 (N3132, N3128, N3011, N658);
and AND4 (N3133, N3129, N1156, N1283, N211);
nor NOR3 (N3134, N3133, N2754, N1247);
not NOT1 (N3135, N3116);
and AND3 (N3136, N3135, N561, N9);
nand NAND4 (N3137, N3134, N1942, N1105, N2304);
buf BUF1 (N3138, N3132);
and AND4 (N3139, N3130, N1124, N2176, N2563);
and AND2 (N3140, N3127, N1308);
buf BUF1 (N3141, N3136);
not NOT1 (N3142, N3117);
xor XOR2 (N3143, N3112, N80);
nand NAND3 (N3144, N3125, N1850, N2689);
and AND3 (N3145, N3143, N568, N1931);
nor NOR4 (N3146, N3139, N2380, N2824, N1107);
and AND3 (N3147, N3131, N2021, N1804);
nor NOR2 (N3148, N3138, N2227);
not NOT1 (N3149, N3148);
nand NAND2 (N3150, N3149, N321);
nor NOR4 (N3151, N3150, N2497, N2533, N2333);
nor NOR2 (N3152, N3147, N459);
or OR3 (N3153, N3124, N2953, N2900);
and AND3 (N3154, N3141, N1458, N2672);
nor NOR4 (N3155, N3146, N2167, N455, N2097);
nor NOR3 (N3156, N3155, N1956, N172);
xor XOR2 (N3157, N3140, N2076);
nand NAND4 (N3158, N3151, N1952, N2859, N2405);
xor XOR2 (N3159, N3154, N1036);
or OR2 (N3160, N3144, N380);
or OR3 (N3161, N3152, N2068, N1244);
nor NOR4 (N3162, N3137, N1828, N863, N1501);
xor XOR2 (N3163, N3153, N2490);
nor NOR2 (N3164, N3161, N986);
xor XOR2 (N3165, N3158, N259);
buf BUF1 (N3166, N3163);
or OR3 (N3167, N3159, N2710, N1614);
and AND3 (N3168, N3167, N2582, N515);
xor XOR2 (N3169, N3168, N182);
and AND3 (N3170, N3142, N3068, N1304);
not NOT1 (N3171, N3170);
buf BUF1 (N3172, N3169);
and AND2 (N3173, N3166, N2071);
xor XOR2 (N3174, N3173, N342);
and AND3 (N3175, N3162, N287, N685);
xor XOR2 (N3176, N3165, N239);
buf BUF1 (N3177, N3157);
nand NAND3 (N3178, N3171, N1532, N225);
or OR3 (N3179, N3174, N32, N2485);
and AND3 (N3180, N3172, N1285, N1667);
and AND4 (N3181, N3176, N282, N2866, N786);
or OR3 (N3182, N3175, N1739, N3);
buf BUF1 (N3183, N3179);
nand NAND2 (N3184, N3182, N2031);
nand NAND2 (N3185, N3181, N2016);
xor XOR2 (N3186, N3178, N2089);
buf BUF1 (N3187, N3183);
xor XOR2 (N3188, N3180, N2514);
nand NAND2 (N3189, N3145, N104);
buf BUF1 (N3190, N3189);
buf BUF1 (N3191, N3164);
buf BUF1 (N3192, N3186);
xor XOR2 (N3193, N3185, N2796);
nor NOR4 (N3194, N3160, N2433, N2365, N3090);
and AND4 (N3195, N3191, N3156, N3087, N2912);
nor NOR3 (N3196, N871, N2795, N2931);
nand NAND2 (N3197, N3194, N1710);
xor XOR2 (N3198, N3195, N2788);
and AND4 (N3199, N3177, N621, N14, N850);
or OR3 (N3200, N3198, N2060, N1706);
xor XOR2 (N3201, N3187, N2237);
not NOT1 (N3202, N3190);
nand NAND4 (N3203, N3196, N961, N1430, N884);
and AND3 (N3204, N3200, N2318, N2111);
nor NOR4 (N3205, N3202, N2960, N2872, N2043);
buf BUF1 (N3206, N3204);
and AND4 (N3207, N3197, N1406, N854, N1726);
not NOT1 (N3208, N3206);
and AND3 (N3209, N3188, N3140, N1251);
not NOT1 (N3210, N3199);
nand NAND4 (N3211, N3208, N2715, N1078, N2710);
nand NAND3 (N3212, N3192, N2347, N2291);
nand NAND4 (N3213, N3205, N1015, N2450, N827);
xor XOR2 (N3214, N3207, N2895);
or OR3 (N3215, N3193, N2992, N2831);
not NOT1 (N3216, N3213);
or OR3 (N3217, N3214, N1961, N607);
not NOT1 (N3218, N3212);
and AND3 (N3219, N3184, N1163, N1171);
and AND4 (N3220, N3217, N1494, N228, N2444);
endmodule