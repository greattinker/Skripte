// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20;

output N300,N307,N316,N313,N312,N308,N304,N317,N319,N320;

nand NAND3 (N21, N19, N11, N17);
not NOT1 (N22, N14);
nor NOR4 (N23, N22, N12, N12, N12);
nor NOR4 (N24, N4, N8, N5, N22);
nand NAND2 (N25, N13, N14);
nor NOR3 (N26, N20, N20, N24);
or OR3 (N27, N10, N2, N11);
nor NOR2 (N28, N15, N9);
and AND3 (N29, N7, N7, N9);
buf BUF1 (N30, N26);
not NOT1 (N31, N8);
nor NOR2 (N32, N17, N18);
and AND2 (N33, N27, N32);
nor NOR2 (N34, N8, N30);
buf BUF1 (N35, N29);
nor NOR3 (N36, N8, N30, N14);
nor NOR2 (N37, N13, N8);
nor NOR2 (N38, N35, N1);
nor NOR3 (N39, N21, N36, N5);
buf BUF1 (N40, N26);
buf BUF1 (N41, N25);
xor XOR2 (N42, N37, N23);
nand NAND2 (N43, N15, N29);
nand NAND3 (N44, N28, N6, N25);
and AND3 (N45, N39, N5, N8);
buf BUF1 (N46, N40);
and AND3 (N47, N45, N2, N6);
buf BUF1 (N48, N34);
nand NAND3 (N49, N41, N44, N44);
not NOT1 (N50, N13);
nor NOR4 (N51, N38, N26, N7, N2);
not NOT1 (N52, N47);
nor NOR3 (N53, N52, N14, N27);
nand NAND3 (N54, N46, N8, N43);
and AND2 (N55, N11, N24);
or OR2 (N56, N33, N31);
buf BUF1 (N57, N5);
or OR2 (N58, N54, N55);
xor XOR2 (N59, N9, N38);
xor XOR2 (N60, N42, N12);
buf BUF1 (N61, N48);
xor XOR2 (N62, N56, N51);
and AND4 (N63, N25, N39, N13, N19);
nor NOR2 (N64, N53, N43);
or OR2 (N65, N49, N2);
and AND3 (N66, N58, N37, N36);
nor NOR4 (N67, N61, N56, N36, N27);
xor XOR2 (N68, N65, N58);
nor NOR3 (N69, N57, N27, N46);
nor NOR2 (N70, N69, N34);
or OR3 (N71, N60, N1, N51);
nand NAND3 (N72, N63, N12, N58);
nor NOR3 (N73, N59, N30, N22);
not NOT1 (N74, N68);
not NOT1 (N75, N70);
or OR3 (N76, N73, N30, N38);
and AND4 (N77, N74, N34, N76, N67);
nor NOR4 (N78, N13, N39, N71, N26);
and AND2 (N79, N33, N26);
nand NAND3 (N80, N15, N76, N58);
not NOT1 (N81, N79);
xor XOR2 (N82, N77, N6);
nor NOR4 (N83, N62, N37, N81, N20);
xor XOR2 (N84, N4, N62);
or OR2 (N85, N80, N18);
buf BUF1 (N86, N85);
and AND3 (N87, N78, N64, N83);
buf BUF1 (N88, N70);
nor NOR4 (N89, N56, N60, N72, N86);
nor NOR4 (N90, N24, N63, N4, N86);
nand NAND3 (N91, N89, N78, N89);
nand NAND2 (N92, N23, N13);
nor NOR3 (N93, N75, N84, N87);
and AND2 (N94, N41, N36);
and AND4 (N95, N71, N65, N62, N69);
nor NOR3 (N96, N92, N17, N89);
or OR4 (N97, N66, N15, N70, N51);
nand NAND3 (N98, N90, N16, N76);
nand NAND3 (N99, N95, N47, N97);
nor NOR3 (N100, N88, N38, N96);
not NOT1 (N101, N17);
xor XOR2 (N102, N71, N95);
or OR4 (N103, N82, N24, N1, N98);
buf BUF1 (N104, N13);
or OR3 (N105, N50, N34, N18);
or OR3 (N106, N93, N81, N87);
xor XOR2 (N107, N106, N73);
nand NAND2 (N108, N91, N48);
buf BUF1 (N109, N94);
xor XOR2 (N110, N103, N37);
not NOT1 (N111, N100);
or OR4 (N112, N102, N6, N41, N66);
nor NOR4 (N113, N112, N33, N87, N94);
xor XOR2 (N114, N104, N45);
nand NAND4 (N115, N107, N41, N107, N51);
buf BUF1 (N116, N114);
and AND3 (N117, N105, N97, N9);
not NOT1 (N118, N110);
not NOT1 (N119, N113);
nand NAND3 (N120, N116, N28, N70);
buf BUF1 (N121, N117);
nand NAND4 (N122, N108, N82, N97, N27);
buf BUF1 (N123, N101);
nand NAND3 (N124, N111, N111, N8);
and AND4 (N125, N119, N26, N36, N33);
buf BUF1 (N126, N123);
buf BUF1 (N127, N126);
not NOT1 (N128, N109);
and AND3 (N129, N128, N3, N101);
or OR2 (N130, N118, N29);
nor NOR2 (N131, N99, N36);
or OR4 (N132, N121, N7, N120, N13);
xor XOR2 (N133, N78, N45);
or OR4 (N134, N132, N113, N32, N48);
not NOT1 (N135, N127);
or OR2 (N136, N124, N7);
not NOT1 (N137, N122);
buf BUF1 (N138, N134);
and AND2 (N139, N125, N124);
nand NAND2 (N140, N136, N3);
or OR2 (N141, N115, N54);
or OR3 (N142, N137, N7, N85);
or OR4 (N143, N142, N72, N125, N7);
nor NOR4 (N144, N138, N32, N143, N100);
buf BUF1 (N145, N87);
nor NOR4 (N146, N140, N143, N2, N102);
or OR4 (N147, N131, N110, N141, N16);
buf BUF1 (N148, N23);
not NOT1 (N149, N135);
and AND2 (N150, N144, N118);
nand NAND2 (N151, N133, N54);
and AND3 (N152, N145, N46, N99);
buf BUF1 (N153, N148);
or OR3 (N154, N146, N139, N67);
buf BUF1 (N155, N31);
buf BUF1 (N156, N153);
nand NAND4 (N157, N156, N11, N20, N49);
and AND3 (N158, N150, N50, N4);
xor XOR2 (N159, N158, N39);
xor XOR2 (N160, N147, N154);
nand NAND2 (N161, N62, N2);
and AND4 (N162, N152, N141, N36, N16);
nor NOR3 (N163, N162, N158, N11);
nand NAND4 (N164, N149, N72, N130, N87);
nand NAND2 (N165, N61, N57);
buf BUF1 (N166, N163);
not NOT1 (N167, N165);
not NOT1 (N168, N129);
and AND4 (N169, N159, N31, N113, N82);
not NOT1 (N170, N169);
buf BUF1 (N171, N166);
not NOT1 (N172, N151);
buf BUF1 (N173, N161);
xor XOR2 (N174, N164, N143);
or OR3 (N175, N172, N89, N69);
not NOT1 (N176, N171);
and AND2 (N177, N174, N84);
buf BUF1 (N178, N155);
or OR4 (N179, N175, N140, N177, N77);
not NOT1 (N180, N114);
nor NOR2 (N181, N178, N132);
or OR3 (N182, N160, N27, N54);
buf BUF1 (N183, N179);
not NOT1 (N184, N168);
nor NOR2 (N185, N170, N80);
buf BUF1 (N186, N173);
xor XOR2 (N187, N186, N141);
or OR3 (N188, N181, N187, N174);
buf BUF1 (N189, N23);
nor NOR2 (N190, N176, N180);
nand NAND4 (N191, N121, N133, N134, N64);
nand NAND2 (N192, N185, N77);
nor NOR4 (N193, N157, N139, N56, N128);
buf BUF1 (N194, N189);
and AND4 (N195, N188, N116, N51, N31);
xor XOR2 (N196, N190, N49);
nor NOR2 (N197, N184, N55);
and AND4 (N198, N182, N48, N64, N87);
xor XOR2 (N199, N167, N1);
or OR2 (N200, N199, N125);
nand NAND2 (N201, N196, N36);
buf BUF1 (N202, N192);
nand NAND3 (N203, N193, N168, N63);
nand NAND3 (N204, N198, N62, N110);
not NOT1 (N205, N183);
xor XOR2 (N206, N204, N199);
nand NAND2 (N207, N200, N103);
nand NAND3 (N208, N201, N130, N155);
or OR3 (N209, N203, N66, N166);
nand NAND2 (N210, N206, N4);
and AND3 (N211, N209, N151, N132);
or OR4 (N212, N202, N17, N197, N93);
nand NAND4 (N213, N159, N149, N210, N171);
or OR3 (N214, N84, N34, N206);
and AND4 (N215, N195, N62, N164, N90);
and AND4 (N216, N213, N8, N211, N118);
buf BUF1 (N217, N128);
nor NOR4 (N218, N207, N149, N87, N207);
xor XOR2 (N219, N208, N30);
xor XOR2 (N220, N218, N46);
or OR2 (N221, N217, N186);
nor NOR4 (N222, N215, N8, N124, N166);
not NOT1 (N223, N212);
nand NAND4 (N224, N214, N53, N33, N210);
nor NOR4 (N225, N223, N179, N149, N74);
or OR3 (N226, N205, N32, N192);
buf BUF1 (N227, N220);
not NOT1 (N228, N221);
xor XOR2 (N229, N224, N196);
xor XOR2 (N230, N226, N97);
and AND4 (N231, N191, N69, N64, N224);
nand NAND3 (N232, N216, N113, N209);
nand NAND2 (N233, N219, N130);
or OR4 (N234, N194, N193, N52, N57);
not NOT1 (N235, N225);
and AND2 (N236, N222, N5);
or OR2 (N237, N227, N123);
xor XOR2 (N238, N235, N19);
xor XOR2 (N239, N228, N42);
and AND4 (N240, N233, N230, N226, N49);
nor NOR2 (N241, N199, N10);
not NOT1 (N242, N240);
not NOT1 (N243, N236);
not NOT1 (N244, N232);
nand NAND2 (N245, N244, N50);
xor XOR2 (N246, N234, N110);
nor NOR2 (N247, N246, N25);
and AND4 (N248, N243, N11, N108, N15);
or OR3 (N249, N242, N109, N90);
nor NOR3 (N250, N237, N213, N241);
and AND4 (N251, N12, N214, N44, N234);
nand NAND4 (N252, N238, N173, N231, N197);
nand NAND2 (N253, N190, N238);
buf BUF1 (N254, N250);
buf BUF1 (N255, N247);
nand NAND2 (N256, N252, N201);
buf BUF1 (N257, N239);
and AND3 (N258, N253, N99, N223);
nand NAND3 (N259, N248, N172, N228);
xor XOR2 (N260, N258, N235);
and AND4 (N261, N260, N161, N163, N37);
not NOT1 (N262, N257);
nand NAND2 (N263, N256, N15);
xor XOR2 (N264, N251, N201);
buf BUF1 (N265, N264);
buf BUF1 (N266, N245);
nand NAND2 (N267, N229, N136);
not NOT1 (N268, N262);
not NOT1 (N269, N263);
nand NAND4 (N270, N261, N77, N57, N30);
buf BUF1 (N271, N249);
nand NAND4 (N272, N267, N100, N54, N34);
buf BUF1 (N273, N268);
not NOT1 (N274, N270);
and AND3 (N275, N269, N274, N226);
not NOT1 (N276, N77);
xor XOR2 (N277, N255, N252);
nor NOR3 (N278, N276, N110, N174);
and AND4 (N279, N271, N232, N28, N74);
buf BUF1 (N280, N278);
xor XOR2 (N281, N272, N65);
or OR4 (N282, N254, N221, N200, N245);
and AND3 (N283, N281, N133, N196);
xor XOR2 (N284, N265, N253);
nor NOR3 (N285, N275, N76, N69);
and AND2 (N286, N282, N32);
xor XOR2 (N287, N279, N202);
buf BUF1 (N288, N283);
buf BUF1 (N289, N280);
and AND4 (N290, N285, N225, N105, N270);
nor NOR3 (N291, N288, N195, N41);
and AND2 (N292, N291, N237);
xor XOR2 (N293, N286, N87);
not NOT1 (N294, N284);
nor NOR3 (N295, N273, N78, N232);
xor XOR2 (N296, N295, N186);
not NOT1 (N297, N259);
buf BUF1 (N298, N296);
buf BUF1 (N299, N277);
and AND3 (N300, N287, N281, N97);
xor XOR2 (N301, N292, N266);
not NOT1 (N302, N235);
xor XOR2 (N303, N290, N171);
xor XOR2 (N304, N301, N206);
and AND2 (N305, N297, N255);
not NOT1 (N306, N303);
or OR2 (N307, N298, N36);
xor XOR2 (N308, N294, N166);
and AND3 (N309, N289, N264, N50);
and AND3 (N310, N293, N94, N276);
or OR2 (N311, N305, N160);
nand NAND3 (N312, N299, N302, N280);
not NOT1 (N313, N85);
or OR3 (N314, N306, N86, N253);
nand NAND4 (N315, N311, N176, N95, N245);
xor XOR2 (N316, N315, N36);
and AND2 (N317, N310, N184);
not NOT1 (N318, N314);
xor XOR2 (N319, N309, N64);
buf BUF1 (N320, N318);
endmodule