// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21;

output N3005,N3007,N3015,N2996,N3014,N3019,N2995,N3020,N3017,N3021;

and AND3 (N22, N4, N3, N13);
xor XOR2 (N23, N18, N6);
nand NAND2 (N24, N13, N1);
and AND4 (N25, N18, N14, N1, N21);
or OR2 (N26, N6, N12);
nand NAND2 (N27, N14, N17);
or OR2 (N28, N6, N5);
xor XOR2 (N29, N3, N2);
nand NAND2 (N30, N3, N22);
not NOT1 (N31, N22);
nand NAND3 (N32, N10, N27, N11);
nor NOR3 (N33, N14, N11, N15);
and AND4 (N34, N32, N16, N24, N6);
buf BUF1 (N35, N7);
not NOT1 (N36, N30);
nand NAND4 (N37, N26, N22, N24, N25);
or OR3 (N38, N15, N29, N29);
xor XOR2 (N39, N9, N34);
nand NAND2 (N40, N1, N16);
nor NOR3 (N41, N37, N2, N36);
not NOT1 (N42, N2);
not NOT1 (N43, N31);
xor XOR2 (N44, N41, N26);
nand NAND2 (N45, N39, N8);
nand NAND3 (N46, N44, N43, N27);
nand NAND3 (N47, N36, N25, N42);
and AND4 (N48, N30, N27, N19, N36);
nand NAND2 (N49, N33, N5);
buf BUF1 (N50, N23);
nor NOR2 (N51, N49, N49);
nor NOR4 (N52, N35, N7, N26, N42);
and AND3 (N53, N47, N7, N42);
buf BUF1 (N54, N38);
not NOT1 (N55, N50);
and AND3 (N56, N53, N20, N5);
nor NOR4 (N57, N55, N37, N31, N18);
or OR4 (N58, N46, N48, N44, N15);
nor NOR4 (N59, N8, N14, N42, N58);
buf BUF1 (N60, N35);
nand NAND3 (N61, N28, N26, N52);
nor NOR2 (N62, N29, N44);
xor XOR2 (N63, N51, N19);
buf BUF1 (N64, N63);
buf BUF1 (N65, N60);
buf BUF1 (N66, N59);
buf BUF1 (N67, N40);
and AND2 (N68, N65, N8);
not NOT1 (N69, N45);
nor NOR3 (N70, N57, N50, N1);
not NOT1 (N71, N62);
buf BUF1 (N72, N54);
and AND4 (N73, N69, N44, N65, N29);
nand NAND3 (N74, N64, N27, N2);
buf BUF1 (N75, N66);
nor NOR4 (N76, N73, N55, N33, N44);
and AND4 (N77, N67, N52, N62, N63);
xor XOR2 (N78, N61, N22);
and AND2 (N79, N68, N54);
buf BUF1 (N80, N72);
and AND4 (N81, N71, N48, N46, N78);
or OR2 (N82, N36, N24);
or OR2 (N83, N76, N63);
xor XOR2 (N84, N56, N28);
xor XOR2 (N85, N75, N21);
nor NOR3 (N86, N85, N78, N17);
and AND3 (N87, N80, N59, N57);
nor NOR2 (N88, N86, N36);
xor XOR2 (N89, N82, N73);
buf BUF1 (N90, N89);
not NOT1 (N91, N74);
not NOT1 (N92, N81);
xor XOR2 (N93, N88, N30);
and AND2 (N94, N92, N9);
nor NOR4 (N95, N84, N7, N6, N11);
buf BUF1 (N96, N95);
or OR4 (N97, N90, N12, N37, N31);
buf BUF1 (N98, N91);
buf BUF1 (N99, N96);
xor XOR2 (N100, N98, N62);
xor XOR2 (N101, N93, N31);
buf BUF1 (N102, N101);
xor XOR2 (N103, N77, N66);
nor NOR3 (N104, N70, N18, N53);
nor NOR3 (N105, N104, N29, N6);
and AND2 (N106, N102, N63);
nor NOR3 (N107, N100, N70, N61);
nor NOR2 (N108, N79, N83);
and AND4 (N109, N5, N84, N61, N5);
not NOT1 (N110, N99);
nand NAND4 (N111, N103, N50, N84, N15);
or OR4 (N112, N109, N24, N89, N109);
xor XOR2 (N113, N110, N27);
or OR4 (N114, N111, N63, N6, N11);
or OR2 (N115, N87, N105);
not NOT1 (N116, N40);
and AND2 (N117, N107, N31);
buf BUF1 (N118, N112);
nor NOR3 (N119, N114, N29, N36);
nand NAND2 (N120, N113, N61);
nor NOR2 (N121, N97, N36);
or OR3 (N122, N121, N83, N30);
not NOT1 (N123, N117);
xor XOR2 (N124, N94, N71);
or OR2 (N125, N124, N96);
not NOT1 (N126, N106);
nand NAND4 (N127, N123, N41, N100, N88);
nand NAND3 (N128, N116, N17, N9);
not NOT1 (N129, N115);
xor XOR2 (N130, N126, N103);
and AND3 (N131, N129, N61, N123);
nand NAND4 (N132, N128, N121, N69, N31);
not NOT1 (N133, N132);
xor XOR2 (N134, N130, N119);
and AND2 (N135, N132, N84);
buf BUF1 (N136, N127);
buf BUF1 (N137, N122);
xor XOR2 (N138, N125, N70);
and AND2 (N139, N135, N103);
nand NAND4 (N140, N134, N27, N3, N60);
nand NAND2 (N141, N120, N64);
and AND2 (N142, N140, N1);
xor XOR2 (N143, N118, N8);
nand NAND2 (N144, N141, N109);
nor NOR3 (N145, N133, N101, N33);
nor NOR3 (N146, N138, N22, N117);
or OR3 (N147, N108, N138, N92);
not NOT1 (N148, N143);
buf BUF1 (N149, N148);
nor NOR4 (N150, N142, N65, N139, N30);
nand NAND4 (N151, N107, N23, N103, N110);
or OR3 (N152, N149, N21, N20);
nor NOR4 (N153, N151, N29, N151, N101);
or OR4 (N154, N152, N56, N37, N34);
and AND4 (N155, N153, N11, N105, N46);
not NOT1 (N156, N146);
and AND3 (N157, N154, N19, N63);
or OR2 (N158, N144, N18);
xor XOR2 (N159, N145, N79);
or OR2 (N160, N157, N71);
nand NAND2 (N161, N136, N20);
not NOT1 (N162, N155);
nand NAND2 (N163, N158, N125);
xor XOR2 (N164, N131, N163);
and AND3 (N165, N65, N161, N58);
not NOT1 (N166, N123);
not NOT1 (N167, N164);
nor NOR2 (N168, N162, N15);
or OR3 (N169, N150, N110, N140);
or OR2 (N170, N159, N21);
and AND2 (N171, N160, N114);
and AND2 (N172, N165, N111);
not NOT1 (N173, N147);
or OR4 (N174, N156, N46, N103, N37);
not NOT1 (N175, N172);
or OR2 (N176, N137, N159);
nor NOR4 (N177, N167, N122, N127, N74);
nand NAND4 (N178, N171, N157, N170, N52);
nand NAND3 (N179, N63, N26, N75);
nor NOR2 (N180, N168, N135);
and AND2 (N181, N179, N129);
and AND2 (N182, N174, N77);
and AND4 (N183, N181, N26, N24, N162);
nand NAND4 (N184, N175, N56, N123, N24);
nand NAND3 (N185, N169, N138, N145);
nor NOR2 (N186, N183, N108);
nand NAND3 (N187, N180, N78, N24);
or OR2 (N188, N185, N173);
and AND3 (N189, N153, N59, N179);
not NOT1 (N190, N178);
nand NAND2 (N191, N184, N85);
nor NOR4 (N192, N187, N102, N121, N28);
and AND4 (N193, N189, N150, N19, N62);
not NOT1 (N194, N193);
nand NAND4 (N195, N191, N171, N31, N84);
and AND2 (N196, N188, N37);
buf BUF1 (N197, N195);
and AND4 (N198, N166, N173, N147, N106);
nor NOR2 (N199, N198, N92);
nand NAND4 (N200, N199, N8, N28, N66);
or OR3 (N201, N182, N123, N172);
nand NAND2 (N202, N201, N132);
and AND3 (N203, N186, N150, N14);
or OR2 (N204, N200, N9);
nand NAND2 (N205, N190, N101);
not NOT1 (N206, N194);
nor NOR2 (N207, N203, N53);
nand NAND2 (N208, N176, N6);
nand NAND4 (N209, N197, N186, N126, N96);
buf BUF1 (N210, N192);
nand NAND2 (N211, N196, N120);
and AND4 (N212, N204, N208, N51, N30);
not NOT1 (N213, N116);
nand NAND2 (N214, N207, N26);
buf BUF1 (N215, N210);
nor NOR2 (N216, N206, N184);
and AND4 (N217, N214, N146, N160, N113);
nor NOR3 (N218, N177, N119, N32);
and AND2 (N219, N218, N138);
xor XOR2 (N220, N219, N74);
not NOT1 (N221, N202);
xor XOR2 (N222, N211, N210);
buf BUF1 (N223, N212);
nor NOR2 (N224, N209, N90);
nand NAND3 (N225, N205, N138, N157);
not NOT1 (N226, N217);
not NOT1 (N227, N223);
nand NAND4 (N228, N213, N128, N57, N27);
not NOT1 (N229, N226);
or OR2 (N230, N220, N133);
nor NOR4 (N231, N229, N121, N127, N121);
buf BUF1 (N232, N215);
nand NAND2 (N233, N221, N145);
buf BUF1 (N234, N232);
nor NOR2 (N235, N227, N122);
and AND2 (N236, N233, N168);
xor XOR2 (N237, N235, N107);
xor XOR2 (N238, N231, N120);
buf BUF1 (N239, N224);
and AND3 (N240, N236, N24, N65);
xor XOR2 (N241, N234, N96);
buf BUF1 (N242, N222);
and AND2 (N243, N230, N36);
xor XOR2 (N244, N243, N43);
nand NAND2 (N245, N237, N218);
and AND3 (N246, N241, N163, N128);
or OR3 (N247, N216, N8, N105);
not NOT1 (N248, N238);
and AND4 (N249, N239, N86, N216, N91);
or OR4 (N250, N247, N218, N246, N242);
nand NAND4 (N251, N94, N136, N151, N49);
buf BUF1 (N252, N202);
xor XOR2 (N253, N248, N230);
or OR2 (N254, N249, N158);
and AND4 (N255, N240, N65, N217, N4);
and AND3 (N256, N254, N21, N57);
nor NOR2 (N257, N245, N83);
not NOT1 (N258, N253);
xor XOR2 (N259, N257, N30);
nor NOR2 (N260, N251, N104);
nand NAND3 (N261, N258, N231, N209);
xor XOR2 (N262, N261, N209);
and AND3 (N263, N259, N19, N126);
nand NAND3 (N264, N228, N82, N258);
nor NOR2 (N265, N263, N52);
nand NAND4 (N266, N260, N6, N121, N83);
and AND4 (N267, N264, N135, N159, N58);
not NOT1 (N268, N252);
xor XOR2 (N269, N265, N9);
not NOT1 (N270, N255);
not NOT1 (N271, N270);
nand NAND2 (N272, N250, N270);
not NOT1 (N273, N267);
nor NOR4 (N274, N271, N267, N253, N187);
buf BUF1 (N275, N272);
and AND3 (N276, N268, N266, N223);
xor XOR2 (N277, N229, N248);
nand NAND4 (N278, N275, N128, N275, N104);
not NOT1 (N279, N262);
not NOT1 (N280, N274);
and AND3 (N281, N225, N68, N271);
buf BUF1 (N282, N279);
or OR2 (N283, N269, N4);
not NOT1 (N284, N256);
nand NAND3 (N285, N283, N264, N70);
nor NOR2 (N286, N244, N268);
nor NOR4 (N287, N273, N152, N49, N13);
buf BUF1 (N288, N276);
nand NAND2 (N289, N288, N182);
buf BUF1 (N290, N286);
nand NAND2 (N291, N278, N209);
xor XOR2 (N292, N281, N211);
nand NAND3 (N293, N277, N165, N204);
and AND3 (N294, N292, N157, N256);
and AND2 (N295, N290, N284);
buf BUF1 (N296, N42);
nand NAND4 (N297, N280, N280, N61, N87);
nor NOR3 (N298, N295, N247, N57);
xor XOR2 (N299, N282, N34);
nor NOR3 (N300, N296, N179, N288);
buf BUF1 (N301, N291);
nor NOR4 (N302, N297, N106, N139, N159);
not NOT1 (N303, N285);
nor NOR4 (N304, N298, N167, N141, N276);
and AND4 (N305, N302, N121, N120, N77);
nand NAND2 (N306, N294, N115);
buf BUF1 (N307, N301);
not NOT1 (N308, N304);
not NOT1 (N309, N300);
buf BUF1 (N310, N287);
buf BUF1 (N311, N306);
not NOT1 (N312, N305);
or OR3 (N313, N307, N182, N211);
and AND4 (N314, N309, N306, N195, N133);
not NOT1 (N315, N311);
buf BUF1 (N316, N308);
xor XOR2 (N317, N316, N224);
nor NOR3 (N318, N289, N268, N108);
and AND2 (N319, N293, N98);
or OR3 (N320, N318, N190, N59);
nand NAND2 (N321, N310, N152);
not NOT1 (N322, N319);
xor XOR2 (N323, N299, N168);
or OR4 (N324, N312, N290, N49, N279);
buf BUF1 (N325, N313);
nor NOR3 (N326, N324, N127, N17);
xor XOR2 (N327, N314, N154);
nor NOR2 (N328, N315, N12);
nand NAND4 (N329, N322, N93, N18, N50);
nand NAND4 (N330, N320, N60, N116, N19);
nand NAND2 (N331, N303, N79);
and AND4 (N332, N325, N86, N299, N189);
nand NAND2 (N333, N323, N179);
buf BUF1 (N334, N333);
buf BUF1 (N335, N329);
nor NOR4 (N336, N331, N180, N72, N87);
and AND2 (N337, N335, N168);
nor NOR4 (N338, N328, N239, N45, N21);
buf BUF1 (N339, N321);
nand NAND2 (N340, N334, N47);
or OR4 (N341, N336, N338, N142, N155);
or OR3 (N342, N321, N221, N13);
and AND2 (N343, N326, N191);
nand NAND3 (N344, N339, N173, N296);
nor NOR3 (N345, N337, N54, N163);
or OR2 (N346, N330, N168);
nand NAND2 (N347, N343, N2);
or OR4 (N348, N344, N217, N183, N144);
nand NAND2 (N349, N317, N156);
nand NAND4 (N350, N342, N18, N78, N94);
xor XOR2 (N351, N346, N207);
nor NOR3 (N352, N348, N231, N147);
nand NAND4 (N353, N347, N266, N41, N150);
or OR3 (N354, N345, N239, N202);
not NOT1 (N355, N352);
and AND2 (N356, N332, N106);
or OR2 (N357, N349, N163);
or OR4 (N358, N354, N187, N110, N21);
or OR3 (N359, N358, N53, N342);
and AND2 (N360, N353, N333);
nor NOR2 (N361, N340, N266);
nor NOR2 (N362, N357, N330);
nor NOR3 (N363, N355, N237, N228);
and AND2 (N364, N361, N49);
buf BUF1 (N365, N364);
and AND4 (N366, N327, N229, N232, N186);
and AND2 (N367, N351, N115);
nand NAND4 (N368, N362, N213, N83, N307);
not NOT1 (N369, N363);
buf BUF1 (N370, N369);
buf BUF1 (N371, N341);
nand NAND2 (N372, N356, N107);
buf BUF1 (N373, N367);
buf BUF1 (N374, N370);
buf BUF1 (N375, N371);
nor NOR3 (N376, N366, N211, N222);
buf BUF1 (N377, N368);
and AND2 (N378, N359, N123);
nor NOR2 (N379, N373, N375);
nand NAND2 (N380, N292, N40);
nand NAND3 (N381, N350, N373, N132);
or OR2 (N382, N360, N97);
not NOT1 (N383, N374);
and AND3 (N384, N382, N197, N76);
nand NAND4 (N385, N384, N97, N143, N285);
buf BUF1 (N386, N385);
xor XOR2 (N387, N377, N27);
xor XOR2 (N388, N381, N214);
buf BUF1 (N389, N376);
xor XOR2 (N390, N372, N168);
buf BUF1 (N391, N390);
nor NOR2 (N392, N365, N294);
or OR3 (N393, N386, N241, N45);
nor NOR2 (N394, N393, N76);
buf BUF1 (N395, N392);
xor XOR2 (N396, N383, N106);
or OR4 (N397, N396, N175, N96, N379);
nand NAND3 (N398, N274, N20, N40);
not NOT1 (N399, N391);
or OR3 (N400, N394, N152, N344);
or OR3 (N401, N400, N120, N341);
or OR2 (N402, N399, N42);
nand NAND3 (N403, N402, N142, N348);
or OR3 (N404, N387, N220, N5);
xor XOR2 (N405, N380, N15);
not NOT1 (N406, N404);
buf BUF1 (N407, N389);
not NOT1 (N408, N406);
xor XOR2 (N409, N395, N169);
buf BUF1 (N410, N407);
xor XOR2 (N411, N378, N384);
nor NOR4 (N412, N411, N330, N273, N181);
and AND4 (N413, N397, N308, N93, N75);
xor XOR2 (N414, N413, N411);
xor XOR2 (N415, N412, N288);
buf BUF1 (N416, N403);
or OR2 (N417, N409, N342);
nor NOR3 (N418, N416, N208, N18);
nor NOR4 (N419, N417, N114, N200, N339);
nor NOR3 (N420, N408, N57, N224);
nand NAND4 (N421, N401, N365, N55, N91);
nand NAND3 (N422, N420, N198, N17);
or OR2 (N423, N419, N131);
nand NAND4 (N424, N418, N268, N24, N42);
xor XOR2 (N425, N388, N35);
not NOT1 (N426, N421);
buf BUF1 (N427, N424);
xor XOR2 (N428, N410, N341);
nor NOR2 (N429, N425, N139);
and AND3 (N430, N427, N81, N260);
not NOT1 (N431, N415);
nor NOR3 (N432, N414, N288, N55);
or OR3 (N433, N422, N139, N348);
buf BUF1 (N434, N398);
and AND3 (N435, N431, N391, N183);
and AND3 (N436, N434, N406, N384);
nand NAND3 (N437, N436, N402, N387);
buf BUF1 (N438, N428);
buf BUF1 (N439, N432);
or OR4 (N440, N439, N329, N142, N364);
xor XOR2 (N441, N437, N315);
or OR3 (N442, N429, N224, N214);
not NOT1 (N443, N435);
or OR2 (N444, N443, N268);
not NOT1 (N445, N430);
nand NAND2 (N446, N445, N4);
or OR3 (N447, N442, N120, N445);
xor XOR2 (N448, N405, N229);
xor XOR2 (N449, N438, N198);
or OR2 (N450, N447, N266);
nand NAND4 (N451, N444, N81, N357, N45);
not NOT1 (N452, N446);
not NOT1 (N453, N440);
or OR2 (N454, N451, N388);
nor NOR4 (N455, N423, N161, N221, N127);
nor NOR2 (N456, N455, N60);
or OR4 (N457, N450, N387, N145, N182);
and AND4 (N458, N456, N249, N230, N12);
nand NAND3 (N459, N458, N282, N284);
nand NAND4 (N460, N459, N113, N57, N241);
buf BUF1 (N461, N449);
buf BUF1 (N462, N460);
and AND4 (N463, N448, N223, N357, N360);
and AND2 (N464, N441, N335);
buf BUF1 (N465, N463);
xor XOR2 (N466, N453, N264);
buf BUF1 (N467, N457);
nor NOR2 (N468, N462, N253);
xor XOR2 (N469, N468, N105);
not NOT1 (N470, N465);
nand NAND2 (N471, N433, N468);
xor XOR2 (N472, N470, N441);
and AND2 (N473, N426, N23);
nor NOR3 (N474, N452, N342, N339);
nand NAND3 (N475, N474, N266, N1);
not NOT1 (N476, N467);
or OR3 (N477, N471, N45, N30);
and AND2 (N478, N461, N390);
and AND4 (N479, N473, N55, N342, N60);
nor NOR2 (N480, N477, N440);
not NOT1 (N481, N476);
and AND3 (N482, N475, N11, N202);
buf BUF1 (N483, N479);
or OR4 (N484, N478, N361, N75, N360);
nor NOR4 (N485, N480, N229, N386, N403);
and AND2 (N486, N466, N482);
xor XOR2 (N487, N253, N9);
nand NAND2 (N488, N486, N90);
nor NOR4 (N489, N484, N170, N352, N132);
or OR4 (N490, N485, N242, N25, N359);
not NOT1 (N491, N481);
or OR2 (N492, N489, N74);
xor XOR2 (N493, N483, N30);
and AND3 (N494, N490, N210, N11);
buf BUF1 (N495, N488);
not NOT1 (N496, N469);
xor XOR2 (N497, N494, N176);
xor XOR2 (N498, N495, N246);
or OR4 (N499, N492, N481, N457, N342);
or OR4 (N500, N487, N104, N106, N75);
xor XOR2 (N501, N493, N204);
xor XOR2 (N502, N491, N163);
nor NOR2 (N503, N499, N136);
xor XOR2 (N504, N501, N413);
and AND2 (N505, N503, N474);
and AND2 (N506, N464, N346);
buf BUF1 (N507, N497);
xor XOR2 (N508, N502, N117);
or OR3 (N509, N505, N103, N277);
not NOT1 (N510, N472);
nand NAND4 (N511, N504, N310, N388, N414);
buf BUF1 (N512, N498);
buf BUF1 (N513, N508);
buf BUF1 (N514, N496);
nand NAND4 (N515, N513, N454, N50, N368);
not NOT1 (N516, N270);
not NOT1 (N517, N516);
nand NAND3 (N518, N514, N296, N366);
buf BUF1 (N519, N517);
and AND3 (N520, N510, N150, N465);
nor NOR4 (N521, N507, N49, N396, N129);
nor NOR2 (N522, N518, N13);
and AND3 (N523, N519, N214, N319);
xor XOR2 (N524, N512, N72);
buf BUF1 (N525, N522);
not NOT1 (N526, N525);
buf BUF1 (N527, N509);
nand NAND2 (N528, N526, N194);
buf BUF1 (N529, N500);
xor XOR2 (N530, N523, N90);
and AND4 (N531, N520, N513, N147, N99);
nor NOR4 (N532, N530, N239, N499, N507);
buf BUF1 (N533, N527);
not NOT1 (N534, N528);
nor NOR2 (N535, N529, N75);
buf BUF1 (N536, N533);
or OR2 (N537, N536, N499);
or OR4 (N538, N532, N18, N195, N168);
and AND4 (N539, N521, N145, N7, N469);
and AND4 (N540, N538, N1, N355, N471);
nand NAND2 (N541, N534, N473);
nor NOR4 (N542, N541, N187, N359, N339);
nor NOR4 (N543, N531, N78, N29, N485);
and AND2 (N544, N537, N109);
or OR3 (N545, N543, N103, N382);
or OR3 (N546, N511, N309, N123);
and AND3 (N547, N546, N10, N111);
not NOT1 (N548, N539);
nand NAND4 (N549, N548, N406, N85, N4);
nand NAND2 (N550, N547, N429);
buf BUF1 (N551, N550);
xor XOR2 (N552, N515, N100);
xor XOR2 (N553, N542, N384);
or OR2 (N554, N551, N187);
xor XOR2 (N555, N544, N207);
not NOT1 (N556, N535);
or OR4 (N557, N554, N34, N523, N66);
or OR3 (N558, N540, N1, N226);
nor NOR3 (N559, N558, N283, N90);
buf BUF1 (N560, N556);
not NOT1 (N561, N557);
nand NAND2 (N562, N553, N513);
not NOT1 (N563, N549);
and AND4 (N564, N524, N497, N154, N204);
xor XOR2 (N565, N555, N317);
nor NOR2 (N566, N561, N284);
nor NOR4 (N567, N566, N456, N555, N221);
buf BUF1 (N568, N560);
or OR3 (N569, N506, N364, N389);
and AND3 (N570, N562, N421, N82);
nor NOR3 (N571, N565, N457, N128);
not NOT1 (N572, N570);
buf BUF1 (N573, N572);
or OR4 (N574, N564, N449, N349, N325);
or OR3 (N575, N573, N264, N18);
buf BUF1 (N576, N559);
nand NAND4 (N577, N569, N355, N154, N155);
buf BUF1 (N578, N571);
nor NOR4 (N579, N563, N275, N393, N188);
nor NOR3 (N580, N578, N133, N380);
nand NAND3 (N581, N577, N143, N253);
buf BUF1 (N582, N552);
nand NAND2 (N583, N545, N409);
nor NOR2 (N584, N579, N535);
nor NOR2 (N585, N580, N237);
nand NAND4 (N586, N567, N237, N377, N529);
not NOT1 (N587, N583);
xor XOR2 (N588, N586, N162);
buf BUF1 (N589, N585);
not NOT1 (N590, N568);
buf BUF1 (N591, N575);
nor NOR3 (N592, N590, N140, N481);
buf BUF1 (N593, N576);
or OR3 (N594, N584, N147, N295);
nor NOR2 (N595, N588, N576);
xor XOR2 (N596, N587, N47);
nor NOR4 (N597, N582, N461, N126, N178);
nor NOR3 (N598, N597, N451, N509);
and AND2 (N599, N595, N145);
or OR3 (N600, N592, N402, N442);
and AND4 (N601, N596, N470, N228, N99);
buf BUF1 (N602, N601);
and AND4 (N603, N598, N372, N153, N98);
nand NAND4 (N604, N599, N182, N523, N130);
xor XOR2 (N605, N594, N100);
and AND3 (N606, N604, N383, N235);
or OR4 (N607, N602, N532, N145, N105);
not NOT1 (N608, N591);
not NOT1 (N609, N574);
buf BUF1 (N610, N593);
not NOT1 (N611, N609);
or OR2 (N612, N581, N146);
and AND4 (N613, N607, N124, N593, N366);
xor XOR2 (N614, N589, N223);
not NOT1 (N615, N614);
buf BUF1 (N616, N615);
and AND2 (N617, N616, N565);
nand NAND2 (N618, N611, N533);
nor NOR2 (N619, N610, N171);
or OR3 (N620, N618, N533, N59);
nand NAND3 (N621, N608, N545, N19);
or OR4 (N622, N620, N66, N121, N605);
nor NOR2 (N623, N485, N37);
xor XOR2 (N624, N600, N396);
nor NOR2 (N625, N603, N225);
buf BUF1 (N626, N617);
and AND2 (N627, N626, N241);
xor XOR2 (N628, N624, N172);
buf BUF1 (N629, N627);
or OR3 (N630, N628, N254, N626);
or OR4 (N631, N623, N383, N444, N330);
and AND4 (N632, N631, N94, N28, N130);
nand NAND2 (N633, N613, N609);
or OR2 (N634, N630, N171);
nand NAND4 (N635, N634, N259, N534, N49);
or OR2 (N636, N622, N51);
nand NAND2 (N637, N629, N262);
xor XOR2 (N638, N612, N470);
not NOT1 (N639, N606);
and AND3 (N640, N635, N367, N27);
or OR2 (N641, N636, N400);
or OR2 (N642, N633, N559);
and AND3 (N643, N621, N43, N249);
nand NAND3 (N644, N619, N632, N52);
nand NAND4 (N645, N328, N135, N82, N88);
or OR4 (N646, N641, N302, N402, N328);
xor XOR2 (N647, N646, N39);
xor XOR2 (N648, N647, N221);
nor NOR4 (N649, N648, N557, N236, N68);
nor NOR3 (N650, N625, N479, N356);
xor XOR2 (N651, N642, N511);
or OR4 (N652, N649, N42, N631, N471);
nor NOR4 (N653, N639, N407, N477, N586);
nor NOR3 (N654, N645, N15, N215);
xor XOR2 (N655, N644, N284);
not NOT1 (N656, N643);
nand NAND4 (N657, N650, N392, N389, N390);
and AND2 (N658, N654, N558);
xor XOR2 (N659, N640, N451);
or OR3 (N660, N659, N146, N177);
xor XOR2 (N661, N652, N214);
nor NOR4 (N662, N657, N51, N141, N519);
nand NAND4 (N663, N651, N523, N590, N36);
buf BUF1 (N664, N662);
nor NOR3 (N665, N663, N656, N615);
nand NAND4 (N666, N471, N190, N382, N497);
and AND4 (N667, N665, N221, N601, N47);
and AND4 (N668, N658, N143, N336, N382);
or OR2 (N669, N638, N590);
nand NAND2 (N670, N667, N487);
nand NAND3 (N671, N653, N565, N146);
not NOT1 (N672, N670);
or OR3 (N673, N664, N320, N575);
not NOT1 (N674, N661);
not NOT1 (N675, N666);
not NOT1 (N676, N655);
nand NAND4 (N677, N674, N47, N73, N589);
xor XOR2 (N678, N676, N255);
not NOT1 (N679, N671);
nor NOR3 (N680, N679, N539, N307);
not NOT1 (N681, N673);
xor XOR2 (N682, N677, N482);
nand NAND4 (N683, N637, N529, N187, N574);
nor NOR2 (N684, N669, N96);
xor XOR2 (N685, N660, N632);
nor NOR4 (N686, N672, N421, N144, N455);
buf BUF1 (N687, N685);
nor NOR3 (N688, N668, N21, N254);
buf BUF1 (N689, N681);
not NOT1 (N690, N680);
or OR3 (N691, N690, N333, N177);
nand NAND4 (N692, N691, N25, N381, N315);
or OR3 (N693, N686, N239, N50);
nand NAND4 (N694, N682, N521, N185, N644);
buf BUF1 (N695, N683);
nand NAND4 (N696, N687, N222, N248, N236);
nand NAND3 (N697, N696, N664, N473);
xor XOR2 (N698, N688, N60);
not NOT1 (N699, N695);
nand NAND4 (N700, N694, N227, N105, N440);
nor NOR4 (N701, N675, N411, N42, N364);
buf BUF1 (N702, N699);
xor XOR2 (N703, N702, N702);
and AND3 (N704, N703, N38, N435);
or OR2 (N705, N701, N234);
nor NOR3 (N706, N684, N97, N292);
not NOT1 (N707, N700);
nor NOR4 (N708, N697, N550, N567, N320);
xor XOR2 (N709, N706, N221);
nor NOR3 (N710, N707, N94, N167);
buf BUF1 (N711, N705);
and AND4 (N712, N693, N548, N376, N74);
not NOT1 (N713, N709);
nand NAND2 (N714, N711, N32);
nor NOR2 (N715, N713, N558);
and AND4 (N716, N708, N694, N294, N453);
and AND4 (N717, N692, N598, N254, N215);
not NOT1 (N718, N712);
or OR4 (N719, N715, N594, N387, N604);
xor XOR2 (N720, N717, N236);
not NOT1 (N721, N698);
not NOT1 (N722, N716);
or OR4 (N723, N678, N156, N614, N644);
and AND3 (N724, N720, N212, N344);
buf BUF1 (N725, N723);
or OR3 (N726, N704, N143, N331);
xor XOR2 (N727, N689, N657);
buf BUF1 (N728, N722);
buf BUF1 (N729, N721);
buf BUF1 (N730, N727);
buf BUF1 (N731, N724);
or OR2 (N732, N730, N597);
and AND3 (N733, N732, N187, N240);
not NOT1 (N734, N718);
not NOT1 (N735, N733);
nand NAND4 (N736, N731, N415, N49, N166);
or OR2 (N737, N728, N138);
not NOT1 (N738, N719);
and AND2 (N739, N710, N41);
buf BUF1 (N740, N739);
not NOT1 (N741, N726);
buf BUF1 (N742, N740);
xor XOR2 (N743, N734, N396);
not NOT1 (N744, N714);
not NOT1 (N745, N742);
or OR3 (N746, N744, N133, N213);
not NOT1 (N747, N745);
and AND3 (N748, N725, N119, N244);
xor XOR2 (N749, N741, N410);
or OR3 (N750, N736, N119, N612);
nor NOR2 (N751, N738, N97);
nor NOR2 (N752, N750, N563);
or OR2 (N753, N743, N161);
and AND4 (N754, N737, N718, N609, N531);
not NOT1 (N755, N751);
not NOT1 (N756, N747);
nor NOR2 (N757, N753, N571);
not NOT1 (N758, N756);
xor XOR2 (N759, N748, N151);
or OR2 (N760, N755, N605);
nor NOR2 (N761, N759, N588);
nor NOR4 (N762, N758, N632, N138, N214);
not NOT1 (N763, N757);
and AND3 (N764, N754, N134, N281);
nor NOR3 (N765, N749, N559, N90);
and AND4 (N766, N735, N199, N113, N191);
xor XOR2 (N767, N762, N606);
xor XOR2 (N768, N767, N599);
not NOT1 (N769, N766);
nand NAND2 (N770, N760, N81);
and AND4 (N771, N763, N5, N541, N316);
buf BUF1 (N772, N746);
and AND3 (N773, N769, N50, N319);
nor NOR3 (N774, N765, N600, N725);
and AND3 (N775, N772, N760, N583);
or OR4 (N776, N768, N28, N134, N418);
xor XOR2 (N777, N774, N42);
not NOT1 (N778, N775);
buf BUF1 (N779, N776);
and AND3 (N780, N779, N395, N772);
not NOT1 (N781, N761);
or OR3 (N782, N778, N107, N463);
xor XOR2 (N783, N781, N215);
nand NAND2 (N784, N771, N318);
buf BUF1 (N785, N729);
xor XOR2 (N786, N773, N47);
buf BUF1 (N787, N770);
nand NAND3 (N788, N780, N250, N311);
and AND2 (N789, N764, N273);
not NOT1 (N790, N782);
or OR2 (N791, N785, N109);
and AND3 (N792, N784, N616, N674);
or OR4 (N793, N788, N300, N164, N110);
and AND2 (N794, N793, N50);
buf BUF1 (N795, N777);
xor XOR2 (N796, N794, N435);
buf BUF1 (N797, N790);
nor NOR3 (N798, N752, N772, N644);
not NOT1 (N799, N787);
xor XOR2 (N800, N797, N662);
and AND3 (N801, N786, N635, N641);
not NOT1 (N802, N801);
xor XOR2 (N803, N800, N657);
not NOT1 (N804, N791);
buf BUF1 (N805, N798);
xor XOR2 (N806, N783, N107);
nor NOR2 (N807, N805, N709);
xor XOR2 (N808, N807, N756);
and AND2 (N809, N795, N461);
buf BUF1 (N810, N808);
xor XOR2 (N811, N796, N138);
or OR2 (N812, N802, N390);
nand NAND2 (N813, N803, N771);
and AND3 (N814, N799, N380, N428);
nor NOR3 (N815, N804, N353, N586);
xor XOR2 (N816, N806, N547);
and AND3 (N817, N810, N387, N16);
nor NOR4 (N818, N814, N189, N315, N405);
and AND4 (N819, N809, N190, N184, N38);
or OR2 (N820, N811, N689);
nand NAND2 (N821, N813, N56);
xor XOR2 (N822, N789, N650);
nor NOR4 (N823, N819, N221, N142, N300);
xor XOR2 (N824, N821, N417);
xor XOR2 (N825, N812, N382);
buf BUF1 (N826, N816);
or OR2 (N827, N815, N79);
or OR2 (N828, N822, N385);
or OR4 (N829, N826, N594, N431, N169);
nor NOR2 (N830, N829, N186);
buf BUF1 (N831, N823);
nor NOR3 (N832, N824, N122, N432);
and AND4 (N833, N792, N270, N301, N536);
buf BUF1 (N834, N828);
buf BUF1 (N835, N832);
not NOT1 (N836, N827);
nor NOR2 (N837, N825, N613);
xor XOR2 (N838, N818, N65);
xor XOR2 (N839, N817, N13);
nand NAND2 (N840, N834, N105);
xor XOR2 (N841, N838, N811);
and AND2 (N842, N836, N91);
not NOT1 (N843, N833);
and AND3 (N844, N842, N625, N817);
nand NAND3 (N845, N830, N716, N282);
nor NOR2 (N846, N844, N493);
buf BUF1 (N847, N845);
and AND4 (N848, N837, N157, N722, N296);
not NOT1 (N849, N820);
and AND3 (N850, N840, N623, N462);
nand NAND4 (N851, N841, N163, N489, N15);
and AND2 (N852, N849, N418);
buf BUF1 (N853, N835);
or OR2 (N854, N850, N759);
or OR3 (N855, N853, N93, N403);
nor NOR2 (N856, N854, N184);
nor NOR2 (N857, N851, N39);
buf BUF1 (N858, N839);
or OR4 (N859, N852, N529, N440, N431);
nor NOR3 (N860, N847, N838, N36);
or OR4 (N861, N831, N826, N202, N434);
buf BUF1 (N862, N857);
xor XOR2 (N863, N846, N59);
xor XOR2 (N864, N861, N796);
nand NAND2 (N865, N859, N815);
buf BUF1 (N866, N855);
nand NAND2 (N867, N863, N522);
buf BUF1 (N868, N864);
buf BUF1 (N869, N866);
and AND2 (N870, N868, N694);
nor NOR4 (N871, N860, N330, N16, N739);
nand NAND4 (N872, N865, N69, N308, N125);
nand NAND2 (N873, N843, N603);
or OR4 (N874, N858, N65, N691, N17);
not NOT1 (N875, N862);
buf BUF1 (N876, N875);
or OR3 (N877, N870, N647, N531);
or OR3 (N878, N848, N750, N232);
nand NAND4 (N879, N867, N125, N722, N210);
and AND4 (N880, N872, N615, N715, N386);
and AND2 (N881, N877, N811);
and AND2 (N882, N874, N869);
not NOT1 (N883, N582);
nor NOR4 (N884, N876, N584, N529, N240);
nor NOR2 (N885, N884, N398);
xor XOR2 (N886, N882, N669);
or OR2 (N887, N885, N581);
nand NAND2 (N888, N879, N851);
nor NOR4 (N889, N883, N259, N201, N426);
xor XOR2 (N890, N878, N286);
nor NOR2 (N891, N887, N95);
nor NOR3 (N892, N886, N42, N795);
nor NOR2 (N893, N881, N69);
and AND3 (N894, N890, N433, N817);
nand NAND3 (N895, N892, N156, N892);
nor NOR4 (N896, N893, N495, N778, N645);
and AND2 (N897, N889, N888);
buf BUF1 (N898, N365);
nor NOR2 (N899, N891, N309);
nor NOR3 (N900, N871, N222, N141);
nand NAND2 (N901, N856, N900);
nor NOR3 (N902, N174, N809, N769);
and AND2 (N903, N902, N791);
nor NOR4 (N904, N903, N814, N374, N200);
and AND2 (N905, N880, N463);
nand NAND4 (N906, N904, N480, N256, N656);
xor XOR2 (N907, N905, N597);
and AND4 (N908, N895, N799, N309, N566);
and AND3 (N909, N899, N642, N595);
or OR4 (N910, N907, N370, N75, N242);
not NOT1 (N911, N908);
nor NOR2 (N912, N901, N217);
nor NOR4 (N913, N906, N533, N144, N608);
xor XOR2 (N914, N894, N597);
nand NAND4 (N915, N910, N126, N464, N737);
nand NAND2 (N916, N915, N570);
nor NOR4 (N917, N896, N80, N579, N732);
buf BUF1 (N918, N914);
and AND3 (N919, N916, N550, N541);
not NOT1 (N920, N918);
xor XOR2 (N921, N909, N252);
or OR2 (N922, N920, N620);
xor XOR2 (N923, N922, N854);
and AND4 (N924, N911, N584, N385, N818);
xor XOR2 (N925, N917, N734);
nor NOR4 (N926, N897, N734, N853, N435);
xor XOR2 (N927, N913, N126);
buf BUF1 (N928, N926);
buf BUF1 (N929, N923);
xor XOR2 (N930, N929, N808);
and AND4 (N931, N927, N567, N587, N322);
nor NOR2 (N932, N925, N692);
or OR2 (N933, N921, N274);
nor NOR3 (N934, N930, N346, N772);
buf BUF1 (N935, N933);
and AND2 (N936, N912, N277);
or OR2 (N937, N931, N689);
and AND2 (N938, N932, N583);
not NOT1 (N939, N919);
xor XOR2 (N940, N924, N532);
xor XOR2 (N941, N936, N267);
or OR3 (N942, N939, N33, N781);
xor XOR2 (N943, N898, N568);
xor XOR2 (N944, N943, N225);
xor XOR2 (N945, N938, N801);
xor XOR2 (N946, N937, N725);
and AND4 (N947, N934, N667, N585, N14);
or OR3 (N948, N942, N87, N594);
or OR3 (N949, N946, N571, N385);
nand NAND2 (N950, N928, N924);
nand NAND4 (N951, N944, N133, N889, N695);
nor NOR2 (N952, N873, N471);
buf BUF1 (N953, N951);
nand NAND2 (N954, N940, N921);
nand NAND4 (N955, N949, N670, N593, N656);
xor XOR2 (N956, N950, N813);
buf BUF1 (N957, N945);
xor XOR2 (N958, N954, N631);
buf BUF1 (N959, N956);
not NOT1 (N960, N955);
not NOT1 (N961, N948);
nor NOR4 (N962, N941, N281, N215, N608);
xor XOR2 (N963, N952, N70);
buf BUF1 (N964, N962);
buf BUF1 (N965, N961);
nor NOR4 (N966, N965, N527, N94, N618);
nand NAND4 (N967, N935, N327, N286, N45);
nor NOR4 (N968, N959, N568, N361, N585);
xor XOR2 (N969, N967, N665);
or OR4 (N970, N963, N622, N247, N176);
not NOT1 (N971, N958);
or OR4 (N972, N957, N935, N184, N737);
nor NOR4 (N973, N966, N790, N297, N8);
buf BUF1 (N974, N953);
not NOT1 (N975, N974);
nor NOR4 (N976, N971, N399, N495, N388);
not NOT1 (N977, N976);
not NOT1 (N978, N973);
xor XOR2 (N979, N964, N681);
xor XOR2 (N980, N947, N721);
buf BUF1 (N981, N960);
nand NAND4 (N982, N978, N1, N451, N34);
not NOT1 (N983, N977);
buf BUF1 (N984, N981);
and AND2 (N985, N972, N956);
xor XOR2 (N986, N970, N188);
or OR2 (N987, N968, N609);
or OR4 (N988, N975, N310, N819, N169);
buf BUF1 (N989, N982);
nand NAND3 (N990, N985, N11, N114);
xor XOR2 (N991, N989, N484);
and AND4 (N992, N988, N804, N321, N90);
xor XOR2 (N993, N979, N219);
not NOT1 (N994, N984);
nand NAND3 (N995, N980, N39, N400);
and AND2 (N996, N990, N503);
and AND3 (N997, N994, N721, N62);
nor NOR4 (N998, N997, N707, N151, N44);
xor XOR2 (N999, N996, N352);
xor XOR2 (N1000, N987, N936);
not NOT1 (N1001, N1000);
buf BUF1 (N1002, N983);
buf BUF1 (N1003, N986);
xor XOR2 (N1004, N999, N370);
xor XOR2 (N1005, N995, N795);
not NOT1 (N1006, N998);
xor XOR2 (N1007, N1006, N984);
nand NAND4 (N1008, N993, N895, N430, N773);
nor NOR4 (N1009, N1003, N552, N292, N155);
nor NOR2 (N1010, N969, N146);
and AND4 (N1011, N992, N2, N18, N211);
or OR3 (N1012, N1001, N56, N148);
not NOT1 (N1013, N991);
not NOT1 (N1014, N1002);
nand NAND4 (N1015, N1010, N84, N825, N377);
buf BUF1 (N1016, N1011);
or OR4 (N1017, N1013, N716, N336, N147);
nand NAND3 (N1018, N1015, N428, N624);
or OR4 (N1019, N1012, N411, N159, N999);
or OR3 (N1020, N1014, N372, N526);
nand NAND2 (N1021, N1017, N543);
not NOT1 (N1022, N1007);
or OR3 (N1023, N1004, N663, N729);
xor XOR2 (N1024, N1005, N52);
nand NAND3 (N1025, N1022, N914, N164);
buf BUF1 (N1026, N1025);
not NOT1 (N1027, N1019);
nor NOR2 (N1028, N1024, N59);
and AND4 (N1029, N1016, N187, N726, N254);
and AND3 (N1030, N1009, N715, N524);
nor NOR2 (N1031, N1021, N974);
xor XOR2 (N1032, N1018, N360);
xor XOR2 (N1033, N1029, N452);
not NOT1 (N1034, N1028);
not NOT1 (N1035, N1033);
nand NAND3 (N1036, N1027, N57, N96);
and AND2 (N1037, N1031, N794);
xor XOR2 (N1038, N1037, N219);
nand NAND2 (N1039, N1036, N800);
buf BUF1 (N1040, N1032);
nand NAND3 (N1041, N1040, N166, N102);
nor NOR2 (N1042, N1034, N711);
or OR3 (N1043, N1038, N522, N350);
nor NOR4 (N1044, N1023, N102, N857, N543);
nand NAND3 (N1045, N1042, N124, N498);
nor NOR2 (N1046, N1039, N705);
buf BUF1 (N1047, N1030);
xor XOR2 (N1048, N1041, N155);
buf BUF1 (N1049, N1044);
or OR2 (N1050, N1008, N11);
nand NAND3 (N1051, N1020, N683, N928);
or OR3 (N1052, N1049, N167, N737);
nand NAND2 (N1053, N1047, N631);
nand NAND2 (N1054, N1048, N161);
nand NAND3 (N1055, N1053, N239, N81);
buf BUF1 (N1056, N1054);
nor NOR4 (N1057, N1055, N781, N631, N921);
and AND4 (N1058, N1043, N816, N83, N604);
buf BUF1 (N1059, N1026);
not NOT1 (N1060, N1051);
and AND2 (N1061, N1045, N734);
and AND4 (N1062, N1056, N313, N156, N1018);
not NOT1 (N1063, N1035);
not NOT1 (N1064, N1061);
and AND3 (N1065, N1060, N193, N119);
buf BUF1 (N1066, N1065);
or OR4 (N1067, N1064, N440, N943, N868);
and AND3 (N1068, N1057, N454, N656);
xor XOR2 (N1069, N1046, N152);
buf BUF1 (N1070, N1063);
or OR3 (N1071, N1066, N885, N212);
and AND4 (N1072, N1071, N818, N1022, N89);
nand NAND3 (N1073, N1069, N726, N549);
and AND4 (N1074, N1073, N774, N382, N268);
nor NOR2 (N1075, N1062, N576);
xor XOR2 (N1076, N1075, N955);
or OR2 (N1077, N1059, N998);
nor NOR2 (N1078, N1074, N712);
buf BUF1 (N1079, N1052);
or OR2 (N1080, N1070, N593);
not NOT1 (N1081, N1078);
or OR4 (N1082, N1081, N702, N370, N952);
or OR2 (N1083, N1050, N39);
not NOT1 (N1084, N1077);
buf BUF1 (N1085, N1080);
and AND2 (N1086, N1082, N620);
and AND4 (N1087, N1086, N450, N1016, N467);
xor XOR2 (N1088, N1087, N883);
buf BUF1 (N1089, N1083);
and AND4 (N1090, N1079, N870, N752, N522);
nand NAND4 (N1091, N1068, N105, N889, N654);
not NOT1 (N1092, N1076);
or OR4 (N1093, N1067, N482, N561, N654);
and AND2 (N1094, N1058, N11);
buf BUF1 (N1095, N1072);
nand NAND3 (N1096, N1089, N1079, N245);
or OR2 (N1097, N1094, N552);
buf BUF1 (N1098, N1084);
or OR3 (N1099, N1088, N70, N913);
and AND2 (N1100, N1093, N337);
buf BUF1 (N1101, N1098);
buf BUF1 (N1102, N1090);
xor XOR2 (N1103, N1095, N127);
and AND2 (N1104, N1092, N201);
xor XOR2 (N1105, N1102, N104);
buf BUF1 (N1106, N1101);
nand NAND4 (N1107, N1104, N839, N265, N537);
and AND2 (N1108, N1106, N679);
not NOT1 (N1109, N1103);
xor XOR2 (N1110, N1105, N540);
nand NAND4 (N1111, N1091, N583, N4, N809);
and AND4 (N1112, N1096, N383, N386, N786);
xor XOR2 (N1113, N1112, N395);
xor XOR2 (N1114, N1110, N756);
xor XOR2 (N1115, N1100, N24);
or OR2 (N1116, N1114, N694);
or OR4 (N1117, N1099, N619, N669, N154);
not NOT1 (N1118, N1115);
not NOT1 (N1119, N1111);
nor NOR3 (N1120, N1117, N1009, N263);
buf BUF1 (N1121, N1120);
nor NOR4 (N1122, N1085, N573, N200, N866);
xor XOR2 (N1123, N1108, N642);
nand NAND2 (N1124, N1119, N988);
and AND4 (N1125, N1123, N799, N97, N388);
not NOT1 (N1126, N1116);
buf BUF1 (N1127, N1107);
not NOT1 (N1128, N1118);
nand NAND3 (N1129, N1097, N658, N712);
or OR2 (N1130, N1113, N43);
buf BUF1 (N1131, N1109);
buf BUF1 (N1132, N1127);
not NOT1 (N1133, N1128);
buf BUF1 (N1134, N1132);
nand NAND2 (N1135, N1130, N1084);
nor NOR4 (N1136, N1134, N1125, N1122, N803);
and AND2 (N1137, N23, N725);
buf BUF1 (N1138, N1113);
buf BUF1 (N1139, N1126);
nand NAND3 (N1140, N1136, N404, N375);
xor XOR2 (N1141, N1124, N114);
or OR2 (N1142, N1137, N1020);
and AND2 (N1143, N1138, N186);
xor XOR2 (N1144, N1129, N519);
buf BUF1 (N1145, N1131);
or OR2 (N1146, N1144, N284);
not NOT1 (N1147, N1145);
or OR4 (N1148, N1133, N670, N552, N633);
buf BUF1 (N1149, N1139);
xor XOR2 (N1150, N1147, N816);
and AND4 (N1151, N1148, N1111, N1069, N544);
nand NAND4 (N1152, N1146, N47, N815, N371);
or OR2 (N1153, N1152, N957);
nand NAND3 (N1154, N1151, N931, N839);
nand NAND2 (N1155, N1143, N297);
and AND4 (N1156, N1135, N1069, N458, N1081);
nor NOR2 (N1157, N1156, N690);
not NOT1 (N1158, N1154);
nor NOR3 (N1159, N1150, N645, N1101);
not NOT1 (N1160, N1159);
and AND3 (N1161, N1121, N846, N176);
not NOT1 (N1162, N1160);
not NOT1 (N1163, N1162);
not NOT1 (N1164, N1141);
or OR2 (N1165, N1157, N525);
xor XOR2 (N1166, N1149, N1145);
buf BUF1 (N1167, N1164);
nand NAND4 (N1168, N1140, N679, N1092, N883);
nand NAND3 (N1169, N1163, N1138, N1066);
not NOT1 (N1170, N1161);
not NOT1 (N1171, N1153);
not NOT1 (N1172, N1171);
nand NAND3 (N1173, N1155, N795, N206);
xor XOR2 (N1174, N1142, N880);
nor NOR4 (N1175, N1170, N322, N901, N292);
nor NOR3 (N1176, N1168, N977, N1045);
nor NOR3 (N1177, N1176, N642, N808);
not NOT1 (N1178, N1166);
buf BUF1 (N1179, N1158);
or OR2 (N1180, N1179, N16);
nand NAND4 (N1181, N1173, N215, N392, N371);
or OR3 (N1182, N1169, N316, N489);
not NOT1 (N1183, N1177);
not NOT1 (N1184, N1181);
nand NAND4 (N1185, N1178, N911, N228, N557);
nor NOR3 (N1186, N1167, N977, N415);
and AND4 (N1187, N1186, N890, N990, N319);
xor XOR2 (N1188, N1182, N28);
or OR4 (N1189, N1185, N1086, N939, N19);
xor XOR2 (N1190, N1175, N704);
not NOT1 (N1191, N1190);
nor NOR3 (N1192, N1174, N427, N38);
nor NOR3 (N1193, N1187, N655, N150);
not NOT1 (N1194, N1192);
not NOT1 (N1195, N1172);
and AND4 (N1196, N1180, N3, N208, N595);
or OR3 (N1197, N1165, N260, N230);
not NOT1 (N1198, N1194);
and AND2 (N1199, N1197, N258);
nand NAND3 (N1200, N1183, N54, N607);
or OR3 (N1201, N1199, N489, N462);
not NOT1 (N1202, N1189);
or OR3 (N1203, N1202, N712, N924);
nor NOR2 (N1204, N1203, N201);
not NOT1 (N1205, N1184);
nand NAND4 (N1206, N1205, N568, N850, N874);
nand NAND2 (N1207, N1188, N137);
and AND3 (N1208, N1204, N179, N841);
xor XOR2 (N1209, N1201, N459);
nor NOR4 (N1210, N1191, N426, N952, N997);
not NOT1 (N1211, N1195);
nand NAND2 (N1212, N1200, N1059);
or OR4 (N1213, N1209, N676, N1127, N12);
or OR2 (N1214, N1206, N1031);
buf BUF1 (N1215, N1212);
nor NOR4 (N1216, N1215, N706, N681, N194);
nand NAND3 (N1217, N1211, N121, N557);
and AND4 (N1218, N1214, N668, N421, N371);
or OR4 (N1219, N1193, N539, N969, N192);
buf BUF1 (N1220, N1216);
and AND2 (N1221, N1219, N1095);
xor XOR2 (N1222, N1220, N10);
nor NOR4 (N1223, N1217, N768, N328, N122);
nand NAND2 (N1224, N1218, N1128);
or OR3 (N1225, N1222, N19, N464);
buf BUF1 (N1226, N1224);
not NOT1 (N1227, N1221);
or OR4 (N1228, N1210, N259, N1124, N160);
nor NOR4 (N1229, N1226, N223, N537, N1087);
or OR2 (N1230, N1227, N1205);
buf BUF1 (N1231, N1198);
xor XOR2 (N1232, N1225, N1181);
or OR3 (N1233, N1231, N1187, N253);
or OR4 (N1234, N1232, N177, N767, N348);
or OR3 (N1235, N1208, N57, N263);
buf BUF1 (N1236, N1213);
xor XOR2 (N1237, N1230, N1212);
xor XOR2 (N1238, N1234, N1016);
buf BUF1 (N1239, N1196);
not NOT1 (N1240, N1237);
buf BUF1 (N1241, N1228);
and AND3 (N1242, N1223, N40, N227);
xor XOR2 (N1243, N1241, N414);
buf BUF1 (N1244, N1240);
nand NAND4 (N1245, N1233, N394, N853, N266);
and AND3 (N1246, N1245, N991, N983);
nand NAND3 (N1247, N1246, N1045, N648);
not NOT1 (N1248, N1229);
buf BUF1 (N1249, N1243);
xor XOR2 (N1250, N1207, N320);
and AND3 (N1251, N1248, N1126, N521);
xor XOR2 (N1252, N1238, N706);
not NOT1 (N1253, N1251);
not NOT1 (N1254, N1247);
not NOT1 (N1255, N1254);
and AND2 (N1256, N1244, N401);
and AND2 (N1257, N1236, N367);
not NOT1 (N1258, N1256);
not NOT1 (N1259, N1242);
not NOT1 (N1260, N1249);
nor NOR3 (N1261, N1235, N1052, N1068);
nor NOR2 (N1262, N1258, N357);
buf BUF1 (N1263, N1250);
nand NAND2 (N1264, N1239, N403);
nor NOR2 (N1265, N1264, N691);
xor XOR2 (N1266, N1252, N1053);
not NOT1 (N1267, N1263);
not NOT1 (N1268, N1253);
xor XOR2 (N1269, N1257, N385);
nor NOR2 (N1270, N1265, N546);
nand NAND2 (N1271, N1259, N716);
buf BUF1 (N1272, N1266);
buf BUF1 (N1273, N1261);
and AND2 (N1274, N1270, N1175);
xor XOR2 (N1275, N1271, N1208);
and AND3 (N1276, N1273, N1138, N735);
xor XOR2 (N1277, N1274, N313);
nor NOR3 (N1278, N1269, N23, N1098);
or OR2 (N1279, N1276, N363);
buf BUF1 (N1280, N1267);
nor NOR4 (N1281, N1268, N445, N1252, N1257);
and AND4 (N1282, N1281, N882, N176, N222);
or OR2 (N1283, N1278, N345);
xor XOR2 (N1284, N1255, N1245);
xor XOR2 (N1285, N1280, N99);
and AND2 (N1286, N1272, N597);
nand NAND4 (N1287, N1260, N279, N759, N361);
and AND3 (N1288, N1286, N501, N482);
nor NOR2 (N1289, N1284, N365);
not NOT1 (N1290, N1279);
or OR4 (N1291, N1283, N240, N1256, N751);
nand NAND3 (N1292, N1290, N497, N317);
nand NAND2 (N1293, N1282, N386);
xor XOR2 (N1294, N1292, N302);
xor XOR2 (N1295, N1275, N666);
nor NOR2 (N1296, N1289, N1183);
nor NOR2 (N1297, N1277, N154);
or OR3 (N1298, N1285, N1005, N748);
xor XOR2 (N1299, N1294, N466);
and AND4 (N1300, N1288, N801, N289, N989);
nor NOR4 (N1301, N1295, N1262, N42, N1210);
and AND3 (N1302, N305, N797, N859);
buf BUF1 (N1303, N1291);
not NOT1 (N1304, N1298);
not NOT1 (N1305, N1304);
not NOT1 (N1306, N1301);
nor NOR4 (N1307, N1302, N623, N1111, N31);
buf BUF1 (N1308, N1305);
nand NAND4 (N1309, N1287, N685, N273, N307);
and AND3 (N1310, N1297, N808, N1305);
buf BUF1 (N1311, N1307);
and AND3 (N1312, N1293, N1222, N293);
and AND4 (N1313, N1312, N1065, N657, N851);
xor XOR2 (N1314, N1311, N973);
buf BUF1 (N1315, N1300);
xor XOR2 (N1316, N1313, N233);
nand NAND2 (N1317, N1303, N995);
buf BUF1 (N1318, N1299);
xor XOR2 (N1319, N1315, N1091);
buf BUF1 (N1320, N1314);
not NOT1 (N1321, N1309);
nand NAND3 (N1322, N1319, N704, N917);
and AND2 (N1323, N1317, N63);
buf BUF1 (N1324, N1321);
buf BUF1 (N1325, N1318);
and AND4 (N1326, N1322, N500, N1269, N675);
and AND2 (N1327, N1306, N634);
nor NOR2 (N1328, N1327, N1148);
buf BUF1 (N1329, N1296);
nand NAND4 (N1330, N1323, N260, N812, N503);
or OR2 (N1331, N1320, N542);
or OR2 (N1332, N1328, N1131);
buf BUF1 (N1333, N1316);
and AND3 (N1334, N1308, N517, N1070);
or OR2 (N1335, N1324, N998);
not NOT1 (N1336, N1330);
nand NAND3 (N1337, N1329, N256, N429);
nor NOR2 (N1338, N1335, N1296);
nor NOR4 (N1339, N1332, N660, N1215, N680);
nor NOR2 (N1340, N1338, N1064);
xor XOR2 (N1341, N1339, N422);
nand NAND2 (N1342, N1334, N793);
nor NOR2 (N1343, N1310, N493);
buf BUF1 (N1344, N1331);
nand NAND4 (N1345, N1326, N924, N882, N893);
not NOT1 (N1346, N1340);
nand NAND4 (N1347, N1344, N1110, N112, N974);
nor NOR2 (N1348, N1343, N404);
or OR2 (N1349, N1333, N1063);
xor XOR2 (N1350, N1325, N118);
xor XOR2 (N1351, N1349, N896);
or OR3 (N1352, N1347, N292, N781);
or OR3 (N1353, N1351, N158, N330);
not NOT1 (N1354, N1337);
and AND4 (N1355, N1342, N840, N1088, N147);
or OR3 (N1356, N1346, N1161, N937);
xor XOR2 (N1357, N1354, N944);
xor XOR2 (N1358, N1345, N260);
nand NAND4 (N1359, N1356, N1023, N695, N123);
xor XOR2 (N1360, N1350, N136);
not NOT1 (N1361, N1348);
xor XOR2 (N1362, N1336, N240);
or OR2 (N1363, N1361, N699);
not NOT1 (N1364, N1360);
nor NOR2 (N1365, N1363, N1214);
buf BUF1 (N1366, N1357);
buf BUF1 (N1367, N1366);
nor NOR2 (N1368, N1352, N128);
xor XOR2 (N1369, N1359, N1168);
nand NAND2 (N1370, N1367, N172);
and AND2 (N1371, N1370, N827);
xor XOR2 (N1372, N1358, N114);
not NOT1 (N1373, N1364);
buf BUF1 (N1374, N1368);
and AND4 (N1375, N1372, N461, N187, N419);
or OR4 (N1376, N1362, N696, N1205, N337);
and AND4 (N1377, N1341, N1139, N311, N750);
and AND3 (N1378, N1355, N20, N1277);
or OR3 (N1379, N1365, N677, N1235);
and AND2 (N1380, N1374, N237);
xor XOR2 (N1381, N1375, N26);
buf BUF1 (N1382, N1380);
and AND2 (N1383, N1379, N84);
buf BUF1 (N1384, N1381);
or OR2 (N1385, N1383, N625);
xor XOR2 (N1386, N1384, N872);
xor XOR2 (N1387, N1386, N722);
xor XOR2 (N1388, N1369, N549);
xor XOR2 (N1389, N1378, N682);
and AND4 (N1390, N1388, N859, N926, N115);
and AND3 (N1391, N1377, N139, N588);
not NOT1 (N1392, N1373);
and AND4 (N1393, N1387, N1184, N72, N768);
xor XOR2 (N1394, N1392, N1266);
or OR4 (N1395, N1382, N746, N85, N678);
and AND4 (N1396, N1389, N751, N229, N56);
nor NOR2 (N1397, N1395, N1074);
not NOT1 (N1398, N1390);
and AND2 (N1399, N1394, N830);
or OR3 (N1400, N1385, N18, N1387);
buf BUF1 (N1401, N1398);
xor XOR2 (N1402, N1376, N292);
buf BUF1 (N1403, N1402);
or OR3 (N1404, N1401, N340, N245);
not NOT1 (N1405, N1400);
xor XOR2 (N1406, N1396, N1033);
nand NAND4 (N1407, N1353, N314, N803, N777);
or OR4 (N1408, N1397, N957, N1163, N943);
nand NAND2 (N1409, N1407, N597);
or OR2 (N1410, N1406, N41);
or OR3 (N1411, N1371, N726, N519);
not NOT1 (N1412, N1393);
nor NOR2 (N1413, N1391, N721);
not NOT1 (N1414, N1410);
and AND4 (N1415, N1408, N939, N1007, N847);
and AND3 (N1416, N1412, N646, N1403);
or OR3 (N1417, N250, N476, N667);
not NOT1 (N1418, N1405);
xor XOR2 (N1419, N1418, N747);
not NOT1 (N1420, N1417);
nand NAND3 (N1421, N1409, N823, N1029);
not NOT1 (N1422, N1414);
and AND3 (N1423, N1399, N975, N10);
nor NOR4 (N1424, N1421, N758, N808, N57);
not NOT1 (N1425, N1424);
nand NAND2 (N1426, N1415, N395);
not NOT1 (N1427, N1411);
xor XOR2 (N1428, N1420, N852);
nor NOR4 (N1429, N1413, N409, N209, N522);
and AND4 (N1430, N1416, N766, N846, N1063);
nor NOR4 (N1431, N1426, N708, N29, N575);
and AND4 (N1432, N1428, N709, N99, N272);
and AND3 (N1433, N1422, N1288, N316);
or OR4 (N1434, N1404, N753, N848, N115);
or OR2 (N1435, N1423, N233);
nand NAND2 (N1436, N1427, N821);
xor XOR2 (N1437, N1434, N8);
and AND4 (N1438, N1433, N800, N565, N227);
not NOT1 (N1439, N1437);
and AND2 (N1440, N1436, N301);
nand NAND2 (N1441, N1438, N176);
nor NOR4 (N1442, N1431, N724, N197, N1192);
or OR2 (N1443, N1442, N1317);
not NOT1 (N1444, N1439);
xor XOR2 (N1445, N1443, N1181);
or OR2 (N1446, N1440, N387);
nand NAND3 (N1447, N1444, N1062, N1383);
and AND2 (N1448, N1441, N788);
and AND3 (N1449, N1419, N1012, N248);
and AND2 (N1450, N1448, N236);
xor XOR2 (N1451, N1447, N1198);
and AND2 (N1452, N1451, N712);
and AND3 (N1453, N1452, N557, N873);
nor NOR2 (N1454, N1429, N708);
and AND4 (N1455, N1425, N606, N1334, N346);
nor NOR3 (N1456, N1449, N172, N1361);
nor NOR3 (N1457, N1456, N277, N1262);
or OR3 (N1458, N1435, N535, N955);
nor NOR2 (N1459, N1445, N839);
nand NAND4 (N1460, N1453, N332, N306, N648);
xor XOR2 (N1461, N1458, N292);
and AND3 (N1462, N1455, N611, N878);
xor XOR2 (N1463, N1454, N621);
xor XOR2 (N1464, N1461, N969);
and AND2 (N1465, N1430, N1074);
or OR3 (N1466, N1462, N953, N230);
and AND4 (N1467, N1450, N795, N2, N1034);
xor XOR2 (N1468, N1459, N1189);
xor XOR2 (N1469, N1467, N146);
or OR3 (N1470, N1465, N871, N1287);
nand NAND3 (N1471, N1432, N1283, N921);
nor NOR2 (N1472, N1466, N536);
and AND3 (N1473, N1469, N659, N438);
buf BUF1 (N1474, N1464);
nand NAND3 (N1475, N1473, N1350, N145);
and AND3 (N1476, N1471, N776, N686);
buf BUF1 (N1477, N1476);
buf BUF1 (N1478, N1474);
and AND4 (N1479, N1478, N69, N232, N1336);
nand NAND2 (N1480, N1479, N951);
buf BUF1 (N1481, N1472);
nand NAND3 (N1482, N1477, N702, N602);
nor NOR3 (N1483, N1446, N894, N569);
and AND2 (N1484, N1460, N621);
and AND4 (N1485, N1470, N715, N985, N1422);
nand NAND2 (N1486, N1481, N802);
buf BUF1 (N1487, N1485);
buf BUF1 (N1488, N1484);
not NOT1 (N1489, N1482);
or OR4 (N1490, N1487, N416, N1462, N961);
xor XOR2 (N1491, N1488, N313);
buf BUF1 (N1492, N1463);
nor NOR4 (N1493, N1468, N370, N33, N768);
or OR4 (N1494, N1486, N426, N86, N810);
or OR4 (N1495, N1483, N409, N44, N785);
buf BUF1 (N1496, N1495);
xor XOR2 (N1497, N1496, N446);
or OR2 (N1498, N1493, N24);
buf BUF1 (N1499, N1491);
xor XOR2 (N1500, N1498, N643);
buf BUF1 (N1501, N1475);
buf BUF1 (N1502, N1497);
buf BUF1 (N1503, N1489);
nor NOR2 (N1504, N1499, N370);
xor XOR2 (N1505, N1494, N422);
or OR3 (N1506, N1505, N82, N1368);
and AND4 (N1507, N1490, N1262, N1345, N952);
buf BUF1 (N1508, N1504);
nor NOR2 (N1509, N1501, N903);
and AND2 (N1510, N1457, N537);
nor NOR2 (N1511, N1492, N638);
not NOT1 (N1512, N1500);
xor XOR2 (N1513, N1508, N1493);
or OR4 (N1514, N1502, N1144, N1007, N505);
buf BUF1 (N1515, N1510);
xor XOR2 (N1516, N1514, N912);
and AND4 (N1517, N1509, N1116, N145, N1138);
buf BUF1 (N1518, N1507);
or OR2 (N1519, N1518, N243);
nor NOR3 (N1520, N1503, N468, N1195);
xor XOR2 (N1521, N1520, N1485);
and AND3 (N1522, N1512, N920, N1055);
and AND3 (N1523, N1480, N867, N465);
not NOT1 (N1524, N1513);
not NOT1 (N1525, N1521);
nand NAND3 (N1526, N1523, N990, N445);
buf BUF1 (N1527, N1519);
and AND4 (N1528, N1511, N551, N1461, N1227);
nand NAND3 (N1529, N1526, N645, N380);
nand NAND2 (N1530, N1515, N841);
nand NAND4 (N1531, N1529, N132, N1529, N1494);
and AND3 (N1532, N1506, N884, N236);
nor NOR3 (N1533, N1530, N737, N764);
xor XOR2 (N1534, N1522, N1115);
xor XOR2 (N1535, N1524, N719);
xor XOR2 (N1536, N1516, N1432);
nor NOR4 (N1537, N1535, N647, N1193, N1476);
buf BUF1 (N1538, N1531);
nor NOR4 (N1539, N1517, N607, N925, N828);
nor NOR2 (N1540, N1539, N823);
xor XOR2 (N1541, N1538, N551);
and AND2 (N1542, N1525, N8);
nand NAND4 (N1543, N1537, N769, N580, N446);
not NOT1 (N1544, N1542);
xor XOR2 (N1545, N1541, N221);
and AND4 (N1546, N1545, N837, N553, N15);
not NOT1 (N1547, N1533);
or OR2 (N1548, N1540, N876);
nor NOR2 (N1549, N1528, N169);
not NOT1 (N1550, N1532);
xor XOR2 (N1551, N1536, N909);
buf BUF1 (N1552, N1534);
nand NAND3 (N1553, N1527, N178, N1294);
nand NAND3 (N1554, N1551, N960, N1003);
and AND2 (N1555, N1547, N719);
xor XOR2 (N1556, N1552, N513);
buf BUF1 (N1557, N1553);
nand NAND2 (N1558, N1548, N794);
and AND4 (N1559, N1543, N710, N1067, N932);
xor XOR2 (N1560, N1558, N1498);
or OR2 (N1561, N1560, N384);
or OR3 (N1562, N1557, N1303, N973);
not NOT1 (N1563, N1556);
buf BUF1 (N1564, N1549);
nor NOR2 (N1565, N1550, N942);
buf BUF1 (N1566, N1561);
not NOT1 (N1567, N1562);
or OR2 (N1568, N1559, N458);
xor XOR2 (N1569, N1565, N217);
and AND2 (N1570, N1563, N721);
nand NAND3 (N1571, N1568, N575, N542);
not NOT1 (N1572, N1569);
not NOT1 (N1573, N1572);
buf BUF1 (N1574, N1555);
xor XOR2 (N1575, N1574, N1359);
or OR3 (N1576, N1566, N913, N1427);
or OR4 (N1577, N1546, N1414, N364, N1368);
nand NAND3 (N1578, N1576, N1566, N1127);
nor NOR3 (N1579, N1573, N355, N1134);
buf BUF1 (N1580, N1567);
not NOT1 (N1581, N1564);
nor NOR2 (N1582, N1577, N339);
and AND3 (N1583, N1578, N1021, N1050);
nor NOR3 (N1584, N1579, N1501, N82);
xor XOR2 (N1585, N1582, N628);
nand NAND2 (N1586, N1570, N1489);
nand NAND4 (N1587, N1581, N1299, N1542, N639);
nand NAND2 (N1588, N1585, N1394);
or OR3 (N1589, N1544, N875, N93);
and AND4 (N1590, N1571, N336, N407, N96);
xor XOR2 (N1591, N1590, N249);
nand NAND4 (N1592, N1580, N373, N539, N1522);
and AND4 (N1593, N1584, N1093, N714, N1177);
and AND2 (N1594, N1589, N1252);
xor XOR2 (N1595, N1594, N337);
nor NOR2 (N1596, N1575, N310);
or OR3 (N1597, N1554, N675, N309);
nor NOR2 (N1598, N1596, N1010);
not NOT1 (N1599, N1593);
nand NAND3 (N1600, N1588, N61, N209);
or OR2 (N1601, N1597, N1101);
xor XOR2 (N1602, N1591, N309);
and AND2 (N1603, N1595, N197);
not NOT1 (N1604, N1603);
nand NAND2 (N1605, N1583, N827);
and AND4 (N1606, N1586, N671, N775, N840);
nand NAND3 (N1607, N1605, N394, N868);
buf BUF1 (N1608, N1600);
and AND2 (N1609, N1598, N318);
and AND4 (N1610, N1609, N228, N1562, N328);
nor NOR3 (N1611, N1602, N906, N1165);
nor NOR4 (N1612, N1610, N1096, N239, N157);
nor NOR3 (N1613, N1592, N867, N533);
and AND4 (N1614, N1606, N1335, N1422, N1215);
and AND4 (N1615, N1612, N1432, N216, N652);
buf BUF1 (N1616, N1601);
not NOT1 (N1617, N1616);
not NOT1 (N1618, N1617);
nand NAND4 (N1619, N1614, N489, N1188, N728);
nor NOR2 (N1620, N1599, N265);
nand NAND4 (N1621, N1620, N1284, N871, N1372);
not NOT1 (N1622, N1608);
not NOT1 (N1623, N1622);
xor XOR2 (N1624, N1587, N795);
nand NAND2 (N1625, N1604, N1565);
nor NOR3 (N1626, N1613, N1404, N883);
nor NOR4 (N1627, N1619, N1575, N1594, N710);
and AND4 (N1628, N1625, N953, N980, N735);
buf BUF1 (N1629, N1611);
nand NAND4 (N1630, N1629, N1210, N1250, N533);
nand NAND2 (N1631, N1626, N336);
nor NOR4 (N1632, N1624, N1393, N1189, N1532);
or OR2 (N1633, N1630, N264);
and AND2 (N1634, N1618, N552);
and AND2 (N1635, N1627, N589);
buf BUF1 (N1636, N1631);
or OR3 (N1637, N1634, N263, N1486);
not NOT1 (N1638, N1623);
or OR4 (N1639, N1635, N29, N1607, N500);
buf BUF1 (N1640, N805);
not NOT1 (N1641, N1636);
or OR2 (N1642, N1621, N500);
and AND2 (N1643, N1641, N1292);
and AND3 (N1644, N1615, N1489, N12);
buf BUF1 (N1645, N1638);
nand NAND2 (N1646, N1639, N994);
nand NAND4 (N1647, N1628, N350, N1487, N1189);
nand NAND4 (N1648, N1637, N209, N632, N639);
or OR3 (N1649, N1647, N656, N586);
buf BUF1 (N1650, N1644);
nor NOR4 (N1651, N1633, N493, N1210, N1012);
xor XOR2 (N1652, N1645, N137);
xor XOR2 (N1653, N1646, N863);
nor NOR4 (N1654, N1642, N848, N107, N1095);
not NOT1 (N1655, N1632);
xor XOR2 (N1656, N1655, N122);
not NOT1 (N1657, N1654);
buf BUF1 (N1658, N1656);
or OR2 (N1659, N1651, N1638);
nand NAND3 (N1660, N1643, N217, N792);
or OR2 (N1661, N1658, N1199);
and AND4 (N1662, N1649, N1079, N1063, N962);
buf BUF1 (N1663, N1650);
nand NAND3 (N1664, N1661, N569, N1528);
nor NOR4 (N1665, N1663, N1135, N1639, N352);
xor XOR2 (N1666, N1660, N1265);
buf BUF1 (N1667, N1664);
or OR2 (N1668, N1652, N390);
nor NOR4 (N1669, N1657, N724, N137, N1236);
not NOT1 (N1670, N1648);
not NOT1 (N1671, N1668);
nand NAND4 (N1672, N1665, N1597, N22, N1619);
not NOT1 (N1673, N1672);
buf BUF1 (N1674, N1667);
buf BUF1 (N1675, N1674);
xor XOR2 (N1676, N1673, N33);
nand NAND3 (N1677, N1675, N1552, N675);
or OR4 (N1678, N1666, N1163, N1458, N1072);
and AND4 (N1679, N1659, N1072, N1420, N784);
or OR3 (N1680, N1669, N316, N776);
xor XOR2 (N1681, N1680, N1265);
xor XOR2 (N1682, N1671, N901);
and AND4 (N1683, N1681, N1146, N1367, N1167);
or OR3 (N1684, N1640, N946, N1597);
and AND3 (N1685, N1678, N977, N1224);
nor NOR2 (N1686, N1676, N1281);
or OR2 (N1687, N1679, N888);
not NOT1 (N1688, N1677);
not NOT1 (N1689, N1682);
nand NAND2 (N1690, N1653, N1505);
nand NAND2 (N1691, N1683, N1685);
or OR2 (N1692, N833, N1645);
nor NOR4 (N1693, N1662, N1289, N990, N1);
and AND3 (N1694, N1687, N326, N697);
or OR3 (N1695, N1686, N952, N1685);
buf BUF1 (N1696, N1695);
xor XOR2 (N1697, N1684, N1342);
not NOT1 (N1698, N1696);
buf BUF1 (N1699, N1697);
xor XOR2 (N1700, N1690, N1173);
xor XOR2 (N1701, N1694, N1251);
nand NAND4 (N1702, N1692, N74, N1640, N729);
xor XOR2 (N1703, N1689, N1422);
not NOT1 (N1704, N1670);
buf BUF1 (N1705, N1704);
and AND4 (N1706, N1688, N1525, N636, N1620);
or OR2 (N1707, N1699, N260);
not NOT1 (N1708, N1701);
buf BUF1 (N1709, N1703);
nor NOR2 (N1710, N1698, N1478);
nor NOR2 (N1711, N1691, N176);
and AND2 (N1712, N1706, N765);
nand NAND2 (N1713, N1711, N1311);
xor XOR2 (N1714, N1700, N437);
nand NAND2 (N1715, N1710, N1620);
or OR2 (N1716, N1715, N952);
or OR2 (N1717, N1716, N982);
nand NAND4 (N1718, N1702, N72, N1222, N1042);
or OR3 (N1719, N1709, N516, N439);
buf BUF1 (N1720, N1714);
xor XOR2 (N1721, N1719, N100);
buf BUF1 (N1722, N1712);
buf BUF1 (N1723, N1705);
xor XOR2 (N1724, N1717, N111);
nand NAND3 (N1725, N1708, N357, N905);
xor XOR2 (N1726, N1693, N127);
or OR2 (N1727, N1713, N1415);
nor NOR4 (N1728, N1707, N104, N886, N1248);
and AND4 (N1729, N1722, N1399, N1030, N1129);
buf BUF1 (N1730, N1723);
buf BUF1 (N1731, N1727);
or OR3 (N1732, N1726, N622, N748);
nor NOR3 (N1733, N1728, N326, N222);
or OR2 (N1734, N1732, N784);
xor XOR2 (N1735, N1731, N625);
or OR4 (N1736, N1725, N655, N638, N539);
buf BUF1 (N1737, N1718);
nor NOR4 (N1738, N1737, N914, N619, N705);
nor NOR2 (N1739, N1736, N1448);
or OR4 (N1740, N1721, N413, N490, N1656);
nor NOR3 (N1741, N1720, N102, N53);
buf BUF1 (N1742, N1733);
buf BUF1 (N1743, N1738);
buf BUF1 (N1744, N1729);
and AND4 (N1745, N1735, N430, N767, N753);
nor NOR4 (N1746, N1739, N248, N819, N1420);
buf BUF1 (N1747, N1743);
buf BUF1 (N1748, N1744);
nand NAND2 (N1749, N1745, N1669);
not NOT1 (N1750, N1749);
or OR4 (N1751, N1730, N469, N329, N1582);
xor XOR2 (N1752, N1750, N211);
and AND2 (N1753, N1724, N1230);
nor NOR4 (N1754, N1752, N1075, N110, N1375);
nor NOR2 (N1755, N1753, N1087);
buf BUF1 (N1756, N1748);
and AND2 (N1757, N1754, N1350);
buf BUF1 (N1758, N1746);
not NOT1 (N1759, N1755);
or OR2 (N1760, N1758, N227);
xor XOR2 (N1761, N1760, N724);
or OR3 (N1762, N1747, N860, N1655);
xor XOR2 (N1763, N1759, N373);
nand NAND4 (N1764, N1734, N327, N372, N572);
or OR3 (N1765, N1763, N336, N1095);
and AND4 (N1766, N1757, N188, N863, N689);
and AND3 (N1767, N1764, N533, N23);
xor XOR2 (N1768, N1767, N531);
nor NOR2 (N1769, N1756, N1635);
and AND4 (N1770, N1762, N940, N636, N238);
not NOT1 (N1771, N1741);
buf BUF1 (N1772, N1768);
and AND3 (N1773, N1771, N1637, N298);
or OR2 (N1774, N1769, N454);
buf BUF1 (N1775, N1751);
and AND2 (N1776, N1761, N5);
not NOT1 (N1777, N1776);
xor XOR2 (N1778, N1775, N356);
and AND2 (N1779, N1742, N1585);
and AND4 (N1780, N1778, N1532, N46, N658);
xor XOR2 (N1781, N1780, N588);
nand NAND2 (N1782, N1766, N1671);
buf BUF1 (N1783, N1777);
and AND2 (N1784, N1781, N638);
buf BUF1 (N1785, N1770);
and AND4 (N1786, N1779, N956, N260, N1748);
xor XOR2 (N1787, N1783, N1752);
or OR4 (N1788, N1740, N1736, N749, N1766);
and AND2 (N1789, N1765, N1552);
or OR2 (N1790, N1784, N830);
buf BUF1 (N1791, N1774);
or OR2 (N1792, N1787, N205);
nand NAND3 (N1793, N1786, N1717, N1697);
not NOT1 (N1794, N1792);
and AND3 (N1795, N1789, N1637, N413);
nor NOR2 (N1796, N1793, N1763);
buf BUF1 (N1797, N1795);
not NOT1 (N1798, N1782);
buf BUF1 (N1799, N1772);
or OR2 (N1800, N1790, N787);
xor XOR2 (N1801, N1788, N903);
not NOT1 (N1802, N1799);
nor NOR4 (N1803, N1794, N922, N1526, N779);
buf BUF1 (N1804, N1785);
buf BUF1 (N1805, N1773);
buf BUF1 (N1806, N1791);
nand NAND3 (N1807, N1797, N1181, N248);
nor NOR2 (N1808, N1803, N1339);
nor NOR3 (N1809, N1801, N1631, N196);
xor XOR2 (N1810, N1809, N1396);
nor NOR2 (N1811, N1805, N874);
not NOT1 (N1812, N1804);
or OR2 (N1813, N1811, N1313);
nor NOR4 (N1814, N1800, N1784, N1369, N281);
xor XOR2 (N1815, N1806, N1650);
nand NAND2 (N1816, N1807, N672);
and AND2 (N1817, N1796, N1060);
xor XOR2 (N1818, N1814, N1193);
not NOT1 (N1819, N1812);
nor NOR2 (N1820, N1819, N28);
and AND3 (N1821, N1810, N450, N244);
buf BUF1 (N1822, N1808);
not NOT1 (N1823, N1813);
not NOT1 (N1824, N1802);
nand NAND2 (N1825, N1817, N482);
and AND3 (N1826, N1822, N1120, N367);
buf BUF1 (N1827, N1820);
xor XOR2 (N1828, N1816, N1232);
buf BUF1 (N1829, N1798);
and AND2 (N1830, N1824, N114);
buf BUF1 (N1831, N1821);
not NOT1 (N1832, N1831);
or OR3 (N1833, N1826, N330, N811);
buf BUF1 (N1834, N1815);
not NOT1 (N1835, N1823);
buf BUF1 (N1836, N1829);
or OR2 (N1837, N1825, N758);
nand NAND3 (N1838, N1828, N990, N326);
or OR3 (N1839, N1833, N915, N610);
buf BUF1 (N1840, N1836);
xor XOR2 (N1841, N1834, N1790);
xor XOR2 (N1842, N1841, N702);
buf BUF1 (N1843, N1837);
xor XOR2 (N1844, N1840, N223);
or OR4 (N1845, N1832, N1182, N362, N900);
xor XOR2 (N1846, N1843, N1402);
not NOT1 (N1847, N1844);
nor NOR4 (N1848, N1827, N934, N374, N57);
xor XOR2 (N1849, N1845, N57);
and AND3 (N1850, N1839, N1135, N855);
and AND4 (N1851, N1850, N1460, N1403, N375);
buf BUF1 (N1852, N1842);
nand NAND3 (N1853, N1846, N936, N382);
or OR2 (N1854, N1852, N900);
not NOT1 (N1855, N1847);
not NOT1 (N1856, N1848);
and AND3 (N1857, N1851, N185, N1784);
and AND3 (N1858, N1854, N966, N1318);
nor NOR2 (N1859, N1835, N1011);
and AND2 (N1860, N1830, N458);
not NOT1 (N1861, N1853);
xor XOR2 (N1862, N1861, N1405);
nand NAND3 (N1863, N1859, N131, N820);
or OR4 (N1864, N1855, N367, N1620, N939);
or OR4 (N1865, N1860, N501, N426, N496);
nand NAND3 (N1866, N1862, N1680, N287);
nand NAND4 (N1867, N1857, N110, N477, N249);
xor XOR2 (N1868, N1818, N876);
or OR3 (N1869, N1867, N4, N319);
xor XOR2 (N1870, N1849, N653);
or OR3 (N1871, N1870, N1084, N983);
buf BUF1 (N1872, N1858);
nand NAND3 (N1873, N1863, N330, N1319);
buf BUF1 (N1874, N1871);
or OR4 (N1875, N1868, N899, N1444, N691);
not NOT1 (N1876, N1856);
not NOT1 (N1877, N1865);
nor NOR3 (N1878, N1874, N1235, N986);
or OR3 (N1879, N1876, N1737, N1063);
xor XOR2 (N1880, N1866, N922);
nand NAND3 (N1881, N1873, N888, N150);
xor XOR2 (N1882, N1864, N353);
not NOT1 (N1883, N1869);
not NOT1 (N1884, N1883);
nand NAND3 (N1885, N1881, N873, N741);
nor NOR4 (N1886, N1872, N492, N58, N1528);
and AND3 (N1887, N1886, N520, N312);
xor XOR2 (N1888, N1882, N153);
xor XOR2 (N1889, N1878, N1548);
buf BUF1 (N1890, N1838);
nand NAND2 (N1891, N1884, N1626);
or OR4 (N1892, N1880, N655, N937, N181);
and AND3 (N1893, N1879, N1056, N1096);
xor XOR2 (N1894, N1892, N937);
and AND4 (N1895, N1885, N201, N1452, N1538);
nor NOR2 (N1896, N1890, N10);
xor XOR2 (N1897, N1896, N124);
and AND2 (N1898, N1875, N1155);
not NOT1 (N1899, N1897);
nor NOR3 (N1900, N1891, N774, N216);
nand NAND4 (N1901, N1889, N476, N526, N1797);
and AND3 (N1902, N1900, N937, N576);
nand NAND2 (N1903, N1901, N600);
not NOT1 (N1904, N1893);
not NOT1 (N1905, N1904);
buf BUF1 (N1906, N1887);
not NOT1 (N1907, N1899);
buf BUF1 (N1908, N1906);
or OR4 (N1909, N1888, N777, N1329, N216);
nor NOR2 (N1910, N1907, N801);
xor XOR2 (N1911, N1910, N972);
nand NAND3 (N1912, N1895, N285, N167);
xor XOR2 (N1913, N1898, N841);
nor NOR3 (N1914, N1911, N889, N1150);
and AND2 (N1915, N1909, N1555);
nor NOR4 (N1916, N1903, N1636, N1871, N528);
buf BUF1 (N1917, N1913);
not NOT1 (N1918, N1877);
nor NOR3 (N1919, N1908, N1645, N558);
not NOT1 (N1920, N1914);
and AND4 (N1921, N1894, N1859, N713, N20);
nand NAND3 (N1922, N1905, N947, N1047);
buf BUF1 (N1923, N1920);
nand NAND4 (N1924, N1916, N1749, N428, N1870);
xor XOR2 (N1925, N1921, N70);
or OR4 (N1926, N1924, N538, N542, N1175);
not NOT1 (N1927, N1902);
nor NOR3 (N1928, N1927, N1667, N1109);
or OR2 (N1929, N1919, N1426);
xor XOR2 (N1930, N1925, N486);
buf BUF1 (N1931, N1918);
not NOT1 (N1932, N1917);
nand NAND3 (N1933, N1915, N644, N795);
not NOT1 (N1934, N1923);
and AND3 (N1935, N1926, N563, N242);
nor NOR3 (N1936, N1935, N130, N1881);
buf BUF1 (N1937, N1931);
or OR2 (N1938, N1937, N1693);
nor NOR2 (N1939, N1912, N33);
or OR3 (N1940, N1934, N1682, N624);
or OR4 (N1941, N1940, N450, N299, N776);
nor NOR2 (N1942, N1933, N400);
not NOT1 (N1943, N1929);
not NOT1 (N1944, N1939);
nand NAND4 (N1945, N1922, N305, N1309, N1716);
buf BUF1 (N1946, N1944);
not NOT1 (N1947, N1943);
and AND2 (N1948, N1932, N1495);
or OR2 (N1949, N1936, N1309);
nor NOR4 (N1950, N1947, N1350, N1753, N757);
nand NAND2 (N1951, N1941, N1294);
or OR2 (N1952, N1948, N1121);
nand NAND2 (N1953, N1950, N705);
and AND4 (N1954, N1942, N841, N1657, N1532);
and AND2 (N1955, N1949, N423);
xor XOR2 (N1956, N1952, N90);
nand NAND2 (N1957, N1946, N230);
or OR2 (N1958, N1951, N1113);
and AND4 (N1959, N1957, N374, N1948, N1351);
nor NOR4 (N1960, N1954, N266, N871, N1589);
nor NOR4 (N1961, N1938, N1866, N1158, N1384);
or OR4 (N1962, N1960, N461, N1263, N880);
nand NAND4 (N1963, N1955, N1556, N1718, N1847);
not NOT1 (N1964, N1930);
nor NOR3 (N1965, N1945, N1387, N732);
xor XOR2 (N1966, N1956, N982);
or OR3 (N1967, N1958, N416, N1048);
not NOT1 (N1968, N1928);
or OR3 (N1969, N1959, N202, N294);
nor NOR4 (N1970, N1966, N1914, N1588, N914);
nor NOR2 (N1971, N1953, N1245);
buf BUF1 (N1972, N1970);
xor XOR2 (N1973, N1972, N1877);
nor NOR3 (N1974, N1962, N378, N820);
or OR2 (N1975, N1974, N533);
nor NOR2 (N1976, N1967, N1904);
or OR3 (N1977, N1976, N228, N394);
xor XOR2 (N1978, N1973, N1562);
or OR3 (N1979, N1971, N1057, N113);
nand NAND2 (N1980, N1978, N656);
buf BUF1 (N1981, N1965);
not NOT1 (N1982, N1963);
not NOT1 (N1983, N1982);
not NOT1 (N1984, N1979);
or OR4 (N1985, N1969, N1030, N186, N327);
nand NAND3 (N1986, N1984, N1546, N396);
nor NOR2 (N1987, N1975, N873);
nor NOR3 (N1988, N1986, N163, N1128);
xor XOR2 (N1989, N1980, N1046);
not NOT1 (N1990, N1977);
nand NAND2 (N1991, N1985, N217);
nor NOR2 (N1992, N1991, N1572);
buf BUF1 (N1993, N1981);
xor XOR2 (N1994, N1983, N140);
nand NAND4 (N1995, N1994, N1300, N1344, N950);
or OR2 (N1996, N1987, N1264);
or OR3 (N1997, N1968, N1375, N122);
xor XOR2 (N1998, N1996, N202);
nand NAND4 (N1999, N1989, N866, N100, N792);
and AND3 (N2000, N1993, N965, N56);
xor XOR2 (N2001, N1992, N1036);
not NOT1 (N2002, N1998);
nand NAND2 (N2003, N1997, N974);
not NOT1 (N2004, N2002);
nor NOR3 (N2005, N1990, N1901, N1030);
and AND3 (N2006, N2005, N1466, N1967);
xor XOR2 (N2007, N1988, N949);
xor XOR2 (N2008, N1964, N969);
and AND2 (N2009, N2006, N967);
nand NAND2 (N2010, N2000, N105);
or OR4 (N2011, N1961, N258, N1903, N955);
or OR4 (N2012, N2011, N633, N1648, N997);
nand NAND3 (N2013, N1999, N1019, N1679);
and AND3 (N2014, N2012, N474, N1319);
and AND2 (N2015, N2007, N413);
buf BUF1 (N2016, N2013);
buf BUF1 (N2017, N2003);
buf BUF1 (N2018, N2001);
nor NOR3 (N2019, N2016, N1276, N1438);
not NOT1 (N2020, N2019);
or OR2 (N2021, N2010, N835);
and AND2 (N2022, N2020, N146);
not NOT1 (N2023, N2014);
nor NOR2 (N2024, N2015, N567);
nor NOR4 (N2025, N2021, N729, N926, N942);
or OR2 (N2026, N2004, N492);
buf BUF1 (N2027, N2025);
nand NAND4 (N2028, N2018, N1497, N972, N1255);
not NOT1 (N2029, N2022);
or OR4 (N2030, N1995, N1539, N1631, N70);
nand NAND2 (N2031, N2027, N1018);
not NOT1 (N2032, N2024);
or OR4 (N2033, N2026, N794, N1551, N1492);
nor NOR2 (N2034, N2033, N775);
nand NAND3 (N2035, N2017, N456, N1103);
xor XOR2 (N2036, N2030, N1973);
nor NOR4 (N2037, N2035, N63, N368, N1013);
nand NAND4 (N2038, N2029, N584, N1807, N655);
or OR2 (N2039, N2037, N646);
or OR4 (N2040, N2036, N138, N509, N273);
nor NOR2 (N2041, N2023, N1876);
or OR3 (N2042, N2031, N1701, N1162);
xor XOR2 (N2043, N2039, N511);
or OR2 (N2044, N2042, N1286);
nor NOR2 (N2045, N2008, N656);
buf BUF1 (N2046, N2032);
and AND2 (N2047, N2044, N1951);
and AND3 (N2048, N2043, N450, N1202);
and AND4 (N2049, N2045, N1876, N894, N313);
not NOT1 (N2050, N2028);
not NOT1 (N2051, N2048);
xor XOR2 (N2052, N2050, N2045);
buf BUF1 (N2053, N2034);
buf BUF1 (N2054, N2051);
not NOT1 (N2055, N2049);
or OR4 (N2056, N2041, N1204, N1298, N393);
xor XOR2 (N2057, N2053, N1332);
buf BUF1 (N2058, N2047);
nor NOR3 (N2059, N2056, N1931, N1244);
xor XOR2 (N2060, N2054, N1547);
xor XOR2 (N2061, N2055, N1013);
or OR2 (N2062, N2061, N1602);
or OR2 (N2063, N2046, N824);
nand NAND3 (N2064, N2057, N1493, N1838);
xor XOR2 (N2065, N2063, N1410);
buf BUF1 (N2066, N2065);
nor NOR2 (N2067, N2060, N51);
buf BUF1 (N2068, N2067);
buf BUF1 (N2069, N2066);
not NOT1 (N2070, N2058);
or OR3 (N2071, N2064, N1132, N81);
not NOT1 (N2072, N2009);
not NOT1 (N2073, N2070);
and AND2 (N2074, N2062, N1135);
buf BUF1 (N2075, N2040);
not NOT1 (N2076, N2052);
nand NAND3 (N2077, N2071, N72, N1088);
xor XOR2 (N2078, N2077, N1558);
and AND4 (N2079, N2078, N1046, N444, N683);
nand NAND2 (N2080, N2074, N438);
nor NOR2 (N2081, N2075, N1283);
or OR4 (N2082, N2068, N318, N1309, N436);
not NOT1 (N2083, N2073);
or OR4 (N2084, N2069, N673, N439, N1680);
and AND4 (N2085, N2082, N389, N276, N234);
buf BUF1 (N2086, N2076);
or OR3 (N2087, N2085, N1780, N1844);
buf BUF1 (N2088, N2038);
nand NAND2 (N2089, N2080, N1709);
not NOT1 (N2090, N2086);
buf BUF1 (N2091, N2083);
or OR2 (N2092, N2087, N831);
nand NAND2 (N2093, N2081, N1124);
or OR3 (N2094, N2079, N1782, N367);
not NOT1 (N2095, N2084);
or OR2 (N2096, N2092, N1847);
and AND2 (N2097, N2090, N799);
not NOT1 (N2098, N2089);
nor NOR4 (N2099, N2072, N1076, N509, N1939);
xor XOR2 (N2100, N2094, N1070);
nor NOR2 (N2101, N2088, N1917);
buf BUF1 (N2102, N2096);
nand NAND3 (N2103, N2091, N2091, N1830);
not NOT1 (N2104, N2101);
not NOT1 (N2105, N2100);
buf BUF1 (N2106, N2098);
nor NOR4 (N2107, N2099, N1641, N883, N771);
not NOT1 (N2108, N2107);
buf BUF1 (N2109, N2106);
or OR4 (N2110, N2097, N75, N1094, N1588);
not NOT1 (N2111, N2109);
nor NOR2 (N2112, N2103, N860);
or OR3 (N2113, N2105, N159, N16);
nand NAND4 (N2114, N2108, N509, N1880, N1511);
nor NOR3 (N2115, N2114, N87, N1920);
not NOT1 (N2116, N2095);
and AND2 (N2117, N2111, N1996);
nand NAND3 (N2118, N2102, N1084, N1996);
not NOT1 (N2119, N2059);
and AND2 (N2120, N2116, N548);
or OR2 (N2121, N2093, N1517);
xor XOR2 (N2122, N2121, N1377);
xor XOR2 (N2123, N2113, N677);
and AND4 (N2124, N2122, N1396, N1681, N854);
nand NAND4 (N2125, N2119, N1790, N1775, N1295);
nand NAND3 (N2126, N2110, N1522, N2039);
buf BUF1 (N2127, N2124);
not NOT1 (N2128, N2104);
and AND4 (N2129, N2126, N1764, N2108, N554);
and AND2 (N2130, N2112, N1393);
xor XOR2 (N2131, N2120, N1023);
nor NOR4 (N2132, N2128, N2003, N446, N1052);
buf BUF1 (N2133, N2127);
not NOT1 (N2134, N2129);
buf BUF1 (N2135, N2131);
not NOT1 (N2136, N2132);
nor NOR4 (N2137, N2118, N1369, N245, N2131);
not NOT1 (N2138, N2123);
nand NAND4 (N2139, N2117, N1878, N1128, N1104);
nand NAND3 (N2140, N2115, N467, N1065);
nand NAND2 (N2141, N2137, N320);
not NOT1 (N2142, N2139);
xor XOR2 (N2143, N2136, N520);
nand NAND4 (N2144, N2142, N409, N1600, N1085);
not NOT1 (N2145, N2133);
and AND4 (N2146, N2135, N210, N1397, N1488);
or OR3 (N2147, N2141, N524, N470);
nand NAND4 (N2148, N2144, N59, N1206, N897);
or OR2 (N2149, N2140, N593);
buf BUF1 (N2150, N2148);
or OR3 (N2151, N2125, N520, N144);
not NOT1 (N2152, N2147);
nor NOR3 (N2153, N2145, N2064, N653);
and AND4 (N2154, N2151, N1505, N2013, N724);
xor XOR2 (N2155, N2150, N325);
buf BUF1 (N2156, N2149);
nor NOR4 (N2157, N2146, N911, N797, N1246);
not NOT1 (N2158, N2157);
nand NAND4 (N2159, N2156, N1378, N324, N945);
or OR2 (N2160, N2143, N1836);
xor XOR2 (N2161, N2154, N1217);
not NOT1 (N2162, N2153);
nand NAND2 (N2163, N2138, N962);
nor NOR3 (N2164, N2158, N1081, N82);
and AND3 (N2165, N2159, N2057, N1954);
nor NOR2 (N2166, N2164, N1829);
nand NAND3 (N2167, N2161, N746, N652);
nand NAND4 (N2168, N2167, N408, N1648, N1962);
nand NAND4 (N2169, N2162, N891, N818, N1346);
and AND3 (N2170, N2134, N1828, N1343);
not NOT1 (N2171, N2169);
nand NAND2 (N2172, N2165, N628);
or OR3 (N2173, N2168, N2134, N2105);
and AND2 (N2174, N2173, N1045);
or OR4 (N2175, N2170, N1198, N242, N394);
or OR4 (N2176, N2166, N714, N87, N180);
nor NOR2 (N2177, N2130, N1075);
nand NAND3 (N2178, N2176, N305, N1314);
and AND3 (N2179, N2152, N215, N314);
nor NOR2 (N2180, N2163, N607);
or OR4 (N2181, N2160, N2098, N87, N1472);
and AND4 (N2182, N2179, N186, N67, N1249);
nand NAND4 (N2183, N2177, N1557, N722, N1663);
xor XOR2 (N2184, N2180, N1227);
not NOT1 (N2185, N2178);
xor XOR2 (N2186, N2171, N758);
xor XOR2 (N2187, N2183, N972);
buf BUF1 (N2188, N2182);
and AND4 (N2189, N2175, N1005, N1474, N1138);
not NOT1 (N2190, N2174);
or OR2 (N2191, N2186, N1505);
or OR2 (N2192, N2188, N756);
and AND4 (N2193, N2189, N816, N201, N1680);
nor NOR3 (N2194, N2181, N1536, N737);
nand NAND2 (N2195, N2190, N1797);
nor NOR3 (N2196, N2172, N1752, N1075);
and AND2 (N2197, N2184, N57);
nor NOR2 (N2198, N2191, N177);
or OR4 (N2199, N2196, N1962, N1987, N1444);
xor XOR2 (N2200, N2192, N56);
nor NOR3 (N2201, N2194, N1047, N1428);
or OR4 (N2202, N2195, N1038, N458, N1374);
nand NAND4 (N2203, N2155, N1766, N1777, N1523);
and AND3 (N2204, N2187, N1191, N902);
nand NAND3 (N2205, N2201, N1346, N343);
xor XOR2 (N2206, N2185, N1560);
not NOT1 (N2207, N2193);
buf BUF1 (N2208, N2203);
or OR2 (N2209, N2200, N461);
or OR4 (N2210, N2208, N1662, N224, N482);
nor NOR3 (N2211, N2207, N1333, N149);
and AND3 (N2212, N2202, N17, N2163);
nand NAND4 (N2213, N2197, N1105, N1736, N1628);
or OR4 (N2214, N2204, N1764, N248, N1991);
nor NOR4 (N2215, N2198, N506, N718, N949);
buf BUF1 (N2216, N2212);
nand NAND4 (N2217, N2213, N245, N1674, N1863);
nor NOR2 (N2218, N2217, N1317);
or OR2 (N2219, N2214, N959);
buf BUF1 (N2220, N2215);
and AND2 (N2221, N2211, N1510);
buf BUF1 (N2222, N2221);
buf BUF1 (N2223, N2209);
buf BUF1 (N2224, N2223);
and AND3 (N2225, N2199, N2089, N689);
nand NAND4 (N2226, N2222, N1685, N1885, N818);
not NOT1 (N2227, N2218);
xor XOR2 (N2228, N2219, N414);
buf BUF1 (N2229, N2227);
xor XOR2 (N2230, N2224, N721);
buf BUF1 (N2231, N2206);
nor NOR4 (N2232, N2231, N1566, N1884, N435);
and AND4 (N2233, N2225, N2044, N421, N888);
and AND4 (N2234, N2230, N1657, N485, N1098);
or OR4 (N2235, N2228, N516, N437, N739);
buf BUF1 (N2236, N2229);
and AND3 (N2237, N2235, N1688, N1936);
and AND4 (N2238, N2233, N1378, N356, N995);
and AND4 (N2239, N2216, N1798, N901, N2196);
and AND4 (N2240, N2237, N1233, N2129, N1136);
not NOT1 (N2241, N2236);
and AND2 (N2242, N2239, N2154);
not NOT1 (N2243, N2210);
or OR3 (N2244, N2234, N1576, N414);
or OR4 (N2245, N2232, N271, N2096, N241);
nand NAND4 (N2246, N2205, N1088, N1655, N754);
nand NAND3 (N2247, N2242, N1116, N2233);
not NOT1 (N2248, N2220);
xor XOR2 (N2249, N2241, N672);
buf BUF1 (N2250, N2247);
or OR4 (N2251, N2245, N1965, N1233, N568);
and AND3 (N2252, N2244, N1993, N1507);
nand NAND3 (N2253, N2240, N290, N771);
or OR4 (N2254, N2250, N1442, N1086, N1560);
not NOT1 (N2255, N2254);
buf BUF1 (N2256, N2243);
not NOT1 (N2257, N2251);
and AND2 (N2258, N2249, N1054);
nand NAND4 (N2259, N2238, N2052, N987, N543);
and AND4 (N2260, N2252, N375, N303, N566);
xor XOR2 (N2261, N2248, N2102);
not NOT1 (N2262, N2246);
xor XOR2 (N2263, N2255, N814);
or OR3 (N2264, N2263, N1118, N2057);
nand NAND3 (N2265, N2256, N1012, N1042);
buf BUF1 (N2266, N2226);
not NOT1 (N2267, N2261);
or OR4 (N2268, N2257, N1000, N2230, N119);
nand NAND3 (N2269, N2259, N1757, N2085);
xor XOR2 (N2270, N2260, N2135);
and AND3 (N2271, N2258, N507, N2012);
not NOT1 (N2272, N2270);
buf BUF1 (N2273, N2269);
buf BUF1 (N2274, N2268);
or OR2 (N2275, N2271, N901);
or OR2 (N2276, N2273, N48);
nor NOR2 (N2277, N2267, N1749);
not NOT1 (N2278, N2276);
or OR3 (N2279, N2277, N1258, N406);
buf BUF1 (N2280, N2262);
xor XOR2 (N2281, N2265, N2097);
not NOT1 (N2282, N2280);
or OR3 (N2283, N2278, N1872, N1908);
or OR2 (N2284, N2279, N485);
nand NAND2 (N2285, N2281, N794);
xor XOR2 (N2286, N2264, N367);
xor XOR2 (N2287, N2283, N582);
nand NAND4 (N2288, N2275, N1188, N971, N968);
and AND3 (N2289, N2272, N173, N1138);
buf BUF1 (N2290, N2288);
nand NAND2 (N2291, N2266, N1253);
xor XOR2 (N2292, N2291, N2103);
buf BUF1 (N2293, N2286);
or OR4 (N2294, N2292, N1459, N642, N2170);
not NOT1 (N2295, N2253);
not NOT1 (N2296, N2295);
xor XOR2 (N2297, N2296, N1809);
xor XOR2 (N2298, N2297, N517);
xor XOR2 (N2299, N2287, N1485);
xor XOR2 (N2300, N2298, N1066);
xor XOR2 (N2301, N2290, N767);
and AND3 (N2302, N2293, N631, N1399);
buf BUF1 (N2303, N2285);
nor NOR3 (N2304, N2289, N1077, N783);
nor NOR3 (N2305, N2302, N1335, N2053);
and AND3 (N2306, N2305, N326, N422);
and AND3 (N2307, N2303, N1627, N193);
or OR3 (N2308, N2306, N100, N349);
nor NOR2 (N2309, N2301, N796);
nor NOR4 (N2310, N2308, N806, N954, N1830);
or OR4 (N2311, N2274, N678, N1947, N1479);
nor NOR4 (N2312, N2307, N1688, N2117, N2303);
or OR4 (N2313, N2299, N1847, N11, N2176);
and AND2 (N2314, N2310, N1661);
xor XOR2 (N2315, N2311, N1992);
and AND4 (N2316, N2309, N745, N1644, N237);
not NOT1 (N2317, N2312);
nand NAND3 (N2318, N2314, N2226, N67);
nor NOR4 (N2319, N2282, N917, N1039, N845);
and AND4 (N2320, N2315, N661, N899, N436);
or OR3 (N2321, N2304, N316, N1225);
buf BUF1 (N2322, N2300);
nand NAND2 (N2323, N2313, N1808);
and AND3 (N2324, N2316, N160, N2078);
nor NOR2 (N2325, N2317, N882);
and AND2 (N2326, N2321, N2308);
and AND2 (N2327, N2320, N1346);
and AND3 (N2328, N2323, N1731, N2112);
nand NAND3 (N2329, N2327, N2143, N878);
xor XOR2 (N2330, N2294, N231);
buf BUF1 (N2331, N2284);
xor XOR2 (N2332, N2329, N2193);
and AND3 (N2333, N2328, N1322, N684);
and AND2 (N2334, N2324, N2005);
nor NOR4 (N2335, N2332, N288, N631, N1799);
nand NAND3 (N2336, N2335, N919, N1512);
and AND4 (N2337, N2319, N603, N2167, N1152);
nor NOR4 (N2338, N2336, N1939, N1182, N919);
not NOT1 (N2339, N2330);
nor NOR2 (N2340, N2325, N1239);
nor NOR3 (N2341, N2322, N207, N1605);
and AND3 (N2342, N2333, N406, N1004);
not NOT1 (N2343, N2341);
not NOT1 (N2344, N2338);
nor NOR4 (N2345, N2343, N1565, N2250, N1655);
xor XOR2 (N2346, N2344, N643);
buf BUF1 (N2347, N2318);
buf BUF1 (N2348, N2326);
buf BUF1 (N2349, N2348);
nor NOR2 (N2350, N2340, N674);
not NOT1 (N2351, N2337);
xor XOR2 (N2352, N2331, N2287);
xor XOR2 (N2353, N2351, N2181);
buf BUF1 (N2354, N2352);
not NOT1 (N2355, N2347);
nor NOR2 (N2356, N2334, N543);
nand NAND2 (N2357, N2345, N1239);
or OR4 (N2358, N2357, N871, N1740, N201);
xor XOR2 (N2359, N2346, N2339);
nor NOR2 (N2360, N2224, N2289);
xor XOR2 (N2361, N2358, N2304);
or OR4 (N2362, N2349, N1365, N1231, N900);
nor NOR3 (N2363, N2342, N669, N1876);
xor XOR2 (N2364, N2350, N1623);
xor XOR2 (N2365, N2364, N323);
buf BUF1 (N2366, N2360);
buf BUF1 (N2367, N2365);
buf BUF1 (N2368, N2362);
nand NAND2 (N2369, N2366, N1250);
not NOT1 (N2370, N2363);
and AND4 (N2371, N2361, N199, N1655, N1927);
not NOT1 (N2372, N2367);
buf BUF1 (N2373, N2356);
or OR3 (N2374, N2371, N1708, N1291);
buf BUF1 (N2375, N2354);
not NOT1 (N2376, N2372);
not NOT1 (N2377, N2374);
nand NAND3 (N2378, N2377, N2370, N257);
buf BUF1 (N2379, N707);
buf BUF1 (N2380, N2369);
nand NAND2 (N2381, N2379, N369);
nor NOR2 (N2382, N2378, N1421);
nor NOR2 (N2383, N2355, N2041);
xor XOR2 (N2384, N2383, N2023);
buf BUF1 (N2385, N2375);
or OR3 (N2386, N2373, N377, N885);
or OR3 (N2387, N2359, N1501, N347);
or OR3 (N2388, N2386, N1395, N1839);
and AND2 (N2389, N2380, N2142);
buf BUF1 (N2390, N2387);
nor NOR4 (N2391, N2384, N1813, N1919, N1270);
and AND4 (N2392, N2382, N798, N2077, N952);
not NOT1 (N2393, N2389);
nand NAND2 (N2394, N2388, N821);
or OR3 (N2395, N2393, N509, N1015);
nand NAND2 (N2396, N2381, N48);
not NOT1 (N2397, N2390);
or OR3 (N2398, N2391, N536, N1725);
or OR3 (N2399, N2392, N330, N2046);
nand NAND2 (N2400, N2368, N2155);
buf BUF1 (N2401, N2400);
xor XOR2 (N2402, N2395, N1517);
or OR3 (N2403, N2376, N2014, N2059);
not NOT1 (N2404, N2402);
not NOT1 (N2405, N2396);
and AND4 (N2406, N2404, N799, N295, N1244);
and AND2 (N2407, N2353, N716);
buf BUF1 (N2408, N2403);
and AND2 (N2409, N2394, N49);
or OR4 (N2410, N2406, N4, N1606, N1034);
xor XOR2 (N2411, N2407, N7);
and AND3 (N2412, N2399, N1138, N2107);
nand NAND2 (N2413, N2408, N1964);
or OR3 (N2414, N2411, N2260, N1281);
not NOT1 (N2415, N2398);
and AND3 (N2416, N2401, N1960, N1148);
nand NAND3 (N2417, N2410, N1230, N2278);
nand NAND2 (N2418, N2405, N1459);
not NOT1 (N2419, N2417);
nand NAND4 (N2420, N2415, N85, N2331, N1812);
xor XOR2 (N2421, N2418, N920);
and AND3 (N2422, N2412, N1494, N594);
buf BUF1 (N2423, N2416);
not NOT1 (N2424, N2421);
and AND4 (N2425, N2413, N1521, N621, N420);
xor XOR2 (N2426, N2422, N1811);
nand NAND2 (N2427, N2424, N1544);
not NOT1 (N2428, N2409);
nor NOR2 (N2429, N2419, N199);
and AND3 (N2430, N2428, N140, N1196);
or OR2 (N2431, N2426, N2195);
not NOT1 (N2432, N2397);
nor NOR3 (N2433, N2423, N108, N529);
nor NOR2 (N2434, N2433, N2100);
xor XOR2 (N2435, N2425, N1376);
nor NOR3 (N2436, N2429, N1491, N1395);
nand NAND2 (N2437, N2436, N657);
or OR3 (N2438, N2430, N1845, N1374);
or OR4 (N2439, N2414, N1359, N1112, N913);
nor NOR4 (N2440, N2420, N998, N1531, N2267);
nor NOR2 (N2441, N2437, N393);
or OR4 (N2442, N2439, N2205, N1076, N1780);
buf BUF1 (N2443, N2434);
nand NAND4 (N2444, N2442, N2083, N1870, N764);
and AND3 (N2445, N2431, N74, N2386);
not NOT1 (N2446, N2432);
and AND2 (N2447, N2385, N343);
and AND2 (N2448, N2445, N630);
xor XOR2 (N2449, N2438, N325);
buf BUF1 (N2450, N2446);
not NOT1 (N2451, N2448);
nand NAND3 (N2452, N2449, N1191, N19);
not NOT1 (N2453, N2443);
not NOT1 (N2454, N2450);
buf BUF1 (N2455, N2454);
buf BUF1 (N2456, N2452);
buf BUF1 (N2457, N2451);
nand NAND3 (N2458, N2456, N698, N251);
nand NAND3 (N2459, N2453, N1885, N1466);
buf BUF1 (N2460, N2427);
nand NAND4 (N2461, N2459, N1814, N895, N589);
nand NAND2 (N2462, N2455, N1452);
and AND2 (N2463, N2461, N1575);
xor XOR2 (N2464, N2444, N1491);
or OR3 (N2465, N2447, N238, N1594);
or OR3 (N2466, N2460, N1975, N106);
or OR3 (N2467, N2440, N2204, N2120);
nor NOR4 (N2468, N2457, N222, N1667, N977);
xor XOR2 (N2469, N2458, N2338);
nor NOR2 (N2470, N2464, N112);
xor XOR2 (N2471, N2468, N1816);
xor XOR2 (N2472, N2465, N1847);
and AND3 (N2473, N2470, N929, N2362);
buf BUF1 (N2474, N2472);
or OR4 (N2475, N2471, N1047, N2156, N192);
buf BUF1 (N2476, N2469);
buf BUF1 (N2477, N2466);
xor XOR2 (N2478, N2441, N1794);
or OR2 (N2479, N2473, N2073);
not NOT1 (N2480, N2478);
or OR4 (N2481, N2462, N2077, N1158, N1345);
not NOT1 (N2482, N2480);
and AND3 (N2483, N2435, N1466, N448);
xor XOR2 (N2484, N2477, N166);
nor NOR3 (N2485, N2476, N908, N2443);
not NOT1 (N2486, N2485);
not NOT1 (N2487, N2475);
not NOT1 (N2488, N2482);
nor NOR2 (N2489, N2463, N1006);
or OR3 (N2490, N2483, N1936, N2477);
and AND3 (N2491, N2467, N1249, N598);
nand NAND2 (N2492, N2481, N645);
and AND4 (N2493, N2474, N876, N2114, N378);
nand NAND2 (N2494, N2487, N1289);
nor NOR4 (N2495, N2490, N1090, N1910, N2165);
and AND2 (N2496, N2491, N1977);
and AND3 (N2497, N2479, N2336, N2141);
or OR4 (N2498, N2494, N1165, N480, N2242);
xor XOR2 (N2499, N2486, N1746);
and AND3 (N2500, N2492, N254, N1480);
and AND3 (N2501, N2500, N1714, N984);
xor XOR2 (N2502, N2498, N824);
nand NAND4 (N2503, N2489, N200, N2343, N407);
buf BUF1 (N2504, N2502);
and AND4 (N2505, N2484, N1264, N1685, N1379);
not NOT1 (N2506, N2496);
buf BUF1 (N2507, N2493);
nor NOR2 (N2508, N2488, N1755);
and AND4 (N2509, N2507, N1925, N1842, N1508);
xor XOR2 (N2510, N2503, N1821);
buf BUF1 (N2511, N2510);
or OR4 (N2512, N2499, N2059, N1207, N2430);
not NOT1 (N2513, N2501);
nor NOR3 (N2514, N2495, N2333, N2512);
xor XOR2 (N2515, N1473, N2096);
xor XOR2 (N2516, N2513, N6);
xor XOR2 (N2517, N2514, N2163);
buf BUF1 (N2518, N2511);
not NOT1 (N2519, N2518);
buf BUF1 (N2520, N2515);
nor NOR3 (N2521, N2519, N1581, N1417);
nor NOR3 (N2522, N2497, N1430, N1916);
nor NOR3 (N2523, N2506, N159, N14);
or OR4 (N2524, N2520, N64, N435, N976);
not NOT1 (N2525, N2505);
nand NAND4 (N2526, N2523, N1379, N283, N1559);
nor NOR3 (N2527, N2516, N558, N1426);
not NOT1 (N2528, N2508);
nor NOR3 (N2529, N2525, N2192, N2086);
or OR2 (N2530, N2509, N1229);
nand NAND2 (N2531, N2530, N1041);
or OR4 (N2532, N2524, N1447, N382, N1345);
buf BUF1 (N2533, N2522);
nor NOR4 (N2534, N2521, N1608, N1817, N992);
nor NOR3 (N2535, N2517, N1532, N2219);
nor NOR2 (N2536, N2531, N873);
or OR2 (N2537, N2504, N1227);
nor NOR2 (N2538, N2536, N1504);
buf BUF1 (N2539, N2526);
or OR2 (N2540, N2538, N1041);
or OR3 (N2541, N2527, N1780, N2424);
xor XOR2 (N2542, N2532, N1567);
and AND3 (N2543, N2537, N1545, N636);
and AND2 (N2544, N2535, N1877);
xor XOR2 (N2545, N2528, N384);
or OR3 (N2546, N2529, N1726, N1201);
not NOT1 (N2547, N2546);
buf BUF1 (N2548, N2533);
buf BUF1 (N2549, N2548);
or OR3 (N2550, N2543, N1701, N764);
buf BUF1 (N2551, N2539);
nand NAND2 (N2552, N2534, N1001);
nand NAND4 (N2553, N2547, N1952, N92, N1725);
nand NAND4 (N2554, N2551, N2135, N1824, N933);
or OR2 (N2555, N2554, N2138);
nand NAND3 (N2556, N2541, N2320, N1734);
nand NAND3 (N2557, N2544, N597, N1385);
xor XOR2 (N2558, N2550, N2323);
nand NAND3 (N2559, N2540, N1547, N1862);
not NOT1 (N2560, N2552);
not NOT1 (N2561, N2545);
buf BUF1 (N2562, N2560);
not NOT1 (N2563, N2553);
buf BUF1 (N2564, N2562);
or OR3 (N2565, N2563, N911, N2481);
xor XOR2 (N2566, N2561, N895);
not NOT1 (N2567, N2549);
xor XOR2 (N2568, N2566, N2514);
nor NOR2 (N2569, N2556, N1797);
not NOT1 (N2570, N2568);
buf BUF1 (N2571, N2555);
not NOT1 (N2572, N2558);
not NOT1 (N2573, N2565);
and AND2 (N2574, N2571, N10);
nor NOR4 (N2575, N2557, N2455, N1353, N859);
xor XOR2 (N2576, N2567, N1560);
buf BUF1 (N2577, N2572);
not NOT1 (N2578, N2559);
xor XOR2 (N2579, N2577, N811);
buf BUF1 (N2580, N2578);
or OR2 (N2581, N2570, N1211);
and AND2 (N2582, N2581, N1272);
nand NAND3 (N2583, N2575, N1682, N384);
and AND4 (N2584, N2573, N876, N1862, N1631);
xor XOR2 (N2585, N2579, N1977);
nor NOR4 (N2586, N2584, N243, N1225, N164);
xor XOR2 (N2587, N2586, N213);
nand NAND4 (N2588, N2569, N1518, N1005, N657);
xor XOR2 (N2589, N2542, N2554);
and AND3 (N2590, N2580, N1908, N62);
or OR3 (N2591, N2574, N277, N32);
nor NOR3 (N2592, N2564, N915, N110);
not NOT1 (N2593, N2583);
not NOT1 (N2594, N2589);
buf BUF1 (N2595, N2594);
nand NAND3 (N2596, N2585, N140, N2519);
nor NOR4 (N2597, N2587, N2536, N2475, N1909);
nor NOR4 (N2598, N2591, N1281, N1570, N2522);
not NOT1 (N2599, N2576);
buf BUF1 (N2600, N2597);
xor XOR2 (N2601, N2595, N2469);
nand NAND2 (N2602, N2598, N1585);
xor XOR2 (N2603, N2596, N2114);
nor NOR2 (N2604, N2592, N1918);
not NOT1 (N2605, N2600);
and AND3 (N2606, N2590, N81, N1335);
nor NOR2 (N2607, N2599, N2210);
and AND4 (N2608, N2593, N31, N1954, N1959);
nand NAND3 (N2609, N2605, N1259, N663);
buf BUF1 (N2610, N2603);
nor NOR2 (N2611, N2606, N1783);
not NOT1 (N2612, N2611);
buf BUF1 (N2613, N2608);
nand NAND3 (N2614, N2604, N1027, N2164);
nand NAND2 (N2615, N2609, N2540);
nand NAND3 (N2616, N2588, N1253, N2590);
or OR4 (N2617, N2601, N1754, N1684, N1584);
or OR2 (N2618, N2615, N2145);
xor XOR2 (N2619, N2612, N1353);
and AND2 (N2620, N2619, N2562);
nor NOR2 (N2621, N2582, N384);
or OR2 (N2622, N2614, N1079);
not NOT1 (N2623, N2616);
nand NAND2 (N2624, N2602, N171);
not NOT1 (N2625, N2618);
xor XOR2 (N2626, N2622, N2024);
buf BUF1 (N2627, N2617);
not NOT1 (N2628, N2613);
or OR4 (N2629, N2628, N864, N39, N1703);
and AND2 (N2630, N2627, N115);
buf BUF1 (N2631, N2623);
and AND4 (N2632, N2630, N1603, N2043, N1140);
or OR2 (N2633, N2631, N340);
not NOT1 (N2634, N2610);
not NOT1 (N2635, N2620);
nor NOR4 (N2636, N2635, N2061, N423, N844);
xor XOR2 (N2637, N2632, N2345);
nor NOR3 (N2638, N2607, N310, N156);
xor XOR2 (N2639, N2625, N2339);
nand NAND3 (N2640, N2639, N1517, N1992);
or OR2 (N2641, N2638, N341);
or OR4 (N2642, N2621, N2304, N303, N2028);
xor XOR2 (N2643, N2637, N2127);
or OR4 (N2644, N2643, N447, N565, N1776);
buf BUF1 (N2645, N2634);
buf BUF1 (N2646, N2636);
nor NOR2 (N2647, N2642, N949);
xor XOR2 (N2648, N2640, N391);
and AND3 (N2649, N2633, N117, N1625);
and AND4 (N2650, N2629, N1602, N2397, N1445);
and AND4 (N2651, N2649, N375, N1575, N770);
not NOT1 (N2652, N2650);
not NOT1 (N2653, N2624);
nand NAND4 (N2654, N2648, N1721, N632, N1455);
buf BUF1 (N2655, N2641);
or OR3 (N2656, N2655, N1744, N1418);
and AND4 (N2657, N2646, N2375, N101, N2239);
not NOT1 (N2658, N2647);
xor XOR2 (N2659, N2658, N1861);
or OR2 (N2660, N2626, N1361);
not NOT1 (N2661, N2656);
and AND3 (N2662, N2644, N1133, N2370);
and AND3 (N2663, N2645, N701, N313);
nand NAND4 (N2664, N2657, N957, N1666, N2536);
and AND2 (N2665, N2661, N93);
buf BUF1 (N2666, N2662);
buf BUF1 (N2667, N2654);
and AND4 (N2668, N2651, N2303, N1847, N1240);
or OR2 (N2669, N2664, N2144);
nor NOR4 (N2670, N2669, N903, N1958, N98);
xor XOR2 (N2671, N2665, N2185);
buf BUF1 (N2672, N2668);
not NOT1 (N2673, N2660);
or OR4 (N2674, N2663, N1641, N540, N1675);
xor XOR2 (N2675, N2666, N2328);
or OR4 (N2676, N2673, N606, N2388, N2504);
buf BUF1 (N2677, N2653);
not NOT1 (N2678, N2670);
or OR2 (N2679, N2659, N1327);
not NOT1 (N2680, N2678);
nand NAND2 (N2681, N2676, N1670);
nor NOR2 (N2682, N2680, N1941);
or OR4 (N2683, N2674, N1417, N1606, N1853);
and AND3 (N2684, N2682, N163, N1524);
buf BUF1 (N2685, N2667);
nand NAND2 (N2686, N2685, N84);
nand NAND3 (N2687, N2652, N1099, N1018);
and AND3 (N2688, N2684, N974, N1647);
xor XOR2 (N2689, N2683, N330);
and AND4 (N2690, N2688, N769, N36, N208);
xor XOR2 (N2691, N2687, N2630);
nor NOR3 (N2692, N2686, N846, N2683);
nor NOR3 (N2693, N2690, N1238, N906);
or OR3 (N2694, N2679, N2474, N651);
and AND2 (N2695, N2694, N435);
xor XOR2 (N2696, N2675, N877);
or OR2 (N2697, N2692, N1157);
or OR3 (N2698, N2671, N718, N1774);
buf BUF1 (N2699, N2696);
buf BUF1 (N2700, N2677);
not NOT1 (N2701, N2697);
buf BUF1 (N2702, N2689);
and AND4 (N2703, N2672, N738, N995, N208);
and AND4 (N2704, N2701, N1877, N828, N1168);
and AND4 (N2705, N2700, N602, N2397, N1475);
nor NOR4 (N2706, N2704, N2163, N185, N2340);
nand NAND2 (N2707, N2699, N418);
or OR4 (N2708, N2695, N1420, N2371, N990);
not NOT1 (N2709, N2708);
and AND4 (N2710, N2703, N1810, N908, N2598);
or OR4 (N2711, N2698, N2588, N1196, N496);
buf BUF1 (N2712, N2705);
buf BUF1 (N2713, N2710);
and AND3 (N2714, N2709, N297, N2559);
xor XOR2 (N2715, N2706, N2251);
not NOT1 (N2716, N2712);
nand NAND4 (N2717, N2716, N2057, N1667, N2705);
nand NAND4 (N2718, N2714, N2067, N2601, N313);
not NOT1 (N2719, N2718);
nand NAND3 (N2720, N2713, N1872, N413);
nor NOR4 (N2721, N2720, N2630, N2006, N251);
not NOT1 (N2722, N2715);
or OR4 (N2723, N2702, N1196, N436, N1577);
nand NAND4 (N2724, N2707, N916, N340, N1058);
and AND3 (N2725, N2721, N1930, N2132);
nand NAND4 (N2726, N2691, N364, N1449, N636);
and AND4 (N2727, N2717, N1532, N453, N1949);
xor XOR2 (N2728, N2693, N1597);
nor NOR3 (N2729, N2726, N533, N1700);
and AND2 (N2730, N2724, N1025);
and AND4 (N2731, N2681, N1920, N748, N1675);
or OR4 (N2732, N2725, N2375, N1195, N1797);
not NOT1 (N2733, N2711);
and AND4 (N2734, N2729, N817, N2215, N2731);
or OR3 (N2735, N237, N1340, N1894);
xor XOR2 (N2736, N2719, N1578);
and AND3 (N2737, N2736, N2712, N2710);
nand NAND3 (N2738, N2730, N119, N272);
nand NAND3 (N2739, N2733, N1798, N1391);
and AND2 (N2740, N2732, N742);
xor XOR2 (N2741, N2722, N1729);
nor NOR4 (N2742, N2734, N2725, N396, N117);
and AND3 (N2743, N2742, N2497, N2282);
and AND3 (N2744, N2740, N2100, N1315);
nor NOR3 (N2745, N2744, N1944, N1663);
xor XOR2 (N2746, N2739, N1611);
nand NAND2 (N2747, N2737, N2339);
or OR3 (N2748, N2741, N81, N2363);
nor NOR3 (N2749, N2735, N2249, N1234);
nor NOR4 (N2750, N2738, N662, N1579, N501);
buf BUF1 (N2751, N2727);
and AND4 (N2752, N2728, N1519, N542, N1383);
xor XOR2 (N2753, N2746, N2053);
xor XOR2 (N2754, N2753, N1693);
not NOT1 (N2755, N2747);
and AND4 (N2756, N2745, N110, N130, N1928);
and AND2 (N2757, N2750, N1992);
not NOT1 (N2758, N2756);
and AND4 (N2759, N2751, N375, N2024, N329);
not NOT1 (N2760, N2754);
or OR3 (N2761, N2759, N2634, N265);
xor XOR2 (N2762, N2743, N805);
not NOT1 (N2763, N2761);
buf BUF1 (N2764, N2723);
not NOT1 (N2765, N2752);
xor XOR2 (N2766, N2764, N605);
and AND3 (N2767, N2763, N673, N49);
or OR4 (N2768, N2767, N2037, N197, N2190);
and AND3 (N2769, N2758, N1762, N962);
not NOT1 (N2770, N2748);
buf BUF1 (N2771, N2766);
xor XOR2 (N2772, N2762, N423);
xor XOR2 (N2773, N2771, N1097);
buf BUF1 (N2774, N2765);
or OR3 (N2775, N2770, N1120, N1444);
nand NAND3 (N2776, N2749, N9, N284);
not NOT1 (N2777, N2772);
buf BUF1 (N2778, N2768);
xor XOR2 (N2779, N2760, N1529);
or OR3 (N2780, N2777, N962, N1633);
and AND2 (N2781, N2778, N1903);
nor NOR2 (N2782, N2779, N582);
xor XOR2 (N2783, N2781, N1749);
and AND3 (N2784, N2757, N2700, N1646);
and AND2 (N2785, N2769, N1179);
xor XOR2 (N2786, N2783, N1480);
or OR3 (N2787, N2773, N2558, N2757);
nand NAND3 (N2788, N2784, N1659, N146);
not NOT1 (N2789, N2776);
not NOT1 (N2790, N2780);
buf BUF1 (N2791, N2782);
not NOT1 (N2792, N2789);
xor XOR2 (N2793, N2792, N286);
not NOT1 (N2794, N2790);
buf BUF1 (N2795, N2793);
not NOT1 (N2796, N2787);
nor NOR2 (N2797, N2795, N2533);
nor NOR3 (N2798, N2785, N2594, N784);
not NOT1 (N2799, N2755);
xor XOR2 (N2800, N2774, N2644);
nor NOR2 (N2801, N2786, N1003);
not NOT1 (N2802, N2799);
or OR4 (N2803, N2800, N704, N2356, N2752);
xor XOR2 (N2804, N2803, N2232);
or OR3 (N2805, N2791, N2716, N1315);
nand NAND4 (N2806, N2797, N881, N2455, N420);
nor NOR3 (N2807, N2806, N1461, N1684);
not NOT1 (N2808, N2794);
and AND2 (N2809, N2775, N103);
xor XOR2 (N2810, N2801, N1721);
or OR2 (N2811, N2796, N1247);
nand NAND4 (N2812, N2807, N177, N2673, N737);
nor NOR2 (N2813, N2812, N1502);
not NOT1 (N2814, N2808);
buf BUF1 (N2815, N2802);
buf BUF1 (N2816, N2809);
nor NOR2 (N2817, N2816, N63);
not NOT1 (N2818, N2788);
nand NAND2 (N2819, N2810, N570);
nor NOR2 (N2820, N2817, N1763);
nand NAND2 (N2821, N2814, N1720);
and AND4 (N2822, N2819, N2430, N2016, N2221);
and AND3 (N2823, N2813, N1225, N2102);
xor XOR2 (N2824, N2805, N2751);
xor XOR2 (N2825, N2804, N433);
buf BUF1 (N2826, N2822);
xor XOR2 (N2827, N2826, N2500);
nand NAND4 (N2828, N2827, N1778, N305, N2646);
not NOT1 (N2829, N2823);
not NOT1 (N2830, N2825);
not NOT1 (N2831, N2818);
nor NOR4 (N2832, N2821, N2276, N425, N1242);
nand NAND4 (N2833, N2811, N1031, N603, N374);
and AND3 (N2834, N2815, N647, N1884);
or OR2 (N2835, N2832, N2823);
xor XOR2 (N2836, N2820, N1695);
nor NOR4 (N2837, N2824, N2540, N2052, N1099);
not NOT1 (N2838, N2837);
nor NOR2 (N2839, N2831, N928);
buf BUF1 (N2840, N2828);
xor XOR2 (N2841, N2830, N1041);
or OR2 (N2842, N2798, N2570);
or OR3 (N2843, N2835, N242, N1679);
or OR3 (N2844, N2839, N1211, N317);
nand NAND3 (N2845, N2843, N2503, N1681);
nor NOR4 (N2846, N2836, N2075, N1643, N2699);
nand NAND2 (N2847, N2841, N2322);
not NOT1 (N2848, N2833);
buf BUF1 (N2849, N2838);
not NOT1 (N2850, N2829);
buf BUF1 (N2851, N2844);
nand NAND2 (N2852, N2834, N135);
and AND3 (N2853, N2849, N1518, N2530);
xor XOR2 (N2854, N2842, N1784);
not NOT1 (N2855, N2851);
and AND2 (N2856, N2840, N178);
nand NAND3 (N2857, N2847, N1842, N974);
nand NAND2 (N2858, N2845, N654);
or OR3 (N2859, N2846, N1957, N1705);
nand NAND4 (N2860, N2857, N2022, N138, N878);
and AND4 (N2861, N2855, N1189, N1399, N2417);
nor NOR3 (N2862, N2854, N388, N1434);
or OR3 (N2863, N2861, N1799, N795);
nor NOR3 (N2864, N2858, N1673, N2258);
and AND3 (N2865, N2864, N439, N1141);
buf BUF1 (N2866, N2860);
nor NOR2 (N2867, N2862, N2339);
or OR4 (N2868, N2866, N928, N1695, N1775);
xor XOR2 (N2869, N2859, N2593);
buf BUF1 (N2870, N2852);
nand NAND4 (N2871, N2869, N1555, N2752, N1605);
nor NOR4 (N2872, N2863, N362, N1665, N2140);
or OR2 (N2873, N2848, N297);
nand NAND3 (N2874, N2867, N2338, N375);
xor XOR2 (N2875, N2874, N1154);
nand NAND4 (N2876, N2870, N1777, N46, N1217);
xor XOR2 (N2877, N2868, N2652);
xor XOR2 (N2878, N2873, N1547);
nor NOR3 (N2879, N2875, N2473, N613);
buf BUF1 (N2880, N2872);
and AND4 (N2881, N2853, N2728, N198, N286);
nor NOR2 (N2882, N2871, N2404);
xor XOR2 (N2883, N2856, N1412);
buf BUF1 (N2884, N2878);
nor NOR4 (N2885, N2880, N1526, N302, N391);
and AND4 (N2886, N2884, N2767, N2828, N462);
not NOT1 (N2887, N2850);
nor NOR2 (N2888, N2885, N1239);
and AND2 (N2889, N2888, N527);
and AND4 (N2890, N2887, N878, N2076, N1683);
not NOT1 (N2891, N2865);
buf BUF1 (N2892, N2886);
not NOT1 (N2893, N2877);
or OR2 (N2894, N2889, N1466);
or OR4 (N2895, N2879, N163, N2859, N1524);
not NOT1 (N2896, N2876);
nand NAND3 (N2897, N2894, N2040, N898);
xor XOR2 (N2898, N2893, N1543);
nand NAND2 (N2899, N2890, N2648);
and AND3 (N2900, N2899, N2522, N1010);
nand NAND3 (N2901, N2897, N2087, N2275);
buf BUF1 (N2902, N2881);
xor XOR2 (N2903, N2891, N662);
or OR4 (N2904, N2902, N170, N1244, N2039);
or OR4 (N2905, N2904, N143, N2611, N2247);
nand NAND2 (N2906, N2882, N2670);
or OR2 (N2907, N2892, N1171);
nand NAND3 (N2908, N2906, N864, N582);
and AND4 (N2909, N2903, N1240, N1556, N2711);
or OR4 (N2910, N2901, N2496, N1431, N819);
not NOT1 (N2911, N2907);
not NOT1 (N2912, N2909);
nand NAND3 (N2913, N2908, N375, N1791);
nor NOR4 (N2914, N2883, N271, N2048, N201);
not NOT1 (N2915, N2910);
xor XOR2 (N2916, N2914, N2449);
and AND3 (N2917, N2898, N1385, N1907);
nand NAND2 (N2918, N2905, N783);
nor NOR4 (N2919, N2895, N2418, N2076, N1707);
or OR4 (N2920, N2915, N2313, N2893, N1452);
not NOT1 (N2921, N2920);
nand NAND4 (N2922, N2912, N1954, N316, N2278);
nor NOR4 (N2923, N2896, N763, N2662, N2841);
not NOT1 (N2924, N2916);
xor XOR2 (N2925, N2923, N50);
buf BUF1 (N2926, N2925);
and AND4 (N2927, N2924, N400, N2562, N423);
not NOT1 (N2928, N2922);
xor XOR2 (N2929, N2911, N2527);
nor NOR4 (N2930, N2919, N2359, N2087, N971);
buf BUF1 (N2931, N2930);
or OR4 (N2932, N2931, N1455, N1443, N1218);
nor NOR4 (N2933, N2928, N1247, N1297, N1197);
nand NAND4 (N2934, N2900, N222, N1225, N591);
xor XOR2 (N2935, N2934, N2859);
nor NOR3 (N2936, N2929, N1235, N194);
or OR3 (N2937, N2926, N2161, N1525);
nand NAND3 (N2938, N2913, N555, N84);
nand NAND3 (N2939, N2932, N924, N360);
and AND2 (N2940, N2939, N2700);
not NOT1 (N2941, N2918);
nor NOR2 (N2942, N2917, N1474);
not NOT1 (N2943, N2942);
or OR2 (N2944, N2921, N1584);
or OR2 (N2945, N2933, N1412);
not NOT1 (N2946, N2936);
or OR3 (N2947, N2927, N1159, N1488);
xor XOR2 (N2948, N2943, N1295);
nand NAND4 (N2949, N2944, N523, N2376, N377);
buf BUF1 (N2950, N2935);
nand NAND2 (N2951, N2947, N83);
and AND3 (N2952, N2948, N2779, N35);
not NOT1 (N2953, N2940);
and AND4 (N2954, N2951, N948, N1813, N606);
or OR4 (N2955, N2946, N2009, N1539, N734);
nand NAND2 (N2956, N2954, N735);
xor XOR2 (N2957, N2937, N2296);
nand NAND3 (N2958, N2938, N197, N597);
buf BUF1 (N2959, N2952);
buf BUF1 (N2960, N2949);
or OR2 (N2961, N2960, N1568);
nand NAND4 (N2962, N2945, N1973, N949, N151);
and AND2 (N2963, N2958, N681);
nand NAND4 (N2964, N2950, N613, N1268, N783);
not NOT1 (N2965, N2956);
and AND2 (N2966, N2957, N2476);
nor NOR4 (N2967, N2959, N476, N354, N320);
nor NOR4 (N2968, N2953, N2700, N1907, N14);
nor NOR4 (N2969, N2964, N2702, N753, N16);
or OR3 (N2970, N2968, N1264, N890);
nand NAND4 (N2971, N2963, N1893, N1515, N1768);
xor XOR2 (N2972, N2955, N2889);
or OR3 (N2973, N2969, N316, N1877);
nor NOR2 (N2974, N2966, N1838);
nor NOR4 (N2975, N2967, N1924, N1046, N2025);
and AND4 (N2976, N2972, N2686, N132, N1405);
not NOT1 (N2977, N2975);
xor XOR2 (N2978, N2961, N245);
nand NAND3 (N2979, N2976, N2084, N251);
or OR4 (N2980, N2974, N562, N1430, N1405);
nor NOR3 (N2981, N2971, N2870, N2226);
xor XOR2 (N2982, N2981, N2212);
not NOT1 (N2983, N2982);
xor XOR2 (N2984, N2978, N668);
buf BUF1 (N2985, N2941);
and AND2 (N2986, N2985, N515);
and AND3 (N2987, N2970, N398, N2534);
nand NAND4 (N2988, N2980, N884, N528, N2310);
or OR4 (N2989, N2988, N2250, N2603, N1043);
nand NAND2 (N2990, N2986, N805);
buf BUF1 (N2991, N2989);
not NOT1 (N2992, N2987);
buf BUF1 (N2993, N2983);
xor XOR2 (N2994, N2973, N1177);
or OR3 (N2995, N2993, N553, N2772);
not NOT1 (N2996, N2962);
nand NAND3 (N2997, N2965, N2346, N852);
or OR4 (N2998, N2991, N722, N91, N794);
or OR4 (N2999, N2984, N147, N299, N861);
xor XOR2 (N3000, N2997, N1173);
not NOT1 (N3001, N2994);
buf BUF1 (N3002, N2998);
or OR2 (N3003, N2990, N1739);
nor NOR2 (N3004, N2992, N165);
not NOT1 (N3005, N2977);
nand NAND4 (N3006, N3000, N183, N983, N409);
not NOT1 (N3007, N3001);
buf BUF1 (N3008, N3004);
or OR2 (N3009, N3006, N2411);
not NOT1 (N3010, N3002);
not NOT1 (N3011, N2999);
or OR2 (N3012, N3009, N1890);
not NOT1 (N3013, N3010);
and AND3 (N3014, N3003, N1622, N561);
and AND4 (N3015, N2979, N340, N867, N854);
xor XOR2 (N3016, N3008, N1387);
or OR4 (N3017, N3012, N76, N586, N2316);
buf BUF1 (N3018, N3013);
nor NOR4 (N3019, N3011, N2492, N2420, N1279);
nor NOR4 (N3020, N3016, N2078, N45, N2236);
xor XOR2 (N3021, N3018, N1374);
endmodule